// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N15963,N16012,N16004,N16009,N16007,N16013,N16011,N16003,N16014,N16015;

buf BUF1 (N16, N12);
and AND2 (N17, N5, N2);
nor NOR2 (N18, N2, N11);
buf BUF1 (N19, N4);
and AND4 (N20, N11, N16, N11, N7);
buf BUF1 (N21, N15);
nand NAND3 (N22, N16, N2, N7);
and AND3 (N23, N20, N1, N20);
nor NOR2 (N24, N20, N13);
nand NAND4 (N25, N11, N16, N24, N12);
buf BUF1 (N26, N8);
or OR4 (N27, N19, N14, N8, N8);
or OR3 (N28, N5, N7, N16);
buf BUF1 (N29, N2);
or OR2 (N30, N29, N4);
nand NAND3 (N31, N25, N6, N29);
buf BUF1 (N32, N26);
nor NOR4 (N33, N28, N18, N6, N28);
not NOT1 (N34, N19);
nand NAND4 (N35, N17, N30, N26, N11);
buf BUF1 (N36, N31);
nor NOR4 (N37, N36, N14, N35, N35);
xor XOR2 (N38, N11, N10);
buf BUF1 (N39, N16);
nor NOR2 (N40, N39, N19);
nor NOR4 (N41, N23, N34, N29, N8);
nand NAND4 (N42, N19, N15, N33, N18);
or OR2 (N43, N1, N15);
buf BUF1 (N44, N37);
nor NOR3 (N45, N32, N33, N15);
nor NOR4 (N46, N43, N14, N33, N3);
nand NAND2 (N47, N40, N33);
or OR3 (N48, N27, N37, N47);
xor XOR2 (N49, N35, N3);
nor NOR2 (N50, N49, N14);
not NOT1 (N51, N41);
xor XOR2 (N52, N46, N5);
xor XOR2 (N53, N52, N12);
nor NOR2 (N54, N21, N29);
buf BUF1 (N55, N38);
not NOT1 (N56, N53);
xor XOR2 (N57, N51, N19);
nor NOR2 (N58, N56, N54);
xor XOR2 (N59, N19, N38);
nand NAND2 (N60, N50, N24);
and AND3 (N61, N48, N47, N46);
nor NOR3 (N62, N61, N18, N44);
or OR2 (N63, N7, N55);
xor XOR2 (N64, N46, N14);
buf BUF1 (N65, N42);
not NOT1 (N66, N64);
xor XOR2 (N67, N59, N13);
xor XOR2 (N68, N58, N6);
not NOT1 (N69, N66);
and AND2 (N70, N63, N16);
nor NOR2 (N71, N22, N24);
not NOT1 (N72, N65);
or OR4 (N73, N71, N13, N70, N27);
nand NAND4 (N74, N46, N46, N40, N45);
nor NOR4 (N75, N43, N38, N44, N34);
nor NOR3 (N76, N68, N8, N58);
nand NAND2 (N77, N62, N34);
and AND4 (N78, N74, N74, N20, N49);
nand NAND2 (N79, N67, N63);
nand NAND2 (N80, N79, N13);
buf BUF1 (N81, N78);
xor XOR2 (N82, N76, N20);
not NOT1 (N83, N69);
or OR2 (N84, N72, N69);
nor NOR4 (N85, N83, N62, N18, N25);
buf BUF1 (N86, N60);
xor XOR2 (N87, N81, N22);
xor XOR2 (N88, N84, N9);
nor NOR4 (N89, N82, N45, N12, N58);
xor XOR2 (N90, N75, N3);
buf BUF1 (N91, N77);
and AND4 (N92, N88, N9, N43, N85);
buf BUF1 (N93, N22);
nand NAND4 (N94, N86, N44, N76, N35);
or OR3 (N95, N80, N75, N8);
nor NOR4 (N96, N90, N47, N26, N83);
xor XOR2 (N97, N73, N70);
nand NAND2 (N98, N96, N26);
xor XOR2 (N99, N89, N79);
and AND4 (N100, N87, N7, N91, N84);
or OR3 (N101, N73, N68, N94);
nor NOR3 (N102, N88, N17, N20);
xor XOR2 (N103, N98, N73);
nor NOR2 (N104, N102, N82);
and AND4 (N105, N103, N34, N76, N74);
buf BUF1 (N106, N57);
xor XOR2 (N107, N97, N13);
buf BUF1 (N108, N93);
buf BUF1 (N109, N104);
nand NAND4 (N110, N101, N101, N41, N65);
nor NOR4 (N111, N95, N62, N68, N31);
nor NOR3 (N112, N99, N105, N43);
xor XOR2 (N113, N68, N31);
and AND4 (N114, N109, N100, N63, N5);
nor NOR4 (N115, N60, N58, N113, N52);
and AND2 (N116, N113, N10);
nor NOR3 (N117, N112, N21, N24);
buf BUF1 (N118, N108);
xor XOR2 (N119, N110, N16);
or OR3 (N120, N119, N29, N20);
nor NOR3 (N121, N120, N103, N42);
and AND4 (N122, N107, N45, N14, N17);
not NOT1 (N123, N115);
nor NOR3 (N124, N122, N23, N122);
buf BUF1 (N125, N114);
buf BUF1 (N126, N117);
nand NAND3 (N127, N106, N32, N23);
and AND2 (N128, N92, N114);
or OR2 (N129, N125, N62);
buf BUF1 (N130, N129);
buf BUF1 (N131, N126);
and AND4 (N132, N127, N42, N34, N58);
buf BUF1 (N133, N123);
not NOT1 (N134, N116);
not NOT1 (N135, N121);
nor NOR4 (N136, N124, N7, N27, N80);
and AND4 (N137, N136, N58, N110, N24);
nand NAND3 (N138, N137, N90, N74);
buf BUF1 (N139, N133);
nand NAND2 (N140, N139, N38);
xor XOR2 (N141, N131, N102);
buf BUF1 (N142, N111);
buf BUF1 (N143, N118);
and AND2 (N144, N128, N128);
and AND4 (N145, N141, N130, N87, N123);
buf BUF1 (N146, N30);
nor NOR4 (N147, N140, N9, N132, N31);
nor NOR3 (N148, N58, N35, N6);
and AND4 (N149, N135, N139, N55, N79);
nor NOR2 (N150, N134, N50);
buf BUF1 (N151, N142);
and AND2 (N152, N149, N103);
buf BUF1 (N153, N147);
not NOT1 (N154, N145);
not NOT1 (N155, N148);
or OR2 (N156, N155, N111);
not NOT1 (N157, N144);
xor XOR2 (N158, N157, N51);
or OR4 (N159, N143, N10, N47, N15);
and AND3 (N160, N138, N61, N94);
xor XOR2 (N161, N153, N76);
not NOT1 (N162, N152);
buf BUF1 (N163, N154);
nor NOR4 (N164, N158, N44, N99, N40);
nand NAND3 (N165, N164, N144, N90);
not NOT1 (N166, N151);
nand NAND2 (N167, N166, N92);
and AND4 (N168, N165, N139, N118, N105);
buf BUF1 (N169, N150);
nor NOR3 (N170, N159, N9, N36);
or OR2 (N171, N168, N145);
and AND2 (N172, N170, N54);
not NOT1 (N173, N146);
or OR4 (N174, N160, N163, N89, N42);
buf BUF1 (N175, N163);
xor XOR2 (N176, N172, N17);
nand NAND4 (N177, N167, N40, N31, N50);
nor NOR3 (N178, N169, N110, N151);
nor NOR4 (N179, N177, N146, N125, N55);
xor XOR2 (N180, N156, N41);
xor XOR2 (N181, N171, N128);
and AND2 (N182, N176, N53);
buf BUF1 (N183, N162);
not NOT1 (N184, N180);
or OR2 (N185, N161, N155);
nor NOR4 (N186, N185, N41, N114, N128);
xor XOR2 (N187, N179, N80);
nor NOR2 (N188, N174, N24);
xor XOR2 (N189, N173, N47);
buf BUF1 (N190, N184);
or OR3 (N191, N189, N127, N45);
nor NOR4 (N192, N181, N44, N102, N11);
buf BUF1 (N193, N182);
xor XOR2 (N194, N192, N103);
or OR3 (N195, N178, N171, N74);
not NOT1 (N196, N188);
nor NOR3 (N197, N186, N77, N178);
not NOT1 (N198, N195);
not NOT1 (N199, N187);
xor XOR2 (N200, N198, N13);
nor NOR3 (N201, N183, N101, N167);
and AND2 (N202, N199, N39);
and AND2 (N203, N193, N62);
not NOT1 (N204, N197);
or OR4 (N205, N190, N152, N168, N78);
or OR3 (N206, N191, N201, N191);
not NOT1 (N207, N77);
nand NAND3 (N208, N175, N165, N186);
nand NAND2 (N209, N203, N62);
or OR4 (N210, N206, N145, N6, N94);
nand NAND2 (N211, N209, N9);
and AND4 (N212, N200, N87, N118, N124);
buf BUF1 (N213, N207);
xor XOR2 (N214, N204, N78);
nor NOR2 (N215, N213, N132);
nand NAND3 (N216, N202, N73, N146);
buf BUF1 (N217, N214);
and AND2 (N218, N217, N16);
xor XOR2 (N219, N210, N43);
and AND4 (N220, N216, N44, N172, N96);
nand NAND2 (N221, N218, N74);
not NOT1 (N222, N211);
not NOT1 (N223, N220);
buf BUF1 (N224, N208);
nor NOR3 (N225, N212, N102, N14);
or OR3 (N226, N196, N140, N86);
and AND3 (N227, N221, N30, N210);
not NOT1 (N228, N222);
buf BUF1 (N229, N226);
or OR3 (N230, N224, N4, N29);
or OR2 (N231, N223, N212);
or OR2 (N232, N225, N205);
nand NAND4 (N233, N216, N24, N77, N173);
nand NAND3 (N234, N229, N224, N14);
not NOT1 (N235, N232);
nand NAND2 (N236, N227, N164);
nor NOR3 (N237, N194, N100, N24);
and AND4 (N238, N219, N154, N215, N173);
and AND3 (N239, N191, N42, N121);
and AND4 (N240, N233, N168, N224, N43);
buf BUF1 (N241, N234);
xor XOR2 (N242, N237, N83);
xor XOR2 (N243, N236, N123);
or OR2 (N244, N242, N8);
nor NOR2 (N245, N244, N199);
not NOT1 (N246, N245);
buf BUF1 (N247, N239);
or OR4 (N248, N235, N86, N225, N214);
or OR3 (N249, N238, N162, N47);
nor NOR4 (N250, N247, N217, N226, N156);
buf BUF1 (N251, N246);
not NOT1 (N252, N250);
and AND2 (N253, N240, N181);
not NOT1 (N254, N248);
xor XOR2 (N255, N253, N135);
nand NAND3 (N256, N228, N165, N22);
xor XOR2 (N257, N255, N95);
nor NOR4 (N258, N249, N31, N57, N14);
and AND3 (N259, N241, N46, N58);
not NOT1 (N260, N258);
nor NOR3 (N261, N256, N116, N256);
or OR3 (N262, N231, N213, N160);
buf BUF1 (N263, N251);
nand NAND3 (N264, N260, N195, N75);
nor NOR4 (N265, N230, N203, N67, N73);
or OR2 (N266, N252, N11);
nor NOR4 (N267, N259, N153, N216, N184);
buf BUF1 (N268, N262);
nor NOR3 (N269, N264, N29, N81);
nor NOR2 (N270, N267, N212);
nand NAND2 (N271, N268, N136);
or OR4 (N272, N266, N230, N7, N229);
buf BUF1 (N273, N270);
or OR4 (N274, N272, N108, N88, N42);
nand NAND4 (N275, N265, N264, N204, N195);
xor XOR2 (N276, N263, N78);
buf BUF1 (N277, N271);
or OR4 (N278, N275, N221, N62, N105);
or OR3 (N279, N243, N183, N173);
nand NAND3 (N280, N279, N169, N95);
xor XOR2 (N281, N261, N223);
buf BUF1 (N282, N277);
nand NAND3 (N283, N281, N114, N108);
nand NAND3 (N284, N257, N152, N27);
not NOT1 (N285, N269);
nor NOR2 (N286, N280, N72);
not NOT1 (N287, N278);
buf BUF1 (N288, N276);
not NOT1 (N289, N274);
nor NOR3 (N290, N287, N163, N240);
xor XOR2 (N291, N286, N121);
and AND3 (N292, N283, N146, N180);
xor XOR2 (N293, N284, N79);
nand NAND2 (N294, N273, N126);
nand NAND3 (N295, N292, N180, N77);
and AND3 (N296, N254, N39, N277);
not NOT1 (N297, N294);
buf BUF1 (N298, N297);
nor NOR4 (N299, N282, N269, N150, N143);
not NOT1 (N300, N289);
nor NOR4 (N301, N296, N277, N263, N259);
buf BUF1 (N302, N299);
not NOT1 (N303, N291);
or OR3 (N304, N300, N287, N236);
not NOT1 (N305, N290);
not NOT1 (N306, N285);
and AND4 (N307, N305, N43, N55, N244);
nor NOR2 (N308, N288, N201);
nand NAND4 (N309, N308, N241, N167, N94);
nand NAND4 (N310, N307, N111, N85, N99);
and AND4 (N311, N310, N126, N176, N310);
and AND2 (N312, N301, N195);
nor NOR3 (N313, N293, N307, N291);
or OR2 (N314, N295, N67);
not NOT1 (N315, N311);
and AND4 (N316, N314, N189, N293, N39);
or OR2 (N317, N306, N22);
buf BUF1 (N318, N315);
nand NAND2 (N319, N303, N51);
not NOT1 (N320, N319);
not NOT1 (N321, N309);
xor XOR2 (N322, N320, N81);
nor NOR4 (N323, N317, N193, N252, N37);
and AND3 (N324, N313, N239, N190);
buf BUF1 (N325, N312);
nor NOR4 (N326, N318, N219, N165, N318);
or OR2 (N327, N302, N20);
buf BUF1 (N328, N304);
and AND4 (N329, N326, N44, N297, N148);
nand NAND2 (N330, N328, N150);
buf BUF1 (N331, N298);
xor XOR2 (N332, N327, N213);
or OR4 (N333, N323, N144, N176, N182);
and AND3 (N334, N322, N275, N159);
buf BUF1 (N335, N316);
xor XOR2 (N336, N321, N286);
not NOT1 (N337, N336);
buf BUF1 (N338, N324);
nor NOR3 (N339, N331, N306, N237);
buf BUF1 (N340, N332);
and AND2 (N341, N333, N175);
nand NAND4 (N342, N329, N311, N197, N119);
xor XOR2 (N343, N334, N220);
buf BUF1 (N344, N341);
buf BUF1 (N345, N338);
nor NOR3 (N346, N337, N62, N210);
buf BUF1 (N347, N345);
nor NOR2 (N348, N335, N108);
buf BUF1 (N349, N343);
nor NOR3 (N350, N339, N304, N347);
not NOT1 (N351, N335);
xor XOR2 (N352, N348, N105);
buf BUF1 (N353, N351);
not NOT1 (N354, N342);
nor NOR3 (N355, N350, N317, N153);
nand NAND3 (N356, N354, N268, N287);
nand NAND2 (N357, N353, N128);
buf BUF1 (N358, N349);
nand NAND3 (N359, N344, N236, N21);
nand NAND4 (N360, N340, N82, N70, N140);
not NOT1 (N361, N325);
not NOT1 (N362, N358);
and AND3 (N363, N352, N135, N358);
buf BUF1 (N364, N361);
nor NOR2 (N365, N363, N228);
or OR4 (N366, N346, N145, N55, N91);
nor NOR2 (N367, N330, N233);
buf BUF1 (N368, N367);
buf BUF1 (N369, N368);
not NOT1 (N370, N359);
buf BUF1 (N371, N357);
xor XOR2 (N372, N356, N234);
nand NAND3 (N373, N366, N362, N291);
nor NOR4 (N374, N163, N138, N130, N91);
buf BUF1 (N375, N369);
xor XOR2 (N376, N365, N216);
nor NOR4 (N377, N372, N15, N50, N366);
and AND3 (N378, N377, N253, N370);
and AND4 (N379, N362, N24, N78, N277);
not NOT1 (N380, N378);
nor NOR3 (N381, N375, N28, N32);
xor XOR2 (N382, N376, N360);
buf BUF1 (N383, N352);
not NOT1 (N384, N355);
nand NAND2 (N385, N364, N97);
and AND2 (N386, N374, N250);
or OR3 (N387, N386, N79, N230);
xor XOR2 (N388, N380, N225);
and AND4 (N389, N387, N108, N58, N191);
buf BUF1 (N390, N382);
nand NAND4 (N391, N385, N14, N175, N236);
nor NOR3 (N392, N391, N289, N297);
nor NOR4 (N393, N381, N229, N60, N105);
or OR3 (N394, N390, N265, N209);
nor NOR2 (N395, N392, N390);
xor XOR2 (N396, N373, N13);
nor NOR3 (N397, N395, N45, N196);
not NOT1 (N398, N397);
and AND2 (N399, N383, N290);
nor NOR3 (N400, N388, N218, N207);
xor XOR2 (N401, N393, N114);
not NOT1 (N402, N384);
not NOT1 (N403, N401);
nand NAND4 (N404, N398, N194, N360, N89);
or OR4 (N405, N396, N87, N325, N53);
xor XOR2 (N406, N405, N147);
nand NAND3 (N407, N404, N332, N403);
nor NOR4 (N408, N405, N176, N229, N208);
nand NAND3 (N409, N407, N402, N388);
and AND3 (N410, N249, N288, N232);
buf BUF1 (N411, N389);
nand NAND3 (N412, N411, N203, N125);
or OR4 (N413, N379, N141, N277, N399);
nor NOR2 (N414, N360, N252);
nand NAND2 (N415, N413, N125);
buf BUF1 (N416, N410);
or OR2 (N417, N409, N339);
nor NOR2 (N418, N400, N78);
or OR4 (N419, N406, N177, N354, N348);
or OR4 (N420, N418, N249, N313, N285);
xor XOR2 (N421, N412, N285);
xor XOR2 (N422, N394, N361);
nor NOR3 (N423, N415, N250, N326);
and AND4 (N424, N371, N245, N317, N334);
xor XOR2 (N425, N421, N147);
nor NOR4 (N426, N425, N330, N10, N52);
buf BUF1 (N427, N417);
and AND3 (N428, N414, N46, N71);
buf BUF1 (N429, N426);
or OR4 (N430, N424, N188, N86, N301);
buf BUF1 (N431, N428);
nor NOR4 (N432, N416, N38, N34, N373);
or OR3 (N433, N430, N186, N327);
xor XOR2 (N434, N422, N298);
and AND3 (N435, N431, N394, N260);
xor XOR2 (N436, N420, N95);
not NOT1 (N437, N423);
and AND2 (N438, N436, N222);
or OR3 (N439, N433, N239, N98);
and AND4 (N440, N427, N410, N424, N180);
xor XOR2 (N441, N408, N409);
buf BUF1 (N442, N432);
and AND3 (N443, N439, N281, N232);
xor XOR2 (N444, N440, N183);
not NOT1 (N445, N442);
or OR4 (N446, N437, N23, N407, N349);
nor NOR2 (N447, N429, N132);
buf BUF1 (N448, N434);
not NOT1 (N449, N446);
buf BUF1 (N450, N447);
buf BUF1 (N451, N449);
and AND3 (N452, N445, N346, N406);
buf BUF1 (N453, N444);
nor NOR3 (N454, N452, N419, N435);
nor NOR3 (N455, N449, N454, N12);
and AND4 (N456, N316, N123, N287, N270);
not NOT1 (N457, N388);
or OR4 (N458, N456, N312, N240, N265);
nor NOR2 (N459, N448, N54);
or OR3 (N460, N453, N200, N68);
or OR3 (N461, N451, N366, N39);
not NOT1 (N462, N458);
and AND2 (N463, N459, N52);
xor XOR2 (N464, N455, N10);
nor NOR3 (N465, N438, N103, N78);
nor NOR4 (N466, N465, N240, N371, N201);
nor NOR3 (N467, N460, N41, N82);
not NOT1 (N468, N466);
nor NOR4 (N469, N462, N6, N465, N157);
and AND4 (N470, N467, N196, N220, N24);
xor XOR2 (N471, N468, N150);
not NOT1 (N472, N450);
not NOT1 (N473, N461);
nor NOR3 (N474, N463, N216, N298);
or OR4 (N475, N470, N452, N225, N180);
or OR4 (N476, N472, N84, N164, N195);
nand NAND3 (N477, N471, N324, N224);
nand NAND4 (N478, N476, N238, N138, N235);
nand NAND4 (N479, N443, N386, N359, N31);
nand NAND2 (N480, N479, N345);
nand NAND2 (N481, N478, N137);
not NOT1 (N482, N481);
nand NAND3 (N483, N469, N441, N253);
nor NOR2 (N484, N34, N305);
not NOT1 (N485, N477);
xor XOR2 (N486, N457, N478);
nand NAND3 (N487, N480, N338, N239);
nor NOR2 (N488, N485, N69);
not NOT1 (N489, N475);
xor XOR2 (N490, N474, N444);
nor NOR3 (N491, N488, N111, N419);
not NOT1 (N492, N473);
xor XOR2 (N493, N487, N282);
and AND3 (N494, N492, N306, N152);
nor NOR3 (N495, N484, N122, N452);
not NOT1 (N496, N489);
buf BUF1 (N497, N490);
nor NOR2 (N498, N495, N458);
buf BUF1 (N499, N493);
nor NOR3 (N500, N464, N5, N384);
or OR3 (N501, N483, N232, N392);
nor NOR3 (N502, N491, N198, N217);
and AND3 (N503, N502, N383, N462);
and AND2 (N504, N486, N127);
buf BUF1 (N505, N501);
nand NAND2 (N506, N505, N52);
and AND2 (N507, N500, N32);
xor XOR2 (N508, N504, N418);
buf BUF1 (N509, N499);
and AND2 (N510, N509, N378);
and AND2 (N511, N510, N506);
nand NAND2 (N512, N394, N64);
xor XOR2 (N513, N494, N304);
nor NOR2 (N514, N507, N127);
or OR2 (N515, N496, N299);
xor XOR2 (N516, N511, N52);
nor NOR3 (N517, N498, N230, N393);
buf BUF1 (N518, N482);
xor XOR2 (N519, N512, N28);
nand NAND4 (N520, N519, N366, N288, N471);
buf BUF1 (N521, N514);
nand NAND2 (N522, N521, N429);
nor NOR3 (N523, N503, N15, N270);
xor XOR2 (N524, N508, N485);
nand NAND4 (N525, N497, N387, N419, N257);
xor XOR2 (N526, N523, N146);
not NOT1 (N527, N516);
nor NOR2 (N528, N517, N284);
nand NAND4 (N529, N526, N89, N286, N189);
nor NOR4 (N530, N525, N286, N455, N191);
buf BUF1 (N531, N528);
xor XOR2 (N532, N522, N401);
or OR3 (N533, N532, N394, N87);
xor XOR2 (N534, N533, N361);
or OR4 (N535, N513, N83, N269, N90);
buf BUF1 (N536, N530);
and AND4 (N537, N534, N401, N112, N198);
xor XOR2 (N538, N531, N276);
or OR2 (N539, N527, N121);
or OR2 (N540, N536, N414);
xor XOR2 (N541, N515, N289);
and AND3 (N542, N540, N520, N72);
nand NAND2 (N543, N537, N472);
nor NOR3 (N544, N459, N531, N233);
xor XOR2 (N545, N518, N335);
and AND2 (N546, N535, N62);
or OR3 (N547, N524, N90, N190);
xor XOR2 (N548, N539, N526);
buf BUF1 (N549, N544);
buf BUF1 (N550, N543);
xor XOR2 (N551, N550, N159);
nand NAND4 (N552, N551, N23, N373, N476);
or OR3 (N553, N549, N88, N546);
buf BUF1 (N554, N364);
nand NAND4 (N555, N529, N321, N95, N429);
xor XOR2 (N556, N545, N272);
buf BUF1 (N557, N556);
or OR4 (N558, N548, N419, N547, N295);
xor XOR2 (N559, N148, N317);
or OR2 (N560, N542, N61);
nor NOR2 (N561, N541, N279);
not NOT1 (N562, N555);
not NOT1 (N563, N558);
and AND2 (N564, N554, N518);
not NOT1 (N565, N563);
not NOT1 (N566, N553);
not NOT1 (N567, N538);
or OR3 (N568, N562, N516, N397);
or OR2 (N569, N559, N531);
nor NOR3 (N570, N560, N371, N526);
buf BUF1 (N571, N569);
or OR4 (N572, N561, N473, N344, N511);
and AND4 (N573, N565, N456, N201, N79);
buf BUF1 (N574, N566);
and AND3 (N575, N564, N128, N280);
and AND3 (N576, N557, N251, N429);
not NOT1 (N577, N568);
or OR3 (N578, N576, N148, N367);
or OR2 (N579, N578, N466);
nor NOR4 (N580, N572, N69, N59, N513);
and AND2 (N581, N577, N529);
nand NAND2 (N582, N581, N220);
buf BUF1 (N583, N582);
nor NOR4 (N584, N552, N480, N289, N43);
nor NOR3 (N585, N580, N133, N539);
and AND3 (N586, N567, N21, N297);
nor NOR2 (N587, N585, N553);
nand NAND2 (N588, N573, N39);
nor NOR2 (N589, N579, N398);
buf BUF1 (N590, N571);
buf BUF1 (N591, N588);
xor XOR2 (N592, N575, N249);
or OR2 (N593, N574, N495);
xor XOR2 (N594, N591, N84);
not NOT1 (N595, N587);
or OR2 (N596, N595, N485);
not NOT1 (N597, N584);
and AND4 (N598, N589, N28, N47, N304);
and AND2 (N599, N590, N493);
buf BUF1 (N600, N596);
buf BUF1 (N601, N586);
xor XOR2 (N602, N593, N404);
or OR3 (N603, N600, N96, N120);
nor NOR4 (N604, N592, N397, N104, N157);
nor NOR3 (N605, N598, N65, N261);
or OR4 (N606, N602, N279, N519, N566);
buf BUF1 (N607, N605);
and AND2 (N608, N594, N466);
nor NOR4 (N609, N583, N397, N541, N222);
not NOT1 (N610, N597);
and AND4 (N611, N601, N485, N492, N346);
nor NOR3 (N612, N608, N518, N75);
or OR3 (N613, N609, N252, N313);
nand NAND2 (N614, N603, N336);
buf BUF1 (N615, N613);
or OR4 (N616, N606, N452, N555, N297);
or OR3 (N617, N607, N273, N187);
not NOT1 (N618, N604);
xor XOR2 (N619, N599, N460);
or OR2 (N620, N617, N23);
xor XOR2 (N621, N618, N186);
xor XOR2 (N622, N614, N328);
or OR4 (N623, N611, N30, N50, N244);
or OR3 (N624, N616, N259, N496);
buf BUF1 (N625, N620);
and AND3 (N626, N624, N33, N490);
buf BUF1 (N627, N612);
nor NOR4 (N628, N627, N106, N133, N502);
or OR3 (N629, N628, N443, N157);
not NOT1 (N630, N610);
nand NAND2 (N631, N619, N480);
nand NAND2 (N632, N629, N83);
or OR2 (N633, N621, N338);
nand NAND4 (N634, N632, N47, N87, N337);
nand NAND2 (N635, N630, N623);
nand NAND3 (N636, N69, N456, N437);
xor XOR2 (N637, N625, N631);
nand NAND3 (N638, N464, N37, N200);
nand NAND4 (N639, N622, N219, N416, N154);
or OR2 (N640, N637, N573);
nand NAND2 (N641, N639, N271);
not NOT1 (N642, N640);
buf BUF1 (N643, N641);
xor XOR2 (N644, N635, N547);
nand NAND2 (N645, N644, N436);
buf BUF1 (N646, N570);
nor NOR4 (N647, N636, N592, N262, N135);
nand NAND2 (N648, N634, N226);
not NOT1 (N649, N647);
xor XOR2 (N650, N649, N4);
buf BUF1 (N651, N648);
or OR2 (N652, N651, N650);
and AND4 (N653, N338, N61, N31, N381);
nor NOR2 (N654, N645, N343);
or OR4 (N655, N633, N287, N483, N595);
not NOT1 (N656, N654);
or OR4 (N657, N646, N291, N333, N411);
not NOT1 (N658, N642);
or OR3 (N659, N657, N332, N251);
or OR4 (N660, N655, N323, N449, N604);
not NOT1 (N661, N653);
buf BUF1 (N662, N656);
xor XOR2 (N663, N652, N605);
buf BUF1 (N664, N658);
buf BUF1 (N665, N659);
or OR3 (N666, N660, N504, N588);
nand NAND2 (N667, N662, N310);
not NOT1 (N668, N667);
buf BUF1 (N669, N666);
buf BUF1 (N670, N668);
buf BUF1 (N671, N665);
nand NAND4 (N672, N643, N254, N503, N88);
buf BUF1 (N673, N671);
or OR3 (N674, N638, N300, N108);
and AND4 (N675, N661, N475, N236, N577);
nor NOR3 (N676, N673, N282, N175);
and AND4 (N677, N670, N266, N203, N167);
xor XOR2 (N678, N672, N110);
not NOT1 (N679, N677);
xor XOR2 (N680, N678, N123);
xor XOR2 (N681, N676, N493);
not NOT1 (N682, N663);
nor NOR2 (N683, N680, N590);
not NOT1 (N684, N682);
and AND4 (N685, N675, N619, N115, N77);
nand NAND4 (N686, N674, N114, N562, N450);
buf BUF1 (N687, N683);
nor NOR2 (N688, N681, N216);
buf BUF1 (N689, N686);
buf BUF1 (N690, N685);
nor NOR3 (N691, N626, N390, N142);
nand NAND4 (N692, N689, N121, N151, N678);
or OR3 (N693, N669, N478, N205);
nand NAND2 (N694, N684, N222);
and AND2 (N695, N694, N523);
nor NOR4 (N696, N688, N274, N335, N595);
buf BUF1 (N697, N664);
nand NAND3 (N698, N696, N89, N347);
or OR2 (N699, N687, N560);
nand NAND3 (N700, N692, N120, N347);
buf BUF1 (N701, N690);
nand NAND3 (N702, N698, N132, N352);
and AND4 (N703, N697, N651, N273, N352);
or OR3 (N704, N699, N304, N397);
buf BUF1 (N705, N703);
nand NAND4 (N706, N695, N245, N574, N249);
xor XOR2 (N707, N706, N557);
xor XOR2 (N708, N704, N643);
or OR4 (N709, N701, N226, N538, N147);
nor NOR3 (N710, N691, N635, N404);
nand NAND3 (N711, N693, N664, N46);
or OR2 (N712, N702, N401);
buf BUF1 (N713, N707);
and AND4 (N714, N710, N339, N219, N33);
or OR3 (N715, N708, N628, N3);
and AND4 (N716, N712, N490, N23, N388);
buf BUF1 (N717, N679);
or OR2 (N718, N709, N300);
not NOT1 (N719, N717);
and AND4 (N720, N615, N202, N146, N182);
not NOT1 (N721, N718);
and AND2 (N722, N720, N299);
buf BUF1 (N723, N716);
buf BUF1 (N724, N721);
not NOT1 (N725, N722);
and AND3 (N726, N725, N617, N157);
xor XOR2 (N727, N719, N674);
nor NOR3 (N728, N705, N674, N691);
and AND4 (N729, N700, N419, N612, N538);
xor XOR2 (N730, N723, N371);
nand NAND4 (N731, N730, N194, N36, N179);
buf BUF1 (N732, N728);
xor XOR2 (N733, N715, N279);
buf BUF1 (N734, N733);
nand NAND2 (N735, N727, N337);
nor NOR4 (N736, N724, N667, N632, N309);
nand NAND2 (N737, N734, N442);
nand NAND2 (N738, N714, N139);
and AND4 (N739, N736, N62, N624, N52);
xor XOR2 (N740, N738, N22);
buf BUF1 (N741, N735);
or OR2 (N742, N732, N706);
or OR3 (N743, N740, N269, N89);
nor NOR3 (N744, N713, N528, N659);
and AND4 (N745, N731, N531, N267, N573);
xor XOR2 (N746, N737, N700);
buf BUF1 (N747, N726);
or OR3 (N748, N747, N584, N392);
buf BUF1 (N749, N748);
nor NOR3 (N750, N746, N491, N590);
and AND4 (N751, N750, N463, N497, N342);
nor NOR2 (N752, N745, N354);
xor XOR2 (N753, N744, N606);
xor XOR2 (N754, N711, N524);
nand NAND2 (N755, N739, N624);
and AND4 (N756, N751, N663, N29, N188);
or OR3 (N757, N754, N540, N457);
not NOT1 (N758, N756);
or OR3 (N759, N742, N680, N88);
nor NOR2 (N760, N743, N218);
and AND2 (N761, N741, N129);
and AND3 (N762, N758, N560, N528);
not NOT1 (N763, N762);
or OR4 (N764, N753, N205, N357, N120);
buf BUF1 (N765, N761);
and AND4 (N766, N749, N311, N580, N137);
nand NAND2 (N767, N755, N156);
buf BUF1 (N768, N752);
not NOT1 (N769, N757);
not NOT1 (N770, N769);
and AND3 (N771, N770, N414, N421);
and AND2 (N772, N771, N573);
not NOT1 (N773, N772);
xor XOR2 (N774, N763, N458);
nor NOR4 (N775, N760, N420, N714, N159);
and AND2 (N776, N765, N94);
not NOT1 (N777, N764);
nand NAND3 (N778, N767, N410, N607);
nand NAND4 (N779, N766, N770, N250, N320);
nor NOR2 (N780, N768, N572);
nand NAND3 (N781, N778, N519, N135);
nor NOR4 (N782, N729, N306, N764, N320);
or OR2 (N783, N779, N623);
not NOT1 (N784, N780);
buf BUF1 (N785, N759);
nor NOR4 (N786, N784, N525, N80, N566);
nor NOR4 (N787, N786, N184, N645, N490);
xor XOR2 (N788, N785, N45);
not NOT1 (N789, N773);
nand NAND3 (N790, N777, N298, N544);
buf BUF1 (N791, N788);
buf BUF1 (N792, N783);
nand NAND4 (N793, N775, N561, N330, N346);
xor XOR2 (N794, N790, N92);
or OR4 (N795, N787, N375, N737, N390);
nor NOR2 (N796, N793, N587);
not NOT1 (N797, N782);
xor XOR2 (N798, N794, N178);
or OR4 (N799, N798, N715, N177, N226);
nor NOR2 (N800, N791, N798);
and AND2 (N801, N796, N750);
nor NOR4 (N802, N801, N786, N8, N264);
or OR3 (N803, N799, N149, N289);
not NOT1 (N804, N792);
xor XOR2 (N805, N789, N95);
buf BUF1 (N806, N804);
and AND2 (N807, N797, N523);
buf BUF1 (N808, N802);
not NOT1 (N809, N781);
nand NAND3 (N810, N774, N589, N445);
xor XOR2 (N811, N776, N485);
nand NAND2 (N812, N807, N605);
not NOT1 (N813, N812);
xor XOR2 (N814, N803, N789);
nor NOR3 (N815, N800, N488, N813);
xor XOR2 (N816, N149, N727);
nor NOR2 (N817, N810, N110);
buf BUF1 (N818, N815);
and AND3 (N819, N805, N150, N191);
xor XOR2 (N820, N817, N620);
and AND4 (N821, N814, N397, N406, N338);
nand NAND4 (N822, N821, N60, N245, N237);
nand NAND2 (N823, N811, N406);
xor XOR2 (N824, N823, N4);
not NOT1 (N825, N818);
not NOT1 (N826, N824);
not NOT1 (N827, N819);
buf BUF1 (N828, N825);
not NOT1 (N829, N822);
or OR4 (N830, N826, N605, N471, N786);
buf BUF1 (N831, N827);
buf BUF1 (N832, N808);
not NOT1 (N833, N830);
nand NAND3 (N834, N833, N559, N221);
buf BUF1 (N835, N809);
xor XOR2 (N836, N835, N279);
nor NOR4 (N837, N836, N503, N219, N357);
and AND3 (N838, N832, N509, N373);
xor XOR2 (N839, N795, N750);
or OR2 (N840, N820, N474);
nand NAND4 (N841, N816, N560, N514, N68);
nand NAND3 (N842, N829, N645, N452);
xor XOR2 (N843, N806, N305);
or OR4 (N844, N834, N701, N305, N105);
buf BUF1 (N845, N839);
xor XOR2 (N846, N845, N590);
or OR4 (N847, N838, N517, N459, N730);
or OR3 (N848, N840, N505, N547);
and AND4 (N849, N841, N651, N775, N467);
not NOT1 (N850, N837);
xor XOR2 (N851, N843, N364);
nand NAND4 (N852, N850, N332, N207, N742);
xor XOR2 (N853, N848, N785);
or OR3 (N854, N847, N719, N509);
nand NAND3 (N855, N842, N172, N198);
buf BUF1 (N856, N844);
buf BUF1 (N857, N852);
nor NOR2 (N858, N857, N387);
buf BUF1 (N859, N853);
nand NAND3 (N860, N851, N305, N742);
nor NOR4 (N861, N855, N435, N432, N660);
nand NAND2 (N862, N846, N202);
or OR2 (N863, N854, N460);
not NOT1 (N864, N856);
or OR2 (N865, N831, N114);
nand NAND2 (N866, N865, N5);
nor NOR4 (N867, N861, N428, N363, N729);
and AND3 (N868, N863, N770, N687);
nor NOR4 (N869, N849, N40, N340, N90);
not NOT1 (N870, N858);
buf BUF1 (N871, N862);
or OR2 (N872, N866, N103);
not NOT1 (N873, N868);
and AND3 (N874, N867, N792, N622);
nor NOR4 (N875, N870, N617, N838, N835);
or OR3 (N876, N869, N290, N447);
not NOT1 (N877, N864);
not NOT1 (N878, N860);
buf BUF1 (N879, N872);
or OR3 (N880, N876, N317, N225);
xor XOR2 (N881, N875, N58);
nor NOR3 (N882, N880, N466, N346);
buf BUF1 (N883, N874);
not NOT1 (N884, N883);
or OR3 (N885, N879, N255, N485);
buf BUF1 (N886, N878);
not NOT1 (N887, N882);
and AND2 (N888, N886, N216);
buf BUF1 (N889, N881);
buf BUF1 (N890, N887);
buf BUF1 (N891, N889);
and AND3 (N892, N890, N333, N797);
nand NAND2 (N893, N891, N117);
and AND4 (N894, N885, N237, N108, N819);
or OR3 (N895, N893, N818, N870);
nand NAND4 (N896, N828, N32, N422, N251);
xor XOR2 (N897, N894, N442);
nand NAND4 (N898, N877, N851, N268, N4);
and AND3 (N899, N896, N474, N470);
nor NOR3 (N900, N899, N477, N101);
and AND2 (N901, N897, N481);
nand NAND3 (N902, N859, N100, N334);
or OR4 (N903, N901, N863, N499, N740);
not NOT1 (N904, N873);
xor XOR2 (N905, N902, N13);
or OR4 (N906, N888, N830, N267, N675);
or OR2 (N907, N906, N593);
or OR3 (N908, N905, N475, N565);
and AND4 (N909, N900, N901, N611, N494);
buf BUF1 (N910, N909);
nor NOR2 (N911, N904, N428);
nand NAND3 (N912, N908, N677, N814);
buf BUF1 (N913, N907);
and AND4 (N914, N912, N846, N405, N532);
buf BUF1 (N915, N884);
and AND2 (N916, N913, N250);
and AND2 (N917, N914, N723);
nor NOR2 (N918, N892, N741);
nand NAND2 (N919, N910, N16);
nand NAND2 (N920, N915, N591);
nand NAND4 (N921, N911, N48, N84, N799);
or OR3 (N922, N918, N481, N525);
or OR3 (N923, N895, N511, N238);
not NOT1 (N924, N920);
not NOT1 (N925, N917);
buf BUF1 (N926, N898);
or OR4 (N927, N871, N508, N214, N902);
buf BUF1 (N928, N903);
not NOT1 (N929, N928);
not NOT1 (N930, N927);
nand NAND2 (N931, N921, N235);
buf BUF1 (N932, N924);
or OR3 (N933, N926, N465, N166);
and AND4 (N934, N922, N473, N26, N656);
and AND3 (N935, N934, N756, N407);
and AND3 (N936, N930, N60, N131);
or OR2 (N937, N932, N268);
xor XOR2 (N938, N916, N928);
nand NAND2 (N939, N938, N501);
and AND4 (N940, N931, N539, N253, N517);
or OR4 (N941, N919, N903, N672, N468);
or OR2 (N942, N936, N920);
nor NOR2 (N943, N925, N873);
not NOT1 (N944, N941);
xor XOR2 (N945, N923, N78);
and AND4 (N946, N933, N703, N92, N314);
xor XOR2 (N947, N942, N295);
not NOT1 (N948, N940);
xor XOR2 (N949, N945, N154);
xor XOR2 (N950, N929, N539);
xor XOR2 (N951, N949, N481);
nand NAND2 (N952, N939, N372);
not NOT1 (N953, N948);
and AND2 (N954, N947, N633);
nand NAND2 (N955, N943, N314);
nand NAND3 (N956, N937, N269, N659);
nand NAND3 (N957, N950, N952, N50);
xor XOR2 (N958, N395, N878);
xor XOR2 (N959, N935, N76);
or OR4 (N960, N954, N662, N950, N141);
nand NAND2 (N961, N944, N892);
nand NAND3 (N962, N961, N129, N406);
nor NOR2 (N963, N960, N662);
xor XOR2 (N964, N955, N421);
nor NOR4 (N965, N946, N25, N414, N799);
buf BUF1 (N966, N963);
not NOT1 (N967, N959);
nor NOR4 (N968, N953, N703, N916, N257);
or OR4 (N969, N967, N248, N300, N32);
xor XOR2 (N970, N962, N253);
not NOT1 (N971, N958);
not NOT1 (N972, N971);
nor NOR2 (N973, N966, N193);
and AND2 (N974, N957, N731);
not NOT1 (N975, N972);
nand NAND4 (N976, N968, N940, N168, N855);
xor XOR2 (N977, N951, N419);
nand NAND2 (N978, N964, N248);
nand NAND4 (N979, N976, N508, N837, N912);
buf BUF1 (N980, N975);
buf BUF1 (N981, N973);
nor NOR4 (N982, N970, N370, N812, N257);
nor NOR4 (N983, N969, N521, N598, N81);
nand NAND2 (N984, N965, N131);
nand NAND4 (N985, N979, N897, N626, N438);
nand NAND4 (N986, N982, N725, N81, N888);
xor XOR2 (N987, N985, N644);
and AND3 (N988, N956, N133, N530);
and AND4 (N989, N988, N846, N392, N277);
and AND4 (N990, N974, N741, N478, N656);
or OR2 (N991, N978, N696);
nand NAND2 (N992, N984, N761);
nor NOR2 (N993, N981, N144);
not NOT1 (N994, N980);
or OR4 (N995, N994, N370, N793, N39);
nor NOR3 (N996, N977, N654, N41);
or OR3 (N997, N987, N489, N796);
nor NOR3 (N998, N997, N182, N831);
nand NAND3 (N999, N986, N140, N979);
buf BUF1 (N1000, N991);
nand NAND3 (N1001, N990, N640, N219);
nor NOR4 (N1002, N983, N677, N975, N80);
xor XOR2 (N1003, N1000, N151);
not NOT1 (N1004, N999);
nor NOR2 (N1005, N1001, N407);
buf BUF1 (N1006, N992);
or OR4 (N1007, N1006, N430, N509, N506);
and AND2 (N1008, N995, N602);
buf BUF1 (N1009, N1007);
buf BUF1 (N1010, N989);
or OR4 (N1011, N1009, N915, N97, N501);
xor XOR2 (N1012, N996, N547);
and AND3 (N1013, N993, N328, N645);
buf BUF1 (N1014, N998);
buf BUF1 (N1015, N1010);
xor XOR2 (N1016, N1015, N816);
xor XOR2 (N1017, N1005, N266);
xor XOR2 (N1018, N1013, N904);
nand NAND2 (N1019, N1012, N376);
xor XOR2 (N1020, N1017, N154);
not NOT1 (N1021, N1020);
or OR4 (N1022, N1021, N50, N448, N919);
xor XOR2 (N1023, N1019, N464);
nand NAND2 (N1024, N1016, N100);
nor NOR4 (N1025, N1004, N673, N615, N772);
or OR2 (N1026, N1002, N323);
and AND3 (N1027, N1023, N663, N854);
not NOT1 (N1028, N1026);
or OR2 (N1029, N1003, N440);
and AND2 (N1030, N1024, N831);
nand NAND3 (N1031, N1011, N79, N5);
not NOT1 (N1032, N1008);
xor XOR2 (N1033, N1018, N16);
nand NAND2 (N1034, N1022, N984);
nor NOR3 (N1035, N1034, N589, N689);
nor NOR2 (N1036, N1035, N345);
xor XOR2 (N1037, N1027, N471);
and AND2 (N1038, N1025, N418);
nand NAND4 (N1039, N1030, N626, N973, N909);
nor NOR2 (N1040, N1037, N545);
or OR2 (N1041, N1028, N379);
buf BUF1 (N1042, N1029);
and AND3 (N1043, N1040, N5, N160);
and AND4 (N1044, N1036, N928, N873, N867);
buf BUF1 (N1045, N1031);
and AND4 (N1046, N1042, N504, N769, N75);
not NOT1 (N1047, N1033);
buf BUF1 (N1048, N1038);
and AND4 (N1049, N1046, N42, N1045, N204);
nor NOR3 (N1050, N437, N506, N34);
or OR3 (N1051, N1014, N400, N774);
and AND4 (N1052, N1032, N183, N746, N211);
or OR2 (N1053, N1052, N673);
or OR4 (N1054, N1053, N666, N1050, N802);
not NOT1 (N1055, N234);
nand NAND3 (N1056, N1044, N273, N214);
nor NOR3 (N1057, N1048, N381, N1000);
nand NAND4 (N1058, N1043, N594, N728, N984);
nand NAND2 (N1059, N1054, N65);
and AND2 (N1060, N1057, N432);
nand NAND2 (N1061, N1039, N632);
or OR4 (N1062, N1058, N830, N137, N211);
or OR3 (N1063, N1059, N464, N171);
and AND3 (N1064, N1060, N468, N876);
and AND4 (N1065, N1047, N687, N109, N1030);
buf BUF1 (N1066, N1055);
and AND3 (N1067, N1065, N687, N254);
nand NAND4 (N1068, N1063, N723, N826, N129);
buf BUF1 (N1069, N1056);
or OR2 (N1070, N1049, N1029);
buf BUF1 (N1071, N1041);
or OR2 (N1072, N1069, N927);
xor XOR2 (N1073, N1068, N453);
nand NAND3 (N1074, N1071, N1053, N308);
not NOT1 (N1075, N1064);
nand NAND2 (N1076, N1072, N316);
nand NAND2 (N1077, N1075, N190);
not NOT1 (N1078, N1077);
not NOT1 (N1079, N1074);
not NOT1 (N1080, N1066);
not NOT1 (N1081, N1062);
buf BUF1 (N1082, N1076);
nand NAND3 (N1083, N1080, N811, N741);
nand NAND2 (N1084, N1067, N657);
buf BUF1 (N1085, N1070);
and AND3 (N1086, N1082, N709, N752);
buf BUF1 (N1087, N1051);
buf BUF1 (N1088, N1085);
nand NAND3 (N1089, N1073, N1011, N659);
or OR4 (N1090, N1079, N721, N938, N683);
nor NOR4 (N1091, N1089, N560, N127, N507);
buf BUF1 (N1092, N1090);
buf BUF1 (N1093, N1061);
buf BUF1 (N1094, N1084);
nand NAND3 (N1095, N1088, N54, N617);
xor XOR2 (N1096, N1083, N746);
nor NOR4 (N1097, N1092, N292, N1049, N204);
nand NAND4 (N1098, N1078, N758, N179, N252);
not NOT1 (N1099, N1081);
xor XOR2 (N1100, N1097, N504);
buf BUF1 (N1101, N1087);
and AND2 (N1102, N1094, N542);
xor XOR2 (N1103, N1100, N599);
and AND4 (N1104, N1101, N829, N44, N773);
nand NAND4 (N1105, N1096, N272, N454, N53);
not NOT1 (N1106, N1093);
xor XOR2 (N1107, N1106, N204);
not NOT1 (N1108, N1107);
nand NAND2 (N1109, N1103, N368);
or OR3 (N1110, N1102, N778, N1002);
nand NAND3 (N1111, N1105, N1093, N612);
nand NAND4 (N1112, N1110, N60, N554, N483);
or OR2 (N1113, N1086, N524);
not NOT1 (N1114, N1113);
xor XOR2 (N1115, N1112, N40);
xor XOR2 (N1116, N1111, N521);
not NOT1 (N1117, N1115);
and AND3 (N1118, N1109, N650, N414);
not NOT1 (N1119, N1118);
nand NAND2 (N1120, N1098, N853);
or OR3 (N1121, N1104, N827, N951);
not NOT1 (N1122, N1114);
or OR4 (N1123, N1119, N372, N658, N338);
or OR2 (N1124, N1122, N800);
buf BUF1 (N1125, N1099);
nand NAND3 (N1126, N1121, N1019, N774);
nand NAND2 (N1127, N1117, N68);
and AND4 (N1128, N1091, N25, N456, N232);
xor XOR2 (N1129, N1124, N98);
or OR2 (N1130, N1128, N925);
xor XOR2 (N1131, N1116, N494);
xor XOR2 (N1132, N1120, N739);
or OR3 (N1133, N1130, N974, N549);
or OR3 (N1134, N1131, N157, N107);
and AND2 (N1135, N1095, N638);
xor XOR2 (N1136, N1132, N267);
nand NAND2 (N1137, N1133, N560);
or OR2 (N1138, N1127, N451);
xor XOR2 (N1139, N1135, N943);
or OR3 (N1140, N1138, N681, N393);
not NOT1 (N1141, N1125);
and AND2 (N1142, N1123, N239);
not NOT1 (N1143, N1142);
nand NAND2 (N1144, N1137, N348);
and AND2 (N1145, N1141, N550);
and AND3 (N1146, N1140, N713, N928);
nand NAND2 (N1147, N1144, N367);
not NOT1 (N1148, N1143);
not NOT1 (N1149, N1126);
and AND2 (N1150, N1108, N200);
nor NOR2 (N1151, N1145, N995);
or OR4 (N1152, N1147, N354, N383, N424);
buf BUF1 (N1153, N1150);
nor NOR4 (N1154, N1134, N803, N365, N664);
not NOT1 (N1155, N1146);
xor XOR2 (N1156, N1136, N777);
xor XOR2 (N1157, N1149, N680);
and AND3 (N1158, N1152, N916, N710);
nand NAND3 (N1159, N1129, N269, N663);
nand NAND4 (N1160, N1148, N386, N970, N680);
nand NAND4 (N1161, N1156, N289, N872, N590);
nor NOR3 (N1162, N1161, N1032, N670);
not NOT1 (N1163, N1139);
buf BUF1 (N1164, N1155);
buf BUF1 (N1165, N1151);
and AND4 (N1166, N1160, N278, N1108, N18);
nor NOR2 (N1167, N1157, N670);
and AND4 (N1168, N1164, N545, N584, N944);
xor XOR2 (N1169, N1167, N586);
and AND2 (N1170, N1158, N948);
xor XOR2 (N1171, N1162, N681);
nor NOR2 (N1172, N1168, N181);
and AND4 (N1173, N1169, N905, N83, N935);
or OR3 (N1174, N1171, N2, N1145);
nand NAND2 (N1175, N1173, N573);
nand NAND3 (N1176, N1172, N203, N267);
and AND3 (N1177, N1175, N693, N42);
and AND4 (N1178, N1153, N616, N10, N16);
xor XOR2 (N1179, N1165, N132);
not NOT1 (N1180, N1170);
nor NOR2 (N1181, N1154, N52);
or OR2 (N1182, N1179, N722);
nor NOR3 (N1183, N1176, N117, N100);
nor NOR3 (N1184, N1183, N424, N637);
not NOT1 (N1185, N1159);
and AND3 (N1186, N1178, N1031, N302);
and AND4 (N1187, N1181, N709, N464, N520);
or OR4 (N1188, N1177, N431, N869, N432);
buf BUF1 (N1189, N1184);
or OR4 (N1190, N1182, N794, N253, N567);
nand NAND4 (N1191, N1180, N1072, N265, N325);
buf BUF1 (N1192, N1174);
and AND2 (N1193, N1185, N1116);
buf BUF1 (N1194, N1191);
nand NAND2 (N1195, N1186, N746);
nand NAND2 (N1196, N1195, N452);
or OR4 (N1197, N1189, N516, N713, N1018);
nand NAND4 (N1198, N1163, N968, N833, N941);
and AND4 (N1199, N1194, N376, N24, N531);
or OR4 (N1200, N1166, N377, N1103, N634);
and AND4 (N1201, N1188, N806, N1050, N382);
or OR2 (N1202, N1192, N485);
or OR2 (N1203, N1190, N31);
nor NOR4 (N1204, N1193, N18, N1203, N248);
not NOT1 (N1205, N774);
and AND3 (N1206, N1204, N578, N522);
and AND3 (N1207, N1198, N654, N762);
buf BUF1 (N1208, N1197);
nor NOR4 (N1209, N1207, N713, N818, N372);
or OR3 (N1210, N1200, N338, N258);
and AND2 (N1211, N1202, N1060);
or OR3 (N1212, N1210, N323, N1066);
nand NAND2 (N1213, N1211, N306);
xor XOR2 (N1214, N1199, N304);
xor XOR2 (N1215, N1206, N220);
xor XOR2 (N1216, N1212, N842);
and AND3 (N1217, N1205, N396, N55);
nor NOR3 (N1218, N1187, N614, N670);
or OR4 (N1219, N1216, N110, N448, N438);
xor XOR2 (N1220, N1201, N1105);
buf BUF1 (N1221, N1220);
nand NAND3 (N1222, N1213, N167, N782);
nand NAND4 (N1223, N1219, N1070, N332, N64);
nor NOR3 (N1224, N1222, N982, N335);
nor NOR2 (N1225, N1224, N739);
nand NAND4 (N1226, N1196, N820, N929, N738);
not NOT1 (N1227, N1209);
nand NAND3 (N1228, N1217, N860, N951);
xor XOR2 (N1229, N1227, N714);
xor XOR2 (N1230, N1214, N303);
or OR4 (N1231, N1223, N705, N583, N298);
xor XOR2 (N1232, N1230, N729);
nor NOR2 (N1233, N1215, N1080);
buf BUF1 (N1234, N1229);
buf BUF1 (N1235, N1231);
buf BUF1 (N1236, N1218);
and AND3 (N1237, N1232, N664, N1175);
nand NAND2 (N1238, N1225, N641);
nor NOR4 (N1239, N1238, N1028, N385, N428);
or OR3 (N1240, N1221, N352, N156);
or OR3 (N1241, N1236, N1032, N589);
not NOT1 (N1242, N1234);
or OR3 (N1243, N1237, N117, N183);
not NOT1 (N1244, N1242);
xor XOR2 (N1245, N1244, N431);
buf BUF1 (N1246, N1240);
not NOT1 (N1247, N1241);
not NOT1 (N1248, N1245);
nand NAND3 (N1249, N1235, N25, N288);
buf BUF1 (N1250, N1228);
not NOT1 (N1251, N1243);
or OR2 (N1252, N1249, N776);
xor XOR2 (N1253, N1247, N1162);
buf BUF1 (N1254, N1250);
not NOT1 (N1255, N1251);
buf BUF1 (N1256, N1239);
or OR3 (N1257, N1233, N734, N864);
buf BUF1 (N1258, N1253);
nand NAND3 (N1259, N1252, N1186, N1240);
and AND3 (N1260, N1246, N180, N1125);
not NOT1 (N1261, N1259);
and AND2 (N1262, N1261, N948);
buf BUF1 (N1263, N1255);
xor XOR2 (N1264, N1258, N573);
and AND4 (N1265, N1256, N618, N401, N186);
not NOT1 (N1266, N1265);
or OR4 (N1267, N1208, N1043, N1214, N21);
nand NAND4 (N1268, N1254, N1266, N733, N835);
nand NAND3 (N1269, N423, N882, N1120);
not NOT1 (N1270, N1268);
not NOT1 (N1271, N1267);
not NOT1 (N1272, N1257);
not NOT1 (N1273, N1271);
and AND3 (N1274, N1273, N836, N683);
not NOT1 (N1275, N1260);
and AND2 (N1276, N1248, N421);
not NOT1 (N1277, N1272);
xor XOR2 (N1278, N1263, N199);
and AND2 (N1279, N1262, N1112);
and AND2 (N1280, N1279, N255);
or OR2 (N1281, N1264, N192);
not NOT1 (N1282, N1270);
and AND4 (N1283, N1276, N810, N1086, N851);
nand NAND2 (N1284, N1226, N1122);
not NOT1 (N1285, N1284);
and AND2 (N1286, N1277, N441);
nand NAND2 (N1287, N1282, N465);
or OR4 (N1288, N1275, N158, N159, N885);
xor XOR2 (N1289, N1285, N878);
or OR2 (N1290, N1283, N896);
or OR4 (N1291, N1274, N1200, N564, N135);
nand NAND2 (N1292, N1288, N858);
nand NAND2 (N1293, N1269, N1276);
nand NAND3 (N1294, N1292, N1114, N288);
nand NAND3 (N1295, N1278, N1128, N460);
buf BUF1 (N1296, N1291);
or OR2 (N1297, N1293, N735);
nand NAND3 (N1298, N1294, N998, N518);
nor NOR2 (N1299, N1297, N743);
xor XOR2 (N1300, N1280, N26);
or OR4 (N1301, N1295, N345, N705, N364);
buf BUF1 (N1302, N1300);
nand NAND2 (N1303, N1301, N119);
buf BUF1 (N1304, N1302);
not NOT1 (N1305, N1299);
not NOT1 (N1306, N1289);
and AND2 (N1307, N1281, N1187);
buf BUF1 (N1308, N1296);
buf BUF1 (N1309, N1287);
nand NAND3 (N1310, N1298, N1285, N413);
xor XOR2 (N1311, N1310, N1094);
nand NAND3 (N1312, N1308, N330, N1134);
xor XOR2 (N1313, N1312, N1008);
buf BUF1 (N1314, N1290);
xor XOR2 (N1315, N1306, N1073);
xor XOR2 (N1316, N1313, N157);
and AND4 (N1317, N1304, N590, N636, N1203);
nand NAND2 (N1318, N1303, N1192);
nor NOR4 (N1319, N1315, N620, N91, N1159);
nand NAND2 (N1320, N1316, N889);
or OR4 (N1321, N1314, N964, N190, N855);
nand NAND3 (N1322, N1318, N416, N58);
not NOT1 (N1323, N1305);
not NOT1 (N1324, N1307);
nand NAND3 (N1325, N1320, N903, N327);
nand NAND4 (N1326, N1321, N1178, N1248, N688);
nand NAND3 (N1327, N1311, N381, N114);
xor XOR2 (N1328, N1286, N426);
nand NAND2 (N1329, N1328, N1289);
not NOT1 (N1330, N1322);
xor XOR2 (N1331, N1329, N360);
not NOT1 (N1332, N1326);
or OR4 (N1333, N1309, N224, N241, N885);
xor XOR2 (N1334, N1319, N210);
xor XOR2 (N1335, N1327, N28);
and AND4 (N1336, N1317, N1194, N1134, N697);
nand NAND3 (N1337, N1323, N999, N1058);
not NOT1 (N1338, N1335);
nand NAND3 (N1339, N1331, N1195, N1324);
or OR4 (N1340, N458, N136, N571, N1122);
or OR4 (N1341, N1330, N563, N574, N905);
nor NOR4 (N1342, N1325, N1302, N983, N733);
or OR4 (N1343, N1333, N799, N359, N947);
not NOT1 (N1344, N1343);
not NOT1 (N1345, N1334);
and AND4 (N1346, N1339, N971, N18, N70);
buf BUF1 (N1347, N1332);
or OR2 (N1348, N1347, N199);
xor XOR2 (N1349, N1348, N161);
nor NOR4 (N1350, N1340, N1168, N25, N1348);
nand NAND3 (N1351, N1338, N14, N718);
buf BUF1 (N1352, N1346);
nor NOR4 (N1353, N1337, N763, N527, N1290);
or OR3 (N1354, N1341, N532, N422);
not NOT1 (N1355, N1353);
or OR4 (N1356, N1344, N495, N188, N423);
buf BUF1 (N1357, N1351);
not NOT1 (N1358, N1336);
nand NAND3 (N1359, N1350, N491, N167);
nor NOR3 (N1360, N1342, N1179, N1058);
xor XOR2 (N1361, N1357, N438);
nor NOR4 (N1362, N1360, N1320, N377, N744);
buf BUF1 (N1363, N1345);
nor NOR2 (N1364, N1354, N685);
not NOT1 (N1365, N1359);
xor XOR2 (N1366, N1365, N425);
nand NAND4 (N1367, N1352, N728, N1126, N1154);
nor NOR4 (N1368, N1363, N418, N502, N1216);
xor XOR2 (N1369, N1358, N909);
buf BUF1 (N1370, N1364);
and AND2 (N1371, N1355, N1321);
not NOT1 (N1372, N1361);
or OR2 (N1373, N1367, N710);
or OR4 (N1374, N1349, N801, N141, N1158);
nor NOR4 (N1375, N1371, N713, N74, N168);
not NOT1 (N1376, N1373);
not NOT1 (N1377, N1376);
buf BUF1 (N1378, N1372);
xor XOR2 (N1379, N1370, N938);
nor NOR2 (N1380, N1379, N276);
buf BUF1 (N1381, N1356);
xor XOR2 (N1382, N1380, N585);
nand NAND3 (N1383, N1369, N937, N161);
buf BUF1 (N1384, N1374);
nor NOR2 (N1385, N1368, N596);
nor NOR4 (N1386, N1362, N615, N191, N347);
nand NAND2 (N1387, N1378, N856);
xor XOR2 (N1388, N1377, N641);
buf BUF1 (N1389, N1383);
nand NAND2 (N1390, N1389, N536);
nand NAND4 (N1391, N1388, N665, N392, N1365);
not NOT1 (N1392, N1366);
buf BUF1 (N1393, N1381);
buf BUF1 (N1394, N1386);
and AND3 (N1395, N1384, N586, N333);
nand NAND4 (N1396, N1390, N717, N966, N495);
buf BUF1 (N1397, N1392);
buf BUF1 (N1398, N1375);
or OR3 (N1399, N1387, N487, N1133);
xor XOR2 (N1400, N1399, N227);
nor NOR4 (N1401, N1400, N10, N683, N259);
nor NOR3 (N1402, N1382, N1210, N322);
and AND3 (N1403, N1398, N775, N706);
nor NOR3 (N1404, N1401, N662, N153);
or OR3 (N1405, N1404, N1111, N699);
nand NAND3 (N1406, N1402, N578, N1337);
buf BUF1 (N1407, N1405);
nand NAND4 (N1408, N1397, N114, N806, N875);
xor XOR2 (N1409, N1408, N1313);
buf BUF1 (N1410, N1396);
nor NOR4 (N1411, N1391, N450, N1200, N754);
nand NAND2 (N1412, N1393, N1339);
and AND2 (N1413, N1409, N91);
or OR3 (N1414, N1407, N1142, N473);
or OR4 (N1415, N1394, N1122, N426, N874);
nand NAND3 (N1416, N1395, N454, N1113);
and AND3 (N1417, N1411, N715, N1118);
and AND2 (N1418, N1413, N409);
nor NOR4 (N1419, N1403, N189, N871, N1089);
xor XOR2 (N1420, N1410, N865);
or OR4 (N1421, N1419, N1319, N1341, N556);
nor NOR3 (N1422, N1417, N774, N631);
nor NOR4 (N1423, N1414, N700, N1368, N1026);
xor XOR2 (N1424, N1406, N927);
nor NOR2 (N1425, N1423, N511);
nor NOR2 (N1426, N1421, N1250);
nor NOR4 (N1427, N1426, N1325, N269, N346);
or OR4 (N1428, N1416, N1323, N1209, N817);
buf BUF1 (N1429, N1424);
buf BUF1 (N1430, N1385);
nand NAND3 (N1431, N1430, N896, N1320);
nor NOR3 (N1432, N1428, N135, N283);
buf BUF1 (N1433, N1425);
buf BUF1 (N1434, N1412);
not NOT1 (N1435, N1431);
nor NOR4 (N1436, N1422, N360, N430, N456);
not NOT1 (N1437, N1429);
nor NOR3 (N1438, N1436, N1119, N188);
nor NOR3 (N1439, N1438, N140, N1284);
nor NOR4 (N1440, N1437, N792, N946, N1356);
and AND4 (N1441, N1415, N233, N145, N508);
nand NAND2 (N1442, N1420, N379);
buf BUF1 (N1443, N1435);
nand NAND2 (N1444, N1443, N1348);
not NOT1 (N1445, N1434);
nand NAND3 (N1446, N1441, N930, N31);
or OR2 (N1447, N1432, N930);
xor XOR2 (N1448, N1440, N1343);
nor NOR2 (N1449, N1418, N950);
not NOT1 (N1450, N1433);
buf BUF1 (N1451, N1447);
and AND2 (N1452, N1445, N724);
nor NOR3 (N1453, N1449, N1007, N523);
xor XOR2 (N1454, N1427, N488);
nand NAND3 (N1455, N1448, N141, N1407);
or OR4 (N1456, N1455, N14, N841, N1411);
and AND4 (N1457, N1439, N227, N826, N21);
xor XOR2 (N1458, N1454, N216);
and AND3 (N1459, N1452, N469, N1321);
buf BUF1 (N1460, N1442);
and AND3 (N1461, N1459, N176, N329);
and AND4 (N1462, N1456, N692, N2, N745);
and AND3 (N1463, N1451, N80, N867);
nor NOR3 (N1464, N1460, N330, N767);
buf BUF1 (N1465, N1462);
not NOT1 (N1466, N1450);
and AND2 (N1467, N1446, N266);
nor NOR2 (N1468, N1461, N832);
or OR4 (N1469, N1465, N1361, N618, N25);
nand NAND3 (N1470, N1444, N1276, N1008);
not NOT1 (N1471, N1457);
and AND3 (N1472, N1468, N255, N1087);
xor XOR2 (N1473, N1453, N932);
not NOT1 (N1474, N1470);
buf BUF1 (N1475, N1474);
buf BUF1 (N1476, N1458);
nor NOR4 (N1477, N1476, N1255, N1032, N1303);
and AND3 (N1478, N1464, N1044, N450);
xor XOR2 (N1479, N1471, N1304);
nor NOR2 (N1480, N1469, N810);
nand NAND3 (N1481, N1479, N941, N1056);
not NOT1 (N1482, N1467);
not NOT1 (N1483, N1480);
nor NOR4 (N1484, N1481, N597, N943, N1203);
and AND4 (N1485, N1478, N1366, N756, N793);
xor XOR2 (N1486, N1482, N1369);
nand NAND2 (N1487, N1463, N94);
or OR2 (N1488, N1487, N831);
xor XOR2 (N1489, N1484, N828);
or OR2 (N1490, N1488, N1272);
nor NOR2 (N1491, N1472, N588);
not NOT1 (N1492, N1466);
nor NOR3 (N1493, N1475, N581, N1187);
nand NAND2 (N1494, N1490, N1158);
not NOT1 (N1495, N1489);
not NOT1 (N1496, N1486);
xor XOR2 (N1497, N1494, N155);
buf BUF1 (N1498, N1483);
and AND2 (N1499, N1498, N1311);
nor NOR3 (N1500, N1491, N460, N638);
nor NOR4 (N1501, N1485, N1155, N1105, N1247);
nand NAND4 (N1502, N1496, N1377, N552, N1418);
or OR4 (N1503, N1502, N476, N685, N324);
nand NAND3 (N1504, N1503, N332, N391);
buf BUF1 (N1505, N1497);
and AND3 (N1506, N1505, N820, N155);
nand NAND2 (N1507, N1473, N345);
not NOT1 (N1508, N1507);
xor XOR2 (N1509, N1493, N372);
or OR4 (N1510, N1501, N1119, N1070, N1172);
buf BUF1 (N1511, N1506);
and AND2 (N1512, N1500, N555);
nor NOR4 (N1513, N1510, N140, N1377, N891);
not NOT1 (N1514, N1513);
or OR3 (N1515, N1511, N907, N822);
buf BUF1 (N1516, N1515);
not NOT1 (N1517, N1495);
xor XOR2 (N1518, N1517, N121);
and AND2 (N1519, N1516, N997);
nand NAND4 (N1520, N1504, N727, N1341, N927);
buf BUF1 (N1521, N1519);
and AND3 (N1522, N1508, N779, N1281);
nand NAND2 (N1523, N1520, N676);
xor XOR2 (N1524, N1492, N583);
nor NOR2 (N1525, N1518, N933);
nand NAND4 (N1526, N1514, N848, N879, N917);
buf BUF1 (N1527, N1477);
and AND3 (N1528, N1512, N832, N528);
nor NOR2 (N1529, N1521, N1065);
buf BUF1 (N1530, N1525);
nor NOR4 (N1531, N1499, N143, N210, N101);
buf BUF1 (N1532, N1526);
and AND3 (N1533, N1522, N976, N941);
xor XOR2 (N1534, N1509, N689);
not NOT1 (N1535, N1530);
nand NAND4 (N1536, N1532, N782, N1249, N756);
not NOT1 (N1537, N1535);
and AND4 (N1538, N1537, N619, N1506, N983);
nand NAND3 (N1539, N1524, N887, N1476);
and AND2 (N1540, N1533, N1407);
nand NAND4 (N1541, N1527, N1498, N1459, N1299);
nor NOR2 (N1542, N1540, N1305);
xor XOR2 (N1543, N1528, N1530);
buf BUF1 (N1544, N1534);
nand NAND2 (N1545, N1541, N1244);
buf BUF1 (N1546, N1538);
nor NOR3 (N1547, N1523, N1488, N1112);
not NOT1 (N1548, N1542);
nor NOR3 (N1549, N1547, N1226, N1292);
xor XOR2 (N1550, N1546, N881);
nor NOR2 (N1551, N1539, N1254);
or OR4 (N1552, N1548, N1035, N1527, N775);
nor NOR4 (N1553, N1549, N1201, N624, N1320);
nor NOR3 (N1554, N1552, N1477, N993);
nand NAND2 (N1555, N1543, N567);
nand NAND2 (N1556, N1531, N164);
nor NOR2 (N1557, N1554, N969);
and AND4 (N1558, N1553, N362, N580, N1494);
not NOT1 (N1559, N1544);
nor NOR2 (N1560, N1529, N1166);
and AND2 (N1561, N1555, N921);
and AND2 (N1562, N1560, N1121);
nor NOR3 (N1563, N1557, N849, N466);
or OR2 (N1564, N1558, N78);
buf BUF1 (N1565, N1550);
not NOT1 (N1566, N1545);
not NOT1 (N1567, N1559);
xor XOR2 (N1568, N1561, N150);
not NOT1 (N1569, N1563);
and AND4 (N1570, N1568, N1288, N16, N749);
nand NAND2 (N1571, N1569, N48);
nand NAND3 (N1572, N1556, N386, N109);
not NOT1 (N1573, N1572);
xor XOR2 (N1574, N1565, N1402);
not NOT1 (N1575, N1562);
not NOT1 (N1576, N1567);
and AND2 (N1577, N1566, N514);
and AND4 (N1578, N1577, N206, N290, N1288);
buf BUF1 (N1579, N1570);
nand NAND2 (N1580, N1551, N473);
nand NAND2 (N1581, N1575, N1561);
or OR2 (N1582, N1581, N526);
nor NOR3 (N1583, N1582, N543, N272);
not NOT1 (N1584, N1571);
or OR3 (N1585, N1536, N569, N74);
not NOT1 (N1586, N1574);
nand NAND2 (N1587, N1585, N575);
xor XOR2 (N1588, N1576, N831);
and AND3 (N1589, N1578, N412, N1579);
nor NOR3 (N1590, N123, N1345, N971);
nor NOR2 (N1591, N1580, N1535);
not NOT1 (N1592, N1586);
xor XOR2 (N1593, N1592, N669);
nor NOR4 (N1594, N1591, N1491, N1479, N294);
nand NAND3 (N1595, N1593, N501, N399);
nor NOR3 (N1596, N1573, N706, N1270);
buf BUF1 (N1597, N1596);
xor XOR2 (N1598, N1584, N1121);
nand NAND4 (N1599, N1594, N1397, N935, N1137);
buf BUF1 (N1600, N1599);
or OR3 (N1601, N1583, N431, N1296);
nand NAND3 (N1602, N1600, N688, N1369);
and AND4 (N1603, N1595, N335, N888, N646);
buf BUF1 (N1604, N1598);
nor NOR4 (N1605, N1597, N1384, N560, N1374);
nand NAND2 (N1606, N1603, N1319);
and AND4 (N1607, N1604, N228, N831, N494);
not NOT1 (N1608, N1590);
and AND4 (N1609, N1608, N1444, N1210, N618);
xor XOR2 (N1610, N1601, N1562);
and AND4 (N1611, N1564, N1150, N1205, N951);
buf BUF1 (N1612, N1611);
or OR4 (N1613, N1602, N1523, N27, N1117);
nand NAND4 (N1614, N1587, N1001, N506, N1220);
and AND3 (N1615, N1589, N221, N469);
nand NAND3 (N1616, N1605, N1487, N563);
buf BUF1 (N1617, N1606);
nor NOR4 (N1618, N1616, N420, N239, N380);
or OR2 (N1619, N1612, N207);
nand NAND2 (N1620, N1618, N896);
not NOT1 (N1621, N1619);
and AND2 (N1622, N1607, N500);
or OR4 (N1623, N1622, N502, N1507, N1172);
nor NOR2 (N1624, N1588, N1237);
not NOT1 (N1625, N1613);
not NOT1 (N1626, N1625);
and AND4 (N1627, N1615, N83, N1420, N109);
nor NOR4 (N1628, N1627, N490, N1295, N1125);
and AND3 (N1629, N1610, N994, N592);
buf BUF1 (N1630, N1626);
xor XOR2 (N1631, N1623, N871);
or OR4 (N1632, N1630, N443, N745, N205);
not NOT1 (N1633, N1621);
and AND2 (N1634, N1629, N1103);
buf BUF1 (N1635, N1609);
and AND2 (N1636, N1628, N970);
buf BUF1 (N1637, N1620);
or OR2 (N1638, N1631, N443);
or OR3 (N1639, N1617, N317, N251);
and AND2 (N1640, N1624, N1608);
buf BUF1 (N1641, N1639);
nor NOR4 (N1642, N1632, N1594, N719, N1448);
not NOT1 (N1643, N1635);
buf BUF1 (N1644, N1642);
not NOT1 (N1645, N1637);
nor NOR3 (N1646, N1645, N792, N570);
buf BUF1 (N1647, N1633);
buf BUF1 (N1648, N1636);
or OR3 (N1649, N1641, N8, N623);
and AND3 (N1650, N1614, N1310, N677);
and AND2 (N1651, N1643, N354);
not NOT1 (N1652, N1638);
and AND2 (N1653, N1650, N41);
xor XOR2 (N1654, N1647, N1489);
buf BUF1 (N1655, N1646);
nor NOR2 (N1656, N1652, N1245);
buf BUF1 (N1657, N1654);
or OR4 (N1658, N1648, N1026, N917, N1625);
or OR4 (N1659, N1649, N1185, N299, N160);
nand NAND2 (N1660, N1651, N38);
nand NAND4 (N1661, N1640, N297, N1546, N261);
not NOT1 (N1662, N1656);
not NOT1 (N1663, N1655);
or OR2 (N1664, N1658, N960);
buf BUF1 (N1665, N1661);
nor NOR4 (N1666, N1657, N720, N1519, N1425);
nand NAND2 (N1667, N1665, N1174);
and AND2 (N1668, N1666, N66);
and AND4 (N1669, N1634, N722, N382, N1281);
xor XOR2 (N1670, N1644, N1390);
xor XOR2 (N1671, N1670, N797);
not NOT1 (N1672, N1663);
not NOT1 (N1673, N1671);
and AND2 (N1674, N1667, N1301);
nand NAND2 (N1675, N1673, N700);
and AND2 (N1676, N1659, N1277);
xor XOR2 (N1677, N1662, N1171);
not NOT1 (N1678, N1676);
not NOT1 (N1679, N1664);
or OR4 (N1680, N1660, N1594, N926, N463);
or OR2 (N1681, N1678, N744);
xor XOR2 (N1682, N1679, N37);
nor NOR4 (N1683, N1682, N973, N1644, N10);
not NOT1 (N1684, N1675);
buf BUF1 (N1685, N1668);
not NOT1 (N1686, N1683);
nor NOR3 (N1687, N1672, N698, N1621);
buf BUF1 (N1688, N1681);
and AND2 (N1689, N1688, N1434);
not NOT1 (N1690, N1669);
nand NAND2 (N1691, N1677, N1469);
and AND3 (N1692, N1674, N863, N848);
and AND3 (N1693, N1687, N34, N1018);
nor NOR2 (N1694, N1690, N222);
buf BUF1 (N1695, N1692);
and AND3 (N1696, N1653, N1206, N625);
xor XOR2 (N1697, N1689, N708);
and AND3 (N1698, N1680, N289, N66);
and AND2 (N1699, N1695, N220);
nor NOR2 (N1700, N1694, N970);
nor NOR4 (N1701, N1685, N639, N67, N1361);
xor XOR2 (N1702, N1701, N644);
not NOT1 (N1703, N1697);
not NOT1 (N1704, N1684);
not NOT1 (N1705, N1691);
xor XOR2 (N1706, N1686, N1616);
buf BUF1 (N1707, N1699);
nand NAND2 (N1708, N1703, N986);
nand NAND3 (N1709, N1698, N1165, N1527);
and AND3 (N1710, N1704, N545, N1633);
and AND3 (N1711, N1709, N1635, N163);
and AND3 (N1712, N1707, N1425, N1543);
buf BUF1 (N1713, N1693);
and AND4 (N1714, N1712, N370, N298, N818);
buf BUF1 (N1715, N1696);
or OR4 (N1716, N1706, N784, N1407, N1192);
or OR3 (N1717, N1715, N174, N1469);
nor NOR2 (N1718, N1710, N314);
xor XOR2 (N1719, N1705, N626);
or OR3 (N1720, N1708, N431, N823);
not NOT1 (N1721, N1702);
nand NAND2 (N1722, N1718, N1213);
not NOT1 (N1723, N1711);
or OR2 (N1724, N1722, N624);
buf BUF1 (N1725, N1717);
buf BUF1 (N1726, N1714);
xor XOR2 (N1727, N1719, N1035);
or OR2 (N1728, N1716, N301);
buf BUF1 (N1729, N1723);
or OR4 (N1730, N1700, N1260, N1289, N627);
buf BUF1 (N1731, N1730);
not NOT1 (N1732, N1713);
buf BUF1 (N1733, N1724);
nand NAND3 (N1734, N1720, N201, N1309);
not NOT1 (N1735, N1725);
or OR3 (N1736, N1734, N38, N845);
nor NOR3 (N1737, N1721, N1567, N992);
or OR3 (N1738, N1736, N1585, N469);
nand NAND4 (N1739, N1728, N357, N1451, N1721);
or OR2 (N1740, N1726, N921);
nand NAND4 (N1741, N1729, N1417, N1387, N239);
xor XOR2 (N1742, N1737, N56);
not NOT1 (N1743, N1735);
nand NAND3 (N1744, N1743, N1480, N1615);
or OR2 (N1745, N1744, N1206);
xor XOR2 (N1746, N1732, N1209);
or OR4 (N1747, N1746, N294, N1308, N717);
nor NOR3 (N1748, N1741, N214, N1045);
nor NOR2 (N1749, N1747, N808);
or OR2 (N1750, N1745, N347);
and AND2 (N1751, N1733, N553);
buf BUF1 (N1752, N1731);
nand NAND3 (N1753, N1739, N976, N1730);
nand NAND4 (N1754, N1742, N1316, N820, N1065);
nor NOR4 (N1755, N1754, N874, N1255, N774);
buf BUF1 (N1756, N1750);
and AND3 (N1757, N1755, N328, N509);
not NOT1 (N1758, N1740);
or OR2 (N1759, N1752, N1232);
nand NAND2 (N1760, N1751, N427);
and AND2 (N1761, N1759, N148);
xor XOR2 (N1762, N1757, N211);
buf BUF1 (N1763, N1727);
xor XOR2 (N1764, N1760, N992);
xor XOR2 (N1765, N1764, N1200);
nand NAND4 (N1766, N1758, N1745, N977, N239);
xor XOR2 (N1767, N1765, N774);
or OR2 (N1768, N1753, N1526);
or OR2 (N1769, N1748, N1303);
nand NAND2 (N1770, N1761, N108);
buf BUF1 (N1771, N1766);
buf BUF1 (N1772, N1756);
nand NAND3 (N1773, N1771, N1066, N1535);
buf BUF1 (N1774, N1762);
and AND4 (N1775, N1774, N1060, N606, N614);
nand NAND2 (N1776, N1738, N903);
and AND4 (N1777, N1763, N1580, N1237, N43);
buf BUF1 (N1778, N1749);
buf BUF1 (N1779, N1768);
and AND3 (N1780, N1776, N420, N329);
xor XOR2 (N1781, N1772, N1482);
buf BUF1 (N1782, N1781);
xor XOR2 (N1783, N1770, N1425);
and AND2 (N1784, N1769, N474);
xor XOR2 (N1785, N1778, N857);
nor NOR3 (N1786, N1785, N261, N472);
not NOT1 (N1787, N1780);
and AND4 (N1788, N1783, N1380, N606, N466);
or OR4 (N1789, N1786, N707, N274, N339);
or OR2 (N1790, N1779, N817);
buf BUF1 (N1791, N1789);
or OR4 (N1792, N1773, N1147, N1257, N1571);
buf BUF1 (N1793, N1791);
or OR3 (N1794, N1782, N1660, N271);
xor XOR2 (N1795, N1793, N1490);
buf BUF1 (N1796, N1787);
xor XOR2 (N1797, N1796, N757);
xor XOR2 (N1798, N1788, N1238);
buf BUF1 (N1799, N1784);
buf BUF1 (N1800, N1797);
buf BUF1 (N1801, N1798);
or OR2 (N1802, N1795, N1154);
and AND4 (N1803, N1802, N1700, N1777, N430);
nand NAND3 (N1804, N1161, N1099, N844);
nor NOR4 (N1805, N1794, N1001, N1367, N1412);
xor XOR2 (N1806, N1801, N436);
nor NOR3 (N1807, N1775, N7, N344);
xor XOR2 (N1808, N1803, N1673);
nor NOR3 (N1809, N1807, N1126, N952);
nand NAND2 (N1810, N1808, N1806);
buf BUF1 (N1811, N713);
not NOT1 (N1812, N1811);
and AND2 (N1813, N1790, N96);
xor XOR2 (N1814, N1792, N1803);
buf BUF1 (N1815, N1809);
buf BUF1 (N1816, N1810);
nand NAND3 (N1817, N1815, N255, N229);
xor XOR2 (N1818, N1813, N553);
and AND4 (N1819, N1816, N1627, N1586, N638);
not NOT1 (N1820, N1819);
or OR4 (N1821, N1767, N48, N506, N544);
nand NAND4 (N1822, N1820, N1398, N331, N1174);
xor XOR2 (N1823, N1822, N1370);
not NOT1 (N1824, N1799);
nand NAND2 (N1825, N1812, N1495);
xor XOR2 (N1826, N1818, N226);
nand NAND4 (N1827, N1804, N1722, N1666, N872);
buf BUF1 (N1828, N1821);
nor NOR4 (N1829, N1826, N539, N379, N1800);
nor NOR2 (N1830, N1427, N714);
nor NOR4 (N1831, N1827, N825, N46, N467);
and AND2 (N1832, N1814, N751);
or OR3 (N1833, N1829, N1534, N38);
xor XOR2 (N1834, N1833, N1092);
buf BUF1 (N1835, N1828);
buf BUF1 (N1836, N1830);
xor XOR2 (N1837, N1831, N93);
or OR4 (N1838, N1835, N1513, N397, N572);
nor NOR2 (N1839, N1838, N25);
nor NOR3 (N1840, N1837, N424, N725);
nor NOR2 (N1841, N1824, N1040);
and AND3 (N1842, N1805, N1265, N1035);
xor XOR2 (N1843, N1825, N5);
not NOT1 (N1844, N1817);
buf BUF1 (N1845, N1841);
xor XOR2 (N1846, N1844, N1507);
and AND3 (N1847, N1832, N802, N46);
xor XOR2 (N1848, N1839, N1767);
xor XOR2 (N1849, N1845, N1495);
xor XOR2 (N1850, N1842, N1280);
nor NOR2 (N1851, N1823, N60);
nor NOR4 (N1852, N1851, N675, N141, N583);
xor XOR2 (N1853, N1836, N1722);
buf BUF1 (N1854, N1846);
and AND2 (N1855, N1848, N1131);
or OR4 (N1856, N1849, N375, N1682, N838);
not NOT1 (N1857, N1850);
xor XOR2 (N1858, N1847, N131);
and AND4 (N1859, N1857, N694, N1804, N1188);
nand NAND2 (N1860, N1856, N327);
or OR4 (N1861, N1858, N535, N426, N470);
xor XOR2 (N1862, N1853, N1635);
and AND3 (N1863, N1859, N1123, N977);
nor NOR4 (N1864, N1861, N18, N1119, N1695);
or OR3 (N1865, N1840, N531, N152);
not NOT1 (N1866, N1865);
not NOT1 (N1867, N1843);
nor NOR3 (N1868, N1866, N1812, N920);
xor XOR2 (N1869, N1863, N1153);
nand NAND2 (N1870, N1862, N592);
buf BUF1 (N1871, N1864);
and AND4 (N1872, N1868, N1063, N1424, N1447);
nor NOR4 (N1873, N1834, N1575, N913, N1069);
or OR3 (N1874, N1872, N825, N1796);
xor XOR2 (N1875, N1855, N304);
xor XOR2 (N1876, N1874, N1574);
not NOT1 (N1877, N1875);
xor XOR2 (N1878, N1852, N1539);
and AND4 (N1879, N1869, N458, N772, N490);
and AND3 (N1880, N1878, N1756, N1752);
nor NOR2 (N1881, N1860, N1162);
nand NAND2 (N1882, N1876, N71);
nand NAND3 (N1883, N1877, N494, N603);
nor NOR4 (N1884, N1881, N1442, N152, N168);
xor XOR2 (N1885, N1871, N637);
not NOT1 (N1886, N1883);
or OR2 (N1887, N1885, N571);
xor XOR2 (N1888, N1867, N1441);
or OR2 (N1889, N1882, N321);
and AND2 (N1890, N1870, N346);
nor NOR2 (N1891, N1884, N654);
not NOT1 (N1892, N1889);
and AND2 (N1893, N1880, N246);
and AND3 (N1894, N1873, N631, N1570);
nor NOR4 (N1895, N1890, N1449, N616, N1754);
or OR3 (N1896, N1892, N770, N106);
nand NAND4 (N1897, N1887, N218, N706, N1080);
xor XOR2 (N1898, N1886, N739);
xor XOR2 (N1899, N1896, N1673);
nand NAND4 (N1900, N1897, N942, N175, N1318);
nor NOR4 (N1901, N1898, N638, N1645, N1530);
or OR2 (N1902, N1894, N1742);
nor NOR2 (N1903, N1902, N743);
and AND4 (N1904, N1899, N1041, N654, N1773);
nor NOR2 (N1905, N1891, N1537);
nand NAND4 (N1906, N1854, N1101, N1600, N1833);
buf BUF1 (N1907, N1893);
nor NOR3 (N1908, N1903, N1540, N575);
xor XOR2 (N1909, N1901, N814);
and AND2 (N1910, N1895, N1463);
or OR4 (N1911, N1904, N273, N1332, N1622);
nand NAND2 (N1912, N1910, N1062);
nor NOR4 (N1913, N1911, N65, N1483, N885);
or OR4 (N1914, N1907, N60, N1430, N1443);
nand NAND3 (N1915, N1909, N1002, N1816);
not NOT1 (N1916, N1908);
nor NOR2 (N1917, N1915, N1349);
xor XOR2 (N1918, N1906, N362);
xor XOR2 (N1919, N1888, N372);
and AND2 (N1920, N1913, N1078);
nor NOR2 (N1921, N1914, N826);
nand NAND3 (N1922, N1920, N1441, N649);
not NOT1 (N1923, N1918);
nand NAND3 (N1924, N1905, N920, N220);
not NOT1 (N1925, N1916);
buf BUF1 (N1926, N1900);
buf BUF1 (N1927, N1922);
nor NOR2 (N1928, N1923, N1791);
nor NOR2 (N1929, N1912, N1349);
xor XOR2 (N1930, N1926, N1019);
xor XOR2 (N1931, N1917, N720);
or OR3 (N1932, N1924, N323, N215);
buf BUF1 (N1933, N1932);
and AND3 (N1934, N1919, N968, N1148);
not NOT1 (N1935, N1931);
xor XOR2 (N1936, N1929, N917);
nor NOR2 (N1937, N1879, N229);
xor XOR2 (N1938, N1933, N658);
not NOT1 (N1939, N1935);
not NOT1 (N1940, N1921);
nand NAND4 (N1941, N1927, N1267, N211, N1797);
not NOT1 (N1942, N1934);
not NOT1 (N1943, N1936);
xor XOR2 (N1944, N1941, N475);
nand NAND3 (N1945, N1937, N766, N163);
and AND2 (N1946, N1925, N497);
buf BUF1 (N1947, N1944);
and AND3 (N1948, N1947, N1297, N103);
and AND3 (N1949, N1938, N1123, N1159);
nor NOR3 (N1950, N1942, N746, N603);
not NOT1 (N1951, N1939);
nand NAND4 (N1952, N1951, N845, N1944, N1486);
xor XOR2 (N1953, N1940, N1017);
nor NOR2 (N1954, N1950, N1803);
xor XOR2 (N1955, N1946, N256);
xor XOR2 (N1956, N1948, N1902);
xor XOR2 (N1957, N1955, N1791);
not NOT1 (N1958, N1945);
not NOT1 (N1959, N1958);
xor XOR2 (N1960, N1957, N232);
xor XOR2 (N1961, N1956, N1100);
and AND4 (N1962, N1953, N869, N1137, N298);
nand NAND4 (N1963, N1930, N1934, N155, N963);
xor XOR2 (N1964, N1959, N472);
nor NOR3 (N1965, N1963, N1407, N112);
not NOT1 (N1966, N1952);
or OR4 (N1967, N1960, N1320, N1916, N973);
or OR2 (N1968, N1961, N30);
buf BUF1 (N1969, N1954);
and AND2 (N1970, N1962, N1812);
xor XOR2 (N1971, N1967, N1678);
or OR2 (N1972, N1969, N1183);
nor NOR4 (N1973, N1970, N1970, N602, N1658);
xor XOR2 (N1974, N1965, N1054);
nor NOR3 (N1975, N1949, N522, N94);
buf BUF1 (N1976, N1968);
xor XOR2 (N1977, N1972, N104);
xor XOR2 (N1978, N1977, N1577);
and AND4 (N1979, N1966, N1156, N1538, N1509);
nor NOR2 (N1980, N1976, N1264);
nand NAND2 (N1981, N1979, N1831);
nor NOR3 (N1982, N1981, N573, N818);
xor XOR2 (N1983, N1964, N323);
xor XOR2 (N1984, N1974, N1524);
nor NOR4 (N1985, N1978, N1662, N898, N552);
or OR3 (N1986, N1985, N282, N260);
and AND4 (N1987, N1928, N377, N433, N1610);
and AND3 (N1988, N1986, N619, N1914);
and AND3 (N1989, N1980, N945, N284);
buf BUF1 (N1990, N1987);
xor XOR2 (N1991, N1971, N110);
xor XOR2 (N1992, N1988, N1781);
buf BUF1 (N1993, N1990);
and AND2 (N1994, N1991, N1907);
buf BUF1 (N1995, N1989);
nor NOR2 (N1996, N1994, N474);
nand NAND3 (N1997, N1984, N641, N457);
xor XOR2 (N1998, N1943, N870);
nor NOR3 (N1999, N1992, N1970, N246);
nor NOR3 (N2000, N1999, N1497, N1405);
buf BUF1 (N2001, N1996);
nor NOR2 (N2002, N2001, N134);
nor NOR4 (N2003, N2000, N1661, N796, N1305);
nor NOR4 (N2004, N1973, N1804, N309, N928);
not NOT1 (N2005, N1993);
nand NAND3 (N2006, N1997, N176, N1867);
and AND2 (N2007, N2002, N557);
or OR2 (N2008, N1998, N88);
buf BUF1 (N2009, N2004);
or OR2 (N2010, N2008, N307);
nand NAND3 (N2011, N1982, N1110, N1779);
xor XOR2 (N2012, N2007, N1771);
xor XOR2 (N2013, N2006, N1418);
or OR4 (N2014, N2005, N458, N1120, N1775);
and AND2 (N2015, N2013, N897);
and AND3 (N2016, N2003, N1831, N622);
nor NOR3 (N2017, N2010, N1469, N1252);
nor NOR3 (N2018, N2017, N281, N728);
or OR3 (N2019, N1983, N1423, N1020);
or OR3 (N2020, N2012, N1696, N659);
xor XOR2 (N2021, N2009, N1681);
nand NAND2 (N2022, N1975, N1023);
xor XOR2 (N2023, N2014, N1143);
nor NOR4 (N2024, N2019, N590, N624, N1284);
nand NAND2 (N2025, N2015, N218);
and AND4 (N2026, N2020, N128, N283, N72);
and AND4 (N2027, N2016, N564, N128, N1390);
not NOT1 (N2028, N2021);
and AND3 (N2029, N1995, N927, N189);
not NOT1 (N2030, N2011);
not NOT1 (N2031, N2029);
nand NAND2 (N2032, N2022, N779);
buf BUF1 (N2033, N2032);
xor XOR2 (N2034, N2026, N919);
nand NAND4 (N2035, N2023, N1784, N1014, N756);
xor XOR2 (N2036, N2024, N1026);
buf BUF1 (N2037, N2033);
xor XOR2 (N2038, N2025, N492);
or OR3 (N2039, N2030, N368, N1950);
buf BUF1 (N2040, N2037);
or OR4 (N2041, N2039, N691, N2016, N1694);
buf BUF1 (N2042, N2034);
nor NOR3 (N2043, N2041, N47, N449);
xor XOR2 (N2044, N2031, N39);
not NOT1 (N2045, N2028);
or OR3 (N2046, N2038, N1514, N775);
xor XOR2 (N2047, N2043, N809);
and AND3 (N2048, N2044, N1781, N478);
buf BUF1 (N2049, N2046);
nor NOR2 (N2050, N2018, N261);
xor XOR2 (N2051, N2042, N1713);
not NOT1 (N2052, N2049);
buf BUF1 (N2053, N2050);
nor NOR3 (N2054, N2040, N1922, N759);
xor XOR2 (N2055, N2035, N1594);
and AND3 (N2056, N2027, N1372, N1326);
and AND2 (N2057, N2052, N874);
nand NAND2 (N2058, N2045, N152);
nor NOR2 (N2059, N2057, N1628);
and AND2 (N2060, N2058, N1758);
buf BUF1 (N2061, N2053);
buf BUF1 (N2062, N2054);
and AND3 (N2063, N2059, N395, N876);
or OR4 (N2064, N2055, N46, N856, N1123);
not NOT1 (N2065, N2048);
nor NOR3 (N2066, N2047, N670, N137);
xor XOR2 (N2067, N2061, N943);
nor NOR2 (N2068, N2036, N1097);
nor NOR2 (N2069, N2064, N1564);
buf BUF1 (N2070, N2051);
or OR4 (N2071, N2063, N1117, N1071, N1601);
and AND3 (N2072, N2065, N523, N1677);
xor XOR2 (N2073, N2071, N2015);
and AND3 (N2074, N2066, N209, N1709);
or OR3 (N2075, N2067, N915, N440);
or OR2 (N2076, N2072, N1367);
and AND3 (N2077, N2056, N1769, N1380);
nor NOR4 (N2078, N2068, N2003, N537, N1615);
and AND3 (N2079, N2062, N1412, N1487);
xor XOR2 (N2080, N2074, N58);
buf BUF1 (N2081, N2070);
nor NOR3 (N2082, N2080, N1047, N1404);
nand NAND2 (N2083, N2076, N1618);
not NOT1 (N2084, N2075);
and AND4 (N2085, N2060, N1697, N1279, N251);
not NOT1 (N2086, N2083);
xor XOR2 (N2087, N2073, N96);
nor NOR2 (N2088, N2078, N1192);
not NOT1 (N2089, N2087);
or OR2 (N2090, N2082, N1351);
or OR2 (N2091, N2084, N569);
nand NAND4 (N2092, N2086, N1748, N1056, N1232);
nand NAND3 (N2093, N2069, N1712, N1834);
nor NOR4 (N2094, N2085, N1336, N1795, N828);
or OR4 (N2095, N2077, N396, N1623, N302);
or OR4 (N2096, N2089, N505, N1312, N542);
buf BUF1 (N2097, N2096);
nand NAND4 (N2098, N2088, N1780, N315, N664);
not NOT1 (N2099, N2098);
nor NOR2 (N2100, N2091, N154);
nor NOR3 (N2101, N2097, N1196, N1731);
not NOT1 (N2102, N2090);
or OR3 (N2103, N2099, N1880, N1927);
xor XOR2 (N2104, N2081, N1699);
or OR4 (N2105, N2103, N1140, N315, N1741);
buf BUF1 (N2106, N2094);
or OR4 (N2107, N2095, N2004, N1339, N134);
or OR4 (N2108, N2100, N1629, N692, N1512);
not NOT1 (N2109, N2104);
xor XOR2 (N2110, N2093, N1357);
buf BUF1 (N2111, N2092);
or OR3 (N2112, N2108, N283, N24);
nor NOR3 (N2113, N2107, N1481, N1754);
nor NOR2 (N2114, N2079, N734);
or OR2 (N2115, N2114, N1495);
buf BUF1 (N2116, N2110);
or OR3 (N2117, N2105, N1619, N1625);
nand NAND3 (N2118, N2101, N1310, N1757);
buf BUF1 (N2119, N2118);
not NOT1 (N2120, N2102);
xor XOR2 (N2121, N2119, N116);
buf BUF1 (N2122, N2109);
nor NOR3 (N2123, N2117, N1771, N2002);
not NOT1 (N2124, N2116);
or OR4 (N2125, N2111, N183, N1790, N1779);
nor NOR4 (N2126, N2120, N52, N600, N503);
xor XOR2 (N2127, N2123, N1085);
or OR2 (N2128, N2127, N996);
buf BUF1 (N2129, N2121);
not NOT1 (N2130, N2122);
and AND3 (N2131, N2113, N1325, N1161);
xor XOR2 (N2132, N2125, N1253);
xor XOR2 (N2133, N2126, N1943);
buf BUF1 (N2134, N2129);
not NOT1 (N2135, N2130);
or OR3 (N2136, N2134, N442, N103);
nand NAND3 (N2137, N2112, N1050, N1898);
xor XOR2 (N2138, N2128, N574);
and AND2 (N2139, N2133, N1717);
not NOT1 (N2140, N2131);
not NOT1 (N2141, N2132);
buf BUF1 (N2142, N2138);
or OR3 (N2143, N2140, N534, N307);
nand NAND3 (N2144, N2137, N1040, N1460);
nor NOR3 (N2145, N2124, N2072, N1552);
xor XOR2 (N2146, N2115, N333);
and AND2 (N2147, N2106, N1402);
xor XOR2 (N2148, N2143, N634);
buf BUF1 (N2149, N2144);
not NOT1 (N2150, N2135);
and AND4 (N2151, N2150, N410, N8, N550);
nand NAND3 (N2152, N2146, N1996, N1590);
and AND3 (N2153, N2148, N534, N1522);
or OR3 (N2154, N2149, N453, N639);
buf BUF1 (N2155, N2142);
nand NAND4 (N2156, N2147, N1138, N169, N292);
nor NOR3 (N2157, N2156, N1266, N1597);
buf BUF1 (N2158, N2141);
or OR4 (N2159, N2151, N1669, N1762, N1775);
and AND3 (N2160, N2154, N209, N1411);
xor XOR2 (N2161, N2145, N1585);
buf BUF1 (N2162, N2136);
not NOT1 (N2163, N2157);
not NOT1 (N2164, N2162);
buf BUF1 (N2165, N2159);
or OR3 (N2166, N2164, N947, N439);
buf BUF1 (N2167, N2152);
not NOT1 (N2168, N2158);
or OR2 (N2169, N2168, N613);
buf BUF1 (N2170, N2153);
and AND2 (N2171, N2161, N1863);
and AND2 (N2172, N2155, N257);
nand NAND4 (N2173, N2166, N1753, N221, N1456);
or OR2 (N2174, N2171, N1716);
buf BUF1 (N2175, N2139);
nor NOR2 (N2176, N2160, N1907);
or OR3 (N2177, N2173, N1658, N1289);
and AND3 (N2178, N2176, N730, N1814);
nor NOR2 (N2179, N2167, N318);
nand NAND4 (N2180, N2169, N243, N63, N1432);
xor XOR2 (N2181, N2178, N762);
nor NOR4 (N2182, N2172, N380, N2151, N1227);
not NOT1 (N2183, N2175);
nor NOR3 (N2184, N2179, N1378, N1120);
buf BUF1 (N2185, N2184);
nor NOR4 (N2186, N2177, N1065, N153, N1169);
or OR4 (N2187, N2180, N17, N847, N207);
xor XOR2 (N2188, N2185, N890);
not NOT1 (N2189, N2188);
and AND3 (N2190, N2174, N1244, N385);
or OR3 (N2191, N2165, N1800, N1745);
or OR2 (N2192, N2187, N944);
nor NOR2 (N2193, N2170, N412);
and AND2 (N2194, N2192, N1294);
buf BUF1 (N2195, N2190);
nor NOR3 (N2196, N2194, N1833, N1144);
and AND4 (N2197, N2189, N1348, N929, N914);
buf BUF1 (N2198, N2195);
xor XOR2 (N2199, N2163, N1097);
nor NOR3 (N2200, N2183, N1961, N425);
nand NAND2 (N2201, N2181, N1533);
or OR2 (N2202, N2196, N1859);
or OR4 (N2203, N2198, N1863, N26, N132);
buf BUF1 (N2204, N2182);
buf BUF1 (N2205, N2201);
nand NAND2 (N2206, N2191, N1384);
buf BUF1 (N2207, N2186);
xor XOR2 (N2208, N2197, N922);
nor NOR4 (N2209, N2200, N1801, N267, N160);
nor NOR3 (N2210, N2203, N263, N1166);
and AND4 (N2211, N2204, N1855, N954, N1987);
nor NOR3 (N2212, N2199, N1375, N1789);
not NOT1 (N2213, N2211);
and AND2 (N2214, N2208, N623);
buf BUF1 (N2215, N2205);
and AND2 (N2216, N2209, N1705);
buf BUF1 (N2217, N2215);
not NOT1 (N2218, N2193);
and AND2 (N2219, N2213, N561);
xor XOR2 (N2220, N2207, N1843);
not NOT1 (N2221, N2202);
or OR3 (N2222, N2210, N2008, N1375);
not NOT1 (N2223, N2222);
and AND2 (N2224, N2221, N1183);
and AND4 (N2225, N2206, N385, N737, N1693);
and AND2 (N2226, N2219, N1627);
not NOT1 (N2227, N2216);
and AND2 (N2228, N2226, N257);
or OR3 (N2229, N2223, N111, N534);
nor NOR4 (N2230, N2212, N1470, N1732, N47);
buf BUF1 (N2231, N2230);
not NOT1 (N2232, N2227);
xor XOR2 (N2233, N2224, N1178);
and AND3 (N2234, N2220, N560, N1192);
nand NAND2 (N2235, N2232, N188);
or OR4 (N2236, N2217, N658, N1001, N2219);
xor XOR2 (N2237, N2214, N219);
or OR2 (N2238, N2233, N1338);
buf BUF1 (N2239, N2236);
or OR4 (N2240, N2225, N914, N289, N1906);
nor NOR3 (N2241, N2228, N2155, N1630);
or OR3 (N2242, N2241, N111, N2049);
buf BUF1 (N2243, N2218);
xor XOR2 (N2244, N2231, N1196);
or OR3 (N2245, N2242, N393, N2102);
and AND3 (N2246, N2245, N1192, N613);
or OR4 (N2247, N2239, N1654, N823, N1358);
not NOT1 (N2248, N2247);
or OR4 (N2249, N2229, N378, N1473, N1514);
nor NOR3 (N2250, N2237, N217, N2149);
nor NOR3 (N2251, N2238, N1661, N2036);
or OR3 (N2252, N2248, N721, N1472);
nor NOR2 (N2253, N2246, N1005);
nand NAND2 (N2254, N2234, N2);
nand NAND4 (N2255, N2240, N1065, N899, N809);
and AND4 (N2256, N2254, N2004, N1718, N1627);
nor NOR3 (N2257, N2256, N2178, N1392);
xor XOR2 (N2258, N2249, N1065);
and AND4 (N2259, N2258, N1520, N941, N1417);
or OR2 (N2260, N2244, N1064);
nand NAND3 (N2261, N2252, N423, N745);
nand NAND2 (N2262, N2235, N1644);
xor XOR2 (N2263, N2255, N567);
buf BUF1 (N2264, N2243);
nand NAND4 (N2265, N2251, N336, N2037, N2106);
nor NOR3 (N2266, N2265, N1394, N1493);
xor XOR2 (N2267, N2253, N1125);
buf BUF1 (N2268, N2261);
xor XOR2 (N2269, N2263, N1054);
nor NOR4 (N2270, N2269, N334, N2240, N780);
xor XOR2 (N2271, N2250, N1525);
xor XOR2 (N2272, N2264, N1555);
nor NOR3 (N2273, N2270, N2181, N317);
and AND4 (N2274, N2259, N1829, N944, N226);
and AND2 (N2275, N2273, N1898);
or OR2 (N2276, N2268, N1367);
and AND3 (N2277, N2271, N129, N760);
xor XOR2 (N2278, N2272, N656);
or OR3 (N2279, N2278, N718, N1558);
nor NOR3 (N2280, N2276, N638, N952);
xor XOR2 (N2281, N2279, N881);
nor NOR3 (N2282, N2275, N2124, N2259);
and AND4 (N2283, N2277, N208, N306, N1769);
and AND2 (N2284, N2280, N2230);
and AND4 (N2285, N2282, N806, N2040, N1948);
nand NAND4 (N2286, N2284, N1779, N536, N493);
not NOT1 (N2287, N2281);
or OR3 (N2288, N2274, N479, N336);
or OR3 (N2289, N2287, N1665, N278);
not NOT1 (N2290, N2283);
xor XOR2 (N2291, N2267, N793);
nand NAND4 (N2292, N2285, N1119, N1687, N1861);
or OR3 (N2293, N2260, N1701, N1610);
buf BUF1 (N2294, N2289);
nor NOR3 (N2295, N2262, N680, N1764);
nand NAND3 (N2296, N2291, N1920, N682);
buf BUF1 (N2297, N2266);
nor NOR3 (N2298, N2295, N1790, N2);
xor XOR2 (N2299, N2297, N165);
xor XOR2 (N2300, N2257, N2284);
nand NAND4 (N2301, N2296, N366, N928, N143);
nand NAND3 (N2302, N2294, N1344, N1817);
buf BUF1 (N2303, N2301);
nand NAND2 (N2304, N2292, N1873);
nor NOR4 (N2305, N2300, N1714, N2019, N1823);
or OR2 (N2306, N2302, N1489);
and AND3 (N2307, N2306, N598, N508);
not NOT1 (N2308, N2307);
not NOT1 (N2309, N2286);
or OR4 (N2310, N2303, N1597, N453, N1314);
nand NAND3 (N2311, N2288, N438, N1100);
not NOT1 (N2312, N2304);
or OR4 (N2313, N2293, N1782, N2125, N1411);
nor NOR2 (N2314, N2312, N1856);
not NOT1 (N2315, N2311);
nand NAND4 (N2316, N2314, N315, N204, N1223);
buf BUF1 (N2317, N2305);
not NOT1 (N2318, N2310);
and AND4 (N2319, N2316, N1, N757, N864);
xor XOR2 (N2320, N2315, N2127);
not NOT1 (N2321, N2308);
xor XOR2 (N2322, N2320, N242);
nor NOR4 (N2323, N2322, N1010, N894, N651);
nand NAND3 (N2324, N2313, N488, N2266);
xor XOR2 (N2325, N2318, N1065);
xor XOR2 (N2326, N2309, N595);
and AND3 (N2327, N2325, N1562, N2185);
and AND4 (N2328, N2324, N764, N1545, N1261);
buf BUF1 (N2329, N2323);
or OR2 (N2330, N2317, N1295);
or OR4 (N2331, N2328, N1339, N965, N1170);
xor XOR2 (N2332, N2321, N1787);
nand NAND4 (N2333, N2332, N1039, N136, N2235);
nor NOR4 (N2334, N2299, N1572, N76, N2194);
xor XOR2 (N2335, N2290, N1329);
not NOT1 (N2336, N2335);
not NOT1 (N2337, N2334);
buf BUF1 (N2338, N2319);
or OR3 (N2339, N2326, N2290, N1634);
not NOT1 (N2340, N2298);
nor NOR4 (N2341, N2339, N693, N34, N1294);
nor NOR2 (N2342, N2327, N205);
and AND2 (N2343, N2340, N405);
or OR2 (N2344, N2331, N296);
buf BUF1 (N2345, N2341);
or OR4 (N2346, N2329, N570, N242, N1824);
and AND3 (N2347, N2338, N2241, N401);
and AND2 (N2348, N2346, N1773);
nand NAND4 (N2349, N2345, N1467, N586, N1938);
nand NAND2 (N2350, N2344, N1288);
or OR2 (N2351, N2336, N476);
and AND4 (N2352, N2337, N513, N430, N2344);
nand NAND4 (N2353, N2347, N825, N1154, N296);
xor XOR2 (N2354, N2350, N1732);
not NOT1 (N2355, N2342);
nand NAND3 (N2356, N2354, N290, N2222);
not NOT1 (N2357, N2352);
nor NOR3 (N2358, N2353, N1302, N1111);
buf BUF1 (N2359, N2356);
not NOT1 (N2360, N2357);
buf BUF1 (N2361, N2343);
or OR4 (N2362, N2359, N1277, N206, N1);
nor NOR4 (N2363, N2330, N445, N1093, N1241);
or OR4 (N2364, N2355, N1638, N827, N2054);
nor NOR4 (N2365, N2358, N1202, N964, N1919);
nor NOR3 (N2366, N2361, N14, N1457);
and AND3 (N2367, N2333, N1620, N2140);
xor XOR2 (N2368, N2351, N1036);
nand NAND4 (N2369, N2363, N2056, N817, N325);
buf BUF1 (N2370, N2369);
buf BUF1 (N2371, N2367);
nor NOR2 (N2372, N2349, N514);
not NOT1 (N2373, N2362);
not NOT1 (N2374, N2372);
xor XOR2 (N2375, N2366, N2320);
xor XOR2 (N2376, N2348, N1378);
not NOT1 (N2377, N2360);
and AND4 (N2378, N2373, N1408, N1466, N7);
or OR4 (N2379, N2370, N2372, N33, N1548);
xor XOR2 (N2380, N2376, N783);
not NOT1 (N2381, N2364);
xor XOR2 (N2382, N2374, N1379);
not NOT1 (N2383, N2365);
buf BUF1 (N2384, N2383);
nand NAND2 (N2385, N2375, N305);
buf BUF1 (N2386, N2378);
nor NOR4 (N2387, N2384, N1964, N860, N752);
xor XOR2 (N2388, N2381, N46);
not NOT1 (N2389, N2371);
nor NOR3 (N2390, N2388, N1220, N862);
nor NOR3 (N2391, N2377, N1468, N354);
not NOT1 (N2392, N2380);
or OR2 (N2393, N2390, N903);
buf BUF1 (N2394, N2385);
nand NAND4 (N2395, N2394, N622, N1079, N1914);
xor XOR2 (N2396, N2392, N423);
and AND4 (N2397, N2368, N2372, N2358, N647);
nand NAND2 (N2398, N2396, N988);
xor XOR2 (N2399, N2391, N165);
nor NOR4 (N2400, N2399, N1073, N1429, N673);
nand NAND4 (N2401, N2395, N1833, N700, N1002);
xor XOR2 (N2402, N2400, N976);
nand NAND4 (N2403, N2393, N1101, N2285, N1601);
not NOT1 (N2404, N2398);
nor NOR2 (N2405, N2382, N1175);
xor XOR2 (N2406, N2387, N681);
and AND2 (N2407, N2404, N437);
nor NOR3 (N2408, N2379, N1175, N1361);
and AND3 (N2409, N2397, N1994, N1524);
buf BUF1 (N2410, N2407);
nand NAND2 (N2411, N2389, N2387);
xor XOR2 (N2412, N2386, N818);
and AND4 (N2413, N2410, N381, N2325, N1682);
and AND4 (N2414, N2406, N1637, N1977, N1075);
xor XOR2 (N2415, N2408, N1207);
nor NOR4 (N2416, N2411, N1691, N2236, N1302);
not NOT1 (N2417, N2401);
or OR2 (N2418, N2403, N870);
xor XOR2 (N2419, N2417, N716);
or OR2 (N2420, N2418, N1000);
xor XOR2 (N2421, N2416, N560);
or OR3 (N2422, N2409, N132, N2128);
buf BUF1 (N2423, N2419);
xor XOR2 (N2424, N2415, N349);
nand NAND4 (N2425, N2421, N2162, N2050, N2088);
not NOT1 (N2426, N2425);
xor XOR2 (N2427, N2420, N262);
or OR2 (N2428, N2412, N1235);
nand NAND3 (N2429, N2424, N2279, N288);
nor NOR4 (N2430, N2428, N2321, N2300, N421);
buf BUF1 (N2431, N2402);
and AND4 (N2432, N2430, N185, N1569, N520);
not NOT1 (N2433, N2405);
nand NAND4 (N2434, N2427, N2008, N868, N1299);
or OR4 (N2435, N2423, N1460, N865, N1194);
not NOT1 (N2436, N2413);
nor NOR4 (N2437, N2436, N1952, N285, N1060);
nor NOR2 (N2438, N2422, N703);
xor XOR2 (N2439, N2433, N652);
nor NOR3 (N2440, N2429, N1152, N845);
xor XOR2 (N2441, N2437, N2410);
buf BUF1 (N2442, N2434);
buf BUF1 (N2443, N2441);
nor NOR2 (N2444, N2414, N504);
nand NAND4 (N2445, N2432, N728, N724, N1525);
or OR4 (N2446, N2442, N1062, N2192, N1746);
buf BUF1 (N2447, N2435);
buf BUF1 (N2448, N2446);
and AND3 (N2449, N2440, N1465, N1995);
or OR3 (N2450, N2443, N615, N618);
and AND2 (N2451, N2426, N1466);
nor NOR3 (N2452, N2445, N255, N221);
or OR2 (N2453, N2451, N1245);
nor NOR3 (N2454, N2449, N940, N1780);
and AND2 (N2455, N2454, N769);
buf BUF1 (N2456, N2455);
nor NOR4 (N2457, N2456, N2196, N2264, N839);
nor NOR2 (N2458, N2431, N2456);
buf BUF1 (N2459, N2444);
nand NAND3 (N2460, N2453, N1337, N1904);
xor XOR2 (N2461, N2457, N965);
nand NAND4 (N2462, N2450, N247, N164, N848);
nor NOR2 (N2463, N2447, N1639);
nor NOR2 (N2464, N2448, N211);
nand NAND4 (N2465, N2460, N2041, N2409, N1511);
nand NAND3 (N2466, N2464, N2216, N1375);
and AND2 (N2467, N2458, N400);
xor XOR2 (N2468, N2465, N883);
not NOT1 (N2469, N2467);
and AND4 (N2470, N2438, N73, N2229, N718);
xor XOR2 (N2471, N2469, N980);
buf BUF1 (N2472, N2471);
nor NOR3 (N2473, N2452, N692, N1659);
nand NAND3 (N2474, N2470, N1134, N1122);
buf BUF1 (N2475, N2463);
nor NOR4 (N2476, N2474, N967, N707, N1323);
or OR2 (N2477, N2439, N1596);
buf BUF1 (N2478, N2466);
xor XOR2 (N2479, N2475, N1081);
or OR2 (N2480, N2478, N797);
buf BUF1 (N2481, N2479);
or OR2 (N2482, N2461, N1258);
not NOT1 (N2483, N2462);
and AND3 (N2484, N2468, N1443, N1272);
xor XOR2 (N2485, N2459, N1059);
buf BUF1 (N2486, N2481);
nor NOR4 (N2487, N2480, N1153, N1635, N1852);
not NOT1 (N2488, N2477);
buf BUF1 (N2489, N2473);
or OR3 (N2490, N2484, N231, N1537);
nand NAND3 (N2491, N2472, N752, N516);
buf BUF1 (N2492, N2476);
or OR2 (N2493, N2491, N299);
or OR4 (N2494, N2492, N440, N2402, N172);
or OR2 (N2495, N2488, N754);
and AND3 (N2496, N2495, N1892, N1161);
and AND4 (N2497, N2485, N2289, N1166, N1513);
or OR2 (N2498, N2494, N2155);
nand NAND2 (N2499, N2496, N386);
nand NAND4 (N2500, N2482, N2423, N1625, N1576);
nor NOR4 (N2501, N2489, N846, N14, N1801);
and AND2 (N2502, N2497, N718);
nand NAND4 (N2503, N2486, N1721, N2198, N2089);
nor NOR4 (N2504, N2501, N2405, N2130, N398);
or OR2 (N2505, N2490, N1543);
nand NAND4 (N2506, N2503, N2185, N103, N2231);
nor NOR4 (N2507, N2505, N2052, N1912, N2352);
xor XOR2 (N2508, N2483, N1368);
nand NAND3 (N2509, N2487, N127, N2329);
xor XOR2 (N2510, N2508, N1432);
or OR3 (N2511, N2507, N413, N358);
nor NOR3 (N2512, N2506, N673, N460);
not NOT1 (N2513, N2512);
buf BUF1 (N2514, N2509);
buf BUF1 (N2515, N2499);
or OR3 (N2516, N2502, N1162, N388);
nor NOR4 (N2517, N2513, N465, N1558, N2492);
or OR2 (N2518, N2500, N1467);
not NOT1 (N2519, N2510);
xor XOR2 (N2520, N2516, N1440);
and AND3 (N2521, N2493, N1979, N434);
nand NAND4 (N2522, N2520, N8, N1087, N2291);
nor NOR4 (N2523, N2504, N1845, N133, N177);
not NOT1 (N2524, N2515);
buf BUF1 (N2525, N2514);
buf BUF1 (N2526, N2518);
nand NAND3 (N2527, N2522, N1500, N2164);
not NOT1 (N2528, N2525);
and AND2 (N2529, N2526, N129);
and AND2 (N2530, N2511, N1551);
and AND4 (N2531, N2528, N1802, N317, N2378);
nor NOR3 (N2532, N2523, N1179, N491);
and AND2 (N2533, N2519, N508);
and AND4 (N2534, N2531, N742, N819, N536);
and AND2 (N2535, N2517, N2146);
and AND3 (N2536, N2534, N1353, N942);
buf BUF1 (N2537, N2535);
and AND4 (N2538, N2533, N232, N2058, N1351);
and AND2 (N2539, N2527, N135);
nand NAND2 (N2540, N2539, N1467);
not NOT1 (N2541, N2530);
nor NOR2 (N2542, N2541, N811);
xor XOR2 (N2543, N2538, N1906);
nor NOR2 (N2544, N2532, N364);
and AND2 (N2545, N2537, N118);
buf BUF1 (N2546, N2545);
or OR3 (N2547, N2546, N2174, N1621);
or OR2 (N2548, N2524, N774);
or OR3 (N2549, N2542, N1938, N476);
nor NOR2 (N2550, N2549, N1096);
buf BUF1 (N2551, N2498);
and AND4 (N2552, N2544, N2304, N1069, N1728);
or OR2 (N2553, N2521, N694);
not NOT1 (N2554, N2536);
nand NAND4 (N2555, N2529, N740, N330, N7);
buf BUF1 (N2556, N2543);
nand NAND3 (N2557, N2547, N1892, N1154);
and AND4 (N2558, N2553, N1836, N808, N2073);
buf BUF1 (N2559, N2551);
xor XOR2 (N2560, N2554, N2319);
not NOT1 (N2561, N2560);
nand NAND4 (N2562, N2550, N1971, N1376, N173);
not NOT1 (N2563, N2557);
xor XOR2 (N2564, N2556, N2478);
nor NOR4 (N2565, N2548, N1405, N303, N1804);
or OR2 (N2566, N2565, N1356);
nand NAND3 (N2567, N2563, N1879, N1750);
nor NOR2 (N2568, N2540, N1940);
and AND3 (N2569, N2566, N1681, N468);
and AND2 (N2570, N2558, N693);
and AND2 (N2571, N2559, N2005);
or OR3 (N2572, N2571, N1261, N2008);
xor XOR2 (N2573, N2561, N1301);
nor NOR2 (N2574, N2567, N421);
or OR4 (N2575, N2570, N826, N361, N2349);
and AND3 (N2576, N2569, N1189, N928);
xor XOR2 (N2577, N2575, N2418);
nor NOR2 (N2578, N2573, N2264);
or OR3 (N2579, N2555, N648, N1742);
nor NOR4 (N2580, N2572, N368, N915, N2277);
nand NAND2 (N2581, N2580, N2205);
buf BUF1 (N2582, N2578);
and AND2 (N2583, N2581, N1500);
not NOT1 (N2584, N2582);
not NOT1 (N2585, N2552);
and AND4 (N2586, N2568, N1540, N2063, N861);
not NOT1 (N2587, N2564);
not NOT1 (N2588, N2584);
xor XOR2 (N2589, N2574, N442);
nand NAND2 (N2590, N2587, N2014);
or OR2 (N2591, N2590, N1040);
and AND3 (N2592, N2583, N2223, N1403);
not NOT1 (N2593, N2577);
xor XOR2 (N2594, N2593, N422);
nand NAND2 (N2595, N2589, N2548);
or OR4 (N2596, N2576, N1139, N557, N713);
not NOT1 (N2597, N2586);
xor XOR2 (N2598, N2591, N1532);
and AND4 (N2599, N2588, N45, N2535, N1646);
xor XOR2 (N2600, N2599, N883);
or OR2 (N2601, N2600, N1005);
not NOT1 (N2602, N2597);
and AND4 (N2603, N2594, N61, N335, N952);
xor XOR2 (N2604, N2602, N2444);
buf BUF1 (N2605, N2585);
or OR4 (N2606, N2562, N594, N1949, N1047);
and AND3 (N2607, N2605, N555, N398);
xor XOR2 (N2608, N2579, N531);
xor XOR2 (N2609, N2607, N953);
xor XOR2 (N2610, N2598, N2580);
nor NOR3 (N2611, N2604, N1798, N2109);
nor NOR2 (N2612, N2603, N472);
not NOT1 (N2613, N2596);
not NOT1 (N2614, N2611);
buf BUF1 (N2615, N2613);
or OR3 (N2616, N2606, N1985, N711);
buf BUF1 (N2617, N2608);
nand NAND3 (N2618, N2616, N1721, N867);
not NOT1 (N2619, N2617);
nand NAND4 (N2620, N2614, N2414, N1723, N810);
or OR2 (N2621, N2620, N2285);
nor NOR3 (N2622, N2618, N676, N2295);
xor XOR2 (N2623, N2610, N1685);
not NOT1 (N2624, N2612);
xor XOR2 (N2625, N2619, N514);
or OR2 (N2626, N2592, N1882);
nor NOR2 (N2627, N2601, N1351);
not NOT1 (N2628, N2625);
not NOT1 (N2629, N2628);
or OR3 (N2630, N2622, N1052, N2337);
nor NOR4 (N2631, N2627, N1107, N1525, N2012);
xor XOR2 (N2632, N2629, N2307);
not NOT1 (N2633, N2632);
and AND2 (N2634, N2621, N1987);
or OR2 (N2635, N2624, N1461);
xor XOR2 (N2636, N2635, N95);
xor XOR2 (N2637, N2615, N1272);
buf BUF1 (N2638, N2626);
buf BUF1 (N2639, N2637);
or OR2 (N2640, N2631, N609);
nand NAND4 (N2641, N2633, N1842, N13, N2553);
xor XOR2 (N2642, N2640, N1199);
not NOT1 (N2643, N2641);
and AND3 (N2644, N2623, N1140, N952);
nand NAND4 (N2645, N2636, N1644, N2560, N2107);
nor NOR3 (N2646, N2609, N2620, N79);
not NOT1 (N2647, N2639);
nand NAND2 (N2648, N2644, N2319);
not NOT1 (N2649, N2595);
buf BUF1 (N2650, N2645);
xor XOR2 (N2651, N2630, N315);
and AND4 (N2652, N2643, N892, N1241, N1954);
xor XOR2 (N2653, N2650, N2569);
or OR3 (N2654, N2653, N1395, N196);
and AND4 (N2655, N2651, N370, N2474, N95);
nand NAND4 (N2656, N2648, N1910, N70, N225);
buf BUF1 (N2657, N2654);
and AND3 (N2658, N2652, N988, N2629);
and AND4 (N2659, N2658, N2656, N1545, N141);
and AND3 (N2660, N2361, N445, N1728);
not NOT1 (N2661, N2647);
or OR2 (N2662, N2659, N1440);
buf BUF1 (N2663, N2638);
or OR3 (N2664, N2662, N919, N2127);
xor XOR2 (N2665, N2634, N1421);
and AND4 (N2666, N2665, N1245, N657, N130);
buf BUF1 (N2667, N2661);
not NOT1 (N2668, N2663);
nor NOR4 (N2669, N2664, N1271, N1426, N1112);
nand NAND3 (N2670, N2666, N1342, N1501);
not NOT1 (N2671, N2667);
and AND2 (N2672, N2671, N1259);
nand NAND3 (N2673, N2642, N60, N167);
not NOT1 (N2674, N2657);
buf BUF1 (N2675, N2673);
nor NOR4 (N2676, N2674, N1235, N1151, N1288);
nand NAND3 (N2677, N2668, N239, N784);
not NOT1 (N2678, N2669);
nor NOR2 (N2679, N2655, N1549);
nor NOR2 (N2680, N2670, N271);
not NOT1 (N2681, N2676);
nand NAND3 (N2682, N2678, N2178, N2033);
or OR3 (N2683, N2680, N147, N558);
buf BUF1 (N2684, N2646);
nor NOR4 (N2685, N2684, N1550, N2062, N1534);
not NOT1 (N2686, N2685);
and AND2 (N2687, N2649, N2438);
buf BUF1 (N2688, N2682);
and AND2 (N2689, N2683, N878);
nor NOR2 (N2690, N2660, N1208);
and AND3 (N2691, N2672, N2138, N1352);
xor XOR2 (N2692, N2686, N39);
or OR4 (N2693, N2679, N1398, N660, N899);
nand NAND4 (N2694, N2692, N1238, N1468, N1127);
and AND3 (N2695, N2688, N1226, N953);
and AND2 (N2696, N2694, N853);
xor XOR2 (N2697, N2677, N120);
or OR4 (N2698, N2693, N1114, N1474, N782);
nor NOR2 (N2699, N2691, N1176);
not NOT1 (N2700, N2689);
not NOT1 (N2701, N2697);
or OR2 (N2702, N2698, N2520);
xor XOR2 (N2703, N2681, N501);
xor XOR2 (N2704, N2699, N1862);
and AND4 (N2705, N2696, N1340, N1252, N160);
buf BUF1 (N2706, N2704);
buf BUF1 (N2707, N2700);
and AND3 (N2708, N2706, N2592, N2599);
not NOT1 (N2709, N2705);
and AND2 (N2710, N2701, N2486);
buf BUF1 (N2711, N2675);
or OR3 (N2712, N2695, N2255, N391);
nor NOR2 (N2713, N2710, N2073);
not NOT1 (N2714, N2702);
nor NOR3 (N2715, N2707, N1299, N2482);
xor XOR2 (N2716, N2687, N820);
nand NAND3 (N2717, N2712, N1646, N264);
and AND4 (N2718, N2711, N206, N1098, N2395);
nor NOR4 (N2719, N2715, N301, N430, N2313);
nor NOR2 (N2720, N2690, N1796);
and AND3 (N2721, N2716, N1152, N1446);
not NOT1 (N2722, N2719);
and AND4 (N2723, N2721, N2275, N2245, N1075);
or OR3 (N2724, N2723, N2419, N1873);
nand NAND3 (N2725, N2722, N1412, N2223);
nor NOR3 (N2726, N2718, N2101, N1258);
xor XOR2 (N2727, N2717, N2353);
and AND4 (N2728, N2720, N161, N1711, N489);
xor XOR2 (N2729, N2713, N190);
or OR2 (N2730, N2724, N576);
not NOT1 (N2731, N2703);
nand NAND3 (N2732, N2729, N1956, N618);
not NOT1 (N2733, N2727);
buf BUF1 (N2734, N2714);
nor NOR3 (N2735, N2733, N1777, N1050);
xor XOR2 (N2736, N2731, N1394);
nand NAND4 (N2737, N2732, N992, N180, N733);
nor NOR4 (N2738, N2734, N31, N1550, N2477);
nand NAND2 (N2739, N2725, N704);
and AND2 (N2740, N2708, N1666);
buf BUF1 (N2741, N2737);
and AND4 (N2742, N2726, N533, N2252, N1302);
buf BUF1 (N2743, N2709);
or OR2 (N2744, N2738, N451);
not NOT1 (N2745, N2735);
xor XOR2 (N2746, N2739, N799);
and AND4 (N2747, N2730, N303, N1123, N1282);
xor XOR2 (N2748, N2744, N313);
xor XOR2 (N2749, N2736, N47);
xor XOR2 (N2750, N2748, N1139);
nor NOR2 (N2751, N2749, N624);
or OR3 (N2752, N2742, N2434, N1271);
and AND2 (N2753, N2746, N882);
buf BUF1 (N2754, N2750);
not NOT1 (N2755, N2753);
or OR3 (N2756, N2751, N2604, N1228);
xor XOR2 (N2757, N2743, N450);
nand NAND4 (N2758, N2740, N1390, N2446, N1709);
buf BUF1 (N2759, N2728);
and AND2 (N2760, N2758, N427);
nand NAND3 (N2761, N2747, N463, N2086);
nand NAND4 (N2762, N2760, N1819, N2326, N1457);
not NOT1 (N2763, N2745);
xor XOR2 (N2764, N2756, N2345);
or OR2 (N2765, N2755, N1661);
or OR2 (N2766, N2757, N951);
nand NAND3 (N2767, N2752, N1181, N60);
and AND4 (N2768, N2764, N2453, N2163, N1934);
xor XOR2 (N2769, N2741, N375);
or OR2 (N2770, N2763, N2244);
and AND2 (N2771, N2769, N2569);
buf BUF1 (N2772, N2766);
nor NOR4 (N2773, N2767, N1260, N2578, N2171);
nand NAND3 (N2774, N2772, N1459, N2248);
xor XOR2 (N2775, N2759, N123);
not NOT1 (N2776, N2768);
not NOT1 (N2777, N2775);
xor XOR2 (N2778, N2765, N133);
buf BUF1 (N2779, N2761);
buf BUF1 (N2780, N2773);
and AND2 (N2781, N2770, N447);
xor XOR2 (N2782, N2777, N102);
and AND4 (N2783, N2779, N1714, N2003, N2545);
and AND3 (N2784, N2781, N61, N1000);
buf BUF1 (N2785, N2783);
xor XOR2 (N2786, N2762, N1289);
xor XOR2 (N2787, N2780, N541);
and AND3 (N2788, N2754, N1213, N416);
or OR4 (N2789, N2782, N1878, N140, N1147);
nand NAND4 (N2790, N2788, N1685, N2231, N1828);
and AND4 (N2791, N2787, N1840, N1814, N2032);
buf BUF1 (N2792, N2784);
buf BUF1 (N2793, N2776);
nand NAND2 (N2794, N2792, N15);
nand NAND2 (N2795, N2786, N2731);
or OR3 (N2796, N2778, N2696, N2605);
or OR2 (N2797, N2790, N1991);
nand NAND4 (N2798, N2791, N2486, N20, N1465);
nor NOR2 (N2799, N2774, N2120);
nand NAND3 (N2800, N2793, N1609, N819);
or OR3 (N2801, N2798, N2777, N1836);
and AND3 (N2802, N2794, N2012, N534);
nor NOR4 (N2803, N2789, N1043, N1647, N1922);
and AND3 (N2804, N2771, N2067, N2066);
not NOT1 (N2805, N2795);
nor NOR3 (N2806, N2802, N710, N1330);
buf BUF1 (N2807, N2804);
or OR4 (N2808, N2797, N938, N2171, N1293);
or OR2 (N2809, N2785, N102);
nand NAND4 (N2810, N2807, N105, N898, N1605);
nand NAND4 (N2811, N2796, N1352, N157, N603);
or OR2 (N2812, N2811, N1250);
nand NAND4 (N2813, N2809, N2373, N1896, N1306);
and AND3 (N2814, N2803, N2389, N886);
and AND3 (N2815, N2813, N1659, N1910);
not NOT1 (N2816, N2812);
buf BUF1 (N2817, N2800);
nor NOR3 (N2818, N2814, N545, N2292);
buf BUF1 (N2819, N2806);
xor XOR2 (N2820, N2799, N707);
not NOT1 (N2821, N2817);
xor XOR2 (N2822, N2816, N410);
or OR4 (N2823, N2801, N1891, N2081, N588);
or OR4 (N2824, N2808, N1794, N2752, N953);
buf BUF1 (N2825, N2823);
buf BUF1 (N2826, N2825);
or OR3 (N2827, N2821, N79, N2108);
nand NAND2 (N2828, N2820, N1560);
or OR2 (N2829, N2819, N2734);
xor XOR2 (N2830, N2824, N906);
and AND3 (N2831, N2805, N1957, N968);
not NOT1 (N2832, N2818);
buf BUF1 (N2833, N2826);
nor NOR4 (N2834, N2832, N147, N2593, N699);
nand NAND4 (N2835, N2829, N1705, N299, N571);
or OR4 (N2836, N2834, N21, N1370, N728);
nand NAND3 (N2837, N2830, N803, N1273);
and AND4 (N2838, N2827, N1788, N896, N2326);
buf BUF1 (N2839, N2831);
not NOT1 (N2840, N2839);
not NOT1 (N2841, N2836);
and AND2 (N2842, N2815, N2359);
and AND2 (N2843, N2822, N706);
buf BUF1 (N2844, N2837);
xor XOR2 (N2845, N2840, N1196);
nor NOR3 (N2846, N2845, N2390, N414);
not NOT1 (N2847, N2842);
or OR2 (N2848, N2847, N1548);
buf BUF1 (N2849, N2833);
xor XOR2 (N2850, N2848, N930);
xor XOR2 (N2851, N2850, N2570);
and AND2 (N2852, N2851, N2024);
xor XOR2 (N2853, N2810, N555);
buf BUF1 (N2854, N2852);
xor XOR2 (N2855, N2828, N1619);
nand NAND3 (N2856, N2849, N206, N2565);
buf BUF1 (N2857, N2856);
nor NOR3 (N2858, N2843, N94, N1582);
and AND2 (N2859, N2841, N1258);
xor XOR2 (N2860, N2854, N868);
nand NAND4 (N2861, N2853, N1363, N1011, N1375);
or OR3 (N2862, N2835, N2570, N2197);
and AND3 (N2863, N2861, N1067, N592);
or OR4 (N2864, N2844, N1445, N1163, N2290);
nand NAND4 (N2865, N2859, N693, N591, N2433);
buf BUF1 (N2866, N2860);
nand NAND3 (N2867, N2855, N2553, N1546);
xor XOR2 (N2868, N2863, N628);
or OR4 (N2869, N2867, N1012, N761, N2287);
nand NAND2 (N2870, N2866, N158);
and AND4 (N2871, N2865, N860, N1655, N1953);
or OR3 (N2872, N2846, N770, N1844);
nor NOR4 (N2873, N2872, N878, N2515, N1783);
buf BUF1 (N2874, N2871);
or OR4 (N2875, N2874, N312, N957, N947);
or OR4 (N2876, N2864, N17, N2196, N1356);
or OR3 (N2877, N2857, N2198, N2213);
nand NAND4 (N2878, N2858, N636, N2490, N39);
buf BUF1 (N2879, N2870);
buf BUF1 (N2880, N2875);
nor NOR3 (N2881, N2877, N956, N2359);
buf BUF1 (N2882, N2879);
or OR4 (N2883, N2838, N1942, N1673, N138);
buf BUF1 (N2884, N2869);
not NOT1 (N2885, N2881);
nor NOR3 (N2886, N2885, N2766, N1818);
xor XOR2 (N2887, N2873, N1710);
nor NOR4 (N2888, N2887, N435, N1956, N1759);
buf BUF1 (N2889, N2862);
xor XOR2 (N2890, N2882, N729);
nand NAND2 (N2891, N2889, N565);
and AND3 (N2892, N2884, N299, N2699);
nand NAND3 (N2893, N2888, N1720, N2600);
nand NAND3 (N2894, N2891, N2185, N1452);
nand NAND3 (N2895, N2868, N2576, N667);
or OR2 (N2896, N2892, N2608);
nor NOR2 (N2897, N2883, N498);
nand NAND4 (N2898, N2878, N1381, N2058, N2559);
not NOT1 (N2899, N2886);
and AND2 (N2900, N2890, N770);
or OR2 (N2901, N2894, N2830);
nor NOR3 (N2902, N2897, N74, N105);
or OR2 (N2903, N2880, N398);
and AND2 (N2904, N2893, N24);
or OR4 (N2905, N2901, N644, N2707, N1529);
not NOT1 (N2906, N2900);
and AND3 (N2907, N2902, N2305, N1148);
and AND3 (N2908, N2903, N497, N2553);
not NOT1 (N2909, N2896);
nand NAND3 (N2910, N2905, N887, N186);
nor NOR4 (N2911, N2904, N2839, N1170, N2840);
nor NOR2 (N2912, N2906, N67);
nor NOR4 (N2913, N2907, N578, N1337, N317);
not NOT1 (N2914, N2895);
buf BUF1 (N2915, N2876);
buf BUF1 (N2916, N2909);
not NOT1 (N2917, N2912);
xor XOR2 (N2918, N2914, N2635);
buf BUF1 (N2919, N2908);
xor XOR2 (N2920, N2918, N2553);
xor XOR2 (N2921, N2920, N1516);
or OR3 (N2922, N2919, N584, N1170);
xor XOR2 (N2923, N2915, N391);
buf BUF1 (N2924, N2910);
nand NAND4 (N2925, N2913, N1350, N1407, N1164);
or OR2 (N2926, N2916, N781);
nor NOR3 (N2927, N2898, N1864, N2881);
and AND4 (N2928, N2922, N1884, N841, N1808);
xor XOR2 (N2929, N2923, N98);
xor XOR2 (N2930, N2926, N835);
not NOT1 (N2931, N2925);
nor NOR2 (N2932, N2921, N2517);
nand NAND2 (N2933, N2930, N558);
or OR3 (N2934, N2932, N2463, N746);
not NOT1 (N2935, N2934);
xor XOR2 (N2936, N2928, N215);
nand NAND2 (N2937, N2924, N2738);
and AND3 (N2938, N2933, N2530, N562);
nand NAND3 (N2939, N2935, N2256, N2027);
not NOT1 (N2940, N2917);
xor XOR2 (N2941, N2927, N2794);
nand NAND2 (N2942, N2911, N166);
not NOT1 (N2943, N2938);
and AND2 (N2944, N2937, N1458);
and AND4 (N2945, N2899, N2035, N953, N1519);
and AND2 (N2946, N2940, N2921);
nor NOR2 (N2947, N2943, N2642);
and AND3 (N2948, N2929, N859, N2766);
not NOT1 (N2949, N2947);
nor NOR3 (N2950, N2945, N1610, N1320);
nand NAND3 (N2951, N2941, N166, N609);
xor XOR2 (N2952, N2951, N966);
nor NOR3 (N2953, N2942, N1207, N1620);
nor NOR3 (N2954, N2939, N1068, N532);
and AND4 (N2955, N2953, N2333, N2289, N2524);
or OR3 (N2956, N2936, N486, N978);
nand NAND2 (N2957, N2946, N1000);
buf BUF1 (N2958, N2944);
xor XOR2 (N2959, N2958, N2072);
xor XOR2 (N2960, N2955, N1402);
or OR4 (N2961, N2948, N705, N199, N2447);
not NOT1 (N2962, N2960);
not NOT1 (N2963, N2952);
buf BUF1 (N2964, N2949);
nand NAND3 (N2965, N2957, N117, N1706);
xor XOR2 (N2966, N2962, N620);
buf BUF1 (N2967, N2965);
nand NAND2 (N2968, N2966, N123);
or OR4 (N2969, N2959, N924, N2845, N258);
or OR2 (N2970, N2963, N2866);
xor XOR2 (N2971, N2961, N1647);
buf BUF1 (N2972, N2964);
or OR4 (N2973, N2931, N2515, N953, N1593);
xor XOR2 (N2974, N2956, N1052);
buf BUF1 (N2975, N2974);
or OR3 (N2976, N2970, N512, N221);
or OR3 (N2977, N2972, N1065, N1904);
not NOT1 (N2978, N2967);
and AND4 (N2979, N2977, N728, N2635, N241);
buf BUF1 (N2980, N2950);
or OR2 (N2981, N2971, N2091);
buf BUF1 (N2982, N2976);
xor XOR2 (N2983, N2981, N1210);
or OR2 (N2984, N2954, N1939);
and AND3 (N2985, N2978, N663, N1476);
nand NAND3 (N2986, N2973, N2238, N521);
nand NAND3 (N2987, N2968, N643, N1994);
or OR2 (N2988, N2979, N2104);
and AND3 (N2989, N2987, N2978, N150);
not NOT1 (N2990, N2975);
nand NAND4 (N2991, N2989, N731, N2887, N1096);
and AND4 (N2992, N2980, N248, N18, N891);
or OR3 (N2993, N2983, N1701, N1159);
nor NOR2 (N2994, N2969, N1436);
nand NAND2 (N2995, N2992, N1677);
xor XOR2 (N2996, N2990, N2799);
xor XOR2 (N2997, N2994, N2959);
buf BUF1 (N2998, N2984);
xor XOR2 (N2999, N2988, N2855);
nand NAND2 (N3000, N2982, N2120);
buf BUF1 (N3001, N2999);
nor NOR2 (N3002, N2985, N1349);
and AND2 (N3003, N3002, N2040);
not NOT1 (N3004, N2998);
and AND2 (N3005, N2993, N2237);
nor NOR2 (N3006, N2997, N2245);
nand NAND4 (N3007, N3006, N2197, N358, N2313);
or OR3 (N3008, N3004, N2382, N2337);
nor NOR2 (N3009, N2995, N510);
or OR4 (N3010, N3001, N2696, N1493, N71);
nor NOR3 (N3011, N3007, N2825, N1483);
buf BUF1 (N3012, N3008);
xor XOR2 (N3013, N3012, N809);
buf BUF1 (N3014, N2996);
not NOT1 (N3015, N3000);
nand NAND3 (N3016, N3010, N2329, N839);
nor NOR4 (N3017, N3014, N2532, N78, N1723);
and AND4 (N3018, N3003, N978, N301, N2869);
xor XOR2 (N3019, N3009, N1502);
nor NOR3 (N3020, N2986, N2851, N394);
nor NOR3 (N3021, N3017, N1591, N2833);
buf BUF1 (N3022, N2991);
not NOT1 (N3023, N3018);
buf BUF1 (N3024, N3023);
buf BUF1 (N3025, N3024);
nand NAND2 (N3026, N3016, N2165);
nor NOR4 (N3027, N3013, N1520, N677, N1578);
not NOT1 (N3028, N3020);
not NOT1 (N3029, N3015);
xor XOR2 (N3030, N3011, N1246);
or OR3 (N3031, N3025, N675, N1681);
nand NAND4 (N3032, N3022, N2950, N789, N2928);
xor XOR2 (N3033, N3032, N850);
or OR2 (N3034, N3026, N2914);
nor NOR4 (N3035, N3033, N1720, N683, N2757);
buf BUF1 (N3036, N3019);
buf BUF1 (N3037, N3021);
buf BUF1 (N3038, N3027);
nor NOR4 (N3039, N3028, N1323, N1493, N287);
xor XOR2 (N3040, N3034, N711);
or OR4 (N3041, N3036, N1061, N1347, N1539);
nor NOR3 (N3042, N3005, N2725, N1305);
nor NOR4 (N3043, N3035, N175, N2947, N867);
nor NOR3 (N3044, N3030, N2055, N1408);
buf BUF1 (N3045, N3037);
nor NOR2 (N3046, N3042, N2586);
buf BUF1 (N3047, N3046);
buf BUF1 (N3048, N3031);
xor XOR2 (N3049, N3043, N610);
not NOT1 (N3050, N3040);
buf BUF1 (N3051, N3048);
nor NOR3 (N3052, N3038, N10, N2084);
or OR3 (N3053, N3049, N1160, N2520);
not NOT1 (N3054, N3039);
and AND2 (N3055, N3054, N809);
and AND3 (N3056, N3047, N983, N511);
or OR2 (N3057, N3051, N763);
and AND4 (N3058, N3053, N1979, N871, N1377);
or OR4 (N3059, N3050, N603, N2097, N2225);
or OR2 (N3060, N3058, N414);
and AND2 (N3061, N3045, N766);
nor NOR4 (N3062, N3057, N2052, N929, N2222);
and AND3 (N3063, N3061, N2305, N2466);
not NOT1 (N3064, N3044);
buf BUF1 (N3065, N3059);
or OR4 (N3066, N3052, N1668, N122, N3033);
or OR3 (N3067, N3041, N1864, N2504);
xor XOR2 (N3068, N3056, N724);
nor NOR2 (N3069, N3055, N2631);
buf BUF1 (N3070, N3068);
nor NOR2 (N3071, N3065, N2238);
or OR3 (N3072, N3029, N736, N2525);
and AND2 (N3073, N3072, N781);
nor NOR3 (N3074, N3062, N2418, N2396);
xor XOR2 (N3075, N3066, N347);
or OR4 (N3076, N3074, N229, N342, N810);
and AND3 (N3077, N3075, N3014, N1878);
not NOT1 (N3078, N3070);
nand NAND3 (N3079, N3064, N1190, N2289);
buf BUF1 (N3080, N3071);
buf BUF1 (N3081, N3069);
buf BUF1 (N3082, N3079);
not NOT1 (N3083, N3063);
buf BUF1 (N3084, N3060);
or OR2 (N3085, N3073, N2976);
or OR3 (N3086, N3084, N2135, N1525);
or OR4 (N3087, N3081, N1823, N2272, N1107);
nand NAND3 (N3088, N3085, N2648, N2907);
nor NOR3 (N3089, N3077, N1246, N2706);
buf BUF1 (N3090, N3067);
nor NOR3 (N3091, N3088, N36, N2694);
or OR2 (N3092, N3090, N821);
buf BUF1 (N3093, N3076);
and AND2 (N3094, N3093, N234);
buf BUF1 (N3095, N3091);
or OR2 (N3096, N3086, N67);
not NOT1 (N3097, N3078);
and AND4 (N3098, N3092, N2837, N2700, N2310);
or OR2 (N3099, N3083, N1963);
not NOT1 (N3100, N3080);
not NOT1 (N3101, N3098);
xor XOR2 (N3102, N3099, N214);
xor XOR2 (N3103, N3089, N837);
not NOT1 (N3104, N3095);
nor NOR4 (N3105, N3102, N2048, N2230, N1045);
buf BUF1 (N3106, N3096);
not NOT1 (N3107, N3097);
xor XOR2 (N3108, N3104, N1569);
and AND2 (N3109, N3107, N564);
not NOT1 (N3110, N3105);
nand NAND4 (N3111, N3082, N453, N543, N2092);
buf BUF1 (N3112, N3109);
nand NAND3 (N3113, N3100, N2336, N1336);
nor NOR3 (N3114, N3106, N1511, N1034);
xor XOR2 (N3115, N3094, N219);
buf BUF1 (N3116, N3115);
not NOT1 (N3117, N3111);
nand NAND2 (N3118, N3110, N2687);
and AND2 (N3119, N3116, N1519);
nor NOR2 (N3120, N3114, N1539);
or OR2 (N3121, N3117, N225);
xor XOR2 (N3122, N3113, N1442);
nand NAND3 (N3123, N3122, N60, N938);
nand NAND2 (N3124, N3121, N3022);
or OR4 (N3125, N3108, N2294, N723, N1308);
or OR3 (N3126, N3125, N1503, N1136);
or OR3 (N3127, N3112, N1579, N1334);
nand NAND3 (N3128, N3127, N980, N505);
nand NAND3 (N3129, N3119, N913, N2445);
and AND3 (N3130, N3101, N2781, N2751);
nand NAND2 (N3131, N3124, N1137);
buf BUF1 (N3132, N3131);
buf BUF1 (N3133, N3126);
buf BUF1 (N3134, N3130);
and AND2 (N3135, N3103, N632);
or OR4 (N3136, N3132, N262, N1664, N117);
nor NOR4 (N3137, N3136, N2795, N308, N2688);
nand NAND3 (N3138, N3137, N1440, N2226);
nor NOR3 (N3139, N3128, N2237, N1313);
nand NAND4 (N3140, N3133, N886, N2600, N126);
or OR3 (N3141, N3134, N2236, N653);
nor NOR4 (N3142, N3123, N2610, N1859, N2338);
and AND3 (N3143, N3139, N16, N574);
or OR2 (N3144, N3140, N2674);
nor NOR3 (N3145, N3138, N1119, N2106);
nand NAND2 (N3146, N3144, N2964);
or OR4 (N3147, N3145, N3138, N1575, N1153);
nand NAND3 (N3148, N3141, N1857, N3021);
nand NAND2 (N3149, N3146, N2847);
or OR4 (N3150, N3129, N985, N2973, N2813);
and AND4 (N3151, N3142, N475, N35, N1906);
or OR3 (N3152, N3135, N166, N1906);
xor XOR2 (N3153, N3151, N2515);
nor NOR2 (N3154, N3148, N1887);
nor NOR4 (N3155, N3147, N231, N3057, N2141);
or OR2 (N3156, N3152, N1640);
not NOT1 (N3157, N3153);
and AND2 (N3158, N3087, N2506);
or OR2 (N3159, N3156, N635);
nor NOR3 (N3160, N3154, N2152, N1377);
xor XOR2 (N3161, N3118, N2095);
and AND4 (N3162, N3161, N2841, N67, N3026);
and AND3 (N3163, N3149, N384, N2576);
buf BUF1 (N3164, N3150);
or OR2 (N3165, N3159, N2280);
nor NOR4 (N3166, N3164, N1161, N1657, N2456);
or OR4 (N3167, N3165, N1524, N1219, N2520);
not NOT1 (N3168, N3120);
or OR3 (N3169, N3160, N1608, N2617);
and AND4 (N3170, N3155, N3006, N2456, N2914);
not NOT1 (N3171, N3158);
or OR2 (N3172, N3171, N1392);
buf BUF1 (N3173, N3162);
buf BUF1 (N3174, N3168);
nor NOR3 (N3175, N3170, N303, N351);
buf BUF1 (N3176, N3157);
nand NAND2 (N3177, N3169, N2203);
or OR3 (N3178, N3176, N495, N2204);
xor XOR2 (N3179, N3178, N2727);
not NOT1 (N3180, N3173);
not NOT1 (N3181, N3177);
nor NOR4 (N3182, N3179, N1475, N1282, N257);
or OR4 (N3183, N3143, N644, N2278, N2180);
not NOT1 (N3184, N3174);
buf BUF1 (N3185, N3175);
nor NOR3 (N3186, N3163, N846, N685);
nand NAND2 (N3187, N3183, N612);
nand NAND4 (N3188, N3172, N224, N40, N3073);
nor NOR3 (N3189, N3180, N561, N2926);
nand NAND3 (N3190, N3187, N2093, N1092);
or OR3 (N3191, N3181, N2778, N889);
buf BUF1 (N3192, N3186);
and AND2 (N3193, N3188, N1202);
or OR2 (N3194, N3167, N1337);
not NOT1 (N3195, N3166);
nor NOR3 (N3196, N3182, N1544, N2733);
not NOT1 (N3197, N3194);
buf BUF1 (N3198, N3193);
or OR4 (N3199, N3184, N3100, N106, N2025);
not NOT1 (N3200, N3195);
or OR3 (N3201, N3189, N2093, N373);
xor XOR2 (N3202, N3190, N1438);
xor XOR2 (N3203, N3197, N1620);
xor XOR2 (N3204, N3191, N996);
buf BUF1 (N3205, N3204);
xor XOR2 (N3206, N3203, N2697);
and AND3 (N3207, N3205, N2098, N1976);
buf BUF1 (N3208, N3192);
xor XOR2 (N3209, N3202, N445);
not NOT1 (N3210, N3201);
nand NAND3 (N3211, N3208, N2757, N388);
buf BUF1 (N3212, N3211);
buf BUF1 (N3213, N3198);
and AND2 (N3214, N3207, N3081);
nand NAND2 (N3215, N3200, N1681);
nand NAND3 (N3216, N3199, N2386, N2162);
or OR4 (N3217, N3215, N1251, N2079, N1783);
nand NAND2 (N3218, N3217, N2593);
nand NAND4 (N3219, N3216, N1933, N1422, N468);
xor XOR2 (N3220, N3218, N3081);
and AND3 (N3221, N3214, N2904, N3141);
xor XOR2 (N3222, N3209, N1820);
or OR3 (N3223, N3220, N1702, N2840);
buf BUF1 (N3224, N3222);
not NOT1 (N3225, N3224);
and AND3 (N3226, N3221, N2836, N36);
or OR2 (N3227, N3206, N2272);
not NOT1 (N3228, N3196);
or OR2 (N3229, N3219, N3132);
nand NAND4 (N3230, N3227, N1623, N1004, N2872);
nand NAND3 (N3231, N3210, N2240, N324);
and AND2 (N3232, N3225, N649);
and AND2 (N3233, N3228, N2761);
xor XOR2 (N3234, N3231, N1803);
xor XOR2 (N3235, N3185, N658);
nand NAND2 (N3236, N3233, N3220);
nand NAND3 (N3237, N3229, N1034, N1706);
xor XOR2 (N3238, N3226, N399);
not NOT1 (N3239, N3238);
not NOT1 (N3240, N3235);
xor XOR2 (N3241, N3230, N3132);
or OR4 (N3242, N3223, N53, N1949, N190);
xor XOR2 (N3243, N3237, N2504);
not NOT1 (N3244, N3242);
or OR2 (N3245, N3236, N1764);
buf BUF1 (N3246, N3245);
nand NAND4 (N3247, N3246, N1052, N444, N1703);
xor XOR2 (N3248, N3240, N2273);
and AND3 (N3249, N3243, N2972, N209);
nor NOR3 (N3250, N3247, N2446, N1061);
and AND2 (N3251, N3248, N908);
and AND3 (N3252, N3249, N2796, N431);
and AND4 (N3253, N3232, N1376, N72, N1385);
and AND2 (N3254, N3239, N911);
xor XOR2 (N3255, N3213, N875);
or OR2 (N3256, N3254, N2467);
xor XOR2 (N3257, N3251, N875);
nand NAND3 (N3258, N3257, N1523, N532);
buf BUF1 (N3259, N3258);
and AND4 (N3260, N3259, N1983, N2295, N198);
nor NOR3 (N3261, N3244, N2836, N2501);
nand NAND2 (N3262, N3212, N1855);
nand NAND4 (N3263, N3253, N2000, N2114, N1114);
nor NOR2 (N3264, N3260, N2091);
xor XOR2 (N3265, N3261, N2653);
and AND2 (N3266, N3263, N1212);
nand NAND4 (N3267, N3256, N1681, N190, N1677);
nor NOR3 (N3268, N3265, N2279, N580);
nand NAND3 (N3269, N3264, N2409, N2257);
buf BUF1 (N3270, N3241);
and AND3 (N3271, N3234, N167, N1995);
not NOT1 (N3272, N3269);
nand NAND2 (N3273, N3272, N385);
nand NAND4 (N3274, N3266, N1629, N1581, N2926);
nor NOR2 (N3275, N3271, N1103);
nand NAND3 (N3276, N3255, N1456, N1244);
nor NOR4 (N3277, N3276, N2962, N87, N3249);
not NOT1 (N3278, N3262);
not NOT1 (N3279, N3278);
xor XOR2 (N3280, N3250, N2659);
buf BUF1 (N3281, N3280);
nor NOR4 (N3282, N3281, N3186, N278, N1526);
not NOT1 (N3283, N3270);
nand NAND3 (N3284, N3252, N2369, N833);
nand NAND3 (N3285, N3282, N2074, N1375);
nand NAND4 (N3286, N3274, N933, N2710, N1101);
nand NAND3 (N3287, N3273, N2422, N2836);
and AND3 (N3288, N3283, N211, N1442);
xor XOR2 (N3289, N3275, N1841);
not NOT1 (N3290, N3284);
nor NOR3 (N3291, N3287, N326, N258);
and AND3 (N3292, N3286, N1838, N1444);
and AND2 (N3293, N3291, N570);
not NOT1 (N3294, N3279);
buf BUF1 (N3295, N3289);
buf BUF1 (N3296, N3295);
nand NAND3 (N3297, N3277, N1997, N2392);
not NOT1 (N3298, N3293);
nand NAND3 (N3299, N3298, N2310, N1516);
buf BUF1 (N3300, N3285);
nor NOR2 (N3301, N3290, N440);
nand NAND2 (N3302, N3267, N223);
buf BUF1 (N3303, N3300);
nor NOR4 (N3304, N3302, N1684, N2829, N3012);
or OR2 (N3305, N3304, N2022);
or OR4 (N3306, N3299, N3019, N576, N1457);
xor XOR2 (N3307, N3306, N2626);
nand NAND2 (N3308, N3303, N2123);
nor NOR2 (N3309, N3308, N2164);
not NOT1 (N3310, N3307);
or OR3 (N3311, N3288, N2927, N3070);
nor NOR4 (N3312, N3301, N1280, N3263, N2030);
not NOT1 (N3313, N3268);
nor NOR2 (N3314, N3297, N1441);
xor XOR2 (N3315, N3294, N3298);
or OR4 (N3316, N3313, N3034, N2854, N2742);
nand NAND4 (N3317, N3296, N295, N554, N2870);
buf BUF1 (N3318, N3312);
buf BUF1 (N3319, N3317);
xor XOR2 (N3320, N3316, N446);
and AND2 (N3321, N3292, N564);
buf BUF1 (N3322, N3314);
or OR2 (N3323, N3321, N2594);
or OR2 (N3324, N3310, N388);
nor NOR3 (N3325, N3305, N1549, N1980);
nand NAND4 (N3326, N3320, N579, N2498, N2148);
buf BUF1 (N3327, N3323);
and AND3 (N3328, N3311, N2101, N560);
nand NAND2 (N3329, N3324, N465);
nand NAND3 (N3330, N3322, N430, N1715);
not NOT1 (N3331, N3327);
not NOT1 (N3332, N3331);
or OR2 (N3333, N3328, N1964);
and AND3 (N3334, N3319, N2974, N2031);
not NOT1 (N3335, N3330);
nand NAND3 (N3336, N3333, N679, N2456);
nor NOR2 (N3337, N3336, N1690);
xor XOR2 (N3338, N3309, N2562);
nand NAND2 (N3339, N3338, N1433);
not NOT1 (N3340, N3337);
nand NAND2 (N3341, N3339, N796);
nor NOR4 (N3342, N3318, N853, N2682, N2074);
nor NOR2 (N3343, N3329, N2632);
nand NAND4 (N3344, N3334, N629, N298, N2807);
nand NAND2 (N3345, N3344, N1153);
not NOT1 (N3346, N3343);
xor XOR2 (N3347, N3332, N1636);
nor NOR2 (N3348, N3345, N383);
nand NAND4 (N3349, N3341, N1780, N827, N2776);
nand NAND4 (N3350, N3346, N952, N1337, N2121);
and AND4 (N3351, N3325, N2990, N3153, N656);
and AND2 (N3352, N3335, N3112);
xor XOR2 (N3353, N3315, N392);
xor XOR2 (N3354, N3353, N2591);
or OR3 (N3355, N3326, N933, N1565);
nor NOR2 (N3356, N3342, N2425);
not NOT1 (N3357, N3349);
nor NOR4 (N3358, N3352, N1824, N1827, N2631);
nand NAND4 (N3359, N3350, N907, N2393, N1882);
nand NAND3 (N3360, N3348, N1411, N1257);
and AND2 (N3361, N3340, N1031);
buf BUF1 (N3362, N3357);
nor NOR4 (N3363, N3351, N2133, N3333, N2059);
or OR2 (N3364, N3361, N2234);
nand NAND3 (N3365, N3354, N1653, N1016);
not NOT1 (N3366, N3355);
not NOT1 (N3367, N3362);
nand NAND3 (N3368, N3367, N223, N2641);
nand NAND3 (N3369, N3360, N2672, N3103);
nor NOR4 (N3370, N3359, N2251, N895, N1673);
nor NOR4 (N3371, N3370, N2418, N144, N2553);
or OR4 (N3372, N3356, N1666, N1938, N2972);
buf BUF1 (N3373, N3347);
and AND4 (N3374, N3371, N2228, N523, N813);
buf BUF1 (N3375, N3364);
nand NAND3 (N3376, N3368, N1009, N2683);
buf BUF1 (N3377, N3358);
not NOT1 (N3378, N3373);
xor XOR2 (N3379, N3374, N2641);
or OR2 (N3380, N3365, N261);
nor NOR4 (N3381, N3379, N1612, N1457, N87);
xor XOR2 (N3382, N3376, N933);
not NOT1 (N3383, N3375);
and AND3 (N3384, N3378, N831, N1723);
and AND3 (N3385, N3366, N926, N2161);
buf BUF1 (N3386, N3363);
buf BUF1 (N3387, N3384);
nor NOR2 (N3388, N3385, N628);
and AND4 (N3389, N3388, N560, N428, N42);
xor XOR2 (N3390, N3383, N324);
nand NAND2 (N3391, N3390, N2897);
not NOT1 (N3392, N3382);
buf BUF1 (N3393, N3391);
and AND3 (N3394, N3386, N1712, N945);
nand NAND3 (N3395, N3392, N2995, N2815);
not NOT1 (N3396, N3372);
xor XOR2 (N3397, N3395, N2533);
or OR2 (N3398, N3380, N2659);
nand NAND2 (N3399, N3387, N2740);
nand NAND3 (N3400, N3398, N2777, N1631);
nor NOR4 (N3401, N3393, N3104, N2914, N3158);
or OR2 (N3402, N3396, N985);
nor NOR3 (N3403, N3402, N3007, N1432);
or OR4 (N3404, N3377, N2433, N1352, N895);
xor XOR2 (N3405, N3397, N2547);
not NOT1 (N3406, N3404);
buf BUF1 (N3407, N3406);
xor XOR2 (N3408, N3400, N2000);
nor NOR4 (N3409, N3405, N3321, N1234, N1324);
or OR2 (N3410, N3399, N1114);
xor XOR2 (N3411, N3381, N410);
nor NOR2 (N3412, N3408, N2793);
buf BUF1 (N3413, N3410);
nand NAND2 (N3414, N3407, N2392);
buf BUF1 (N3415, N3403);
and AND4 (N3416, N3413, N2186, N1439, N3104);
xor XOR2 (N3417, N3414, N2302);
and AND2 (N3418, N3411, N2136);
nor NOR4 (N3419, N3401, N165, N1130, N2714);
xor XOR2 (N3420, N3369, N2413);
xor XOR2 (N3421, N3419, N1167);
xor XOR2 (N3422, N3409, N3373);
nand NAND4 (N3423, N3422, N301, N760, N2580);
buf BUF1 (N3424, N3418);
or OR3 (N3425, N3420, N700, N2474);
nor NOR4 (N3426, N3415, N2625, N3393, N548);
not NOT1 (N3427, N3425);
nor NOR3 (N3428, N3423, N636, N1611);
buf BUF1 (N3429, N3421);
xor XOR2 (N3430, N3394, N2589);
and AND2 (N3431, N3417, N1931);
nand NAND2 (N3432, N3424, N3000);
not NOT1 (N3433, N3431);
or OR2 (N3434, N3429, N2856);
and AND4 (N3435, N3426, N668, N1059, N2907);
xor XOR2 (N3436, N3416, N1546);
or OR2 (N3437, N3412, N371);
or OR2 (N3438, N3427, N1908);
or OR2 (N3439, N3437, N167);
nor NOR4 (N3440, N3434, N3380, N3255, N1587);
xor XOR2 (N3441, N3436, N3437);
nor NOR3 (N3442, N3435, N2313, N3032);
or OR3 (N3443, N3441, N2585, N457);
not NOT1 (N3444, N3438);
nand NAND2 (N3445, N3442, N1524);
xor XOR2 (N3446, N3428, N1989);
xor XOR2 (N3447, N3439, N836);
nand NAND3 (N3448, N3430, N3272, N1564);
xor XOR2 (N3449, N3447, N2143);
nor NOR4 (N3450, N3444, N2258, N1072, N732);
nand NAND4 (N3451, N3432, N1800, N1575, N2794);
not NOT1 (N3452, N3449);
and AND3 (N3453, N3451, N2004, N305);
buf BUF1 (N3454, N3452);
nand NAND4 (N3455, N3454, N2893, N1162, N3204);
buf BUF1 (N3456, N3440);
buf BUF1 (N3457, N3443);
nor NOR3 (N3458, N3448, N3337, N3449);
nor NOR2 (N3459, N3453, N3068);
and AND3 (N3460, N3456, N2105, N2729);
nor NOR3 (N3461, N3389, N1122, N1296);
nor NOR2 (N3462, N3446, N1932);
not NOT1 (N3463, N3433);
or OR2 (N3464, N3457, N1480);
and AND2 (N3465, N3461, N2445);
or OR2 (N3466, N3445, N226);
nand NAND2 (N3467, N3459, N2327);
nor NOR3 (N3468, N3458, N1591, N1353);
xor XOR2 (N3469, N3465, N2077);
nor NOR3 (N3470, N3462, N1452, N3199);
and AND4 (N3471, N3468, N3393, N709, N1200);
and AND4 (N3472, N3471, N3375, N2363, N1048);
xor XOR2 (N3473, N3467, N1370);
and AND2 (N3474, N3460, N1562);
not NOT1 (N3475, N3450);
xor XOR2 (N3476, N3473, N1185);
nor NOR2 (N3477, N3469, N2828);
buf BUF1 (N3478, N3466);
and AND4 (N3479, N3472, N3163, N3085, N2682);
nand NAND2 (N3480, N3463, N457);
or OR3 (N3481, N3455, N3177, N1548);
not NOT1 (N3482, N3479);
not NOT1 (N3483, N3481);
not NOT1 (N3484, N3478);
not NOT1 (N3485, N3470);
buf BUF1 (N3486, N3483);
not NOT1 (N3487, N3476);
or OR3 (N3488, N3480, N1679, N2711);
not NOT1 (N3489, N3487);
nand NAND2 (N3490, N3484, N327);
or OR3 (N3491, N3475, N1930, N2423);
xor XOR2 (N3492, N3485, N1413);
buf BUF1 (N3493, N3491);
buf BUF1 (N3494, N3482);
nor NOR4 (N3495, N3474, N2842, N3218, N75);
and AND3 (N3496, N3464, N1681, N3105);
xor XOR2 (N3497, N3493, N1497);
buf BUF1 (N3498, N3490);
nor NOR4 (N3499, N3494, N613, N2431, N2395);
nand NAND3 (N3500, N3496, N839, N124);
xor XOR2 (N3501, N3498, N3376);
nand NAND2 (N3502, N3488, N105);
and AND2 (N3503, N3497, N878);
xor XOR2 (N3504, N3500, N1311);
buf BUF1 (N3505, N3477);
or OR2 (N3506, N3504, N2137);
xor XOR2 (N3507, N3499, N1349);
not NOT1 (N3508, N3486);
nand NAND4 (N3509, N3502, N1014, N2730, N843);
nand NAND4 (N3510, N3505, N3014, N544, N2540);
buf BUF1 (N3511, N3501);
or OR3 (N3512, N3492, N3454, N2844);
and AND2 (N3513, N3489, N1305);
and AND2 (N3514, N3507, N2947);
nand NAND2 (N3515, N3506, N2349);
xor XOR2 (N3516, N3513, N2669);
nor NOR3 (N3517, N3508, N1291, N1134);
or OR2 (N3518, N3511, N914);
not NOT1 (N3519, N3512);
nor NOR4 (N3520, N3509, N2725, N1350, N1267);
not NOT1 (N3521, N3517);
or OR3 (N3522, N3514, N1520, N1470);
or OR3 (N3523, N3521, N2984, N2435);
not NOT1 (N3524, N3510);
or OR4 (N3525, N3519, N3345, N3173, N2020);
buf BUF1 (N3526, N3522);
and AND4 (N3527, N3495, N1314, N1971, N2642);
not NOT1 (N3528, N3516);
or OR2 (N3529, N3520, N3106);
xor XOR2 (N3530, N3529, N1412);
or OR2 (N3531, N3526, N480);
and AND3 (N3532, N3518, N1009, N279);
xor XOR2 (N3533, N3515, N2704);
not NOT1 (N3534, N3527);
nor NOR3 (N3535, N3532, N1023, N1003);
or OR4 (N3536, N3525, N2559, N1260, N3413);
not NOT1 (N3537, N3503);
or OR2 (N3538, N3535, N663);
xor XOR2 (N3539, N3537, N168);
xor XOR2 (N3540, N3539, N3212);
nor NOR3 (N3541, N3528, N3397, N1834);
buf BUF1 (N3542, N3523);
xor XOR2 (N3543, N3540, N320);
nand NAND2 (N3544, N3533, N3285);
xor XOR2 (N3545, N3538, N850);
nand NAND3 (N3546, N3524, N3251, N1510);
buf BUF1 (N3547, N3534);
and AND4 (N3548, N3546, N256, N1358, N1707);
xor XOR2 (N3549, N3545, N735);
not NOT1 (N3550, N3547);
or OR3 (N3551, N3550, N1044, N1383);
buf BUF1 (N3552, N3531);
not NOT1 (N3553, N3548);
not NOT1 (N3554, N3553);
xor XOR2 (N3555, N3549, N2143);
nor NOR4 (N3556, N3555, N2841, N1645, N2119);
nand NAND3 (N3557, N3544, N1817, N1150);
or OR3 (N3558, N3556, N1458, N3205);
or OR2 (N3559, N3530, N1740);
not NOT1 (N3560, N3542);
nor NOR2 (N3561, N3551, N3363);
nand NAND3 (N3562, N3560, N642, N423);
xor XOR2 (N3563, N3541, N1340);
not NOT1 (N3564, N3557);
and AND4 (N3565, N3536, N2905, N1917, N3002);
nor NOR3 (N3566, N3543, N2700, N200);
and AND3 (N3567, N3562, N1312, N2327);
and AND3 (N3568, N3554, N3181, N1583);
not NOT1 (N3569, N3568);
buf BUF1 (N3570, N3566);
nand NAND2 (N3571, N3552, N1691);
and AND4 (N3572, N3567, N902, N1817, N3499);
or OR4 (N3573, N3559, N2112, N2802, N2972);
nand NAND2 (N3574, N3571, N1364);
nor NOR3 (N3575, N3565, N2806, N3230);
not NOT1 (N3576, N3575);
nor NOR4 (N3577, N3563, N1907, N2575, N421);
not NOT1 (N3578, N3572);
nor NOR3 (N3579, N3564, N2123, N2007);
buf BUF1 (N3580, N3579);
nor NOR4 (N3581, N3580, N676, N372, N1361);
not NOT1 (N3582, N3581);
nand NAND3 (N3583, N3577, N3228, N724);
and AND2 (N3584, N3570, N639);
and AND2 (N3585, N3582, N2837);
nor NOR3 (N3586, N3561, N303, N2900);
nand NAND3 (N3587, N3573, N2524, N2098);
xor XOR2 (N3588, N3578, N1515);
not NOT1 (N3589, N3574);
and AND4 (N3590, N3569, N1018, N3174, N2977);
nand NAND4 (N3591, N3586, N3461, N1513, N2370);
and AND4 (N3592, N3558, N1286, N2980, N987);
or OR4 (N3593, N3592, N3060, N950, N1603);
and AND2 (N3594, N3591, N1820);
not NOT1 (N3595, N3594);
xor XOR2 (N3596, N3576, N153);
and AND2 (N3597, N3589, N3442);
nor NOR4 (N3598, N3583, N854, N2055, N2251);
or OR2 (N3599, N3587, N2557);
xor XOR2 (N3600, N3593, N1768);
not NOT1 (N3601, N3598);
nand NAND2 (N3602, N3597, N39);
xor XOR2 (N3603, N3590, N1696);
and AND4 (N3604, N3601, N2318, N1160, N2288);
or OR4 (N3605, N3603, N3594, N740, N2392);
or OR4 (N3606, N3585, N1688, N1060, N3180);
nand NAND4 (N3607, N3584, N682, N2804, N2609);
not NOT1 (N3608, N3599);
not NOT1 (N3609, N3605);
xor XOR2 (N3610, N3608, N899);
not NOT1 (N3611, N3606);
nor NOR3 (N3612, N3611, N1659, N6);
xor XOR2 (N3613, N3596, N371);
not NOT1 (N3614, N3600);
buf BUF1 (N3615, N3595);
or OR2 (N3616, N3612, N3344);
and AND3 (N3617, N3604, N190, N646);
xor XOR2 (N3618, N3614, N3549);
and AND4 (N3619, N3607, N2148, N641, N3002);
buf BUF1 (N3620, N3609);
xor XOR2 (N3621, N3619, N545);
buf BUF1 (N3622, N3620);
not NOT1 (N3623, N3602);
not NOT1 (N3624, N3615);
not NOT1 (N3625, N3624);
and AND3 (N3626, N3610, N3451, N1725);
xor XOR2 (N3627, N3588, N890);
or OR3 (N3628, N3626, N1360, N765);
or OR4 (N3629, N3613, N1678, N1038, N370);
not NOT1 (N3630, N3616);
nand NAND4 (N3631, N3621, N1209, N1951, N2592);
buf BUF1 (N3632, N3630);
or OR3 (N3633, N3618, N2052, N555);
buf BUF1 (N3634, N3633);
xor XOR2 (N3635, N3631, N286);
buf BUF1 (N3636, N3627);
nor NOR2 (N3637, N3636, N2866);
xor XOR2 (N3638, N3628, N1105);
not NOT1 (N3639, N3632);
xor XOR2 (N3640, N3635, N1898);
xor XOR2 (N3641, N3622, N2588);
nand NAND3 (N3642, N3637, N1088, N2562);
not NOT1 (N3643, N3625);
not NOT1 (N3644, N3623);
not NOT1 (N3645, N3634);
xor XOR2 (N3646, N3642, N1152);
xor XOR2 (N3647, N3639, N406);
xor XOR2 (N3648, N3645, N2622);
not NOT1 (N3649, N3617);
nor NOR3 (N3650, N3649, N1885, N602);
nor NOR3 (N3651, N3629, N2287, N1727);
and AND2 (N3652, N3644, N6);
nand NAND3 (N3653, N3640, N3017, N776);
not NOT1 (N3654, N3641);
buf BUF1 (N3655, N3653);
buf BUF1 (N3656, N3647);
not NOT1 (N3657, N3646);
xor XOR2 (N3658, N3643, N2350);
not NOT1 (N3659, N3658);
not NOT1 (N3660, N3638);
nor NOR3 (N3661, N3648, N2255, N50);
or OR3 (N3662, N3650, N3510, N1887);
buf BUF1 (N3663, N3651);
buf BUF1 (N3664, N3663);
buf BUF1 (N3665, N3662);
not NOT1 (N3666, N3652);
nor NOR2 (N3667, N3664, N192);
not NOT1 (N3668, N3659);
buf BUF1 (N3669, N3660);
nand NAND3 (N3670, N3666, N2852, N3656);
nand NAND2 (N3671, N905, N2969);
or OR4 (N3672, N3655, N3640, N1854, N1288);
xor XOR2 (N3673, N3668, N669);
buf BUF1 (N3674, N3654);
nor NOR4 (N3675, N3672, N2151, N907, N317);
buf BUF1 (N3676, N3675);
buf BUF1 (N3677, N3671);
xor XOR2 (N3678, N3677, N2401);
not NOT1 (N3679, N3661);
or OR2 (N3680, N3679, N1442);
nand NAND4 (N3681, N3665, N3021, N1474, N702);
xor XOR2 (N3682, N3674, N1740);
or OR4 (N3683, N3678, N1382, N2042, N2123);
xor XOR2 (N3684, N3669, N368);
or OR2 (N3685, N3681, N1347);
not NOT1 (N3686, N3683);
and AND2 (N3687, N3673, N671);
nor NOR2 (N3688, N3657, N650);
nor NOR2 (N3689, N3687, N1980);
nor NOR2 (N3690, N3688, N1504);
xor XOR2 (N3691, N3682, N3560);
and AND2 (N3692, N3691, N2268);
and AND3 (N3693, N3676, N1377, N1177);
nand NAND4 (N3694, N3693, N576, N2029, N854);
nand NAND2 (N3695, N3689, N2813);
nor NOR2 (N3696, N3694, N3360);
nor NOR4 (N3697, N3680, N3364, N3324, N2043);
not NOT1 (N3698, N3692);
nor NOR4 (N3699, N3696, N2576, N58, N798);
or OR2 (N3700, N3684, N2183);
nand NAND4 (N3701, N3699, N1862, N1778, N2607);
or OR3 (N3702, N3701, N1495, N3683);
nor NOR3 (N3703, N3670, N3536, N844);
or OR4 (N3704, N3695, N1707, N2108, N948);
and AND3 (N3705, N3697, N2549, N771);
xor XOR2 (N3706, N3703, N3190);
not NOT1 (N3707, N3690);
xor XOR2 (N3708, N3700, N1790);
and AND2 (N3709, N3706, N1291);
or OR3 (N3710, N3686, N3494, N3348);
xor XOR2 (N3711, N3710, N1141);
and AND2 (N3712, N3667, N1523);
not NOT1 (N3713, N3702);
or OR4 (N3714, N3705, N3469, N2294, N44);
or OR4 (N3715, N3698, N209, N1346, N1022);
not NOT1 (N3716, N3709);
buf BUF1 (N3717, N3715);
nand NAND2 (N3718, N3713, N2875);
or OR3 (N3719, N3704, N2384, N1065);
nand NAND2 (N3720, N3712, N898);
or OR4 (N3721, N3720, N779, N1347, N2375);
buf BUF1 (N3722, N3707);
xor XOR2 (N3723, N3711, N2396);
nor NOR4 (N3724, N3719, N2668, N1156, N2621);
nor NOR3 (N3725, N3708, N3577, N3270);
or OR4 (N3726, N3685, N3368, N3674, N1951);
nand NAND4 (N3727, N3726, N272, N2901, N1283);
not NOT1 (N3728, N3723);
buf BUF1 (N3729, N3724);
nor NOR4 (N3730, N3718, N3251, N2983, N2471);
buf BUF1 (N3731, N3727);
xor XOR2 (N3732, N3717, N717);
and AND2 (N3733, N3728, N2874);
or OR3 (N3734, N3722, N1145, N158);
nor NOR2 (N3735, N3731, N2805);
buf BUF1 (N3736, N3721);
or OR3 (N3737, N3734, N3358, N2199);
and AND3 (N3738, N3725, N1047, N1399);
nand NAND3 (N3739, N3736, N506, N2180);
nand NAND2 (N3740, N3738, N1286);
not NOT1 (N3741, N3733);
not NOT1 (N3742, N3732);
and AND4 (N3743, N3739, N2471, N2647, N2401);
buf BUF1 (N3744, N3714);
and AND3 (N3745, N3741, N2686, N2774);
xor XOR2 (N3746, N3745, N2423);
buf BUF1 (N3747, N3740);
or OR3 (N3748, N3737, N1596, N1327);
and AND3 (N3749, N3747, N1196, N3239);
or OR2 (N3750, N3744, N1782);
not NOT1 (N3751, N3742);
or OR2 (N3752, N3748, N922);
buf BUF1 (N3753, N3743);
not NOT1 (N3754, N3730);
buf BUF1 (N3755, N3751);
nand NAND2 (N3756, N3754, N501);
or OR3 (N3757, N3755, N1879, N272);
buf BUF1 (N3758, N3752);
xor XOR2 (N3759, N3756, N2878);
nor NOR4 (N3760, N3729, N1855, N1509, N3473);
buf BUF1 (N3761, N3758);
xor XOR2 (N3762, N3750, N370);
not NOT1 (N3763, N3757);
buf BUF1 (N3764, N3746);
xor XOR2 (N3765, N3764, N1244);
and AND4 (N3766, N3759, N2086, N1803, N829);
nand NAND4 (N3767, N3762, N45, N1175, N1468);
and AND2 (N3768, N3765, N1588);
buf BUF1 (N3769, N3753);
buf BUF1 (N3770, N3767);
not NOT1 (N3771, N3749);
buf BUF1 (N3772, N3766);
nand NAND4 (N3773, N3770, N2974, N2440, N1508);
or OR4 (N3774, N3760, N3521, N3535, N3030);
or OR3 (N3775, N3773, N653, N389);
nor NOR2 (N3776, N3771, N357);
nor NOR2 (N3777, N3774, N2204);
buf BUF1 (N3778, N3761);
not NOT1 (N3779, N3735);
nand NAND2 (N3780, N3779, N3159);
buf BUF1 (N3781, N3775);
nor NOR3 (N3782, N3778, N3245, N2390);
and AND4 (N3783, N3763, N1962, N3178, N1078);
xor XOR2 (N3784, N3783, N2717);
not NOT1 (N3785, N3784);
or OR2 (N3786, N3782, N1031);
xor XOR2 (N3787, N3785, N2961);
nor NOR2 (N3788, N3772, N2468);
or OR2 (N3789, N3781, N238);
or OR2 (N3790, N3786, N3212);
buf BUF1 (N3791, N3716);
nand NAND2 (N3792, N3788, N3388);
nand NAND2 (N3793, N3776, N3536);
xor XOR2 (N3794, N3777, N2224);
and AND4 (N3795, N3769, N3643, N3243, N76);
xor XOR2 (N3796, N3780, N2031);
buf BUF1 (N3797, N3787);
or OR4 (N3798, N3797, N1367, N1347, N1968);
and AND4 (N3799, N3796, N1551, N843, N1162);
nor NOR3 (N3800, N3792, N1277, N3408);
nand NAND4 (N3801, N3799, N2259, N98, N801);
nand NAND4 (N3802, N3800, N1555, N2695, N2403);
and AND4 (N3803, N3768, N943, N2055, N1500);
nand NAND4 (N3804, N3801, N1817, N3763, N2623);
xor XOR2 (N3805, N3803, N2310);
nand NAND4 (N3806, N3798, N2405, N512, N2062);
and AND2 (N3807, N3804, N2454);
nand NAND4 (N3808, N3794, N135, N3265, N998);
nor NOR2 (N3809, N3807, N3397);
nand NAND2 (N3810, N3789, N1157);
nor NOR2 (N3811, N3808, N1379);
or OR4 (N3812, N3809, N1240, N1444, N526);
nand NAND4 (N3813, N3793, N2650, N1097, N2799);
and AND2 (N3814, N3811, N1811);
not NOT1 (N3815, N3805);
or OR4 (N3816, N3795, N2715, N1562, N2000);
nand NAND3 (N3817, N3802, N3726, N1043);
and AND4 (N3818, N3817, N2825, N2837, N1447);
xor XOR2 (N3819, N3812, N3667);
and AND3 (N3820, N3813, N1706, N1448);
or OR4 (N3821, N3818, N182, N2877, N244);
not NOT1 (N3822, N3791);
nand NAND4 (N3823, N3819, N1092, N772, N3169);
buf BUF1 (N3824, N3823);
not NOT1 (N3825, N3806);
not NOT1 (N3826, N3820);
nor NOR3 (N3827, N3790, N587, N1822);
nor NOR4 (N3828, N3810, N1231, N3581, N1814);
or OR3 (N3829, N3826, N3456, N2925);
and AND3 (N3830, N3814, N1758, N472);
or OR4 (N3831, N3822, N1234, N2568, N1343);
nand NAND2 (N3832, N3827, N3342);
buf BUF1 (N3833, N3816);
not NOT1 (N3834, N3829);
nand NAND4 (N3835, N3824, N1011, N3771, N3631);
and AND3 (N3836, N3833, N2948, N1696);
buf BUF1 (N3837, N3825);
buf BUF1 (N3838, N3821);
nand NAND4 (N3839, N3836, N3409, N3141, N355);
not NOT1 (N3840, N3831);
not NOT1 (N3841, N3834);
nand NAND2 (N3842, N3830, N1525);
buf BUF1 (N3843, N3837);
nor NOR2 (N3844, N3832, N2639);
nor NOR3 (N3845, N3835, N2867, N274);
and AND2 (N3846, N3839, N3030);
buf BUF1 (N3847, N3846);
xor XOR2 (N3848, N3815, N3345);
nand NAND3 (N3849, N3841, N2976, N3419);
nor NOR2 (N3850, N3845, N3293);
buf BUF1 (N3851, N3843);
or OR2 (N3852, N3848, N2332);
nor NOR2 (N3853, N3844, N3614);
or OR2 (N3854, N3853, N1845);
or OR2 (N3855, N3849, N1839);
not NOT1 (N3856, N3850);
buf BUF1 (N3857, N3852);
nor NOR2 (N3858, N3838, N1924);
nor NOR2 (N3859, N3857, N513);
xor XOR2 (N3860, N3854, N1714);
buf BUF1 (N3861, N3859);
or OR4 (N3862, N3861, N3041, N2083, N3312);
nand NAND4 (N3863, N3842, N2680, N3775, N137);
and AND3 (N3864, N3840, N2281, N3376);
nand NAND3 (N3865, N3862, N3567, N2055);
xor XOR2 (N3866, N3858, N577);
not NOT1 (N3867, N3847);
or OR3 (N3868, N3828, N3622, N1911);
nor NOR2 (N3869, N3856, N3604);
nand NAND2 (N3870, N3864, N240);
xor XOR2 (N3871, N3867, N1815);
xor XOR2 (N3872, N3869, N3420);
xor XOR2 (N3873, N3870, N2449);
buf BUF1 (N3874, N3866);
xor XOR2 (N3875, N3871, N78);
xor XOR2 (N3876, N3860, N214);
nor NOR4 (N3877, N3865, N223, N1686, N3671);
and AND2 (N3878, N3874, N3342);
nor NOR3 (N3879, N3855, N168, N3777);
and AND4 (N3880, N3868, N319, N131, N2678);
xor XOR2 (N3881, N3878, N47);
buf BUF1 (N3882, N3863);
and AND2 (N3883, N3880, N68);
nor NOR3 (N3884, N3881, N3357, N3607);
or OR4 (N3885, N3872, N3713, N3878, N3381);
and AND4 (N3886, N3882, N1243, N3651, N113);
nand NAND4 (N3887, N3885, N157, N2014, N3458);
nand NAND2 (N3888, N3884, N1506);
buf BUF1 (N3889, N3887);
nand NAND3 (N3890, N3851, N3629, N87);
or OR3 (N3891, N3876, N3719, N3806);
buf BUF1 (N3892, N3877);
not NOT1 (N3893, N3873);
xor XOR2 (N3894, N3879, N1126);
buf BUF1 (N3895, N3892);
not NOT1 (N3896, N3889);
nand NAND3 (N3897, N3886, N880, N608);
not NOT1 (N3898, N3894);
nor NOR4 (N3899, N3890, N622, N606, N3886);
xor XOR2 (N3900, N3883, N1605);
and AND2 (N3901, N3899, N2009);
and AND3 (N3902, N3897, N359, N1534);
xor XOR2 (N3903, N3888, N2416);
xor XOR2 (N3904, N3893, N60);
buf BUF1 (N3905, N3891);
nand NAND2 (N3906, N3902, N3266);
or OR4 (N3907, N3905, N1138, N714, N3317);
xor XOR2 (N3908, N3875, N299);
buf BUF1 (N3909, N3898);
nor NOR4 (N3910, N3907, N1515, N1780, N3066);
xor XOR2 (N3911, N3901, N1295);
xor XOR2 (N3912, N3903, N1270);
and AND3 (N3913, N3909, N103, N3186);
nand NAND4 (N3914, N3896, N1289, N2635, N507);
not NOT1 (N3915, N3900);
nor NOR4 (N3916, N3912, N497, N1190, N3618);
nor NOR2 (N3917, N3910, N81);
or OR2 (N3918, N3895, N517);
nand NAND2 (N3919, N3911, N1570);
nor NOR4 (N3920, N3914, N3831, N2859, N697);
nand NAND3 (N3921, N3916, N1893, N954);
buf BUF1 (N3922, N3919);
and AND4 (N3923, N3913, N910, N2364, N2985);
or OR3 (N3924, N3918, N530, N2203);
or OR4 (N3925, N3906, N1985, N3310, N1582);
xor XOR2 (N3926, N3922, N2850);
buf BUF1 (N3927, N3920);
xor XOR2 (N3928, N3921, N3420);
and AND3 (N3929, N3924, N1944, N18);
buf BUF1 (N3930, N3923);
and AND2 (N3931, N3930, N3142);
nor NOR4 (N3932, N3931, N1750, N301, N882);
buf BUF1 (N3933, N3927);
not NOT1 (N3934, N3908);
buf BUF1 (N3935, N3915);
or OR4 (N3936, N3932, N3247, N3111, N1484);
buf BUF1 (N3937, N3933);
xor XOR2 (N3938, N3929, N1690);
or OR4 (N3939, N3917, N3912, N675, N341);
nor NOR4 (N3940, N3928, N2231, N1170, N2271);
and AND2 (N3941, N3939, N461);
not NOT1 (N3942, N3936);
nand NAND3 (N3943, N3940, N3246, N1092);
and AND2 (N3944, N3935, N2449);
nor NOR3 (N3945, N3942, N3847, N95);
nand NAND2 (N3946, N3926, N3620);
or OR3 (N3947, N3904, N2270, N820);
buf BUF1 (N3948, N3941);
and AND4 (N3949, N3937, N2724, N3010, N788);
xor XOR2 (N3950, N3948, N1760);
nand NAND2 (N3951, N3947, N3576);
xor XOR2 (N3952, N3945, N3724);
xor XOR2 (N3953, N3946, N1507);
nor NOR3 (N3954, N3934, N2759, N1584);
nand NAND2 (N3955, N3954, N1421);
and AND3 (N3956, N3950, N249, N2741);
nor NOR3 (N3957, N3949, N2598, N2910);
xor XOR2 (N3958, N3952, N1822);
or OR2 (N3959, N3958, N3677);
or OR4 (N3960, N3956, N1976, N2580, N3858);
not NOT1 (N3961, N3957);
buf BUF1 (N3962, N3961);
and AND4 (N3963, N3953, N2467, N1556, N3353);
or OR2 (N3964, N3960, N2728);
nand NAND4 (N3965, N3955, N3497, N722, N383);
xor XOR2 (N3966, N3943, N165);
buf BUF1 (N3967, N3963);
nand NAND3 (N3968, N3944, N3315, N2839);
and AND3 (N3969, N3967, N3624, N2566);
xor XOR2 (N3970, N3959, N2568);
buf BUF1 (N3971, N3965);
or OR2 (N3972, N3970, N2297);
buf BUF1 (N3973, N3925);
or OR2 (N3974, N3966, N2253);
xor XOR2 (N3975, N3962, N2088);
not NOT1 (N3976, N3975);
or OR2 (N3977, N3951, N878);
xor XOR2 (N3978, N3938, N618);
and AND3 (N3979, N3969, N897, N1265);
nand NAND2 (N3980, N3973, N2918);
or OR4 (N3981, N3971, N3381, N2958, N2319);
nor NOR2 (N3982, N3981, N1933);
nor NOR3 (N3983, N3979, N453, N3857);
xor XOR2 (N3984, N3972, N2355);
xor XOR2 (N3985, N3983, N1180);
nand NAND4 (N3986, N3964, N463, N263, N1677);
not NOT1 (N3987, N3984);
and AND4 (N3988, N3987, N3880, N2578, N3838);
xor XOR2 (N3989, N3980, N787);
xor XOR2 (N3990, N3968, N970);
nand NAND4 (N3991, N3974, N3786, N2809, N3646);
buf BUF1 (N3992, N3991);
nand NAND3 (N3993, N3990, N1958, N3709);
nand NAND4 (N3994, N3978, N854, N2773, N1518);
and AND3 (N3995, N3977, N513, N132);
and AND3 (N3996, N3989, N2663, N2442);
nand NAND2 (N3997, N3996, N1883);
buf BUF1 (N3998, N3995);
or OR2 (N3999, N3993, N632);
or OR4 (N4000, N3998, N2898, N1518, N1109);
nor NOR2 (N4001, N3994, N895);
or OR2 (N4002, N3976, N3835);
nor NOR3 (N4003, N3982, N739, N1241);
or OR3 (N4004, N4001, N3286, N1546);
not NOT1 (N4005, N3985);
or OR2 (N4006, N3986, N2966);
or OR2 (N4007, N4006, N3030);
buf BUF1 (N4008, N4000);
and AND3 (N4009, N4005, N1142, N3578);
not NOT1 (N4010, N3992);
buf BUF1 (N4011, N3997);
buf BUF1 (N4012, N4008);
or OR4 (N4013, N4009, N1412, N2892, N3052);
or OR2 (N4014, N4002, N2090);
xor XOR2 (N4015, N4012, N3696);
buf BUF1 (N4016, N3999);
nand NAND3 (N4017, N4007, N2195, N1955);
nand NAND3 (N4018, N4003, N2481, N414);
or OR4 (N4019, N4015, N2507, N3027, N764);
and AND2 (N4020, N4019, N258);
nand NAND3 (N4021, N4014, N1519, N2909);
buf BUF1 (N4022, N4011);
buf BUF1 (N4023, N3988);
buf BUF1 (N4024, N4016);
or OR3 (N4025, N4017, N2576, N3995);
buf BUF1 (N4026, N4021);
and AND4 (N4027, N4025, N1434, N1107, N2085);
not NOT1 (N4028, N4022);
buf BUF1 (N4029, N4028);
nand NAND2 (N4030, N4010, N1070);
buf BUF1 (N4031, N4004);
nand NAND4 (N4032, N4020, N3335, N769, N3993);
or OR2 (N4033, N4030, N3021);
xor XOR2 (N4034, N4029, N1528);
or OR2 (N4035, N4027, N2974);
buf BUF1 (N4036, N4023);
nor NOR2 (N4037, N4034, N779);
and AND3 (N4038, N4026, N3351, N3033);
or OR2 (N4039, N4038, N3708);
buf BUF1 (N4040, N4018);
xor XOR2 (N4041, N4035, N1251);
nand NAND4 (N4042, N4036, N645, N987, N2493);
nand NAND2 (N4043, N4013, N1067);
or OR4 (N4044, N4024, N857, N3096, N1090);
xor XOR2 (N4045, N4041, N3819);
not NOT1 (N4046, N4040);
buf BUF1 (N4047, N4044);
xor XOR2 (N4048, N4047, N3515);
and AND3 (N4049, N4046, N3737, N290);
nand NAND3 (N4050, N4049, N973, N794);
nand NAND3 (N4051, N4048, N383, N3745);
buf BUF1 (N4052, N4045);
or OR4 (N4053, N4033, N1826, N1467, N3160);
xor XOR2 (N4054, N4031, N2868);
buf BUF1 (N4055, N4039);
and AND4 (N4056, N4053, N1927, N3072, N2361);
xor XOR2 (N4057, N4043, N2812);
nor NOR2 (N4058, N4051, N2032);
not NOT1 (N4059, N4056);
or OR4 (N4060, N4042, N575, N54, N3130);
buf BUF1 (N4061, N4050);
buf BUF1 (N4062, N4037);
and AND4 (N4063, N4061, N1699, N724, N2283);
xor XOR2 (N4064, N4060, N379);
xor XOR2 (N4065, N4059, N2597);
nand NAND3 (N4066, N4058, N2003, N2156);
xor XOR2 (N4067, N4055, N699);
nor NOR3 (N4068, N4057, N301, N281);
not NOT1 (N4069, N4068);
or OR3 (N4070, N4066, N4040, N245);
not NOT1 (N4071, N4052);
and AND2 (N4072, N4065, N3961);
nand NAND3 (N4073, N4032, N105, N1372);
nor NOR4 (N4074, N4071, N1407, N2444, N2433);
or OR4 (N4075, N4062, N740, N3706, N2745);
not NOT1 (N4076, N4072);
nor NOR4 (N4077, N4069, N1573, N2108, N3525);
nor NOR3 (N4078, N4054, N3856, N640);
nor NOR2 (N4079, N4075, N1873);
and AND3 (N4080, N4076, N2080, N1767);
and AND4 (N4081, N4079, N981, N3798, N611);
or OR4 (N4082, N4073, N3828, N2285, N1535);
and AND4 (N4083, N4070, N3652, N1589, N1710);
xor XOR2 (N4084, N4063, N2531);
or OR2 (N4085, N4064, N764);
or OR4 (N4086, N4080, N3951, N507, N819);
buf BUF1 (N4087, N4081);
not NOT1 (N4088, N4077);
nor NOR4 (N4089, N4088, N3568, N3018, N3344);
nand NAND3 (N4090, N4082, N2687, N2446);
buf BUF1 (N4091, N4086);
buf BUF1 (N4092, N4085);
not NOT1 (N4093, N4078);
or OR4 (N4094, N4087, N3488, N3250, N2784);
not NOT1 (N4095, N4084);
or OR2 (N4096, N4092, N2325);
nor NOR2 (N4097, N4096, N2652);
and AND2 (N4098, N4091, N154);
or OR3 (N4099, N4067, N870, N2296);
and AND4 (N4100, N4089, N2119, N685, N2198);
buf BUF1 (N4101, N4093);
not NOT1 (N4102, N4098);
and AND4 (N4103, N4074, N2456, N189, N1116);
xor XOR2 (N4104, N4101, N2258);
nor NOR3 (N4105, N4083, N2600, N807);
xor XOR2 (N4106, N4105, N3286);
xor XOR2 (N4107, N4099, N2992);
and AND4 (N4108, N4103, N3182, N957, N191);
nor NOR3 (N4109, N4108, N3973, N3884);
nand NAND4 (N4110, N4100, N1633, N3470, N323);
not NOT1 (N4111, N4102);
nor NOR4 (N4112, N4094, N2652, N2039, N2663);
nand NAND2 (N4113, N4095, N354);
xor XOR2 (N4114, N4104, N3635);
xor XOR2 (N4115, N4111, N1352);
not NOT1 (N4116, N4114);
and AND3 (N4117, N4090, N2763, N3098);
not NOT1 (N4118, N4110);
and AND3 (N4119, N4115, N142, N2688);
or OR3 (N4120, N4109, N2886, N155);
not NOT1 (N4121, N4112);
xor XOR2 (N4122, N4107, N1981);
nand NAND2 (N4123, N4118, N1082);
or OR2 (N4124, N4117, N271);
or OR3 (N4125, N4122, N2264, N2558);
buf BUF1 (N4126, N4097);
nor NOR3 (N4127, N4113, N3495, N2026);
nor NOR4 (N4128, N4126, N557, N2567, N820);
not NOT1 (N4129, N4124);
or OR3 (N4130, N4125, N3547, N3301);
and AND3 (N4131, N4130, N1270, N1502);
nand NAND2 (N4132, N4121, N994);
not NOT1 (N4133, N4106);
xor XOR2 (N4134, N4123, N283);
and AND2 (N4135, N4131, N2807);
xor XOR2 (N4136, N4134, N348);
not NOT1 (N4137, N4133);
nand NAND3 (N4138, N4136, N3581, N2034);
xor XOR2 (N4139, N4132, N4081);
buf BUF1 (N4140, N4127);
nand NAND4 (N4141, N4137, N3581, N2357, N748);
buf BUF1 (N4142, N4120);
buf BUF1 (N4143, N4140);
nor NOR3 (N4144, N4143, N426, N516);
xor XOR2 (N4145, N4144, N241);
buf BUF1 (N4146, N4128);
nor NOR3 (N4147, N4142, N2717, N3620);
nand NAND4 (N4148, N4138, N3010, N469, N434);
nand NAND3 (N4149, N4147, N390, N826);
nand NAND2 (N4150, N4135, N3915);
nor NOR2 (N4151, N4141, N1156);
nand NAND4 (N4152, N4149, N1473, N958, N552);
nand NAND3 (N4153, N4150, N3347, N928);
buf BUF1 (N4154, N4151);
nor NOR4 (N4155, N4152, N2996, N994, N1640);
nor NOR2 (N4156, N4129, N2459);
or OR4 (N4157, N4145, N1563, N3964, N406);
or OR4 (N4158, N4116, N961, N1427, N3018);
xor XOR2 (N4159, N4156, N877);
nand NAND3 (N4160, N4146, N1924, N71);
nand NAND4 (N4161, N4157, N3159, N3545, N2390);
and AND4 (N4162, N4158, N377, N3531, N1147);
nor NOR3 (N4163, N4162, N147, N1581);
nand NAND2 (N4164, N4161, N716);
buf BUF1 (N4165, N4164);
not NOT1 (N4166, N4165);
not NOT1 (N4167, N4139);
not NOT1 (N4168, N4159);
xor XOR2 (N4169, N4155, N3451);
buf BUF1 (N4170, N4154);
or OR4 (N4171, N4163, N2898, N1577, N2792);
nor NOR3 (N4172, N4119, N3285, N2543);
not NOT1 (N4173, N4171);
buf BUF1 (N4174, N4172);
nand NAND4 (N4175, N4148, N3679, N1117, N1782);
not NOT1 (N4176, N4173);
or OR2 (N4177, N4170, N3898);
not NOT1 (N4178, N4160);
xor XOR2 (N4179, N4169, N3223);
or OR2 (N4180, N4166, N687);
not NOT1 (N4181, N4176);
not NOT1 (N4182, N4179);
xor XOR2 (N4183, N4175, N3894);
nor NOR4 (N4184, N4174, N1316, N976, N2311);
nand NAND2 (N4185, N4182, N72);
and AND3 (N4186, N4181, N3459, N2147);
nand NAND2 (N4187, N4167, N681);
and AND2 (N4188, N4177, N878);
not NOT1 (N4189, N4184);
or OR4 (N4190, N4153, N101, N1329, N3183);
nor NOR4 (N4191, N4190, N2079, N637, N1738);
xor XOR2 (N4192, N4168, N2228);
not NOT1 (N4193, N4191);
nor NOR3 (N4194, N4193, N3825, N1787);
and AND2 (N4195, N4194, N1625);
or OR3 (N4196, N4187, N3723, N3845);
buf BUF1 (N4197, N4192);
buf BUF1 (N4198, N4196);
and AND4 (N4199, N4189, N3330, N354, N475);
xor XOR2 (N4200, N4185, N649);
or OR2 (N4201, N4180, N213);
xor XOR2 (N4202, N4201, N1253);
or OR2 (N4203, N4195, N879);
nor NOR3 (N4204, N4197, N3201, N51);
nor NOR2 (N4205, N4178, N3922);
not NOT1 (N4206, N4200);
nor NOR4 (N4207, N4206, N2650, N1029, N4081);
not NOT1 (N4208, N4188);
nor NOR2 (N4209, N4199, N735);
buf BUF1 (N4210, N4202);
not NOT1 (N4211, N4183);
buf BUF1 (N4212, N4207);
nand NAND4 (N4213, N4212, N3737, N896, N2683);
buf BUF1 (N4214, N4211);
not NOT1 (N4215, N4205);
xor XOR2 (N4216, N4210, N244);
or OR3 (N4217, N4214, N3572, N1280);
or OR2 (N4218, N4204, N1166);
buf BUF1 (N4219, N4216);
buf BUF1 (N4220, N4215);
nand NAND2 (N4221, N4213, N4013);
or OR2 (N4222, N4208, N990);
nand NAND3 (N4223, N4219, N2564, N4001);
xor XOR2 (N4224, N4223, N1403);
and AND4 (N4225, N4186, N767, N4096, N2375);
xor XOR2 (N4226, N4198, N4128);
and AND4 (N4227, N4220, N1027, N195, N1093);
or OR4 (N4228, N4224, N371, N3349, N3484);
nor NOR4 (N4229, N4227, N3421, N3797, N1624);
nor NOR2 (N4230, N4225, N3907);
xor XOR2 (N4231, N4209, N2197);
or OR2 (N4232, N4222, N1921);
or OR4 (N4233, N4231, N4200, N3520, N1710);
xor XOR2 (N4234, N4217, N3342);
nand NAND3 (N4235, N4230, N2507, N1861);
or OR3 (N4236, N4229, N3553, N598);
nor NOR2 (N4237, N4226, N1554);
nand NAND4 (N4238, N4233, N3325, N1184, N4156);
not NOT1 (N4239, N4237);
not NOT1 (N4240, N4218);
nor NOR2 (N4241, N4236, N1180);
xor XOR2 (N4242, N4239, N1098);
nor NOR2 (N4243, N4228, N3429);
and AND3 (N4244, N4232, N1509, N2596);
or OR4 (N4245, N4234, N2718, N885, N2681);
xor XOR2 (N4246, N4242, N2314);
nand NAND2 (N4247, N4243, N51);
or OR4 (N4248, N4235, N949, N725, N3045);
not NOT1 (N4249, N4241);
not NOT1 (N4250, N4221);
nor NOR4 (N4251, N4246, N1560, N2318, N307);
or OR3 (N4252, N4249, N2375, N3170);
and AND2 (N4253, N4250, N1425);
nor NOR3 (N4254, N4247, N2117, N170);
nor NOR3 (N4255, N4245, N529, N2810);
not NOT1 (N4256, N4254);
not NOT1 (N4257, N4238);
buf BUF1 (N4258, N4240);
and AND3 (N4259, N4258, N3703, N1435);
buf BUF1 (N4260, N4252);
or OR2 (N4261, N4253, N2793);
or OR2 (N4262, N4251, N4126);
nor NOR3 (N4263, N4261, N3409, N3339);
not NOT1 (N4264, N4257);
nor NOR2 (N4265, N4256, N1840);
buf BUF1 (N4266, N4264);
nor NOR4 (N4267, N4266, N4171, N2971, N1774);
nor NOR2 (N4268, N4255, N2265);
not NOT1 (N4269, N4263);
or OR4 (N4270, N4269, N482, N2466, N404);
nand NAND3 (N4271, N4244, N975, N2690);
buf BUF1 (N4272, N4270);
not NOT1 (N4273, N4265);
buf BUF1 (N4274, N4273);
nor NOR4 (N4275, N4267, N1732, N1537, N2130);
nand NAND3 (N4276, N4274, N824, N318);
nand NAND4 (N4277, N4271, N334, N3971, N1429);
or OR2 (N4278, N4277, N2120);
xor XOR2 (N4279, N4248, N553);
and AND4 (N4280, N4262, N1474, N359, N582);
and AND3 (N4281, N4278, N1551, N2796);
and AND2 (N4282, N4259, N1914);
nor NOR4 (N4283, N4279, N2475, N334, N669);
buf BUF1 (N4284, N4280);
xor XOR2 (N4285, N4283, N360);
nand NAND2 (N4286, N4281, N506);
nor NOR4 (N4287, N4285, N3483, N1306, N774);
nand NAND4 (N4288, N4275, N982, N738, N2937);
buf BUF1 (N4289, N4272);
nor NOR4 (N4290, N4286, N2905, N1346, N4117);
buf BUF1 (N4291, N4289);
nor NOR3 (N4292, N4260, N2424, N1707);
or OR4 (N4293, N4287, N4170, N3026, N1788);
xor XOR2 (N4294, N4291, N456);
buf BUF1 (N4295, N4276);
xor XOR2 (N4296, N4203, N1329);
buf BUF1 (N4297, N4284);
buf BUF1 (N4298, N4296);
buf BUF1 (N4299, N4292);
buf BUF1 (N4300, N4295);
xor XOR2 (N4301, N4294, N3683);
xor XOR2 (N4302, N4301, N311);
and AND4 (N4303, N4302, N1155, N3598, N1506);
and AND3 (N4304, N4282, N340, N2875);
buf BUF1 (N4305, N4297);
xor XOR2 (N4306, N4305, N460);
or OR2 (N4307, N4268, N4075);
or OR4 (N4308, N4299, N1559, N2384, N3780);
nor NOR3 (N4309, N4304, N2903, N1466);
and AND3 (N4310, N4288, N2397, N1856);
not NOT1 (N4311, N4290);
and AND2 (N4312, N4307, N1131);
xor XOR2 (N4313, N4298, N4177);
xor XOR2 (N4314, N4311, N2671);
buf BUF1 (N4315, N4303);
and AND3 (N4316, N4313, N3066, N1134);
nand NAND3 (N4317, N4300, N2582, N1963);
buf BUF1 (N4318, N4306);
xor XOR2 (N4319, N4309, N1718);
nor NOR3 (N4320, N4308, N1255, N3312);
or OR3 (N4321, N4312, N736, N2277);
nand NAND4 (N4322, N4319, N771, N4242, N587);
and AND4 (N4323, N4315, N4038, N1218, N465);
nand NAND2 (N4324, N4321, N2823);
xor XOR2 (N4325, N4324, N666);
nor NOR2 (N4326, N4325, N3735);
xor XOR2 (N4327, N4326, N22);
nand NAND3 (N4328, N4327, N1640, N2014);
not NOT1 (N4329, N4310);
or OR3 (N4330, N4328, N1310, N2400);
or OR3 (N4331, N4317, N3211, N3768);
xor XOR2 (N4332, N4320, N957);
not NOT1 (N4333, N4331);
and AND2 (N4334, N4314, N877);
nand NAND3 (N4335, N4332, N1044, N3663);
and AND3 (N4336, N4329, N1614, N773);
and AND2 (N4337, N4330, N735);
or OR4 (N4338, N4322, N749, N3593, N1533);
or OR4 (N4339, N4323, N2470, N456, N2610);
nor NOR2 (N4340, N4334, N2361);
not NOT1 (N4341, N4335);
buf BUF1 (N4342, N4338);
nor NOR3 (N4343, N4341, N3626, N46);
buf BUF1 (N4344, N4342);
nor NOR4 (N4345, N4316, N997, N2847, N3824);
buf BUF1 (N4346, N4345);
xor XOR2 (N4347, N4346, N1850);
not NOT1 (N4348, N4343);
nand NAND2 (N4349, N4337, N743);
buf BUF1 (N4350, N4339);
and AND3 (N4351, N4336, N3278, N3733);
not NOT1 (N4352, N4350);
nand NAND2 (N4353, N4340, N2864);
nand NAND3 (N4354, N4348, N4018, N84);
or OR3 (N4355, N4354, N765, N615);
and AND3 (N4356, N4349, N190, N4145);
or OR4 (N4357, N4347, N3820, N2530, N3444);
or OR2 (N4358, N4352, N2764);
xor XOR2 (N4359, N4344, N2822);
not NOT1 (N4360, N4357);
buf BUF1 (N4361, N4351);
nor NOR4 (N4362, N4356, N3999, N1286, N1006);
buf BUF1 (N4363, N4362);
xor XOR2 (N4364, N4333, N939);
nor NOR4 (N4365, N4355, N994, N1031, N1902);
buf BUF1 (N4366, N4361);
nor NOR3 (N4367, N4358, N336, N1932);
and AND4 (N4368, N4359, N4320, N1553, N2247);
buf BUF1 (N4369, N4367);
buf BUF1 (N4370, N4365);
buf BUF1 (N4371, N4366);
or OR3 (N4372, N4363, N2128, N407);
or OR2 (N4373, N4372, N1901);
not NOT1 (N4374, N4353);
and AND2 (N4375, N4374, N4162);
nand NAND2 (N4376, N4370, N2819);
not NOT1 (N4377, N4371);
not NOT1 (N4378, N4369);
xor XOR2 (N4379, N4377, N2924);
not NOT1 (N4380, N4375);
nor NOR2 (N4381, N4360, N3445);
or OR3 (N4382, N4368, N2925, N2263);
xor XOR2 (N4383, N4293, N2240);
and AND3 (N4384, N4373, N255, N2061);
nor NOR3 (N4385, N4382, N1179, N136);
not NOT1 (N4386, N4384);
nand NAND2 (N4387, N4379, N3127);
not NOT1 (N4388, N4378);
buf BUF1 (N4389, N4386);
xor XOR2 (N4390, N4385, N732);
nor NOR4 (N4391, N4381, N1851, N535, N290);
xor XOR2 (N4392, N4387, N2998);
or OR4 (N4393, N4380, N378, N3309, N3633);
buf BUF1 (N4394, N4392);
nor NOR4 (N4395, N4389, N1087, N3048, N2823);
buf BUF1 (N4396, N4376);
or OR4 (N4397, N4388, N2812, N1776, N2799);
xor XOR2 (N4398, N4383, N3913);
buf BUF1 (N4399, N4391);
nand NAND4 (N4400, N4318, N3225, N1527, N1608);
and AND2 (N4401, N4397, N3849);
nand NAND3 (N4402, N4390, N1014, N2307);
xor XOR2 (N4403, N4399, N549);
nand NAND3 (N4404, N4398, N1771, N379);
nand NAND2 (N4405, N4404, N3894);
nand NAND3 (N4406, N4402, N3296, N2981);
xor XOR2 (N4407, N4401, N3809);
xor XOR2 (N4408, N4405, N2986);
xor XOR2 (N4409, N4395, N2828);
not NOT1 (N4410, N4403);
not NOT1 (N4411, N4394);
or OR4 (N4412, N4408, N4252, N1965, N3017);
nand NAND4 (N4413, N4412, N948, N50, N4223);
nor NOR3 (N4414, N4410, N3147, N3965);
not NOT1 (N4415, N4414);
nor NOR3 (N4416, N4364, N3642, N2584);
xor XOR2 (N4417, N4396, N1144);
or OR4 (N4418, N4409, N1267, N3908, N3592);
nand NAND3 (N4419, N4418, N709, N2228);
and AND2 (N4420, N4407, N324);
or OR4 (N4421, N4420, N1385, N1473, N3914);
nand NAND3 (N4422, N4413, N3657, N2850);
nor NOR4 (N4423, N4416, N1886, N977, N3266);
xor XOR2 (N4424, N4411, N3733);
or OR4 (N4425, N4419, N366, N3848, N2648);
or OR4 (N4426, N4415, N4199, N4097, N725);
buf BUF1 (N4427, N4423);
and AND4 (N4428, N4406, N376, N2398, N77);
buf BUF1 (N4429, N4426);
nand NAND4 (N4430, N4417, N2344, N2540, N2805);
buf BUF1 (N4431, N4427);
xor XOR2 (N4432, N4430, N2641);
buf BUF1 (N4433, N4400);
xor XOR2 (N4434, N4428, N443);
or OR3 (N4435, N4434, N3258, N585);
buf BUF1 (N4436, N4421);
not NOT1 (N4437, N4436);
nand NAND4 (N4438, N4424, N1522, N1917, N2316);
buf BUF1 (N4439, N4437);
and AND3 (N4440, N4432, N3232, N3841);
buf BUF1 (N4441, N4431);
buf BUF1 (N4442, N4433);
nor NOR4 (N4443, N4440, N1276, N799, N3838);
xor XOR2 (N4444, N4443, N1709);
or OR4 (N4445, N4438, N2215, N1099, N3626);
not NOT1 (N4446, N4422);
or OR3 (N4447, N4439, N2437, N2223);
xor XOR2 (N4448, N4446, N29);
and AND2 (N4449, N4445, N636);
nand NAND3 (N4450, N4429, N1034, N2759);
nor NOR3 (N4451, N4435, N1048, N999);
and AND4 (N4452, N4444, N178, N4047, N1697);
xor XOR2 (N4453, N4425, N2373);
not NOT1 (N4454, N4451);
nor NOR2 (N4455, N4441, N119);
nand NAND3 (N4456, N4450, N1340, N1136);
buf BUF1 (N4457, N4448);
nor NOR3 (N4458, N4457, N6, N3186);
or OR4 (N4459, N4456, N2912, N4202, N4362);
nor NOR3 (N4460, N4442, N952, N12);
or OR4 (N4461, N4460, N2342, N662, N951);
nor NOR3 (N4462, N4461, N913, N3722);
nor NOR3 (N4463, N4459, N2283, N2916);
buf BUF1 (N4464, N4462);
nor NOR4 (N4465, N4447, N2988, N1309, N2108);
and AND4 (N4466, N4464, N3504, N1624, N3211);
buf BUF1 (N4467, N4454);
buf BUF1 (N4468, N4455);
and AND3 (N4469, N4466, N4038, N4375);
buf BUF1 (N4470, N4452);
and AND4 (N4471, N4465, N1345, N2625, N412);
buf BUF1 (N4472, N4467);
nor NOR2 (N4473, N4472, N2364);
xor XOR2 (N4474, N4470, N594);
buf BUF1 (N4475, N4393);
or OR4 (N4476, N4475, N4015, N3835, N4128);
buf BUF1 (N4477, N4471);
nand NAND2 (N4478, N4473, N1581);
nand NAND3 (N4479, N4477, N1991, N263);
not NOT1 (N4480, N4449);
nor NOR2 (N4481, N4453, N3337);
nor NOR2 (N4482, N4474, N660);
not NOT1 (N4483, N4481);
or OR4 (N4484, N4476, N1196, N195, N213);
nor NOR2 (N4485, N4484, N4098);
not NOT1 (N4486, N4468);
xor XOR2 (N4487, N4483, N208);
or OR4 (N4488, N4478, N1906, N430, N4228);
and AND3 (N4489, N4485, N2472, N1979);
nor NOR2 (N4490, N4479, N3300);
nor NOR4 (N4491, N4469, N1179, N4103, N553);
not NOT1 (N4492, N4488);
buf BUF1 (N4493, N4480);
not NOT1 (N4494, N4482);
or OR4 (N4495, N4494, N3089, N4205, N2557);
or OR3 (N4496, N4486, N3993, N4169);
or OR3 (N4497, N4489, N1920, N1697);
and AND3 (N4498, N4492, N4160, N2250);
or OR3 (N4499, N4496, N1625, N2601);
or OR3 (N4500, N4497, N941, N638);
nand NAND4 (N4501, N4500, N416, N1879, N739);
nor NOR2 (N4502, N4487, N537);
buf BUF1 (N4503, N4463);
or OR4 (N4504, N4495, N2897, N692, N2770);
or OR4 (N4505, N4504, N1385, N3081, N3913);
nor NOR2 (N4506, N4503, N2747);
xor XOR2 (N4507, N4491, N1044);
not NOT1 (N4508, N4490);
and AND4 (N4509, N4499, N4201, N305, N22);
not NOT1 (N4510, N4498);
nand NAND2 (N4511, N4505, N3800);
xor XOR2 (N4512, N4507, N1224);
buf BUF1 (N4513, N4511);
and AND3 (N4514, N4502, N857, N844);
xor XOR2 (N4515, N4513, N3249);
not NOT1 (N4516, N4501);
not NOT1 (N4517, N4510);
or OR2 (N4518, N4458, N944);
buf BUF1 (N4519, N4516);
or OR2 (N4520, N4514, N1464);
nand NAND2 (N4521, N4517, N685);
nor NOR2 (N4522, N4520, N1333);
not NOT1 (N4523, N4512);
or OR3 (N4524, N4493, N3218, N2849);
xor XOR2 (N4525, N4508, N652);
nand NAND4 (N4526, N4519, N2191, N1320, N2490);
nor NOR2 (N4527, N4526, N2507);
and AND2 (N4528, N4525, N2849);
not NOT1 (N4529, N4515);
nor NOR4 (N4530, N4509, N3492, N3942, N1334);
xor XOR2 (N4531, N4527, N4432);
buf BUF1 (N4532, N4521);
and AND3 (N4533, N4518, N3322, N3889);
buf BUF1 (N4534, N4528);
or OR3 (N4535, N4524, N3169, N2371);
xor XOR2 (N4536, N4523, N1398);
not NOT1 (N4537, N4522);
xor XOR2 (N4538, N4531, N2964);
nand NAND2 (N4539, N4532, N2739);
nand NAND3 (N4540, N4530, N3362, N3419);
and AND4 (N4541, N4536, N1143, N992, N4160);
not NOT1 (N4542, N4533);
xor XOR2 (N4543, N4540, N4047);
nor NOR4 (N4544, N4541, N3460, N328, N3140);
nand NAND2 (N4545, N4538, N2230);
not NOT1 (N4546, N4539);
buf BUF1 (N4547, N4529);
not NOT1 (N4548, N4542);
nand NAND3 (N4549, N4547, N2406, N463);
not NOT1 (N4550, N4544);
or OR2 (N4551, N4537, N2999);
not NOT1 (N4552, N4551);
not NOT1 (N4553, N4550);
not NOT1 (N4554, N4546);
nand NAND4 (N4555, N4506, N4497, N1970, N2445);
not NOT1 (N4556, N4534);
nand NAND2 (N4557, N4553, N4121);
or OR3 (N4558, N4552, N3268, N4090);
buf BUF1 (N4559, N4557);
buf BUF1 (N4560, N4549);
buf BUF1 (N4561, N4548);
not NOT1 (N4562, N4555);
nand NAND4 (N4563, N4543, N2633, N716, N1650);
buf BUF1 (N4564, N4560);
and AND2 (N4565, N4559, N4508);
and AND3 (N4566, N4561, N746, N213);
xor XOR2 (N4567, N4563, N2100);
nand NAND4 (N4568, N4565, N1162, N4294, N161);
not NOT1 (N4569, N4564);
xor XOR2 (N4570, N4545, N427);
not NOT1 (N4571, N4570);
not NOT1 (N4572, N4554);
not NOT1 (N4573, N4572);
nor NOR2 (N4574, N4562, N2117);
xor XOR2 (N4575, N4556, N4077);
nor NOR4 (N4576, N4558, N2980, N2877, N2359);
and AND2 (N4577, N4566, N800);
xor XOR2 (N4578, N4535, N20);
xor XOR2 (N4579, N4567, N4104);
xor XOR2 (N4580, N4579, N3507);
and AND3 (N4581, N4574, N2710, N1669);
and AND3 (N4582, N4577, N1545, N1776);
not NOT1 (N4583, N4568);
xor XOR2 (N4584, N4580, N3031);
nor NOR2 (N4585, N4571, N2033);
nor NOR4 (N4586, N4578, N583, N3542, N1029);
buf BUF1 (N4587, N4575);
not NOT1 (N4588, N4583);
xor XOR2 (N4589, N4576, N4212);
xor XOR2 (N4590, N4589, N2723);
or OR2 (N4591, N4590, N2173);
buf BUF1 (N4592, N4584);
not NOT1 (N4593, N4587);
or OR4 (N4594, N4593, N1027, N3043, N4198);
nand NAND3 (N4595, N4573, N4509, N2500);
xor XOR2 (N4596, N4582, N2254);
and AND2 (N4597, N4591, N1620);
not NOT1 (N4598, N4569);
nand NAND3 (N4599, N4581, N860, N21);
nor NOR2 (N4600, N4597, N1292);
nor NOR4 (N4601, N4594, N2891, N2959, N1630);
not NOT1 (N4602, N4596);
or OR2 (N4603, N4592, N998);
nor NOR3 (N4604, N4595, N3967, N2049);
buf BUF1 (N4605, N4586);
xor XOR2 (N4606, N4598, N2541);
xor XOR2 (N4607, N4588, N65);
nor NOR3 (N4608, N4601, N115, N1986);
and AND4 (N4609, N4608, N1223, N1218, N1952);
and AND4 (N4610, N4600, N3913, N4170, N1537);
buf BUF1 (N4611, N4606);
nor NOR4 (N4612, N4599, N2561, N487, N138);
and AND2 (N4613, N4603, N4232);
not NOT1 (N4614, N4605);
xor XOR2 (N4615, N4609, N2129);
or OR2 (N4616, N4613, N3672);
and AND2 (N4617, N4615, N3096);
and AND2 (N4618, N4585, N3736);
nand NAND4 (N4619, N4610, N1000, N2471, N790);
or OR3 (N4620, N4611, N1584, N2384);
xor XOR2 (N4621, N4619, N3046);
not NOT1 (N4622, N4612);
nor NOR2 (N4623, N4604, N2358);
and AND3 (N4624, N4607, N228, N241);
buf BUF1 (N4625, N4623);
nor NOR2 (N4626, N4622, N3960);
nor NOR2 (N4627, N4617, N1862);
nor NOR2 (N4628, N4616, N104);
or OR2 (N4629, N4624, N1161);
not NOT1 (N4630, N4620);
xor XOR2 (N4631, N4630, N59);
nor NOR4 (N4632, N4614, N3255, N1784, N1322);
not NOT1 (N4633, N4625);
or OR3 (N4634, N4628, N4116, N2663);
nand NAND2 (N4635, N4627, N629);
not NOT1 (N4636, N4626);
and AND4 (N4637, N4618, N557, N172, N1140);
xor XOR2 (N4638, N4633, N1316);
or OR3 (N4639, N4635, N913, N1834);
xor XOR2 (N4640, N4631, N899);
nand NAND2 (N4641, N4640, N4281);
not NOT1 (N4642, N4621);
nor NOR2 (N4643, N4637, N1316);
not NOT1 (N4644, N4641);
nand NAND4 (N4645, N4638, N3622, N2822, N37);
nor NOR2 (N4646, N4634, N2348);
nand NAND4 (N4647, N4629, N313, N204, N569);
nand NAND4 (N4648, N4639, N4103, N1741, N2673);
nor NOR2 (N4649, N4647, N3085);
or OR3 (N4650, N4632, N2985, N1657);
buf BUF1 (N4651, N4644);
buf BUF1 (N4652, N4602);
and AND2 (N4653, N4651, N73);
nor NOR3 (N4654, N4636, N2091, N3695);
buf BUF1 (N4655, N4649);
nor NOR4 (N4656, N4655, N2807, N3626, N1316);
nor NOR2 (N4657, N4654, N672);
and AND3 (N4658, N4642, N981, N3107);
and AND4 (N4659, N4645, N1759, N2747, N2916);
not NOT1 (N4660, N4646);
and AND3 (N4661, N4653, N1787, N371);
or OR3 (N4662, N4660, N1287, N2198);
and AND3 (N4663, N4661, N3508, N1215);
buf BUF1 (N4664, N4659);
nor NOR2 (N4665, N4663, N1520);
xor XOR2 (N4666, N4648, N802);
xor XOR2 (N4667, N4666, N4528);
or OR3 (N4668, N4664, N3466, N4067);
and AND2 (N4669, N4665, N823);
and AND2 (N4670, N4662, N717);
nor NOR4 (N4671, N4643, N2958, N2309, N1854);
nor NOR3 (N4672, N4656, N2190, N2139);
nor NOR2 (N4673, N4652, N3269);
nand NAND2 (N4674, N4657, N4228);
and AND4 (N4675, N4670, N428, N3627, N3439);
nor NOR3 (N4676, N4672, N2417, N4190);
buf BUF1 (N4677, N4650);
buf BUF1 (N4678, N4677);
nand NAND4 (N4679, N4669, N4543, N4365, N976);
nand NAND2 (N4680, N4673, N3068);
and AND3 (N4681, N4675, N568, N1542);
nand NAND2 (N4682, N4668, N728);
not NOT1 (N4683, N4676);
nor NOR3 (N4684, N4671, N3259, N3042);
xor XOR2 (N4685, N4680, N4276);
nor NOR4 (N4686, N4685, N2636, N2663, N2113);
xor XOR2 (N4687, N4674, N3546);
nand NAND4 (N4688, N4687, N3839, N2247, N320);
or OR2 (N4689, N4686, N4287);
xor XOR2 (N4690, N4684, N3326);
buf BUF1 (N4691, N4688);
nor NOR4 (N4692, N4667, N1285, N725, N3711);
and AND3 (N4693, N4658, N1281, N3003);
not NOT1 (N4694, N4693);
and AND4 (N4695, N4691, N1578, N3572, N1190);
xor XOR2 (N4696, N4682, N405);
xor XOR2 (N4697, N4683, N2859);
xor XOR2 (N4698, N4697, N2394);
not NOT1 (N4699, N4689);
and AND2 (N4700, N4679, N4638);
xor XOR2 (N4701, N4690, N42);
nor NOR4 (N4702, N4698, N3692, N923, N4380);
buf BUF1 (N4703, N4702);
and AND4 (N4704, N4678, N4230, N77, N1419);
nor NOR3 (N4705, N4699, N4214, N1788);
and AND3 (N4706, N4695, N4689, N680);
nand NAND4 (N4707, N4704, N1635, N3740, N4126);
nand NAND2 (N4708, N4692, N2325);
nand NAND3 (N4709, N4703, N3021, N370);
buf BUF1 (N4710, N4696);
buf BUF1 (N4711, N4681);
nand NAND2 (N4712, N4707, N3426);
or OR2 (N4713, N4706, N2424);
nand NAND4 (N4714, N4700, N902, N2233, N3839);
or OR4 (N4715, N4701, N2581, N3474, N681);
xor XOR2 (N4716, N4710, N4633);
or OR4 (N4717, N4708, N3655, N3323, N1406);
buf BUF1 (N4718, N4714);
xor XOR2 (N4719, N4717, N2493);
and AND2 (N4720, N4709, N4633);
nand NAND2 (N4721, N4719, N4509);
not NOT1 (N4722, N4694);
or OR2 (N4723, N4705, N506);
and AND3 (N4724, N4720, N2516, N4378);
xor XOR2 (N4725, N4721, N588);
xor XOR2 (N4726, N4718, N3149);
or OR3 (N4727, N4726, N3644, N973);
nor NOR4 (N4728, N4722, N3644, N4311, N4084);
not NOT1 (N4729, N4728);
buf BUF1 (N4730, N4724);
not NOT1 (N4731, N4713);
not NOT1 (N4732, N4729);
or OR3 (N4733, N4711, N2089, N3251);
nor NOR3 (N4734, N4727, N432, N2040);
nor NOR3 (N4735, N4715, N3484, N2966);
or OR3 (N4736, N4716, N3617, N349);
not NOT1 (N4737, N4732);
or OR2 (N4738, N4723, N4325);
not NOT1 (N4739, N4738);
nor NOR2 (N4740, N4712, N1647);
xor XOR2 (N4741, N4735, N2629);
nand NAND4 (N4742, N4733, N3894, N3369, N1490);
nor NOR4 (N4743, N4741, N1661, N2678, N1862);
or OR2 (N4744, N4737, N4400);
xor XOR2 (N4745, N4736, N2990);
nand NAND2 (N4746, N4740, N3889);
nand NAND4 (N4747, N4743, N2806, N2574, N679);
nand NAND2 (N4748, N4744, N1640);
not NOT1 (N4749, N4746);
not NOT1 (N4750, N4739);
and AND4 (N4751, N4730, N3380, N3695, N1207);
and AND3 (N4752, N4734, N828, N3172);
not NOT1 (N4753, N4749);
not NOT1 (N4754, N4748);
nor NOR4 (N4755, N4725, N2504, N3244, N799);
nor NOR2 (N4756, N4755, N678);
xor XOR2 (N4757, N4742, N2202);
buf BUF1 (N4758, N4745);
or OR3 (N4759, N4757, N1520, N2840);
buf BUF1 (N4760, N4753);
not NOT1 (N4761, N4758);
xor XOR2 (N4762, N4747, N154);
or OR4 (N4763, N4750, N790, N1289, N3342);
or OR4 (N4764, N4752, N150, N3513, N1810);
and AND3 (N4765, N4764, N3602, N3504);
or OR2 (N4766, N4760, N4123);
nand NAND2 (N4767, N4756, N2772);
nor NOR2 (N4768, N4765, N4484);
or OR2 (N4769, N4768, N4331);
and AND2 (N4770, N4763, N907);
buf BUF1 (N4771, N4751);
nor NOR2 (N4772, N4769, N3753);
nand NAND3 (N4773, N4770, N4483, N2904);
buf BUF1 (N4774, N4767);
nor NOR2 (N4775, N4762, N3829);
or OR3 (N4776, N4731, N1093, N733);
or OR3 (N4777, N4754, N4240, N3482);
not NOT1 (N4778, N4771);
nand NAND3 (N4779, N4766, N44, N959);
buf BUF1 (N4780, N4761);
and AND3 (N4781, N4776, N172, N3383);
xor XOR2 (N4782, N4772, N4437);
nand NAND3 (N4783, N4759, N511, N2270);
buf BUF1 (N4784, N4778);
nor NOR3 (N4785, N4777, N4777, N4393);
xor XOR2 (N4786, N4779, N1851);
buf BUF1 (N4787, N4784);
and AND2 (N4788, N4773, N3862);
or OR2 (N4789, N4780, N3314);
xor XOR2 (N4790, N4788, N830);
or OR4 (N4791, N4790, N1711, N1113, N4220);
xor XOR2 (N4792, N4781, N4731);
xor XOR2 (N4793, N4775, N4716);
not NOT1 (N4794, N4793);
and AND3 (N4795, N4785, N2097, N4501);
nor NOR3 (N4796, N4794, N4211, N1774);
not NOT1 (N4797, N4774);
and AND3 (N4798, N4792, N1058, N1858);
and AND2 (N4799, N4789, N2590);
nor NOR4 (N4800, N4795, N2231, N1894, N2428);
xor XOR2 (N4801, N4791, N3585);
xor XOR2 (N4802, N4787, N614);
xor XOR2 (N4803, N4799, N3664);
xor XOR2 (N4804, N4786, N801);
and AND3 (N4805, N4804, N2754, N2520);
or OR4 (N4806, N4798, N2392, N4805, N24);
or OR4 (N4807, N4338, N4078, N100, N1978);
and AND3 (N4808, N4800, N1392, N4467);
nand NAND4 (N4809, N4807, N485, N4378, N4193);
xor XOR2 (N4810, N4783, N3685);
nor NOR4 (N4811, N4808, N3197, N206, N4310);
not NOT1 (N4812, N4782);
nor NOR3 (N4813, N4806, N971, N2973);
and AND2 (N4814, N4809, N932);
or OR3 (N4815, N4813, N3191, N3516);
not NOT1 (N4816, N4812);
nor NOR3 (N4817, N4803, N1970, N3732);
nand NAND4 (N4818, N4801, N2196, N2950, N3305);
buf BUF1 (N4819, N4810);
nor NOR4 (N4820, N4818, N4572, N1595, N3380);
buf BUF1 (N4821, N4815);
xor XOR2 (N4822, N4811, N2913);
or OR2 (N4823, N4821, N291);
or OR4 (N4824, N4814, N3969, N4353, N1007);
or OR4 (N4825, N4823, N24, N1472, N2107);
not NOT1 (N4826, N4820);
not NOT1 (N4827, N4819);
nand NAND3 (N4828, N4827, N3096, N1661);
buf BUF1 (N4829, N4797);
or OR3 (N4830, N4817, N4598, N1533);
or OR3 (N4831, N4802, N4133, N3043);
nor NOR4 (N4832, N4826, N2745, N764, N2930);
and AND2 (N4833, N4830, N1957);
nand NAND2 (N4834, N4828, N3848);
nor NOR4 (N4835, N4831, N1807, N1244, N3666);
or OR2 (N4836, N4834, N4455);
and AND2 (N4837, N4832, N166);
nand NAND2 (N4838, N4837, N3236);
nor NOR4 (N4839, N4835, N4112, N3722, N4072);
xor XOR2 (N4840, N4796, N1197);
nor NOR3 (N4841, N4838, N429, N4594);
buf BUF1 (N4842, N4825);
not NOT1 (N4843, N4829);
buf BUF1 (N4844, N4836);
or OR4 (N4845, N4844, N3939, N135, N1476);
nor NOR2 (N4846, N4824, N1558);
nor NOR3 (N4847, N4816, N4084, N1854);
xor XOR2 (N4848, N4842, N1419);
nand NAND3 (N4849, N4847, N4227, N3948);
buf BUF1 (N4850, N4841);
xor XOR2 (N4851, N4822, N34);
or OR2 (N4852, N4849, N2173);
not NOT1 (N4853, N4833);
not NOT1 (N4854, N4843);
or OR2 (N4855, N4848, N1039);
or OR4 (N4856, N4854, N1142, N641, N1173);
and AND4 (N4857, N4855, N3930, N1300, N1947);
and AND4 (N4858, N4853, N2435, N4790, N2337);
buf BUF1 (N4859, N4851);
and AND3 (N4860, N4858, N1013, N1467);
or OR2 (N4861, N4850, N4154);
or OR3 (N4862, N4840, N4595, N3607);
nor NOR4 (N4863, N4852, N2118, N1586, N1120);
and AND2 (N4864, N4862, N1035);
buf BUF1 (N4865, N4859);
nor NOR4 (N4866, N4861, N3864, N2802, N4828);
xor XOR2 (N4867, N4863, N642);
and AND3 (N4868, N4846, N4634, N2472);
or OR2 (N4869, N4839, N3131);
nand NAND4 (N4870, N4845, N475, N2407, N2667);
or OR4 (N4871, N4866, N1054, N3269, N452);
or OR4 (N4872, N4867, N19, N2990, N2154);
nor NOR4 (N4873, N4860, N2952, N987, N490);
buf BUF1 (N4874, N4864);
or OR2 (N4875, N4872, N2510);
not NOT1 (N4876, N4857);
buf BUF1 (N4877, N4869);
and AND3 (N4878, N4865, N4668, N3595);
xor XOR2 (N4879, N4868, N2560);
nor NOR3 (N4880, N4874, N1121, N1154);
buf BUF1 (N4881, N4856);
buf BUF1 (N4882, N4873);
not NOT1 (N4883, N4880);
nor NOR2 (N4884, N4870, N193);
nor NOR4 (N4885, N4871, N2929, N840, N1247);
not NOT1 (N4886, N4878);
nor NOR3 (N4887, N4881, N2, N3471);
or OR2 (N4888, N4875, N1949);
nor NOR4 (N4889, N4887, N3977, N4351, N948);
buf BUF1 (N4890, N4888);
xor XOR2 (N4891, N4886, N2787);
nand NAND3 (N4892, N4891, N2375, N2111);
xor XOR2 (N4893, N4884, N4222);
nor NOR4 (N4894, N4893, N2434, N2578, N3618);
or OR3 (N4895, N4885, N1997, N4760);
nor NOR2 (N4896, N4879, N3025);
not NOT1 (N4897, N4877);
buf BUF1 (N4898, N4896);
and AND3 (N4899, N4883, N3951, N855);
or OR4 (N4900, N4897, N2772, N2678, N4544);
buf BUF1 (N4901, N4882);
or OR3 (N4902, N4889, N4617, N563);
xor XOR2 (N4903, N4902, N4863);
not NOT1 (N4904, N4901);
or OR2 (N4905, N4894, N1349);
not NOT1 (N4906, N4892);
or OR3 (N4907, N4899, N22, N2936);
buf BUF1 (N4908, N4907);
not NOT1 (N4909, N4895);
not NOT1 (N4910, N4904);
buf BUF1 (N4911, N4906);
not NOT1 (N4912, N4890);
xor XOR2 (N4913, N4912, N2091);
nor NOR3 (N4914, N4908, N3847, N2743);
nand NAND2 (N4915, N4876, N256);
not NOT1 (N4916, N4903);
xor XOR2 (N4917, N4916, N2230);
and AND2 (N4918, N4898, N4382);
not NOT1 (N4919, N4918);
or OR2 (N4920, N4915, N4152);
or OR2 (N4921, N4911, N3337);
xor XOR2 (N4922, N4900, N4501);
nor NOR4 (N4923, N4917, N4010, N4655, N4066);
buf BUF1 (N4924, N4921);
or OR2 (N4925, N4922, N940);
buf BUF1 (N4926, N4919);
xor XOR2 (N4927, N4923, N2091);
xor XOR2 (N4928, N4910, N3748);
or OR3 (N4929, N4905, N3809, N947);
and AND2 (N4930, N4927, N4401);
nor NOR4 (N4931, N4926, N4048, N3681, N3899);
xor XOR2 (N4932, N4929, N970);
or OR4 (N4933, N4914, N3451, N1616, N1868);
nand NAND2 (N4934, N4930, N1157);
buf BUF1 (N4935, N4909);
not NOT1 (N4936, N4933);
buf BUF1 (N4937, N4928);
or OR2 (N4938, N4931, N2219);
nand NAND2 (N4939, N4937, N4815);
buf BUF1 (N4940, N4936);
buf BUF1 (N4941, N4925);
or OR4 (N4942, N4940, N588, N1935, N534);
nand NAND3 (N4943, N4934, N4440, N2593);
not NOT1 (N4944, N4935);
and AND4 (N4945, N4920, N601, N906, N1223);
buf BUF1 (N4946, N4943);
xor XOR2 (N4947, N4938, N2476);
not NOT1 (N4948, N4932);
or OR2 (N4949, N4944, N2039);
nor NOR4 (N4950, N4942, N1788, N394, N4112);
xor XOR2 (N4951, N4941, N1075);
not NOT1 (N4952, N4951);
nor NOR2 (N4953, N4924, N2374);
xor XOR2 (N4954, N4945, N1610);
or OR4 (N4955, N4913, N1974, N3707, N1291);
nor NOR4 (N4956, N4947, N1477, N4532, N1314);
nand NAND4 (N4957, N4954, N3720, N4937, N1873);
and AND4 (N4958, N4955, N2476, N1424, N1340);
xor XOR2 (N4959, N4949, N1013);
xor XOR2 (N4960, N4950, N4055);
or OR4 (N4961, N4957, N2059, N2001, N765);
buf BUF1 (N4962, N4958);
xor XOR2 (N4963, N4956, N306);
buf BUF1 (N4964, N4963);
and AND2 (N4965, N4948, N4881);
and AND4 (N4966, N4959, N3215, N2493, N4696);
not NOT1 (N4967, N4952);
and AND3 (N4968, N4962, N2798, N2094);
nor NOR4 (N4969, N4966, N117, N328, N2340);
nand NAND2 (N4970, N4965, N282);
and AND4 (N4971, N4953, N3307, N1364, N2671);
not NOT1 (N4972, N4939);
not NOT1 (N4973, N4967);
xor XOR2 (N4974, N4946, N2256);
nor NOR3 (N4975, N4973, N3460, N4079);
nand NAND3 (N4976, N4971, N3489, N169);
nand NAND4 (N4977, N4961, N173, N482, N3166);
xor XOR2 (N4978, N4977, N3367);
nor NOR3 (N4979, N4968, N1752, N1761);
nor NOR2 (N4980, N4976, N4562);
nor NOR2 (N4981, N4975, N1299);
not NOT1 (N4982, N4970);
not NOT1 (N4983, N4980);
nor NOR3 (N4984, N4960, N490, N1839);
xor XOR2 (N4985, N4972, N4392);
or OR3 (N4986, N4969, N3709, N4767);
and AND3 (N4987, N4986, N1360, N4812);
and AND4 (N4988, N4964, N3290, N3207, N318);
and AND2 (N4989, N4983, N2043);
nand NAND4 (N4990, N4981, N4339, N2130, N2603);
xor XOR2 (N4991, N4990, N4033);
and AND3 (N4992, N4982, N4559, N3861);
nand NAND2 (N4993, N4984, N2569);
buf BUF1 (N4994, N4993);
xor XOR2 (N4995, N4989, N1412);
xor XOR2 (N4996, N4979, N2310);
nand NAND3 (N4997, N4991, N395, N3479);
nor NOR2 (N4998, N4997, N713);
not NOT1 (N4999, N4995);
buf BUF1 (N5000, N4988);
nand NAND3 (N5001, N4978, N2453, N3777);
xor XOR2 (N5002, N4974, N3756);
buf BUF1 (N5003, N4992);
buf BUF1 (N5004, N4987);
xor XOR2 (N5005, N5003, N406);
and AND3 (N5006, N5001, N1042, N849);
xor XOR2 (N5007, N4985, N64);
and AND4 (N5008, N5005, N1908, N3185, N4786);
nor NOR2 (N5009, N4994, N1883);
nor NOR3 (N5010, N4998, N2069, N565);
nand NAND2 (N5011, N5009, N4221);
buf BUF1 (N5012, N5008);
nand NAND3 (N5013, N5002, N4375, N399);
or OR4 (N5014, N4996, N707, N796, N3510);
nand NAND4 (N5015, N5006, N2799, N1799, N4451);
buf BUF1 (N5016, N4999);
and AND3 (N5017, N5015, N4948, N846);
not NOT1 (N5018, N5013);
not NOT1 (N5019, N5012);
or OR4 (N5020, N5000, N3209, N784, N3038);
and AND4 (N5021, N5016, N1050, N1048, N1571);
and AND4 (N5022, N5018, N2470, N3245, N1021);
nand NAND2 (N5023, N5022, N4906);
or OR4 (N5024, N5004, N4638, N2789, N4973);
not NOT1 (N5025, N5023);
nand NAND3 (N5026, N5020, N1492, N3900);
xor XOR2 (N5027, N5026, N2844);
buf BUF1 (N5028, N5019);
nor NOR3 (N5029, N5028, N556, N4226);
not NOT1 (N5030, N5024);
nand NAND4 (N5031, N5011, N2446, N3663, N2002);
buf BUF1 (N5032, N5029);
and AND3 (N5033, N5025, N321, N2658);
buf BUF1 (N5034, N5033);
buf BUF1 (N5035, N5032);
nor NOR2 (N5036, N5034, N460);
or OR4 (N5037, N5027, N128, N1337, N634);
nand NAND4 (N5038, N5007, N3443, N4256, N2281);
not NOT1 (N5039, N5036);
and AND4 (N5040, N5037, N1153, N1813, N4205);
buf BUF1 (N5041, N5038);
buf BUF1 (N5042, N5039);
nand NAND4 (N5043, N5040, N671, N3662, N3902);
xor XOR2 (N5044, N5014, N343);
nor NOR2 (N5045, N5031, N3847);
or OR3 (N5046, N5035, N4006, N4586);
nand NAND2 (N5047, N5044, N2249);
buf BUF1 (N5048, N5041);
nand NAND4 (N5049, N5030, N1786, N3602, N2109);
buf BUF1 (N5050, N5046);
nor NOR4 (N5051, N5017, N2754, N191, N120);
buf BUF1 (N5052, N5042);
and AND2 (N5053, N5051, N2010);
xor XOR2 (N5054, N5043, N412);
nor NOR4 (N5055, N5048, N3486, N1975, N3214);
nor NOR2 (N5056, N5052, N2678);
or OR3 (N5057, N5053, N4029, N4344);
or OR4 (N5058, N5057, N2564, N544, N3622);
not NOT1 (N5059, N5047);
or OR3 (N5060, N5010, N2298, N3547);
or OR4 (N5061, N5049, N4845, N195, N484);
and AND2 (N5062, N5056, N2474);
buf BUF1 (N5063, N5045);
or OR3 (N5064, N5059, N4988, N4529);
nand NAND4 (N5065, N5061, N2060, N2785, N962);
buf BUF1 (N5066, N5054);
and AND4 (N5067, N5066, N1011, N3065, N4908);
buf BUF1 (N5068, N5050);
nand NAND2 (N5069, N5058, N959);
or OR4 (N5070, N5068, N2812, N3928, N304);
or OR2 (N5071, N5055, N3290);
or OR3 (N5072, N5067, N2828, N1196);
nand NAND4 (N5073, N5064, N49, N3501, N1368);
not NOT1 (N5074, N5070);
buf BUF1 (N5075, N5072);
nand NAND2 (N5076, N5065, N4809);
and AND2 (N5077, N5063, N4433);
or OR4 (N5078, N5077, N4995, N2344, N1409);
nand NAND4 (N5079, N5074, N2163, N1895, N4321);
xor XOR2 (N5080, N5079, N270);
xor XOR2 (N5081, N5078, N3808);
not NOT1 (N5082, N5060);
and AND3 (N5083, N5082, N1299, N4125);
nand NAND2 (N5084, N5062, N4562);
buf BUF1 (N5085, N5081);
nor NOR4 (N5086, N5084, N1783, N4, N3131);
or OR3 (N5087, N5021, N914, N3072);
nand NAND2 (N5088, N5085, N3898);
xor XOR2 (N5089, N5071, N2539);
and AND3 (N5090, N5083, N2224, N1013);
nor NOR4 (N5091, N5089, N1470, N1910, N618);
nand NAND3 (N5092, N5073, N4006, N2523);
not NOT1 (N5093, N5090);
xor XOR2 (N5094, N5080, N1852);
buf BUF1 (N5095, N5087);
buf BUF1 (N5096, N5093);
xor XOR2 (N5097, N5094, N5061);
xor XOR2 (N5098, N5092, N4780);
xor XOR2 (N5099, N5075, N2120);
or OR3 (N5100, N5076, N2101, N2998);
and AND4 (N5101, N5091, N4918, N1065, N4364);
buf BUF1 (N5102, N5088);
and AND3 (N5103, N5097, N4387, N4598);
and AND2 (N5104, N5098, N2574);
not NOT1 (N5105, N5103);
and AND3 (N5106, N5086, N1395, N2814);
not NOT1 (N5107, N5106);
nand NAND3 (N5108, N5102, N2038, N3144);
nor NOR3 (N5109, N5105, N2918, N4729);
nand NAND3 (N5110, N5104, N1780, N4263);
nand NAND3 (N5111, N5100, N2854, N4887);
nor NOR3 (N5112, N5096, N2887, N742);
nor NOR3 (N5113, N5101, N2258, N1156);
nor NOR4 (N5114, N5107, N1972, N361, N1874);
nor NOR4 (N5115, N5099, N1043, N2599, N4774);
nor NOR2 (N5116, N5111, N2679);
nand NAND3 (N5117, N5108, N2214, N3415);
or OR4 (N5118, N5110, N3969, N2043, N1888);
buf BUF1 (N5119, N5115);
not NOT1 (N5120, N5118);
buf BUF1 (N5121, N5117);
xor XOR2 (N5122, N5119, N1312);
xor XOR2 (N5123, N5121, N2486);
xor XOR2 (N5124, N5114, N2571);
nor NOR4 (N5125, N5124, N4455, N555, N2371);
and AND4 (N5126, N5112, N3183, N4817, N2405);
or OR4 (N5127, N5126, N2611, N2270, N2940);
xor XOR2 (N5128, N5125, N3247);
xor XOR2 (N5129, N5128, N3713);
nand NAND3 (N5130, N5113, N3166, N4830);
not NOT1 (N5131, N5127);
nand NAND2 (N5132, N5131, N3524);
and AND3 (N5133, N5123, N1988, N282);
nand NAND2 (N5134, N5095, N3642);
and AND3 (N5135, N5069, N2289, N175);
buf BUF1 (N5136, N5135);
buf BUF1 (N5137, N5120);
xor XOR2 (N5138, N5116, N1191);
or OR2 (N5139, N5136, N3034);
nand NAND3 (N5140, N5138, N2782, N4020);
or OR3 (N5141, N5134, N3976, N3604);
xor XOR2 (N5142, N5122, N3028);
nand NAND4 (N5143, N5129, N3999, N2359, N4462);
nor NOR3 (N5144, N5130, N2146, N3728);
nand NAND4 (N5145, N5133, N4077, N1282, N3396);
and AND4 (N5146, N5143, N2585, N1682, N911);
nor NOR4 (N5147, N5109, N714, N4956, N817);
or OR2 (N5148, N5142, N2590);
or OR2 (N5149, N5132, N4949);
not NOT1 (N5150, N5146);
nand NAND4 (N5151, N5148, N4389, N502, N3528);
buf BUF1 (N5152, N5145);
nor NOR2 (N5153, N5139, N1422);
or OR2 (N5154, N5151, N4506);
not NOT1 (N5155, N5150);
xor XOR2 (N5156, N5152, N3654);
xor XOR2 (N5157, N5140, N5097);
or OR2 (N5158, N5141, N893);
buf BUF1 (N5159, N5156);
nor NOR4 (N5160, N5144, N899, N1134, N1728);
xor XOR2 (N5161, N5157, N238);
nand NAND4 (N5162, N5160, N2874, N541, N1445);
nor NOR2 (N5163, N5159, N1325);
and AND2 (N5164, N5162, N4141);
xor XOR2 (N5165, N5164, N1555);
nor NOR4 (N5166, N5137, N334, N2860, N3402);
and AND4 (N5167, N5161, N2559, N1411, N169);
nand NAND4 (N5168, N5154, N930, N3370, N5055);
nand NAND2 (N5169, N5166, N2209);
or OR4 (N5170, N5158, N881, N5136, N1919);
buf BUF1 (N5171, N5168);
or OR2 (N5172, N5167, N3867);
or OR2 (N5173, N5155, N671);
and AND3 (N5174, N5147, N1186, N3178);
and AND3 (N5175, N5169, N4578, N2897);
or OR3 (N5176, N5149, N3927, N1602);
not NOT1 (N5177, N5163);
xor XOR2 (N5178, N5172, N3795);
and AND3 (N5179, N5171, N4151, N3813);
and AND4 (N5180, N5165, N2374, N4182, N1448);
or OR4 (N5181, N5179, N1997, N3315, N521);
buf BUF1 (N5182, N5177);
or OR4 (N5183, N5181, N966, N4772, N4844);
nand NAND2 (N5184, N5153, N290);
buf BUF1 (N5185, N5176);
and AND2 (N5186, N5184, N216);
not NOT1 (N5187, N5174);
and AND2 (N5188, N5178, N1341);
nor NOR4 (N5189, N5187, N4045, N4425, N2302);
or OR2 (N5190, N5175, N2891);
nor NOR2 (N5191, N5185, N3297);
and AND3 (N5192, N5170, N1131, N808);
nand NAND4 (N5193, N5173, N588, N3523, N2123);
or OR4 (N5194, N5193, N3570, N4370, N3616);
nor NOR2 (N5195, N5192, N3369);
buf BUF1 (N5196, N5189);
and AND3 (N5197, N5180, N4301, N2695);
and AND3 (N5198, N5190, N2606, N3688);
not NOT1 (N5199, N5195);
and AND2 (N5200, N5199, N2358);
buf BUF1 (N5201, N5200);
nand NAND2 (N5202, N5183, N3944);
nor NOR2 (N5203, N5191, N4489);
buf BUF1 (N5204, N5196);
nor NOR2 (N5205, N5203, N638);
nand NAND3 (N5206, N5197, N2267, N2162);
nand NAND4 (N5207, N5186, N3760, N3915, N1858);
or OR4 (N5208, N5201, N4918, N1587, N2440);
nor NOR2 (N5209, N5194, N5018);
nor NOR4 (N5210, N5208, N685, N2600, N5015);
nand NAND2 (N5211, N5210, N4743);
xor XOR2 (N5212, N5207, N1961);
and AND2 (N5213, N5205, N1379);
nor NOR4 (N5214, N5206, N1751, N4973, N1960);
nand NAND3 (N5215, N5211, N4450, N911);
and AND2 (N5216, N5204, N4177);
buf BUF1 (N5217, N5198);
or OR3 (N5218, N5209, N4737, N3492);
xor XOR2 (N5219, N5212, N3621);
nor NOR2 (N5220, N5216, N3364);
xor XOR2 (N5221, N5217, N4466);
nor NOR4 (N5222, N5202, N4912, N2553, N2044);
xor XOR2 (N5223, N5215, N1059);
buf BUF1 (N5224, N5218);
not NOT1 (N5225, N5222);
not NOT1 (N5226, N5188);
not NOT1 (N5227, N5226);
buf BUF1 (N5228, N5223);
or OR3 (N5229, N5213, N3653, N3942);
and AND3 (N5230, N5219, N4788, N963);
not NOT1 (N5231, N5214);
nor NOR3 (N5232, N5224, N3480, N1440);
nor NOR4 (N5233, N5229, N4705, N673, N1547);
buf BUF1 (N5234, N5221);
nand NAND2 (N5235, N5234, N1535);
nor NOR3 (N5236, N5228, N3055, N3074);
not NOT1 (N5237, N5235);
nor NOR4 (N5238, N5233, N4825, N1526, N98);
not NOT1 (N5239, N5237);
nor NOR4 (N5240, N5231, N4772, N752, N3064);
or OR2 (N5241, N5230, N4928);
nand NAND4 (N5242, N5241, N686, N2989, N294);
or OR3 (N5243, N5240, N1643, N3899);
buf BUF1 (N5244, N5238);
xor XOR2 (N5245, N5232, N1978);
xor XOR2 (N5246, N5225, N3044);
not NOT1 (N5247, N5227);
or OR2 (N5248, N5220, N509);
not NOT1 (N5249, N5246);
nand NAND3 (N5250, N5247, N1035, N1363);
and AND4 (N5251, N5242, N2848, N1143, N4249);
nor NOR4 (N5252, N5248, N2259, N3878, N3357);
and AND3 (N5253, N5236, N3376, N1593);
buf BUF1 (N5254, N5249);
not NOT1 (N5255, N5252);
nand NAND2 (N5256, N5182, N1725);
nand NAND3 (N5257, N5253, N1976, N4983);
or OR4 (N5258, N5255, N2467, N3111, N957);
buf BUF1 (N5259, N5256);
nand NAND3 (N5260, N5250, N2858, N4487);
and AND4 (N5261, N5259, N3751, N3295, N2284);
buf BUF1 (N5262, N5260);
or OR3 (N5263, N5244, N1612, N4772);
not NOT1 (N5264, N5261);
buf BUF1 (N5265, N5245);
nand NAND3 (N5266, N5265, N3550, N5171);
and AND4 (N5267, N5263, N2669, N1015, N3357);
and AND4 (N5268, N5251, N170, N1047, N1391);
and AND3 (N5269, N5254, N2004, N131);
or OR3 (N5270, N5239, N4842, N693);
nand NAND3 (N5271, N5267, N5042, N1479);
or OR3 (N5272, N5268, N1648, N1263);
nor NOR2 (N5273, N5258, N745);
and AND4 (N5274, N5270, N3650, N2733, N1257);
nand NAND4 (N5275, N5272, N3146, N3654, N4120);
buf BUF1 (N5276, N5273);
or OR3 (N5277, N5274, N5214, N4715);
not NOT1 (N5278, N5262);
buf BUF1 (N5279, N5276);
nand NAND2 (N5280, N5243, N3481);
buf BUF1 (N5281, N5264);
or OR3 (N5282, N5275, N1716, N4459);
buf BUF1 (N5283, N5280);
buf BUF1 (N5284, N5283);
not NOT1 (N5285, N5266);
nand NAND4 (N5286, N5257, N3975, N4493, N37);
nor NOR2 (N5287, N5271, N333);
or OR2 (N5288, N5281, N3000);
not NOT1 (N5289, N5287);
buf BUF1 (N5290, N5269);
nor NOR2 (N5291, N5288, N3535);
xor XOR2 (N5292, N5282, N392);
nand NAND3 (N5293, N5292, N3512, N712);
xor XOR2 (N5294, N5289, N1994);
not NOT1 (N5295, N5286);
or OR3 (N5296, N5291, N1846, N3698);
or OR4 (N5297, N5294, N2474, N4851, N2789);
xor XOR2 (N5298, N5284, N285);
nand NAND4 (N5299, N5296, N2861, N2, N2478);
xor XOR2 (N5300, N5290, N1616);
not NOT1 (N5301, N5297);
or OR2 (N5302, N5277, N1824);
and AND3 (N5303, N5293, N2519, N1878);
and AND3 (N5304, N5298, N2231, N4286);
not NOT1 (N5305, N5279);
xor XOR2 (N5306, N5301, N2342);
buf BUF1 (N5307, N5303);
xor XOR2 (N5308, N5304, N5147);
buf BUF1 (N5309, N5295);
or OR4 (N5310, N5305, N409, N492, N2312);
buf BUF1 (N5311, N5302);
or OR3 (N5312, N5308, N5072, N2860);
buf BUF1 (N5313, N5311);
nand NAND2 (N5314, N5299, N4744);
or OR2 (N5315, N5309, N3432);
and AND4 (N5316, N5312, N909, N3626, N2602);
xor XOR2 (N5317, N5316, N347);
nand NAND3 (N5318, N5310, N2573, N2808);
nor NOR2 (N5319, N5307, N3219);
nor NOR4 (N5320, N5319, N1648, N1314, N328);
nor NOR2 (N5321, N5313, N817);
nor NOR3 (N5322, N5321, N1788, N4797);
xor XOR2 (N5323, N5278, N3830);
not NOT1 (N5324, N5320);
not NOT1 (N5325, N5322);
not NOT1 (N5326, N5306);
buf BUF1 (N5327, N5314);
nand NAND3 (N5328, N5323, N1023, N2686);
xor XOR2 (N5329, N5285, N3575);
buf BUF1 (N5330, N5315);
or OR4 (N5331, N5300, N465, N1906, N149);
xor XOR2 (N5332, N5331, N145);
nor NOR2 (N5333, N5326, N640);
nand NAND3 (N5334, N5329, N267, N466);
and AND3 (N5335, N5324, N4130, N2469);
nor NOR3 (N5336, N5330, N2078, N1265);
not NOT1 (N5337, N5327);
buf BUF1 (N5338, N5328);
nand NAND4 (N5339, N5325, N5222, N1000, N4002);
nand NAND4 (N5340, N5333, N4563, N5042, N4777);
nand NAND4 (N5341, N5338, N5032, N1436, N1044);
buf BUF1 (N5342, N5335);
nor NOR4 (N5343, N5341, N1425, N2635, N2964);
or OR2 (N5344, N5339, N1971);
xor XOR2 (N5345, N5342, N1499);
nor NOR4 (N5346, N5344, N1598, N5019, N2944);
buf BUF1 (N5347, N5340);
buf BUF1 (N5348, N5343);
nor NOR2 (N5349, N5336, N409);
and AND3 (N5350, N5337, N1365, N1392);
buf BUF1 (N5351, N5345);
not NOT1 (N5352, N5348);
buf BUF1 (N5353, N5349);
nor NOR4 (N5354, N5332, N5343, N2124, N1559);
and AND4 (N5355, N5351, N1676, N5197, N3670);
nand NAND4 (N5356, N5346, N3483, N3506, N410);
not NOT1 (N5357, N5356);
nor NOR3 (N5358, N5352, N221, N480);
buf BUF1 (N5359, N5347);
nor NOR2 (N5360, N5317, N1375);
or OR2 (N5361, N5354, N1248);
nand NAND3 (N5362, N5358, N3599, N3297);
not NOT1 (N5363, N5361);
not NOT1 (N5364, N5359);
xor XOR2 (N5365, N5334, N4121);
buf BUF1 (N5366, N5318);
xor XOR2 (N5367, N5350, N412);
nor NOR3 (N5368, N5363, N2845, N2432);
or OR4 (N5369, N5360, N2403, N648, N4119);
or OR3 (N5370, N5355, N357, N2521);
or OR4 (N5371, N5369, N601, N1881, N1723);
and AND3 (N5372, N5365, N3394, N277);
buf BUF1 (N5373, N5372);
buf BUF1 (N5374, N5366);
buf BUF1 (N5375, N5353);
nor NOR2 (N5376, N5357, N3135);
or OR2 (N5377, N5367, N1981);
buf BUF1 (N5378, N5362);
and AND2 (N5379, N5364, N3486);
xor XOR2 (N5380, N5378, N536);
or OR4 (N5381, N5371, N2563, N1567, N1338);
nand NAND3 (N5382, N5373, N3249, N3665);
or OR2 (N5383, N5374, N127);
xor XOR2 (N5384, N5377, N4388);
nand NAND2 (N5385, N5383, N3227);
xor XOR2 (N5386, N5382, N1258);
buf BUF1 (N5387, N5376);
or OR3 (N5388, N5386, N3276, N1214);
xor XOR2 (N5389, N5375, N3444);
buf BUF1 (N5390, N5380);
not NOT1 (N5391, N5379);
xor XOR2 (N5392, N5391, N3311);
xor XOR2 (N5393, N5384, N3573);
xor XOR2 (N5394, N5381, N1784);
xor XOR2 (N5395, N5393, N3018);
xor XOR2 (N5396, N5389, N1084);
not NOT1 (N5397, N5385);
nor NOR3 (N5398, N5388, N604, N4598);
not NOT1 (N5399, N5394);
nor NOR4 (N5400, N5398, N4455, N438, N4821);
buf BUF1 (N5401, N5395);
not NOT1 (N5402, N5397);
nor NOR3 (N5403, N5399, N4573, N141);
not NOT1 (N5404, N5390);
not NOT1 (N5405, N5396);
not NOT1 (N5406, N5402);
xor XOR2 (N5407, N5401, N4935);
or OR2 (N5408, N5368, N3472);
and AND4 (N5409, N5406, N674, N135, N1511);
nand NAND3 (N5410, N5400, N4525, N1547);
nor NOR2 (N5411, N5405, N4639);
buf BUF1 (N5412, N5408);
nand NAND3 (N5413, N5403, N5344, N5163);
nor NOR4 (N5414, N5392, N3614, N620, N4956);
buf BUF1 (N5415, N5404);
buf BUF1 (N5416, N5387);
buf BUF1 (N5417, N5414);
xor XOR2 (N5418, N5409, N4568);
nand NAND2 (N5419, N5411, N1419);
nor NOR3 (N5420, N5410, N4283, N3076);
buf BUF1 (N5421, N5420);
xor XOR2 (N5422, N5421, N5034);
and AND2 (N5423, N5415, N2236);
not NOT1 (N5424, N5416);
nand NAND3 (N5425, N5423, N1237, N3217);
and AND2 (N5426, N5424, N4784);
nor NOR3 (N5427, N5418, N644, N2919);
and AND3 (N5428, N5422, N2104, N2305);
nand NAND2 (N5429, N5419, N3750);
or OR2 (N5430, N5425, N2960);
nand NAND2 (N5431, N5429, N4521);
nand NAND4 (N5432, N5430, N427, N3947, N2918);
nand NAND4 (N5433, N5426, N4733, N3196, N1123);
not NOT1 (N5434, N5417);
nand NAND2 (N5435, N5433, N1698);
buf BUF1 (N5436, N5427);
or OR3 (N5437, N5407, N2890, N1044);
not NOT1 (N5438, N5435);
nand NAND3 (N5439, N5438, N1847, N5269);
not NOT1 (N5440, N5413);
not NOT1 (N5441, N5428);
xor XOR2 (N5442, N5436, N3051);
and AND2 (N5443, N5437, N824);
not NOT1 (N5444, N5370);
xor XOR2 (N5445, N5434, N319);
or OR2 (N5446, N5445, N5344);
and AND2 (N5447, N5412, N4531);
or OR4 (N5448, N5442, N4778, N4872, N3967);
nor NOR2 (N5449, N5440, N3780);
nand NAND4 (N5450, N5441, N4135, N4799, N612);
nor NOR4 (N5451, N5444, N250, N4665, N4461);
and AND3 (N5452, N5451, N1454, N3215);
nor NOR3 (N5453, N5443, N3931, N4884);
and AND2 (N5454, N5453, N149);
and AND2 (N5455, N5439, N5449);
not NOT1 (N5456, N3247);
or OR4 (N5457, N5455, N4172, N2850, N2874);
not NOT1 (N5458, N5447);
buf BUF1 (N5459, N5446);
xor XOR2 (N5460, N5452, N5269);
buf BUF1 (N5461, N5459);
xor XOR2 (N5462, N5454, N1777);
nand NAND4 (N5463, N5462, N2830, N2584, N293);
buf BUF1 (N5464, N5458);
or OR3 (N5465, N5461, N2040, N405);
not NOT1 (N5466, N5457);
not NOT1 (N5467, N5450);
or OR4 (N5468, N5463, N4714, N651, N2574);
not NOT1 (N5469, N5431);
nand NAND2 (N5470, N5460, N2080);
and AND4 (N5471, N5469, N3490, N1462, N5417);
xor XOR2 (N5472, N5464, N2240);
buf BUF1 (N5473, N5471);
not NOT1 (N5474, N5466);
and AND4 (N5475, N5473, N402, N766, N4829);
nor NOR2 (N5476, N5475, N844);
and AND4 (N5477, N5467, N3886, N1066, N2048);
not NOT1 (N5478, N5468);
or OR4 (N5479, N5472, N1170, N459, N2225);
xor XOR2 (N5480, N5448, N1036);
xor XOR2 (N5481, N5480, N3690);
nand NAND2 (N5482, N5476, N626);
buf BUF1 (N5483, N5432);
or OR4 (N5484, N5479, N922, N4431, N3303);
nor NOR4 (N5485, N5482, N1577, N209, N768);
not NOT1 (N5486, N5483);
xor XOR2 (N5487, N5470, N3473);
buf BUF1 (N5488, N5456);
and AND3 (N5489, N5481, N1661, N2553);
not NOT1 (N5490, N5488);
and AND3 (N5491, N5489, N1631, N1238);
nor NOR2 (N5492, N5491, N860);
nand NAND4 (N5493, N5492, N3582, N5130, N1418);
not NOT1 (N5494, N5493);
buf BUF1 (N5495, N5485);
and AND4 (N5496, N5494, N5384, N1977, N1657);
xor XOR2 (N5497, N5496, N1667);
buf BUF1 (N5498, N5484);
nor NOR2 (N5499, N5498, N525);
xor XOR2 (N5500, N5499, N3458);
or OR2 (N5501, N5486, N4936);
and AND3 (N5502, N5495, N5465, N4384);
nand NAND4 (N5503, N1673, N4769, N1739, N1221);
or OR3 (N5504, N5502, N1500, N3497);
or OR4 (N5505, N5487, N1464, N4516, N2463);
xor XOR2 (N5506, N5504, N2911);
xor XOR2 (N5507, N5505, N1809);
not NOT1 (N5508, N5503);
nor NOR2 (N5509, N5497, N3056);
or OR3 (N5510, N5478, N2894, N4087);
not NOT1 (N5511, N5477);
and AND2 (N5512, N5474, N3389);
nor NOR3 (N5513, N5509, N897, N918);
nand NAND3 (N5514, N5512, N471, N3311);
and AND2 (N5515, N5510, N1812);
buf BUF1 (N5516, N5490);
nand NAND3 (N5517, N5511, N524, N1178);
nand NAND3 (N5518, N5516, N1434, N3287);
and AND4 (N5519, N5513, N67, N2368, N1539);
nor NOR2 (N5520, N5506, N4631);
and AND2 (N5521, N5508, N4219);
nand NAND3 (N5522, N5519, N4093, N4685);
nand NAND2 (N5523, N5515, N2577);
not NOT1 (N5524, N5517);
nor NOR3 (N5525, N5501, N2047, N3313);
nand NAND4 (N5526, N5524, N4284, N4681, N2892);
and AND3 (N5527, N5523, N4145, N4236);
nor NOR2 (N5528, N5518, N101);
xor XOR2 (N5529, N5525, N411);
nor NOR4 (N5530, N5514, N1336, N2185, N1415);
and AND4 (N5531, N5500, N2545, N3523, N5105);
buf BUF1 (N5532, N5507);
nor NOR4 (N5533, N5521, N475, N3199, N4);
and AND3 (N5534, N5529, N4066, N4110);
xor XOR2 (N5535, N5528, N4684);
and AND3 (N5536, N5532, N4803, N4450);
nand NAND2 (N5537, N5531, N5291);
nand NAND3 (N5538, N5535, N2643, N3510);
nand NAND3 (N5539, N5520, N2347, N3404);
xor XOR2 (N5540, N5538, N286);
nand NAND4 (N5541, N5540, N5081, N2046, N5155);
nand NAND4 (N5542, N5526, N3266, N726, N849);
nor NOR4 (N5543, N5537, N3339, N2498, N4081);
not NOT1 (N5544, N5541);
xor XOR2 (N5545, N5533, N2522);
nand NAND2 (N5546, N5534, N5289);
nand NAND2 (N5547, N5530, N1967);
and AND2 (N5548, N5546, N1827);
buf BUF1 (N5549, N5544);
nand NAND3 (N5550, N5545, N2219, N2650);
and AND2 (N5551, N5536, N4355);
and AND4 (N5552, N5543, N498, N3498, N3689);
nand NAND2 (N5553, N5539, N3973);
nor NOR2 (N5554, N5551, N1873);
xor XOR2 (N5555, N5554, N2161);
not NOT1 (N5556, N5549);
and AND2 (N5557, N5522, N1868);
not NOT1 (N5558, N5557);
nor NOR3 (N5559, N5542, N3429, N1922);
nand NAND2 (N5560, N5556, N4481);
buf BUF1 (N5561, N5548);
buf BUF1 (N5562, N5550);
or OR3 (N5563, N5561, N2632, N5112);
and AND2 (N5564, N5559, N1600);
and AND3 (N5565, N5560, N3321, N3245);
or OR3 (N5566, N5563, N582, N1468);
nand NAND3 (N5567, N5566, N5178, N1847);
xor XOR2 (N5568, N5552, N3924);
nor NOR2 (N5569, N5564, N5123);
nand NAND3 (N5570, N5562, N5022, N4166);
nor NOR3 (N5571, N5569, N566, N1288);
and AND2 (N5572, N5570, N2128);
or OR3 (N5573, N5571, N543, N2835);
buf BUF1 (N5574, N5553);
xor XOR2 (N5575, N5527, N2393);
or OR2 (N5576, N5547, N3318);
not NOT1 (N5577, N5575);
nand NAND3 (N5578, N5573, N3615, N4795);
not NOT1 (N5579, N5578);
nand NAND4 (N5580, N5577, N3243, N996, N680);
nand NAND2 (N5581, N5576, N5000);
xor XOR2 (N5582, N5579, N3765);
nor NOR4 (N5583, N5580, N2725, N201, N4606);
not NOT1 (N5584, N5574);
and AND4 (N5585, N5582, N5220, N2646, N2425);
not NOT1 (N5586, N5585);
not NOT1 (N5587, N5586);
xor XOR2 (N5588, N5558, N1106);
not NOT1 (N5589, N5567);
not NOT1 (N5590, N5568);
nor NOR2 (N5591, N5588, N4151);
and AND3 (N5592, N5581, N666, N667);
nor NOR2 (N5593, N5572, N401);
or OR3 (N5594, N5555, N646, N1733);
not NOT1 (N5595, N5591);
nor NOR2 (N5596, N5589, N3706);
and AND2 (N5597, N5595, N1749);
not NOT1 (N5598, N5565);
and AND4 (N5599, N5596, N2726, N645, N2368);
nor NOR3 (N5600, N5583, N2621, N2408);
or OR4 (N5601, N5597, N2826, N1364, N4602);
xor XOR2 (N5602, N5590, N4304);
not NOT1 (N5603, N5592);
nand NAND3 (N5604, N5599, N5464, N1680);
nor NOR2 (N5605, N5584, N732);
nand NAND3 (N5606, N5587, N5418, N4153);
nor NOR2 (N5607, N5605, N4890);
and AND3 (N5608, N5604, N1914, N3855);
or OR2 (N5609, N5603, N5363);
or OR3 (N5610, N5602, N1299, N2161);
nand NAND2 (N5611, N5607, N785);
xor XOR2 (N5612, N5609, N1944);
nand NAND3 (N5613, N5600, N838, N622);
xor XOR2 (N5614, N5594, N1298);
nor NOR4 (N5615, N5613, N2715, N3301, N2045);
not NOT1 (N5616, N5612);
xor XOR2 (N5617, N5615, N650);
buf BUF1 (N5618, N5601);
buf BUF1 (N5619, N5617);
or OR3 (N5620, N5593, N801, N2549);
not NOT1 (N5621, N5606);
and AND4 (N5622, N5611, N566, N5, N3827);
xor XOR2 (N5623, N5608, N1143);
buf BUF1 (N5624, N5618);
nand NAND2 (N5625, N5616, N1506);
nand NAND3 (N5626, N5610, N1357, N3447);
xor XOR2 (N5627, N5598, N191);
nor NOR2 (N5628, N5620, N3650);
nor NOR2 (N5629, N5621, N2098);
nor NOR4 (N5630, N5626, N4547, N3564, N4505);
xor XOR2 (N5631, N5625, N1579);
buf BUF1 (N5632, N5622);
nand NAND3 (N5633, N5619, N499, N3051);
not NOT1 (N5634, N5632);
not NOT1 (N5635, N5614);
nand NAND4 (N5636, N5635, N2052, N2215, N1106);
not NOT1 (N5637, N5623);
nand NAND4 (N5638, N5630, N3377, N2233, N868);
or OR3 (N5639, N5628, N2819, N3076);
xor XOR2 (N5640, N5629, N2677);
or OR2 (N5641, N5640, N2526);
and AND4 (N5642, N5627, N2210, N1344, N4618);
and AND4 (N5643, N5633, N1814, N4194, N2607);
xor XOR2 (N5644, N5637, N2513);
nor NOR2 (N5645, N5634, N2711);
nand NAND4 (N5646, N5631, N5547, N1159, N386);
buf BUF1 (N5647, N5646);
not NOT1 (N5648, N5636);
xor XOR2 (N5649, N5638, N5166);
nor NOR2 (N5650, N5649, N827);
and AND2 (N5651, N5643, N871);
nand NAND3 (N5652, N5644, N4695, N2377);
not NOT1 (N5653, N5651);
nor NOR3 (N5654, N5639, N4002, N1306);
buf BUF1 (N5655, N5645);
and AND3 (N5656, N5641, N4288, N5223);
or OR2 (N5657, N5653, N1668);
nor NOR4 (N5658, N5642, N4289, N2879, N384);
xor XOR2 (N5659, N5624, N635);
nand NAND4 (N5660, N5659, N5334, N4121, N2243);
or OR3 (N5661, N5650, N1746, N3655);
nor NOR3 (N5662, N5657, N3113, N2915);
xor XOR2 (N5663, N5656, N3380);
or OR4 (N5664, N5662, N1490, N3134, N922);
nor NOR3 (N5665, N5652, N5213, N2216);
not NOT1 (N5666, N5664);
or OR3 (N5667, N5660, N4325, N801);
nor NOR3 (N5668, N5658, N1092, N2463);
and AND4 (N5669, N5663, N4606, N1932, N5338);
and AND4 (N5670, N5655, N3119, N829, N4449);
and AND2 (N5671, N5654, N429);
buf BUF1 (N5672, N5668);
nand NAND2 (N5673, N5661, N1939);
buf BUF1 (N5674, N5672);
or OR3 (N5675, N5647, N2523, N1432);
xor XOR2 (N5676, N5648, N662);
nor NOR3 (N5677, N5669, N3572, N66);
or OR4 (N5678, N5676, N4978, N191, N1665);
and AND2 (N5679, N5667, N4770);
and AND3 (N5680, N5679, N3857, N2856);
nor NOR4 (N5681, N5674, N4921, N2487, N4875);
or OR3 (N5682, N5666, N4291, N467);
or OR3 (N5683, N5673, N4202, N4197);
xor XOR2 (N5684, N5681, N834);
or OR4 (N5685, N5675, N1027, N4626, N2623);
buf BUF1 (N5686, N5682);
nor NOR2 (N5687, N5665, N5129);
nand NAND4 (N5688, N5670, N1050, N2471, N1653);
not NOT1 (N5689, N5686);
nor NOR4 (N5690, N5683, N5558, N3263, N2959);
nor NOR3 (N5691, N5685, N1910, N630);
not NOT1 (N5692, N5689);
and AND4 (N5693, N5692, N567, N3823, N1583);
and AND3 (N5694, N5688, N3898, N3758);
nand NAND4 (N5695, N5690, N3947, N254, N1709);
nand NAND4 (N5696, N5677, N2146, N2331, N4157);
xor XOR2 (N5697, N5691, N1965);
or OR2 (N5698, N5671, N601);
and AND4 (N5699, N5696, N4255, N1003, N3697);
nor NOR4 (N5700, N5693, N79, N1505, N4460);
or OR2 (N5701, N5695, N21);
xor XOR2 (N5702, N5701, N5106);
and AND4 (N5703, N5698, N3377, N3158, N1556);
nor NOR4 (N5704, N5684, N1065, N4593, N599);
xor XOR2 (N5705, N5700, N4421);
not NOT1 (N5706, N5687);
nor NOR3 (N5707, N5699, N3201, N756);
buf BUF1 (N5708, N5680);
nand NAND2 (N5709, N5703, N70);
and AND3 (N5710, N5697, N5634, N4650);
buf BUF1 (N5711, N5702);
nor NOR3 (N5712, N5711, N3058, N2030);
buf BUF1 (N5713, N5706);
or OR4 (N5714, N5705, N2093, N3906, N4947);
or OR4 (N5715, N5704, N5094, N384, N2843);
buf BUF1 (N5716, N5710);
nand NAND2 (N5717, N5713, N4091);
nor NOR4 (N5718, N5717, N948, N580, N5555);
nand NAND2 (N5719, N5707, N4942);
not NOT1 (N5720, N5678);
nand NAND3 (N5721, N5709, N4864, N1462);
and AND3 (N5722, N5720, N1253, N2069);
nor NOR3 (N5723, N5719, N3701, N1795);
nor NOR4 (N5724, N5723, N3933, N145, N382);
buf BUF1 (N5725, N5716);
and AND2 (N5726, N5725, N901);
and AND2 (N5727, N5712, N3354);
or OR4 (N5728, N5694, N2368, N1289, N1915);
nand NAND2 (N5729, N5722, N4820);
buf BUF1 (N5730, N5727);
and AND4 (N5731, N5708, N5026, N5349, N4980);
nor NOR4 (N5732, N5718, N692, N1147, N131);
xor XOR2 (N5733, N5726, N3911);
and AND3 (N5734, N5721, N4589, N344);
xor XOR2 (N5735, N5724, N4294);
buf BUF1 (N5736, N5734);
nor NOR3 (N5737, N5735, N2663, N278);
buf BUF1 (N5738, N5728);
nor NOR4 (N5739, N5731, N5636, N3447, N4901);
xor XOR2 (N5740, N5714, N4371);
or OR4 (N5741, N5733, N3955, N33, N4535);
not NOT1 (N5742, N5738);
nand NAND3 (N5743, N5729, N3164, N4336);
nand NAND3 (N5744, N5737, N929, N3380);
or OR3 (N5745, N5736, N3047, N2432);
or OR4 (N5746, N5730, N71, N1308, N5485);
xor XOR2 (N5747, N5742, N687);
not NOT1 (N5748, N5746);
xor XOR2 (N5749, N5741, N4088);
xor XOR2 (N5750, N5732, N1581);
xor XOR2 (N5751, N5740, N3020);
not NOT1 (N5752, N5748);
xor XOR2 (N5753, N5739, N4884);
not NOT1 (N5754, N5743);
not NOT1 (N5755, N5744);
or OR3 (N5756, N5715, N5066, N3397);
or OR3 (N5757, N5753, N3844, N1863);
or OR4 (N5758, N5747, N5099, N5296, N3235);
or OR2 (N5759, N5756, N5421);
or OR2 (N5760, N5745, N623);
nand NAND4 (N5761, N5759, N424, N2179, N4250);
nor NOR4 (N5762, N5754, N4887, N4434, N58);
and AND4 (N5763, N5762, N3698, N2221, N4820);
or OR3 (N5764, N5755, N4241, N3023);
not NOT1 (N5765, N5750);
not NOT1 (N5766, N5765);
nand NAND3 (N5767, N5761, N5684, N3293);
and AND4 (N5768, N5763, N1060, N2035, N4094);
nor NOR2 (N5769, N5752, N594);
nor NOR4 (N5770, N5749, N5679, N2511, N4629);
nor NOR2 (N5771, N5767, N3131);
or OR2 (N5772, N5770, N5579);
xor XOR2 (N5773, N5772, N4414);
buf BUF1 (N5774, N5757);
or OR4 (N5775, N5771, N2892, N2796, N350);
and AND2 (N5776, N5764, N5561);
not NOT1 (N5777, N5768);
nor NOR4 (N5778, N5777, N2071, N4837, N738);
and AND2 (N5779, N5751, N1639);
nor NOR2 (N5780, N5758, N4400);
buf BUF1 (N5781, N5778);
nand NAND3 (N5782, N5781, N590, N5781);
xor XOR2 (N5783, N5775, N4561);
not NOT1 (N5784, N5774);
nor NOR4 (N5785, N5782, N5547, N425, N3550);
xor XOR2 (N5786, N5773, N823);
xor XOR2 (N5787, N5760, N4684);
or OR2 (N5788, N5766, N3164);
not NOT1 (N5789, N5783);
buf BUF1 (N5790, N5776);
nand NAND2 (N5791, N5779, N4094);
nor NOR2 (N5792, N5769, N824);
and AND4 (N5793, N5791, N1334, N344, N4433);
nor NOR4 (N5794, N5787, N4463, N4893, N1461);
nand NAND3 (N5795, N5784, N3117, N106);
xor XOR2 (N5796, N5793, N1791);
or OR3 (N5797, N5795, N820, N2127);
nand NAND2 (N5798, N5780, N941);
or OR4 (N5799, N5790, N5177, N5332, N4451);
and AND3 (N5800, N5785, N5207, N5208);
not NOT1 (N5801, N5798);
and AND2 (N5802, N5801, N3948);
nor NOR4 (N5803, N5802, N1725, N5766, N3108);
xor XOR2 (N5804, N5792, N1770);
nand NAND4 (N5805, N5800, N3325, N4826, N2896);
and AND2 (N5806, N5788, N235);
nand NAND2 (N5807, N5806, N5475);
nor NOR2 (N5808, N5794, N2855);
buf BUF1 (N5809, N5804);
or OR2 (N5810, N5789, N5146);
nor NOR4 (N5811, N5796, N1940, N202, N810);
and AND3 (N5812, N5810, N4663, N2479);
not NOT1 (N5813, N5812);
nor NOR2 (N5814, N5799, N5316);
nor NOR4 (N5815, N5814, N4528, N4630, N3918);
xor XOR2 (N5816, N5805, N705);
and AND4 (N5817, N5797, N5571, N450, N4261);
or OR2 (N5818, N5807, N2431);
nand NAND4 (N5819, N5816, N527, N4798, N4681);
not NOT1 (N5820, N5815);
nand NAND4 (N5821, N5809, N375, N420, N5612);
nor NOR2 (N5822, N5818, N5781);
buf BUF1 (N5823, N5821);
nand NAND4 (N5824, N5786, N1506, N1903, N5098);
xor XOR2 (N5825, N5823, N5773);
and AND3 (N5826, N5819, N56, N4019);
and AND4 (N5827, N5825, N5247, N5269, N3919);
nor NOR4 (N5828, N5813, N662, N5434, N1747);
nor NOR2 (N5829, N5824, N3906);
or OR4 (N5830, N5817, N1310, N3880, N581);
nand NAND4 (N5831, N5827, N591, N4568, N2643);
not NOT1 (N5832, N5828);
nor NOR4 (N5833, N5811, N1984, N2991, N5558);
or OR3 (N5834, N5831, N2437, N3176);
xor XOR2 (N5835, N5808, N4212);
or OR4 (N5836, N5834, N4050, N883, N4365);
or OR4 (N5837, N5822, N5568, N5558, N1096);
not NOT1 (N5838, N5833);
nor NOR2 (N5839, N5838, N2211);
nor NOR4 (N5840, N5820, N4415, N2115, N3067);
nand NAND3 (N5841, N5840, N5784, N5235);
xor XOR2 (N5842, N5803, N4889);
not NOT1 (N5843, N5835);
and AND2 (N5844, N5842, N4391);
xor XOR2 (N5845, N5839, N2343);
nor NOR2 (N5846, N5844, N5571);
or OR2 (N5847, N5829, N4612);
and AND3 (N5848, N5841, N2336, N1434);
or OR3 (N5849, N5848, N3463, N19);
or OR4 (N5850, N5849, N486, N3952, N4676);
not NOT1 (N5851, N5850);
xor XOR2 (N5852, N5826, N4030);
buf BUF1 (N5853, N5846);
xor XOR2 (N5854, N5836, N142);
or OR4 (N5855, N5843, N4024, N408, N2750);
and AND3 (N5856, N5851, N2273, N690);
nand NAND4 (N5857, N5845, N917, N5357, N3642);
xor XOR2 (N5858, N5852, N5515);
nor NOR4 (N5859, N5857, N1646, N4159, N2929);
and AND2 (N5860, N5832, N3925);
nand NAND3 (N5861, N5859, N3949, N4167);
xor XOR2 (N5862, N5858, N2285);
xor XOR2 (N5863, N5855, N4563);
buf BUF1 (N5864, N5830);
or OR2 (N5865, N5864, N1335);
xor XOR2 (N5866, N5861, N4807);
nand NAND4 (N5867, N5854, N4721, N4559, N5077);
nor NOR2 (N5868, N5837, N1395);
nor NOR3 (N5869, N5860, N4076, N518);
or OR4 (N5870, N5856, N5467, N675, N2902);
nor NOR3 (N5871, N5847, N4042, N1957);
buf BUF1 (N5872, N5863);
nand NAND2 (N5873, N5872, N666);
buf BUF1 (N5874, N5868);
or OR2 (N5875, N5866, N115);
not NOT1 (N5876, N5862);
nand NAND3 (N5877, N5867, N1135, N1817);
or OR2 (N5878, N5870, N37);
nand NAND3 (N5879, N5871, N4112, N2635);
xor XOR2 (N5880, N5869, N2016);
and AND4 (N5881, N5877, N1982, N4028, N4365);
buf BUF1 (N5882, N5865);
nand NAND4 (N5883, N5875, N3402, N3926, N4502);
or OR4 (N5884, N5853, N3926, N2090, N2750);
nor NOR2 (N5885, N5883, N3119);
nor NOR4 (N5886, N5880, N3277, N3068, N832);
or OR4 (N5887, N5882, N2244, N1604, N5786);
or OR4 (N5888, N5886, N2953, N2098, N2189);
buf BUF1 (N5889, N5876);
not NOT1 (N5890, N5889);
nor NOR3 (N5891, N5884, N764, N3018);
and AND2 (N5892, N5874, N3030);
or OR2 (N5893, N5888, N1826);
or OR2 (N5894, N5885, N5459);
or OR3 (N5895, N5881, N1755, N4650);
or OR4 (N5896, N5891, N5699, N5786, N5728);
or OR2 (N5897, N5879, N5609);
buf BUF1 (N5898, N5873);
or OR4 (N5899, N5897, N3637, N1773, N5324);
buf BUF1 (N5900, N5896);
buf BUF1 (N5901, N5887);
or OR3 (N5902, N5894, N2021, N1770);
xor XOR2 (N5903, N5895, N5876);
and AND3 (N5904, N5900, N3891, N3622);
nand NAND4 (N5905, N5901, N5128, N936, N3497);
nor NOR3 (N5906, N5892, N5407, N189);
and AND3 (N5907, N5902, N4053, N3448);
nand NAND4 (N5908, N5906, N4532, N3336, N3932);
not NOT1 (N5909, N5908);
and AND4 (N5910, N5893, N2274, N289, N4930);
nor NOR3 (N5911, N5904, N5114, N1114);
nor NOR2 (N5912, N5911, N4871);
nand NAND4 (N5913, N5905, N1549, N3241, N3436);
or OR3 (N5914, N5899, N2423, N4302);
or OR2 (N5915, N5903, N136);
or OR2 (N5916, N5913, N403);
not NOT1 (N5917, N5910);
xor XOR2 (N5918, N5915, N249);
not NOT1 (N5919, N5912);
buf BUF1 (N5920, N5914);
or OR2 (N5921, N5878, N5734);
not NOT1 (N5922, N5898);
buf BUF1 (N5923, N5907);
nand NAND2 (N5924, N5920, N3831);
xor XOR2 (N5925, N5916, N1675);
nand NAND3 (N5926, N5917, N261, N5216);
and AND4 (N5927, N5922, N3934, N298, N3600);
or OR3 (N5928, N5918, N1924, N2634);
nor NOR2 (N5929, N5927, N1469);
xor XOR2 (N5930, N5919, N1596);
xor XOR2 (N5931, N5923, N2261);
and AND4 (N5932, N5926, N4985, N4112, N3448);
nand NAND3 (N5933, N5909, N2715, N3625);
xor XOR2 (N5934, N5932, N3304);
xor XOR2 (N5935, N5933, N4617);
nand NAND2 (N5936, N5928, N4852);
and AND3 (N5937, N5925, N2642, N5921);
nor NOR4 (N5938, N4829, N5678, N175, N4089);
xor XOR2 (N5939, N5890, N3808);
and AND2 (N5940, N5931, N253);
xor XOR2 (N5941, N5930, N2852);
nor NOR3 (N5942, N5941, N1430, N5422);
or OR3 (N5943, N5924, N5486, N2345);
nor NOR4 (N5944, N5935, N5851, N1560, N913);
nor NOR2 (N5945, N5936, N2746);
xor XOR2 (N5946, N5937, N3933);
or OR2 (N5947, N5929, N1710);
or OR2 (N5948, N5942, N3366);
nand NAND3 (N5949, N5944, N3359, N5740);
and AND2 (N5950, N5940, N3814);
nor NOR4 (N5951, N5934, N2420, N3353, N332);
not NOT1 (N5952, N5939);
xor XOR2 (N5953, N5949, N3735);
nor NOR4 (N5954, N5946, N5510, N714, N583);
nand NAND4 (N5955, N5951, N5632, N543, N1687);
xor XOR2 (N5956, N5950, N582);
buf BUF1 (N5957, N5943);
buf BUF1 (N5958, N5952);
buf BUF1 (N5959, N5953);
xor XOR2 (N5960, N5938, N3272);
buf BUF1 (N5961, N5955);
and AND4 (N5962, N5959, N51, N3867, N2664);
and AND2 (N5963, N5948, N275);
nand NAND2 (N5964, N5957, N4011);
nor NOR4 (N5965, N5958, N738, N1793, N2422);
or OR3 (N5966, N5960, N2848, N125);
and AND4 (N5967, N5954, N4009, N696, N2704);
or OR3 (N5968, N5966, N1730, N2820);
nor NOR3 (N5969, N5964, N761, N1809);
buf BUF1 (N5970, N5965);
nor NOR4 (N5971, N5945, N439, N2698, N2731);
nand NAND2 (N5972, N5962, N4110);
xor XOR2 (N5973, N5947, N1314);
nand NAND3 (N5974, N5971, N4153, N1704);
buf BUF1 (N5975, N5974);
not NOT1 (N5976, N5967);
nor NOR2 (N5977, N5970, N3029);
nand NAND4 (N5978, N5969, N467, N2181, N1607);
and AND4 (N5979, N5978, N4218, N5142, N2772);
not NOT1 (N5980, N5963);
nor NOR4 (N5981, N5961, N5056, N2485, N5838);
not NOT1 (N5982, N5979);
not NOT1 (N5983, N5956);
buf BUF1 (N5984, N5975);
xor XOR2 (N5985, N5984, N1616);
xor XOR2 (N5986, N5976, N4289);
and AND4 (N5987, N5972, N5240, N1827, N2480);
xor XOR2 (N5988, N5968, N5790);
nor NOR4 (N5989, N5980, N3407, N1981, N3378);
nor NOR3 (N5990, N5986, N5106, N4085);
nor NOR4 (N5991, N5982, N5138, N5751, N4081);
or OR2 (N5992, N5983, N3472);
and AND3 (N5993, N5989, N4076, N2592);
xor XOR2 (N5994, N5985, N2035);
and AND2 (N5995, N5981, N906);
and AND3 (N5996, N5973, N4345, N1280);
xor XOR2 (N5997, N5977, N5504);
nand NAND3 (N5998, N5991, N2442, N2259);
and AND2 (N5999, N5993, N5553);
nand NAND3 (N6000, N5990, N4337, N830);
not NOT1 (N6001, N5999);
not NOT1 (N6002, N5994);
nand NAND3 (N6003, N5988, N2637, N706);
nor NOR2 (N6004, N5995, N949);
not NOT1 (N6005, N5992);
nand NAND2 (N6006, N6004, N841);
nor NOR2 (N6007, N6002, N5069);
not NOT1 (N6008, N5997);
nor NOR4 (N6009, N5996, N1526, N1296, N2074);
and AND2 (N6010, N6007, N503);
xor XOR2 (N6011, N6008, N1052);
not NOT1 (N6012, N6010);
not NOT1 (N6013, N6012);
xor XOR2 (N6014, N6000, N948);
xor XOR2 (N6015, N5998, N725);
nand NAND4 (N6016, N5987, N4476, N3785, N4657);
and AND2 (N6017, N6001, N4992);
nor NOR4 (N6018, N6009, N1350, N2334, N5384);
buf BUF1 (N6019, N6011);
or OR3 (N6020, N6018, N2883, N1068);
buf BUF1 (N6021, N6016);
not NOT1 (N6022, N6014);
buf BUF1 (N6023, N6020);
xor XOR2 (N6024, N6019, N4474);
not NOT1 (N6025, N6017);
nand NAND2 (N6026, N6006, N2519);
not NOT1 (N6027, N6024);
not NOT1 (N6028, N6025);
not NOT1 (N6029, N6013);
xor XOR2 (N6030, N6021, N1844);
or OR3 (N6031, N6003, N5015, N4377);
nor NOR4 (N6032, N6031, N5117, N2865, N4376);
buf BUF1 (N6033, N6030);
nand NAND3 (N6034, N6026, N2037, N754);
nor NOR2 (N6035, N6022, N4528);
buf BUF1 (N6036, N6034);
xor XOR2 (N6037, N6035, N812);
nor NOR3 (N6038, N6015, N5406, N1785);
and AND3 (N6039, N6028, N5653, N1175);
and AND3 (N6040, N6027, N4509, N5003);
buf BUF1 (N6041, N6037);
xor XOR2 (N6042, N6036, N5785);
buf BUF1 (N6043, N6039);
and AND3 (N6044, N6040, N3850, N1063);
not NOT1 (N6045, N6033);
or OR4 (N6046, N6045, N307, N1247, N4839);
not NOT1 (N6047, N6042);
nand NAND2 (N6048, N6005, N3169);
nor NOR2 (N6049, N6023, N4057);
not NOT1 (N6050, N6043);
xor XOR2 (N6051, N6047, N5110);
nand NAND3 (N6052, N6050, N2076, N1672);
and AND2 (N6053, N6041, N4444);
or OR4 (N6054, N6044, N2195, N6012, N4351);
buf BUF1 (N6055, N6051);
nor NOR2 (N6056, N6038, N2217);
buf BUF1 (N6057, N6029);
nor NOR4 (N6058, N6054, N1579, N3865, N3365);
not NOT1 (N6059, N6056);
and AND4 (N6060, N6032, N5740, N2790, N5572);
xor XOR2 (N6061, N6049, N171);
not NOT1 (N6062, N6061);
xor XOR2 (N6063, N6057, N3500);
xor XOR2 (N6064, N6053, N3666);
or OR4 (N6065, N6063, N5422, N2900, N826);
or OR3 (N6066, N6046, N449, N3468);
nor NOR3 (N6067, N6064, N3681, N1648);
buf BUF1 (N6068, N6065);
and AND4 (N6069, N6062, N2059, N846, N4579);
nand NAND4 (N6070, N6068, N3698, N5222, N2052);
not NOT1 (N6071, N6067);
and AND2 (N6072, N6058, N1919);
xor XOR2 (N6073, N6069, N343);
nor NOR2 (N6074, N6072, N5408);
not NOT1 (N6075, N6048);
not NOT1 (N6076, N6070);
and AND4 (N6077, N6076, N284, N3781, N4992);
or OR2 (N6078, N6060, N4016);
xor XOR2 (N6079, N6078, N5604);
buf BUF1 (N6080, N6059);
nor NOR2 (N6081, N6079, N2064);
nor NOR2 (N6082, N6077, N2392);
nand NAND4 (N6083, N6082, N5881, N3241, N757);
not NOT1 (N6084, N6071);
or OR4 (N6085, N6052, N144, N4782, N2221);
nor NOR3 (N6086, N6073, N4923, N5182);
nand NAND2 (N6087, N6066, N4798);
and AND3 (N6088, N6083, N403, N195);
and AND3 (N6089, N6088, N4680, N3195);
nand NAND4 (N6090, N6074, N690, N5518, N1393);
buf BUF1 (N6091, N6075);
nor NOR4 (N6092, N6055, N2464, N3017, N1694);
and AND3 (N6093, N6090, N2517, N69);
xor XOR2 (N6094, N6081, N4126);
and AND2 (N6095, N6087, N28);
or OR3 (N6096, N6080, N5798, N3920);
xor XOR2 (N6097, N6095, N1885);
nand NAND3 (N6098, N6085, N475, N4819);
nand NAND3 (N6099, N6098, N1004, N4802);
or OR3 (N6100, N6091, N4969, N1114);
or OR4 (N6101, N6089, N5791, N4178, N2842);
xor XOR2 (N6102, N6099, N614);
and AND4 (N6103, N6093, N1841, N3200, N5347);
nand NAND4 (N6104, N6097, N668, N4401, N2500);
not NOT1 (N6105, N6094);
xor XOR2 (N6106, N6104, N3462);
buf BUF1 (N6107, N6084);
buf BUF1 (N6108, N6105);
or OR3 (N6109, N6096, N1215, N4848);
or OR4 (N6110, N6108, N761, N632, N4265);
not NOT1 (N6111, N6107);
nand NAND3 (N6112, N6092, N1574, N2014);
and AND2 (N6113, N6110, N5893);
or OR4 (N6114, N6109, N2525, N2421, N627);
or OR3 (N6115, N6111, N1280, N46);
not NOT1 (N6116, N6106);
not NOT1 (N6117, N6101);
buf BUF1 (N6118, N6113);
xor XOR2 (N6119, N6116, N5541);
not NOT1 (N6120, N6114);
and AND2 (N6121, N6119, N4133);
and AND3 (N6122, N6112, N607, N3497);
nor NOR4 (N6123, N6117, N3237, N158, N2234);
xor XOR2 (N6124, N6115, N5540);
nand NAND3 (N6125, N6122, N3719, N1540);
and AND2 (N6126, N6124, N3796);
not NOT1 (N6127, N6086);
and AND4 (N6128, N6100, N4609, N3607, N4959);
buf BUF1 (N6129, N6127);
and AND3 (N6130, N6129, N4327, N5266);
and AND4 (N6131, N6125, N5378, N2495, N991);
buf BUF1 (N6132, N6130);
or OR4 (N6133, N6118, N2022, N2776, N3103);
not NOT1 (N6134, N6131);
buf BUF1 (N6135, N6132);
xor XOR2 (N6136, N6123, N5740);
and AND3 (N6137, N6136, N2676, N3616);
buf BUF1 (N6138, N6103);
or OR3 (N6139, N6133, N3363, N3743);
buf BUF1 (N6140, N6128);
xor XOR2 (N6141, N6140, N5968);
nand NAND2 (N6142, N6121, N2979);
not NOT1 (N6143, N6137);
or OR4 (N6144, N6141, N4291, N1539, N984);
nor NOR4 (N6145, N6144, N1096, N1364, N2433);
nor NOR3 (N6146, N6102, N5215, N3622);
xor XOR2 (N6147, N6120, N4225);
xor XOR2 (N6148, N6126, N3599);
xor XOR2 (N6149, N6143, N3159);
nand NAND2 (N6150, N6134, N713);
and AND3 (N6151, N6146, N5037, N2964);
and AND3 (N6152, N6142, N5842, N2383);
nor NOR4 (N6153, N6147, N3914, N1408, N3109);
buf BUF1 (N6154, N6148);
and AND4 (N6155, N6145, N3443, N3561, N821);
nor NOR2 (N6156, N6152, N787);
and AND4 (N6157, N6151, N3179, N4372, N3725);
nand NAND2 (N6158, N6135, N2740);
xor XOR2 (N6159, N6150, N3035);
buf BUF1 (N6160, N6158);
nand NAND2 (N6161, N6138, N6005);
nand NAND4 (N6162, N6149, N3677, N1022, N2267);
and AND3 (N6163, N6155, N4220, N1349);
nand NAND4 (N6164, N6157, N3818, N1386, N5461);
nand NAND4 (N6165, N6164, N4946, N5292, N293);
nor NOR3 (N6166, N6153, N5099, N2310);
not NOT1 (N6167, N6166);
nor NOR2 (N6168, N6154, N5714);
or OR4 (N6169, N6167, N5454, N3455, N4609);
buf BUF1 (N6170, N6169);
xor XOR2 (N6171, N6165, N2107);
xor XOR2 (N6172, N6156, N175);
nor NOR2 (N6173, N6160, N3356);
nand NAND3 (N6174, N6168, N5359, N336);
or OR3 (N6175, N6174, N4163, N850);
or OR3 (N6176, N6162, N6025, N5345);
nand NAND3 (N6177, N6161, N5225, N836);
buf BUF1 (N6178, N6163);
not NOT1 (N6179, N6172);
xor XOR2 (N6180, N6176, N5689);
nand NAND4 (N6181, N6170, N4573, N5660, N1586);
not NOT1 (N6182, N6171);
and AND2 (N6183, N6179, N721);
buf BUF1 (N6184, N6182);
not NOT1 (N6185, N6175);
and AND4 (N6186, N6181, N2774, N5282, N5197);
not NOT1 (N6187, N6185);
buf BUF1 (N6188, N6183);
nand NAND2 (N6189, N6184, N4144);
buf BUF1 (N6190, N6189);
nand NAND2 (N6191, N6177, N761);
not NOT1 (N6192, N6180);
xor XOR2 (N6193, N6178, N5177);
not NOT1 (N6194, N6159);
and AND2 (N6195, N6192, N855);
nand NAND4 (N6196, N6194, N2056, N3459, N5227);
nand NAND2 (N6197, N6186, N4190);
and AND2 (N6198, N6195, N1813);
not NOT1 (N6199, N6193);
nor NOR4 (N6200, N6191, N6163, N2631, N923);
or OR3 (N6201, N6198, N367, N3327);
not NOT1 (N6202, N6173);
or OR2 (N6203, N6190, N2681);
not NOT1 (N6204, N6199);
xor XOR2 (N6205, N6187, N1062);
nand NAND3 (N6206, N6205, N5338, N3184);
xor XOR2 (N6207, N6203, N651);
xor XOR2 (N6208, N6139, N2188);
or OR3 (N6209, N6201, N4950, N3419);
nor NOR2 (N6210, N6206, N3923);
and AND2 (N6211, N6200, N2458);
nor NOR3 (N6212, N6209, N4211, N1692);
xor XOR2 (N6213, N6207, N776);
not NOT1 (N6214, N6196);
buf BUF1 (N6215, N6188);
and AND4 (N6216, N6204, N5820, N3540, N3273);
or OR2 (N6217, N6197, N3887);
and AND4 (N6218, N6208, N2871, N4505, N5305);
and AND2 (N6219, N6211, N2139);
and AND2 (N6220, N6216, N913);
or OR2 (N6221, N6212, N3706);
buf BUF1 (N6222, N6213);
xor XOR2 (N6223, N6210, N5190);
nor NOR2 (N6224, N6214, N1018);
or OR4 (N6225, N6215, N5414, N2845, N4973);
buf BUF1 (N6226, N6224);
not NOT1 (N6227, N6222);
buf BUF1 (N6228, N6202);
not NOT1 (N6229, N6223);
xor XOR2 (N6230, N6217, N6138);
or OR3 (N6231, N6227, N6182, N6022);
nand NAND4 (N6232, N6219, N488, N3246, N2001);
or OR3 (N6233, N6221, N4929, N1361);
and AND4 (N6234, N6225, N4154, N5941, N4353);
nand NAND4 (N6235, N6234, N2936, N6207, N6058);
nor NOR2 (N6236, N6228, N4559);
or OR2 (N6237, N6230, N3664);
or OR2 (N6238, N6237, N4354);
or OR4 (N6239, N6238, N1308, N1648, N5790);
nor NOR4 (N6240, N6233, N3544, N2055, N5068);
buf BUF1 (N6241, N6231);
or OR4 (N6242, N6226, N1685, N958, N2533);
nor NOR2 (N6243, N6241, N5552);
nand NAND4 (N6244, N6240, N2984, N2735, N2045);
or OR4 (N6245, N6236, N1092, N1917, N3542);
and AND4 (N6246, N6239, N4108, N3700, N3593);
not NOT1 (N6247, N6235);
buf BUF1 (N6248, N6242);
not NOT1 (N6249, N6232);
or OR4 (N6250, N6229, N5412, N3326, N5933);
nor NOR3 (N6251, N6243, N718, N358);
nand NAND3 (N6252, N6248, N1832, N2845);
and AND4 (N6253, N6249, N491, N2249, N2417);
nand NAND4 (N6254, N6253, N4435, N667, N572);
not NOT1 (N6255, N6245);
or OR3 (N6256, N6246, N3015, N2666);
nor NOR4 (N6257, N6220, N4374, N1274, N1958);
nand NAND3 (N6258, N6257, N6163, N4196);
nor NOR3 (N6259, N6244, N891, N739);
not NOT1 (N6260, N6254);
or OR4 (N6261, N6258, N2261, N625, N2927);
or OR3 (N6262, N6261, N4457, N4992);
nor NOR2 (N6263, N6252, N2983);
and AND3 (N6264, N6250, N3860, N4902);
and AND4 (N6265, N6218, N3936, N5940, N3884);
xor XOR2 (N6266, N6264, N4709);
buf BUF1 (N6267, N6247);
nor NOR4 (N6268, N6260, N1834, N5665, N5807);
buf BUF1 (N6269, N6265);
xor XOR2 (N6270, N6251, N931);
xor XOR2 (N6271, N6270, N1559);
or OR3 (N6272, N6266, N173, N3541);
xor XOR2 (N6273, N6259, N3901);
nor NOR2 (N6274, N6256, N1837);
xor XOR2 (N6275, N6268, N760);
xor XOR2 (N6276, N6263, N708);
not NOT1 (N6277, N6275);
and AND3 (N6278, N6255, N4494, N6170);
or OR2 (N6279, N6276, N2795);
or OR3 (N6280, N6274, N5106, N4678);
nand NAND3 (N6281, N6269, N795, N377);
and AND3 (N6282, N6273, N4159, N3054);
not NOT1 (N6283, N6281);
nand NAND3 (N6284, N6279, N1786, N3531);
nand NAND3 (N6285, N6262, N574, N528);
xor XOR2 (N6286, N6267, N3459);
nand NAND2 (N6287, N6272, N4753);
not NOT1 (N6288, N6283);
or OR4 (N6289, N6277, N969, N4668, N3773);
xor XOR2 (N6290, N6287, N2653);
buf BUF1 (N6291, N6280);
or OR3 (N6292, N6291, N495, N3392);
and AND4 (N6293, N6290, N1110, N1750, N2322);
not NOT1 (N6294, N6278);
not NOT1 (N6295, N6292);
and AND2 (N6296, N6282, N465);
and AND2 (N6297, N6288, N552);
or OR4 (N6298, N6271, N4298, N919, N1460);
xor XOR2 (N6299, N6285, N3335);
not NOT1 (N6300, N6295);
nor NOR4 (N6301, N6284, N4119, N3516, N624);
not NOT1 (N6302, N6297);
nor NOR3 (N6303, N6298, N3252, N620);
nand NAND3 (N6304, N6299, N4671, N1468);
not NOT1 (N6305, N6294);
or OR2 (N6306, N6286, N3019);
xor XOR2 (N6307, N6304, N396);
nor NOR3 (N6308, N6306, N2231, N214);
nor NOR2 (N6309, N6293, N492);
xor XOR2 (N6310, N6289, N178);
nand NAND4 (N6311, N6308, N3205, N5506, N4263);
not NOT1 (N6312, N6307);
or OR3 (N6313, N6303, N3981, N1943);
not NOT1 (N6314, N6300);
or OR4 (N6315, N6313, N5016, N4441, N4591);
not NOT1 (N6316, N6312);
or OR2 (N6317, N6301, N3309);
or OR3 (N6318, N6317, N2055, N5979);
or OR3 (N6319, N6310, N4035, N4119);
xor XOR2 (N6320, N6309, N3523);
or OR4 (N6321, N6305, N3964, N5060, N3850);
nand NAND4 (N6322, N6315, N5753, N4190, N1817);
xor XOR2 (N6323, N6321, N1542);
buf BUF1 (N6324, N6311);
or OR2 (N6325, N6318, N536);
nand NAND4 (N6326, N6319, N1951, N2137, N5198);
and AND2 (N6327, N6296, N3957);
not NOT1 (N6328, N6323);
nor NOR2 (N6329, N6316, N2091);
or OR4 (N6330, N6326, N4744, N1785, N5241);
buf BUF1 (N6331, N6328);
not NOT1 (N6332, N6322);
nor NOR3 (N6333, N6324, N3270, N6031);
not NOT1 (N6334, N6331);
nand NAND3 (N6335, N6325, N5764, N4020);
nand NAND4 (N6336, N6302, N3597, N406, N1467);
xor XOR2 (N6337, N6330, N3115);
or OR4 (N6338, N6327, N4099, N1996, N528);
or OR4 (N6339, N6333, N5391, N5107, N2482);
xor XOR2 (N6340, N6329, N276);
and AND3 (N6341, N6335, N3862, N1337);
not NOT1 (N6342, N6334);
nor NOR3 (N6343, N6340, N5055, N2186);
nand NAND4 (N6344, N6341, N140, N3490, N6148);
nand NAND2 (N6345, N6336, N3938);
or OR3 (N6346, N6339, N86, N1969);
and AND4 (N6347, N6332, N2444, N5060, N5818);
not NOT1 (N6348, N6314);
and AND4 (N6349, N6345, N3338, N4992, N4983);
nor NOR4 (N6350, N6342, N248, N5967, N1460);
nand NAND2 (N6351, N6343, N3423);
or OR4 (N6352, N6349, N40, N4949, N3851);
not NOT1 (N6353, N6352);
nand NAND2 (N6354, N6320, N2948);
and AND4 (N6355, N6351, N2426, N474, N4169);
or OR4 (N6356, N6348, N3917, N5264, N3970);
xor XOR2 (N6357, N6355, N3219);
not NOT1 (N6358, N6350);
xor XOR2 (N6359, N6338, N5717);
not NOT1 (N6360, N6347);
nor NOR4 (N6361, N6344, N3979, N354, N4125);
not NOT1 (N6362, N6337);
buf BUF1 (N6363, N6353);
or OR4 (N6364, N6360, N6077, N3569, N2997);
or OR4 (N6365, N6356, N2562, N164, N16);
xor XOR2 (N6366, N6346, N6043);
nor NOR2 (N6367, N6359, N5198);
nand NAND2 (N6368, N6363, N2048);
or OR4 (N6369, N6367, N4813, N4396, N2592);
and AND4 (N6370, N6362, N5421, N1701, N2015);
buf BUF1 (N6371, N6357);
buf BUF1 (N6372, N6370);
not NOT1 (N6373, N6361);
not NOT1 (N6374, N6364);
buf BUF1 (N6375, N6354);
and AND3 (N6376, N6372, N1240, N696);
buf BUF1 (N6377, N6375);
or OR2 (N6378, N6376, N5882);
nor NOR3 (N6379, N6371, N1543, N1800);
or OR2 (N6380, N6379, N631);
or OR4 (N6381, N6366, N3928, N30, N285);
or OR2 (N6382, N6369, N4563);
buf BUF1 (N6383, N6382);
or OR2 (N6384, N6380, N1280);
xor XOR2 (N6385, N6373, N4938);
and AND3 (N6386, N6365, N5384, N3723);
buf BUF1 (N6387, N6368);
not NOT1 (N6388, N6378);
buf BUF1 (N6389, N6383);
not NOT1 (N6390, N6374);
or OR3 (N6391, N6389, N3761, N16);
xor XOR2 (N6392, N6381, N4815);
and AND4 (N6393, N6392, N666, N1407, N305);
and AND4 (N6394, N6391, N4429, N4923, N4653);
nor NOR3 (N6395, N6390, N3193, N6252);
xor XOR2 (N6396, N6393, N185);
and AND4 (N6397, N6396, N747, N3670, N2305);
buf BUF1 (N6398, N6395);
not NOT1 (N6399, N6397);
xor XOR2 (N6400, N6358, N2246);
nand NAND2 (N6401, N6394, N2766);
xor XOR2 (N6402, N6386, N2621);
xor XOR2 (N6403, N6399, N2533);
nand NAND2 (N6404, N6400, N5531);
and AND4 (N6405, N6404, N6219, N1449, N5933);
nor NOR2 (N6406, N6405, N6253);
not NOT1 (N6407, N6401);
xor XOR2 (N6408, N6377, N2459);
not NOT1 (N6409, N6407);
nor NOR3 (N6410, N6408, N5436, N4412);
xor XOR2 (N6411, N6403, N157);
nor NOR4 (N6412, N6398, N5852, N5380, N4398);
not NOT1 (N6413, N6410);
xor XOR2 (N6414, N6384, N1365);
and AND4 (N6415, N6387, N3169, N4304, N5791);
not NOT1 (N6416, N6413);
xor XOR2 (N6417, N6406, N4771);
buf BUF1 (N6418, N6385);
or OR3 (N6419, N6402, N4364, N53);
and AND2 (N6420, N6415, N1301);
or OR3 (N6421, N6412, N2045, N2402);
buf BUF1 (N6422, N6409);
not NOT1 (N6423, N6416);
and AND3 (N6424, N6420, N412, N5571);
nor NOR2 (N6425, N6423, N2154);
and AND4 (N6426, N6414, N3137, N2190, N5048);
not NOT1 (N6427, N6388);
not NOT1 (N6428, N6422);
not NOT1 (N6429, N6425);
or OR4 (N6430, N6424, N2369, N2633, N2616);
nor NOR4 (N6431, N6428, N4742, N4296, N2827);
xor XOR2 (N6432, N6429, N5567);
not NOT1 (N6433, N6426);
xor XOR2 (N6434, N6433, N3691);
nand NAND4 (N6435, N6421, N606, N5252, N5558);
nor NOR2 (N6436, N6434, N1997);
buf BUF1 (N6437, N6427);
nor NOR2 (N6438, N6417, N2637);
not NOT1 (N6439, N6431);
nand NAND2 (N6440, N6411, N4831);
nor NOR4 (N6441, N6432, N811, N1010, N1275);
and AND3 (N6442, N6419, N3124, N2304);
nor NOR4 (N6443, N6439, N4478, N4479, N1113);
buf BUF1 (N6444, N6418);
nand NAND3 (N6445, N6440, N2341, N286);
not NOT1 (N6446, N6442);
not NOT1 (N6447, N6430);
or OR4 (N6448, N6436, N843, N6439, N716);
nor NOR4 (N6449, N6448, N2628, N6326, N5038);
nor NOR3 (N6450, N6449, N658, N4432);
not NOT1 (N6451, N6446);
not NOT1 (N6452, N6437);
not NOT1 (N6453, N6450);
nor NOR2 (N6454, N6444, N4870);
xor XOR2 (N6455, N6454, N6383);
and AND3 (N6456, N6438, N5891, N3057);
or OR3 (N6457, N6452, N2844, N2900);
nand NAND2 (N6458, N6435, N6092);
nor NOR2 (N6459, N6455, N4942);
nand NAND4 (N6460, N6456, N6177, N3407, N2250);
nand NAND4 (N6461, N6441, N3832, N3559, N4487);
buf BUF1 (N6462, N6461);
and AND3 (N6463, N6460, N231, N401);
nor NOR4 (N6464, N6447, N2198, N667, N2049);
buf BUF1 (N6465, N6459);
and AND2 (N6466, N6463, N3930);
nor NOR3 (N6467, N6464, N5410, N3300);
buf BUF1 (N6468, N6467);
nand NAND4 (N6469, N6468, N3824, N1000, N415);
xor XOR2 (N6470, N6462, N5634);
xor XOR2 (N6471, N6443, N6280);
and AND4 (N6472, N6465, N3660, N5948, N2348);
nor NOR3 (N6473, N6457, N1014, N2290);
or OR4 (N6474, N6472, N5490, N4936, N6469);
and AND2 (N6475, N5601, N3319);
xor XOR2 (N6476, N6473, N5358);
buf BUF1 (N6477, N6445);
and AND3 (N6478, N6476, N6387, N6177);
xor XOR2 (N6479, N6474, N5763);
not NOT1 (N6480, N6470);
nand NAND2 (N6481, N6451, N2406);
or OR3 (N6482, N6466, N6341, N5919);
or OR2 (N6483, N6482, N4023);
not NOT1 (N6484, N6475);
nor NOR2 (N6485, N6480, N1460);
xor XOR2 (N6486, N6478, N3248);
or OR2 (N6487, N6479, N604);
not NOT1 (N6488, N6477);
buf BUF1 (N6489, N6485);
or OR3 (N6490, N6481, N3521, N377);
nand NAND4 (N6491, N6458, N4901, N5653, N4352);
xor XOR2 (N6492, N6453, N5595);
xor XOR2 (N6493, N6487, N3122);
not NOT1 (N6494, N6491);
not NOT1 (N6495, N6484);
xor XOR2 (N6496, N6486, N113);
xor XOR2 (N6497, N6496, N2957);
nor NOR3 (N6498, N6497, N938, N4786);
or OR4 (N6499, N6489, N298, N2970, N2982);
xor XOR2 (N6500, N6498, N5396);
xor XOR2 (N6501, N6471, N5728);
or OR2 (N6502, N6499, N5125);
buf BUF1 (N6503, N6492);
nor NOR2 (N6504, N6483, N2630);
xor XOR2 (N6505, N6502, N2213);
xor XOR2 (N6506, N6503, N2306);
or OR4 (N6507, N6501, N5041, N209, N5705);
nor NOR3 (N6508, N6507, N3557, N2826);
xor XOR2 (N6509, N6500, N3814);
nor NOR2 (N6510, N6509, N550);
nor NOR4 (N6511, N6506, N4641, N5138, N756);
xor XOR2 (N6512, N6494, N6143);
not NOT1 (N6513, N6505);
or OR4 (N6514, N6504, N756, N3861, N1612);
buf BUF1 (N6515, N6495);
or OR2 (N6516, N6515, N2947);
nor NOR4 (N6517, N6490, N1771, N4706, N2300);
or OR4 (N6518, N6510, N729, N1633, N4530);
xor XOR2 (N6519, N6493, N3254);
xor XOR2 (N6520, N6488, N715);
and AND3 (N6521, N6519, N3554, N4569);
or OR3 (N6522, N6516, N4781, N4562);
buf BUF1 (N6523, N6514);
xor XOR2 (N6524, N6520, N291);
buf BUF1 (N6525, N6512);
or OR4 (N6526, N6523, N6018, N4756, N2475);
and AND3 (N6527, N6518, N2174, N2262);
nor NOR4 (N6528, N6527, N5898, N2102, N1229);
xor XOR2 (N6529, N6522, N4929);
nor NOR3 (N6530, N6526, N4607, N2247);
not NOT1 (N6531, N6521);
and AND3 (N6532, N6517, N2433, N3699);
or OR3 (N6533, N6513, N6261, N920);
nand NAND4 (N6534, N6531, N5805, N237, N4242);
not NOT1 (N6535, N6511);
xor XOR2 (N6536, N6535, N2782);
nor NOR3 (N6537, N6524, N3795, N4285);
and AND2 (N6538, N6532, N6379);
nand NAND2 (N6539, N6508, N6197);
buf BUF1 (N6540, N6534);
xor XOR2 (N6541, N6540, N5859);
and AND2 (N6542, N6536, N3172);
or OR3 (N6543, N6525, N6019, N2897);
buf BUF1 (N6544, N6541);
nor NOR4 (N6545, N6528, N3615, N4698, N3780);
or OR3 (N6546, N6529, N2157, N6415);
nor NOR4 (N6547, N6537, N6286, N4869, N3403);
not NOT1 (N6548, N6530);
and AND3 (N6549, N6543, N1836, N2348);
not NOT1 (N6550, N6542);
buf BUF1 (N6551, N6544);
and AND4 (N6552, N6545, N5082, N1748, N3140);
xor XOR2 (N6553, N6538, N3591);
and AND3 (N6554, N6547, N364, N410);
and AND3 (N6555, N6533, N1999, N32);
not NOT1 (N6556, N6549);
xor XOR2 (N6557, N6539, N1215);
buf BUF1 (N6558, N6551);
xor XOR2 (N6559, N6555, N1047);
nor NOR2 (N6560, N6556, N3715);
or OR3 (N6561, N6550, N5262, N370);
nor NOR2 (N6562, N6558, N1805);
and AND3 (N6563, N6561, N109, N5480);
xor XOR2 (N6564, N6554, N6390);
not NOT1 (N6565, N6553);
nor NOR2 (N6566, N6564, N1638);
or OR2 (N6567, N6565, N636);
xor XOR2 (N6568, N6560, N218);
not NOT1 (N6569, N6568);
xor XOR2 (N6570, N6563, N5);
nand NAND2 (N6571, N6567, N3111);
and AND2 (N6572, N6557, N4021);
nor NOR3 (N6573, N6546, N3726, N2927);
xor XOR2 (N6574, N6570, N415);
nand NAND4 (N6575, N6562, N614, N4842, N1230);
xor XOR2 (N6576, N6571, N6324);
buf BUF1 (N6577, N6573);
xor XOR2 (N6578, N6566, N5543);
not NOT1 (N6579, N6569);
not NOT1 (N6580, N6576);
and AND4 (N6581, N6572, N4727, N4052, N800);
nand NAND2 (N6582, N6578, N4239);
or OR3 (N6583, N6559, N5832, N1426);
not NOT1 (N6584, N6581);
nand NAND2 (N6585, N6579, N78);
or OR2 (N6586, N6583, N2004);
buf BUF1 (N6587, N6584);
buf BUF1 (N6588, N6582);
nand NAND3 (N6589, N6585, N3475, N2928);
buf BUF1 (N6590, N6588);
xor XOR2 (N6591, N6587, N4914);
or OR4 (N6592, N6580, N3489, N71, N6098);
nor NOR4 (N6593, N6591, N3274, N2948, N1297);
buf BUF1 (N6594, N6574);
nand NAND4 (N6595, N6589, N5579, N5293, N2353);
nor NOR3 (N6596, N6575, N6185, N5633);
not NOT1 (N6597, N6595);
not NOT1 (N6598, N6590);
not NOT1 (N6599, N6593);
and AND3 (N6600, N6577, N4456, N842);
and AND4 (N6601, N6596, N2141, N2594, N6036);
nand NAND3 (N6602, N6598, N6360, N5018);
and AND4 (N6603, N6594, N3903, N5016, N455);
xor XOR2 (N6604, N6586, N509);
xor XOR2 (N6605, N6552, N199);
and AND3 (N6606, N6605, N3620, N5880);
not NOT1 (N6607, N6597);
xor XOR2 (N6608, N6600, N2607);
nand NAND4 (N6609, N6601, N2392, N2832, N4628);
nand NAND4 (N6610, N6604, N4152, N3391, N106);
and AND2 (N6611, N6607, N2391);
not NOT1 (N6612, N6611);
and AND3 (N6613, N6602, N3421, N580);
nand NAND3 (N6614, N6606, N697, N4413);
nand NAND3 (N6615, N6592, N357, N6208);
not NOT1 (N6616, N6548);
or OR4 (N6617, N6615, N6175, N4184, N3498);
nand NAND3 (N6618, N6613, N1840, N773);
xor XOR2 (N6619, N6617, N5073);
not NOT1 (N6620, N6609);
nor NOR2 (N6621, N6612, N3467);
nor NOR4 (N6622, N6621, N1799, N6324, N3205);
nand NAND4 (N6623, N6622, N2582, N5819, N6583);
not NOT1 (N6624, N6610);
not NOT1 (N6625, N6608);
buf BUF1 (N6626, N6619);
nor NOR3 (N6627, N6623, N4268, N4190);
nor NOR3 (N6628, N6614, N5293, N1182);
nor NOR2 (N6629, N6616, N146);
nand NAND2 (N6630, N6628, N1282);
nor NOR4 (N6631, N6629, N3305, N1025, N143);
nor NOR2 (N6632, N6627, N4768);
buf BUF1 (N6633, N6631);
nand NAND4 (N6634, N6630, N5609, N506, N42);
nand NAND2 (N6635, N6603, N1510);
not NOT1 (N6636, N6632);
not NOT1 (N6637, N6626);
nor NOR2 (N6638, N6633, N764);
nand NAND4 (N6639, N6618, N3527, N715, N5278);
buf BUF1 (N6640, N6625);
nor NOR4 (N6641, N6634, N4762, N219, N124);
xor XOR2 (N6642, N6636, N441);
xor XOR2 (N6643, N6620, N1014);
xor XOR2 (N6644, N6640, N5206);
buf BUF1 (N6645, N6642);
nor NOR3 (N6646, N6635, N2382, N2247);
xor XOR2 (N6647, N6644, N2710);
nor NOR4 (N6648, N6638, N5841, N1068, N1228);
not NOT1 (N6649, N6624);
nor NOR2 (N6650, N6647, N1682);
or OR4 (N6651, N6639, N4078, N6077, N5154);
buf BUF1 (N6652, N6649);
not NOT1 (N6653, N6645);
and AND4 (N6654, N6641, N5233, N5232, N2872);
and AND4 (N6655, N6651, N5475, N1068, N2885);
or OR4 (N6656, N6648, N4660, N2686, N2569);
xor XOR2 (N6657, N6637, N6642);
xor XOR2 (N6658, N6653, N6041);
nand NAND2 (N6659, N6654, N26);
and AND3 (N6660, N6655, N2950, N6252);
or OR3 (N6661, N6652, N518, N2888);
not NOT1 (N6662, N6660);
or OR4 (N6663, N6650, N6065, N72, N6108);
nor NOR3 (N6664, N6643, N6529, N5432);
and AND2 (N6665, N6661, N983);
xor XOR2 (N6666, N6657, N4652);
nor NOR2 (N6667, N6646, N1730);
not NOT1 (N6668, N6599);
and AND2 (N6669, N6664, N285);
or OR4 (N6670, N6666, N4389, N4299, N3808);
xor XOR2 (N6671, N6663, N1065);
buf BUF1 (N6672, N6669);
buf BUF1 (N6673, N6656);
nor NOR4 (N6674, N6667, N1569, N3395, N1052);
nor NOR4 (N6675, N6674, N3378, N5407, N3749);
xor XOR2 (N6676, N6675, N1507);
buf BUF1 (N6677, N6668);
not NOT1 (N6678, N6673);
nor NOR2 (N6679, N6659, N1811);
xor XOR2 (N6680, N6658, N3130);
or OR3 (N6681, N6678, N6060, N1630);
not NOT1 (N6682, N6672);
xor XOR2 (N6683, N6671, N4925);
nor NOR4 (N6684, N6682, N3133, N2993, N6494);
xor XOR2 (N6685, N6680, N6122);
not NOT1 (N6686, N6681);
buf BUF1 (N6687, N6686);
buf BUF1 (N6688, N6679);
buf BUF1 (N6689, N6688);
or OR3 (N6690, N6687, N5686, N1829);
buf BUF1 (N6691, N6690);
and AND2 (N6692, N6665, N3805);
nor NOR2 (N6693, N6685, N1128);
and AND2 (N6694, N6693, N5577);
and AND4 (N6695, N6689, N5986, N753, N21);
nor NOR4 (N6696, N6677, N112, N3429, N5108);
and AND2 (N6697, N6696, N1418);
and AND3 (N6698, N6684, N3583, N6665);
not NOT1 (N6699, N6676);
not NOT1 (N6700, N6691);
nor NOR4 (N6701, N6670, N3556, N1747, N1844);
nand NAND2 (N6702, N6695, N6309);
nor NOR2 (N6703, N6702, N2510);
nand NAND2 (N6704, N6662, N327);
not NOT1 (N6705, N6683);
and AND2 (N6706, N6694, N2731);
and AND4 (N6707, N6705, N1685, N6275, N2214);
nor NOR3 (N6708, N6701, N3908, N4404);
buf BUF1 (N6709, N6704);
buf BUF1 (N6710, N6692);
nand NAND4 (N6711, N6706, N1151, N539, N5089);
xor XOR2 (N6712, N6703, N1099);
or OR4 (N6713, N6700, N1884, N4572, N5910);
nor NOR4 (N6714, N6707, N1133, N1917, N3376);
nand NAND4 (N6715, N6699, N2326, N76, N3753);
or OR3 (N6716, N6711, N1315, N323);
buf BUF1 (N6717, N6698);
buf BUF1 (N6718, N6697);
nor NOR3 (N6719, N6718, N4668, N5248);
xor XOR2 (N6720, N6713, N2350);
and AND4 (N6721, N6716, N3370, N2945, N5808);
nand NAND3 (N6722, N6720, N3820, N5515);
nand NAND2 (N6723, N6717, N2124);
nand NAND2 (N6724, N6709, N5582);
xor XOR2 (N6725, N6722, N1675);
and AND4 (N6726, N6715, N4867, N3035, N1856);
nand NAND4 (N6727, N6725, N2015, N2876, N1089);
not NOT1 (N6728, N6708);
nor NOR3 (N6729, N6727, N2946, N2516);
nor NOR4 (N6730, N6714, N394, N1294, N3627);
buf BUF1 (N6731, N6710);
or OR3 (N6732, N6728, N1647, N3729);
or OR3 (N6733, N6726, N2499, N2812);
buf BUF1 (N6734, N6721);
xor XOR2 (N6735, N6723, N5846);
or OR3 (N6736, N6729, N4562, N1298);
xor XOR2 (N6737, N6719, N345);
not NOT1 (N6738, N6735);
and AND2 (N6739, N6738, N5799);
or OR2 (N6740, N6724, N27);
or OR2 (N6741, N6733, N6049);
nand NAND2 (N6742, N6737, N4896);
xor XOR2 (N6743, N6712, N4849);
xor XOR2 (N6744, N6739, N1732);
buf BUF1 (N6745, N6734);
nand NAND2 (N6746, N6741, N4145);
and AND4 (N6747, N6746, N2785, N831, N5973);
and AND4 (N6748, N6742, N6116, N1033, N6697);
nor NOR2 (N6749, N6744, N5755);
nor NOR2 (N6750, N6731, N1774);
not NOT1 (N6751, N6749);
nor NOR3 (N6752, N6751, N2603, N5700);
or OR4 (N6753, N6732, N335, N652, N3292);
nand NAND4 (N6754, N6747, N4610, N3128, N5552);
nor NOR3 (N6755, N6745, N2441, N6531);
buf BUF1 (N6756, N6754);
or OR3 (N6757, N6752, N5014, N3912);
and AND2 (N6758, N6748, N2580);
not NOT1 (N6759, N6753);
buf BUF1 (N6760, N6759);
not NOT1 (N6761, N6736);
and AND3 (N6762, N6761, N590, N3046);
not NOT1 (N6763, N6750);
buf BUF1 (N6764, N6762);
nand NAND2 (N6765, N6758, N1850);
nand NAND2 (N6766, N6763, N1420);
xor XOR2 (N6767, N6756, N5037);
nor NOR3 (N6768, N6765, N1228, N3924);
not NOT1 (N6769, N6740);
nor NOR2 (N6770, N6743, N4207);
not NOT1 (N6771, N6768);
xor XOR2 (N6772, N6771, N3551);
xor XOR2 (N6773, N6757, N3428);
or OR2 (N6774, N6766, N704);
or OR2 (N6775, N6770, N1315);
and AND2 (N6776, N6760, N2551);
not NOT1 (N6777, N6776);
buf BUF1 (N6778, N6773);
not NOT1 (N6779, N6730);
xor XOR2 (N6780, N6772, N2332);
and AND4 (N6781, N6769, N4669, N6581, N5234);
xor XOR2 (N6782, N6777, N1489);
nor NOR3 (N6783, N6781, N2516, N4604);
not NOT1 (N6784, N6774);
xor XOR2 (N6785, N6780, N6340);
xor XOR2 (N6786, N6775, N6479);
and AND3 (N6787, N6785, N2727, N1391);
nand NAND3 (N6788, N6787, N3595, N2161);
nor NOR3 (N6789, N6764, N2979, N3);
xor XOR2 (N6790, N6783, N1059);
nor NOR4 (N6791, N6767, N3967, N5735, N6611);
not NOT1 (N6792, N6778);
not NOT1 (N6793, N6791);
nand NAND2 (N6794, N6782, N2911);
and AND4 (N6795, N6792, N2487, N430, N18);
nor NOR3 (N6796, N6779, N2376, N4974);
nand NAND3 (N6797, N6793, N5649, N1218);
and AND2 (N6798, N6796, N1707);
not NOT1 (N6799, N6755);
xor XOR2 (N6800, N6797, N2202);
buf BUF1 (N6801, N6800);
nand NAND3 (N6802, N6801, N1193, N5419);
not NOT1 (N6803, N6789);
not NOT1 (N6804, N6802);
and AND3 (N6805, N6786, N374, N1971);
and AND4 (N6806, N6795, N4852, N3210, N621);
and AND4 (N6807, N6799, N4138, N6492, N2063);
xor XOR2 (N6808, N6803, N5973);
and AND4 (N6809, N6805, N5849, N3636, N4378);
and AND4 (N6810, N6809, N5991, N1252, N3724);
nor NOR2 (N6811, N6807, N4377);
nand NAND2 (N6812, N6794, N6324);
nor NOR2 (N6813, N6810, N4832);
nor NOR2 (N6814, N6811, N6257);
not NOT1 (N6815, N6784);
not NOT1 (N6816, N6812);
or OR4 (N6817, N6788, N5112, N2491, N4494);
nor NOR2 (N6818, N6814, N1481);
xor XOR2 (N6819, N6808, N2832);
and AND2 (N6820, N6817, N4694);
or OR4 (N6821, N6790, N6114, N3708, N1834);
and AND2 (N6822, N6820, N2629);
and AND4 (N6823, N6813, N3469, N4919, N707);
and AND2 (N6824, N6798, N69);
or OR3 (N6825, N6818, N1781, N5209);
nand NAND3 (N6826, N6806, N1086, N4364);
or OR2 (N6827, N6819, N1390);
nor NOR3 (N6828, N6825, N1534, N14);
nor NOR3 (N6829, N6816, N5421, N591);
or OR2 (N6830, N6824, N4486);
buf BUF1 (N6831, N6830);
nor NOR3 (N6832, N6822, N3452, N3223);
nand NAND2 (N6833, N6829, N5609);
nand NAND2 (N6834, N6833, N619);
not NOT1 (N6835, N6831);
buf BUF1 (N6836, N6834);
xor XOR2 (N6837, N6815, N57);
xor XOR2 (N6838, N6836, N3586);
buf BUF1 (N6839, N6804);
xor XOR2 (N6840, N6838, N4638);
and AND2 (N6841, N6827, N2571);
buf BUF1 (N6842, N6821);
not NOT1 (N6843, N6823);
xor XOR2 (N6844, N6835, N6674);
xor XOR2 (N6845, N6837, N6580);
nor NOR3 (N6846, N6841, N5822, N4168);
xor XOR2 (N6847, N6839, N512);
nor NOR4 (N6848, N6832, N844, N5605, N4011);
nand NAND4 (N6849, N6843, N3817, N5887, N5317);
not NOT1 (N6850, N6847);
xor XOR2 (N6851, N6846, N6231);
and AND3 (N6852, N6844, N4058, N3705);
not NOT1 (N6853, N6851);
or OR3 (N6854, N6848, N134, N5498);
not NOT1 (N6855, N6849);
and AND4 (N6856, N6826, N2496, N1836, N5657);
buf BUF1 (N6857, N6842);
or OR2 (N6858, N6828, N5363);
or OR4 (N6859, N6852, N161, N2143, N1907);
buf BUF1 (N6860, N6859);
not NOT1 (N6861, N6860);
and AND4 (N6862, N6857, N3849, N5222, N2443);
xor XOR2 (N6863, N6856, N5684);
or OR3 (N6864, N6858, N912, N75);
xor XOR2 (N6865, N6861, N749);
or OR4 (N6866, N6855, N5700, N3067, N1785);
nand NAND2 (N6867, N6865, N3801);
or OR3 (N6868, N6845, N3044, N1157);
not NOT1 (N6869, N6854);
not NOT1 (N6870, N6863);
nand NAND4 (N6871, N6867, N1343, N6150, N6819);
not NOT1 (N6872, N6868);
nor NOR4 (N6873, N6869, N6332, N2767, N3828);
and AND3 (N6874, N6871, N6292, N5007);
and AND2 (N6875, N6862, N6781);
nand NAND4 (N6876, N6866, N4559, N6646, N1916);
nand NAND4 (N6877, N6850, N6613, N4476, N462);
or OR3 (N6878, N6872, N5721, N5027);
nand NAND3 (N6879, N6876, N5422, N474);
buf BUF1 (N6880, N6840);
and AND3 (N6881, N6875, N689, N3559);
buf BUF1 (N6882, N6880);
and AND3 (N6883, N6877, N2532, N4887);
buf BUF1 (N6884, N6874);
and AND3 (N6885, N6873, N3281, N3119);
not NOT1 (N6886, N6882);
and AND4 (N6887, N6881, N3096, N1034, N4070);
and AND2 (N6888, N6885, N3296);
nand NAND3 (N6889, N6886, N3269, N5257);
or OR4 (N6890, N6889, N3042, N1683, N3876);
buf BUF1 (N6891, N6878);
and AND4 (N6892, N6883, N6865, N714, N2903);
xor XOR2 (N6893, N6892, N11);
nand NAND2 (N6894, N6870, N5948);
xor XOR2 (N6895, N6891, N6772);
buf BUF1 (N6896, N6890);
buf BUF1 (N6897, N6888);
and AND2 (N6898, N6893, N5672);
buf BUF1 (N6899, N6897);
and AND2 (N6900, N6879, N6631);
nor NOR3 (N6901, N6887, N5784, N2274);
buf BUF1 (N6902, N6900);
not NOT1 (N6903, N6864);
xor XOR2 (N6904, N6895, N2990);
and AND4 (N6905, N6902, N3916, N4163, N3420);
buf BUF1 (N6906, N6904);
nor NOR2 (N6907, N6894, N1250);
buf BUF1 (N6908, N6905);
nand NAND4 (N6909, N6901, N157, N5243, N3493);
buf BUF1 (N6910, N6903);
nand NAND3 (N6911, N6906, N2129, N504);
nand NAND3 (N6912, N6911, N6319, N412);
and AND2 (N6913, N6898, N5543);
not NOT1 (N6914, N6910);
and AND2 (N6915, N6908, N4734);
xor XOR2 (N6916, N6915, N6598);
buf BUF1 (N6917, N6909);
xor XOR2 (N6918, N6899, N22);
not NOT1 (N6919, N6884);
nor NOR2 (N6920, N6916, N295);
or OR2 (N6921, N6913, N1459);
nor NOR3 (N6922, N6914, N6866, N2265);
nor NOR4 (N6923, N6918, N3480, N6175, N4298);
nand NAND3 (N6924, N6919, N5264, N337);
not NOT1 (N6925, N6907);
nand NAND3 (N6926, N6920, N4607, N2068);
xor XOR2 (N6927, N6912, N4053);
or OR3 (N6928, N6925, N841, N1694);
or OR4 (N6929, N6921, N4213, N252, N6587);
not NOT1 (N6930, N6929);
buf BUF1 (N6931, N6923);
nand NAND2 (N6932, N6926, N1690);
and AND2 (N6933, N6928, N6858);
not NOT1 (N6934, N6927);
nor NOR3 (N6935, N6934, N42, N4846);
nor NOR4 (N6936, N6933, N3732, N979, N5826);
buf BUF1 (N6937, N6924);
or OR2 (N6938, N6932, N2858);
nor NOR3 (N6939, N6938, N4947, N79);
xor XOR2 (N6940, N6853, N1045);
nor NOR2 (N6941, N6930, N4481);
nor NOR3 (N6942, N6939, N1918, N2106);
nand NAND4 (N6943, N6896, N5815, N1454, N4873);
and AND2 (N6944, N6931, N2440);
or OR2 (N6945, N6917, N5912);
or OR2 (N6946, N6940, N6430);
and AND3 (N6947, N6942, N4907, N6042);
or OR2 (N6948, N6922, N1608);
nand NAND2 (N6949, N6935, N4869);
buf BUF1 (N6950, N6945);
nand NAND4 (N6951, N6946, N1666, N5895, N1294);
nand NAND2 (N6952, N6944, N2222);
nor NOR4 (N6953, N6952, N1353, N1757, N4766);
nor NOR4 (N6954, N6936, N6616, N2681, N33);
xor XOR2 (N6955, N6949, N1865);
nor NOR2 (N6956, N6955, N2337);
nor NOR3 (N6957, N6941, N5649, N2477);
nand NAND3 (N6958, N6957, N4213, N1082);
and AND3 (N6959, N6950, N4656, N6401);
or OR3 (N6960, N6943, N2591, N1166);
nand NAND2 (N6961, N6954, N3978);
nor NOR2 (N6962, N6953, N333);
nand NAND2 (N6963, N6962, N5909);
xor XOR2 (N6964, N6961, N6083);
nand NAND3 (N6965, N6964, N5274, N2503);
and AND4 (N6966, N6948, N1255, N2895, N3483);
or OR3 (N6967, N6951, N4985, N5755);
xor XOR2 (N6968, N6956, N3195);
buf BUF1 (N6969, N6966);
buf BUF1 (N6970, N6967);
and AND4 (N6971, N6958, N3938, N5059, N212);
xor XOR2 (N6972, N6969, N5910);
xor XOR2 (N6973, N6937, N1622);
and AND4 (N6974, N6947, N180, N2436, N1402);
not NOT1 (N6975, N6968);
buf BUF1 (N6976, N6960);
xor XOR2 (N6977, N6971, N3495);
and AND3 (N6978, N6974, N4965, N2479);
or OR2 (N6979, N6973, N6523);
nand NAND2 (N6980, N6975, N5772);
and AND4 (N6981, N6977, N2924, N937, N5116);
not NOT1 (N6982, N6972);
and AND4 (N6983, N6981, N585, N3872, N4150);
and AND3 (N6984, N6982, N740, N5383);
nor NOR2 (N6985, N6983, N4682);
buf BUF1 (N6986, N6980);
nand NAND4 (N6987, N6985, N1331, N838, N5646);
buf BUF1 (N6988, N6976);
nand NAND3 (N6989, N6970, N4190, N781);
and AND2 (N6990, N6986, N455);
xor XOR2 (N6991, N6959, N387);
and AND4 (N6992, N6965, N5401, N2903, N2521);
buf BUF1 (N6993, N6990);
not NOT1 (N6994, N6992);
or OR2 (N6995, N6994, N6419);
and AND3 (N6996, N6978, N5178, N1484);
buf BUF1 (N6997, N6989);
or OR4 (N6998, N6995, N2763, N36, N137);
xor XOR2 (N6999, N6993, N2374);
buf BUF1 (N7000, N6991);
or OR3 (N7001, N6997, N5566, N5173);
buf BUF1 (N7002, N6998);
nor NOR4 (N7003, N6963, N2062, N3435, N1669);
nor NOR3 (N7004, N6984, N3162, N4001);
xor XOR2 (N7005, N6988, N4985);
buf BUF1 (N7006, N6996);
or OR4 (N7007, N6999, N2121, N493, N1101);
and AND3 (N7008, N7007, N6078, N3212);
or OR4 (N7009, N6979, N4317, N6531, N4560);
or OR4 (N7010, N7001, N2295, N6430, N199);
or OR3 (N7011, N7004, N522, N6053);
nand NAND3 (N7012, N7011, N3250, N3961);
xor XOR2 (N7013, N7006, N2884);
buf BUF1 (N7014, N7002);
and AND3 (N7015, N7013, N4036, N1536);
not NOT1 (N7016, N7003);
nor NOR2 (N7017, N7016, N1739);
or OR2 (N7018, N7000, N5016);
or OR3 (N7019, N7018, N3299, N5553);
or OR4 (N7020, N7017, N6448, N2249, N376);
or OR4 (N7021, N7019, N2220, N1009, N4620);
nor NOR4 (N7022, N7021, N745, N2009, N5793);
nand NAND2 (N7023, N7008, N6515);
nand NAND2 (N7024, N7022, N4786);
nand NAND2 (N7025, N7015, N6599);
not NOT1 (N7026, N7023);
nand NAND2 (N7027, N7012, N5959);
or OR4 (N7028, N7026, N1796, N6446, N2609);
nor NOR2 (N7029, N7025, N3715);
nand NAND2 (N7030, N7009, N6041);
nand NAND4 (N7031, N7024, N6758, N4276, N436);
nand NAND3 (N7032, N6987, N6060, N4031);
xor XOR2 (N7033, N7029, N4004);
xor XOR2 (N7034, N7014, N6561);
xor XOR2 (N7035, N7030, N1443);
or OR2 (N7036, N7034, N74);
not NOT1 (N7037, N7005);
not NOT1 (N7038, N7036);
xor XOR2 (N7039, N7038, N6427);
not NOT1 (N7040, N7035);
nand NAND4 (N7041, N7031, N1030, N4765, N4077);
nand NAND3 (N7042, N7040, N6200, N1232);
nor NOR2 (N7043, N7037, N3123);
and AND4 (N7044, N7033, N5794, N4047, N3577);
nand NAND3 (N7045, N7043, N7015, N290);
or OR4 (N7046, N7032, N6009, N5046, N6153);
or OR2 (N7047, N7042, N2655);
and AND2 (N7048, N7047, N1611);
xor XOR2 (N7049, N7027, N4492);
nor NOR4 (N7050, N7044, N6136, N6575, N6540);
nor NOR2 (N7051, N7039, N2884);
or OR2 (N7052, N7048, N3705);
nand NAND4 (N7053, N7020, N2578, N4686, N1408);
nor NOR3 (N7054, N7010, N6093, N2011);
not NOT1 (N7055, N7050);
nand NAND4 (N7056, N7045, N6873, N823, N3567);
not NOT1 (N7057, N7054);
xor XOR2 (N7058, N7057, N5336);
nand NAND2 (N7059, N7049, N1845);
buf BUF1 (N7060, N7053);
or OR4 (N7061, N7055, N5574, N2856, N4511);
or OR4 (N7062, N7046, N1808, N1646, N4582);
not NOT1 (N7063, N7060);
not NOT1 (N7064, N7051);
or OR3 (N7065, N7062, N7055, N4492);
nand NAND3 (N7066, N7058, N5531, N4105);
nor NOR3 (N7067, N7041, N6032, N1685);
buf BUF1 (N7068, N7061);
or OR4 (N7069, N7063, N3184, N3981, N2925);
and AND2 (N7070, N7056, N5632);
buf BUF1 (N7071, N7052);
nor NOR3 (N7072, N7066, N2821, N6492);
not NOT1 (N7073, N7070);
or OR4 (N7074, N7068, N5130, N4476, N6190);
or OR2 (N7075, N7071, N2106);
nand NAND4 (N7076, N7069, N1924, N3897, N4869);
xor XOR2 (N7077, N7065, N581);
and AND2 (N7078, N7075, N4154);
xor XOR2 (N7079, N7074, N4554);
xor XOR2 (N7080, N7076, N711);
and AND3 (N7081, N7072, N5788, N6343);
nor NOR2 (N7082, N7079, N1338);
and AND4 (N7083, N7073, N1107, N2909, N3625);
nor NOR2 (N7084, N7064, N3158);
nand NAND3 (N7085, N7028, N6741, N450);
not NOT1 (N7086, N7081);
buf BUF1 (N7087, N7082);
and AND3 (N7088, N7077, N215, N3607);
buf BUF1 (N7089, N7085);
or OR3 (N7090, N7067, N856, N5645);
xor XOR2 (N7091, N7083, N1850);
xor XOR2 (N7092, N7086, N5308);
nor NOR3 (N7093, N7091, N4923, N5767);
buf BUF1 (N7094, N7089);
nand NAND3 (N7095, N7092, N3870, N4401);
buf BUF1 (N7096, N7080);
xor XOR2 (N7097, N7078, N5199);
nor NOR4 (N7098, N7084, N1894, N2137, N6170);
or OR2 (N7099, N7090, N675);
and AND2 (N7100, N7096, N3688);
buf BUF1 (N7101, N7094);
buf BUF1 (N7102, N7059);
and AND4 (N7103, N7098, N6488, N6299, N417);
or OR2 (N7104, N7099, N343);
xor XOR2 (N7105, N7093, N1091);
buf BUF1 (N7106, N7088);
nand NAND4 (N7107, N7104, N3994, N3806, N5855);
buf BUF1 (N7108, N7107);
and AND2 (N7109, N7101, N4669);
not NOT1 (N7110, N7105);
nor NOR3 (N7111, N7106, N900, N2231);
xor XOR2 (N7112, N7111, N3861);
and AND3 (N7113, N7100, N1398, N6206);
xor XOR2 (N7114, N7109, N373);
xor XOR2 (N7115, N7087, N4624);
not NOT1 (N7116, N7103);
xor XOR2 (N7117, N7110, N4322);
or OR2 (N7118, N7114, N2621);
nor NOR3 (N7119, N7113, N4824, N2812);
nor NOR4 (N7120, N7119, N557, N7071, N1097);
nor NOR4 (N7121, N7118, N5514, N6851, N6610);
not NOT1 (N7122, N7112);
and AND4 (N7123, N7095, N582, N1172, N3208);
xor XOR2 (N7124, N7108, N4581);
not NOT1 (N7125, N7116);
buf BUF1 (N7126, N7123);
nor NOR3 (N7127, N7117, N5696, N5790);
not NOT1 (N7128, N7124);
xor XOR2 (N7129, N7128, N685);
buf BUF1 (N7130, N7115);
or OR3 (N7131, N7121, N5488, N3721);
nand NAND4 (N7132, N7126, N1037, N5873, N4554);
not NOT1 (N7133, N7122);
xor XOR2 (N7134, N7127, N5206);
xor XOR2 (N7135, N7102, N2278);
or OR3 (N7136, N7134, N1544, N1461);
and AND4 (N7137, N7131, N633, N6277, N4720);
buf BUF1 (N7138, N7133);
nor NOR3 (N7139, N7125, N5138, N4324);
xor XOR2 (N7140, N7132, N2472);
xor XOR2 (N7141, N7139, N1285);
xor XOR2 (N7142, N7138, N5367);
xor XOR2 (N7143, N7141, N4703);
and AND3 (N7144, N7129, N6066, N3196);
buf BUF1 (N7145, N7140);
buf BUF1 (N7146, N7137);
not NOT1 (N7147, N7136);
nor NOR4 (N7148, N7146, N1853, N595, N584);
nand NAND3 (N7149, N7120, N6826, N5666);
or OR3 (N7150, N7145, N3241, N2616);
buf BUF1 (N7151, N7097);
buf BUF1 (N7152, N7149);
or OR3 (N7153, N7148, N3839, N1983);
nand NAND2 (N7154, N7147, N3458);
and AND3 (N7155, N7152, N391, N3380);
or OR4 (N7156, N7150, N4133, N6896, N1694);
nand NAND4 (N7157, N7153, N1236, N1052, N6521);
buf BUF1 (N7158, N7144);
buf BUF1 (N7159, N7157);
nand NAND2 (N7160, N7130, N6929);
nor NOR4 (N7161, N7159, N7110, N985, N5956);
xor XOR2 (N7162, N7161, N4165);
or OR2 (N7163, N7158, N7060);
nor NOR2 (N7164, N7155, N6499);
nor NOR4 (N7165, N7143, N4013, N3214, N6381);
and AND4 (N7166, N7160, N6161, N3363, N6687);
xor XOR2 (N7167, N7164, N3434);
xor XOR2 (N7168, N7135, N4341);
nor NOR4 (N7169, N7163, N5091, N5633, N118);
nor NOR3 (N7170, N7167, N5349, N334);
or OR4 (N7171, N7151, N719, N6435, N6006);
buf BUF1 (N7172, N7166);
and AND2 (N7173, N7169, N2553);
and AND2 (N7174, N7170, N2665);
not NOT1 (N7175, N7174);
nand NAND3 (N7176, N7173, N3126, N3698);
not NOT1 (N7177, N7162);
xor XOR2 (N7178, N7168, N566);
or OR3 (N7179, N7142, N4715, N5712);
nor NOR3 (N7180, N7172, N3517, N577);
xor XOR2 (N7181, N7154, N3179);
nand NAND3 (N7182, N7181, N497, N2923);
buf BUF1 (N7183, N7177);
not NOT1 (N7184, N7175);
xor XOR2 (N7185, N7184, N6603);
and AND3 (N7186, N7165, N4375, N3739);
or OR3 (N7187, N7186, N3622, N5102);
nor NOR4 (N7188, N7171, N105, N5701, N6490);
nor NOR4 (N7189, N7188, N7088, N5355, N1889);
or OR2 (N7190, N7185, N149);
buf BUF1 (N7191, N7176);
nand NAND2 (N7192, N7187, N295);
xor XOR2 (N7193, N7178, N615);
and AND3 (N7194, N7190, N4893, N4694);
or OR4 (N7195, N7183, N2297, N3009, N1740);
and AND3 (N7196, N7192, N390, N1415);
not NOT1 (N7197, N7182);
nand NAND4 (N7198, N7195, N4123, N4912, N1355);
nand NAND4 (N7199, N7189, N3729, N1359, N4434);
or OR2 (N7200, N7191, N835);
xor XOR2 (N7201, N7179, N968);
nand NAND4 (N7202, N7197, N1130, N6031, N5565);
not NOT1 (N7203, N7202);
not NOT1 (N7204, N7199);
or OR4 (N7205, N7204, N3772, N1891, N5056);
not NOT1 (N7206, N7156);
buf BUF1 (N7207, N7180);
xor XOR2 (N7208, N7198, N1328);
nand NAND3 (N7209, N7194, N6059, N4951);
xor XOR2 (N7210, N7205, N5754);
not NOT1 (N7211, N7208);
or OR3 (N7212, N7209, N5755, N5273);
or OR2 (N7213, N7212, N4933);
not NOT1 (N7214, N7201);
nor NOR3 (N7215, N7207, N6616, N1897);
xor XOR2 (N7216, N7206, N6992);
xor XOR2 (N7217, N7216, N4802);
xor XOR2 (N7218, N7196, N6848);
or OR3 (N7219, N7193, N1278, N705);
and AND4 (N7220, N7214, N5897, N3143, N6553);
or OR3 (N7221, N7211, N3806, N837);
or OR4 (N7222, N7213, N2356, N5909, N4271);
and AND2 (N7223, N7210, N4802);
buf BUF1 (N7224, N7200);
not NOT1 (N7225, N7215);
nand NAND2 (N7226, N7222, N6692);
or OR4 (N7227, N7221, N3072, N1930, N355);
nor NOR2 (N7228, N7226, N3115);
xor XOR2 (N7229, N7203, N3875);
buf BUF1 (N7230, N7228);
and AND4 (N7231, N7218, N3011, N1792, N2548);
xor XOR2 (N7232, N7217, N5764);
nand NAND4 (N7233, N7220, N1696, N737, N5725);
buf BUF1 (N7234, N7231);
buf BUF1 (N7235, N7232);
not NOT1 (N7236, N7225);
xor XOR2 (N7237, N7233, N3740);
xor XOR2 (N7238, N7227, N3249);
and AND4 (N7239, N7235, N6856, N1760, N1535);
buf BUF1 (N7240, N7237);
xor XOR2 (N7241, N7229, N1846);
nor NOR3 (N7242, N7240, N5488, N2452);
or OR4 (N7243, N7230, N5567, N1587, N5167);
nand NAND4 (N7244, N7243, N6290, N5619, N3814);
not NOT1 (N7245, N7242);
nor NOR4 (N7246, N7224, N2554, N5733, N266);
and AND2 (N7247, N7223, N3823);
buf BUF1 (N7248, N7234);
nand NAND3 (N7249, N7244, N3351, N5017);
buf BUF1 (N7250, N7247);
nand NAND2 (N7251, N7245, N7194);
buf BUF1 (N7252, N7239);
not NOT1 (N7253, N7248);
and AND2 (N7254, N7253, N5844);
nand NAND2 (N7255, N7219, N1963);
nand NAND3 (N7256, N7250, N6698, N3844);
xor XOR2 (N7257, N7252, N1424);
buf BUF1 (N7258, N7238);
nor NOR4 (N7259, N7251, N2702, N4394, N3528);
xor XOR2 (N7260, N7257, N5501);
buf BUF1 (N7261, N7254);
xor XOR2 (N7262, N7258, N7013);
nor NOR4 (N7263, N7246, N255, N5796, N5372);
xor XOR2 (N7264, N7236, N7071);
nand NAND2 (N7265, N7263, N270);
buf BUF1 (N7266, N7261);
not NOT1 (N7267, N7256);
or OR2 (N7268, N7267, N456);
buf BUF1 (N7269, N7255);
and AND2 (N7270, N7249, N6761);
and AND2 (N7271, N7241, N3207);
and AND4 (N7272, N7264, N1838, N8, N6446);
and AND4 (N7273, N7272, N3217, N1456, N6150);
and AND2 (N7274, N7260, N2255);
nor NOR3 (N7275, N7266, N5200, N3440);
not NOT1 (N7276, N7262);
not NOT1 (N7277, N7270);
not NOT1 (N7278, N7276);
nand NAND3 (N7279, N7278, N5466, N3008);
buf BUF1 (N7280, N7277);
buf BUF1 (N7281, N7279);
xor XOR2 (N7282, N7274, N6585);
buf BUF1 (N7283, N7269);
nand NAND3 (N7284, N7275, N80, N3257);
not NOT1 (N7285, N7281);
nand NAND2 (N7286, N7259, N2198);
not NOT1 (N7287, N7273);
not NOT1 (N7288, N7280);
buf BUF1 (N7289, N7265);
not NOT1 (N7290, N7282);
nor NOR4 (N7291, N7289, N5337, N3911, N3915);
nand NAND3 (N7292, N7284, N928, N6271);
buf BUF1 (N7293, N7288);
and AND3 (N7294, N7287, N874, N2114);
buf BUF1 (N7295, N7293);
xor XOR2 (N7296, N7294, N4452);
not NOT1 (N7297, N7295);
not NOT1 (N7298, N7291);
buf BUF1 (N7299, N7283);
nand NAND4 (N7300, N7297, N2687, N3863, N3874);
nor NOR4 (N7301, N7299, N6324, N3520, N3237);
not NOT1 (N7302, N7268);
not NOT1 (N7303, N7298);
nand NAND3 (N7304, N7300, N2228, N3996);
buf BUF1 (N7305, N7271);
or OR2 (N7306, N7301, N6671);
xor XOR2 (N7307, N7285, N6255);
and AND3 (N7308, N7304, N4670, N357);
and AND2 (N7309, N7302, N4670);
not NOT1 (N7310, N7303);
xor XOR2 (N7311, N7290, N2294);
nor NOR4 (N7312, N7308, N5785, N2373, N797);
buf BUF1 (N7313, N7292);
nand NAND2 (N7314, N7313, N2435);
or OR4 (N7315, N7312, N6020, N2265, N619);
buf BUF1 (N7316, N7310);
nor NOR4 (N7317, N7306, N1859, N3391, N4288);
not NOT1 (N7318, N7314);
not NOT1 (N7319, N7296);
or OR2 (N7320, N7309, N6326);
xor XOR2 (N7321, N7315, N4563);
and AND4 (N7322, N7316, N2625, N4005, N2276);
or OR4 (N7323, N7321, N4810, N4971, N4450);
and AND4 (N7324, N7307, N4451, N5999, N2565);
nand NAND4 (N7325, N7324, N4025, N2358, N2175);
and AND3 (N7326, N7318, N5346, N5880);
nand NAND2 (N7327, N7325, N5117);
or OR2 (N7328, N7286, N5952);
nor NOR2 (N7329, N7327, N137);
xor XOR2 (N7330, N7319, N2018);
and AND2 (N7331, N7311, N745);
and AND3 (N7332, N7317, N6619, N1151);
or OR3 (N7333, N7305, N2156, N6374);
not NOT1 (N7334, N7333);
nor NOR3 (N7335, N7331, N6374, N3767);
nor NOR2 (N7336, N7330, N2558);
buf BUF1 (N7337, N7334);
or OR3 (N7338, N7326, N688, N5346);
buf BUF1 (N7339, N7320);
or OR2 (N7340, N7329, N2161);
nand NAND2 (N7341, N7337, N5291);
nor NOR4 (N7342, N7341, N6815, N5511, N6206);
nor NOR4 (N7343, N7339, N2837, N2279, N5388);
xor XOR2 (N7344, N7328, N862);
xor XOR2 (N7345, N7342, N1793);
nand NAND4 (N7346, N7322, N6943, N4122, N3542);
buf BUF1 (N7347, N7335);
buf BUF1 (N7348, N7347);
nor NOR4 (N7349, N7344, N525, N3112, N4838);
or OR4 (N7350, N7332, N3573, N7223, N4537);
not NOT1 (N7351, N7343);
or OR2 (N7352, N7348, N1444);
and AND4 (N7353, N7340, N2577, N3716, N1134);
or OR3 (N7354, N7346, N6705, N4734);
xor XOR2 (N7355, N7353, N7140);
nand NAND2 (N7356, N7338, N2990);
and AND3 (N7357, N7336, N1662, N6076);
not NOT1 (N7358, N7351);
nor NOR2 (N7359, N7357, N1712);
nor NOR2 (N7360, N7349, N6306);
and AND3 (N7361, N7350, N856, N6867);
nor NOR4 (N7362, N7354, N5192, N6192, N6658);
nand NAND4 (N7363, N7345, N6358, N4669, N6122);
nand NAND3 (N7364, N7360, N2450, N3159);
not NOT1 (N7365, N7362);
nor NOR2 (N7366, N7358, N1259);
and AND3 (N7367, N7364, N2019, N2287);
nor NOR3 (N7368, N7355, N72, N1294);
buf BUF1 (N7369, N7352);
xor XOR2 (N7370, N7368, N1036);
and AND3 (N7371, N7323, N5732, N867);
or OR3 (N7372, N7367, N5112, N4054);
not NOT1 (N7373, N7369);
xor XOR2 (N7374, N7365, N7269);
nor NOR3 (N7375, N7366, N5493, N6394);
not NOT1 (N7376, N7363);
nor NOR4 (N7377, N7370, N1816, N5301, N459);
buf BUF1 (N7378, N7372);
xor XOR2 (N7379, N7376, N6706);
and AND2 (N7380, N7361, N5590);
nor NOR4 (N7381, N7356, N3487, N6608, N5601);
xor XOR2 (N7382, N7380, N5845);
nand NAND2 (N7383, N7374, N3921);
nand NAND4 (N7384, N7378, N71, N4926, N6221);
nand NAND2 (N7385, N7379, N375);
nor NOR2 (N7386, N7383, N2463);
and AND3 (N7387, N7373, N5884, N6337);
or OR2 (N7388, N7384, N5949);
xor XOR2 (N7389, N7385, N6712);
nor NOR3 (N7390, N7375, N818, N6571);
xor XOR2 (N7391, N7387, N4003);
nand NAND3 (N7392, N7389, N4721, N1798);
xor XOR2 (N7393, N7388, N3552);
buf BUF1 (N7394, N7386);
xor XOR2 (N7395, N7377, N7131);
nor NOR4 (N7396, N7371, N5999, N5378, N3804);
not NOT1 (N7397, N7390);
not NOT1 (N7398, N7393);
nand NAND4 (N7399, N7397, N1373, N639, N2836);
or OR3 (N7400, N7394, N3671, N5448);
buf BUF1 (N7401, N7395);
nor NOR2 (N7402, N7382, N359);
not NOT1 (N7403, N7359);
buf BUF1 (N7404, N7398);
buf BUF1 (N7405, N7399);
nor NOR2 (N7406, N7403, N372);
and AND4 (N7407, N7381, N5037, N6795, N3618);
nor NOR3 (N7408, N7405, N3960, N6033);
not NOT1 (N7409, N7408);
buf BUF1 (N7410, N7404);
not NOT1 (N7411, N7407);
buf BUF1 (N7412, N7400);
buf BUF1 (N7413, N7410);
nor NOR2 (N7414, N7396, N3425);
and AND4 (N7415, N7411, N2258, N1201, N6538);
nand NAND2 (N7416, N7402, N7232);
nand NAND4 (N7417, N7409, N1319, N3180, N5205);
nand NAND2 (N7418, N7416, N467);
buf BUF1 (N7419, N7413);
nor NOR2 (N7420, N7392, N2590);
not NOT1 (N7421, N7415);
and AND2 (N7422, N7420, N2981);
buf BUF1 (N7423, N7391);
and AND2 (N7424, N7401, N6796);
nor NOR3 (N7425, N7414, N3850, N282);
buf BUF1 (N7426, N7424);
nand NAND3 (N7427, N7425, N1039, N349);
xor XOR2 (N7428, N7406, N1520);
nor NOR4 (N7429, N7422, N7402, N3072, N6061);
xor XOR2 (N7430, N7428, N121);
nor NOR4 (N7431, N7421, N4817, N1663, N2706);
and AND2 (N7432, N7412, N3161);
buf BUF1 (N7433, N7418);
not NOT1 (N7434, N7419);
buf BUF1 (N7435, N7431);
not NOT1 (N7436, N7429);
or OR2 (N7437, N7427, N3430);
buf BUF1 (N7438, N7435);
not NOT1 (N7439, N7430);
and AND4 (N7440, N7432, N4486, N5260, N3848);
xor XOR2 (N7441, N7434, N6517);
and AND2 (N7442, N7426, N6410);
xor XOR2 (N7443, N7438, N435);
and AND2 (N7444, N7433, N5372);
xor XOR2 (N7445, N7442, N2825);
not NOT1 (N7446, N7443);
xor XOR2 (N7447, N7439, N3904);
buf BUF1 (N7448, N7444);
not NOT1 (N7449, N7436);
nand NAND2 (N7450, N7440, N5784);
buf BUF1 (N7451, N7445);
nand NAND4 (N7452, N7441, N1863, N4110, N4608);
nand NAND4 (N7453, N7423, N5686, N5597, N65);
and AND2 (N7454, N7452, N1227);
buf BUF1 (N7455, N7454);
not NOT1 (N7456, N7446);
buf BUF1 (N7457, N7455);
nand NAND2 (N7458, N7417, N6957);
nand NAND4 (N7459, N7437, N6888, N6899, N5388);
xor XOR2 (N7460, N7449, N3423);
nand NAND2 (N7461, N7460, N6666);
and AND4 (N7462, N7457, N7216, N1392, N297);
nor NOR4 (N7463, N7450, N3046, N2436, N147);
nor NOR4 (N7464, N7462, N6319, N1968, N3431);
buf BUF1 (N7465, N7453);
xor XOR2 (N7466, N7458, N2320);
or OR3 (N7467, N7448, N5609, N6535);
and AND3 (N7468, N7466, N5185, N794);
or OR4 (N7469, N7468, N6718, N605, N6559);
or OR2 (N7470, N7459, N1573);
nand NAND3 (N7471, N7461, N458, N4270);
nor NOR4 (N7472, N7469, N6238, N2027, N2449);
and AND2 (N7473, N7464, N3700);
and AND3 (N7474, N7456, N2469, N1819);
xor XOR2 (N7475, N7472, N3728);
nand NAND2 (N7476, N7465, N2640);
nand NAND2 (N7477, N7471, N3462);
or OR3 (N7478, N7470, N5634, N7404);
xor XOR2 (N7479, N7475, N2075);
and AND3 (N7480, N7476, N4034, N561);
or OR3 (N7481, N7463, N5852, N4053);
xor XOR2 (N7482, N7447, N6941);
nand NAND4 (N7483, N7480, N2958, N69, N5084);
or OR3 (N7484, N7478, N5555, N6314);
xor XOR2 (N7485, N7483, N478);
buf BUF1 (N7486, N7477);
buf BUF1 (N7487, N7473);
and AND4 (N7488, N7479, N3145, N3663, N743);
xor XOR2 (N7489, N7482, N2293);
nand NAND2 (N7490, N7489, N2183);
xor XOR2 (N7491, N7451, N5233);
not NOT1 (N7492, N7491);
and AND2 (N7493, N7474, N3098);
xor XOR2 (N7494, N7467, N2990);
nor NOR4 (N7495, N7481, N681, N2575, N6678);
buf BUF1 (N7496, N7492);
and AND2 (N7497, N7485, N7078);
not NOT1 (N7498, N7497);
nand NAND2 (N7499, N7490, N5934);
xor XOR2 (N7500, N7498, N4097);
and AND2 (N7501, N7488, N375);
nor NOR3 (N7502, N7493, N153, N7373);
not NOT1 (N7503, N7499);
xor XOR2 (N7504, N7484, N4795);
xor XOR2 (N7505, N7496, N3457);
buf BUF1 (N7506, N7487);
or OR4 (N7507, N7486, N3821, N5620, N3539);
and AND2 (N7508, N7506, N4434);
not NOT1 (N7509, N7504);
nor NOR2 (N7510, N7494, N4065);
xor XOR2 (N7511, N7508, N2737);
nor NOR3 (N7512, N7495, N6952, N231);
or OR2 (N7513, N7507, N1827);
buf BUF1 (N7514, N7513);
xor XOR2 (N7515, N7511, N3374);
not NOT1 (N7516, N7501);
xor XOR2 (N7517, N7512, N5295);
or OR2 (N7518, N7509, N1356);
buf BUF1 (N7519, N7503);
buf BUF1 (N7520, N7518);
or OR4 (N7521, N7520, N4702, N7212, N6785);
nand NAND3 (N7522, N7502, N672, N1377);
or OR4 (N7523, N7515, N6887, N2097, N248);
and AND4 (N7524, N7500, N7411, N506, N3223);
or OR2 (N7525, N7523, N3782);
nand NAND3 (N7526, N7519, N6445, N2932);
nor NOR3 (N7527, N7522, N1418, N5525);
or OR3 (N7528, N7517, N5264, N2324);
nor NOR2 (N7529, N7524, N5619);
xor XOR2 (N7530, N7516, N6545);
nor NOR2 (N7531, N7527, N5788);
and AND3 (N7532, N7514, N1470, N3814);
buf BUF1 (N7533, N7521);
nand NAND3 (N7534, N7532, N6559, N3269);
nand NAND2 (N7535, N7531, N1016);
nand NAND4 (N7536, N7505, N4723, N5150, N960);
or OR3 (N7537, N7528, N7049, N6556);
nor NOR2 (N7538, N7535, N2485);
or OR4 (N7539, N7538, N6739, N3340, N866);
or OR4 (N7540, N7510, N3421, N6173, N7314);
and AND3 (N7541, N7525, N3556, N369);
nand NAND3 (N7542, N7537, N230, N7382);
nand NAND4 (N7543, N7526, N4764, N4421, N6756);
nand NAND3 (N7544, N7533, N6346, N319);
not NOT1 (N7545, N7534);
nor NOR3 (N7546, N7539, N1889, N5744);
nand NAND4 (N7547, N7546, N4048, N6590, N1674);
and AND3 (N7548, N7547, N1204, N5032);
buf BUF1 (N7549, N7543);
or OR3 (N7550, N7529, N1769, N3633);
not NOT1 (N7551, N7530);
nor NOR4 (N7552, N7536, N5328, N1489, N6464);
buf BUF1 (N7553, N7545);
or OR3 (N7554, N7548, N6948, N3647);
nor NOR2 (N7555, N7542, N1629);
or OR2 (N7556, N7554, N3848);
nand NAND3 (N7557, N7552, N841, N1725);
nor NOR4 (N7558, N7556, N7115, N1559, N6689);
xor XOR2 (N7559, N7549, N4848);
buf BUF1 (N7560, N7544);
nand NAND4 (N7561, N7551, N800, N5343, N4102);
nor NOR4 (N7562, N7559, N2193, N6533, N6690);
or OR2 (N7563, N7558, N3444);
nor NOR3 (N7564, N7560, N2276, N1751);
or OR3 (N7565, N7555, N2370, N95);
nand NAND3 (N7566, N7561, N3519, N2876);
nor NOR3 (N7567, N7566, N5350, N1086);
nand NAND2 (N7568, N7541, N1155);
or OR3 (N7569, N7550, N2299, N1453);
or OR2 (N7570, N7568, N3999);
xor XOR2 (N7571, N7553, N65);
nor NOR3 (N7572, N7570, N5393, N6410);
and AND2 (N7573, N7557, N307);
not NOT1 (N7574, N7571);
nor NOR4 (N7575, N7540, N6774, N4096, N5031);
not NOT1 (N7576, N7565);
buf BUF1 (N7577, N7569);
buf BUF1 (N7578, N7572);
and AND2 (N7579, N7563, N539);
and AND4 (N7580, N7577, N7168, N7567, N1745);
not NOT1 (N7581, N5835);
nand NAND3 (N7582, N7578, N4414, N2170);
nand NAND4 (N7583, N7574, N3297, N940, N5678);
nand NAND3 (N7584, N7579, N2509, N6560);
xor XOR2 (N7585, N7582, N682);
not NOT1 (N7586, N7576);
not NOT1 (N7587, N7585);
not NOT1 (N7588, N7584);
nand NAND3 (N7589, N7580, N749, N4237);
and AND2 (N7590, N7583, N5516);
not NOT1 (N7591, N7562);
and AND2 (N7592, N7586, N1476);
or OR4 (N7593, N7573, N4838, N5019, N4346);
buf BUF1 (N7594, N7564);
or OR3 (N7595, N7593, N1689, N7534);
and AND2 (N7596, N7575, N340);
or OR3 (N7597, N7591, N312, N6804);
nor NOR4 (N7598, N7581, N1290, N7401, N1127);
nor NOR2 (N7599, N7589, N617);
nor NOR2 (N7600, N7592, N4741);
or OR3 (N7601, N7588, N1859, N2714);
xor XOR2 (N7602, N7598, N7278);
not NOT1 (N7603, N7600);
or OR2 (N7604, N7595, N4163);
nand NAND4 (N7605, N7599, N7233, N5149, N4489);
not NOT1 (N7606, N7590);
nand NAND2 (N7607, N7605, N2811);
and AND2 (N7608, N7601, N7287);
nor NOR3 (N7609, N7608, N7077, N6311);
not NOT1 (N7610, N7587);
or OR3 (N7611, N7602, N7360, N4160);
xor XOR2 (N7612, N7607, N7336);
xor XOR2 (N7613, N7606, N4157);
buf BUF1 (N7614, N7609);
buf BUF1 (N7615, N7597);
not NOT1 (N7616, N7603);
xor XOR2 (N7617, N7615, N4366);
and AND3 (N7618, N7594, N6114, N6513);
nand NAND2 (N7619, N7613, N1829);
xor XOR2 (N7620, N7612, N100);
nand NAND4 (N7621, N7611, N4886, N1930, N3318);
buf BUF1 (N7622, N7610);
xor XOR2 (N7623, N7616, N1761);
buf BUF1 (N7624, N7617);
nor NOR3 (N7625, N7604, N6930, N3366);
and AND2 (N7626, N7623, N405);
nand NAND3 (N7627, N7619, N113, N7261);
or OR3 (N7628, N7622, N4510, N7172);
nand NAND2 (N7629, N7628, N4869);
or OR2 (N7630, N7626, N5041);
and AND4 (N7631, N7624, N5724, N4302, N2797);
xor XOR2 (N7632, N7620, N7247);
buf BUF1 (N7633, N7629);
buf BUF1 (N7634, N7633);
and AND4 (N7635, N7634, N1669, N4293, N2736);
nor NOR2 (N7636, N7631, N3168);
nand NAND2 (N7637, N7621, N212);
and AND4 (N7638, N7596, N530, N3176, N4451);
not NOT1 (N7639, N7635);
nand NAND4 (N7640, N7638, N1996, N6635, N1056);
nor NOR4 (N7641, N7630, N2773, N2518, N3943);
nor NOR4 (N7642, N7639, N5529, N4230, N6833);
xor XOR2 (N7643, N7618, N6107);
and AND3 (N7644, N7642, N3060, N1621);
buf BUF1 (N7645, N7614);
not NOT1 (N7646, N7627);
or OR2 (N7647, N7636, N6913);
or OR3 (N7648, N7641, N4557, N4843);
not NOT1 (N7649, N7646);
and AND4 (N7650, N7637, N5826, N2016, N2091);
buf BUF1 (N7651, N7632);
and AND2 (N7652, N7644, N3883);
and AND2 (N7653, N7650, N3211);
buf BUF1 (N7654, N7625);
buf BUF1 (N7655, N7640);
not NOT1 (N7656, N7648);
nor NOR3 (N7657, N7645, N2357, N1984);
nand NAND2 (N7658, N7653, N7177);
not NOT1 (N7659, N7654);
buf BUF1 (N7660, N7657);
buf BUF1 (N7661, N7658);
not NOT1 (N7662, N7643);
nor NOR4 (N7663, N7660, N4289, N7230, N5724);
nand NAND2 (N7664, N7647, N4313);
not NOT1 (N7665, N7664);
not NOT1 (N7666, N7655);
not NOT1 (N7667, N7662);
xor XOR2 (N7668, N7666, N6772);
and AND3 (N7669, N7665, N4931, N5605);
buf BUF1 (N7670, N7663);
xor XOR2 (N7671, N7661, N5331);
and AND3 (N7672, N7651, N2702, N662);
buf BUF1 (N7673, N7669);
nor NOR4 (N7674, N7656, N4860, N1538, N3401);
or OR4 (N7675, N7649, N204, N2655, N6457);
nand NAND4 (N7676, N7671, N6198, N7482, N3317);
and AND3 (N7677, N7670, N1548, N5161);
nand NAND4 (N7678, N7667, N7238, N4642, N2769);
and AND3 (N7679, N7659, N1432, N2849);
nor NOR3 (N7680, N7677, N5130, N332);
and AND4 (N7681, N7668, N5545, N4781, N6620);
nor NOR4 (N7682, N7681, N509, N2370, N4522);
nand NAND2 (N7683, N7676, N943);
or OR3 (N7684, N7672, N5260, N7098);
not NOT1 (N7685, N7673);
xor XOR2 (N7686, N7674, N2737);
not NOT1 (N7687, N7678);
buf BUF1 (N7688, N7686);
xor XOR2 (N7689, N7679, N2749);
and AND4 (N7690, N7682, N3762, N5150, N5287);
nand NAND3 (N7691, N7685, N3551, N6506);
or OR4 (N7692, N7680, N639, N6847, N1156);
xor XOR2 (N7693, N7690, N6753);
not NOT1 (N7694, N7684);
nor NOR4 (N7695, N7683, N4952, N5617, N2681);
nand NAND3 (N7696, N7694, N4519, N6194);
not NOT1 (N7697, N7688);
or OR4 (N7698, N7675, N2716, N2220, N2649);
buf BUF1 (N7699, N7691);
buf BUF1 (N7700, N7697);
or OR3 (N7701, N7693, N5030, N5619);
or OR2 (N7702, N7689, N4059);
or OR2 (N7703, N7692, N2949);
xor XOR2 (N7704, N7701, N4516);
xor XOR2 (N7705, N7652, N5465);
and AND4 (N7706, N7702, N3763, N4868, N5570);
not NOT1 (N7707, N7706);
nand NAND4 (N7708, N7707, N2829, N5703, N517);
not NOT1 (N7709, N7705);
nor NOR3 (N7710, N7699, N3685, N3899);
buf BUF1 (N7711, N7704);
buf BUF1 (N7712, N7696);
xor XOR2 (N7713, N7698, N4798);
not NOT1 (N7714, N7695);
and AND2 (N7715, N7703, N4524);
nor NOR2 (N7716, N7714, N3852);
xor XOR2 (N7717, N7709, N7686);
xor XOR2 (N7718, N7713, N2138);
nand NAND3 (N7719, N7687, N2955, N7367);
buf BUF1 (N7720, N7710);
not NOT1 (N7721, N7708);
nand NAND3 (N7722, N7700, N3146, N1570);
nand NAND2 (N7723, N7716, N7678);
buf BUF1 (N7724, N7717);
nor NOR4 (N7725, N7724, N5490, N6202, N6166);
or OR4 (N7726, N7722, N1737, N2063, N6924);
xor XOR2 (N7727, N7718, N620);
nand NAND4 (N7728, N7719, N499, N7017, N4381);
buf BUF1 (N7729, N7711);
buf BUF1 (N7730, N7712);
nand NAND4 (N7731, N7720, N4774, N3284, N1295);
nand NAND3 (N7732, N7726, N7550, N3222);
nor NOR4 (N7733, N7723, N4725, N5821, N4129);
and AND2 (N7734, N7715, N1444);
buf BUF1 (N7735, N7728);
and AND3 (N7736, N7729, N6302, N1527);
and AND3 (N7737, N7730, N262, N1828);
or OR2 (N7738, N7732, N4191);
and AND3 (N7739, N7721, N1812, N2002);
xor XOR2 (N7740, N7727, N7072);
and AND4 (N7741, N7731, N6955, N6422, N7016);
nor NOR2 (N7742, N7734, N6479);
nor NOR2 (N7743, N7725, N898);
or OR2 (N7744, N7739, N53);
and AND2 (N7745, N7733, N5833);
nor NOR4 (N7746, N7740, N1092, N3941, N339);
buf BUF1 (N7747, N7743);
not NOT1 (N7748, N7737);
nor NOR3 (N7749, N7745, N4438, N3007);
nand NAND2 (N7750, N7746, N4890);
nand NAND2 (N7751, N7747, N7216);
and AND3 (N7752, N7751, N3757, N2804);
nor NOR3 (N7753, N7744, N6044, N1722);
nand NAND4 (N7754, N7752, N4596, N4150, N6710);
nor NOR3 (N7755, N7738, N1163, N4862);
buf BUF1 (N7756, N7754);
nor NOR2 (N7757, N7750, N4945);
nor NOR3 (N7758, N7736, N355, N406);
nor NOR2 (N7759, N7748, N6562);
nand NAND4 (N7760, N7742, N7319, N2536, N7159);
nand NAND4 (N7761, N7758, N4723, N5907, N5199);
nor NOR2 (N7762, N7753, N1623);
and AND4 (N7763, N7761, N3885, N2434, N5076);
or OR2 (N7764, N7757, N3975);
nand NAND4 (N7765, N7741, N5828, N4640, N7711);
xor XOR2 (N7766, N7764, N497);
not NOT1 (N7767, N7755);
not NOT1 (N7768, N7765);
or OR3 (N7769, N7756, N6732, N543);
not NOT1 (N7770, N7766);
and AND4 (N7771, N7763, N2073, N3237, N5722);
not NOT1 (N7772, N7769);
nand NAND3 (N7773, N7767, N2081, N6407);
and AND2 (N7774, N7768, N4121);
or OR4 (N7775, N7760, N6592, N5242, N3568);
not NOT1 (N7776, N7774);
buf BUF1 (N7777, N7771);
or OR4 (N7778, N7775, N1983, N431, N3916);
and AND4 (N7779, N7776, N6144, N947, N4629);
or OR2 (N7780, N7735, N7367);
not NOT1 (N7781, N7778);
nand NAND2 (N7782, N7773, N4789);
nor NOR2 (N7783, N7782, N7533);
nor NOR3 (N7784, N7777, N4113, N5667);
and AND3 (N7785, N7749, N7567, N5416);
nor NOR2 (N7786, N7780, N5365);
nand NAND4 (N7787, N7770, N896, N4336, N6088);
nor NOR3 (N7788, N7785, N5208, N1287);
nand NAND2 (N7789, N7783, N4154);
nand NAND3 (N7790, N7762, N5272, N3666);
xor XOR2 (N7791, N7788, N2794);
and AND3 (N7792, N7789, N816, N6701);
not NOT1 (N7793, N7779);
not NOT1 (N7794, N7792);
and AND2 (N7795, N7759, N2230);
or OR2 (N7796, N7784, N7058);
or OR4 (N7797, N7791, N7127, N4670, N5391);
or OR3 (N7798, N7797, N3265, N5004);
nand NAND3 (N7799, N7787, N1869, N4441);
nor NOR4 (N7800, N7798, N4815, N2538, N2546);
or OR2 (N7801, N7781, N5210);
nor NOR4 (N7802, N7795, N6001, N3473, N1469);
xor XOR2 (N7803, N7802, N837);
nor NOR4 (N7804, N7796, N745, N6871, N7266);
xor XOR2 (N7805, N7800, N6122);
not NOT1 (N7806, N7799);
not NOT1 (N7807, N7794);
nor NOR3 (N7808, N7793, N1076, N1664);
nor NOR2 (N7809, N7772, N3439);
xor XOR2 (N7810, N7803, N4316);
and AND4 (N7811, N7805, N2544, N5875, N277);
or OR2 (N7812, N7790, N1487);
not NOT1 (N7813, N7812);
and AND2 (N7814, N7809, N5873);
buf BUF1 (N7815, N7807);
xor XOR2 (N7816, N7815, N169);
buf BUF1 (N7817, N7816);
not NOT1 (N7818, N7808);
and AND2 (N7819, N7804, N6839);
nor NOR3 (N7820, N7811, N4348, N1005);
xor XOR2 (N7821, N7806, N3769);
not NOT1 (N7822, N7821);
buf BUF1 (N7823, N7818);
nand NAND2 (N7824, N7786, N7686);
or OR4 (N7825, N7820, N7702, N2493, N3941);
nor NOR2 (N7826, N7810, N2242);
nor NOR3 (N7827, N7824, N7244, N3673);
nor NOR4 (N7828, N7826, N4556, N1531, N4155);
buf BUF1 (N7829, N7801);
not NOT1 (N7830, N7814);
or OR3 (N7831, N7823, N7803, N293);
or OR4 (N7832, N7825, N2948, N5746, N7293);
nand NAND2 (N7833, N7829, N48);
xor XOR2 (N7834, N7827, N4213);
or OR3 (N7835, N7833, N83, N3345);
buf BUF1 (N7836, N7830);
and AND3 (N7837, N7832, N2840, N97);
or OR4 (N7838, N7831, N5006, N7655, N1613);
buf BUF1 (N7839, N7834);
or OR4 (N7840, N7836, N3562, N6383, N5938);
or OR3 (N7841, N7822, N1899, N3338);
nor NOR3 (N7842, N7841, N5448, N3806);
nor NOR3 (N7843, N7837, N7692, N1659);
xor XOR2 (N7844, N7819, N7501);
or OR4 (N7845, N7828, N942, N7626, N7836);
not NOT1 (N7846, N7835);
nand NAND3 (N7847, N7839, N2745, N2423);
and AND4 (N7848, N7813, N6392, N308, N2242);
xor XOR2 (N7849, N7840, N6278);
or OR3 (N7850, N7843, N1487, N6616);
buf BUF1 (N7851, N7846);
not NOT1 (N7852, N7817);
nand NAND2 (N7853, N7851, N6899);
or OR2 (N7854, N7852, N4988);
nor NOR2 (N7855, N7844, N1213);
and AND3 (N7856, N7849, N4666, N4241);
xor XOR2 (N7857, N7856, N7131);
nand NAND3 (N7858, N7838, N3624, N3357);
not NOT1 (N7859, N7855);
not NOT1 (N7860, N7858);
and AND4 (N7861, N7859, N2755, N5244, N7157);
xor XOR2 (N7862, N7848, N1269);
not NOT1 (N7863, N7861);
nand NAND3 (N7864, N7847, N7359, N5690);
nor NOR3 (N7865, N7850, N3740, N933);
buf BUF1 (N7866, N7862);
or OR3 (N7867, N7863, N7675, N5226);
and AND2 (N7868, N7845, N6886);
nand NAND2 (N7869, N7866, N5477);
or OR4 (N7870, N7867, N6010, N22, N4189);
buf BUF1 (N7871, N7865);
and AND4 (N7872, N7871, N3153, N6137, N3518);
or OR3 (N7873, N7872, N469, N1324);
xor XOR2 (N7874, N7873, N866);
not NOT1 (N7875, N7864);
buf BUF1 (N7876, N7874);
buf BUF1 (N7877, N7854);
xor XOR2 (N7878, N7853, N4900);
not NOT1 (N7879, N7878);
nand NAND2 (N7880, N7842, N1977);
not NOT1 (N7881, N7869);
xor XOR2 (N7882, N7857, N5851);
buf BUF1 (N7883, N7868);
xor XOR2 (N7884, N7877, N3851);
xor XOR2 (N7885, N7880, N2940);
or OR3 (N7886, N7884, N3857, N2237);
not NOT1 (N7887, N7885);
xor XOR2 (N7888, N7876, N6184);
nor NOR4 (N7889, N7875, N7276, N3036, N2495);
not NOT1 (N7890, N7889);
xor XOR2 (N7891, N7890, N6378);
nand NAND2 (N7892, N7879, N1821);
buf BUF1 (N7893, N7886);
not NOT1 (N7894, N7860);
and AND2 (N7895, N7888, N461);
buf BUF1 (N7896, N7893);
buf BUF1 (N7897, N7881);
nand NAND2 (N7898, N7892, N1344);
nand NAND3 (N7899, N7895, N4207, N3100);
or OR3 (N7900, N7891, N4744, N5395);
or OR2 (N7901, N7899, N1949);
xor XOR2 (N7902, N7882, N2815);
nor NOR3 (N7903, N7887, N6747, N2836);
xor XOR2 (N7904, N7870, N7540);
nor NOR3 (N7905, N7883, N4182, N974);
xor XOR2 (N7906, N7903, N769);
buf BUF1 (N7907, N7897);
nor NOR4 (N7908, N7906, N1365, N489, N4837);
not NOT1 (N7909, N7908);
nor NOR4 (N7910, N7900, N3735, N2025, N4307);
not NOT1 (N7911, N7894);
xor XOR2 (N7912, N7896, N5203);
nand NAND3 (N7913, N7905, N4526, N3413);
nand NAND2 (N7914, N7898, N910);
xor XOR2 (N7915, N7902, N7677);
nor NOR4 (N7916, N7901, N7814, N7115, N764);
nand NAND2 (N7917, N7913, N4570);
xor XOR2 (N7918, N7914, N6822);
buf BUF1 (N7919, N7904);
xor XOR2 (N7920, N7909, N5922);
not NOT1 (N7921, N7918);
nor NOR3 (N7922, N7910, N4058, N1452);
xor XOR2 (N7923, N7915, N2135);
nand NAND4 (N7924, N7920, N3145, N7438, N2991);
and AND3 (N7925, N7924, N2180, N2294);
nor NOR4 (N7926, N7916, N4948, N1383, N6367);
nand NAND2 (N7927, N7921, N6067);
nand NAND2 (N7928, N7927, N6654);
and AND4 (N7929, N7923, N2845, N2763, N7723);
buf BUF1 (N7930, N7926);
nand NAND4 (N7931, N7919, N2019, N5697, N1534);
nor NOR3 (N7932, N7925, N5828, N336);
not NOT1 (N7933, N7928);
nor NOR4 (N7934, N7922, N7581, N1254, N3591);
buf BUF1 (N7935, N7911);
and AND4 (N7936, N7934, N1093, N1505, N6235);
nor NOR4 (N7937, N7930, N1689, N6670, N2468);
nand NAND3 (N7938, N7912, N2642, N7325);
nor NOR3 (N7939, N7917, N6445, N1088);
and AND2 (N7940, N7939, N5174);
nand NAND3 (N7941, N7937, N919, N7880);
nand NAND4 (N7942, N7907, N903, N7697, N4741);
nor NOR3 (N7943, N7938, N3823, N2869);
or OR2 (N7944, N7935, N3837);
nand NAND2 (N7945, N7941, N5828);
and AND3 (N7946, N7943, N7699, N5616);
nand NAND3 (N7947, N7931, N5699, N1679);
and AND2 (N7948, N7929, N5966);
and AND2 (N7949, N7942, N2560);
and AND2 (N7950, N7933, N1108);
not NOT1 (N7951, N7949);
xor XOR2 (N7952, N7950, N510);
nor NOR4 (N7953, N7932, N1509, N2874, N1950);
or OR2 (N7954, N7951, N5629);
xor XOR2 (N7955, N7944, N3110);
nor NOR4 (N7956, N7936, N5900, N4794, N6989);
nand NAND3 (N7957, N7940, N42, N342);
and AND2 (N7958, N7954, N3694);
not NOT1 (N7959, N7947);
or OR2 (N7960, N7956, N2021);
buf BUF1 (N7961, N7960);
nor NOR4 (N7962, N7958, N4135, N5891, N139);
or OR4 (N7963, N7953, N7242, N5322, N1393);
nand NAND4 (N7964, N7961, N3337, N3380, N7090);
xor XOR2 (N7965, N7952, N7642);
nand NAND3 (N7966, N7946, N1473, N3945);
xor XOR2 (N7967, N7948, N1104);
nor NOR3 (N7968, N7963, N2601, N474);
nand NAND3 (N7969, N7965, N3117, N4778);
and AND2 (N7970, N7957, N5384);
xor XOR2 (N7971, N7968, N3264);
not NOT1 (N7972, N7971);
nor NOR3 (N7973, N7945, N6374, N7690);
buf BUF1 (N7974, N7955);
xor XOR2 (N7975, N7959, N5657);
xor XOR2 (N7976, N7975, N4708);
buf BUF1 (N7977, N7962);
buf BUF1 (N7978, N7966);
or OR2 (N7979, N7978, N1983);
nor NOR2 (N7980, N7973, N3833);
buf BUF1 (N7981, N7976);
xor XOR2 (N7982, N7981, N4510);
buf BUF1 (N7983, N7977);
nor NOR3 (N7984, N7972, N7810, N6618);
buf BUF1 (N7985, N7974);
nand NAND3 (N7986, N7980, N6773, N601);
and AND2 (N7987, N7970, N5705);
or OR4 (N7988, N7979, N1374, N6210, N5287);
nand NAND3 (N7989, N7984, N3930, N3230);
and AND3 (N7990, N7985, N5807, N7436);
and AND3 (N7991, N7969, N3357, N5766);
xor XOR2 (N7992, N7982, N5339);
xor XOR2 (N7993, N7988, N5586);
not NOT1 (N7994, N7991);
and AND4 (N7995, N7990, N1336, N146, N2545);
nand NAND2 (N7996, N7992, N466);
nand NAND2 (N7997, N7993, N2871);
nor NOR3 (N7998, N7996, N5569, N587);
or OR4 (N7999, N7967, N5150, N5921, N706);
or OR4 (N8000, N7998, N6394, N5927, N6597);
buf BUF1 (N8001, N7994);
or OR2 (N8002, N7999, N367);
not NOT1 (N8003, N7986);
not NOT1 (N8004, N7964);
buf BUF1 (N8005, N8004);
nor NOR2 (N8006, N7995, N2993);
buf BUF1 (N8007, N8003);
not NOT1 (N8008, N7997);
nor NOR2 (N8009, N7989, N3587);
nand NAND2 (N8010, N8009, N4975);
not NOT1 (N8011, N8001);
nand NAND3 (N8012, N8002, N613, N1695);
and AND4 (N8013, N8010, N4191, N947, N5235);
nand NAND3 (N8014, N8012, N496, N7848);
nor NOR3 (N8015, N8005, N7959, N1685);
xor XOR2 (N8016, N8011, N991);
not NOT1 (N8017, N7983);
nand NAND2 (N8018, N8008, N1936);
and AND3 (N8019, N8007, N4551, N2728);
not NOT1 (N8020, N8000);
or OR4 (N8021, N8018, N2614, N3483, N6835);
not NOT1 (N8022, N7987);
or OR3 (N8023, N8021, N7200, N353);
xor XOR2 (N8024, N8023, N3185);
not NOT1 (N8025, N8013);
not NOT1 (N8026, N8016);
xor XOR2 (N8027, N8019, N2926);
and AND2 (N8028, N8006, N1038);
and AND4 (N8029, N8024, N3774, N4526, N5435);
buf BUF1 (N8030, N8015);
buf BUF1 (N8031, N8028);
not NOT1 (N8032, N8020);
or OR4 (N8033, N8032, N339, N5025, N2611);
nand NAND4 (N8034, N8031, N4292, N3426, N6980);
buf BUF1 (N8035, N8025);
buf BUF1 (N8036, N8014);
or OR3 (N8037, N8017, N5144, N4988);
nand NAND3 (N8038, N8022, N3024, N7448);
xor XOR2 (N8039, N8037, N7201);
nand NAND3 (N8040, N8030, N4756, N7203);
buf BUF1 (N8041, N8034);
not NOT1 (N8042, N8027);
not NOT1 (N8043, N8035);
and AND3 (N8044, N8040, N3801, N7319);
nor NOR4 (N8045, N8026, N931, N2868, N6593);
and AND3 (N8046, N8041, N7987, N5087);
nor NOR3 (N8047, N8039, N3201, N6477);
nor NOR3 (N8048, N8033, N6027, N526);
buf BUF1 (N8049, N8042);
nand NAND4 (N8050, N8045, N1084, N3535, N7945);
buf BUF1 (N8051, N8048);
buf BUF1 (N8052, N8047);
buf BUF1 (N8053, N8050);
buf BUF1 (N8054, N8046);
nand NAND3 (N8055, N8054, N1014, N5264);
xor XOR2 (N8056, N8052, N394);
buf BUF1 (N8057, N8051);
nor NOR4 (N8058, N8044, N2350, N5258, N6393);
nand NAND4 (N8059, N8056, N1610, N5816, N559);
xor XOR2 (N8060, N8055, N1853);
nor NOR3 (N8061, N8058, N880, N2468);
not NOT1 (N8062, N8059);
buf BUF1 (N8063, N8057);
or OR4 (N8064, N8053, N6339, N7593, N6903);
buf BUF1 (N8065, N8038);
nor NOR3 (N8066, N8043, N5343, N620);
buf BUF1 (N8067, N8066);
xor XOR2 (N8068, N8065, N6058);
and AND2 (N8069, N8067, N4870);
and AND2 (N8070, N8049, N4232);
not NOT1 (N8071, N8036);
and AND2 (N8072, N8071, N1854);
or OR2 (N8073, N8063, N2911);
nand NAND4 (N8074, N8072, N5021, N1636, N5039);
and AND4 (N8075, N8073, N6873, N441, N5411);
not NOT1 (N8076, N8070);
nor NOR2 (N8077, N8029, N3968);
nand NAND3 (N8078, N8068, N6308, N3127);
nand NAND2 (N8079, N8060, N3534);
buf BUF1 (N8080, N8077);
not NOT1 (N8081, N8078);
and AND2 (N8082, N8080, N1533);
buf BUF1 (N8083, N8081);
nor NOR4 (N8084, N8075, N7143, N5449, N6210);
nand NAND4 (N8085, N8062, N4423, N3470, N608);
not NOT1 (N8086, N8074);
buf BUF1 (N8087, N8086);
and AND2 (N8088, N8064, N2182);
and AND4 (N8089, N8088, N3896, N1187, N7174);
buf BUF1 (N8090, N8061);
nor NOR3 (N8091, N8079, N6183, N2713);
nor NOR3 (N8092, N8087, N1219, N2513);
or OR4 (N8093, N8083, N7858, N7546, N6897);
nor NOR3 (N8094, N8076, N7434, N7529);
nor NOR2 (N8095, N8091, N4508);
not NOT1 (N8096, N8089);
nor NOR4 (N8097, N8094, N7790, N1369, N4659);
buf BUF1 (N8098, N8095);
buf BUF1 (N8099, N8097);
buf BUF1 (N8100, N8099);
and AND4 (N8101, N8093, N4173, N1337, N1725);
nand NAND2 (N8102, N8085, N2273);
and AND2 (N8103, N8098, N5754);
nand NAND4 (N8104, N8082, N3160, N1892, N3815);
or OR4 (N8105, N8100, N1183, N873, N1769);
buf BUF1 (N8106, N8069);
xor XOR2 (N8107, N8105, N6868);
buf BUF1 (N8108, N8103);
not NOT1 (N8109, N8096);
nand NAND4 (N8110, N8102, N3810, N7165, N2139);
not NOT1 (N8111, N8108);
and AND4 (N8112, N8109, N4375, N4163, N3437);
or OR4 (N8113, N8112, N711, N7302, N6499);
xor XOR2 (N8114, N8104, N8046);
or OR4 (N8115, N8084, N2812, N3697, N906);
and AND4 (N8116, N8111, N5122, N7484, N7739);
nand NAND2 (N8117, N8115, N505);
nand NAND4 (N8118, N8114, N19, N5088, N5291);
xor XOR2 (N8119, N8107, N7697);
and AND2 (N8120, N8101, N171);
nand NAND3 (N8121, N8119, N4071, N67);
nor NOR2 (N8122, N8113, N5616);
nor NOR3 (N8123, N8116, N2301, N3582);
xor XOR2 (N8124, N8092, N4839);
buf BUF1 (N8125, N8120);
not NOT1 (N8126, N8118);
nand NAND4 (N8127, N8122, N1164, N5945, N5664);
xor XOR2 (N8128, N8110, N7802);
and AND4 (N8129, N8123, N95, N2452, N7691);
not NOT1 (N8130, N8126);
nor NOR2 (N8131, N8117, N1926);
and AND4 (N8132, N8127, N4684, N7013, N252);
or OR4 (N8133, N8090, N1515, N1463, N2419);
xor XOR2 (N8134, N8128, N4957);
xor XOR2 (N8135, N8132, N5645);
xor XOR2 (N8136, N8129, N3136);
not NOT1 (N8137, N8124);
or OR4 (N8138, N8130, N5571, N1968, N4830);
nand NAND4 (N8139, N8133, N501, N1419, N4472);
or OR3 (N8140, N8134, N6512, N5305);
buf BUF1 (N8141, N8136);
xor XOR2 (N8142, N8139, N7942);
or OR2 (N8143, N8121, N1905);
or OR2 (N8144, N8140, N541);
and AND4 (N8145, N8142, N3704, N6771, N1591);
not NOT1 (N8146, N8125);
not NOT1 (N8147, N8131);
and AND3 (N8148, N8145, N7171, N3653);
not NOT1 (N8149, N8147);
xor XOR2 (N8150, N8146, N2283);
not NOT1 (N8151, N8148);
xor XOR2 (N8152, N8106, N328);
not NOT1 (N8153, N8141);
xor XOR2 (N8154, N8149, N2142);
or OR2 (N8155, N8151, N3809);
nor NOR4 (N8156, N8153, N6058, N7257, N7179);
or OR3 (N8157, N8156, N4018, N7007);
nor NOR2 (N8158, N8152, N360);
buf BUF1 (N8159, N8154);
nand NAND4 (N8160, N8155, N2364, N6656, N3181);
xor XOR2 (N8161, N8144, N1183);
buf BUF1 (N8162, N8160);
xor XOR2 (N8163, N8138, N6371);
not NOT1 (N8164, N8161);
xor XOR2 (N8165, N8135, N4895);
not NOT1 (N8166, N8162);
and AND3 (N8167, N8158, N1114, N3118);
buf BUF1 (N8168, N8163);
xor XOR2 (N8169, N8159, N1995);
nand NAND3 (N8170, N8169, N3061, N3391);
nor NOR3 (N8171, N8157, N892, N1506);
or OR2 (N8172, N8168, N3508);
or OR3 (N8173, N8137, N5671, N2962);
and AND3 (N8174, N8167, N1464, N5983);
xor XOR2 (N8175, N8166, N4541);
and AND3 (N8176, N8174, N6724, N6463);
xor XOR2 (N8177, N8165, N1658);
and AND4 (N8178, N8150, N4716, N3712, N2351);
xor XOR2 (N8179, N8170, N1864);
nand NAND3 (N8180, N8172, N5836, N4901);
nor NOR2 (N8181, N8176, N3041);
nor NOR4 (N8182, N8173, N1972, N6370, N1250);
or OR4 (N8183, N8180, N2045, N729, N7976);
xor XOR2 (N8184, N8164, N4598);
xor XOR2 (N8185, N8182, N557);
and AND4 (N8186, N8171, N707, N6593, N3303);
nand NAND2 (N8187, N8185, N5572);
nand NAND4 (N8188, N8143, N4146, N447, N5643);
not NOT1 (N8189, N8183);
not NOT1 (N8190, N8179);
nor NOR3 (N8191, N8188, N2953, N6579);
not NOT1 (N8192, N8178);
buf BUF1 (N8193, N8192);
not NOT1 (N8194, N8187);
xor XOR2 (N8195, N8190, N3687);
xor XOR2 (N8196, N8189, N6825);
buf BUF1 (N8197, N8194);
buf BUF1 (N8198, N8197);
and AND2 (N8199, N8193, N4975);
not NOT1 (N8200, N8196);
and AND4 (N8201, N8195, N5283, N3837, N484);
or OR2 (N8202, N8177, N6071);
nand NAND2 (N8203, N8184, N2289);
or OR3 (N8204, N8198, N148, N7978);
xor XOR2 (N8205, N8203, N2412);
and AND4 (N8206, N8201, N6221, N6261, N3418);
or OR3 (N8207, N8205, N4601, N6580);
or OR4 (N8208, N8175, N3536, N6921, N8048);
buf BUF1 (N8209, N8202);
nand NAND3 (N8210, N8191, N4999, N252);
nor NOR3 (N8211, N8206, N3163, N2760);
nor NOR3 (N8212, N8210, N416, N1821);
not NOT1 (N8213, N8181);
and AND3 (N8214, N8212, N7794, N7350);
xor XOR2 (N8215, N8208, N7847);
buf BUF1 (N8216, N8207);
buf BUF1 (N8217, N8213);
nor NOR3 (N8218, N8200, N4973, N5067);
and AND2 (N8219, N8214, N6657);
and AND3 (N8220, N8216, N2719, N509);
and AND3 (N8221, N8219, N3971, N6073);
or OR4 (N8222, N8186, N7112, N2911, N1257);
and AND2 (N8223, N8220, N8054);
nand NAND3 (N8224, N8211, N6209, N6283);
nor NOR4 (N8225, N8217, N1934, N7848, N4677);
or OR4 (N8226, N8199, N1411, N5093, N889);
and AND2 (N8227, N8223, N1720);
nand NAND4 (N8228, N8221, N50, N6133, N1038);
nand NAND3 (N8229, N8225, N6878, N4933);
or OR2 (N8230, N8224, N34);
and AND2 (N8231, N8229, N3137);
nor NOR3 (N8232, N8218, N6012, N2100);
buf BUF1 (N8233, N8230);
and AND4 (N8234, N8228, N8083, N7796, N5242);
not NOT1 (N8235, N8227);
xor XOR2 (N8236, N8235, N4063);
nor NOR4 (N8237, N8233, N1842, N362, N3062);
not NOT1 (N8238, N8234);
and AND4 (N8239, N8222, N6952, N39, N6403);
buf BUF1 (N8240, N8231);
and AND3 (N8241, N8239, N2959, N5671);
and AND4 (N8242, N8232, N1004, N4079, N3621);
buf BUF1 (N8243, N8209);
not NOT1 (N8244, N8240);
nor NOR2 (N8245, N8215, N2646);
not NOT1 (N8246, N8243);
xor XOR2 (N8247, N8242, N3356);
xor XOR2 (N8248, N8246, N7509);
buf BUF1 (N8249, N8226);
xor XOR2 (N8250, N8238, N7074);
xor XOR2 (N8251, N8248, N393);
nor NOR4 (N8252, N8247, N5807, N2619, N7426);
xor XOR2 (N8253, N8252, N5566);
and AND4 (N8254, N8249, N1778, N2018, N1789);
not NOT1 (N8255, N8250);
nor NOR2 (N8256, N8204, N622);
and AND4 (N8257, N8253, N7671, N2314, N6059);
buf BUF1 (N8258, N8257);
or OR2 (N8259, N8255, N330);
buf BUF1 (N8260, N8258);
buf BUF1 (N8261, N8251);
nor NOR2 (N8262, N8259, N5068);
xor XOR2 (N8263, N8244, N5939);
buf BUF1 (N8264, N8263);
nor NOR3 (N8265, N8262, N6457, N7628);
and AND4 (N8266, N8241, N5481, N84, N908);
buf BUF1 (N8267, N8245);
buf BUF1 (N8268, N8236);
and AND2 (N8269, N8265, N926);
nand NAND2 (N8270, N8261, N5799);
nor NOR4 (N8271, N8264, N8138, N2413, N4612);
xor XOR2 (N8272, N8267, N593);
nand NAND2 (N8273, N8271, N5998);
or OR2 (N8274, N8272, N1803);
nand NAND2 (N8275, N8273, N1305);
nor NOR4 (N8276, N8254, N2024, N167, N3116);
and AND3 (N8277, N8256, N641, N5992);
and AND3 (N8278, N8277, N3385, N1563);
nor NOR4 (N8279, N8237, N7253, N4994, N6222);
buf BUF1 (N8280, N8268);
or OR4 (N8281, N8260, N4450, N5666, N7502);
and AND2 (N8282, N8269, N557);
not NOT1 (N8283, N8282);
buf BUF1 (N8284, N8280);
buf BUF1 (N8285, N8278);
or OR2 (N8286, N8285, N6732);
not NOT1 (N8287, N8281);
not NOT1 (N8288, N8283);
not NOT1 (N8289, N8275);
nor NOR4 (N8290, N8279, N5113, N3224, N7540);
buf BUF1 (N8291, N8288);
xor XOR2 (N8292, N8274, N4324);
buf BUF1 (N8293, N8276);
not NOT1 (N8294, N8292);
not NOT1 (N8295, N8270);
not NOT1 (N8296, N8295);
nand NAND3 (N8297, N8290, N482, N7781);
buf BUF1 (N8298, N8297);
or OR4 (N8299, N8294, N5797, N8009, N1940);
or OR4 (N8300, N8293, N1344, N7113, N939);
or OR3 (N8301, N8286, N5905, N4163);
nand NAND3 (N8302, N8284, N1865, N5418);
xor XOR2 (N8303, N8287, N7259);
nand NAND2 (N8304, N8299, N4921);
buf BUF1 (N8305, N8303);
and AND4 (N8306, N8298, N990, N598, N4747);
nand NAND4 (N8307, N8306, N3446, N1988, N7285);
and AND2 (N8308, N8289, N6045);
not NOT1 (N8309, N8302);
or OR4 (N8310, N8300, N4018, N4350, N7182);
not NOT1 (N8311, N8310);
not NOT1 (N8312, N8311);
nor NOR2 (N8313, N8296, N343);
not NOT1 (N8314, N8307);
nand NAND2 (N8315, N8308, N930);
buf BUF1 (N8316, N8301);
xor XOR2 (N8317, N8314, N1595);
xor XOR2 (N8318, N8309, N5419);
buf BUF1 (N8319, N8312);
nor NOR2 (N8320, N8316, N817);
and AND2 (N8321, N8291, N6696);
or OR3 (N8322, N8313, N5829, N1128);
not NOT1 (N8323, N8322);
nor NOR2 (N8324, N8305, N699);
and AND4 (N8325, N8315, N76, N7798, N2182);
or OR2 (N8326, N8323, N62);
xor XOR2 (N8327, N8304, N1865);
nand NAND2 (N8328, N8325, N242);
nand NAND3 (N8329, N8326, N1320, N7485);
and AND2 (N8330, N8324, N6253);
not NOT1 (N8331, N8327);
buf BUF1 (N8332, N8319);
and AND4 (N8333, N8266, N1849, N1803, N5321);
nor NOR4 (N8334, N8329, N7267, N5065, N3400);
buf BUF1 (N8335, N8320);
or OR3 (N8336, N8331, N7467, N7925);
xor XOR2 (N8337, N8334, N7146);
nand NAND2 (N8338, N8318, N2149);
xor XOR2 (N8339, N8335, N5996);
not NOT1 (N8340, N8339);
not NOT1 (N8341, N8317);
and AND4 (N8342, N8337, N815, N1816, N4327);
buf BUF1 (N8343, N8328);
or OR4 (N8344, N8330, N6904, N4876, N6167);
and AND2 (N8345, N8333, N467);
xor XOR2 (N8346, N8345, N8075);
buf BUF1 (N8347, N8338);
buf BUF1 (N8348, N8336);
xor XOR2 (N8349, N8341, N1580);
or OR3 (N8350, N8342, N7580, N1226);
buf BUF1 (N8351, N8347);
not NOT1 (N8352, N8344);
nor NOR4 (N8353, N8349, N2409, N6110, N7791);
nand NAND4 (N8354, N8343, N2859, N4647, N4835);
nor NOR3 (N8355, N8346, N2958, N516);
buf BUF1 (N8356, N8354);
xor XOR2 (N8357, N8348, N3913);
nor NOR4 (N8358, N8321, N2281, N3345, N3841);
and AND3 (N8359, N8356, N6911, N2110);
xor XOR2 (N8360, N8351, N4636);
nand NAND2 (N8361, N8357, N1476);
not NOT1 (N8362, N8360);
xor XOR2 (N8363, N8332, N2333);
xor XOR2 (N8364, N8340, N1664);
buf BUF1 (N8365, N8358);
nand NAND4 (N8366, N8352, N3491, N6304, N5553);
xor XOR2 (N8367, N8355, N7387);
nand NAND3 (N8368, N8363, N912, N2403);
not NOT1 (N8369, N8367);
not NOT1 (N8370, N8361);
nand NAND4 (N8371, N8359, N7351, N1629, N7129);
not NOT1 (N8372, N8364);
or OR3 (N8373, N8369, N7535, N202);
or OR4 (N8374, N8373, N4423, N39, N1857);
nand NAND2 (N8375, N8368, N8095);
or OR4 (N8376, N8372, N6940, N5974, N2191);
xor XOR2 (N8377, N8375, N7050);
and AND3 (N8378, N8370, N8038, N7383);
not NOT1 (N8379, N8365);
or OR4 (N8380, N8371, N2826, N2376, N7461);
nand NAND3 (N8381, N8379, N1707, N49);
buf BUF1 (N8382, N8353);
not NOT1 (N8383, N8380);
not NOT1 (N8384, N8366);
nor NOR4 (N8385, N8381, N5283, N2857, N4550);
buf BUF1 (N8386, N8384);
or OR3 (N8387, N8350, N6114, N6950);
nand NAND4 (N8388, N8378, N3325, N7807, N5146);
and AND2 (N8389, N8385, N7908);
not NOT1 (N8390, N8374);
or OR4 (N8391, N8389, N7687, N2980, N437);
or OR3 (N8392, N8390, N1701, N6997);
nand NAND4 (N8393, N8392, N4544, N2895, N6643);
xor XOR2 (N8394, N8362, N1371);
not NOT1 (N8395, N8383);
and AND4 (N8396, N8394, N7608, N382, N2937);
xor XOR2 (N8397, N8386, N6552);
and AND2 (N8398, N8397, N8305);
xor XOR2 (N8399, N8393, N4085);
nor NOR2 (N8400, N8382, N5089);
and AND3 (N8401, N8398, N2959, N2696);
xor XOR2 (N8402, N8388, N4854);
not NOT1 (N8403, N8402);
buf BUF1 (N8404, N8403);
buf BUF1 (N8405, N8400);
or OR3 (N8406, N8376, N3436, N6612);
nand NAND3 (N8407, N8405, N3004, N3668);
nor NOR2 (N8408, N8395, N5552);
xor XOR2 (N8409, N8387, N6669);
nor NOR4 (N8410, N8406, N5934, N2900, N7350);
not NOT1 (N8411, N8399);
nor NOR2 (N8412, N8404, N6326);
and AND4 (N8413, N8401, N2894, N5797, N5175);
buf BUF1 (N8414, N8413);
buf BUF1 (N8415, N8396);
xor XOR2 (N8416, N8412, N4256);
nand NAND3 (N8417, N8416, N5427, N2812);
not NOT1 (N8418, N8407);
buf BUF1 (N8419, N8417);
nor NOR2 (N8420, N8418, N344);
or OR3 (N8421, N8415, N156, N1058);
not NOT1 (N8422, N8377);
not NOT1 (N8423, N8411);
buf BUF1 (N8424, N8419);
not NOT1 (N8425, N8408);
buf BUF1 (N8426, N8410);
not NOT1 (N8427, N8420);
xor XOR2 (N8428, N8424, N409);
buf BUF1 (N8429, N8421);
or OR4 (N8430, N8428, N5737, N8389, N6472);
and AND3 (N8431, N8414, N3973, N6412);
xor XOR2 (N8432, N8429, N1523);
xor XOR2 (N8433, N8409, N2974);
buf BUF1 (N8434, N8426);
and AND4 (N8435, N8391, N3756, N1719, N7802);
nand NAND3 (N8436, N8432, N3174, N5279);
and AND2 (N8437, N8431, N188);
not NOT1 (N8438, N8437);
buf BUF1 (N8439, N8427);
nand NAND2 (N8440, N8438, N5022);
or OR3 (N8441, N8440, N207, N6933);
nand NAND2 (N8442, N8433, N7604);
and AND2 (N8443, N8436, N3508);
and AND4 (N8444, N8443, N8363, N7011, N8032);
nor NOR4 (N8445, N8422, N3521, N5859, N617);
and AND4 (N8446, N8439, N4346, N1660, N7193);
not NOT1 (N8447, N8434);
nand NAND2 (N8448, N8446, N5779);
not NOT1 (N8449, N8442);
nor NOR3 (N8450, N8447, N6335, N7716);
nand NAND3 (N8451, N8435, N809, N5794);
buf BUF1 (N8452, N8423);
nand NAND2 (N8453, N8449, N5652);
nand NAND3 (N8454, N8425, N7731, N4642);
buf BUF1 (N8455, N8451);
nor NOR2 (N8456, N8430, N7726);
nand NAND2 (N8457, N8453, N5838);
or OR3 (N8458, N8441, N44, N4332);
not NOT1 (N8459, N8455);
buf BUF1 (N8460, N8459);
xor XOR2 (N8461, N8458, N3481);
xor XOR2 (N8462, N8461, N1228);
buf BUF1 (N8463, N8452);
and AND4 (N8464, N8456, N8434, N97, N6713);
buf BUF1 (N8465, N8445);
not NOT1 (N8466, N8463);
nor NOR3 (N8467, N8462, N2700, N2042);
or OR3 (N8468, N8466, N7103, N1696);
xor XOR2 (N8469, N8468, N6794);
nor NOR3 (N8470, N8454, N7139, N4480);
xor XOR2 (N8471, N8450, N7144);
and AND3 (N8472, N8469, N2973, N1651);
and AND4 (N8473, N8465, N2591, N1495, N1492);
buf BUF1 (N8474, N8471);
nand NAND2 (N8475, N8448, N7217);
not NOT1 (N8476, N8467);
and AND3 (N8477, N8473, N4243, N2831);
not NOT1 (N8478, N8472);
buf BUF1 (N8479, N8457);
buf BUF1 (N8480, N8444);
or OR2 (N8481, N8478, N3143);
buf BUF1 (N8482, N8480);
nor NOR3 (N8483, N8476, N5125, N2010);
and AND2 (N8484, N8482, N942);
buf BUF1 (N8485, N8479);
or OR2 (N8486, N8474, N4181);
and AND2 (N8487, N8481, N5363);
not NOT1 (N8488, N8464);
not NOT1 (N8489, N8486);
buf BUF1 (N8490, N8485);
nand NAND4 (N8491, N8475, N3114, N2184, N3960);
nand NAND3 (N8492, N8460, N813, N4830);
and AND2 (N8493, N8492, N1240);
xor XOR2 (N8494, N8470, N1794);
or OR2 (N8495, N8491, N2445);
nor NOR4 (N8496, N8493, N3660, N7500, N318);
buf BUF1 (N8497, N8483);
xor XOR2 (N8498, N8494, N4503);
xor XOR2 (N8499, N8488, N6774);
xor XOR2 (N8500, N8477, N1990);
nand NAND3 (N8501, N8497, N6495, N4652);
and AND4 (N8502, N8500, N5691, N3100, N7778);
nor NOR3 (N8503, N8501, N4622, N7921);
not NOT1 (N8504, N8503);
nand NAND2 (N8505, N8504, N7967);
nand NAND2 (N8506, N8499, N5810);
xor XOR2 (N8507, N8505, N1741);
not NOT1 (N8508, N8502);
not NOT1 (N8509, N8484);
and AND2 (N8510, N8498, N3660);
xor XOR2 (N8511, N8490, N3034);
buf BUF1 (N8512, N8495);
and AND3 (N8513, N8489, N6686, N1781);
nor NOR4 (N8514, N8506, N4207, N3764, N5120);
xor XOR2 (N8515, N8511, N4437);
xor XOR2 (N8516, N8509, N6145);
buf BUF1 (N8517, N8512);
buf BUF1 (N8518, N8487);
and AND3 (N8519, N8510, N4281, N3119);
nor NOR2 (N8520, N8496, N7544);
buf BUF1 (N8521, N8513);
xor XOR2 (N8522, N8521, N6522);
buf BUF1 (N8523, N8518);
or OR3 (N8524, N8515, N5872, N1808);
nor NOR2 (N8525, N8524, N6155);
and AND3 (N8526, N8519, N1878, N1297);
nor NOR3 (N8527, N8526, N215, N1694);
or OR2 (N8528, N8520, N3779);
and AND3 (N8529, N8523, N7075, N3163);
nand NAND4 (N8530, N8517, N1330, N1112, N4551);
not NOT1 (N8531, N8514);
buf BUF1 (N8532, N8527);
not NOT1 (N8533, N8525);
nand NAND2 (N8534, N8530, N3433);
xor XOR2 (N8535, N8534, N3905);
buf BUF1 (N8536, N8531);
xor XOR2 (N8537, N8507, N7676);
nand NAND2 (N8538, N8536, N387);
nand NAND2 (N8539, N8516, N6186);
nor NOR4 (N8540, N8539, N2995, N5789, N4319);
or OR3 (N8541, N8529, N2694, N6120);
buf BUF1 (N8542, N8532);
or OR4 (N8543, N8528, N737, N4563, N6823);
nor NOR4 (N8544, N8542, N2195, N4905, N6065);
or OR2 (N8545, N8538, N4453);
xor XOR2 (N8546, N8540, N4592);
nor NOR2 (N8547, N8544, N4884);
buf BUF1 (N8548, N8543);
xor XOR2 (N8549, N8508, N3810);
not NOT1 (N8550, N8522);
buf BUF1 (N8551, N8548);
nand NAND3 (N8552, N8547, N6838, N3033);
not NOT1 (N8553, N8549);
or OR2 (N8554, N8541, N5818);
or OR4 (N8555, N8552, N4388, N6775, N1018);
nor NOR4 (N8556, N8554, N3138, N5402, N6050);
nor NOR2 (N8557, N8555, N6986);
and AND4 (N8558, N8533, N2383, N4796, N7048);
buf BUF1 (N8559, N8535);
not NOT1 (N8560, N8556);
or OR2 (N8561, N8560, N5643);
and AND2 (N8562, N8550, N2350);
xor XOR2 (N8563, N8557, N300);
xor XOR2 (N8564, N8553, N7889);
buf BUF1 (N8565, N8551);
nand NAND3 (N8566, N8545, N3383, N88);
or OR3 (N8567, N8537, N806, N914);
or OR4 (N8568, N8562, N6562, N4294, N4727);
xor XOR2 (N8569, N8558, N5980);
xor XOR2 (N8570, N8564, N8260);
or OR2 (N8571, N8559, N103);
xor XOR2 (N8572, N8569, N1466);
or OR3 (N8573, N8571, N5424, N5510);
xor XOR2 (N8574, N8565, N595);
and AND4 (N8575, N8567, N2753, N1208, N6060);
buf BUF1 (N8576, N8563);
nand NAND3 (N8577, N8568, N1633, N325);
buf BUF1 (N8578, N8576);
or OR2 (N8579, N8572, N3549);
xor XOR2 (N8580, N8570, N4081);
not NOT1 (N8581, N8580);
nand NAND4 (N8582, N8579, N7123, N5992, N1267);
buf BUF1 (N8583, N8575);
nand NAND4 (N8584, N8546, N5923, N7911, N3895);
not NOT1 (N8585, N8573);
nand NAND4 (N8586, N8577, N3251, N819, N2737);
nor NOR2 (N8587, N8586, N2636);
nand NAND3 (N8588, N8561, N7383, N1265);
and AND3 (N8589, N8587, N6331, N6065);
or OR4 (N8590, N8574, N2477, N4456, N5237);
and AND2 (N8591, N8584, N1996);
not NOT1 (N8592, N8589);
and AND3 (N8593, N8582, N495, N2964);
xor XOR2 (N8594, N8583, N8447);
and AND2 (N8595, N8594, N7969);
xor XOR2 (N8596, N8595, N5189);
not NOT1 (N8597, N8588);
nor NOR4 (N8598, N8591, N2590, N860, N6539);
nor NOR4 (N8599, N8598, N1202, N4220, N6447);
nand NAND4 (N8600, N8593, N1576, N47, N4131);
nand NAND4 (N8601, N8566, N2501, N2167, N340);
nor NOR2 (N8602, N8601, N3633);
xor XOR2 (N8603, N8597, N2272);
or OR2 (N8604, N8596, N8422);
nor NOR4 (N8605, N8599, N7629, N6486, N2670);
buf BUF1 (N8606, N8585);
xor XOR2 (N8607, N8581, N187);
not NOT1 (N8608, N8607);
nor NOR4 (N8609, N8604, N2116, N4969, N4630);
xor XOR2 (N8610, N8602, N8088);
not NOT1 (N8611, N8605);
not NOT1 (N8612, N8600);
nand NAND4 (N8613, N8590, N7509, N5303, N8202);
nor NOR3 (N8614, N8592, N3859, N2149);
not NOT1 (N8615, N8578);
nor NOR2 (N8616, N8606, N6850);
and AND4 (N8617, N8611, N6931, N2238, N1705);
and AND2 (N8618, N8612, N835);
nand NAND3 (N8619, N8617, N1008, N140);
xor XOR2 (N8620, N8608, N8383);
not NOT1 (N8621, N8620);
and AND4 (N8622, N8618, N4331, N7243, N4934);
not NOT1 (N8623, N8609);
not NOT1 (N8624, N8621);
or OR2 (N8625, N8624, N872);
xor XOR2 (N8626, N8622, N6784);
nor NOR2 (N8627, N8614, N3151);
or OR3 (N8628, N8627, N5980, N697);
nor NOR4 (N8629, N8613, N7832, N2809, N7053);
xor XOR2 (N8630, N8603, N1792);
nor NOR4 (N8631, N8623, N2622, N3641, N543);
or OR3 (N8632, N8625, N6319, N71);
xor XOR2 (N8633, N8616, N1624);
buf BUF1 (N8634, N8619);
buf BUF1 (N8635, N8628);
nand NAND4 (N8636, N8610, N418, N6684, N2737);
nor NOR3 (N8637, N8635, N2547, N7976);
xor XOR2 (N8638, N8631, N688);
nand NAND3 (N8639, N8634, N2040, N4434);
or OR4 (N8640, N8636, N1579, N583, N6901);
not NOT1 (N8641, N8639);
nor NOR2 (N8642, N8626, N6217);
and AND2 (N8643, N8629, N2782);
not NOT1 (N8644, N8632);
nand NAND3 (N8645, N8640, N5530, N731);
or OR3 (N8646, N8638, N4016, N8407);
buf BUF1 (N8647, N8646);
xor XOR2 (N8648, N8615, N3280);
nand NAND4 (N8649, N8641, N1628, N1964, N5649);
buf BUF1 (N8650, N8643);
not NOT1 (N8651, N8649);
not NOT1 (N8652, N8650);
nor NOR3 (N8653, N8648, N7589, N3025);
and AND2 (N8654, N8644, N1904);
xor XOR2 (N8655, N8637, N2977);
xor XOR2 (N8656, N8651, N4852);
not NOT1 (N8657, N8642);
xor XOR2 (N8658, N8657, N4488);
nand NAND3 (N8659, N8658, N7358, N4517);
nand NAND4 (N8660, N8645, N7345, N7530, N8202);
buf BUF1 (N8661, N8660);
xor XOR2 (N8662, N8630, N2127);
buf BUF1 (N8663, N8647);
nand NAND2 (N8664, N8663, N3537);
or OR4 (N8665, N8633, N6021, N4544, N8232);
not NOT1 (N8666, N8661);
and AND2 (N8667, N8656, N3943);
nand NAND2 (N8668, N8653, N3563);
nor NOR4 (N8669, N8652, N423, N4135, N6405);
not NOT1 (N8670, N8654);
not NOT1 (N8671, N8664);
not NOT1 (N8672, N8667);
nand NAND3 (N8673, N8671, N1398, N5);
buf BUF1 (N8674, N8673);
and AND2 (N8675, N8666, N518);
nand NAND2 (N8676, N8655, N2910);
xor XOR2 (N8677, N8672, N7307);
nand NAND2 (N8678, N8670, N5277);
nor NOR4 (N8679, N8674, N4349, N1113, N5113);
or OR3 (N8680, N8659, N4283, N2732);
xor XOR2 (N8681, N8662, N1405);
buf BUF1 (N8682, N8681);
not NOT1 (N8683, N8668);
nand NAND2 (N8684, N8677, N7031);
nor NOR4 (N8685, N8682, N6933, N1512, N807);
buf BUF1 (N8686, N8683);
or OR4 (N8687, N8665, N1975, N1157, N6169);
buf BUF1 (N8688, N8680);
and AND3 (N8689, N8676, N2672, N8445);
nand NAND2 (N8690, N8687, N2859);
nor NOR3 (N8691, N8675, N6795, N8662);
and AND3 (N8692, N8686, N3698, N2469);
or OR2 (N8693, N8679, N7127);
xor XOR2 (N8694, N8689, N8432);
and AND4 (N8695, N8688, N5587, N1840, N2339);
xor XOR2 (N8696, N8691, N6570);
buf BUF1 (N8697, N8669);
nor NOR4 (N8698, N8692, N7658, N7313, N5793);
not NOT1 (N8699, N8693);
or OR3 (N8700, N8678, N6524, N1337);
buf BUF1 (N8701, N8695);
and AND3 (N8702, N8694, N2321, N1374);
and AND2 (N8703, N8684, N3224);
nand NAND4 (N8704, N8703, N8610, N4971, N2718);
xor XOR2 (N8705, N8701, N4557);
not NOT1 (N8706, N8698);
or OR3 (N8707, N8697, N4235, N7123);
nand NAND4 (N8708, N8707, N6988, N8008, N981);
not NOT1 (N8709, N8704);
and AND4 (N8710, N8709, N5431, N2404, N4371);
and AND4 (N8711, N8690, N7373, N15, N398);
xor XOR2 (N8712, N8710, N7273);
or OR4 (N8713, N8700, N1967, N2531, N213);
or OR3 (N8714, N8708, N363, N383);
buf BUF1 (N8715, N8702);
or OR2 (N8716, N8706, N3181);
buf BUF1 (N8717, N8713);
nand NAND3 (N8718, N8696, N6691, N8682);
buf BUF1 (N8719, N8716);
not NOT1 (N8720, N8719);
or OR2 (N8721, N8711, N5600);
xor XOR2 (N8722, N8717, N8721);
not NOT1 (N8723, N6812);
or OR3 (N8724, N8685, N5076, N6468);
nor NOR3 (N8725, N8718, N1326, N5749);
nand NAND2 (N8726, N8724, N4104);
not NOT1 (N8727, N8715);
or OR2 (N8728, N8714, N4769);
and AND4 (N8729, N8723, N5568, N3346, N7043);
xor XOR2 (N8730, N8720, N4029);
nor NOR4 (N8731, N8726, N154, N1100, N959);
xor XOR2 (N8732, N8727, N1783);
buf BUF1 (N8733, N8712);
nand NAND2 (N8734, N8733, N7194);
and AND3 (N8735, N8699, N8654, N358);
xor XOR2 (N8736, N8705, N8084);
not NOT1 (N8737, N8732);
xor XOR2 (N8738, N8735, N3833);
buf BUF1 (N8739, N8736);
buf BUF1 (N8740, N8739);
not NOT1 (N8741, N8731);
nand NAND2 (N8742, N8725, N5551);
buf BUF1 (N8743, N8737);
or OR3 (N8744, N8740, N2131, N4263);
and AND4 (N8745, N8742, N7127, N22, N3990);
nand NAND2 (N8746, N8744, N117);
not NOT1 (N8747, N8734);
or OR4 (N8748, N8722, N7528, N146, N7218);
nor NOR3 (N8749, N8728, N4589, N594);
not NOT1 (N8750, N8729);
nor NOR2 (N8751, N8747, N1383);
or OR3 (N8752, N8749, N6917, N5375);
buf BUF1 (N8753, N8746);
and AND4 (N8754, N8751, N2223, N7346, N4437);
or OR3 (N8755, N8745, N970, N4655);
nor NOR2 (N8756, N8750, N7309);
xor XOR2 (N8757, N8756, N3835);
nand NAND2 (N8758, N8754, N2825);
xor XOR2 (N8759, N8758, N3539);
xor XOR2 (N8760, N8755, N7412);
nor NOR4 (N8761, N8741, N2692, N3064, N1378);
buf BUF1 (N8762, N8743);
and AND3 (N8763, N8753, N4267, N6202);
not NOT1 (N8764, N8759);
buf BUF1 (N8765, N8748);
and AND3 (N8766, N8764, N1837, N3583);
and AND3 (N8767, N8766, N1727, N1063);
nand NAND3 (N8768, N8763, N41, N4016);
xor XOR2 (N8769, N8760, N7495);
nor NOR3 (N8770, N8761, N2470, N7864);
xor XOR2 (N8771, N8757, N2385);
nor NOR3 (N8772, N8752, N1515, N1150);
or OR2 (N8773, N8772, N5879);
buf BUF1 (N8774, N8730);
buf BUF1 (N8775, N8767);
nor NOR3 (N8776, N8774, N1035, N8408);
not NOT1 (N8777, N8773);
not NOT1 (N8778, N8771);
and AND2 (N8779, N8765, N1240);
nor NOR4 (N8780, N8768, N8004, N8051, N4480);
xor XOR2 (N8781, N8778, N5497);
xor XOR2 (N8782, N8780, N541);
nand NAND4 (N8783, N8762, N2267, N8391, N1150);
buf BUF1 (N8784, N8781);
or OR3 (N8785, N8770, N5630, N8348);
nor NOR4 (N8786, N8776, N7953, N1664, N8437);
not NOT1 (N8787, N8738);
and AND2 (N8788, N8775, N5553);
nor NOR4 (N8789, N8786, N3897, N2341, N5210);
nand NAND3 (N8790, N8789, N5065, N792);
and AND4 (N8791, N8785, N5345, N3188, N8321);
xor XOR2 (N8792, N8790, N8125);
or OR3 (N8793, N8777, N3450, N8312);
xor XOR2 (N8794, N8787, N7098);
nor NOR2 (N8795, N8784, N381);
and AND4 (N8796, N8783, N852, N687, N3092);
and AND2 (N8797, N8793, N4511);
xor XOR2 (N8798, N8791, N7165);
xor XOR2 (N8799, N8794, N4736);
xor XOR2 (N8800, N8795, N3736);
or OR3 (N8801, N8796, N5041, N115);
xor XOR2 (N8802, N8782, N5085);
not NOT1 (N8803, N8779);
buf BUF1 (N8804, N8788);
nand NAND3 (N8805, N8802, N5442, N2235);
xor XOR2 (N8806, N8792, N2792);
xor XOR2 (N8807, N8804, N3324);
and AND3 (N8808, N8801, N103, N8712);
buf BUF1 (N8809, N8797);
buf BUF1 (N8810, N8803);
nand NAND3 (N8811, N8798, N8409, N201);
buf BUF1 (N8812, N8809);
nand NAND3 (N8813, N8769, N3622, N419);
nor NOR4 (N8814, N8800, N193, N3381, N6919);
not NOT1 (N8815, N8810);
not NOT1 (N8816, N8813);
buf BUF1 (N8817, N8816);
not NOT1 (N8818, N8817);
nor NOR4 (N8819, N8818, N918, N852, N8426);
nor NOR2 (N8820, N8807, N6912);
not NOT1 (N8821, N8805);
not NOT1 (N8822, N8814);
and AND2 (N8823, N8820, N1840);
xor XOR2 (N8824, N8812, N469);
buf BUF1 (N8825, N8821);
nor NOR3 (N8826, N8825, N4602, N4306);
nand NAND4 (N8827, N8815, N5590, N642, N7523);
or OR4 (N8828, N8826, N6460, N6115, N7274);
nand NAND2 (N8829, N8806, N6821);
not NOT1 (N8830, N8823);
xor XOR2 (N8831, N8828, N551);
xor XOR2 (N8832, N8827, N1302);
and AND2 (N8833, N8811, N5724);
and AND3 (N8834, N8833, N126, N291);
buf BUF1 (N8835, N8822);
not NOT1 (N8836, N8824);
not NOT1 (N8837, N8834);
or OR2 (N8838, N8835, N3010);
or OR2 (N8839, N8830, N8576);
or OR4 (N8840, N8832, N4624, N1261, N1764);
nand NAND3 (N8841, N8808, N7099, N7764);
not NOT1 (N8842, N8841);
not NOT1 (N8843, N8836);
or OR4 (N8844, N8840, N7067, N6998, N5392);
not NOT1 (N8845, N8829);
not NOT1 (N8846, N8831);
not NOT1 (N8847, N8844);
and AND2 (N8848, N8839, N3410);
or OR3 (N8849, N8837, N6709, N7904);
not NOT1 (N8850, N8849);
not NOT1 (N8851, N8846);
not NOT1 (N8852, N8845);
not NOT1 (N8853, N8850);
nand NAND3 (N8854, N8851, N7804, N6319);
nor NOR4 (N8855, N8854, N6929, N3473, N2192);
xor XOR2 (N8856, N8848, N472);
xor XOR2 (N8857, N8852, N6825);
and AND3 (N8858, N8857, N4119, N5873);
and AND4 (N8859, N8842, N7528, N1333, N8168);
nand NAND4 (N8860, N8856, N4380, N6790, N7339);
or OR3 (N8861, N8838, N2494, N7765);
or OR3 (N8862, N8859, N1959, N3428);
or OR2 (N8863, N8855, N8114);
and AND4 (N8864, N8819, N7129, N7249, N5753);
buf BUF1 (N8865, N8862);
not NOT1 (N8866, N8843);
not NOT1 (N8867, N8858);
nor NOR2 (N8868, N8847, N3486);
buf BUF1 (N8869, N8866);
nor NOR4 (N8870, N8861, N4822, N5009, N6981);
nand NAND2 (N8871, N8867, N3911);
and AND3 (N8872, N8864, N6572, N3456);
not NOT1 (N8873, N8871);
and AND3 (N8874, N8799, N1339, N8270);
and AND3 (N8875, N8874, N1090, N1307);
or OR4 (N8876, N8865, N6838, N5940, N6564);
and AND3 (N8877, N8853, N7212, N7935);
not NOT1 (N8878, N8873);
xor XOR2 (N8879, N8872, N3583);
and AND2 (N8880, N8868, N8198);
nor NOR4 (N8881, N8863, N8263, N1132, N3099);
buf BUF1 (N8882, N8875);
not NOT1 (N8883, N8860);
nor NOR2 (N8884, N8876, N5565);
nand NAND2 (N8885, N8882, N6808);
buf BUF1 (N8886, N8881);
or OR3 (N8887, N8877, N4364, N7503);
buf BUF1 (N8888, N8887);
buf BUF1 (N8889, N8886);
or OR2 (N8890, N8869, N4773);
or OR4 (N8891, N8878, N5906, N5036, N1470);
and AND3 (N8892, N8884, N91, N2529);
not NOT1 (N8893, N8891);
or OR2 (N8894, N8870, N537);
and AND4 (N8895, N8890, N2451, N8406, N5786);
xor XOR2 (N8896, N8892, N3084);
not NOT1 (N8897, N8889);
nor NOR3 (N8898, N8880, N2338, N3277);
buf BUF1 (N8899, N8898);
buf BUF1 (N8900, N8894);
buf BUF1 (N8901, N8883);
buf BUF1 (N8902, N8901);
and AND3 (N8903, N8899, N3707, N4143);
not NOT1 (N8904, N8895);
nor NOR4 (N8905, N8879, N8356, N4127, N7155);
nand NAND2 (N8906, N8903, N1171);
buf BUF1 (N8907, N8906);
xor XOR2 (N8908, N8902, N809);
or OR2 (N8909, N8885, N741);
buf BUF1 (N8910, N8905);
and AND3 (N8911, N8904, N7189, N6038);
not NOT1 (N8912, N8908);
nand NAND2 (N8913, N8910, N3743);
nor NOR3 (N8914, N8900, N8276, N3355);
xor XOR2 (N8915, N8909, N4698);
nor NOR2 (N8916, N8915, N1680);
and AND3 (N8917, N8893, N1321, N4491);
buf BUF1 (N8918, N8888);
and AND2 (N8919, N8916, N1932);
and AND4 (N8920, N8897, N4221, N5005, N1288);
or OR3 (N8921, N8914, N8474, N611);
not NOT1 (N8922, N8918);
nor NOR4 (N8923, N8912, N46, N6891, N8810);
and AND4 (N8924, N8917, N3600, N6029, N4026);
buf BUF1 (N8925, N8907);
or OR4 (N8926, N8911, N1795, N3331, N2581);
nand NAND4 (N8927, N8919, N3375, N1645, N5327);
nand NAND4 (N8928, N8920, N2570, N7666, N1130);
xor XOR2 (N8929, N8926, N1661);
xor XOR2 (N8930, N8922, N3648);
not NOT1 (N8931, N8927);
nand NAND4 (N8932, N8925, N178, N3861, N8194);
or OR4 (N8933, N8923, N1355, N3406, N118);
nand NAND2 (N8934, N8932, N1898);
and AND4 (N8935, N8931, N7451, N8689, N117);
nand NAND3 (N8936, N8896, N1305, N5710);
buf BUF1 (N8937, N8935);
and AND3 (N8938, N8928, N1532, N8007);
or OR3 (N8939, N8913, N1453, N8620);
nand NAND3 (N8940, N8930, N671, N1986);
and AND4 (N8941, N8937, N7154, N4558, N3919);
buf BUF1 (N8942, N8941);
xor XOR2 (N8943, N8936, N4295);
and AND2 (N8944, N8943, N571);
nor NOR4 (N8945, N8933, N4745, N7996, N439);
xor XOR2 (N8946, N8944, N2378);
nand NAND3 (N8947, N8921, N1568, N2066);
and AND2 (N8948, N8946, N4905);
xor XOR2 (N8949, N8942, N8904);
nand NAND3 (N8950, N8924, N6490, N280);
nor NOR2 (N8951, N8950, N1729);
buf BUF1 (N8952, N8948);
buf BUF1 (N8953, N8952);
not NOT1 (N8954, N8945);
and AND4 (N8955, N8947, N2265, N5456, N2961);
and AND3 (N8956, N8940, N6212, N690);
nand NAND4 (N8957, N8939, N1771, N317, N8567);
buf BUF1 (N8958, N8949);
nand NAND4 (N8959, N8929, N8503, N1759, N8732);
and AND2 (N8960, N8956, N2066);
buf BUF1 (N8961, N8954);
xor XOR2 (N8962, N8957, N8301);
not NOT1 (N8963, N8934);
or OR3 (N8964, N8962, N6298, N7670);
nor NOR4 (N8965, N8953, N1304, N1772, N5568);
xor XOR2 (N8966, N8964, N3340);
buf BUF1 (N8967, N8965);
xor XOR2 (N8968, N8938, N4179);
not NOT1 (N8969, N8967);
or OR3 (N8970, N8961, N5125, N1021);
buf BUF1 (N8971, N8970);
xor XOR2 (N8972, N8959, N3094);
buf BUF1 (N8973, N8971);
xor XOR2 (N8974, N8960, N4524);
nor NOR3 (N8975, N8958, N168, N6937);
not NOT1 (N8976, N8975);
nor NOR3 (N8977, N8966, N6721, N3524);
buf BUF1 (N8978, N8973);
not NOT1 (N8979, N8976);
not NOT1 (N8980, N8972);
buf BUF1 (N8981, N8980);
xor XOR2 (N8982, N8969, N4722);
nor NOR3 (N8983, N8982, N5376, N2984);
and AND4 (N8984, N8977, N5827, N7859, N7326);
and AND3 (N8985, N8981, N6939, N5407);
nand NAND3 (N8986, N8963, N3605, N6753);
and AND4 (N8987, N8985, N1425, N4155, N6977);
or OR2 (N8988, N8974, N756);
buf BUF1 (N8989, N8986);
nor NOR4 (N8990, N8984, N466, N1237, N6049);
nor NOR4 (N8991, N8979, N8301, N758, N5758);
xor XOR2 (N8992, N8951, N2080);
buf BUF1 (N8993, N8978);
nor NOR2 (N8994, N8988, N3824);
not NOT1 (N8995, N8968);
nor NOR2 (N8996, N8990, N8245);
buf BUF1 (N8997, N8993);
buf BUF1 (N8998, N8983);
and AND3 (N8999, N8997, N8955, N4317);
nand NAND3 (N9000, N8872, N2678, N7486);
xor XOR2 (N9001, N8998, N3953);
buf BUF1 (N9002, N8996);
nand NAND4 (N9003, N8991, N4567, N614, N7736);
or OR3 (N9004, N9001, N6262, N5002);
or OR3 (N9005, N9000, N1840, N441);
xor XOR2 (N9006, N8999, N3537);
not NOT1 (N9007, N9004);
and AND3 (N9008, N9006, N1335, N1175);
nand NAND4 (N9009, N8992, N4047, N2973, N4416);
nand NAND2 (N9010, N9005, N4622);
buf BUF1 (N9011, N8995);
nand NAND2 (N9012, N9008, N5905);
xor XOR2 (N9013, N9003, N3837);
buf BUF1 (N9014, N8994);
nor NOR4 (N9015, N8987, N3185, N4012, N6713);
nor NOR3 (N9016, N9011, N239, N670);
or OR2 (N9017, N9012, N2611);
nor NOR2 (N9018, N8989, N975);
not NOT1 (N9019, N9002);
or OR2 (N9020, N9018, N5274);
buf BUF1 (N9021, N9020);
not NOT1 (N9022, N9010);
buf BUF1 (N9023, N9007);
and AND2 (N9024, N9019, N4211);
and AND2 (N9025, N9014, N1726);
not NOT1 (N9026, N9021);
buf BUF1 (N9027, N9017);
nand NAND4 (N9028, N9027, N1229, N5610, N7733);
not NOT1 (N9029, N9024);
and AND2 (N9030, N9023, N7728);
not NOT1 (N9031, N9013);
or OR2 (N9032, N9031, N4443);
buf BUF1 (N9033, N9030);
nand NAND3 (N9034, N9025, N4768, N3898);
or OR4 (N9035, N9026, N2273, N7767, N781);
and AND2 (N9036, N9028, N7816);
not NOT1 (N9037, N9034);
buf BUF1 (N9038, N9033);
or OR4 (N9039, N9035, N3693, N3023, N3844);
xor XOR2 (N9040, N9029, N1030);
buf BUF1 (N9041, N9038);
xor XOR2 (N9042, N9009, N2600);
xor XOR2 (N9043, N9039, N596);
xor XOR2 (N9044, N9015, N4912);
or OR4 (N9045, N9016, N5504, N5355, N2356);
buf BUF1 (N9046, N9032);
and AND3 (N9047, N9046, N6303, N8092);
xor XOR2 (N9048, N9042, N1324);
buf BUF1 (N9049, N9047);
xor XOR2 (N9050, N9041, N4788);
nand NAND2 (N9051, N9036, N8670);
not NOT1 (N9052, N9049);
nor NOR2 (N9053, N9040, N4754);
nand NAND2 (N9054, N9052, N5898);
xor XOR2 (N9055, N9022, N4320);
or OR2 (N9056, N9050, N2227);
xor XOR2 (N9057, N9044, N2862);
or OR3 (N9058, N9055, N2607, N4840);
or OR2 (N9059, N9053, N4836);
not NOT1 (N9060, N9056);
not NOT1 (N9061, N9054);
nor NOR3 (N9062, N9045, N9011, N6232);
or OR4 (N9063, N9060, N6410, N2644, N542);
nand NAND3 (N9064, N9061, N2022, N2046);
or OR4 (N9065, N9048, N4846, N6808, N5769);
nor NOR4 (N9066, N9043, N61, N4078, N3359);
buf BUF1 (N9067, N9062);
xor XOR2 (N9068, N9057, N4241);
nand NAND4 (N9069, N9037, N4596, N4437, N5049);
nand NAND2 (N9070, N9063, N4254);
buf BUF1 (N9071, N9067);
xor XOR2 (N9072, N9064, N341);
xor XOR2 (N9073, N9072, N8818);
not NOT1 (N9074, N9068);
and AND4 (N9075, N9059, N2289, N7305, N4458);
xor XOR2 (N9076, N9073, N1897);
and AND3 (N9077, N9051, N1716, N3783);
nand NAND4 (N9078, N9066, N719, N345, N2273);
nor NOR4 (N9079, N9074, N6517, N6535, N6292);
xor XOR2 (N9080, N9071, N9029);
xor XOR2 (N9081, N9058, N1535);
nand NAND2 (N9082, N9077, N249);
or OR2 (N9083, N9079, N2991);
not NOT1 (N9084, N9078);
nor NOR2 (N9085, N9081, N7546);
and AND3 (N9086, N9070, N3828, N7722);
buf BUF1 (N9087, N9083);
and AND2 (N9088, N9084, N4459);
buf BUF1 (N9089, N9088);
and AND3 (N9090, N9085, N1777, N4539);
and AND4 (N9091, N9069, N5205, N840, N5587);
nor NOR2 (N9092, N9089, N6167);
not NOT1 (N9093, N9091);
not NOT1 (N9094, N9092);
nor NOR3 (N9095, N9065, N1474, N5590);
nor NOR2 (N9096, N9095, N452);
nor NOR2 (N9097, N9082, N8920);
nor NOR3 (N9098, N9086, N2670, N7620);
xor XOR2 (N9099, N9094, N4374);
xor XOR2 (N9100, N9099, N5860);
and AND2 (N9101, N9093, N7909);
nand NAND3 (N9102, N9098, N1943, N6121);
buf BUF1 (N9103, N9075);
and AND2 (N9104, N9076, N5856);
nand NAND3 (N9105, N9101, N1353, N3569);
buf BUF1 (N9106, N9100);
or OR2 (N9107, N9105, N7477);
and AND3 (N9108, N9087, N5568, N7638);
or OR4 (N9109, N9103, N483, N3422, N2367);
xor XOR2 (N9110, N9090, N8157);
buf BUF1 (N9111, N9104);
nand NAND2 (N9112, N9107, N6949);
nor NOR4 (N9113, N9102, N2045, N3368, N3319);
buf BUF1 (N9114, N9111);
nor NOR2 (N9115, N9096, N3044);
nand NAND3 (N9116, N9080, N8360, N1275);
or OR3 (N9117, N9114, N2239, N2894);
or OR2 (N9118, N9106, N3293);
and AND3 (N9119, N9115, N7314, N4418);
and AND3 (N9120, N9118, N7507, N4468);
and AND4 (N9121, N9119, N2318, N4661, N3549);
nor NOR2 (N9122, N9112, N820);
or OR3 (N9123, N9120, N1405, N7045);
not NOT1 (N9124, N9110);
and AND4 (N9125, N9121, N5612, N2932, N7021);
or OR2 (N9126, N9108, N134);
and AND4 (N9127, N9125, N3770, N3946, N4995);
buf BUF1 (N9128, N9123);
nor NOR3 (N9129, N9122, N1498, N3280);
not NOT1 (N9130, N9124);
nor NOR3 (N9131, N9130, N8087, N7867);
xor XOR2 (N9132, N9126, N1595);
buf BUF1 (N9133, N9132);
nand NAND2 (N9134, N9131, N3466);
and AND3 (N9135, N9127, N9110, N8434);
nand NAND4 (N9136, N9113, N8790, N1447, N2712);
or OR2 (N9137, N9116, N5136);
or OR4 (N9138, N9133, N5737, N7008, N6754);
nand NAND2 (N9139, N9129, N7728);
nor NOR4 (N9140, N9137, N3162, N6700, N2742);
or OR2 (N9141, N9134, N4616);
xor XOR2 (N9142, N9135, N7585);
nand NAND3 (N9143, N9097, N527, N4299);
xor XOR2 (N9144, N9117, N6880);
and AND2 (N9145, N9143, N7248);
and AND4 (N9146, N9142, N882, N1377, N7150);
buf BUF1 (N9147, N9109);
or OR3 (N9148, N9139, N4392, N3211);
buf BUF1 (N9149, N9138);
or OR2 (N9150, N9145, N2221);
or OR3 (N9151, N9149, N1777, N1622);
nand NAND2 (N9152, N9144, N1547);
or OR2 (N9153, N9150, N2815);
nand NAND2 (N9154, N9136, N7914);
buf BUF1 (N9155, N9128);
not NOT1 (N9156, N9152);
buf BUF1 (N9157, N9155);
xor XOR2 (N9158, N9153, N4858);
not NOT1 (N9159, N9141);
nand NAND2 (N9160, N9156, N168);
and AND4 (N9161, N9160, N6560, N56, N6551);
xor XOR2 (N9162, N9148, N7457);
buf BUF1 (N9163, N9146);
xor XOR2 (N9164, N9162, N2751);
nand NAND2 (N9165, N9159, N2187);
not NOT1 (N9166, N9154);
or OR4 (N9167, N9166, N4339, N7029, N7378);
nor NOR4 (N9168, N9161, N6214, N7065, N2721);
buf BUF1 (N9169, N9164);
nand NAND4 (N9170, N9158, N2163, N2362, N5703);
or OR3 (N9171, N9169, N7377, N792);
nand NAND4 (N9172, N9170, N2718, N5813, N953);
nor NOR2 (N9173, N9151, N1436);
xor XOR2 (N9174, N9171, N384);
xor XOR2 (N9175, N9174, N8815);
or OR2 (N9176, N9165, N653);
and AND3 (N9177, N9168, N1758, N2586);
xor XOR2 (N9178, N9157, N6803);
nand NAND4 (N9179, N9167, N2939, N4258, N9069);
buf BUF1 (N9180, N9175);
nand NAND2 (N9181, N9180, N2789);
buf BUF1 (N9182, N9163);
or OR4 (N9183, N9176, N7145, N5267, N7034);
nand NAND4 (N9184, N9182, N3835, N4872, N5402);
nand NAND4 (N9185, N9178, N549, N8093, N9017);
nand NAND2 (N9186, N9177, N4765);
not NOT1 (N9187, N9173);
and AND3 (N9188, N9172, N1632, N141);
buf BUF1 (N9189, N9183);
and AND2 (N9190, N9147, N3901);
xor XOR2 (N9191, N9181, N7440);
xor XOR2 (N9192, N9186, N7230);
and AND2 (N9193, N9184, N953);
nor NOR3 (N9194, N9190, N1050, N4537);
or OR2 (N9195, N9179, N4012);
nand NAND4 (N9196, N9193, N5112, N8613, N6677);
xor XOR2 (N9197, N9140, N719);
and AND2 (N9198, N9195, N2984);
not NOT1 (N9199, N9185);
nor NOR4 (N9200, N9192, N4072, N4477, N2592);
nor NOR2 (N9201, N9187, N778);
nor NOR4 (N9202, N9194, N8173, N8513, N1304);
buf BUF1 (N9203, N9200);
buf BUF1 (N9204, N9196);
xor XOR2 (N9205, N9201, N6821);
or OR2 (N9206, N9188, N579);
or OR2 (N9207, N9206, N1713);
xor XOR2 (N9208, N9197, N2073);
nand NAND4 (N9209, N9191, N3589, N2357, N7612);
nand NAND3 (N9210, N9209, N1321, N2683);
nand NAND3 (N9211, N9203, N3327, N6987);
nand NAND2 (N9212, N9202, N5170);
not NOT1 (N9213, N9199);
nor NOR2 (N9214, N9212, N620);
buf BUF1 (N9215, N9207);
not NOT1 (N9216, N9189);
nor NOR2 (N9217, N9213, N3046);
nand NAND2 (N9218, N9215, N7113);
not NOT1 (N9219, N9205);
not NOT1 (N9220, N9214);
xor XOR2 (N9221, N9216, N8720);
xor XOR2 (N9222, N9217, N915);
nor NOR3 (N9223, N9220, N4343, N8986);
buf BUF1 (N9224, N9222);
not NOT1 (N9225, N9198);
xor XOR2 (N9226, N9204, N2071);
and AND2 (N9227, N9211, N7497);
or OR4 (N9228, N9224, N5263, N6788, N8597);
xor XOR2 (N9229, N9219, N9061);
or OR2 (N9230, N9229, N8871);
and AND3 (N9231, N9208, N5536, N3595);
nand NAND3 (N9232, N9210, N6744, N7824);
xor XOR2 (N9233, N9221, N6836);
not NOT1 (N9234, N9218);
and AND2 (N9235, N9230, N3806);
xor XOR2 (N9236, N9233, N3332);
nand NAND4 (N9237, N9227, N961, N8346, N1704);
nand NAND3 (N9238, N9231, N2500, N3586);
xor XOR2 (N9239, N9228, N45);
nor NOR2 (N9240, N9232, N5347);
nor NOR3 (N9241, N9236, N8301, N2676);
not NOT1 (N9242, N9240);
buf BUF1 (N9243, N9223);
nand NAND3 (N9244, N9226, N1649, N1158);
nand NAND4 (N9245, N9242, N7341, N7968, N8529);
or OR4 (N9246, N9244, N7261, N3726, N6749);
nand NAND4 (N9247, N9239, N3740, N5522, N710);
buf BUF1 (N9248, N9237);
nand NAND3 (N9249, N9243, N6241, N9018);
nor NOR3 (N9250, N9249, N667, N8565);
xor XOR2 (N9251, N9247, N8697);
xor XOR2 (N9252, N9235, N22);
xor XOR2 (N9253, N9225, N5933);
nor NOR3 (N9254, N9241, N7368, N5272);
nor NOR2 (N9255, N9246, N5423);
xor XOR2 (N9256, N9252, N4024);
and AND4 (N9257, N9251, N4779, N3300, N6578);
or OR2 (N9258, N9253, N8906);
xor XOR2 (N9259, N9248, N8256);
nand NAND2 (N9260, N9254, N3927);
or OR2 (N9261, N9259, N1525);
and AND2 (N9262, N9256, N2044);
or OR3 (N9263, N9238, N6089, N2313);
nor NOR2 (N9264, N9255, N1387);
buf BUF1 (N9265, N9263);
buf BUF1 (N9266, N9260);
xor XOR2 (N9267, N9234, N6737);
not NOT1 (N9268, N9264);
not NOT1 (N9269, N9266);
or OR2 (N9270, N9262, N3365);
nor NOR2 (N9271, N9270, N3104);
not NOT1 (N9272, N9250);
and AND4 (N9273, N9265, N1390, N2036, N1943);
nor NOR4 (N9274, N9267, N3070, N6434, N4706);
nor NOR4 (N9275, N9274, N364, N8239, N1690);
buf BUF1 (N9276, N9258);
and AND4 (N9277, N9272, N1992, N8877, N1604);
and AND2 (N9278, N9245, N3808);
xor XOR2 (N9279, N9273, N3203);
nand NAND2 (N9280, N9261, N4607);
or OR2 (N9281, N9278, N8130);
nor NOR3 (N9282, N9271, N2624, N7569);
nor NOR2 (N9283, N9280, N4751);
or OR2 (N9284, N9268, N4863);
not NOT1 (N9285, N9275);
nor NOR3 (N9286, N9281, N8863, N8679);
nand NAND2 (N9287, N9276, N1142);
buf BUF1 (N9288, N9284);
not NOT1 (N9289, N9283);
xor XOR2 (N9290, N9288, N1710);
not NOT1 (N9291, N9289);
buf BUF1 (N9292, N9257);
buf BUF1 (N9293, N9277);
and AND3 (N9294, N9269, N337, N5647);
xor XOR2 (N9295, N9293, N6524);
xor XOR2 (N9296, N9294, N4770);
xor XOR2 (N9297, N9282, N4349);
nand NAND3 (N9298, N9279, N7699, N7291);
not NOT1 (N9299, N9291);
and AND4 (N9300, N9292, N8795, N4401, N8225);
nor NOR4 (N9301, N9290, N3031, N1996, N4607);
nor NOR4 (N9302, N9298, N5315, N7765, N97);
xor XOR2 (N9303, N9295, N1458);
not NOT1 (N9304, N9299);
buf BUF1 (N9305, N9296);
nor NOR4 (N9306, N9303, N5202, N579, N2308);
nand NAND3 (N9307, N9301, N2712, N1782);
and AND2 (N9308, N9300, N4472);
nand NAND2 (N9309, N9287, N5075);
or OR4 (N9310, N9302, N7841, N4283, N3044);
nand NAND2 (N9311, N9286, N3502);
xor XOR2 (N9312, N9307, N4302);
nor NOR2 (N9313, N9304, N45);
buf BUF1 (N9314, N9310);
not NOT1 (N9315, N9305);
not NOT1 (N9316, N9285);
not NOT1 (N9317, N9315);
nor NOR3 (N9318, N9314, N5476, N1322);
and AND3 (N9319, N9313, N2778, N8549);
and AND4 (N9320, N9319, N520, N2627, N1028);
xor XOR2 (N9321, N9316, N5336);
and AND4 (N9322, N9306, N2657, N7751, N2478);
and AND2 (N9323, N9309, N8602);
xor XOR2 (N9324, N9312, N7368);
or OR2 (N9325, N9320, N4187);
nor NOR3 (N9326, N9297, N1169, N7922);
buf BUF1 (N9327, N9321);
and AND4 (N9328, N9311, N3244, N3995, N5021);
xor XOR2 (N9329, N9328, N6889);
xor XOR2 (N9330, N9329, N7313);
nor NOR4 (N9331, N9323, N6078, N3687, N9159);
not NOT1 (N9332, N9308);
xor XOR2 (N9333, N9327, N1899);
buf BUF1 (N9334, N9331);
or OR4 (N9335, N9326, N3531, N645, N2325);
buf BUF1 (N9336, N9322);
xor XOR2 (N9337, N9330, N2538);
nand NAND2 (N9338, N9333, N137);
not NOT1 (N9339, N9324);
and AND4 (N9340, N9325, N2656, N4654, N3690);
nor NOR3 (N9341, N9335, N3806, N3583);
buf BUF1 (N9342, N9337);
xor XOR2 (N9343, N9334, N2409);
buf BUF1 (N9344, N9336);
not NOT1 (N9345, N9318);
xor XOR2 (N9346, N9332, N6534);
nand NAND4 (N9347, N9339, N4835, N4830, N2360);
buf BUF1 (N9348, N9347);
nand NAND2 (N9349, N9348, N2279);
and AND4 (N9350, N9340, N8272, N8219, N2359);
nand NAND3 (N9351, N9350, N2243, N6620);
nor NOR3 (N9352, N9349, N381, N6162);
not NOT1 (N9353, N9342);
and AND3 (N9354, N9344, N6094, N540);
nor NOR3 (N9355, N9346, N2713, N7247);
xor XOR2 (N9356, N9317, N1669);
or OR4 (N9357, N9352, N6737, N3718, N624);
xor XOR2 (N9358, N9343, N7298);
and AND3 (N9359, N9351, N1556, N580);
or OR2 (N9360, N9357, N651);
nand NAND4 (N9361, N9355, N5467, N2763, N2818);
and AND3 (N9362, N9361, N931, N1289);
xor XOR2 (N9363, N9356, N1967);
xor XOR2 (N9364, N9341, N345);
or OR3 (N9365, N9354, N6423, N6050);
nor NOR4 (N9366, N9362, N2005, N5100, N4335);
or OR2 (N9367, N9366, N6943);
xor XOR2 (N9368, N9363, N2905);
buf BUF1 (N9369, N9364);
xor XOR2 (N9370, N9367, N2492);
and AND3 (N9371, N9360, N2432, N9351);
nand NAND2 (N9372, N9338, N7990);
xor XOR2 (N9373, N9372, N593);
buf BUF1 (N9374, N9369);
nor NOR4 (N9375, N9374, N5506, N8076, N7166);
xor XOR2 (N9376, N9353, N3445);
nor NOR4 (N9377, N9345, N6201, N9065, N4855);
not NOT1 (N9378, N9375);
and AND3 (N9379, N9358, N5889, N2741);
and AND3 (N9380, N9378, N7962, N7228);
buf BUF1 (N9381, N9359);
nor NOR3 (N9382, N9373, N2761, N5066);
nand NAND4 (N9383, N9365, N5782, N7079, N2096);
buf BUF1 (N9384, N9383);
not NOT1 (N9385, N9377);
xor XOR2 (N9386, N9370, N2947);
and AND3 (N9387, N9368, N8748, N346);
buf BUF1 (N9388, N9387);
nand NAND4 (N9389, N9379, N1784, N7980, N7144);
and AND4 (N9390, N9381, N2325, N9264, N1153);
not NOT1 (N9391, N9388);
buf BUF1 (N9392, N9391);
or OR3 (N9393, N9371, N6470, N846);
buf BUF1 (N9394, N9386);
and AND4 (N9395, N9392, N4214, N1763, N9281);
not NOT1 (N9396, N9395);
nand NAND3 (N9397, N9393, N1074, N7747);
not NOT1 (N9398, N9382);
or OR4 (N9399, N9398, N7031, N1705, N9218);
buf BUF1 (N9400, N9396);
or OR3 (N9401, N9380, N2175, N8586);
and AND4 (N9402, N9390, N6662, N1102, N4623);
buf BUF1 (N9403, N9385);
xor XOR2 (N9404, N9400, N3738);
not NOT1 (N9405, N9399);
not NOT1 (N9406, N9403);
not NOT1 (N9407, N9402);
xor XOR2 (N9408, N9405, N2466);
buf BUF1 (N9409, N9407);
xor XOR2 (N9410, N9409, N3400);
buf BUF1 (N9411, N9406);
xor XOR2 (N9412, N9401, N8573);
not NOT1 (N9413, N9376);
buf BUF1 (N9414, N9384);
not NOT1 (N9415, N9411);
xor XOR2 (N9416, N9412, N450);
nor NOR3 (N9417, N9389, N2131, N2072);
xor XOR2 (N9418, N9415, N2993);
and AND4 (N9419, N9410, N9080, N2022, N4781);
xor XOR2 (N9420, N9417, N795);
and AND3 (N9421, N9419, N4815, N1591);
xor XOR2 (N9422, N9408, N4445);
nor NOR3 (N9423, N9420, N281, N6048);
or OR2 (N9424, N9423, N1122);
buf BUF1 (N9425, N9422);
buf BUF1 (N9426, N9397);
not NOT1 (N9427, N9413);
nand NAND3 (N9428, N9394, N735, N1680);
or OR4 (N9429, N9425, N6903, N2355, N8875);
nand NAND2 (N9430, N9404, N7425);
not NOT1 (N9431, N9427);
xor XOR2 (N9432, N9421, N7406);
and AND3 (N9433, N9432, N842, N7003);
or OR3 (N9434, N9414, N9377, N846);
not NOT1 (N9435, N9418);
buf BUF1 (N9436, N9429);
nand NAND3 (N9437, N9416, N1464, N8741);
not NOT1 (N9438, N9424);
or OR3 (N9439, N9437, N2960, N7859);
not NOT1 (N9440, N9426);
buf BUF1 (N9441, N9433);
and AND4 (N9442, N9435, N3097, N5741, N724);
or OR4 (N9443, N9440, N4573, N4021, N6223);
not NOT1 (N9444, N9428);
nand NAND4 (N9445, N9444, N8614, N7408, N3706);
nor NOR4 (N9446, N9443, N2564, N8164, N6331);
xor XOR2 (N9447, N9430, N56);
nand NAND2 (N9448, N9445, N7730);
or OR4 (N9449, N9438, N6197, N1881, N3233);
or OR3 (N9450, N9448, N7819, N2062);
nand NAND2 (N9451, N9436, N3745);
not NOT1 (N9452, N9442);
nand NAND2 (N9453, N9439, N2622);
nor NOR2 (N9454, N9431, N6574);
not NOT1 (N9455, N9441);
nor NOR3 (N9456, N9451, N580, N18);
buf BUF1 (N9457, N9446);
buf BUF1 (N9458, N9454);
xor XOR2 (N9459, N9456, N6620);
and AND2 (N9460, N9457, N9427);
and AND4 (N9461, N9450, N5012, N1686, N1489);
nor NOR3 (N9462, N9447, N6320, N7100);
and AND2 (N9463, N9459, N3189);
nand NAND3 (N9464, N9460, N7993, N5942);
or OR4 (N9465, N9455, N9455, N1087, N2438);
or OR2 (N9466, N9452, N9097);
or OR3 (N9467, N9462, N5318, N3575);
buf BUF1 (N9468, N9453);
not NOT1 (N9469, N9458);
not NOT1 (N9470, N9466);
not NOT1 (N9471, N9470);
nand NAND3 (N9472, N9471, N2744, N1623);
xor XOR2 (N9473, N9449, N7794);
and AND2 (N9474, N9465, N6582);
and AND3 (N9475, N9473, N5769, N4985);
buf BUF1 (N9476, N9461);
xor XOR2 (N9477, N9464, N2814);
nand NAND4 (N9478, N9463, N9188, N9477, N8173);
and AND4 (N9479, N8674, N8117, N1861, N8853);
or OR4 (N9480, N9467, N2999, N7547, N225);
or OR2 (N9481, N9478, N9324);
or OR4 (N9482, N9480, N5454, N6521, N9145);
not NOT1 (N9483, N9472);
or OR3 (N9484, N9434, N2186, N7569);
buf BUF1 (N9485, N9468);
nand NAND2 (N9486, N9474, N5045);
nand NAND3 (N9487, N9483, N4808, N7163);
not NOT1 (N9488, N9487);
nor NOR2 (N9489, N9475, N7132);
nand NAND2 (N9490, N9476, N2248);
buf BUF1 (N9491, N9488);
or OR3 (N9492, N9469, N5468, N6903);
not NOT1 (N9493, N9481);
not NOT1 (N9494, N9482);
not NOT1 (N9495, N9492);
and AND3 (N9496, N9490, N2053, N623);
not NOT1 (N9497, N9493);
and AND4 (N9498, N9491, N7111, N3730, N8841);
not NOT1 (N9499, N9494);
not NOT1 (N9500, N9489);
nand NAND3 (N9501, N9479, N2333, N9301);
nor NOR4 (N9502, N9500, N450, N4994, N5209);
and AND4 (N9503, N9496, N7932, N6316, N4972);
nor NOR2 (N9504, N9501, N8254);
xor XOR2 (N9505, N9499, N3848);
nor NOR4 (N9506, N9495, N1248, N2657, N1172);
nor NOR2 (N9507, N9502, N1425);
nand NAND4 (N9508, N9506, N9341, N318, N5940);
or OR2 (N9509, N9508, N3444);
or OR4 (N9510, N9507, N4453, N7603, N66);
not NOT1 (N9511, N9509);
not NOT1 (N9512, N9485);
or OR4 (N9513, N9505, N266, N1576, N3022);
nor NOR3 (N9514, N9497, N6420, N2801);
or OR2 (N9515, N9510, N3262);
buf BUF1 (N9516, N9486);
buf BUF1 (N9517, N9498);
xor XOR2 (N9518, N9513, N8565);
not NOT1 (N9519, N9516);
or OR3 (N9520, N9518, N5377, N8260);
nand NAND3 (N9521, N9504, N2062, N6581);
not NOT1 (N9522, N9512);
or OR4 (N9523, N9511, N1823, N2628, N420);
or OR2 (N9524, N9503, N266);
buf BUF1 (N9525, N9520);
not NOT1 (N9526, N9521);
and AND2 (N9527, N9515, N7063);
nand NAND3 (N9528, N9519, N6045, N3658);
buf BUF1 (N9529, N9523);
nand NAND4 (N9530, N9528, N7347, N7590, N8663);
buf BUF1 (N9531, N9530);
not NOT1 (N9532, N9484);
and AND2 (N9533, N9531, N9061);
buf BUF1 (N9534, N9533);
nor NOR3 (N9535, N9527, N4363, N362);
nor NOR3 (N9536, N9514, N1846, N7303);
nor NOR4 (N9537, N9529, N2663, N2938, N3452);
and AND4 (N9538, N9526, N7296, N4436, N2428);
nand NAND2 (N9539, N9532, N2092);
xor XOR2 (N9540, N9522, N240);
nand NAND2 (N9541, N9535, N3838);
buf BUF1 (N9542, N9525);
and AND3 (N9543, N9537, N8154, N1836);
not NOT1 (N9544, N9541);
and AND2 (N9545, N9524, N5138);
nor NOR3 (N9546, N9540, N8705, N4074);
and AND4 (N9547, N9545, N2200, N8138, N8568);
not NOT1 (N9548, N9534);
nor NOR3 (N9549, N9538, N7286, N8079);
and AND2 (N9550, N9543, N2075);
xor XOR2 (N9551, N9550, N6616);
and AND3 (N9552, N9548, N1217, N3171);
xor XOR2 (N9553, N9542, N4283);
nand NAND3 (N9554, N9539, N1806, N163);
not NOT1 (N9555, N9546);
xor XOR2 (N9556, N9551, N2261);
not NOT1 (N9557, N9552);
nand NAND3 (N9558, N9554, N9552, N8970);
nor NOR3 (N9559, N9555, N6333, N9105);
not NOT1 (N9560, N9517);
nor NOR3 (N9561, N9553, N76, N5115);
buf BUF1 (N9562, N9560);
and AND4 (N9563, N9556, N9453, N9072, N1521);
nand NAND2 (N9564, N9563, N4766);
nand NAND2 (N9565, N9557, N2505);
nand NAND3 (N9566, N9547, N2264, N4449);
nand NAND4 (N9567, N9558, N3137, N8478, N6114);
nand NAND3 (N9568, N9544, N4670, N4582);
or OR3 (N9569, N9568, N6688, N6150);
xor XOR2 (N9570, N9561, N2668);
nor NOR3 (N9571, N9565, N8844, N4629);
xor XOR2 (N9572, N9569, N7753);
xor XOR2 (N9573, N9570, N6783);
nor NOR2 (N9574, N9566, N7531);
or OR3 (N9575, N9536, N9467, N6605);
or OR4 (N9576, N9575, N2584, N4451, N613);
not NOT1 (N9577, N9574);
or OR4 (N9578, N9573, N4514, N7156, N4333);
nor NOR2 (N9579, N9577, N6997);
and AND4 (N9580, N9572, N7842, N3219, N3249);
and AND2 (N9581, N9562, N7716);
buf BUF1 (N9582, N9578);
not NOT1 (N9583, N9580);
not NOT1 (N9584, N9583);
nor NOR4 (N9585, N9549, N2827, N4000, N964);
or OR2 (N9586, N9576, N75);
xor XOR2 (N9587, N9586, N1700);
nor NOR3 (N9588, N9571, N3407, N2950);
xor XOR2 (N9589, N9559, N8108);
buf BUF1 (N9590, N9585);
and AND3 (N9591, N9587, N5457, N2180);
not NOT1 (N9592, N9567);
nor NOR3 (N9593, N9582, N6647, N4733);
and AND2 (N9594, N9589, N6132);
or OR3 (N9595, N9564, N9458, N6982);
nor NOR4 (N9596, N9584, N4614, N7717, N6428);
xor XOR2 (N9597, N9579, N85);
and AND2 (N9598, N9597, N3073);
nor NOR2 (N9599, N9593, N2822);
nand NAND4 (N9600, N9595, N177, N3981, N9497);
xor XOR2 (N9601, N9581, N8033);
nand NAND4 (N9602, N9600, N5013, N9506, N3748);
xor XOR2 (N9603, N9590, N8259);
nand NAND2 (N9604, N9603, N8597);
nor NOR4 (N9605, N9592, N8720, N8979, N303);
buf BUF1 (N9606, N9605);
buf BUF1 (N9607, N9598);
buf BUF1 (N9608, N9606);
nand NAND2 (N9609, N9588, N5214);
nand NAND4 (N9610, N9596, N3224, N2050, N4817);
or OR2 (N9611, N9604, N6948);
buf BUF1 (N9612, N9608);
not NOT1 (N9613, N9609);
buf BUF1 (N9614, N9612);
not NOT1 (N9615, N9591);
buf BUF1 (N9616, N9611);
nor NOR4 (N9617, N9594, N4791, N7224, N3522);
or OR3 (N9618, N9616, N5592, N8374);
nand NAND3 (N9619, N9610, N7944, N6466);
xor XOR2 (N9620, N9601, N6623);
xor XOR2 (N9621, N9619, N5191);
buf BUF1 (N9622, N9607);
or OR2 (N9623, N9615, N3141);
or OR2 (N9624, N9614, N177);
or OR4 (N9625, N9621, N7126, N7581, N8585);
buf BUF1 (N9626, N9618);
nor NOR3 (N9627, N9623, N3686, N2043);
nand NAND2 (N9628, N9627, N8988);
nand NAND2 (N9629, N9622, N1291);
or OR3 (N9630, N9617, N2650, N8002);
nor NOR2 (N9631, N9626, N3911);
not NOT1 (N9632, N9630);
nor NOR3 (N9633, N9632, N7575, N5447);
buf BUF1 (N9634, N9620);
or OR2 (N9635, N9634, N1914);
buf BUF1 (N9636, N9602);
xor XOR2 (N9637, N9628, N5056);
and AND3 (N9638, N9599, N6366, N2749);
not NOT1 (N9639, N9613);
or OR4 (N9640, N9625, N3880, N6853, N9637);
not NOT1 (N9641, N1938);
not NOT1 (N9642, N9633);
xor XOR2 (N9643, N9636, N4410);
and AND4 (N9644, N9638, N2124, N6040, N688);
xor XOR2 (N9645, N9643, N3594);
xor XOR2 (N9646, N9640, N8311);
and AND4 (N9647, N9624, N7506, N4150, N8087);
or OR3 (N9648, N9644, N3214, N7852);
nand NAND2 (N9649, N9631, N7769);
nor NOR3 (N9650, N9641, N4855, N196);
not NOT1 (N9651, N9629);
nand NAND4 (N9652, N9651, N219, N8339, N9074);
buf BUF1 (N9653, N9649);
buf BUF1 (N9654, N9653);
and AND2 (N9655, N9639, N4043);
or OR2 (N9656, N9642, N4508);
nor NOR4 (N9657, N9655, N5400, N205, N4101);
buf BUF1 (N9658, N9635);
not NOT1 (N9659, N9656);
not NOT1 (N9660, N9659);
nand NAND4 (N9661, N9645, N1660, N7999, N3483);
xor XOR2 (N9662, N9648, N5001);
buf BUF1 (N9663, N9646);
not NOT1 (N9664, N9660);
nor NOR3 (N9665, N9652, N1058, N3117);
nand NAND3 (N9666, N9647, N203, N5228);
buf BUF1 (N9667, N9654);
buf BUF1 (N9668, N9663);
nand NAND4 (N9669, N9650, N2878, N2542, N6956);
nand NAND3 (N9670, N9669, N6689, N5505);
buf BUF1 (N9671, N9665);
xor XOR2 (N9672, N9668, N8243);
or OR3 (N9673, N9664, N1783, N4773);
buf BUF1 (N9674, N9670);
nor NOR3 (N9675, N9662, N2763, N8041);
nand NAND3 (N9676, N9673, N525, N6466);
buf BUF1 (N9677, N9661);
xor XOR2 (N9678, N9666, N7253);
or OR3 (N9679, N9676, N1435, N4637);
or OR3 (N9680, N9678, N3050, N8834);
nand NAND4 (N9681, N9671, N7542, N8227, N4160);
not NOT1 (N9682, N9672);
buf BUF1 (N9683, N9674);
not NOT1 (N9684, N9681);
nand NAND2 (N9685, N9675, N6818);
buf BUF1 (N9686, N9685);
or OR2 (N9687, N9667, N7945);
not NOT1 (N9688, N9657);
not NOT1 (N9689, N9686);
and AND3 (N9690, N9680, N6360, N3708);
not NOT1 (N9691, N9682);
and AND2 (N9692, N9684, N4209);
nor NOR3 (N9693, N9692, N8316, N2303);
xor XOR2 (N9694, N9690, N770);
and AND4 (N9695, N9691, N3471, N6012, N6508);
and AND2 (N9696, N9683, N4055);
or OR2 (N9697, N9694, N4027);
buf BUF1 (N9698, N9687);
nand NAND3 (N9699, N9698, N192, N4094);
or OR3 (N9700, N9693, N1998, N5898);
not NOT1 (N9701, N9689);
not NOT1 (N9702, N9688);
and AND2 (N9703, N9679, N5399);
or OR3 (N9704, N9699, N769, N5795);
buf BUF1 (N9705, N9658);
or OR4 (N9706, N9697, N7792, N5583, N4029);
or OR2 (N9707, N9677, N4470);
and AND3 (N9708, N9696, N8627, N9203);
nor NOR3 (N9709, N9695, N8504, N2502);
nand NAND4 (N9710, N9704, N1303, N7201, N4897);
nand NAND4 (N9711, N9707, N7398, N4796, N8784);
or OR3 (N9712, N9705, N9325, N1554);
not NOT1 (N9713, N9711);
not NOT1 (N9714, N9708);
nor NOR4 (N9715, N9701, N4120, N3006, N860);
nor NOR2 (N9716, N9703, N1160);
buf BUF1 (N9717, N9709);
not NOT1 (N9718, N9710);
nand NAND2 (N9719, N9713, N753);
xor XOR2 (N9720, N9719, N6848);
and AND3 (N9721, N9716, N800, N1546);
and AND4 (N9722, N9720, N2270, N1749, N1222);
not NOT1 (N9723, N9721);
not NOT1 (N9724, N9706);
buf BUF1 (N9725, N9712);
and AND2 (N9726, N9715, N2936);
xor XOR2 (N9727, N9702, N8460);
buf BUF1 (N9728, N9717);
buf BUF1 (N9729, N9723);
nand NAND3 (N9730, N9714, N6911, N7476);
nor NOR3 (N9731, N9727, N7901, N5069);
buf BUF1 (N9732, N9728);
not NOT1 (N9733, N9732);
buf BUF1 (N9734, N9733);
nor NOR4 (N9735, N9718, N7298, N3863, N6449);
buf BUF1 (N9736, N9724);
nand NAND4 (N9737, N9736, N2568, N1366, N6761);
not NOT1 (N9738, N9700);
nor NOR3 (N9739, N9734, N7754, N9432);
nand NAND2 (N9740, N9726, N4644);
buf BUF1 (N9741, N9738);
nor NOR2 (N9742, N9741, N8139);
and AND3 (N9743, N9740, N9418, N906);
buf BUF1 (N9744, N9729);
not NOT1 (N9745, N9730);
buf BUF1 (N9746, N9725);
nand NAND4 (N9747, N9722, N6374, N5868, N4954);
nand NAND2 (N9748, N9743, N6152);
nor NOR2 (N9749, N9731, N7106);
xor XOR2 (N9750, N9746, N9724);
and AND3 (N9751, N9737, N1512, N3736);
buf BUF1 (N9752, N9747);
nand NAND2 (N9753, N9749, N1554);
buf BUF1 (N9754, N9739);
not NOT1 (N9755, N9751);
and AND4 (N9756, N9744, N3540, N3295, N1130);
or OR4 (N9757, N9748, N8646, N1505, N6406);
and AND3 (N9758, N9754, N6091, N1046);
nand NAND3 (N9759, N9745, N7819, N7173);
and AND4 (N9760, N9742, N9018, N4757, N7378);
and AND4 (N9761, N9756, N1570, N3468, N6426);
nand NAND4 (N9762, N9735, N1114, N763, N5513);
and AND2 (N9763, N9753, N3511);
not NOT1 (N9764, N9758);
xor XOR2 (N9765, N9761, N643);
not NOT1 (N9766, N9762);
nand NAND3 (N9767, N9755, N4676, N8138);
and AND3 (N9768, N9760, N9462, N1440);
and AND4 (N9769, N9767, N8375, N1978, N6039);
and AND3 (N9770, N9766, N1450, N8715);
buf BUF1 (N9771, N9750);
xor XOR2 (N9772, N9752, N3386);
or OR4 (N9773, N9765, N7238, N4888, N2995);
nor NOR4 (N9774, N9763, N3131, N1681, N2969);
or OR4 (N9775, N9757, N8552, N4981, N9344);
nor NOR4 (N9776, N9769, N7941, N6172, N8774);
not NOT1 (N9777, N9776);
xor XOR2 (N9778, N9771, N5065);
xor XOR2 (N9779, N9759, N8342);
nor NOR3 (N9780, N9772, N5279, N5295);
nor NOR2 (N9781, N9778, N1506);
buf BUF1 (N9782, N9781);
and AND4 (N9783, N9770, N2588, N9639, N8085);
not NOT1 (N9784, N9774);
xor XOR2 (N9785, N9768, N4346);
nand NAND2 (N9786, N9764, N7259);
nand NAND4 (N9787, N9779, N4990, N3684, N3823);
nor NOR3 (N9788, N9787, N4787, N4523);
not NOT1 (N9789, N9775);
xor XOR2 (N9790, N9786, N7093);
or OR2 (N9791, N9780, N6284);
or OR3 (N9792, N9784, N9622, N7557);
or OR2 (N9793, N9791, N2934);
xor XOR2 (N9794, N9782, N1088);
or OR2 (N9795, N9793, N8380);
buf BUF1 (N9796, N9777);
buf BUF1 (N9797, N9790);
not NOT1 (N9798, N9783);
and AND4 (N9799, N9785, N5809, N4521, N228);
buf BUF1 (N9800, N9789);
buf BUF1 (N9801, N9798);
xor XOR2 (N9802, N9792, N5078);
xor XOR2 (N9803, N9800, N943);
buf BUF1 (N9804, N9799);
not NOT1 (N9805, N9804);
xor XOR2 (N9806, N9794, N657);
not NOT1 (N9807, N9796);
and AND4 (N9808, N9788, N2761, N1181, N1973);
and AND4 (N9809, N9806, N6629, N3753, N179);
nor NOR3 (N9810, N9795, N1391, N6485);
nand NAND2 (N9811, N9803, N9473);
buf BUF1 (N9812, N9810);
nand NAND3 (N9813, N9808, N1703, N8632);
or OR4 (N9814, N9813, N5991, N2910, N9136);
or OR4 (N9815, N9809, N2541, N2808, N4742);
nand NAND2 (N9816, N9812, N5510);
buf BUF1 (N9817, N9802);
nand NAND2 (N9818, N9816, N3327);
xor XOR2 (N9819, N9815, N8101);
and AND4 (N9820, N9801, N2686, N6420, N6185);
nand NAND4 (N9821, N9811, N8821, N8623, N2287);
nor NOR4 (N9822, N9819, N2435, N4365, N596);
nor NOR4 (N9823, N9820, N8229, N5725, N1953);
not NOT1 (N9824, N9805);
and AND3 (N9825, N9821, N4041, N8054);
nor NOR2 (N9826, N9817, N377);
not NOT1 (N9827, N9797);
xor XOR2 (N9828, N9823, N1890);
buf BUF1 (N9829, N9814);
or OR2 (N9830, N9822, N5515);
or OR4 (N9831, N9825, N1268, N8298, N6329);
nor NOR2 (N9832, N9826, N6561);
or OR3 (N9833, N9807, N7626, N1240);
or OR4 (N9834, N9831, N849, N5640, N7026);
nand NAND2 (N9835, N9830, N4690);
xor XOR2 (N9836, N9833, N8960);
xor XOR2 (N9837, N9828, N2449);
nor NOR2 (N9838, N9827, N9040);
buf BUF1 (N9839, N9818);
buf BUF1 (N9840, N9834);
buf BUF1 (N9841, N9839);
and AND4 (N9842, N9837, N9043, N4279, N7996);
xor XOR2 (N9843, N9842, N4994);
not NOT1 (N9844, N9832);
not NOT1 (N9845, N9844);
xor XOR2 (N9846, N9836, N6259);
or OR2 (N9847, N9829, N8299);
and AND3 (N9848, N9843, N4121, N7977);
and AND2 (N9849, N9773, N7240);
buf BUF1 (N9850, N9824);
xor XOR2 (N9851, N9838, N2226);
nand NAND4 (N9852, N9835, N1213, N4489, N1486);
xor XOR2 (N9853, N9846, N6055);
and AND2 (N9854, N9840, N60);
buf BUF1 (N9855, N9849);
nor NOR2 (N9856, N9855, N5885);
or OR2 (N9857, N9853, N274);
nor NOR4 (N9858, N9847, N1405, N168, N4850);
buf BUF1 (N9859, N9856);
and AND4 (N9860, N9858, N6574, N374, N8795);
not NOT1 (N9861, N9857);
nand NAND2 (N9862, N9848, N9746);
nor NOR4 (N9863, N9854, N2667, N9241, N7672);
and AND3 (N9864, N9851, N9391, N4299);
nand NAND4 (N9865, N9850, N968, N963, N6990);
buf BUF1 (N9866, N9865);
and AND3 (N9867, N9845, N9685, N5949);
not NOT1 (N9868, N9863);
and AND4 (N9869, N9852, N5241, N5870, N6712);
buf BUF1 (N9870, N9867);
buf BUF1 (N9871, N9870);
not NOT1 (N9872, N9871);
not NOT1 (N9873, N9860);
and AND4 (N9874, N9862, N9629, N138, N8849);
nor NOR4 (N9875, N9861, N6919, N6666, N7696);
not NOT1 (N9876, N9841);
not NOT1 (N9877, N9873);
or OR3 (N9878, N9868, N4828, N1237);
or OR3 (N9879, N9874, N5146, N3571);
xor XOR2 (N9880, N9869, N5123);
nand NAND3 (N9881, N9864, N4363, N8416);
xor XOR2 (N9882, N9872, N7779);
or OR3 (N9883, N9875, N4884, N2609);
and AND3 (N9884, N9883, N3268, N8247);
not NOT1 (N9885, N9884);
nor NOR4 (N9886, N9881, N5092, N1971, N3304);
not NOT1 (N9887, N9876);
and AND4 (N9888, N9887, N2737, N1967, N290);
nand NAND2 (N9889, N9885, N8598);
buf BUF1 (N9890, N9878);
nand NAND4 (N9891, N9890, N2615, N7189, N9224);
nand NAND4 (N9892, N9882, N243, N1062, N7604);
or OR4 (N9893, N9879, N8288, N9092, N7254);
nor NOR4 (N9894, N9880, N5495, N6911, N6313);
nor NOR4 (N9895, N9889, N5431, N1752, N3919);
nor NOR3 (N9896, N9891, N5414, N7640);
nand NAND3 (N9897, N9892, N2082, N8639);
or OR4 (N9898, N9896, N3553, N7324, N3784);
and AND3 (N9899, N9898, N9689, N2908);
nand NAND4 (N9900, N9893, N6657, N3674, N6239);
and AND3 (N9901, N9897, N6252, N8323);
xor XOR2 (N9902, N9895, N6270);
nor NOR4 (N9903, N9866, N6719, N7203, N2723);
and AND4 (N9904, N9901, N1651, N3535, N4201);
nand NAND4 (N9905, N9904, N6799, N2680, N5165);
xor XOR2 (N9906, N9903, N3467);
or OR4 (N9907, N9900, N9204, N5486, N1531);
nor NOR3 (N9908, N9886, N4354, N4608);
nor NOR3 (N9909, N9907, N9206, N6229);
buf BUF1 (N9910, N9877);
buf BUF1 (N9911, N9888);
nor NOR4 (N9912, N9902, N3952, N3495, N6087);
nor NOR3 (N9913, N9899, N9287, N9004);
nand NAND4 (N9914, N9859, N3562, N709, N2157);
not NOT1 (N9915, N9913);
buf BUF1 (N9916, N9912);
not NOT1 (N9917, N9908);
buf BUF1 (N9918, N9915);
nand NAND3 (N9919, N9918, N9427, N2145);
not NOT1 (N9920, N9911);
nor NOR3 (N9921, N9917, N3332, N205);
nor NOR3 (N9922, N9905, N3408, N3250);
not NOT1 (N9923, N9909);
nor NOR4 (N9924, N9906, N9151, N5475, N9908);
xor XOR2 (N9925, N9914, N9438);
nor NOR3 (N9926, N9925, N7515, N6012);
buf BUF1 (N9927, N9921);
not NOT1 (N9928, N9923);
not NOT1 (N9929, N9926);
nor NOR3 (N9930, N9894, N5182, N3922);
xor XOR2 (N9931, N9927, N6339);
and AND2 (N9932, N9931, N5415);
xor XOR2 (N9933, N9910, N4163);
and AND3 (N9934, N9929, N3289, N3006);
xor XOR2 (N9935, N9922, N724);
not NOT1 (N9936, N9919);
not NOT1 (N9937, N9930);
xor XOR2 (N9938, N9935, N5994);
or OR4 (N9939, N9932, N7482, N8410, N4172);
or OR4 (N9940, N9938, N1418, N2722, N3941);
buf BUF1 (N9941, N9939);
nand NAND3 (N9942, N9933, N7858, N3172);
and AND3 (N9943, N9928, N8526, N923);
not NOT1 (N9944, N9924);
not NOT1 (N9945, N9937);
and AND4 (N9946, N9941, N4305, N6956, N4615);
buf BUF1 (N9947, N9916);
or OR2 (N9948, N9920, N8925);
or OR2 (N9949, N9942, N7261);
not NOT1 (N9950, N9944);
buf BUF1 (N9951, N9946);
and AND4 (N9952, N9950, N3452, N4679, N1309);
buf BUF1 (N9953, N9952);
nand NAND4 (N9954, N9951, N157, N2159, N4680);
nand NAND3 (N9955, N9936, N7646, N9246);
and AND2 (N9956, N9943, N7311);
nand NAND4 (N9957, N9934, N8429, N1616, N3796);
buf BUF1 (N9958, N9957);
nand NAND3 (N9959, N9953, N834, N7783);
or OR2 (N9960, N9945, N7740);
xor XOR2 (N9961, N9956, N97);
xor XOR2 (N9962, N9959, N7222);
nand NAND3 (N9963, N9960, N9766, N9676);
nor NOR4 (N9964, N9955, N1829, N7027, N3684);
or OR2 (N9965, N9958, N5097);
nor NOR3 (N9966, N9947, N7985, N9363);
buf BUF1 (N9967, N9963);
nand NAND4 (N9968, N9949, N2215, N4696, N7191);
xor XOR2 (N9969, N9962, N38);
or OR3 (N9970, N9965, N128, N7078);
nand NAND3 (N9971, N9940, N3141, N2072);
buf BUF1 (N9972, N9966);
nor NOR3 (N9973, N9972, N1245, N2638);
xor XOR2 (N9974, N9961, N8760);
and AND4 (N9975, N9974, N7890, N7073, N3859);
not NOT1 (N9976, N9971);
and AND4 (N9977, N9970, N3789, N1600, N7625);
not NOT1 (N9978, N9964);
or OR4 (N9979, N9948, N6455, N205, N1761);
nor NOR2 (N9980, N9976, N5541);
or OR3 (N9981, N9968, N4960, N2047);
buf BUF1 (N9982, N9975);
not NOT1 (N9983, N9973);
buf BUF1 (N9984, N9977);
or OR3 (N9985, N9981, N3777, N1246);
or OR3 (N9986, N9980, N5347, N7175);
not NOT1 (N9987, N9984);
buf BUF1 (N9988, N9983);
not NOT1 (N9989, N9978);
and AND2 (N9990, N9982, N5873);
nand NAND4 (N9991, N9990, N5195, N230, N378);
or OR2 (N9992, N9967, N1173);
not NOT1 (N9993, N9989);
or OR2 (N9994, N9991, N677);
or OR2 (N9995, N9993, N3268);
xor XOR2 (N9996, N9954, N3824);
not NOT1 (N9997, N9988);
buf BUF1 (N9998, N9997);
or OR3 (N9999, N9987, N5523, N8874);
nand NAND2 (N10000, N9998, N5326);
buf BUF1 (N10001, N9994);
buf BUF1 (N10002, N9986);
xor XOR2 (N10003, N9999, N920);
xor XOR2 (N10004, N10001, N3663);
or OR3 (N10005, N9996, N7301, N4041);
and AND2 (N10006, N9995, N920);
buf BUF1 (N10007, N10004);
nor NOR3 (N10008, N9985, N5925, N2084);
nand NAND3 (N10009, N10000, N3833, N8739);
nand NAND2 (N10010, N9969, N1723);
nor NOR3 (N10011, N10006, N336, N2248);
nand NAND2 (N10012, N10007, N9708);
xor XOR2 (N10013, N9979, N8405);
not NOT1 (N10014, N10010);
xor XOR2 (N10015, N10008, N8632);
buf BUF1 (N10016, N10003);
xor XOR2 (N10017, N10009, N5709);
xor XOR2 (N10018, N10016, N4980);
and AND4 (N10019, N10002, N744, N509, N3386);
buf BUF1 (N10020, N10018);
nor NOR2 (N10021, N10013, N2758);
nor NOR2 (N10022, N10014, N1221);
or OR3 (N10023, N10015, N967, N379);
buf BUF1 (N10024, N10020);
xor XOR2 (N10025, N10023, N4207);
nor NOR2 (N10026, N10019, N2952);
or OR4 (N10027, N10022, N1431, N1570, N3609);
or OR2 (N10028, N10026, N6868);
or OR2 (N10029, N10011, N5378);
nand NAND3 (N10030, N10024, N9000, N1124);
buf BUF1 (N10031, N10012);
xor XOR2 (N10032, N10025, N7183);
buf BUF1 (N10033, N10028);
nand NAND4 (N10034, N10029, N5975, N9983, N8752);
nor NOR3 (N10035, N10034, N4330, N5940);
and AND3 (N10036, N10030, N8669, N3530);
buf BUF1 (N10037, N10031);
buf BUF1 (N10038, N10037);
nand NAND2 (N10039, N10035, N4355);
buf BUF1 (N10040, N10036);
or OR3 (N10041, N10032, N364, N4422);
and AND3 (N10042, N10027, N9514, N7942);
or OR2 (N10043, N10005, N6514);
nand NAND3 (N10044, N10017, N5269, N7166);
nor NOR2 (N10045, N10041, N7010);
buf BUF1 (N10046, N10039);
buf BUF1 (N10047, N10042);
buf BUF1 (N10048, N10045);
buf BUF1 (N10049, N10038);
nor NOR4 (N10050, N10048, N5619, N9273, N219);
and AND2 (N10051, N10050, N7848);
or OR4 (N10052, N10033, N5158, N6581, N5395);
or OR2 (N10053, N10051, N8506);
xor XOR2 (N10054, N10052, N3033);
xor XOR2 (N10055, N10046, N2212);
and AND2 (N10056, N10021, N3010);
or OR4 (N10057, N10043, N9199, N7255, N6836);
not NOT1 (N10058, N10054);
buf BUF1 (N10059, N10049);
or OR4 (N10060, N10056, N2233, N872, N7356);
nor NOR2 (N10061, N9992, N8942);
nand NAND3 (N10062, N10053, N8066, N4841);
xor XOR2 (N10063, N10047, N4391);
nor NOR4 (N10064, N10063, N1376, N2763, N1611);
or OR3 (N10065, N10059, N1226, N3899);
or OR2 (N10066, N10057, N255);
nor NOR4 (N10067, N10060, N5588, N9216, N7551);
and AND2 (N10068, N10062, N9073);
xor XOR2 (N10069, N10055, N9898);
or OR4 (N10070, N10061, N5731, N668, N4752);
nand NAND2 (N10071, N10066, N3024);
not NOT1 (N10072, N10068);
nand NAND2 (N10073, N10069, N3337);
nand NAND3 (N10074, N10040, N7555, N1099);
nor NOR4 (N10075, N10072, N702, N583, N8132);
buf BUF1 (N10076, N10075);
nor NOR4 (N10077, N10074, N7535, N8619, N95);
nor NOR4 (N10078, N10044, N39, N6007, N8971);
nor NOR4 (N10079, N10064, N4106, N4973, N9359);
xor XOR2 (N10080, N10071, N3824);
not NOT1 (N10081, N10078);
nor NOR3 (N10082, N10077, N6971, N6754);
nand NAND2 (N10083, N10080, N2155);
xor XOR2 (N10084, N10079, N8516);
or OR2 (N10085, N10070, N5687);
nand NAND2 (N10086, N10084, N6905);
or OR3 (N10087, N10076, N3837, N8942);
nor NOR4 (N10088, N10086, N4179, N79, N6792);
buf BUF1 (N10089, N10087);
nor NOR4 (N10090, N10067, N4013, N1092, N1894);
buf BUF1 (N10091, N10073);
and AND4 (N10092, N10091, N364, N9400, N5209);
nor NOR4 (N10093, N10082, N6880, N194, N9002);
not NOT1 (N10094, N10085);
not NOT1 (N10095, N10083);
or OR4 (N10096, N10089, N7595, N2029, N5274);
nand NAND2 (N10097, N10095, N7459);
and AND2 (N10098, N10088, N9346);
and AND4 (N10099, N10092, N312, N7427, N3502);
not NOT1 (N10100, N10081);
and AND2 (N10101, N10098, N7104);
and AND3 (N10102, N10058, N8577, N3666);
nor NOR4 (N10103, N10065, N3403, N4351, N5446);
not NOT1 (N10104, N10102);
and AND4 (N10105, N10090, N3185, N826, N2791);
nand NAND4 (N10106, N10093, N9260, N3993, N3781);
not NOT1 (N10107, N10099);
nor NOR2 (N10108, N10103, N2217);
xor XOR2 (N10109, N10104, N2901);
and AND2 (N10110, N10100, N1598);
xor XOR2 (N10111, N10101, N8576);
buf BUF1 (N10112, N10109);
buf BUF1 (N10113, N10108);
or OR2 (N10114, N10105, N2428);
not NOT1 (N10115, N10113);
xor XOR2 (N10116, N10114, N8322);
buf BUF1 (N10117, N10107);
xor XOR2 (N10118, N10111, N2036);
xor XOR2 (N10119, N10115, N9378);
and AND3 (N10120, N10097, N481, N7878);
not NOT1 (N10121, N10106);
and AND3 (N10122, N10118, N6319, N3125);
xor XOR2 (N10123, N10120, N2447);
nand NAND3 (N10124, N10117, N8492, N7269);
nor NOR3 (N10125, N10119, N8901, N8905);
xor XOR2 (N10126, N10123, N6274);
or OR3 (N10127, N10126, N6989, N4088);
or OR3 (N10128, N10116, N5498, N3566);
buf BUF1 (N10129, N10096);
buf BUF1 (N10130, N10121);
nand NAND2 (N10131, N10128, N6219);
xor XOR2 (N10132, N10122, N4670);
nand NAND3 (N10133, N10094, N2332, N7090);
xor XOR2 (N10134, N10129, N4757);
nand NAND2 (N10135, N10131, N204);
nor NOR2 (N10136, N10125, N5289);
not NOT1 (N10137, N10135);
nand NAND4 (N10138, N10127, N4364, N5829, N7686);
nand NAND2 (N10139, N10134, N8601);
xor XOR2 (N10140, N10132, N3411);
and AND2 (N10141, N10136, N7846);
xor XOR2 (N10142, N10130, N96);
xor XOR2 (N10143, N10124, N7817);
xor XOR2 (N10144, N10137, N9001);
xor XOR2 (N10145, N10143, N7866);
nand NAND3 (N10146, N10138, N3638, N6087);
not NOT1 (N10147, N10144);
nor NOR2 (N10148, N10110, N3351);
or OR2 (N10149, N10145, N5320);
and AND2 (N10150, N10140, N9442);
not NOT1 (N10151, N10142);
buf BUF1 (N10152, N10150);
nand NAND3 (N10153, N10149, N4093, N2077);
nand NAND4 (N10154, N10139, N2813, N9340, N4983);
and AND2 (N10155, N10152, N1745);
nand NAND3 (N10156, N10146, N8254, N9856);
not NOT1 (N10157, N10147);
buf BUF1 (N10158, N10155);
or OR2 (N10159, N10157, N3603);
xor XOR2 (N10160, N10148, N3462);
xor XOR2 (N10161, N10133, N5398);
buf BUF1 (N10162, N10151);
buf BUF1 (N10163, N10112);
or OR2 (N10164, N10141, N5058);
buf BUF1 (N10165, N10160);
or OR2 (N10166, N10162, N9584);
xor XOR2 (N10167, N10156, N6875);
and AND2 (N10168, N10167, N4742);
xor XOR2 (N10169, N10153, N6097);
nand NAND4 (N10170, N10159, N4022, N4706, N2483);
and AND4 (N10171, N10161, N7855, N2187, N5009);
or OR4 (N10172, N10170, N9380, N1989, N3017);
not NOT1 (N10173, N10158);
xor XOR2 (N10174, N10169, N4883);
and AND4 (N10175, N10163, N3057, N5620, N5564);
and AND4 (N10176, N10171, N9882, N1183, N1811);
or OR2 (N10177, N10172, N5552);
nand NAND3 (N10178, N10154, N862, N9296);
and AND4 (N10179, N10168, N9479, N5809, N3720);
or OR3 (N10180, N10179, N4999, N9875);
buf BUF1 (N10181, N10178);
not NOT1 (N10182, N10176);
and AND3 (N10183, N10182, N2439, N1047);
nand NAND2 (N10184, N10164, N9370);
and AND2 (N10185, N10175, N5914);
and AND4 (N10186, N10180, N8206, N944, N6716);
or OR3 (N10187, N10186, N2219, N1652);
not NOT1 (N10188, N10166);
nand NAND3 (N10189, N10187, N7295, N1468);
xor XOR2 (N10190, N10185, N121);
nand NAND2 (N10191, N10177, N5583);
xor XOR2 (N10192, N10183, N9324);
or OR2 (N10193, N10191, N475);
or OR3 (N10194, N10193, N6347, N5840);
buf BUF1 (N10195, N10184);
xor XOR2 (N10196, N10173, N943);
nor NOR4 (N10197, N10189, N4395, N4065, N1875);
nand NAND3 (N10198, N10190, N8942, N9383);
nor NOR4 (N10199, N10181, N3365, N2101, N8194);
nor NOR3 (N10200, N10194, N977, N9158);
nand NAND3 (N10201, N10197, N5651, N369);
nand NAND2 (N10202, N10199, N3682);
and AND3 (N10203, N10200, N6427, N5780);
not NOT1 (N10204, N10192);
xor XOR2 (N10205, N10204, N9494);
and AND4 (N10206, N10196, N3336, N6096, N6381);
or OR4 (N10207, N10203, N715, N5315, N4268);
or OR2 (N10208, N10207, N5846);
or OR3 (N10209, N10205, N10131, N6845);
not NOT1 (N10210, N10174);
not NOT1 (N10211, N10202);
buf BUF1 (N10212, N10195);
buf BUF1 (N10213, N10212);
xor XOR2 (N10214, N10201, N3844);
and AND4 (N10215, N10188, N9470, N6800, N6540);
nand NAND2 (N10216, N10198, N9347);
buf BUF1 (N10217, N10165);
or OR2 (N10218, N10210, N7602);
or OR3 (N10219, N10214, N3114, N8828);
nand NAND3 (N10220, N10217, N7266, N1237);
nand NAND3 (N10221, N10219, N5993, N2383);
not NOT1 (N10222, N10220);
or OR2 (N10223, N10218, N4772);
buf BUF1 (N10224, N10222);
nor NOR4 (N10225, N10209, N4776, N7492, N9576);
buf BUF1 (N10226, N10224);
xor XOR2 (N10227, N10211, N2272);
xor XOR2 (N10228, N10221, N2795);
not NOT1 (N10229, N10225);
xor XOR2 (N10230, N10216, N2219);
xor XOR2 (N10231, N10208, N4098);
or OR3 (N10232, N10206, N2474, N8496);
buf BUF1 (N10233, N10230);
nand NAND4 (N10234, N10223, N2596, N2174, N7155);
nor NOR4 (N10235, N10213, N4173, N6424, N4586);
not NOT1 (N10236, N10235);
or OR4 (N10237, N10236, N3553, N4288, N2096);
nand NAND4 (N10238, N10227, N4186, N5357, N8992);
not NOT1 (N10239, N10237);
nor NOR2 (N10240, N10231, N6082);
nor NOR4 (N10241, N10228, N9688, N5126, N4038);
not NOT1 (N10242, N10239);
xor XOR2 (N10243, N10226, N7983);
not NOT1 (N10244, N10242);
nand NAND4 (N10245, N10215, N3060, N9336, N1262);
not NOT1 (N10246, N10244);
or OR2 (N10247, N10240, N2866);
not NOT1 (N10248, N10246);
or OR2 (N10249, N10243, N3488);
or OR2 (N10250, N10234, N5007);
or OR3 (N10251, N10238, N2814, N9751);
not NOT1 (N10252, N10233);
or OR2 (N10253, N10251, N5105);
nand NAND4 (N10254, N10229, N1960, N7525, N6046);
or OR3 (N10255, N10250, N5445, N9205);
and AND3 (N10256, N10252, N1470, N8741);
and AND4 (N10257, N10249, N248, N1933, N7536);
not NOT1 (N10258, N10247);
buf BUF1 (N10259, N10232);
nor NOR3 (N10260, N10253, N6716, N3544);
not NOT1 (N10261, N10260);
nand NAND2 (N10262, N10248, N2761);
buf BUF1 (N10263, N10256);
not NOT1 (N10264, N10259);
nor NOR4 (N10265, N10255, N8126, N2055, N1886);
nor NOR3 (N10266, N10265, N8039, N8534);
nor NOR3 (N10267, N10266, N1463, N3750);
xor XOR2 (N10268, N10257, N9141);
nor NOR3 (N10269, N10258, N97, N1085);
nand NAND3 (N10270, N10261, N7471, N7343);
not NOT1 (N10271, N10262);
buf BUF1 (N10272, N10254);
nand NAND3 (N10273, N10245, N3109, N10117);
and AND4 (N10274, N10241, N3116, N5999, N5161);
nand NAND4 (N10275, N10264, N2612, N3348, N3718);
not NOT1 (N10276, N10271);
buf BUF1 (N10277, N10263);
buf BUF1 (N10278, N10272);
not NOT1 (N10279, N10269);
xor XOR2 (N10280, N10267, N6948);
buf BUF1 (N10281, N10273);
xor XOR2 (N10282, N10279, N1179);
or OR3 (N10283, N10268, N3668, N766);
xor XOR2 (N10284, N10275, N4009);
or OR2 (N10285, N10283, N4755);
nor NOR2 (N10286, N10270, N7537);
not NOT1 (N10287, N10274);
nand NAND2 (N10288, N10276, N7227);
buf BUF1 (N10289, N10282);
xor XOR2 (N10290, N10280, N1114);
or OR2 (N10291, N10290, N4882);
nor NOR2 (N10292, N10284, N5968);
xor XOR2 (N10293, N10285, N4738);
and AND4 (N10294, N10281, N9158, N1076, N9615);
xor XOR2 (N10295, N10291, N8232);
nor NOR2 (N10296, N10277, N4077);
not NOT1 (N10297, N10287);
not NOT1 (N10298, N10286);
or OR3 (N10299, N10297, N342, N5074);
buf BUF1 (N10300, N10288);
buf BUF1 (N10301, N10299);
buf BUF1 (N10302, N10300);
not NOT1 (N10303, N10302);
nor NOR2 (N10304, N10289, N8640);
buf BUF1 (N10305, N10278);
not NOT1 (N10306, N10303);
nor NOR2 (N10307, N10292, N4365);
xor XOR2 (N10308, N10307, N7517);
xor XOR2 (N10309, N10295, N2369);
xor XOR2 (N10310, N10296, N890);
buf BUF1 (N10311, N10304);
xor XOR2 (N10312, N10308, N2684);
nor NOR2 (N10313, N10310, N1359);
or OR2 (N10314, N10301, N953);
or OR2 (N10315, N10305, N3384);
or OR4 (N10316, N10309, N1854, N3315, N9446);
xor XOR2 (N10317, N10293, N6735);
or OR4 (N10318, N10298, N4662, N8150, N5530);
nand NAND3 (N10319, N10317, N1976, N1667);
buf BUF1 (N10320, N10312);
and AND2 (N10321, N10316, N4491);
nor NOR2 (N10322, N10321, N4596);
or OR4 (N10323, N10320, N590, N9621, N9440);
buf BUF1 (N10324, N10319);
buf BUF1 (N10325, N10313);
and AND4 (N10326, N10323, N207, N7024, N3697);
and AND4 (N10327, N10314, N5784, N8521, N9063);
and AND3 (N10328, N10311, N508, N2803);
buf BUF1 (N10329, N10325);
nor NOR4 (N10330, N10318, N5650, N933, N5523);
nor NOR2 (N10331, N10324, N9103);
and AND4 (N10332, N10315, N1965, N8175, N5448);
or OR3 (N10333, N10294, N2651, N1817);
nor NOR2 (N10334, N10332, N3898);
xor XOR2 (N10335, N10306, N9625);
xor XOR2 (N10336, N10326, N6419);
nor NOR3 (N10337, N10334, N1618, N8804);
buf BUF1 (N10338, N10335);
buf BUF1 (N10339, N10331);
buf BUF1 (N10340, N10329);
xor XOR2 (N10341, N10330, N2123);
nand NAND2 (N10342, N10337, N2672);
nor NOR3 (N10343, N10340, N1368, N1648);
buf BUF1 (N10344, N10322);
not NOT1 (N10345, N10343);
nor NOR2 (N10346, N10341, N2266);
and AND4 (N10347, N10333, N8741, N4414, N6424);
nand NAND2 (N10348, N10347, N3525);
and AND3 (N10349, N10336, N1284, N8569);
nor NOR2 (N10350, N10345, N7220);
nor NOR2 (N10351, N10344, N5477);
and AND2 (N10352, N10327, N10003);
or OR3 (N10353, N10342, N7617, N10230);
nand NAND2 (N10354, N10348, N6593);
nor NOR2 (N10355, N10352, N7603);
nand NAND4 (N10356, N10339, N6925, N7557, N3243);
nor NOR2 (N10357, N10346, N4228);
buf BUF1 (N10358, N10328);
or OR4 (N10359, N10350, N8606, N3074, N1918);
nor NOR2 (N10360, N10359, N2203);
nor NOR4 (N10361, N10355, N3622, N8666, N8227);
xor XOR2 (N10362, N10357, N9539);
and AND4 (N10363, N10338, N2321, N6763, N7194);
nor NOR2 (N10364, N10353, N851);
buf BUF1 (N10365, N10351);
nor NOR4 (N10366, N10356, N5759, N327, N7364);
and AND2 (N10367, N10365, N6732);
buf BUF1 (N10368, N10360);
xor XOR2 (N10369, N10364, N3109);
buf BUF1 (N10370, N10358);
buf BUF1 (N10371, N10368);
and AND2 (N10372, N10367, N4899);
xor XOR2 (N10373, N10349, N4219);
buf BUF1 (N10374, N10369);
buf BUF1 (N10375, N10373);
or OR4 (N10376, N10362, N3566, N10214, N2360);
and AND2 (N10377, N10354, N10288);
and AND3 (N10378, N10374, N9180, N1948);
buf BUF1 (N10379, N10361);
nor NOR2 (N10380, N10375, N2679);
or OR4 (N10381, N10366, N4953, N510, N2979);
or OR4 (N10382, N10379, N4356, N2296, N5732);
xor XOR2 (N10383, N10363, N3020);
nand NAND2 (N10384, N10376, N3295);
and AND3 (N10385, N10384, N7609, N2776);
and AND2 (N10386, N10370, N261);
nor NOR2 (N10387, N10385, N3600);
buf BUF1 (N10388, N10377);
nand NAND4 (N10389, N10387, N2088, N539, N1588);
nand NAND3 (N10390, N10378, N8456, N8519);
or OR3 (N10391, N10371, N9379, N5536);
buf BUF1 (N10392, N10388);
xor XOR2 (N10393, N10389, N8494);
nor NOR2 (N10394, N10391, N9412);
nand NAND4 (N10395, N10381, N2556, N3811, N4550);
and AND2 (N10396, N10393, N10208);
nand NAND4 (N10397, N10380, N6464, N191, N3051);
not NOT1 (N10398, N10395);
buf BUF1 (N10399, N10392);
not NOT1 (N10400, N10382);
xor XOR2 (N10401, N10399, N5978);
not NOT1 (N10402, N10390);
nand NAND2 (N10403, N10383, N3316);
and AND2 (N10404, N10398, N6699);
and AND4 (N10405, N10402, N3317, N10092, N356);
nand NAND2 (N10406, N10396, N6164);
not NOT1 (N10407, N10404);
xor XOR2 (N10408, N10401, N7705);
xor XOR2 (N10409, N10407, N2879);
nor NOR2 (N10410, N10400, N2952);
nor NOR2 (N10411, N10372, N2281);
xor XOR2 (N10412, N10405, N9350);
not NOT1 (N10413, N10409);
and AND3 (N10414, N10411, N1688, N6594);
or OR2 (N10415, N10408, N5491);
and AND3 (N10416, N10406, N1172, N5858);
nor NOR3 (N10417, N10386, N6525, N4140);
buf BUF1 (N10418, N10415);
nor NOR4 (N10419, N10418, N6360, N9712, N8267);
nor NOR3 (N10420, N10397, N6717, N1499);
not NOT1 (N10421, N10394);
nor NOR4 (N10422, N10420, N4055, N8543, N1897);
not NOT1 (N10423, N10416);
and AND3 (N10424, N10414, N9910, N10086);
xor XOR2 (N10425, N10403, N2442);
and AND2 (N10426, N10425, N1957);
buf BUF1 (N10427, N10417);
nand NAND3 (N10428, N10421, N3852, N6411);
nor NOR4 (N10429, N10426, N4967, N7498, N2820);
or OR4 (N10430, N10413, N7786, N5792, N4410);
or OR4 (N10431, N10422, N10206, N9534, N7198);
not NOT1 (N10432, N10429);
buf BUF1 (N10433, N10424);
nand NAND4 (N10434, N10430, N1204, N9881, N2063);
not NOT1 (N10435, N10433);
not NOT1 (N10436, N10431);
buf BUF1 (N10437, N10432);
nor NOR3 (N10438, N10423, N1607, N8023);
xor XOR2 (N10439, N10434, N5984);
and AND3 (N10440, N10428, N8285, N7266);
and AND4 (N10441, N10439, N9812, N9324, N2293);
buf BUF1 (N10442, N10435);
xor XOR2 (N10443, N10441, N8813);
not NOT1 (N10444, N10442);
xor XOR2 (N10445, N10444, N4853);
not NOT1 (N10446, N10440);
not NOT1 (N10447, N10436);
or OR2 (N10448, N10438, N8530);
buf BUF1 (N10449, N10443);
nor NOR3 (N10450, N10419, N1802, N6095);
not NOT1 (N10451, N10448);
xor XOR2 (N10452, N10445, N3269);
xor XOR2 (N10453, N10451, N1476);
or OR4 (N10454, N10427, N7753, N3801, N8057);
and AND2 (N10455, N10412, N5119);
nand NAND2 (N10456, N10452, N7673);
and AND4 (N10457, N10447, N2379, N4574, N9929);
buf BUF1 (N10458, N10410);
nor NOR3 (N10459, N10446, N6681, N4381);
nand NAND3 (N10460, N10437, N3112, N9228);
nand NAND2 (N10461, N10454, N4286);
buf BUF1 (N10462, N10457);
buf BUF1 (N10463, N10449);
nand NAND4 (N10464, N10461, N2083, N3156, N7935);
xor XOR2 (N10465, N10453, N7698);
not NOT1 (N10466, N10463);
nand NAND4 (N10467, N10466, N8235, N6632, N10196);
or OR3 (N10468, N10450, N6647, N10415);
not NOT1 (N10469, N10458);
nor NOR3 (N10470, N10459, N7501, N3990);
and AND2 (N10471, N10456, N6044);
xor XOR2 (N10472, N10468, N3296);
not NOT1 (N10473, N10462);
xor XOR2 (N10474, N10465, N3261);
buf BUF1 (N10475, N10455);
or OR2 (N10476, N10475, N201);
xor XOR2 (N10477, N10472, N5049);
nor NOR2 (N10478, N10476, N4068);
nor NOR4 (N10479, N10474, N9050, N8580, N5404);
not NOT1 (N10480, N10464);
not NOT1 (N10481, N10479);
or OR4 (N10482, N10477, N1535, N5207, N10268);
xor XOR2 (N10483, N10481, N6970);
xor XOR2 (N10484, N10480, N4496);
nand NAND2 (N10485, N10483, N5601);
buf BUF1 (N10486, N10485);
nand NAND3 (N10487, N10478, N9564, N6131);
nor NOR4 (N10488, N10471, N1623, N9425, N4463);
buf BUF1 (N10489, N10467);
and AND4 (N10490, N10473, N996, N5542, N8043);
and AND2 (N10491, N10482, N5378);
or OR4 (N10492, N10486, N3378, N3379, N55);
not NOT1 (N10493, N10489);
nand NAND2 (N10494, N10484, N5362);
nor NOR4 (N10495, N10494, N6862, N7917, N6739);
and AND3 (N10496, N10491, N9392, N1261);
buf BUF1 (N10497, N10488);
and AND3 (N10498, N10487, N2428, N1695);
and AND2 (N10499, N10495, N8604);
and AND4 (N10500, N10469, N2836, N1026, N991);
xor XOR2 (N10501, N10499, N3903);
not NOT1 (N10502, N10498);
and AND3 (N10503, N10492, N6065, N1655);
nor NOR2 (N10504, N10493, N3802);
not NOT1 (N10505, N10460);
xor XOR2 (N10506, N10505, N6720);
not NOT1 (N10507, N10470);
and AND2 (N10508, N10500, N5543);
buf BUF1 (N10509, N10497);
xor XOR2 (N10510, N10501, N6377);
nor NOR2 (N10511, N10496, N9611);
nor NOR4 (N10512, N10503, N2008, N9553, N2042);
xor XOR2 (N10513, N10508, N5763);
nand NAND3 (N10514, N10506, N7967, N7322);
nand NAND4 (N10515, N10509, N3945, N9084, N6101);
nor NOR4 (N10516, N10502, N8006, N808, N4094);
xor XOR2 (N10517, N10515, N5934);
xor XOR2 (N10518, N10513, N3941);
nor NOR4 (N10519, N10490, N2906, N4669, N4049);
not NOT1 (N10520, N10504);
nor NOR3 (N10521, N10519, N8927, N607);
and AND2 (N10522, N10514, N1377);
nand NAND3 (N10523, N10517, N2313, N4437);
buf BUF1 (N10524, N10507);
nand NAND2 (N10525, N10523, N1370);
nor NOR3 (N10526, N10524, N4617, N6585);
and AND2 (N10527, N10518, N3364);
xor XOR2 (N10528, N10520, N10169);
buf BUF1 (N10529, N10516);
not NOT1 (N10530, N10525);
xor XOR2 (N10531, N10527, N3228);
and AND2 (N10532, N10521, N2886);
xor XOR2 (N10533, N10531, N6738);
xor XOR2 (N10534, N10532, N4552);
buf BUF1 (N10535, N10530);
and AND3 (N10536, N10511, N5206, N7892);
nor NOR2 (N10537, N10526, N2492);
and AND3 (N10538, N10529, N7795, N2531);
and AND3 (N10539, N10538, N10447, N5277);
buf BUF1 (N10540, N10534);
nor NOR3 (N10541, N10512, N4232, N3529);
nor NOR4 (N10542, N10522, N7353, N553, N10006);
buf BUF1 (N10543, N10533);
nor NOR3 (N10544, N10535, N10064, N4264);
and AND2 (N10545, N10539, N1924);
nor NOR3 (N10546, N10543, N4529, N6884);
and AND3 (N10547, N10546, N1356, N6057);
or OR4 (N10548, N10545, N560, N4668, N7965);
not NOT1 (N10549, N10547);
xor XOR2 (N10550, N10540, N481);
or OR2 (N10551, N10544, N5389);
nand NAND2 (N10552, N10550, N980);
or OR2 (N10553, N10537, N7753);
buf BUF1 (N10554, N10552);
and AND2 (N10555, N10542, N21);
and AND3 (N10556, N10549, N4416, N6497);
and AND3 (N10557, N10556, N4854, N839);
nand NAND2 (N10558, N10528, N9295);
nand NAND2 (N10559, N10541, N2948);
and AND3 (N10560, N10536, N5317, N297);
and AND2 (N10561, N10551, N2460);
buf BUF1 (N10562, N10555);
nand NAND4 (N10563, N10558, N6002, N7726, N3582);
buf BUF1 (N10564, N10553);
nor NOR3 (N10565, N10548, N3325, N3894);
not NOT1 (N10566, N10561);
nor NOR3 (N10567, N10564, N3270, N7791);
not NOT1 (N10568, N10554);
and AND4 (N10569, N10510, N9219, N2457, N5517);
xor XOR2 (N10570, N10566, N4618);
buf BUF1 (N10571, N10560);
nor NOR3 (N10572, N10567, N3891, N2181);
nor NOR4 (N10573, N10562, N3706, N3056, N4849);
nand NAND3 (N10574, N10571, N7458, N6221);
or OR3 (N10575, N10574, N3129, N9012);
not NOT1 (N10576, N10572);
and AND4 (N10577, N10569, N6205, N5412, N2808);
xor XOR2 (N10578, N10570, N5252);
nand NAND3 (N10579, N10573, N2140, N519);
not NOT1 (N10580, N10575);
nand NAND4 (N10581, N10576, N6999, N8358, N7952);
xor XOR2 (N10582, N10581, N4985);
xor XOR2 (N10583, N10578, N3349);
not NOT1 (N10584, N10579);
and AND4 (N10585, N10563, N308, N7370, N3132);
nor NOR4 (N10586, N10584, N8293, N1239, N8998);
not NOT1 (N10587, N10580);
not NOT1 (N10588, N10565);
xor XOR2 (N10589, N10559, N4012);
or OR2 (N10590, N10568, N2624);
xor XOR2 (N10591, N10585, N4862);
buf BUF1 (N10592, N10557);
buf BUF1 (N10593, N10591);
nor NOR4 (N10594, N10587, N5261, N3141, N1080);
not NOT1 (N10595, N10593);
nor NOR2 (N10596, N10588, N1345);
xor XOR2 (N10597, N10589, N6642);
and AND4 (N10598, N10582, N9684, N5280, N6523);
and AND3 (N10599, N10577, N7138, N8434);
and AND3 (N10600, N10595, N10407, N1998);
or OR3 (N10601, N10598, N1643, N9838);
or OR4 (N10602, N10597, N204, N2751, N6562);
xor XOR2 (N10603, N10596, N2431);
and AND3 (N10604, N10583, N5982, N8823);
nor NOR4 (N10605, N10603, N9205, N8975, N1913);
or OR4 (N10606, N10605, N2413, N1480, N829);
nand NAND3 (N10607, N10592, N6331, N2040);
xor XOR2 (N10608, N10602, N4347);
buf BUF1 (N10609, N10594);
nor NOR2 (N10610, N10604, N6829);
or OR2 (N10611, N10608, N3758);
buf BUF1 (N10612, N10600);
buf BUF1 (N10613, N10607);
nand NAND3 (N10614, N10610, N2318, N3006);
nand NAND3 (N10615, N10599, N8411, N8865);
nand NAND4 (N10616, N10611, N569, N5807, N933);
not NOT1 (N10617, N10586);
not NOT1 (N10618, N10614);
nor NOR3 (N10619, N10601, N9566, N2837);
or OR2 (N10620, N10619, N5897);
nand NAND2 (N10621, N10620, N8391);
and AND3 (N10622, N10615, N7165, N2551);
xor XOR2 (N10623, N10612, N8323);
xor XOR2 (N10624, N10609, N10106);
not NOT1 (N10625, N10622);
nor NOR2 (N10626, N10617, N5155);
buf BUF1 (N10627, N10616);
buf BUF1 (N10628, N10618);
and AND2 (N10629, N10606, N9653);
nand NAND3 (N10630, N10626, N7637, N573);
or OR4 (N10631, N10621, N9403, N1727, N3161);
and AND2 (N10632, N10631, N900);
nor NOR3 (N10633, N10623, N1418, N2616);
not NOT1 (N10634, N10632);
xor XOR2 (N10635, N10625, N6890);
xor XOR2 (N10636, N10633, N27);
not NOT1 (N10637, N10613);
xor XOR2 (N10638, N10635, N7620);
and AND4 (N10639, N10637, N5829, N5831, N5602);
xor XOR2 (N10640, N10639, N6664);
buf BUF1 (N10641, N10630);
xor XOR2 (N10642, N10641, N9657);
nand NAND3 (N10643, N10638, N2747, N8481);
xor XOR2 (N10644, N10643, N778);
and AND3 (N10645, N10590, N6475, N10412);
nor NOR3 (N10646, N10634, N5066, N551);
buf BUF1 (N10647, N10645);
not NOT1 (N10648, N10627);
not NOT1 (N10649, N10628);
xor XOR2 (N10650, N10629, N9636);
xor XOR2 (N10651, N10642, N6337);
nand NAND3 (N10652, N10649, N6554, N4892);
nand NAND3 (N10653, N10648, N6153, N6982);
or OR3 (N10654, N10624, N81, N1971);
not NOT1 (N10655, N10651);
nand NAND3 (N10656, N10654, N5235, N9643);
xor XOR2 (N10657, N10646, N9649);
nand NAND2 (N10658, N10655, N2861);
xor XOR2 (N10659, N10650, N638);
nor NOR2 (N10660, N10657, N7491);
not NOT1 (N10661, N10644);
or OR2 (N10662, N10658, N8101);
nor NOR3 (N10663, N10647, N7398, N9456);
and AND4 (N10664, N10662, N5019, N1532, N8172);
xor XOR2 (N10665, N10661, N6528);
nand NAND3 (N10666, N10640, N3466, N3304);
nand NAND4 (N10667, N10664, N7231, N6289, N6856);
xor XOR2 (N10668, N10636, N3091);
nand NAND3 (N10669, N10652, N8047, N4201);
nor NOR2 (N10670, N10667, N5663);
xor XOR2 (N10671, N10659, N2168);
buf BUF1 (N10672, N10656);
or OR4 (N10673, N10671, N7750, N1784, N5117);
xor XOR2 (N10674, N10668, N10345);
buf BUF1 (N10675, N10660);
and AND3 (N10676, N10672, N4256, N4214);
or OR2 (N10677, N10665, N74);
buf BUF1 (N10678, N10670);
xor XOR2 (N10679, N10663, N5269);
nand NAND4 (N10680, N10666, N10318, N5075, N8954);
buf BUF1 (N10681, N10677);
xor XOR2 (N10682, N10675, N2915);
or OR4 (N10683, N10678, N8996, N8360, N8629);
nand NAND4 (N10684, N10679, N1448, N1849, N3549);
or OR4 (N10685, N10681, N430, N8477, N8958);
nand NAND4 (N10686, N10684, N8753, N10627, N2383);
or OR3 (N10687, N10685, N297, N941);
nor NOR3 (N10688, N10674, N1625, N3489);
or OR4 (N10689, N10680, N9554, N5818, N6261);
or OR3 (N10690, N10676, N3704, N3205);
nor NOR3 (N10691, N10669, N314, N2265);
xor XOR2 (N10692, N10653, N3983);
buf BUF1 (N10693, N10691);
xor XOR2 (N10694, N10689, N6965);
buf BUF1 (N10695, N10693);
buf BUF1 (N10696, N10686);
nor NOR3 (N10697, N10683, N4803, N2811);
nor NOR2 (N10698, N10694, N1946);
or OR2 (N10699, N10696, N8094);
and AND4 (N10700, N10673, N737, N5700, N8214);
xor XOR2 (N10701, N10687, N3278);
buf BUF1 (N10702, N10695);
not NOT1 (N10703, N10697);
xor XOR2 (N10704, N10700, N1391);
nor NOR2 (N10705, N10692, N8424);
or OR3 (N10706, N10705, N4324, N979);
not NOT1 (N10707, N10690);
nand NAND4 (N10708, N10703, N272, N7441, N9686);
xor XOR2 (N10709, N10701, N182);
and AND4 (N10710, N10688, N5692, N9239, N3785);
not NOT1 (N10711, N10709);
not NOT1 (N10712, N10704);
buf BUF1 (N10713, N10706);
nand NAND2 (N10714, N10702, N6386);
or OR2 (N10715, N10711, N4680);
nand NAND2 (N10716, N10698, N3551);
buf BUF1 (N10717, N10707);
buf BUF1 (N10718, N10682);
nand NAND3 (N10719, N10718, N2366, N2458);
xor XOR2 (N10720, N10717, N3833);
xor XOR2 (N10721, N10713, N5949);
xor XOR2 (N10722, N10699, N10569);
buf BUF1 (N10723, N10722);
xor XOR2 (N10724, N10719, N5117);
nand NAND3 (N10725, N10720, N9160, N8196);
nor NOR2 (N10726, N10714, N7707);
buf BUF1 (N10727, N10724);
nand NAND2 (N10728, N10723, N6637);
buf BUF1 (N10729, N10715);
xor XOR2 (N10730, N10725, N6965);
xor XOR2 (N10731, N10727, N9816);
nand NAND2 (N10732, N10728, N1392);
xor XOR2 (N10733, N10716, N9107);
not NOT1 (N10734, N10721);
or OR2 (N10735, N10731, N5424);
not NOT1 (N10736, N10708);
xor XOR2 (N10737, N10710, N9881);
nand NAND2 (N10738, N10726, N9236);
not NOT1 (N10739, N10734);
not NOT1 (N10740, N10735);
nand NAND4 (N10741, N10740, N2553, N9252, N3878);
xor XOR2 (N10742, N10730, N8349);
nor NOR4 (N10743, N10737, N8658, N885, N481);
not NOT1 (N10744, N10712);
not NOT1 (N10745, N10744);
buf BUF1 (N10746, N10743);
nand NAND2 (N10747, N10733, N2312);
buf BUF1 (N10748, N10738);
xor XOR2 (N10749, N10739, N85);
nand NAND3 (N10750, N10748, N7849, N7602);
buf BUF1 (N10751, N10750);
nor NOR2 (N10752, N10751, N6277);
or OR2 (N10753, N10747, N5331);
or OR2 (N10754, N10741, N6500);
and AND3 (N10755, N10729, N7923, N5891);
nor NOR3 (N10756, N10753, N8107, N5782);
xor XOR2 (N10757, N10755, N6346);
xor XOR2 (N10758, N10757, N8994);
not NOT1 (N10759, N10756);
not NOT1 (N10760, N10758);
nor NOR2 (N10761, N10749, N3410);
and AND4 (N10762, N10754, N931, N7234, N3667);
not NOT1 (N10763, N10742);
nor NOR4 (N10764, N10746, N10537, N6562, N4766);
nor NOR2 (N10765, N10764, N7325);
and AND4 (N10766, N10745, N7582, N316, N3807);
nand NAND2 (N10767, N10732, N2317);
xor XOR2 (N10768, N10763, N1185);
xor XOR2 (N10769, N10768, N8360);
or OR4 (N10770, N10762, N7586, N10740, N7716);
not NOT1 (N10771, N10766);
or OR2 (N10772, N10770, N8893);
or OR4 (N10773, N10767, N8978, N8483, N7852);
xor XOR2 (N10774, N10765, N691);
nor NOR3 (N10775, N10772, N2593, N33);
nor NOR2 (N10776, N10761, N3636);
buf BUF1 (N10777, N10759);
not NOT1 (N10778, N10760);
xor XOR2 (N10779, N10736, N9331);
not NOT1 (N10780, N10771);
or OR3 (N10781, N10780, N5627, N1646);
xor XOR2 (N10782, N10781, N5372);
nor NOR3 (N10783, N10769, N7069, N5085);
nor NOR4 (N10784, N10778, N2601, N6475, N8216);
xor XOR2 (N10785, N10773, N1883);
xor XOR2 (N10786, N10776, N681);
and AND4 (N10787, N10785, N646, N9702, N7230);
and AND4 (N10788, N10784, N6090, N6147, N7204);
and AND4 (N10789, N10777, N4576, N6353, N5352);
not NOT1 (N10790, N10783);
nor NOR2 (N10791, N10790, N8327);
nor NOR4 (N10792, N10752, N3152, N4923, N6395);
not NOT1 (N10793, N10792);
and AND2 (N10794, N10793, N3866);
nand NAND2 (N10795, N10789, N10506);
not NOT1 (N10796, N10791);
xor XOR2 (N10797, N10779, N4058);
and AND2 (N10798, N10787, N1495);
nor NOR2 (N10799, N10794, N3734);
and AND3 (N10800, N10782, N4484, N8051);
and AND3 (N10801, N10796, N6372, N3723);
nand NAND4 (N10802, N10800, N7332, N6528, N2420);
not NOT1 (N10803, N10774);
nor NOR2 (N10804, N10775, N1574);
not NOT1 (N10805, N10801);
xor XOR2 (N10806, N10804, N4348);
and AND4 (N10807, N10788, N2429, N8582, N7739);
nor NOR2 (N10808, N10795, N7145);
not NOT1 (N10809, N10799);
not NOT1 (N10810, N10809);
not NOT1 (N10811, N10806);
not NOT1 (N10812, N10802);
buf BUF1 (N10813, N10810);
nor NOR3 (N10814, N10797, N6716, N1661);
and AND4 (N10815, N10812, N7110, N3679, N813);
nand NAND3 (N10816, N10786, N3577, N2113);
or OR4 (N10817, N10805, N10007, N10293, N1535);
or OR2 (N10818, N10798, N1645);
xor XOR2 (N10819, N10814, N4827);
nor NOR4 (N10820, N10816, N8870, N10432, N2827);
or OR2 (N10821, N10813, N3723);
not NOT1 (N10822, N10815);
nand NAND4 (N10823, N10820, N4576, N1857, N8351);
nor NOR4 (N10824, N10819, N586, N1799, N3786);
and AND3 (N10825, N10803, N2141, N6462);
buf BUF1 (N10826, N10808);
nor NOR3 (N10827, N10818, N8208, N8447);
not NOT1 (N10828, N10821);
not NOT1 (N10829, N10817);
or OR3 (N10830, N10826, N7220, N10237);
buf BUF1 (N10831, N10828);
and AND2 (N10832, N10823, N6249);
buf BUF1 (N10833, N10824);
and AND3 (N10834, N10832, N9544, N3462);
or OR4 (N10835, N10831, N9018, N773, N4428);
xor XOR2 (N10836, N10833, N8827);
nor NOR2 (N10837, N10807, N3862);
nand NAND3 (N10838, N10811, N1222, N9712);
and AND2 (N10839, N10838, N3320);
xor XOR2 (N10840, N10829, N4813);
nand NAND4 (N10841, N10822, N5775, N9765, N3108);
and AND3 (N10842, N10825, N10757, N3042);
or OR3 (N10843, N10836, N7845, N7541);
not NOT1 (N10844, N10835);
nor NOR3 (N10845, N10834, N2947, N6357);
nor NOR2 (N10846, N10830, N1129);
and AND4 (N10847, N10837, N7303, N5052, N3283);
xor XOR2 (N10848, N10827, N7407);
not NOT1 (N10849, N10844);
nor NOR2 (N10850, N10845, N10621);
or OR3 (N10851, N10846, N6857, N4817);
not NOT1 (N10852, N10843);
or OR3 (N10853, N10848, N8275, N3802);
nand NAND3 (N10854, N10847, N7842, N7544);
buf BUF1 (N10855, N10851);
nor NOR2 (N10856, N10841, N513);
nor NOR3 (N10857, N10854, N451, N5948);
buf BUF1 (N10858, N10853);
buf BUF1 (N10859, N10842);
buf BUF1 (N10860, N10858);
buf BUF1 (N10861, N10849);
nand NAND4 (N10862, N10855, N6853, N7094, N2309);
xor XOR2 (N10863, N10850, N5967);
not NOT1 (N10864, N10852);
or OR3 (N10865, N10861, N8112, N6686);
or OR4 (N10866, N10865, N4736, N10500, N7905);
xor XOR2 (N10867, N10840, N2928);
nand NAND3 (N10868, N10867, N7708, N10814);
nor NOR3 (N10869, N10859, N6758, N5253);
and AND3 (N10870, N10864, N597, N1929);
nor NOR4 (N10871, N10870, N10088, N9927, N5507);
buf BUF1 (N10872, N10869);
not NOT1 (N10873, N10862);
not NOT1 (N10874, N10839);
nand NAND3 (N10875, N10866, N921, N9420);
and AND3 (N10876, N10856, N1909, N7800);
nor NOR3 (N10877, N10872, N4446, N8983);
xor XOR2 (N10878, N10874, N1251);
and AND4 (N10879, N10875, N8562, N9871, N6460);
nand NAND3 (N10880, N10877, N3170, N7738);
not NOT1 (N10881, N10871);
buf BUF1 (N10882, N10879);
not NOT1 (N10883, N10868);
and AND3 (N10884, N10857, N3898, N2134);
or OR2 (N10885, N10882, N10365);
and AND4 (N10886, N10881, N8660, N654, N7965);
nor NOR3 (N10887, N10863, N3547, N5221);
nand NAND4 (N10888, N10878, N10706, N9181, N7093);
not NOT1 (N10889, N10860);
nor NOR3 (N10890, N10880, N257, N9171);
buf BUF1 (N10891, N10889);
and AND4 (N10892, N10887, N3047, N2654, N6717);
xor XOR2 (N10893, N10873, N7593);
not NOT1 (N10894, N10884);
and AND4 (N10895, N10892, N995, N596, N528);
xor XOR2 (N10896, N10876, N4651);
nor NOR4 (N10897, N10891, N781, N1602, N28);
xor XOR2 (N10898, N10885, N9098);
and AND2 (N10899, N10888, N3077);
or OR4 (N10900, N10895, N8926, N5502, N6704);
and AND2 (N10901, N10899, N10098);
xor XOR2 (N10902, N10893, N3340);
or OR4 (N10903, N10901, N9182, N5234, N1862);
nor NOR3 (N10904, N10886, N8445, N9619);
xor XOR2 (N10905, N10900, N7657);
or OR2 (N10906, N10894, N8095);
nand NAND3 (N10907, N10890, N4093, N6437);
nand NAND3 (N10908, N10903, N5410, N762);
nor NOR4 (N10909, N10904, N723, N391, N4637);
and AND4 (N10910, N10907, N10451, N7090, N4519);
or OR3 (N10911, N10908, N9249, N2170);
not NOT1 (N10912, N10910);
or OR2 (N10913, N10902, N3723);
not NOT1 (N10914, N10896);
and AND2 (N10915, N10906, N1706);
buf BUF1 (N10916, N10912);
nor NOR3 (N10917, N10905, N7909, N9173);
nor NOR4 (N10918, N10909, N8006, N8952, N635);
and AND4 (N10919, N10916, N9158, N10288, N1590);
xor XOR2 (N10920, N10917, N10710);
not NOT1 (N10921, N10883);
and AND2 (N10922, N10914, N1699);
not NOT1 (N10923, N10915);
nand NAND4 (N10924, N10922, N3277, N9851, N2507);
xor XOR2 (N10925, N10913, N1874);
not NOT1 (N10926, N10923);
nor NOR4 (N10927, N10921, N1946, N7442, N10027);
and AND2 (N10928, N10924, N9810);
buf BUF1 (N10929, N10928);
xor XOR2 (N10930, N10898, N9430);
or OR4 (N10931, N10926, N3578, N5219, N8687);
nor NOR2 (N10932, N10897, N2623);
xor XOR2 (N10933, N10925, N4786);
not NOT1 (N10934, N10930);
nor NOR4 (N10935, N10932, N10136, N10679, N1602);
or OR3 (N10936, N10929, N4945, N10454);
nand NAND2 (N10937, N10919, N7926);
and AND2 (N10938, N10937, N846);
and AND2 (N10939, N10927, N2771);
nor NOR4 (N10940, N10936, N328, N6056, N10464);
or OR3 (N10941, N10931, N2967, N6215);
xor XOR2 (N10942, N10918, N2096);
xor XOR2 (N10943, N10941, N7925);
and AND2 (N10944, N10911, N3518);
xor XOR2 (N10945, N10938, N4975);
not NOT1 (N10946, N10944);
or OR2 (N10947, N10943, N8555);
not NOT1 (N10948, N10940);
and AND2 (N10949, N10947, N4813);
or OR2 (N10950, N10939, N3921);
buf BUF1 (N10951, N10946);
nor NOR4 (N10952, N10933, N1620, N5556, N1195);
buf BUF1 (N10953, N10945);
not NOT1 (N10954, N10935);
nand NAND3 (N10955, N10954, N3495, N5348);
not NOT1 (N10956, N10942);
and AND2 (N10957, N10951, N5751);
nor NOR3 (N10958, N10952, N5742, N1261);
or OR4 (N10959, N10956, N4417, N5937, N5288);
or OR3 (N10960, N10950, N8449, N10754);
nand NAND4 (N10961, N10958, N3079, N5301, N9406);
xor XOR2 (N10962, N10949, N6436);
nor NOR3 (N10963, N10920, N977, N3650);
xor XOR2 (N10964, N10934, N7007);
buf BUF1 (N10965, N10961);
nand NAND2 (N10966, N10953, N131);
nand NAND3 (N10967, N10965, N9177, N1588);
or OR2 (N10968, N10963, N922);
nor NOR2 (N10969, N10960, N1971);
not NOT1 (N10970, N10969);
xor XOR2 (N10971, N10964, N8747);
and AND2 (N10972, N10948, N4875);
nor NOR4 (N10973, N10967, N9233, N241, N5500);
nand NAND3 (N10974, N10959, N4397, N548);
nor NOR4 (N10975, N10974, N6192, N6356, N7287);
or OR3 (N10976, N10972, N1254, N3104);
and AND2 (N10977, N10966, N4837);
nor NOR4 (N10978, N10955, N7287, N5921, N4387);
not NOT1 (N10979, N10976);
nor NOR2 (N10980, N10970, N9550);
not NOT1 (N10981, N10971);
and AND3 (N10982, N10962, N1046, N7778);
nand NAND2 (N10983, N10977, N9215);
or OR4 (N10984, N10979, N732, N4278, N5886);
nand NAND3 (N10985, N10980, N752, N8418);
nand NAND3 (N10986, N10984, N934, N5545);
xor XOR2 (N10987, N10957, N8927);
not NOT1 (N10988, N10978);
not NOT1 (N10989, N10973);
nor NOR3 (N10990, N10983, N4147, N9294);
xor XOR2 (N10991, N10989, N9072);
xor XOR2 (N10992, N10986, N10289);
nand NAND2 (N10993, N10990, N7386);
or OR4 (N10994, N10991, N9616, N9486, N10303);
nand NAND2 (N10995, N10988, N9547);
nand NAND2 (N10996, N10982, N8219);
xor XOR2 (N10997, N10985, N848);
not NOT1 (N10998, N10987);
and AND4 (N10999, N10996, N6296, N1526, N1070);
and AND2 (N11000, N10997, N6503);
or OR2 (N11001, N11000, N4116);
buf BUF1 (N11002, N10968);
xor XOR2 (N11003, N10992, N9249);
not NOT1 (N11004, N10975);
not NOT1 (N11005, N11002);
nand NAND3 (N11006, N10981, N1752, N10919);
nand NAND3 (N11007, N11003, N3085, N7965);
xor XOR2 (N11008, N11001, N1773);
not NOT1 (N11009, N11006);
xor XOR2 (N11010, N11004, N2649);
buf BUF1 (N11011, N10995);
and AND2 (N11012, N11011, N4822);
nor NOR4 (N11013, N10999, N4755, N10047, N6067);
xor XOR2 (N11014, N10998, N3352);
xor XOR2 (N11015, N11005, N3500);
buf BUF1 (N11016, N10994);
buf BUF1 (N11017, N11016);
not NOT1 (N11018, N11015);
xor XOR2 (N11019, N11013, N6607);
nor NOR2 (N11020, N11017, N6872);
xor XOR2 (N11021, N11007, N7067);
and AND4 (N11022, N11014, N1818, N5904, N9987);
buf BUF1 (N11023, N11012);
and AND2 (N11024, N11023, N1281);
not NOT1 (N11025, N10993);
and AND4 (N11026, N11010, N6918, N10674, N9100);
not NOT1 (N11027, N11022);
buf BUF1 (N11028, N11021);
buf BUF1 (N11029, N11027);
nand NAND3 (N11030, N11029, N10313, N10373);
nor NOR2 (N11031, N11019, N607);
xor XOR2 (N11032, N11008, N6039);
nand NAND3 (N11033, N11026, N3299, N10521);
not NOT1 (N11034, N11033);
not NOT1 (N11035, N11032);
nand NAND2 (N11036, N11009, N5629);
nand NAND3 (N11037, N11020, N10964, N67);
xor XOR2 (N11038, N11024, N5794);
nor NOR3 (N11039, N11018, N10086, N1912);
xor XOR2 (N11040, N11035, N10106);
and AND2 (N11041, N11030, N10044);
nor NOR2 (N11042, N11025, N7794);
buf BUF1 (N11043, N11031);
nand NAND4 (N11044, N11028, N4770, N7085, N1185);
buf BUF1 (N11045, N11044);
buf BUF1 (N11046, N11045);
nand NAND4 (N11047, N11040, N5917, N4875, N7168);
not NOT1 (N11048, N11034);
buf BUF1 (N11049, N11043);
nor NOR2 (N11050, N11041, N8211);
nor NOR3 (N11051, N11046, N2156, N8828);
nor NOR4 (N11052, N11047, N2857, N2844, N10864);
or OR4 (N11053, N11050, N64, N10819, N74);
xor XOR2 (N11054, N11042, N10741);
buf BUF1 (N11055, N11038);
xor XOR2 (N11056, N11037, N8137);
nand NAND2 (N11057, N11048, N2800);
nand NAND2 (N11058, N11051, N2106);
not NOT1 (N11059, N11052);
buf BUF1 (N11060, N11058);
nand NAND3 (N11061, N11056, N4010, N10211);
xor XOR2 (N11062, N11053, N3384);
nor NOR3 (N11063, N11059, N4865, N9503);
xor XOR2 (N11064, N11055, N3939);
or OR4 (N11065, N11054, N114, N3753, N3307);
nor NOR3 (N11066, N11063, N1718, N10877);
or OR2 (N11067, N11064, N8919);
nand NAND2 (N11068, N11062, N8016);
nand NAND4 (N11069, N11067, N7370, N8935, N8935);
xor XOR2 (N11070, N11066, N4571);
or OR2 (N11071, N11061, N6800);
and AND4 (N11072, N11070, N1719, N3797, N8281);
or OR2 (N11073, N11065, N3567);
or OR4 (N11074, N11060, N7015, N1088, N5985);
nand NAND2 (N11075, N11049, N2911);
or OR2 (N11076, N11057, N5599);
or OR2 (N11077, N11075, N5999);
xor XOR2 (N11078, N11069, N6015);
or OR2 (N11079, N11068, N4672);
buf BUF1 (N11080, N11073);
not NOT1 (N11081, N11036);
xor XOR2 (N11082, N11081, N2560);
nand NAND3 (N11083, N11074, N8309, N10050);
and AND4 (N11084, N11078, N2423, N6243, N10848);
buf BUF1 (N11085, N11072);
not NOT1 (N11086, N11079);
nor NOR3 (N11087, N11071, N6747, N5714);
xor XOR2 (N11088, N11076, N5742);
not NOT1 (N11089, N11083);
or OR2 (N11090, N11077, N2109);
nor NOR2 (N11091, N11088, N3397);
nor NOR2 (N11092, N11090, N7978);
xor XOR2 (N11093, N11091, N5127);
nand NAND2 (N11094, N11080, N3954);
nand NAND3 (N11095, N11084, N2152, N9422);
buf BUF1 (N11096, N11094);
nor NOR2 (N11097, N11086, N6830);
nor NOR2 (N11098, N11096, N7286);
and AND3 (N11099, N11092, N6135, N5083);
nor NOR4 (N11100, N11099, N4591, N5720, N8230);
buf BUF1 (N11101, N11087);
xor XOR2 (N11102, N11101, N9586);
buf BUF1 (N11103, N11093);
nor NOR4 (N11104, N11039, N4115, N6576, N3819);
and AND3 (N11105, N11102, N242, N1510);
buf BUF1 (N11106, N11103);
nor NOR4 (N11107, N11082, N8047, N10901, N712);
not NOT1 (N11108, N11095);
not NOT1 (N11109, N11104);
xor XOR2 (N11110, N11098, N11049);
not NOT1 (N11111, N11108);
nor NOR2 (N11112, N11100, N5220);
nand NAND3 (N11113, N11106, N10404, N8514);
nor NOR3 (N11114, N11109, N814, N10840);
or OR2 (N11115, N11114, N1721);
and AND4 (N11116, N11107, N6973, N8274, N5484);
and AND2 (N11117, N11089, N7700);
nor NOR4 (N11118, N11085, N10848, N683, N1479);
nand NAND2 (N11119, N11115, N2504);
and AND2 (N11120, N11097, N3791);
xor XOR2 (N11121, N11116, N6919);
buf BUF1 (N11122, N11110);
nand NAND2 (N11123, N11118, N2116);
buf BUF1 (N11124, N11111);
and AND3 (N11125, N11112, N7892, N6514);
not NOT1 (N11126, N11105);
xor XOR2 (N11127, N11124, N9683);
or OR3 (N11128, N11117, N9308, N8225);
not NOT1 (N11129, N11122);
xor XOR2 (N11130, N11129, N10337);
nand NAND4 (N11131, N11125, N5328, N3727, N273);
not NOT1 (N11132, N11130);
not NOT1 (N11133, N11127);
or OR4 (N11134, N11120, N991, N9706, N9808);
not NOT1 (N11135, N11121);
nand NAND3 (N11136, N11135, N9352, N304);
or OR4 (N11137, N11128, N8718, N9320, N2196);
xor XOR2 (N11138, N11123, N7887);
or OR4 (N11139, N11138, N8802, N10820, N6297);
nand NAND2 (N11140, N11133, N10789);
and AND4 (N11141, N11136, N9385, N7917, N4430);
nand NAND4 (N11142, N11141, N40, N1591, N7465);
and AND4 (N11143, N11137, N9601, N5180, N4726);
nand NAND3 (N11144, N11142, N4625, N6592);
xor XOR2 (N11145, N11131, N1984);
or OR3 (N11146, N11144, N8870, N6297);
nor NOR4 (N11147, N11126, N4812, N630, N11123);
nand NAND2 (N11148, N11147, N684);
and AND3 (N11149, N11113, N10510, N3804);
nand NAND2 (N11150, N11148, N7507);
or OR2 (N11151, N11139, N232);
or OR2 (N11152, N11140, N8715);
or OR2 (N11153, N11152, N361);
xor XOR2 (N11154, N11143, N6372);
xor XOR2 (N11155, N11149, N2849);
buf BUF1 (N11156, N11132);
xor XOR2 (N11157, N11145, N9914);
or OR3 (N11158, N11119, N8317, N11106);
or OR3 (N11159, N11155, N5646, N6134);
not NOT1 (N11160, N11134);
not NOT1 (N11161, N11150);
nor NOR3 (N11162, N11156, N5651, N8634);
not NOT1 (N11163, N11162);
not NOT1 (N11164, N11163);
and AND2 (N11165, N11154, N5777);
buf BUF1 (N11166, N11157);
not NOT1 (N11167, N11153);
xor XOR2 (N11168, N11159, N1674);
or OR4 (N11169, N11166, N6069, N2978, N5349);
xor XOR2 (N11170, N11146, N6838);
xor XOR2 (N11171, N11167, N2545);
not NOT1 (N11172, N11158);
nor NOR4 (N11173, N11168, N10307, N776, N243);
nor NOR2 (N11174, N11171, N5266);
not NOT1 (N11175, N11164);
nor NOR3 (N11176, N11174, N6818, N7128);
buf BUF1 (N11177, N11176);
nand NAND4 (N11178, N11175, N6437, N8160, N6565);
xor XOR2 (N11179, N11172, N2915);
and AND4 (N11180, N11178, N3306, N6969, N3355);
xor XOR2 (N11181, N11180, N8769);
not NOT1 (N11182, N11181);
not NOT1 (N11183, N11169);
and AND4 (N11184, N11183, N4366, N2225, N1833);
and AND2 (N11185, N11165, N9741);
or OR3 (N11186, N11185, N6750, N7510);
or OR4 (N11187, N11182, N9255, N10728, N4509);
buf BUF1 (N11188, N11161);
nand NAND3 (N11189, N11184, N4083, N10162);
or OR3 (N11190, N11187, N2345, N3884);
xor XOR2 (N11191, N11170, N9034);
buf BUF1 (N11192, N11151);
not NOT1 (N11193, N11177);
nand NAND2 (N11194, N11193, N2259);
nand NAND2 (N11195, N11192, N6701);
or OR2 (N11196, N11160, N1403);
buf BUF1 (N11197, N11173);
nand NAND2 (N11198, N11188, N4929);
nand NAND3 (N11199, N11194, N6657, N2709);
xor XOR2 (N11200, N11198, N3808);
xor XOR2 (N11201, N11196, N7618);
xor XOR2 (N11202, N11199, N2208);
or OR4 (N11203, N11189, N554, N1177, N4768);
nand NAND4 (N11204, N11203, N4572, N7682, N413);
nand NAND4 (N11205, N11200, N7323, N10227, N5854);
not NOT1 (N11206, N11197);
and AND3 (N11207, N11206, N10233, N9707);
xor XOR2 (N11208, N11201, N8954);
or OR3 (N11209, N11191, N9140, N1417);
xor XOR2 (N11210, N11202, N4984);
or OR3 (N11211, N11208, N9719, N6449);
nor NOR4 (N11212, N11207, N6426, N3157, N3757);
or OR2 (N11213, N11212, N3875);
buf BUF1 (N11214, N11210);
buf BUF1 (N11215, N11205);
xor XOR2 (N11216, N11186, N5531);
not NOT1 (N11217, N11214);
buf BUF1 (N11218, N11217);
nor NOR3 (N11219, N11195, N9678, N8825);
xor XOR2 (N11220, N11190, N3104);
or OR4 (N11221, N11204, N7554, N1197, N4396);
xor XOR2 (N11222, N11221, N6670);
and AND4 (N11223, N11215, N9659, N5868, N10261);
not NOT1 (N11224, N11222);
nor NOR2 (N11225, N11223, N7188);
nand NAND2 (N11226, N11216, N2345);
not NOT1 (N11227, N11213);
nand NAND2 (N11228, N11220, N3080);
not NOT1 (N11229, N11218);
xor XOR2 (N11230, N11179, N10673);
nor NOR4 (N11231, N11219, N8857, N1414, N10189);
not NOT1 (N11232, N11230);
buf BUF1 (N11233, N11211);
buf BUF1 (N11234, N11209);
buf BUF1 (N11235, N11229);
nand NAND3 (N11236, N11228, N1089, N7982);
not NOT1 (N11237, N11236);
and AND3 (N11238, N11235, N10413, N912);
nor NOR3 (N11239, N11227, N4293, N8650);
buf BUF1 (N11240, N11238);
and AND3 (N11241, N11232, N10163, N251);
nand NAND2 (N11242, N11226, N7267);
not NOT1 (N11243, N11233);
nor NOR3 (N11244, N11243, N10728, N6367);
not NOT1 (N11245, N11244);
nand NAND2 (N11246, N11234, N9713);
or OR3 (N11247, N11239, N7227, N9509);
not NOT1 (N11248, N11247);
and AND2 (N11249, N11246, N1810);
nand NAND4 (N11250, N11237, N1832, N9763, N5293);
nor NOR3 (N11251, N11224, N384, N3275);
nand NAND3 (N11252, N11241, N5327, N66);
nor NOR4 (N11253, N11249, N2687, N6416, N7815);
xor XOR2 (N11254, N11250, N4038);
or OR4 (N11255, N11240, N3237, N10308, N8006);
or OR4 (N11256, N11254, N4159, N2368, N10467);
xor XOR2 (N11257, N11252, N10393);
nand NAND2 (N11258, N11256, N8491);
nor NOR3 (N11259, N11248, N4068, N10542);
or OR2 (N11260, N11245, N4937);
nor NOR2 (N11261, N11225, N3343);
xor XOR2 (N11262, N11251, N7692);
nor NOR2 (N11263, N11253, N5702);
or OR3 (N11264, N11257, N6286, N1300);
not NOT1 (N11265, N11258);
nand NAND2 (N11266, N11264, N3736);
or OR3 (N11267, N11263, N4989, N4293);
nand NAND4 (N11268, N11262, N10605, N506, N10437);
and AND4 (N11269, N11259, N11258, N10051, N771);
nor NOR4 (N11270, N11260, N7174, N10874, N6090);
buf BUF1 (N11271, N11265);
xor XOR2 (N11272, N11242, N8425);
buf BUF1 (N11273, N11271);
xor XOR2 (N11274, N11269, N9525);
or OR4 (N11275, N11274, N1371, N6482, N5692);
buf BUF1 (N11276, N11255);
and AND3 (N11277, N11268, N5815, N9275);
xor XOR2 (N11278, N11277, N9125);
nor NOR3 (N11279, N11275, N4005, N9236);
not NOT1 (N11280, N11276);
not NOT1 (N11281, N11267);
and AND3 (N11282, N11281, N7626, N434);
not NOT1 (N11283, N11280);
buf BUF1 (N11284, N11283);
nor NOR3 (N11285, N11270, N113, N1390);
buf BUF1 (N11286, N11278);
nand NAND3 (N11287, N11284, N8751, N9057);
or OR2 (N11288, N11273, N9633);
or OR3 (N11289, N11287, N4471, N467);
nand NAND3 (N11290, N11285, N1082, N3106);
xor XOR2 (N11291, N11261, N37);
not NOT1 (N11292, N11282);
xor XOR2 (N11293, N11279, N7948);
xor XOR2 (N11294, N11293, N1737);
buf BUF1 (N11295, N11286);
and AND3 (N11296, N11294, N897, N4395);
buf BUF1 (N11297, N11272);
buf BUF1 (N11298, N11288);
buf BUF1 (N11299, N11295);
not NOT1 (N11300, N11296);
nor NOR4 (N11301, N11299, N5703, N11231, N10437);
xor XOR2 (N11302, N294, N5735);
buf BUF1 (N11303, N11292);
buf BUF1 (N11304, N11291);
xor XOR2 (N11305, N11301, N1804);
not NOT1 (N11306, N11297);
or OR3 (N11307, N11300, N10802, N4793);
and AND4 (N11308, N11266, N3900, N4241, N3554);
buf BUF1 (N11309, N11308);
nor NOR4 (N11310, N11298, N5620, N926, N10381);
buf BUF1 (N11311, N11310);
and AND2 (N11312, N11305, N7821);
or OR4 (N11313, N11290, N7627, N3172, N9664);
or OR2 (N11314, N11309, N5401);
nand NAND3 (N11315, N11306, N11110, N3414);
xor XOR2 (N11316, N11311, N2689);
nand NAND2 (N11317, N11289, N2523);
buf BUF1 (N11318, N11315);
nand NAND2 (N11319, N11318, N4544);
xor XOR2 (N11320, N11302, N8139);
nor NOR2 (N11321, N11317, N10835);
not NOT1 (N11322, N11321);
buf BUF1 (N11323, N11303);
xor XOR2 (N11324, N11316, N3131);
xor XOR2 (N11325, N11319, N1605);
not NOT1 (N11326, N11304);
xor XOR2 (N11327, N11325, N10540);
and AND4 (N11328, N11322, N8658, N8134, N7062);
nand NAND4 (N11329, N11314, N6434, N10495, N5542);
nor NOR3 (N11330, N11312, N11171, N4843);
not NOT1 (N11331, N11330);
xor XOR2 (N11332, N11326, N8990);
nor NOR2 (N11333, N11328, N9316);
or OR3 (N11334, N11332, N1780, N5527);
xor XOR2 (N11335, N11313, N9468);
xor XOR2 (N11336, N11334, N6876);
and AND3 (N11337, N11327, N8613, N8431);
or OR2 (N11338, N11335, N4419);
or OR4 (N11339, N11320, N7546, N9181, N170);
nand NAND3 (N11340, N11338, N9057, N9967);
and AND4 (N11341, N11336, N7080, N4221, N7957);
buf BUF1 (N11342, N11323);
nand NAND4 (N11343, N11324, N7630, N8891, N3993);
nor NOR2 (N11344, N11342, N8687);
and AND2 (N11345, N11340, N5656);
and AND4 (N11346, N11331, N5960, N11186, N260);
not NOT1 (N11347, N11307);
and AND4 (N11348, N11333, N8105, N6434, N4414);
xor XOR2 (N11349, N11339, N10127);
nand NAND2 (N11350, N11345, N10759);
or OR4 (N11351, N11350, N3612, N8589, N1479);
nand NAND4 (N11352, N11344, N9735, N687, N7957);
xor XOR2 (N11353, N11337, N6703);
buf BUF1 (N11354, N11351);
not NOT1 (N11355, N11329);
xor XOR2 (N11356, N11352, N10667);
xor XOR2 (N11357, N11343, N3162);
xor XOR2 (N11358, N11355, N6284);
nor NOR3 (N11359, N11353, N11182, N4812);
or OR3 (N11360, N11359, N2794, N3110);
buf BUF1 (N11361, N11354);
nand NAND2 (N11362, N11349, N1916);
nand NAND3 (N11363, N11346, N6599, N4520);
and AND3 (N11364, N11357, N2529, N8290);
nor NOR4 (N11365, N11341, N4586, N8837, N9992);
nor NOR3 (N11366, N11358, N3189, N9918);
and AND3 (N11367, N11356, N7852, N9647);
nor NOR2 (N11368, N11367, N2198);
not NOT1 (N11369, N11348);
nand NAND2 (N11370, N11362, N1885);
or OR3 (N11371, N11360, N2533, N6270);
and AND2 (N11372, N11365, N3125);
or OR3 (N11373, N11371, N7515, N5832);
or OR3 (N11374, N11370, N4009, N5152);
xor XOR2 (N11375, N11368, N8785);
not NOT1 (N11376, N11373);
xor XOR2 (N11377, N11376, N5771);
nand NAND3 (N11378, N11363, N3573, N2825);
nor NOR2 (N11379, N11347, N4565);
xor XOR2 (N11380, N11379, N5390);
and AND4 (N11381, N11378, N6408, N325, N11272);
nor NOR4 (N11382, N11366, N7252, N7374, N8281);
buf BUF1 (N11383, N11381);
or OR2 (N11384, N11361, N9827);
xor XOR2 (N11385, N11369, N3259);
nand NAND3 (N11386, N11372, N7875, N1034);
nand NAND4 (N11387, N11384, N10329, N4034, N9571);
and AND2 (N11388, N11364, N393);
buf BUF1 (N11389, N11377);
and AND2 (N11390, N11385, N3079);
not NOT1 (N11391, N11380);
xor XOR2 (N11392, N11386, N1364);
nor NOR4 (N11393, N11374, N1555, N3309, N5539);
nor NOR4 (N11394, N11383, N3810, N11277, N4732);
buf BUF1 (N11395, N11390);
nand NAND3 (N11396, N11387, N1932, N10138);
not NOT1 (N11397, N11394);
and AND2 (N11398, N11382, N448);
nor NOR3 (N11399, N11397, N10944, N20);
nor NOR4 (N11400, N11393, N10439, N7075, N10142);
and AND4 (N11401, N11391, N5716, N3394, N4645);
xor XOR2 (N11402, N11401, N11117);
buf BUF1 (N11403, N11399);
or OR4 (N11404, N11389, N10145, N10457, N9259);
nor NOR2 (N11405, N11388, N4863);
buf BUF1 (N11406, N11398);
nor NOR4 (N11407, N11405, N2197, N9875, N6673);
buf BUF1 (N11408, N11407);
and AND2 (N11409, N11408, N10571);
nor NOR3 (N11410, N11403, N1996, N1030);
nand NAND2 (N11411, N11392, N1077);
and AND4 (N11412, N11409, N7246, N477, N7472);
not NOT1 (N11413, N11404);
and AND3 (N11414, N11411, N10907, N6696);
nand NAND2 (N11415, N11400, N4971);
nor NOR4 (N11416, N11375, N323, N10593, N11382);
and AND4 (N11417, N11395, N9133, N743, N2067);
xor XOR2 (N11418, N11396, N1389);
or OR2 (N11419, N11412, N2554);
xor XOR2 (N11420, N11414, N10645);
not NOT1 (N11421, N11415);
or OR3 (N11422, N11419, N9113, N3652);
nor NOR3 (N11423, N11418, N2640, N9976);
xor XOR2 (N11424, N11416, N9261);
xor XOR2 (N11425, N11421, N6723);
or OR3 (N11426, N11417, N601, N1618);
nand NAND2 (N11427, N11424, N3858);
or OR2 (N11428, N11423, N3563);
nor NOR4 (N11429, N11428, N10311, N4277, N10176);
not NOT1 (N11430, N11422);
nor NOR3 (N11431, N11427, N942, N8310);
nand NAND2 (N11432, N11431, N2583);
or OR3 (N11433, N11406, N810, N2956);
or OR4 (N11434, N11420, N979, N682, N10811);
buf BUF1 (N11435, N11430);
buf BUF1 (N11436, N11402);
buf BUF1 (N11437, N11434);
nand NAND3 (N11438, N11432, N6522, N3587);
or OR2 (N11439, N11426, N6963);
xor XOR2 (N11440, N11410, N3904);
buf BUF1 (N11441, N11435);
nor NOR2 (N11442, N11438, N3424);
not NOT1 (N11443, N11442);
xor XOR2 (N11444, N11429, N423);
or OR3 (N11445, N11433, N10218, N5416);
or OR2 (N11446, N11439, N5124);
xor XOR2 (N11447, N11446, N1861);
buf BUF1 (N11448, N11413);
nor NOR3 (N11449, N11440, N10984, N10192);
buf BUF1 (N11450, N11448);
nor NOR3 (N11451, N11447, N3703, N563);
buf BUF1 (N11452, N11449);
or OR3 (N11453, N11451, N7263, N11109);
nand NAND2 (N11454, N11445, N5368);
nor NOR4 (N11455, N11436, N3219, N4445, N2758);
not NOT1 (N11456, N11452);
and AND2 (N11457, N11455, N2560);
nand NAND3 (N11458, N11457, N6092, N10695);
and AND3 (N11459, N11425, N157, N4548);
not NOT1 (N11460, N11441);
nand NAND2 (N11461, N11458, N7998);
nor NOR2 (N11462, N11461, N8320);
buf BUF1 (N11463, N11454);
nand NAND4 (N11464, N11453, N10721, N8469, N4690);
nand NAND2 (N11465, N11444, N14);
and AND2 (N11466, N11464, N8387);
xor XOR2 (N11467, N11443, N8534);
nor NOR4 (N11468, N11460, N9302, N1896, N878);
nor NOR2 (N11469, N11437, N5367);
nor NOR2 (N11470, N11466, N4710);
not NOT1 (N11471, N11463);
nand NAND3 (N11472, N11469, N10303, N223);
nand NAND4 (N11473, N11456, N5355, N6036, N4020);
nor NOR3 (N11474, N11468, N10001, N1351);
nor NOR3 (N11475, N11467, N7283, N8182);
not NOT1 (N11476, N11470);
xor XOR2 (N11477, N11459, N9725);
nand NAND3 (N11478, N11471, N8618, N5859);
and AND4 (N11479, N11476, N7770, N2464, N9638);
not NOT1 (N11480, N11475);
nand NAND2 (N11481, N11473, N9930);
not NOT1 (N11482, N11480);
nand NAND2 (N11483, N11474, N7595);
or OR3 (N11484, N11477, N9357, N6607);
nor NOR3 (N11485, N11481, N2562, N6529);
nand NAND4 (N11486, N11484, N8396, N6928, N10907);
and AND3 (N11487, N11479, N7901, N2702);
nand NAND2 (N11488, N11485, N1561);
nor NOR3 (N11489, N11486, N1753, N11026);
and AND4 (N11490, N11488, N5540, N1438, N7056);
nand NAND2 (N11491, N11450, N7140);
buf BUF1 (N11492, N11465);
or OR4 (N11493, N11487, N8152, N7938, N9729);
or OR3 (N11494, N11482, N6132, N4669);
xor XOR2 (N11495, N11478, N10381);
or OR4 (N11496, N11472, N10815, N6305, N775);
and AND4 (N11497, N11489, N1217, N5594, N6159);
xor XOR2 (N11498, N11483, N557);
nor NOR4 (N11499, N11492, N583, N9550, N7312);
buf BUF1 (N11500, N11493);
buf BUF1 (N11501, N11490);
nand NAND2 (N11502, N11494, N6933);
nand NAND4 (N11503, N11498, N11144, N10006, N11134);
or OR2 (N11504, N11499, N7047);
and AND3 (N11505, N11503, N9382, N7754);
not NOT1 (N11506, N11497);
not NOT1 (N11507, N11496);
nor NOR3 (N11508, N11506, N7208, N4270);
nand NAND4 (N11509, N11491, N10269, N10834, N4234);
or OR3 (N11510, N11509, N3719, N3780);
nor NOR4 (N11511, N11505, N779, N8305, N232);
not NOT1 (N11512, N11495);
nand NAND4 (N11513, N11502, N9438, N8906, N913);
xor XOR2 (N11514, N11512, N2416);
nor NOR3 (N11515, N11501, N6373, N7467);
or OR4 (N11516, N11500, N8536, N3146, N6351);
buf BUF1 (N11517, N11513);
xor XOR2 (N11518, N11517, N2940);
not NOT1 (N11519, N11511);
not NOT1 (N11520, N11514);
nor NOR2 (N11521, N11510, N4764);
not NOT1 (N11522, N11518);
or OR4 (N11523, N11515, N5657, N7139, N9611);
or OR4 (N11524, N11462, N1051, N1759, N1682);
buf BUF1 (N11525, N11504);
nor NOR2 (N11526, N11525, N9171);
xor XOR2 (N11527, N11524, N7444);
nor NOR2 (N11528, N11519, N1892);
nand NAND3 (N11529, N11527, N2752, N8195);
buf BUF1 (N11530, N11522);
not NOT1 (N11531, N11528);
buf BUF1 (N11532, N11520);
or OR2 (N11533, N11521, N1474);
not NOT1 (N11534, N11507);
nor NOR3 (N11535, N11523, N4485, N5545);
nor NOR4 (N11536, N11535, N8253, N1633, N2251);
nor NOR2 (N11537, N11534, N3573);
nor NOR4 (N11538, N11532, N8246, N8177, N10832);
nor NOR2 (N11539, N11538, N6392);
and AND3 (N11540, N11516, N934, N9842);
not NOT1 (N11541, N11530);
and AND2 (N11542, N11508, N4680);
nor NOR4 (N11543, N11531, N8526, N7478, N4912);
or OR2 (N11544, N11540, N437);
nor NOR2 (N11545, N11536, N44);
or OR4 (N11546, N11541, N10545, N1219, N5016);
nand NAND3 (N11547, N11545, N5876, N10977);
nor NOR3 (N11548, N11543, N9819, N5168);
nor NOR3 (N11549, N11542, N11361, N1897);
and AND4 (N11550, N11537, N11263, N5172, N4610);
buf BUF1 (N11551, N11548);
or OR4 (N11552, N11549, N10423, N4401, N5366);
xor XOR2 (N11553, N11529, N2930);
nor NOR4 (N11554, N11547, N5406, N3871, N4137);
not NOT1 (N11555, N11551);
not NOT1 (N11556, N11526);
or OR4 (N11557, N11550, N6397, N6713, N8067);
not NOT1 (N11558, N11557);
and AND3 (N11559, N11552, N5321, N6191);
or OR3 (N11560, N11533, N4968, N1363);
or OR4 (N11561, N11560, N9672, N7882, N6746);
nand NAND4 (N11562, N11553, N7490, N10404, N10099);
xor XOR2 (N11563, N11558, N7519);
or OR4 (N11564, N11563, N6084, N7894, N10218);
and AND3 (N11565, N11539, N909, N1731);
not NOT1 (N11566, N11556);
nand NAND2 (N11567, N11566, N5204);
xor XOR2 (N11568, N11562, N6947);
not NOT1 (N11569, N11555);
and AND2 (N11570, N11564, N2635);
nor NOR4 (N11571, N11565, N9239, N1850, N3893);
buf BUF1 (N11572, N11568);
nand NAND2 (N11573, N11569, N5546);
and AND4 (N11574, N11572, N8608, N9442, N5994);
buf BUF1 (N11575, N11567);
buf BUF1 (N11576, N11573);
not NOT1 (N11577, N11570);
and AND3 (N11578, N11574, N2233, N10575);
and AND4 (N11579, N11578, N468, N2701, N9754);
nand NAND2 (N11580, N11561, N10914);
or OR4 (N11581, N11576, N4228, N1841, N131);
and AND2 (N11582, N11577, N1029);
nand NAND3 (N11583, N11559, N10264, N7319);
or OR4 (N11584, N11546, N1022, N3413, N7893);
xor XOR2 (N11585, N11544, N6711);
nand NAND3 (N11586, N11580, N10409, N882);
not NOT1 (N11587, N11586);
xor XOR2 (N11588, N11581, N11036);
nand NAND3 (N11589, N11579, N8113, N7971);
or OR2 (N11590, N11584, N3970);
nor NOR2 (N11591, N11583, N4962);
buf BUF1 (N11592, N11588);
or OR3 (N11593, N11575, N6409, N11562);
nand NAND3 (N11594, N11592, N3217, N964);
not NOT1 (N11595, N11587);
nand NAND3 (N11596, N11594, N9601, N9404);
or OR3 (N11597, N11554, N7101, N534);
buf BUF1 (N11598, N11582);
xor XOR2 (N11599, N11571, N4386);
and AND3 (N11600, N11590, N7871, N6605);
or OR2 (N11601, N11598, N430);
nand NAND4 (N11602, N11597, N4084, N11021, N5560);
nand NAND4 (N11603, N11591, N9043, N11332, N8560);
buf BUF1 (N11604, N11599);
nand NAND2 (N11605, N11603, N2369);
nand NAND2 (N11606, N11604, N4614);
or OR3 (N11607, N11605, N5882, N4014);
nor NOR3 (N11608, N11595, N6695, N662);
xor XOR2 (N11609, N11593, N4438);
nor NOR2 (N11610, N11589, N2619);
buf BUF1 (N11611, N11608);
buf BUF1 (N11612, N11610);
nor NOR2 (N11613, N11609, N10228);
buf BUF1 (N11614, N11600);
xor XOR2 (N11615, N11607, N3287);
or OR4 (N11616, N11585, N4000, N7283, N3189);
buf BUF1 (N11617, N11602);
buf BUF1 (N11618, N11611);
xor XOR2 (N11619, N11606, N10522);
nor NOR4 (N11620, N11596, N8638, N8257, N9104);
not NOT1 (N11621, N11616);
and AND2 (N11622, N11614, N9108);
and AND4 (N11623, N11612, N540, N9059, N2921);
and AND2 (N11624, N11613, N2788);
xor XOR2 (N11625, N11615, N9729);
nand NAND4 (N11626, N11619, N9987, N6455, N858);
buf BUF1 (N11627, N11618);
nand NAND2 (N11628, N11620, N1166);
not NOT1 (N11629, N11621);
nand NAND3 (N11630, N11627, N1957, N9644);
and AND4 (N11631, N11623, N815, N5517, N5391);
nor NOR2 (N11632, N11601, N10842);
xor XOR2 (N11633, N11630, N3877);
nand NAND2 (N11634, N11625, N621);
nor NOR3 (N11635, N11624, N1650, N5903);
xor XOR2 (N11636, N11631, N8869);
or OR3 (N11637, N11628, N3217, N2519);
xor XOR2 (N11638, N11636, N3404);
buf BUF1 (N11639, N11626);
not NOT1 (N11640, N11639);
nor NOR4 (N11641, N11634, N2215, N7660, N666);
not NOT1 (N11642, N11635);
not NOT1 (N11643, N11641);
not NOT1 (N11644, N11633);
nor NOR2 (N11645, N11640, N214);
or OR4 (N11646, N11632, N1753, N10446, N11036);
nand NAND4 (N11647, N11617, N7659, N11479, N10397);
not NOT1 (N11648, N11637);
not NOT1 (N11649, N11629);
and AND2 (N11650, N11648, N4912);
and AND4 (N11651, N11647, N11062, N2880, N5582);
and AND3 (N11652, N11643, N6737, N193);
nand NAND3 (N11653, N11650, N2580, N8896);
and AND4 (N11654, N11653, N10773, N3633, N9986);
xor XOR2 (N11655, N11638, N6616);
xor XOR2 (N11656, N11622, N1888);
nor NOR2 (N11657, N11654, N9158);
buf BUF1 (N11658, N11652);
nand NAND4 (N11659, N11642, N5318, N11582, N6215);
buf BUF1 (N11660, N11655);
xor XOR2 (N11661, N11649, N10223);
and AND2 (N11662, N11645, N457);
nand NAND3 (N11663, N11656, N11224, N6780);
buf BUF1 (N11664, N11660);
or OR4 (N11665, N11661, N3550, N10647, N7749);
or OR3 (N11666, N11646, N10127, N4712);
buf BUF1 (N11667, N11651);
nor NOR4 (N11668, N11662, N6050, N11323, N8630);
nor NOR2 (N11669, N11644, N3488);
and AND2 (N11670, N11667, N8105);
buf BUF1 (N11671, N11657);
nand NAND2 (N11672, N11671, N5509);
xor XOR2 (N11673, N11670, N7587);
and AND4 (N11674, N11663, N7605, N5797, N4701);
or OR3 (N11675, N11669, N5708, N9465);
and AND3 (N11676, N11658, N11469, N3178);
not NOT1 (N11677, N11674);
nor NOR4 (N11678, N11672, N8614, N517, N6232);
xor XOR2 (N11679, N11664, N11199);
or OR3 (N11680, N11678, N11024, N8409);
buf BUF1 (N11681, N11676);
or OR2 (N11682, N11675, N519);
nor NOR4 (N11683, N11680, N1586, N7329, N1814);
nor NOR4 (N11684, N11665, N8590, N8440, N3449);
and AND4 (N11685, N11677, N7590, N9523, N5385);
nor NOR4 (N11686, N11681, N5251, N6675, N5328);
nand NAND2 (N11687, N11668, N6750);
xor XOR2 (N11688, N11666, N1220);
or OR3 (N11689, N11688, N5462, N3588);
buf BUF1 (N11690, N11689);
nor NOR3 (N11691, N11685, N111, N7815);
nand NAND3 (N11692, N11673, N2351, N5590);
nor NOR2 (N11693, N11684, N2123);
xor XOR2 (N11694, N11659, N10652);
nor NOR3 (N11695, N11690, N1813, N8842);
and AND3 (N11696, N11693, N8882, N4742);
and AND3 (N11697, N11679, N1783, N5747);
or OR4 (N11698, N11683, N5736, N9089, N2700);
nand NAND2 (N11699, N11694, N1451);
and AND4 (N11700, N11697, N5765, N10996, N7692);
and AND4 (N11701, N11700, N4571, N7469, N3674);
not NOT1 (N11702, N11682);
nand NAND2 (N11703, N11699, N11647);
nor NOR4 (N11704, N11695, N9066, N5007, N8591);
or OR4 (N11705, N11696, N3711, N6178, N3614);
buf BUF1 (N11706, N11702);
and AND2 (N11707, N11687, N9171);
xor XOR2 (N11708, N11704, N992);
or OR3 (N11709, N11692, N1118, N7185);
or OR2 (N11710, N11708, N11640);
nor NOR3 (N11711, N11706, N2232, N9707);
and AND2 (N11712, N11701, N9522);
nor NOR3 (N11713, N11710, N6907, N2287);
nor NOR2 (N11714, N11711, N351);
not NOT1 (N11715, N11705);
or OR4 (N11716, N11714, N1085, N3111, N1315);
not NOT1 (N11717, N11713);
xor XOR2 (N11718, N11709, N843);
or OR2 (N11719, N11703, N11593);
or OR2 (N11720, N11715, N8444);
xor XOR2 (N11721, N11716, N221);
xor XOR2 (N11722, N11718, N6664);
and AND2 (N11723, N11722, N10710);
nand NAND3 (N11724, N11707, N3651, N4790);
xor XOR2 (N11725, N11720, N8638);
or OR4 (N11726, N11698, N1812, N9221, N3723);
and AND2 (N11727, N11723, N3328);
nand NAND3 (N11728, N11712, N5852, N10419);
nor NOR3 (N11729, N11727, N5160, N4504);
buf BUF1 (N11730, N11726);
nor NOR4 (N11731, N11721, N8659, N8369, N5824);
nor NOR2 (N11732, N11691, N5561);
or OR2 (N11733, N11730, N9170);
nor NOR4 (N11734, N11686, N3293, N4244, N6246);
nand NAND2 (N11735, N11729, N4731);
or OR4 (N11736, N11735, N8642, N277, N6089);
nand NAND2 (N11737, N11734, N6433);
buf BUF1 (N11738, N11728);
buf BUF1 (N11739, N11724);
not NOT1 (N11740, N11733);
xor XOR2 (N11741, N11725, N6047);
xor XOR2 (N11742, N11739, N6323);
or OR4 (N11743, N11717, N3702, N127, N10351);
or OR3 (N11744, N11731, N7035, N2690);
or OR3 (N11745, N11738, N1857, N7466);
nor NOR3 (N11746, N11737, N8647, N325);
buf BUF1 (N11747, N11732);
and AND4 (N11748, N11719, N2201, N1036, N765);
nand NAND2 (N11749, N11740, N1605);
xor XOR2 (N11750, N11748, N3436);
not NOT1 (N11751, N11743);
nor NOR2 (N11752, N11745, N3828);
nor NOR2 (N11753, N11736, N7601);
not NOT1 (N11754, N11753);
xor XOR2 (N11755, N11749, N10496);
xor XOR2 (N11756, N11742, N8171);
nor NOR3 (N11757, N11756, N2445, N2197);
nor NOR2 (N11758, N11752, N2962);
and AND3 (N11759, N11755, N6997, N3153);
and AND3 (N11760, N11758, N11434, N159);
nand NAND2 (N11761, N11757, N4384);
xor XOR2 (N11762, N11760, N1111);
or OR3 (N11763, N11741, N2469, N7702);
nor NOR3 (N11764, N11750, N6937, N9119);
xor XOR2 (N11765, N11759, N9133);
nand NAND3 (N11766, N11764, N3739, N3174);
nor NOR4 (N11767, N11746, N2981, N11009, N1630);
xor XOR2 (N11768, N11744, N258);
and AND2 (N11769, N11763, N868);
xor XOR2 (N11770, N11769, N11410);
buf BUF1 (N11771, N11765);
and AND4 (N11772, N11754, N2539, N8294, N3427);
nand NAND3 (N11773, N11771, N5915, N7148);
buf BUF1 (N11774, N11767);
xor XOR2 (N11775, N11761, N1859);
nor NOR4 (N11776, N11773, N11620, N10606, N2645);
and AND3 (N11777, N11776, N9256, N219);
nor NOR4 (N11778, N11766, N7070, N3669, N8155);
nor NOR2 (N11779, N11775, N7417);
buf BUF1 (N11780, N11751);
or OR3 (N11781, N11778, N10768, N4896);
nand NAND2 (N11782, N11781, N1987);
and AND3 (N11783, N11747, N146, N8034);
nor NOR3 (N11784, N11768, N7422, N7914);
nor NOR4 (N11785, N11777, N11516, N5201, N3006);
xor XOR2 (N11786, N11782, N3799);
or OR2 (N11787, N11783, N11434);
and AND4 (N11788, N11779, N7253, N8293, N10395);
or OR3 (N11789, N11762, N5118, N6675);
buf BUF1 (N11790, N11786);
not NOT1 (N11791, N11784);
nor NOR4 (N11792, N11787, N3505, N144, N875);
not NOT1 (N11793, N11790);
nand NAND3 (N11794, N11793, N1956, N5907);
or OR4 (N11795, N11780, N8097, N8249, N9110);
nor NOR2 (N11796, N11788, N6084);
nand NAND2 (N11797, N11785, N5309);
and AND4 (N11798, N11770, N7061, N7433, N1628);
nor NOR2 (N11799, N11789, N5153);
not NOT1 (N11800, N11774);
buf BUF1 (N11801, N11796);
not NOT1 (N11802, N11799);
and AND3 (N11803, N11772, N5715, N10074);
or OR2 (N11804, N11797, N11538);
nand NAND4 (N11805, N11791, N7240, N39, N2871);
buf BUF1 (N11806, N11804);
xor XOR2 (N11807, N11795, N3905);
buf BUF1 (N11808, N11802);
nand NAND2 (N11809, N11807, N10392);
xor XOR2 (N11810, N11794, N444);
not NOT1 (N11811, N11798);
not NOT1 (N11812, N11806);
not NOT1 (N11813, N11812);
or OR4 (N11814, N11792, N9659, N6929, N7102);
nand NAND2 (N11815, N11809, N11075);
nand NAND3 (N11816, N11801, N772, N9884);
not NOT1 (N11817, N11814);
nand NAND4 (N11818, N11816, N2957, N2115, N6800);
nor NOR4 (N11819, N11805, N6340, N6088, N2485);
buf BUF1 (N11820, N11818);
nor NOR4 (N11821, N11815, N5350, N6707, N3496);
xor XOR2 (N11822, N11811, N5922);
or OR3 (N11823, N11821, N1468, N4590);
and AND2 (N11824, N11808, N6722);
buf BUF1 (N11825, N11817);
or OR2 (N11826, N11813, N11695);
nor NOR4 (N11827, N11823, N9793, N7310, N1843);
xor XOR2 (N11828, N11810, N7689);
and AND4 (N11829, N11820, N8905, N8372, N624);
not NOT1 (N11830, N11803);
xor XOR2 (N11831, N11824, N5933);
not NOT1 (N11832, N11830);
or OR3 (N11833, N11829, N1501, N10652);
xor XOR2 (N11834, N11826, N9862);
or OR4 (N11835, N11825, N926, N11455, N11299);
not NOT1 (N11836, N11832);
and AND3 (N11837, N11828, N2050, N9757);
buf BUF1 (N11838, N11833);
nand NAND3 (N11839, N11819, N4532, N4683);
nor NOR2 (N11840, N11836, N4434);
not NOT1 (N11841, N11837);
buf BUF1 (N11842, N11839);
nor NOR4 (N11843, N11840, N4100, N6318, N4564);
not NOT1 (N11844, N11835);
xor XOR2 (N11845, N11844, N5442);
and AND4 (N11846, N11800, N4940, N7935, N821);
nand NAND4 (N11847, N11822, N7463, N2741, N2130);
nand NAND2 (N11848, N11846, N6092);
nand NAND4 (N11849, N11841, N4104, N8038, N9819);
nand NAND3 (N11850, N11838, N3462, N9315);
nand NAND3 (N11851, N11848, N7152, N8033);
xor XOR2 (N11852, N11851, N5088);
xor XOR2 (N11853, N11850, N11515);
and AND4 (N11854, N11842, N11454, N5669, N5965);
xor XOR2 (N11855, N11847, N5089);
or OR2 (N11856, N11854, N11674);
buf BUF1 (N11857, N11827);
and AND4 (N11858, N11857, N2056, N5519, N3630);
not NOT1 (N11859, N11858);
nand NAND4 (N11860, N11853, N11626, N9249, N6732);
nand NAND3 (N11861, N11859, N436, N59);
or OR3 (N11862, N11852, N6262, N2835);
and AND4 (N11863, N11831, N2580, N7557, N9816);
nand NAND3 (N11864, N11860, N9710, N7803);
nor NOR3 (N11865, N11845, N11070, N2788);
and AND4 (N11866, N11834, N3650, N6532, N11157);
nor NOR3 (N11867, N11862, N8858, N104);
and AND2 (N11868, N11866, N8738);
and AND2 (N11869, N11867, N10769);
or OR2 (N11870, N11869, N4482);
not NOT1 (N11871, N11855);
not NOT1 (N11872, N11870);
buf BUF1 (N11873, N11872);
buf BUF1 (N11874, N11871);
xor XOR2 (N11875, N11856, N824);
buf BUF1 (N11876, N11873);
nand NAND2 (N11877, N11868, N8688);
nand NAND2 (N11878, N11865, N4172);
nand NAND3 (N11879, N11863, N7580, N6973);
not NOT1 (N11880, N11877);
xor XOR2 (N11881, N11843, N7918);
nor NOR4 (N11882, N11881, N3881, N3618, N3139);
not NOT1 (N11883, N11879);
nor NOR4 (N11884, N11864, N4766, N7399, N5408);
or OR3 (N11885, N11883, N5434, N6212);
buf BUF1 (N11886, N11882);
xor XOR2 (N11887, N11874, N7296);
xor XOR2 (N11888, N11876, N3087);
xor XOR2 (N11889, N11888, N6716);
xor XOR2 (N11890, N11884, N3626);
and AND3 (N11891, N11880, N8196, N3237);
not NOT1 (N11892, N11889);
not NOT1 (N11893, N11878);
nor NOR2 (N11894, N11887, N2751);
nand NAND3 (N11895, N11893, N118, N6803);
nor NOR4 (N11896, N11891, N1578, N11671, N10426);
nand NAND2 (N11897, N11894, N1436);
or OR4 (N11898, N11885, N11855, N7766, N6825);
nor NOR4 (N11899, N11849, N10913, N3946, N9228);
buf BUF1 (N11900, N11892);
nor NOR4 (N11901, N11861, N4508, N806, N3582);
or OR4 (N11902, N11890, N6081, N4117, N2989);
nor NOR2 (N11903, N11896, N7892);
and AND2 (N11904, N11900, N9557);
not NOT1 (N11905, N11903);
or OR4 (N11906, N11897, N5860, N6975, N11639);
and AND2 (N11907, N11901, N7873);
not NOT1 (N11908, N11875);
not NOT1 (N11909, N11886);
nor NOR3 (N11910, N11907, N5407, N10291);
not NOT1 (N11911, N11905);
xor XOR2 (N11912, N11899, N8276);
nor NOR4 (N11913, N11895, N3668, N9681, N736);
xor XOR2 (N11914, N11912, N10891);
or OR3 (N11915, N11902, N7343, N9367);
nor NOR3 (N11916, N11909, N3405, N11644);
buf BUF1 (N11917, N11910);
and AND2 (N11918, N11917, N1819);
xor XOR2 (N11919, N11911, N10036);
and AND4 (N11920, N11906, N2636, N3671, N10795);
nor NOR2 (N11921, N11918, N2694);
xor XOR2 (N11922, N11898, N5458);
nand NAND2 (N11923, N11914, N7793);
and AND4 (N11924, N11920, N4783, N6917, N1413);
and AND2 (N11925, N11913, N4579);
not NOT1 (N11926, N11904);
xor XOR2 (N11927, N11919, N10775);
buf BUF1 (N11928, N11908);
nor NOR3 (N11929, N11925, N8463, N4652);
nand NAND2 (N11930, N11929, N1864);
not NOT1 (N11931, N11921);
xor XOR2 (N11932, N11915, N1518);
and AND2 (N11933, N11923, N9810);
and AND2 (N11934, N11916, N3606);
nor NOR2 (N11935, N11924, N10666);
and AND2 (N11936, N11922, N5961);
nand NAND2 (N11937, N11930, N4616);
nor NOR3 (N11938, N11934, N7681, N5134);
xor XOR2 (N11939, N11933, N11151);
and AND2 (N11940, N11939, N6935);
and AND2 (N11941, N11928, N10515);
nor NOR4 (N11942, N11932, N11724, N6757, N5686);
not NOT1 (N11943, N11942);
or OR4 (N11944, N11927, N6940, N1464, N3012);
and AND3 (N11945, N11941, N6227, N4100);
xor XOR2 (N11946, N11940, N9573);
buf BUF1 (N11947, N11926);
nand NAND2 (N11948, N11945, N6501);
xor XOR2 (N11949, N11947, N335);
and AND3 (N11950, N11944, N6135, N7330);
nand NAND4 (N11951, N11949, N1646, N10644, N5910);
nand NAND3 (N11952, N11950, N1860, N5447);
nand NAND3 (N11953, N11931, N4701, N11116);
or OR4 (N11954, N11951, N4121, N1777, N5138);
nor NOR3 (N11955, N11954, N2473, N4017);
and AND4 (N11956, N11938, N6865, N10990, N9373);
and AND3 (N11957, N11946, N9785, N544);
nor NOR4 (N11958, N11955, N717, N4105, N7729);
or OR2 (N11959, N11937, N9528);
and AND4 (N11960, N11958, N3525, N8711, N5296);
xor XOR2 (N11961, N11948, N310);
nor NOR2 (N11962, N11952, N6951);
not NOT1 (N11963, N11960);
xor XOR2 (N11964, N11936, N7561);
xor XOR2 (N11965, N11959, N4052);
nand NAND3 (N11966, N11961, N11951, N10393);
not NOT1 (N11967, N11963);
or OR4 (N11968, N11956, N9422, N5312, N9069);
nor NOR2 (N11969, N11953, N3155);
and AND2 (N11970, N11957, N11231);
buf BUF1 (N11971, N11962);
nor NOR2 (N11972, N11935, N1741);
or OR4 (N11973, N11971, N3736, N9627, N1579);
nand NAND3 (N11974, N11968, N11271, N455);
xor XOR2 (N11975, N11969, N1231);
nor NOR2 (N11976, N11975, N8796);
and AND4 (N11977, N11964, N6669, N933, N11886);
nor NOR2 (N11978, N11972, N4647);
not NOT1 (N11979, N11976);
xor XOR2 (N11980, N11970, N9349);
nand NAND2 (N11981, N11977, N3258);
buf BUF1 (N11982, N11965);
nand NAND3 (N11983, N11967, N5955, N8693);
not NOT1 (N11984, N11973);
or OR4 (N11985, N11983, N10546, N2631, N5923);
not NOT1 (N11986, N11985);
or OR2 (N11987, N11980, N9862);
and AND2 (N11988, N11984, N11952);
buf BUF1 (N11989, N11987);
nand NAND3 (N11990, N11974, N3501, N8495);
xor XOR2 (N11991, N11981, N242);
xor XOR2 (N11992, N11966, N10318);
xor XOR2 (N11993, N11982, N4658);
and AND3 (N11994, N11988, N11680, N6318);
buf BUF1 (N11995, N11986);
not NOT1 (N11996, N11994);
nor NOR3 (N11997, N11943, N10154, N9419);
nand NAND2 (N11998, N11995, N6116);
xor XOR2 (N11999, N11990, N9768);
not NOT1 (N12000, N11993);
xor XOR2 (N12001, N11989, N929);
and AND3 (N12002, N11997, N9870, N9479);
xor XOR2 (N12003, N12002, N3345);
and AND2 (N12004, N12001, N2500);
not NOT1 (N12005, N11979);
not NOT1 (N12006, N11999);
nand NAND3 (N12007, N12006, N11891, N5682);
xor XOR2 (N12008, N12004, N5295);
buf BUF1 (N12009, N11992);
xor XOR2 (N12010, N12003, N1301);
nor NOR2 (N12011, N12000, N11846);
not NOT1 (N12012, N12007);
and AND4 (N12013, N12012, N7573, N7483, N8369);
or OR2 (N12014, N12005, N4250);
buf BUF1 (N12015, N12008);
nand NAND3 (N12016, N12011, N7482, N371);
buf BUF1 (N12017, N12014);
or OR2 (N12018, N12013, N6159);
or OR2 (N12019, N11978, N3238);
or OR3 (N12020, N11991, N11888, N1114);
nand NAND2 (N12021, N12009, N5944);
or OR3 (N12022, N12017, N3644, N7691);
or OR2 (N12023, N12016, N9232);
buf BUF1 (N12024, N12021);
xor XOR2 (N12025, N12018, N657);
or OR2 (N12026, N12010, N10066);
not NOT1 (N12027, N12015);
or OR4 (N12028, N12020, N11363, N8844, N3016);
not NOT1 (N12029, N12028);
buf BUF1 (N12030, N12019);
xor XOR2 (N12031, N11998, N10706);
or OR4 (N12032, N11996, N10143, N11819, N9330);
nand NAND2 (N12033, N12022, N10827);
not NOT1 (N12034, N12027);
nor NOR2 (N12035, N12030, N1578);
nor NOR3 (N12036, N12032, N4269, N11809);
or OR2 (N12037, N12031, N4989);
xor XOR2 (N12038, N12025, N2370);
nand NAND2 (N12039, N12029, N10335);
xor XOR2 (N12040, N12039, N9374);
or OR2 (N12041, N12023, N10142);
nor NOR3 (N12042, N12033, N2711, N7727);
or OR2 (N12043, N12038, N116);
or OR2 (N12044, N12040, N398);
xor XOR2 (N12045, N12037, N5909);
nand NAND3 (N12046, N12024, N7250, N1659);
and AND3 (N12047, N12041, N2000, N7088);
nand NAND4 (N12048, N12034, N8001, N6545, N11818);
nor NOR3 (N12049, N12043, N10062, N2185);
buf BUF1 (N12050, N12047);
not NOT1 (N12051, N12046);
xor XOR2 (N12052, N12026, N7295);
nand NAND4 (N12053, N12035, N1487, N1739, N9180);
xor XOR2 (N12054, N12048, N4566);
nand NAND2 (N12055, N12045, N1159);
not NOT1 (N12056, N12050);
not NOT1 (N12057, N12055);
or OR3 (N12058, N12057, N11331, N5128);
or OR4 (N12059, N12054, N1025, N8898, N11238);
xor XOR2 (N12060, N12051, N10871);
nand NAND4 (N12061, N12044, N1260, N3904, N7997);
or OR3 (N12062, N12061, N792, N6469);
nor NOR3 (N12063, N12052, N7972, N3898);
nor NOR2 (N12064, N12062, N3336);
and AND2 (N12065, N12058, N11037);
buf BUF1 (N12066, N12059);
nand NAND2 (N12067, N12049, N1306);
or OR4 (N12068, N12036, N6123, N11990, N5798);
nand NAND4 (N12069, N12065, N9699, N8399, N7179);
buf BUF1 (N12070, N12066);
nand NAND2 (N12071, N12056, N8385);
nand NAND4 (N12072, N12071, N11525, N2230, N5778);
buf BUF1 (N12073, N12060);
nand NAND2 (N12074, N12067, N11949);
not NOT1 (N12075, N12070);
xor XOR2 (N12076, N12072, N1082);
buf BUF1 (N12077, N12074);
nand NAND4 (N12078, N12073, N3449, N3889, N3639);
nor NOR4 (N12079, N12078, N10019, N6000, N7499);
and AND3 (N12080, N12075, N11472, N1385);
nor NOR2 (N12081, N12079, N9276);
or OR3 (N12082, N12064, N7149, N10515);
nor NOR2 (N12083, N12076, N10600);
nand NAND4 (N12084, N12083, N11834, N11746, N5455);
xor XOR2 (N12085, N12077, N9170);
or OR2 (N12086, N12063, N1383);
and AND3 (N12087, N12085, N2454, N7669);
nor NOR2 (N12088, N12068, N894);
xor XOR2 (N12089, N12087, N2077);
and AND4 (N12090, N12080, N3856, N70, N11890);
nor NOR3 (N12091, N12053, N9656, N9188);
or OR2 (N12092, N12091, N3360);
and AND4 (N12093, N12082, N11005, N6994, N11029);
and AND2 (N12094, N12042, N2166);
not NOT1 (N12095, N12094);
buf BUF1 (N12096, N12069);
and AND4 (N12097, N12095, N8534, N4678, N495);
not NOT1 (N12098, N12089);
nor NOR3 (N12099, N12081, N8028, N5818);
nor NOR4 (N12100, N12092, N11434, N5548, N8181);
and AND2 (N12101, N12090, N6713);
xor XOR2 (N12102, N12088, N389);
not NOT1 (N12103, N12101);
or OR4 (N12104, N12093, N2387, N2222, N8307);
nand NAND4 (N12105, N12104, N9305, N4245, N11607);
xor XOR2 (N12106, N12105, N8813);
xor XOR2 (N12107, N12086, N2020);
not NOT1 (N12108, N12096);
nor NOR4 (N12109, N12084, N3195, N1385, N8473);
or OR2 (N12110, N12106, N1616);
xor XOR2 (N12111, N12107, N1454);
nand NAND3 (N12112, N12098, N10748, N8344);
not NOT1 (N12113, N12102);
nand NAND4 (N12114, N12109, N5163, N3427, N5452);
not NOT1 (N12115, N12113);
or OR3 (N12116, N12108, N3470, N4085);
and AND4 (N12117, N12097, N9912, N10369, N4826);
nor NOR2 (N12118, N12110, N5747);
or OR4 (N12119, N12112, N9746, N8363, N9127);
nor NOR4 (N12120, N12100, N368, N7066, N6968);
not NOT1 (N12121, N12103);
and AND2 (N12122, N12120, N1391);
xor XOR2 (N12123, N12114, N1441);
nor NOR3 (N12124, N12117, N9000, N7300);
nor NOR3 (N12125, N12116, N8776, N5211);
not NOT1 (N12126, N12115);
or OR2 (N12127, N12123, N8001);
or OR3 (N12128, N12111, N5955, N11941);
nand NAND4 (N12129, N12119, N6898, N10797, N9248);
xor XOR2 (N12130, N12125, N6101);
nor NOR3 (N12131, N12099, N11732, N6010);
and AND3 (N12132, N12129, N6632, N6411);
buf BUF1 (N12133, N12124);
not NOT1 (N12134, N12118);
nor NOR4 (N12135, N12134, N10169, N1956, N515);
nand NAND4 (N12136, N12135, N2950, N3571, N11442);
or OR4 (N12137, N12127, N11739, N11741, N4507);
xor XOR2 (N12138, N12133, N6185);
xor XOR2 (N12139, N12138, N4528);
not NOT1 (N12140, N12122);
and AND4 (N12141, N12137, N2575, N4293, N637);
xor XOR2 (N12142, N12131, N6039);
xor XOR2 (N12143, N12141, N2543);
buf BUF1 (N12144, N12142);
nand NAND2 (N12145, N12128, N11481);
nor NOR2 (N12146, N12130, N9153);
nand NAND2 (N12147, N12121, N459);
nor NOR3 (N12148, N12140, N4083, N9363);
buf BUF1 (N12149, N12132);
not NOT1 (N12150, N12149);
and AND2 (N12151, N12126, N3595);
not NOT1 (N12152, N12143);
buf BUF1 (N12153, N12136);
nor NOR2 (N12154, N12144, N4547);
nand NAND4 (N12155, N12152, N3604, N2324, N408);
xor XOR2 (N12156, N12148, N5265);
or OR4 (N12157, N12156, N3729, N4165, N10184);
xor XOR2 (N12158, N12139, N187);
or OR3 (N12159, N12158, N11016, N8508);
nor NOR2 (N12160, N12153, N1243);
buf BUF1 (N12161, N12159);
xor XOR2 (N12162, N12147, N8678);
nor NOR3 (N12163, N12154, N11084, N7539);
nor NOR3 (N12164, N12161, N10587, N6250);
xor XOR2 (N12165, N12151, N6794);
xor XOR2 (N12166, N12163, N87);
buf BUF1 (N12167, N12145);
buf BUF1 (N12168, N12157);
xor XOR2 (N12169, N12150, N3199);
nand NAND3 (N12170, N12166, N2929, N6);
nand NAND3 (N12171, N12169, N8109, N283);
not NOT1 (N12172, N12170);
not NOT1 (N12173, N12160);
not NOT1 (N12174, N12162);
nand NAND4 (N12175, N12171, N4767, N3754, N6106);
buf BUF1 (N12176, N12165);
not NOT1 (N12177, N12173);
xor XOR2 (N12178, N12176, N165);
nor NOR3 (N12179, N12164, N5263, N6261);
xor XOR2 (N12180, N12167, N2027);
not NOT1 (N12181, N12180);
nor NOR3 (N12182, N12172, N9696, N12089);
or OR4 (N12183, N12168, N9438, N7409, N2989);
or OR3 (N12184, N12174, N5307, N6152);
nand NAND4 (N12185, N12179, N10677, N1615, N2821);
xor XOR2 (N12186, N12181, N7847);
or OR3 (N12187, N12186, N10401, N1309);
nand NAND4 (N12188, N12182, N11206, N5027, N5674);
or OR4 (N12189, N12178, N6246, N6447, N1036);
or OR4 (N12190, N12189, N9544, N3833, N1488);
nor NOR4 (N12191, N12146, N5670, N2640, N6036);
and AND2 (N12192, N12187, N10472);
and AND2 (N12193, N12177, N241);
or OR2 (N12194, N12188, N6641);
and AND3 (N12195, N12194, N1674, N805);
and AND3 (N12196, N12155, N8931, N9909);
nor NOR3 (N12197, N12190, N8147, N881);
not NOT1 (N12198, N12185);
or OR2 (N12199, N12191, N7203);
nand NAND4 (N12200, N12192, N1607, N9616, N2832);
buf BUF1 (N12201, N12198);
buf BUF1 (N12202, N12175);
xor XOR2 (N12203, N12193, N11021);
and AND2 (N12204, N12199, N11110);
nor NOR2 (N12205, N12204, N4999);
or OR2 (N12206, N12184, N11996);
or OR4 (N12207, N12205, N1529, N7993, N5707);
nand NAND4 (N12208, N12207, N7860, N303, N1744);
or OR2 (N12209, N12201, N8587);
not NOT1 (N12210, N12203);
nand NAND2 (N12211, N12195, N7773);
nand NAND4 (N12212, N12183, N9024, N10733, N7230);
not NOT1 (N12213, N12206);
buf BUF1 (N12214, N12200);
and AND3 (N12215, N12208, N2896, N12050);
and AND4 (N12216, N12215, N7738, N10018, N5732);
xor XOR2 (N12217, N12202, N5995);
nand NAND2 (N12218, N12213, N9536);
nand NAND2 (N12219, N12210, N10410);
xor XOR2 (N12220, N12196, N9259);
or OR4 (N12221, N12209, N6824, N5747, N5980);
or OR4 (N12222, N12216, N6328, N10242, N4442);
nand NAND3 (N12223, N12211, N9385, N12217);
nor NOR4 (N12224, N1254, N6848, N4727, N25);
and AND2 (N12225, N12224, N1780);
or OR4 (N12226, N12219, N4070, N3427, N4907);
xor XOR2 (N12227, N12226, N6450);
or OR4 (N12228, N12220, N9864, N7190, N7961);
and AND4 (N12229, N12227, N9667, N921, N8998);
not NOT1 (N12230, N12214);
xor XOR2 (N12231, N12221, N2805);
buf BUF1 (N12232, N12229);
nor NOR3 (N12233, N12223, N2068, N8500);
not NOT1 (N12234, N12212);
nand NAND4 (N12235, N12230, N3543, N7239, N6520);
not NOT1 (N12236, N12228);
or OR3 (N12237, N12218, N1237, N11829);
nor NOR2 (N12238, N12222, N2235);
or OR2 (N12239, N12237, N5296);
nand NAND2 (N12240, N12233, N7746);
xor XOR2 (N12241, N12238, N1721);
and AND3 (N12242, N12241, N10098, N3307);
buf BUF1 (N12243, N12235);
xor XOR2 (N12244, N12232, N7839);
not NOT1 (N12245, N12244);
nor NOR3 (N12246, N12240, N9029, N1686);
not NOT1 (N12247, N12242);
and AND4 (N12248, N12197, N4212, N4265, N1701);
buf BUF1 (N12249, N12236);
and AND4 (N12250, N12246, N7025, N9216, N6022);
buf BUF1 (N12251, N12248);
xor XOR2 (N12252, N12251, N1287);
or OR3 (N12253, N12245, N2756, N4877);
xor XOR2 (N12254, N12243, N7958);
or OR3 (N12255, N12249, N10184, N4230);
nor NOR3 (N12256, N12252, N2941, N3217);
or OR3 (N12257, N12234, N6190, N779);
xor XOR2 (N12258, N12254, N10512);
xor XOR2 (N12259, N12258, N10761);
or OR3 (N12260, N12250, N6329, N2055);
nand NAND3 (N12261, N12225, N8936, N2351);
xor XOR2 (N12262, N12247, N2360);
not NOT1 (N12263, N12262);
nor NOR4 (N12264, N12239, N7621, N4434, N5170);
or OR3 (N12265, N12264, N10336, N11267);
nand NAND4 (N12266, N12261, N1007, N10289, N5404);
not NOT1 (N12267, N12257);
and AND4 (N12268, N12260, N12092, N10033, N672);
not NOT1 (N12269, N12266);
xor XOR2 (N12270, N12256, N2486);
and AND4 (N12271, N12263, N8887, N8994, N4589);
nand NAND4 (N12272, N12269, N1334, N8606, N8565);
buf BUF1 (N12273, N12270);
or OR4 (N12274, N12273, N5091, N3069, N2944);
and AND3 (N12275, N12274, N10924, N7219);
nor NOR3 (N12276, N12272, N1391, N11866);
or OR3 (N12277, N12253, N3941, N3618);
and AND3 (N12278, N12275, N6682, N2908);
nor NOR4 (N12279, N12271, N10083, N10970, N10181);
buf BUF1 (N12280, N12265);
not NOT1 (N12281, N12278);
or OR2 (N12282, N12231, N9887);
nand NAND4 (N12283, N12281, N3973, N8792, N3211);
xor XOR2 (N12284, N12279, N4795);
or OR3 (N12285, N12267, N10878, N112);
or OR3 (N12286, N12280, N7839, N11588);
nor NOR2 (N12287, N12259, N6272);
not NOT1 (N12288, N12283);
xor XOR2 (N12289, N12277, N5401);
not NOT1 (N12290, N12286);
nor NOR4 (N12291, N12285, N3805, N546, N8130);
buf BUF1 (N12292, N12288);
nand NAND2 (N12293, N12284, N11175);
xor XOR2 (N12294, N12276, N9337);
xor XOR2 (N12295, N12294, N5598);
nor NOR4 (N12296, N12289, N11345, N4778, N12087);
nor NOR2 (N12297, N12268, N6575);
nor NOR4 (N12298, N12282, N8005, N7450, N9987);
not NOT1 (N12299, N12297);
nand NAND3 (N12300, N12291, N6962, N9124);
xor XOR2 (N12301, N12298, N2608);
and AND2 (N12302, N12296, N5130);
nor NOR3 (N12303, N12299, N4820, N3747);
buf BUF1 (N12304, N12302);
nor NOR4 (N12305, N12303, N10683, N4681, N4999);
or OR2 (N12306, N12305, N4978);
or OR2 (N12307, N12287, N254);
buf BUF1 (N12308, N12292);
xor XOR2 (N12309, N12304, N4033);
nand NAND4 (N12310, N12255, N6126, N12304, N8190);
and AND4 (N12311, N12295, N4904, N4670, N11568);
nand NAND3 (N12312, N12308, N45, N5076);
xor XOR2 (N12313, N12300, N604);
or OR2 (N12314, N12310, N5952);
xor XOR2 (N12315, N12290, N1008);
or OR3 (N12316, N12312, N10548, N1694);
xor XOR2 (N12317, N12314, N10690);
buf BUF1 (N12318, N12293);
buf BUF1 (N12319, N12309);
or OR2 (N12320, N12318, N9219);
nor NOR3 (N12321, N12313, N1063, N12142);
xor XOR2 (N12322, N12307, N11839);
not NOT1 (N12323, N12317);
nor NOR4 (N12324, N12306, N4542, N9880, N8416);
buf BUF1 (N12325, N12319);
and AND3 (N12326, N12324, N5488, N5637);
buf BUF1 (N12327, N12322);
nand NAND2 (N12328, N12301, N3716);
nor NOR3 (N12329, N12323, N7807, N3352);
xor XOR2 (N12330, N12315, N9713);
not NOT1 (N12331, N12326);
or OR4 (N12332, N12325, N7534, N1698, N8124);
xor XOR2 (N12333, N12330, N11152);
buf BUF1 (N12334, N12331);
xor XOR2 (N12335, N12320, N3623);
nand NAND3 (N12336, N12327, N8530, N9662);
and AND3 (N12337, N12336, N10694, N7559);
or OR2 (N12338, N12316, N6775);
or OR3 (N12339, N12321, N7750, N10594);
nor NOR2 (N12340, N12328, N10611);
xor XOR2 (N12341, N12340, N2935);
nor NOR3 (N12342, N12334, N9170, N7574);
not NOT1 (N12343, N12337);
xor XOR2 (N12344, N12343, N6461);
xor XOR2 (N12345, N12342, N3675);
not NOT1 (N12346, N12311);
nand NAND4 (N12347, N12333, N2166, N5324, N10220);
or OR2 (N12348, N12339, N9658);
xor XOR2 (N12349, N12335, N7949);
and AND3 (N12350, N12346, N8947, N11434);
nor NOR3 (N12351, N12348, N1903, N7860);
nor NOR2 (N12352, N12332, N10400);
buf BUF1 (N12353, N12352);
buf BUF1 (N12354, N12345);
xor XOR2 (N12355, N12344, N11201);
and AND2 (N12356, N12347, N425);
not NOT1 (N12357, N12338);
buf BUF1 (N12358, N12349);
not NOT1 (N12359, N12354);
and AND4 (N12360, N12350, N11884, N1372, N6125);
nand NAND4 (N12361, N12360, N4092, N1808, N2297);
and AND4 (N12362, N12351, N1622, N8961, N4524);
and AND4 (N12363, N12358, N3874, N2282, N12216);
buf BUF1 (N12364, N12356);
not NOT1 (N12365, N12353);
or OR4 (N12366, N12364, N4769, N9736, N12089);
or OR3 (N12367, N12359, N6022, N8299);
xor XOR2 (N12368, N12363, N10032);
xor XOR2 (N12369, N12368, N11725);
xor XOR2 (N12370, N12361, N2485);
nand NAND3 (N12371, N12370, N2437, N5375);
nor NOR2 (N12372, N12367, N11953);
buf BUF1 (N12373, N12362);
and AND4 (N12374, N12357, N6530, N10281, N5851);
nor NOR3 (N12375, N12355, N7340, N11281);
or OR2 (N12376, N12371, N2961);
xor XOR2 (N12377, N12366, N8076);
and AND4 (N12378, N12341, N8240, N8679, N9467);
not NOT1 (N12379, N12373);
nor NOR3 (N12380, N12369, N2777, N3043);
not NOT1 (N12381, N12329);
buf BUF1 (N12382, N12374);
buf BUF1 (N12383, N12378);
buf BUF1 (N12384, N12380);
not NOT1 (N12385, N12379);
buf BUF1 (N12386, N12376);
buf BUF1 (N12387, N12386);
xor XOR2 (N12388, N12387, N2449);
not NOT1 (N12389, N12381);
or OR2 (N12390, N12382, N8110);
nor NOR4 (N12391, N12375, N3760, N5117, N2536);
or OR3 (N12392, N12383, N5105, N3143);
buf BUF1 (N12393, N12389);
nand NAND2 (N12394, N12391, N3282);
nand NAND2 (N12395, N12384, N6190);
xor XOR2 (N12396, N12395, N7702);
nand NAND4 (N12397, N12396, N12346, N2799, N3499);
not NOT1 (N12398, N12388);
buf BUF1 (N12399, N12372);
not NOT1 (N12400, N12385);
xor XOR2 (N12401, N12400, N6744);
or OR4 (N12402, N12398, N3491, N5662, N12056);
nand NAND2 (N12403, N12397, N8405);
xor XOR2 (N12404, N12365, N5214);
nand NAND3 (N12405, N12401, N5560, N5724);
or OR3 (N12406, N12403, N5349, N12326);
and AND3 (N12407, N12377, N7050, N9176);
buf BUF1 (N12408, N12393);
nor NOR4 (N12409, N12399, N7621, N5743, N3618);
or OR2 (N12410, N12392, N7856);
nand NAND4 (N12411, N12390, N7948, N9040, N1977);
nand NAND4 (N12412, N12407, N12396, N10570, N4339);
not NOT1 (N12413, N12406);
not NOT1 (N12414, N12413);
or OR2 (N12415, N12411, N7134);
nor NOR2 (N12416, N12410, N109);
buf BUF1 (N12417, N12415);
not NOT1 (N12418, N12408);
nor NOR4 (N12419, N12402, N6682, N9035, N10682);
or OR4 (N12420, N12419, N4308, N4583, N10795);
buf BUF1 (N12421, N12418);
buf BUF1 (N12422, N12404);
nand NAND4 (N12423, N12414, N6842, N7738, N4878);
xor XOR2 (N12424, N12423, N11585);
not NOT1 (N12425, N12394);
and AND3 (N12426, N12420, N2409, N4805);
not NOT1 (N12427, N12409);
not NOT1 (N12428, N12421);
nand NAND3 (N12429, N12412, N6674, N6351);
and AND2 (N12430, N12427, N7698);
not NOT1 (N12431, N12425);
buf BUF1 (N12432, N12417);
xor XOR2 (N12433, N12432, N4512);
xor XOR2 (N12434, N12426, N4742);
nand NAND2 (N12435, N12416, N6006);
not NOT1 (N12436, N12430);
or OR3 (N12437, N12435, N1755, N1402);
nor NOR3 (N12438, N12428, N10332, N5479);
nor NOR2 (N12439, N12422, N1449);
or OR4 (N12440, N12424, N8920, N8765, N23);
nor NOR4 (N12441, N12405, N8507, N6968, N10807);
nand NAND4 (N12442, N12441, N11021, N10320, N849);
or OR2 (N12443, N12433, N9335);
nor NOR3 (N12444, N12442, N10512, N1235);
buf BUF1 (N12445, N12438);
buf BUF1 (N12446, N12440);
nor NOR3 (N12447, N12437, N9121, N10569);
xor XOR2 (N12448, N12439, N6049);
nor NOR3 (N12449, N12436, N1520, N419);
or OR4 (N12450, N12448, N4558, N9159, N5249);
or OR4 (N12451, N12449, N11670, N7366, N7423);
or OR4 (N12452, N12434, N5549, N7955, N11424);
or OR4 (N12453, N12452, N5119, N7752, N9650);
nor NOR3 (N12454, N12444, N4463, N3837);
nor NOR2 (N12455, N12450, N11482);
buf BUF1 (N12456, N12446);
nor NOR3 (N12457, N12454, N10788, N3308);
nor NOR2 (N12458, N12457, N8821);
and AND4 (N12459, N12451, N8852, N6385, N8178);
not NOT1 (N12460, N12455);
and AND3 (N12461, N12458, N1563, N320);
nor NOR4 (N12462, N12443, N2345, N8564, N11410);
not NOT1 (N12463, N12429);
xor XOR2 (N12464, N12463, N7517);
or OR3 (N12465, N12462, N5375, N7966);
or OR4 (N12466, N12460, N11819, N227, N12133);
xor XOR2 (N12467, N12465, N704);
nand NAND4 (N12468, N12461, N12175, N6704, N2304);
and AND4 (N12469, N12447, N6651, N1201, N2575);
xor XOR2 (N12470, N12469, N23);
nand NAND4 (N12471, N12431, N4554, N3856, N1921);
or OR2 (N12472, N12445, N8718);
nand NAND3 (N12473, N12459, N12311, N11260);
not NOT1 (N12474, N12467);
xor XOR2 (N12475, N12453, N2893);
nand NAND4 (N12476, N12468, N523, N1467, N9159);
nand NAND2 (N12477, N12470, N9985);
or OR3 (N12478, N12474, N11172, N6635);
xor XOR2 (N12479, N12475, N953);
buf BUF1 (N12480, N12479);
buf BUF1 (N12481, N12480);
or OR3 (N12482, N12471, N8599, N4521);
xor XOR2 (N12483, N12481, N1425);
nor NOR2 (N12484, N12477, N9107);
xor XOR2 (N12485, N12472, N10404);
and AND2 (N12486, N12466, N10791);
buf BUF1 (N12487, N12485);
nand NAND3 (N12488, N12464, N853, N5420);
nor NOR3 (N12489, N12486, N1740, N10099);
not NOT1 (N12490, N12489);
and AND2 (N12491, N12484, N7593);
xor XOR2 (N12492, N12491, N5368);
not NOT1 (N12493, N12488);
and AND4 (N12494, N12476, N10278, N9381, N11243);
and AND4 (N12495, N12483, N2924, N810, N9761);
buf BUF1 (N12496, N12478);
buf BUF1 (N12497, N12487);
nand NAND3 (N12498, N12492, N2299, N2078);
not NOT1 (N12499, N12497);
and AND4 (N12500, N12456, N4218, N736, N7283);
or OR2 (N12501, N12500, N7929);
and AND4 (N12502, N12501, N5326, N9945, N3014);
nand NAND2 (N12503, N12490, N4061);
not NOT1 (N12504, N12496);
buf BUF1 (N12505, N12498);
nor NOR2 (N12506, N12473, N3361);
xor XOR2 (N12507, N12505, N3117);
buf BUF1 (N12508, N12504);
and AND3 (N12509, N12499, N3655, N3564);
buf BUF1 (N12510, N12509);
nand NAND4 (N12511, N12510, N10895, N12078, N1129);
xor XOR2 (N12512, N12503, N11916);
or OR4 (N12513, N12495, N4073, N7469, N4857);
and AND3 (N12514, N12507, N1841, N10025);
or OR2 (N12515, N12513, N10400);
buf BUF1 (N12516, N12512);
and AND3 (N12517, N12514, N9392, N433);
nand NAND3 (N12518, N12517, N11799, N5429);
nor NOR3 (N12519, N12502, N3036, N163);
not NOT1 (N12520, N12508);
or OR2 (N12521, N12515, N11636);
nand NAND2 (N12522, N12521, N5550);
nor NOR4 (N12523, N12511, N10400, N1319, N4637);
xor XOR2 (N12524, N12482, N5206);
not NOT1 (N12525, N12520);
and AND4 (N12526, N12522, N5817, N12353, N899);
buf BUF1 (N12527, N12525);
buf BUF1 (N12528, N12518);
or OR3 (N12529, N12516, N10182, N460);
nand NAND3 (N12530, N12506, N1, N3971);
buf BUF1 (N12531, N12519);
nand NAND2 (N12532, N12493, N10992);
not NOT1 (N12533, N12523);
xor XOR2 (N12534, N12527, N10223);
buf BUF1 (N12535, N12526);
or OR4 (N12536, N12532, N1673, N10965, N2933);
nand NAND2 (N12537, N12494, N3085);
buf BUF1 (N12538, N12529);
nand NAND2 (N12539, N12530, N9420);
buf BUF1 (N12540, N12537);
and AND2 (N12541, N12535, N4899);
nor NOR3 (N12542, N12524, N2106, N4864);
buf BUF1 (N12543, N12533);
nor NOR2 (N12544, N12528, N11397);
and AND2 (N12545, N12543, N11595);
not NOT1 (N12546, N12542);
nor NOR2 (N12547, N12540, N4434);
nand NAND3 (N12548, N12544, N4536, N4431);
nand NAND2 (N12549, N12541, N1811);
nand NAND2 (N12550, N12545, N6992);
nor NOR3 (N12551, N12549, N1745, N11358);
nand NAND4 (N12552, N12551, N268, N8044, N7088);
xor XOR2 (N12553, N12547, N10575);
not NOT1 (N12554, N12536);
nor NOR4 (N12555, N12534, N4977, N9170, N856);
and AND4 (N12556, N12552, N7274, N3224, N6050);
nor NOR3 (N12557, N12548, N5807, N7716);
and AND4 (N12558, N12550, N7080, N6859, N9421);
and AND4 (N12559, N12555, N6757, N2972, N10197);
and AND4 (N12560, N12546, N6271, N10955, N5652);
or OR3 (N12561, N12556, N11530, N8190);
or OR4 (N12562, N12557, N6340, N12542, N4726);
or OR2 (N12563, N12554, N10538);
buf BUF1 (N12564, N12539);
and AND3 (N12565, N12562, N9616, N10848);
nand NAND4 (N12566, N12559, N3932, N9357, N1640);
and AND4 (N12567, N12566, N8544, N1210, N2358);
not NOT1 (N12568, N12558);
not NOT1 (N12569, N12553);
or OR3 (N12570, N12563, N5881, N1095);
xor XOR2 (N12571, N12531, N12396);
xor XOR2 (N12572, N12570, N1412);
buf BUF1 (N12573, N12571);
xor XOR2 (N12574, N12538, N5561);
or OR4 (N12575, N12568, N2082, N4553, N6920);
nor NOR3 (N12576, N12565, N7750, N4146);
or OR3 (N12577, N12560, N2729, N6917);
nand NAND4 (N12578, N12577, N2720, N9500, N4962);
xor XOR2 (N12579, N12575, N2905);
nor NOR3 (N12580, N12564, N173, N6132);
xor XOR2 (N12581, N12574, N3249);
nor NOR3 (N12582, N12573, N1267, N10909);
not NOT1 (N12583, N12579);
xor XOR2 (N12584, N12581, N12184);
nand NAND2 (N12585, N12576, N251);
buf BUF1 (N12586, N12561);
and AND3 (N12587, N12569, N6702, N3807);
not NOT1 (N12588, N12584);
xor XOR2 (N12589, N12578, N6221);
not NOT1 (N12590, N12572);
or OR4 (N12591, N12567, N418, N11980, N2853);
or OR2 (N12592, N12589, N202);
nor NOR4 (N12593, N12591, N2891, N3004, N4331);
buf BUF1 (N12594, N12590);
xor XOR2 (N12595, N12580, N5074);
not NOT1 (N12596, N12593);
xor XOR2 (N12597, N12585, N165);
not NOT1 (N12598, N12592);
or OR2 (N12599, N12588, N12480);
nand NAND2 (N12600, N12596, N3858);
buf BUF1 (N12601, N12597);
or OR2 (N12602, N12587, N8139);
or OR2 (N12603, N12599, N12504);
not NOT1 (N12604, N12594);
and AND4 (N12605, N12586, N10418, N3532, N10890);
not NOT1 (N12606, N12595);
nor NOR2 (N12607, N12582, N11805);
or OR3 (N12608, N12607, N6140, N1711);
and AND4 (N12609, N12604, N427, N2803, N9442);
or OR3 (N12610, N12608, N1261, N9991);
nand NAND3 (N12611, N12610, N9434, N9348);
nor NOR2 (N12612, N12611, N12311);
or OR2 (N12613, N12601, N9970);
nor NOR2 (N12614, N12605, N4740);
nor NOR4 (N12615, N12598, N8757, N3833, N4497);
and AND4 (N12616, N12606, N7343, N607, N7071);
not NOT1 (N12617, N12612);
xor XOR2 (N12618, N12617, N11664);
and AND3 (N12619, N12613, N7029, N1230);
xor XOR2 (N12620, N12583, N941);
not NOT1 (N12621, N12618);
nor NOR3 (N12622, N12615, N4304, N6127);
buf BUF1 (N12623, N12622);
buf BUF1 (N12624, N12619);
nand NAND3 (N12625, N12603, N4520, N5638);
buf BUF1 (N12626, N12621);
or OR2 (N12627, N12609, N6874);
and AND4 (N12628, N12626, N6826, N8161, N4009);
or OR2 (N12629, N12628, N10250);
nand NAND2 (N12630, N12620, N5478);
or OR4 (N12631, N12602, N10974, N1105, N5746);
xor XOR2 (N12632, N12627, N9142);
buf BUF1 (N12633, N12616);
and AND3 (N12634, N12633, N12365, N6730);
or OR3 (N12635, N12625, N545, N11128);
xor XOR2 (N12636, N12631, N8956);
xor XOR2 (N12637, N12630, N6936);
buf BUF1 (N12638, N12634);
or OR4 (N12639, N12636, N8733, N8759, N10740);
not NOT1 (N12640, N12639);
nand NAND4 (N12641, N12637, N7019, N3401, N10212);
buf BUF1 (N12642, N12629);
buf BUF1 (N12643, N12614);
nor NOR3 (N12644, N12641, N5062, N4185);
not NOT1 (N12645, N12642);
nand NAND4 (N12646, N12640, N10465, N7291, N8145);
nand NAND4 (N12647, N12646, N5585, N6143, N6755);
buf BUF1 (N12648, N12623);
buf BUF1 (N12649, N12632);
xor XOR2 (N12650, N12638, N4349);
nor NOR2 (N12651, N12635, N9533);
or OR4 (N12652, N12647, N8533, N11617, N5515);
nor NOR2 (N12653, N12650, N6917);
not NOT1 (N12654, N12624);
buf BUF1 (N12655, N12600);
nor NOR3 (N12656, N12652, N1015, N1051);
and AND2 (N12657, N12648, N9560);
or OR4 (N12658, N12644, N7910, N4262, N2597);
nor NOR3 (N12659, N12658, N6892, N5284);
and AND2 (N12660, N12659, N5661);
nor NOR3 (N12661, N12656, N6835, N2463);
buf BUF1 (N12662, N12649);
and AND2 (N12663, N12645, N11013);
and AND3 (N12664, N12657, N2125, N5662);
not NOT1 (N12665, N12664);
not NOT1 (N12666, N12662);
or OR3 (N12667, N12643, N4528, N592);
or OR2 (N12668, N12653, N5608);
xor XOR2 (N12669, N12661, N5018);
and AND2 (N12670, N12660, N12615);
not NOT1 (N12671, N12665);
xor XOR2 (N12672, N12671, N8301);
nor NOR4 (N12673, N12672, N8925, N7880, N4316);
not NOT1 (N12674, N12655);
nor NOR2 (N12675, N12663, N9256);
or OR3 (N12676, N12674, N10172, N1934);
nor NOR4 (N12677, N12673, N4424, N10918, N9623);
not NOT1 (N12678, N12668);
or OR3 (N12679, N12670, N5181, N6760);
xor XOR2 (N12680, N12651, N6674);
nand NAND2 (N12681, N12667, N9832);
buf BUF1 (N12682, N12676);
buf BUF1 (N12683, N12682);
or OR3 (N12684, N12666, N8553, N2665);
nand NAND4 (N12685, N12684, N8154, N6438, N5237);
nor NOR2 (N12686, N12678, N7733);
nand NAND4 (N12687, N12680, N4791, N10181, N7723);
and AND4 (N12688, N12654, N852, N5694, N3840);
nor NOR4 (N12689, N12685, N2085, N6077, N7999);
and AND3 (N12690, N12681, N558, N7577);
nor NOR2 (N12691, N12677, N9718);
or OR2 (N12692, N12688, N10140);
nand NAND3 (N12693, N12687, N1922, N4556);
buf BUF1 (N12694, N12692);
and AND2 (N12695, N12690, N3931);
not NOT1 (N12696, N12694);
nor NOR4 (N12697, N12683, N544, N3491, N9674);
nor NOR3 (N12698, N12697, N146, N11372);
xor XOR2 (N12699, N12698, N10307);
or OR4 (N12700, N12675, N7859, N2703, N3863);
or OR2 (N12701, N12679, N3564);
or OR4 (N12702, N12695, N9411, N2405, N10305);
and AND3 (N12703, N12686, N2362, N19);
buf BUF1 (N12704, N12699);
nor NOR2 (N12705, N12703, N12183);
or OR3 (N12706, N12700, N7246, N9861);
nand NAND3 (N12707, N12701, N7533, N4359);
and AND3 (N12708, N12707, N11868, N6664);
not NOT1 (N12709, N12702);
xor XOR2 (N12710, N12693, N4430);
buf BUF1 (N12711, N12691);
nor NOR3 (N12712, N12696, N9960, N2454);
xor XOR2 (N12713, N12706, N6800);
and AND2 (N12714, N12669, N6605);
or OR3 (N12715, N12705, N745, N6571);
not NOT1 (N12716, N12713);
and AND2 (N12717, N12714, N4969);
or OR4 (N12718, N12712, N4621, N4333, N11316);
or OR4 (N12719, N12717, N226, N3188, N7309);
nor NOR3 (N12720, N12719, N10280, N7061);
and AND4 (N12721, N12708, N4084, N1384, N10547);
or OR4 (N12722, N12704, N11192, N2724, N12376);
nor NOR3 (N12723, N12716, N11549, N1965);
nor NOR3 (N12724, N12711, N2429, N6759);
nand NAND3 (N12725, N12721, N4909, N968);
not NOT1 (N12726, N12715);
nor NOR4 (N12727, N12709, N734, N6315, N6092);
buf BUF1 (N12728, N12710);
xor XOR2 (N12729, N12728, N10740);
xor XOR2 (N12730, N12725, N6614);
nor NOR4 (N12731, N12689, N3927, N9556, N920);
buf BUF1 (N12732, N12727);
or OR4 (N12733, N12723, N4260, N1911, N12233);
xor XOR2 (N12734, N12732, N4760);
not NOT1 (N12735, N12724);
nand NAND4 (N12736, N12718, N9598, N9330, N10585);
not NOT1 (N12737, N12726);
nor NOR2 (N12738, N12722, N12366);
nor NOR3 (N12739, N12733, N9069, N1640);
nand NAND2 (N12740, N12731, N1461);
nand NAND2 (N12741, N12729, N2279);
not NOT1 (N12742, N12720);
not NOT1 (N12743, N12738);
and AND4 (N12744, N12742, N4709, N7224, N8703);
nor NOR2 (N12745, N12735, N964);
not NOT1 (N12746, N12736);
buf BUF1 (N12747, N12746);
or OR2 (N12748, N12740, N7128);
xor XOR2 (N12749, N12741, N10698);
nand NAND4 (N12750, N12734, N8717, N11275, N6187);
nor NOR2 (N12751, N12749, N1079);
and AND3 (N12752, N12737, N10431, N8657);
xor XOR2 (N12753, N12744, N589);
not NOT1 (N12754, N12739);
buf BUF1 (N12755, N12747);
not NOT1 (N12756, N12750);
not NOT1 (N12757, N12745);
and AND4 (N12758, N12756, N17, N11356, N6480);
and AND2 (N12759, N12730, N1949);
or OR2 (N12760, N12754, N9479);
buf BUF1 (N12761, N12752);
nor NOR2 (N12762, N12757, N5649);
xor XOR2 (N12763, N12751, N3954);
xor XOR2 (N12764, N12760, N8298);
and AND3 (N12765, N12764, N8734, N7517);
xor XOR2 (N12766, N12762, N4605);
and AND3 (N12767, N12743, N10109, N8648);
and AND4 (N12768, N12763, N1427, N58, N11490);
and AND2 (N12769, N12748, N5051);
nor NOR4 (N12770, N12766, N9589, N9231, N7758);
not NOT1 (N12771, N12769);
nand NAND4 (N12772, N12765, N10799, N11026, N4363);
buf BUF1 (N12773, N12772);
and AND4 (N12774, N12755, N10846, N8927, N10251);
or OR3 (N12775, N12774, N8422, N11135);
nand NAND4 (N12776, N12771, N2368, N7815, N2904);
and AND2 (N12777, N12768, N9050);
buf BUF1 (N12778, N12759);
nand NAND4 (N12779, N12776, N9197, N6623, N7816);
not NOT1 (N12780, N12777);
nand NAND4 (N12781, N12761, N7153, N8927, N909);
nor NOR2 (N12782, N12773, N1266);
buf BUF1 (N12783, N12782);
buf BUF1 (N12784, N12758);
and AND4 (N12785, N12783, N9769, N5410, N2206);
nor NOR3 (N12786, N12753, N8952, N48);
xor XOR2 (N12787, N12770, N2043);
nand NAND3 (N12788, N12780, N2969, N7748);
buf BUF1 (N12789, N12778);
or OR4 (N12790, N12787, N9673, N9522, N10465);
nand NAND3 (N12791, N12779, N4887, N5456);
and AND3 (N12792, N12786, N2433, N12412);
nand NAND2 (N12793, N12789, N11771);
not NOT1 (N12794, N12775);
nor NOR4 (N12795, N12785, N6731, N1263, N364);
nor NOR4 (N12796, N12788, N3295, N274, N7441);
or OR3 (N12797, N12793, N8368, N5995);
buf BUF1 (N12798, N12784);
nand NAND2 (N12799, N12792, N7914);
xor XOR2 (N12800, N12781, N1267);
nor NOR4 (N12801, N12796, N5292, N11520, N5436);
nor NOR3 (N12802, N12767, N3518, N7201);
or OR2 (N12803, N12801, N12329);
nand NAND2 (N12804, N12803, N10856);
not NOT1 (N12805, N12795);
nor NOR2 (N12806, N12805, N6537);
and AND2 (N12807, N12799, N8578);
nor NOR3 (N12808, N12790, N818, N9900);
and AND4 (N12809, N12800, N10683, N901, N2740);
not NOT1 (N12810, N12804);
xor XOR2 (N12811, N12810, N5128);
nor NOR3 (N12812, N12809, N7034, N5376);
nor NOR4 (N12813, N12808, N131, N4342, N8415);
not NOT1 (N12814, N12791);
or OR4 (N12815, N12794, N7208, N5111, N6842);
not NOT1 (N12816, N12813);
nor NOR2 (N12817, N12815, N8860);
or OR4 (N12818, N12797, N11759, N5826, N2338);
nand NAND4 (N12819, N12806, N12368, N4378, N9451);
xor XOR2 (N12820, N12802, N7900);
not NOT1 (N12821, N12816);
and AND4 (N12822, N12821, N3958, N7399, N11981);
buf BUF1 (N12823, N12807);
nor NOR2 (N12824, N12819, N10589);
nand NAND2 (N12825, N12818, N11788);
not NOT1 (N12826, N12798);
or OR3 (N12827, N12822, N2795, N4326);
nand NAND4 (N12828, N12827, N1114, N6408, N2178);
and AND4 (N12829, N12825, N9908, N5005, N8375);
and AND2 (N12830, N12817, N8411);
nor NOR3 (N12831, N12828, N6776, N1260);
buf BUF1 (N12832, N12811);
and AND3 (N12833, N12829, N1191, N2280);
not NOT1 (N12834, N12824);
or OR4 (N12835, N12833, N5487, N9940, N10337);
and AND3 (N12836, N12820, N7088, N190);
buf BUF1 (N12837, N12832);
and AND4 (N12838, N12837, N6383, N313, N8161);
buf BUF1 (N12839, N12812);
buf BUF1 (N12840, N12835);
and AND2 (N12841, N12834, N3300);
or OR2 (N12842, N12839, N8143);
xor XOR2 (N12843, N12814, N12108);
xor XOR2 (N12844, N12840, N10036);
xor XOR2 (N12845, N12843, N2203);
xor XOR2 (N12846, N12845, N10860);
buf BUF1 (N12847, N12844);
and AND2 (N12848, N12826, N12148);
or OR2 (N12849, N12836, N7823);
xor XOR2 (N12850, N12831, N2607);
not NOT1 (N12851, N12830);
nor NOR3 (N12852, N12851, N8860, N7354);
buf BUF1 (N12853, N12846);
buf BUF1 (N12854, N12838);
buf BUF1 (N12855, N12849);
buf BUF1 (N12856, N12855);
buf BUF1 (N12857, N12856);
nor NOR2 (N12858, N12823, N1906);
and AND2 (N12859, N12841, N5093);
buf BUF1 (N12860, N12854);
or OR3 (N12861, N12850, N4833, N3590);
and AND2 (N12862, N12847, N4002);
buf BUF1 (N12863, N12853);
or OR3 (N12864, N12852, N12441, N6559);
and AND3 (N12865, N12863, N9918, N8159);
or OR2 (N12866, N12842, N4744);
buf BUF1 (N12867, N12857);
and AND4 (N12868, N12866, N5606, N4250, N2111);
not NOT1 (N12869, N12867);
nor NOR2 (N12870, N12869, N4402);
nor NOR3 (N12871, N12864, N1571, N4196);
xor XOR2 (N12872, N12858, N9550);
buf BUF1 (N12873, N12872);
or OR3 (N12874, N12862, N4608, N1798);
or OR4 (N12875, N12873, N11213, N5612, N10742);
buf BUF1 (N12876, N12868);
or OR4 (N12877, N12859, N10117, N10583, N8146);
not NOT1 (N12878, N12874);
nor NOR2 (N12879, N12860, N3863);
nand NAND2 (N12880, N12876, N2547);
or OR4 (N12881, N12880, N4688, N11066, N5597);
not NOT1 (N12882, N12870);
nand NAND4 (N12883, N12875, N10981, N12878, N5457);
xor XOR2 (N12884, N9759, N7169);
buf BUF1 (N12885, N12883);
or OR3 (N12886, N12882, N9159, N12863);
nand NAND2 (N12887, N12865, N6853);
and AND2 (N12888, N12871, N6053);
not NOT1 (N12889, N12888);
and AND3 (N12890, N12881, N1452, N2783);
nor NOR2 (N12891, N12877, N1302);
nand NAND4 (N12892, N12848, N9504, N3516, N11466);
nor NOR4 (N12893, N12892, N6364, N12759, N98);
buf BUF1 (N12894, N12879);
nand NAND2 (N12895, N12885, N7226);
not NOT1 (N12896, N12891);
nor NOR2 (N12897, N12861, N9972);
nor NOR4 (N12898, N12897, N80, N2205, N6225);
or OR3 (N12899, N12890, N2569, N6306);
not NOT1 (N12900, N12896);
nor NOR3 (N12901, N12898, N1508, N9607);
and AND3 (N12902, N12893, N1639, N3612);
or OR2 (N12903, N12901, N11089);
nor NOR3 (N12904, N12884, N7789, N5171);
xor XOR2 (N12905, N12899, N2786);
not NOT1 (N12906, N12902);
and AND2 (N12907, N12895, N10242);
not NOT1 (N12908, N12887);
and AND2 (N12909, N12907, N12226);
xor XOR2 (N12910, N12900, N7176);
or OR4 (N12911, N12905, N9791, N2280, N86);
xor XOR2 (N12912, N12903, N5464);
not NOT1 (N12913, N12889);
or OR2 (N12914, N12910, N4834);
nor NOR3 (N12915, N12906, N9810, N11864);
xor XOR2 (N12916, N12913, N8045);
nor NOR4 (N12917, N12894, N5223, N10006, N7716);
not NOT1 (N12918, N12909);
xor XOR2 (N12919, N12918, N8498);
nand NAND4 (N12920, N12919, N4721, N12734, N5188);
not NOT1 (N12921, N12915);
and AND4 (N12922, N12908, N10901, N9690, N11936);
nand NAND3 (N12923, N12911, N11075, N3915);
nand NAND3 (N12924, N12904, N9081, N6912);
and AND3 (N12925, N12924, N6001, N11457);
nor NOR3 (N12926, N12920, N10730, N8797);
xor XOR2 (N12927, N12912, N9192);
not NOT1 (N12928, N12921);
and AND2 (N12929, N12925, N7602);
not NOT1 (N12930, N12922);
xor XOR2 (N12931, N12928, N10248);
xor XOR2 (N12932, N12917, N5895);
or OR3 (N12933, N12916, N7084, N11403);
xor XOR2 (N12934, N12929, N5656);
or OR4 (N12935, N12923, N5661, N1695, N11173);
or OR2 (N12936, N12931, N3080);
nor NOR4 (N12937, N12930, N12328, N4297, N1850);
nand NAND3 (N12938, N12886, N5813, N6087);
or OR3 (N12939, N12933, N188, N67);
buf BUF1 (N12940, N12926);
xor XOR2 (N12941, N12927, N3846);
buf BUF1 (N12942, N12936);
nand NAND3 (N12943, N12941, N2072, N8846);
xor XOR2 (N12944, N12943, N12921);
buf BUF1 (N12945, N12937);
or OR3 (N12946, N12935, N6484, N2762);
and AND3 (N12947, N12946, N5505, N344);
not NOT1 (N12948, N12942);
and AND3 (N12949, N12940, N12908, N10715);
xor XOR2 (N12950, N12939, N2530);
nor NOR4 (N12951, N12914, N2981, N4573, N1022);
and AND4 (N12952, N12950, N656, N10026, N5944);
nand NAND2 (N12953, N12938, N5186);
nand NAND4 (N12954, N12944, N5403, N3282, N2683);
buf BUF1 (N12955, N12949);
not NOT1 (N12956, N12951);
not NOT1 (N12957, N12954);
nand NAND2 (N12958, N12957, N2478);
nor NOR3 (N12959, N12952, N921, N11325);
or OR2 (N12960, N12947, N3315);
or OR3 (N12961, N12956, N6281, N7247);
and AND3 (N12962, N12958, N10020, N12386);
and AND3 (N12963, N12945, N3231, N404);
xor XOR2 (N12964, N12962, N2706);
nor NOR4 (N12965, N12932, N934, N12079, N4577);
xor XOR2 (N12966, N12955, N6087);
nand NAND3 (N12967, N12965, N5561, N186);
buf BUF1 (N12968, N12953);
buf BUF1 (N12969, N12959);
and AND2 (N12970, N12968, N9932);
and AND2 (N12971, N12969, N1846);
buf BUF1 (N12972, N12967);
nand NAND4 (N12973, N12972, N7151, N12068, N1279);
xor XOR2 (N12974, N12971, N12718);
and AND3 (N12975, N12948, N2678, N5174);
or OR2 (N12976, N12960, N3346);
nand NAND3 (N12977, N12963, N11351, N1836);
or OR3 (N12978, N12975, N12444, N4001);
xor XOR2 (N12979, N12970, N7992);
buf BUF1 (N12980, N12977);
or OR3 (N12981, N12966, N8369, N10256);
not NOT1 (N12982, N12974);
nand NAND3 (N12983, N12982, N10279, N5623);
xor XOR2 (N12984, N12979, N11276);
and AND3 (N12985, N12934, N8660, N12718);
xor XOR2 (N12986, N12983, N1726);
not NOT1 (N12987, N12986);
buf BUF1 (N12988, N12978);
or OR2 (N12989, N12981, N16);
xor XOR2 (N12990, N12988, N2909);
buf BUF1 (N12991, N12984);
or OR4 (N12992, N12964, N5284, N2011, N3982);
xor XOR2 (N12993, N12991, N8996);
and AND3 (N12994, N12987, N1157, N9840);
and AND2 (N12995, N12993, N12012);
and AND3 (N12996, N12995, N8195, N1045);
buf BUF1 (N12997, N12961);
xor XOR2 (N12998, N12985, N1916);
nor NOR3 (N12999, N12990, N8638, N5552);
nor NOR4 (N13000, N12999, N12210, N8274, N2839);
buf BUF1 (N13001, N12996);
nand NAND2 (N13002, N12976, N4985);
not NOT1 (N13003, N12989);
xor XOR2 (N13004, N13000, N3983);
or OR3 (N13005, N12992, N11278, N804);
nand NAND3 (N13006, N13001, N9112, N11824);
nor NOR3 (N13007, N12980, N2832, N5834);
or OR2 (N13008, N13005, N4100);
and AND3 (N13009, N12994, N12048, N1191);
or OR2 (N13010, N13007, N734);
buf BUF1 (N13011, N12998);
and AND3 (N13012, N13010, N5377, N11801);
xor XOR2 (N13013, N13011, N5196);
or OR3 (N13014, N12997, N1918, N1133);
nand NAND2 (N13015, N12973, N3727);
or OR4 (N13016, N13004, N6382, N12632, N1273);
buf BUF1 (N13017, N13003);
xor XOR2 (N13018, N13009, N8634);
nand NAND3 (N13019, N13017, N4180, N7149);
nor NOR2 (N13020, N13019, N5831);
nand NAND2 (N13021, N13015, N826);
not NOT1 (N13022, N13021);
xor XOR2 (N13023, N13006, N6007);
nor NOR3 (N13024, N13016, N7848, N9963);
or OR3 (N13025, N13013, N4146, N3436);
and AND2 (N13026, N13008, N8721);
nor NOR3 (N13027, N13024, N5389, N1007);
and AND4 (N13028, N13026, N2753, N8997, N831);
and AND4 (N13029, N13023, N7325, N5141, N4988);
or OR3 (N13030, N13028, N5912, N5480);
nand NAND4 (N13031, N13022, N5684, N8642, N11586);
not NOT1 (N13032, N13018);
and AND4 (N13033, N13002, N10278, N1792, N33);
or OR3 (N13034, N13012, N6399, N3996);
not NOT1 (N13035, N13027);
and AND3 (N13036, N13014, N6090, N9345);
or OR4 (N13037, N13032, N2582, N6311, N9911);
not NOT1 (N13038, N13037);
and AND2 (N13039, N13029, N12569);
nand NAND4 (N13040, N13039, N8901, N7355, N4852);
nor NOR4 (N13041, N13036, N796, N2369, N8513);
nand NAND4 (N13042, N13034, N10240, N7182, N6903);
nand NAND2 (N13043, N13038, N10793);
nor NOR2 (N13044, N13031, N10760);
nor NOR2 (N13045, N13030, N10933);
or OR2 (N13046, N13044, N12461);
not NOT1 (N13047, N13020);
nor NOR4 (N13048, N13045, N11615, N9703, N1929);
or OR2 (N13049, N13047, N3923);
buf BUF1 (N13050, N13042);
and AND2 (N13051, N13041, N5659);
or OR2 (N13052, N13046, N3268);
not NOT1 (N13053, N13025);
buf BUF1 (N13054, N13043);
not NOT1 (N13055, N13051);
buf BUF1 (N13056, N13049);
nand NAND3 (N13057, N13055, N9262, N8698);
buf BUF1 (N13058, N13048);
or OR2 (N13059, N13040, N124);
not NOT1 (N13060, N13058);
xor XOR2 (N13061, N13057, N9082);
buf BUF1 (N13062, N13035);
nor NOR4 (N13063, N13056, N10815, N4797, N5368);
buf BUF1 (N13064, N13053);
xor XOR2 (N13065, N13033, N1470);
not NOT1 (N13066, N13052);
nand NAND3 (N13067, N13054, N12108, N10443);
nor NOR2 (N13068, N13064, N5758);
and AND4 (N13069, N13061, N3929, N7561, N3616);
and AND4 (N13070, N13067, N5839, N5987, N3199);
nor NOR2 (N13071, N13059, N8597);
nand NAND2 (N13072, N13063, N8549);
buf BUF1 (N13073, N13070);
and AND3 (N13074, N13060, N9138, N2305);
and AND2 (N13075, N13068, N7061);
buf BUF1 (N13076, N13073);
nand NAND4 (N13077, N13072, N9740, N4704, N8015);
nor NOR3 (N13078, N13071, N12399, N5409);
and AND4 (N13079, N13062, N5318, N3851, N312);
or OR4 (N13080, N13078, N7161, N3219, N3431);
buf BUF1 (N13081, N13065);
nand NAND3 (N13082, N13081, N5276, N355);
nand NAND4 (N13083, N13077, N10788, N3309, N4706);
xor XOR2 (N13084, N13080, N8049);
nand NAND2 (N13085, N13069, N11536);
not NOT1 (N13086, N13076);
nand NAND2 (N13087, N13050, N6573);
not NOT1 (N13088, N13074);
or OR2 (N13089, N13066, N7420);
buf BUF1 (N13090, N13088);
not NOT1 (N13091, N13090);
and AND2 (N13092, N13084, N9125);
not NOT1 (N13093, N13087);
and AND3 (N13094, N13075, N4316, N4226);
or OR4 (N13095, N13094, N1985, N7972, N1824);
and AND4 (N13096, N13091, N8704, N4580, N12009);
xor XOR2 (N13097, N13095, N10711);
not NOT1 (N13098, N13083);
xor XOR2 (N13099, N13085, N10563);
nor NOR2 (N13100, N13098, N11230);
or OR3 (N13101, N13093, N8635, N5256);
not NOT1 (N13102, N13082);
nand NAND4 (N13103, N13092, N3587, N12336, N3597);
buf BUF1 (N13104, N13103);
buf BUF1 (N13105, N13079);
xor XOR2 (N13106, N13104, N2926);
buf BUF1 (N13107, N13086);
xor XOR2 (N13108, N13102, N1499);
xor XOR2 (N13109, N13106, N7424);
xor XOR2 (N13110, N13107, N12430);
not NOT1 (N13111, N13089);
buf BUF1 (N13112, N13096);
buf BUF1 (N13113, N13110);
or OR3 (N13114, N13100, N3889, N8131);
and AND2 (N13115, N13099, N6115);
xor XOR2 (N13116, N13112, N688);
not NOT1 (N13117, N13111);
or OR2 (N13118, N13115, N3046);
xor XOR2 (N13119, N13097, N1290);
not NOT1 (N13120, N13105);
xor XOR2 (N13121, N13120, N3626);
buf BUF1 (N13122, N13118);
nor NOR2 (N13123, N13101, N8043);
nor NOR2 (N13124, N13109, N1872);
or OR4 (N13125, N13122, N7843, N3446, N2015);
xor XOR2 (N13126, N13117, N5200);
not NOT1 (N13127, N13121);
or OR2 (N13128, N13116, N6759);
buf BUF1 (N13129, N13124);
or OR3 (N13130, N13129, N9595, N9462);
nor NOR4 (N13131, N13114, N3864, N12546, N10418);
buf BUF1 (N13132, N13126);
not NOT1 (N13133, N13130);
or OR4 (N13134, N13128, N4681, N1307, N5203);
and AND4 (N13135, N13134, N99, N8184, N1337);
or OR3 (N13136, N13127, N577, N8089);
nor NOR2 (N13137, N13125, N1129);
or OR4 (N13138, N13113, N13048, N3814, N10932);
not NOT1 (N13139, N13135);
not NOT1 (N13140, N13132);
nand NAND4 (N13141, N13131, N11053, N12240, N13054);
xor XOR2 (N13142, N13141, N7362);
buf BUF1 (N13143, N13108);
and AND4 (N13144, N13123, N1169, N7964, N5779);
xor XOR2 (N13145, N13136, N4293);
buf BUF1 (N13146, N13140);
not NOT1 (N13147, N13142);
buf BUF1 (N13148, N13143);
nand NAND4 (N13149, N13144, N7048, N11096, N8720);
not NOT1 (N13150, N13138);
nand NAND2 (N13151, N13149, N6282);
xor XOR2 (N13152, N13139, N1805);
not NOT1 (N13153, N13152);
nor NOR3 (N13154, N13146, N9150, N6683);
not NOT1 (N13155, N13154);
nand NAND3 (N13156, N13145, N4498, N11587);
xor XOR2 (N13157, N13148, N2133);
nand NAND4 (N13158, N13155, N2314, N623, N12651);
not NOT1 (N13159, N13151);
or OR2 (N13160, N13150, N8387);
buf BUF1 (N13161, N13159);
nand NAND2 (N13162, N13153, N10597);
nand NAND2 (N13163, N13119, N12047);
xor XOR2 (N13164, N13162, N9588);
nand NAND4 (N13165, N13160, N9244, N8317, N11026);
and AND4 (N13166, N13165, N6933, N5744, N6398);
nor NOR3 (N13167, N13163, N10263, N2244);
not NOT1 (N13168, N13133);
and AND2 (N13169, N13158, N1653);
or OR4 (N13170, N13161, N4257, N1025, N7618);
not NOT1 (N13171, N13156);
not NOT1 (N13172, N13170);
or OR2 (N13173, N13137, N11986);
nor NOR4 (N13174, N13172, N12425, N12363, N11202);
nor NOR3 (N13175, N13168, N2764, N10747);
or OR3 (N13176, N13164, N454, N1134);
xor XOR2 (N13177, N13147, N8477);
nand NAND3 (N13178, N13175, N6276, N950);
or OR4 (N13179, N13173, N12432, N2913, N5353);
buf BUF1 (N13180, N13179);
not NOT1 (N13181, N13166);
nand NAND3 (N13182, N13178, N12791, N4170);
and AND3 (N13183, N13171, N7944, N3487);
and AND3 (N13184, N13180, N6197, N6483);
xor XOR2 (N13185, N13182, N10824);
nor NOR2 (N13186, N13167, N8677);
nor NOR3 (N13187, N13176, N7745, N141);
buf BUF1 (N13188, N13186);
xor XOR2 (N13189, N13174, N11768);
nand NAND4 (N13190, N13185, N9085, N6482, N3181);
or OR4 (N13191, N13169, N5997, N9597, N7842);
nand NAND2 (N13192, N13190, N4543);
not NOT1 (N13193, N13189);
buf BUF1 (N13194, N13183);
xor XOR2 (N13195, N13177, N5538);
not NOT1 (N13196, N13157);
or OR4 (N13197, N13184, N1021, N12184, N10250);
not NOT1 (N13198, N13187);
xor XOR2 (N13199, N13193, N10354);
buf BUF1 (N13200, N13194);
or OR3 (N13201, N13192, N8502, N11017);
nor NOR4 (N13202, N13196, N6359, N8956, N4903);
nand NAND4 (N13203, N13191, N1453, N11206, N3066);
xor XOR2 (N13204, N13202, N1103);
and AND3 (N13205, N13197, N3227, N2360);
nor NOR3 (N13206, N13205, N10947, N605);
buf BUF1 (N13207, N13204);
xor XOR2 (N13208, N13181, N5754);
not NOT1 (N13209, N13201);
xor XOR2 (N13210, N13206, N11163);
nand NAND2 (N13211, N13210, N9694);
not NOT1 (N13212, N13188);
nand NAND4 (N13213, N13198, N3775, N116, N261);
nor NOR2 (N13214, N13211, N6158);
nand NAND4 (N13215, N13203, N9898, N5240, N4515);
not NOT1 (N13216, N13200);
or OR2 (N13217, N13208, N5768);
not NOT1 (N13218, N13216);
nand NAND2 (N13219, N13215, N2256);
buf BUF1 (N13220, N13219);
not NOT1 (N13221, N13220);
nor NOR2 (N13222, N13209, N862);
not NOT1 (N13223, N13195);
or OR2 (N13224, N13217, N8368);
nand NAND3 (N13225, N13223, N2291, N3014);
or OR4 (N13226, N13221, N8284, N3354, N1843);
not NOT1 (N13227, N13226);
nand NAND4 (N13228, N13225, N4765, N12240, N3509);
not NOT1 (N13229, N13212);
nand NAND3 (N13230, N13222, N1687, N2055);
not NOT1 (N13231, N13228);
or OR4 (N13232, N13231, N3011, N290, N7746);
buf BUF1 (N13233, N13230);
xor XOR2 (N13234, N13218, N11641);
or OR2 (N13235, N13232, N10903);
buf BUF1 (N13236, N13213);
xor XOR2 (N13237, N13236, N12971);
not NOT1 (N13238, N13233);
buf BUF1 (N13239, N13235);
buf BUF1 (N13240, N13224);
buf BUF1 (N13241, N13207);
buf BUF1 (N13242, N13214);
and AND3 (N13243, N13242, N11683, N10809);
and AND2 (N13244, N13229, N1464);
not NOT1 (N13245, N13243);
nand NAND2 (N13246, N13238, N5760);
nand NAND4 (N13247, N13240, N4693, N695, N843);
not NOT1 (N13248, N13246);
or OR4 (N13249, N13247, N7057, N7217, N6922);
nor NOR4 (N13250, N13248, N4032, N7156, N12933);
or OR3 (N13251, N13227, N6141, N6652);
nor NOR2 (N13252, N13234, N10242);
nor NOR2 (N13253, N13241, N300);
nor NOR2 (N13254, N13249, N1668);
not NOT1 (N13255, N13254);
or OR2 (N13256, N13239, N2146);
and AND4 (N13257, N13237, N3006, N12261, N7412);
nand NAND2 (N13258, N13245, N3417);
nand NAND4 (N13259, N13255, N10278, N6681, N11156);
buf BUF1 (N13260, N13252);
buf BUF1 (N13261, N13256);
nor NOR4 (N13262, N13257, N5927, N955, N8937);
nor NOR3 (N13263, N13244, N13124, N4452);
and AND3 (N13264, N13250, N11759, N11980);
not NOT1 (N13265, N13199);
buf BUF1 (N13266, N13263);
xor XOR2 (N13267, N13261, N12967);
or OR2 (N13268, N13251, N11956);
buf BUF1 (N13269, N13267);
nand NAND3 (N13270, N13264, N9352, N12797);
and AND4 (N13271, N13262, N5551, N2310, N8214);
xor XOR2 (N13272, N13253, N422);
xor XOR2 (N13273, N13268, N13010);
nor NOR2 (N13274, N13270, N11332);
not NOT1 (N13275, N13260);
or OR2 (N13276, N13266, N6531);
nor NOR2 (N13277, N13265, N6256);
xor XOR2 (N13278, N13276, N3642);
and AND3 (N13279, N13259, N4390, N998);
buf BUF1 (N13280, N13272);
nand NAND2 (N13281, N13275, N2683);
or OR3 (N13282, N13258, N479, N8729);
nor NOR3 (N13283, N13273, N9289, N12868);
xor XOR2 (N13284, N13279, N2809);
nand NAND4 (N13285, N13284, N12331, N5567, N10300);
nand NAND4 (N13286, N13269, N3296, N765, N11446);
xor XOR2 (N13287, N13274, N1473);
not NOT1 (N13288, N13287);
buf BUF1 (N13289, N13281);
not NOT1 (N13290, N13283);
nand NAND4 (N13291, N13280, N12339, N4654, N497);
not NOT1 (N13292, N13286);
xor XOR2 (N13293, N13290, N3780);
nor NOR3 (N13294, N13282, N13269, N11458);
not NOT1 (N13295, N13278);
xor XOR2 (N13296, N13293, N9332);
or OR4 (N13297, N13289, N3434, N335, N4378);
and AND2 (N13298, N13294, N3103);
and AND4 (N13299, N13295, N9006, N9728, N6608);
nor NOR3 (N13300, N13298, N11815, N36);
and AND3 (N13301, N13296, N2064, N6483);
xor XOR2 (N13302, N13285, N316);
xor XOR2 (N13303, N13291, N556);
buf BUF1 (N13304, N13301);
buf BUF1 (N13305, N13288);
or OR4 (N13306, N13271, N9918, N652, N7436);
and AND2 (N13307, N13300, N311);
buf BUF1 (N13308, N13304);
not NOT1 (N13309, N13302);
buf BUF1 (N13310, N13306);
buf BUF1 (N13311, N13307);
xor XOR2 (N13312, N13277, N899);
or OR2 (N13313, N13312, N10616);
nand NAND3 (N13314, N13305, N1566, N11616);
xor XOR2 (N13315, N13297, N3802);
not NOT1 (N13316, N13313);
buf BUF1 (N13317, N13311);
and AND2 (N13318, N13317, N1201);
or OR4 (N13319, N13314, N11034, N10087, N7290);
xor XOR2 (N13320, N13292, N10596);
not NOT1 (N13321, N13309);
or OR3 (N13322, N13310, N8702, N2528);
not NOT1 (N13323, N13316);
nor NOR3 (N13324, N13318, N12317, N304);
xor XOR2 (N13325, N13315, N11391);
nand NAND3 (N13326, N13320, N2704, N6390);
not NOT1 (N13327, N13303);
buf BUF1 (N13328, N13327);
xor XOR2 (N13329, N13322, N295);
xor XOR2 (N13330, N13323, N4165);
xor XOR2 (N13331, N13330, N10513);
not NOT1 (N13332, N13331);
or OR4 (N13333, N13321, N12174, N8227, N169);
nand NAND3 (N13334, N13325, N11536, N9460);
nor NOR3 (N13335, N13332, N1255, N2774);
nor NOR4 (N13336, N13335, N2989, N8084, N1595);
nor NOR2 (N13337, N13336, N10283);
nand NAND4 (N13338, N13329, N11008, N2431, N8149);
nor NOR3 (N13339, N13328, N9064, N10525);
nand NAND4 (N13340, N13334, N7453, N4892, N11905);
nor NOR2 (N13341, N13337, N12273);
buf BUF1 (N13342, N13339);
and AND3 (N13343, N13326, N7010, N8932);
or OR4 (N13344, N13343, N3577, N13246, N7021);
buf BUF1 (N13345, N13308);
buf BUF1 (N13346, N13342);
nor NOR4 (N13347, N13338, N12205, N1021, N9762);
xor XOR2 (N13348, N13319, N5501);
nand NAND2 (N13349, N13346, N1038);
or OR3 (N13350, N13299, N2016, N2098);
nor NOR2 (N13351, N13324, N11051);
buf BUF1 (N13352, N13340);
nor NOR4 (N13353, N13348, N5836, N11439, N2240);
or OR2 (N13354, N13345, N6299);
xor XOR2 (N13355, N13349, N11488);
buf BUF1 (N13356, N13354);
nand NAND3 (N13357, N13347, N9257, N8772);
or OR3 (N13358, N13351, N1677, N5295);
not NOT1 (N13359, N13344);
nor NOR4 (N13360, N13357, N1041, N8562, N11459);
and AND4 (N13361, N13355, N6435, N10575, N12092);
nor NOR4 (N13362, N13358, N6511, N5987, N6603);
nor NOR2 (N13363, N13341, N12013);
xor XOR2 (N13364, N13353, N11584);
or OR2 (N13365, N13352, N5290);
or OR4 (N13366, N13362, N2824, N9582, N6280);
and AND2 (N13367, N13363, N9763);
nand NAND3 (N13368, N13361, N1254, N792);
nor NOR3 (N13369, N13365, N8926, N8490);
nor NOR2 (N13370, N13359, N564);
nor NOR4 (N13371, N13368, N10055, N4661, N12946);
and AND3 (N13372, N13366, N8942, N11288);
not NOT1 (N13373, N13360);
nand NAND3 (N13374, N13372, N9026, N11416);
nand NAND3 (N13375, N13374, N11283, N3036);
not NOT1 (N13376, N13369);
and AND4 (N13377, N13364, N5184, N11642, N175);
and AND3 (N13378, N13373, N12795, N7730);
and AND2 (N13379, N13375, N13009);
and AND3 (N13380, N13376, N10616, N10555);
not NOT1 (N13381, N13379);
buf BUF1 (N13382, N13377);
not NOT1 (N13383, N13370);
nor NOR4 (N13384, N13333, N5938, N3975, N2278);
and AND3 (N13385, N13371, N8454, N8954);
buf BUF1 (N13386, N13381);
nand NAND3 (N13387, N13386, N165, N272);
buf BUF1 (N13388, N13383);
buf BUF1 (N13389, N13380);
nand NAND2 (N13390, N13387, N7542);
xor XOR2 (N13391, N13389, N11460);
buf BUF1 (N13392, N13367);
nor NOR3 (N13393, N13392, N9470, N11081);
nor NOR3 (N13394, N13382, N7587, N5688);
and AND2 (N13395, N13390, N8696);
nand NAND2 (N13396, N13350, N1347);
and AND2 (N13397, N13385, N8812);
xor XOR2 (N13398, N13388, N5439);
nand NAND2 (N13399, N13395, N4161);
buf BUF1 (N13400, N13399);
xor XOR2 (N13401, N13356, N8658);
nand NAND4 (N13402, N13393, N1440, N11567, N9019);
not NOT1 (N13403, N13398);
nand NAND3 (N13404, N13394, N1663, N11787);
nand NAND4 (N13405, N13401, N8142, N11642, N12098);
nand NAND2 (N13406, N13400, N6004);
nand NAND2 (N13407, N13403, N11457);
nor NOR4 (N13408, N13402, N12860, N3393, N9888);
buf BUF1 (N13409, N13396);
xor XOR2 (N13410, N13404, N3502);
nand NAND2 (N13411, N13409, N5860);
nand NAND3 (N13412, N13411, N6065, N13159);
or OR2 (N13413, N13407, N5128);
nand NAND3 (N13414, N13397, N3357, N4305);
nor NOR3 (N13415, N13410, N9077, N2641);
nor NOR3 (N13416, N13413, N10390, N8702);
nor NOR2 (N13417, N13384, N12021);
nand NAND2 (N13418, N13408, N6286);
and AND2 (N13419, N13414, N1826);
nand NAND2 (N13420, N13416, N3430);
or OR4 (N13421, N13420, N621, N2068, N572);
buf BUF1 (N13422, N13421);
not NOT1 (N13423, N13415);
nand NAND2 (N13424, N13422, N3095);
buf BUF1 (N13425, N13406);
nor NOR3 (N13426, N13419, N5307, N13330);
buf BUF1 (N13427, N13412);
not NOT1 (N13428, N13405);
nand NAND4 (N13429, N13418, N5638, N8683, N11317);
or OR3 (N13430, N13425, N9100, N12468);
nand NAND4 (N13431, N13391, N6324, N6995, N1934);
and AND3 (N13432, N13429, N7731, N328);
buf BUF1 (N13433, N13417);
nand NAND3 (N13434, N13432, N5237, N170);
and AND2 (N13435, N13431, N6668);
buf BUF1 (N13436, N13423);
buf BUF1 (N13437, N13435);
or OR2 (N13438, N13434, N3943);
buf BUF1 (N13439, N13424);
not NOT1 (N13440, N13433);
and AND3 (N13441, N13437, N7781, N4882);
and AND4 (N13442, N13427, N8361, N3522, N11124);
xor XOR2 (N13443, N13428, N12534);
nor NOR4 (N13444, N13441, N2478, N4687, N8944);
not NOT1 (N13445, N13378);
xor XOR2 (N13446, N13430, N7665);
nor NOR3 (N13447, N13442, N3991, N4521);
or OR2 (N13448, N13445, N12538);
xor XOR2 (N13449, N13436, N8392);
and AND3 (N13450, N13448, N3227, N12447);
or OR3 (N13451, N13447, N2735, N9702);
and AND4 (N13452, N13451, N3559, N8516, N6569);
and AND2 (N13453, N13438, N9426);
nand NAND2 (N13454, N13444, N11839);
nand NAND3 (N13455, N13440, N7898, N10091);
not NOT1 (N13456, N13455);
xor XOR2 (N13457, N13456, N6047);
buf BUF1 (N13458, N13452);
and AND2 (N13459, N13450, N7241);
not NOT1 (N13460, N13449);
xor XOR2 (N13461, N13460, N11594);
xor XOR2 (N13462, N13446, N1510);
and AND3 (N13463, N13458, N3410, N8895);
xor XOR2 (N13464, N13443, N12198);
and AND4 (N13465, N13454, N9472, N4427, N12852);
not NOT1 (N13466, N13439);
nand NAND3 (N13467, N13465, N13241, N2916);
not NOT1 (N13468, N13426);
nor NOR2 (N13469, N13461, N9765);
or OR4 (N13470, N13459, N3364, N10884, N9069);
nor NOR4 (N13471, N13469, N13029, N2877, N2718);
not NOT1 (N13472, N13462);
or OR3 (N13473, N13463, N12704, N3849);
or OR2 (N13474, N13468, N11473);
or OR4 (N13475, N13464, N12083, N7223, N10244);
xor XOR2 (N13476, N13453, N13452);
and AND3 (N13477, N13474, N3395, N10247);
nand NAND2 (N13478, N13466, N8525);
or OR3 (N13479, N13475, N8261, N2189);
nand NAND2 (N13480, N13479, N3679);
not NOT1 (N13481, N13471);
or OR2 (N13482, N13467, N1906);
nor NOR4 (N13483, N13481, N4533, N6431, N10470);
xor XOR2 (N13484, N13482, N3251);
xor XOR2 (N13485, N13484, N11310);
nand NAND2 (N13486, N13473, N9823);
xor XOR2 (N13487, N13480, N7253);
buf BUF1 (N13488, N13457);
nor NOR3 (N13489, N13476, N8483, N932);
or OR4 (N13490, N13488, N13019, N2027, N1522);
nand NAND2 (N13491, N13489, N12346);
nand NAND2 (N13492, N13472, N3632);
not NOT1 (N13493, N13485);
nand NAND2 (N13494, N13491, N12395);
buf BUF1 (N13495, N13494);
nor NOR4 (N13496, N13478, N1688, N7705, N7848);
nand NAND3 (N13497, N13493, N6930, N8131);
nand NAND3 (N13498, N13486, N679, N13420);
and AND3 (N13499, N13477, N12232, N8463);
or OR4 (N13500, N13499, N12211, N7485, N6688);
buf BUF1 (N13501, N13487);
buf BUF1 (N13502, N13483);
nor NOR2 (N13503, N13496, N6210);
nor NOR2 (N13504, N13495, N12265);
and AND4 (N13505, N13502, N12918, N11664, N12821);
or OR2 (N13506, N13501, N12272);
and AND4 (N13507, N13503, N4528, N12894, N10904);
buf BUF1 (N13508, N13497);
or OR2 (N13509, N13470, N8848);
or OR3 (N13510, N13492, N5307, N11650);
buf BUF1 (N13511, N13506);
not NOT1 (N13512, N13500);
buf BUF1 (N13513, N13512);
and AND3 (N13514, N13490, N7505, N11395);
xor XOR2 (N13515, N13514, N11455);
not NOT1 (N13516, N13507);
or OR2 (N13517, N13511, N8845);
buf BUF1 (N13518, N13516);
nor NOR3 (N13519, N13508, N6634, N276);
nor NOR3 (N13520, N13504, N5271, N6158);
nor NOR2 (N13521, N13515, N13214);
nand NAND2 (N13522, N13498, N4115);
buf BUF1 (N13523, N13513);
and AND3 (N13524, N13510, N6733, N4350);
nand NAND2 (N13525, N13521, N5316);
xor XOR2 (N13526, N13509, N1976);
not NOT1 (N13527, N13523);
buf BUF1 (N13528, N13520);
xor XOR2 (N13529, N13528, N6027);
not NOT1 (N13530, N13526);
nand NAND4 (N13531, N13529, N1098, N1240, N13284);
nand NAND2 (N13532, N13505, N3530);
buf BUF1 (N13533, N13524);
or OR4 (N13534, N13518, N6539, N9258, N9619);
not NOT1 (N13535, N13525);
nand NAND3 (N13536, N13532, N4862, N3457);
or OR4 (N13537, N13535, N2283, N3716, N5509);
not NOT1 (N13538, N13517);
xor XOR2 (N13539, N13519, N425);
and AND3 (N13540, N13531, N9051, N7091);
xor XOR2 (N13541, N13534, N2390);
xor XOR2 (N13542, N13538, N11939);
nand NAND3 (N13543, N13522, N12181, N3715);
buf BUF1 (N13544, N13536);
xor XOR2 (N13545, N13537, N387);
nand NAND3 (N13546, N13545, N1544, N4232);
buf BUF1 (N13547, N13541);
or OR3 (N13548, N13544, N3902, N3588);
or OR2 (N13549, N13527, N2062);
buf BUF1 (N13550, N13548);
nand NAND4 (N13551, N13530, N8581, N1435, N12880);
nor NOR4 (N13552, N13547, N11065, N10323, N7299);
nand NAND3 (N13553, N13546, N6562, N7815);
not NOT1 (N13554, N13553);
not NOT1 (N13555, N13533);
not NOT1 (N13556, N13554);
buf BUF1 (N13557, N13549);
buf BUF1 (N13558, N13542);
or OR2 (N13559, N13558, N8744);
nor NOR3 (N13560, N13550, N2683, N13495);
not NOT1 (N13561, N13557);
nand NAND4 (N13562, N13559, N7192, N7797, N5503);
nor NOR4 (N13563, N13543, N9637, N2479, N2297);
not NOT1 (N13564, N13560);
not NOT1 (N13565, N13561);
nor NOR2 (N13566, N13555, N9911);
not NOT1 (N13567, N13556);
nand NAND4 (N13568, N13565, N7318, N7655, N3885);
and AND2 (N13569, N13552, N12231);
xor XOR2 (N13570, N13568, N9716);
or OR3 (N13571, N13551, N1627, N7751);
not NOT1 (N13572, N13569);
nor NOR2 (N13573, N13563, N697);
xor XOR2 (N13574, N13564, N717);
or OR3 (N13575, N13539, N737, N9652);
not NOT1 (N13576, N13567);
and AND4 (N13577, N13540, N827, N10370, N11342);
nor NOR2 (N13578, N13562, N10663);
or OR4 (N13579, N13570, N11786, N12446, N1115);
not NOT1 (N13580, N13579);
buf BUF1 (N13581, N13575);
nand NAND2 (N13582, N13577, N9978);
nor NOR4 (N13583, N13571, N11412, N1964, N11996);
not NOT1 (N13584, N13582);
nand NAND2 (N13585, N13573, N3698);
xor XOR2 (N13586, N13583, N12957);
or OR2 (N13587, N13586, N10524);
buf BUF1 (N13588, N13581);
xor XOR2 (N13589, N13574, N13467);
or OR4 (N13590, N13566, N786, N1509, N3253);
nor NOR2 (N13591, N13584, N10112);
or OR3 (N13592, N13587, N11304, N9997);
nor NOR4 (N13593, N13592, N6906, N8024, N9823);
buf BUF1 (N13594, N13580);
or OR4 (N13595, N13578, N12591, N2943, N439);
not NOT1 (N13596, N13594);
nand NAND3 (N13597, N13596, N853, N11483);
nor NOR4 (N13598, N13589, N4390, N13004, N12031);
not NOT1 (N13599, N13591);
xor XOR2 (N13600, N13597, N4758);
nor NOR3 (N13601, N13595, N13228, N2868);
nor NOR3 (N13602, N13588, N8715, N3029);
xor XOR2 (N13603, N13593, N5299);
not NOT1 (N13604, N13600);
xor XOR2 (N13605, N13598, N12225);
nor NOR4 (N13606, N13605, N10833, N9822, N8070);
nor NOR2 (N13607, N13585, N11879);
not NOT1 (N13608, N13604);
or OR4 (N13609, N13607, N2653, N4117, N7704);
buf BUF1 (N13610, N13603);
buf BUF1 (N13611, N13601);
buf BUF1 (N13612, N13572);
nand NAND2 (N13613, N13602, N1881);
buf BUF1 (N13614, N13612);
not NOT1 (N13615, N13590);
or OR3 (N13616, N13606, N8971, N4170);
not NOT1 (N13617, N13576);
not NOT1 (N13618, N13608);
or OR2 (N13619, N13617, N7726);
not NOT1 (N13620, N13609);
nor NOR2 (N13621, N13614, N11348);
buf BUF1 (N13622, N13616);
or OR2 (N13623, N13619, N6586);
or OR2 (N13624, N13621, N4959);
xor XOR2 (N13625, N13610, N2005);
buf BUF1 (N13626, N13611);
nor NOR2 (N13627, N13620, N4935);
nand NAND2 (N13628, N13623, N11813);
and AND4 (N13629, N13613, N13103, N9889, N3938);
xor XOR2 (N13630, N13626, N3881);
or OR2 (N13631, N13628, N2047);
not NOT1 (N13632, N13624);
and AND4 (N13633, N13631, N7500, N5849, N9902);
not NOT1 (N13634, N13629);
xor XOR2 (N13635, N13627, N11152);
xor XOR2 (N13636, N13625, N4595);
or OR2 (N13637, N13615, N11115);
xor XOR2 (N13638, N13634, N13174);
xor XOR2 (N13639, N13599, N6609);
and AND2 (N13640, N13632, N1733);
or OR3 (N13641, N13622, N5490, N8154);
xor XOR2 (N13642, N13638, N11992);
buf BUF1 (N13643, N13640);
nor NOR2 (N13644, N13641, N5876);
or OR4 (N13645, N13635, N12062, N9096, N12503);
xor XOR2 (N13646, N13645, N9710);
and AND2 (N13647, N13618, N10595);
xor XOR2 (N13648, N13636, N6539);
buf BUF1 (N13649, N13642);
xor XOR2 (N13650, N13647, N8117);
not NOT1 (N13651, N13650);
nand NAND2 (N13652, N13643, N10499);
or OR2 (N13653, N13630, N2682);
or OR3 (N13654, N13652, N1787, N5983);
or OR2 (N13655, N13653, N2160);
and AND3 (N13656, N13639, N9514, N49);
xor XOR2 (N13657, N13649, N5445);
nand NAND3 (N13658, N13633, N8516, N11364);
or OR2 (N13659, N13658, N11318);
nor NOR3 (N13660, N13659, N4845, N4752);
and AND2 (N13661, N13660, N12689);
buf BUF1 (N13662, N13654);
buf BUF1 (N13663, N13655);
nor NOR2 (N13664, N13657, N8912);
nand NAND2 (N13665, N13637, N9407);
xor XOR2 (N13666, N13656, N8467);
not NOT1 (N13667, N13664);
nor NOR3 (N13668, N13651, N2906, N2086);
not NOT1 (N13669, N13668);
or OR4 (N13670, N13661, N151, N5061, N6877);
and AND4 (N13671, N13646, N216, N3354, N11451);
xor XOR2 (N13672, N13663, N12380);
buf BUF1 (N13673, N13671);
or OR3 (N13674, N13672, N10581, N10508);
buf BUF1 (N13675, N13670);
buf BUF1 (N13676, N13667);
nor NOR2 (N13677, N13674, N1721);
nor NOR4 (N13678, N13644, N2192, N9789, N7502);
not NOT1 (N13679, N13669);
not NOT1 (N13680, N13666);
not NOT1 (N13681, N13673);
nand NAND3 (N13682, N13678, N9519, N660);
nand NAND2 (N13683, N13676, N5916);
nand NAND3 (N13684, N13662, N3949, N720);
and AND2 (N13685, N13680, N13672);
not NOT1 (N13686, N13683);
xor XOR2 (N13687, N13665, N10697);
xor XOR2 (N13688, N13686, N7580);
nor NOR2 (N13689, N13684, N3088);
or OR4 (N13690, N13675, N612, N11287, N1288);
and AND2 (N13691, N13679, N1325);
nand NAND2 (N13692, N13685, N13150);
xor XOR2 (N13693, N13687, N13525);
xor XOR2 (N13694, N13682, N6767);
buf BUF1 (N13695, N13688);
xor XOR2 (N13696, N13681, N7470);
nand NAND4 (N13697, N13696, N9216, N1256, N11279);
xor XOR2 (N13698, N13694, N8334);
nor NOR4 (N13699, N13695, N2143, N1067, N3946);
or OR2 (N13700, N13689, N12999);
nor NOR2 (N13701, N13648, N7163);
buf BUF1 (N13702, N13693);
and AND3 (N13703, N13701, N1350, N11891);
buf BUF1 (N13704, N13677);
and AND4 (N13705, N13697, N75, N1355, N1483);
not NOT1 (N13706, N13702);
nand NAND4 (N13707, N13692, N4753, N4202, N332);
or OR3 (N13708, N13705, N640, N12451);
xor XOR2 (N13709, N13704, N5966);
or OR4 (N13710, N13703, N10331, N2641, N3362);
not NOT1 (N13711, N13709);
nand NAND2 (N13712, N13691, N6652);
or OR2 (N13713, N13698, N9610);
nand NAND3 (N13714, N13710, N549, N12205);
xor XOR2 (N13715, N13706, N2681);
nor NOR4 (N13716, N13707, N4539, N13353, N1446);
buf BUF1 (N13717, N13711);
nor NOR2 (N13718, N13717, N711);
buf BUF1 (N13719, N13714);
xor XOR2 (N13720, N13708, N7700);
not NOT1 (N13721, N13718);
buf BUF1 (N13722, N13700);
buf BUF1 (N13723, N13690);
or OR4 (N13724, N13716, N8925, N3101, N4071);
not NOT1 (N13725, N13724);
nand NAND3 (N13726, N13723, N1228, N2675);
xor XOR2 (N13727, N13722, N10147);
xor XOR2 (N13728, N13721, N11943);
and AND3 (N13729, N13713, N11434, N1912);
nor NOR2 (N13730, N13720, N2805);
nand NAND4 (N13731, N13725, N12843, N2599, N25);
and AND4 (N13732, N13719, N12289, N2019, N6472);
buf BUF1 (N13733, N13699);
nand NAND2 (N13734, N13731, N8597);
xor XOR2 (N13735, N13726, N869);
nor NOR4 (N13736, N13733, N7915, N8128, N3149);
nor NOR2 (N13737, N13715, N1673);
nand NAND3 (N13738, N13737, N6918, N5207);
xor XOR2 (N13739, N13732, N10886);
buf BUF1 (N13740, N13738);
buf BUF1 (N13741, N13740);
and AND2 (N13742, N13730, N3121);
or OR3 (N13743, N13728, N12570, N7193);
or OR3 (N13744, N13742, N2304, N3572);
nor NOR2 (N13745, N13727, N8045);
nor NOR4 (N13746, N13734, N4027, N7911, N2730);
nand NAND4 (N13747, N13746, N202, N5409, N3698);
buf BUF1 (N13748, N13743);
and AND2 (N13749, N13741, N12155);
xor XOR2 (N13750, N13747, N7970);
buf BUF1 (N13751, N13744);
nor NOR3 (N13752, N13729, N7441, N2595);
and AND2 (N13753, N13739, N5467);
buf BUF1 (N13754, N13750);
nor NOR4 (N13755, N13749, N5318, N12922, N12497);
or OR3 (N13756, N13745, N12326, N3176);
xor XOR2 (N13757, N13753, N9317);
buf BUF1 (N13758, N13736);
not NOT1 (N13759, N13735);
not NOT1 (N13760, N13712);
or OR4 (N13761, N13754, N6742, N4008, N1287);
buf BUF1 (N13762, N13751);
nor NOR2 (N13763, N13762, N8250);
and AND2 (N13764, N13760, N6034);
not NOT1 (N13765, N13748);
nand NAND4 (N13766, N13755, N3604, N13442, N8845);
nand NAND3 (N13767, N13756, N2344, N5644);
not NOT1 (N13768, N13765);
nor NOR4 (N13769, N13768, N13010, N2419, N12469);
not NOT1 (N13770, N13769);
not NOT1 (N13771, N13758);
nor NOR2 (N13772, N13763, N8658);
or OR3 (N13773, N13759, N8863, N1933);
not NOT1 (N13774, N13771);
buf BUF1 (N13775, N13774);
and AND3 (N13776, N13766, N12742, N2053);
nand NAND4 (N13777, N13772, N2314, N1521, N11017);
nand NAND4 (N13778, N13770, N4935, N7892, N6737);
xor XOR2 (N13779, N13761, N2064);
xor XOR2 (N13780, N13767, N4164);
not NOT1 (N13781, N13780);
xor XOR2 (N13782, N13775, N1555);
or OR3 (N13783, N13782, N2197, N11200);
nor NOR4 (N13784, N13779, N5794, N2441, N4234);
not NOT1 (N13785, N13783);
buf BUF1 (N13786, N13781);
or OR3 (N13787, N13777, N9026, N9503);
buf BUF1 (N13788, N13778);
xor XOR2 (N13789, N13757, N23);
nand NAND3 (N13790, N13752, N2198, N12070);
and AND4 (N13791, N13776, N11953, N10337, N5247);
not NOT1 (N13792, N13788);
xor XOR2 (N13793, N13792, N7884);
nor NOR4 (N13794, N13785, N9332, N5553, N12688);
nand NAND2 (N13795, N13793, N33);
nor NOR4 (N13796, N13795, N6069, N8807, N12303);
or OR4 (N13797, N13789, N11900, N13544, N2384);
xor XOR2 (N13798, N13790, N6694);
xor XOR2 (N13799, N13794, N736);
xor XOR2 (N13800, N13798, N10057);
buf BUF1 (N13801, N13787);
and AND4 (N13802, N13801, N2250, N5527, N11213);
or OR3 (N13803, N13799, N8774, N4680);
nor NOR4 (N13804, N13791, N2923, N12285, N4346);
nor NOR3 (N13805, N13804, N5784, N8577);
nand NAND2 (N13806, N13784, N3280);
nor NOR2 (N13807, N13805, N10858);
xor XOR2 (N13808, N13802, N193);
or OR2 (N13809, N13808, N10881);
buf BUF1 (N13810, N13809);
buf BUF1 (N13811, N13786);
nand NAND3 (N13812, N13806, N2012, N7796);
not NOT1 (N13813, N13773);
buf BUF1 (N13814, N13797);
nand NAND3 (N13815, N13810, N5465, N5769);
buf BUF1 (N13816, N13812);
nor NOR3 (N13817, N13796, N198, N6119);
nor NOR2 (N13818, N13800, N11921);
not NOT1 (N13819, N13815);
and AND3 (N13820, N13807, N9802, N2407);
or OR4 (N13821, N13803, N7481, N8800, N3359);
xor XOR2 (N13822, N13817, N5648);
xor XOR2 (N13823, N13822, N2679);
nor NOR2 (N13824, N13821, N9694);
and AND4 (N13825, N13814, N8818, N7039, N8641);
xor XOR2 (N13826, N13811, N1153);
not NOT1 (N13827, N13818);
xor XOR2 (N13828, N13764, N11366);
nand NAND2 (N13829, N13813, N8943);
nor NOR4 (N13830, N13819, N8450, N7506, N2464);
nand NAND3 (N13831, N13828, N8648, N2657);
nor NOR3 (N13832, N13816, N5517, N843);
nor NOR3 (N13833, N13829, N9688, N3790);
buf BUF1 (N13834, N13827);
not NOT1 (N13835, N13825);
nor NOR2 (N13836, N13823, N6054);
not NOT1 (N13837, N13832);
buf BUF1 (N13838, N13833);
xor XOR2 (N13839, N13830, N10958);
nor NOR4 (N13840, N13834, N9448, N2111, N3866);
and AND4 (N13841, N13826, N6102, N8916, N6245);
nand NAND4 (N13842, N13838, N607, N2417, N1270);
nor NOR2 (N13843, N13831, N4449);
or OR2 (N13844, N13820, N6602);
and AND3 (N13845, N13836, N1774, N12421);
buf BUF1 (N13846, N13835);
nor NOR3 (N13847, N13843, N5976, N8961);
xor XOR2 (N13848, N13842, N2239);
nand NAND2 (N13849, N13841, N11698);
xor XOR2 (N13850, N13846, N3391);
or OR4 (N13851, N13837, N487, N7793, N10529);
not NOT1 (N13852, N13851);
and AND2 (N13853, N13824, N10830);
not NOT1 (N13854, N13849);
not NOT1 (N13855, N13845);
and AND3 (N13856, N13853, N12752, N8297);
xor XOR2 (N13857, N13840, N5170);
nand NAND4 (N13858, N13839, N10020, N1902, N2861);
nand NAND3 (N13859, N13854, N3255, N8339);
xor XOR2 (N13860, N13856, N1330);
not NOT1 (N13861, N13847);
nor NOR3 (N13862, N13852, N1582, N2522);
buf BUF1 (N13863, N13860);
nor NOR3 (N13864, N13855, N3097, N8361);
or OR4 (N13865, N13857, N7499, N7292, N10347);
and AND3 (N13866, N13863, N6233, N8574);
nor NOR3 (N13867, N13861, N4729, N7291);
and AND4 (N13868, N13859, N9666, N2390, N4538);
nor NOR3 (N13869, N13866, N8388, N11471);
xor XOR2 (N13870, N13862, N9785);
xor XOR2 (N13871, N13865, N2846);
or OR2 (N13872, N13858, N106);
and AND4 (N13873, N13867, N9696, N4291, N3403);
and AND4 (N13874, N13848, N1609, N2887, N3911);
not NOT1 (N13875, N13868);
xor XOR2 (N13876, N13869, N8194);
xor XOR2 (N13877, N13864, N2789);
xor XOR2 (N13878, N13876, N5113);
or OR3 (N13879, N13877, N1149, N10606);
nand NAND2 (N13880, N13874, N8339);
or OR3 (N13881, N13879, N9535, N7160);
and AND3 (N13882, N13850, N228, N7077);
buf BUF1 (N13883, N13881);
not NOT1 (N13884, N13882);
nor NOR3 (N13885, N13870, N12421, N12140);
xor XOR2 (N13886, N13875, N2934);
xor XOR2 (N13887, N13883, N4361);
buf BUF1 (N13888, N13887);
nor NOR3 (N13889, N13878, N4049, N6062);
and AND4 (N13890, N13886, N13165, N5096, N1517);
nor NOR2 (N13891, N13871, N7738);
not NOT1 (N13892, N13880);
nand NAND4 (N13893, N13884, N4470, N3415, N3761);
or OR4 (N13894, N13892, N4943, N2062, N2906);
nor NOR4 (N13895, N13891, N7547, N10706, N8268);
nor NOR3 (N13896, N13895, N8148, N5801);
and AND2 (N13897, N13896, N145);
nand NAND4 (N13898, N13873, N7966, N13198, N7657);
and AND4 (N13899, N13888, N2168, N2437, N9461);
xor XOR2 (N13900, N13893, N3362);
buf BUF1 (N13901, N13872);
buf BUF1 (N13902, N13901);
or OR4 (N13903, N13899, N1327, N8680, N7524);
not NOT1 (N13904, N13903);
not NOT1 (N13905, N13900);
nand NAND3 (N13906, N13890, N11099, N5710);
not NOT1 (N13907, N13906);
nor NOR2 (N13908, N13898, N6721);
nand NAND3 (N13909, N13897, N11110, N11163);
nand NAND3 (N13910, N13902, N9134, N9898);
or OR4 (N13911, N13908, N7537, N8354, N3860);
buf BUF1 (N13912, N13911);
nor NOR3 (N13913, N13909, N3130, N3192);
nand NAND4 (N13914, N13905, N4618, N1477, N2560);
and AND3 (N13915, N13913, N1836, N9008);
not NOT1 (N13916, N13889);
or OR3 (N13917, N13907, N3806, N7832);
xor XOR2 (N13918, N13912, N6614);
nand NAND4 (N13919, N13904, N1105, N4052, N4259);
and AND3 (N13920, N13917, N12275, N12303);
or OR2 (N13921, N13894, N6383);
nor NOR2 (N13922, N13919, N6906);
and AND4 (N13923, N13910, N6548, N1352, N12650);
not NOT1 (N13924, N13918);
and AND4 (N13925, N13923, N10181, N13017, N8658);
buf BUF1 (N13926, N13920);
nor NOR4 (N13927, N13915, N3660, N12769, N9577);
not NOT1 (N13928, N13927);
not NOT1 (N13929, N13925);
or OR4 (N13930, N13929, N157, N10653, N10226);
or OR4 (N13931, N13921, N10999, N5785, N10717);
xor XOR2 (N13932, N13914, N7378);
or OR3 (N13933, N13924, N3902, N9140);
or OR4 (N13934, N13932, N4325, N9524, N12163);
xor XOR2 (N13935, N13916, N10506);
not NOT1 (N13936, N13926);
and AND2 (N13937, N13931, N2066);
xor XOR2 (N13938, N13937, N11778);
or OR3 (N13939, N13928, N3232, N4505);
not NOT1 (N13940, N13844);
nor NOR2 (N13941, N13930, N3149);
nand NAND4 (N13942, N13936, N1815, N3608, N12351);
buf BUF1 (N13943, N13938);
xor XOR2 (N13944, N13935, N12606);
or OR4 (N13945, N13944, N5133, N6173, N418);
not NOT1 (N13946, N13939);
buf BUF1 (N13947, N13922);
or OR3 (N13948, N13940, N2795, N3390);
not NOT1 (N13949, N13941);
nor NOR3 (N13950, N13945, N8266, N3828);
not NOT1 (N13951, N13948);
and AND2 (N13952, N13933, N9082);
nand NAND2 (N13953, N13947, N12878);
not NOT1 (N13954, N13942);
buf BUF1 (N13955, N13934);
or OR4 (N13956, N13955, N10949, N8249, N6451);
and AND4 (N13957, N13953, N10300, N7247, N539);
buf BUF1 (N13958, N13943);
not NOT1 (N13959, N13954);
buf BUF1 (N13960, N13958);
nor NOR4 (N13961, N13885, N2141, N4050, N4722);
nor NOR2 (N13962, N13952, N10649);
buf BUF1 (N13963, N13960);
xor XOR2 (N13964, N13962, N10301);
nand NAND4 (N13965, N13950, N13323, N3332, N7301);
not NOT1 (N13966, N13965);
not NOT1 (N13967, N13966);
and AND2 (N13968, N13946, N3584);
and AND4 (N13969, N13959, N9378, N775, N12591);
nand NAND4 (N13970, N13951, N3781, N1606, N5344);
nor NOR4 (N13971, N13969, N8981, N13568, N9110);
not NOT1 (N13972, N13968);
nor NOR2 (N13973, N13972, N13638);
not NOT1 (N13974, N13967);
and AND3 (N13975, N13961, N6487, N2063);
not NOT1 (N13976, N13949);
xor XOR2 (N13977, N13964, N8524);
nor NOR2 (N13978, N13970, N10870);
xor XOR2 (N13979, N13973, N9945);
not NOT1 (N13980, N13963);
not NOT1 (N13981, N13980);
buf BUF1 (N13982, N13979);
buf BUF1 (N13983, N13956);
or OR2 (N13984, N13977, N12661);
or OR2 (N13985, N13982, N8585);
or OR3 (N13986, N13984, N8187, N5264);
buf BUF1 (N13987, N13971);
nor NOR2 (N13988, N13987, N3004);
or OR2 (N13989, N13957, N11888);
or OR3 (N13990, N13988, N5291, N13517);
and AND3 (N13991, N13989, N11869, N9791);
nor NOR2 (N13992, N13990, N5146);
or OR3 (N13993, N13975, N3280, N5687);
nand NAND4 (N13994, N13978, N10673, N7393, N154);
xor XOR2 (N13995, N13993, N8983);
xor XOR2 (N13996, N13981, N1072);
xor XOR2 (N13997, N13974, N2850);
not NOT1 (N13998, N13997);
nor NOR3 (N13999, N13991, N7681, N6894);
xor XOR2 (N14000, N13998, N7912);
or OR2 (N14001, N13999, N11249);
nand NAND2 (N14002, N13986, N7493);
and AND3 (N14003, N14002, N500, N6609);
buf BUF1 (N14004, N13983);
buf BUF1 (N14005, N14003);
nor NOR2 (N14006, N13992, N12183);
nor NOR3 (N14007, N13976, N11675, N8507);
buf BUF1 (N14008, N14007);
nand NAND3 (N14009, N14008, N7492, N7534);
nand NAND3 (N14010, N13994, N10094, N10167);
not NOT1 (N14011, N14005);
nand NAND4 (N14012, N13985, N10408, N4779, N11024);
nand NAND2 (N14013, N14006, N109);
buf BUF1 (N14014, N14010);
and AND2 (N14015, N14001, N9634);
nand NAND3 (N14016, N14012, N9437, N6890);
or OR3 (N14017, N14000, N12451, N8054);
nand NAND2 (N14018, N14015, N6137);
buf BUF1 (N14019, N14013);
and AND4 (N14020, N13996, N8574, N5558, N687);
or OR2 (N14021, N14018, N12164);
nor NOR3 (N14022, N14020, N10829, N5004);
and AND4 (N14023, N14011, N8037, N53, N2964);
not NOT1 (N14024, N14021);
and AND3 (N14025, N14019, N11084, N5045);
nor NOR3 (N14026, N14017, N6834, N7318);
nor NOR3 (N14027, N14004, N4296, N11676);
xor XOR2 (N14028, N13995, N13923);
and AND3 (N14029, N14022, N6679, N9391);
nor NOR4 (N14030, N14014, N13586, N10317, N6931);
and AND2 (N14031, N14025, N1030);
and AND3 (N14032, N14027, N2338, N8882);
nand NAND2 (N14033, N14023, N13862);
buf BUF1 (N14034, N14032);
not NOT1 (N14035, N14029);
nand NAND4 (N14036, N14034, N654, N137, N4615);
and AND4 (N14037, N14028, N3878, N4500, N7292);
or OR3 (N14038, N14026, N12669, N5548);
or OR4 (N14039, N14035, N1979, N480, N5030);
nand NAND2 (N14040, N14038, N2018);
xor XOR2 (N14041, N14030, N490);
nand NAND4 (N14042, N14039, N661, N8998, N6264);
and AND4 (N14043, N14037, N1998, N5313, N7164);
and AND3 (N14044, N14036, N10679, N4914);
or OR3 (N14045, N14009, N7929, N10588);
and AND4 (N14046, N14045, N10731, N1600, N5871);
not NOT1 (N14047, N14046);
nand NAND2 (N14048, N14043, N9891);
xor XOR2 (N14049, N14047, N9223);
buf BUF1 (N14050, N14044);
not NOT1 (N14051, N14041);
nor NOR4 (N14052, N14051, N8808, N8768, N9661);
buf BUF1 (N14053, N14048);
nor NOR3 (N14054, N14050, N4147, N13857);
buf BUF1 (N14055, N14054);
not NOT1 (N14056, N14049);
or OR4 (N14057, N14040, N7444, N6426, N12539);
or OR2 (N14058, N14042, N8696);
buf BUF1 (N14059, N14057);
or OR2 (N14060, N14055, N11218);
nor NOR3 (N14061, N14060, N11455, N7957);
xor XOR2 (N14062, N14033, N11979);
xor XOR2 (N14063, N14016, N6680);
xor XOR2 (N14064, N14031, N2933);
and AND2 (N14065, N14056, N6194);
and AND2 (N14066, N14064, N11451);
buf BUF1 (N14067, N14063);
buf BUF1 (N14068, N14067);
and AND2 (N14069, N14058, N3125);
and AND2 (N14070, N14061, N386);
not NOT1 (N14071, N14068);
xor XOR2 (N14072, N14062, N12735);
nor NOR3 (N14073, N14069, N7225, N3274);
nor NOR3 (N14074, N14065, N7602, N8252);
nand NAND4 (N14075, N14066, N170, N9765, N13271);
not NOT1 (N14076, N14071);
buf BUF1 (N14077, N14024);
and AND4 (N14078, N14072, N12100, N1852, N10237);
and AND4 (N14079, N14078, N1629, N4819, N12214);
nor NOR4 (N14080, N14070, N9667, N2198, N180);
nor NOR3 (N14081, N14073, N10187, N7954);
nand NAND2 (N14082, N14076, N5394);
buf BUF1 (N14083, N14059);
xor XOR2 (N14084, N14083, N3092);
not NOT1 (N14085, N14081);
xor XOR2 (N14086, N14082, N8945);
nand NAND4 (N14087, N14053, N207, N5598, N10467);
xor XOR2 (N14088, N14084, N13107);
xor XOR2 (N14089, N14075, N9669);
buf BUF1 (N14090, N14088);
buf BUF1 (N14091, N14085);
and AND4 (N14092, N14087, N1013, N2285, N13680);
or OR4 (N14093, N14074, N6674, N8061, N864);
buf BUF1 (N14094, N14091);
nor NOR2 (N14095, N14080, N4001);
not NOT1 (N14096, N14093);
not NOT1 (N14097, N14089);
buf BUF1 (N14098, N14096);
not NOT1 (N14099, N14095);
nand NAND3 (N14100, N14098, N5589, N3690);
buf BUF1 (N14101, N14090);
nand NAND2 (N14102, N14099, N4709);
nand NAND3 (N14103, N14086, N2319, N11848);
nand NAND3 (N14104, N14103, N7670, N14022);
buf BUF1 (N14105, N14094);
and AND4 (N14106, N14077, N2586, N546, N13803);
xor XOR2 (N14107, N14102, N3742);
and AND2 (N14108, N14106, N12735);
and AND2 (N14109, N14100, N1216);
or OR3 (N14110, N14107, N3839, N753);
nand NAND3 (N14111, N14097, N941, N9181);
nor NOR2 (N14112, N14111, N7907);
or OR3 (N14113, N14112, N5623, N856);
xor XOR2 (N14114, N14105, N9244);
or OR4 (N14115, N14113, N586, N8563, N5637);
buf BUF1 (N14116, N14114);
nand NAND4 (N14117, N14079, N6820, N1477, N13812);
or OR3 (N14118, N14101, N5331, N8879);
and AND4 (N14119, N14118, N12371, N1795, N8150);
or OR4 (N14120, N14108, N1563, N2195, N9739);
not NOT1 (N14121, N14119);
nand NAND4 (N14122, N14121, N5858, N11808, N6877);
or OR4 (N14123, N14116, N3033, N4163, N11100);
not NOT1 (N14124, N14104);
or OR3 (N14125, N14124, N13603, N5295);
nor NOR3 (N14126, N14123, N2660, N10558);
buf BUF1 (N14127, N14115);
and AND2 (N14128, N14052, N8816);
and AND2 (N14129, N14128, N9328);
xor XOR2 (N14130, N14127, N10244);
and AND2 (N14131, N14126, N10663);
nand NAND4 (N14132, N14092, N2983, N9739, N3986);
xor XOR2 (N14133, N14110, N7872);
or OR2 (N14134, N14117, N245);
xor XOR2 (N14135, N14131, N9131);
nor NOR4 (N14136, N14133, N3324, N6637, N11099);
buf BUF1 (N14137, N14130);
xor XOR2 (N14138, N14134, N2670);
and AND3 (N14139, N14129, N8827, N7564);
buf BUF1 (N14140, N14138);
or OR3 (N14141, N14139, N4501, N3318);
and AND4 (N14142, N14122, N10560, N10715, N7756);
nor NOR3 (N14143, N14141, N1410, N6866);
nand NAND4 (N14144, N14135, N8436, N3937, N9506);
not NOT1 (N14145, N14136);
nand NAND2 (N14146, N14144, N5759);
buf BUF1 (N14147, N14145);
or OR2 (N14148, N14147, N4485);
buf BUF1 (N14149, N14146);
nor NOR4 (N14150, N14149, N5575, N8417, N11300);
not NOT1 (N14151, N14109);
nor NOR3 (N14152, N14137, N6188, N12585);
nor NOR3 (N14153, N14148, N2764, N5520);
nand NAND4 (N14154, N14153, N9731, N9550, N9441);
xor XOR2 (N14155, N14143, N7502);
not NOT1 (N14156, N14132);
and AND4 (N14157, N14154, N931, N2552, N3853);
xor XOR2 (N14158, N14142, N10837);
and AND3 (N14159, N14140, N3739, N6629);
or OR3 (N14160, N14152, N868, N7383);
or OR2 (N14161, N14151, N9979);
buf BUF1 (N14162, N14155);
nand NAND2 (N14163, N14125, N10671);
xor XOR2 (N14164, N14156, N13366);
buf BUF1 (N14165, N14162);
and AND3 (N14166, N14150, N7174, N12682);
nand NAND2 (N14167, N14160, N2764);
and AND4 (N14168, N14163, N1810, N11996, N12842);
or OR4 (N14169, N14159, N8350, N11333, N2216);
nand NAND2 (N14170, N14158, N3592);
nor NOR3 (N14171, N14167, N12997, N9743);
not NOT1 (N14172, N14166);
not NOT1 (N14173, N14165);
or OR4 (N14174, N14170, N13658, N8169, N2140);
nor NOR2 (N14175, N14174, N3410);
nand NAND2 (N14176, N14171, N12854);
xor XOR2 (N14177, N14172, N9321);
buf BUF1 (N14178, N14120);
nand NAND2 (N14179, N14177, N6666);
xor XOR2 (N14180, N14175, N4913);
not NOT1 (N14181, N14176);
not NOT1 (N14182, N14173);
nand NAND2 (N14183, N14178, N6127);
nand NAND4 (N14184, N14164, N7898, N4584, N8101);
or OR4 (N14185, N14168, N11269, N8844, N12887);
nor NOR4 (N14186, N14180, N2341, N4715, N12270);
not NOT1 (N14187, N14179);
and AND2 (N14188, N14185, N7052);
and AND3 (N14189, N14186, N1732, N4405);
or OR3 (N14190, N14181, N7050, N1349);
buf BUF1 (N14191, N14190);
nand NAND2 (N14192, N14157, N8595);
or OR4 (N14193, N14184, N5644, N9127, N13212);
nor NOR3 (N14194, N14189, N14148, N7260);
not NOT1 (N14195, N14188);
not NOT1 (N14196, N14187);
and AND3 (N14197, N14183, N13031, N4107);
or OR3 (N14198, N14192, N10499, N2699);
and AND4 (N14199, N14193, N780, N13731, N13900);
xor XOR2 (N14200, N14194, N32);
and AND3 (N14201, N14198, N804, N865);
not NOT1 (N14202, N14161);
or OR3 (N14203, N14182, N10715, N8988);
buf BUF1 (N14204, N14201);
or OR2 (N14205, N14200, N5593);
nand NAND4 (N14206, N14196, N7375, N925, N12463);
and AND3 (N14207, N14169, N6137, N362);
nor NOR4 (N14208, N14206, N4045, N7235, N11326);
xor XOR2 (N14209, N14207, N2699);
xor XOR2 (N14210, N14197, N951);
not NOT1 (N14211, N14203);
buf BUF1 (N14212, N14210);
nand NAND3 (N14213, N14212, N12656, N3580);
buf BUF1 (N14214, N14209);
xor XOR2 (N14215, N14214, N11561);
nand NAND3 (N14216, N14215, N12985, N5206);
nor NOR3 (N14217, N14208, N587, N4353);
and AND4 (N14218, N14195, N4509, N10198, N3997);
and AND3 (N14219, N14216, N8037, N6076);
buf BUF1 (N14220, N14218);
not NOT1 (N14221, N14199);
or OR3 (N14222, N14202, N12056, N2988);
nand NAND3 (N14223, N14191, N8695, N4251);
nand NAND2 (N14224, N14219, N7762);
and AND3 (N14225, N14224, N271, N4086);
nor NOR3 (N14226, N14204, N8222, N147);
nand NAND2 (N14227, N14222, N10300);
nand NAND3 (N14228, N14213, N11794, N7702);
nor NOR4 (N14229, N14217, N6206, N13946, N5340);
xor XOR2 (N14230, N14223, N11350);
xor XOR2 (N14231, N14230, N3392);
and AND3 (N14232, N14227, N2352, N8197);
or OR2 (N14233, N14226, N221);
or OR4 (N14234, N14211, N6816, N11254, N10537);
xor XOR2 (N14235, N14228, N7064);
nand NAND3 (N14236, N14221, N11857, N873);
or OR3 (N14237, N14231, N13868, N1911);
nor NOR4 (N14238, N14236, N938, N10225, N6469);
nand NAND3 (N14239, N14234, N4196, N11610);
and AND4 (N14240, N14232, N11204, N9164, N216);
not NOT1 (N14241, N14240);
or OR3 (N14242, N14225, N10203, N1218);
nor NOR2 (N14243, N14239, N4787);
xor XOR2 (N14244, N14229, N2559);
nand NAND4 (N14245, N14205, N3044, N7273, N13665);
and AND4 (N14246, N14235, N5650, N2738, N4075);
nand NAND3 (N14247, N14220, N10663, N7607);
not NOT1 (N14248, N14238);
nand NAND4 (N14249, N14237, N8341, N12976, N13103);
xor XOR2 (N14250, N14243, N7762);
nor NOR4 (N14251, N14233, N9831, N14104, N12797);
xor XOR2 (N14252, N14248, N4572);
xor XOR2 (N14253, N14252, N8939);
xor XOR2 (N14254, N14249, N5473);
xor XOR2 (N14255, N14250, N2502);
nor NOR2 (N14256, N14241, N10119);
and AND3 (N14257, N14245, N1271, N783);
nor NOR4 (N14258, N14246, N3435, N6812, N6763);
buf BUF1 (N14259, N14254);
or OR3 (N14260, N14255, N1086, N5615);
buf BUF1 (N14261, N14242);
buf BUF1 (N14262, N14247);
nand NAND2 (N14263, N14260, N6782);
not NOT1 (N14264, N14253);
nand NAND3 (N14265, N14257, N7137, N4371);
not NOT1 (N14266, N14259);
xor XOR2 (N14267, N14261, N11179);
nor NOR4 (N14268, N14251, N2371, N8297, N13675);
or OR2 (N14269, N14263, N7113);
buf BUF1 (N14270, N14256);
xor XOR2 (N14271, N14265, N1039);
not NOT1 (N14272, N14270);
nor NOR3 (N14273, N14269, N5718, N7038);
or OR3 (N14274, N14268, N5065, N1155);
buf BUF1 (N14275, N14244);
xor XOR2 (N14276, N14267, N2750);
and AND2 (N14277, N14272, N6381);
xor XOR2 (N14278, N14274, N2637);
buf BUF1 (N14279, N14262);
nand NAND4 (N14280, N14264, N10287, N2693, N9406);
or OR4 (N14281, N14273, N3116, N5724, N11174);
nor NOR4 (N14282, N14271, N8610, N1204, N12431);
nand NAND2 (N14283, N14266, N7720);
nand NAND4 (N14284, N14278, N5683, N3649, N2464);
or OR2 (N14285, N14279, N6513);
nand NAND3 (N14286, N14275, N13670, N5585);
buf BUF1 (N14287, N14284);
buf BUF1 (N14288, N14258);
not NOT1 (N14289, N14282);
buf BUF1 (N14290, N14288);
nand NAND4 (N14291, N14283, N926, N11630, N493);
and AND2 (N14292, N14291, N2518);
or OR2 (N14293, N14287, N2774);
or OR3 (N14294, N14289, N1661, N4426);
buf BUF1 (N14295, N14292);
and AND3 (N14296, N14286, N8636, N7889);
buf BUF1 (N14297, N14295);
buf BUF1 (N14298, N14276);
buf BUF1 (N14299, N14290);
nor NOR4 (N14300, N14296, N8335, N1838, N302);
nand NAND3 (N14301, N14277, N4523, N12114);
buf BUF1 (N14302, N14285);
nand NAND3 (N14303, N14297, N7777, N11436);
nand NAND3 (N14304, N14300, N5625, N7656);
nor NOR4 (N14305, N14281, N9233, N4078, N679);
not NOT1 (N14306, N14299);
xor XOR2 (N14307, N14305, N13689);
nor NOR4 (N14308, N14307, N5444, N3366, N2482);
nand NAND4 (N14309, N14304, N3543, N1185, N3230);
buf BUF1 (N14310, N14306);
nor NOR2 (N14311, N14303, N12772);
or OR3 (N14312, N14309, N687, N8689);
and AND2 (N14313, N14310, N51);
nor NOR4 (N14314, N14280, N12513, N3759, N10642);
buf BUF1 (N14315, N14312);
nand NAND4 (N14316, N14315, N8996, N14058, N6019);
and AND3 (N14317, N14311, N13278, N7765);
and AND3 (N14318, N14317, N8799, N12412);
nand NAND3 (N14319, N14298, N6259, N4223);
or OR2 (N14320, N14302, N11423);
not NOT1 (N14321, N14320);
xor XOR2 (N14322, N14308, N9805);
buf BUF1 (N14323, N14293);
nand NAND4 (N14324, N14322, N171, N3459, N6124);
and AND2 (N14325, N14319, N6181);
xor XOR2 (N14326, N14321, N5909);
nand NAND4 (N14327, N14294, N12582, N2015, N7234);
nand NAND4 (N14328, N14318, N1669, N10763, N13019);
buf BUF1 (N14329, N14327);
or OR3 (N14330, N14324, N8868, N9190);
buf BUF1 (N14331, N14326);
not NOT1 (N14332, N14329);
nand NAND4 (N14333, N14330, N2760, N2980, N5544);
nor NOR3 (N14334, N14328, N149, N7493);
not NOT1 (N14335, N14333);
not NOT1 (N14336, N14301);
and AND2 (N14337, N14332, N645);
buf BUF1 (N14338, N14323);
nor NOR4 (N14339, N14316, N8497, N8684, N3747);
not NOT1 (N14340, N14336);
xor XOR2 (N14341, N14338, N10834);
nand NAND2 (N14342, N14339, N12200);
buf BUF1 (N14343, N14341);
nor NOR4 (N14344, N14343, N3379, N4238, N9472);
xor XOR2 (N14345, N14334, N315);
xor XOR2 (N14346, N14314, N7259);
nand NAND2 (N14347, N14345, N7105);
and AND3 (N14348, N14337, N5163, N7147);
xor XOR2 (N14349, N14325, N13271);
and AND2 (N14350, N14346, N1734);
nor NOR3 (N14351, N14349, N1670, N11050);
xor XOR2 (N14352, N14344, N5018);
xor XOR2 (N14353, N14347, N9600);
or OR3 (N14354, N14313, N13849, N10010);
not NOT1 (N14355, N14348);
not NOT1 (N14356, N14351);
nor NOR2 (N14357, N14342, N13989);
or OR4 (N14358, N14352, N10351, N11493, N5857);
not NOT1 (N14359, N14331);
and AND3 (N14360, N14356, N1719, N8909);
nor NOR2 (N14361, N14358, N4185);
or OR4 (N14362, N14335, N12815, N1386, N5529);
nor NOR4 (N14363, N14353, N3283, N8482, N10124);
buf BUF1 (N14364, N14362);
nand NAND2 (N14365, N14355, N10474);
and AND2 (N14366, N14365, N12529);
nor NOR2 (N14367, N14359, N3333);
or OR3 (N14368, N14366, N8836, N5912);
xor XOR2 (N14369, N14364, N13198);
nand NAND3 (N14370, N14354, N105, N7976);
or OR2 (N14371, N14340, N4225);
xor XOR2 (N14372, N14369, N2946);
and AND3 (N14373, N14368, N5738, N2545);
xor XOR2 (N14374, N14370, N7564);
nor NOR4 (N14375, N14350, N1138, N11784, N8935);
nor NOR2 (N14376, N14367, N9467);
or OR2 (N14377, N14376, N1873);
and AND4 (N14378, N14372, N8955, N14239, N2639);
or OR2 (N14379, N14371, N12784);
xor XOR2 (N14380, N14361, N12148);
or OR4 (N14381, N14375, N3992, N13795, N12365);
and AND2 (N14382, N14377, N1176);
or OR2 (N14383, N14357, N10698);
not NOT1 (N14384, N14380);
buf BUF1 (N14385, N14379);
buf BUF1 (N14386, N14373);
or OR3 (N14387, N14363, N1477, N6377);
not NOT1 (N14388, N14378);
or OR2 (N14389, N14385, N8776);
buf BUF1 (N14390, N14382);
and AND4 (N14391, N14384, N7226, N3637, N11575);
xor XOR2 (N14392, N14386, N7689);
buf BUF1 (N14393, N14383);
nand NAND4 (N14394, N14360, N13148, N2118, N816);
nor NOR4 (N14395, N14390, N13680, N13873, N4171);
or OR4 (N14396, N14392, N3670, N12821, N3290);
xor XOR2 (N14397, N14389, N4121);
buf BUF1 (N14398, N14397);
and AND2 (N14399, N14394, N10634);
nor NOR2 (N14400, N14393, N5304);
nand NAND2 (N14401, N14388, N11077);
buf BUF1 (N14402, N14374);
and AND2 (N14403, N14387, N12041);
nand NAND3 (N14404, N14403, N13664, N9313);
not NOT1 (N14405, N14381);
buf BUF1 (N14406, N14399);
not NOT1 (N14407, N14398);
not NOT1 (N14408, N14404);
buf BUF1 (N14409, N14408);
buf BUF1 (N14410, N14400);
buf BUF1 (N14411, N14391);
not NOT1 (N14412, N14409);
nand NAND2 (N14413, N14411, N8589);
nand NAND3 (N14414, N14402, N6502, N7227);
nand NAND3 (N14415, N14407, N4432, N9402);
buf BUF1 (N14416, N14410);
and AND4 (N14417, N14415, N305, N6567, N13075);
nand NAND4 (N14418, N14395, N2279, N2220, N7344);
nand NAND3 (N14419, N14401, N2129, N8999);
and AND4 (N14420, N14414, N7758, N579, N2907);
and AND4 (N14421, N14412, N5416, N3414, N12955);
buf BUF1 (N14422, N14421);
or OR3 (N14423, N14419, N4705, N10031);
not NOT1 (N14424, N14418);
buf BUF1 (N14425, N14396);
not NOT1 (N14426, N14425);
buf BUF1 (N14427, N14424);
nor NOR4 (N14428, N14417, N9462, N12870, N8499);
and AND4 (N14429, N14427, N9643, N9040, N5457);
nor NOR2 (N14430, N14416, N6867);
and AND2 (N14431, N14406, N14223);
buf BUF1 (N14432, N14428);
buf BUF1 (N14433, N14426);
nor NOR4 (N14434, N14405, N11026, N4224, N11863);
not NOT1 (N14435, N14430);
nor NOR4 (N14436, N14429, N8642, N12636, N531);
not NOT1 (N14437, N14434);
xor XOR2 (N14438, N14436, N971);
buf BUF1 (N14439, N14433);
not NOT1 (N14440, N14423);
and AND4 (N14441, N14435, N6531, N6612, N8854);
nor NOR4 (N14442, N14437, N4305, N2332, N5116);
nor NOR4 (N14443, N14413, N5495, N4785, N6381);
nor NOR4 (N14444, N14431, N672, N3851, N4044);
xor XOR2 (N14445, N14444, N6882);
and AND4 (N14446, N14443, N9148, N8491, N10409);
not NOT1 (N14447, N14446);
buf BUF1 (N14448, N14440);
not NOT1 (N14449, N14438);
buf BUF1 (N14450, N14422);
nand NAND3 (N14451, N14420, N5931, N6841);
buf BUF1 (N14452, N14448);
or OR3 (N14453, N14441, N13994, N3451);
nand NAND4 (N14454, N14452, N6974, N10028, N10180);
buf BUF1 (N14455, N14442);
not NOT1 (N14456, N14432);
nand NAND4 (N14457, N14451, N4929, N3237, N2920);
xor XOR2 (N14458, N14456, N5152);
xor XOR2 (N14459, N14450, N4859);
nor NOR3 (N14460, N14449, N3057, N4847);
not NOT1 (N14461, N14454);
xor XOR2 (N14462, N14458, N3308);
not NOT1 (N14463, N14460);
xor XOR2 (N14464, N14462, N13490);
xor XOR2 (N14465, N14459, N5350);
nand NAND4 (N14466, N14439, N3691, N13208, N8321);
nand NAND4 (N14467, N14461, N952, N14010, N12055);
or OR2 (N14468, N14445, N14357);
or OR3 (N14469, N14465, N11030, N12229);
or OR2 (N14470, N14453, N5316);
buf BUF1 (N14471, N14457);
or OR3 (N14472, N14463, N3111, N8852);
or OR3 (N14473, N14469, N2297, N5392);
nand NAND3 (N14474, N14455, N5909, N10067);
or OR3 (N14475, N14447, N13897, N5947);
not NOT1 (N14476, N14467);
or OR3 (N14477, N14466, N1743, N3368);
nand NAND3 (N14478, N14473, N9442, N10078);
buf BUF1 (N14479, N14471);
or OR2 (N14480, N14478, N2647);
or OR2 (N14481, N14464, N6324);
and AND4 (N14482, N14472, N9646, N12133, N5494);
or OR2 (N14483, N14474, N8373);
or OR3 (N14484, N14480, N6007, N9662);
xor XOR2 (N14485, N14475, N9419);
not NOT1 (N14486, N14482);
not NOT1 (N14487, N14484);
not NOT1 (N14488, N14483);
nand NAND3 (N14489, N14479, N1754, N14475);
xor XOR2 (N14490, N14486, N10828);
or OR4 (N14491, N14489, N14392, N3219, N6585);
buf BUF1 (N14492, N14468);
not NOT1 (N14493, N14481);
nor NOR3 (N14494, N14490, N10401, N790);
not NOT1 (N14495, N14488);
buf BUF1 (N14496, N14492);
nand NAND3 (N14497, N14494, N8715, N5538);
and AND4 (N14498, N14493, N4363, N452, N2286);
xor XOR2 (N14499, N14497, N3213);
buf BUF1 (N14500, N14470);
buf BUF1 (N14501, N14500);
buf BUF1 (N14502, N14501);
not NOT1 (N14503, N14499);
and AND4 (N14504, N14487, N12522, N4855, N7668);
buf BUF1 (N14505, N14496);
and AND4 (N14506, N14477, N1526, N12344, N9206);
or OR4 (N14507, N14498, N7037, N10178, N9425);
and AND4 (N14508, N14505, N13482, N2047, N12518);
buf BUF1 (N14509, N14502);
nor NOR4 (N14510, N14476, N4643, N2540, N7822);
nor NOR3 (N14511, N14506, N12547, N13459);
nand NAND2 (N14512, N14504, N14109);
xor XOR2 (N14513, N14491, N10887);
buf BUF1 (N14514, N14485);
nor NOR4 (N14515, N14510, N6866, N2349, N12248);
buf BUF1 (N14516, N14513);
or OR4 (N14517, N14507, N10458, N13048, N14057);
nor NOR4 (N14518, N14495, N14236, N6038, N1744);
buf BUF1 (N14519, N14518);
and AND2 (N14520, N14514, N8232);
not NOT1 (N14521, N14503);
or OR4 (N14522, N14515, N2531, N11584, N934);
not NOT1 (N14523, N14517);
or OR3 (N14524, N14508, N796, N14500);
nand NAND3 (N14525, N14509, N6941, N7470);
nor NOR2 (N14526, N14519, N4239);
nand NAND4 (N14527, N14525, N5332, N10030, N8704);
and AND2 (N14528, N14526, N13486);
buf BUF1 (N14529, N14516);
buf BUF1 (N14530, N14523);
nor NOR4 (N14531, N14511, N4541, N4964, N11709);
nor NOR2 (N14532, N14520, N10862);
and AND2 (N14533, N14521, N8688);
xor XOR2 (N14534, N14531, N10218);
xor XOR2 (N14535, N14527, N7427);
nor NOR4 (N14536, N14535, N8566, N1977, N6619);
not NOT1 (N14537, N14533);
nor NOR4 (N14538, N14524, N131, N9054, N3940);
xor XOR2 (N14539, N14528, N5322);
or OR3 (N14540, N14534, N4061, N13112);
nand NAND4 (N14541, N14512, N5052, N5994, N4997);
not NOT1 (N14542, N14537);
nand NAND4 (N14543, N14542, N7785, N2511, N2076);
and AND3 (N14544, N14536, N12742, N8848);
xor XOR2 (N14545, N14538, N376);
buf BUF1 (N14546, N14541);
nand NAND3 (N14547, N14532, N2327, N7678);
nand NAND3 (N14548, N14547, N13179, N4303);
and AND4 (N14549, N14545, N7098, N13690, N1398);
not NOT1 (N14550, N14529);
not NOT1 (N14551, N14544);
not NOT1 (N14552, N14543);
buf BUF1 (N14553, N14522);
xor XOR2 (N14554, N14550, N10396);
nand NAND4 (N14555, N14549, N8357, N11373, N1841);
not NOT1 (N14556, N14554);
buf BUF1 (N14557, N14546);
xor XOR2 (N14558, N14539, N14385);
xor XOR2 (N14559, N14548, N6257);
and AND3 (N14560, N14558, N10441, N6223);
nand NAND3 (N14561, N14556, N9217, N9109);
or OR2 (N14562, N14553, N3622);
nand NAND3 (N14563, N14540, N348, N9445);
nor NOR2 (N14564, N14562, N4421);
xor XOR2 (N14565, N14563, N12086);
buf BUF1 (N14566, N14555);
nor NOR3 (N14567, N14559, N12377, N3154);
and AND3 (N14568, N14565, N6946, N2285);
and AND2 (N14569, N14557, N3879);
or OR3 (N14570, N14560, N3429, N14278);
or OR3 (N14571, N14530, N11019, N4293);
or OR3 (N14572, N14551, N4293, N39);
nor NOR3 (N14573, N14564, N12180, N913);
buf BUF1 (N14574, N14552);
nor NOR2 (N14575, N14568, N8908);
and AND4 (N14576, N14572, N8464, N13728, N7221);
not NOT1 (N14577, N14570);
or OR3 (N14578, N14561, N10476, N4028);
xor XOR2 (N14579, N14566, N8010);
or OR2 (N14580, N14567, N7134);
nand NAND2 (N14581, N14569, N1351);
and AND3 (N14582, N14579, N2046, N209);
or OR4 (N14583, N14580, N4048, N9465, N6615);
xor XOR2 (N14584, N14573, N4376);
buf BUF1 (N14585, N14576);
or OR2 (N14586, N14575, N6790);
and AND2 (N14587, N14578, N2651);
xor XOR2 (N14588, N14571, N12696);
or OR4 (N14589, N14584, N1896, N14574, N7016);
not NOT1 (N14590, N8035);
not NOT1 (N14591, N14590);
or OR4 (N14592, N14581, N703, N2631, N1004);
not NOT1 (N14593, N14588);
and AND3 (N14594, N14593, N7425, N1070);
and AND3 (N14595, N14592, N6286, N233);
xor XOR2 (N14596, N14587, N7363);
xor XOR2 (N14597, N14585, N4237);
nand NAND3 (N14598, N14582, N4594, N12294);
or OR2 (N14599, N14598, N4181);
nand NAND2 (N14600, N14591, N13810);
or OR4 (N14601, N14599, N11058, N14260, N176);
xor XOR2 (N14602, N14596, N2397);
nor NOR3 (N14603, N14600, N8659, N1954);
not NOT1 (N14604, N14577);
nor NOR2 (N14605, N14595, N1044);
buf BUF1 (N14606, N14594);
and AND3 (N14607, N14602, N13355, N5991);
not NOT1 (N14608, N14603);
or OR2 (N14609, N14589, N3775);
buf BUF1 (N14610, N14605);
xor XOR2 (N14611, N14583, N9376);
xor XOR2 (N14612, N14604, N885);
xor XOR2 (N14613, N14607, N9986);
nor NOR2 (N14614, N14611, N6089);
nor NOR3 (N14615, N14586, N6501, N3550);
not NOT1 (N14616, N14597);
nor NOR3 (N14617, N14608, N5322, N7550);
xor XOR2 (N14618, N14612, N5143);
or OR2 (N14619, N14606, N3859);
nand NAND2 (N14620, N14618, N1242);
buf BUF1 (N14621, N14620);
xor XOR2 (N14622, N14613, N8344);
nand NAND2 (N14623, N14601, N7111);
not NOT1 (N14624, N14619);
not NOT1 (N14625, N14610);
xor XOR2 (N14626, N14615, N4679);
not NOT1 (N14627, N14614);
nor NOR3 (N14628, N14626, N12439, N3065);
buf BUF1 (N14629, N14624);
and AND4 (N14630, N14628, N1213, N3926, N6273);
nand NAND3 (N14631, N14622, N4514, N12925);
or OR2 (N14632, N14631, N9087);
nand NAND4 (N14633, N14617, N2595, N5825, N6887);
xor XOR2 (N14634, N14632, N4980);
and AND2 (N14635, N14609, N284);
or OR3 (N14636, N14634, N8491, N10479);
nand NAND3 (N14637, N14630, N11679, N9867);
nor NOR2 (N14638, N14623, N9709);
xor XOR2 (N14639, N14637, N8426);
and AND2 (N14640, N14638, N7437);
and AND2 (N14641, N14625, N12395);
nand NAND4 (N14642, N14616, N10649, N10819, N1384);
buf BUF1 (N14643, N14636);
xor XOR2 (N14644, N14639, N11821);
or OR4 (N14645, N14640, N13005, N1497, N12070);
nor NOR3 (N14646, N14643, N14257, N8971);
xor XOR2 (N14647, N14633, N8548);
xor XOR2 (N14648, N14645, N7368);
xor XOR2 (N14649, N14647, N1531);
buf BUF1 (N14650, N14648);
or OR4 (N14651, N14635, N6947, N1184, N7007);
nor NOR4 (N14652, N14642, N666, N13539, N14445);
nand NAND3 (N14653, N14649, N1427, N9971);
nor NOR3 (N14654, N14650, N3389, N2610);
nand NAND4 (N14655, N14652, N6722, N1182, N9399);
not NOT1 (N14656, N14627);
xor XOR2 (N14657, N14655, N12229);
nor NOR4 (N14658, N14657, N14218, N1459, N2168);
buf BUF1 (N14659, N14656);
nor NOR2 (N14660, N14646, N6972);
nand NAND4 (N14661, N14653, N2897, N10123, N9795);
buf BUF1 (N14662, N14654);
or OR3 (N14663, N14660, N7391, N872);
xor XOR2 (N14664, N14651, N4611);
nor NOR4 (N14665, N14629, N9094, N9268, N3340);
xor XOR2 (N14666, N14665, N6044);
buf BUF1 (N14667, N14662);
not NOT1 (N14668, N14658);
xor XOR2 (N14669, N14664, N789);
buf BUF1 (N14670, N14666);
nor NOR4 (N14671, N14641, N11248, N2780, N3498);
buf BUF1 (N14672, N14667);
nand NAND4 (N14673, N14659, N5656, N12278, N6149);
nand NAND3 (N14674, N14671, N9548, N174);
nor NOR3 (N14675, N14669, N1528, N14101);
and AND2 (N14676, N14621, N699);
or OR4 (N14677, N14644, N11869, N8572, N14628);
not NOT1 (N14678, N14674);
nor NOR3 (N14679, N14678, N11759, N12423);
nand NAND3 (N14680, N14668, N3520, N10017);
not NOT1 (N14681, N14676);
or OR4 (N14682, N14675, N12994, N2832, N6116);
nor NOR3 (N14683, N14682, N4046, N1293);
not NOT1 (N14684, N14673);
xor XOR2 (N14685, N14679, N10970);
and AND4 (N14686, N14684, N11320, N14182, N1330);
buf BUF1 (N14687, N14686);
and AND2 (N14688, N14687, N443);
buf BUF1 (N14689, N14685);
buf BUF1 (N14690, N14689);
nor NOR4 (N14691, N14672, N7561, N2015, N13789);
nand NAND2 (N14692, N14691, N296);
and AND3 (N14693, N14670, N11706, N14597);
not NOT1 (N14694, N14677);
xor XOR2 (N14695, N14683, N13723);
nor NOR3 (N14696, N14663, N752, N1332);
nand NAND3 (N14697, N14688, N10835, N8507);
nand NAND2 (N14698, N14695, N13939);
xor XOR2 (N14699, N14693, N1798);
nand NAND4 (N14700, N14696, N3854, N9012, N7047);
nor NOR2 (N14701, N14680, N9460);
not NOT1 (N14702, N14681);
xor XOR2 (N14703, N14697, N9304);
nand NAND3 (N14704, N14699, N7331, N7617);
buf BUF1 (N14705, N14690);
or OR3 (N14706, N14703, N8311, N12439);
nand NAND3 (N14707, N14701, N3198, N2097);
nor NOR4 (N14708, N14700, N11261, N4606, N14119);
not NOT1 (N14709, N14661);
nand NAND3 (N14710, N14707, N3327, N522);
nor NOR2 (N14711, N14702, N4240);
buf BUF1 (N14712, N14706);
and AND3 (N14713, N14709, N8773, N7139);
or OR2 (N14714, N14694, N1885);
or OR4 (N14715, N14713, N10089, N5419, N11427);
and AND3 (N14716, N14704, N4174, N14208);
not NOT1 (N14717, N14714);
and AND4 (N14718, N14710, N245, N9841, N9811);
nor NOR2 (N14719, N14712, N13481);
or OR4 (N14720, N14705, N10988, N4039, N1793);
not NOT1 (N14721, N14717);
not NOT1 (N14722, N14716);
buf BUF1 (N14723, N14721);
nand NAND3 (N14724, N14720, N3751, N9642);
buf BUF1 (N14725, N14698);
xor XOR2 (N14726, N14715, N1038);
nand NAND2 (N14727, N14708, N1617);
buf BUF1 (N14728, N14727);
and AND3 (N14729, N14725, N7450, N14358);
or OR3 (N14730, N14724, N11294, N9541);
not NOT1 (N14731, N14711);
xor XOR2 (N14732, N14728, N3128);
nor NOR3 (N14733, N14726, N10692, N4146);
and AND2 (N14734, N14729, N12789);
not NOT1 (N14735, N14734);
not NOT1 (N14736, N14732);
xor XOR2 (N14737, N14719, N889);
nor NOR4 (N14738, N14733, N9524, N13347, N2136);
and AND4 (N14739, N14723, N4912, N10847, N5494);
buf BUF1 (N14740, N14722);
and AND3 (N14741, N14718, N14740, N7333);
not NOT1 (N14742, N8970);
not NOT1 (N14743, N14739);
buf BUF1 (N14744, N14731);
nand NAND3 (N14745, N14744, N7465, N262);
buf BUF1 (N14746, N14737);
nor NOR2 (N14747, N14738, N5540);
nor NOR4 (N14748, N14745, N10231, N1060, N10015);
xor XOR2 (N14749, N14736, N7858);
not NOT1 (N14750, N14749);
nand NAND3 (N14751, N14747, N13717, N3949);
xor XOR2 (N14752, N14748, N6722);
nor NOR3 (N14753, N14735, N14138, N1020);
not NOT1 (N14754, N14753);
xor XOR2 (N14755, N14742, N7349);
not NOT1 (N14756, N14755);
or OR4 (N14757, N14743, N1957, N6764, N10427);
and AND3 (N14758, N14757, N4629, N7421);
nor NOR3 (N14759, N14751, N14440, N12089);
xor XOR2 (N14760, N14741, N11936);
buf BUF1 (N14761, N14746);
buf BUF1 (N14762, N14692);
and AND3 (N14763, N14761, N9651, N2492);
or OR4 (N14764, N14750, N12908, N10260, N8768);
nand NAND3 (N14765, N14752, N5852, N9931);
xor XOR2 (N14766, N14762, N3564);
or OR4 (N14767, N14758, N5814, N3813, N9626);
xor XOR2 (N14768, N14759, N11361);
or OR4 (N14769, N14768, N6319, N14754, N5363);
nor NOR3 (N14770, N567, N4125, N2417);
not NOT1 (N14771, N14730);
not NOT1 (N14772, N14760);
xor XOR2 (N14773, N14767, N11483);
xor XOR2 (N14774, N14766, N786);
not NOT1 (N14775, N14763);
not NOT1 (N14776, N14772);
buf BUF1 (N14777, N14756);
nand NAND2 (N14778, N14771, N300);
xor XOR2 (N14779, N14774, N3665);
nor NOR3 (N14780, N14777, N2070, N1181);
xor XOR2 (N14781, N14770, N682);
not NOT1 (N14782, N14775);
not NOT1 (N14783, N14773);
xor XOR2 (N14784, N14769, N10787);
or OR4 (N14785, N14780, N1135, N7794, N9497);
nor NOR3 (N14786, N14782, N12488, N7820);
not NOT1 (N14787, N14781);
not NOT1 (N14788, N14783);
xor XOR2 (N14789, N14788, N11434);
nand NAND3 (N14790, N14787, N9455, N8248);
nand NAND3 (N14791, N14786, N8620, N5754);
not NOT1 (N14792, N14765);
and AND4 (N14793, N14778, N6, N8789, N1946);
or OR4 (N14794, N14785, N9351, N10426, N6695);
nand NAND3 (N14795, N14790, N3766, N6980);
and AND2 (N14796, N14791, N954);
and AND3 (N14797, N14789, N14121, N11548);
and AND3 (N14798, N14797, N8984, N14434);
and AND2 (N14799, N14795, N1596);
and AND4 (N14800, N14796, N1365, N6703, N6592);
and AND2 (N14801, N14776, N9826);
nand NAND4 (N14802, N14793, N3658, N2390, N4883);
xor XOR2 (N14803, N14798, N2424);
xor XOR2 (N14804, N14784, N8576);
nand NAND2 (N14805, N14804, N13324);
nand NAND4 (N14806, N14805, N8508, N11340, N13082);
buf BUF1 (N14807, N14802);
buf BUF1 (N14808, N14779);
or OR3 (N14809, N14801, N476, N3983);
xor XOR2 (N14810, N14806, N8822);
and AND2 (N14811, N14803, N6520);
not NOT1 (N14812, N14764);
nand NAND4 (N14813, N14808, N13941, N13219, N8934);
or OR2 (N14814, N14800, N6848);
xor XOR2 (N14815, N14810, N6467);
not NOT1 (N14816, N14799);
nor NOR2 (N14817, N14813, N12516);
xor XOR2 (N14818, N14807, N5229);
not NOT1 (N14819, N14817);
buf BUF1 (N14820, N14792);
and AND3 (N14821, N14814, N7364, N4612);
buf BUF1 (N14822, N14821);
xor XOR2 (N14823, N14820, N12143);
xor XOR2 (N14824, N14819, N11664);
not NOT1 (N14825, N14811);
or OR3 (N14826, N14825, N1872, N4978);
and AND2 (N14827, N14818, N12238);
nor NOR2 (N14828, N14816, N12600);
nor NOR4 (N14829, N14826, N4676, N10277, N956);
nand NAND2 (N14830, N14824, N1903);
buf BUF1 (N14831, N14815);
not NOT1 (N14832, N14809);
nand NAND4 (N14833, N14794, N7837, N13407, N4301);
nand NAND3 (N14834, N14832, N1135, N12059);
xor XOR2 (N14835, N14830, N8074);
nor NOR2 (N14836, N14834, N6180);
or OR4 (N14837, N14827, N7833, N6376, N9512);
or OR4 (N14838, N14812, N2698, N7730, N6880);
or OR2 (N14839, N14828, N9197);
nand NAND2 (N14840, N14837, N6682);
or OR2 (N14841, N14839, N7801);
nand NAND4 (N14842, N14835, N2517, N13921, N1057);
xor XOR2 (N14843, N14836, N5854);
and AND3 (N14844, N14831, N9081, N1301);
nand NAND4 (N14845, N14842, N1319, N7993, N7903);
nand NAND4 (N14846, N14833, N11191, N2051, N620);
and AND2 (N14847, N14846, N3356);
not NOT1 (N14848, N14847);
nor NOR3 (N14849, N14829, N6160, N2397);
nor NOR2 (N14850, N14848, N8976);
nand NAND2 (N14851, N14843, N3796);
nor NOR2 (N14852, N14840, N1936);
and AND3 (N14853, N14841, N4256, N13987);
buf BUF1 (N14854, N14823);
xor XOR2 (N14855, N14849, N12451);
not NOT1 (N14856, N14855);
nand NAND3 (N14857, N14838, N2939, N145);
not NOT1 (N14858, N14853);
or OR4 (N14859, N14851, N7145, N6996, N8042);
nor NOR2 (N14860, N14854, N10540);
and AND2 (N14861, N14845, N11164);
not NOT1 (N14862, N14850);
xor XOR2 (N14863, N14822, N9815);
nand NAND2 (N14864, N14863, N7660);
or OR2 (N14865, N14844, N6442);
and AND3 (N14866, N14861, N369, N6995);
xor XOR2 (N14867, N14857, N6086);
nand NAND4 (N14868, N14867, N6533, N2438, N9197);
xor XOR2 (N14869, N14856, N13578);
xor XOR2 (N14870, N14852, N2217);
buf BUF1 (N14871, N14869);
or OR2 (N14872, N14866, N1161);
and AND4 (N14873, N14859, N14138, N245, N5470);
nor NOR3 (N14874, N14864, N6899, N4154);
or OR3 (N14875, N14858, N10127, N5237);
xor XOR2 (N14876, N14871, N8039);
buf BUF1 (N14877, N14876);
xor XOR2 (N14878, N14877, N3345);
and AND4 (N14879, N14870, N14093, N10435, N8714);
nand NAND4 (N14880, N14862, N12982, N7294, N192);
buf BUF1 (N14881, N14878);
nand NAND4 (N14882, N14879, N14705, N7849, N12670);
buf BUF1 (N14883, N14873);
not NOT1 (N14884, N14875);
not NOT1 (N14885, N14868);
or OR3 (N14886, N14874, N7197, N9281);
not NOT1 (N14887, N14865);
not NOT1 (N14888, N14883);
nand NAND4 (N14889, N14884, N12462, N5545, N7031);
or OR2 (N14890, N14887, N14531);
buf BUF1 (N14891, N14890);
buf BUF1 (N14892, N14882);
nand NAND3 (N14893, N14880, N5932, N595);
or OR2 (N14894, N14891, N2346);
nand NAND2 (N14895, N14886, N832);
not NOT1 (N14896, N14893);
nand NAND3 (N14897, N14896, N9178, N8484);
not NOT1 (N14898, N14894);
nand NAND3 (N14899, N14892, N3477, N2646);
nand NAND2 (N14900, N14885, N12992);
buf BUF1 (N14901, N14898);
and AND3 (N14902, N14899, N3032, N1123);
and AND2 (N14903, N14889, N1615);
nor NOR4 (N14904, N14872, N10525, N2717, N13626);
buf BUF1 (N14905, N14901);
not NOT1 (N14906, N14905);
and AND3 (N14907, N14904, N368, N4298);
xor XOR2 (N14908, N14881, N6197);
and AND3 (N14909, N14906, N10796, N2533);
nand NAND2 (N14910, N14888, N4301);
not NOT1 (N14911, N14907);
and AND4 (N14912, N14902, N10059, N937, N3429);
buf BUF1 (N14913, N14912);
not NOT1 (N14914, N14913);
not NOT1 (N14915, N14897);
and AND3 (N14916, N14915, N7461, N11110);
or OR4 (N14917, N14910, N320, N298, N8511);
nand NAND3 (N14918, N14914, N3390, N193);
nand NAND4 (N14919, N14916, N8262, N2695, N12483);
or OR4 (N14920, N14911, N3679, N7164, N6213);
buf BUF1 (N14921, N14919);
xor XOR2 (N14922, N14917, N9137);
or OR4 (N14923, N14903, N5457, N5075, N8686);
or OR2 (N14924, N14920, N1042);
or OR3 (N14925, N14908, N8717, N7443);
not NOT1 (N14926, N14924);
and AND3 (N14927, N14923, N4607, N12297);
not NOT1 (N14928, N14900);
buf BUF1 (N14929, N14928);
nand NAND4 (N14930, N14929, N1953, N9550, N3787);
nor NOR2 (N14931, N14918, N9425);
buf BUF1 (N14932, N14895);
not NOT1 (N14933, N14922);
not NOT1 (N14934, N14933);
nand NAND2 (N14935, N14921, N11863);
or OR3 (N14936, N14927, N1041, N10535);
buf BUF1 (N14937, N14931);
xor XOR2 (N14938, N14930, N9541);
xor XOR2 (N14939, N14935, N3760);
xor XOR2 (N14940, N14860, N4950);
buf BUF1 (N14941, N14926);
or OR4 (N14942, N14940, N5579, N3252, N2405);
xor XOR2 (N14943, N14942, N6653);
buf BUF1 (N14944, N14932);
buf BUF1 (N14945, N14944);
buf BUF1 (N14946, N14939);
nand NAND4 (N14947, N14941, N9931, N13312, N12340);
nand NAND4 (N14948, N14937, N5763, N11639, N8836);
buf BUF1 (N14949, N14946);
not NOT1 (N14950, N14949);
buf BUF1 (N14951, N14950);
nor NOR3 (N14952, N14945, N14885, N353);
nor NOR4 (N14953, N14934, N241, N13320, N10081);
nor NOR2 (N14954, N14938, N672);
and AND2 (N14955, N14947, N4480);
nand NAND2 (N14956, N14936, N12691);
nor NOR4 (N14957, N14952, N1017, N5745, N14375);
or OR4 (N14958, N14909, N2732, N814, N1266);
xor XOR2 (N14959, N14943, N864);
not NOT1 (N14960, N14951);
buf BUF1 (N14961, N14957);
or OR3 (N14962, N14958, N11205, N11911);
buf BUF1 (N14963, N14953);
or OR4 (N14964, N14955, N9756, N1640, N1993);
and AND2 (N14965, N14964, N14570);
or OR3 (N14966, N14948, N12667, N7195);
xor XOR2 (N14967, N14960, N9172);
not NOT1 (N14968, N14925);
buf BUF1 (N14969, N14962);
or OR4 (N14970, N14954, N9244, N14025, N13711);
xor XOR2 (N14971, N14959, N3033);
buf BUF1 (N14972, N14966);
buf BUF1 (N14973, N14963);
or OR3 (N14974, N14972, N13127, N5162);
not NOT1 (N14975, N14961);
nand NAND4 (N14976, N14974, N12979, N276, N9499);
xor XOR2 (N14977, N14969, N940);
nand NAND4 (N14978, N14977, N7623, N488, N12181);
or OR3 (N14979, N14968, N11849, N11636);
nand NAND3 (N14980, N14967, N3164, N12192);
not NOT1 (N14981, N14980);
not NOT1 (N14982, N14971);
or OR3 (N14983, N14981, N7760, N11045);
buf BUF1 (N14984, N14973);
nand NAND4 (N14985, N14965, N9636, N12344, N3264);
and AND2 (N14986, N14970, N6826);
or OR4 (N14987, N14956, N1900, N13018, N4183);
xor XOR2 (N14988, N14978, N5061);
buf BUF1 (N14989, N14985);
buf BUF1 (N14990, N14988);
or OR3 (N14991, N14982, N4006, N7709);
buf BUF1 (N14992, N14975);
and AND3 (N14993, N14987, N700, N7812);
xor XOR2 (N14994, N14984, N4028);
nand NAND4 (N14995, N14992, N5884, N6268, N13889);
nand NAND2 (N14996, N14995, N6205);
nand NAND3 (N14997, N14990, N8384, N12241);
nor NOR3 (N14998, N14979, N6493, N1883);
and AND3 (N14999, N14997, N4018, N1654);
or OR2 (N15000, N14989, N12910);
or OR4 (N15001, N14986, N8062, N7166, N4600);
not NOT1 (N15002, N14976);
buf BUF1 (N15003, N14983);
or OR4 (N15004, N15001, N11941, N6559, N9742);
nor NOR4 (N15005, N14998, N13629, N135, N12789);
or OR4 (N15006, N14996, N2382, N110, N3081);
nor NOR4 (N15007, N14991, N11911, N5396, N5197);
nand NAND3 (N15008, N15005, N905, N206);
buf BUF1 (N15009, N14999);
nand NAND4 (N15010, N15003, N13962, N9497, N410);
buf BUF1 (N15011, N15008);
or OR4 (N15012, N15002, N2979, N5723, N1306);
not NOT1 (N15013, N15004);
xor XOR2 (N15014, N15012, N6521);
and AND2 (N15015, N15014, N10774);
and AND3 (N15016, N15011, N8147, N8293);
xor XOR2 (N15017, N15013, N1688);
and AND3 (N15018, N15016, N768, N1695);
buf BUF1 (N15019, N15017);
nand NAND2 (N15020, N15006, N2068);
nand NAND2 (N15021, N15018, N9622);
and AND3 (N15022, N15021, N8194, N12279);
nand NAND4 (N15023, N15022, N12885, N10809, N4187);
buf BUF1 (N15024, N15009);
and AND3 (N15025, N15020, N13980, N5969);
or OR2 (N15026, N15024, N5737);
and AND4 (N15027, N14993, N1921, N11388, N7768);
nor NOR4 (N15028, N15000, N11853, N11589, N7469);
buf BUF1 (N15029, N15023);
nand NAND4 (N15030, N15029, N13197, N13954, N6059);
buf BUF1 (N15031, N15027);
nand NAND4 (N15032, N15030, N1074, N3408, N12293);
nand NAND2 (N15033, N15028, N5482);
and AND2 (N15034, N15033, N925);
buf BUF1 (N15035, N15031);
xor XOR2 (N15036, N15035, N12922);
nand NAND3 (N15037, N15010, N11647, N11248);
or OR4 (N15038, N15025, N7750, N1993, N296);
and AND4 (N15039, N15036, N11885, N555, N6678);
and AND3 (N15040, N15007, N13626, N8114);
nand NAND2 (N15041, N15015, N33);
or OR3 (N15042, N15040, N13579, N7749);
nand NAND4 (N15043, N15037, N3580, N7378, N2255);
buf BUF1 (N15044, N14994);
or OR3 (N15045, N15041, N6584, N3594);
nand NAND4 (N15046, N15039, N5220, N1049, N8014);
xor XOR2 (N15047, N15043, N9521);
nand NAND3 (N15048, N15047, N6647, N6038);
or OR2 (N15049, N15046, N6109);
not NOT1 (N15050, N15038);
nor NOR3 (N15051, N15044, N14286, N13857);
buf BUF1 (N15052, N15026);
buf BUF1 (N15053, N15052);
or OR2 (N15054, N15048, N2888);
nand NAND3 (N15055, N15019, N14195, N4532);
or OR4 (N15056, N15051, N1630, N12056, N1276);
nor NOR2 (N15057, N15049, N751);
buf BUF1 (N15058, N15056);
xor XOR2 (N15059, N15055, N6814);
buf BUF1 (N15060, N15050);
buf BUF1 (N15061, N15034);
nand NAND3 (N15062, N15053, N3712, N2618);
not NOT1 (N15063, N15032);
nor NOR3 (N15064, N15058, N2665, N7606);
not NOT1 (N15065, N15059);
buf BUF1 (N15066, N15054);
or OR4 (N15067, N15063, N10677, N4433, N9859);
and AND4 (N15068, N15061, N13557, N5805, N6525);
not NOT1 (N15069, N15045);
buf BUF1 (N15070, N15065);
and AND3 (N15071, N15064, N9136, N3744);
nor NOR3 (N15072, N15069, N1113, N4803);
not NOT1 (N15073, N15068);
buf BUF1 (N15074, N15062);
nand NAND3 (N15075, N15070, N9695, N1443);
not NOT1 (N15076, N15060);
not NOT1 (N15077, N15042);
xor XOR2 (N15078, N15057, N2617);
xor XOR2 (N15079, N15072, N10776);
and AND4 (N15080, N15078, N14857, N3300, N7104);
not NOT1 (N15081, N15074);
and AND3 (N15082, N15077, N9225, N3103);
not NOT1 (N15083, N15066);
nor NOR4 (N15084, N15082, N1011, N5982, N5182);
not NOT1 (N15085, N15079);
or OR3 (N15086, N15084, N7483, N4210);
xor XOR2 (N15087, N15083, N5961);
nand NAND3 (N15088, N15081, N4075, N14633);
nand NAND4 (N15089, N15073, N4258, N2247, N45);
and AND2 (N15090, N15076, N9352);
or OR3 (N15091, N15086, N11553, N4940);
nor NOR4 (N15092, N15087, N10919, N11576, N6638);
and AND3 (N15093, N15075, N14040, N4804);
nor NOR4 (N15094, N15067, N2781, N12581, N11035);
or OR2 (N15095, N15089, N11160);
buf BUF1 (N15096, N15092);
buf BUF1 (N15097, N15094);
or OR2 (N15098, N15080, N10474);
nor NOR4 (N15099, N15088, N14257, N12416, N6602);
xor XOR2 (N15100, N15097, N7371);
buf BUF1 (N15101, N15099);
buf BUF1 (N15102, N15095);
xor XOR2 (N15103, N15085, N2935);
buf BUF1 (N15104, N15093);
nor NOR4 (N15105, N15102, N11160, N14424, N8705);
buf BUF1 (N15106, N15104);
not NOT1 (N15107, N15106);
not NOT1 (N15108, N15090);
or OR3 (N15109, N15100, N2679, N817);
nor NOR4 (N15110, N15071, N2033, N604, N15044);
xor XOR2 (N15111, N15108, N14314);
nand NAND3 (N15112, N15110, N8683, N7210);
nand NAND3 (N15113, N15107, N5436, N11199);
nor NOR2 (N15114, N15096, N4360);
and AND4 (N15115, N15103, N2617, N33, N3133);
not NOT1 (N15116, N15109);
buf BUF1 (N15117, N15113);
nor NOR4 (N15118, N15101, N10446, N10822, N8025);
nor NOR4 (N15119, N15112, N3526, N5829, N2129);
xor XOR2 (N15120, N15117, N14479);
or OR3 (N15121, N15118, N12005, N4958);
nand NAND4 (N15122, N15105, N14442, N15010, N6461);
buf BUF1 (N15123, N15114);
xor XOR2 (N15124, N15091, N10293);
not NOT1 (N15125, N15124);
nor NOR4 (N15126, N15125, N9423, N8657, N8740);
xor XOR2 (N15127, N15115, N9082);
or OR4 (N15128, N15120, N9666, N10387, N13087);
nor NOR2 (N15129, N15123, N2705);
not NOT1 (N15130, N15121);
or OR3 (N15131, N15126, N9483, N499);
nor NOR4 (N15132, N15111, N9647, N3273, N5817);
nor NOR2 (N15133, N15128, N10425);
nand NAND2 (N15134, N15130, N9172);
nor NOR2 (N15135, N15131, N13472);
xor XOR2 (N15136, N15116, N8718);
or OR4 (N15137, N15119, N3641, N11965, N534);
nand NAND3 (N15138, N15134, N7746, N8665);
not NOT1 (N15139, N15137);
xor XOR2 (N15140, N15132, N10029);
or OR4 (N15141, N15133, N3400, N7604, N14442);
or OR3 (N15142, N15139, N13992, N13782);
nand NAND3 (N15143, N15142, N12923, N7468);
xor XOR2 (N15144, N15141, N5539);
nand NAND3 (N15145, N15143, N11366, N1647);
not NOT1 (N15146, N15145);
and AND4 (N15147, N15122, N3410, N9308, N9029);
or OR4 (N15148, N15140, N575, N8956, N6574);
nand NAND2 (N15149, N15135, N697);
not NOT1 (N15150, N15098);
not NOT1 (N15151, N15148);
and AND3 (N15152, N15129, N1612, N10363);
xor XOR2 (N15153, N15150, N14191);
xor XOR2 (N15154, N15147, N10903);
nor NOR4 (N15155, N15127, N8635, N3437, N12409);
xor XOR2 (N15156, N15136, N12675);
and AND3 (N15157, N15144, N13769, N7802);
nand NAND3 (N15158, N15149, N13753, N1815);
nor NOR4 (N15159, N15154, N12451, N9957, N13659);
or OR3 (N15160, N15159, N9765, N3074);
and AND2 (N15161, N15157, N12813);
nor NOR3 (N15162, N15151, N14743, N3766);
and AND4 (N15163, N15155, N1954, N12635, N12953);
or OR3 (N15164, N15138, N2069, N5805);
nor NOR2 (N15165, N15160, N4121);
nand NAND2 (N15166, N15161, N3855);
and AND2 (N15167, N15152, N2770);
not NOT1 (N15168, N15164);
nand NAND4 (N15169, N15156, N9390, N14342, N10384);
nor NOR2 (N15170, N15166, N13638);
not NOT1 (N15171, N15163);
or OR4 (N15172, N15171, N11809, N1413, N7269);
and AND2 (N15173, N15172, N3784);
xor XOR2 (N15174, N15162, N15092);
nor NOR2 (N15175, N15153, N8188);
not NOT1 (N15176, N15174);
nand NAND3 (N15177, N15167, N14355, N14571);
nand NAND4 (N15178, N15168, N14646, N14872, N12684);
xor XOR2 (N15179, N15146, N12367);
xor XOR2 (N15180, N15177, N619);
buf BUF1 (N15181, N15180);
xor XOR2 (N15182, N15165, N1285);
not NOT1 (N15183, N15170);
xor XOR2 (N15184, N15175, N13320);
nand NAND4 (N15185, N15158, N592, N14678, N13533);
xor XOR2 (N15186, N15173, N6105);
and AND2 (N15187, N15182, N15093);
buf BUF1 (N15188, N15181);
buf BUF1 (N15189, N15183);
not NOT1 (N15190, N15178);
xor XOR2 (N15191, N15186, N2173);
not NOT1 (N15192, N15188);
buf BUF1 (N15193, N15189);
xor XOR2 (N15194, N15192, N3697);
nor NOR2 (N15195, N15185, N13159);
xor XOR2 (N15196, N15176, N4089);
buf BUF1 (N15197, N15184);
xor XOR2 (N15198, N15196, N6365);
buf BUF1 (N15199, N15191);
buf BUF1 (N15200, N15193);
not NOT1 (N15201, N15187);
xor XOR2 (N15202, N15179, N5548);
buf BUF1 (N15203, N15198);
xor XOR2 (N15204, N15195, N1044);
xor XOR2 (N15205, N15201, N5788);
not NOT1 (N15206, N15203);
not NOT1 (N15207, N15200);
nor NOR2 (N15208, N15199, N2324);
and AND3 (N15209, N15206, N13591, N4821);
buf BUF1 (N15210, N15197);
buf BUF1 (N15211, N15207);
nand NAND3 (N15212, N15210, N15104, N13325);
nor NOR4 (N15213, N15194, N1714, N14294, N4422);
not NOT1 (N15214, N15208);
and AND2 (N15215, N15204, N11338);
and AND3 (N15216, N15209, N3573, N4462);
nand NAND4 (N15217, N15205, N3250, N3028, N75);
buf BUF1 (N15218, N15213);
buf BUF1 (N15219, N15218);
not NOT1 (N15220, N15219);
or OR4 (N15221, N15212, N10673, N2018, N14566);
and AND3 (N15222, N15215, N11969, N15020);
nand NAND4 (N15223, N15222, N7189, N14479, N8173);
buf BUF1 (N15224, N15217);
not NOT1 (N15225, N15223);
not NOT1 (N15226, N15169);
xor XOR2 (N15227, N15224, N113);
not NOT1 (N15228, N15190);
buf BUF1 (N15229, N15202);
nand NAND2 (N15230, N15220, N5211);
nand NAND2 (N15231, N15227, N13961);
nor NOR4 (N15232, N15221, N14876, N6914, N8842);
nand NAND2 (N15233, N15230, N2928);
xor XOR2 (N15234, N15233, N1017);
not NOT1 (N15235, N15216);
xor XOR2 (N15236, N15234, N6295);
and AND4 (N15237, N15226, N6656, N7280, N5935);
not NOT1 (N15238, N15232);
buf BUF1 (N15239, N15231);
or OR4 (N15240, N15239, N10295, N8029, N1700);
and AND4 (N15241, N15237, N12109, N4836, N6490);
nand NAND3 (N15242, N15236, N12740, N6144);
xor XOR2 (N15243, N15242, N4642);
nor NOR4 (N15244, N15229, N4908, N4930, N10622);
buf BUF1 (N15245, N15244);
or OR3 (N15246, N15211, N972, N6487);
nor NOR3 (N15247, N15243, N7545, N13005);
xor XOR2 (N15248, N15240, N12572);
or OR4 (N15249, N15247, N7298, N13607, N5988);
and AND3 (N15250, N15225, N3919, N6415);
or OR4 (N15251, N15214, N11364, N4840, N4557);
xor XOR2 (N15252, N15250, N6418);
or OR4 (N15253, N15241, N4663, N10581, N3309);
xor XOR2 (N15254, N15246, N9681);
nor NOR4 (N15255, N15251, N2343, N9624, N7473);
nor NOR4 (N15256, N15238, N800, N3522, N6665);
xor XOR2 (N15257, N15245, N9144);
nand NAND3 (N15258, N15256, N5759, N1291);
nand NAND4 (N15259, N15252, N7987, N10685, N4630);
not NOT1 (N15260, N15248);
xor XOR2 (N15261, N15253, N3083);
buf BUF1 (N15262, N15259);
not NOT1 (N15263, N15258);
buf BUF1 (N15264, N15262);
not NOT1 (N15265, N15235);
buf BUF1 (N15266, N15254);
buf BUF1 (N15267, N15260);
or OR2 (N15268, N15266, N1157);
nor NOR2 (N15269, N15267, N5787);
buf BUF1 (N15270, N15261);
or OR3 (N15271, N15268, N880, N7175);
or OR2 (N15272, N15257, N2826);
nor NOR4 (N15273, N15228, N4429, N3150, N11278);
and AND2 (N15274, N15264, N3409);
nand NAND4 (N15275, N15255, N9880, N3060, N6200);
nor NOR2 (N15276, N15275, N5943);
not NOT1 (N15277, N15273);
nand NAND3 (N15278, N15263, N11043, N10505);
buf BUF1 (N15279, N15277);
or OR4 (N15280, N15278, N7026, N2171, N1166);
buf BUF1 (N15281, N15279);
or OR4 (N15282, N15280, N14095, N8917, N14268);
not NOT1 (N15283, N15272);
nand NAND3 (N15284, N15274, N13348, N5504);
and AND4 (N15285, N15249, N3997, N8418, N7872);
or OR4 (N15286, N15284, N14606, N6667, N12969);
nand NAND3 (N15287, N15286, N14285, N6816);
buf BUF1 (N15288, N15282);
xor XOR2 (N15289, N15281, N10177);
nand NAND4 (N15290, N15289, N7946, N7235, N7440);
and AND4 (N15291, N15290, N9171, N385, N6586);
and AND2 (N15292, N15276, N9591);
buf BUF1 (N15293, N15288);
buf BUF1 (N15294, N15293);
and AND4 (N15295, N15265, N5350, N2804, N5698);
nor NOR2 (N15296, N15295, N6237);
nor NOR4 (N15297, N15283, N11324, N13229, N6660);
or OR2 (N15298, N15292, N9966);
and AND2 (N15299, N15296, N13907);
not NOT1 (N15300, N15270);
not NOT1 (N15301, N15285);
xor XOR2 (N15302, N15300, N10421);
and AND4 (N15303, N15298, N166, N4872, N43);
xor XOR2 (N15304, N15271, N13467);
not NOT1 (N15305, N15303);
xor XOR2 (N15306, N15299, N739);
or OR4 (N15307, N15294, N2745, N12641, N2609);
buf BUF1 (N15308, N15306);
buf BUF1 (N15309, N15305);
nor NOR3 (N15310, N15291, N13045, N11024);
not NOT1 (N15311, N15310);
or OR4 (N15312, N15302, N3884, N7661, N12370);
and AND3 (N15313, N15309, N12221, N4687);
or OR2 (N15314, N15287, N8063);
nor NOR2 (N15315, N15314, N3551);
not NOT1 (N15316, N15311);
nor NOR2 (N15317, N15312, N8845);
and AND2 (N15318, N15317, N409);
buf BUF1 (N15319, N15316);
or OR3 (N15320, N15308, N4919, N6074);
not NOT1 (N15321, N15315);
nand NAND4 (N15322, N15321, N8788, N4560, N8598);
and AND4 (N15323, N15318, N1422, N807, N3358);
or OR2 (N15324, N15301, N7741);
xor XOR2 (N15325, N15297, N2620);
or OR3 (N15326, N15304, N14446, N10411);
xor XOR2 (N15327, N15320, N9548);
buf BUF1 (N15328, N15327);
buf BUF1 (N15329, N15307);
nor NOR4 (N15330, N15323, N8622, N8791, N2645);
nand NAND3 (N15331, N15269, N6848, N8100);
or OR3 (N15332, N15326, N5379, N1403);
or OR3 (N15333, N15331, N13448, N1092);
nor NOR4 (N15334, N15330, N13308, N3457, N7298);
nand NAND2 (N15335, N15325, N14943);
xor XOR2 (N15336, N15313, N2558);
nor NOR3 (N15337, N15324, N519, N396);
nand NAND4 (N15338, N15322, N10411, N9778, N13683);
nor NOR2 (N15339, N15336, N4536);
or OR3 (N15340, N15334, N4128, N11376);
nor NOR4 (N15341, N15319, N7681, N1705, N1360);
buf BUF1 (N15342, N15337);
xor XOR2 (N15343, N15339, N14587);
buf BUF1 (N15344, N15340);
nand NAND3 (N15345, N15338, N15001, N12949);
nor NOR3 (N15346, N15329, N6524, N887);
xor XOR2 (N15347, N15346, N10585);
nor NOR4 (N15348, N15347, N13044, N7976, N7878);
and AND2 (N15349, N15344, N9919);
xor XOR2 (N15350, N15345, N14764);
buf BUF1 (N15351, N15350);
buf BUF1 (N15352, N15349);
not NOT1 (N15353, N15335);
nor NOR2 (N15354, N15343, N1604);
or OR2 (N15355, N15332, N1364);
xor XOR2 (N15356, N15355, N2039);
xor XOR2 (N15357, N15341, N5619);
or OR2 (N15358, N15354, N7236);
or OR4 (N15359, N15348, N7007, N10431, N10241);
nor NOR4 (N15360, N15328, N5807, N5683, N1945);
buf BUF1 (N15361, N15353);
nor NOR3 (N15362, N15359, N4001, N9171);
nor NOR4 (N15363, N15360, N13498, N3443, N373);
and AND3 (N15364, N15361, N4477, N12730);
buf BUF1 (N15365, N15356);
or OR3 (N15366, N15333, N13268, N4605);
not NOT1 (N15367, N15352);
buf BUF1 (N15368, N15358);
buf BUF1 (N15369, N15368);
buf BUF1 (N15370, N15369);
buf BUF1 (N15371, N15363);
not NOT1 (N15372, N15365);
xor XOR2 (N15373, N15357, N11962);
buf BUF1 (N15374, N15351);
or OR3 (N15375, N15370, N8713, N15131);
buf BUF1 (N15376, N15372);
xor XOR2 (N15377, N15374, N1054);
xor XOR2 (N15378, N15364, N2928);
nand NAND2 (N15379, N15373, N8088);
nand NAND2 (N15380, N15367, N6324);
and AND3 (N15381, N15375, N2429, N8510);
buf BUF1 (N15382, N15371);
nor NOR4 (N15383, N15382, N9413, N13789, N14178);
not NOT1 (N15384, N15362);
nand NAND2 (N15385, N15378, N9571);
not NOT1 (N15386, N15384);
not NOT1 (N15387, N15342);
nand NAND2 (N15388, N15379, N14042);
buf BUF1 (N15389, N15376);
nand NAND2 (N15390, N15388, N12078);
not NOT1 (N15391, N15390);
nor NOR4 (N15392, N15380, N14318, N5175, N14797);
nand NAND3 (N15393, N15387, N6013, N14016);
or OR4 (N15394, N15381, N1504, N5792, N6388);
nor NOR4 (N15395, N15393, N10729, N13645, N9395);
nor NOR2 (N15396, N15392, N13522);
and AND3 (N15397, N15386, N14842, N10222);
not NOT1 (N15398, N15397);
buf BUF1 (N15399, N15366);
and AND2 (N15400, N15383, N5325);
nor NOR4 (N15401, N15400, N15257, N4804, N3380);
nor NOR2 (N15402, N15398, N13003);
nand NAND3 (N15403, N15394, N3116, N10321);
buf BUF1 (N15404, N15385);
not NOT1 (N15405, N15403);
buf BUF1 (N15406, N15395);
or OR2 (N15407, N15399, N15310);
buf BUF1 (N15408, N15402);
or OR3 (N15409, N15391, N8824, N1381);
buf BUF1 (N15410, N15408);
xor XOR2 (N15411, N15377, N9190);
xor XOR2 (N15412, N15396, N14634);
xor XOR2 (N15413, N15389, N15022);
or OR4 (N15414, N15404, N1237, N3896, N8281);
or OR3 (N15415, N15411, N3698, N2714);
xor XOR2 (N15416, N15406, N5233);
and AND3 (N15417, N15416, N3732, N15401);
xor XOR2 (N15418, N3008, N9388);
and AND4 (N15419, N15415, N10660, N10724, N10362);
not NOT1 (N15420, N15410);
nor NOR3 (N15421, N15412, N398, N4856);
xor XOR2 (N15422, N15407, N11645);
and AND3 (N15423, N15421, N6750, N1647);
and AND4 (N15424, N15420, N12423, N3002, N12346);
nor NOR4 (N15425, N15423, N3997, N12695, N4212);
and AND2 (N15426, N15409, N9584);
xor XOR2 (N15427, N15418, N5362);
and AND3 (N15428, N15414, N13419, N9937);
and AND3 (N15429, N15405, N3441, N5252);
not NOT1 (N15430, N15419);
nor NOR2 (N15431, N15422, N8407);
or OR2 (N15432, N15413, N12181);
or OR3 (N15433, N15425, N13412, N12912);
or OR4 (N15434, N15430, N14447, N3886, N850);
nor NOR2 (N15435, N15428, N3657);
or OR4 (N15436, N15434, N634, N12779, N2721);
not NOT1 (N15437, N15436);
xor XOR2 (N15438, N15424, N4350);
buf BUF1 (N15439, N15437);
or OR3 (N15440, N15431, N12953, N1475);
nor NOR4 (N15441, N15439, N6528, N11508, N4266);
nand NAND3 (N15442, N15440, N7665, N964);
or OR3 (N15443, N15435, N1130, N11395);
or OR3 (N15444, N15417, N618, N1050);
or OR4 (N15445, N15438, N7482, N2380, N4274);
or OR2 (N15446, N15444, N12213);
xor XOR2 (N15447, N15433, N5279);
nor NOR2 (N15448, N15445, N13858);
buf BUF1 (N15449, N15429);
xor XOR2 (N15450, N15427, N13180);
xor XOR2 (N15451, N15432, N2997);
nor NOR2 (N15452, N15451, N12263);
xor XOR2 (N15453, N15443, N5878);
or OR4 (N15454, N15442, N5266, N3196, N11913);
nand NAND3 (N15455, N15449, N8580, N11891);
and AND3 (N15456, N15455, N10168, N1779);
nor NOR4 (N15457, N15452, N9033, N2912, N3154);
nor NOR3 (N15458, N15426, N14924, N14119);
and AND2 (N15459, N15453, N6063);
buf BUF1 (N15460, N15458);
not NOT1 (N15461, N15456);
nand NAND2 (N15462, N15441, N8208);
buf BUF1 (N15463, N15454);
nor NOR4 (N15464, N15461, N2218, N3827, N1612);
xor XOR2 (N15465, N15457, N11435);
and AND3 (N15466, N15446, N4349, N11089);
nor NOR3 (N15467, N15460, N10358, N450);
xor XOR2 (N15468, N15466, N6371);
nor NOR2 (N15469, N15468, N13291);
not NOT1 (N15470, N15459);
xor XOR2 (N15471, N15447, N2881);
nor NOR2 (N15472, N15462, N13752);
or OR3 (N15473, N15467, N791, N13285);
nor NOR3 (N15474, N15464, N7246, N7297);
xor XOR2 (N15475, N15463, N3046);
and AND3 (N15476, N15475, N9657, N876);
xor XOR2 (N15477, N15450, N3147);
or OR2 (N15478, N15477, N5798);
nand NAND4 (N15479, N15465, N1606, N9432, N7651);
or OR4 (N15480, N15471, N8607, N11130, N5068);
xor XOR2 (N15481, N15474, N10095);
nor NOR2 (N15482, N15470, N7843);
not NOT1 (N15483, N15448);
and AND2 (N15484, N15482, N10836);
and AND3 (N15485, N15483, N13556, N459);
nor NOR3 (N15486, N15481, N4696, N11316);
xor XOR2 (N15487, N15472, N11711);
buf BUF1 (N15488, N15479);
or OR2 (N15489, N15478, N2162);
xor XOR2 (N15490, N15489, N2900);
buf BUF1 (N15491, N15469);
nand NAND2 (N15492, N15473, N9981);
nor NOR4 (N15493, N15492, N7450, N7091, N13513);
nor NOR3 (N15494, N15480, N10960, N671);
and AND2 (N15495, N15484, N14719);
buf BUF1 (N15496, N15476);
and AND2 (N15497, N15488, N11733);
nor NOR3 (N15498, N15496, N10599, N2803);
buf BUF1 (N15499, N15494);
and AND3 (N15500, N15495, N3916, N15252);
nand NAND4 (N15501, N15499, N3121, N7785, N9808);
nor NOR2 (N15502, N15500, N4421);
nor NOR4 (N15503, N15501, N1345, N7249, N15225);
nand NAND2 (N15504, N15485, N13610);
xor XOR2 (N15505, N15504, N7414);
xor XOR2 (N15506, N15490, N15132);
nand NAND2 (N15507, N15486, N6764);
not NOT1 (N15508, N15502);
xor XOR2 (N15509, N15493, N11111);
nand NAND3 (N15510, N15497, N127, N400);
xor XOR2 (N15511, N15508, N8216);
nor NOR3 (N15512, N15506, N14022, N5154);
or OR3 (N15513, N15507, N7795, N13569);
nand NAND2 (N15514, N15498, N3732);
xor XOR2 (N15515, N15512, N15141);
buf BUF1 (N15516, N15505);
nor NOR3 (N15517, N15487, N9012, N2676);
not NOT1 (N15518, N15511);
not NOT1 (N15519, N15503);
nand NAND3 (N15520, N15509, N3331, N14653);
nand NAND2 (N15521, N15491, N5109);
buf BUF1 (N15522, N15520);
nand NAND3 (N15523, N15515, N1571, N14973);
not NOT1 (N15524, N15519);
xor XOR2 (N15525, N15514, N14773);
xor XOR2 (N15526, N15521, N4525);
xor XOR2 (N15527, N15518, N4606);
not NOT1 (N15528, N15516);
nor NOR2 (N15529, N15510, N5408);
not NOT1 (N15530, N15513);
not NOT1 (N15531, N15522);
or OR4 (N15532, N15531, N9296, N3264, N9574);
xor XOR2 (N15533, N15524, N12680);
nand NAND2 (N15534, N15517, N13519);
nor NOR2 (N15535, N15534, N6592);
not NOT1 (N15536, N15529);
or OR4 (N15537, N15533, N11478, N8042, N15268);
or OR2 (N15538, N15536, N6282);
nor NOR3 (N15539, N15535, N533, N4196);
or OR3 (N15540, N15537, N3570, N964);
not NOT1 (N15541, N15538);
and AND4 (N15542, N15523, N7344, N2318, N378);
xor XOR2 (N15543, N15530, N15054);
nor NOR2 (N15544, N15532, N14254);
and AND2 (N15545, N15525, N6170);
xor XOR2 (N15546, N15544, N12092);
nor NOR2 (N15547, N15539, N876);
buf BUF1 (N15548, N15541);
xor XOR2 (N15549, N15528, N12823);
and AND3 (N15550, N15546, N4435, N1024);
buf BUF1 (N15551, N15548);
and AND4 (N15552, N15527, N9474, N1851, N7464);
xor XOR2 (N15553, N15551, N8749);
buf BUF1 (N15554, N15550);
buf BUF1 (N15555, N15545);
xor XOR2 (N15556, N15540, N4967);
buf BUF1 (N15557, N15542);
or OR4 (N15558, N15543, N14419, N10340, N13585);
xor XOR2 (N15559, N15547, N13928);
not NOT1 (N15560, N15526);
not NOT1 (N15561, N15556);
or OR4 (N15562, N15559, N8905, N5685, N13330);
and AND4 (N15563, N15560, N7460, N11619, N2316);
nand NAND2 (N15564, N15554, N3525);
or OR4 (N15565, N15557, N9827, N8999, N7058);
not NOT1 (N15566, N15555);
not NOT1 (N15567, N15563);
nor NOR3 (N15568, N15561, N15367, N14148);
nand NAND3 (N15569, N15552, N2924, N12956);
or OR4 (N15570, N15564, N3241, N12070, N8668);
xor XOR2 (N15571, N15568, N14719);
xor XOR2 (N15572, N15565, N10433);
or OR3 (N15573, N15549, N11204, N5883);
nand NAND3 (N15574, N15573, N8736, N3928);
nand NAND4 (N15575, N15571, N13490, N9711, N9572);
nor NOR3 (N15576, N15570, N13650, N536);
or OR3 (N15577, N15576, N249, N11881);
nand NAND4 (N15578, N15569, N9557, N10689, N11463);
buf BUF1 (N15579, N15574);
xor XOR2 (N15580, N15575, N15158);
nand NAND4 (N15581, N15567, N7179, N8431, N4689);
xor XOR2 (N15582, N15572, N11439);
and AND3 (N15583, N15558, N3858, N14629);
nor NOR2 (N15584, N15580, N7031);
nand NAND3 (N15585, N15579, N3630, N8115);
nor NOR2 (N15586, N15577, N1804);
or OR4 (N15587, N15583, N9599, N3752, N10407);
xor XOR2 (N15588, N15582, N15546);
xor XOR2 (N15589, N15588, N11899);
buf BUF1 (N15590, N15578);
and AND4 (N15591, N15566, N4727, N10318, N13620);
buf BUF1 (N15592, N15584);
and AND2 (N15593, N15592, N15380);
xor XOR2 (N15594, N15586, N12752);
and AND2 (N15595, N15587, N979);
nor NOR3 (N15596, N15562, N4179, N13976);
nand NAND3 (N15597, N15596, N6600, N12363);
buf BUF1 (N15598, N15553);
or OR4 (N15599, N15590, N4233, N800, N14382);
nand NAND3 (N15600, N15591, N7291, N14503);
buf BUF1 (N15601, N15581);
xor XOR2 (N15602, N15601, N2985);
and AND4 (N15603, N15593, N3399, N3545, N15395);
nor NOR2 (N15604, N15600, N7284);
xor XOR2 (N15605, N15589, N4029);
not NOT1 (N15606, N15585);
nor NOR3 (N15607, N15595, N10526, N4910);
xor XOR2 (N15608, N15594, N8830);
or OR2 (N15609, N15607, N7601);
nand NAND4 (N15610, N15597, N2858, N3438, N11120);
not NOT1 (N15611, N15598);
xor XOR2 (N15612, N15604, N14289);
nor NOR4 (N15613, N15609, N11237, N11088, N11264);
buf BUF1 (N15614, N15611);
nor NOR3 (N15615, N15599, N2416, N6633);
nand NAND3 (N15616, N15608, N1798, N7995);
buf BUF1 (N15617, N15612);
not NOT1 (N15618, N15606);
buf BUF1 (N15619, N15613);
xor XOR2 (N15620, N15616, N2666);
buf BUF1 (N15621, N15614);
or OR2 (N15622, N15603, N1983);
xor XOR2 (N15623, N15618, N3660);
xor XOR2 (N15624, N15617, N3703);
nor NOR3 (N15625, N15620, N8846, N4611);
nor NOR3 (N15626, N15624, N13535, N4656);
buf BUF1 (N15627, N15626);
not NOT1 (N15628, N15605);
not NOT1 (N15629, N15625);
xor XOR2 (N15630, N15623, N14839);
and AND4 (N15631, N15610, N9857, N13553, N1576);
not NOT1 (N15632, N15627);
xor XOR2 (N15633, N15602, N3486);
xor XOR2 (N15634, N15628, N9728);
nand NAND2 (N15635, N15615, N7862);
or OR3 (N15636, N15619, N7213, N12056);
not NOT1 (N15637, N15633);
nand NAND4 (N15638, N15634, N10128, N10308, N11364);
nand NAND4 (N15639, N15636, N12079, N2880, N10025);
not NOT1 (N15640, N15635);
xor XOR2 (N15641, N15637, N2226);
and AND3 (N15642, N15641, N10264, N7792);
and AND2 (N15643, N15642, N14359);
and AND4 (N15644, N15632, N9796, N7187, N8775);
nand NAND3 (N15645, N15640, N6244, N9920);
xor XOR2 (N15646, N15644, N7822);
nor NOR3 (N15647, N15631, N7420, N8294);
and AND4 (N15648, N15647, N5848, N2755, N6077);
xor XOR2 (N15649, N15629, N4336);
nand NAND4 (N15650, N15649, N5015, N5900, N10068);
or OR3 (N15651, N15646, N14717, N3920);
not NOT1 (N15652, N15651);
and AND4 (N15653, N15650, N8654, N8156, N3414);
or OR3 (N15654, N15652, N4922, N1184);
nor NOR2 (N15655, N15648, N13970);
nor NOR4 (N15656, N15654, N15372, N1500, N1693);
xor XOR2 (N15657, N15656, N5452);
and AND2 (N15658, N15655, N10283);
buf BUF1 (N15659, N15639);
and AND3 (N15660, N15659, N13678, N8450);
not NOT1 (N15661, N15660);
nand NAND4 (N15662, N15622, N5643, N14013, N14030);
nand NAND4 (N15663, N15645, N1117, N11583, N9825);
xor XOR2 (N15664, N15630, N13949);
and AND4 (N15665, N15657, N12050, N15619, N12294);
and AND4 (N15666, N15638, N3962, N10952, N3944);
xor XOR2 (N15667, N15662, N924);
buf BUF1 (N15668, N15643);
nand NAND4 (N15669, N15661, N7827, N13428, N11732);
xor XOR2 (N15670, N15653, N8190);
not NOT1 (N15671, N15668);
or OR4 (N15672, N15669, N3252, N15287, N14081);
xor XOR2 (N15673, N15667, N8760);
not NOT1 (N15674, N15621);
nand NAND2 (N15675, N15670, N7628);
nor NOR3 (N15676, N15675, N9100, N5619);
buf BUF1 (N15677, N15658);
buf BUF1 (N15678, N15666);
nor NOR4 (N15679, N15665, N6622, N246, N6910);
not NOT1 (N15680, N15677);
nand NAND3 (N15681, N15678, N962, N7481);
not NOT1 (N15682, N15664);
buf BUF1 (N15683, N15672);
or OR2 (N15684, N15674, N61);
xor XOR2 (N15685, N15671, N2694);
not NOT1 (N15686, N15676);
nor NOR3 (N15687, N15683, N9989, N2047);
or OR2 (N15688, N15685, N9608);
not NOT1 (N15689, N15684);
buf BUF1 (N15690, N15688);
buf BUF1 (N15691, N15680);
not NOT1 (N15692, N15687);
xor XOR2 (N15693, N15673, N6725);
not NOT1 (N15694, N15692);
nand NAND4 (N15695, N15693, N3029, N14437, N6999);
nand NAND4 (N15696, N15691, N14854, N14664, N10567);
buf BUF1 (N15697, N15681);
nor NOR4 (N15698, N15697, N8369, N11894, N14552);
xor XOR2 (N15699, N15698, N10222);
nand NAND3 (N15700, N15699, N529, N2689);
nor NOR3 (N15701, N15682, N5252, N13387);
nand NAND3 (N15702, N15689, N13883, N4212);
not NOT1 (N15703, N15686);
and AND4 (N15704, N15703, N375, N3635, N15684);
and AND3 (N15705, N15679, N10754, N12152);
nand NAND3 (N15706, N15702, N13845, N4569);
nand NAND4 (N15707, N15700, N9468, N11138, N7358);
nor NOR4 (N15708, N15701, N11626, N6458, N13098);
xor XOR2 (N15709, N15690, N11847);
or OR2 (N15710, N15709, N4717);
nor NOR3 (N15711, N15705, N9626, N292);
buf BUF1 (N15712, N15663);
or OR4 (N15713, N15694, N15633, N802, N5809);
not NOT1 (N15714, N15696);
and AND3 (N15715, N15704, N14605, N12097);
nand NAND2 (N15716, N15695, N1753);
and AND3 (N15717, N15706, N9628, N823);
buf BUF1 (N15718, N15708);
nand NAND4 (N15719, N15717, N3360, N2905, N2992);
or OR2 (N15720, N15719, N4573);
not NOT1 (N15721, N15716);
not NOT1 (N15722, N15710);
nand NAND3 (N15723, N15721, N14178, N9576);
nand NAND4 (N15724, N15713, N12750, N12177, N1713);
xor XOR2 (N15725, N15714, N14314);
not NOT1 (N15726, N15724);
and AND3 (N15727, N15726, N8879, N13881);
buf BUF1 (N15728, N15712);
or OR4 (N15729, N15707, N1705, N12849, N15517);
nand NAND3 (N15730, N15722, N14009, N12664);
xor XOR2 (N15731, N15730, N14164);
buf BUF1 (N15732, N15729);
xor XOR2 (N15733, N15731, N15461);
nor NOR2 (N15734, N15723, N6730);
not NOT1 (N15735, N15725);
nor NOR2 (N15736, N15728, N5526);
nor NOR3 (N15737, N15733, N2201, N3121);
not NOT1 (N15738, N15727);
xor XOR2 (N15739, N15732, N14916);
nand NAND3 (N15740, N15738, N7130, N14196);
and AND4 (N15741, N15735, N6882, N8686, N10694);
nor NOR3 (N15742, N15736, N483, N5967);
not NOT1 (N15743, N15741);
xor XOR2 (N15744, N15740, N12831);
and AND2 (N15745, N15715, N10714);
nand NAND3 (N15746, N15744, N10212, N6707);
or OR2 (N15747, N15737, N5317);
or OR4 (N15748, N15739, N15287, N794, N8173);
and AND4 (N15749, N15720, N15270, N5446, N13278);
or OR3 (N15750, N15745, N666, N9484);
nor NOR3 (N15751, N15718, N12784, N5020);
or OR3 (N15752, N15748, N4075, N15551);
and AND3 (N15753, N15742, N10443, N13919);
and AND2 (N15754, N15734, N4686);
or OR4 (N15755, N15746, N9792, N12207, N7648);
nor NOR3 (N15756, N15750, N2296, N10083);
buf BUF1 (N15757, N15752);
nor NOR2 (N15758, N15754, N13935);
nand NAND2 (N15759, N15747, N7659);
nor NOR2 (N15760, N15743, N6217);
nand NAND2 (N15761, N15759, N7117);
buf BUF1 (N15762, N15757);
and AND3 (N15763, N15760, N4853, N12891);
nand NAND4 (N15764, N15762, N7510, N11179, N6346);
xor XOR2 (N15765, N15756, N13839);
xor XOR2 (N15766, N15763, N1732);
not NOT1 (N15767, N15765);
nor NOR3 (N15768, N15758, N3211, N4551);
not NOT1 (N15769, N15768);
nand NAND2 (N15770, N15753, N5056);
xor XOR2 (N15771, N15711, N753);
nand NAND3 (N15772, N15749, N13684, N13004);
or OR2 (N15773, N15761, N8597);
and AND2 (N15774, N15767, N1633);
nand NAND4 (N15775, N15766, N5607, N13755, N14968);
and AND4 (N15776, N15772, N3922, N6029, N10854);
nand NAND3 (N15777, N15755, N12532, N11080);
nor NOR4 (N15778, N15777, N2179, N12814, N10450);
xor XOR2 (N15779, N15774, N5065);
buf BUF1 (N15780, N15770);
not NOT1 (N15781, N15779);
xor XOR2 (N15782, N15776, N2380);
and AND3 (N15783, N15778, N15162, N14773);
buf BUF1 (N15784, N15781);
xor XOR2 (N15785, N15769, N6828);
nor NOR3 (N15786, N15780, N6096, N7975);
not NOT1 (N15787, N15751);
buf BUF1 (N15788, N15783);
nand NAND2 (N15789, N15764, N15358);
and AND3 (N15790, N15788, N15397, N12645);
nor NOR4 (N15791, N15786, N2287, N2909, N8463);
xor XOR2 (N15792, N15782, N8660);
or OR3 (N15793, N15792, N14340, N9121);
and AND2 (N15794, N15785, N14017);
not NOT1 (N15795, N15771);
xor XOR2 (N15796, N15794, N9307);
xor XOR2 (N15797, N15784, N8115);
nand NAND4 (N15798, N15793, N14441, N12702, N3442);
nand NAND2 (N15799, N15790, N9735);
or OR2 (N15800, N15798, N7130);
buf BUF1 (N15801, N15795);
nand NAND2 (N15802, N15775, N10832);
buf BUF1 (N15803, N15773);
or OR4 (N15804, N15789, N9118, N4188, N104);
nand NAND3 (N15805, N15801, N5590, N6582);
or OR2 (N15806, N15787, N12122);
buf BUF1 (N15807, N15803);
and AND2 (N15808, N15797, N7218);
buf BUF1 (N15809, N15804);
not NOT1 (N15810, N15807);
nor NOR2 (N15811, N15800, N10488);
buf BUF1 (N15812, N15811);
not NOT1 (N15813, N15810);
buf BUF1 (N15814, N15813);
nand NAND4 (N15815, N15796, N15171, N14727, N11035);
not NOT1 (N15816, N15802);
xor XOR2 (N15817, N15815, N3630);
not NOT1 (N15818, N15816);
and AND2 (N15819, N15799, N4013);
or OR3 (N15820, N15809, N11953, N7675);
not NOT1 (N15821, N15820);
buf BUF1 (N15822, N15812);
not NOT1 (N15823, N15808);
xor XOR2 (N15824, N15791, N14848);
nand NAND4 (N15825, N15821, N12720, N946, N11910);
nor NOR3 (N15826, N15818, N9843, N13029);
nor NOR2 (N15827, N15814, N12329);
buf BUF1 (N15828, N15819);
nand NAND3 (N15829, N15825, N11537, N9763);
buf BUF1 (N15830, N15828);
xor XOR2 (N15831, N15824, N14817);
and AND2 (N15832, N15805, N14678);
not NOT1 (N15833, N15826);
nand NAND2 (N15834, N15833, N6676);
xor XOR2 (N15835, N15834, N10980);
or OR3 (N15836, N15829, N5206, N4735);
nand NAND3 (N15837, N15806, N10286, N12271);
nand NAND3 (N15838, N15830, N11859, N11984);
nand NAND3 (N15839, N15832, N360, N10011);
nand NAND3 (N15840, N15817, N6523, N14110);
not NOT1 (N15841, N15840);
nand NAND4 (N15842, N15822, N7310, N12056, N1047);
and AND4 (N15843, N15823, N6938, N7824, N9637);
and AND2 (N15844, N15842, N7885);
buf BUF1 (N15845, N15837);
and AND2 (N15846, N15838, N5984);
nor NOR3 (N15847, N15835, N15325, N14333);
not NOT1 (N15848, N15846);
buf BUF1 (N15849, N15848);
nor NOR4 (N15850, N15839, N6188, N9061, N11215);
nor NOR3 (N15851, N15850, N13071, N3356);
nand NAND2 (N15852, N15831, N2572);
not NOT1 (N15853, N15849);
and AND4 (N15854, N15852, N3737, N7360, N11490);
nor NOR3 (N15855, N15841, N10561, N12226);
or OR4 (N15856, N15847, N374, N11225, N12790);
or OR3 (N15857, N15856, N9923, N11282);
xor XOR2 (N15858, N15845, N423);
nand NAND2 (N15859, N15851, N13480);
not NOT1 (N15860, N15855);
nor NOR2 (N15861, N15844, N7068);
xor XOR2 (N15862, N15861, N10078);
not NOT1 (N15863, N15836);
nand NAND2 (N15864, N15862, N9793);
not NOT1 (N15865, N15854);
or OR2 (N15866, N15858, N740);
nand NAND3 (N15867, N15865, N1745, N228);
not NOT1 (N15868, N15867);
nor NOR3 (N15869, N15827, N7615, N8525);
not NOT1 (N15870, N15863);
and AND2 (N15871, N15866, N7970);
buf BUF1 (N15872, N15857);
not NOT1 (N15873, N15859);
xor XOR2 (N15874, N15853, N15486);
nand NAND2 (N15875, N15868, N11394);
or OR4 (N15876, N15870, N3427, N25, N643);
xor XOR2 (N15877, N15874, N4030);
or OR4 (N15878, N15877, N727, N8951, N6856);
xor XOR2 (N15879, N15878, N1981);
not NOT1 (N15880, N15875);
not NOT1 (N15881, N15876);
nand NAND4 (N15882, N15871, N7333, N7462, N5613);
buf BUF1 (N15883, N15882);
nor NOR3 (N15884, N15872, N9823, N7113);
nor NOR2 (N15885, N15843, N10917);
and AND3 (N15886, N15881, N5992, N15169);
or OR2 (N15887, N15884, N2572);
nand NAND3 (N15888, N15879, N12382, N1562);
nor NOR4 (N15889, N15883, N290, N7805, N14429);
or OR4 (N15890, N15885, N1835, N11647, N2664);
or OR2 (N15891, N15860, N14303);
not NOT1 (N15892, N15873);
buf BUF1 (N15893, N15891);
or OR2 (N15894, N15889, N1293);
and AND3 (N15895, N15890, N8159, N7196);
or OR4 (N15896, N15886, N953, N1236, N92);
nand NAND4 (N15897, N15896, N10582, N9745, N2367);
nor NOR2 (N15898, N15880, N691);
or OR4 (N15899, N15893, N15657, N8807, N7283);
buf BUF1 (N15900, N15894);
and AND4 (N15901, N15895, N12570, N2016, N4580);
buf BUF1 (N15902, N15900);
not NOT1 (N15903, N15897);
or OR4 (N15904, N15869, N2602, N3209, N13059);
not NOT1 (N15905, N15898);
buf BUF1 (N15906, N15902);
buf BUF1 (N15907, N15906);
and AND2 (N15908, N15864, N6407);
or OR3 (N15909, N15901, N15112, N4806);
xor XOR2 (N15910, N15887, N6561);
nand NAND3 (N15911, N15908, N13006, N1361);
buf BUF1 (N15912, N15892);
xor XOR2 (N15913, N15912, N497);
nand NAND3 (N15914, N15909, N13084, N4243);
nand NAND2 (N15915, N15911, N3452);
buf BUF1 (N15916, N15905);
buf BUF1 (N15917, N15910);
nor NOR2 (N15918, N15916, N6210);
and AND2 (N15919, N15904, N11133);
nand NAND4 (N15920, N15917, N5743, N447, N1359);
and AND3 (N15921, N15919, N11080, N11776);
xor XOR2 (N15922, N15921, N1527);
xor XOR2 (N15923, N15918, N3335);
xor XOR2 (N15924, N15913, N3418);
not NOT1 (N15925, N15903);
or OR4 (N15926, N15888, N6222, N1513, N14015);
or OR3 (N15927, N15914, N10772, N3718);
nand NAND2 (N15928, N15924, N10351);
buf BUF1 (N15929, N15926);
not NOT1 (N15930, N15922);
nor NOR4 (N15931, N15915, N13318, N10201, N10183);
not NOT1 (N15932, N15923);
or OR3 (N15933, N15930, N8742, N14681);
nor NOR4 (N15934, N15925, N15764, N5751, N8626);
or OR2 (N15935, N15934, N3902);
and AND2 (N15936, N15907, N11931);
not NOT1 (N15937, N15932);
or OR4 (N15938, N15920, N14137, N13183, N6011);
buf BUF1 (N15939, N15931);
buf BUF1 (N15940, N15939);
xor XOR2 (N15941, N15940, N8882);
xor XOR2 (N15942, N15933, N10049);
buf BUF1 (N15943, N15936);
nand NAND3 (N15944, N15941, N11296, N11273);
and AND3 (N15945, N15938, N6685, N15000);
xor XOR2 (N15946, N15942, N65);
buf BUF1 (N15947, N15945);
nand NAND3 (N15948, N15943, N8197, N2343);
or OR3 (N15949, N15944, N73, N806);
buf BUF1 (N15950, N15928);
xor XOR2 (N15951, N15935, N11599);
and AND4 (N15952, N15948, N10205, N4007, N7326);
or OR2 (N15953, N15899, N2347);
buf BUF1 (N15954, N15950);
or OR4 (N15955, N15929, N13366, N14687, N1206);
not NOT1 (N15956, N15955);
buf BUF1 (N15957, N15946);
nand NAND4 (N15958, N15954, N14587, N9539, N6961);
nand NAND4 (N15959, N15957, N9249, N1380, N371);
or OR3 (N15960, N15927, N9466, N2541);
nand NAND3 (N15961, N15953, N14079, N4151);
buf BUF1 (N15962, N15947);
or OR2 (N15963, N15959, N4597);
and AND3 (N15964, N15958, N6285, N15155);
and AND4 (N15965, N15949, N7985, N2596, N10459);
nor NOR3 (N15966, N15961, N15013, N4303);
nor NOR4 (N15967, N15952, N10595, N5293, N14869);
and AND3 (N15968, N15962, N7051, N2035);
nor NOR3 (N15969, N15937, N15327, N4252);
xor XOR2 (N15970, N15960, N5066);
buf BUF1 (N15971, N15965);
and AND4 (N15972, N15951, N3544, N12145, N3664);
buf BUF1 (N15973, N15964);
nor NOR4 (N15974, N15970, N2215, N7959, N15944);
not NOT1 (N15975, N15969);
or OR4 (N15976, N15975, N3936, N363, N3038);
nor NOR4 (N15977, N15967, N4920, N6970, N8594);
nor NOR4 (N15978, N15972, N11522, N8789, N8075);
not NOT1 (N15979, N15968);
nor NOR3 (N15980, N15976, N3400, N28);
nor NOR3 (N15981, N15977, N7012, N15276);
not NOT1 (N15982, N15980);
nand NAND2 (N15983, N15966, N2615);
not NOT1 (N15984, N15979);
nand NAND4 (N15985, N15971, N3354, N4329, N6619);
or OR4 (N15986, N15981, N11320, N5841, N14581);
or OR3 (N15987, N15956, N10464, N6986);
and AND2 (N15988, N15985, N218);
and AND2 (N15989, N15983, N14173);
nand NAND3 (N15990, N15986, N13914, N3671);
xor XOR2 (N15991, N15988, N9410);
not NOT1 (N15992, N15982);
or OR4 (N15993, N15990, N9637, N2094, N5146);
and AND4 (N15994, N15973, N13097, N13946, N2163);
buf BUF1 (N15995, N15987);
nor NOR3 (N15996, N15995, N9040, N11993);
buf BUF1 (N15997, N15992);
buf BUF1 (N15998, N15978);
nand NAND2 (N15999, N15994, N7023);
xor XOR2 (N16000, N15999, N1623);
nor NOR3 (N16001, N15993, N14569, N2200);
xor XOR2 (N16002, N15989, N454);
xor XOR2 (N16003, N15997, N889);
xor XOR2 (N16004, N16001, N4335);
nand NAND2 (N16005, N15996, N10804);
nand NAND4 (N16006, N15984, N5007, N9993, N605);
or OR3 (N16007, N16005, N4926, N9809);
or OR4 (N16008, N16006, N9193, N971, N1165);
not NOT1 (N16009, N16002);
not NOT1 (N16010, N15998);
or OR4 (N16011, N16000, N378, N6883, N6238);
nor NOR3 (N16012, N15974, N12419, N6329);
and AND2 (N16013, N15991, N2678);
not NOT1 (N16014, N16008);
nand NAND3 (N16015, N16010, N9247, N4563);
endmodule