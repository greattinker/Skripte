// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N2517,N2510,N2499,N2513,N2504,N2522,N2451,N2521,N2519,N2523;

and AND4 (N24, N17, N19, N23, N9);
nor NOR2 (N25, N5, N9);
nor NOR4 (N26, N21, N7, N16, N18);
xor XOR2 (N27, N21, N9);
nor NOR3 (N28, N4, N3, N16);
not NOT1 (N29, N3);
or OR4 (N30, N10, N19, N18, N2);
not NOT1 (N31, N19);
buf BUF1 (N32, N4);
nand NAND3 (N33, N17, N2, N27);
nand NAND2 (N34, N31, N27);
buf BUF1 (N35, N1);
nand NAND4 (N36, N28, N24, N7, N29);
nor NOR4 (N37, N31, N22, N20, N10);
nand NAND2 (N38, N23, N11);
and AND4 (N39, N26, N21, N34, N38);
nand NAND3 (N40, N20, N23, N24);
nor NOR4 (N41, N38, N21, N18, N1);
or OR4 (N42, N35, N33, N26, N29);
not NOT1 (N43, N7);
not NOT1 (N44, N32);
buf BUF1 (N45, N39);
and AND2 (N46, N44, N19);
nand NAND4 (N47, N41, N29, N37, N16);
nand NAND2 (N48, N44, N34);
buf BUF1 (N49, N36);
nand NAND2 (N50, N47, N19);
and AND2 (N51, N30, N47);
nand NAND3 (N52, N51, N30, N43);
xor XOR2 (N53, N27, N21);
nand NAND3 (N54, N45, N21, N6);
or OR4 (N55, N50, N10, N54, N3);
xor XOR2 (N56, N39, N21);
and AND2 (N57, N48, N39);
nor NOR2 (N58, N40, N48);
or OR3 (N59, N52, N3, N22);
nor NOR2 (N60, N56, N54);
nor NOR4 (N61, N49, N35, N17, N48);
not NOT1 (N62, N55);
not NOT1 (N63, N61);
xor XOR2 (N64, N59, N5);
nor NOR2 (N65, N46, N47);
and AND3 (N66, N65, N39, N4);
xor XOR2 (N67, N60, N51);
xor XOR2 (N68, N57, N22);
buf BUF1 (N69, N53);
and AND3 (N70, N69, N61, N69);
nor NOR2 (N71, N68, N21);
and AND4 (N72, N62, N50, N19, N40);
and AND4 (N73, N63, N15, N11, N22);
or OR3 (N74, N72, N25, N5);
or OR3 (N75, N11, N52, N18);
and AND4 (N76, N74, N20, N3, N18);
nor NOR4 (N77, N67, N63, N26, N22);
nor NOR4 (N78, N73, N53, N30, N76);
not NOT1 (N79, N21);
and AND4 (N80, N75, N29, N6, N9);
xor XOR2 (N81, N58, N11);
xor XOR2 (N82, N77, N78);
not NOT1 (N83, N12);
xor XOR2 (N84, N83, N50);
or OR3 (N85, N66, N68, N75);
not NOT1 (N86, N81);
nor NOR3 (N87, N71, N21, N35);
and AND4 (N88, N85, N71, N75, N82);
xor XOR2 (N89, N32, N68);
and AND3 (N90, N79, N49, N12);
or OR3 (N91, N90, N25, N1);
or OR3 (N92, N89, N35, N46);
xor XOR2 (N93, N80, N59);
not NOT1 (N94, N92);
nor NOR3 (N95, N42, N70, N38);
nor NOR4 (N96, N81, N32, N20, N50);
and AND2 (N97, N94, N58);
not NOT1 (N98, N86);
nand NAND4 (N99, N93, N92, N94, N48);
not NOT1 (N100, N87);
nand NAND2 (N101, N91, N84);
nor NOR3 (N102, N31, N73, N14);
nor NOR2 (N103, N88, N42);
buf BUF1 (N104, N102);
nor NOR2 (N105, N100, N48);
nor NOR4 (N106, N97, N20, N67, N75);
nand NAND3 (N107, N96, N37, N64);
or OR2 (N108, N46, N98);
and AND2 (N109, N86, N55);
nor NOR3 (N110, N105, N37, N31);
nor NOR4 (N111, N95, N41, N29, N78);
and AND3 (N112, N111, N40, N6);
nor NOR2 (N113, N99, N15);
or OR2 (N114, N106, N13);
or OR4 (N115, N114, N87, N55, N30);
or OR2 (N116, N101, N75);
nand NAND3 (N117, N116, N14, N20);
nand NAND4 (N118, N115, N92, N109, N69);
or OR3 (N119, N15, N60, N75);
buf BUF1 (N120, N112);
nor NOR4 (N121, N118, N75, N19, N14);
nor NOR2 (N122, N120, N39);
xor XOR2 (N123, N117, N61);
buf BUF1 (N124, N119);
nor NOR2 (N125, N121, N62);
nor NOR3 (N126, N125, N104, N121);
xor XOR2 (N127, N66, N88);
and AND4 (N128, N113, N33, N48, N100);
nand NAND3 (N129, N110, N51, N83);
not NOT1 (N130, N108);
xor XOR2 (N131, N103, N58);
and AND2 (N132, N107, N63);
and AND2 (N133, N127, N33);
nand NAND2 (N134, N128, N23);
or OR3 (N135, N130, N66, N44);
and AND2 (N136, N133, N11);
xor XOR2 (N137, N134, N86);
not NOT1 (N138, N132);
not NOT1 (N139, N136);
nand NAND4 (N140, N138, N31, N135, N59);
buf BUF1 (N141, N6);
buf BUF1 (N142, N126);
nand NAND3 (N143, N137, N72, N133);
buf BUF1 (N144, N142);
or OR4 (N145, N131, N26, N8, N109);
and AND2 (N146, N124, N131);
or OR4 (N147, N122, N85, N15, N98);
not NOT1 (N148, N139);
nand NAND4 (N149, N140, N18, N61, N61);
buf BUF1 (N150, N144);
buf BUF1 (N151, N148);
nand NAND3 (N152, N146, N110, N22);
xor XOR2 (N153, N143, N63);
nand NAND3 (N154, N150, N29, N95);
nor NOR4 (N155, N147, N130, N24, N5);
buf BUF1 (N156, N153);
and AND4 (N157, N123, N83, N118, N19);
xor XOR2 (N158, N157, N66);
nor NOR2 (N159, N151, N94);
nor NOR4 (N160, N145, N77, N100, N45);
nand NAND4 (N161, N149, N68, N44, N154);
xor XOR2 (N162, N147, N29);
not NOT1 (N163, N141);
nor NOR2 (N164, N161, N70);
buf BUF1 (N165, N159);
buf BUF1 (N166, N156);
buf BUF1 (N167, N158);
or OR2 (N168, N164, N4);
or OR2 (N169, N165, N42);
nand NAND3 (N170, N168, N13, N25);
nand NAND3 (N171, N166, N88, N55);
xor XOR2 (N172, N169, N170);
and AND3 (N173, N95, N12, N38);
or OR4 (N174, N129, N98, N60, N24);
buf BUF1 (N175, N171);
not NOT1 (N176, N163);
nor NOR4 (N177, N155, N119, N166, N52);
xor XOR2 (N178, N162, N66);
or OR2 (N179, N172, N143);
nand NAND4 (N180, N177, N41, N105, N52);
buf BUF1 (N181, N175);
or OR4 (N182, N173, N122, N159, N23);
nand NAND3 (N183, N174, N135, N149);
and AND3 (N184, N152, N10, N78);
buf BUF1 (N185, N178);
and AND2 (N186, N183, N173);
and AND3 (N187, N180, N74, N149);
nor NOR3 (N188, N184, N44, N171);
nand NAND4 (N189, N176, N10, N135, N156);
and AND2 (N190, N167, N2);
not NOT1 (N191, N187);
nor NOR2 (N192, N182, N124);
nor NOR2 (N193, N189, N157);
nand NAND4 (N194, N160, N186, N187, N177);
nor NOR3 (N195, N21, N32, N41);
xor XOR2 (N196, N185, N167);
nor NOR4 (N197, N181, N154, N87, N58);
nor NOR3 (N198, N179, N4, N5);
not NOT1 (N199, N196);
nand NAND3 (N200, N197, N99, N166);
not NOT1 (N201, N188);
buf BUF1 (N202, N199);
and AND3 (N203, N201, N142, N186);
and AND4 (N204, N202, N88, N103, N88);
or OR3 (N205, N200, N48, N67);
and AND3 (N206, N205, N62, N123);
not NOT1 (N207, N195);
nor NOR2 (N208, N207, N97);
buf BUF1 (N209, N193);
nand NAND4 (N210, N204, N109, N199, N7);
nand NAND3 (N211, N203, N137, N203);
not NOT1 (N212, N198);
and AND2 (N213, N212, N200);
or OR2 (N214, N208, N46);
buf BUF1 (N215, N191);
nand NAND2 (N216, N213, N80);
not NOT1 (N217, N209);
nor NOR4 (N218, N192, N164, N91, N119);
or OR2 (N219, N214, N63);
xor XOR2 (N220, N190, N102);
buf BUF1 (N221, N217);
and AND3 (N222, N219, N10, N129);
nor NOR4 (N223, N211, N168, N61, N151);
not NOT1 (N224, N194);
nand NAND4 (N225, N224, N172, N215, N172);
nor NOR3 (N226, N41, N107, N108);
xor XOR2 (N227, N226, N139);
xor XOR2 (N228, N221, N197);
and AND3 (N229, N220, N80, N140);
xor XOR2 (N230, N225, N211);
nand NAND4 (N231, N223, N118, N209, N161);
nor NOR4 (N232, N227, N43, N113, N161);
and AND2 (N233, N231, N117);
nand NAND2 (N234, N222, N159);
nor NOR4 (N235, N206, N163, N74, N34);
nand NAND2 (N236, N234, N37);
xor XOR2 (N237, N216, N132);
xor XOR2 (N238, N232, N34);
nand NAND2 (N239, N237, N27);
xor XOR2 (N240, N238, N82);
and AND2 (N241, N210, N65);
xor XOR2 (N242, N240, N63);
not NOT1 (N243, N228);
not NOT1 (N244, N233);
and AND3 (N245, N239, N32, N27);
or OR3 (N246, N230, N224, N68);
nor NOR2 (N247, N235, N99);
buf BUF1 (N248, N241);
not NOT1 (N249, N247);
nor NOR2 (N250, N249, N216);
nor NOR2 (N251, N245, N164);
xor XOR2 (N252, N243, N189);
nand NAND2 (N253, N236, N104);
nand NAND2 (N254, N250, N165);
xor XOR2 (N255, N246, N73);
nand NAND4 (N256, N244, N244, N111, N26);
buf BUF1 (N257, N253);
nor NOR2 (N258, N257, N117);
xor XOR2 (N259, N256, N84);
xor XOR2 (N260, N259, N118);
buf BUF1 (N261, N255);
xor XOR2 (N262, N261, N102);
and AND3 (N263, N242, N86, N42);
xor XOR2 (N264, N252, N255);
nand NAND3 (N265, N229, N198, N13);
or OR3 (N266, N258, N127, N238);
not NOT1 (N267, N248);
not NOT1 (N268, N264);
and AND4 (N269, N218, N35, N148, N34);
nor NOR2 (N270, N269, N107);
buf BUF1 (N271, N262);
nand NAND4 (N272, N260, N171, N183, N258);
buf BUF1 (N273, N270);
and AND2 (N274, N266, N12);
nor NOR3 (N275, N273, N16, N3);
nor NOR3 (N276, N272, N181, N3);
nor NOR4 (N277, N254, N101, N87, N160);
buf BUF1 (N278, N267);
and AND3 (N279, N278, N243, N228);
or OR2 (N280, N251, N197);
xor XOR2 (N281, N280, N142);
nor NOR4 (N282, N268, N176, N266, N11);
nand NAND4 (N283, N279, N268, N156, N206);
or OR3 (N284, N281, N135, N108);
nand NAND4 (N285, N283, N33, N166, N76);
nor NOR2 (N286, N263, N131);
xor XOR2 (N287, N265, N113);
not NOT1 (N288, N284);
not NOT1 (N289, N271);
xor XOR2 (N290, N277, N178);
nand NAND4 (N291, N275, N171, N116, N144);
not NOT1 (N292, N274);
xor XOR2 (N293, N289, N222);
xor XOR2 (N294, N276, N83);
nor NOR3 (N295, N282, N77, N260);
nor NOR3 (N296, N294, N81, N53);
or OR3 (N297, N293, N287, N22);
nor NOR3 (N298, N10, N113, N221);
and AND3 (N299, N297, N208, N114);
nor NOR3 (N300, N290, N72, N192);
not NOT1 (N301, N300);
not NOT1 (N302, N285);
nor NOR2 (N303, N292, N138);
not NOT1 (N304, N295);
not NOT1 (N305, N304);
not NOT1 (N306, N299);
xor XOR2 (N307, N306, N265);
xor XOR2 (N308, N298, N9);
or OR2 (N309, N305, N199);
and AND3 (N310, N307, N213, N145);
and AND4 (N311, N303, N185, N25, N48);
or OR2 (N312, N288, N204);
and AND4 (N313, N302, N28, N104, N1);
buf BUF1 (N314, N310);
nor NOR4 (N315, N311, N13, N80, N250);
nand NAND2 (N316, N296, N263);
nor NOR2 (N317, N286, N255);
not NOT1 (N318, N317);
and AND4 (N319, N309, N11, N84, N249);
not NOT1 (N320, N319);
nand NAND3 (N321, N301, N234, N203);
not NOT1 (N322, N313);
nor NOR2 (N323, N316, N277);
or OR3 (N324, N322, N111, N282);
not NOT1 (N325, N314);
xor XOR2 (N326, N325, N137);
or OR4 (N327, N321, N299, N75, N83);
and AND3 (N328, N308, N171, N263);
and AND3 (N329, N327, N116, N208);
or OR2 (N330, N323, N219);
and AND2 (N331, N328, N72);
buf BUF1 (N332, N315);
buf BUF1 (N333, N318);
and AND3 (N334, N326, N141, N246);
nand NAND2 (N335, N332, N207);
and AND3 (N336, N331, N320, N138);
or OR3 (N337, N76, N284, N185);
nand NAND2 (N338, N334, N135);
nor NOR3 (N339, N329, N182, N136);
xor XOR2 (N340, N333, N181);
xor XOR2 (N341, N335, N285);
buf BUF1 (N342, N337);
xor XOR2 (N343, N330, N141);
and AND2 (N344, N312, N165);
or OR3 (N345, N342, N187, N223);
nor NOR2 (N346, N336, N219);
buf BUF1 (N347, N345);
nor NOR4 (N348, N338, N265, N7, N198);
nand NAND4 (N349, N344, N238, N195, N147);
not NOT1 (N350, N291);
nand NAND2 (N351, N348, N265);
not NOT1 (N352, N341);
buf BUF1 (N353, N340);
xor XOR2 (N354, N351, N159);
nand NAND3 (N355, N349, N213, N208);
not NOT1 (N356, N353);
not NOT1 (N357, N324);
xor XOR2 (N358, N352, N118);
xor XOR2 (N359, N358, N156);
nand NAND4 (N360, N343, N325, N156, N135);
nand NAND4 (N361, N359, N263, N18, N313);
xor XOR2 (N362, N339, N193);
or OR2 (N363, N350, N131);
or OR3 (N364, N362, N89, N202);
or OR3 (N365, N361, N126, N267);
and AND2 (N366, N357, N161);
or OR3 (N367, N366, N332, N171);
buf BUF1 (N368, N363);
buf BUF1 (N369, N364);
nand NAND2 (N370, N369, N246);
and AND4 (N371, N367, N175, N345, N134);
or OR2 (N372, N355, N213);
not NOT1 (N373, N356);
or OR2 (N374, N365, N281);
not NOT1 (N375, N346);
xor XOR2 (N376, N370, N369);
xor XOR2 (N377, N372, N4);
nor NOR2 (N378, N376, N73);
and AND2 (N379, N368, N189);
nor NOR4 (N380, N371, N285, N170, N174);
and AND4 (N381, N377, N296, N213, N63);
nand NAND4 (N382, N379, N143, N267, N343);
buf BUF1 (N383, N382);
buf BUF1 (N384, N373);
not NOT1 (N385, N375);
and AND4 (N386, N354, N229, N304, N86);
and AND4 (N387, N347, N155, N204, N256);
nand NAND3 (N388, N360, N149, N42);
xor XOR2 (N389, N378, N101);
nand NAND2 (N390, N374, N36);
and AND2 (N391, N388, N333);
not NOT1 (N392, N390);
not NOT1 (N393, N383);
nand NAND3 (N394, N381, N159, N202);
not NOT1 (N395, N384);
not NOT1 (N396, N386);
buf BUF1 (N397, N394);
nor NOR2 (N398, N385, N25);
nor NOR4 (N399, N397, N343, N201, N44);
nand NAND3 (N400, N392, N191, N181);
buf BUF1 (N401, N400);
xor XOR2 (N402, N396, N263);
nand NAND4 (N403, N399, N224, N345, N286);
not NOT1 (N404, N402);
and AND2 (N405, N404, N195);
xor XOR2 (N406, N398, N163);
not NOT1 (N407, N380);
nand NAND4 (N408, N406, N358, N367, N69);
not NOT1 (N409, N389);
xor XOR2 (N410, N393, N377);
xor XOR2 (N411, N401, N362);
buf BUF1 (N412, N395);
or OR2 (N413, N408, N211);
nor NOR2 (N414, N409, N174);
nand NAND3 (N415, N387, N196, N183);
nor NOR2 (N416, N411, N357);
and AND4 (N417, N413, N186, N75, N87);
and AND4 (N418, N415, N4, N173, N292);
buf BUF1 (N419, N416);
nand NAND3 (N420, N405, N127, N147);
buf BUF1 (N421, N418);
nand NAND4 (N422, N419, N151, N380, N260);
xor XOR2 (N423, N410, N138);
not NOT1 (N424, N412);
xor XOR2 (N425, N424, N85);
buf BUF1 (N426, N417);
nand NAND2 (N427, N414, N139);
buf BUF1 (N428, N421);
not NOT1 (N429, N425);
xor XOR2 (N430, N403, N419);
nand NAND2 (N431, N430, N168);
buf BUF1 (N432, N420);
and AND3 (N433, N426, N5, N98);
nand NAND3 (N434, N422, N371, N322);
not NOT1 (N435, N427);
not NOT1 (N436, N435);
or OR2 (N437, N429, N407);
buf BUF1 (N438, N414);
nor NOR3 (N439, N433, N381, N382);
or OR3 (N440, N428, N271, N398);
and AND4 (N441, N440, N399, N363, N236);
nand NAND3 (N442, N439, N122, N432);
or OR3 (N443, N416, N82, N56);
not NOT1 (N444, N436);
buf BUF1 (N445, N391);
or OR3 (N446, N438, N245, N128);
buf BUF1 (N447, N444);
not NOT1 (N448, N443);
nand NAND3 (N449, N437, N401, N12);
nor NOR2 (N450, N445, N357);
buf BUF1 (N451, N446);
and AND3 (N452, N442, N449, N448);
or OR4 (N453, N211, N430, N305, N58);
nor NOR2 (N454, N253, N285);
and AND3 (N455, N452, N376, N362);
and AND4 (N456, N431, N176, N64, N432);
and AND2 (N457, N454, N364);
nor NOR2 (N458, N453, N255);
nand NAND4 (N459, N450, N335, N278, N183);
not NOT1 (N460, N441);
nor NOR2 (N461, N460, N371);
buf BUF1 (N462, N423);
not NOT1 (N463, N455);
buf BUF1 (N464, N447);
nand NAND4 (N465, N462, N269, N197, N314);
nor NOR2 (N466, N465, N203);
not NOT1 (N467, N466);
and AND4 (N468, N451, N466, N313, N250);
or OR2 (N469, N434, N379);
not NOT1 (N470, N457);
nand NAND4 (N471, N463, N152, N374, N192);
and AND3 (N472, N459, N56, N36);
nand NAND2 (N473, N458, N414);
buf BUF1 (N474, N472);
nor NOR3 (N475, N471, N436, N140);
buf BUF1 (N476, N469);
not NOT1 (N477, N476);
not NOT1 (N478, N477);
nand NAND4 (N479, N468, N422, N148, N191);
nand NAND3 (N480, N461, N473, N62);
or OR3 (N481, N216, N76, N261);
and AND3 (N482, N467, N282, N75);
not NOT1 (N483, N482);
buf BUF1 (N484, N483);
or OR2 (N485, N474, N173);
or OR3 (N486, N470, N481, N393);
nand NAND3 (N487, N237, N4, N482);
not NOT1 (N488, N487);
or OR4 (N489, N486, N125, N462, N59);
nor NOR3 (N490, N475, N89, N231);
not NOT1 (N491, N456);
buf BUF1 (N492, N488);
nand NAND4 (N493, N492, N389, N492, N344);
not NOT1 (N494, N489);
and AND4 (N495, N491, N31, N254, N199);
or OR2 (N496, N478, N158);
nor NOR3 (N497, N494, N428, N269);
not NOT1 (N498, N496);
or OR4 (N499, N480, N4, N68, N104);
or OR4 (N500, N499, N86, N260, N134);
xor XOR2 (N501, N497, N466);
nor NOR2 (N502, N464, N41);
and AND3 (N503, N479, N77, N327);
or OR4 (N504, N498, N413, N341, N330);
not NOT1 (N505, N484);
or OR2 (N506, N504, N451);
nand NAND4 (N507, N485, N477, N116, N250);
or OR4 (N508, N505, N12, N349, N378);
nand NAND3 (N509, N493, N199, N252);
and AND2 (N510, N500, N231);
nor NOR2 (N511, N508, N502);
xor XOR2 (N512, N423, N59);
not NOT1 (N513, N510);
nand NAND4 (N514, N503, N422, N320, N353);
buf BUF1 (N515, N511);
nand NAND4 (N516, N513, N477, N148, N428);
xor XOR2 (N517, N506, N36);
xor XOR2 (N518, N490, N328);
nor NOR3 (N519, N507, N172, N249);
nand NAND4 (N520, N495, N275, N361, N64);
not NOT1 (N521, N514);
or OR4 (N522, N519, N421, N348, N89);
nand NAND4 (N523, N516, N227, N47, N351);
and AND2 (N524, N522, N280);
or OR2 (N525, N517, N80);
buf BUF1 (N526, N515);
nand NAND4 (N527, N524, N491, N510, N70);
nor NOR2 (N528, N527, N53);
xor XOR2 (N529, N501, N317);
or OR3 (N530, N526, N214, N421);
nor NOR3 (N531, N518, N463, N243);
not NOT1 (N532, N531);
nand NAND3 (N533, N525, N338, N506);
nor NOR2 (N534, N532, N214);
or OR2 (N535, N533, N324);
or OR4 (N536, N535, N29, N505, N447);
xor XOR2 (N537, N523, N2);
buf BUF1 (N538, N509);
not NOT1 (N539, N534);
and AND2 (N540, N537, N366);
or OR3 (N541, N520, N440, N399);
and AND4 (N542, N540, N395, N458, N287);
xor XOR2 (N543, N539, N6);
nand NAND4 (N544, N528, N297, N381, N327);
and AND2 (N545, N530, N152);
or OR4 (N546, N536, N541, N23, N532);
and AND2 (N547, N498, N43);
buf BUF1 (N548, N512);
nor NOR3 (N549, N545, N436, N21);
xor XOR2 (N550, N529, N217);
nand NAND4 (N551, N550, N65, N529, N76);
nand NAND4 (N552, N549, N230, N429, N52);
not NOT1 (N553, N543);
xor XOR2 (N554, N521, N159);
or OR3 (N555, N552, N478, N223);
xor XOR2 (N556, N538, N506);
and AND4 (N557, N553, N124, N482, N2);
nand NAND4 (N558, N546, N214, N335, N201);
not NOT1 (N559, N551);
or OR4 (N560, N547, N29, N168, N486);
nor NOR2 (N561, N555, N414);
not NOT1 (N562, N542);
not NOT1 (N563, N556);
buf BUF1 (N564, N562);
or OR3 (N565, N554, N398, N290);
nand NAND3 (N566, N544, N129, N287);
nand NAND4 (N567, N559, N154, N368, N134);
not NOT1 (N568, N567);
not NOT1 (N569, N560);
or OR4 (N570, N568, N472, N549, N441);
buf BUF1 (N571, N569);
or OR2 (N572, N565, N462);
and AND3 (N573, N563, N82, N179);
xor XOR2 (N574, N572, N486);
buf BUF1 (N575, N570);
xor XOR2 (N576, N571, N99);
not NOT1 (N577, N558);
nor NOR3 (N578, N548, N46, N568);
nor NOR2 (N579, N574, N474);
buf BUF1 (N580, N573);
and AND2 (N581, N576, N292);
and AND2 (N582, N577, N200);
and AND4 (N583, N580, N252, N522, N124);
and AND2 (N584, N566, N194);
nand NAND2 (N585, N564, N528);
or OR3 (N586, N579, N338, N96);
buf BUF1 (N587, N557);
not NOT1 (N588, N581);
nand NAND4 (N589, N584, N575, N483, N3);
or OR4 (N590, N568, N502, N172, N106);
buf BUF1 (N591, N588);
nor NOR3 (N592, N591, N141, N445);
nor NOR2 (N593, N592, N301);
nand NAND2 (N594, N587, N98);
xor XOR2 (N595, N561, N461);
not NOT1 (N596, N595);
not NOT1 (N597, N590);
and AND4 (N598, N583, N336, N187, N432);
or OR3 (N599, N597, N432, N73);
nor NOR4 (N600, N586, N112, N33, N567);
or OR4 (N601, N578, N188, N268, N23);
and AND3 (N602, N598, N85, N365);
and AND4 (N603, N600, N211, N499, N480);
not NOT1 (N604, N599);
or OR3 (N605, N601, N454, N415);
nor NOR2 (N606, N593, N27);
xor XOR2 (N607, N606, N127);
or OR3 (N608, N607, N409, N441);
xor XOR2 (N609, N582, N85);
or OR4 (N610, N608, N435, N405, N93);
xor XOR2 (N611, N603, N91);
not NOT1 (N612, N585);
buf BUF1 (N613, N596);
nand NAND3 (N614, N589, N151, N373);
not NOT1 (N615, N594);
nand NAND3 (N616, N615, N278, N24);
nor NOR2 (N617, N609, N239);
not NOT1 (N618, N614);
xor XOR2 (N619, N618, N447);
or OR2 (N620, N602, N134);
or OR2 (N621, N611, N264);
and AND4 (N622, N620, N537, N220, N66);
not NOT1 (N623, N610);
xor XOR2 (N624, N619, N565);
nor NOR2 (N625, N616, N493);
and AND2 (N626, N604, N477);
xor XOR2 (N627, N605, N317);
not NOT1 (N628, N621);
xor XOR2 (N629, N622, N477);
or OR4 (N630, N623, N449, N129, N383);
not NOT1 (N631, N625);
nor NOR4 (N632, N617, N152, N385, N99);
nor NOR4 (N633, N624, N71, N495, N151);
buf BUF1 (N634, N613);
nand NAND3 (N635, N630, N184, N391);
or OR2 (N636, N626, N173);
and AND3 (N637, N612, N209, N520);
xor XOR2 (N638, N632, N472);
nor NOR3 (N639, N635, N517, N523);
and AND2 (N640, N636, N137);
not NOT1 (N641, N629);
buf BUF1 (N642, N641);
or OR4 (N643, N633, N125, N14, N99);
not NOT1 (N644, N637);
and AND3 (N645, N640, N606, N491);
not NOT1 (N646, N638);
and AND3 (N647, N644, N430, N340);
buf BUF1 (N648, N628);
or OR4 (N649, N648, N603, N97, N356);
nand NAND3 (N650, N634, N410, N536);
and AND4 (N651, N631, N327, N554, N294);
or OR3 (N652, N650, N434, N632);
and AND2 (N653, N627, N644);
and AND2 (N654, N646, N246);
not NOT1 (N655, N649);
or OR4 (N656, N651, N384, N216, N265);
buf BUF1 (N657, N639);
not NOT1 (N658, N652);
nand NAND4 (N659, N645, N483, N600, N494);
and AND4 (N660, N655, N28, N25, N61);
nand NAND4 (N661, N658, N540, N215, N79);
xor XOR2 (N662, N643, N22);
and AND3 (N663, N659, N580, N497);
or OR3 (N664, N653, N478, N136);
not NOT1 (N665, N657);
and AND3 (N666, N654, N179, N565);
nand NAND3 (N667, N664, N147, N164);
buf BUF1 (N668, N666);
nand NAND2 (N669, N667, N356);
not NOT1 (N670, N662);
xor XOR2 (N671, N656, N296);
nor NOR4 (N672, N660, N142, N410, N390);
or OR2 (N673, N642, N672);
not NOT1 (N674, N110);
buf BUF1 (N675, N674);
buf BUF1 (N676, N671);
buf BUF1 (N677, N668);
or OR3 (N678, N670, N72, N94);
buf BUF1 (N679, N663);
or OR4 (N680, N661, N171, N298, N274);
or OR3 (N681, N676, N431, N567);
nor NOR3 (N682, N665, N594, N610);
or OR2 (N683, N673, N385);
buf BUF1 (N684, N682);
nor NOR4 (N685, N669, N195, N315, N580);
nand NAND2 (N686, N647, N455);
nor NOR3 (N687, N684, N300, N283);
or OR2 (N688, N675, N603);
buf BUF1 (N689, N685);
xor XOR2 (N690, N688, N249);
and AND3 (N691, N687, N55, N97);
nand NAND3 (N692, N677, N328, N371);
buf BUF1 (N693, N686);
nand NAND2 (N694, N693, N430);
and AND4 (N695, N678, N410, N145, N107);
nor NOR3 (N696, N694, N652, N395);
nor NOR3 (N697, N695, N417, N149);
nor NOR4 (N698, N683, N463, N161, N128);
xor XOR2 (N699, N698, N469);
not NOT1 (N700, N691);
xor XOR2 (N701, N697, N375);
buf BUF1 (N702, N701);
not NOT1 (N703, N699);
and AND2 (N704, N689, N26);
nor NOR2 (N705, N692, N683);
xor XOR2 (N706, N704, N179);
or OR2 (N707, N705, N10);
not NOT1 (N708, N681);
nor NOR2 (N709, N700, N375);
buf BUF1 (N710, N702);
not NOT1 (N711, N690);
buf BUF1 (N712, N709);
nand NAND4 (N713, N712, N496, N369, N9);
not NOT1 (N714, N706);
or OR3 (N715, N711, N410, N67);
and AND3 (N716, N708, N606, N468);
nor NOR2 (N717, N714, N325);
or OR3 (N718, N680, N202, N619);
nor NOR4 (N719, N715, N147, N335, N637);
xor XOR2 (N720, N717, N458);
not NOT1 (N721, N679);
and AND2 (N722, N721, N314);
nand NAND4 (N723, N703, N617, N322, N665);
not NOT1 (N724, N722);
or OR2 (N725, N718, N367);
or OR3 (N726, N724, N517, N7);
or OR3 (N727, N707, N163, N64);
and AND2 (N728, N723, N360);
or OR2 (N729, N713, N670);
not NOT1 (N730, N725);
or OR4 (N731, N727, N589, N432, N345);
or OR3 (N732, N720, N393, N314);
or OR2 (N733, N719, N313);
nand NAND3 (N734, N726, N139, N287);
and AND3 (N735, N733, N637, N436);
and AND2 (N736, N731, N96);
xor XOR2 (N737, N729, N158);
buf BUF1 (N738, N716);
nand NAND2 (N739, N730, N649);
buf BUF1 (N740, N732);
or OR3 (N741, N736, N265, N110);
nand NAND3 (N742, N734, N273, N711);
nand NAND4 (N743, N739, N177, N257, N116);
buf BUF1 (N744, N738);
not NOT1 (N745, N737);
nor NOR3 (N746, N696, N115, N131);
or OR2 (N747, N746, N430);
or OR4 (N748, N743, N653, N522, N521);
nor NOR2 (N749, N710, N745);
xor XOR2 (N750, N275, N50);
nor NOR2 (N751, N728, N539);
nor NOR3 (N752, N740, N630, N605);
buf BUF1 (N753, N741);
not NOT1 (N754, N744);
buf BUF1 (N755, N751);
not NOT1 (N756, N753);
nor NOR4 (N757, N755, N74, N252, N78);
not NOT1 (N758, N750);
nor NOR3 (N759, N758, N529, N454);
and AND4 (N760, N735, N679, N16, N486);
or OR4 (N761, N749, N459, N16, N78);
buf BUF1 (N762, N757);
buf BUF1 (N763, N754);
xor XOR2 (N764, N756, N577);
xor XOR2 (N765, N762, N245);
or OR4 (N766, N765, N263, N251, N611);
xor XOR2 (N767, N760, N730);
xor XOR2 (N768, N752, N534);
or OR3 (N769, N764, N130, N685);
buf BUF1 (N770, N759);
and AND4 (N771, N768, N347, N502, N467);
or OR2 (N772, N747, N393);
nor NOR3 (N773, N748, N505, N554);
or OR4 (N774, N767, N436, N637, N374);
buf BUF1 (N775, N772);
nand NAND4 (N776, N742, N434, N405, N337);
or OR3 (N777, N773, N104, N55);
xor XOR2 (N778, N763, N510);
buf BUF1 (N779, N775);
nand NAND2 (N780, N771, N485);
nand NAND4 (N781, N776, N533, N412, N558);
nor NOR2 (N782, N770, N327);
not NOT1 (N783, N777);
or OR4 (N784, N783, N235, N286, N52);
or OR4 (N785, N781, N615, N403, N138);
and AND3 (N786, N778, N148, N236);
or OR4 (N787, N782, N610, N202, N108);
buf BUF1 (N788, N785);
nand NAND3 (N789, N787, N85, N321);
or OR4 (N790, N766, N531, N709, N185);
buf BUF1 (N791, N780);
not NOT1 (N792, N784);
buf BUF1 (N793, N769);
nor NOR2 (N794, N779, N707);
nor NOR2 (N795, N774, N358);
xor XOR2 (N796, N786, N564);
nand NAND4 (N797, N792, N122, N178, N542);
buf BUF1 (N798, N789);
not NOT1 (N799, N793);
nor NOR4 (N800, N791, N522, N377, N135);
nor NOR2 (N801, N790, N464);
nor NOR4 (N802, N798, N779, N450, N573);
buf BUF1 (N803, N802);
xor XOR2 (N804, N761, N399);
or OR2 (N805, N799, N169);
nor NOR4 (N806, N796, N400, N759, N67);
xor XOR2 (N807, N788, N55);
not NOT1 (N808, N806);
xor XOR2 (N809, N797, N337);
xor XOR2 (N810, N809, N726);
buf BUF1 (N811, N808);
xor XOR2 (N812, N804, N24);
or OR4 (N813, N803, N491, N677, N227);
nor NOR3 (N814, N805, N94, N785);
not NOT1 (N815, N801);
nand NAND4 (N816, N813, N259, N808, N230);
not NOT1 (N817, N795);
xor XOR2 (N818, N815, N37);
buf BUF1 (N819, N817);
and AND4 (N820, N818, N226, N610, N321);
and AND4 (N821, N800, N451, N553, N637);
not NOT1 (N822, N820);
nor NOR2 (N823, N811, N296);
and AND3 (N824, N819, N139, N599);
or OR2 (N825, N807, N40);
xor XOR2 (N826, N824, N101);
not NOT1 (N827, N826);
nand NAND3 (N828, N822, N278, N68);
buf BUF1 (N829, N814);
xor XOR2 (N830, N823, N165);
nand NAND4 (N831, N829, N722, N402, N290);
not NOT1 (N832, N810);
buf BUF1 (N833, N794);
and AND4 (N834, N812, N82, N199, N514);
and AND2 (N835, N833, N340);
nand NAND4 (N836, N832, N576, N758, N436);
not NOT1 (N837, N835);
nor NOR2 (N838, N825, N31);
xor XOR2 (N839, N830, N371);
and AND2 (N840, N836, N458);
not NOT1 (N841, N840);
not NOT1 (N842, N827);
buf BUF1 (N843, N821);
xor XOR2 (N844, N842, N342);
buf BUF1 (N845, N831);
not NOT1 (N846, N844);
not NOT1 (N847, N841);
buf BUF1 (N848, N847);
buf BUF1 (N849, N837);
nand NAND2 (N850, N848, N334);
or OR2 (N851, N828, N114);
xor XOR2 (N852, N850, N597);
nor NOR2 (N853, N846, N570);
not NOT1 (N854, N839);
nor NOR3 (N855, N816, N246, N125);
xor XOR2 (N856, N849, N656);
not NOT1 (N857, N843);
xor XOR2 (N858, N853, N675);
nand NAND4 (N859, N858, N354, N670, N224);
buf BUF1 (N860, N854);
nor NOR4 (N861, N859, N153, N102, N817);
and AND4 (N862, N857, N313, N666, N313);
not NOT1 (N863, N852);
not NOT1 (N864, N860);
and AND2 (N865, N862, N485);
xor XOR2 (N866, N838, N435);
buf BUF1 (N867, N865);
or OR4 (N868, N863, N331, N394, N477);
xor XOR2 (N869, N834, N373);
nor NOR3 (N870, N868, N464, N554);
and AND3 (N871, N845, N813, N310);
buf BUF1 (N872, N864);
nand NAND2 (N873, N870, N122);
not NOT1 (N874, N866);
and AND2 (N875, N874, N419);
nand NAND2 (N876, N851, N569);
or OR2 (N877, N876, N757);
not NOT1 (N878, N867);
nand NAND3 (N879, N856, N280, N398);
not NOT1 (N880, N877);
nand NAND4 (N881, N879, N154, N392, N612);
and AND4 (N882, N872, N653, N601, N759);
not NOT1 (N883, N880);
buf BUF1 (N884, N882);
xor XOR2 (N885, N873, N274);
and AND4 (N886, N878, N486, N540, N655);
xor XOR2 (N887, N861, N153);
nand NAND2 (N888, N884, N310);
and AND4 (N889, N881, N497, N398, N844);
xor XOR2 (N890, N883, N233);
buf BUF1 (N891, N875);
nor NOR2 (N892, N871, N158);
buf BUF1 (N893, N889);
buf BUF1 (N894, N869);
buf BUF1 (N895, N888);
xor XOR2 (N896, N885, N290);
nand NAND2 (N897, N887, N739);
buf BUF1 (N898, N895);
and AND4 (N899, N896, N520, N865, N161);
xor XOR2 (N900, N893, N288);
xor XOR2 (N901, N892, N103);
nor NOR4 (N902, N894, N528, N537, N425);
or OR2 (N903, N886, N536);
buf BUF1 (N904, N890);
or OR2 (N905, N903, N387);
or OR2 (N906, N901, N74);
not NOT1 (N907, N899);
not NOT1 (N908, N855);
nor NOR3 (N909, N906, N60, N600);
or OR4 (N910, N904, N835, N605, N352);
not NOT1 (N911, N908);
and AND3 (N912, N897, N781, N878);
nand NAND2 (N913, N909, N532);
xor XOR2 (N914, N910, N412);
xor XOR2 (N915, N914, N388);
xor XOR2 (N916, N891, N411);
and AND2 (N917, N916, N43);
nand NAND4 (N918, N917, N567, N850, N260);
and AND2 (N919, N898, N318);
xor XOR2 (N920, N902, N806);
buf BUF1 (N921, N918);
or OR2 (N922, N920, N563);
xor XOR2 (N923, N921, N641);
nor NOR2 (N924, N915, N169);
nor NOR3 (N925, N907, N317, N304);
not NOT1 (N926, N923);
nor NOR4 (N927, N924, N148, N294, N276);
nand NAND3 (N928, N926, N407, N439);
buf BUF1 (N929, N912);
nor NOR3 (N930, N927, N68, N260);
xor XOR2 (N931, N900, N865);
or OR4 (N932, N930, N541, N12, N94);
and AND4 (N933, N913, N723, N144, N766);
buf BUF1 (N934, N929);
xor XOR2 (N935, N922, N389);
buf BUF1 (N936, N925);
or OR4 (N937, N932, N205, N886, N772);
not NOT1 (N938, N905);
nor NOR2 (N939, N919, N474);
nand NAND3 (N940, N935, N792, N443);
and AND4 (N941, N911, N114, N719, N632);
buf BUF1 (N942, N937);
and AND4 (N943, N939, N461, N542, N237);
and AND3 (N944, N942, N867, N647);
and AND4 (N945, N943, N827, N269, N268);
nand NAND3 (N946, N931, N448, N364);
nor NOR4 (N947, N936, N826, N904, N756);
and AND4 (N948, N934, N295, N788, N609);
xor XOR2 (N949, N928, N651);
nor NOR3 (N950, N945, N851, N631);
nand NAND3 (N951, N944, N93, N656);
and AND2 (N952, N940, N258);
buf BUF1 (N953, N952);
nand NAND2 (N954, N941, N755);
nand NAND2 (N955, N938, N228);
or OR3 (N956, N955, N164, N122);
or OR4 (N957, N946, N903, N244, N452);
xor XOR2 (N958, N951, N343);
or OR3 (N959, N933, N537, N832);
nor NOR3 (N960, N959, N728, N703);
buf BUF1 (N961, N949);
buf BUF1 (N962, N956);
not NOT1 (N963, N961);
and AND4 (N964, N963, N830, N590, N676);
nand NAND2 (N965, N962, N247);
and AND2 (N966, N954, N802);
buf BUF1 (N967, N947);
or OR4 (N968, N953, N374, N45, N263);
and AND4 (N969, N965, N273, N616, N444);
and AND4 (N970, N968, N80, N483, N459);
not NOT1 (N971, N960);
nor NOR4 (N972, N958, N753, N355, N107);
and AND3 (N973, N970, N687, N481);
nand NAND4 (N974, N964, N358, N43, N625);
or OR4 (N975, N974, N126, N283, N840);
and AND3 (N976, N950, N830, N463);
not NOT1 (N977, N966);
buf BUF1 (N978, N973);
or OR4 (N979, N948, N22, N943, N53);
nand NAND2 (N980, N957, N399);
nor NOR2 (N981, N972, N272);
nand NAND2 (N982, N977, N797);
and AND4 (N983, N975, N893, N713, N127);
nor NOR4 (N984, N981, N942, N351, N525);
not NOT1 (N985, N982);
nand NAND2 (N986, N967, N420);
buf BUF1 (N987, N984);
not NOT1 (N988, N978);
and AND2 (N989, N980, N718);
not NOT1 (N990, N985);
or OR4 (N991, N990, N567, N154, N145);
xor XOR2 (N992, N986, N807);
nand NAND2 (N993, N992, N618);
xor XOR2 (N994, N991, N143);
xor XOR2 (N995, N983, N279);
nand NAND4 (N996, N971, N84, N837, N36);
nand NAND4 (N997, N993, N776, N305, N517);
nor NOR2 (N998, N969, N318);
nor NOR4 (N999, N976, N6, N208, N440);
xor XOR2 (N1000, N989, N167);
and AND4 (N1001, N996, N622, N606, N11);
or OR3 (N1002, N988, N284, N639);
or OR3 (N1003, N987, N109, N529);
xor XOR2 (N1004, N994, N16);
xor XOR2 (N1005, N997, N721);
and AND4 (N1006, N1001, N485, N771, N794);
nand NAND3 (N1007, N995, N318, N562);
nand NAND2 (N1008, N1003, N42);
xor XOR2 (N1009, N999, N458);
and AND4 (N1010, N1007, N620, N99, N848);
or OR4 (N1011, N1004, N774, N160, N374);
or OR3 (N1012, N1000, N916, N464);
not NOT1 (N1013, N1009);
xor XOR2 (N1014, N998, N325);
not NOT1 (N1015, N1002);
and AND3 (N1016, N1006, N554, N278);
buf BUF1 (N1017, N1013);
not NOT1 (N1018, N1014);
and AND4 (N1019, N1005, N905, N372, N91);
buf BUF1 (N1020, N1019);
nand NAND2 (N1021, N1008, N574);
and AND3 (N1022, N1017, N193, N566);
and AND2 (N1023, N979, N864);
xor XOR2 (N1024, N1021, N469);
nand NAND2 (N1025, N1010, N146);
nor NOR2 (N1026, N1025, N198);
nand NAND3 (N1027, N1020, N552, N512);
xor XOR2 (N1028, N1024, N390);
xor XOR2 (N1029, N1027, N1015);
nand NAND3 (N1030, N467, N528, N452);
buf BUF1 (N1031, N1016);
or OR4 (N1032, N1028, N730, N907, N1030);
and AND2 (N1033, N650, N905);
nand NAND2 (N1034, N1011, N131);
buf BUF1 (N1035, N1012);
buf BUF1 (N1036, N1026);
or OR2 (N1037, N1018, N832);
buf BUF1 (N1038, N1032);
buf BUF1 (N1039, N1038);
buf BUF1 (N1040, N1031);
buf BUF1 (N1041, N1040);
nand NAND2 (N1042, N1035, N68);
not NOT1 (N1043, N1023);
buf BUF1 (N1044, N1034);
or OR3 (N1045, N1029, N165, N540);
nand NAND2 (N1046, N1045, N855);
xor XOR2 (N1047, N1022, N1002);
not NOT1 (N1048, N1033);
nand NAND2 (N1049, N1044, N225);
and AND4 (N1050, N1039, N214, N853, N332);
nand NAND2 (N1051, N1036, N763);
and AND3 (N1052, N1037, N885, N988);
nor NOR4 (N1053, N1052, N783, N254, N227);
buf BUF1 (N1054, N1049);
or OR2 (N1055, N1050, N732);
nand NAND3 (N1056, N1047, N210, N930);
nor NOR4 (N1057, N1042, N630, N664, N569);
nand NAND3 (N1058, N1041, N412, N1051);
and AND3 (N1059, N657, N60, N318);
or OR3 (N1060, N1059, N843, N249);
buf BUF1 (N1061, N1056);
not NOT1 (N1062, N1055);
or OR4 (N1063, N1048, N887, N721, N523);
buf BUF1 (N1064, N1046);
or OR2 (N1065, N1043, N67);
buf BUF1 (N1066, N1058);
nand NAND2 (N1067, N1062, N872);
buf BUF1 (N1068, N1063);
buf BUF1 (N1069, N1067);
nand NAND4 (N1070, N1060, N43, N512, N599);
not NOT1 (N1071, N1061);
nand NAND2 (N1072, N1053, N29);
or OR2 (N1073, N1070, N530);
buf BUF1 (N1074, N1064);
not NOT1 (N1075, N1072);
or OR4 (N1076, N1071, N520, N143, N1074);
and AND2 (N1077, N230, N290);
and AND3 (N1078, N1075, N834, N539);
nor NOR3 (N1079, N1065, N745, N658);
or OR4 (N1080, N1054, N579, N731, N404);
and AND3 (N1081, N1077, N794, N521);
or OR3 (N1082, N1069, N304, N703);
xor XOR2 (N1083, N1079, N101);
xor XOR2 (N1084, N1083, N1053);
not NOT1 (N1085, N1082);
xor XOR2 (N1086, N1068, N689);
and AND3 (N1087, N1057, N304, N762);
and AND4 (N1088, N1076, N422, N448, N624);
not NOT1 (N1089, N1078);
or OR3 (N1090, N1081, N930, N227);
nand NAND4 (N1091, N1073, N361, N395, N1021);
or OR3 (N1092, N1066, N471, N825);
not NOT1 (N1093, N1090);
nand NAND3 (N1094, N1085, N562, N396);
xor XOR2 (N1095, N1092, N807);
nor NOR3 (N1096, N1094, N793, N756);
not NOT1 (N1097, N1096);
and AND2 (N1098, N1093, N70);
and AND2 (N1099, N1095, N798);
not NOT1 (N1100, N1087);
and AND4 (N1101, N1100, N140, N405, N926);
buf BUF1 (N1102, N1097);
nor NOR4 (N1103, N1080, N574, N391, N1024);
nand NAND4 (N1104, N1102, N309, N380, N580);
or OR2 (N1105, N1098, N793);
nand NAND4 (N1106, N1088, N1080, N564, N611);
not NOT1 (N1107, N1091);
nor NOR2 (N1108, N1101, N147);
nand NAND3 (N1109, N1104, N894, N859);
not NOT1 (N1110, N1105);
and AND3 (N1111, N1110, N50, N656);
or OR3 (N1112, N1106, N1056, N285);
xor XOR2 (N1113, N1084, N287);
buf BUF1 (N1114, N1108);
or OR4 (N1115, N1107, N161, N105, N994);
nor NOR4 (N1116, N1113, N1047, N333, N103);
nand NAND2 (N1117, N1086, N460);
xor XOR2 (N1118, N1117, N775);
and AND2 (N1119, N1111, N1099);
nand NAND2 (N1120, N1112, N405);
not NOT1 (N1121, N55);
buf BUF1 (N1122, N1119);
buf BUF1 (N1123, N1109);
xor XOR2 (N1124, N1121, N629);
buf BUF1 (N1125, N1120);
buf BUF1 (N1126, N1116);
nor NOR3 (N1127, N1123, N1103, N711);
and AND2 (N1128, N597, N163);
or OR2 (N1129, N1126, N1093);
xor XOR2 (N1130, N1129, N523);
nor NOR4 (N1131, N1130, N832, N733, N599);
nor NOR4 (N1132, N1115, N953, N608, N775);
nand NAND4 (N1133, N1124, N841, N10, N977);
or OR2 (N1134, N1127, N473);
xor XOR2 (N1135, N1114, N827);
buf BUF1 (N1136, N1122);
and AND2 (N1137, N1128, N464);
and AND2 (N1138, N1136, N188);
or OR3 (N1139, N1131, N1079, N818);
or OR4 (N1140, N1135, N119, N456, N390);
buf BUF1 (N1141, N1125);
xor XOR2 (N1142, N1133, N510);
nor NOR4 (N1143, N1089, N965, N232, N872);
nand NAND2 (N1144, N1118, N302);
xor XOR2 (N1145, N1144, N10);
not NOT1 (N1146, N1138);
or OR4 (N1147, N1132, N807, N455, N227);
nand NAND4 (N1148, N1142, N1010, N733, N810);
nor NOR2 (N1149, N1134, N888);
nand NAND3 (N1150, N1147, N618, N559);
xor XOR2 (N1151, N1140, N213);
and AND4 (N1152, N1141, N245, N1074, N735);
and AND3 (N1153, N1151, N927, N1100);
and AND4 (N1154, N1153, N954, N638, N25);
nand NAND3 (N1155, N1152, N92, N94);
and AND3 (N1156, N1154, N785, N478);
buf BUF1 (N1157, N1150);
and AND3 (N1158, N1149, N777, N552);
buf BUF1 (N1159, N1148);
xor XOR2 (N1160, N1146, N584);
nand NAND3 (N1161, N1145, N543, N367);
not NOT1 (N1162, N1137);
nor NOR3 (N1163, N1160, N134, N1067);
not NOT1 (N1164, N1163);
or OR3 (N1165, N1158, N1030, N721);
or OR2 (N1166, N1165, N194);
buf BUF1 (N1167, N1155);
buf BUF1 (N1168, N1159);
xor XOR2 (N1169, N1143, N74);
xor XOR2 (N1170, N1139, N469);
and AND2 (N1171, N1162, N502);
and AND4 (N1172, N1170, N1030, N676, N117);
and AND4 (N1173, N1157, N209, N328, N608);
and AND4 (N1174, N1164, N797, N300, N607);
not NOT1 (N1175, N1167);
and AND2 (N1176, N1168, N272);
buf BUF1 (N1177, N1176);
nand NAND3 (N1178, N1166, N1049, N207);
nand NAND2 (N1179, N1172, N92);
nor NOR4 (N1180, N1156, N746, N875, N649);
and AND4 (N1181, N1175, N48, N100, N173);
and AND3 (N1182, N1180, N1056, N641);
not NOT1 (N1183, N1171);
buf BUF1 (N1184, N1181);
nor NOR3 (N1185, N1178, N77, N776);
nand NAND3 (N1186, N1173, N1163, N926);
not NOT1 (N1187, N1182);
not NOT1 (N1188, N1177);
or OR4 (N1189, N1184, N67, N985, N363);
xor XOR2 (N1190, N1187, N910);
or OR2 (N1191, N1169, N762);
and AND2 (N1192, N1188, N969);
not NOT1 (N1193, N1192);
nor NOR2 (N1194, N1193, N145);
not NOT1 (N1195, N1194);
nor NOR3 (N1196, N1183, N454, N295);
nand NAND4 (N1197, N1195, N598, N1013, N618);
not NOT1 (N1198, N1191);
not NOT1 (N1199, N1174);
xor XOR2 (N1200, N1190, N1194);
nand NAND2 (N1201, N1196, N442);
not NOT1 (N1202, N1198);
not NOT1 (N1203, N1189);
nand NAND3 (N1204, N1197, N366, N585);
nor NOR4 (N1205, N1203, N1103, N726, N139);
and AND3 (N1206, N1161, N516, N1140);
xor XOR2 (N1207, N1206, N1026);
xor XOR2 (N1208, N1200, N1051);
buf BUF1 (N1209, N1205);
nand NAND2 (N1210, N1179, N253);
nor NOR3 (N1211, N1202, N996, N695);
or OR4 (N1212, N1204, N1041, N84, N916);
nand NAND2 (N1213, N1185, N86);
xor XOR2 (N1214, N1209, N238);
not NOT1 (N1215, N1211);
or OR4 (N1216, N1212, N175, N1057, N51);
nand NAND2 (N1217, N1216, N861);
and AND3 (N1218, N1217, N585, N414);
buf BUF1 (N1219, N1210);
and AND3 (N1220, N1186, N610, N731);
nand NAND2 (N1221, N1213, N1028);
or OR3 (N1222, N1208, N547, N411);
nor NOR4 (N1223, N1219, N792, N1197, N810);
or OR2 (N1224, N1207, N229);
xor XOR2 (N1225, N1201, N235);
and AND4 (N1226, N1221, N919, N575, N1180);
buf BUF1 (N1227, N1225);
xor XOR2 (N1228, N1222, N443);
nand NAND2 (N1229, N1227, N374);
and AND2 (N1230, N1228, N722);
and AND2 (N1231, N1229, N1093);
not NOT1 (N1232, N1230);
nand NAND4 (N1233, N1220, N394, N765, N1119);
or OR2 (N1234, N1223, N972);
and AND3 (N1235, N1224, N1164, N1079);
nor NOR4 (N1236, N1232, N192, N1108, N589);
nor NOR2 (N1237, N1226, N946);
nand NAND3 (N1238, N1199, N1169, N1082);
nand NAND2 (N1239, N1236, N864);
or OR3 (N1240, N1233, N428, N101);
and AND2 (N1241, N1215, N645);
nor NOR2 (N1242, N1214, N46);
nand NAND2 (N1243, N1240, N802);
not NOT1 (N1244, N1241);
xor XOR2 (N1245, N1231, N204);
nor NOR4 (N1246, N1244, N1127, N602, N134);
buf BUF1 (N1247, N1242);
xor XOR2 (N1248, N1245, N259);
buf BUF1 (N1249, N1237);
xor XOR2 (N1250, N1243, N648);
buf BUF1 (N1251, N1239);
nand NAND4 (N1252, N1218, N642, N13, N886);
or OR4 (N1253, N1234, N507, N492, N296);
nand NAND3 (N1254, N1252, N523, N901);
xor XOR2 (N1255, N1247, N124);
buf BUF1 (N1256, N1255);
and AND4 (N1257, N1235, N337, N92, N367);
nor NOR3 (N1258, N1248, N1172, N1063);
nand NAND3 (N1259, N1256, N486, N739);
xor XOR2 (N1260, N1246, N1257);
nor NOR2 (N1261, N1124, N295);
not NOT1 (N1262, N1261);
nand NAND4 (N1263, N1258, N1217, N786, N901);
not NOT1 (N1264, N1249);
buf BUF1 (N1265, N1254);
buf BUF1 (N1266, N1265);
nor NOR2 (N1267, N1250, N1236);
or OR2 (N1268, N1238, N338);
buf BUF1 (N1269, N1266);
and AND4 (N1270, N1269, N1205, N995, N1130);
or OR2 (N1271, N1253, N525);
not NOT1 (N1272, N1264);
or OR2 (N1273, N1268, N373);
nor NOR3 (N1274, N1251, N471, N857);
not NOT1 (N1275, N1263);
nand NAND4 (N1276, N1271, N525, N24, N265);
buf BUF1 (N1277, N1260);
buf BUF1 (N1278, N1267);
nand NAND3 (N1279, N1262, N164, N483);
not NOT1 (N1280, N1274);
nand NAND4 (N1281, N1273, N604, N439, N811);
and AND2 (N1282, N1275, N1165);
and AND3 (N1283, N1272, N294, N1124);
nor NOR2 (N1284, N1280, N311);
nor NOR3 (N1285, N1278, N1217, N551);
buf BUF1 (N1286, N1276);
buf BUF1 (N1287, N1284);
or OR3 (N1288, N1279, N461, N111);
or OR4 (N1289, N1282, N1113, N373, N932);
not NOT1 (N1290, N1259);
xor XOR2 (N1291, N1290, N587);
xor XOR2 (N1292, N1286, N1118);
and AND3 (N1293, N1287, N1108, N1094);
nand NAND4 (N1294, N1277, N1142, N344, N185);
not NOT1 (N1295, N1291);
xor XOR2 (N1296, N1288, N645);
xor XOR2 (N1297, N1283, N1192);
not NOT1 (N1298, N1295);
xor XOR2 (N1299, N1293, N542);
or OR4 (N1300, N1292, N345, N1197, N1059);
not NOT1 (N1301, N1294);
nor NOR2 (N1302, N1296, N559);
nor NOR2 (N1303, N1270, N1064);
xor XOR2 (N1304, N1297, N1186);
or OR2 (N1305, N1298, N498);
not NOT1 (N1306, N1300);
nand NAND2 (N1307, N1304, N1280);
xor XOR2 (N1308, N1281, N446);
nand NAND4 (N1309, N1301, N435, N172, N91);
and AND4 (N1310, N1306, N1069, N189, N358);
buf BUF1 (N1311, N1299);
or OR4 (N1312, N1310, N194, N546, N1302);
nand NAND4 (N1313, N1170, N982, N1064, N1034);
nor NOR4 (N1314, N1311, N146, N1023, N1295);
nand NAND2 (N1315, N1314, N913);
nor NOR3 (N1316, N1305, N410, N621);
buf BUF1 (N1317, N1303);
nand NAND2 (N1318, N1285, N377);
not NOT1 (N1319, N1309);
nand NAND2 (N1320, N1289, N969);
not NOT1 (N1321, N1315);
buf BUF1 (N1322, N1317);
xor XOR2 (N1323, N1321, N59);
or OR2 (N1324, N1307, N545);
buf BUF1 (N1325, N1319);
buf BUF1 (N1326, N1320);
xor XOR2 (N1327, N1312, N373);
not NOT1 (N1328, N1327);
and AND3 (N1329, N1328, N710, N677);
xor XOR2 (N1330, N1323, N815);
not NOT1 (N1331, N1318);
nand NAND2 (N1332, N1329, N788);
nand NAND3 (N1333, N1316, N330, N719);
not NOT1 (N1334, N1332);
nor NOR4 (N1335, N1330, N738, N703, N517);
not NOT1 (N1336, N1331);
and AND3 (N1337, N1333, N1180, N1139);
and AND3 (N1338, N1325, N468, N1201);
or OR4 (N1339, N1322, N394, N1010, N1200);
nand NAND4 (N1340, N1335, N737, N1310, N1216);
nor NOR2 (N1341, N1326, N643);
or OR4 (N1342, N1324, N113, N166, N154);
and AND4 (N1343, N1334, N1131, N1335, N637);
not NOT1 (N1344, N1313);
or OR4 (N1345, N1344, N268, N313, N1174);
xor XOR2 (N1346, N1339, N583);
nor NOR2 (N1347, N1337, N831);
not NOT1 (N1348, N1346);
xor XOR2 (N1349, N1347, N1165);
buf BUF1 (N1350, N1345);
nand NAND3 (N1351, N1343, N162, N478);
nand NAND4 (N1352, N1336, N523, N784, N775);
or OR4 (N1353, N1352, N563, N1291, N430);
nand NAND4 (N1354, N1338, N486, N632, N1331);
not NOT1 (N1355, N1351);
or OR3 (N1356, N1340, N558, N387);
nand NAND4 (N1357, N1355, N943, N894, N1079);
not NOT1 (N1358, N1308);
nand NAND3 (N1359, N1356, N905, N206);
nor NOR4 (N1360, N1348, N243, N219, N1001);
xor XOR2 (N1361, N1354, N699);
or OR4 (N1362, N1360, N1057, N764, N248);
nand NAND2 (N1363, N1341, N1337);
buf BUF1 (N1364, N1359);
or OR4 (N1365, N1357, N196, N1056, N767);
nand NAND4 (N1366, N1363, N233, N956, N742);
or OR3 (N1367, N1349, N250, N1269);
buf BUF1 (N1368, N1365);
or OR3 (N1369, N1342, N967, N1053);
buf BUF1 (N1370, N1362);
or OR3 (N1371, N1361, N509, N616);
and AND3 (N1372, N1369, N980, N1041);
nand NAND3 (N1373, N1372, N938, N259);
xor XOR2 (N1374, N1368, N346);
nor NOR4 (N1375, N1358, N1237, N342, N1150);
buf BUF1 (N1376, N1367);
not NOT1 (N1377, N1350);
and AND3 (N1378, N1376, N443, N380);
not NOT1 (N1379, N1366);
and AND3 (N1380, N1371, N453, N1019);
xor XOR2 (N1381, N1378, N433);
or OR4 (N1382, N1370, N1111, N893, N1214);
nand NAND3 (N1383, N1381, N162, N334);
not NOT1 (N1384, N1379);
buf BUF1 (N1385, N1377);
nand NAND2 (N1386, N1375, N950);
nor NOR3 (N1387, N1380, N47, N644);
not NOT1 (N1388, N1384);
nand NAND4 (N1389, N1374, N210, N25, N104);
or OR4 (N1390, N1383, N736, N340, N798);
or OR3 (N1391, N1388, N1156, N495);
nor NOR2 (N1392, N1373, N1148);
buf BUF1 (N1393, N1382);
xor XOR2 (N1394, N1392, N724);
nand NAND4 (N1395, N1385, N760, N277, N456);
and AND4 (N1396, N1389, N1261, N1044, N632);
buf BUF1 (N1397, N1393);
nand NAND2 (N1398, N1397, N148);
or OR3 (N1399, N1396, N800, N1147);
and AND4 (N1400, N1398, N576, N609, N1354);
not NOT1 (N1401, N1387);
xor XOR2 (N1402, N1391, N389);
nor NOR3 (N1403, N1399, N757, N1367);
or OR2 (N1404, N1401, N239);
nand NAND4 (N1405, N1402, N1341, N1384, N527);
not NOT1 (N1406, N1404);
buf BUF1 (N1407, N1353);
buf BUF1 (N1408, N1394);
nand NAND3 (N1409, N1405, N748, N1311);
or OR2 (N1410, N1408, N68);
xor XOR2 (N1411, N1364, N1326);
buf BUF1 (N1412, N1386);
nor NOR3 (N1413, N1411, N957, N1103);
not NOT1 (N1414, N1395);
or OR2 (N1415, N1412, N943);
nor NOR4 (N1416, N1409, N848, N927, N1162);
buf BUF1 (N1417, N1416);
and AND2 (N1418, N1407, N1049);
or OR4 (N1419, N1417, N727, N249, N126);
not NOT1 (N1420, N1413);
not NOT1 (N1421, N1390);
xor XOR2 (N1422, N1421, N467);
buf BUF1 (N1423, N1406);
and AND4 (N1424, N1414, N1213, N1293, N1232);
not NOT1 (N1425, N1424);
not NOT1 (N1426, N1418);
not NOT1 (N1427, N1423);
and AND4 (N1428, N1400, N331, N975, N958);
nand NAND2 (N1429, N1422, N1415);
xor XOR2 (N1430, N724, N284);
xor XOR2 (N1431, N1426, N810);
and AND2 (N1432, N1428, N187);
buf BUF1 (N1433, N1432);
xor XOR2 (N1434, N1403, N585);
xor XOR2 (N1435, N1420, N1056);
xor XOR2 (N1436, N1425, N1210);
nor NOR4 (N1437, N1431, N498, N689, N1379);
and AND3 (N1438, N1437, N1355, N578);
and AND2 (N1439, N1410, N1231);
or OR4 (N1440, N1439, N621, N176, N607);
nand NAND2 (N1441, N1430, N1278);
buf BUF1 (N1442, N1419);
xor XOR2 (N1443, N1438, N253);
nand NAND2 (N1444, N1441, N1287);
not NOT1 (N1445, N1434);
or OR4 (N1446, N1442, N415, N335, N921);
xor XOR2 (N1447, N1440, N130);
or OR4 (N1448, N1443, N229, N1010, N656);
buf BUF1 (N1449, N1436);
xor XOR2 (N1450, N1448, N1026);
and AND2 (N1451, N1446, N902);
xor XOR2 (N1452, N1449, N1042);
or OR2 (N1453, N1450, N1090);
buf BUF1 (N1454, N1447);
and AND2 (N1455, N1452, N547);
not NOT1 (N1456, N1455);
nand NAND4 (N1457, N1453, N613, N1035, N1021);
nor NOR3 (N1458, N1444, N1338, N16);
xor XOR2 (N1459, N1433, N718);
buf BUF1 (N1460, N1451);
or OR3 (N1461, N1427, N816, N645);
and AND3 (N1462, N1459, N1015, N466);
or OR4 (N1463, N1445, N392, N611, N589);
buf BUF1 (N1464, N1454);
buf BUF1 (N1465, N1463);
and AND4 (N1466, N1457, N1218, N1174, N267);
not NOT1 (N1467, N1464);
xor XOR2 (N1468, N1461, N213);
nor NOR3 (N1469, N1465, N203, N418);
and AND4 (N1470, N1435, N1043, N1385, N345);
buf BUF1 (N1471, N1462);
buf BUF1 (N1472, N1456);
xor XOR2 (N1473, N1471, N867);
or OR4 (N1474, N1473, N96, N882, N1097);
nand NAND4 (N1475, N1458, N953, N383, N1465);
nand NAND4 (N1476, N1475, N1070, N329, N504);
or OR3 (N1477, N1429, N727, N609);
nand NAND2 (N1478, N1474, N1436);
buf BUF1 (N1479, N1469);
not NOT1 (N1480, N1476);
nor NOR4 (N1481, N1479, N1380, N450, N604);
buf BUF1 (N1482, N1478);
nand NAND2 (N1483, N1468, N1061);
xor XOR2 (N1484, N1460, N429);
buf BUF1 (N1485, N1472);
buf BUF1 (N1486, N1480);
xor XOR2 (N1487, N1470, N775);
nand NAND2 (N1488, N1467, N775);
buf BUF1 (N1489, N1482);
xor XOR2 (N1490, N1477, N25);
xor XOR2 (N1491, N1484, N347);
not NOT1 (N1492, N1490);
not NOT1 (N1493, N1486);
nor NOR4 (N1494, N1466, N857, N354, N733);
nand NAND2 (N1495, N1491, N881);
nor NOR4 (N1496, N1487, N89, N1465, N1393);
and AND3 (N1497, N1489, N687, N972);
or OR3 (N1498, N1497, N834, N1153);
buf BUF1 (N1499, N1495);
not NOT1 (N1500, N1496);
nand NAND2 (N1501, N1498, N997);
xor XOR2 (N1502, N1494, N710);
or OR3 (N1503, N1488, N722, N1028);
nand NAND2 (N1504, N1492, N658);
not NOT1 (N1505, N1485);
and AND3 (N1506, N1483, N366, N994);
xor XOR2 (N1507, N1501, N867);
xor XOR2 (N1508, N1502, N1063);
or OR2 (N1509, N1481, N99);
nand NAND3 (N1510, N1505, N948, N370);
or OR3 (N1511, N1503, N1498, N1370);
or OR4 (N1512, N1510, N809, N607, N504);
or OR4 (N1513, N1499, N768, N1159, N804);
xor XOR2 (N1514, N1493, N151);
not NOT1 (N1515, N1512);
and AND3 (N1516, N1511, N1275, N319);
buf BUF1 (N1517, N1513);
nor NOR4 (N1518, N1516, N608, N1490, N439);
not NOT1 (N1519, N1508);
buf BUF1 (N1520, N1519);
nand NAND2 (N1521, N1509, N992);
or OR2 (N1522, N1500, N577);
nor NOR2 (N1523, N1517, N1039);
and AND4 (N1524, N1515, N908, N562, N814);
buf BUF1 (N1525, N1518);
nand NAND3 (N1526, N1521, N1430, N838);
nand NAND2 (N1527, N1504, N233);
or OR2 (N1528, N1522, N1420);
and AND2 (N1529, N1527, N849);
nor NOR3 (N1530, N1526, N1348, N52);
nand NAND3 (N1531, N1506, N1423, N1419);
xor XOR2 (N1532, N1524, N1033);
nor NOR3 (N1533, N1531, N939, N376);
nor NOR2 (N1534, N1523, N1201);
nor NOR4 (N1535, N1528, N1082, N601, N930);
nor NOR2 (N1536, N1533, N1240);
nand NAND3 (N1537, N1520, N576, N174);
and AND4 (N1538, N1525, N982, N456, N402);
or OR3 (N1539, N1532, N506, N1031);
or OR3 (N1540, N1536, N959, N178);
not NOT1 (N1541, N1530);
xor XOR2 (N1542, N1535, N3);
and AND3 (N1543, N1539, N941, N1288);
and AND2 (N1544, N1507, N85);
buf BUF1 (N1545, N1538);
nor NOR2 (N1546, N1544, N460);
and AND3 (N1547, N1541, N1293, N761);
nor NOR3 (N1548, N1546, N261, N484);
and AND4 (N1549, N1537, N982, N1193, N283);
nor NOR4 (N1550, N1543, N10, N1047, N324);
nand NAND3 (N1551, N1550, N1079, N385);
or OR3 (N1552, N1548, N1299, N650);
xor XOR2 (N1553, N1552, N648);
not NOT1 (N1554, N1540);
buf BUF1 (N1555, N1551);
not NOT1 (N1556, N1549);
buf BUF1 (N1557, N1555);
nand NAND4 (N1558, N1542, N1055, N1001, N153);
buf BUF1 (N1559, N1529);
and AND3 (N1560, N1554, N833, N461);
and AND3 (N1561, N1553, N1208, N544);
not NOT1 (N1562, N1557);
nand NAND4 (N1563, N1558, N75, N338, N355);
nor NOR2 (N1564, N1561, N740);
buf BUF1 (N1565, N1545);
not NOT1 (N1566, N1559);
buf BUF1 (N1567, N1534);
nor NOR3 (N1568, N1556, N1204, N283);
not NOT1 (N1569, N1563);
xor XOR2 (N1570, N1565, N122);
or OR3 (N1571, N1562, N1433, N258);
and AND2 (N1572, N1570, N425);
or OR3 (N1573, N1514, N959, N1534);
buf BUF1 (N1574, N1573);
not NOT1 (N1575, N1560);
xor XOR2 (N1576, N1564, N986);
and AND3 (N1577, N1572, N1297, N887);
or OR4 (N1578, N1577, N1282, N741, N118);
xor XOR2 (N1579, N1547, N22);
and AND2 (N1580, N1568, N1038);
nand NAND3 (N1581, N1576, N1389, N1475);
xor XOR2 (N1582, N1578, N1332);
not NOT1 (N1583, N1575);
and AND3 (N1584, N1574, N677, N4);
nand NAND2 (N1585, N1579, N485);
xor XOR2 (N1586, N1581, N1502);
not NOT1 (N1587, N1585);
xor XOR2 (N1588, N1567, N1165);
or OR3 (N1589, N1583, N231, N228);
nand NAND4 (N1590, N1588, N1039, N615, N1085);
or OR2 (N1591, N1584, N1567);
xor XOR2 (N1592, N1590, N1309);
nor NOR2 (N1593, N1569, N648);
or OR4 (N1594, N1580, N631, N66, N890);
buf BUF1 (N1595, N1566);
xor XOR2 (N1596, N1589, N800);
buf BUF1 (N1597, N1591);
buf BUF1 (N1598, N1592);
xor XOR2 (N1599, N1571, N1560);
buf BUF1 (N1600, N1599);
not NOT1 (N1601, N1597);
nand NAND3 (N1602, N1598, N491, N1565);
nand NAND2 (N1603, N1582, N1602);
nor NOR3 (N1604, N1160, N146, N185);
nor NOR3 (N1605, N1603, N512, N1190);
nor NOR2 (N1606, N1605, N916);
xor XOR2 (N1607, N1595, N1299);
nor NOR2 (N1608, N1586, N858);
nand NAND2 (N1609, N1596, N1446);
buf BUF1 (N1610, N1606);
not NOT1 (N1611, N1600);
not NOT1 (N1612, N1604);
or OR4 (N1613, N1612, N804, N1208, N850);
buf BUF1 (N1614, N1608);
xor XOR2 (N1615, N1593, N1328);
or OR2 (N1616, N1615, N308);
or OR2 (N1617, N1607, N423);
xor XOR2 (N1618, N1613, N34);
nor NOR4 (N1619, N1616, N246, N553, N987);
and AND4 (N1620, N1619, N578, N62, N994);
buf BUF1 (N1621, N1587);
or OR4 (N1622, N1601, N585, N366, N77);
not NOT1 (N1623, N1622);
and AND3 (N1624, N1617, N532, N561);
or OR3 (N1625, N1618, N234, N710);
nand NAND2 (N1626, N1621, N1533);
or OR2 (N1627, N1625, N1277);
or OR3 (N1628, N1623, N1119, N24);
and AND2 (N1629, N1624, N154);
nor NOR2 (N1630, N1594, N1173);
and AND3 (N1631, N1609, N66, N957);
not NOT1 (N1632, N1611);
xor XOR2 (N1633, N1632, N1383);
buf BUF1 (N1634, N1631);
xor XOR2 (N1635, N1620, N1292);
and AND2 (N1636, N1633, N716);
xor XOR2 (N1637, N1634, N233);
or OR2 (N1638, N1627, N926);
xor XOR2 (N1639, N1636, N782);
xor XOR2 (N1640, N1628, N550);
xor XOR2 (N1641, N1626, N869);
buf BUF1 (N1642, N1637);
not NOT1 (N1643, N1635);
xor XOR2 (N1644, N1641, N585);
not NOT1 (N1645, N1610);
not NOT1 (N1646, N1630);
or OR4 (N1647, N1642, N817, N467, N817);
xor XOR2 (N1648, N1644, N1152);
or OR3 (N1649, N1614, N169, N22);
xor XOR2 (N1650, N1639, N307);
nand NAND2 (N1651, N1649, N1329);
xor XOR2 (N1652, N1645, N1336);
nand NAND3 (N1653, N1651, N820, N1125);
nor NOR4 (N1654, N1640, N351, N11, N1136);
nand NAND2 (N1655, N1652, N659);
or OR4 (N1656, N1629, N1, N1114, N644);
or OR4 (N1657, N1653, N1543, N1202, N389);
nand NAND2 (N1658, N1654, N722);
nand NAND4 (N1659, N1643, N1298, N1559, N594);
and AND4 (N1660, N1655, N174, N452, N509);
or OR4 (N1661, N1656, N1469, N1365, N1574);
not NOT1 (N1662, N1648);
buf BUF1 (N1663, N1638);
or OR2 (N1664, N1657, N1225);
and AND3 (N1665, N1650, N929, N1406);
and AND4 (N1666, N1659, N1037, N542, N1288);
buf BUF1 (N1667, N1662);
nor NOR4 (N1668, N1660, N945, N690, N1374);
nor NOR4 (N1669, N1647, N273, N462, N1413);
nand NAND3 (N1670, N1661, N1090, N755);
xor XOR2 (N1671, N1646, N940);
buf BUF1 (N1672, N1663);
buf BUF1 (N1673, N1667);
buf BUF1 (N1674, N1658);
buf BUF1 (N1675, N1668);
buf BUF1 (N1676, N1671);
or OR3 (N1677, N1669, N127, N741);
not NOT1 (N1678, N1666);
buf BUF1 (N1679, N1677);
nand NAND2 (N1680, N1678, N1109);
nand NAND3 (N1681, N1676, N953, N1658);
buf BUF1 (N1682, N1680);
not NOT1 (N1683, N1673);
nor NOR3 (N1684, N1674, N380, N730);
xor XOR2 (N1685, N1682, N1498);
xor XOR2 (N1686, N1664, N1435);
and AND4 (N1687, N1685, N1018, N804, N1294);
or OR3 (N1688, N1687, N1665, N406);
and AND3 (N1689, N915, N254, N304);
nor NOR3 (N1690, N1688, N1313, N1503);
or OR4 (N1691, N1684, N1099, N172, N1011);
nor NOR2 (N1692, N1679, N148);
not NOT1 (N1693, N1681);
buf BUF1 (N1694, N1683);
nand NAND4 (N1695, N1690, N841, N772, N1281);
nand NAND4 (N1696, N1686, N275, N412, N427);
buf BUF1 (N1697, N1689);
nor NOR2 (N1698, N1695, N1408);
and AND4 (N1699, N1698, N1158, N147, N1619);
not NOT1 (N1700, N1694);
and AND3 (N1701, N1672, N168, N158);
nor NOR2 (N1702, N1701, N69);
and AND3 (N1703, N1697, N1291, N935);
nor NOR3 (N1704, N1692, N1333, N923);
or OR3 (N1705, N1702, N1650, N1692);
not NOT1 (N1706, N1703);
buf BUF1 (N1707, N1706);
nor NOR4 (N1708, N1704, N973, N702, N1317);
buf BUF1 (N1709, N1699);
and AND4 (N1710, N1691, N1348, N1424, N619);
or OR2 (N1711, N1709, N382);
nor NOR3 (N1712, N1675, N943, N1149);
or OR2 (N1713, N1708, N1236);
nand NAND2 (N1714, N1707, N149);
nor NOR3 (N1715, N1670, N1501, N208);
and AND2 (N1716, N1711, N315);
nor NOR3 (N1717, N1710, N1308, N1062);
nor NOR2 (N1718, N1714, N1077);
and AND3 (N1719, N1700, N231, N681);
and AND4 (N1720, N1713, N662, N971, N1335);
buf BUF1 (N1721, N1718);
not NOT1 (N1722, N1693);
nor NOR3 (N1723, N1721, N412, N681);
buf BUF1 (N1724, N1715);
and AND3 (N1725, N1722, N1275, N1433);
not NOT1 (N1726, N1717);
not NOT1 (N1727, N1720);
and AND3 (N1728, N1723, N192, N703);
not NOT1 (N1729, N1719);
xor XOR2 (N1730, N1729, N329);
and AND3 (N1731, N1696, N1725, N1201);
nor NOR4 (N1732, N1406, N887, N1417, N366);
and AND4 (N1733, N1716, N973, N607, N1204);
nor NOR4 (N1734, N1733, N835, N1422, N1385);
nor NOR4 (N1735, N1712, N340, N361, N688);
and AND3 (N1736, N1732, N1649, N981);
or OR3 (N1737, N1735, N881, N828);
or OR3 (N1738, N1731, N1646, N678);
and AND4 (N1739, N1724, N1485, N73, N1651);
nand NAND2 (N1740, N1705, N254);
nand NAND3 (N1741, N1730, N1550, N359);
nand NAND4 (N1742, N1736, N565, N4, N384);
buf BUF1 (N1743, N1739);
and AND3 (N1744, N1734, N319, N1062);
and AND4 (N1745, N1740, N645, N970, N637);
buf BUF1 (N1746, N1737);
xor XOR2 (N1747, N1741, N985);
and AND3 (N1748, N1738, N446, N1576);
nand NAND2 (N1749, N1728, N780);
nand NAND4 (N1750, N1748, N450, N806, N1071);
and AND4 (N1751, N1749, N1511, N651, N862);
buf BUF1 (N1752, N1743);
not NOT1 (N1753, N1746);
and AND2 (N1754, N1744, N730);
nor NOR2 (N1755, N1754, N595);
buf BUF1 (N1756, N1752);
and AND4 (N1757, N1756, N1329, N425, N235);
xor XOR2 (N1758, N1757, N1058);
buf BUF1 (N1759, N1750);
or OR3 (N1760, N1753, N102, N1552);
buf BUF1 (N1761, N1759);
nand NAND4 (N1762, N1761, N499, N1243, N1137);
not NOT1 (N1763, N1747);
nand NAND2 (N1764, N1755, N1136);
or OR4 (N1765, N1745, N1118, N493, N709);
and AND3 (N1766, N1742, N1073, N1039);
xor XOR2 (N1767, N1765, N1695);
buf BUF1 (N1768, N1726);
or OR4 (N1769, N1767, N1662, N527, N7);
nand NAND4 (N1770, N1764, N1288, N55, N101);
nor NOR3 (N1771, N1770, N1020, N1270);
nor NOR2 (N1772, N1758, N619);
nor NOR3 (N1773, N1727, N861, N56);
and AND4 (N1774, N1763, N1334, N1138, N882);
or OR2 (N1775, N1769, N217);
and AND4 (N1776, N1766, N1206, N902, N1668);
or OR2 (N1777, N1760, N69);
xor XOR2 (N1778, N1768, N211);
not NOT1 (N1779, N1776);
nor NOR2 (N1780, N1762, N1012);
buf BUF1 (N1781, N1780);
and AND3 (N1782, N1751, N763, N809);
nor NOR3 (N1783, N1777, N1069, N811);
not NOT1 (N1784, N1783);
or OR4 (N1785, N1772, N211, N1485, N1346);
not NOT1 (N1786, N1785);
and AND3 (N1787, N1775, N705, N1024);
or OR3 (N1788, N1779, N472, N721);
nand NAND4 (N1789, N1778, N82, N145, N1159);
xor XOR2 (N1790, N1788, N1612);
nor NOR4 (N1791, N1771, N335, N448, N1168);
not NOT1 (N1792, N1791);
xor XOR2 (N1793, N1774, N856);
and AND2 (N1794, N1792, N1668);
nor NOR2 (N1795, N1789, N462);
nand NAND2 (N1796, N1782, N950);
nor NOR4 (N1797, N1784, N875, N948, N1179);
or OR3 (N1798, N1773, N89, N226);
nor NOR4 (N1799, N1794, N1123, N1556, N1302);
nand NAND2 (N1800, N1798, N1104);
buf BUF1 (N1801, N1781);
not NOT1 (N1802, N1793);
and AND2 (N1803, N1796, N740);
nand NAND4 (N1804, N1801, N540, N1668, N1688);
buf BUF1 (N1805, N1790);
not NOT1 (N1806, N1802);
nand NAND3 (N1807, N1795, N259, N722);
nand NAND2 (N1808, N1806, N475);
xor XOR2 (N1809, N1787, N1026);
nand NAND3 (N1810, N1808, N1002, N977);
nand NAND4 (N1811, N1804, N16, N904, N296);
and AND2 (N1812, N1803, N1149);
and AND3 (N1813, N1805, N421, N645);
xor XOR2 (N1814, N1809, N322);
nand NAND4 (N1815, N1786, N1559, N521, N1205);
or OR4 (N1816, N1812, N1636, N320, N1309);
buf BUF1 (N1817, N1815);
or OR3 (N1818, N1817, N1558, N1468);
and AND2 (N1819, N1813, N50);
nand NAND4 (N1820, N1807, N1736, N931, N597);
and AND2 (N1821, N1810, N1055);
or OR4 (N1822, N1814, N1454, N1773, N1674);
or OR4 (N1823, N1797, N1134, N1389, N376);
nand NAND2 (N1824, N1799, N1704);
or OR2 (N1825, N1822, N1140);
buf BUF1 (N1826, N1821);
or OR4 (N1827, N1823, N1411, N784, N85);
and AND3 (N1828, N1800, N1076, N301);
or OR3 (N1829, N1811, N1344, N305);
buf BUF1 (N1830, N1829);
buf BUF1 (N1831, N1824);
and AND2 (N1832, N1831, N47);
or OR4 (N1833, N1825, N661, N150, N1504);
xor XOR2 (N1834, N1828, N1687);
not NOT1 (N1835, N1826);
nor NOR4 (N1836, N1833, N1402, N700, N609);
or OR3 (N1837, N1835, N1730, N1012);
not NOT1 (N1838, N1818);
buf BUF1 (N1839, N1834);
and AND2 (N1840, N1836, N92);
and AND4 (N1841, N1827, N1000, N213, N548);
or OR2 (N1842, N1838, N740);
buf BUF1 (N1843, N1832);
and AND4 (N1844, N1830, N1786, N588, N963);
and AND3 (N1845, N1844, N248, N23);
not NOT1 (N1846, N1842);
or OR4 (N1847, N1820, N421, N1044, N1700);
or OR2 (N1848, N1847, N1526);
nor NOR2 (N1849, N1846, N1037);
nand NAND3 (N1850, N1819, N300, N1040);
not NOT1 (N1851, N1837);
not NOT1 (N1852, N1848);
and AND2 (N1853, N1843, N1406);
not NOT1 (N1854, N1851);
buf BUF1 (N1855, N1849);
buf BUF1 (N1856, N1852);
nand NAND4 (N1857, N1856, N1392, N1800, N673);
buf BUF1 (N1858, N1839);
not NOT1 (N1859, N1816);
buf BUF1 (N1860, N1853);
nand NAND4 (N1861, N1859, N586, N450, N1283);
buf BUF1 (N1862, N1861);
xor XOR2 (N1863, N1862, N622);
not NOT1 (N1864, N1841);
or OR2 (N1865, N1855, N1702);
buf BUF1 (N1866, N1865);
and AND3 (N1867, N1860, N1488, N614);
or OR2 (N1868, N1850, N1811);
buf BUF1 (N1869, N1857);
or OR4 (N1870, N1840, N685, N1233, N1292);
or OR2 (N1871, N1870, N249);
nor NOR3 (N1872, N1864, N1510, N1811);
nand NAND3 (N1873, N1872, N690, N1050);
xor XOR2 (N1874, N1854, N1779);
not NOT1 (N1875, N1873);
buf BUF1 (N1876, N1874);
nor NOR2 (N1877, N1863, N676);
nor NOR3 (N1878, N1867, N1308, N634);
nand NAND4 (N1879, N1858, N187, N1377, N35);
nand NAND4 (N1880, N1877, N399, N711, N771);
or OR4 (N1881, N1868, N466, N829, N760);
nand NAND3 (N1882, N1878, N71, N150);
buf BUF1 (N1883, N1871);
or OR2 (N1884, N1876, N393);
and AND4 (N1885, N1845, N215, N869, N57);
nor NOR4 (N1886, N1883, N1230, N187, N626);
or OR4 (N1887, N1866, N1090, N1858, N798);
nand NAND2 (N1888, N1884, N111);
xor XOR2 (N1889, N1888, N1555);
or OR2 (N1890, N1880, N1036);
nand NAND3 (N1891, N1890, N1005, N1433);
and AND3 (N1892, N1875, N942, N401);
xor XOR2 (N1893, N1879, N1730);
nor NOR2 (N1894, N1887, N1323);
or OR3 (N1895, N1891, N637, N1385);
not NOT1 (N1896, N1881);
or OR4 (N1897, N1895, N1778, N69, N1099);
xor XOR2 (N1898, N1893, N380);
or OR3 (N1899, N1886, N743, N1727);
buf BUF1 (N1900, N1897);
or OR3 (N1901, N1892, N11, N260);
nand NAND3 (N1902, N1885, N348, N825);
nand NAND4 (N1903, N1889, N1840, N1237, N1873);
not NOT1 (N1904, N1903);
and AND4 (N1905, N1904, N363, N1224, N1516);
nor NOR4 (N1906, N1899, N988, N632, N401);
or OR2 (N1907, N1900, N1016);
not NOT1 (N1908, N1869);
buf BUF1 (N1909, N1905);
or OR3 (N1910, N1908, N1393, N777);
nor NOR3 (N1911, N1882, N591, N1664);
xor XOR2 (N1912, N1894, N1091);
buf BUF1 (N1913, N1909);
nand NAND2 (N1914, N1912, N298);
buf BUF1 (N1915, N1907);
and AND2 (N1916, N1902, N1704);
nor NOR4 (N1917, N1910, N1784, N935, N1349);
and AND3 (N1918, N1911, N1856, N252);
not NOT1 (N1919, N1913);
nor NOR3 (N1920, N1917, N1351, N706);
xor XOR2 (N1921, N1915, N1687);
and AND3 (N1922, N1916, N305, N769);
or OR4 (N1923, N1920, N795, N574, N406);
nand NAND3 (N1924, N1906, N263, N1346);
not NOT1 (N1925, N1919);
not NOT1 (N1926, N1925);
not NOT1 (N1927, N1921);
or OR4 (N1928, N1923, N1673, N1132, N466);
not NOT1 (N1929, N1927);
xor XOR2 (N1930, N1896, N1093);
or OR3 (N1931, N1930, N102, N178);
nor NOR3 (N1932, N1928, N1646, N1517);
buf BUF1 (N1933, N1929);
xor XOR2 (N1934, N1924, N1314);
nand NAND3 (N1935, N1901, N771, N1521);
or OR2 (N1936, N1933, N152);
nand NAND3 (N1937, N1935, N1700, N81);
not NOT1 (N1938, N1937);
nor NOR4 (N1939, N1926, N968, N849, N403);
buf BUF1 (N1940, N1914);
or OR2 (N1941, N1936, N1687);
or OR2 (N1942, N1932, N827);
not NOT1 (N1943, N1931);
or OR2 (N1944, N1940, N76);
not NOT1 (N1945, N1938);
buf BUF1 (N1946, N1943);
or OR3 (N1947, N1898, N729, N1193);
not NOT1 (N1948, N1945);
xor XOR2 (N1949, N1946, N591);
nand NAND4 (N1950, N1942, N1514, N794, N476);
nand NAND3 (N1951, N1949, N850, N1274);
and AND4 (N1952, N1934, N963, N1740, N328);
xor XOR2 (N1953, N1939, N1031);
nor NOR2 (N1954, N1944, N715);
not NOT1 (N1955, N1918);
buf BUF1 (N1956, N1948);
nor NOR3 (N1957, N1955, N366, N1096);
buf BUF1 (N1958, N1954);
xor XOR2 (N1959, N1951, N1063);
or OR2 (N1960, N1952, N392);
nand NAND2 (N1961, N1957, N1566);
nand NAND4 (N1962, N1953, N1866, N1668, N1958);
or OR3 (N1963, N1400, N11, N1390);
buf BUF1 (N1964, N1961);
not NOT1 (N1965, N1941);
xor XOR2 (N1966, N1956, N1962);
not NOT1 (N1967, N556);
nor NOR2 (N1968, N1966, N1630);
not NOT1 (N1969, N1963);
buf BUF1 (N1970, N1960);
xor XOR2 (N1971, N1967, N10);
xor XOR2 (N1972, N1969, N764);
xor XOR2 (N1973, N1968, N919);
not NOT1 (N1974, N1950);
nor NOR4 (N1975, N1947, N213, N1414, N239);
xor XOR2 (N1976, N1972, N400);
and AND4 (N1977, N1970, N348, N343, N1904);
nand NAND4 (N1978, N1922, N926, N1164, N112);
xor XOR2 (N1979, N1964, N1878);
nand NAND4 (N1980, N1979, N298, N257, N138);
buf BUF1 (N1981, N1977);
xor XOR2 (N1982, N1971, N133);
nor NOR4 (N1983, N1980, N1728, N1925, N254);
xor XOR2 (N1984, N1976, N1442);
and AND2 (N1985, N1984, N1153);
nand NAND4 (N1986, N1959, N1340, N587, N199);
xor XOR2 (N1987, N1985, N194);
xor XOR2 (N1988, N1973, N228);
not NOT1 (N1989, N1986);
xor XOR2 (N1990, N1988, N1164);
nand NAND4 (N1991, N1975, N1041, N479, N283);
nor NOR2 (N1992, N1989, N333);
and AND4 (N1993, N1965, N624, N1576, N997);
not NOT1 (N1994, N1990);
nand NAND2 (N1995, N1983, N1957);
buf BUF1 (N1996, N1992);
nor NOR2 (N1997, N1981, N177);
not NOT1 (N1998, N1995);
and AND2 (N1999, N1991, N494);
not NOT1 (N2000, N1982);
xor XOR2 (N2001, N1999, N1896);
and AND3 (N2002, N1974, N799, N1732);
not NOT1 (N2003, N1997);
or OR4 (N2004, N1978, N1480, N850, N1300);
nor NOR3 (N2005, N2004, N637, N1135);
or OR2 (N2006, N2002, N402);
and AND4 (N2007, N1987, N186, N881, N1337);
xor XOR2 (N2008, N2006, N1861);
or OR3 (N2009, N2001, N550, N712);
not NOT1 (N2010, N1994);
nand NAND2 (N2011, N1993, N924);
buf BUF1 (N2012, N2005);
xor XOR2 (N2013, N2000, N37);
buf BUF1 (N2014, N2011);
xor XOR2 (N2015, N2013, N195);
or OR4 (N2016, N2008, N43, N57, N12);
xor XOR2 (N2017, N2003, N1931);
buf BUF1 (N2018, N2017);
or OR2 (N2019, N2018, N730);
nand NAND4 (N2020, N1998, N1819, N1514, N669);
or OR3 (N2021, N2009, N292, N686);
and AND4 (N2022, N1996, N117, N115, N1152);
not NOT1 (N2023, N2016);
xor XOR2 (N2024, N2012, N315);
buf BUF1 (N2025, N2019);
xor XOR2 (N2026, N2020, N1299);
xor XOR2 (N2027, N2014, N742);
and AND3 (N2028, N2010, N603, N1094);
buf BUF1 (N2029, N2024);
nand NAND3 (N2030, N2007, N1642, N216);
xor XOR2 (N2031, N2026, N928);
xor XOR2 (N2032, N2031, N1008);
nand NAND2 (N2033, N2015, N874);
nand NAND3 (N2034, N2027, N223, N1650);
buf BUF1 (N2035, N2022);
not NOT1 (N2036, N2034);
buf BUF1 (N2037, N2032);
nor NOR3 (N2038, N2035, N547, N491);
not NOT1 (N2039, N2038);
or OR2 (N2040, N2029, N1445);
or OR4 (N2041, N2037, N623, N1894, N1559);
xor XOR2 (N2042, N2021, N741);
xor XOR2 (N2043, N2036, N578);
nand NAND2 (N2044, N2043, N1700);
not NOT1 (N2045, N2033);
xor XOR2 (N2046, N2030, N173);
nand NAND2 (N2047, N2046, N200);
not NOT1 (N2048, N2039);
and AND2 (N2049, N2045, N1119);
not NOT1 (N2050, N2025);
xor XOR2 (N2051, N2050, N1607);
nor NOR3 (N2052, N2028, N233, N529);
xor XOR2 (N2053, N2049, N880);
or OR3 (N2054, N2044, N1627, N891);
xor XOR2 (N2055, N2053, N1378);
or OR3 (N2056, N2040, N801, N324);
not NOT1 (N2057, N2054);
nor NOR4 (N2058, N2047, N1864, N788, N1483);
xor XOR2 (N2059, N2041, N1411);
or OR2 (N2060, N2056, N1139);
xor XOR2 (N2061, N2057, N1682);
and AND2 (N2062, N2042, N1037);
xor XOR2 (N2063, N2062, N1250);
nor NOR3 (N2064, N2061, N1620, N5);
buf BUF1 (N2065, N2058);
xor XOR2 (N2066, N2052, N1269);
not NOT1 (N2067, N2059);
or OR4 (N2068, N2051, N1754, N2033, N1635);
nor NOR4 (N2069, N2065, N1870, N5, N1959);
nand NAND2 (N2070, N2060, N553);
not NOT1 (N2071, N2063);
buf BUF1 (N2072, N2070);
not NOT1 (N2073, N2072);
xor XOR2 (N2074, N2073, N753);
not NOT1 (N2075, N2067);
nor NOR4 (N2076, N2075, N261, N513, N298);
not NOT1 (N2077, N2023);
nor NOR3 (N2078, N2066, N358, N1936);
nand NAND4 (N2079, N2077, N1400, N768, N613);
and AND2 (N2080, N2071, N2033);
nor NOR4 (N2081, N2048, N1515, N133, N1452);
buf BUF1 (N2082, N2074);
xor XOR2 (N2083, N2069, N1724);
nor NOR3 (N2084, N2064, N284, N732);
nand NAND2 (N2085, N2076, N956);
nor NOR2 (N2086, N2055, N521);
nand NAND3 (N2087, N2068, N910, N897);
xor XOR2 (N2088, N2085, N584);
nor NOR2 (N2089, N2088, N884);
nand NAND4 (N2090, N2089, N1267, N1313, N1574);
or OR2 (N2091, N2080, N614);
not NOT1 (N2092, N2078);
buf BUF1 (N2093, N2086);
and AND2 (N2094, N2084, N568);
and AND3 (N2095, N2090, N294, N1189);
or OR2 (N2096, N2082, N610);
nand NAND3 (N2097, N2091, N1043, N1517);
xor XOR2 (N2098, N2093, N447);
not NOT1 (N2099, N2081);
not NOT1 (N2100, N2095);
not NOT1 (N2101, N2098);
and AND4 (N2102, N2099, N445, N1767, N633);
not NOT1 (N2103, N2087);
not NOT1 (N2104, N2103);
nor NOR4 (N2105, N2102, N631, N1465, N1187);
and AND4 (N2106, N2083, N1680, N1406, N1152);
not NOT1 (N2107, N2094);
and AND3 (N2108, N2079, N427, N1300);
buf BUF1 (N2109, N2108);
nand NAND2 (N2110, N2097, N1248);
buf BUF1 (N2111, N2096);
or OR2 (N2112, N2111, N1770);
not NOT1 (N2113, N2107);
xor XOR2 (N2114, N2110, N1190);
nand NAND3 (N2115, N2105, N152, N1737);
not NOT1 (N2116, N2115);
nand NAND4 (N2117, N2116, N305, N2009, N1890);
and AND3 (N2118, N2106, N1694, N767);
nor NOR2 (N2119, N2092, N263);
xor XOR2 (N2120, N2104, N1789);
xor XOR2 (N2121, N2100, N234);
and AND3 (N2122, N2118, N1263, N205);
and AND2 (N2123, N2121, N474);
xor XOR2 (N2124, N2120, N1486);
nor NOR3 (N2125, N2101, N19, N2064);
or OR3 (N2126, N2117, N1620, N1016);
xor XOR2 (N2127, N2109, N380);
buf BUF1 (N2128, N2125);
or OR3 (N2129, N2112, N1622, N2091);
or OR4 (N2130, N2127, N1654, N1587, N983);
and AND3 (N2131, N2113, N1721, N1376);
nand NAND2 (N2132, N2123, N918);
nor NOR3 (N2133, N2114, N717, N1425);
buf BUF1 (N2134, N2132);
nor NOR2 (N2135, N2131, N1995);
or OR4 (N2136, N2133, N1751, N557, N536);
nand NAND3 (N2137, N2130, N1215, N925);
nor NOR2 (N2138, N2129, N1238);
buf BUF1 (N2139, N2128);
nand NAND3 (N2140, N2134, N972, N1710);
buf BUF1 (N2141, N2124);
not NOT1 (N2142, N2137);
not NOT1 (N2143, N2142);
xor XOR2 (N2144, N2140, N1049);
nor NOR3 (N2145, N2144, N2081, N1295);
not NOT1 (N2146, N2143);
buf BUF1 (N2147, N2145);
xor XOR2 (N2148, N2147, N1932);
not NOT1 (N2149, N2148);
buf BUF1 (N2150, N2126);
nor NOR4 (N2151, N2138, N994, N1659, N968);
not NOT1 (N2152, N2136);
not NOT1 (N2153, N2151);
nand NAND3 (N2154, N2152, N1965, N1174);
not NOT1 (N2155, N2154);
nor NOR4 (N2156, N2141, N1626, N1036, N1066);
nor NOR3 (N2157, N2119, N1183, N857);
and AND2 (N2158, N2153, N1070);
nand NAND4 (N2159, N2157, N1612, N583, N793);
nor NOR3 (N2160, N2156, N1857, N595);
not NOT1 (N2161, N2149);
nor NOR4 (N2162, N2161, N1071, N1128, N2109);
buf BUF1 (N2163, N2150);
buf BUF1 (N2164, N2163);
nor NOR3 (N2165, N2158, N1886, N49);
nor NOR3 (N2166, N2146, N1194, N1856);
buf BUF1 (N2167, N2139);
or OR3 (N2168, N2155, N256, N1901);
xor XOR2 (N2169, N2162, N513);
nor NOR3 (N2170, N2166, N377, N1268);
nand NAND4 (N2171, N2135, N835, N1347, N869);
nor NOR3 (N2172, N2167, N546, N1341);
not NOT1 (N2173, N2170);
xor XOR2 (N2174, N2169, N827);
or OR2 (N2175, N2122, N1557);
nand NAND2 (N2176, N2160, N299);
and AND2 (N2177, N2165, N1267);
nand NAND4 (N2178, N2174, N1641, N591, N101);
and AND2 (N2179, N2176, N636);
not NOT1 (N2180, N2159);
nor NOR2 (N2181, N2173, N2101);
and AND4 (N2182, N2181, N768, N1593, N798);
buf BUF1 (N2183, N2164);
buf BUF1 (N2184, N2182);
or OR2 (N2185, N2178, N1914);
nor NOR2 (N2186, N2172, N1557);
and AND4 (N2187, N2177, N2055, N1388, N90);
buf BUF1 (N2188, N2185);
or OR3 (N2189, N2188, N952, N1902);
and AND3 (N2190, N2184, N1184, N1396);
buf BUF1 (N2191, N2171);
nor NOR3 (N2192, N2190, N452, N919);
not NOT1 (N2193, N2175);
nor NOR4 (N2194, N2186, N1284, N659, N693);
nand NAND2 (N2195, N2191, N1637);
xor XOR2 (N2196, N2183, N1826);
nor NOR3 (N2197, N2180, N423, N2093);
and AND4 (N2198, N2192, N1336, N1707, N807);
buf BUF1 (N2199, N2189);
buf BUF1 (N2200, N2195);
or OR3 (N2201, N2197, N2094, N495);
xor XOR2 (N2202, N2168, N1891);
nor NOR4 (N2203, N2198, N275, N1270, N1747);
xor XOR2 (N2204, N2193, N20);
xor XOR2 (N2205, N2194, N121);
or OR2 (N2206, N2196, N2202);
not NOT1 (N2207, N317);
not NOT1 (N2208, N2205);
nor NOR3 (N2209, N2187, N1813, N152);
not NOT1 (N2210, N2179);
xor XOR2 (N2211, N2210, N1396);
not NOT1 (N2212, N2206);
not NOT1 (N2213, N2209);
buf BUF1 (N2214, N2211);
or OR2 (N2215, N2212, N1072);
or OR2 (N2216, N2207, N421);
nand NAND3 (N2217, N2213, N2154, N310);
buf BUF1 (N2218, N2204);
buf BUF1 (N2219, N2217);
and AND4 (N2220, N2203, N694, N96, N2193);
not NOT1 (N2221, N2216);
nand NAND4 (N2222, N2199, N109, N908, N2144);
not NOT1 (N2223, N2215);
or OR4 (N2224, N2218, N708, N1615, N124);
or OR2 (N2225, N2220, N2035);
xor XOR2 (N2226, N2222, N2042);
xor XOR2 (N2227, N2224, N161);
xor XOR2 (N2228, N2225, N1142);
not NOT1 (N2229, N2223);
or OR2 (N2230, N2200, N1699);
or OR4 (N2231, N2226, N634, N208, N821);
nand NAND2 (N2232, N2228, N730);
xor XOR2 (N2233, N2221, N299);
and AND3 (N2234, N2219, N158, N1035);
buf BUF1 (N2235, N2233);
nand NAND4 (N2236, N2234, N126, N689, N2234);
nand NAND4 (N2237, N2227, N209, N91, N2163);
nor NOR3 (N2238, N2230, N37, N1985);
xor XOR2 (N2239, N2208, N1590);
not NOT1 (N2240, N2236);
or OR2 (N2241, N2238, N2188);
xor XOR2 (N2242, N2232, N1765);
nand NAND4 (N2243, N2201, N27, N1503, N1280);
xor XOR2 (N2244, N2229, N1476);
not NOT1 (N2245, N2235);
or OR4 (N2246, N2240, N2212, N1709, N761);
and AND4 (N2247, N2246, N1549, N59, N1609);
or OR2 (N2248, N2231, N858);
xor XOR2 (N2249, N2242, N1886);
xor XOR2 (N2250, N2247, N1327);
buf BUF1 (N2251, N2249);
and AND4 (N2252, N2248, N45, N2170, N1925);
and AND2 (N2253, N2214, N1949);
nor NOR2 (N2254, N2239, N1766);
and AND4 (N2255, N2252, N411, N1336, N1310);
or OR3 (N2256, N2251, N1286, N1470);
or OR4 (N2257, N2250, N2230, N1644, N1669);
nor NOR3 (N2258, N2255, N1912, N797);
not NOT1 (N2259, N2237);
xor XOR2 (N2260, N2258, N1991);
nor NOR3 (N2261, N2243, N1057, N165);
and AND4 (N2262, N2257, N1659, N940, N990);
not NOT1 (N2263, N2261);
and AND3 (N2264, N2263, N1055, N1670);
nor NOR4 (N2265, N2260, N1572, N1968, N349);
nor NOR4 (N2266, N2259, N198, N140, N8);
or OR3 (N2267, N2244, N1621, N1778);
nand NAND3 (N2268, N2245, N627, N337);
xor XOR2 (N2269, N2253, N1956);
nand NAND3 (N2270, N2266, N489, N580);
buf BUF1 (N2271, N2270);
buf BUF1 (N2272, N2271);
not NOT1 (N2273, N2264);
xor XOR2 (N2274, N2273, N2123);
and AND2 (N2275, N2267, N1895);
buf BUF1 (N2276, N2275);
nand NAND4 (N2277, N2276, N2204, N114, N811);
and AND2 (N2278, N2268, N2231);
not NOT1 (N2279, N2274);
nor NOR4 (N2280, N2254, N2189, N1472, N1888);
xor XOR2 (N2281, N2262, N1806);
buf BUF1 (N2282, N2272);
buf BUF1 (N2283, N2277);
nor NOR4 (N2284, N2265, N1189, N613, N222);
buf BUF1 (N2285, N2280);
nand NAND2 (N2286, N2278, N2189);
or OR3 (N2287, N2282, N312, N1427);
and AND2 (N2288, N2256, N2272);
nor NOR4 (N2289, N2287, N2073, N481, N1426);
and AND2 (N2290, N2285, N257);
xor XOR2 (N2291, N2283, N2198);
or OR3 (N2292, N2291, N328, N718);
nand NAND4 (N2293, N2241, N1293, N703, N753);
xor XOR2 (N2294, N2286, N46);
nand NAND3 (N2295, N2279, N1488, N1186);
and AND2 (N2296, N2281, N20);
buf BUF1 (N2297, N2288);
xor XOR2 (N2298, N2297, N1883);
buf BUF1 (N2299, N2298);
and AND3 (N2300, N2294, N979, N1800);
nand NAND4 (N2301, N2289, N217, N2111, N46);
buf BUF1 (N2302, N2292);
buf BUF1 (N2303, N2301);
xor XOR2 (N2304, N2303, N794);
nand NAND2 (N2305, N2295, N1458);
not NOT1 (N2306, N2296);
and AND4 (N2307, N2302, N2013, N1909, N1725);
nor NOR4 (N2308, N2307, N1150, N1171, N2055);
xor XOR2 (N2309, N2269, N1611);
or OR4 (N2310, N2305, N2219, N2040, N196);
nand NAND2 (N2311, N2293, N2270);
not NOT1 (N2312, N2310);
or OR3 (N2313, N2304, N1943, N59);
or OR3 (N2314, N2308, N369, N1580);
nor NOR4 (N2315, N2300, N1667, N768, N1797);
xor XOR2 (N2316, N2299, N2298);
not NOT1 (N2317, N2312);
or OR3 (N2318, N2309, N629, N1379);
nand NAND3 (N2319, N2318, N896, N947);
not NOT1 (N2320, N2317);
nor NOR2 (N2321, N2313, N1783);
not NOT1 (N2322, N2306);
xor XOR2 (N2323, N2321, N475);
and AND2 (N2324, N2322, N1070);
and AND2 (N2325, N2320, N1343);
or OR2 (N2326, N2325, N1068);
nor NOR4 (N2327, N2319, N1594, N630, N798);
nand NAND2 (N2328, N2327, N1806);
xor XOR2 (N2329, N2328, N2257);
and AND4 (N2330, N2324, N1609, N1192, N1457);
xor XOR2 (N2331, N2311, N805);
not NOT1 (N2332, N2315);
nand NAND4 (N2333, N2323, N1967, N1169, N1711);
not NOT1 (N2334, N2329);
and AND2 (N2335, N2333, N2323);
or OR2 (N2336, N2284, N1089);
xor XOR2 (N2337, N2332, N870);
and AND3 (N2338, N2326, N1501, N1837);
nor NOR3 (N2339, N2337, N2095, N358);
and AND4 (N2340, N2338, N1240, N304, N1982);
or OR2 (N2341, N2335, N1035);
buf BUF1 (N2342, N2314);
or OR2 (N2343, N2330, N1093);
nand NAND2 (N2344, N2334, N20);
buf BUF1 (N2345, N2344);
or OR3 (N2346, N2331, N633, N1083);
and AND2 (N2347, N2316, N377);
nor NOR4 (N2348, N2347, N1307, N1879, N561);
not NOT1 (N2349, N2346);
or OR2 (N2350, N2342, N1225);
and AND3 (N2351, N2350, N785, N211);
nand NAND3 (N2352, N2290, N909, N868);
buf BUF1 (N2353, N2351);
or OR4 (N2354, N2353, N2005, N1387, N1291);
and AND3 (N2355, N2349, N18, N1305);
and AND3 (N2356, N2348, N422, N1770);
nand NAND3 (N2357, N2345, N1462, N15);
and AND3 (N2358, N2356, N1980, N1555);
or OR4 (N2359, N2358, N1110, N543, N931);
nor NOR3 (N2360, N2355, N1479, N2234);
xor XOR2 (N2361, N2343, N102);
nor NOR3 (N2362, N2341, N2038, N1274);
not NOT1 (N2363, N2339);
nor NOR3 (N2364, N2359, N1298, N994);
nand NAND3 (N2365, N2336, N1837, N1879);
and AND3 (N2366, N2360, N2329, N702);
and AND2 (N2367, N2352, N2197);
and AND3 (N2368, N2366, N750, N2323);
or OR2 (N2369, N2357, N2033);
nor NOR4 (N2370, N2354, N248, N432, N2368);
and AND3 (N2371, N1973, N1262, N1461);
nand NAND3 (N2372, N2365, N308, N544);
nand NAND4 (N2373, N2370, N843, N1216, N1446);
buf BUF1 (N2374, N2369);
not NOT1 (N2375, N2372);
buf BUF1 (N2376, N2362);
nor NOR2 (N2377, N2363, N1509);
nor NOR4 (N2378, N2340, N1224, N2011, N2087);
and AND4 (N2379, N2367, N143, N1291, N2257);
and AND2 (N2380, N2378, N874);
or OR4 (N2381, N2377, N1144, N1595, N696);
and AND2 (N2382, N2373, N1739);
or OR4 (N2383, N2382, N1292, N913, N2345);
nor NOR4 (N2384, N2374, N2366, N1205, N964);
xor XOR2 (N2385, N2383, N650);
and AND4 (N2386, N2379, N1948, N45, N386);
nor NOR4 (N2387, N2364, N1368, N698, N1142);
not NOT1 (N2388, N2375);
nor NOR2 (N2389, N2388, N1065);
nand NAND4 (N2390, N2384, N629, N705, N785);
not NOT1 (N2391, N2389);
nor NOR3 (N2392, N2386, N1289, N1059);
not NOT1 (N2393, N2380);
nor NOR3 (N2394, N2391, N485, N1213);
xor XOR2 (N2395, N2390, N75);
and AND4 (N2396, N2361, N1812, N512, N2149);
nand NAND4 (N2397, N2376, N530, N271, N38);
nand NAND2 (N2398, N2396, N1756);
and AND2 (N2399, N2392, N758);
nand NAND3 (N2400, N2394, N2152, N707);
not NOT1 (N2401, N2398);
xor XOR2 (N2402, N2400, N1292);
buf BUF1 (N2403, N2381);
nor NOR2 (N2404, N2385, N18);
not NOT1 (N2405, N2402);
xor XOR2 (N2406, N2371, N2364);
and AND3 (N2407, N2393, N1730, N572);
xor XOR2 (N2408, N2407, N1796);
nor NOR3 (N2409, N2395, N999, N551);
nor NOR4 (N2410, N2408, N757, N800, N1840);
xor XOR2 (N2411, N2403, N945);
not NOT1 (N2412, N2409);
buf BUF1 (N2413, N2410);
and AND4 (N2414, N2413, N2133, N1028, N567);
or OR4 (N2415, N2399, N2398, N998, N1276);
and AND4 (N2416, N2411, N129, N1948, N1992);
not NOT1 (N2417, N2397);
xor XOR2 (N2418, N2406, N1134);
and AND4 (N2419, N2404, N883, N134, N1641);
xor XOR2 (N2420, N2415, N528);
or OR4 (N2421, N2387, N567, N1255, N984);
or OR4 (N2422, N2419, N1674, N697, N2278);
and AND4 (N2423, N2416, N475, N423, N2395);
or OR3 (N2424, N2421, N308, N1270);
xor XOR2 (N2425, N2424, N1381);
or OR4 (N2426, N2425, N2059, N498, N1469);
or OR2 (N2427, N2426, N1249);
xor XOR2 (N2428, N2417, N969);
nor NOR2 (N2429, N2428, N2210);
nand NAND4 (N2430, N2405, N326, N2406, N2094);
not NOT1 (N2431, N2427);
not NOT1 (N2432, N2418);
buf BUF1 (N2433, N2414);
not NOT1 (N2434, N2423);
nor NOR3 (N2435, N2433, N832, N283);
nor NOR2 (N2436, N2430, N2014);
nor NOR2 (N2437, N2432, N1181);
or OR3 (N2438, N2437, N330, N369);
xor XOR2 (N2439, N2431, N2059);
nand NAND3 (N2440, N2401, N549, N1087);
xor XOR2 (N2441, N2439, N2063);
not NOT1 (N2442, N2434);
nor NOR2 (N2443, N2412, N1954);
xor XOR2 (N2444, N2442, N863);
and AND4 (N2445, N2420, N1936, N2013, N243);
or OR3 (N2446, N2440, N221, N2286);
nand NAND4 (N2447, N2446, N1106, N2434, N623);
xor XOR2 (N2448, N2443, N903);
nor NOR3 (N2449, N2444, N1981, N564);
xor XOR2 (N2450, N2441, N2223);
not NOT1 (N2451, N2438);
and AND3 (N2452, N2449, N2069, N1075);
nor NOR4 (N2453, N2429, N2239, N1843, N400);
xor XOR2 (N2454, N2450, N1259);
and AND3 (N2455, N2435, N2178, N1910);
buf BUF1 (N2456, N2447);
and AND3 (N2457, N2454, N2352, N2253);
xor XOR2 (N2458, N2445, N1739);
nor NOR3 (N2459, N2458, N2283, N1806);
not NOT1 (N2460, N2422);
nor NOR3 (N2461, N2459, N1665, N1535);
nand NAND2 (N2462, N2460, N945);
or OR4 (N2463, N2452, N95, N189, N1651);
nor NOR2 (N2464, N2462, N335);
xor XOR2 (N2465, N2453, N2114);
nor NOR4 (N2466, N2456, N2008, N866, N63);
buf BUF1 (N2467, N2436);
xor XOR2 (N2468, N2465, N849);
not NOT1 (N2469, N2455);
not NOT1 (N2470, N2448);
not NOT1 (N2471, N2466);
or OR2 (N2472, N2457, N1321);
and AND3 (N2473, N2467, N2458, N317);
or OR2 (N2474, N2461, N1815);
and AND4 (N2475, N2464, N2440, N324, N1563);
not NOT1 (N2476, N2463);
nor NOR2 (N2477, N2469, N2128);
and AND4 (N2478, N2475, N2284, N1101, N827);
and AND3 (N2479, N2468, N2096, N391);
xor XOR2 (N2480, N2474, N560);
nand NAND2 (N2481, N2470, N2108);
nand NAND4 (N2482, N2478, N143, N1421, N611);
not NOT1 (N2483, N2480);
nand NAND4 (N2484, N2476, N2003, N1585, N1702);
or OR4 (N2485, N2477, N1963, N1647, N1350);
nand NAND2 (N2486, N2479, N2310);
and AND2 (N2487, N2473, N2246);
buf BUF1 (N2488, N2483);
or OR4 (N2489, N2481, N688, N778, N610);
nand NAND2 (N2490, N2485, N2329);
nor NOR2 (N2491, N2486, N1753);
nor NOR2 (N2492, N2489, N2252);
and AND2 (N2493, N2492, N2270);
or OR2 (N2494, N2490, N1303);
not NOT1 (N2495, N2472);
not NOT1 (N2496, N2487);
nand NAND2 (N2497, N2484, N1303);
xor XOR2 (N2498, N2494, N1777);
not NOT1 (N2499, N2495);
buf BUF1 (N2500, N2471);
nor NOR4 (N2501, N2496, N47, N398, N2043);
nand NAND2 (N2502, N2497, N448);
and AND3 (N2503, N2493, N2429, N460);
or OR4 (N2504, N2498, N1016, N192, N1314);
xor XOR2 (N2505, N2501, N1547);
and AND4 (N2506, N2503, N146, N2272, N1347);
xor XOR2 (N2507, N2500, N150);
buf BUF1 (N2508, N2491);
or OR4 (N2509, N2505, N677, N125, N110);
buf BUF1 (N2510, N2488);
xor XOR2 (N2511, N2509, N1985);
nor NOR2 (N2512, N2508, N1338);
not NOT1 (N2513, N2502);
nand NAND4 (N2514, N2507, N1528, N552, N430);
not NOT1 (N2515, N2512);
buf BUF1 (N2516, N2511);
xor XOR2 (N2517, N2482, N552);
buf BUF1 (N2518, N2514);
nor NOR4 (N2519, N2518, N2087, N2145, N820);
nor NOR3 (N2520, N2506, N295, N1955);
or OR3 (N2521, N2516, N187, N1169);
and AND2 (N2522, N2515, N1210);
xor XOR2 (N2523, N2520, N1974);
endmodule