// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N12798,N12814,N12812,N12813,N12808,N12817,N12810,N12816,N12788,N12818;

and AND4 (N19, N8, N15, N9, N18);
and AND2 (N20, N17, N12);
nor NOR4 (N21, N7, N19, N12, N13);
xor XOR2 (N22, N18, N15);
nor NOR2 (N23, N3, N19);
xor XOR2 (N24, N6, N15);
or OR4 (N25, N20, N17, N23, N10);
not NOT1 (N26, N19);
or OR3 (N27, N24, N14, N22);
xor XOR2 (N28, N10, N15);
nor NOR2 (N29, N20, N14);
nand NAND2 (N30, N24, N2);
not NOT1 (N31, N5);
not NOT1 (N32, N25);
and AND2 (N33, N4, N2);
xor XOR2 (N34, N4, N13);
and AND3 (N35, N31, N1, N13);
nor NOR3 (N36, N28, N35, N1);
and AND2 (N37, N19, N18);
nor NOR2 (N38, N33, N2);
and AND3 (N39, N32, N13, N16);
buf BUF1 (N40, N36);
or OR2 (N41, N21, N40);
or OR4 (N42, N11, N12, N36, N37);
or OR2 (N43, N17, N38);
and AND2 (N44, N4, N21);
xor XOR2 (N45, N27, N24);
nor NOR3 (N46, N34, N2, N15);
nor NOR2 (N47, N29, N23);
and AND4 (N48, N44, N14, N21, N21);
buf BUF1 (N49, N42);
not NOT1 (N50, N49);
nor NOR3 (N51, N48, N31, N31);
and AND2 (N52, N45, N14);
or OR4 (N53, N43, N49, N45, N20);
not NOT1 (N54, N52);
or OR2 (N55, N51, N41);
or OR3 (N56, N55, N17, N10);
or OR3 (N57, N19, N25, N17);
buf BUF1 (N58, N56);
nand NAND2 (N59, N26, N24);
nor NOR2 (N60, N53, N45);
nor NOR2 (N61, N60, N38);
not NOT1 (N62, N61);
nor NOR4 (N63, N46, N1, N17, N47);
nand NAND4 (N64, N63, N55, N49, N40);
xor XOR2 (N65, N61, N51);
xor XOR2 (N66, N57, N57);
and AND4 (N67, N30, N21, N2, N59);
and AND4 (N68, N41, N14, N10, N29);
nor NOR3 (N69, N66, N8, N50);
and AND3 (N70, N30, N50, N51);
and AND4 (N71, N70, N66, N15, N28);
not NOT1 (N72, N54);
not NOT1 (N73, N65);
not NOT1 (N74, N39);
xor XOR2 (N75, N67, N20);
or OR2 (N76, N58, N58);
xor XOR2 (N77, N75, N53);
and AND2 (N78, N69, N10);
nand NAND4 (N79, N74, N72, N7, N25);
or OR3 (N80, N61, N50, N18);
xor XOR2 (N81, N76, N54);
and AND3 (N82, N73, N62, N70);
and AND3 (N83, N71, N31, N27);
or OR4 (N84, N53, N78, N43, N49);
or OR4 (N85, N25, N8, N51, N60);
not NOT1 (N86, N82);
nand NAND3 (N87, N80, N84, N39);
and AND4 (N88, N80, N47, N16, N36);
buf BUF1 (N89, N86);
and AND3 (N90, N87, N66, N43);
nand NAND4 (N91, N85, N13, N12, N15);
and AND4 (N92, N81, N21, N46, N49);
buf BUF1 (N93, N83);
or OR4 (N94, N91, N76, N30, N1);
buf BUF1 (N95, N68);
xor XOR2 (N96, N90, N82);
or OR2 (N97, N95, N26);
or OR2 (N98, N92, N18);
and AND2 (N99, N98, N70);
and AND4 (N100, N77, N14, N98, N76);
and AND4 (N101, N99, N65, N83, N23);
nand NAND3 (N102, N96, N16, N29);
xor XOR2 (N103, N93, N65);
and AND2 (N104, N79, N64);
nor NOR4 (N105, N47, N89, N77, N34);
buf BUF1 (N106, N30);
and AND4 (N107, N105, N16, N45, N88);
or OR2 (N108, N23, N67);
nand NAND3 (N109, N94, N83, N34);
nand NAND2 (N110, N100, N104);
xor XOR2 (N111, N67, N95);
not NOT1 (N112, N110);
buf BUF1 (N113, N102);
nand NAND3 (N114, N101, N113, N23);
or OR3 (N115, N26, N19, N54);
and AND3 (N116, N97, N81, N65);
not NOT1 (N117, N108);
xor XOR2 (N118, N107, N36);
nor NOR4 (N119, N115, N28, N86, N92);
nor NOR3 (N120, N119, N86, N22);
not NOT1 (N121, N114);
nand NAND3 (N122, N117, N27, N56);
nor NOR4 (N123, N111, N120, N4, N80);
nand NAND2 (N124, N42, N23);
nand NAND4 (N125, N124, N44, N23, N8);
nand NAND3 (N126, N116, N41, N32);
xor XOR2 (N127, N126, N117);
buf BUF1 (N128, N112);
nor NOR3 (N129, N118, N106, N106);
buf BUF1 (N130, N93);
xor XOR2 (N131, N109, N65);
buf BUF1 (N132, N127);
nor NOR4 (N133, N132, N47, N132, N113);
nand NAND4 (N134, N133, N81, N20, N12);
not NOT1 (N135, N103);
nor NOR4 (N136, N129, N10, N111, N61);
or OR4 (N137, N121, N49, N6, N112);
buf BUF1 (N138, N136);
buf BUF1 (N139, N137);
not NOT1 (N140, N138);
nor NOR4 (N141, N140, N76, N33, N87);
or OR3 (N142, N128, N62, N32);
xor XOR2 (N143, N139, N54);
nand NAND2 (N144, N141, N121);
xor XOR2 (N145, N135, N7);
not NOT1 (N146, N145);
xor XOR2 (N147, N144, N56);
nor NOR2 (N148, N146, N26);
nand NAND4 (N149, N123, N59, N79, N53);
buf BUF1 (N150, N142);
not NOT1 (N151, N134);
buf BUF1 (N152, N147);
xor XOR2 (N153, N143, N151);
or OR2 (N154, N149, N35);
xor XOR2 (N155, N20, N102);
or OR3 (N156, N150, N48, N9);
xor XOR2 (N157, N131, N99);
or OR3 (N158, N157, N49, N78);
nand NAND3 (N159, N156, N43, N135);
buf BUF1 (N160, N154);
nor NOR4 (N161, N125, N28, N149, N2);
xor XOR2 (N162, N122, N82);
or OR2 (N163, N158, N122);
or OR3 (N164, N163, N48, N104);
xor XOR2 (N165, N130, N157);
nor NOR3 (N166, N155, N44, N164);
and AND3 (N167, N49, N60, N14);
nor NOR3 (N168, N148, N61, N82);
buf BUF1 (N169, N153);
nand NAND3 (N170, N162, N5, N25);
not NOT1 (N171, N169);
nor NOR2 (N172, N170, N76);
xor XOR2 (N173, N159, N116);
nor NOR2 (N174, N160, N29);
buf BUF1 (N175, N161);
buf BUF1 (N176, N167);
xor XOR2 (N177, N166, N26);
and AND3 (N178, N173, N99, N146);
nand NAND4 (N179, N152, N30, N81, N121);
not NOT1 (N180, N176);
or OR3 (N181, N180, N77, N145);
or OR4 (N182, N171, N99, N165, N41);
buf BUF1 (N183, N98);
nor NOR3 (N184, N181, N165, N128);
nand NAND3 (N185, N174, N142, N1);
buf BUF1 (N186, N182);
nor NOR3 (N187, N183, N35, N62);
xor XOR2 (N188, N178, N15);
not NOT1 (N189, N172);
not NOT1 (N190, N177);
nor NOR3 (N191, N185, N167, N64);
xor XOR2 (N192, N189, N128);
and AND4 (N193, N191, N45, N50, N110);
and AND4 (N194, N188, N161, N75, N39);
xor XOR2 (N195, N168, N52);
buf BUF1 (N196, N187);
or OR4 (N197, N196, N149, N15, N51);
xor XOR2 (N198, N186, N126);
and AND3 (N199, N184, N70, N115);
nor NOR4 (N200, N194, N108, N65, N98);
not NOT1 (N201, N179);
nand NAND2 (N202, N193, N112);
or OR2 (N203, N200, N107);
or OR2 (N204, N197, N102);
not NOT1 (N205, N203);
not NOT1 (N206, N175);
not NOT1 (N207, N206);
not NOT1 (N208, N198);
not NOT1 (N209, N195);
nor NOR2 (N210, N209, N199);
not NOT1 (N211, N118);
nand NAND3 (N212, N211, N32, N133);
nand NAND2 (N213, N208, N193);
not NOT1 (N214, N190);
nor NOR3 (N215, N192, N199, N138);
nor NOR2 (N216, N213, N18);
xor XOR2 (N217, N212, N171);
nand NAND2 (N218, N201, N92);
not NOT1 (N219, N218);
xor XOR2 (N220, N210, N36);
buf BUF1 (N221, N202);
nor NOR4 (N222, N204, N156, N193, N60);
not NOT1 (N223, N217);
buf BUF1 (N224, N220);
or OR4 (N225, N207, N81, N76, N13);
not NOT1 (N226, N223);
not NOT1 (N227, N222);
or OR3 (N228, N205, N137, N197);
and AND2 (N229, N216, N111);
xor XOR2 (N230, N215, N205);
not NOT1 (N231, N228);
nand NAND4 (N232, N214, N188, N64, N71);
nand NAND3 (N233, N226, N54, N9);
xor XOR2 (N234, N224, N37);
not NOT1 (N235, N225);
xor XOR2 (N236, N221, N77);
xor XOR2 (N237, N231, N219);
nand NAND2 (N238, N223, N113);
xor XOR2 (N239, N238, N70);
not NOT1 (N240, N236);
nor NOR4 (N241, N232, N60, N214, N223);
not NOT1 (N242, N240);
and AND2 (N243, N229, N126);
and AND3 (N244, N237, N159, N97);
not NOT1 (N245, N234);
or OR2 (N246, N241, N44);
nor NOR3 (N247, N245, N184, N224);
and AND4 (N248, N227, N85, N205, N200);
or OR4 (N249, N233, N14, N61, N222);
xor XOR2 (N250, N235, N98);
nor NOR3 (N251, N244, N200, N49);
nor NOR4 (N252, N242, N80, N110, N113);
nor NOR4 (N253, N251, N235, N172, N66);
nor NOR4 (N254, N230, N155, N54, N123);
or OR3 (N255, N246, N245, N223);
buf BUF1 (N256, N250);
not NOT1 (N257, N254);
nor NOR2 (N258, N243, N13);
nor NOR4 (N259, N248, N47, N54, N78);
xor XOR2 (N260, N253, N73);
buf BUF1 (N261, N259);
or OR4 (N262, N257, N40, N4, N85);
nand NAND2 (N263, N258, N215);
nor NOR2 (N264, N247, N50);
not NOT1 (N265, N255);
not NOT1 (N266, N256);
nor NOR3 (N267, N239, N2, N99);
and AND2 (N268, N262, N258);
and AND3 (N269, N267, N67, N178);
buf BUF1 (N270, N269);
and AND4 (N271, N266, N213, N162, N162);
not NOT1 (N272, N263);
xor XOR2 (N273, N272, N42);
not NOT1 (N274, N271);
nor NOR4 (N275, N265, N228, N125, N74);
or OR4 (N276, N252, N128, N236, N157);
and AND3 (N277, N268, N218, N190);
nor NOR3 (N278, N260, N262, N168);
xor XOR2 (N279, N278, N258);
or OR3 (N280, N275, N277, N268);
nand NAND2 (N281, N248, N277);
nand NAND2 (N282, N281, N106);
nand NAND4 (N283, N249, N197, N195, N38);
and AND3 (N284, N274, N163, N123);
nand NAND4 (N285, N270, N11, N231, N279);
not NOT1 (N286, N217);
xor XOR2 (N287, N283, N108);
or OR3 (N288, N264, N64, N38);
not NOT1 (N289, N285);
nor NOR2 (N290, N282, N167);
or OR3 (N291, N286, N272, N142);
nand NAND3 (N292, N261, N288, N171);
nand NAND3 (N293, N174, N129, N70);
and AND2 (N294, N287, N189);
xor XOR2 (N295, N290, N89);
or OR3 (N296, N276, N280, N150);
not NOT1 (N297, N101);
and AND2 (N298, N297, N136);
nor NOR4 (N299, N292, N234, N115, N250);
and AND3 (N300, N299, N132, N64);
or OR3 (N301, N295, N251, N117);
nor NOR4 (N302, N273, N2, N215, N116);
not NOT1 (N303, N301);
buf BUF1 (N304, N296);
or OR3 (N305, N294, N151, N207);
nand NAND3 (N306, N304, N286, N50);
nand NAND3 (N307, N289, N229, N86);
nand NAND2 (N308, N305, N119);
not NOT1 (N309, N300);
and AND4 (N310, N308, N177, N215, N169);
not NOT1 (N311, N309);
not NOT1 (N312, N310);
nand NAND3 (N313, N302, N280, N68);
not NOT1 (N314, N298);
not NOT1 (N315, N307);
nand NAND3 (N316, N303, N148, N129);
nor NOR3 (N317, N315, N161, N56);
xor XOR2 (N318, N312, N237);
nand NAND4 (N319, N293, N117, N213, N197);
and AND4 (N320, N316, N89, N255, N67);
xor XOR2 (N321, N311, N202);
nand NAND4 (N322, N313, N189, N166, N180);
xor XOR2 (N323, N284, N169);
or OR2 (N324, N322, N78);
xor XOR2 (N325, N324, N151);
or OR2 (N326, N314, N183);
buf BUF1 (N327, N306);
xor XOR2 (N328, N326, N277);
nand NAND4 (N329, N319, N306, N198, N167);
nor NOR3 (N330, N320, N173, N129);
not NOT1 (N331, N291);
buf BUF1 (N332, N325);
nand NAND3 (N333, N327, N69, N85);
nor NOR4 (N334, N331, N194, N238, N19);
xor XOR2 (N335, N334, N278);
nand NAND3 (N336, N333, N218, N245);
xor XOR2 (N337, N336, N310);
nor NOR4 (N338, N321, N31, N315, N322);
nand NAND3 (N339, N328, N42, N71);
buf BUF1 (N340, N337);
or OR3 (N341, N330, N9, N210);
buf BUF1 (N342, N318);
buf BUF1 (N343, N323);
and AND4 (N344, N335, N163, N319, N262);
xor XOR2 (N345, N338, N121);
and AND2 (N346, N342, N128);
xor XOR2 (N347, N317, N72);
xor XOR2 (N348, N339, N49);
not NOT1 (N349, N332);
not NOT1 (N350, N329);
nand NAND4 (N351, N350, N273, N275, N344);
not NOT1 (N352, N108);
not NOT1 (N353, N340);
and AND2 (N354, N352, N266);
xor XOR2 (N355, N348, N96);
nand NAND3 (N356, N343, N304, N324);
not NOT1 (N357, N349);
and AND3 (N358, N354, N106, N20);
nand NAND4 (N359, N341, N342, N319, N66);
nor NOR3 (N360, N355, N150, N297);
nand NAND4 (N361, N357, N179, N255, N132);
nor NOR4 (N362, N356, N327, N332, N341);
not NOT1 (N363, N351);
and AND4 (N364, N353, N87, N340, N189);
and AND3 (N365, N363, N67, N278);
buf BUF1 (N366, N345);
buf BUF1 (N367, N361);
not NOT1 (N368, N358);
nand NAND4 (N369, N366, N206, N69, N217);
xor XOR2 (N370, N364, N244);
or OR4 (N371, N346, N256, N326, N354);
or OR4 (N372, N359, N105, N153, N3);
and AND4 (N373, N367, N245, N347, N171);
buf BUF1 (N374, N30);
nand NAND4 (N375, N365, N295, N356, N178);
nor NOR4 (N376, N362, N122, N286, N231);
nor NOR4 (N377, N360, N55, N83, N248);
xor XOR2 (N378, N370, N133);
and AND3 (N379, N372, N65, N290);
nand NAND3 (N380, N376, N13, N300);
not NOT1 (N381, N378);
or OR4 (N382, N369, N92, N166, N3);
or OR3 (N383, N375, N250, N160);
buf BUF1 (N384, N377);
and AND2 (N385, N371, N354);
or OR2 (N386, N374, N336);
buf BUF1 (N387, N383);
nand NAND2 (N388, N386, N302);
and AND3 (N389, N373, N49, N64);
nand NAND4 (N390, N384, N273, N267, N175);
or OR2 (N391, N389, N23);
nand NAND3 (N392, N385, N374, N14);
or OR2 (N393, N379, N16);
or OR3 (N394, N390, N240, N171);
or OR3 (N395, N394, N348, N50);
xor XOR2 (N396, N380, N19);
nand NAND3 (N397, N382, N344, N167);
not NOT1 (N398, N387);
nor NOR2 (N399, N395, N170);
nor NOR4 (N400, N398, N148, N172, N18);
nand NAND2 (N401, N368, N229);
nor NOR2 (N402, N401, N82);
xor XOR2 (N403, N393, N268);
and AND4 (N404, N392, N94, N386, N98);
xor XOR2 (N405, N391, N336);
buf BUF1 (N406, N396);
not NOT1 (N407, N403);
or OR2 (N408, N407, N109);
buf BUF1 (N409, N408);
xor XOR2 (N410, N404, N153);
buf BUF1 (N411, N402);
nand NAND3 (N412, N406, N71, N242);
xor XOR2 (N413, N399, N265);
nor NOR4 (N414, N412, N285, N138, N262);
buf BUF1 (N415, N388);
buf BUF1 (N416, N409);
xor XOR2 (N417, N397, N268);
and AND3 (N418, N400, N76, N386);
xor XOR2 (N419, N381, N404);
buf BUF1 (N420, N411);
not NOT1 (N421, N415);
nor NOR3 (N422, N421, N209, N294);
nand NAND2 (N423, N422, N109);
nand NAND2 (N424, N413, N387);
nor NOR2 (N425, N423, N174);
not NOT1 (N426, N420);
or OR2 (N427, N424, N310);
nand NAND4 (N428, N410, N376, N5, N80);
not NOT1 (N429, N428);
not NOT1 (N430, N417);
nor NOR4 (N431, N418, N198, N87, N336);
not NOT1 (N432, N427);
not NOT1 (N433, N432);
nand NAND2 (N434, N430, N275);
or OR2 (N435, N416, N391);
xor XOR2 (N436, N405, N402);
nor NOR2 (N437, N426, N257);
buf BUF1 (N438, N435);
nand NAND4 (N439, N438, N201, N203, N268);
xor XOR2 (N440, N437, N409);
xor XOR2 (N441, N429, N173);
nand NAND2 (N442, N431, N22);
not NOT1 (N443, N436);
or OR2 (N444, N414, N375);
or OR3 (N445, N419, N422, N108);
nor NOR4 (N446, N440, N196, N89, N209);
buf BUF1 (N447, N433);
not NOT1 (N448, N442);
nor NOR3 (N449, N443, N34, N245);
xor XOR2 (N450, N439, N198);
not NOT1 (N451, N447);
nor NOR2 (N452, N445, N389);
not NOT1 (N453, N452);
or OR3 (N454, N449, N223, N255);
buf BUF1 (N455, N446);
not NOT1 (N456, N454);
nor NOR4 (N457, N434, N235, N157, N148);
nor NOR2 (N458, N441, N369);
and AND3 (N459, N456, N59, N45);
nand NAND4 (N460, N450, N244, N97, N450);
xor XOR2 (N461, N455, N138);
nand NAND3 (N462, N459, N255, N325);
or OR3 (N463, N457, N343, N310);
not NOT1 (N464, N448);
and AND3 (N465, N460, N12, N6);
or OR3 (N466, N462, N118, N197);
or OR2 (N467, N464, N108);
or OR4 (N468, N425, N322, N141, N202);
and AND3 (N469, N468, N65, N326);
nor NOR4 (N470, N461, N365, N410, N395);
nand NAND4 (N471, N458, N225, N49, N402);
or OR2 (N472, N463, N228);
xor XOR2 (N473, N444, N101);
or OR3 (N474, N473, N251, N28);
and AND2 (N475, N451, N224);
nand NAND3 (N476, N472, N134, N293);
not NOT1 (N477, N471);
and AND3 (N478, N475, N75, N271);
nand NAND3 (N479, N478, N441, N288);
nor NOR4 (N480, N477, N446, N162, N262);
xor XOR2 (N481, N480, N319);
buf BUF1 (N482, N474);
nand NAND2 (N483, N469, N207);
nor NOR3 (N484, N453, N76, N340);
not NOT1 (N485, N483);
xor XOR2 (N486, N479, N47);
buf BUF1 (N487, N476);
nor NOR4 (N488, N487, N191, N61, N398);
xor XOR2 (N489, N484, N280);
buf BUF1 (N490, N485);
nor NOR3 (N491, N482, N232, N251);
buf BUF1 (N492, N466);
nand NAND4 (N493, N488, N290, N21, N447);
nor NOR3 (N494, N465, N242, N297);
buf BUF1 (N495, N494);
and AND3 (N496, N486, N448, N30);
buf BUF1 (N497, N470);
or OR3 (N498, N467, N414, N134);
or OR3 (N499, N493, N373, N442);
nor NOR4 (N500, N481, N184, N94, N334);
xor XOR2 (N501, N490, N154);
buf BUF1 (N502, N496);
buf BUF1 (N503, N498);
buf BUF1 (N504, N491);
buf BUF1 (N505, N500);
or OR4 (N506, N501, N454, N475, N413);
or OR3 (N507, N497, N1, N155);
xor XOR2 (N508, N505, N474);
nor NOR3 (N509, N489, N374, N359);
buf BUF1 (N510, N492);
and AND4 (N511, N499, N203, N248, N296);
not NOT1 (N512, N511);
buf BUF1 (N513, N506);
buf BUF1 (N514, N509);
nand NAND3 (N515, N503, N273, N92);
nor NOR3 (N516, N515, N454, N245);
and AND3 (N517, N514, N322, N367);
buf BUF1 (N518, N510);
and AND4 (N519, N508, N267, N471, N400);
or OR3 (N520, N495, N414, N430);
xor XOR2 (N521, N512, N117);
or OR2 (N522, N520, N22);
nand NAND3 (N523, N513, N271, N222);
buf BUF1 (N524, N517);
nor NOR3 (N525, N516, N469, N479);
nor NOR2 (N526, N525, N492);
and AND2 (N527, N518, N91);
buf BUF1 (N528, N521);
nand NAND3 (N529, N522, N120, N133);
xor XOR2 (N530, N524, N57);
xor XOR2 (N531, N528, N267);
not NOT1 (N532, N527);
xor XOR2 (N533, N502, N139);
nor NOR2 (N534, N507, N253);
or OR3 (N535, N530, N210, N211);
and AND3 (N536, N533, N312, N517);
nand NAND3 (N537, N532, N374, N59);
nand NAND2 (N538, N504, N231);
xor XOR2 (N539, N535, N462);
buf BUF1 (N540, N538);
buf BUF1 (N541, N523);
buf BUF1 (N542, N529);
nand NAND2 (N543, N526, N152);
not NOT1 (N544, N539);
xor XOR2 (N545, N531, N529);
or OR2 (N546, N534, N326);
nand NAND3 (N547, N537, N409, N184);
or OR3 (N548, N545, N405, N431);
xor XOR2 (N549, N546, N80);
and AND4 (N550, N544, N505, N493, N118);
nand NAND3 (N551, N550, N534, N40);
and AND3 (N552, N536, N46, N407);
not NOT1 (N553, N547);
nor NOR3 (N554, N553, N136, N308);
buf BUF1 (N555, N519);
xor XOR2 (N556, N552, N456);
or OR3 (N557, N541, N183, N276);
and AND2 (N558, N551, N100);
nand NAND3 (N559, N557, N134, N347);
or OR3 (N560, N543, N275, N404);
buf BUF1 (N561, N560);
xor XOR2 (N562, N555, N120);
or OR4 (N563, N562, N3, N143, N504);
nor NOR2 (N564, N549, N195);
and AND2 (N565, N548, N434);
buf BUF1 (N566, N565);
xor XOR2 (N567, N542, N210);
and AND4 (N568, N556, N51, N294, N316);
buf BUF1 (N569, N566);
nor NOR4 (N570, N563, N569, N267, N543);
xor XOR2 (N571, N259, N410);
buf BUF1 (N572, N554);
not NOT1 (N573, N570);
nor NOR2 (N574, N540, N355);
nor NOR4 (N575, N558, N279, N558, N270);
or OR4 (N576, N572, N273, N210, N569);
and AND2 (N577, N575, N399);
not NOT1 (N578, N574);
xor XOR2 (N579, N573, N347);
and AND2 (N580, N578, N264);
buf BUF1 (N581, N564);
buf BUF1 (N582, N571);
not NOT1 (N583, N567);
and AND3 (N584, N582, N498, N195);
nor NOR3 (N585, N581, N431, N381);
not NOT1 (N586, N568);
and AND3 (N587, N576, N82, N299);
nor NOR4 (N588, N584, N316, N265, N368);
and AND3 (N589, N579, N235, N552);
xor XOR2 (N590, N583, N116);
or OR3 (N591, N559, N170, N320);
nor NOR4 (N592, N561, N447, N588, N265);
xor XOR2 (N593, N532, N201);
nor NOR4 (N594, N593, N489, N343, N541);
and AND4 (N595, N589, N154, N3, N297);
not NOT1 (N596, N594);
nor NOR3 (N597, N587, N458, N161);
nand NAND4 (N598, N577, N16, N79, N445);
or OR3 (N599, N586, N246, N207);
and AND3 (N600, N580, N27, N503);
nor NOR4 (N601, N596, N105, N203, N62);
buf BUF1 (N602, N585);
nand NAND3 (N603, N600, N89, N414);
xor XOR2 (N604, N591, N370);
buf BUF1 (N605, N592);
nor NOR2 (N606, N598, N581);
not NOT1 (N607, N604);
buf BUF1 (N608, N601);
not NOT1 (N609, N590);
buf BUF1 (N610, N595);
not NOT1 (N611, N605);
nor NOR2 (N612, N597, N374);
xor XOR2 (N613, N610, N391);
xor XOR2 (N614, N611, N411);
not NOT1 (N615, N599);
buf BUF1 (N616, N603);
xor XOR2 (N617, N613, N611);
nand NAND4 (N618, N609, N611, N569, N45);
and AND2 (N619, N614, N485);
not NOT1 (N620, N602);
nor NOR4 (N621, N607, N145, N572, N458);
nand NAND2 (N622, N619, N426);
nand NAND4 (N623, N615, N609, N485, N219);
buf BUF1 (N624, N623);
buf BUF1 (N625, N617);
nand NAND3 (N626, N608, N103, N365);
xor XOR2 (N627, N616, N165);
nor NOR2 (N628, N621, N347);
nand NAND3 (N629, N626, N353, N430);
and AND3 (N630, N627, N622, N220);
nand NAND3 (N631, N509, N280, N242);
and AND3 (N632, N618, N9, N263);
or OR2 (N633, N632, N430);
or OR4 (N634, N630, N414, N221, N176);
not NOT1 (N635, N624);
nand NAND3 (N636, N628, N335, N267);
not NOT1 (N637, N620);
nand NAND3 (N638, N637, N433, N230);
buf BUF1 (N639, N612);
nand NAND3 (N640, N638, N557, N204);
nand NAND4 (N641, N633, N81, N62, N506);
nand NAND4 (N642, N634, N211, N288, N328);
and AND2 (N643, N641, N602);
nor NOR4 (N644, N606, N297, N607, N378);
buf BUF1 (N645, N644);
or OR4 (N646, N640, N376, N420, N519);
buf BUF1 (N647, N646);
buf BUF1 (N648, N625);
not NOT1 (N649, N639);
and AND2 (N650, N647, N224);
nor NOR2 (N651, N643, N80);
and AND4 (N652, N642, N651, N599, N436);
buf BUF1 (N653, N111);
buf BUF1 (N654, N650);
or OR2 (N655, N654, N129);
and AND4 (N656, N645, N326, N330, N489);
xor XOR2 (N657, N653, N248);
nor NOR4 (N658, N657, N11, N69, N154);
xor XOR2 (N659, N649, N551);
and AND4 (N660, N652, N107, N310, N625);
nor NOR3 (N661, N658, N479, N528);
and AND2 (N662, N660, N203);
buf BUF1 (N663, N648);
and AND4 (N664, N656, N26, N181, N526);
or OR3 (N665, N663, N507, N215);
nand NAND3 (N666, N661, N9, N303);
and AND2 (N667, N629, N535);
nor NOR3 (N668, N664, N584, N136);
or OR3 (N669, N635, N554, N550);
nand NAND3 (N670, N662, N304, N180);
xor XOR2 (N671, N659, N384);
or OR2 (N672, N665, N331);
xor XOR2 (N673, N668, N77);
nand NAND4 (N674, N669, N343, N54, N305);
nor NOR3 (N675, N670, N204, N215);
xor XOR2 (N676, N666, N365);
buf BUF1 (N677, N673);
and AND2 (N678, N671, N123);
or OR4 (N679, N667, N329, N458, N523);
and AND2 (N680, N672, N463);
and AND2 (N681, N675, N629);
xor XOR2 (N682, N681, N47);
or OR4 (N683, N631, N109, N93, N120);
xor XOR2 (N684, N655, N24);
nor NOR3 (N685, N676, N516, N147);
nor NOR3 (N686, N677, N281, N137);
buf BUF1 (N687, N678);
xor XOR2 (N688, N683, N275);
buf BUF1 (N689, N679);
or OR4 (N690, N687, N197, N285, N137);
nor NOR4 (N691, N674, N681, N270, N362);
or OR3 (N692, N682, N121, N612);
xor XOR2 (N693, N690, N189);
buf BUF1 (N694, N688);
or OR4 (N695, N684, N492, N29, N53);
buf BUF1 (N696, N695);
not NOT1 (N697, N693);
not NOT1 (N698, N685);
buf BUF1 (N699, N689);
or OR4 (N700, N680, N429, N431, N34);
buf BUF1 (N701, N691);
nor NOR3 (N702, N697, N639, N241);
xor XOR2 (N703, N698, N586);
and AND2 (N704, N699, N333);
xor XOR2 (N705, N694, N336);
and AND4 (N706, N703, N24, N162, N647);
xor XOR2 (N707, N696, N271);
and AND3 (N708, N636, N573, N173);
and AND2 (N709, N704, N331);
and AND2 (N710, N706, N561);
nor NOR4 (N711, N708, N344, N220, N404);
or OR3 (N712, N709, N700, N10);
not NOT1 (N713, N452);
buf BUF1 (N714, N705);
nor NOR3 (N715, N714, N658, N186);
or OR4 (N716, N712, N655, N241, N499);
nor NOR2 (N717, N711, N667);
xor XOR2 (N718, N707, N217);
nand NAND4 (N719, N717, N287, N387, N556);
or OR3 (N720, N686, N332, N656);
or OR2 (N721, N692, N353);
xor XOR2 (N722, N719, N719);
xor XOR2 (N723, N718, N219);
nand NAND3 (N724, N723, N706, N291);
or OR2 (N725, N720, N451);
and AND4 (N726, N702, N144, N233, N81);
xor XOR2 (N727, N726, N672);
or OR3 (N728, N724, N192, N105);
nand NAND2 (N729, N716, N249);
and AND4 (N730, N722, N670, N310, N690);
and AND4 (N731, N728, N92, N411, N639);
or OR4 (N732, N710, N552, N228, N489);
buf BUF1 (N733, N731);
nand NAND2 (N734, N701, N316);
and AND2 (N735, N734, N361);
xor XOR2 (N736, N727, N58);
and AND2 (N737, N713, N583);
xor XOR2 (N738, N732, N185);
xor XOR2 (N739, N735, N735);
nand NAND2 (N740, N737, N137);
nor NOR2 (N741, N739, N566);
not NOT1 (N742, N729);
and AND4 (N743, N715, N542, N71, N636);
and AND2 (N744, N721, N70);
not NOT1 (N745, N738);
not NOT1 (N746, N743);
buf BUF1 (N747, N745);
or OR4 (N748, N736, N59, N377, N289);
nand NAND4 (N749, N746, N350, N138, N441);
nand NAND2 (N750, N748, N480);
and AND4 (N751, N740, N556, N121, N365);
and AND4 (N752, N749, N349, N323, N554);
nand NAND3 (N753, N752, N96, N687);
nor NOR3 (N754, N744, N41, N707);
xor XOR2 (N755, N725, N682);
or OR4 (N756, N747, N349, N666, N350);
buf BUF1 (N757, N753);
nand NAND3 (N758, N756, N442, N567);
nand NAND2 (N759, N757, N559);
xor XOR2 (N760, N755, N350);
not NOT1 (N761, N758);
nor NOR2 (N762, N751, N31);
or OR3 (N763, N760, N528, N281);
nor NOR3 (N764, N761, N538, N550);
or OR3 (N765, N733, N443, N496);
or OR2 (N766, N754, N704);
nand NAND4 (N767, N765, N364, N203, N544);
not NOT1 (N768, N759);
buf BUF1 (N769, N730);
not NOT1 (N770, N764);
nor NOR2 (N771, N750, N281);
nor NOR3 (N772, N763, N138, N699);
not NOT1 (N773, N770);
and AND2 (N774, N771, N169);
or OR3 (N775, N774, N271, N63);
xor XOR2 (N776, N772, N188);
nor NOR3 (N777, N742, N632, N133);
nor NOR3 (N778, N766, N68, N5);
nand NAND4 (N779, N775, N633, N29, N660);
and AND3 (N780, N768, N160, N386);
not NOT1 (N781, N776);
nand NAND4 (N782, N779, N568, N185, N188);
buf BUF1 (N783, N778);
and AND2 (N784, N741, N645);
nor NOR4 (N785, N767, N66, N97, N547);
nor NOR3 (N786, N782, N751, N345);
buf BUF1 (N787, N786);
and AND3 (N788, N784, N199, N227);
nor NOR4 (N789, N773, N1, N62, N318);
nor NOR3 (N790, N781, N766, N80);
or OR4 (N791, N788, N688, N75, N739);
buf BUF1 (N792, N787);
nand NAND3 (N793, N783, N213, N366);
not NOT1 (N794, N780);
buf BUF1 (N795, N790);
nor NOR4 (N796, N792, N711, N234, N689);
or OR2 (N797, N795, N693);
and AND2 (N798, N762, N43);
nor NOR4 (N799, N793, N514, N740, N587);
and AND3 (N800, N796, N775, N131);
nand NAND3 (N801, N777, N637, N56);
nor NOR2 (N802, N797, N663);
or OR4 (N803, N801, N677, N518, N123);
xor XOR2 (N804, N791, N423);
not NOT1 (N805, N799);
or OR2 (N806, N805, N570);
and AND4 (N807, N789, N79, N508, N449);
and AND4 (N808, N794, N138, N46, N345);
or OR3 (N809, N803, N204, N598);
or OR4 (N810, N785, N258, N454, N362);
and AND4 (N811, N798, N555, N16, N41);
or OR2 (N812, N806, N251);
xor XOR2 (N813, N809, N233);
buf BUF1 (N814, N808);
and AND4 (N815, N802, N559, N382, N550);
xor XOR2 (N816, N810, N188);
buf BUF1 (N817, N804);
or OR2 (N818, N816, N371);
nand NAND3 (N819, N800, N249, N500);
or OR2 (N820, N815, N786);
and AND4 (N821, N807, N761, N549, N742);
xor XOR2 (N822, N818, N579);
not NOT1 (N823, N817);
xor XOR2 (N824, N769, N342);
or OR2 (N825, N812, N440);
nor NOR3 (N826, N820, N194, N785);
and AND4 (N827, N813, N621, N701, N445);
nor NOR4 (N828, N821, N534, N156, N349);
nand NAND4 (N829, N823, N709, N460, N488);
nand NAND4 (N830, N825, N322, N781, N403);
buf BUF1 (N831, N811);
nor NOR3 (N832, N814, N352, N661);
or OR3 (N833, N830, N93, N1);
and AND4 (N834, N829, N327, N572, N490);
or OR2 (N835, N826, N776);
xor XOR2 (N836, N832, N241);
not NOT1 (N837, N833);
not NOT1 (N838, N836);
nor NOR3 (N839, N828, N298, N479);
not NOT1 (N840, N824);
and AND4 (N841, N831, N674, N237, N652);
and AND3 (N842, N819, N516, N516);
not NOT1 (N843, N834);
and AND2 (N844, N835, N493);
buf BUF1 (N845, N822);
buf BUF1 (N846, N844);
not NOT1 (N847, N838);
or OR3 (N848, N845, N287, N307);
or OR3 (N849, N837, N152, N668);
not NOT1 (N850, N843);
not NOT1 (N851, N827);
or OR2 (N852, N841, N603);
or OR4 (N853, N848, N428, N751, N290);
not NOT1 (N854, N839);
buf BUF1 (N855, N854);
or OR3 (N856, N849, N830, N691);
buf BUF1 (N857, N842);
and AND3 (N858, N853, N207, N615);
nor NOR2 (N859, N856, N162);
and AND2 (N860, N847, N515);
nand NAND3 (N861, N857, N46, N790);
nand NAND4 (N862, N861, N462, N301, N758);
nand NAND3 (N863, N859, N762, N257);
and AND4 (N864, N863, N267, N708, N752);
nor NOR4 (N865, N862, N319, N680, N431);
nor NOR2 (N866, N858, N330);
and AND4 (N867, N865, N267, N299, N607);
not NOT1 (N868, N866);
buf BUF1 (N869, N855);
or OR4 (N870, N852, N401, N481, N323);
and AND2 (N871, N869, N100);
xor XOR2 (N872, N867, N191);
not NOT1 (N873, N872);
xor XOR2 (N874, N850, N350);
buf BUF1 (N875, N860);
xor XOR2 (N876, N874, N137);
nand NAND4 (N877, N873, N59, N448, N468);
not NOT1 (N878, N877);
nand NAND3 (N879, N868, N37, N127);
buf BUF1 (N880, N876);
and AND4 (N881, N879, N569, N313, N591);
or OR3 (N882, N871, N434, N254);
nand NAND3 (N883, N851, N517, N710);
nor NOR4 (N884, N880, N49, N729, N106);
and AND4 (N885, N840, N238, N75, N678);
nor NOR4 (N886, N881, N835, N345, N706);
and AND2 (N887, N875, N615);
not NOT1 (N888, N884);
buf BUF1 (N889, N882);
and AND2 (N890, N889, N228);
xor XOR2 (N891, N890, N807);
nor NOR3 (N892, N883, N175, N597);
not NOT1 (N893, N846);
and AND2 (N894, N887, N605);
buf BUF1 (N895, N892);
not NOT1 (N896, N893);
or OR4 (N897, N895, N202, N357, N348);
not NOT1 (N898, N894);
or OR2 (N899, N870, N297);
nand NAND3 (N900, N896, N579, N737);
xor XOR2 (N901, N891, N876);
and AND4 (N902, N886, N384, N764, N109);
nor NOR3 (N903, N901, N368, N568);
and AND2 (N904, N888, N322);
or OR4 (N905, N878, N334, N685, N524);
nor NOR2 (N906, N897, N398);
xor XOR2 (N907, N864, N660);
and AND4 (N908, N904, N799, N645, N366);
xor XOR2 (N909, N906, N102);
nand NAND3 (N910, N909, N482, N773);
or OR2 (N911, N898, N699);
or OR2 (N912, N900, N705);
nor NOR3 (N913, N903, N37, N336);
or OR2 (N914, N885, N149);
buf BUF1 (N915, N905);
and AND2 (N916, N914, N747);
buf BUF1 (N917, N912);
nor NOR4 (N918, N915, N852, N394, N194);
not NOT1 (N919, N916);
nor NOR3 (N920, N902, N758, N573);
or OR4 (N921, N911, N896, N458, N283);
or OR2 (N922, N919, N568);
not NOT1 (N923, N907);
buf BUF1 (N924, N918);
nor NOR4 (N925, N899, N228, N837, N277);
nand NAND2 (N926, N922, N613);
not NOT1 (N927, N908);
xor XOR2 (N928, N921, N252);
nand NAND4 (N929, N920, N272, N254, N890);
nor NOR4 (N930, N928, N661, N71, N245);
nor NOR4 (N931, N913, N117, N418, N171);
not NOT1 (N932, N929);
buf BUF1 (N933, N932);
buf BUF1 (N934, N924);
xor XOR2 (N935, N917, N897);
not NOT1 (N936, N923);
nand NAND2 (N937, N935, N477);
nand NAND3 (N938, N934, N648, N925);
xor XOR2 (N939, N414, N469);
nand NAND4 (N940, N931, N432, N516, N888);
xor XOR2 (N941, N930, N119);
or OR4 (N942, N910, N739, N500, N804);
nor NOR4 (N943, N936, N388, N559, N408);
nor NOR4 (N944, N926, N665, N275, N661);
not NOT1 (N945, N944);
buf BUF1 (N946, N933);
buf BUF1 (N947, N938);
xor XOR2 (N948, N945, N73);
buf BUF1 (N949, N927);
xor XOR2 (N950, N947, N372);
xor XOR2 (N951, N939, N877);
xor XOR2 (N952, N951, N744);
nand NAND4 (N953, N948, N492, N35, N4);
nand NAND3 (N954, N943, N409, N644);
nor NOR4 (N955, N952, N71, N92, N243);
and AND4 (N956, N954, N213, N891, N240);
nand NAND4 (N957, N949, N285, N846, N153);
xor XOR2 (N958, N956, N907);
and AND4 (N959, N957, N559, N610, N744);
or OR4 (N960, N937, N881, N37, N283);
or OR4 (N961, N946, N932, N648, N450);
buf BUF1 (N962, N958);
nor NOR3 (N963, N961, N418, N615);
nor NOR4 (N964, N942, N144, N772, N42);
xor XOR2 (N965, N962, N656);
or OR2 (N966, N964, N749);
nor NOR4 (N967, N950, N806, N402, N59);
or OR4 (N968, N953, N668, N43, N66);
or OR2 (N969, N965, N821);
buf BUF1 (N970, N940);
nor NOR2 (N971, N963, N71);
nand NAND4 (N972, N966, N944, N407, N545);
and AND3 (N973, N967, N731, N761);
nand NAND3 (N974, N969, N634, N429);
nand NAND4 (N975, N972, N953, N133, N288);
buf BUF1 (N976, N955);
not NOT1 (N977, N960);
or OR4 (N978, N968, N372, N567, N888);
and AND4 (N979, N971, N233, N654, N547);
not NOT1 (N980, N979);
nor NOR4 (N981, N974, N772, N387, N36);
nand NAND2 (N982, N973, N661);
nor NOR2 (N983, N980, N542);
xor XOR2 (N984, N977, N520);
nor NOR3 (N985, N975, N136, N383);
not NOT1 (N986, N976);
xor XOR2 (N987, N983, N505);
nand NAND3 (N988, N981, N202, N469);
nor NOR4 (N989, N988, N474, N974, N644);
nand NAND3 (N990, N970, N154, N417);
or OR4 (N991, N959, N396, N842, N785);
xor XOR2 (N992, N986, N468);
or OR2 (N993, N984, N351);
buf BUF1 (N994, N993);
not NOT1 (N995, N992);
not NOT1 (N996, N989);
xor XOR2 (N997, N996, N921);
nand NAND2 (N998, N995, N550);
nand NAND2 (N999, N985, N282);
nor NOR3 (N1000, N997, N959, N110);
and AND4 (N1001, N987, N401, N64, N301);
and AND3 (N1002, N994, N992, N751);
or OR4 (N1003, N998, N149, N923, N792);
nor NOR2 (N1004, N999, N414);
nand NAND4 (N1005, N990, N96, N705, N168);
or OR2 (N1006, N982, N434);
and AND2 (N1007, N1004, N365);
not NOT1 (N1008, N978);
not NOT1 (N1009, N1008);
xor XOR2 (N1010, N1000, N22);
xor XOR2 (N1011, N1003, N44);
buf BUF1 (N1012, N1001);
nand NAND3 (N1013, N991, N511, N180);
nand NAND3 (N1014, N1011, N802, N110);
nand NAND3 (N1015, N1013, N525, N170);
not NOT1 (N1016, N1014);
or OR2 (N1017, N1010, N575);
buf BUF1 (N1018, N941);
buf BUF1 (N1019, N1002);
nand NAND2 (N1020, N1005, N800);
not NOT1 (N1021, N1019);
or OR4 (N1022, N1006, N219, N726, N761);
or OR3 (N1023, N1012, N693, N791);
and AND3 (N1024, N1020, N18, N879);
nor NOR4 (N1025, N1023, N1023, N896, N191);
nand NAND4 (N1026, N1016, N676, N157, N715);
xor XOR2 (N1027, N1018, N700);
nor NOR4 (N1028, N1017, N940, N1027, N807);
not NOT1 (N1029, N848);
not NOT1 (N1030, N1015);
nand NAND3 (N1031, N1028, N400, N352);
not NOT1 (N1032, N1029);
nor NOR2 (N1033, N1009, N488);
or OR2 (N1034, N1030, N705);
buf BUF1 (N1035, N1022);
or OR3 (N1036, N1024, N421, N789);
nand NAND4 (N1037, N1033, N393, N646, N404);
nor NOR2 (N1038, N1034, N990);
nor NOR2 (N1039, N1031, N548);
nand NAND4 (N1040, N1021, N737, N238, N229);
or OR3 (N1041, N1032, N308, N677);
and AND4 (N1042, N1025, N995, N367, N420);
nor NOR3 (N1043, N1042, N893, N393);
or OR3 (N1044, N1038, N57, N977);
nand NAND2 (N1045, N1026, N90);
nand NAND3 (N1046, N1045, N812, N856);
buf BUF1 (N1047, N1043);
and AND2 (N1048, N1040, N1045);
buf BUF1 (N1049, N1044);
nand NAND4 (N1050, N1047, N127, N956, N508);
not NOT1 (N1051, N1039);
nand NAND2 (N1052, N1035, N17);
or OR2 (N1053, N1049, N1028);
not NOT1 (N1054, N1041);
not NOT1 (N1055, N1036);
buf BUF1 (N1056, N1050);
xor XOR2 (N1057, N1053, N202);
or OR2 (N1058, N1037, N392);
and AND4 (N1059, N1054, N575, N560, N403);
or OR3 (N1060, N1051, N55, N800);
and AND4 (N1061, N1057, N749, N672, N546);
or OR4 (N1062, N1059, N675, N858, N208);
buf BUF1 (N1063, N1061);
or OR4 (N1064, N1056, N978, N584, N539);
buf BUF1 (N1065, N1058);
buf BUF1 (N1066, N1064);
nand NAND4 (N1067, N1048, N601, N849, N405);
and AND3 (N1068, N1007, N537, N500);
buf BUF1 (N1069, N1066);
not NOT1 (N1070, N1046);
or OR3 (N1071, N1052, N222, N738);
and AND4 (N1072, N1062, N885, N358, N588);
not NOT1 (N1073, N1070);
nor NOR4 (N1074, N1065, N259, N516, N1002);
buf BUF1 (N1075, N1068);
and AND4 (N1076, N1071, N806, N329, N559);
not NOT1 (N1077, N1072);
or OR4 (N1078, N1060, N601, N215, N946);
not NOT1 (N1079, N1073);
nand NAND4 (N1080, N1074, N434, N567, N379);
and AND2 (N1081, N1055, N806);
not NOT1 (N1082, N1081);
nor NOR2 (N1083, N1076, N1038);
buf BUF1 (N1084, N1078);
or OR2 (N1085, N1082, N916);
xor XOR2 (N1086, N1063, N563);
buf BUF1 (N1087, N1086);
nor NOR4 (N1088, N1075, N148, N1011, N206);
buf BUF1 (N1089, N1084);
nor NOR2 (N1090, N1069, N583);
buf BUF1 (N1091, N1067);
and AND4 (N1092, N1091, N285, N118, N538);
or OR2 (N1093, N1079, N137);
nor NOR4 (N1094, N1087, N1050, N40, N606);
xor XOR2 (N1095, N1089, N239);
buf BUF1 (N1096, N1093);
or OR3 (N1097, N1092, N787, N133);
nor NOR3 (N1098, N1088, N1071, N193);
xor XOR2 (N1099, N1096, N966);
xor XOR2 (N1100, N1099, N991);
nand NAND4 (N1101, N1097, N485, N80, N456);
nand NAND2 (N1102, N1094, N382);
buf BUF1 (N1103, N1080);
nor NOR2 (N1104, N1103, N157);
or OR2 (N1105, N1098, N897);
not NOT1 (N1106, N1083);
or OR3 (N1107, N1090, N183, N918);
nor NOR3 (N1108, N1104, N389, N220);
nor NOR4 (N1109, N1106, N25, N773, N459);
buf BUF1 (N1110, N1077);
nand NAND4 (N1111, N1107, N881, N854, N540);
buf BUF1 (N1112, N1108);
nor NOR3 (N1113, N1085, N931, N1029);
not NOT1 (N1114, N1109);
xor XOR2 (N1115, N1111, N307);
xor XOR2 (N1116, N1095, N423);
buf BUF1 (N1117, N1110);
nand NAND2 (N1118, N1101, N1052);
xor XOR2 (N1119, N1116, N687);
or OR3 (N1120, N1102, N352, N814);
not NOT1 (N1121, N1120);
buf BUF1 (N1122, N1114);
nand NAND3 (N1123, N1122, N885, N502);
nor NOR2 (N1124, N1123, N845);
nor NOR2 (N1125, N1117, N465);
buf BUF1 (N1126, N1125);
buf BUF1 (N1127, N1126);
or OR3 (N1128, N1113, N28, N168);
nand NAND3 (N1129, N1128, N1022, N735);
not NOT1 (N1130, N1121);
nand NAND4 (N1131, N1130, N1022, N426, N363);
nand NAND3 (N1132, N1100, N781, N272);
not NOT1 (N1133, N1119);
and AND4 (N1134, N1133, N395, N991, N1045);
and AND4 (N1135, N1129, N951, N310, N674);
nand NAND3 (N1136, N1112, N617, N807);
nor NOR4 (N1137, N1135, N880, N809, N304);
nor NOR2 (N1138, N1131, N396);
buf BUF1 (N1139, N1137);
or OR3 (N1140, N1134, N310, N434);
nor NOR2 (N1141, N1127, N8);
buf BUF1 (N1142, N1139);
buf BUF1 (N1143, N1124);
nor NOR3 (N1144, N1105, N248, N49);
buf BUF1 (N1145, N1136);
and AND4 (N1146, N1115, N788, N954, N1102);
buf BUF1 (N1147, N1143);
nor NOR4 (N1148, N1140, N798, N391, N884);
not NOT1 (N1149, N1138);
nor NOR4 (N1150, N1148, N61, N579, N18);
buf BUF1 (N1151, N1150);
and AND4 (N1152, N1149, N811, N742, N263);
and AND2 (N1153, N1118, N386);
or OR2 (N1154, N1151, N1014);
not NOT1 (N1155, N1154);
not NOT1 (N1156, N1146);
not NOT1 (N1157, N1145);
or OR3 (N1158, N1156, N1109, N185);
buf BUF1 (N1159, N1158);
buf BUF1 (N1160, N1159);
not NOT1 (N1161, N1160);
not NOT1 (N1162, N1141);
buf BUF1 (N1163, N1152);
nand NAND3 (N1164, N1155, N272, N219);
or OR3 (N1165, N1164, N112, N1138);
not NOT1 (N1166, N1144);
nand NAND2 (N1167, N1157, N343);
or OR3 (N1168, N1132, N601, N1109);
nand NAND3 (N1169, N1147, N941, N674);
or OR3 (N1170, N1168, N969, N368);
nor NOR3 (N1171, N1166, N616, N914);
nand NAND2 (N1172, N1167, N680);
nand NAND3 (N1173, N1165, N1134, N713);
buf BUF1 (N1174, N1162);
not NOT1 (N1175, N1153);
not NOT1 (N1176, N1170);
nand NAND3 (N1177, N1176, N971, N360);
buf BUF1 (N1178, N1174);
or OR3 (N1179, N1175, N134, N1044);
nand NAND2 (N1180, N1171, N675);
nor NOR2 (N1181, N1178, N1044);
and AND4 (N1182, N1179, N666, N830, N954);
buf BUF1 (N1183, N1172);
or OR3 (N1184, N1142, N562, N948);
and AND2 (N1185, N1181, N52);
or OR3 (N1186, N1184, N872, N430);
buf BUF1 (N1187, N1185);
buf BUF1 (N1188, N1161);
buf BUF1 (N1189, N1188);
buf BUF1 (N1190, N1180);
buf BUF1 (N1191, N1186);
not NOT1 (N1192, N1189);
not NOT1 (N1193, N1182);
xor XOR2 (N1194, N1192, N1022);
xor XOR2 (N1195, N1173, N604);
buf BUF1 (N1196, N1183);
or OR4 (N1197, N1187, N1007, N287, N408);
xor XOR2 (N1198, N1197, N389);
not NOT1 (N1199, N1177);
nand NAND3 (N1200, N1193, N1018, N858);
nor NOR3 (N1201, N1195, N747, N434);
or OR2 (N1202, N1163, N332);
and AND2 (N1203, N1194, N1166);
buf BUF1 (N1204, N1190);
nor NOR3 (N1205, N1198, N89, N809);
or OR3 (N1206, N1201, N528, N774);
xor XOR2 (N1207, N1199, N512);
and AND3 (N1208, N1204, N781, N127);
xor XOR2 (N1209, N1207, N523);
xor XOR2 (N1210, N1203, N708);
nand NAND4 (N1211, N1209, N745, N381, N978);
and AND2 (N1212, N1169, N182);
not NOT1 (N1213, N1211);
buf BUF1 (N1214, N1213);
nand NAND4 (N1215, N1214, N25, N4, N549);
xor XOR2 (N1216, N1212, N357);
buf BUF1 (N1217, N1216);
not NOT1 (N1218, N1215);
nor NOR4 (N1219, N1205, N521, N1139, N832);
nor NOR3 (N1220, N1210, N256, N339);
nand NAND3 (N1221, N1220, N800, N415);
not NOT1 (N1222, N1221);
not NOT1 (N1223, N1200);
buf BUF1 (N1224, N1223);
xor XOR2 (N1225, N1206, N589);
nand NAND4 (N1226, N1218, N534, N340, N189);
or OR4 (N1227, N1191, N334, N610, N800);
xor XOR2 (N1228, N1196, N861);
buf BUF1 (N1229, N1226);
nor NOR4 (N1230, N1227, N1126, N684, N356);
nand NAND3 (N1231, N1208, N1073, N508);
or OR2 (N1232, N1230, N801);
buf BUF1 (N1233, N1232);
nor NOR4 (N1234, N1219, N1038, N1211, N287);
and AND2 (N1235, N1233, N316);
not NOT1 (N1236, N1234);
nand NAND4 (N1237, N1222, N539, N543, N422);
buf BUF1 (N1238, N1202);
or OR4 (N1239, N1229, N592, N228, N762);
nand NAND2 (N1240, N1231, N19);
buf BUF1 (N1241, N1224);
or OR2 (N1242, N1239, N841);
buf BUF1 (N1243, N1236);
buf BUF1 (N1244, N1237);
buf BUF1 (N1245, N1243);
or OR4 (N1246, N1240, N887, N518, N67);
nor NOR2 (N1247, N1225, N844);
nor NOR3 (N1248, N1244, N643, N88);
or OR4 (N1249, N1245, N399, N113, N940);
not NOT1 (N1250, N1247);
nor NOR4 (N1251, N1249, N758, N1045, N1069);
not NOT1 (N1252, N1217);
nand NAND2 (N1253, N1238, N878);
nor NOR2 (N1254, N1251, N192);
buf BUF1 (N1255, N1241);
buf BUF1 (N1256, N1254);
nand NAND4 (N1257, N1252, N788, N755, N910);
buf BUF1 (N1258, N1228);
nand NAND2 (N1259, N1253, N790);
nand NAND2 (N1260, N1246, N43);
xor XOR2 (N1261, N1235, N1234);
nor NOR3 (N1262, N1257, N1200, N216);
and AND2 (N1263, N1248, N1243);
or OR4 (N1264, N1250, N538, N1218, N1100);
nand NAND2 (N1265, N1261, N969);
buf BUF1 (N1266, N1263);
xor XOR2 (N1267, N1262, N470);
buf BUF1 (N1268, N1256);
xor XOR2 (N1269, N1259, N272);
or OR2 (N1270, N1258, N792);
nor NOR3 (N1271, N1266, N478, N895);
nand NAND2 (N1272, N1268, N133);
or OR2 (N1273, N1242, N1204);
nand NAND3 (N1274, N1255, N80, N526);
xor XOR2 (N1275, N1272, N285);
buf BUF1 (N1276, N1269);
or OR4 (N1277, N1273, N1068, N884, N766);
buf BUF1 (N1278, N1264);
buf BUF1 (N1279, N1267);
and AND2 (N1280, N1276, N788);
not NOT1 (N1281, N1278);
and AND3 (N1282, N1274, N242, N188);
nor NOR4 (N1283, N1281, N154, N427, N1260);
and AND3 (N1284, N583, N893, N370);
buf BUF1 (N1285, N1275);
nand NAND4 (N1286, N1277, N972, N257, N975);
or OR2 (N1287, N1270, N871);
xor XOR2 (N1288, N1282, N90);
xor XOR2 (N1289, N1279, N688);
and AND3 (N1290, N1284, N917, N1075);
or OR2 (N1291, N1289, N732);
not NOT1 (N1292, N1291);
xor XOR2 (N1293, N1290, N339);
and AND3 (N1294, N1286, N143, N639);
not NOT1 (N1295, N1265);
not NOT1 (N1296, N1292);
or OR4 (N1297, N1271, N697, N494, N1031);
xor XOR2 (N1298, N1283, N131);
xor XOR2 (N1299, N1296, N1020);
xor XOR2 (N1300, N1298, N649);
nor NOR4 (N1301, N1293, N780, N526, N1282);
buf BUF1 (N1302, N1294);
nand NAND4 (N1303, N1299, N1251, N898, N920);
or OR3 (N1304, N1302, N242, N340);
buf BUF1 (N1305, N1301);
and AND3 (N1306, N1285, N395, N34);
or OR4 (N1307, N1305, N115, N624, N371);
xor XOR2 (N1308, N1297, N1091);
nand NAND3 (N1309, N1300, N391, N390);
buf BUF1 (N1310, N1307);
not NOT1 (N1311, N1306);
nor NOR3 (N1312, N1280, N1050, N1306);
nor NOR2 (N1313, N1304, N888);
not NOT1 (N1314, N1303);
not NOT1 (N1315, N1311);
or OR3 (N1316, N1309, N1023, N421);
buf BUF1 (N1317, N1287);
not NOT1 (N1318, N1312);
not NOT1 (N1319, N1313);
nor NOR4 (N1320, N1315, N1315, N294, N1297);
not NOT1 (N1321, N1314);
xor XOR2 (N1322, N1308, N1210);
not NOT1 (N1323, N1318);
xor XOR2 (N1324, N1295, N979);
or OR3 (N1325, N1323, N764, N338);
nor NOR2 (N1326, N1310, N88);
and AND4 (N1327, N1319, N636, N508, N1002);
nor NOR2 (N1328, N1288, N220);
nand NAND3 (N1329, N1320, N67, N604);
and AND4 (N1330, N1329, N301, N873, N765);
nor NOR3 (N1331, N1321, N1122, N980);
buf BUF1 (N1332, N1331);
nand NAND3 (N1333, N1324, N1305, N673);
xor XOR2 (N1334, N1333, N530);
nor NOR2 (N1335, N1316, N603);
or OR3 (N1336, N1335, N879, N81);
buf BUF1 (N1337, N1327);
nand NAND3 (N1338, N1317, N1261, N1264);
and AND4 (N1339, N1332, N937, N430, N485);
nand NAND2 (N1340, N1325, N1142);
or OR2 (N1341, N1338, N551);
nand NAND3 (N1342, N1337, N1235, N1293);
nand NAND3 (N1343, N1326, N648, N1067);
not NOT1 (N1344, N1339);
nand NAND2 (N1345, N1342, N262);
nand NAND2 (N1346, N1336, N1148);
and AND4 (N1347, N1344, N54, N226, N168);
nand NAND3 (N1348, N1347, N1309, N219);
nor NOR3 (N1349, N1346, N1248, N567);
or OR4 (N1350, N1334, N97, N720, N807);
xor XOR2 (N1351, N1341, N1315);
xor XOR2 (N1352, N1343, N1);
or OR3 (N1353, N1350, N1121, N183);
xor XOR2 (N1354, N1330, N575);
not NOT1 (N1355, N1351);
xor XOR2 (N1356, N1352, N621);
buf BUF1 (N1357, N1355);
and AND3 (N1358, N1345, N137, N1281);
buf BUF1 (N1359, N1349);
nor NOR2 (N1360, N1322, N295);
buf BUF1 (N1361, N1328);
nand NAND4 (N1362, N1361, N724, N324, N996);
xor XOR2 (N1363, N1354, N316);
nand NAND2 (N1364, N1362, N1094);
nand NAND3 (N1365, N1360, N854, N178);
and AND4 (N1366, N1365, N1226, N1156, N1316);
buf BUF1 (N1367, N1353);
nand NAND2 (N1368, N1357, N719);
buf BUF1 (N1369, N1368);
not NOT1 (N1370, N1369);
xor XOR2 (N1371, N1358, N157);
not NOT1 (N1372, N1371);
nor NOR3 (N1373, N1348, N417, N1276);
or OR3 (N1374, N1359, N278, N687);
buf BUF1 (N1375, N1366);
not NOT1 (N1376, N1375);
nor NOR3 (N1377, N1376, N301, N58);
not NOT1 (N1378, N1373);
xor XOR2 (N1379, N1377, N134);
and AND4 (N1380, N1363, N633, N652, N1022);
or OR3 (N1381, N1340, N183, N1069);
buf BUF1 (N1382, N1381);
not NOT1 (N1383, N1374);
or OR3 (N1384, N1379, N269, N961);
not NOT1 (N1385, N1356);
nor NOR3 (N1386, N1367, N867, N955);
not NOT1 (N1387, N1378);
xor XOR2 (N1388, N1382, N1172);
nor NOR2 (N1389, N1383, N118);
buf BUF1 (N1390, N1389);
or OR4 (N1391, N1370, N749, N533, N306);
nor NOR3 (N1392, N1391, N828, N1363);
not NOT1 (N1393, N1384);
nand NAND3 (N1394, N1392, N78, N1092);
or OR4 (N1395, N1380, N122, N682, N1143);
not NOT1 (N1396, N1372);
or OR4 (N1397, N1390, N107, N468, N1321);
nor NOR4 (N1398, N1396, N1198, N751, N1256);
buf BUF1 (N1399, N1394);
or OR4 (N1400, N1395, N1056, N884, N16);
buf BUF1 (N1401, N1397);
and AND2 (N1402, N1399, N312);
buf BUF1 (N1403, N1387);
xor XOR2 (N1404, N1401, N54);
xor XOR2 (N1405, N1403, N653);
not NOT1 (N1406, N1364);
nand NAND3 (N1407, N1405, N1333, N467);
nor NOR2 (N1408, N1400, N760);
not NOT1 (N1409, N1385);
buf BUF1 (N1410, N1386);
nor NOR4 (N1411, N1410, N207, N158, N542);
buf BUF1 (N1412, N1406);
nor NOR2 (N1413, N1388, N801);
buf BUF1 (N1414, N1413);
not NOT1 (N1415, N1408);
xor XOR2 (N1416, N1411, N620);
nor NOR4 (N1417, N1404, N1364, N318, N1009);
or OR2 (N1418, N1417, N2);
buf BUF1 (N1419, N1412);
nand NAND2 (N1420, N1419, N509);
and AND3 (N1421, N1402, N1402, N1409);
xor XOR2 (N1422, N329, N83);
buf BUF1 (N1423, N1393);
and AND3 (N1424, N1423, N368, N176);
xor XOR2 (N1425, N1422, N1177);
nand NAND3 (N1426, N1421, N58, N822);
buf BUF1 (N1427, N1420);
xor XOR2 (N1428, N1427, N1129);
not NOT1 (N1429, N1428);
buf BUF1 (N1430, N1415);
or OR2 (N1431, N1426, N301);
nor NOR4 (N1432, N1429, N1083, N724, N398);
buf BUF1 (N1433, N1416);
or OR4 (N1434, N1424, N240, N271, N199);
buf BUF1 (N1435, N1425);
not NOT1 (N1436, N1432);
nor NOR4 (N1437, N1430, N94, N451, N964);
or OR2 (N1438, N1434, N1094);
not NOT1 (N1439, N1414);
and AND4 (N1440, N1435, N138, N812, N49);
nor NOR3 (N1441, N1431, N118, N921);
and AND3 (N1442, N1441, N753, N484);
buf BUF1 (N1443, N1439);
and AND4 (N1444, N1443, N841, N597, N142);
and AND4 (N1445, N1407, N992, N578, N637);
not NOT1 (N1446, N1437);
and AND2 (N1447, N1398, N189);
nand NAND3 (N1448, N1440, N1407, N236);
xor XOR2 (N1449, N1446, N587);
xor XOR2 (N1450, N1433, N138);
nand NAND4 (N1451, N1447, N875, N1174, N356);
and AND2 (N1452, N1444, N57);
not NOT1 (N1453, N1448);
or OR3 (N1454, N1442, N56, N1255);
and AND4 (N1455, N1454, N1115, N520, N1018);
not NOT1 (N1456, N1453);
xor XOR2 (N1457, N1455, N943);
xor XOR2 (N1458, N1449, N1291);
and AND3 (N1459, N1418, N467, N696);
nor NOR3 (N1460, N1458, N319, N581);
nand NAND2 (N1461, N1452, N361);
nand NAND3 (N1462, N1459, N1314, N607);
or OR4 (N1463, N1460, N846, N866, N1145);
not NOT1 (N1464, N1461);
and AND2 (N1465, N1451, N61);
nor NOR3 (N1466, N1436, N1168, N1136);
xor XOR2 (N1467, N1464, N300);
not NOT1 (N1468, N1450);
nand NAND4 (N1469, N1468, N507, N851, N1052);
nand NAND3 (N1470, N1465, N1289, N247);
not NOT1 (N1471, N1466);
xor XOR2 (N1472, N1470, N405);
and AND2 (N1473, N1438, N112);
or OR2 (N1474, N1457, N527);
xor XOR2 (N1475, N1456, N697);
nor NOR2 (N1476, N1471, N352);
and AND3 (N1477, N1463, N164, N1414);
or OR2 (N1478, N1462, N1366);
buf BUF1 (N1479, N1475);
or OR4 (N1480, N1476, N242, N1204, N14);
and AND4 (N1481, N1472, N129, N380, N1085);
nor NOR4 (N1482, N1445, N893, N655, N1194);
not NOT1 (N1483, N1482);
not NOT1 (N1484, N1477);
nand NAND3 (N1485, N1483, N1097, N1232);
and AND2 (N1486, N1478, N1073);
buf BUF1 (N1487, N1486);
and AND4 (N1488, N1484, N810, N1115, N229);
and AND4 (N1489, N1481, N747, N549, N502);
buf BUF1 (N1490, N1485);
xor XOR2 (N1491, N1488, N233);
nand NAND4 (N1492, N1474, N430, N261, N740);
and AND3 (N1493, N1487, N321, N195);
xor XOR2 (N1494, N1473, N430);
nor NOR4 (N1495, N1467, N494, N133, N793);
or OR2 (N1496, N1492, N1270);
not NOT1 (N1497, N1480);
xor XOR2 (N1498, N1469, N1053);
nand NAND2 (N1499, N1493, N417);
and AND3 (N1500, N1496, N380, N911);
not NOT1 (N1501, N1497);
nand NAND3 (N1502, N1490, N506, N1098);
or OR4 (N1503, N1502, N72, N1148, N108);
xor XOR2 (N1504, N1498, N379);
nand NAND4 (N1505, N1504, N680, N600, N1440);
and AND3 (N1506, N1499, N292, N297);
xor XOR2 (N1507, N1505, N1483);
or OR3 (N1508, N1495, N1016, N1469);
nand NAND4 (N1509, N1500, N867, N422, N285);
xor XOR2 (N1510, N1506, N1016);
xor XOR2 (N1511, N1494, N1039);
nor NOR3 (N1512, N1479, N854, N784);
nor NOR3 (N1513, N1503, N375, N1169);
and AND3 (N1514, N1511, N529, N787);
nor NOR2 (N1515, N1514, N647);
not NOT1 (N1516, N1513);
buf BUF1 (N1517, N1501);
xor XOR2 (N1518, N1491, N1116);
not NOT1 (N1519, N1512);
or OR3 (N1520, N1517, N476, N849);
buf BUF1 (N1521, N1518);
nand NAND4 (N1522, N1508, N584, N51, N100);
or OR4 (N1523, N1516, N974, N1515, N1456);
or OR2 (N1524, N936, N891);
and AND2 (N1525, N1509, N1307);
nand NAND4 (N1526, N1522, N377, N1237, N1040);
nand NAND2 (N1527, N1489, N287);
not NOT1 (N1528, N1526);
nand NAND3 (N1529, N1527, N556, N57);
not NOT1 (N1530, N1528);
not NOT1 (N1531, N1524);
xor XOR2 (N1532, N1521, N111);
and AND2 (N1533, N1519, N775);
not NOT1 (N1534, N1520);
nor NOR2 (N1535, N1507, N726);
not NOT1 (N1536, N1532);
or OR4 (N1537, N1523, N1294, N801, N1029);
not NOT1 (N1538, N1533);
xor XOR2 (N1539, N1538, N353);
nand NAND3 (N1540, N1529, N881, N601);
not NOT1 (N1541, N1525);
nor NOR2 (N1542, N1541, N49);
nand NAND3 (N1543, N1542, N1509, N1318);
nor NOR3 (N1544, N1543, N396, N1453);
and AND2 (N1545, N1531, N973);
not NOT1 (N1546, N1537);
xor XOR2 (N1547, N1544, N1211);
xor XOR2 (N1548, N1540, N929);
xor XOR2 (N1549, N1510, N1220);
and AND4 (N1550, N1546, N471, N1249, N563);
and AND2 (N1551, N1535, N356);
xor XOR2 (N1552, N1548, N280);
and AND4 (N1553, N1534, N738, N1438, N335);
or OR2 (N1554, N1550, N1183);
buf BUF1 (N1555, N1530);
and AND3 (N1556, N1539, N970, N393);
buf BUF1 (N1557, N1536);
nor NOR3 (N1558, N1549, N1101, N880);
nand NAND2 (N1559, N1555, N69);
nor NOR4 (N1560, N1557, N1071, N879, N267);
not NOT1 (N1561, N1551);
and AND2 (N1562, N1561, N674);
or OR2 (N1563, N1560, N18);
not NOT1 (N1564, N1553);
or OR3 (N1565, N1552, N511, N586);
buf BUF1 (N1566, N1545);
buf BUF1 (N1567, N1556);
buf BUF1 (N1568, N1565);
and AND4 (N1569, N1562, N512, N237, N1521);
buf BUF1 (N1570, N1554);
not NOT1 (N1571, N1567);
nor NOR3 (N1572, N1566, N939, N1130);
nand NAND2 (N1573, N1571, N771);
nor NOR2 (N1574, N1572, N982);
or OR2 (N1575, N1569, N1518);
nor NOR2 (N1576, N1558, N1005);
buf BUF1 (N1577, N1570);
or OR3 (N1578, N1563, N619, N693);
or OR2 (N1579, N1578, N480);
and AND4 (N1580, N1547, N294, N776, N1203);
or OR3 (N1581, N1575, N346, N666);
not NOT1 (N1582, N1568);
or OR2 (N1583, N1564, N547);
buf BUF1 (N1584, N1583);
nand NAND2 (N1585, N1577, N148);
nand NAND3 (N1586, N1582, N911, N1238);
nor NOR4 (N1587, N1574, N1179, N1171, N1563);
xor XOR2 (N1588, N1573, N782);
not NOT1 (N1589, N1585);
not NOT1 (N1590, N1576);
nor NOR3 (N1591, N1586, N1419, N9);
nor NOR2 (N1592, N1590, N57);
nor NOR4 (N1593, N1592, N376, N1027, N195);
xor XOR2 (N1594, N1591, N155);
not NOT1 (N1595, N1584);
or OR2 (N1596, N1559, N662);
xor XOR2 (N1597, N1579, N1287);
and AND3 (N1598, N1588, N846, N75);
or OR4 (N1599, N1597, N691, N940, N1137);
nand NAND4 (N1600, N1580, N204, N1444, N186);
buf BUF1 (N1601, N1594);
buf BUF1 (N1602, N1599);
not NOT1 (N1603, N1595);
xor XOR2 (N1604, N1601, N262);
not NOT1 (N1605, N1600);
and AND3 (N1606, N1598, N1355, N475);
buf BUF1 (N1607, N1581);
and AND4 (N1608, N1593, N651, N1243, N175);
buf BUF1 (N1609, N1589);
and AND2 (N1610, N1587, N997);
and AND2 (N1611, N1603, N1075);
or OR4 (N1612, N1606, N1357, N381, N1198);
or OR2 (N1613, N1608, N1219);
not NOT1 (N1614, N1612);
xor XOR2 (N1615, N1602, N1245);
or OR2 (N1616, N1610, N132);
nor NOR2 (N1617, N1616, N433);
nand NAND3 (N1618, N1617, N1172, N1320);
not NOT1 (N1619, N1614);
nor NOR2 (N1620, N1605, N1539);
and AND3 (N1621, N1620, N419, N232);
nor NOR2 (N1622, N1619, N407);
nand NAND2 (N1623, N1618, N388);
and AND3 (N1624, N1613, N1345, N405);
or OR2 (N1625, N1623, N1488);
and AND2 (N1626, N1609, N456);
and AND4 (N1627, N1622, N1334, N1267, N1080);
nand NAND2 (N1628, N1607, N521);
not NOT1 (N1629, N1627);
and AND4 (N1630, N1626, N441, N318, N489);
nor NOR4 (N1631, N1628, N698, N1380, N1518);
not NOT1 (N1632, N1625);
xor XOR2 (N1633, N1611, N303);
and AND2 (N1634, N1624, N42);
nor NOR2 (N1635, N1631, N392);
buf BUF1 (N1636, N1621);
xor XOR2 (N1637, N1604, N716);
nor NOR4 (N1638, N1596, N1080, N1222, N737);
nand NAND3 (N1639, N1629, N827, N976);
xor XOR2 (N1640, N1615, N105);
nand NAND2 (N1641, N1632, N1548);
and AND3 (N1642, N1641, N480, N468);
xor XOR2 (N1643, N1633, N352);
or OR2 (N1644, N1637, N485);
buf BUF1 (N1645, N1635);
nand NAND2 (N1646, N1642, N1466);
not NOT1 (N1647, N1634);
nor NOR3 (N1648, N1646, N676, N643);
or OR2 (N1649, N1644, N1246);
xor XOR2 (N1650, N1630, N34);
xor XOR2 (N1651, N1636, N977);
and AND2 (N1652, N1638, N1254);
nor NOR2 (N1653, N1643, N625);
nor NOR2 (N1654, N1647, N1594);
and AND3 (N1655, N1640, N471, N511);
or OR4 (N1656, N1655, N236, N42, N1043);
and AND2 (N1657, N1654, N1399);
buf BUF1 (N1658, N1656);
buf BUF1 (N1659, N1648);
xor XOR2 (N1660, N1652, N1565);
xor XOR2 (N1661, N1645, N130);
or OR4 (N1662, N1650, N239, N38, N1124);
or OR2 (N1663, N1649, N604);
buf BUF1 (N1664, N1661);
not NOT1 (N1665, N1662);
nor NOR3 (N1666, N1660, N995, N1253);
nand NAND3 (N1667, N1658, N303, N986);
not NOT1 (N1668, N1639);
xor XOR2 (N1669, N1659, N34);
nand NAND4 (N1670, N1657, N1272, N1446, N1041);
not NOT1 (N1671, N1667);
or OR4 (N1672, N1664, N554, N1036, N1133);
nor NOR2 (N1673, N1666, N1011);
buf BUF1 (N1674, N1651);
or OR2 (N1675, N1672, N1063);
nand NAND4 (N1676, N1675, N76, N94, N1155);
nor NOR4 (N1677, N1668, N1418, N789, N37);
or OR2 (N1678, N1674, N385);
nor NOR4 (N1679, N1678, N132, N449, N756);
buf BUF1 (N1680, N1670);
nor NOR2 (N1681, N1671, N1209);
or OR4 (N1682, N1665, N1498, N1300, N411);
nand NAND3 (N1683, N1682, N1193, N328);
nor NOR3 (N1684, N1676, N1302, N476);
buf BUF1 (N1685, N1683);
and AND2 (N1686, N1680, N141);
buf BUF1 (N1687, N1677);
and AND3 (N1688, N1653, N711, N914);
nand NAND2 (N1689, N1681, N1556);
nor NOR3 (N1690, N1669, N716, N1166);
and AND3 (N1691, N1689, N585, N1064);
and AND2 (N1692, N1673, N1506);
not NOT1 (N1693, N1679);
or OR2 (N1694, N1693, N330);
nor NOR2 (N1695, N1687, N1167);
xor XOR2 (N1696, N1686, N1637);
and AND3 (N1697, N1691, N905, N352);
nand NAND3 (N1698, N1694, N56, N1302);
nor NOR3 (N1699, N1697, N955, N763);
buf BUF1 (N1700, N1685);
nor NOR2 (N1701, N1699, N474);
or OR3 (N1702, N1690, N1193, N1173);
or OR3 (N1703, N1696, N519, N1346);
nand NAND3 (N1704, N1701, N346, N1406);
and AND3 (N1705, N1684, N617, N435);
nand NAND2 (N1706, N1663, N1536);
xor XOR2 (N1707, N1688, N644);
or OR2 (N1708, N1698, N1697);
and AND3 (N1709, N1702, N793, N1512);
nand NAND4 (N1710, N1692, N1230, N1530, N954);
xor XOR2 (N1711, N1703, N631);
nand NAND2 (N1712, N1704, N1579);
or OR2 (N1713, N1707, N970);
or OR4 (N1714, N1708, N606, N940, N768);
nor NOR3 (N1715, N1709, N168, N1227);
and AND2 (N1716, N1713, N653);
buf BUF1 (N1717, N1706);
or OR3 (N1718, N1716, N149, N1248);
and AND4 (N1719, N1715, N361, N115, N1544);
nand NAND2 (N1720, N1714, N1685);
or OR3 (N1721, N1712, N1113, N325);
nand NAND2 (N1722, N1695, N1357);
buf BUF1 (N1723, N1717);
nor NOR4 (N1724, N1721, N1091, N424, N1247);
not NOT1 (N1725, N1700);
xor XOR2 (N1726, N1720, N1135);
or OR2 (N1727, N1726, N780);
nor NOR2 (N1728, N1711, N1519);
nor NOR4 (N1729, N1710, N277, N972, N552);
nor NOR2 (N1730, N1729, N1492);
xor XOR2 (N1731, N1728, N100);
nor NOR4 (N1732, N1725, N16, N1706, N1456);
xor XOR2 (N1733, N1724, N1414);
and AND2 (N1734, N1730, N742);
nand NAND2 (N1735, N1734, N50);
nand NAND2 (N1736, N1723, N1045);
nand NAND3 (N1737, N1705, N44, N1142);
buf BUF1 (N1738, N1736);
buf BUF1 (N1739, N1718);
nand NAND3 (N1740, N1738, N686, N1690);
buf BUF1 (N1741, N1737);
and AND2 (N1742, N1727, N1282);
and AND3 (N1743, N1722, N355, N926);
nor NOR4 (N1744, N1731, N635, N1352, N830);
nor NOR3 (N1745, N1719, N412, N706);
nand NAND2 (N1746, N1743, N867);
xor XOR2 (N1747, N1742, N940);
or OR2 (N1748, N1745, N1489);
xor XOR2 (N1749, N1746, N1293);
nor NOR2 (N1750, N1735, N471);
not NOT1 (N1751, N1750);
not NOT1 (N1752, N1732);
nor NOR3 (N1753, N1747, N436, N597);
not NOT1 (N1754, N1749);
xor XOR2 (N1755, N1741, N670);
nand NAND4 (N1756, N1751, N468, N998, N1041);
or OR4 (N1757, N1739, N1416, N924, N118);
nand NAND3 (N1758, N1756, N1728, N1179);
and AND4 (N1759, N1755, N912, N236, N1407);
nand NAND3 (N1760, N1752, N1341, N932);
and AND3 (N1761, N1740, N1573, N1392);
not NOT1 (N1762, N1761);
nor NOR3 (N1763, N1757, N111, N820);
nand NAND4 (N1764, N1762, N1109, N840, N352);
or OR4 (N1765, N1754, N375, N1532, N103);
or OR2 (N1766, N1759, N1095);
and AND3 (N1767, N1760, N661, N161);
nand NAND4 (N1768, N1763, N193, N1276, N850);
nand NAND2 (N1769, N1758, N317);
buf BUF1 (N1770, N1768);
nor NOR4 (N1771, N1766, N140, N1351, N727);
not NOT1 (N1772, N1765);
buf BUF1 (N1773, N1748);
buf BUF1 (N1774, N1773);
xor XOR2 (N1775, N1771, N1043);
xor XOR2 (N1776, N1769, N1145);
buf BUF1 (N1777, N1767);
and AND3 (N1778, N1774, N1199, N995);
or OR3 (N1779, N1777, N251, N504);
and AND3 (N1780, N1753, N1266, N1622);
and AND4 (N1781, N1770, N633, N1204, N957);
xor XOR2 (N1782, N1781, N1474);
buf BUF1 (N1783, N1764);
nand NAND2 (N1784, N1744, N1358);
or OR2 (N1785, N1778, N591);
xor XOR2 (N1786, N1776, N751);
and AND2 (N1787, N1786, N1025);
buf BUF1 (N1788, N1780);
buf BUF1 (N1789, N1733);
nor NOR4 (N1790, N1787, N218, N1343, N1514);
or OR3 (N1791, N1779, N1585, N674);
xor XOR2 (N1792, N1785, N1586);
or OR3 (N1793, N1792, N178, N1058);
nand NAND3 (N1794, N1784, N541, N192);
and AND2 (N1795, N1790, N101);
and AND4 (N1796, N1775, N625, N585, N704);
nor NOR4 (N1797, N1796, N220, N911, N756);
nand NAND3 (N1798, N1772, N5, N850);
xor XOR2 (N1799, N1782, N1786);
or OR4 (N1800, N1797, N1662, N1454, N1565);
and AND3 (N1801, N1783, N343, N897);
nor NOR2 (N1802, N1800, N1655);
xor XOR2 (N1803, N1801, N582);
not NOT1 (N1804, N1793);
xor XOR2 (N1805, N1794, N561);
or OR4 (N1806, N1788, N1313, N934, N1087);
nand NAND3 (N1807, N1799, N928, N135);
buf BUF1 (N1808, N1798);
buf BUF1 (N1809, N1802);
xor XOR2 (N1810, N1791, N67);
and AND4 (N1811, N1805, N1622, N292, N1443);
not NOT1 (N1812, N1803);
buf BUF1 (N1813, N1804);
buf BUF1 (N1814, N1811);
nand NAND3 (N1815, N1810, N837, N55);
buf BUF1 (N1816, N1789);
nor NOR3 (N1817, N1807, N106, N1540);
not NOT1 (N1818, N1813);
xor XOR2 (N1819, N1806, N1605);
not NOT1 (N1820, N1815);
and AND3 (N1821, N1795, N107, N969);
buf BUF1 (N1822, N1821);
nand NAND2 (N1823, N1809, N160);
xor XOR2 (N1824, N1823, N811);
xor XOR2 (N1825, N1817, N1491);
buf BUF1 (N1826, N1818);
nor NOR4 (N1827, N1816, N1793, N1423, N616);
not NOT1 (N1828, N1826);
nor NOR3 (N1829, N1822, N649, N1093);
and AND4 (N1830, N1820, N434, N531, N355);
xor XOR2 (N1831, N1819, N161);
not NOT1 (N1832, N1812);
buf BUF1 (N1833, N1828);
nand NAND3 (N1834, N1829, N1098, N230);
not NOT1 (N1835, N1825);
nand NAND2 (N1836, N1834, N1427);
nand NAND2 (N1837, N1827, N465);
or OR3 (N1838, N1836, N1432, N689);
buf BUF1 (N1839, N1814);
nor NOR4 (N1840, N1833, N437, N871, N1739);
not NOT1 (N1841, N1840);
and AND4 (N1842, N1835, N203, N1084, N544);
nor NOR2 (N1843, N1832, N1683);
buf BUF1 (N1844, N1808);
nand NAND2 (N1845, N1842, N1294);
or OR4 (N1846, N1845, N848, N217, N22);
not NOT1 (N1847, N1831);
not NOT1 (N1848, N1844);
buf BUF1 (N1849, N1824);
xor XOR2 (N1850, N1849, N366);
and AND2 (N1851, N1848, N736);
buf BUF1 (N1852, N1839);
xor XOR2 (N1853, N1838, N533);
xor XOR2 (N1854, N1853, N512);
nand NAND2 (N1855, N1854, N119);
and AND3 (N1856, N1837, N1803, N1164);
xor XOR2 (N1857, N1843, N836);
nor NOR4 (N1858, N1830, N107, N289, N1374);
not NOT1 (N1859, N1855);
nor NOR4 (N1860, N1841, N183, N1676, N871);
and AND4 (N1861, N1847, N840, N103, N769);
nand NAND4 (N1862, N1858, N435, N200, N1329);
buf BUF1 (N1863, N1856);
nor NOR4 (N1864, N1851, N151, N1570, N1236);
and AND3 (N1865, N1846, N1268, N343);
nand NAND4 (N1866, N1865, N1551, N541, N1536);
nand NAND3 (N1867, N1852, N1658, N929);
not NOT1 (N1868, N1850);
not NOT1 (N1869, N1866);
xor XOR2 (N1870, N1863, N178);
not NOT1 (N1871, N1861);
not NOT1 (N1872, N1859);
xor XOR2 (N1873, N1872, N420);
nand NAND3 (N1874, N1862, N181, N900);
nor NOR3 (N1875, N1869, N571, N669);
buf BUF1 (N1876, N1867);
not NOT1 (N1877, N1857);
and AND2 (N1878, N1871, N1359);
or OR2 (N1879, N1876, N263);
not NOT1 (N1880, N1879);
xor XOR2 (N1881, N1868, N38);
buf BUF1 (N1882, N1878);
nor NOR2 (N1883, N1864, N34);
nand NAND3 (N1884, N1883, N1160, N1560);
or OR2 (N1885, N1874, N752);
not NOT1 (N1886, N1881);
xor XOR2 (N1887, N1877, N1166);
nand NAND3 (N1888, N1887, N1612, N48);
nand NAND2 (N1889, N1884, N1729);
xor XOR2 (N1890, N1870, N326);
or OR2 (N1891, N1888, N1461);
or OR2 (N1892, N1860, N459);
or OR3 (N1893, N1875, N1675, N1374);
xor XOR2 (N1894, N1873, N1017);
not NOT1 (N1895, N1890);
not NOT1 (N1896, N1882);
or OR3 (N1897, N1885, N1800, N42);
nor NOR2 (N1898, N1895, N158);
nand NAND2 (N1899, N1896, N304);
xor XOR2 (N1900, N1894, N1452);
nand NAND4 (N1901, N1886, N740, N912, N714);
or OR4 (N1902, N1889, N1176, N597, N1141);
not NOT1 (N1903, N1900);
nor NOR3 (N1904, N1897, N805, N1737);
nand NAND4 (N1905, N1898, N113, N404, N1880);
xor XOR2 (N1906, N775, N1794);
buf BUF1 (N1907, N1902);
not NOT1 (N1908, N1903);
nor NOR3 (N1909, N1891, N1711, N527);
buf BUF1 (N1910, N1893);
buf BUF1 (N1911, N1899);
not NOT1 (N1912, N1910);
buf BUF1 (N1913, N1901);
buf BUF1 (N1914, N1892);
nor NOR4 (N1915, N1908, N304, N1252, N598);
nand NAND4 (N1916, N1914, N1615, N209, N1420);
nand NAND3 (N1917, N1909, N1158, N1693);
buf BUF1 (N1918, N1913);
nor NOR2 (N1919, N1912, N476);
or OR2 (N1920, N1905, N1525);
not NOT1 (N1921, N1917);
buf BUF1 (N1922, N1906);
nand NAND4 (N1923, N1916, N260, N309, N1823);
nand NAND3 (N1924, N1918, N1454, N806);
or OR4 (N1925, N1911, N701, N1793, N771);
nor NOR4 (N1926, N1904, N1741, N322, N40);
nand NAND4 (N1927, N1925, N98, N263, N314);
and AND4 (N1928, N1920, N679, N1164, N1803);
nand NAND3 (N1929, N1928, N43, N533);
and AND4 (N1930, N1907, N689, N1610, N356);
nor NOR4 (N1931, N1924, N1448, N1321, N6);
or OR3 (N1932, N1926, N561, N106);
not NOT1 (N1933, N1929);
xor XOR2 (N1934, N1919, N1243);
not NOT1 (N1935, N1927);
or OR3 (N1936, N1921, N1360, N1077);
nand NAND3 (N1937, N1932, N1091, N115);
buf BUF1 (N1938, N1936);
nand NAND3 (N1939, N1923, N1909, N875);
not NOT1 (N1940, N1922);
buf BUF1 (N1941, N1935);
not NOT1 (N1942, N1938);
xor XOR2 (N1943, N1937, N1334);
nor NOR2 (N1944, N1934, N460);
not NOT1 (N1945, N1940);
not NOT1 (N1946, N1931);
nor NOR2 (N1947, N1941, N600);
nor NOR3 (N1948, N1945, N704, N1528);
nand NAND2 (N1949, N1930, N1171);
and AND3 (N1950, N1946, N1106, N787);
nand NAND2 (N1951, N1948, N1393);
nand NAND2 (N1952, N1939, N305);
and AND4 (N1953, N1951, N350, N1495, N1225);
nor NOR3 (N1954, N1942, N222, N861);
or OR4 (N1955, N1950, N1134, N1047, N250);
or OR3 (N1956, N1947, N1340, N904);
not NOT1 (N1957, N1952);
nand NAND4 (N1958, N1915, N106, N677, N1409);
or OR3 (N1959, N1933, N784, N887);
and AND4 (N1960, N1958, N1584, N835, N1416);
not NOT1 (N1961, N1960);
not NOT1 (N1962, N1943);
buf BUF1 (N1963, N1962);
or OR2 (N1964, N1953, N1206);
nand NAND3 (N1965, N1944, N1813, N1357);
xor XOR2 (N1966, N1965, N426);
and AND3 (N1967, N1963, N199, N984);
not NOT1 (N1968, N1957);
and AND3 (N1969, N1949, N1353, N22);
buf BUF1 (N1970, N1968);
buf BUF1 (N1971, N1954);
or OR4 (N1972, N1961, N1258, N1262, N1044);
nor NOR4 (N1973, N1972, N998, N1404, N553);
nand NAND2 (N1974, N1955, N1609);
or OR4 (N1975, N1974, N910, N500, N1054);
nor NOR2 (N1976, N1970, N928);
buf BUF1 (N1977, N1959);
and AND3 (N1978, N1956, N1367, N1037);
nor NOR4 (N1979, N1971, N847, N1638, N1101);
nand NAND3 (N1980, N1976, N473, N1564);
xor XOR2 (N1981, N1969, N86);
buf BUF1 (N1982, N1973);
and AND2 (N1983, N1964, N523);
buf BUF1 (N1984, N1979);
xor XOR2 (N1985, N1983, N170);
not NOT1 (N1986, N1978);
and AND3 (N1987, N1985, N1779, N12);
nor NOR3 (N1988, N1966, N1387, N762);
xor XOR2 (N1989, N1986, N1226);
buf BUF1 (N1990, N1980);
or OR2 (N1991, N1977, N1675);
xor XOR2 (N1992, N1981, N1148);
nand NAND3 (N1993, N1987, N599, N1534);
nor NOR2 (N1994, N1984, N455);
nand NAND2 (N1995, N1989, N46);
nand NAND2 (N1996, N1967, N1688);
buf BUF1 (N1997, N1992);
nor NOR2 (N1998, N1996, N884);
xor XOR2 (N1999, N1991, N387);
xor XOR2 (N2000, N1998, N1320);
nor NOR2 (N2001, N2000, N1074);
not NOT1 (N2002, N1988);
not NOT1 (N2003, N1999);
xor XOR2 (N2004, N1993, N1425);
not NOT1 (N2005, N2004);
and AND3 (N2006, N1994, N936, N934);
xor XOR2 (N2007, N1990, N1360);
buf BUF1 (N2008, N1982);
nand NAND3 (N2009, N2005, N779, N1254);
nor NOR3 (N2010, N2006, N250, N1483);
not NOT1 (N2011, N2010);
or OR2 (N2012, N2001, N1945);
nand NAND2 (N2013, N1975, N860);
not NOT1 (N2014, N1995);
nand NAND2 (N2015, N2011, N19);
or OR4 (N2016, N2007, N598, N438, N974);
or OR4 (N2017, N2016, N1517, N1106, N1814);
or OR2 (N2018, N2003, N1432);
or OR2 (N2019, N2012, N1061);
buf BUF1 (N2020, N2015);
nor NOR4 (N2021, N2008, N1406, N843, N1461);
not NOT1 (N2022, N2002);
nor NOR3 (N2023, N2017, N240, N160);
nand NAND2 (N2024, N2021, N31);
nand NAND3 (N2025, N2022, N272, N1502);
xor XOR2 (N2026, N2014, N1416);
nand NAND2 (N2027, N2026, N902);
xor XOR2 (N2028, N2018, N206);
and AND4 (N2029, N2028, N1728, N1183, N146);
xor XOR2 (N2030, N2019, N1651);
nor NOR3 (N2031, N2030, N1676, N71);
buf BUF1 (N2032, N2013);
buf BUF1 (N2033, N2024);
nor NOR3 (N2034, N2027, N1074, N1088);
xor XOR2 (N2035, N1997, N1564);
buf BUF1 (N2036, N2034);
nor NOR2 (N2037, N2031, N204);
nor NOR2 (N2038, N2020, N2019);
or OR3 (N2039, N2009, N1142, N86);
and AND2 (N2040, N2039, N2022);
nand NAND2 (N2041, N2035, N580);
nand NAND3 (N2042, N2032, N848, N539);
not NOT1 (N2043, N2040);
nand NAND3 (N2044, N2029, N760, N592);
nor NOR2 (N2045, N2041, N208);
buf BUF1 (N2046, N2033);
nor NOR3 (N2047, N2038, N1836, N292);
buf BUF1 (N2048, N2037);
nor NOR4 (N2049, N2043, N1737, N265, N1896);
not NOT1 (N2050, N2047);
not NOT1 (N2051, N2036);
xor XOR2 (N2052, N2025, N1397);
and AND3 (N2053, N2044, N1386, N1623);
and AND4 (N2054, N2050, N1803, N925, N875);
xor XOR2 (N2055, N2045, N149);
buf BUF1 (N2056, N2046);
nor NOR4 (N2057, N2052, N1896, N708, N1450);
nand NAND2 (N2058, N2057, N1372);
not NOT1 (N2059, N2023);
nand NAND2 (N2060, N2059, N974);
not NOT1 (N2061, N2056);
buf BUF1 (N2062, N2053);
nor NOR2 (N2063, N2058, N1113);
nor NOR4 (N2064, N2042, N1180, N1091, N243);
and AND2 (N2065, N2048, N1467);
or OR3 (N2066, N2062, N167, N1694);
buf BUF1 (N2067, N2061);
nor NOR2 (N2068, N2054, N994);
or OR3 (N2069, N2065, N1422, N637);
nor NOR4 (N2070, N2051, N441, N1255, N32);
xor XOR2 (N2071, N2063, N841);
buf BUF1 (N2072, N2070);
xor XOR2 (N2073, N2060, N1364);
not NOT1 (N2074, N2064);
nor NOR2 (N2075, N2071, N208);
not NOT1 (N2076, N2072);
nor NOR4 (N2077, N2068, N1264, N520, N477);
nor NOR3 (N2078, N2075, N808, N23);
or OR3 (N2079, N2055, N1513, N1966);
nor NOR4 (N2080, N2073, N180, N1800, N29);
and AND4 (N2081, N2067, N47, N1076, N952);
and AND3 (N2082, N2076, N553, N1070);
buf BUF1 (N2083, N2066);
buf BUF1 (N2084, N2081);
buf BUF1 (N2085, N2049);
not NOT1 (N2086, N2069);
nand NAND2 (N2087, N2078, N799);
nand NAND2 (N2088, N2086, N721);
and AND3 (N2089, N2084, N443, N934);
buf BUF1 (N2090, N2087);
xor XOR2 (N2091, N2074, N548);
or OR3 (N2092, N2091, N201, N2049);
nand NAND3 (N2093, N2079, N399, N1616);
xor XOR2 (N2094, N2082, N433);
not NOT1 (N2095, N2080);
or OR3 (N2096, N2092, N1301, N1331);
nor NOR4 (N2097, N2089, N186, N1179, N790);
nand NAND3 (N2098, N2097, N1361, N467);
not NOT1 (N2099, N2093);
xor XOR2 (N2100, N2077, N878);
xor XOR2 (N2101, N2096, N1202);
nor NOR4 (N2102, N2094, N692, N715, N1341);
and AND4 (N2103, N2085, N364, N616, N2058);
nand NAND4 (N2104, N2090, N1751, N2022, N1210);
not NOT1 (N2105, N2102);
nor NOR3 (N2106, N2104, N765, N587);
or OR3 (N2107, N2099, N163, N1340);
nor NOR2 (N2108, N2105, N2054);
not NOT1 (N2109, N2088);
nor NOR3 (N2110, N2100, N1836, N804);
buf BUF1 (N2111, N2107);
nand NAND4 (N2112, N2083, N870, N1039, N2031);
nand NAND3 (N2113, N2110, N290, N1359);
nand NAND3 (N2114, N2103, N1105, N1239);
xor XOR2 (N2115, N2113, N896);
nand NAND4 (N2116, N2112, N503, N1741, N1236);
buf BUF1 (N2117, N2109);
and AND2 (N2118, N2101, N1332);
nor NOR3 (N2119, N2114, N661, N1484);
nor NOR4 (N2120, N2111, N78, N676, N1145);
nor NOR2 (N2121, N2116, N2023);
not NOT1 (N2122, N2118);
or OR4 (N2123, N2115, N953, N307, N1518);
and AND4 (N2124, N2123, N266, N1108, N963);
not NOT1 (N2125, N2121);
buf BUF1 (N2126, N2106);
buf BUF1 (N2127, N2108);
not NOT1 (N2128, N2117);
buf BUF1 (N2129, N2127);
buf BUF1 (N2130, N2120);
or OR2 (N2131, N2119, N1141);
nor NOR4 (N2132, N2129, N1466, N1839, N1117);
buf BUF1 (N2133, N2130);
not NOT1 (N2134, N2128);
and AND3 (N2135, N2122, N1877, N586);
or OR3 (N2136, N2132, N523, N1998);
xor XOR2 (N2137, N2134, N1123);
not NOT1 (N2138, N2137);
nand NAND3 (N2139, N2136, N1300, N1814);
buf BUF1 (N2140, N2139);
xor XOR2 (N2141, N2131, N430);
not NOT1 (N2142, N2098);
nor NOR4 (N2143, N2140, N990, N1441, N1988);
xor XOR2 (N2144, N2133, N1047);
xor XOR2 (N2145, N2138, N1660);
xor XOR2 (N2146, N2145, N519);
or OR3 (N2147, N2124, N904, N2090);
nor NOR3 (N2148, N2126, N2101, N767);
nand NAND2 (N2149, N2141, N1943);
nand NAND4 (N2150, N2146, N1276, N696, N984);
and AND4 (N2151, N2150, N226, N1668, N150);
nand NAND2 (N2152, N2149, N858);
or OR4 (N2153, N2147, N1493, N218, N1819);
not NOT1 (N2154, N2151);
nand NAND2 (N2155, N2144, N1739);
nand NAND3 (N2156, N2143, N1761, N1928);
nand NAND3 (N2157, N2148, N1007, N530);
buf BUF1 (N2158, N2155);
not NOT1 (N2159, N2153);
nor NOR2 (N2160, N2125, N298);
nand NAND4 (N2161, N2159, N1158, N1762, N675);
xor XOR2 (N2162, N2157, N401);
or OR2 (N2163, N2135, N1929);
buf BUF1 (N2164, N2158);
xor XOR2 (N2165, N2095, N992);
nand NAND3 (N2166, N2160, N766, N1138);
nand NAND2 (N2167, N2164, N1474);
or OR3 (N2168, N2152, N1293, N1342);
nand NAND2 (N2169, N2167, N784);
or OR2 (N2170, N2169, N1275);
and AND3 (N2171, N2154, N1161, N39);
nand NAND4 (N2172, N2166, N1760, N305, N1812);
buf BUF1 (N2173, N2165);
xor XOR2 (N2174, N2168, N1045);
nand NAND3 (N2175, N2142, N851, N169);
buf BUF1 (N2176, N2173);
or OR2 (N2177, N2172, N1278);
and AND2 (N2178, N2170, N581);
nand NAND4 (N2179, N2162, N1262, N1812, N480);
buf BUF1 (N2180, N2179);
xor XOR2 (N2181, N2177, N562);
nand NAND4 (N2182, N2171, N1622, N1405, N794);
nand NAND4 (N2183, N2176, N72, N544, N1222);
or OR2 (N2184, N2181, N2008);
not NOT1 (N2185, N2184);
or OR3 (N2186, N2178, N1490, N271);
buf BUF1 (N2187, N2161);
or OR2 (N2188, N2174, N736);
nor NOR2 (N2189, N2188, N848);
and AND2 (N2190, N2182, N1966);
xor XOR2 (N2191, N2180, N1234);
nand NAND2 (N2192, N2156, N2112);
not NOT1 (N2193, N2175);
and AND4 (N2194, N2186, N1892, N461, N256);
or OR3 (N2195, N2193, N166, N1577);
buf BUF1 (N2196, N2163);
or OR3 (N2197, N2195, N1262, N811);
nand NAND3 (N2198, N2197, N1195, N1451);
nor NOR2 (N2199, N2194, N1174);
or OR4 (N2200, N2196, N1686, N1444, N1025);
and AND2 (N2201, N2191, N1658);
xor XOR2 (N2202, N2192, N1460);
nand NAND4 (N2203, N2185, N737, N1795, N1144);
xor XOR2 (N2204, N2190, N905);
or OR2 (N2205, N2187, N908);
or OR4 (N2206, N2199, N874, N808, N705);
and AND4 (N2207, N2202, N176, N2007, N2103);
xor XOR2 (N2208, N2206, N951);
and AND3 (N2209, N2198, N1964, N518);
xor XOR2 (N2210, N2189, N76);
buf BUF1 (N2211, N2205);
nor NOR3 (N2212, N2208, N1790, N1466);
nand NAND3 (N2213, N2204, N1761, N1739);
or OR4 (N2214, N2212, N98, N299, N1381);
nor NOR3 (N2215, N2183, N279, N1677);
or OR3 (N2216, N2215, N1569, N1687);
or OR3 (N2217, N2210, N1012, N1666);
and AND3 (N2218, N2203, N2121, N665);
xor XOR2 (N2219, N2214, N1225);
xor XOR2 (N2220, N2216, N1891);
not NOT1 (N2221, N2217);
and AND4 (N2222, N2213, N2203, N555, N282);
not NOT1 (N2223, N2221);
nor NOR3 (N2224, N2220, N446, N2023);
buf BUF1 (N2225, N2211);
and AND4 (N2226, N2225, N1596, N1839, N35);
and AND2 (N2227, N2209, N1022);
buf BUF1 (N2228, N2226);
and AND2 (N2229, N2218, N193);
nor NOR2 (N2230, N2224, N746);
nand NAND4 (N2231, N2229, N176, N684, N1420);
buf BUF1 (N2232, N2219);
and AND3 (N2233, N2230, N836, N1415);
nand NAND2 (N2234, N2227, N1369);
xor XOR2 (N2235, N2222, N875);
and AND2 (N2236, N2200, N1372);
nor NOR3 (N2237, N2232, N1382, N207);
xor XOR2 (N2238, N2231, N549);
nand NAND2 (N2239, N2236, N2219);
xor XOR2 (N2240, N2235, N1709);
and AND3 (N2241, N2228, N2092, N1436);
nand NAND2 (N2242, N2233, N253);
and AND2 (N2243, N2238, N1190);
xor XOR2 (N2244, N2223, N398);
xor XOR2 (N2245, N2207, N245);
buf BUF1 (N2246, N2241);
or OR2 (N2247, N2245, N913);
and AND3 (N2248, N2239, N584, N516);
xor XOR2 (N2249, N2201, N2248);
or OR3 (N2250, N123, N666, N194);
xor XOR2 (N2251, N2247, N1801);
nor NOR4 (N2252, N2240, N2039, N28, N929);
or OR2 (N2253, N2234, N1550);
nor NOR3 (N2254, N2237, N147, N212);
buf BUF1 (N2255, N2244);
buf BUF1 (N2256, N2242);
buf BUF1 (N2257, N2250);
xor XOR2 (N2258, N2243, N746);
xor XOR2 (N2259, N2253, N514);
xor XOR2 (N2260, N2255, N1655);
nand NAND4 (N2261, N2259, N685, N531, N1844);
or OR3 (N2262, N2260, N805, N546);
or OR4 (N2263, N2246, N60, N1123, N1113);
not NOT1 (N2264, N2257);
xor XOR2 (N2265, N2254, N890);
or OR4 (N2266, N2261, N906, N1082, N1541);
nand NAND2 (N2267, N2249, N504);
or OR2 (N2268, N2263, N1084);
xor XOR2 (N2269, N2256, N436);
nand NAND4 (N2270, N2252, N484, N1997, N1171);
nand NAND3 (N2271, N2267, N1948, N118);
xor XOR2 (N2272, N2268, N1105);
not NOT1 (N2273, N2264);
nor NOR2 (N2274, N2266, N2190);
not NOT1 (N2275, N2273);
nor NOR4 (N2276, N2269, N1240, N313, N2135);
not NOT1 (N2277, N2272);
and AND4 (N2278, N2275, N2238, N904, N605);
buf BUF1 (N2279, N2278);
not NOT1 (N2280, N2265);
nor NOR2 (N2281, N2277, N2060);
or OR4 (N2282, N2258, N716, N559, N1590);
nor NOR3 (N2283, N2281, N540, N2270);
buf BUF1 (N2284, N1293);
or OR2 (N2285, N2280, N681);
buf BUF1 (N2286, N2262);
xor XOR2 (N2287, N2276, N1439);
nor NOR2 (N2288, N2284, N346);
or OR3 (N2289, N2279, N2137, N514);
or OR2 (N2290, N2288, N1464);
not NOT1 (N2291, N2287);
buf BUF1 (N2292, N2271);
nor NOR4 (N2293, N2290, N1919, N295, N731);
nand NAND4 (N2294, N2285, N533, N1339, N1101);
xor XOR2 (N2295, N2293, N2229);
and AND2 (N2296, N2282, N569);
not NOT1 (N2297, N2289);
nand NAND3 (N2298, N2274, N42, N345);
xor XOR2 (N2299, N2251, N1648);
buf BUF1 (N2300, N2291);
not NOT1 (N2301, N2297);
buf BUF1 (N2302, N2295);
not NOT1 (N2303, N2286);
buf BUF1 (N2304, N2292);
buf BUF1 (N2305, N2304);
nor NOR4 (N2306, N2303, N377, N139, N538);
or OR2 (N2307, N2305, N1354);
nor NOR4 (N2308, N2296, N945, N2009, N1820);
or OR4 (N2309, N2283, N2161, N2070, N878);
and AND4 (N2310, N2307, N1915, N669, N700);
nand NAND4 (N2311, N2298, N1664, N1819, N720);
or OR4 (N2312, N2301, N1916, N300, N1245);
nand NAND3 (N2313, N2300, N2065, N1282);
or OR3 (N2314, N2311, N1197, N1743);
xor XOR2 (N2315, N2294, N1554);
buf BUF1 (N2316, N2315);
buf BUF1 (N2317, N2309);
not NOT1 (N2318, N2312);
xor XOR2 (N2319, N2310, N1537);
nor NOR3 (N2320, N2308, N1754, N822);
or OR4 (N2321, N2318, N1637, N1001, N8);
xor XOR2 (N2322, N2314, N749);
and AND3 (N2323, N2320, N1146, N905);
not NOT1 (N2324, N2323);
nand NAND2 (N2325, N2316, N1426);
xor XOR2 (N2326, N2302, N2085);
nand NAND2 (N2327, N2324, N49);
xor XOR2 (N2328, N2321, N2070);
buf BUF1 (N2329, N2322);
nor NOR3 (N2330, N2306, N1042, N934);
not NOT1 (N2331, N2313);
not NOT1 (N2332, N2317);
not NOT1 (N2333, N2299);
not NOT1 (N2334, N2326);
buf BUF1 (N2335, N2332);
or OR3 (N2336, N2334, N649, N2267);
nor NOR4 (N2337, N2333, N365, N691, N429);
or OR4 (N2338, N2335, N142, N323, N2087);
nor NOR3 (N2339, N2331, N940, N711);
xor XOR2 (N2340, N2337, N757);
and AND4 (N2341, N2330, N917, N899, N190);
and AND2 (N2342, N2341, N1321);
or OR3 (N2343, N2327, N920, N431);
buf BUF1 (N2344, N2336);
or OR3 (N2345, N2338, N1183, N1904);
or OR4 (N2346, N2325, N2332, N919, N2060);
xor XOR2 (N2347, N2339, N866);
xor XOR2 (N2348, N2345, N2171);
buf BUF1 (N2349, N2342);
xor XOR2 (N2350, N2329, N2308);
xor XOR2 (N2351, N2346, N245);
buf BUF1 (N2352, N2319);
nand NAND3 (N2353, N2351, N692, N1662);
and AND3 (N2354, N2347, N1235, N205);
buf BUF1 (N2355, N2352);
not NOT1 (N2356, N2348);
and AND3 (N2357, N2349, N1635, N65);
not NOT1 (N2358, N2350);
and AND3 (N2359, N2355, N1882, N2113);
or OR4 (N2360, N2340, N1249, N550, N1771);
not NOT1 (N2361, N2344);
not NOT1 (N2362, N2356);
buf BUF1 (N2363, N2359);
not NOT1 (N2364, N2354);
nand NAND2 (N2365, N2358, N1467);
not NOT1 (N2366, N2360);
not NOT1 (N2367, N2357);
nand NAND2 (N2368, N2361, N695);
nand NAND4 (N2369, N2367, N259, N342, N469);
buf BUF1 (N2370, N2364);
buf BUF1 (N2371, N2366);
and AND4 (N2372, N2363, N2023, N2365, N305);
not NOT1 (N2373, N2244);
xor XOR2 (N2374, N2370, N2163);
xor XOR2 (N2375, N2368, N2011);
and AND2 (N2376, N2369, N1242);
and AND2 (N2377, N2362, N1901);
and AND4 (N2378, N2372, N1677, N89, N1068);
not NOT1 (N2379, N2343);
nor NOR3 (N2380, N2373, N752, N882);
buf BUF1 (N2381, N2378);
or OR2 (N2382, N2371, N1436);
and AND2 (N2383, N2380, N1910);
nor NOR3 (N2384, N2379, N456, N511);
or OR2 (N2385, N2376, N994);
xor XOR2 (N2386, N2328, N1273);
or OR4 (N2387, N2382, N1224, N113, N861);
and AND2 (N2388, N2381, N154);
xor XOR2 (N2389, N2385, N2224);
or OR3 (N2390, N2375, N146, N2067);
nand NAND3 (N2391, N2387, N1085, N1446);
buf BUF1 (N2392, N2386);
nand NAND3 (N2393, N2392, N101, N1022);
and AND3 (N2394, N2377, N1387, N504);
or OR2 (N2395, N2374, N1520);
buf BUF1 (N2396, N2394);
not NOT1 (N2397, N2389);
nor NOR4 (N2398, N2395, N82, N1466, N2019);
and AND3 (N2399, N2390, N960, N1991);
nand NAND2 (N2400, N2384, N741);
buf BUF1 (N2401, N2388);
nor NOR4 (N2402, N2401, N1916, N1159, N811);
nand NAND3 (N2403, N2399, N2148, N2261);
not NOT1 (N2404, N2383);
and AND2 (N2405, N2391, N605);
nand NAND4 (N2406, N2403, N838, N1315, N1937);
nor NOR3 (N2407, N2353, N1868, N1777);
nor NOR4 (N2408, N2400, N2292, N811, N2107);
nand NAND3 (N2409, N2402, N1849, N812);
or OR4 (N2410, N2407, N103, N1384, N115);
nor NOR4 (N2411, N2406, N1884, N2356, N2270);
nand NAND4 (N2412, N2397, N882, N1532, N222);
xor XOR2 (N2413, N2393, N1392);
and AND2 (N2414, N2413, N476);
or OR3 (N2415, N2408, N141, N1218);
xor XOR2 (N2416, N2409, N2264);
or OR2 (N2417, N2416, N150);
not NOT1 (N2418, N2396);
and AND4 (N2419, N2410, N1486, N1476, N409);
or OR3 (N2420, N2419, N1092, N2102);
or OR2 (N2421, N2398, N1522);
nand NAND4 (N2422, N2415, N202, N2105, N32);
buf BUF1 (N2423, N2421);
buf BUF1 (N2424, N2405);
buf BUF1 (N2425, N2404);
not NOT1 (N2426, N2411);
and AND2 (N2427, N2418, N2182);
nand NAND3 (N2428, N2424, N2180, N663);
buf BUF1 (N2429, N2412);
or OR4 (N2430, N2427, N1010, N287, N2);
xor XOR2 (N2431, N2414, N1291);
nand NAND4 (N2432, N2417, N1818, N2413, N850);
and AND4 (N2433, N2423, N292, N2389, N371);
xor XOR2 (N2434, N2420, N569);
buf BUF1 (N2435, N2432);
buf BUF1 (N2436, N2433);
buf BUF1 (N2437, N2425);
or OR4 (N2438, N2436, N1673, N2376, N868);
nand NAND3 (N2439, N2428, N728, N1370);
nor NOR3 (N2440, N2422, N1822, N1210);
or OR2 (N2441, N2437, N733);
and AND2 (N2442, N2440, N2199);
buf BUF1 (N2443, N2434);
buf BUF1 (N2444, N2430);
and AND3 (N2445, N2444, N744, N10);
nand NAND2 (N2446, N2439, N1271);
not NOT1 (N2447, N2445);
nor NOR4 (N2448, N2441, N1168, N2133, N28);
not NOT1 (N2449, N2442);
buf BUF1 (N2450, N2429);
not NOT1 (N2451, N2431);
and AND2 (N2452, N2426, N1514);
nand NAND2 (N2453, N2449, N1862);
not NOT1 (N2454, N2447);
or OR2 (N2455, N2454, N2052);
nand NAND2 (N2456, N2450, N1049);
not NOT1 (N2457, N2448);
nor NOR2 (N2458, N2438, N1120);
nor NOR4 (N2459, N2457, N1890, N2442, N153);
nor NOR3 (N2460, N2456, N740, N198);
buf BUF1 (N2461, N2443);
nand NAND2 (N2462, N2458, N2191);
buf BUF1 (N2463, N2451);
nand NAND4 (N2464, N2460, N1364, N2126, N1861);
buf BUF1 (N2465, N2459);
not NOT1 (N2466, N2465);
or OR3 (N2467, N2464, N804, N879);
nand NAND2 (N2468, N2455, N1060);
nor NOR3 (N2469, N2435, N1480, N931);
or OR2 (N2470, N2468, N14);
buf BUF1 (N2471, N2462);
or OR3 (N2472, N2453, N1704, N1732);
xor XOR2 (N2473, N2471, N2438);
buf BUF1 (N2474, N2469);
xor XOR2 (N2475, N2452, N1974);
and AND4 (N2476, N2466, N2028, N2180, N234);
nand NAND3 (N2477, N2461, N1748, N1206);
not NOT1 (N2478, N2467);
and AND2 (N2479, N2475, N978);
not NOT1 (N2480, N2474);
nor NOR3 (N2481, N2446, N468, N105);
nor NOR2 (N2482, N2480, N227);
not NOT1 (N2483, N2476);
nor NOR2 (N2484, N2483, N1185);
buf BUF1 (N2485, N2473);
nand NAND3 (N2486, N2479, N2224, N934);
nand NAND3 (N2487, N2485, N1279, N983);
nor NOR2 (N2488, N2484, N1022);
nand NAND3 (N2489, N2477, N37, N1968);
or OR4 (N2490, N2481, N2417, N1755, N861);
xor XOR2 (N2491, N2486, N1134);
nor NOR3 (N2492, N2482, N727, N2463);
buf BUF1 (N2493, N1193);
xor XOR2 (N2494, N2489, N1665);
buf BUF1 (N2495, N2470);
nor NOR3 (N2496, N2490, N167, N2035);
buf BUF1 (N2497, N2472);
or OR3 (N2498, N2478, N53, N997);
nand NAND2 (N2499, N2488, N257);
and AND3 (N2500, N2496, N1975, N330);
and AND3 (N2501, N2497, N1242, N1871);
buf BUF1 (N2502, N2495);
nor NOR4 (N2503, N2501, N1959, N1634, N1402);
not NOT1 (N2504, N2500);
and AND4 (N2505, N2491, N2397, N792, N1740);
nand NAND2 (N2506, N2492, N1188);
not NOT1 (N2507, N2506);
or OR3 (N2508, N2504, N2502, N2201);
buf BUF1 (N2509, N1883);
buf BUF1 (N2510, N2503);
nand NAND2 (N2511, N2510, N626);
buf BUF1 (N2512, N2487);
buf BUF1 (N2513, N2498);
xor XOR2 (N2514, N2511, N2068);
xor XOR2 (N2515, N2512, N360);
and AND4 (N2516, N2509, N1164, N1322, N1882);
xor XOR2 (N2517, N2494, N847);
nor NOR2 (N2518, N2514, N2374);
not NOT1 (N2519, N2517);
not NOT1 (N2520, N2518);
nor NOR4 (N2521, N2507, N389, N902, N1324);
nor NOR4 (N2522, N2493, N410, N1549, N2255);
nand NAND2 (N2523, N2508, N2091);
not NOT1 (N2524, N2522);
nand NAND3 (N2525, N2519, N876, N2038);
or OR3 (N2526, N2516, N235, N1175);
xor XOR2 (N2527, N2523, N1696);
xor XOR2 (N2528, N2499, N1922);
and AND3 (N2529, N2527, N1356, N1276);
not NOT1 (N2530, N2525);
nand NAND2 (N2531, N2521, N2078);
nor NOR2 (N2532, N2530, N1899);
buf BUF1 (N2533, N2520);
xor XOR2 (N2534, N2529, N1530);
buf BUF1 (N2535, N2513);
nor NOR4 (N2536, N2526, N1541, N1636, N554);
xor XOR2 (N2537, N2528, N430);
or OR4 (N2538, N2524, N55, N1047, N1877);
or OR4 (N2539, N2532, N1624, N645, N2354);
nor NOR3 (N2540, N2535, N1727, N2430);
and AND3 (N2541, N2538, N1476, N839);
or OR4 (N2542, N2515, N2371, N1834, N2167);
not NOT1 (N2543, N2539);
buf BUF1 (N2544, N2541);
nand NAND3 (N2545, N2542, N2327, N946);
or OR2 (N2546, N2533, N591);
and AND3 (N2547, N2537, N1696, N765);
and AND2 (N2548, N2543, N1135);
or OR2 (N2549, N2544, N299);
and AND2 (N2550, N2548, N1492);
nand NAND3 (N2551, N2505, N1332, N1718);
not NOT1 (N2552, N2545);
buf BUF1 (N2553, N2531);
nand NAND2 (N2554, N2540, N922);
not NOT1 (N2555, N2546);
or OR2 (N2556, N2549, N2007);
buf BUF1 (N2557, N2547);
not NOT1 (N2558, N2556);
and AND2 (N2559, N2551, N647);
not NOT1 (N2560, N2552);
not NOT1 (N2561, N2554);
not NOT1 (N2562, N2560);
nor NOR2 (N2563, N2561, N568);
and AND3 (N2564, N2536, N808, N492);
and AND4 (N2565, N2558, N569, N991, N685);
or OR3 (N2566, N2564, N1008, N1421);
xor XOR2 (N2567, N2534, N1408);
nor NOR2 (N2568, N2555, N1501);
or OR4 (N2569, N2568, N170, N1764, N1556);
or OR4 (N2570, N2559, N1657, N439, N1930);
nand NAND2 (N2571, N2569, N2250);
or OR2 (N2572, N2570, N2243);
or OR2 (N2573, N2550, N372);
nor NOR2 (N2574, N2563, N1617);
buf BUF1 (N2575, N2571);
nand NAND4 (N2576, N2574, N194, N2279, N622);
buf BUF1 (N2577, N2572);
or OR3 (N2578, N2565, N710, N1072);
nand NAND4 (N2579, N2553, N1693, N2547, N2425);
or OR2 (N2580, N2579, N1055);
and AND4 (N2581, N2573, N1451, N136, N2335);
buf BUF1 (N2582, N2580);
or OR4 (N2583, N2576, N824, N2004, N798);
buf BUF1 (N2584, N2577);
buf BUF1 (N2585, N2578);
nand NAND3 (N2586, N2584, N1189, N2452);
xor XOR2 (N2587, N2583, N1220);
not NOT1 (N2588, N2581);
xor XOR2 (N2589, N2588, N133);
nor NOR4 (N2590, N2586, N2474, N1348, N771);
or OR3 (N2591, N2582, N1691, N1383);
or OR4 (N2592, N2591, N1041, N1333, N90);
nor NOR2 (N2593, N2566, N2544);
nand NAND2 (N2594, N2562, N1488);
not NOT1 (N2595, N2592);
or OR2 (N2596, N2567, N1232);
not NOT1 (N2597, N2589);
buf BUF1 (N2598, N2587);
nand NAND4 (N2599, N2590, N2409, N2296, N1134);
nand NAND4 (N2600, N2585, N1061, N2329, N1381);
or OR3 (N2601, N2600, N1706, N1048);
nand NAND3 (N2602, N2594, N91, N873);
not NOT1 (N2603, N2602);
nand NAND4 (N2604, N2575, N2384, N1112, N2311);
buf BUF1 (N2605, N2603);
buf BUF1 (N2606, N2595);
xor XOR2 (N2607, N2598, N1699);
nand NAND2 (N2608, N2607, N2245);
buf BUF1 (N2609, N2593);
or OR4 (N2610, N2605, N99, N1978, N2351);
and AND3 (N2611, N2610, N2033, N1407);
nor NOR4 (N2612, N2604, N478, N207, N794);
xor XOR2 (N2613, N2596, N75);
not NOT1 (N2614, N2599);
xor XOR2 (N2615, N2608, N1330);
or OR4 (N2616, N2611, N47, N2522, N2047);
xor XOR2 (N2617, N2609, N339);
and AND4 (N2618, N2557, N1554, N460, N772);
or OR2 (N2619, N2616, N588);
nor NOR4 (N2620, N2597, N85, N1069, N1889);
xor XOR2 (N2621, N2617, N17);
not NOT1 (N2622, N2619);
buf BUF1 (N2623, N2618);
xor XOR2 (N2624, N2622, N777);
or OR4 (N2625, N2620, N188, N1351, N1444);
nand NAND4 (N2626, N2601, N1409, N1561, N2619);
nor NOR2 (N2627, N2615, N124);
and AND2 (N2628, N2612, N103);
not NOT1 (N2629, N2621);
xor XOR2 (N2630, N2613, N1540);
nand NAND3 (N2631, N2626, N1386, N1093);
or OR2 (N2632, N2631, N1738);
nand NAND2 (N2633, N2627, N1165);
nor NOR2 (N2634, N2629, N81);
nand NAND3 (N2635, N2606, N917, N160);
xor XOR2 (N2636, N2632, N1954);
buf BUF1 (N2637, N2633);
xor XOR2 (N2638, N2624, N118);
and AND2 (N2639, N2614, N659);
buf BUF1 (N2640, N2638);
nor NOR2 (N2641, N2630, N309);
nor NOR3 (N2642, N2641, N1530, N1593);
nand NAND2 (N2643, N2636, N2245);
xor XOR2 (N2644, N2637, N1088);
nor NOR4 (N2645, N2642, N2443, N1006, N2099);
xor XOR2 (N2646, N2639, N1754);
xor XOR2 (N2647, N2628, N1615);
xor XOR2 (N2648, N2645, N1291);
nand NAND4 (N2649, N2634, N2236, N530, N2092);
nor NOR2 (N2650, N2625, N1953);
or OR4 (N2651, N2649, N2124, N1107, N435);
and AND3 (N2652, N2623, N248, N1445);
xor XOR2 (N2653, N2650, N814);
not NOT1 (N2654, N2644);
nor NOR2 (N2655, N2653, N650);
xor XOR2 (N2656, N2654, N1081);
nand NAND2 (N2657, N2643, N537);
and AND2 (N2658, N2646, N908);
not NOT1 (N2659, N2657);
nand NAND2 (N2660, N2647, N2435);
and AND2 (N2661, N2635, N666);
or OR4 (N2662, N2648, N2005, N1856, N1577);
not NOT1 (N2663, N2662);
nand NAND4 (N2664, N2660, N1422, N1706, N1136);
and AND3 (N2665, N2659, N2620, N2445);
or OR4 (N2666, N2655, N67, N1862, N1179);
nor NOR4 (N2667, N2665, N2064, N676, N2442);
or OR4 (N2668, N2661, N1561, N2410, N1356);
and AND2 (N2669, N2667, N66);
nor NOR2 (N2670, N2656, N2076);
and AND3 (N2671, N2658, N2657, N726);
and AND2 (N2672, N2663, N1749);
nand NAND3 (N2673, N2671, N438, N1763);
nor NOR3 (N2674, N2664, N2337, N1289);
buf BUF1 (N2675, N2640);
and AND4 (N2676, N2672, N609, N2444, N986);
and AND4 (N2677, N2652, N1549, N2381, N2214);
and AND3 (N2678, N2677, N305, N1797);
or OR4 (N2679, N2669, N1982, N327, N2583);
nand NAND2 (N2680, N2675, N151);
xor XOR2 (N2681, N2666, N2625);
or OR3 (N2682, N2651, N2553, N944);
nor NOR4 (N2683, N2680, N287, N431, N2351);
and AND4 (N2684, N2679, N2145, N1951, N1299);
nand NAND3 (N2685, N2683, N1389, N1079);
and AND2 (N2686, N2668, N1132);
or OR4 (N2687, N2681, N1575, N1335, N185);
nand NAND3 (N2688, N2678, N1707, N2614);
nor NOR2 (N2689, N2684, N232);
xor XOR2 (N2690, N2674, N1967);
and AND2 (N2691, N2670, N1642);
and AND3 (N2692, N2690, N319, N2075);
nand NAND2 (N2693, N2685, N2644);
or OR3 (N2694, N2686, N2208, N2083);
and AND4 (N2695, N2694, N2253, N331, N547);
or OR4 (N2696, N2676, N1997, N209, N389);
or OR4 (N2697, N2696, N884, N2671, N745);
nand NAND4 (N2698, N2689, N414, N1862, N2208);
or OR2 (N2699, N2682, N940);
or OR2 (N2700, N2688, N1655);
and AND2 (N2701, N2697, N1911);
buf BUF1 (N2702, N2687);
xor XOR2 (N2703, N2693, N2685);
not NOT1 (N2704, N2702);
nor NOR4 (N2705, N2692, N284, N2438, N172);
and AND2 (N2706, N2704, N2320);
or OR4 (N2707, N2706, N871, N2606, N518);
and AND3 (N2708, N2699, N2459, N1171);
xor XOR2 (N2709, N2691, N2456);
not NOT1 (N2710, N2698);
buf BUF1 (N2711, N2703);
nand NAND4 (N2712, N2708, N220, N548, N957);
not NOT1 (N2713, N2701);
or OR4 (N2714, N2711, N1386, N2064, N1394);
not NOT1 (N2715, N2673);
not NOT1 (N2716, N2709);
not NOT1 (N2717, N2714);
buf BUF1 (N2718, N2707);
nor NOR4 (N2719, N2713, N2584, N1588, N2684);
nand NAND4 (N2720, N2719, N449, N2685, N699);
xor XOR2 (N2721, N2718, N1679);
nand NAND2 (N2722, N2710, N2632);
nor NOR2 (N2723, N2721, N1560);
buf BUF1 (N2724, N2720);
nand NAND2 (N2725, N2700, N1271);
or OR2 (N2726, N2716, N1459);
nor NOR4 (N2727, N2726, N128, N837, N1145);
nand NAND2 (N2728, N2712, N2536);
not NOT1 (N2729, N2695);
and AND4 (N2730, N2723, N1999, N1103, N2407);
nor NOR3 (N2731, N2724, N85, N2143);
and AND4 (N2732, N2717, N2357, N999, N2242);
and AND2 (N2733, N2731, N1723);
xor XOR2 (N2734, N2722, N517);
not NOT1 (N2735, N2715);
or OR3 (N2736, N2729, N503, N811);
not NOT1 (N2737, N2732);
and AND2 (N2738, N2725, N1122);
and AND4 (N2739, N2738, N2630, N1899, N1248);
xor XOR2 (N2740, N2736, N1567);
xor XOR2 (N2741, N2705, N1358);
xor XOR2 (N2742, N2728, N2419);
buf BUF1 (N2743, N2741);
not NOT1 (N2744, N2730);
and AND2 (N2745, N2744, N316);
not NOT1 (N2746, N2740);
nor NOR4 (N2747, N2745, N303, N527, N365);
xor XOR2 (N2748, N2733, N693);
nor NOR3 (N2749, N2727, N165, N1666);
buf BUF1 (N2750, N2742);
or OR3 (N2751, N2747, N508, N1072);
xor XOR2 (N2752, N2735, N908);
or OR3 (N2753, N2734, N2222, N1643);
or OR2 (N2754, N2752, N1112);
buf BUF1 (N2755, N2743);
xor XOR2 (N2756, N2737, N1534);
nand NAND3 (N2757, N2739, N2744, N1834);
buf BUF1 (N2758, N2753);
xor XOR2 (N2759, N2749, N1050);
or OR3 (N2760, N2751, N370, N2559);
not NOT1 (N2761, N2748);
not NOT1 (N2762, N2746);
buf BUF1 (N2763, N2754);
nor NOR2 (N2764, N2761, N1967);
nand NAND4 (N2765, N2750, N886, N1771, N1464);
or OR3 (N2766, N2759, N1363, N2190);
nor NOR4 (N2767, N2755, N2480, N1796, N2246);
nor NOR3 (N2768, N2758, N1609, N2766);
nand NAND3 (N2769, N256, N844, N810);
or OR3 (N2770, N2767, N509, N803);
nor NOR2 (N2771, N2762, N1414);
and AND4 (N2772, N2763, N1025, N958, N1453);
not NOT1 (N2773, N2768);
xor XOR2 (N2774, N2772, N184);
or OR3 (N2775, N2756, N275, N1795);
xor XOR2 (N2776, N2771, N1564);
not NOT1 (N2777, N2770);
buf BUF1 (N2778, N2775);
nand NAND2 (N2779, N2765, N1574);
and AND4 (N2780, N2773, N2742, N1832, N1018);
not NOT1 (N2781, N2774);
and AND4 (N2782, N2779, N349, N348, N2662);
buf BUF1 (N2783, N2778);
and AND3 (N2784, N2757, N38, N1092);
xor XOR2 (N2785, N2780, N1045);
nor NOR4 (N2786, N2784, N2486, N2327, N2454);
nor NOR4 (N2787, N2769, N288, N2555, N974);
not NOT1 (N2788, N2764);
and AND3 (N2789, N2760, N459, N622);
buf BUF1 (N2790, N2782);
nor NOR3 (N2791, N2777, N601, N2329);
nand NAND3 (N2792, N2781, N713, N692);
xor XOR2 (N2793, N2776, N1389);
nand NAND4 (N2794, N2783, N72, N1245, N2468);
nor NOR3 (N2795, N2790, N2094, N380);
nor NOR2 (N2796, N2787, N92);
or OR3 (N2797, N2796, N855, N1155);
buf BUF1 (N2798, N2794);
not NOT1 (N2799, N2793);
and AND2 (N2800, N2795, N2532);
buf BUF1 (N2801, N2791);
xor XOR2 (N2802, N2785, N1529);
xor XOR2 (N2803, N2797, N127);
nor NOR2 (N2804, N2786, N714);
xor XOR2 (N2805, N2804, N21);
nor NOR3 (N2806, N2789, N663, N1667);
buf BUF1 (N2807, N2805);
and AND4 (N2808, N2807, N2425, N1894, N2425);
nor NOR4 (N2809, N2803, N1519, N105, N2228);
buf BUF1 (N2810, N2800);
not NOT1 (N2811, N2808);
buf BUF1 (N2812, N2801);
nor NOR2 (N2813, N2810, N394);
xor XOR2 (N2814, N2806, N1915);
buf BUF1 (N2815, N2809);
xor XOR2 (N2816, N2812, N2597);
not NOT1 (N2817, N2811);
and AND2 (N2818, N2814, N788);
nor NOR2 (N2819, N2798, N1623);
and AND3 (N2820, N2799, N1997, N1472);
nand NAND3 (N2821, N2820, N570, N641);
nor NOR3 (N2822, N2802, N2701, N1859);
nand NAND3 (N2823, N2818, N2058, N1521);
xor XOR2 (N2824, N2788, N1444);
or OR4 (N2825, N2815, N2339, N2007, N2568);
or OR2 (N2826, N2823, N164);
buf BUF1 (N2827, N2822);
buf BUF1 (N2828, N2819);
and AND4 (N2829, N2813, N342, N1237, N63);
or OR4 (N2830, N2821, N2822, N1365, N293);
xor XOR2 (N2831, N2824, N2577);
not NOT1 (N2832, N2829);
nand NAND4 (N2833, N2792, N1693, N1713, N984);
or OR4 (N2834, N2825, N254, N2627, N1500);
nor NOR2 (N2835, N2828, N710);
not NOT1 (N2836, N2830);
nor NOR3 (N2837, N2826, N2542, N1745);
or OR2 (N2838, N2834, N918);
or OR4 (N2839, N2817, N729, N1766, N1787);
or OR4 (N2840, N2836, N1057, N2615, N1514);
nand NAND2 (N2841, N2837, N1759);
xor XOR2 (N2842, N2840, N1869);
or OR4 (N2843, N2831, N1899, N1375, N1031);
and AND2 (N2844, N2832, N2133);
buf BUF1 (N2845, N2844);
buf BUF1 (N2846, N2827);
not NOT1 (N2847, N2846);
not NOT1 (N2848, N2845);
nand NAND4 (N2849, N2842, N1813, N1916, N2146);
buf BUF1 (N2850, N2833);
nor NOR3 (N2851, N2849, N1248, N2430);
nand NAND2 (N2852, N2816, N1846);
nor NOR3 (N2853, N2850, N2415, N1940);
not NOT1 (N2854, N2852);
and AND2 (N2855, N2835, N2049);
or OR4 (N2856, N2855, N581, N718, N1742);
and AND2 (N2857, N2839, N523);
and AND3 (N2858, N2851, N802, N1127);
or OR2 (N2859, N2857, N1500);
buf BUF1 (N2860, N2838);
nor NOR3 (N2861, N2843, N2295, N1481);
nor NOR4 (N2862, N2859, N149, N2347, N2524);
not NOT1 (N2863, N2856);
not NOT1 (N2864, N2854);
buf BUF1 (N2865, N2863);
not NOT1 (N2866, N2862);
nand NAND4 (N2867, N2847, N2182, N1045, N2299);
not NOT1 (N2868, N2867);
nor NOR4 (N2869, N2848, N1982, N2574, N1924);
xor XOR2 (N2870, N2858, N312);
xor XOR2 (N2871, N2853, N192);
and AND3 (N2872, N2864, N1646, N2149);
nor NOR4 (N2873, N2861, N9, N471, N33);
nor NOR3 (N2874, N2865, N2170, N1111);
not NOT1 (N2875, N2874);
not NOT1 (N2876, N2875);
nand NAND4 (N2877, N2866, N1657, N1007, N2280);
not NOT1 (N2878, N2871);
and AND4 (N2879, N2876, N666, N1962, N1114);
and AND2 (N2880, N2870, N1797);
nand NAND4 (N2881, N2878, N25, N1543, N290);
xor XOR2 (N2882, N2877, N1268);
nand NAND4 (N2883, N2881, N1714, N2017, N1826);
nor NOR2 (N2884, N2873, N1245);
or OR4 (N2885, N2869, N821, N173, N1975);
nor NOR4 (N2886, N2885, N1243, N2876, N1091);
xor XOR2 (N2887, N2841, N2589);
not NOT1 (N2888, N2872);
nand NAND2 (N2889, N2883, N2869);
nor NOR3 (N2890, N2886, N1116, N771);
or OR2 (N2891, N2880, N2382);
nand NAND2 (N2892, N2888, N1235);
and AND4 (N2893, N2890, N645, N2650, N1212);
xor XOR2 (N2894, N2882, N2698);
nand NAND3 (N2895, N2887, N2087, N458);
nor NOR2 (N2896, N2891, N736);
not NOT1 (N2897, N2868);
nor NOR4 (N2898, N2889, N1091, N2770, N77);
buf BUF1 (N2899, N2894);
buf BUF1 (N2900, N2897);
nor NOR4 (N2901, N2892, N1028, N1825, N1308);
not NOT1 (N2902, N2879);
and AND4 (N2903, N2895, N1673, N293, N1918);
nor NOR2 (N2904, N2896, N1143);
xor XOR2 (N2905, N2901, N2141);
and AND4 (N2906, N2904, N1892, N2244, N2596);
nand NAND2 (N2907, N2893, N1210);
nand NAND3 (N2908, N2906, N2481, N119);
or OR2 (N2909, N2902, N2749);
buf BUF1 (N2910, N2903);
not NOT1 (N2911, N2884);
and AND4 (N2912, N2907, N1677, N2645, N1480);
xor XOR2 (N2913, N2911, N2472);
nor NOR4 (N2914, N2909, N459, N1465, N260);
not NOT1 (N2915, N2910);
not NOT1 (N2916, N2913);
and AND4 (N2917, N2898, N924, N24, N2582);
and AND4 (N2918, N2916, N1233, N1011, N782);
nand NAND2 (N2919, N2900, N2001);
nand NAND2 (N2920, N2860, N251);
nor NOR4 (N2921, N2914, N1714, N112, N46);
not NOT1 (N2922, N2912);
buf BUF1 (N2923, N2899);
and AND2 (N2924, N2920, N1634);
xor XOR2 (N2925, N2915, N2117);
nor NOR3 (N2926, N2919, N500, N1141);
or OR3 (N2927, N2922, N612, N41);
nand NAND4 (N2928, N2918, N2846, N523, N1141);
xor XOR2 (N2929, N2924, N1119);
xor XOR2 (N2930, N2927, N629);
not NOT1 (N2931, N2930);
and AND4 (N2932, N2931, N175, N643, N2832);
not NOT1 (N2933, N2932);
nor NOR2 (N2934, N2926, N2577);
and AND2 (N2935, N2934, N2482);
xor XOR2 (N2936, N2905, N1370);
or OR4 (N2937, N2908, N2629, N2633, N1597);
nand NAND2 (N2938, N2921, N2937);
and AND4 (N2939, N359, N1017, N7, N1646);
nor NOR2 (N2940, N2929, N54);
or OR2 (N2941, N2933, N1952);
xor XOR2 (N2942, N2939, N1057);
nand NAND3 (N2943, N2938, N314, N221);
or OR4 (N2944, N2936, N1961, N2728, N1723);
nor NOR3 (N2945, N2941, N1560, N1935);
buf BUF1 (N2946, N2940);
not NOT1 (N2947, N2917);
xor XOR2 (N2948, N2935, N902);
nor NOR2 (N2949, N2942, N2944);
buf BUF1 (N2950, N1879);
or OR3 (N2951, N2950, N2561, N534);
xor XOR2 (N2952, N2945, N589);
nand NAND2 (N2953, N2948, N1009);
buf BUF1 (N2954, N2923);
and AND3 (N2955, N2943, N86, N2667);
nor NOR2 (N2956, N2925, N255);
nand NAND3 (N2957, N2946, N2371, N20);
xor XOR2 (N2958, N2954, N2266);
nand NAND4 (N2959, N2957, N452, N2633, N2464);
or OR2 (N2960, N2958, N2289);
and AND3 (N2961, N2952, N1204, N1766);
xor XOR2 (N2962, N2947, N1751);
nor NOR3 (N2963, N2949, N1636, N2579);
and AND3 (N2964, N2960, N1388, N937);
xor XOR2 (N2965, N2955, N2811);
xor XOR2 (N2966, N2959, N2274);
nor NOR2 (N2967, N2951, N1335);
not NOT1 (N2968, N2965);
nor NOR2 (N2969, N2956, N47);
xor XOR2 (N2970, N2928, N2750);
nand NAND3 (N2971, N2966, N2469, N1217);
and AND3 (N2972, N2970, N1348, N2681);
xor XOR2 (N2973, N2972, N1218);
xor XOR2 (N2974, N2963, N2433);
xor XOR2 (N2975, N2969, N1343);
and AND3 (N2976, N2971, N1379, N2379);
xor XOR2 (N2977, N2964, N2935);
and AND3 (N2978, N2968, N2764, N2883);
and AND2 (N2979, N2962, N1288);
xor XOR2 (N2980, N2973, N657);
buf BUF1 (N2981, N2953);
or OR4 (N2982, N2980, N351, N2305, N2835);
and AND3 (N2983, N2975, N1840, N12);
and AND2 (N2984, N2961, N2010);
buf BUF1 (N2985, N2979);
and AND4 (N2986, N2978, N521, N2829, N606);
and AND2 (N2987, N2984, N1667);
xor XOR2 (N2988, N2967, N1264);
xor XOR2 (N2989, N2977, N1428);
and AND4 (N2990, N2981, N2443, N228, N1024);
xor XOR2 (N2991, N2976, N2702);
or OR3 (N2992, N2985, N895, N2507);
or OR2 (N2993, N2987, N574);
nand NAND4 (N2994, N2993, N1916, N1748, N2547);
or OR3 (N2995, N2988, N2206, N1080);
nor NOR4 (N2996, N2974, N1599, N2133, N1137);
nand NAND3 (N2997, N2994, N2838, N1492);
or OR2 (N2998, N2989, N2210);
nand NAND2 (N2999, N2998, N2934);
xor XOR2 (N3000, N2992, N280);
nand NAND3 (N3001, N3000, N2151, N2026);
or OR3 (N3002, N2983, N1695, N207);
nand NAND2 (N3003, N2996, N2843);
or OR3 (N3004, N2990, N2457, N2767);
not NOT1 (N3005, N3003);
xor XOR2 (N3006, N2986, N2297);
or OR4 (N3007, N2991, N2052, N1073, N1981);
nor NOR2 (N3008, N3002, N1221);
nand NAND2 (N3009, N2995, N316);
nor NOR2 (N3010, N2999, N931);
xor XOR2 (N3011, N3006, N2859);
buf BUF1 (N3012, N2982);
and AND2 (N3013, N3008, N3005);
buf BUF1 (N3014, N1371);
not NOT1 (N3015, N3012);
nor NOR2 (N3016, N3011, N1955);
xor XOR2 (N3017, N3015, N2249);
nor NOR4 (N3018, N3007, N296, N2245, N1749);
or OR3 (N3019, N3001, N1593, N2094);
not NOT1 (N3020, N3013);
buf BUF1 (N3021, N3020);
xor XOR2 (N3022, N3010, N157);
or OR3 (N3023, N3016, N1088, N446);
nor NOR2 (N3024, N3021, N2111);
nor NOR4 (N3025, N3004, N694, N1639, N1849);
xor XOR2 (N3026, N3019, N1347);
nand NAND3 (N3027, N3009, N237, N2252);
or OR4 (N3028, N3018, N2469, N2839, N85);
and AND2 (N3029, N3025, N1956);
or OR4 (N3030, N3027, N558, N2839, N2859);
nor NOR2 (N3031, N3030, N2237);
and AND3 (N3032, N3014, N2969, N958);
buf BUF1 (N3033, N3022);
and AND3 (N3034, N3032, N465, N370);
xor XOR2 (N3035, N3033, N143);
not NOT1 (N3036, N3017);
buf BUF1 (N3037, N3028);
and AND4 (N3038, N3031, N2248, N1660, N86);
or OR3 (N3039, N3029, N2266, N1339);
buf BUF1 (N3040, N3034);
and AND3 (N3041, N2997, N2326, N809);
not NOT1 (N3042, N3036);
nor NOR2 (N3043, N3042, N1274);
buf BUF1 (N3044, N3035);
not NOT1 (N3045, N3038);
or OR4 (N3046, N3041, N1441, N1620, N1003);
nor NOR4 (N3047, N3045, N2444, N1140, N2899);
nor NOR3 (N3048, N3037, N2084, N298);
buf BUF1 (N3049, N3046);
or OR4 (N3050, N3023, N2792, N2781, N2134);
nand NAND4 (N3051, N3044, N618, N369, N1197);
nand NAND3 (N3052, N3047, N789, N174);
buf BUF1 (N3053, N3026);
xor XOR2 (N3054, N3052, N1428);
nand NAND3 (N3055, N3051, N980, N2987);
not NOT1 (N3056, N3053);
nand NAND4 (N3057, N3055, N2443, N2793, N1322);
nand NAND4 (N3058, N3043, N979, N2764, N90);
and AND2 (N3059, N3039, N678);
not NOT1 (N3060, N3054);
not NOT1 (N3061, N3059);
nand NAND2 (N3062, N3057, N1805);
xor XOR2 (N3063, N3049, N2536);
nand NAND3 (N3064, N3050, N1923, N1244);
buf BUF1 (N3065, N3024);
xor XOR2 (N3066, N3063, N2675);
xor XOR2 (N3067, N3061, N2686);
and AND4 (N3068, N3040, N2952, N1804, N615);
nand NAND3 (N3069, N3067, N1433, N90);
or OR2 (N3070, N3048, N2081);
buf BUF1 (N3071, N3062);
and AND4 (N3072, N3065, N2353, N2858, N831);
buf BUF1 (N3073, N3058);
nor NOR3 (N3074, N3060, N1414, N668);
xor XOR2 (N3075, N3066, N2001);
buf BUF1 (N3076, N3064);
and AND4 (N3077, N3070, N2996, N1998, N269);
or OR2 (N3078, N3074, N811);
and AND2 (N3079, N3072, N1309);
nand NAND2 (N3080, N3068, N1710);
or OR3 (N3081, N3071, N1499, N1147);
nand NAND2 (N3082, N3081, N164);
or OR3 (N3083, N3079, N2296, N258);
xor XOR2 (N3084, N3075, N2845);
xor XOR2 (N3085, N3073, N1915);
nor NOR3 (N3086, N3069, N128, N1231);
not NOT1 (N3087, N3085);
and AND2 (N3088, N3087, N2821);
buf BUF1 (N3089, N3076);
xor XOR2 (N3090, N3084, N1302);
buf BUF1 (N3091, N3088);
nand NAND4 (N3092, N3056, N339, N355, N243);
buf BUF1 (N3093, N3080);
or OR2 (N3094, N3090, N675);
and AND2 (N3095, N3082, N1712);
or OR2 (N3096, N3091, N32);
buf BUF1 (N3097, N3083);
not NOT1 (N3098, N3086);
or OR2 (N3099, N3093, N567);
and AND2 (N3100, N3096, N2980);
nor NOR3 (N3101, N3100, N1241, N1892);
or OR2 (N3102, N3099, N2965);
nand NAND3 (N3103, N3097, N258, N485);
not NOT1 (N3104, N3102);
or OR4 (N3105, N3104, N2599, N252, N3102);
not NOT1 (N3106, N3089);
nor NOR3 (N3107, N3095, N215, N885);
and AND4 (N3108, N3078, N2321, N829, N1097);
and AND4 (N3109, N3108, N1116, N254, N102);
nand NAND2 (N3110, N3077, N492);
or OR2 (N3111, N3098, N177);
and AND3 (N3112, N3092, N766, N900);
nor NOR4 (N3113, N3106, N1669, N503, N2020);
not NOT1 (N3114, N3101);
buf BUF1 (N3115, N3094);
nand NAND4 (N3116, N3115, N2402, N486, N1985);
xor XOR2 (N3117, N3107, N3018);
buf BUF1 (N3118, N3110);
nand NAND4 (N3119, N3117, N2383, N1328, N622);
xor XOR2 (N3120, N3109, N922);
xor XOR2 (N3121, N3113, N1693);
buf BUF1 (N3122, N3120);
buf BUF1 (N3123, N3121);
and AND3 (N3124, N3118, N1759, N1586);
or OR3 (N3125, N3124, N2306, N1595);
or OR2 (N3126, N3125, N180);
not NOT1 (N3127, N3111);
nand NAND2 (N3128, N3122, N2869);
and AND3 (N3129, N3126, N2294, N1429);
nor NOR3 (N3130, N3129, N840, N2457);
or OR2 (N3131, N3130, N1324);
or OR3 (N3132, N3123, N842, N2764);
xor XOR2 (N3133, N3132, N3116);
xor XOR2 (N3134, N715, N2829);
not NOT1 (N3135, N3131);
or OR3 (N3136, N3119, N1857, N645);
or OR2 (N3137, N3136, N890);
and AND2 (N3138, N3133, N1471);
or OR2 (N3139, N3135, N587);
buf BUF1 (N3140, N3105);
buf BUF1 (N3141, N3138);
buf BUF1 (N3142, N3140);
and AND3 (N3143, N3112, N1907, N2407);
xor XOR2 (N3144, N3143, N653);
xor XOR2 (N3145, N3103, N754);
buf BUF1 (N3146, N3134);
and AND4 (N3147, N3127, N419, N43, N3050);
and AND4 (N3148, N3145, N6, N1500, N1555);
not NOT1 (N3149, N3141);
buf BUF1 (N3150, N3147);
not NOT1 (N3151, N3137);
not NOT1 (N3152, N3139);
nand NAND3 (N3153, N3128, N636, N2723);
nor NOR2 (N3154, N3142, N328);
not NOT1 (N3155, N3152);
nand NAND2 (N3156, N3148, N1808);
or OR2 (N3157, N3144, N1617);
or OR3 (N3158, N3146, N955, N1570);
buf BUF1 (N3159, N3151);
and AND3 (N3160, N3157, N433, N2566);
nor NOR3 (N3161, N3149, N2228, N949);
or OR4 (N3162, N3160, N1881, N582, N33);
buf BUF1 (N3163, N3114);
and AND2 (N3164, N3158, N2751);
buf BUF1 (N3165, N3155);
buf BUF1 (N3166, N3159);
or OR3 (N3167, N3156, N509, N2373);
nor NOR2 (N3168, N3154, N2424);
nor NOR3 (N3169, N3150, N71, N674);
and AND2 (N3170, N3153, N701);
nand NAND2 (N3171, N3169, N1162);
nor NOR3 (N3172, N3166, N793, N549);
nand NAND2 (N3173, N3167, N1620);
nand NAND4 (N3174, N3170, N157, N826, N2831);
xor XOR2 (N3175, N3165, N2188);
or OR4 (N3176, N3173, N3081, N2183, N1548);
nand NAND3 (N3177, N3172, N1319, N2631);
and AND3 (N3178, N3177, N2523, N604);
and AND3 (N3179, N3163, N954, N3056);
nand NAND4 (N3180, N3161, N1822, N397, N1745);
or OR2 (N3181, N3162, N2639);
buf BUF1 (N3182, N3179);
nand NAND3 (N3183, N3176, N2212, N1802);
buf BUF1 (N3184, N3180);
not NOT1 (N3185, N3164);
nand NAND4 (N3186, N3184, N2926, N111, N360);
and AND4 (N3187, N3175, N739, N1534, N1822);
not NOT1 (N3188, N3183);
nand NAND2 (N3189, N3185, N2910);
nor NOR4 (N3190, N3182, N2590, N2371, N1438);
not NOT1 (N3191, N3168);
xor XOR2 (N3192, N3190, N2180);
xor XOR2 (N3193, N3181, N1648);
or OR2 (N3194, N3191, N2059);
or OR4 (N3195, N3187, N2381, N216, N1225);
buf BUF1 (N3196, N3192);
and AND2 (N3197, N3194, N292);
xor XOR2 (N3198, N3178, N2412);
or OR4 (N3199, N3198, N44, N2415, N1130);
not NOT1 (N3200, N3195);
and AND2 (N3201, N3186, N2489);
xor XOR2 (N3202, N3200, N692);
nand NAND2 (N3203, N3193, N3066);
not NOT1 (N3204, N3171);
or OR2 (N3205, N3202, N543);
buf BUF1 (N3206, N3201);
nor NOR3 (N3207, N3206, N1936, N90);
or OR4 (N3208, N3205, N44, N2565, N1780);
nand NAND3 (N3209, N3189, N2338, N1526);
not NOT1 (N3210, N3196);
buf BUF1 (N3211, N3174);
nand NAND2 (N3212, N3208, N1704);
or OR3 (N3213, N3197, N2330, N2434);
nand NAND3 (N3214, N3199, N1755, N1327);
xor XOR2 (N3215, N3209, N1707);
or OR4 (N3216, N3212, N1456, N2574, N1228);
buf BUF1 (N3217, N3203);
nand NAND4 (N3218, N3210, N1274, N3177, N1082);
buf BUF1 (N3219, N3214);
xor XOR2 (N3220, N3207, N1891);
or OR4 (N3221, N3216, N1187, N1394, N578);
nor NOR3 (N3222, N3218, N2738, N1363);
nor NOR4 (N3223, N3215, N1312, N213, N915);
and AND3 (N3224, N3213, N2771, N928);
buf BUF1 (N3225, N3221);
or OR2 (N3226, N3219, N2857);
buf BUF1 (N3227, N3204);
and AND3 (N3228, N3226, N2359, N1489);
nor NOR4 (N3229, N3220, N2836, N3106, N1344);
xor XOR2 (N3230, N3225, N1068);
nor NOR4 (N3231, N3228, N166, N1813, N2379);
nand NAND2 (N3232, N3217, N580);
or OR3 (N3233, N3188, N282, N854);
or OR2 (N3234, N3211, N1840);
xor XOR2 (N3235, N3233, N1632);
not NOT1 (N3236, N3235);
and AND2 (N3237, N3229, N336);
nor NOR4 (N3238, N3230, N860, N2580, N11);
nor NOR3 (N3239, N3231, N669, N2507);
or OR3 (N3240, N3223, N12, N2196);
not NOT1 (N3241, N3238);
not NOT1 (N3242, N3239);
nand NAND3 (N3243, N3236, N1739, N846);
or OR3 (N3244, N3243, N1397, N3162);
and AND2 (N3245, N3234, N1181);
buf BUF1 (N3246, N3227);
xor XOR2 (N3247, N3242, N2072);
not NOT1 (N3248, N3237);
buf BUF1 (N3249, N3245);
buf BUF1 (N3250, N3248);
nor NOR4 (N3251, N3247, N1747, N633, N2998);
xor XOR2 (N3252, N3250, N1102);
or OR4 (N3253, N3244, N478, N1549, N2220);
buf BUF1 (N3254, N3240);
not NOT1 (N3255, N3253);
and AND2 (N3256, N3252, N1337);
not NOT1 (N3257, N3255);
or OR3 (N3258, N3224, N1866, N894);
not NOT1 (N3259, N3256);
buf BUF1 (N3260, N3249);
and AND2 (N3261, N3251, N2241);
buf BUF1 (N3262, N3241);
and AND4 (N3263, N3260, N2192, N1086, N3250);
not NOT1 (N3264, N3262);
nor NOR3 (N3265, N3232, N2139, N2366);
nor NOR4 (N3266, N3222, N1447, N930, N1466);
or OR4 (N3267, N3259, N1985, N1527, N2887);
or OR2 (N3268, N3264, N653);
nand NAND3 (N3269, N3261, N140, N2012);
not NOT1 (N3270, N3266);
not NOT1 (N3271, N3265);
and AND2 (N3272, N3267, N1643);
not NOT1 (N3273, N3271);
nand NAND2 (N3274, N3258, N47);
or OR3 (N3275, N3270, N2426, N243);
nor NOR4 (N3276, N3263, N2981, N644, N961);
xor XOR2 (N3277, N3274, N2135);
buf BUF1 (N3278, N3276);
nand NAND2 (N3279, N3273, N727);
xor XOR2 (N3280, N3272, N561);
or OR4 (N3281, N3257, N793, N792, N1770);
and AND2 (N3282, N3277, N2802);
nand NAND4 (N3283, N3275, N3197, N2499, N903);
or OR2 (N3284, N3282, N765);
xor XOR2 (N3285, N3246, N710);
buf BUF1 (N3286, N3281);
nor NOR4 (N3287, N3283, N2608, N2820, N877);
not NOT1 (N3288, N3280);
not NOT1 (N3289, N3287);
or OR4 (N3290, N3286, N2493, N1277, N491);
xor XOR2 (N3291, N3254, N1960);
xor XOR2 (N3292, N3289, N2908);
nor NOR2 (N3293, N3269, N1098);
xor XOR2 (N3294, N3268, N2086);
not NOT1 (N3295, N3278);
xor XOR2 (N3296, N3284, N708);
buf BUF1 (N3297, N3291);
xor XOR2 (N3298, N3297, N2752);
xor XOR2 (N3299, N3296, N536);
not NOT1 (N3300, N3293);
or OR2 (N3301, N3295, N1150);
buf BUF1 (N3302, N3301);
or OR4 (N3303, N3288, N2100, N1381, N2566);
not NOT1 (N3304, N3285);
nand NAND2 (N3305, N3279, N2165);
nand NAND2 (N3306, N3292, N85);
or OR2 (N3307, N3298, N259);
not NOT1 (N3308, N3302);
xor XOR2 (N3309, N3294, N1894);
or OR2 (N3310, N3304, N1952);
not NOT1 (N3311, N3290);
buf BUF1 (N3312, N3300);
xor XOR2 (N3313, N3307, N2463);
not NOT1 (N3314, N3313);
buf BUF1 (N3315, N3305);
or OR2 (N3316, N3315, N2958);
xor XOR2 (N3317, N3312, N580);
not NOT1 (N3318, N3317);
buf BUF1 (N3319, N3306);
xor XOR2 (N3320, N3316, N1222);
or OR3 (N3321, N3310, N1773, N183);
or OR3 (N3322, N3320, N3024, N2811);
and AND2 (N3323, N3322, N2608);
xor XOR2 (N3324, N3319, N3306);
nor NOR3 (N3325, N3324, N2098, N2367);
and AND3 (N3326, N3303, N1214, N2227);
or OR3 (N3327, N3326, N1868, N1289);
not NOT1 (N3328, N3318);
and AND3 (N3329, N3314, N102, N2081);
and AND3 (N3330, N3323, N1910, N891);
or OR4 (N3331, N3325, N1083, N837, N287);
not NOT1 (N3332, N3308);
nand NAND4 (N3333, N3327, N2290, N266, N719);
nand NAND3 (N3334, N3311, N3329, N2252);
and AND4 (N3335, N2495, N2371, N614, N3325);
or OR2 (N3336, N3299, N1605);
not NOT1 (N3337, N3334);
nor NOR2 (N3338, N3331, N3226);
xor XOR2 (N3339, N3338, N899);
or OR2 (N3340, N3339, N617);
buf BUF1 (N3341, N3321);
and AND4 (N3342, N3340, N125, N3206, N725);
nor NOR3 (N3343, N3333, N789, N2591);
not NOT1 (N3344, N3337);
not NOT1 (N3345, N3335);
nor NOR3 (N3346, N3342, N2278, N2583);
buf BUF1 (N3347, N3309);
nand NAND4 (N3348, N3343, N2785, N3065, N3294);
nand NAND3 (N3349, N3341, N2541, N2902);
or OR3 (N3350, N3347, N1628, N476);
nor NOR2 (N3351, N3350, N1565);
not NOT1 (N3352, N3330);
and AND4 (N3353, N3336, N1989, N1898, N1864);
nand NAND3 (N3354, N3346, N3251, N3095);
buf BUF1 (N3355, N3344);
buf BUF1 (N3356, N3328);
nand NAND4 (N3357, N3354, N1721, N1822, N199);
or OR3 (N3358, N3349, N1445, N224);
nor NOR2 (N3359, N3345, N104);
nand NAND4 (N3360, N3359, N1648, N2565, N3274);
xor XOR2 (N3361, N3357, N2448);
not NOT1 (N3362, N3332);
and AND4 (N3363, N3351, N1074, N2293, N3179);
and AND3 (N3364, N3361, N2040, N1307);
or OR3 (N3365, N3353, N1266, N644);
xor XOR2 (N3366, N3356, N3077);
and AND3 (N3367, N3365, N1394, N2027);
or OR3 (N3368, N3364, N1537, N1290);
nor NOR3 (N3369, N3368, N903, N3113);
buf BUF1 (N3370, N3369);
buf BUF1 (N3371, N3367);
nor NOR3 (N3372, N3362, N1500, N967);
and AND2 (N3373, N3355, N2782);
nor NOR4 (N3374, N3358, N3370, N2060, N2539);
nand NAND2 (N3375, N2235, N2012);
and AND4 (N3376, N3375, N2675, N2791, N3311);
or OR3 (N3377, N3372, N864, N1025);
nor NOR4 (N3378, N3348, N1464, N429, N1194);
or OR3 (N3379, N3378, N1042, N108);
nand NAND3 (N3380, N3373, N3020, N2252);
xor XOR2 (N3381, N3371, N2459);
not NOT1 (N3382, N3374);
nor NOR4 (N3383, N3363, N2604, N2066, N1586);
nor NOR3 (N3384, N3383, N687, N1548);
nand NAND2 (N3385, N3360, N2060);
not NOT1 (N3386, N3384);
nor NOR2 (N3387, N3382, N1996);
not NOT1 (N3388, N3352);
and AND4 (N3389, N3379, N1801, N1131, N1597);
nand NAND4 (N3390, N3381, N212, N1449, N2993);
buf BUF1 (N3391, N3388);
not NOT1 (N3392, N3389);
and AND2 (N3393, N3366, N882);
or OR4 (N3394, N3386, N3019, N1741, N1020);
xor XOR2 (N3395, N3376, N163);
or OR3 (N3396, N3392, N1358, N1627);
buf BUF1 (N3397, N3391);
not NOT1 (N3398, N3393);
and AND3 (N3399, N3396, N1032, N1745);
nand NAND2 (N3400, N3397, N2825);
nor NOR4 (N3401, N3398, N1346, N205, N1340);
and AND2 (N3402, N3401, N3142);
not NOT1 (N3403, N3387);
nand NAND4 (N3404, N3394, N2137, N1681, N1459);
or OR2 (N3405, N3399, N2316);
not NOT1 (N3406, N3380);
not NOT1 (N3407, N3395);
nand NAND3 (N3408, N3377, N86, N1500);
nand NAND2 (N3409, N3408, N1317);
nand NAND2 (N3410, N3403, N1822);
nor NOR2 (N3411, N3405, N1958);
not NOT1 (N3412, N3402);
not NOT1 (N3413, N3400);
nand NAND4 (N3414, N3409, N2107, N1557, N1152);
nand NAND3 (N3415, N3411, N2524, N244);
nor NOR4 (N3416, N3407, N1519, N288, N227);
nand NAND2 (N3417, N3390, N2800);
buf BUF1 (N3418, N3385);
buf BUF1 (N3419, N3414);
buf BUF1 (N3420, N3406);
nor NOR2 (N3421, N3415, N875);
nor NOR3 (N3422, N3417, N62, N387);
nor NOR4 (N3423, N3410, N612, N1544, N2373);
or OR4 (N3424, N3419, N2433, N2460, N169);
nand NAND4 (N3425, N3420, N620, N1579, N2285);
buf BUF1 (N3426, N3418);
nor NOR4 (N3427, N3422, N1544, N1018, N302);
nor NOR4 (N3428, N3412, N1150, N153, N2966);
and AND3 (N3429, N3423, N844, N3408);
not NOT1 (N3430, N3427);
nor NOR3 (N3431, N3425, N2916, N139);
not NOT1 (N3432, N3421);
xor XOR2 (N3433, N3430, N2228);
not NOT1 (N3434, N3426);
or OR3 (N3435, N3429, N897, N954);
buf BUF1 (N3436, N3432);
xor XOR2 (N3437, N3413, N2332);
nand NAND3 (N3438, N3437, N1858, N2953);
or OR3 (N3439, N3436, N727, N1265);
and AND2 (N3440, N3424, N1818);
buf BUF1 (N3441, N3439);
buf BUF1 (N3442, N3438);
xor XOR2 (N3443, N3433, N2477);
or OR4 (N3444, N3442, N2191, N960, N2656);
nand NAND4 (N3445, N3404, N778, N2286, N374);
buf BUF1 (N3446, N3431);
xor XOR2 (N3447, N3444, N1381);
and AND4 (N3448, N3435, N2667, N2058, N1491);
nor NOR4 (N3449, N3434, N845, N894, N2297);
or OR3 (N3450, N3449, N499, N3141);
xor XOR2 (N3451, N3440, N2096);
and AND2 (N3452, N3446, N3250);
buf BUF1 (N3453, N3452);
xor XOR2 (N3454, N3451, N1619);
xor XOR2 (N3455, N3453, N3132);
and AND2 (N3456, N3454, N74);
and AND4 (N3457, N3455, N3088, N2125, N2563);
nor NOR2 (N3458, N3457, N3000);
not NOT1 (N3459, N3456);
buf BUF1 (N3460, N3459);
and AND2 (N3461, N3460, N851);
and AND2 (N3462, N3428, N1960);
nor NOR3 (N3463, N3447, N1514, N1118);
buf BUF1 (N3464, N3461);
buf BUF1 (N3465, N3445);
buf BUF1 (N3466, N3465);
buf BUF1 (N3467, N3443);
not NOT1 (N3468, N3463);
or OR3 (N3469, N3448, N1648, N1965);
not NOT1 (N3470, N3466);
nand NAND3 (N3471, N3462, N1209, N1454);
and AND2 (N3472, N3471, N1448);
not NOT1 (N3473, N3469);
nand NAND2 (N3474, N3472, N509);
nand NAND4 (N3475, N3416, N917, N149, N111);
buf BUF1 (N3476, N3450);
nor NOR2 (N3477, N3473, N1394);
xor XOR2 (N3478, N3474, N1319);
nand NAND2 (N3479, N3441, N96);
buf BUF1 (N3480, N3467);
or OR3 (N3481, N3479, N1171, N1907);
or OR3 (N3482, N3470, N32, N722);
or OR2 (N3483, N3458, N1214);
buf BUF1 (N3484, N3468);
buf BUF1 (N3485, N3480);
buf BUF1 (N3486, N3484);
nand NAND2 (N3487, N3482, N3236);
nand NAND4 (N3488, N3485, N1091, N2595, N2235);
or OR2 (N3489, N3475, N1038);
nand NAND2 (N3490, N3487, N1746);
buf BUF1 (N3491, N3488);
or OR2 (N3492, N3476, N1480);
and AND2 (N3493, N3478, N1420);
or OR2 (N3494, N3490, N2563);
nor NOR3 (N3495, N3494, N230, N2802);
or OR2 (N3496, N3492, N1061);
not NOT1 (N3497, N3496);
not NOT1 (N3498, N3483);
xor XOR2 (N3499, N3464, N1138);
nand NAND3 (N3500, N3499, N447, N29);
or OR3 (N3501, N3500, N1039, N2621);
not NOT1 (N3502, N3486);
and AND3 (N3503, N3502, N1070, N1585);
buf BUF1 (N3504, N3477);
buf BUF1 (N3505, N3498);
xor XOR2 (N3506, N3493, N1889);
and AND2 (N3507, N3506, N1441);
xor XOR2 (N3508, N3505, N246);
not NOT1 (N3509, N3491);
or OR3 (N3510, N3503, N3409, N3398);
xor XOR2 (N3511, N3508, N1980);
nand NAND4 (N3512, N3501, N835, N1268, N959);
or OR4 (N3513, N3495, N188, N3480, N1221);
or OR4 (N3514, N3497, N2346, N1125, N1245);
and AND4 (N3515, N3514, N1109, N3466, N3035);
xor XOR2 (N3516, N3507, N243);
nand NAND2 (N3517, N3489, N2522);
buf BUF1 (N3518, N3513);
not NOT1 (N3519, N3481);
or OR2 (N3520, N3510, N1174);
nor NOR3 (N3521, N3504, N1968, N3095);
not NOT1 (N3522, N3511);
or OR3 (N3523, N3512, N862, N3243);
buf BUF1 (N3524, N3522);
or OR3 (N3525, N3520, N2484, N2205);
xor XOR2 (N3526, N3516, N1533);
and AND3 (N3527, N3521, N1385, N900);
or OR2 (N3528, N3527, N209);
buf BUF1 (N3529, N3528);
nand NAND3 (N3530, N3515, N1955, N284);
not NOT1 (N3531, N3518);
xor XOR2 (N3532, N3519, N2503);
or OR3 (N3533, N3524, N2210, N1077);
xor XOR2 (N3534, N3533, N2472);
buf BUF1 (N3535, N3526);
nand NAND4 (N3536, N3525, N3096, N2444, N2353);
and AND3 (N3537, N3529, N1075, N227);
not NOT1 (N3538, N3517);
or OR2 (N3539, N3531, N3070);
nand NAND4 (N3540, N3523, N1532, N577, N3457);
or OR3 (N3541, N3538, N2928, N2063);
buf BUF1 (N3542, N3540);
buf BUF1 (N3543, N3536);
xor XOR2 (N3544, N3543, N1910);
or OR3 (N3545, N3539, N2400, N2360);
buf BUF1 (N3546, N3535);
buf BUF1 (N3547, N3541);
and AND2 (N3548, N3534, N507);
nand NAND2 (N3549, N3544, N869);
xor XOR2 (N3550, N3546, N1398);
nand NAND3 (N3551, N3549, N996, N380);
buf BUF1 (N3552, N3509);
buf BUF1 (N3553, N3537);
or OR2 (N3554, N3545, N3232);
and AND3 (N3555, N3550, N816, N428);
and AND4 (N3556, N3553, N681, N621, N2206);
nand NAND2 (N3557, N3542, N2020);
nor NOR3 (N3558, N3530, N749, N1274);
buf BUF1 (N3559, N3548);
and AND3 (N3560, N3558, N2144, N3291);
nor NOR2 (N3561, N3555, N3211);
buf BUF1 (N3562, N3556);
nor NOR2 (N3563, N3562, N1859);
xor XOR2 (N3564, N3532, N3539);
not NOT1 (N3565, N3563);
nand NAND4 (N3566, N3547, N1930, N880, N2823);
not NOT1 (N3567, N3561);
nand NAND2 (N3568, N3559, N2529);
buf BUF1 (N3569, N3552);
xor XOR2 (N3570, N3551, N2062);
xor XOR2 (N3571, N3565, N609);
not NOT1 (N3572, N3554);
and AND4 (N3573, N3570, N2664, N3290, N1670);
nor NOR4 (N3574, N3557, N2540, N78, N2743);
buf BUF1 (N3575, N3571);
xor XOR2 (N3576, N3568, N47);
or OR3 (N3577, N3567, N15, N1364);
nand NAND4 (N3578, N3577, N3370, N575, N896);
buf BUF1 (N3579, N3578);
not NOT1 (N3580, N3560);
nor NOR4 (N3581, N3579, N1070, N623, N728);
not NOT1 (N3582, N3575);
nor NOR2 (N3583, N3580, N2629);
or OR2 (N3584, N3564, N1799);
buf BUF1 (N3585, N3581);
xor XOR2 (N3586, N3566, N2287);
buf BUF1 (N3587, N3576);
nor NOR2 (N3588, N3572, N3228);
xor XOR2 (N3589, N3583, N1320);
nor NOR3 (N3590, N3585, N1952, N1474);
nor NOR2 (N3591, N3590, N2213);
not NOT1 (N3592, N3582);
and AND3 (N3593, N3574, N1205, N968);
buf BUF1 (N3594, N3573);
xor XOR2 (N3595, N3589, N2699);
not NOT1 (N3596, N3588);
and AND2 (N3597, N3596, N2873);
nand NAND4 (N3598, N3592, N559, N1029, N2189);
and AND4 (N3599, N3597, N1550, N2550, N2399);
buf BUF1 (N3600, N3593);
buf BUF1 (N3601, N3569);
buf BUF1 (N3602, N3600);
buf BUF1 (N3603, N3587);
not NOT1 (N3604, N3598);
buf BUF1 (N3605, N3601);
and AND2 (N3606, N3595, N1563);
buf BUF1 (N3607, N3606);
nand NAND4 (N3608, N3604, N2869, N1789, N1707);
or OR4 (N3609, N3608, N1236, N91, N1796);
buf BUF1 (N3610, N3607);
buf BUF1 (N3611, N3594);
or OR3 (N3612, N3586, N1127, N675);
nor NOR2 (N3613, N3610, N3175);
nor NOR2 (N3614, N3611, N111);
or OR3 (N3615, N3603, N1527, N2146);
or OR4 (N3616, N3612, N1683, N191, N1342);
nor NOR2 (N3617, N3605, N1376);
or OR3 (N3618, N3614, N138, N2585);
buf BUF1 (N3619, N3599);
xor XOR2 (N3620, N3602, N2517);
xor XOR2 (N3621, N3619, N574);
not NOT1 (N3622, N3616);
nand NAND2 (N3623, N3617, N2715);
nand NAND4 (N3624, N3591, N1635, N2930, N2829);
and AND2 (N3625, N3622, N3149);
buf BUF1 (N3626, N3624);
nor NOR2 (N3627, N3613, N2118);
xor XOR2 (N3628, N3623, N1854);
xor XOR2 (N3629, N3628, N2687);
nand NAND3 (N3630, N3618, N3555, N1464);
buf BUF1 (N3631, N3609);
or OR2 (N3632, N3630, N2173);
buf BUF1 (N3633, N3584);
nand NAND2 (N3634, N3621, N3487);
nor NOR3 (N3635, N3632, N2367, N566);
xor XOR2 (N3636, N3620, N956);
and AND2 (N3637, N3633, N1590);
not NOT1 (N3638, N3625);
nor NOR2 (N3639, N3615, N2405);
not NOT1 (N3640, N3637);
not NOT1 (N3641, N3631);
and AND3 (N3642, N3635, N2110, N192);
nor NOR2 (N3643, N3636, N1214);
xor XOR2 (N3644, N3639, N295);
not NOT1 (N3645, N3638);
and AND4 (N3646, N3643, N1604, N3510, N2112);
and AND3 (N3647, N3629, N1150, N2681);
nor NOR3 (N3648, N3640, N2152, N915);
and AND3 (N3649, N3646, N1786, N2251);
xor XOR2 (N3650, N3642, N1232);
buf BUF1 (N3651, N3650);
buf BUF1 (N3652, N3634);
nor NOR2 (N3653, N3648, N3080);
nand NAND3 (N3654, N3651, N1559, N2464);
or OR2 (N3655, N3626, N2588);
not NOT1 (N3656, N3641);
nand NAND4 (N3657, N3627, N3028, N2361, N2983);
xor XOR2 (N3658, N3656, N2926);
not NOT1 (N3659, N3653);
not NOT1 (N3660, N3652);
not NOT1 (N3661, N3660);
nor NOR4 (N3662, N3645, N734, N3310, N2920);
not NOT1 (N3663, N3659);
buf BUF1 (N3664, N3649);
buf BUF1 (N3665, N3662);
nand NAND3 (N3666, N3644, N1339, N1531);
nand NAND2 (N3667, N3647, N1856);
xor XOR2 (N3668, N3664, N3535);
buf BUF1 (N3669, N3658);
xor XOR2 (N3670, N3669, N303);
buf BUF1 (N3671, N3667);
or OR2 (N3672, N3663, N1350);
and AND4 (N3673, N3670, N1970, N3161, N1906);
buf BUF1 (N3674, N3657);
nor NOR2 (N3675, N3674, N2011);
and AND3 (N3676, N3666, N468, N1622);
not NOT1 (N3677, N3672);
buf BUF1 (N3678, N3665);
buf BUF1 (N3679, N3661);
and AND2 (N3680, N3679, N2592);
nand NAND2 (N3681, N3668, N3235);
nand NAND2 (N3682, N3671, N3560);
buf BUF1 (N3683, N3681);
or OR2 (N3684, N3676, N2890);
buf BUF1 (N3685, N3655);
xor XOR2 (N3686, N3678, N11);
not NOT1 (N3687, N3685);
nor NOR4 (N3688, N3682, N3168, N2084, N1835);
not NOT1 (N3689, N3677);
xor XOR2 (N3690, N3684, N3432);
not NOT1 (N3691, N3683);
and AND2 (N3692, N3673, N1828);
xor XOR2 (N3693, N3690, N2827);
buf BUF1 (N3694, N3654);
xor XOR2 (N3695, N3693, N1186);
nor NOR3 (N3696, N3688, N804, N1218);
nand NAND2 (N3697, N3689, N1932);
nor NOR2 (N3698, N3695, N1486);
xor XOR2 (N3699, N3687, N2838);
nand NAND3 (N3700, N3680, N2935, N3132);
buf BUF1 (N3701, N3696);
not NOT1 (N3702, N3697);
or OR4 (N3703, N3694, N3657, N2545, N1956);
not NOT1 (N3704, N3686);
xor XOR2 (N3705, N3675, N2838);
not NOT1 (N3706, N3700);
nand NAND3 (N3707, N3701, N2681, N590);
xor XOR2 (N3708, N3699, N1441);
xor XOR2 (N3709, N3707, N2396);
and AND4 (N3710, N3706, N3696, N2670, N1909);
xor XOR2 (N3711, N3692, N3541);
or OR4 (N3712, N3691, N3261, N74, N125);
nor NOR2 (N3713, N3711, N1893);
buf BUF1 (N3714, N3704);
buf BUF1 (N3715, N3703);
nand NAND3 (N3716, N3702, N1630, N86);
buf BUF1 (N3717, N3712);
not NOT1 (N3718, N3698);
or OR3 (N3719, N3708, N1765, N914);
buf BUF1 (N3720, N3705);
nand NAND4 (N3721, N3719, N576, N2664, N1008);
nor NOR2 (N3722, N3715, N2592);
nand NAND4 (N3723, N3717, N3551, N1700, N1965);
buf BUF1 (N3724, N3723);
and AND2 (N3725, N3722, N1930);
nor NOR2 (N3726, N3716, N3692);
and AND4 (N3727, N3714, N325, N667, N2966);
and AND4 (N3728, N3718, N1985, N2386, N786);
buf BUF1 (N3729, N3709);
xor XOR2 (N3730, N3726, N1052);
xor XOR2 (N3731, N3725, N2063);
or OR2 (N3732, N3731, N1911);
xor XOR2 (N3733, N3729, N166);
or OR4 (N3734, N3727, N98, N440, N1976);
nand NAND2 (N3735, N3728, N3341);
xor XOR2 (N3736, N3721, N2000);
and AND4 (N3737, N3735, N1778, N55, N2784);
buf BUF1 (N3738, N3720);
xor XOR2 (N3739, N3737, N3531);
nor NOR2 (N3740, N3734, N2664);
and AND2 (N3741, N3740, N2976);
or OR2 (N3742, N3733, N2347);
and AND3 (N3743, N3739, N1038, N1706);
nor NOR4 (N3744, N3742, N2698, N1292, N1981);
and AND4 (N3745, N3736, N130, N289, N3648);
nor NOR2 (N3746, N3738, N3486);
and AND4 (N3747, N3732, N1155, N3431, N156);
nand NAND2 (N3748, N3741, N716);
or OR4 (N3749, N3710, N3638, N1856, N516);
and AND4 (N3750, N3747, N1377, N1450, N167);
xor XOR2 (N3751, N3744, N2098);
and AND3 (N3752, N3724, N138, N3313);
not NOT1 (N3753, N3749);
nor NOR2 (N3754, N3753, N2253);
xor XOR2 (N3755, N3746, N128);
nand NAND4 (N3756, N3751, N641, N764, N265);
not NOT1 (N3757, N3750);
nor NOR3 (N3758, N3713, N958, N1531);
nor NOR3 (N3759, N3754, N2910, N2015);
nand NAND2 (N3760, N3752, N2932);
buf BUF1 (N3761, N3757);
nand NAND2 (N3762, N3743, N2469);
not NOT1 (N3763, N3755);
nor NOR4 (N3764, N3745, N326, N2404, N3760);
nand NAND2 (N3765, N2824, N411);
xor XOR2 (N3766, N3764, N2430);
buf BUF1 (N3767, N3762);
nand NAND3 (N3768, N3759, N414, N955);
buf BUF1 (N3769, N3748);
nor NOR4 (N3770, N3761, N2924, N3322, N3617);
nand NAND4 (N3771, N3730, N2028, N653, N1523);
xor XOR2 (N3772, N3765, N2849);
not NOT1 (N3773, N3770);
buf BUF1 (N3774, N3763);
not NOT1 (N3775, N3774);
and AND3 (N3776, N3756, N1809, N1453);
xor XOR2 (N3777, N3771, N3016);
buf BUF1 (N3778, N3776);
xor XOR2 (N3779, N3768, N896);
nand NAND3 (N3780, N3767, N3264, N2746);
and AND4 (N3781, N3780, N725, N3768, N2576);
nor NOR3 (N3782, N3766, N2276, N1569);
buf BUF1 (N3783, N3781);
not NOT1 (N3784, N3772);
or OR3 (N3785, N3784, N1886, N1045);
not NOT1 (N3786, N3777);
xor XOR2 (N3787, N3786, N1833);
not NOT1 (N3788, N3785);
nand NAND3 (N3789, N3758, N998, N3472);
nand NAND2 (N3790, N3779, N1921);
nand NAND2 (N3791, N3787, N1307);
buf BUF1 (N3792, N3775);
and AND2 (N3793, N3789, N592);
or OR3 (N3794, N3783, N1371, N1455);
buf BUF1 (N3795, N3793);
and AND2 (N3796, N3788, N472);
or OR2 (N3797, N3791, N1489);
not NOT1 (N3798, N3790);
buf BUF1 (N3799, N3795);
or OR3 (N3800, N3798, N3215, N1951);
buf BUF1 (N3801, N3778);
and AND4 (N3802, N3797, N59, N2364, N659);
or OR3 (N3803, N3800, N1507, N1598);
or OR2 (N3804, N3769, N605);
nor NOR4 (N3805, N3773, N3187, N209, N1561);
xor XOR2 (N3806, N3805, N3443);
xor XOR2 (N3807, N3796, N1419);
buf BUF1 (N3808, N3803);
nor NOR4 (N3809, N3799, N3064, N2417, N752);
or OR3 (N3810, N3794, N3685, N604);
or OR2 (N3811, N3807, N1763);
nand NAND3 (N3812, N3810, N2123, N3618);
nor NOR2 (N3813, N3812, N3055);
xor XOR2 (N3814, N3782, N2376);
not NOT1 (N3815, N3801);
buf BUF1 (N3816, N3802);
and AND4 (N3817, N3816, N78, N2245, N802);
not NOT1 (N3818, N3815);
xor XOR2 (N3819, N3808, N353);
buf BUF1 (N3820, N3817);
buf BUF1 (N3821, N3813);
nand NAND2 (N3822, N3820, N672);
xor XOR2 (N3823, N3822, N3822);
nand NAND3 (N3824, N3819, N3054, N2257);
xor XOR2 (N3825, N3823, N2628);
nor NOR4 (N3826, N3824, N3161, N17, N3602);
xor XOR2 (N3827, N3814, N1240);
not NOT1 (N3828, N3821);
nand NAND3 (N3829, N3827, N3788, N3235);
xor XOR2 (N3830, N3828, N1912);
nand NAND4 (N3831, N3806, N2476, N3052, N1019);
or OR2 (N3832, N3818, N2357);
or OR2 (N3833, N3792, N3345);
nand NAND3 (N3834, N3825, N104, N2708);
or OR2 (N3835, N3831, N2485);
xor XOR2 (N3836, N3811, N587);
xor XOR2 (N3837, N3829, N2922);
nand NAND3 (N3838, N3830, N1816, N255);
nand NAND4 (N3839, N3809, N1431, N3489, N261);
and AND4 (N3840, N3836, N2702, N3390, N2318);
not NOT1 (N3841, N3826);
buf BUF1 (N3842, N3841);
nor NOR2 (N3843, N3837, N3380);
or OR3 (N3844, N3838, N2407, N162);
nor NOR4 (N3845, N3833, N1777, N1382, N3195);
or OR2 (N3846, N3843, N3833);
nor NOR4 (N3847, N3845, N2792, N1413, N584);
nand NAND2 (N3848, N3842, N1642);
not NOT1 (N3849, N3835);
nor NOR4 (N3850, N3847, N222, N1772, N506);
xor XOR2 (N3851, N3804, N2410);
xor XOR2 (N3852, N3848, N740);
buf BUF1 (N3853, N3832);
nand NAND2 (N3854, N3839, N2277);
not NOT1 (N3855, N3840);
nand NAND4 (N3856, N3855, N1720, N2268, N2040);
and AND4 (N3857, N3846, N306, N1358, N289);
nor NOR3 (N3858, N3834, N997, N313);
not NOT1 (N3859, N3854);
nand NAND3 (N3860, N3849, N138, N1763);
not NOT1 (N3861, N3857);
xor XOR2 (N3862, N3861, N1517);
and AND2 (N3863, N3858, N1986);
and AND4 (N3864, N3852, N1862, N3558, N2335);
nor NOR2 (N3865, N3856, N2813);
and AND3 (N3866, N3862, N339, N106);
buf BUF1 (N3867, N3864);
xor XOR2 (N3868, N3844, N1657);
nor NOR3 (N3869, N3860, N3651, N3672);
xor XOR2 (N3870, N3859, N1246);
and AND2 (N3871, N3853, N2006);
or OR4 (N3872, N3865, N2212, N424, N2186);
nor NOR4 (N3873, N3851, N1071, N652, N1554);
xor XOR2 (N3874, N3867, N613);
xor XOR2 (N3875, N3871, N102);
and AND4 (N3876, N3863, N1677, N1665, N2635);
nand NAND3 (N3877, N3869, N1029, N2340);
or OR2 (N3878, N3874, N2359);
nand NAND4 (N3879, N3875, N658, N2144, N2498);
nor NOR3 (N3880, N3872, N2145, N1506);
nor NOR2 (N3881, N3868, N3417);
nand NAND3 (N3882, N3850, N1146, N2261);
nor NOR3 (N3883, N3870, N1700, N62);
nand NAND3 (N3884, N3882, N778, N21);
xor XOR2 (N3885, N3877, N288);
or OR4 (N3886, N3876, N547, N2792, N1059);
nor NOR2 (N3887, N3881, N3061);
nor NOR2 (N3888, N3883, N1129);
not NOT1 (N3889, N3878);
nand NAND3 (N3890, N3880, N65, N2671);
xor XOR2 (N3891, N3885, N2621);
and AND3 (N3892, N3873, N1761, N2530);
buf BUF1 (N3893, N3892);
nor NOR3 (N3894, N3887, N3587, N189);
nor NOR2 (N3895, N3866, N2362);
or OR4 (N3896, N3895, N2144, N1005, N3001);
not NOT1 (N3897, N3884);
nand NAND3 (N3898, N3890, N673, N1530);
xor XOR2 (N3899, N3896, N2081);
xor XOR2 (N3900, N3891, N2165);
or OR2 (N3901, N3898, N2621);
nor NOR3 (N3902, N3899, N2169, N3611);
or OR4 (N3903, N3893, N3701, N1090, N3374);
not NOT1 (N3904, N3902);
nand NAND2 (N3905, N3904, N2120);
buf BUF1 (N3906, N3894);
nor NOR3 (N3907, N3906, N1152, N2760);
nor NOR4 (N3908, N3907, N2930, N1575, N1221);
xor XOR2 (N3909, N3901, N2059);
buf BUF1 (N3910, N3905);
buf BUF1 (N3911, N3908);
nor NOR2 (N3912, N3909, N1661);
buf BUF1 (N3913, N3886);
or OR4 (N3914, N3913, N761, N3561, N3837);
buf BUF1 (N3915, N3888);
xor XOR2 (N3916, N3910, N1653);
nor NOR2 (N3917, N3879, N2557);
nor NOR4 (N3918, N3915, N783, N645, N347);
xor XOR2 (N3919, N3903, N183);
and AND4 (N3920, N3912, N2364, N972, N2721);
xor XOR2 (N3921, N3920, N2666);
nor NOR2 (N3922, N3921, N3339);
or OR2 (N3923, N3922, N942);
not NOT1 (N3924, N3919);
and AND4 (N3925, N3889, N828, N3721, N1165);
and AND2 (N3926, N3900, N2098);
not NOT1 (N3927, N3917);
nor NOR4 (N3928, N3916, N2817, N1010, N1915);
buf BUF1 (N3929, N3897);
nand NAND2 (N3930, N3927, N1926);
and AND2 (N3931, N3911, N2903);
xor XOR2 (N3932, N3926, N1384);
nor NOR2 (N3933, N3923, N2150);
not NOT1 (N3934, N3929);
and AND2 (N3935, N3932, N560);
xor XOR2 (N3936, N3930, N2412);
nor NOR4 (N3937, N3936, N590, N741, N1675);
nand NAND2 (N3938, N3931, N560);
or OR2 (N3939, N3924, N1910);
not NOT1 (N3940, N3938);
and AND3 (N3941, N3939, N389, N400);
xor XOR2 (N3942, N3914, N3546);
not NOT1 (N3943, N3933);
buf BUF1 (N3944, N3940);
and AND2 (N3945, N3928, N3122);
nor NOR4 (N3946, N3925, N726, N937, N3849);
nand NAND2 (N3947, N3945, N3466);
nand NAND3 (N3948, N3947, N465, N1609);
or OR2 (N3949, N3934, N1860);
nor NOR2 (N3950, N3937, N3608);
not NOT1 (N3951, N3944);
buf BUF1 (N3952, N3943);
nor NOR3 (N3953, N3948, N3949, N1515);
and AND2 (N3954, N1445, N981);
buf BUF1 (N3955, N3946);
buf BUF1 (N3956, N3955);
nand NAND3 (N3957, N3941, N2797, N1223);
buf BUF1 (N3958, N3950);
and AND2 (N3959, N3954, N1497);
nor NOR3 (N3960, N3959, N3951, N2039);
nor NOR4 (N3961, N3089, N2188, N3673, N761);
not NOT1 (N3962, N3958);
xor XOR2 (N3963, N3957, N1371);
or OR4 (N3964, N3942, N404, N2455, N1092);
and AND2 (N3965, N3935, N1869);
and AND4 (N3966, N3964, N2750, N3288, N3908);
buf BUF1 (N3967, N3965);
nand NAND2 (N3968, N3953, N3525);
nand NAND2 (N3969, N3963, N3634);
buf BUF1 (N3970, N3918);
buf BUF1 (N3971, N3956);
or OR2 (N3972, N3961, N2952);
nor NOR4 (N3973, N3970, N1860, N3041, N707);
or OR4 (N3974, N3967, N2915, N3623, N3697);
nor NOR2 (N3975, N3968, N2775);
and AND4 (N3976, N3974, N101, N2803, N2722);
or OR3 (N3977, N3952, N447, N1422);
xor XOR2 (N3978, N3975, N981);
buf BUF1 (N3979, N3966);
xor XOR2 (N3980, N3977, N2777);
or OR3 (N3981, N3976, N125, N198);
xor XOR2 (N3982, N3971, N326);
and AND2 (N3983, N3978, N2441);
and AND2 (N3984, N3973, N324);
xor XOR2 (N3985, N3972, N1077);
nand NAND3 (N3986, N3979, N277, N2329);
or OR4 (N3987, N3962, N2298, N774, N2441);
nor NOR3 (N3988, N3986, N2461, N3122);
and AND2 (N3989, N3985, N3422);
or OR4 (N3990, N3989, N3816, N785, N2164);
nor NOR4 (N3991, N3990, N2206, N3089, N3659);
nand NAND4 (N3992, N3983, N2090, N3205, N3854);
buf BUF1 (N3993, N3980);
not NOT1 (N3994, N3981);
buf BUF1 (N3995, N3984);
or OR4 (N3996, N3960, N1440, N1244, N2810);
and AND4 (N3997, N3993, N2352, N669, N321);
and AND2 (N3998, N3997, N2399);
and AND3 (N3999, N3991, N3680, N3302);
and AND2 (N4000, N3988, N1135);
not NOT1 (N4001, N3995);
xor XOR2 (N4002, N3982, N2642);
not NOT1 (N4003, N3999);
xor XOR2 (N4004, N4000, N3162);
nor NOR2 (N4005, N4002, N2014);
nor NOR3 (N4006, N3996, N837, N3663);
and AND3 (N4007, N4003, N2042, N1934);
buf BUF1 (N4008, N3994);
or OR2 (N4009, N3992, N3422);
buf BUF1 (N4010, N3969);
xor XOR2 (N4011, N4006, N2133);
or OR2 (N4012, N3987, N1772);
not NOT1 (N4013, N4007);
nand NAND4 (N4014, N4011, N828, N2042, N1750);
buf BUF1 (N4015, N4014);
xor XOR2 (N4016, N4010, N893);
xor XOR2 (N4017, N4005, N2652);
or OR4 (N4018, N4015, N2283, N1571, N3012);
nand NAND4 (N4019, N4009, N473, N1744, N2394);
xor XOR2 (N4020, N3998, N1332);
nor NOR2 (N4021, N4016, N223);
nor NOR2 (N4022, N4012, N897);
nand NAND2 (N4023, N4017, N2566);
and AND2 (N4024, N4022, N246);
buf BUF1 (N4025, N4021);
nor NOR3 (N4026, N4024, N3904, N1309);
nor NOR2 (N4027, N4025, N1100);
nand NAND3 (N4028, N4004, N2732, N1886);
and AND2 (N4029, N4019, N2320);
nor NOR4 (N4030, N4008, N3655, N1584, N2950);
or OR3 (N4031, N4028, N1500, N3519);
not NOT1 (N4032, N4001);
nand NAND3 (N4033, N4026, N1199, N2313);
not NOT1 (N4034, N4018);
not NOT1 (N4035, N4027);
not NOT1 (N4036, N4034);
xor XOR2 (N4037, N4023, N3530);
and AND2 (N4038, N4020, N2303);
nor NOR3 (N4039, N4033, N2238, N2974);
nand NAND4 (N4040, N4031, N1645, N2877, N3978);
and AND4 (N4041, N4029, N3052, N3946, N1799);
or OR2 (N4042, N4013, N387);
nor NOR2 (N4043, N4030, N3589);
xor XOR2 (N4044, N4041, N3673);
nand NAND3 (N4045, N4036, N3780, N977);
buf BUF1 (N4046, N4038);
and AND3 (N4047, N4035, N3193, N3483);
or OR3 (N4048, N4037, N606, N381);
not NOT1 (N4049, N4039);
nand NAND2 (N4050, N4044, N725);
not NOT1 (N4051, N4040);
and AND2 (N4052, N4047, N3929);
or OR3 (N4053, N4042, N2373, N3587);
nand NAND2 (N4054, N4051, N2138);
xor XOR2 (N4055, N4050, N3536);
or OR4 (N4056, N4048, N4004, N1780, N1165);
and AND4 (N4057, N4032, N3981, N2175, N1924);
or OR3 (N4058, N4045, N2505, N216);
and AND2 (N4059, N4046, N946);
not NOT1 (N4060, N4056);
not NOT1 (N4061, N4052);
xor XOR2 (N4062, N4060, N706);
not NOT1 (N4063, N4054);
nor NOR3 (N4064, N4062, N2546, N367);
or OR4 (N4065, N4053, N1339, N3329, N2233);
or OR4 (N4066, N4058, N2310, N1865, N2992);
not NOT1 (N4067, N4059);
xor XOR2 (N4068, N4043, N1140);
nor NOR3 (N4069, N4065, N3194, N1350);
or OR3 (N4070, N4057, N1360, N2274);
and AND4 (N4071, N4067, N114, N1179, N956);
or OR2 (N4072, N4070, N1462);
or OR4 (N4073, N4061, N1348, N2146, N3200);
and AND2 (N4074, N4063, N3825);
nand NAND4 (N4075, N4066, N774, N1433, N3913);
nor NOR2 (N4076, N4064, N879);
buf BUF1 (N4077, N4075);
nor NOR2 (N4078, N4055, N3956);
nand NAND4 (N4079, N4077, N1477, N3123, N2706);
not NOT1 (N4080, N4078);
or OR4 (N4081, N4071, N3373, N624, N2456);
nor NOR2 (N4082, N4079, N484);
or OR4 (N4083, N4069, N2959, N1853, N963);
not NOT1 (N4084, N4080);
buf BUF1 (N4085, N4076);
xor XOR2 (N4086, N4083, N3233);
nor NOR2 (N4087, N4068, N3442);
or OR4 (N4088, N4049, N2914, N2258, N1645);
xor XOR2 (N4089, N4087, N1806);
and AND2 (N4090, N4074, N243);
buf BUF1 (N4091, N4085);
nor NOR4 (N4092, N4081, N1554, N3752, N1875);
not NOT1 (N4093, N4090);
nor NOR3 (N4094, N4089, N4034, N3933);
nor NOR3 (N4095, N4086, N1808, N2632);
and AND3 (N4096, N4084, N359, N920);
and AND4 (N4097, N4088, N797, N1666, N2880);
nand NAND3 (N4098, N4082, N3002, N3189);
nand NAND2 (N4099, N4091, N2394);
xor XOR2 (N4100, N4098, N721);
xor XOR2 (N4101, N4093, N1928);
nor NOR3 (N4102, N4096, N1607, N1330);
buf BUF1 (N4103, N4092);
buf BUF1 (N4104, N4099);
or OR4 (N4105, N4102, N2561, N286, N1584);
xor XOR2 (N4106, N4104, N3592);
nor NOR4 (N4107, N4101, N1139, N1959, N1903);
or OR4 (N4108, N4095, N261, N1715, N1776);
xor XOR2 (N4109, N4103, N2945);
nand NAND3 (N4110, N4108, N785, N1723);
xor XOR2 (N4111, N4107, N1322);
and AND2 (N4112, N4111, N2782);
xor XOR2 (N4113, N4094, N2039);
and AND2 (N4114, N4110, N1442);
and AND2 (N4115, N4113, N3758);
nor NOR4 (N4116, N4097, N1622, N871, N4009);
buf BUF1 (N4117, N4105);
nand NAND2 (N4118, N4100, N1859);
or OR3 (N4119, N4116, N798, N3301);
and AND3 (N4120, N4114, N1863, N2658);
or OR4 (N4121, N4117, N59, N3656, N490);
not NOT1 (N4122, N4072);
and AND2 (N4123, N4106, N3198);
xor XOR2 (N4124, N4120, N2095);
buf BUF1 (N4125, N4118);
nor NOR3 (N4126, N4115, N2960, N2368);
nand NAND2 (N4127, N4122, N947);
or OR2 (N4128, N4121, N3249);
not NOT1 (N4129, N4123);
buf BUF1 (N4130, N4129);
xor XOR2 (N4131, N4109, N2712);
xor XOR2 (N4132, N4128, N267);
nand NAND2 (N4133, N4119, N4117);
buf BUF1 (N4134, N4073);
nor NOR2 (N4135, N4112, N1160);
nand NAND3 (N4136, N4132, N2064, N2178);
nor NOR2 (N4137, N4125, N515);
xor XOR2 (N4138, N4133, N1505);
buf BUF1 (N4139, N4131);
nor NOR2 (N4140, N4136, N3500);
nand NAND4 (N4141, N4127, N3856, N3910, N3249);
and AND3 (N4142, N4139, N2009, N450);
xor XOR2 (N4143, N4141, N1921);
or OR2 (N4144, N4130, N2813);
or OR3 (N4145, N4144, N1049, N522);
not NOT1 (N4146, N4135);
and AND2 (N4147, N4142, N1420);
or OR4 (N4148, N4145, N1425, N1950, N119);
nor NOR3 (N4149, N4124, N3264, N1293);
nand NAND4 (N4150, N4140, N2017, N516, N1002);
nand NAND2 (N4151, N4146, N3700);
not NOT1 (N4152, N4137);
nand NAND4 (N4153, N4126, N396, N1640, N2882);
and AND3 (N4154, N4147, N614, N989);
xor XOR2 (N4155, N4138, N2986);
and AND2 (N4156, N4148, N462);
buf BUF1 (N4157, N4151);
not NOT1 (N4158, N4143);
not NOT1 (N4159, N4156);
and AND3 (N4160, N4155, N1046, N4073);
xor XOR2 (N4161, N4157, N2460);
xor XOR2 (N4162, N4152, N3868);
not NOT1 (N4163, N4153);
buf BUF1 (N4164, N4154);
not NOT1 (N4165, N4164);
buf BUF1 (N4166, N4161);
and AND2 (N4167, N4163, N1759);
nand NAND3 (N4168, N4150, N2533, N3190);
and AND3 (N4169, N4167, N2147, N1484);
and AND2 (N4170, N4168, N1411);
xor XOR2 (N4171, N4162, N442);
not NOT1 (N4172, N4170);
xor XOR2 (N4173, N4134, N69);
not NOT1 (N4174, N4169);
and AND3 (N4175, N4159, N815, N596);
nand NAND4 (N4176, N4149, N1043, N1518, N2193);
or OR3 (N4177, N4172, N3705, N1182);
or OR3 (N4178, N4174, N1923, N3645);
or OR2 (N4179, N4178, N1588);
and AND3 (N4180, N4177, N3014, N2413);
or OR4 (N4181, N4166, N859, N2047, N1559);
buf BUF1 (N4182, N4165);
xor XOR2 (N4183, N4175, N1293);
xor XOR2 (N4184, N4171, N1765);
xor XOR2 (N4185, N4181, N1085);
nand NAND3 (N4186, N4183, N2552, N2670);
xor XOR2 (N4187, N4185, N3959);
or OR2 (N4188, N4158, N2276);
xor XOR2 (N4189, N4160, N587);
or OR3 (N4190, N4187, N2536, N1699);
not NOT1 (N4191, N4173);
buf BUF1 (N4192, N4176);
nor NOR3 (N4193, N4179, N853, N2033);
not NOT1 (N4194, N4188);
xor XOR2 (N4195, N4180, N3455);
not NOT1 (N4196, N4193);
xor XOR2 (N4197, N4190, N2474);
nand NAND2 (N4198, N4182, N4105);
or OR2 (N4199, N4184, N1929);
xor XOR2 (N4200, N4192, N3753);
or OR2 (N4201, N4200, N182);
and AND2 (N4202, N4199, N1585);
nand NAND2 (N4203, N4195, N1648);
nand NAND2 (N4204, N4197, N506);
or OR4 (N4205, N4191, N1873, N1843, N48);
and AND4 (N4206, N4198, N551, N2952, N3925);
nand NAND3 (N4207, N4194, N3919, N1437);
nor NOR4 (N4208, N4202, N3867, N2985, N1016);
xor XOR2 (N4209, N4206, N3623);
xor XOR2 (N4210, N4186, N1018);
nor NOR4 (N4211, N4203, N2748, N269, N2313);
and AND2 (N4212, N4208, N1438);
buf BUF1 (N4213, N4209);
not NOT1 (N4214, N4211);
nor NOR3 (N4215, N4207, N2001, N4003);
or OR3 (N4216, N4205, N447, N2098);
xor XOR2 (N4217, N4210, N807);
buf BUF1 (N4218, N4204);
buf BUF1 (N4219, N4216);
or OR4 (N4220, N4213, N1393, N600, N2462);
or OR4 (N4221, N4189, N1632, N1518, N3484);
not NOT1 (N4222, N4201);
buf BUF1 (N4223, N4218);
nor NOR2 (N4224, N4196, N317);
or OR3 (N4225, N4217, N1489, N1906);
buf BUF1 (N4226, N4222);
not NOT1 (N4227, N4215);
and AND3 (N4228, N4212, N3186, N1362);
nand NAND4 (N4229, N4219, N119, N1603, N122);
xor XOR2 (N4230, N4224, N3124);
buf BUF1 (N4231, N4229);
nand NAND2 (N4232, N4227, N801);
nand NAND2 (N4233, N4230, N773);
not NOT1 (N4234, N4220);
nor NOR4 (N4235, N4232, N3942, N3064, N2114);
or OR4 (N4236, N4234, N978, N544, N1335);
nor NOR2 (N4237, N4221, N2282);
nor NOR4 (N4238, N4233, N1971, N1417, N4150);
or OR2 (N4239, N4231, N29);
nand NAND3 (N4240, N4237, N2071, N603);
buf BUF1 (N4241, N4238);
or OR3 (N4242, N4241, N3436, N3796);
buf BUF1 (N4243, N4223);
xor XOR2 (N4244, N4214, N2447);
nor NOR3 (N4245, N4240, N1374, N382);
not NOT1 (N4246, N4236);
or OR2 (N4247, N4244, N1902);
nand NAND4 (N4248, N4239, N3210, N1914, N1665);
nand NAND2 (N4249, N4245, N1206);
nor NOR2 (N4250, N4249, N2315);
nand NAND3 (N4251, N4247, N306, N450);
xor XOR2 (N4252, N4248, N2502);
nor NOR4 (N4253, N4226, N1829, N3110, N899);
not NOT1 (N4254, N4225);
and AND4 (N4255, N4250, N2644, N148, N1277);
nor NOR2 (N4256, N4254, N3232);
buf BUF1 (N4257, N4242);
buf BUF1 (N4258, N4256);
not NOT1 (N4259, N4258);
nor NOR4 (N4260, N4252, N1518, N178, N4079);
buf BUF1 (N4261, N4257);
or OR3 (N4262, N4246, N3583, N1529);
and AND4 (N4263, N4260, N3132, N2349, N2425);
buf BUF1 (N4264, N4255);
nand NAND2 (N4265, N4235, N3732);
not NOT1 (N4266, N4262);
and AND4 (N4267, N4251, N3209, N1797, N2589);
not NOT1 (N4268, N4261);
nand NAND4 (N4269, N4268, N196, N1940, N1425);
nand NAND3 (N4270, N4269, N1174, N783);
and AND4 (N4271, N4228, N1832, N4015, N3019);
or OR4 (N4272, N4266, N1916, N2343, N3874);
or OR3 (N4273, N4243, N3654, N4180);
nand NAND2 (N4274, N4267, N261);
xor XOR2 (N4275, N4265, N1198);
buf BUF1 (N4276, N4275);
not NOT1 (N4277, N4274);
and AND3 (N4278, N4276, N1650, N2025);
or OR2 (N4279, N4253, N2557);
not NOT1 (N4280, N4278);
nand NAND4 (N4281, N4264, N1992, N810, N1291);
not NOT1 (N4282, N4259);
nand NAND3 (N4283, N4277, N115, N282);
nand NAND3 (N4284, N4279, N390, N3815);
not NOT1 (N4285, N4280);
and AND2 (N4286, N4272, N2494);
not NOT1 (N4287, N4263);
or OR4 (N4288, N4285, N3376, N4156, N2600);
not NOT1 (N4289, N4287);
not NOT1 (N4290, N4270);
xor XOR2 (N4291, N4271, N3876);
not NOT1 (N4292, N4286);
and AND4 (N4293, N4288, N3552, N3630, N2275);
nor NOR4 (N4294, N4281, N4221, N1856, N3325);
not NOT1 (N4295, N4292);
nand NAND3 (N4296, N4283, N912, N735);
nand NAND3 (N4297, N4284, N3214, N2636);
buf BUF1 (N4298, N4290);
not NOT1 (N4299, N4294);
not NOT1 (N4300, N4293);
nand NAND4 (N4301, N4289, N2981, N624, N1957);
nor NOR4 (N4302, N4299, N2073, N3134, N3282);
not NOT1 (N4303, N4302);
nor NOR2 (N4304, N4303, N2365);
and AND4 (N4305, N4296, N2354, N3113, N3040);
and AND3 (N4306, N4297, N862, N3489);
nor NOR2 (N4307, N4304, N1632);
not NOT1 (N4308, N4307);
nand NAND4 (N4309, N4305, N987, N2069, N843);
or OR3 (N4310, N4273, N442, N3818);
and AND2 (N4311, N4309, N509);
nor NOR2 (N4312, N4308, N1024);
nand NAND4 (N4313, N4295, N211, N406, N4114);
nor NOR2 (N4314, N4282, N346);
not NOT1 (N4315, N4301);
and AND3 (N4316, N4311, N3785, N4151);
xor XOR2 (N4317, N4298, N682);
nand NAND4 (N4318, N4300, N3707, N3742, N2019);
buf BUF1 (N4319, N4317);
nand NAND2 (N4320, N4310, N724);
or OR4 (N4321, N4314, N2049, N2209, N2284);
nor NOR2 (N4322, N4291, N2037);
nand NAND2 (N4323, N4313, N518);
xor XOR2 (N4324, N4322, N4309);
buf BUF1 (N4325, N4316);
and AND4 (N4326, N4318, N3267, N549, N496);
nand NAND3 (N4327, N4321, N1831, N830);
nor NOR2 (N4328, N4312, N2464);
buf BUF1 (N4329, N4324);
xor XOR2 (N4330, N4326, N588);
and AND4 (N4331, N4319, N3580, N3581, N43);
and AND4 (N4332, N4330, N4111, N3618, N1663);
and AND4 (N4333, N4325, N2950, N3410, N2613);
not NOT1 (N4334, N4323);
not NOT1 (N4335, N4315);
and AND2 (N4336, N4328, N1703);
not NOT1 (N4337, N4329);
nor NOR3 (N4338, N4335, N33, N4128);
xor XOR2 (N4339, N4332, N4316);
or OR2 (N4340, N4334, N3301);
not NOT1 (N4341, N4338);
and AND2 (N4342, N4320, N2119);
nor NOR3 (N4343, N4342, N4254, N1999);
or OR4 (N4344, N4339, N1959, N1034, N4162);
xor XOR2 (N4345, N4331, N1350);
not NOT1 (N4346, N4336);
or OR2 (N4347, N4337, N652);
xor XOR2 (N4348, N4344, N2147);
not NOT1 (N4349, N4327);
nor NOR4 (N4350, N4306, N861, N2663, N633);
not NOT1 (N4351, N4341);
and AND2 (N4352, N4351, N1575);
not NOT1 (N4353, N4348);
or OR4 (N4354, N4347, N1983, N2164, N3897);
or OR2 (N4355, N4343, N172);
xor XOR2 (N4356, N4354, N3283);
nor NOR3 (N4357, N4345, N1357, N532);
and AND4 (N4358, N4355, N4249, N1835, N4028);
nor NOR3 (N4359, N4350, N314, N3642);
not NOT1 (N4360, N4333);
not NOT1 (N4361, N4340);
buf BUF1 (N4362, N4352);
nand NAND4 (N4363, N4361, N2895, N1482, N3495);
not NOT1 (N4364, N4360);
buf BUF1 (N4365, N4362);
nand NAND2 (N4366, N4359, N45);
xor XOR2 (N4367, N4365, N3236);
nand NAND3 (N4368, N4346, N2917, N3849);
xor XOR2 (N4369, N4368, N4054);
buf BUF1 (N4370, N4353);
buf BUF1 (N4371, N4357);
buf BUF1 (N4372, N4370);
nor NOR3 (N4373, N4363, N3458, N1966);
buf BUF1 (N4374, N4373);
buf BUF1 (N4375, N4349);
not NOT1 (N4376, N4367);
buf BUF1 (N4377, N4375);
buf BUF1 (N4378, N4374);
and AND3 (N4379, N4376, N2047, N107);
xor XOR2 (N4380, N4372, N4092);
or OR3 (N4381, N4364, N3435, N1148);
or OR4 (N4382, N4381, N373, N2403, N3333);
and AND3 (N4383, N4356, N877, N1151);
buf BUF1 (N4384, N4369);
buf BUF1 (N4385, N4358);
nor NOR3 (N4386, N4371, N3348, N1413);
and AND4 (N4387, N4382, N2244, N1679, N3152);
or OR3 (N4388, N4386, N296, N2433);
nor NOR4 (N4389, N4380, N602, N2294, N1266);
buf BUF1 (N4390, N4379);
buf BUF1 (N4391, N4390);
nand NAND3 (N4392, N4385, N164, N1888);
nand NAND2 (N4393, N4388, N287);
and AND4 (N4394, N4366, N3672, N26, N220);
buf BUF1 (N4395, N4389);
xor XOR2 (N4396, N4393, N1104);
buf BUF1 (N4397, N4377);
nor NOR2 (N4398, N4378, N3767);
buf BUF1 (N4399, N4398);
xor XOR2 (N4400, N4396, N1941);
nand NAND3 (N4401, N4387, N1291, N3430);
buf BUF1 (N4402, N4400);
not NOT1 (N4403, N4395);
or OR4 (N4404, N4391, N2511, N3176, N3875);
buf BUF1 (N4405, N4383);
buf BUF1 (N4406, N4405);
nand NAND3 (N4407, N4403, N929, N1592);
buf BUF1 (N4408, N4402);
nor NOR3 (N4409, N4384, N3602, N287);
not NOT1 (N4410, N4407);
nand NAND2 (N4411, N4401, N3393);
buf BUF1 (N4412, N4394);
nor NOR2 (N4413, N4399, N3456);
not NOT1 (N4414, N4409);
not NOT1 (N4415, N4397);
not NOT1 (N4416, N4404);
or OR2 (N4417, N4406, N180);
nand NAND3 (N4418, N4411, N4248, N971);
nand NAND4 (N4419, N4412, N602, N4216, N4097);
buf BUF1 (N4420, N4413);
and AND3 (N4421, N4418, N4293, N4333);
xor XOR2 (N4422, N4392, N2050);
buf BUF1 (N4423, N4415);
buf BUF1 (N4424, N4417);
nand NAND3 (N4425, N4416, N2826, N2095);
or OR2 (N4426, N4408, N3498);
and AND2 (N4427, N4424, N4120);
not NOT1 (N4428, N4423);
or OR3 (N4429, N4427, N3584, N2344);
nand NAND3 (N4430, N4428, N2393, N2208);
buf BUF1 (N4431, N4429);
nand NAND2 (N4432, N4422, N3966);
nand NAND3 (N4433, N4421, N3853, N1511);
not NOT1 (N4434, N4419);
xor XOR2 (N4435, N4433, N1684);
or OR3 (N4436, N4420, N1805, N1496);
or OR4 (N4437, N4410, N3514, N2060, N2897);
nor NOR2 (N4438, N4425, N3857);
and AND2 (N4439, N4435, N2447);
buf BUF1 (N4440, N4414);
buf BUF1 (N4441, N4434);
and AND3 (N4442, N4436, N1027, N1616);
nand NAND4 (N4443, N4442, N2194, N1074, N1191);
or OR4 (N4444, N4432, N2358, N2848, N1103);
not NOT1 (N4445, N4444);
not NOT1 (N4446, N4445);
nor NOR2 (N4447, N4439, N729);
xor XOR2 (N4448, N4441, N1251);
or OR2 (N4449, N4437, N3285);
not NOT1 (N4450, N4446);
nand NAND3 (N4451, N4448, N3383, N3725);
not NOT1 (N4452, N4443);
and AND4 (N4453, N4452, N4371, N878, N2779);
nand NAND3 (N4454, N4426, N3348, N4);
buf BUF1 (N4455, N4454);
and AND4 (N4456, N4447, N1280, N2033, N3648);
nor NOR3 (N4457, N4440, N1570, N1967);
buf BUF1 (N4458, N4453);
or OR2 (N4459, N4451, N1993);
nor NOR3 (N4460, N4455, N727, N3118);
or OR4 (N4461, N4438, N2436, N1028, N1126);
xor XOR2 (N4462, N4459, N158);
or OR2 (N4463, N4449, N1566);
nand NAND2 (N4464, N4430, N3595);
not NOT1 (N4465, N4431);
buf BUF1 (N4466, N4457);
not NOT1 (N4467, N4464);
or OR2 (N4468, N4456, N3774);
or OR3 (N4469, N4450, N3563, N2213);
buf BUF1 (N4470, N4461);
xor XOR2 (N4471, N4469, N135);
buf BUF1 (N4472, N4471);
xor XOR2 (N4473, N4460, N1301);
or OR4 (N4474, N4468, N587, N7, N3845);
not NOT1 (N4475, N4463);
nand NAND2 (N4476, N4472, N2570);
or OR2 (N4477, N4476, N1006);
buf BUF1 (N4478, N4465);
xor XOR2 (N4479, N4467, N1702);
or OR4 (N4480, N4474, N1016, N2153, N3492);
or OR4 (N4481, N4478, N3584, N1069, N468);
or OR3 (N4482, N4479, N1884, N2750);
not NOT1 (N4483, N4480);
nor NOR3 (N4484, N4462, N3541, N3004);
nor NOR2 (N4485, N4470, N4115);
nand NAND4 (N4486, N4481, N4215, N2034, N397);
and AND4 (N4487, N4483, N3322, N1970, N1883);
or OR3 (N4488, N4484, N4046, N3699);
and AND4 (N4489, N4482, N2576, N2484, N3088);
or OR3 (N4490, N4487, N1336, N183);
not NOT1 (N4491, N4475);
or OR3 (N4492, N4473, N2703, N721);
or OR4 (N4493, N4491, N3152, N442, N706);
buf BUF1 (N4494, N4466);
not NOT1 (N4495, N4494);
buf BUF1 (N4496, N4488);
buf BUF1 (N4497, N4489);
nor NOR3 (N4498, N4458, N213, N3671);
or OR3 (N4499, N4490, N2321, N109);
or OR2 (N4500, N4495, N3775);
or OR3 (N4501, N4498, N1495, N1912);
nor NOR4 (N4502, N4493, N484, N742, N2256);
buf BUF1 (N4503, N4477);
and AND4 (N4504, N4496, N3686, N2979, N3001);
nor NOR2 (N4505, N4499, N3473);
nand NAND2 (N4506, N4504, N3428);
or OR2 (N4507, N4502, N2544);
xor XOR2 (N4508, N4507, N3781);
nor NOR2 (N4509, N4506, N1872);
xor XOR2 (N4510, N4505, N3779);
or OR3 (N4511, N4508, N1504, N2043);
buf BUF1 (N4512, N4503);
and AND3 (N4513, N4485, N319, N751);
buf BUF1 (N4514, N4513);
buf BUF1 (N4515, N4509);
and AND4 (N4516, N4514, N491, N3481, N24);
and AND2 (N4517, N4511, N2330);
nand NAND3 (N4518, N4510, N3042, N2381);
not NOT1 (N4519, N4500);
nor NOR4 (N4520, N4492, N587, N3440, N4262);
and AND2 (N4521, N4518, N404);
nor NOR3 (N4522, N4512, N2560, N4323);
and AND2 (N4523, N4522, N493);
xor XOR2 (N4524, N4516, N3490);
or OR2 (N4525, N4520, N2388);
xor XOR2 (N4526, N4525, N2782);
not NOT1 (N4527, N4501);
nor NOR4 (N4528, N4519, N587, N3844, N1336);
not NOT1 (N4529, N4523);
xor XOR2 (N4530, N4527, N553);
nand NAND3 (N4531, N4529, N926, N3216);
and AND2 (N4532, N4486, N1794);
not NOT1 (N4533, N4530);
or OR2 (N4534, N4533, N2229);
buf BUF1 (N4535, N4515);
xor XOR2 (N4536, N4517, N2795);
and AND2 (N4537, N4526, N138);
not NOT1 (N4538, N4528);
nor NOR4 (N4539, N4497, N504, N674, N2188);
or OR4 (N4540, N4536, N1381, N4526, N526);
not NOT1 (N4541, N4521);
xor XOR2 (N4542, N4534, N1073);
and AND2 (N4543, N4538, N1075);
not NOT1 (N4544, N4540);
or OR4 (N4545, N4542, N4333, N2369, N4259);
or OR4 (N4546, N4524, N2932, N3204, N168);
nand NAND2 (N4547, N4532, N2478);
nand NAND3 (N4548, N4545, N2189, N222);
nor NOR4 (N4549, N4546, N3445, N3162, N4372);
or OR4 (N4550, N4549, N340, N2962, N4021);
nand NAND3 (N4551, N4548, N1925, N2488);
and AND3 (N4552, N4550, N2489, N1134);
nand NAND4 (N4553, N4539, N2264, N3207, N4054);
buf BUF1 (N4554, N4551);
and AND4 (N4555, N4547, N863, N1, N1857);
xor XOR2 (N4556, N4552, N1465);
and AND4 (N4557, N4535, N699, N1542, N3090);
nor NOR4 (N4558, N4541, N3524, N1308, N4220);
not NOT1 (N4559, N4553);
and AND2 (N4560, N4543, N1968);
or OR2 (N4561, N4560, N1553);
xor XOR2 (N4562, N4556, N4296);
and AND3 (N4563, N4531, N3579, N298);
xor XOR2 (N4564, N4554, N764);
buf BUF1 (N4565, N4557);
or OR4 (N4566, N4559, N449, N2123, N3894);
buf BUF1 (N4567, N4555);
not NOT1 (N4568, N4565);
and AND3 (N4569, N4544, N678, N4037);
and AND2 (N4570, N4561, N395);
nand NAND4 (N4571, N4568, N1455, N2369, N1991);
not NOT1 (N4572, N4569);
or OR3 (N4573, N4571, N2604, N3060);
nor NOR2 (N4574, N4572, N846);
nor NOR3 (N4575, N4558, N3712, N389);
not NOT1 (N4576, N4566);
not NOT1 (N4577, N4576);
nor NOR3 (N4578, N4575, N2400, N2865);
not NOT1 (N4579, N4564);
nand NAND3 (N4580, N4574, N4466, N2176);
nor NOR3 (N4581, N4563, N3725, N448);
or OR4 (N4582, N4573, N1834, N752, N3764);
nor NOR4 (N4583, N4562, N623, N4187, N1674);
and AND4 (N4584, N4580, N2419, N3668, N15);
or OR4 (N4585, N4584, N1303, N1563, N1743);
nand NAND4 (N4586, N4537, N1039, N583, N3172);
not NOT1 (N4587, N4577);
or OR2 (N4588, N4585, N1663);
nor NOR2 (N4589, N4587, N1902);
and AND2 (N4590, N4579, N1976);
nand NAND2 (N4591, N4590, N1275);
nand NAND3 (N4592, N4586, N3933, N3960);
xor XOR2 (N4593, N4570, N2108);
not NOT1 (N4594, N4567);
nand NAND3 (N4595, N4593, N547, N966);
nand NAND3 (N4596, N4582, N54, N4480);
or OR2 (N4597, N4592, N4040);
nand NAND2 (N4598, N4581, N1094);
nor NOR3 (N4599, N4594, N3879, N3915);
buf BUF1 (N4600, N4589);
or OR2 (N4601, N4591, N2859);
or OR2 (N4602, N4597, N1803);
nor NOR3 (N4603, N4595, N2417, N3184);
not NOT1 (N4604, N4596);
or OR3 (N4605, N4603, N825, N4345);
nand NAND4 (N4606, N4578, N2673, N2614, N19);
xor XOR2 (N4607, N4598, N3814);
and AND3 (N4608, N4600, N2101, N928);
nor NOR2 (N4609, N4604, N2639);
nand NAND4 (N4610, N4599, N1987, N252, N1376);
nand NAND3 (N4611, N4609, N1011, N2847);
buf BUF1 (N4612, N4602);
buf BUF1 (N4613, N4588);
and AND2 (N4614, N4612, N360);
not NOT1 (N4615, N4610);
or OR2 (N4616, N4608, N1299);
xor XOR2 (N4617, N4583, N806);
nor NOR3 (N4618, N4601, N1047, N2285);
not NOT1 (N4619, N4615);
nor NOR3 (N4620, N4611, N264, N2550);
and AND3 (N4621, N4619, N1766, N3341);
and AND2 (N4622, N4613, N3447);
nor NOR4 (N4623, N4618, N1559, N2572, N3360);
nand NAND2 (N4624, N4617, N1190);
nand NAND4 (N4625, N4616, N842, N4225, N4534);
xor XOR2 (N4626, N4623, N158);
or OR3 (N4627, N4607, N2094, N2818);
nor NOR4 (N4628, N4624, N636, N307, N4566);
or OR2 (N4629, N4606, N1206);
and AND4 (N4630, N4626, N372, N250, N566);
nor NOR4 (N4631, N4630, N4496, N2178, N3198);
nand NAND3 (N4632, N4631, N3928, N1541);
not NOT1 (N4633, N4620);
xor XOR2 (N4634, N4605, N298);
xor XOR2 (N4635, N4614, N1956);
or OR3 (N4636, N4628, N511, N2158);
not NOT1 (N4637, N4636);
and AND3 (N4638, N4621, N1708, N3702);
or OR4 (N4639, N4622, N4176, N4463, N3731);
and AND2 (N4640, N4635, N1356);
or OR4 (N4641, N4627, N660, N3430, N4166);
and AND4 (N4642, N4637, N2772, N878, N4579);
and AND2 (N4643, N4632, N1684);
xor XOR2 (N4644, N4629, N1017);
xor XOR2 (N4645, N4640, N4618);
xor XOR2 (N4646, N4634, N2471);
and AND2 (N4647, N4641, N2127);
buf BUF1 (N4648, N4646);
or OR4 (N4649, N4639, N3494, N512, N1062);
not NOT1 (N4650, N4645);
or OR2 (N4651, N4648, N4262);
xor XOR2 (N4652, N4642, N65);
nor NOR4 (N4653, N4643, N400, N2736, N1576);
or OR3 (N4654, N4652, N119, N784);
nor NOR2 (N4655, N4650, N150);
buf BUF1 (N4656, N4625);
and AND3 (N4657, N4653, N2324, N3471);
nand NAND4 (N4658, N4638, N3075, N414, N809);
buf BUF1 (N4659, N4658);
not NOT1 (N4660, N4654);
and AND4 (N4661, N4660, N1707, N379, N1436);
not NOT1 (N4662, N4657);
xor XOR2 (N4663, N4662, N3257);
buf BUF1 (N4664, N4655);
nor NOR2 (N4665, N4647, N3236);
not NOT1 (N4666, N4644);
xor XOR2 (N4667, N4666, N3257);
and AND4 (N4668, N4633, N429, N1497, N3105);
not NOT1 (N4669, N4661);
buf BUF1 (N4670, N4656);
nor NOR3 (N4671, N4664, N3684, N2368);
nand NAND3 (N4672, N4663, N2663, N1068);
nand NAND3 (N4673, N4667, N230, N3306);
not NOT1 (N4674, N4671);
buf BUF1 (N4675, N4674);
nand NAND4 (N4676, N4669, N483, N2966, N232);
xor XOR2 (N4677, N4649, N4291);
and AND2 (N4678, N4659, N1118);
nor NOR2 (N4679, N4672, N2651);
buf BUF1 (N4680, N4679);
xor XOR2 (N4681, N4673, N2068);
xor XOR2 (N4682, N4676, N3610);
nand NAND4 (N4683, N4651, N998, N1069, N1658);
xor XOR2 (N4684, N4680, N4344);
nor NOR3 (N4685, N4684, N2546, N3308);
xor XOR2 (N4686, N4668, N2267);
nor NOR2 (N4687, N4685, N3403);
nor NOR4 (N4688, N4665, N2987, N4427, N1455);
nor NOR2 (N4689, N4687, N2423);
or OR2 (N4690, N4688, N615);
and AND3 (N4691, N4690, N1288, N2054);
buf BUF1 (N4692, N4691);
nand NAND3 (N4693, N4686, N2934, N3183);
xor XOR2 (N4694, N4670, N232);
and AND4 (N4695, N4677, N2250, N679, N4439);
not NOT1 (N4696, N4692);
nand NAND2 (N4697, N4689, N3318);
nand NAND2 (N4698, N4678, N1811);
nor NOR2 (N4699, N4693, N4041);
and AND3 (N4700, N4694, N230, N3034);
or OR4 (N4701, N4675, N817, N129, N2592);
xor XOR2 (N4702, N4695, N486);
and AND4 (N4703, N4700, N2813, N4146, N4324);
and AND4 (N4704, N4697, N3901, N3233, N2525);
nand NAND4 (N4705, N4682, N1952, N2075, N560);
not NOT1 (N4706, N4701);
buf BUF1 (N4707, N4699);
or OR3 (N4708, N4702, N1833, N2013);
nor NOR4 (N4709, N4703, N3240, N479, N1788);
and AND4 (N4710, N4696, N2247, N2390, N123);
nor NOR2 (N4711, N4681, N1780);
or OR2 (N4712, N4709, N4248);
xor XOR2 (N4713, N4706, N1785);
nand NAND3 (N4714, N4711, N282, N2910);
nand NAND4 (N4715, N4712, N3049, N4012, N4693);
buf BUF1 (N4716, N4715);
not NOT1 (N4717, N4698);
buf BUF1 (N4718, N4717);
buf BUF1 (N4719, N4713);
or OR3 (N4720, N4707, N4251, N968);
buf BUF1 (N4721, N4718);
nor NOR4 (N4722, N4708, N1756, N2895, N4146);
xor XOR2 (N4723, N4714, N3884);
or OR2 (N4724, N4705, N3546);
buf BUF1 (N4725, N4720);
nor NOR4 (N4726, N4725, N4336, N2324, N1180);
or OR3 (N4727, N4721, N1726, N2292);
buf BUF1 (N4728, N4719);
nand NAND2 (N4729, N4723, N4032);
not NOT1 (N4730, N4710);
not NOT1 (N4731, N4729);
or OR2 (N4732, N4730, N2814);
buf BUF1 (N4733, N4726);
nor NOR2 (N4734, N4716, N1183);
nand NAND4 (N4735, N4733, N4696, N2694, N3164);
or OR2 (N4736, N4683, N2580);
xor XOR2 (N4737, N4724, N4347);
nor NOR4 (N4738, N4704, N3741, N2696, N728);
xor XOR2 (N4739, N4737, N3253);
buf BUF1 (N4740, N4731);
and AND4 (N4741, N4732, N3041, N1060, N3138);
nand NAND3 (N4742, N4741, N1741, N3176);
and AND4 (N4743, N4736, N1800, N2341, N4561);
buf BUF1 (N4744, N4742);
nor NOR2 (N4745, N4740, N2865);
buf BUF1 (N4746, N4727);
buf BUF1 (N4747, N4738);
or OR2 (N4748, N4743, N1231);
xor XOR2 (N4749, N4722, N593);
buf BUF1 (N4750, N4744);
nor NOR2 (N4751, N4745, N3765);
xor XOR2 (N4752, N4728, N984);
and AND3 (N4753, N4746, N1677, N3717);
not NOT1 (N4754, N4751);
not NOT1 (N4755, N4748);
xor XOR2 (N4756, N4750, N2204);
nor NOR4 (N4757, N4755, N4600, N2322, N20);
nor NOR2 (N4758, N4752, N4034);
nand NAND4 (N4759, N4747, N4755, N1504, N1465);
nand NAND3 (N4760, N4734, N2482, N2209);
nor NOR3 (N4761, N4758, N1223, N3022);
and AND3 (N4762, N4761, N628, N241);
nor NOR2 (N4763, N4735, N2219);
nand NAND3 (N4764, N4762, N2873, N3971);
xor XOR2 (N4765, N4753, N4679);
xor XOR2 (N4766, N4749, N3372);
xor XOR2 (N4767, N4756, N1310);
nand NAND3 (N4768, N4759, N1709, N887);
xor XOR2 (N4769, N4765, N3210);
buf BUF1 (N4770, N4754);
buf BUF1 (N4771, N4766);
and AND3 (N4772, N4764, N1085, N77);
and AND2 (N4773, N4757, N1673);
nand NAND2 (N4774, N4770, N4763);
nor NOR3 (N4775, N32, N566, N2157);
xor XOR2 (N4776, N4774, N3259);
nand NAND2 (N4777, N4760, N1583);
or OR2 (N4778, N4767, N1602);
buf BUF1 (N4779, N4739);
or OR4 (N4780, N4768, N2575, N2560, N2230);
and AND2 (N4781, N4775, N2351);
and AND4 (N4782, N4772, N3404, N3958, N4614);
not NOT1 (N4783, N4781);
xor XOR2 (N4784, N4779, N871);
and AND2 (N4785, N4777, N2157);
nor NOR3 (N4786, N4776, N456, N3796);
buf BUF1 (N4787, N4784);
buf BUF1 (N4788, N4787);
buf BUF1 (N4789, N4778);
and AND2 (N4790, N4773, N4288);
or OR3 (N4791, N4790, N1832, N792);
not NOT1 (N4792, N4771);
or OR2 (N4793, N4788, N3606);
xor XOR2 (N4794, N4785, N494);
xor XOR2 (N4795, N4794, N3818);
or OR2 (N4796, N4793, N1460);
nand NAND3 (N4797, N4769, N2740, N1187);
not NOT1 (N4798, N4795);
not NOT1 (N4799, N4783);
nor NOR4 (N4800, N4792, N1165, N2988, N4329);
nand NAND4 (N4801, N4799, N3326, N1424, N4486);
and AND3 (N4802, N4797, N3193, N1193);
nand NAND2 (N4803, N4782, N2307);
or OR4 (N4804, N4791, N1095, N1659, N3050);
not NOT1 (N4805, N4786);
not NOT1 (N4806, N4780);
or OR3 (N4807, N4804, N2128, N1062);
xor XOR2 (N4808, N4807, N632);
buf BUF1 (N4809, N4801);
nor NOR4 (N4810, N4796, N3725, N2871, N1284);
buf BUF1 (N4811, N4803);
or OR2 (N4812, N4806, N1943);
or OR4 (N4813, N4789, N1743, N918, N1853);
buf BUF1 (N4814, N4802);
and AND4 (N4815, N4809, N2954, N1448, N4657);
not NOT1 (N4816, N4808);
buf BUF1 (N4817, N4800);
not NOT1 (N4818, N4812);
xor XOR2 (N4819, N4817, N2331);
and AND4 (N4820, N4816, N2338, N2787, N2443);
not NOT1 (N4821, N4819);
xor XOR2 (N4822, N4811, N3197);
xor XOR2 (N4823, N4814, N2823);
and AND2 (N4824, N4798, N1954);
not NOT1 (N4825, N4821);
nand NAND4 (N4826, N4820, N2659, N810, N1109);
nand NAND3 (N4827, N4826, N3237, N2426);
and AND2 (N4828, N4815, N3241);
nand NAND3 (N4829, N4828, N2995, N3056);
nand NAND4 (N4830, N4823, N33, N1574, N2341);
or OR2 (N4831, N4824, N563);
not NOT1 (N4832, N4805);
xor XOR2 (N4833, N4830, N1055);
or OR3 (N4834, N4831, N1529, N3992);
xor XOR2 (N4835, N4818, N313);
nor NOR3 (N4836, N4835, N2045, N1427);
xor XOR2 (N4837, N4810, N2342);
xor XOR2 (N4838, N4837, N1497);
or OR2 (N4839, N4825, N3644);
nor NOR3 (N4840, N4827, N3165, N4496);
nand NAND3 (N4841, N4838, N2129, N1441);
not NOT1 (N4842, N4839);
nand NAND3 (N4843, N4829, N1774, N4039);
or OR4 (N4844, N4842, N2765, N691, N95);
buf BUF1 (N4845, N4813);
and AND2 (N4846, N4840, N857);
xor XOR2 (N4847, N4844, N3318);
not NOT1 (N4848, N4822);
nand NAND2 (N4849, N4833, N1104);
and AND4 (N4850, N4836, N3279, N4322, N1967);
and AND4 (N4851, N4849, N1281, N3424, N2467);
nor NOR3 (N4852, N4846, N4320, N1333);
nor NOR4 (N4853, N4841, N3706, N2838, N3047);
nand NAND4 (N4854, N4853, N2940, N1681, N4046);
xor XOR2 (N4855, N4850, N827);
nor NOR3 (N4856, N4843, N2406, N2908);
or OR3 (N4857, N4856, N2917, N1913);
and AND2 (N4858, N4848, N3630);
and AND2 (N4859, N4854, N2701);
and AND3 (N4860, N4834, N1273, N3236);
xor XOR2 (N4861, N4845, N4358);
and AND4 (N4862, N4859, N966, N3979, N2265);
nor NOR4 (N4863, N4860, N4240, N4801, N4366);
buf BUF1 (N4864, N4855);
nand NAND4 (N4865, N4861, N854, N563, N2315);
not NOT1 (N4866, N4857);
nor NOR3 (N4867, N4852, N3312, N247);
nand NAND3 (N4868, N4866, N2335, N4187);
xor XOR2 (N4869, N4864, N2596);
nand NAND2 (N4870, N4869, N4268);
nand NAND4 (N4871, N4863, N811, N716, N1591);
nand NAND4 (N4872, N4868, N1611, N1490, N1083);
or OR2 (N4873, N4832, N4274);
nand NAND3 (N4874, N4847, N455, N1050);
or OR3 (N4875, N4872, N3492, N168);
nand NAND4 (N4876, N4871, N988, N194, N13);
not NOT1 (N4877, N4876);
or OR3 (N4878, N4867, N1066, N638);
not NOT1 (N4879, N4870);
nor NOR4 (N4880, N4858, N2770, N1346, N3604);
nand NAND2 (N4881, N4851, N619);
nor NOR3 (N4882, N4873, N3886, N764);
or OR4 (N4883, N4865, N1007, N4836, N4568);
xor XOR2 (N4884, N4877, N3176);
xor XOR2 (N4885, N4880, N3905);
xor XOR2 (N4886, N4881, N2990);
not NOT1 (N4887, N4862);
xor XOR2 (N4888, N4883, N300);
not NOT1 (N4889, N4886);
nor NOR4 (N4890, N4882, N2895, N1623, N3483);
and AND4 (N4891, N4887, N1462, N386, N77);
nand NAND4 (N4892, N4891, N189, N1775, N3227);
nor NOR3 (N4893, N4884, N2299, N155);
or OR3 (N4894, N4879, N1437, N3047);
xor XOR2 (N4895, N4890, N2032);
buf BUF1 (N4896, N4894);
not NOT1 (N4897, N4885);
nor NOR2 (N4898, N4893, N3696);
buf BUF1 (N4899, N4897);
nand NAND2 (N4900, N4899, N764);
not NOT1 (N4901, N4875);
or OR3 (N4902, N4874, N1598, N4678);
xor XOR2 (N4903, N4895, N1661);
nand NAND2 (N4904, N4892, N3644);
nor NOR3 (N4905, N4904, N1164, N3433);
nand NAND2 (N4906, N4905, N3234);
buf BUF1 (N4907, N4906);
nor NOR2 (N4908, N4903, N2569);
nor NOR4 (N4909, N4896, N1626, N2992, N434);
nand NAND3 (N4910, N4878, N288, N4579);
or OR3 (N4911, N4901, N3913, N2655);
buf BUF1 (N4912, N4902);
not NOT1 (N4913, N4912);
buf BUF1 (N4914, N4913);
nor NOR2 (N4915, N4900, N2576);
xor XOR2 (N4916, N4910, N63);
nor NOR4 (N4917, N4909, N2176, N1751, N4132);
xor XOR2 (N4918, N4908, N1653);
nand NAND4 (N4919, N4911, N3852, N3584, N2993);
and AND2 (N4920, N4898, N608);
or OR3 (N4921, N4907, N3242, N2462);
and AND3 (N4922, N4889, N1733, N1340);
nor NOR2 (N4923, N4918, N2975);
and AND2 (N4924, N4922, N1166);
not NOT1 (N4925, N4888);
not NOT1 (N4926, N4917);
nand NAND2 (N4927, N4920, N2534);
nor NOR3 (N4928, N4919, N2870, N2770);
xor XOR2 (N4929, N4916, N4094);
not NOT1 (N4930, N4926);
nand NAND4 (N4931, N4921, N3784, N3577, N4573);
or OR3 (N4932, N4915, N1879, N4089);
buf BUF1 (N4933, N4924);
or OR4 (N4934, N4930, N3478, N4915, N345);
buf BUF1 (N4935, N4927);
buf BUF1 (N4936, N4928);
buf BUF1 (N4937, N4936);
xor XOR2 (N4938, N4914, N1019);
not NOT1 (N4939, N4925);
and AND2 (N4940, N4931, N2846);
nor NOR3 (N4941, N4940, N1040, N3706);
not NOT1 (N4942, N4941);
xor XOR2 (N4943, N4939, N2744);
buf BUF1 (N4944, N4938);
nand NAND2 (N4945, N4944, N2304);
buf BUF1 (N4946, N4932);
nand NAND3 (N4947, N4929, N4004, N2920);
not NOT1 (N4948, N4947);
or OR2 (N4949, N4943, N3112);
buf BUF1 (N4950, N4933);
nor NOR4 (N4951, N4934, N4060, N4245, N541);
buf BUF1 (N4952, N4949);
buf BUF1 (N4953, N4945);
and AND2 (N4954, N4946, N169);
or OR2 (N4955, N4923, N705);
nor NOR3 (N4956, N4942, N2672, N4020);
xor XOR2 (N4957, N4951, N2247);
nor NOR4 (N4958, N4948, N4578, N615, N4893);
not NOT1 (N4959, N4953);
buf BUF1 (N4960, N4957);
nor NOR4 (N4961, N4958, N308, N1785, N947);
nand NAND4 (N4962, N4961, N3284, N4867, N1508);
and AND3 (N4963, N4952, N4096, N3570);
nand NAND2 (N4964, N4937, N288);
nand NAND4 (N4965, N4954, N2537, N2348, N2231);
nor NOR2 (N4966, N4956, N2868);
nand NAND4 (N4967, N4964, N2748, N1640, N3128);
buf BUF1 (N4968, N4955);
buf BUF1 (N4969, N4935);
nor NOR4 (N4970, N4969, N4349, N4944, N4807);
nand NAND2 (N4971, N4959, N3235);
buf BUF1 (N4972, N4962);
nor NOR2 (N4973, N4950, N677);
buf BUF1 (N4974, N4960);
nand NAND4 (N4975, N4971, N826, N2285, N74);
not NOT1 (N4976, N4965);
nor NOR4 (N4977, N4968, N2906, N936, N4655);
not NOT1 (N4978, N4974);
buf BUF1 (N4979, N4970);
not NOT1 (N4980, N4963);
not NOT1 (N4981, N4978);
and AND3 (N4982, N4972, N3173, N4352);
or OR4 (N4983, N4980, N3086, N1542, N1602);
nand NAND2 (N4984, N4981, N2376);
nor NOR4 (N4985, N4973, N2923, N4159, N569);
xor XOR2 (N4986, N4985, N3058);
or OR3 (N4987, N4977, N1934, N4169);
nand NAND4 (N4988, N4982, N61, N4850, N1162);
nand NAND4 (N4989, N4987, N3111, N4367, N4499);
nor NOR2 (N4990, N4989, N1623);
and AND2 (N4991, N4975, N4353);
not NOT1 (N4992, N4986);
and AND4 (N4993, N4992, N2314, N1648, N1667);
nor NOR3 (N4994, N4990, N557, N3317);
or OR2 (N4995, N4967, N1599);
nor NOR2 (N4996, N4979, N3180);
not NOT1 (N4997, N4996);
buf BUF1 (N4998, N4997);
and AND3 (N4999, N4991, N4224, N937);
nor NOR4 (N5000, N4994, N1821, N1928, N2989);
xor XOR2 (N5001, N4995, N3151);
nor NOR4 (N5002, N4993, N1961, N1302, N1863);
buf BUF1 (N5003, N4999);
not NOT1 (N5004, N4998);
xor XOR2 (N5005, N4976, N4999);
buf BUF1 (N5006, N5001);
or OR3 (N5007, N5000, N2262, N4537);
not NOT1 (N5008, N5003);
or OR3 (N5009, N5004, N1982, N3050);
xor XOR2 (N5010, N4983, N1394);
not NOT1 (N5011, N4984);
xor XOR2 (N5012, N5006, N4842);
and AND4 (N5013, N4988, N4294, N4869, N3538);
and AND3 (N5014, N4966, N212, N4519);
not NOT1 (N5015, N5005);
nand NAND4 (N5016, N5014, N4888, N1166, N889);
buf BUF1 (N5017, N5015);
buf BUF1 (N5018, N5012);
xor XOR2 (N5019, N5010, N4446);
and AND3 (N5020, N5002, N1114, N4496);
buf BUF1 (N5021, N5013);
not NOT1 (N5022, N5007);
not NOT1 (N5023, N5009);
xor XOR2 (N5024, N5008, N2474);
xor XOR2 (N5025, N5023, N3511);
not NOT1 (N5026, N5020);
buf BUF1 (N5027, N5011);
nand NAND3 (N5028, N5027, N1521, N2464);
or OR3 (N5029, N5028, N3708, N4325);
xor XOR2 (N5030, N5017, N4632);
xor XOR2 (N5031, N5024, N150);
or OR2 (N5032, N5031, N942);
xor XOR2 (N5033, N5025, N2208);
xor XOR2 (N5034, N5019, N2177);
and AND3 (N5035, N5033, N4635, N1071);
nand NAND4 (N5036, N5021, N3740, N1700, N2290);
and AND2 (N5037, N5029, N1228);
xor XOR2 (N5038, N5022, N2032);
or OR2 (N5039, N5034, N89);
or OR2 (N5040, N5032, N4496);
buf BUF1 (N5041, N5035);
buf BUF1 (N5042, N5041);
or OR3 (N5043, N5030, N3705, N3589);
buf BUF1 (N5044, N5038);
and AND4 (N5045, N5043, N4442, N1158, N4906);
nand NAND4 (N5046, N5044, N626, N2978, N659);
and AND3 (N5047, N5036, N1686, N1938);
nand NAND4 (N5048, N5026, N1225, N3892, N3776);
or OR2 (N5049, N5039, N2649);
or OR4 (N5050, N5042, N1817, N4093, N2167);
xor XOR2 (N5051, N5048, N4999);
nand NAND4 (N5052, N5046, N244, N4521, N3453);
nor NOR3 (N5053, N5040, N1309, N4924);
and AND4 (N5054, N5049, N604, N1544, N3041);
buf BUF1 (N5055, N5054);
nand NAND4 (N5056, N5053, N993, N4525, N4266);
buf BUF1 (N5057, N5037);
and AND2 (N5058, N5018, N2003);
nor NOR4 (N5059, N5057, N383, N3531, N2394);
nand NAND4 (N5060, N5045, N1336, N161, N3819);
not NOT1 (N5061, N5056);
buf BUF1 (N5062, N5047);
nor NOR4 (N5063, N5052, N4746, N4534, N3009);
nand NAND3 (N5064, N5050, N3209, N3681);
and AND3 (N5065, N5051, N2749, N1768);
nor NOR4 (N5066, N5064, N3062, N1574, N2149);
or OR2 (N5067, N5061, N3990);
nand NAND4 (N5068, N5062, N3311, N3226, N2372);
or OR2 (N5069, N5055, N3488);
nand NAND4 (N5070, N5063, N4363, N2110, N1260);
nor NOR3 (N5071, N5065, N2403, N1935);
and AND2 (N5072, N5071, N4806);
and AND4 (N5073, N5067, N886, N1246, N3781);
nor NOR4 (N5074, N5066, N230, N3160, N3532);
buf BUF1 (N5075, N5058);
or OR2 (N5076, N5072, N979);
and AND2 (N5077, N5060, N1458);
not NOT1 (N5078, N5073);
or OR3 (N5079, N5077, N924, N1811);
not NOT1 (N5080, N5068);
and AND3 (N5081, N5080, N3495, N3922);
nand NAND3 (N5082, N5059, N4902, N3373);
and AND4 (N5083, N5082, N4351, N784, N107);
buf BUF1 (N5084, N5081);
or OR4 (N5085, N5074, N1732, N4794, N1753);
and AND2 (N5086, N5083, N1575);
not NOT1 (N5087, N5076);
nand NAND4 (N5088, N5084, N363, N3384, N2647);
and AND2 (N5089, N5079, N3712);
and AND4 (N5090, N5069, N3065, N4167, N1635);
or OR4 (N5091, N5078, N1485, N1920, N354);
and AND2 (N5092, N5085, N3567);
and AND4 (N5093, N5090, N4182, N1616, N3965);
nor NOR4 (N5094, N5092, N2596, N3874, N1153);
nand NAND2 (N5095, N5075, N2140);
not NOT1 (N5096, N5091);
or OR2 (N5097, N5095, N4077);
xor XOR2 (N5098, N5070, N3059);
buf BUF1 (N5099, N5016);
nand NAND4 (N5100, N5099, N161, N294, N513);
xor XOR2 (N5101, N5096, N3588);
buf BUF1 (N5102, N5093);
buf BUF1 (N5103, N5101);
not NOT1 (N5104, N5100);
xor XOR2 (N5105, N5104, N719);
or OR4 (N5106, N5087, N74, N2420, N3273);
or OR2 (N5107, N5103, N4344);
xor XOR2 (N5108, N5094, N4913);
xor XOR2 (N5109, N5088, N1388);
nor NOR4 (N5110, N5089, N510, N2187, N3866);
or OR4 (N5111, N5109, N4062, N630, N4770);
not NOT1 (N5112, N5111);
xor XOR2 (N5113, N5105, N2533);
nor NOR2 (N5114, N5102, N4480);
nand NAND4 (N5115, N5098, N4391, N3895, N5058);
not NOT1 (N5116, N5097);
buf BUF1 (N5117, N5107);
xor XOR2 (N5118, N5115, N140);
xor XOR2 (N5119, N5110, N3886);
and AND4 (N5120, N5119, N738, N2142, N4493);
not NOT1 (N5121, N5117);
nor NOR2 (N5122, N5108, N245);
not NOT1 (N5123, N5118);
or OR2 (N5124, N5116, N4219);
buf BUF1 (N5125, N5113);
nor NOR4 (N5126, N5120, N1428, N3742, N552);
nor NOR2 (N5127, N5112, N4038);
nor NOR3 (N5128, N5127, N1443, N3720);
and AND2 (N5129, N5114, N4585);
and AND2 (N5130, N5128, N689);
nor NOR2 (N5131, N5124, N1815);
and AND3 (N5132, N5125, N4306, N3976);
xor XOR2 (N5133, N5130, N2904);
nor NOR3 (N5134, N5086, N250, N1030);
nand NAND2 (N5135, N5123, N4774);
nor NOR3 (N5136, N5131, N3323, N1170);
not NOT1 (N5137, N5126);
nor NOR3 (N5138, N5135, N4099, N1972);
nand NAND3 (N5139, N5138, N4202, N167);
xor XOR2 (N5140, N5139, N1837);
nor NOR4 (N5141, N5137, N762, N1849, N1794);
xor XOR2 (N5142, N5132, N3665);
or OR4 (N5143, N5122, N2413, N599, N81);
nand NAND2 (N5144, N5140, N3579);
xor XOR2 (N5145, N5134, N1958);
buf BUF1 (N5146, N5129);
xor XOR2 (N5147, N5141, N4927);
nor NOR4 (N5148, N5106, N803, N1557, N1532);
xor XOR2 (N5149, N5148, N5139);
nor NOR4 (N5150, N5143, N2353, N3871, N4503);
nand NAND3 (N5151, N5144, N4479, N1341);
nor NOR2 (N5152, N5146, N4722);
and AND4 (N5153, N5145, N1428, N456, N4962);
nand NAND3 (N5154, N5149, N2771, N3062);
nor NOR4 (N5155, N5142, N1646, N3909, N4733);
xor XOR2 (N5156, N5150, N1963);
or OR2 (N5157, N5152, N4250);
buf BUF1 (N5158, N5147);
nand NAND3 (N5159, N5156, N4082, N752);
and AND2 (N5160, N5158, N1942);
not NOT1 (N5161, N5157);
buf BUF1 (N5162, N5151);
not NOT1 (N5163, N5133);
buf BUF1 (N5164, N5162);
and AND4 (N5165, N5154, N4440, N2549, N1263);
or OR3 (N5166, N5153, N4781, N3035);
xor XOR2 (N5167, N5159, N678);
or OR2 (N5168, N5155, N3663);
nor NOR3 (N5169, N5166, N571, N1004);
nor NOR4 (N5170, N5160, N1420, N684, N593);
or OR3 (N5171, N5163, N70, N3098);
nor NOR2 (N5172, N5161, N3009);
or OR3 (N5173, N5168, N1814, N1703);
and AND3 (N5174, N5173, N1724, N3434);
buf BUF1 (N5175, N5172);
buf BUF1 (N5176, N5165);
nor NOR2 (N5177, N5164, N2503);
not NOT1 (N5178, N5174);
or OR3 (N5179, N5121, N2728, N120);
nand NAND4 (N5180, N5169, N84, N4254, N3792);
not NOT1 (N5181, N5167);
nand NAND3 (N5182, N5180, N3662, N182);
or OR2 (N5183, N5136, N4934);
xor XOR2 (N5184, N5170, N2338);
buf BUF1 (N5185, N5184);
and AND4 (N5186, N5175, N3582, N4064, N674);
or OR2 (N5187, N5177, N1986);
and AND4 (N5188, N5187, N4754, N1286, N2029);
xor XOR2 (N5189, N5178, N4499);
not NOT1 (N5190, N5185);
or OR3 (N5191, N5182, N1515, N5017);
nand NAND4 (N5192, N5191, N157, N560, N1484);
not NOT1 (N5193, N5189);
nor NOR4 (N5194, N5183, N2534, N3139, N609);
buf BUF1 (N5195, N5171);
nand NAND3 (N5196, N5186, N2163, N3343);
buf BUF1 (N5197, N5181);
or OR2 (N5198, N5196, N2321);
xor XOR2 (N5199, N5193, N1328);
and AND3 (N5200, N5190, N3791, N2579);
nor NOR2 (N5201, N5195, N3442);
and AND3 (N5202, N5176, N5033, N1908);
buf BUF1 (N5203, N5198);
nor NOR3 (N5204, N5200, N3690, N2306);
nor NOR4 (N5205, N5194, N2038, N2303, N4904);
buf BUF1 (N5206, N5202);
and AND3 (N5207, N5192, N1200, N4357);
and AND2 (N5208, N5205, N4192);
and AND3 (N5209, N5188, N4814, N126);
and AND2 (N5210, N5209, N3213);
xor XOR2 (N5211, N5199, N3010);
and AND4 (N5212, N5210, N4721, N4035, N343);
xor XOR2 (N5213, N5203, N4958);
nor NOR3 (N5214, N5179, N5059, N4727);
nand NAND4 (N5215, N5211, N1271, N1378, N1868);
nand NAND4 (N5216, N5201, N941, N2647, N4357);
nor NOR4 (N5217, N5206, N5036, N3671, N2135);
not NOT1 (N5218, N5204);
buf BUF1 (N5219, N5207);
or OR3 (N5220, N5197, N1733, N3642);
not NOT1 (N5221, N5212);
buf BUF1 (N5222, N5213);
or OR4 (N5223, N5220, N273, N4702, N1906);
buf BUF1 (N5224, N5214);
or OR4 (N5225, N5221, N2022, N3214, N2856);
nand NAND2 (N5226, N5215, N3600);
xor XOR2 (N5227, N5216, N2768);
nor NOR2 (N5228, N5227, N1741);
not NOT1 (N5229, N5219);
nand NAND3 (N5230, N5208, N174, N4419);
and AND2 (N5231, N5224, N4157);
buf BUF1 (N5232, N5231);
xor XOR2 (N5233, N5218, N2482);
xor XOR2 (N5234, N5233, N459);
xor XOR2 (N5235, N5217, N596);
not NOT1 (N5236, N5223);
and AND3 (N5237, N5229, N2137, N1279);
xor XOR2 (N5238, N5236, N987);
xor XOR2 (N5239, N5235, N814);
or OR2 (N5240, N5239, N578);
and AND2 (N5241, N5228, N5178);
nor NOR4 (N5242, N5225, N3577, N3824, N561);
xor XOR2 (N5243, N5232, N4412);
not NOT1 (N5244, N5238);
nand NAND2 (N5245, N5242, N1827);
buf BUF1 (N5246, N5222);
not NOT1 (N5247, N5244);
not NOT1 (N5248, N5246);
nand NAND2 (N5249, N5247, N4219);
buf BUF1 (N5250, N5243);
nand NAND2 (N5251, N5250, N979);
and AND4 (N5252, N5251, N3719, N3990, N949);
xor XOR2 (N5253, N5249, N1137);
nor NOR2 (N5254, N5252, N4282);
xor XOR2 (N5255, N5230, N1995);
nand NAND3 (N5256, N5245, N2454, N2998);
or OR2 (N5257, N5240, N1065);
xor XOR2 (N5258, N5257, N2045);
nand NAND3 (N5259, N5255, N3923, N3345);
nor NOR3 (N5260, N5254, N1424, N3402);
xor XOR2 (N5261, N5260, N737);
not NOT1 (N5262, N5234);
or OR3 (N5263, N5248, N3870, N801);
or OR4 (N5264, N5256, N491, N1921, N2652);
or OR3 (N5265, N5226, N1070, N3902);
nand NAND4 (N5266, N5237, N462, N186, N434);
not NOT1 (N5267, N5261);
xor XOR2 (N5268, N5253, N4864);
not NOT1 (N5269, N5265);
and AND2 (N5270, N5267, N3844);
xor XOR2 (N5271, N5269, N2807);
or OR2 (N5272, N5268, N1932);
or OR4 (N5273, N5263, N2370, N4835, N4137);
xor XOR2 (N5274, N5266, N1928);
not NOT1 (N5275, N5258);
not NOT1 (N5276, N5262);
and AND2 (N5277, N5274, N487);
or OR2 (N5278, N5270, N1324);
nor NOR3 (N5279, N5272, N3563, N3276);
nor NOR3 (N5280, N5259, N5047, N3832);
nand NAND3 (N5281, N5278, N1978, N3505);
and AND3 (N5282, N5264, N4131, N3487);
or OR4 (N5283, N5275, N2319, N5187, N4111);
not NOT1 (N5284, N5277);
or OR4 (N5285, N5271, N1308, N4244, N1815);
or OR4 (N5286, N5283, N2597, N1788, N4129);
or OR4 (N5287, N5273, N1150, N3790, N25);
and AND4 (N5288, N5282, N1949, N3926, N1457);
xor XOR2 (N5289, N5241, N4444);
xor XOR2 (N5290, N5289, N3028);
or OR2 (N5291, N5286, N4049);
not NOT1 (N5292, N5284);
nor NOR2 (N5293, N5280, N3264);
and AND4 (N5294, N5287, N679, N1225, N4549);
nor NOR3 (N5295, N5293, N3374, N1780);
buf BUF1 (N5296, N5292);
buf BUF1 (N5297, N5285);
not NOT1 (N5298, N5279);
not NOT1 (N5299, N5296);
nand NAND3 (N5300, N5288, N2672, N3825);
or OR3 (N5301, N5298, N4781, N4957);
xor XOR2 (N5302, N5297, N5144);
and AND4 (N5303, N5300, N4282, N4898, N3812);
and AND3 (N5304, N5301, N4011, N1960);
xor XOR2 (N5305, N5303, N1864);
and AND2 (N5306, N5302, N2097);
not NOT1 (N5307, N5276);
nor NOR2 (N5308, N5294, N1201);
nor NOR3 (N5309, N5306, N67, N3512);
and AND3 (N5310, N5309, N3949, N218);
and AND3 (N5311, N5291, N552, N533);
or OR4 (N5312, N5281, N3802, N1493, N4738);
not NOT1 (N5313, N5305);
and AND3 (N5314, N5310, N788, N4561);
xor XOR2 (N5315, N5295, N213);
nor NOR3 (N5316, N5299, N692, N4817);
nand NAND2 (N5317, N5316, N3623);
xor XOR2 (N5318, N5304, N4485);
or OR3 (N5319, N5314, N4653, N1653);
and AND3 (N5320, N5311, N4839, N2330);
nor NOR4 (N5321, N5290, N1600, N5259, N300);
xor XOR2 (N5322, N5308, N2694);
not NOT1 (N5323, N5315);
xor XOR2 (N5324, N5323, N1854);
buf BUF1 (N5325, N5318);
buf BUF1 (N5326, N5325);
xor XOR2 (N5327, N5320, N2594);
nor NOR2 (N5328, N5307, N4475);
or OR4 (N5329, N5328, N4874, N4086, N4511);
and AND4 (N5330, N5317, N1374, N2882, N4030);
or OR4 (N5331, N5327, N3300, N2133, N907);
or OR2 (N5332, N5319, N2676);
xor XOR2 (N5333, N5331, N876);
nand NAND3 (N5334, N5313, N3810, N2192);
buf BUF1 (N5335, N5332);
xor XOR2 (N5336, N5324, N1189);
xor XOR2 (N5337, N5312, N3187);
nand NAND3 (N5338, N5334, N3533, N3996);
nand NAND2 (N5339, N5329, N699);
not NOT1 (N5340, N5337);
nor NOR4 (N5341, N5330, N500, N2306, N551);
nor NOR2 (N5342, N5340, N4546);
nand NAND3 (N5343, N5336, N3870, N3448);
nor NOR3 (N5344, N5335, N1175, N939);
or OR3 (N5345, N5343, N4627, N4631);
and AND3 (N5346, N5321, N3000, N4011);
nor NOR3 (N5347, N5339, N2512, N4381);
nand NAND2 (N5348, N5333, N4825);
and AND2 (N5349, N5345, N350);
xor XOR2 (N5350, N5344, N1924);
or OR4 (N5351, N5348, N2263, N2984, N4985);
xor XOR2 (N5352, N5350, N1749);
nor NOR2 (N5353, N5341, N591);
or OR2 (N5354, N5349, N708);
nand NAND2 (N5355, N5347, N1145);
not NOT1 (N5356, N5352);
buf BUF1 (N5357, N5355);
not NOT1 (N5358, N5354);
or OR2 (N5359, N5338, N4445);
xor XOR2 (N5360, N5346, N1489);
not NOT1 (N5361, N5342);
buf BUF1 (N5362, N5361);
xor XOR2 (N5363, N5360, N4887);
nor NOR3 (N5364, N5362, N4045, N4942);
and AND2 (N5365, N5357, N1295);
buf BUF1 (N5366, N5326);
nor NOR4 (N5367, N5365, N2494, N3546, N4282);
or OR4 (N5368, N5367, N3935, N4451, N974);
buf BUF1 (N5369, N5356);
or OR2 (N5370, N5368, N2111);
not NOT1 (N5371, N5364);
nand NAND3 (N5372, N5322, N3933, N4384);
buf BUF1 (N5373, N5351);
not NOT1 (N5374, N5373);
xor XOR2 (N5375, N5363, N3583);
nor NOR2 (N5376, N5358, N1653);
or OR4 (N5377, N5375, N2718, N2613, N3455);
buf BUF1 (N5378, N5366);
and AND4 (N5379, N5377, N5001, N4837, N3935);
xor XOR2 (N5380, N5378, N36);
nand NAND3 (N5381, N5376, N1474, N318);
buf BUF1 (N5382, N5370);
buf BUF1 (N5383, N5379);
nor NOR4 (N5384, N5359, N3709, N848, N5306);
nand NAND3 (N5385, N5382, N1473, N918);
or OR3 (N5386, N5383, N796, N2199);
or OR2 (N5387, N5353, N2072);
not NOT1 (N5388, N5387);
buf BUF1 (N5389, N5380);
xor XOR2 (N5390, N5388, N1050);
and AND2 (N5391, N5372, N483);
and AND3 (N5392, N5386, N620, N5254);
buf BUF1 (N5393, N5369);
not NOT1 (N5394, N5390);
buf BUF1 (N5395, N5394);
xor XOR2 (N5396, N5392, N776);
and AND2 (N5397, N5389, N1053);
buf BUF1 (N5398, N5396);
xor XOR2 (N5399, N5397, N5122);
buf BUF1 (N5400, N5371);
xor XOR2 (N5401, N5374, N4522);
xor XOR2 (N5402, N5399, N292);
or OR2 (N5403, N5402, N3182);
buf BUF1 (N5404, N5398);
or OR2 (N5405, N5391, N1859);
or OR2 (N5406, N5395, N918);
and AND3 (N5407, N5401, N150, N5390);
buf BUF1 (N5408, N5381);
nand NAND3 (N5409, N5384, N1511, N4890);
nand NAND2 (N5410, N5403, N3753);
or OR4 (N5411, N5405, N153, N4951, N2354);
nor NOR4 (N5412, N5393, N3344, N2703, N901);
and AND4 (N5413, N5412, N4424, N4919, N2192);
nor NOR4 (N5414, N5410, N5212, N3286, N2235);
buf BUF1 (N5415, N5408);
buf BUF1 (N5416, N5406);
buf BUF1 (N5417, N5413);
not NOT1 (N5418, N5407);
not NOT1 (N5419, N5415);
xor XOR2 (N5420, N5400, N3824);
buf BUF1 (N5421, N5409);
not NOT1 (N5422, N5414);
and AND3 (N5423, N5419, N3555, N1669);
or OR2 (N5424, N5385, N3860);
not NOT1 (N5425, N5424);
nor NOR3 (N5426, N5404, N3895, N426);
nand NAND2 (N5427, N5418, N420);
and AND2 (N5428, N5411, N2735);
nor NOR2 (N5429, N5428, N4947);
xor XOR2 (N5430, N5425, N4713);
not NOT1 (N5431, N5426);
nand NAND2 (N5432, N5430, N3887);
xor XOR2 (N5433, N5420, N5140);
nand NAND2 (N5434, N5417, N4637);
buf BUF1 (N5435, N5431);
or OR4 (N5436, N5432, N178, N342, N3041);
and AND3 (N5437, N5429, N2311, N3966);
nor NOR4 (N5438, N5437, N754, N1314, N4257);
nand NAND4 (N5439, N5416, N2391, N3326, N670);
nand NAND2 (N5440, N5439, N1632);
nand NAND2 (N5441, N5423, N5217);
buf BUF1 (N5442, N5438);
buf BUF1 (N5443, N5442);
xor XOR2 (N5444, N5422, N1196);
xor XOR2 (N5445, N5441, N1116);
nand NAND3 (N5446, N5433, N2690, N606);
not NOT1 (N5447, N5445);
or OR3 (N5448, N5444, N1129, N4928);
nor NOR4 (N5449, N5446, N5264, N4565, N4821);
not NOT1 (N5450, N5421);
xor XOR2 (N5451, N5450, N3966);
nor NOR2 (N5452, N5427, N2062);
or OR2 (N5453, N5451, N5417);
nand NAND4 (N5454, N5449, N1128, N2340, N2662);
buf BUF1 (N5455, N5454);
or OR4 (N5456, N5448, N864, N850, N4871);
and AND4 (N5457, N5452, N587, N4031, N1458);
not NOT1 (N5458, N5453);
xor XOR2 (N5459, N5458, N5009);
buf BUF1 (N5460, N5436);
buf BUF1 (N5461, N5459);
xor XOR2 (N5462, N5455, N3947);
buf BUF1 (N5463, N5456);
nand NAND2 (N5464, N5461, N1696);
nand NAND4 (N5465, N5462, N2500, N2108, N4005);
nand NAND2 (N5466, N5465, N1030);
or OR3 (N5467, N5463, N2649, N1031);
buf BUF1 (N5468, N5467);
xor XOR2 (N5469, N5468, N5201);
nand NAND4 (N5470, N5443, N1965, N3377, N1288);
buf BUF1 (N5471, N5470);
nand NAND3 (N5472, N5447, N579, N1268);
not NOT1 (N5473, N5471);
buf BUF1 (N5474, N5469);
not NOT1 (N5475, N5440);
buf BUF1 (N5476, N5472);
xor XOR2 (N5477, N5464, N4017);
nand NAND3 (N5478, N5477, N805, N3070);
xor XOR2 (N5479, N5473, N4668);
not NOT1 (N5480, N5466);
not NOT1 (N5481, N5460);
xor XOR2 (N5482, N5481, N2607);
not NOT1 (N5483, N5474);
and AND4 (N5484, N5434, N2690, N4299, N15);
nand NAND2 (N5485, N5457, N483);
and AND3 (N5486, N5478, N943, N4139);
and AND2 (N5487, N5486, N491);
not NOT1 (N5488, N5485);
nor NOR4 (N5489, N5435, N121, N722, N468);
and AND3 (N5490, N5488, N460, N942);
not NOT1 (N5491, N5482);
nor NOR4 (N5492, N5483, N1572, N5407, N5417);
nor NOR2 (N5493, N5484, N4008);
or OR4 (N5494, N5479, N2747, N2851, N3771);
buf BUF1 (N5495, N5491);
buf BUF1 (N5496, N5493);
nand NAND3 (N5497, N5496, N395, N2370);
buf BUF1 (N5498, N5476);
xor XOR2 (N5499, N5498, N5325);
not NOT1 (N5500, N5480);
nand NAND2 (N5501, N5497, N2326);
and AND2 (N5502, N5492, N1992);
nand NAND4 (N5503, N5501, N3790, N2260, N685);
or OR4 (N5504, N5494, N1159, N5153, N1266);
nand NAND3 (N5505, N5495, N3015, N5277);
buf BUF1 (N5506, N5499);
or OR4 (N5507, N5502, N5100, N3483, N3131);
or OR4 (N5508, N5500, N1586, N4200, N1084);
not NOT1 (N5509, N5475);
nor NOR3 (N5510, N5487, N190, N3587);
buf BUF1 (N5511, N5489);
nand NAND3 (N5512, N5510, N3348, N82);
buf BUF1 (N5513, N5504);
nor NOR2 (N5514, N5490, N733);
or OR3 (N5515, N5505, N1187, N461);
buf BUF1 (N5516, N5509);
nand NAND3 (N5517, N5511, N463, N2684);
buf BUF1 (N5518, N5508);
or OR2 (N5519, N5515, N2247);
or OR2 (N5520, N5518, N5019);
and AND4 (N5521, N5519, N3493, N2944, N3883);
nand NAND2 (N5522, N5521, N118);
nand NAND4 (N5523, N5513, N163, N2855, N528);
and AND3 (N5524, N5514, N5240, N3158);
or OR3 (N5525, N5503, N735, N723);
xor XOR2 (N5526, N5512, N4594);
nand NAND2 (N5527, N5523, N2358);
nand NAND4 (N5528, N5524, N1410, N3081, N1788);
nand NAND4 (N5529, N5526, N4906, N3117, N3859);
nand NAND3 (N5530, N5529, N1206, N2425);
xor XOR2 (N5531, N5516, N4932);
or OR3 (N5532, N5528, N5101, N3701);
not NOT1 (N5533, N5517);
buf BUF1 (N5534, N5506);
and AND3 (N5535, N5534, N2062, N1556);
nor NOR3 (N5536, N5533, N5064, N1410);
nand NAND4 (N5537, N5535, N1882, N515, N4638);
xor XOR2 (N5538, N5536, N3646);
or OR2 (N5539, N5538, N3835);
nor NOR2 (N5540, N5530, N1381);
and AND3 (N5541, N5537, N868, N1265);
buf BUF1 (N5542, N5520);
or OR4 (N5543, N5531, N2431, N585, N493);
or OR3 (N5544, N5527, N2585, N5434);
buf BUF1 (N5545, N5507);
not NOT1 (N5546, N5541);
nor NOR3 (N5547, N5539, N2365, N4011);
or OR2 (N5548, N5542, N4072);
or OR2 (N5549, N5532, N2635);
and AND4 (N5550, N5549, N3089, N4257, N4987);
and AND4 (N5551, N5540, N2677, N2787, N791);
nor NOR3 (N5552, N5548, N5438, N1038);
and AND2 (N5553, N5543, N5168);
xor XOR2 (N5554, N5551, N3151);
or OR3 (N5555, N5553, N1179, N4212);
not NOT1 (N5556, N5554);
and AND2 (N5557, N5552, N3766);
buf BUF1 (N5558, N5522);
xor XOR2 (N5559, N5557, N3905);
and AND2 (N5560, N5556, N226);
xor XOR2 (N5561, N5546, N2761);
or OR2 (N5562, N5561, N147);
not NOT1 (N5563, N5558);
nor NOR2 (N5564, N5545, N1748);
nand NAND4 (N5565, N5547, N543, N4026, N2727);
or OR4 (N5566, N5555, N1965, N4011, N1790);
and AND4 (N5567, N5550, N849, N4804, N3055);
not NOT1 (N5568, N5560);
xor XOR2 (N5569, N5559, N120);
or OR4 (N5570, N5544, N2266, N3626, N2204);
xor XOR2 (N5571, N5562, N3113);
xor XOR2 (N5572, N5564, N674);
not NOT1 (N5573, N5569);
nor NOR4 (N5574, N5571, N1486, N3786, N3485);
nand NAND2 (N5575, N5573, N4569);
xor XOR2 (N5576, N5565, N4147);
nor NOR4 (N5577, N5563, N5320, N3201, N2003);
or OR2 (N5578, N5576, N4343);
and AND3 (N5579, N5567, N4389, N3077);
or OR3 (N5580, N5568, N3367, N4140);
and AND2 (N5581, N5579, N1439);
xor XOR2 (N5582, N5577, N1773);
nand NAND3 (N5583, N5578, N4079, N1549);
or OR4 (N5584, N5574, N3325, N2391, N729);
nand NAND4 (N5585, N5581, N3643, N2911, N350);
nor NOR4 (N5586, N5525, N5561, N2039, N4277);
buf BUF1 (N5587, N5585);
nand NAND4 (N5588, N5587, N1357, N4961, N2855);
nor NOR2 (N5589, N5580, N4669);
xor XOR2 (N5590, N5584, N2069);
nand NAND4 (N5591, N5586, N579, N4686, N973);
and AND2 (N5592, N5570, N1395);
nand NAND2 (N5593, N5588, N2262);
or OR2 (N5594, N5590, N1702);
not NOT1 (N5595, N5593);
nor NOR3 (N5596, N5566, N5382, N5312);
nor NOR3 (N5597, N5594, N1949, N3634);
nor NOR2 (N5598, N5572, N4555);
nor NOR2 (N5599, N5575, N4483);
and AND2 (N5600, N5596, N1928);
not NOT1 (N5601, N5582);
xor XOR2 (N5602, N5597, N5070);
nand NAND2 (N5603, N5595, N2166);
and AND3 (N5604, N5599, N3185, N4964);
xor XOR2 (N5605, N5602, N5155);
not NOT1 (N5606, N5601);
nor NOR3 (N5607, N5606, N5584, N4509);
nand NAND2 (N5608, N5603, N1898);
or OR4 (N5609, N5598, N2059, N2084, N1242);
nor NOR3 (N5610, N5605, N2992, N1489);
xor XOR2 (N5611, N5608, N5245);
or OR2 (N5612, N5604, N3452);
nand NAND4 (N5613, N5592, N3593, N4691, N4550);
and AND2 (N5614, N5611, N5152);
or OR3 (N5615, N5607, N3824, N2821);
xor XOR2 (N5616, N5610, N666);
xor XOR2 (N5617, N5612, N1494);
and AND2 (N5618, N5615, N894);
or OR4 (N5619, N5583, N859, N4280, N4433);
or OR4 (N5620, N5614, N2029, N3631, N2197);
and AND2 (N5621, N5619, N1388);
nand NAND2 (N5622, N5617, N3513);
not NOT1 (N5623, N5591);
xor XOR2 (N5624, N5620, N4416);
and AND2 (N5625, N5613, N2);
and AND4 (N5626, N5622, N405, N1675, N4653);
and AND3 (N5627, N5623, N1113, N1669);
nor NOR2 (N5628, N5625, N2009);
and AND3 (N5629, N5618, N4738, N553);
xor XOR2 (N5630, N5609, N2531);
and AND4 (N5631, N5600, N4427, N2759, N2501);
and AND3 (N5632, N5616, N999, N2482);
nor NOR4 (N5633, N5624, N3014, N836, N87);
xor XOR2 (N5634, N5630, N5043);
or OR4 (N5635, N5627, N462, N5491, N3632);
buf BUF1 (N5636, N5635);
not NOT1 (N5637, N5631);
nand NAND4 (N5638, N5628, N3096, N2500, N3849);
nor NOR2 (N5639, N5633, N3941);
not NOT1 (N5640, N5629);
xor XOR2 (N5641, N5634, N3209);
not NOT1 (N5642, N5641);
buf BUF1 (N5643, N5632);
buf BUF1 (N5644, N5589);
or OR2 (N5645, N5636, N3835);
not NOT1 (N5646, N5642);
nand NAND4 (N5647, N5639, N914, N1193, N3223);
buf BUF1 (N5648, N5626);
and AND2 (N5649, N5646, N1687);
not NOT1 (N5650, N5648);
or OR4 (N5651, N5638, N1223, N4566, N1210);
or OR2 (N5652, N5643, N1705);
or OR4 (N5653, N5652, N4658, N2792, N1524);
and AND3 (N5654, N5649, N3408, N5570);
nand NAND4 (N5655, N5654, N3465, N1934, N4040);
xor XOR2 (N5656, N5645, N3116);
xor XOR2 (N5657, N5637, N4628);
and AND3 (N5658, N5647, N1533, N3820);
and AND2 (N5659, N5640, N121);
and AND3 (N5660, N5621, N930, N2975);
buf BUF1 (N5661, N5657);
xor XOR2 (N5662, N5651, N3665);
and AND4 (N5663, N5658, N4162, N5453, N490);
xor XOR2 (N5664, N5655, N3398);
buf BUF1 (N5665, N5663);
buf BUF1 (N5666, N5656);
not NOT1 (N5667, N5650);
and AND3 (N5668, N5653, N5318, N2895);
not NOT1 (N5669, N5662);
nor NOR3 (N5670, N5661, N2257, N5114);
and AND4 (N5671, N5670, N4577, N2861, N2570);
nor NOR4 (N5672, N5667, N686, N4429, N5516);
nor NOR4 (N5673, N5659, N4280, N3662, N1540);
buf BUF1 (N5674, N5672);
nand NAND4 (N5675, N5666, N3805, N1090, N2431);
nand NAND3 (N5676, N5665, N921, N4465);
nand NAND2 (N5677, N5668, N4893);
not NOT1 (N5678, N5675);
xor XOR2 (N5679, N5673, N1682);
or OR3 (N5680, N5674, N4980, N662);
and AND3 (N5681, N5679, N5444, N4318);
xor XOR2 (N5682, N5669, N2601);
nand NAND2 (N5683, N5644, N1535);
or OR4 (N5684, N5664, N2939, N1581, N2912);
nand NAND3 (N5685, N5680, N2190, N452);
xor XOR2 (N5686, N5678, N1743);
and AND3 (N5687, N5660, N4480, N3218);
buf BUF1 (N5688, N5677);
buf BUF1 (N5689, N5685);
nor NOR3 (N5690, N5671, N3615, N2778);
not NOT1 (N5691, N5687);
and AND2 (N5692, N5686, N5223);
and AND3 (N5693, N5689, N3341, N3713);
or OR4 (N5694, N5684, N1728, N1975, N1026);
xor XOR2 (N5695, N5682, N2249);
nand NAND2 (N5696, N5694, N1546);
or OR4 (N5697, N5688, N1403, N2499, N4993);
nand NAND4 (N5698, N5676, N4821, N3741, N4157);
xor XOR2 (N5699, N5690, N1824);
xor XOR2 (N5700, N5683, N3892);
nand NAND2 (N5701, N5692, N1655);
buf BUF1 (N5702, N5700);
buf BUF1 (N5703, N5697);
xor XOR2 (N5704, N5701, N1208);
nand NAND2 (N5705, N5681, N2012);
or OR3 (N5706, N5698, N513, N3098);
xor XOR2 (N5707, N5691, N4181);
nor NOR2 (N5708, N5706, N3139);
or OR2 (N5709, N5702, N2832);
buf BUF1 (N5710, N5709);
or OR2 (N5711, N5710, N2009);
and AND4 (N5712, N5711, N5614, N1135, N3902);
nand NAND3 (N5713, N5712, N3768, N5592);
xor XOR2 (N5714, N5707, N4624);
nor NOR3 (N5715, N5714, N425, N1810);
buf BUF1 (N5716, N5713);
nor NOR2 (N5717, N5708, N2228);
and AND2 (N5718, N5716, N4473);
nor NOR4 (N5719, N5704, N4490, N1826, N3528);
xor XOR2 (N5720, N5695, N1714);
not NOT1 (N5721, N5720);
xor XOR2 (N5722, N5715, N2793);
nand NAND2 (N5723, N5718, N5405);
nor NOR2 (N5724, N5723, N4134);
xor XOR2 (N5725, N5703, N4556);
buf BUF1 (N5726, N5699);
or OR2 (N5727, N5719, N875);
or OR2 (N5728, N5727, N1798);
or OR3 (N5729, N5722, N5290, N1394);
xor XOR2 (N5730, N5726, N3074);
nor NOR4 (N5731, N5721, N1717, N1870, N362);
and AND2 (N5732, N5730, N3021);
nor NOR3 (N5733, N5717, N973, N64);
xor XOR2 (N5734, N5705, N5422);
or OR2 (N5735, N5729, N1474);
nor NOR2 (N5736, N5731, N4252);
or OR4 (N5737, N5696, N3132, N2065, N4415);
buf BUF1 (N5738, N5728);
nand NAND3 (N5739, N5733, N2528, N4937);
buf BUF1 (N5740, N5736);
buf BUF1 (N5741, N5737);
not NOT1 (N5742, N5725);
not NOT1 (N5743, N5732);
and AND2 (N5744, N5724, N1361);
not NOT1 (N5745, N5743);
nor NOR2 (N5746, N5734, N5228);
and AND2 (N5747, N5740, N3809);
buf BUF1 (N5748, N5735);
and AND2 (N5749, N5739, N5624);
buf BUF1 (N5750, N5742);
nor NOR4 (N5751, N5744, N1195, N5656, N4010);
or OR4 (N5752, N5741, N5420, N4716, N1049);
and AND2 (N5753, N5751, N5002);
not NOT1 (N5754, N5750);
or OR3 (N5755, N5747, N2269, N1319);
xor XOR2 (N5756, N5693, N145);
and AND2 (N5757, N5745, N3266);
or OR2 (N5758, N5738, N3801);
xor XOR2 (N5759, N5748, N5451);
and AND4 (N5760, N5753, N1611, N2239, N4011);
xor XOR2 (N5761, N5759, N4958);
not NOT1 (N5762, N5756);
xor XOR2 (N5763, N5746, N5732);
nand NAND2 (N5764, N5749, N1688);
or OR2 (N5765, N5755, N2022);
buf BUF1 (N5766, N5762);
and AND4 (N5767, N5758, N5166, N1418, N860);
or OR2 (N5768, N5757, N2612);
buf BUF1 (N5769, N5760);
and AND4 (N5770, N5752, N3431, N4997, N1833);
or OR2 (N5771, N5766, N3650);
nand NAND3 (N5772, N5767, N636, N4012);
and AND3 (N5773, N5765, N4037, N818);
and AND4 (N5774, N5770, N4803, N1623, N2689);
nand NAND3 (N5775, N5772, N1196, N740);
xor XOR2 (N5776, N5754, N4021);
xor XOR2 (N5777, N5771, N1312);
and AND3 (N5778, N5768, N2591, N1470);
xor XOR2 (N5779, N5775, N4270);
buf BUF1 (N5780, N5778);
and AND4 (N5781, N5773, N2948, N2815, N1797);
or OR2 (N5782, N5761, N3552);
and AND3 (N5783, N5763, N1008, N3863);
not NOT1 (N5784, N5782);
nor NOR4 (N5785, N5779, N2654, N3361, N1176);
xor XOR2 (N5786, N5776, N1447);
and AND3 (N5787, N5785, N2394, N2724);
not NOT1 (N5788, N5787);
nand NAND3 (N5789, N5777, N2729, N2465);
or OR2 (N5790, N5780, N658);
xor XOR2 (N5791, N5764, N2996);
nand NAND3 (N5792, N5783, N1079, N150);
nor NOR2 (N5793, N5790, N4608);
xor XOR2 (N5794, N5788, N3792);
nor NOR3 (N5795, N5781, N3719, N3728);
buf BUF1 (N5796, N5789);
nor NOR3 (N5797, N5774, N3731, N269);
nor NOR4 (N5798, N5794, N2558, N4113, N4198);
not NOT1 (N5799, N5797);
nand NAND4 (N5800, N5791, N5714, N3635, N4017);
nand NAND2 (N5801, N5786, N2317);
buf BUF1 (N5802, N5769);
not NOT1 (N5803, N5800);
nor NOR3 (N5804, N5795, N2476, N2092);
xor XOR2 (N5805, N5793, N394);
nand NAND4 (N5806, N5804, N4024, N764, N2667);
nand NAND3 (N5807, N5803, N5437, N1353);
and AND4 (N5808, N5798, N1935, N856, N1140);
or OR4 (N5809, N5792, N4090, N3645, N892);
and AND2 (N5810, N5802, N5705);
and AND2 (N5811, N5796, N3793);
and AND3 (N5812, N5801, N1770, N4875);
nor NOR2 (N5813, N5809, N3122);
nor NOR3 (N5814, N5808, N3732, N2942);
or OR3 (N5815, N5811, N2980, N1256);
nand NAND3 (N5816, N5805, N3441, N1401);
and AND3 (N5817, N5806, N3515, N763);
buf BUF1 (N5818, N5813);
not NOT1 (N5819, N5814);
nor NOR3 (N5820, N5819, N321, N938);
or OR2 (N5821, N5815, N156);
buf BUF1 (N5822, N5820);
nand NAND4 (N5823, N5799, N4812, N209, N4330);
and AND2 (N5824, N5784, N5197);
and AND3 (N5825, N5812, N912, N3141);
and AND4 (N5826, N5821, N3668, N1910, N2027);
nand NAND4 (N5827, N5826, N3345, N3706, N180);
xor XOR2 (N5828, N5825, N4058);
xor XOR2 (N5829, N5822, N4994);
buf BUF1 (N5830, N5810);
and AND2 (N5831, N5816, N4781);
not NOT1 (N5832, N5829);
buf BUF1 (N5833, N5832);
xor XOR2 (N5834, N5827, N5364);
not NOT1 (N5835, N5823);
not NOT1 (N5836, N5818);
xor XOR2 (N5837, N5807, N1112);
and AND2 (N5838, N5833, N3090);
or OR3 (N5839, N5828, N2396, N4686);
or OR3 (N5840, N5837, N4082, N2766);
buf BUF1 (N5841, N5835);
nand NAND4 (N5842, N5838, N5386, N3156, N4157);
not NOT1 (N5843, N5839);
buf BUF1 (N5844, N5842);
not NOT1 (N5845, N5836);
nand NAND2 (N5846, N5834, N2133);
or OR2 (N5847, N5830, N1924);
and AND3 (N5848, N5846, N1419, N4452);
nand NAND3 (N5849, N5817, N43, N5078);
xor XOR2 (N5850, N5845, N2763);
and AND4 (N5851, N5840, N2373, N55, N1264);
buf BUF1 (N5852, N5848);
and AND4 (N5853, N5844, N3578, N5768, N4358);
nor NOR3 (N5854, N5852, N4725, N5664);
nand NAND2 (N5855, N5854, N1414);
not NOT1 (N5856, N5847);
nor NOR2 (N5857, N5850, N5289);
nand NAND3 (N5858, N5824, N4863, N2237);
not NOT1 (N5859, N5841);
buf BUF1 (N5860, N5843);
nand NAND3 (N5861, N5858, N2297, N5192);
and AND3 (N5862, N5855, N1676, N234);
nand NAND4 (N5863, N5853, N5164, N5763, N4848);
buf BUF1 (N5864, N5860);
or OR2 (N5865, N5851, N2985);
or OR2 (N5866, N5861, N2540);
or OR4 (N5867, N5864, N1141, N1941, N1920);
not NOT1 (N5868, N5831);
nand NAND4 (N5869, N5866, N399, N3588, N4220);
xor XOR2 (N5870, N5849, N4591);
nor NOR3 (N5871, N5857, N935, N4918);
not NOT1 (N5872, N5868);
xor XOR2 (N5873, N5856, N1120);
xor XOR2 (N5874, N5871, N3328);
nand NAND3 (N5875, N5873, N5483, N3108);
or OR2 (N5876, N5872, N1388);
nand NAND3 (N5877, N5870, N1142, N5121);
nor NOR2 (N5878, N5865, N5662);
and AND4 (N5879, N5874, N2915, N5288, N1928);
buf BUF1 (N5880, N5878);
not NOT1 (N5881, N5869);
not NOT1 (N5882, N5877);
nand NAND3 (N5883, N5881, N1125, N5076);
or OR3 (N5884, N5883, N4447, N5255);
nand NAND4 (N5885, N5875, N3681, N1557, N3465);
nor NOR4 (N5886, N5880, N2222, N1406, N570);
nor NOR4 (N5887, N5862, N2434, N2298, N2718);
or OR4 (N5888, N5885, N5321, N1988, N965);
nand NAND2 (N5889, N5867, N3363);
and AND2 (N5890, N5886, N3881);
nand NAND2 (N5891, N5884, N156);
nor NOR3 (N5892, N5879, N610, N169);
or OR4 (N5893, N5876, N4985, N4101, N3635);
buf BUF1 (N5894, N5882);
and AND3 (N5895, N5859, N1865, N1590);
or OR3 (N5896, N5894, N1190, N1825);
buf BUF1 (N5897, N5889);
or OR3 (N5898, N5892, N4526, N276);
buf BUF1 (N5899, N5893);
nand NAND2 (N5900, N5898, N3541);
buf BUF1 (N5901, N5863);
xor XOR2 (N5902, N5895, N5032);
buf BUF1 (N5903, N5891);
not NOT1 (N5904, N5887);
buf BUF1 (N5905, N5902);
and AND4 (N5906, N5901, N3916, N4631, N3592);
and AND4 (N5907, N5890, N325, N2349, N2226);
nand NAND2 (N5908, N5906, N5501);
not NOT1 (N5909, N5896);
or OR2 (N5910, N5907, N3066);
not NOT1 (N5911, N5904);
buf BUF1 (N5912, N5900);
buf BUF1 (N5913, N5903);
xor XOR2 (N5914, N5905, N214);
or OR4 (N5915, N5913, N5280, N3823, N73);
buf BUF1 (N5916, N5915);
nand NAND2 (N5917, N5909, N4752);
buf BUF1 (N5918, N5917);
or OR2 (N5919, N5911, N770);
xor XOR2 (N5920, N5888, N4346);
not NOT1 (N5921, N5916);
nor NOR3 (N5922, N5899, N1871, N419);
buf BUF1 (N5923, N5897);
buf BUF1 (N5924, N5922);
or OR4 (N5925, N5914, N2512, N4440, N3863);
nand NAND3 (N5926, N5925, N4293, N4838);
nor NOR2 (N5927, N5912, N5231);
not NOT1 (N5928, N5923);
and AND4 (N5929, N5924, N591, N3087, N2014);
buf BUF1 (N5930, N5920);
nor NOR4 (N5931, N5927, N1832, N3850, N200);
and AND4 (N5932, N5908, N249, N4890, N3569);
not NOT1 (N5933, N5931);
buf BUF1 (N5934, N5932);
and AND4 (N5935, N5910, N2761, N4163, N1300);
not NOT1 (N5936, N5934);
and AND3 (N5937, N5926, N1610, N5396);
nor NOR4 (N5938, N5937, N4092, N1642, N1781);
or OR3 (N5939, N5929, N5691, N3726);
not NOT1 (N5940, N5939);
nor NOR2 (N5941, N5918, N5167);
nor NOR2 (N5942, N5938, N1746);
not NOT1 (N5943, N5930);
not NOT1 (N5944, N5921);
nand NAND2 (N5945, N5919, N1836);
nor NOR3 (N5946, N5936, N1447, N5420);
nand NAND2 (N5947, N5940, N5080);
or OR4 (N5948, N5942, N2178, N3072, N75);
xor XOR2 (N5949, N5933, N2577);
nand NAND3 (N5950, N5944, N397, N5406);
nor NOR3 (N5951, N5943, N3812, N600);
xor XOR2 (N5952, N5951, N984);
nor NOR3 (N5953, N5928, N4060, N764);
nor NOR2 (N5954, N5947, N136);
nand NAND2 (N5955, N5948, N2748);
nor NOR4 (N5956, N5952, N5692, N5610, N5728);
nor NOR3 (N5957, N5949, N3269, N676);
or OR2 (N5958, N5957, N4208);
not NOT1 (N5959, N5945);
nor NOR3 (N5960, N5946, N3646, N2566);
buf BUF1 (N5961, N5958);
not NOT1 (N5962, N5955);
and AND2 (N5963, N5962, N107);
and AND3 (N5964, N5941, N312, N4577);
buf BUF1 (N5965, N5964);
xor XOR2 (N5966, N5954, N2400);
nor NOR4 (N5967, N5956, N4305, N135, N5085);
buf BUF1 (N5968, N5966);
and AND4 (N5969, N5967, N3868, N2519, N5855);
and AND4 (N5970, N5960, N466, N4343, N4398);
and AND3 (N5971, N5961, N1468, N958);
or OR4 (N5972, N5950, N1480, N1006, N690);
nand NAND2 (N5973, N5972, N1651);
xor XOR2 (N5974, N5970, N2466);
nand NAND3 (N5975, N5959, N5085, N369);
nand NAND2 (N5976, N5969, N2633);
xor XOR2 (N5977, N5975, N4349);
not NOT1 (N5978, N5963);
and AND3 (N5979, N5974, N3596, N235);
nand NAND4 (N5980, N5971, N147, N1682, N4964);
nand NAND4 (N5981, N5973, N5967, N256, N599);
not NOT1 (N5982, N5935);
not NOT1 (N5983, N5977);
or OR3 (N5984, N5983, N3615, N3073);
nand NAND2 (N5985, N5968, N4501);
xor XOR2 (N5986, N5976, N1181);
and AND3 (N5987, N5980, N2108, N5459);
nand NAND2 (N5988, N5978, N3637);
buf BUF1 (N5989, N5979);
and AND4 (N5990, N5985, N557, N394, N2355);
buf BUF1 (N5991, N5981);
nor NOR2 (N5992, N5991, N1348);
and AND4 (N5993, N5989, N1394, N1423, N3264);
not NOT1 (N5994, N5993);
xor XOR2 (N5995, N5988, N43);
and AND2 (N5996, N5995, N4438);
buf BUF1 (N5997, N5994);
nand NAND2 (N5998, N5986, N5991);
nand NAND3 (N5999, N5953, N3127, N1415);
buf BUF1 (N6000, N5987);
and AND2 (N6001, N5984, N865);
not NOT1 (N6002, N5992);
buf BUF1 (N6003, N5998);
and AND4 (N6004, N5990, N3730, N3632, N5055);
buf BUF1 (N6005, N5999);
not NOT1 (N6006, N5996);
buf BUF1 (N6007, N6001);
xor XOR2 (N6008, N6003, N3504);
xor XOR2 (N6009, N6006, N4176);
or OR2 (N6010, N6009, N1521);
nor NOR2 (N6011, N6008, N2444);
nor NOR3 (N6012, N6005, N4491, N1720);
nand NAND3 (N6013, N6007, N1047, N62);
buf BUF1 (N6014, N6002);
not NOT1 (N6015, N6011);
buf BUF1 (N6016, N6004);
buf BUF1 (N6017, N5965);
buf BUF1 (N6018, N6016);
nor NOR3 (N6019, N5997, N4661, N1512);
not NOT1 (N6020, N5982);
nand NAND3 (N6021, N6018, N3376, N4085);
not NOT1 (N6022, N6000);
nand NAND4 (N6023, N6019, N5327, N3959, N4543);
or OR2 (N6024, N6013, N1580);
and AND4 (N6025, N6012, N896, N2617, N2652);
nor NOR4 (N6026, N6017, N1010, N2880, N5744);
not NOT1 (N6027, N6021);
xor XOR2 (N6028, N6022, N4188);
nor NOR2 (N6029, N6014, N4689);
buf BUF1 (N6030, N6024);
xor XOR2 (N6031, N6025, N1194);
xor XOR2 (N6032, N6020, N513);
xor XOR2 (N6033, N6027, N594);
xor XOR2 (N6034, N6030, N1726);
xor XOR2 (N6035, N6029, N2305);
and AND3 (N6036, N6033, N5379, N578);
not NOT1 (N6037, N6028);
or OR4 (N6038, N6034, N2370, N232, N2566);
not NOT1 (N6039, N6010);
nand NAND2 (N6040, N6032, N3236);
and AND3 (N6041, N6039, N874, N4236);
and AND4 (N6042, N6031, N1411, N4545, N4058);
buf BUF1 (N6043, N6026);
buf BUF1 (N6044, N6043);
or OR2 (N6045, N6035, N2798);
and AND2 (N6046, N6038, N2710);
and AND3 (N6047, N6044, N2033, N2919);
or OR3 (N6048, N6023, N4585, N2612);
nor NOR3 (N6049, N6047, N4051, N4914);
or OR4 (N6050, N6041, N1684, N1889, N5044);
buf BUF1 (N6051, N6045);
nand NAND4 (N6052, N6042, N4, N608, N1791);
not NOT1 (N6053, N6048);
and AND3 (N6054, N6050, N1661, N3595);
buf BUF1 (N6055, N6015);
and AND4 (N6056, N6054, N4955, N3495, N4274);
nand NAND3 (N6057, N6051, N1856, N2818);
and AND2 (N6058, N6046, N1118);
or OR3 (N6059, N6040, N4670, N3329);
not NOT1 (N6060, N6055);
nor NOR4 (N6061, N6057, N358, N5961, N5820);
or OR4 (N6062, N6053, N4469, N1698, N4338);
and AND2 (N6063, N6036, N213);
not NOT1 (N6064, N6059);
buf BUF1 (N6065, N6037);
xor XOR2 (N6066, N6065, N1004);
nand NAND2 (N6067, N6056, N2758);
nand NAND3 (N6068, N6061, N3598, N3627);
or OR3 (N6069, N6062, N2625, N3527);
or OR2 (N6070, N6060, N1701);
and AND4 (N6071, N6064, N3940, N4187, N4696);
nand NAND3 (N6072, N6063, N2667, N455);
xor XOR2 (N6073, N6058, N2444);
nor NOR3 (N6074, N6070, N3707, N2790);
buf BUF1 (N6075, N6052);
nor NOR3 (N6076, N6067, N3185, N478);
buf BUF1 (N6077, N6073);
buf BUF1 (N6078, N6077);
or OR3 (N6079, N6049, N3196, N1958);
and AND2 (N6080, N6071, N5066);
and AND2 (N6081, N6079, N5960);
buf BUF1 (N6082, N6074);
xor XOR2 (N6083, N6069, N2110);
and AND2 (N6084, N6081, N446);
xor XOR2 (N6085, N6076, N4325);
and AND2 (N6086, N6075, N2063);
xor XOR2 (N6087, N6083, N1841);
nor NOR2 (N6088, N6082, N3064);
nor NOR4 (N6089, N6066, N3793, N5370, N1635);
not NOT1 (N6090, N6086);
nand NAND2 (N6091, N6085, N5900);
xor XOR2 (N6092, N6087, N3703);
not NOT1 (N6093, N6091);
or OR4 (N6094, N6068, N2073, N5054, N4797);
xor XOR2 (N6095, N6078, N3396);
and AND4 (N6096, N6089, N992, N1579, N5323);
nand NAND4 (N6097, N6088, N826, N165, N3572);
xor XOR2 (N6098, N6090, N5544);
or OR3 (N6099, N6080, N3309, N4805);
or OR4 (N6100, N6094, N1720, N6014, N2349);
or OR4 (N6101, N6072, N4952, N2559, N5367);
not NOT1 (N6102, N6084);
nor NOR4 (N6103, N6101, N5793, N4665, N1454);
buf BUF1 (N6104, N6098);
not NOT1 (N6105, N6100);
xor XOR2 (N6106, N6099, N392);
xor XOR2 (N6107, N6092, N2860);
nor NOR2 (N6108, N6095, N5762);
nand NAND3 (N6109, N6093, N2146, N4318);
and AND3 (N6110, N6103, N1097, N5943);
nor NOR4 (N6111, N6109, N2051, N4734, N5576);
nand NAND4 (N6112, N6096, N5056, N1196, N1847);
nor NOR3 (N6113, N6110, N2079, N3705);
nand NAND4 (N6114, N6106, N5418, N453, N3832);
nor NOR3 (N6115, N6114, N2700, N5022);
nand NAND2 (N6116, N6102, N1549);
xor XOR2 (N6117, N6105, N5845);
or OR4 (N6118, N6116, N4118, N2411, N482);
not NOT1 (N6119, N6104);
xor XOR2 (N6120, N6119, N4949);
buf BUF1 (N6121, N6111);
nor NOR2 (N6122, N6113, N3047);
xor XOR2 (N6123, N6118, N4369);
and AND2 (N6124, N6121, N5007);
or OR2 (N6125, N6107, N1091);
nor NOR2 (N6126, N6108, N5081);
and AND2 (N6127, N6120, N2263);
xor XOR2 (N6128, N6097, N228);
not NOT1 (N6129, N6125);
not NOT1 (N6130, N6115);
and AND3 (N6131, N6112, N508, N509);
nor NOR2 (N6132, N6122, N3286);
nand NAND4 (N6133, N6131, N5399, N652, N3390);
xor XOR2 (N6134, N6124, N4412);
nor NOR3 (N6135, N6129, N4880, N2908);
and AND4 (N6136, N6127, N3665, N946, N4752);
nor NOR2 (N6137, N6132, N2116);
buf BUF1 (N6138, N6137);
buf BUF1 (N6139, N6123);
and AND4 (N6140, N6135, N4293, N3802, N4002);
and AND3 (N6141, N6133, N4640, N667);
nor NOR4 (N6142, N6128, N2270, N2191, N1234);
buf BUF1 (N6143, N6126);
and AND4 (N6144, N6143, N3685, N5532, N6131);
nor NOR3 (N6145, N6144, N5770, N2158);
xor XOR2 (N6146, N6141, N2248);
buf BUF1 (N6147, N6117);
not NOT1 (N6148, N6145);
not NOT1 (N6149, N6142);
nor NOR2 (N6150, N6140, N3107);
buf BUF1 (N6151, N6148);
not NOT1 (N6152, N6138);
nor NOR2 (N6153, N6146, N4274);
buf BUF1 (N6154, N6151);
nor NOR2 (N6155, N6153, N81);
buf BUF1 (N6156, N6139);
not NOT1 (N6157, N6147);
buf BUF1 (N6158, N6152);
not NOT1 (N6159, N6157);
nor NOR4 (N6160, N6150, N2293, N4570, N2626);
or OR4 (N6161, N6160, N1367, N6142, N2222);
or OR4 (N6162, N6136, N5107, N1205, N3436);
and AND4 (N6163, N6159, N5384, N1025, N5590);
buf BUF1 (N6164, N6134);
buf BUF1 (N6165, N6130);
nand NAND3 (N6166, N6163, N3698, N3701);
and AND2 (N6167, N6158, N2702);
buf BUF1 (N6168, N6162);
and AND3 (N6169, N6154, N4050, N2200);
and AND4 (N6170, N6161, N5409, N1332, N4292);
not NOT1 (N6171, N6167);
not NOT1 (N6172, N6149);
nand NAND2 (N6173, N6169, N2722);
and AND4 (N6174, N6164, N5402, N6141, N2810);
nor NOR3 (N6175, N6173, N478, N5823);
nand NAND2 (N6176, N6170, N3739);
nor NOR4 (N6177, N6174, N5200, N2819, N1041);
nor NOR4 (N6178, N6165, N1413, N3713, N4389);
nand NAND2 (N6179, N6172, N5481);
xor XOR2 (N6180, N6155, N3307);
xor XOR2 (N6181, N6156, N587);
or OR3 (N6182, N6166, N2380, N5083);
or OR4 (N6183, N6175, N5213, N3585, N6056);
or OR2 (N6184, N6181, N1460);
not NOT1 (N6185, N6179);
and AND4 (N6186, N6183, N4929, N657, N1668);
nand NAND3 (N6187, N6184, N1328, N4665);
xor XOR2 (N6188, N6182, N4672);
and AND3 (N6189, N6186, N5116, N1300);
or OR2 (N6190, N6168, N5320);
nor NOR3 (N6191, N6189, N3903, N951);
or OR2 (N6192, N6191, N2234);
nor NOR3 (N6193, N6187, N2684, N622);
xor XOR2 (N6194, N6192, N3602);
not NOT1 (N6195, N6171);
not NOT1 (N6196, N6177);
not NOT1 (N6197, N6180);
nor NOR4 (N6198, N6194, N3156, N2337, N2494);
xor XOR2 (N6199, N6197, N2048);
buf BUF1 (N6200, N6199);
not NOT1 (N6201, N6190);
and AND3 (N6202, N6178, N3244, N1019);
buf BUF1 (N6203, N6200);
not NOT1 (N6204, N6202);
nand NAND4 (N6205, N6195, N5206, N815, N568);
nand NAND3 (N6206, N6176, N1936, N2846);
nand NAND3 (N6207, N6205, N1126, N4226);
buf BUF1 (N6208, N6198);
not NOT1 (N6209, N6188);
and AND2 (N6210, N6201, N5097);
and AND4 (N6211, N6203, N2090, N3721, N1791);
and AND4 (N6212, N6204, N794, N3272, N2906);
not NOT1 (N6213, N6212);
xor XOR2 (N6214, N6207, N266);
nor NOR2 (N6215, N6213, N196);
not NOT1 (N6216, N6211);
nand NAND2 (N6217, N6206, N4950);
xor XOR2 (N6218, N6209, N4527);
and AND2 (N6219, N6218, N671);
not NOT1 (N6220, N6219);
buf BUF1 (N6221, N6220);
xor XOR2 (N6222, N6193, N4771);
xor XOR2 (N6223, N6196, N5501);
and AND2 (N6224, N6216, N1183);
nand NAND2 (N6225, N6214, N5214);
not NOT1 (N6226, N6185);
or OR4 (N6227, N6224, N1878, N6149, N1054);
not NOT1 (N6228, N6208);
not NOT1 (N6229, N6217);
and AND4 (N6230, N6210, N2792, N1917, N5727);
not NOT1 (N6231, N6222);
xor XOR2 (N6232, N6229, N462);
nor NOR2 (N6233, N6231, N1840);
nand NAND4 (N6234, N6233, N5675, N4319, N1085);
buf BUF1 (N6235, N6223);
buf BUF1 (N6236, N6227);
nand NAND2 (N6237, N6232, N5312);
not NOT1 (N6238, N6237);
buf BUF1 (N6239, N6225);
xor XOR2 (N6240, N6228, N3326);
and AND2 (N6241, N6230, N5924);
not NOT1 (N6242, N6239);
and AND2 (N6243, N6226, N6170);
nor NOR2 (N6244, N6242, N6198);
nand NAND3 (N6245, N6241, N811, N237);
or OR3 (N6246, N6244, N984, N684);
and AND3 (N6247, N6236, N1004, N1060);
nor NOR3 (N6248, N6238, N941, N5785);
and AND2 (N6249, N6240, N2718);
not NOT1 (N6250, N6249);
nand NAND4 (N6251, N6221, N1825, N347, N1384);
and AND4 (N6252, N6215, N5208, N1608, N4045);
and AND3 (N6253, N6247, N3884, N713);
not NOT1 (N6254, N6235);
or OR3 (N6255, N6234, N2087, N4551);
nor NOR3 (N6256, N6243, N5209, N5404);
and AND2 (N6257, N6256, N5634);
and AND4 (N6258, N6254, N1436, N4334, N2815);
not NOT1 (N6259, N6246);
nand NAND3 (N6260, N6251, N3064, N661);
buf BUF1 (N6261, N6260);
or OR2 (N6262, N6261, N3495);
nor NOR4 (N6263, N6255, N2424, N5438, N2105);
nand NAND2 (N6264, N6253, N5856);
nand NAND3 (N6265, N6248, N2488, N1924);
xor XOR2 (N6266, N6250, N4194);
nor NOR3 (N6267, N6265, N1056, N1953);
nand NAND2 (N6268, N6262, N4659);
nand NAND3 (N6269, N6252, N5313, N1870);
nor NOR3 (N6270, N6264, N3127, N3172);
xor XOR2 (N6271, N6266, N1307);
or OR3 (N6272, N6259, N4161, N333);
nand NAND2 (N6273, N6245, N748);
nor NOR3 (N6274, N6270, N3814, N5089);
or OR2 (N6275, N6257, N2330);
not NOT1 (N6276, N6274);
xor XOR2 (N6277, N6275, N1326);
buf BUF1 (N6278, N6258);
nand NAND2 (N6279, N6269, N4604);
or OR2 (N6280, N6277, N2143);
not NOT1 (N6281, N6279);
buf BUF1 (N6282, N6276);
not NOT1 (N6283, N6271);
and AND4 (N6284, N6263, N3136, N5623, N1495);
buf BUF1 (N6285, N6282);
or OR2 (N6286, N6283, N459);
xor XOR2 (N6287, N6280, N5859);
nor NOR3 (N6288, N6285, N5142, N1566);
nor NOR2 (N6289, N6272, N4166);
nand NAND3 (N6290, N6284, N2562, N1142);
nand NAND3 (N6291, N6281, N3211, N1727);
and AND2 (N6292, N6278, N2878);
or OR2 (N6293, N6273, N2668);
and AND2 (N6294, N6291, N5411);
buf BUF1 (N6295, N6290);
and AND4 (N6296, N6288, N904, N4085, N2485);
nand NAND2 (N6297, N6286, N4479);
xor XOR2 (N6298, N6292, N4175);
nand NAND3 (N6299, N6267, N3477, N6106);
xor XOR2 (N6300, N6289, N5702);
buf BUF1 (N6301, N6298);
not NOT1 (N6302, N6287);
xor XOR2 (N6303, N6297, N3786);
nor NOR2 (N6304, N6268, N4490);
not NOT1 (N6305, N6300);
not NOT1 (N6306, N6299);
nand NAND2 (N6307, N6301, N6142);
buf BUF1 (N6308, N6306);
and AND3 (N6309, N6304, N2485, N2146);
buf BUF1 (N6310, N6294);
nor NOR4 (N6311, N6309, N6157, N168, N5557);
not NOT1 (N6312, N6302);
and AND3 (N6313, N6308, N2315, N3377);
nand NAND4 (N6314, N6307, N707, N5085, N680);
or OR4 (N6315, N6293, N4733, N194, N5242);
nand NAND3 (N6316, N6305, N4200, N2408);
buf BUF1 (N6317, N6315);
and AND2 (N6318, N6314, N3199);
and AND3 (N6319, N6295, N4869, N1900);
or OR3 (N6320, N6311, N3866, N3966);
xor XOR2 (N6321, N6312, N2068);
nor NOR3 (N6322, N6303, N4864, N4258);
buf BUF1 (N6323, N6316);
xor XOR2 (N6324, N6313, N5291);
and AND4 (N6325, N6319, N2883, N5144, N31);
nand NAND3 (N6326, N6318, N5465, N2959);
nor NOR4 (N6327, N6326, N1163, N3028, N4539);
xor XOR2 (N6328, N6317, N2145);
and AND2 (N6329, N6325, N3448);
or OR4 (N6330, N6296, N3755, N194, N3002);
nor NOR4 (N6331, N6327, N3179, N4247, N4227);
nor NOR3 (N6332, N6320, N1335, N3653);
and AND4 (N6333, N6323, N5526, N2882, N3375);
or OR4 (N6334, N6324, N3191, N4975, N646);
and AND3 (N6335, N6321, N1623, N6140);
nor NOR2 (N6336, N6328, N1056);
nor NOR2 (N6337, N6331, N2948);
buf BUF1 (N6338, N6330);
nor NOR4 (N6339, N6334, N915, N5954, N3772);
nand NAND2 (N6340, N6329, N1332);
buf BUF1 (N6341, N6333);
nor NOR4 (N6342, N6335, N5104, N1821, N795);
not NOT1 (N6343, N6340);
and AND4 (N6344, N6332, N3467, N3915, N1630);
or OR3 (N6345, N6342, N3186, N2095);
buf BUF1 (N6346, N6310);
not NOT1 (N6347, N6339);
nor NOR4 (N6348, N6341, N2036, N2027, N3885);
buf BUF1 (N6349, N6322);
nor NOR3 (N6350, N6348, N4059, N372);
and AND2 (N6351, N6344, N3726);
or OR4 (N6352, N6343, N6016, N3292, N2237);
nand NAND2 (N6353, N6352, N4242);
or OR3 (N6354, N6350, N2959, N696);
xor XOR2 (N6355, N6336, N4556);
nor NOR2 (N6356, N6346, N4310);
xor XOR2 (N6357, N6338, N2780);
not NOT1 (N6358, N6345);
not NOT1 (N6359, N6358);
nand NAND3 (N6360, N6353, N6048, N5581);
buf BUF1 (N6361, N6360);
nor NOR3 (N6362, N6356, N2857, N3924);
not NOT1 (N6363, N6349);
nand NAND4 (N6364, N6347, N6168, N2864, N163);
buf BUF1 (N6365, N6354);
not NOT1 (N6366, N6364);
and AND2 (N6367, N6362, N3981);
not NOT1 (N6368, N6366);
and AND3 (N6369, N6368, N110, N6261);
xor XOR2 (N6370, N6351, N897);
buf BUF1 (N6371, N6365);
nor NOR4 (N6372, N6363, N5409, N3593, N1418);
buf BUF1 (N6373, N6371);
xor XOR2 (N6374, N6369, N101);
or OR4 (N6375, N6357, N4214, N974, N3251);
xor XOR2 (N6376, N6337, N5216);
buf BUF1 (N6377, N6375);
not NOT1 (N6378, N6376);
xor XOR2 (N6379, N6361, N1165);
nor NOR4 (N6380, N6378, N5233, N1359, N626);
not NOT1 (N6381, N6373);
xor XOR2 (N6382, N6370, N2024);
not NOT1 (N6383, N6355);
or OR2 (N6384, N6367, N6037);
nand NAND2 (N6385, N6372, N5156);
and AND4 (N6386, N6359, N2396, N2224, N2074);
and AND3 (N6387, N6377, N4922, N3787);
nor NOR4 (N6388, N6385, N2743, N5052, N556);
or OR4 (N6389, N6388, N4411, N5398, N1395);
nor NOR2 (N6390, N6382, N2869);
and AND2 (N6391, N6387, N2012);
nand NAND3 (N6392, N6390, N3380, N1856);
nand NAND3 (N6393, N6392, N4606, N3753);
and AND2 (N6394, N6391, N3264);
xor XOR2 (N6395, N6379, N3071);
not NOT1 (N6396, N6380);
xor XOR2 (N6397, N6389, N1221);
and AND4 (N6398, N6384, N3465, N5757, N1764);
buf BUF1 (N6399, N6395);
nor NOR4 (N6400, N6386, N5795, N2251, N3057);
and AND4 (N6401, N6398, N3631, N788, N5618);
not NOT1 (N6402, N6400);
and AND4 (N6403, N6397, N4152, N1071, N745);
nand NAND2 (N6404, N6374, N2247);
not NOT1 (N6405, N6401);
not NOT1 (N6406, N6396);
xor XOR2 (N6407, N6393, N190);
not NOT1 (N6408, N6404);
and AND4 (N6409, N6394, N4687, N4433, N6154);
and AND3 (N6410, N6408, N3353, N1607);
nor NOR4 (N6411, N6406, N5613, N979, N4748);
buf BUF1 (N6412, N6405);
xor XOR2 (N6413, N6399, N2181);
not NOT1 (N6414, N6410);
nor NOR3 (N6415, N6381, N1693, N5973);
nand NAND3 (N6416, N6407, N3575, N278);
xor XOR2 (N6417, N6415, N3063);
and AND4 (N6418, N6413, N1355, N261, N3746);
or OR2 (N6419, N6416, N2799);
buf BUF1 (N6420, N6383);
or OR2 (N6421, N6403, N1674);
nor NOR3 (N6422, N6419, N652, N3729);
not NOT1 (N6423, N6414);
xor XOR2 (N6424, N6409, N256);
xor XOR2 (N6425, N6424, N5918);
nor NOR3 (N6426, N6412, N2086, N5427);
or OR4 (N6427, N6418, N4668, N2879, N1845);
xor XOR2 (N6428, N6417, N3158);
buf BUF1 (N6429, N6411);
xor XOR2 (N6430, N6429, N1036);
and AND4 (N6431, N6402, N946, N6337, N2304);
or OR3 (N6432, N6428, N2679, N360);
nor NOR2 (N6433, N6431, N4697);
not NOT1 (N6434, N6423);
nor NOR4 (N6435, N6426, N5395, N1210, N1538);
nor NOR3 (N6436, N6434, N4044, N3595);
nor NOR4 (N6437, N6435, N739, N4932, N5436);
nand NAND2 (N6438, N6430, N4247);
not NOT1 (N6439, N6427);
buf BUF1 (N6440, N6433);
xor XOR2 (N6441, N6432, N4415);
xor XOR2 (N6442, N6420, N3460);
or OR4 (N6443, N6436, N2785, N4777, N1963);
and AND2 (N6444, N6437, N371);
xor XOR2 (N6445, N6438, N4033);
nand NAND3 (N6446, N6421, N5240, N5902);
buf BUF1 (N6447, N6446);
nor NOR3 (N6448, N6440, N2092, N3470);
not NOT1 (N6449, N6447);
xor XOR2 (N6450, N6422, N535);
nor NOR3 (N6451, N6439, N3851, N2683);
xor XOR2 (N6452, N6444, N4028);
and AND4 (N6453, N6450, N609, N3073, N5422);
xor XOR2 (N6454, N6449, N1012);
xor XOR2 (N6455, N6451, N4389);
not NOT1 (N6456, N6445);
or OR3 (N6457, N6455, N3680, N1916);
or OR2 (N6458, N6448, N3810);
and AND2 (N6459, N6443, N5854);
xor XOR2 (N6460, N6452, N4628);
or OR2 (N6461, N6454, N637);
not NOT1 (N6462, N6460);
and AND4 (N6463, N6441, N3727, N446, N4733);
xor XOR2 (N6464, N6456, N877);
not NOT1 (N6465, N6457);
not NOT1 (N6466, N6461);
nand NAND3 (N6467, N6442, N5072, N2927);
nand NAND3 (N6468, N6464, N396, N1748);
and AND4 (N6469, N6425, N512, N401, N725);
buf BUF1 (N6470, N6453);
or OR4 (N6471, N6469, N5493, N209, N4510);
or OR4 (N6472, N6465, N1509, N2581, N1153);
xor XOR2 (N6473, N6462, N4929);
nand NAND4 (N6474, N6468, N918, N3181, N809);
xor XOR2 (N6475, N6474, N1027);
nand NAND3 (N6476, N6458, N4798, N1034);
or OR2 (N6477, N6463, N3511);
or OR4 (N6478, N6473, N2335, N695, N2450);
and AND3 (N6479, N6476, N4035, N6214);
or OR3 (N6480, N6467, N590, N5022);
nor NOR4 (N6481, N6459, N2855, N1113, N4096);
nand NAND3 (N6482, N6480, N3489, N1848);
buf BUF1 (N6483, N6481);
buf BUF1 (N6484, N6478);
not NOT1 (N6485, N6479);
nor NOR3 (N6486, N6472, N1534, N4901);
xor XOR2 (N6487, N6486, N3149);
buf BUF1 (N6488, N6477);
and AND2 (N6489, N6471, N2856);
buf BUF1 (N6490, N6489);
and AND3 (N6491, N6483, N3391, N2333);
nand NAND4 (N6492, N6466, N4765, N3171, N730);
nor NOR4 (N6493, N6488, N6162, N2029, N3257);
not NOT1 (N6494, N6482);
nand NAND4 (N6495, N6484, N3650, N5159, N6453);
not NOT1 (N6496, N6493);
or OR4 (N6497, N6475, N439, N4413, N2161);
not NOT1 (N6498, N6490);
nand NAND3 (N6499, N6498, N1776, N302);
and AND2 (N6500, N6487, N3743);
xor XOR2 (N6501, N6500, N2258);
and AND4 (N6502, N6495, N3424, N2756, N5081);
not NOT1 (N6503, N6491);
nand NAND3 (N6504, N6502, N3236, N169);
buf BUF1 (N6505, N6470);
xor XOR2 (N6506, N6505, N2237);
and AND4 (N6507, N6499, N1978, N4870, N4049);
buf BUF1 (N6508, N6506);
nor NOR3 (N6509, N6503, N5225, N4894);
buf BUF1 (N6510, N6492);
buf BUF1 (N6511, N6497);
xor XOR2 (N6512, N6501, N2610);
or OR2 (N6513, N6508, N505);
buf BUF1 (N6514, N6510);
and AND4 (N6515, N6514, N3761, N1565, N5934);
nand NAND3 (N6516, N6515, N2830, N4528);
nand NAND4 (N6517, N6512, N1110, N1443, N4958);
and AND2 (N6518, N6516, N5724);
not NOT1 (N6519, N6494);
nand NAND3 (N6520, N6485, N4209, N6400);
and AND3 (N6521, N6511, N3968, N525);
and AND2 (N6522, N6518, N449);
or OR3 (N6523, N6509, N540, N232);
and AND4 (N6524, N6521, N4332, N2516, N869);
xor XOR2 (N6525, N6517, N5652);
buf BUF1 (N6526, N6504);
nand NAND2 (N6527, N6507, N4705);
or OR2 (N6528, N6522, N4787);
xor XOR2 (N6529, N6523, N4617);
or OR3 (N6530, N6528, N3554, N1343);
nor NOR3 (N6531, N6526, N2735, N2631);
and AND4 (N6532, N6520, N2340, N2291, N1417);
xor XOR2 (N6533, N6513, N125);
nand NAND4 (N6534, N6524, N597, N2814, N5223);
or OR3 (N6535, N6530, N637, N3859);
not NOT1 (N6536, N6496);
or OR4 (N6537, N6525, N3824, N2580, N4726);
nor NOR2 (N6538, N6531, N712);
nor NOR3 (N6539, N6519, N1374, N3190);
nand NAND2 (N6540, N6536, N1182);
and AND4 (N6541, N6529, N6129, N962, N6253);
or OR4 (N6542, N6537, N3096, N4628, N396);
nor NOR4 (N6543, N6534, N4764, N4057, N5871);
xor XOR2 (N6544, N6535, N1915);
or OR3 (N6545, N6539, N5882, N1289);
nand NAND4 (N6546, N6532, N3468, N960, N5728);
not NOT1 (N6547, N6538);
or OR2 (N6548, N6542, N1869);
or OR3 (N6549, N6544, N2940, N5945);
buf BUF1 (N6550, N6549);
nand NAND3 (N6551, N6546, N4478, N3170);
or OR4 (N6552, N6545, N2232, N3530, N3501);
xor XOR2 (N6553, N6550, N488);
or OR4 (N6554, N6527, N961, N5755, N5967);
not NOT1 (N6555, N6547);
nand NAND3 (N6556, N6541, N2149, N795);
and AND3 (N6557, N6533, N685, N1957);
nand NAND2 (N6558, N6551, N2826);
nor NOR2 (N6559, N6553, N3096);
nand NAND4 (N6560, N6548, N865, N4150, N2962);
nand NAND3 (N6561, N6560, N1417, N3508);
nand NAND4 (N6562, N6543, N4523, N584, N155);
buf BUF1 (N6563, N6556);
xor XOR2 (N6564, N6557, N2396);
and AND3 (N6565, N6558, N2674, N656);
not NOT1 (N6566, N6540);
nor NOR3 (N6567, N6566, N5248, N2144);
nor NOR3 (N6568, N6563, N791, N1294);
nand NAND2 (N6569, N6567, N4045);
nor NOR4 (N6570, N6562, N3071, N3725, N6493);
xor XOR2 (N6571, N6569, N4560);
nand NAND4 (N6572, N6555, N3478, N4952, N3547);
xor XOR2 (N6573, N6554, N1344);
nor NOR3 (N6574, N6565, N1973, N937);
xor XOR2 (N6575, N6571, N4965);
and AND3 (N6576, N6573, N5320, N3997);
buf BUF1 (N6577, N6576);
and AND2 (N6578, N6568, N1202);
not NOT1 (N6579, N6561);
buf BUF1 (N6580, N6579);
buf BUF1 (N6581, N6574);
and AND3 (N6582, N6552, N1861, N147);
or OR4 (N6583, N6582, N681, N4730, N4441);
nand NAND3 (N6584, N6578, N909, N3977);
nor NOR3 (N6585, N6577, N3466, N5366);
not NOT1 (N6586, N6559);
nand NAND2 (N6587, N6583, N2243);
nand NAND4 (N6588, N6585, N5663, N3054, N2182);
nor NOR2 (N6589, N6581, N275);
nand NAND3 (N6590, N6588, N5425, N2028);
and AND2 (N6591, N6586, N2809);
buf BUF1 (N6592, N6590);
or OR3 (N6593, N6575, N5532, N5036);
nand NAND3 (N6594, N6593, N5692, N6129);
not NOT1 (N6595, N6594);
xor XOR2 (N6596, N6595, N2077);
or OR2 (N6597, N6591, N1892);
nor NOR2 (N6598, N6597, N977);
buf BUF1 (N6599, N6584);
or OR2 (N6600, N6570, N4858);
nor NOR2 (N6601, N6596, N4744);
or OR4 (N6602, N6592, N706, N1430, N988);
nand NAND3 (N6603, N6602, N3297, N1603);
buf BUF1 (N6604, N6603);
nand NAND3 (N6605, N6599, N5656, N1207);
buf BUF1 (N6606, N6604);
not NOT1 (N6607, N6572);
buf BUF1 (N6608, N6606);
buf BUF1 (N6609, N6580);
or OR2 (N6610, N6605, N3192);
or OR4 (N6611, N6607, N5234, N2028, N2611);
not NOT1 (N6612, N6589);
buf BUF1 (N6613, N6611);
not NOT1 (N6614, N6600);
buf BUF1 (N6615, N6608);
and AND3 (N6616, N6613, N5091, N4692);
and AND4 (N6617, N6564, N4738, N872, N2541);
buf BUF1 (N6618, N6610);
xor XOR2 (N6619, N6617, N5859);
not NOT1 (N6620, N6619);
or OR2 (N6621, N6620, N111);
nand NAND3 (N6622, N6609, N1831, N2570);
nor NOR3 (N6623, N6622, N1595, N984);
xor XOR2 (N6624, N6598, N6358);
or OR2 (N6625, N6624, N5604);
xor XOR2 (N6626, N6616, N1294);
nand NAND2 (N6627, N6612, N402);
and AND3 (N6628, N6621, N2266, N3510);
and AND4 (N6629, N6601, N3870, N1232, N1785);
and AND2 (N6630, N6629, N2949);
buf BUF1 (N6631, N6626);
not NOT1 (N6632, N6587);
or OR2 (N6633, N6632, N6420);
nand NAND3 (N6634, N6614, N5948, N4159);
xor XOR2 (N6635, N6630, N3319);
buf BUF1 (N6636, N6628);
not NOT1 (N6637, N6623);
nor NOR2 (N6638, N6633, N4373);
and AND4 (N6639, N6635, N4789, N4771, N3335);
and AND2 (N6640, N6615, N1306);
not NOT1 (N6641, N6639);
nand NAND2 (N6642, N6641, N717);
xor XOR2 (N6643, N6637, N4334);
and AND4 (N6644, N6636, N3258, N5116, N3190);
nor NOR2 (N6645, N6644, N1024);
buf BUF1 (N6646, N6638);
xor XOR2 (N6647, N6643, N4771);
buf BUF1 (N6648, N6618);
xor XOR2 (N6649, N6647, N4481);
or OR4 (N6650, N6648, N181, N3061, N452);
xor XOR2 (N6651, N6642, N817);
nor NOR4 (N6652, N6634, N2950, N2542, N306);
and AND2 (N6653, N6652, N2728);
nor NOR3 (N6654, N6646, N1098, N1242);
buf BUF1 (N6655, N6631);
xor XOR2 (N6656, N6627, N4354);
buf BUF1 (N6657, N6654);
nor NOR3 (N6658, N6657, N747, N1641);
nand NAND2 (N6659, N6649, N5238);
nor NOR2 (N6660, N6645, N5128);
buf BUF1 (N6661, N6650);
not NOT1 (N6662, N6655);
nand NAND2 (N6663, N6658, N965);
xor XOR2 (N6664, N6653, N3551);
and AND2 (N6665, N6625, N4519);
and AND3 (N6666, N6661, N3779, N2832);
xor XOR2 (N6667, N6663, N1051);
xor XOR2 (N6668, N6660, N297);
and AND2 (N6669, N6640, N3260);
xor XOR2 (N6670, N6665, N1061);
buf BUF1 (N6671, N6670);
buf BUF1 (N6672, N6668);
not NOT1 (N6673, N6651);
buf BUF1 (N6674, N6662);
buf BUF1 (N6675, N6664);
nor NOR4 (N6676, N6671, N672, N5406, N6490);
nand NAND2 (N6677, N6666, N3748);
nand NAND4 (N6678, N6674, N4283, N3174, N3808);
or OR3 (N6679, N6667, N21, N3257);
or OR4 (N6680, N6659, N3147, N3934, N3726);
buf BUF1 (N6681, N6677);
and AND3 (N6682, N6678, N5714, N1232);
and AND4 (N6683, N6682, N6632, N5213, N3964);
and AND2 (N6684, N6681, N2461);
or OR3 (N6685, N6656, N862, N6519);
and AND4 (N6686, N6684, N521, N4288, N6114);
nand NAND3 (N6687, N6679, N646, N5706);
nor NOR2 (N6688, N6687, N3985);
nor NOR2 (N6689, N6685, N2785);
and AND3 (N6690, N6686, N1254, N6447);
buf BUF1 (N6691, N6683);
xor XOR2 (N6692, N6690, N2793);
xor XOR2 (N6693, N6691, N6383);
xor XOR2 (N6694, N6675, N5050);
nand NAND2 (N6695, N6672, N5225);
or OR4 (N6696, N6688, N1234, N842, N47);
nand NAND3 (N6697, N6673, N3918, N6368);
nand NAND3 (N6698, N6697, N1490, N5537);
xor XOR2 (N6699, N6696, N4241);
nand NAND2 (N6700, N6699, N3284);
and AND2 (N6701, N6700, N2863);
not NOT1 (N6702, N6694);
nor NOR2 (N6703, N6695, N2379);
buf BUF1 (N6704, N6693);
or OR2 (N6705, N6702, N4122);
nor NOR4 (N6706, N6680, N4820, N488, N280);
nand NAND4 (N6707, N6698, N6119, N3652, N3787);
not NOT1 (N6708, N6701);
nor NOR2 (N6709, N6689, N5281);
or OR3 (N6710, N6669, N3722, N3853);
not NOT1 (N6711, N6704);
and AND3 (N6712, N6706, N1674, N4810);
xor XOR2 (N6713, N6703, N4271);
xor XOR2 (N6714, N6711, N3064);
buf BUF1 (N6715, N6707);
not NOT1 (N6716, N6676);
not NOT1 (N6717, N6710);
not NOT1 (N6718, N6717);
and AND2 (N6719, N6692, N4430);
buf BUF1 (N6720, N6719);
not NOT1 (N6721, N6708);
or OR4 (N6722, N6720, N4072, N251, N3422);
not NOT1 (N6723, N6722);
or OR2 (N6724, N6718, N2260);
xor XOR2 (N6725, N6716, N4068);
and AND4 (N6726, N6709, N3068, N377, N2471);
not NOT1 (N6727, N6705);
not NOT1 (N6728, N6714);
or OR2 (N6729, N6723, N4640);
xor XOR2 (N6730, N6727, N5737);
buf BUF1 (N6731, N6721);
or OR3 (N6732, N6730, N4348, N1048);
nand NAND4 (N6733, N6729, N3310, N3571, N731);
xor XOR2 (N6734, N6726, N3755);
not NOT1 (N6735, N6734);
and AND4 (N6736, N6713, N1065, N5380, N5534);
or OR4 (N6737, N6715, N6285, N2602, N2105);
and AND2 (N6738, N6736, N3987);
not NOT1 (N6739, N6728);
not NOT1 (N6740, N6725);
not NOT1 (N6741, N6739);
or OR3 (N6742, N6740, N4820, N4533);
nand NAND3 (N6743, N6738, N2748, N2554);
nor NOR3 (N6744, N6724, N2232, N3742);
and AND3 (N6745, N6737, N5135, N1266);
xor XOR2 (N6746, N6731, N237);
and AND3 (N6747, N6746, N5672, N3055);
nor NOR2 (N6748, N6741, N6337);
and AND2 (N6749, N6742, N2434);
or OR4 (N6750, N6747, N4880, N2208, N16);
and AND3 (N6751, N6712, N3919, N1338);
nor NOR3 (N6752, N6748, N4174, N101);
buf BUF1 (N6753, N6751);
nand NAND4 (N6754, N6732, N164, N591, N3125);
buf BUF1 (N6755, N6745);
not NOT1 (N6756, N6744);
nand NAND4 (N6757, N6749, N2368, N3972, N2577);
nand NAND4 (N6758, N6754, N2385, N4670, N2740);
xor XOR2 (N6759, N6756, N248);
not NOT1 (N6760, N6733);
buf BUF1 (N6761, N6757);
not NOT1 (N6762, N6735);
xor XOR2 (N6763, N6758, N6183);
or OR2 (N6764, N6750, N5020);
xor XOR2 (N6765, N6764, N2672);
xor XOR2 (N6766, N6762, N2896);
xor XOR2 (N6767, N6743, N598);
not NOT1 (N6768, N6752);
and AND3 (N6769, N6753, N5242, N1662);
buf BUF1 (N6770, N6759);
or OR3 (N6771, N6766, N4499, N5343);
nor NOR4 (N6772, N6761, N1879, N4770, N5492);
nor NOR2 (N6773, N6769, N5599);
or OR2 (N6774, N6765, N6010);
nand NAND2 (N6775, N6771, N4723);
buf BUF1 (N6776, N6763);
and AND4 (N6777, N6773, N4550, N2138, N2234);
buf BUF1 (N6778, N6768);
xor XOR2 (N6779, N6767, N4120);
xor XOR2 (N6780, N6775, N140);
nand NAND3 (N6781, N6755, N914, N3066);
not NOT1 (N6782, N6778);
and AND4 (N6783, N6782, N2476, N1215, N3611);
not NOT1 (N6784, N6779);
nor NOR4 (N6785, N6784, N6649, N1010, N5701);
xor XOR2 (N6786, N6772, N1047);
buf BUF1 (N6787, N6774);
nand NAND3 (N6788, N6777, N5238, N837);
nand NAND4 (N6789, N6760, N868, N2813, N3929);
xor XOR2 (N6790, N6776, N4921);
not NOT1 (N6791, N6788);
xor XOR2 (N6792, N6780, N6096);
xor XOR2 (N6793, N6783, N770);
xor XOR2 (N6794, N6790, N2015);
xor XOR2 (N6795, N6787, N6049);
or OR4 (N6796, N6794, N1419, N1892, N3143);
or OR4 (N6797, N6770, N4283, N57, N4170);
nor NOR4 (N6798, N6793, N5449, N5274, N5519);
nor NOR4 (N6799, N6797, N1804, N3888, N2614);
and AND2 (N6800, N6791, N2330);
buf BUF1 (N6801, N6796);
not NOT1 (N6802, N6801);
and AND4 (N6803, N6785, N5160, N5496, N1869);
not NOT1 (N6804, N6802);
not NOT1 (N6805, N6804);
nor NOR3 (N6806, N6781, N5529, N1066);
nand NAND4 (N6807, N6789, N5471, N4893, N6767);
not NOT1 (N6808, N6806);
not NOT1 (N6809, N6805);
buf BUF1 (N6810, N6799);
nand NAND2 (N6811, N6807, N1382);
nor NOR2 (N6812, N6786, N5529);
xor XOR2 (N6813, N6795, N760);
xor XOR2 (N6814, N6792, N2084);
nor NOR4 (N6815, N6812, N6103, N1583, N3451);
xor XOR2 (N6816, N6813, N1157);
nor NOR3 (N6817, N6808, N2522, N122);
xor XOR2 (N6818, N6815, N425);
xor XOR2 (N6819, N6798, N502);
and AND3 (N6820, N6818, N5121, N4936);
nor NOR2 (N6821, N6817, N2474);
and AND2 (N6822, N6816, N4588);
or OR4 (N6823, N6809, N559, N1252, N2536);
nand NAND3 (N6824, N6810, N428, N3181);
nor NOR3 (N6825, N6824, N5482, N6613);
xor XOR2 (N6826, N6823, N3862);
nor NOR2 (N6827, N6826, N1885);
buf BUF1 (N6828, N6820);
nor NOR4 (N6829, N6803, N2238, N5688, N4411);
not NOT1 (N6830, N6825);
buf BUF1 (N6831, N6828);
nand NAND2 (N6832, N6827, N6056);
nor NOR4 (N6833, N6831, N6690, N5380, N2478);
not NOT1 (N6834, N6800);
or OR2 (N6835, N6822, N6803);
xor XOR2 (N6836, N6834, N3785);
buf BUF1 (N6837, N6819);
xor XOR2 (N6838, N6837, N5547);
xor XOR2 (N6839, N6836, N3396);
xor XOR2 (N6840, N6838, N3073);
nand NAND3 (N6841, N6830, N2467, N1086);
nand NAND4 (N6842, N6840, N2148, N4531, N4125);
or OR3 (N6843, N6842, N31, N1560);
buf BUF1 (N6844, N6832);
or OR2 (N6845, N6843, N163);
buf BUF1 (N6846, N6839);
buf BUF1 (N6847, N6811);
buf BUF1 (N6848, N6833);
or OR2 (N6849, N6829, N4464);
and AND4 (N6850, N6841, N5033, N3679, N4310);
buf BUF1 (N6851, N6850);
nand NAND2 (N6852, N6849, N5345);
nor NOR4 (N6853, N6847, N4596, N5627, N4066);
not NOT1 (N6854, N6846);
nand NAND4 (N6855, N6853, N2109, N4892, N2409);
xor XOR2 (N6856, N6845, N5198);
and AND3 (N6857, N6821, N6782, N4014);
or OR2 (N6858, N6814, N5174);
nand NAND2 (N6859, N6856, N6627);
xor XOR2 (N6860, N6855, N3656);
and AND4 (N6861, N6859, N823, N1921, N988);
nor NOR2 (N6862, N6860, N3076);
nand NAND4 (N6863, N6854, N558, N3459, N4135);
and AND3 (N6864, N6858, N6560, N6324);
or OR3 (N6865, N6835, N4669, N847);
buf BUF1 (N6866, N6844);
nor NOR2 (N6867, N6864, N3694);
not NOT1 (N6868, N6861);
nor NOR2 (N6869, N6863, N4140);
and AND3 (N6870, N6868, N5224, N4701);
xor XOR2 (N6871, N6851, N4570);
and AND2 (N6872, N6852, N919);
and AND3 (N6873, N6848, N4246, N4357);
or OR4 (N6874, N6872, N6520, N6818, N4975);
xor XOR2 (N6875, N6871, N2306);
not NOT1 (N6876, N6874);
buf BUF1 (N6877, N6870);
nor NOR2 (N6878, N6867, N5242);
and AND4 (N6879, N6866, N2754, N3010, N4623);
xor XOR2 (N6880, N6869, N2511);
and AND2 (N6881, N6879, N5487);
nor NOR3 (N6882, N6873, N2982, N3748);
xor XOR2 (N6883, N6878, N2603);
and AND2 (N6884, N6883, N660);
xor XOR2 (N6885, N6865, N2045);
nor NOR3 (N6886, N6862, N3269, N6773);
xor XOR2 (N6887, N6876, N1610);
xor XOR2 (N6888, N6885, N943);
or OR3 (N6889, N6857, N3728, N6292);
and AND3 (N6890, N6889, N1014, N6309);
nand NAND3 (N6891, N6890, N2807, N4097);
and AND2 (N6892, N6875, N3868);
or OR4 (N6893, N6886, N5036, N3490, N2896);
not NOT1 (N6894, N6891);
not NOT1 (N6895, N6881);
nor NOR3 (N6896, N6894, N6054, N1079);
not NOT1 (N6897, N6888);
xor XOR2 (N6898, N6895, N312);
nand NAND3 (N6899, N6892, N4941, N1069);
nand NAND3 (N6900, N6896, N5263, N3652);
and AND2 (N6901, N6880, N4633);
nor NOR2 (N6902, N6884, N889);
or OR3 (N6903, N6887, N3025, N4938);
and AND3 (N6904, N6877, N805, N6523);
or OR2 (N6905, N6893, N3044);
and AND3 (N6906, N6902, N4706, N3153);
not NOT1 (N6907, N6901);
buf BUF1 (N6908, N6900);
and AND4 (N6909, N6882, N6275, N1581, N3731);
not NOT1 (N6910, N6897);
nand NAND3 (N6911, N6903, N27, N1709);
not NOT1 (N6912, N6907);
xor XOR2 (N6913, N6906, N718);
and AND3 (N6914, N6908, N445, N5136);
nor NOR2 (N6915, N6898, N4398);
not NOT1 (N6916, N6910);
nand NAND3 (N6917, N6909, N3597, N208);
buf BUF1 (N6918, N6899);
nor NOR2 (N6919, N6913, N4694);
and AND3 (N6920, N6917, N1602, N2610);
xor XOR2 (N6921, N6912, N6589);
or OR2 (N6922, N6919, N970);
nor NOR2 (N6923, N6914, N195);
or OR4 (N6924, N6923, N3223, N2279, N6618);
buf BUF1 (N6925, N6921);
not NOT1 (N6926, N6920);
buf BUF1 (N6927, N6904);
buf BUF1 (N6928, N6926);
or OR3 (N6929, N6918, N818, N5785);
nand NAND3 (N6930, N6905, N519, N2875);
or OR2 (N6931, N6927, N3573);
buf BUF1 (N6932, N6928);
nor NOR2 (N6933, N6911, N1896);
or OR2 (N6934, N6931, N186);
and AND2 (N6935, N6924, N5045);
buf BUF1 (N6936, N6932);
or OR4 (N6937, N6929, N5438, N5820, N2062);
nand NAND2 (N6938, N6930, N2713);
not NOT1 (N6939, N6938);
xor XOR2 (N6940, N6937, N1469);
nand NAND2 (N6941, N6933, N4247);
and AND2 (N6942, N6925, N3486);
not NOT1 (N6943, N6922);
xor XOR2 (N6944, N6942, N1839);
and AND3 (N6945, N6916, N6636, N3692);
and AND2 (N6946, N6943, N4651);
nor NOR2 (N6947, N6940, N6613);
and AND2 (N6948, N6915, N3281);
xor XOR2 (N6949, N6944, N1932);
nor NOR2 (N6950, N6939, N273);
or OR4 (N6951, N6945, N4165, N879, N4998);
not NOT1 (N6952, N6936);
buf BUF1 (N6953, N6949);
xor XOR2 (N6954, N6941, N1763);
or OR2 (N6955, N6950, N5258);
xor XOR2 (N6956, N6948, N265);
nor NOR3 (N6957, N6946, N4003, N2481);
xor XOR2 (N6958, N6951, N1832);
xor XOR2 (N6959, N6952, N4325);
not NOT1 (N6960, N6953);
not NOT1 (N6961, N6935);
buf BUF1 (N6962, N6960);
not NOT1 (N6963, N6954);
not NOT1 (N6964, N6956);
xor XOR2 (N6965, N6934, N3846);
not NOT1 (N6966, N6947);
nor NOR3 (N6967, N6958, N4835, N511);
buf BUF1 (N6968, N6962);
or OR3 (N6969, N6961, N1346, N4783);
xor XOR2 (N6970, N6957, N3518);
nor NOR4 (N6971, N6964, N5306, N1134, N4020);
nor NOR4 (N6972, N6967, N610, N4178, N3759);
or OR4 (N6973, N6955, N1672, N2040, N1311);
or OR2 (N6974, N6965, N4948);
xor XOR2 (N6975, N6970, N273);
nand NAND4 (N6976, N6973, N771, N1669, N3139);
buf BUF1 (N6977, N6969);
and AND4 (N6978, N6959, N1839, N3203, N5331);
nor NOR4 (N6979, N6976, N4898, N1073, N6941);
nor NOR2 (N6980, N6975, N3456);
or OR3 (N6981, N6980, N5885, N2000);
or OR2 (N6982, N6974, N2559);
xor XOR2 (N6983, N6977, N5785);
nand NAND2 (N6984, N6968, N6684);
nor NOR3 (N6985, N6966, N6288, N4296);
xor XOR2 (N6986, N6985, N466);
xor XOR2 (N6987, N6981, N2680);
xor XOR2 (N6988, N6971, N3052);
or OR2 (N6989, N6982, N2750);
or OR3 (N6990, N6988, N6738, N2468);
and AND2 (N6991, N6986, N6835);
nor NOR4 (N6992, N6972, N1888, N3828, N35);
buf BUF1 (N6993, N6990);
buf BUF1 (N6994, N6978);
or OR4 (N6995, N6984, N1887, N1, N3163);
xor XOR2 (N6996, N6989, N3209);
xor XOR2 (N6997, N6979, N6777);
nor NOR4 (N6998, N6997, N1929, N6915, N5762);
or OR4 (N6999, N6998, N1326, N700, N3367);
not NOT1 (N7000, N6963);
or OR2 (N7001, N7000, N245);
xor XOR2 (N7002, N6992, N1762);
or OR2 (N7003, N6987, N6471);
nor NOR4 (N7004, N7003, N6413, N428, N1587);
and AND2 (N7005, N7001, N3434);
nor NOR3 (N7006, N6991, N4434, N2302);
nand NAND2 (N7007, N6996, N774);
xor XOR2 (N7008, N7002, N3198);
or OR4 (N7009, N7006, N1259, N5778, N5616);
not NOT1 (N7010, N7005);
buf BUF1 (N7011, N7004);
and AND4 (N7012, N7011, N2105, N1609, N4140);
nor NOR4 (N7013, N7012, N2059, N5780, N6496);
or OR4 (N7014, N6994, N4836, N2311, N1473);
buf BUF1 (N7015, N7007);
nand NAND3 (N7016, N6983, N1524, N5275);
not NOT1 (N7017, N7008);
nand NAND2 (N7018, N7009, N1932);
nand NAND2 (N7019, N7015, N4339);
xor XOR2 (N7020, N6999, N5605);
not NOT1 (N7021, N7017);
nand NAND4 (N7022, N6993, N1079, N3798, N2872);
and AND3 (N7023, N7018, N3127, N3131);
or OR3 (N7024, N7019, N6181, N6395);
not NOT1 (N7025, N7022);
nor NOR4 (N7026, N6995, N2754, N1032, N244);
xor XOR2 (N7027, N7026, N4473);
and AND4 (N7028, N7021, N1813, N1381, N4899);
and AND2 (N7029, N7014, N985);
xor XOR2 (N7030, N7027, N5342);
xor XOR2 (N7031, N7024, N4144);
nor NOR3 (N7032, N7031, N3548, N2978);
nand NAND4 (N7033, N7025, N6896, N2216, N3585);
buf BUF1 (N7034, N7029);
and AND3 (N7035, N7033, N4550, N4357);
buf BUF1 (N7036, N7020);
nand NAND3 (N7037, N7035, N5205, N2447);
and AND3 (N7038, N7023, N1595, N1224);
nand NAND2 (N7039, N7034, N6562);
nor NOR4 (N7040, N7028, N3392, N217, N6285);
nor NOR4 (N7041, N7037, N4440, N5820, N303);
buf BUF1 (N7042, N7016);
not NOT1 (N7043, N7042);
not NOT1 (N7044, N7038);
xor XOR2 (N7045, N7039, N4602);
or OR3 (N7046, N7044, N6745, N5958);
xor XOR2 (N7047, N7046, N2823);
not NOT1 (N7048, N7041);
xor XOR2 (N7049, N7043, N2169);
or OR3 (N7050, N7013, N3340, N4982);
or OR2 (N7051, N7045, N6473);
nor NOR4 (N7052, N7030, N1028, N343, N6816);
nor NOR2 (N7053, N7048, N886);
nand NAND3 (N7054, N7010, N686, N1818);
and AND2 (N7055, N7053, N4816);
or OR4 (N7056, N7055, N2130, N1524, N3322);
and AND4 (N7057, N7051, N4392, N5541, N4507);
buf BUF1 (N7058, N7047);
or OR4 (N7059, N7036, N6608, N5711, N5447);
or OR4 (N7060, N7057, N2487, N5177, N4390);
buf BUF1 (N7061, N7052);
and AND3 (N7062, N7060, N4619, N4755);
and AND2 (N7063, N7032, N4733);
buf BUF1 (N7064, N7063);
not NOT1 (N7065, N7050);
not NOT1 (N7066, N7049);
not NOT1 (N7067, N7040);
nor NOR3 (N7068, N7064, N379, N1176);
not NOT1 (N7069, N7066);
nand NAND3 (N7070, N7056, N2271, N2001);
buf BUF1 (N7071, N7054);
and AND4 (N7072, N7070, N3349, N4529, N873);
buf BUF1 (N7073, N7068);
not NOT1 (N7074, N7073);
nor NOR2 (N7075, N7062, N4288);
xor XOR2 (N7076, N7075, N6324);
and AND3 (N7077, N7076, N3752, N1508);
xor XOR2 (N7078, N7061, N1996);
and AND4 (N7079, N7074, N1957, N4783, N2830);
xor XOR2 (N7080, N7077, N435);
nand NAND4 (N7081, N7067, N3789, N3687, N6492);
not NOT1 (N7082, N7081);
nand NAND4 (N7083, N7059, N6865, N5177, N5006);
buf BUF1 (N7084, N7080);
buf BUF1 (N7085, N7078);
or OR3 (N7086, N7084, N3158, N1071);
not NOT1 (N7087, N7071);
nand NAND4 (N7088, N7058, N318, N4821, N2494);
nand NAND4 (N7089, N7072, N6733, N2768, N3800);
xor XOR2 (N7090, N7088, N4208);
xor XOR2 (N7091, N7090, N4469);
or OR4 (N7092, N7086, N6281, N2226, N1595);
xor XOR2 (N7093, N7079, N1490);
buf BUF1 (N7094, N7087);
nand NAND2 (N7095, N7085, N508);
xor XOR2 (N7096, N7095, N520);
xor XOR2 (N7097, N7094, N2498);
nand NAND2 (N7098, N7069, N4129);
xor XOR2 (N7099, N7083, N3807);
and AND2 (N7100, N7092, N5930);
or OR4 (N7101, N7091, N1705, N2977, N5029);
xor XOR2 (N7102, N7089, N4067);
buf BUF1 (N7103, N7097);
buf BUF1 (N7104, N7101);
nand NAND2 (N7105, N7100, N2432);
nand NAND4 (N7106, N7093, N7085, N5743, N5375);
and AND3 (N7107, N7106, N6530, N2448);
or OR3 (N7108, N7107, N973, N1770);
not NOT1 (N7109, N7102);
nand NAND3 (N7110, N7096, N5275, N4223);
buf BUF1 (N7111, N7082);
nand NAND4 (N7112, N7109, N3097, N6879, N884);
nand NAND2 (N7113, N7111, N4934);
and AND4 (N7114, N7112, N2324, N6284, N5535);
buf BUF1 (N7115, N7105);
not NOT1 (N7116, N7115);
nor NOR2 (N7117, N7108, N2393);
or OR2 (N7118, N7116, N4493);
xor XOR2 (N7119, N7110, N6010);
nand NAND2 (N7120, N7098, N5315);
not NOT1 (N7121, N7117);
and AND2 (N7122, N7121, N5898);
and AND2 (N7123, N7114, N684);
xor XOR2 (N7124, N7104, N4320);
xor XOR2 (N7125, N7118, N3119);
nor NOR2 (N7126, N7065, N5125);
xor XOR2 (N7127, N7125, N2543);
and AND4 (N7128, N7103, N3443, N1348, N3532);
nor NOR2 (N7129, N7127, N6228);
not NOT1 (N7130, N7123);
buf BUF1 (N7131, N7119);
and AND2 (N7132, N7128, N2021);
xor XOR2 (N7133, N7129, N5744);
not NOT1 (N7134, N7133);
buf BUF1 (N7135, N7122);
or OR2 (N7136, N7099, N1478);
xor XOR2 (N7137, N7124, N3706);
nor NOR2 (N7138, N7126, N815);
nor NOR4 (N7139, N7136, N5495, N1060, N3177);
xor XOR2 (N7140, N7134, N3998);
and AND3 (N7141, N7132, N2797, N52);
or OR2 (N7142, N7137, N202);
and AND4 (N7143, N7138, N4477, N4267, N5082);
or OR4 (N7144, N7142, N5664, N4469, N3123);
or OR3 (N7145, N7141, N3307, N86);
and AND2 (N7146, N7135, N6180);
and AND3 (N7147, N7139, N6657, N37);
nand NAND3 (N7148, N7120, N3793, N231);
not NOT1 (N7149, N7145);
and AND2 (N7150, N7143, N4480);
or OR2 (N7151, N7140, N526);
or OR2 (N7152, N7144, N1104);
or OR2 (N7153, N7152, N963);
nor NOR3 (N7154, N7146, N1340, N6073);
nand NAND4 (N7155, N7150, N2649, N681, N2918);
and AND2 (N7156, N7149, N6708);
or OR2 (N7157, N7153, N397);
not NOT1 (N7158, N7148);
and AND4 (N7159, N7130, N3994, N4162, N6481);
or OR2 (N7160, N7151, N2845);
and AND3 (N7161, N7155, N7155, N931);
buf BUF1 (N7162, N7154);
or OR3 (N7163, N7161, N5569, N1628);
nand NAND4 (N7164, N7131, N2747, N3779, N4846);
and AND3 (N7165, N7162, N793, N160);
and AND2 (N7166, N7158, N568);
nor NOR3 (N7167, N7160, N893, N4846);
xor XOR2 (N7168, N7166, N5482);
nor NOR3 (N7169, N7163, N5116, N709);
or OR4 (N7170, N7156, N4450, N5617, N2910);
buf BUF1 (N7171, N7164);
nand NAND2 (N7172, N7113, N1061);
not NOT1 (N7173, N7167);
buf BUF1 (N7174, N7165);
buf BUF1 (N7175, N7157);
nor NOR3 (N7176, N7174, N3945, N3531);
or OR3 (N7177, N7173, N3951, N6612);
and AND2 (N7178, N7147, N6971);
xor XOR2 (N7179, N7176, N6074);
not NOT1 (N7180, N7159);
buf BUF1 (N7181, N7171);
and AND3 (N7182, N7168, N3130, N3548);
nor NOR4 (N7183, N7172, N937, N1980, N5815);
xor XOR2 (N7184, N7170, N6134);
nor NOR2 (N7185, N7169, N194);
nor NOR4 (N7186, N7178, N2691, N3009, N4470);
nor NOR4 (N7187, N7184, N1006, N4927, N3420);
nand NAND4 (N7188, N7177, N2713, N1074, N6520);
nor NOR3 (N7189, N7183, N3726, N3263);
nand NAND4 (N7190, N7185, N6532, N4542, N3720);
nand NAND2 (N7191, N7179, N7122);
not NOT1 (N7192, N7175);
buf BUF1 (N7193, N7188);
xor XOR2 (N7194, N7181, N6460);
buf BUF1 (N7195, N7194);
not NOT1 (N7196, N7195);
nor NOR3 (N7197, N7192, N1071, N3192);
nand NAND3 (N7198, N7197, N4763, N6953);
xor XOR2 (N7199, N7193, N2513);
not NOT1 (N7200, N7182);
or OR4 (N7201, N7189, N6687, N2443, N510);
and AND4 (N7202, N7190, N300, N698, N685);
buf BUF1 (N7203, N7202);
buf BUF1 (N7204, N7203);
buf BUF1 (N7205, N7191);
nand NAND4 (N7206, N7199, N4389, N2606, N4501);
nor NOR3 (N7207, N7186, N279, N5216);
and AND2 (N7208, N7187, N2820);
or OR3 (N7209, N7201, N2392, N3391);
buf BUF1 (N7210, N7198);
nand NAND4 (N7211, N7209, N358, N1315, N4684);
nand NAND2 (N7212, N7210, N6461);
nand NAND4 (N7213, N7207, N942, N6970, N4669);
nand NAND2 (N7214, N7204, N3639);
nor NOR2 (N7215, N7212, N3329);
nand NAND4 (N7216, N7214, N2596, N6872, N3713);
nand NAND4 (N7217, N7215, N5842, N2726, N1443);
xor XOR2 (N7218, N7206, N1463);
nand NAND2 (N7219, N7180, N1766);
nor NOR2 (N7220, N7211, N5091);
buf BUF1 (N7221, N7218);
nand NAND2 (N7222, N7200, N5721);
xor XOR2 (N7223, N7208, N2111);
nand NAND3 (N7224, N7213, N5744, N6406);
or OR2 (N7225, N7221, N5196);
nand NAND3 (N7226, N7220, N6406, N2962);
or OR3 (N7227, N7219, N1316, N6786);
buf BUF1 (N7228, N7217);
and AND2 (N7229, N7227, N6226);
nand NAND3 (N7230, N7196, N22, N2826);
nand NAND2 (N7231, N7230, N1706);
and AND4 (N7232, N7229, N1228, N1233, N4403);
buf BUF1 (N7233, N7216);
xor XOR2 (N7234, N7225, N6554);
or OR2 (N7235, N7228, N3651);
and AND3 (N7236, N7234, N693, N2966);
and AND3 (N7237, N7222, N1781, N2098);
and AND4 (N7238, N7205, N169, N5352, N5997);
nand NAND2 (N7239, N7231, N1256);
not NOT1 (N7240, N7238);
or OR4 (N7241, N7236, N4937, N3752, N502);
buf BUF1 (N7242, N7237);
nand NAND3 (N7243, N7241, N1770, N1516);
xor XOR2 (N7244, N7223, N2433);
and AND2 (N7245, N7239, N5002);
not NOT1 (N7246, N7240);
and AND3 (N7247, N7224, N1743, N2361);
nor NOR4 (N7248, N7246, N437, N2263, N667);
and AND3 (N7249, N7243, N4502, N2038);
not NOT1 (N7250, N7247);
or OR3 (N7251, N7242, N785, N2974);
and AND3 (N7252, N7232, N3311, N6555);
not NOT1 (N7253, N7252);
or OR4 (N7254, N7248, N3834, N1935, N2265);
not NOT1 (N7255, N7233);
or OR4 (N7256, N7251, N6226, N6329, N804);
buf BUF1 (N7257, N7253);
buf BUF1 (N7258, N7245);
nor NOR4 (N7259, N7244, N6537, N5283, N4294);
buf BUF1 (N7260, N7257);
buf BUF1 (N7261, N7258);
and AND4 (N7262, N7259, N4229, N482, N4534);
not NOT1 (N7263, N7250);
not NOT1 (N7264, N7263);
nor NOR3 (N7265, N7261, N5300, N2779);
and AND4 (N7266, N7264, N5595, N5845, N6972);
or OR4 (N7267, N7266, N5108, N1507, N442);
buf BUF1 (N7268, N7235);
buf BUF1 (N7269, N7260);
buf BUF1 (N7270, N7226);
or OR3 (N7271, N7268, N4374, N1843);
xor XOR2 (N7272, N7270, N30);
not NOT1 (N7273, N7262);
nand NAND3 (N7274, N7255, N4611, N295);
xor XOR2 (N7275, N7271, N6677);
and AND2 (N7276, N7249, N1114);
buf BUF1 (N7277, N7274);
xor XOR2 (N7278, N7256, N2184);
or OR2 (N7279, N7269, N6843);
buf BUF1 (N7280, N7265);
and AND3 (N7281, N7254, N6717, N4074);
and AND3 (N7282, N7272, N5617, N854);
or OR3 (N7283, N7280, N6197, N892);
nand NAND4 (N7284, N7275, N7165, N5708, N5359);
or OR3 (N7285, N7273, N4974, N3920);
nand NAND2 (N7286, N7276, N5639);
buf BUF1 (N7287, N7282);
nor NOR4 (N7288, N7278, N2, N1654, N929);
and AND3 (N7289, N7284, N1917, N1550);
buf BUF1 (N7290, N7289);
xor XOR2 (N7291, N7279, N2969);
nand NAND4 (N7292, N7277, N7239, N5516, N2961);
nand NAND2 (N7293, N7288, N635);
buf BUF1 (N7294, N7292);
not NOT1 (N7295, N7285);
buf BUF1 (N7296, N7291);
not NOT1 (N7297, N7293);
nand NAND4 (N7298, N7297, N1623, N4500, N895);
and AND4 (N7299, N7286, N3302, N5455, N1752);
buf BUF1 (N7300, N7283);
nand NAND2 (N7301, N7299, N2682);
nor NOR4 (N7302, N7298, N5940, N6567, N5018);
and AND3 (N7303, N7295, N5579, N2240);
nand NAND4 (N7304, N7290, N2442, N6660, N7208);
nor NOR2 (N7305, N7296, N4083);
or OR3 (N7306, N7302, N7038, N2111);
nand NAND3 (N7307, N7267, N4278, N2171);
nor NOR2 (N7308, N7281, N6554);
and AND4 (N7309, N7300, N5077, N4033, N2416);
or OR3 (N7310, N7303, N5421, N7298);
nand NAND3 (N7311, N7304, N5723, N2108);
nand NAND2 (N7312, N7308, N5189);
nor NOR3 (N7313, N7307, N784, N2828);
xor XOR2 (N7314, N7313, N4179);
nor NOR2 (N7315, N7310, N3205);
xor XOR2 (N7316, N7315, N5319);
nand NAND3 (N7317, N7316, N2463, N5576);
or OR2 (N7318, N7305, N4435);
nor NOR4 (N7319, N7301, N2705, N5058, N1889);
nor NOR2 (N7320, N7311, N4476);
or OR3 (N7321, N7319, N1488, N6740);
and AND4 (N7322, N7321, N921, N4116, N5928);
or OR2 (N7323, N7287, N4927);
not NOT1 (N7324, N7312);
or OR2 (N7325, N7317, N5610);
and AND2 (N7326, N7294, N47);
or OR2 (N7327, N7325, N5149);
or OR2 (N7328, N7320, N5653);
xor XOR2 (N7329, N7309, N797);
not NOT1 (N7330, N7328);
not NOT1 (N7331, N7327);
and AND3 (N7332, N7324, N4619, N142);
or OR2 (N7333, N7330, N4994);
not NOT1 (N7334, N7322);
nor NOR4 (N7335, N7323, N371, N265, N3457);
nand NAND2 (N7336, N7329, N700);
nand NAND2 (N7337, N7306, N4360);
nor NOR4 (N7338, N7326, N6889, N4203, N2627);
and AND2 (N7339, N7335, N280);
not NOT1 (N7340, N7332);
nand NAND4 (N7341, N7334, N4767, N4822, N2367);
or OR4 (N7342, N7339, N2115, N2425, N1025);
nand NAND3 (N7343, N7336, N1680, N4140);
xor XOR2 (N7344, N7340, N5297);
xor XOR2 (N7345, N7341, N937);
buf BUF1 (N7346, N7338);
and AND3 (N7347, N7318, N6710, N2878);
and AND3 (N7348, N7333, N2857, N1879);
xor XOR2 (N7349, N7344, N6520);
nor NOR4 (N7350, N7349, N447, N3970, N2185);
nor NOR4 (N7351, N7348, N1058, N5490, N3405);
nor NOR2 (N7352, N7314, N2072);
nand NAND4 (N7353, N7346, N2754, N7276, N6301);
buf BUF1 (N7354, N7342);
or OR2 (N7355, N7343, N3314);
not NOT1 (N7356, N7347);
xor XOR2 (N7357, N7356, N2118);
nand NAND4 (N7358, N7337, N1492, N887, N6366);
or OR3 (N7359, N7355, N7358, N2395);
not NOT1 (N7360, N3606);
and AND3 (N7361, N7345, N6947, N1577);
nor NOR3 (N7362, N7361, N410, N6766);
or OR3 (N7363, N7354, N3373, N3111);
and AND4 (N7364, N7360, N1823, N6931, N767);
buf BUF1 (N7365, N7364);
nor NOR4 (N7366, N7363, N3591, N1697, N7288);
and AND2 (N7367, N7359, N6869);
buf BUF1 (N7368, N7365);
xor XOR2 (N7369, N7331, N2251);
buf BUF1 (N7370, N7367);
and AND3 (N7371, N7362, N7291, N6854);
buf BUF1 (N7372, N7351);
not NOT1 (N7373, N7350);
buf BUF1 (N7374, N7372);
buf BUF1 (N7375, N7357);
and AND3 (N7376, N7371, N6515, N1118);
nor NOR4 (N7377, N7375, N2604, N6589, N5138);
and AND2 (N7378, N7373, N55);
xor XOR2 (N7379, N7352, N1207);
or OR3 (N7380, N7374, N3452, N4429);
nand NAND3 (N7381, N7370, N772, N6943);
buf BUF1 (N7382, N7378);
and AND3 (N7383, N7381, N5185, N6265);
xor XOR2 (N7384, N7368, N6414);
nor NOR2 (N7385, N7380, N704);
not NOT1 (N7386, N7384);
nor NOR3 (N7387, N7353, N2608, N4908);
xor XOR2 (N7388, N7379, N3837);
buf BUF1 (N7389, N7388);
not NOT1 (N7390, N7385);
xor XOR2 (N7391, N7376, N1603);
or OR2 (N7392, N7387, N3789);
and AND2 (N7393, N7390, N5533);
xor XOR2 (N7394, N7369, N1829);
or OR3 (N7395, N7394, N2126, N3268);
buf BUF1 (N7396, N7393);
buf BUF1 (N7397, N7391);
or OR3 (N7398, N7383, N6769, N706);
not NOT1 (N7399, N7392);
nor NOR3 (N7400, N7386, N501, N3588);
and AND3 (N7401, N7382, N4704, N2220);
or OR4 (N7402, N7400, N2767, N3990, N3794);
buf BUF1 (N7403, N7395);
and AND4 (N7404, N7398, N63, N4828, N2597);
nor NOR3 (N7405, N7404, N2049, N6502);
and AND4 (N7406, N7405, N6620, N6852, N6545);
nand NAND2 (N7407, N7399, N3167);
nand NAND2 (N7408, N7366, N4734);
xor XOR2 (N7409, N7408, N3267);
buf BUF1 (N7410, N7406);
and AND4 (N7411, N7410, N5588, N510, N3821);
not NOT1 (N7412, N7397);
nand NAND2 (N7413, N7412, N4113);
nand NAND2 (N7414, N7403, N334);
and AND3 (N7415, N7402, N5759, N2238);
not NOT1 (N7416, N7413);
and AND3 (N7417, N7389, N516, N288);
not NOT1 (N7418, N7377);
buf BUF1 (N7419, N7401);
not NOT1 (N7420, N7418);
not NOT1 (N7421, N7407);
xor XOR2 (N7422, N7420, N1506);
nor NOR4 (N7423, N7396, N7238, N585, N2909);
or OR4 (N7424, N7419, N2205, N5082, N3551);
or OR4 (N7425, N7424, N431, N6663, N4399);
and AND3 (N7426, N7414, N6034, N6261);
not NOT1 (N7427, N7409);
and AND4 (N7428, N7427, N1833, N4926, N5512);
and AND3 (N7429, N7423, N4389, N1722);
nand NAND2 (N7430, N7417, N3968);
not NOT1 (N7431, N7422);
or OR3 (N7432, N7426, N7391, N1353);
xor XOR2 (N7433, N7425, N3533);
nor NOR4 (N7434, N7429, N2774, N4001, N2352);
buf BUF1 (N7435, N7431);
nand NAND4 (N7436, N7430, N37, N5439, N3438);
not NOT1 (N7437, N7434);
xor XOR2 (N7438, N7436, N3058);
nor NOR3 (N7439, N7428, N4991, N686);
xor XOR2 (N7440, N7421, N3129);
nand NAND4 (N7441, N7440, N4449, N7093, N4123);
or OR4 (N7442, N7411, N3831, N4539, N3717);
buf BUF1 (N7443, N7442);
not NOT1 (N7444, N7438);
nor NOR4 (N7445, N7415, N5655, N4931, N3274);
or OR3 (N7446, N7444, N5533, N2669);
or OR2 (N7447, N7432, N6519);
and AND3 (N7448, N7416, N6354, N2840);
nor NOR4 (N7449, N7446, N3750, N706, N1024);
nor NOR2 (N7450, N7443, N7446);
or OR3 (N7451, N7450, N4618, N763);
and AND2 (N7452, N7433, N5745);
xor XOR2 (N7453, N7451, N3672);
or OR3 (N7454, N7453, N5591, N2848);
not NOT1 (N7455, N7454);
and AND2 (N7456, N7452, N6565);
or OR3 (N7457, N7435, N5186, N4388);
nand NAND2 (N7458, N7457, N5115);
and AND3 (N7459, N7437, N6277, N148);
and AND2 (N7460, N7449, N7129);
xor XOR2 (N7461, N7458, N4514);
or OR3 (N7462, N7459, N1415, N6390);
and AND3 (N7463, N7439, N4410, N5215);
nor NOR4 (N7464, N7463, N4253, N4825, N5153);
and AND4 (N7465, N7445, N554, N6429, N1771);
and AND3 (N7466, N7455, N1426, N6968);
xor XOR2 (N7467, N7466, N7080);
and AND4 (N7468, N7461, N3555, N1196, N2511);
nand NAND4 (N7469, N7448, N5010, N4297, N1263);
xor XOR2 (N7470, N7462, N3790);
nand NAND4 (N7471, N7465, N865, N7376, N6676);
buf BUF1 (N7472, N7471);
and AND4 (N7473, N7460, N1980, N4745, N1457);
nor NOR4 (N7474, N7456, N5717, N866, N3285);
or OR2 (N7475, N7468, N3648);
nor NOR3 (N7476, N7469, N5692, N4223);
nand NAND2 (N7477, N7475, N5774);
and AND4 (N7478, N7473, N5246, N2440, N4476);
nor NOR3 (N7479, N7476, N5378, N5101);
buf BUF1 (N7480, N7472);
nand NAND3 (N7481, N7447, N696, N4722);
not NOT1 (N7482, N7480);
or OR2 (N7483, N7467, N1456);
not NOT1 (N7484, N7470);
xor XOR2 (N7485, N7484, N2717);
buf BUF1 (N7486, N7483);
or OR3 (N7487, N7479, N5087, N2953);
or OR2 (N7488, N7481, N3163);
or OR2 (N7489, N7487, N1460);
and AND4 (N7490, N7478, N6505, N3639, N3529);
xor XOR2 (N7491, N7441, N2434);
xor XOR2 (N7492, N7477, N1637);
not NOT1 (N7493, N7488);
xor XOR2 (N7494, N7485, N466);
xor XOR2 (N7495, N7493, N4986);
nor NOR4 (N7496, N7495, N637, N5367, N2303);
and AND2 (N7497, N7492, N6063);
buf BUF1 (N7498, N7494);
not NOT1 (N7499, N7489);
and AND3 (N7500, N7464, N2298, N930);
nor NOR3 (N7501, N7491, N2663, N2606);
buf BUF1 (N7502, N7499);
xor XOR2 (N7503, N7486, N518);
xor XOR2 (N7504, N7490, N3568);
and AND4 (N7505, N7503, N7333, N7021, N7348);
or OR3 (N7506, N7500, N727, N1909);
and AND2 (N7507, N7482, N1154);
xor XOR2 (N7508, N7497, N7374);
or OR3 (N7509, N7507, N5654, N3696);
nor NOR2 (N7510, N7502, N6465);
xor XOR2 (N7511, N7508, N7500);
xor XOR2 (N7512, N7509, N6934);
xor XOR2 (N7513, N7474, N1054);
and AND2 (N7514, N7505, N1771);
nor NOR4 (N7515, N7510, N4278, N1193, N1433);
xor XOR2 (N7516, N7498, N3779);
and AND3 (N7517, N7506, N241, N3321);
or OR2 (N7518, N7514, N3522);
nor NOR4 (N7519, N7496, N7297, N1350, N572);
and AND2 (N7520, N7518, N7354);
not NOT1 (N7521, N7512);
buf BUF1 (N7522, N7511);
and AND2 (N7523, N7516, N4372);
or OR3 (N7524, N7523, N6117, N2979);
xor XOR2 (N7525, N7501, N3627);
nor NOR3 (N7526, N7519, N3749, N1856);
buf BUF1 (N7527, N7504);
or OR3 (N7528, N7517, N1752, N471);
or OR2 (N7529, N7524, N3525);
not NOT1 (N7530, N7528);
xor XOR2 (N7531, N7520, N5943);
nor NOR4 (N7532, N7515, N6175, N2498, N1683);
not NOT1 (N7533, N7532);
nor NOR3 (N7534, N7533, N5381, N2299);
buf BUF1 (N7535, N7530);
buf BUF1 (N7536, N7535);
and AND3 (N7537, N7536, N6969, N2614);
buf BUF1 (N7538, N7521);
not NOT1 (N7539, N7531);
nor NOR2 (N7540, N7522, N1269);
not NOT1 (N7541, N7527);
nor NOR3 (N7542, N7539, N6642, N2624);
buf BUF1 (N7543, N7537);
buf BUF1 (N7544, N7526);
nor NOR4 (N7545, N7544, N6851, N6736, N5243);
or OR2 (N7546, N7513, N5532);
nor NOR4 (N7547, N7529, N569, N6812, N491);
not NOT1 (N7548, N7540);
and AND4 (N7549, N7545, N2725, N7500, N355);
or OR4 (N7550, N7542, N487, N3980, N7369);
not NOT1 (N7551, N7547);
and AND4 (N7552, N7546, N5054, N4828, N1896);
or OR4 (N7553, N7549, N7176, N5843, N640);
buf BUF1 (N7554, N7525);
not NOT1 (N7555, N7553);
xor XOR2 (N7556, N7548, N2291);
nand NAND2 (N7557, N7550, N4462);
or OR4 (N7558, N7552, N3183, N6025, N3975);
or OR2 (N7559, N7538, N7349);
nor NOR4 (N7560, N7551, N1441, N1860, N2477);
nor NOR2 (N7561, N7554, N4482);
nor NOR3 (N7562, N7541, N7061, N3458);
nor NOR3 (N7563, N7555, N1237, N4202);
nand NAND4 (N7564, N7557, N3440, N346, N4539);
xor XOR2 (N7565, N7563, N424);
or OR3 (N7566, N7543, N2013, N4190);
and AND3 (N7567, N7534, N517, N134);
buf BUF1 (N7568, N7564);
buf BUF1 (N7569, N7565);
xor XOR2 (N7570, N7556, N3963);
buf BUF1 (N7571, N7567);
buf BUF1 (N7572, N7571);
nor NOR2 (N7573, N7569, N413);
nand NAND2 (N7574, N7566, N3834);
buf BUF1 (N7575, N7572);
xor XOR2 (N7576, N7575, N340);
or OR2 (N7577, N7559, N703);
or OR2 (N7578, N7568, N3418);
nor NOR3 (N7579, N7562, N4632, N19);
and AND2 (N7580, N7578, N6800);
not NOT1 (N7581, N7561);
nand NAND3 (N7582, N7570, N2500, N1013);
xor XOR2 (N7583, N7574, N5664);
nor NOR2 (N7584, N7576, N214);
nand NAND2 (N7585, N7580, N1163);
or OR4 (N7586, N7581, N1643, N5220, N5468);
xor XOR2 (N7587, N7583, N7204);
nand NAND4 (N7588, N7573, N778, N7288, N151);
nand NAND2 (N7589, N7560, N6022);
xor XOR2 (N7590, N7582, N6686);
nor NOR4 (N7591, N7587, N934, N2323, N5636);
nand NAND4 (N7592, N7577, N1190, N7246, N6806);
or OR4 (N7593, N7589, N258, N1448, N335);
nand NAND2 (N7594, N7584, N3692);
nor NOR4 (N7595, N7558, N253, N2846, N2682);
nand NAND2 (N7596, N7588, N3462);
nand NAND3 (N7597, N7593, N1950, N642);
and AND2 (N7598, N7585, N413);
not NOT1 (N7599, N7594);
nand NAND3 (N7600, N7586, N691, N6061);
or OR2 (N7601, N7597, N2952);
nand NAND3 (N7602, N7601, N4437, N4001);
xor XOR2 (N7603, N7598, N1025);
nand NAND2 (N7604, N7579, N7209);
xor XOR2 (N7605, N7604, N213);
and AND4 (N7606, N7605, N1839, N5666, N7166);
or OR3 (N7607, N7600, N4858, N2442);
nor NOR2 (N7608, N7595, N93);
not NOT1 (N7609, N7607);
and AND2 (N7610, N7592, N330);
not NOT1 (N7611, N7590);
or OR2 (N7612, N7602, N1080);
and AND3 (N7613, N7603, N1790, N7148);
buf BUF1 (N7614, N7596);
and AND4 (N7615, N7611, N5306, N6882, N1004);
nor NOR4 (N7616, N7599, N5917, N1250, N553);
xor XOR2 (N7617, N7615, N6025);
not NOT1 (N7618, N7610);
and AND4 (N7619, N7606, N417, N2137, N6137);
nor NOR2 (N7620, N7612, N5394);
buf BUF1 (N7621, N7620);
xor XOR2 (N7622, N7591, N5082);
xor XOR2 (N7623, N7622, N5182);
xor XOR2 (N7624, N7613, N6226);
nand NAND2 (N7625, N7624, N4811);
not NOT1 (N7626, N7625);
xor XOR2 (N7627, N7621, N767);
xor XOR2 (N7628, N7616, N1588);
nand NAND2 (N7629, N7614, N3652);
not NOT1 (N7630, N7623);
buf BUF1 (N7631, N7627);
and AND4 (N7632, N7619, N6753, N7166, N2243);
or OR2 (N7633, N7618, N2435);
buf BUF1 (N7634, N7626);
not NOT1 (N7635, N7628);
not NOT1 (N7636, N7633);
and AND4 (N7637, N7630, N4775, N478, N3734);
buf BUF1 (N7638, N7634);
xor XOR2 (N7639, N7636, N3705);
nor NOR4 (N7640, N7609, N1770, N6678, N1105);
nor NOR3 (N7641, N7617, N5962, N4269);
not NOT1 (N7642, N7632);
nand NAND3 (N7643, N7629, N3753, N5573);
xor XOR2 (N7644, N7637, N3207);
or OR4 (N7645, N7608, N5216, N6174, N6453);
nor NOR2 (N7646, N7631, N6129);
xor XOR2 (N7647, N7640, N5201);
xor XOR2 (N7648, N7635, N4637);
nor NOR3 (N7649, N7647, N55, N4263);
buf BUF1 (N7650, N7639);
buf BUF1 (N7651, N7645);
or OR2 (N7652, N7649, N5779);
and AND4 (N7653, N7646, N7561, N4586, N4643);
xor XOR2 (N7654, N7650, N2007);
buf BUF1 (N7655, N7641);
nor NOR3 (N7656, N7644, N3505, N2427);
and AND2 (N7657, N7654, N5754);
nor NOR4 (N7658, N7648, N7430, N366, N485);
not NOT1 (N7659, N7651);
and AND2 (N7660, N7655, N5580);
nor NOR3 (N7661, N7659, N3341, N1739);
xor XOR2 (N7662, N7660, N3302);
and AND4 (N7663, N7653, N3525, N583, N6565);
nand NAND4 (N7664, N7652, N2688, N6781, N3708);
nor NOR2 (N7665, N7656, N2766);
xor XOR2 (N7666, N7664, N2063);
and AND2 (N7667, N7643, N1563);
xor XOR2 (N7668, N7663, N5309);
buf BUF1 (N7669, N7662);
xor XOR2 (N7670, N7669, N1875);
and AND2 (N7671, N7638, N5980);
not NOT1 (N7672, N7668);
nor NOR4 (N7673, N7667, N6656, N1536, N1348);
and AND2 (N7674, N7665, N1892);
nand NAND2 (N7675, N7670, N3713);
or OR3 (N7676, N7674, N3589, N36);
xor XOR2 (N7677, N7666, N2558);
nor NOR3 (N7678, N7658, N1677, N5315);
or OR3 (N7679, N7671, N1770, N2693);
not NOT1 (N7680, N7676);
not NOT1 (N7681, N7675);
and AND3 (N7682, N7680, N5819, N2612);
nor NOR3 (N7683, N7679, N3424, N6876);
buf BUF1 (N7684, N7642);
buf BUF1 (N7685, N7657);
nor NOR3 (N7686, N7682, N3593, N188);
or OR3 (N7687, N7686, N1859, N3834);
xor XOR2 (N7688, N7684, N7270);
and AND3 (N7689, N7683, N2224, N5062);
xor XOR2 (N7690, N7681, N6246);
not NOT1 (N7691, N7688);
or OR4 (N7692, N7677, N4280, N975, N6759);
or OR2 (N7693, N7689, N5456);
nor NOR2 (N7694, N7690, N2824);
not NOT1 (N7695, N7685);
not NOT1 (N7696, N7693);
nor NOR2 (N7697, N7661, N4819);
and AND2 (N7698, N7694, N6767);
or OR4 (N7699, N7673, N5237, N3272, N4795);
buf BUF1 (N7700, N7696);
or OR3 (N7701, N7698, N133, N3767);
nand NAND3 (N7702, N7699, N1484, N865);
buf BUF1 (N7703, N7701);
nand NAND3 (N7704, N7691, N4936, N4622);
and AND4 (N7705, N7704, N2684, N6109, N6195);
or OR3 (N7706, N7678, N5790, N3066);
xor XOR2 (N7707, N7687, N96);
not NOT1 (N7708, N7697);
or OR3 (N7709, N7708, N437, N1062);
nor NOR2 (N7710, N7705, N1336);
nand NAND3 (N7711, N7702, N4816, N5006);
nor NOR2 (N7712, N7710, N6956);
xor XOR2 (N7713, N7712, N5800);
xor XOR2 (N7714, N7700, N5114);
xor XOR2 (N7715, N7706, N4629);
nor NOR4 (N7716, N7703, N2871, N4229, N1379);
nor NOR2 (N7717, N7715, N909);
or OR2 (N7718, N7714, N7715);
nor NOR4 (N7719, N7707, N6559, N4866, N1814);
nor NOR3 (N7720, N7711, N3643, N5317);
nor NOR2 (N7721, N7692, N7638);
or OR2 (N7722, N7721, N3574);
buf BUF1 (N7723, N7695);
xor XOR2 (N7724, N7723, N4978);
or OR2 (N7725, N7719, N759);
nor NOR2 (N7726, N7716, N3071);
not NOT1 (N7727, N7713);
buf BUF1 (N7728, N7724);
not NOT1 (N7729, N7709);
nand NAND2 (N7730, N7725, N73);
nand NAND3 (N7731, N7717, N1391, N4884);
buf BUF1 (N7732, N7730);
or OR2 (N7733, N7728, N2883);
nand NAND3 (N7734, N7731, N6746, N1401);
and AND4 (N7735, N7726, N3064, N3261, N1824);
xor XOR2 (N7736, N7727, N6868);
and AND4 (N7737, N7672, N4116, N5985, N4445);
xor XOR2 (N7738, N7718, N1512);
not NOT1 (N7739, N7720);
xor XOR2 (N7740, N7722, N1175);
or OR2 (N7741, N7732, N2748);
or OR4 (N7742, N7741, N281, N5312, N7260);
and AND4 (N7743, N7739, N5699, N6850, N5458);
and AND3 (N7744, N7743, N1398, N5847);
xor XOR2 (N7745, N7735, N5816);
nor NOR4 (N7746, N7745, N415, N4744, N5084);
or OR3 (N7747, N7729, N6256, N335);
and AND3 (N7748, N7747, N1926, N5138);
or OR3 (N7749, N7738, N666, N4789);
and AND3 (N7750, N7744, N7494, N5265);
nand NAND4 (N7751, N7750, N6101, N4610, N207);
xor XOR2 (N7752, N7742, N1355);
and AND4 (N7753, N7734, N3729, N1048, N5878);
not NOT1 (N7754, N7751);
or OR2 (N7755, N7746, N4143);
xor XOR2 (N7756, N7740, N3810);
nor NOR3 (N7757, N7748, N3826, N786);
or OR2 (N7758, N7733, N5042);
and AND3 (N7759, N7757, N6719, N849);
nand NAND4 (N7760, N7758, N7639, N7336, N1830);
nor NOR3 (N7761, N7759, N2800, N4718);
buf BUF1 (N7762, N7737);
xor XOR2 (N7763, N7753, N4436);
nand NAND3 (N7764, N7736, N793, N6763);
nor NOR3 (N7765, N7763, N2127, N3373);
nand NAND2 (N7766, N7749, N1463);
not NOT1 (N7767, N7766);
buf BUF1 (N7768, N7760);
xor XOR2 (N7769, N7764, N3446);
and AND4 (N7770, N7765, N2909, N1508, N5687);
and AND3 (N7771, N7752, N5773, N7172);
and AND3 (N7772, N7762, N344, N1329);
not NOT1 (N7773, N7756);
nor NOR3 (N7774, N7768, N2028, N6536);
xor XOR2 (N7775, N7754, N780);
nand NAND4 (N7776, N7769, N2204, N492, N4334);
xor XOR2 (N7777, N7767, N2621);
xor XOR2 (N7778, N7772, N481);
buf BUF1 (N7779, N7778);
or OR2 (N7780, N7779, N7115);
or OR3 (N7781, N7773, N1412, N1782);
nor NOR3 (N7782, N7774, N1048, N7552);
nand NAND2 (N7783, N7781, N1105);
buf BUF1 (N7784, N7775);
not NOT1 (N7785, N7783);
buf BUF1 (N7786, N7785);
nor NOR2 (N7787, N7755, N4240);
and AND4 (N7788, N7761, N6644, N2161, N6474);
and AND3 (N7789, N7787, N6500, N1917);
nand NAND2 (N7790, N7770, N3520);
nor NOR3 (N7791, N7789, N6718, N697);
xor XOR2 (N7792, N7782, N4761);
xor XOR2 (N7793, N7780, N6605);
not NOT1 (N7794, N7784);
nand NAND3 (N7795, N7786, N1698, N4441);
or OR3 (N7796, N7771, N3660, N1421);
or OR2 (N7797, N7795, N7615);
xor XOR2 (N7798, N7791, N7114);
nor NOR2 (N7799, N7793, N5185);
or OR4 (N7800, N7796, N697, N6926, N6523);
or OR3 (N7801, N7794, N7123, N2748);
or OR3 (N7802, N7798, N7670, N7701);
xor XOR2 (N7803, N7777, N5528);
or OR3 (N7804, N7801, N2797, N3078);
xor XOR2 (N7805, N7797, N6022);
buf BUF1 (N7806, N7800);
nor NOR2 (N7807, N7805, N3625);
nor NOR4 (N7808, N7806, N6382, N6077, N4485);
xor XOR2 (N7809, N7799, N3889);
xor XOR2 (N7810, N7792, N4587);
not NOT1 (N7811, N7803);
nor NOR2 (N7812, N7804, N2353);
xor XOR2 (N7813, N7809, N5959);
xor XOR2 (N7814, N7807, N6146);
buf BUF1 (N7815, N7790);
buf BUF1 (N7816, N7811);
not NOT1 (N7817, N7802);
buf BUF1 (N7818, N7815);
nand NAND3 (N7819, N7812, N5058, N7817);
not NOT1 (N7820, N7331);
nor NOR4 (N7821, N7776, N5966, N2199, N5934);
nand NAND2 (N7822, N7813, N1687);
xor XOR2 (N7823, N7788, N6453);
or OR3 (N7824, N7821, N1510, N6461);
xor XOR2 (N7825, N7820, N5845);
buf BUF1 (N7826, N7814);
xor XOR2 (N7827, N7825, N1944);
buf BUF1 (N7828, N7826);
or OR3 (N7829, N7818, N1350, N5147);
nor NOR4 (N7830, N7824, N6076, N2392, N1553);
buf BUF1 (N7831, N7829);
nor NOR4 (N7832, N7810, N402, N5507, N6275);
nand NAND4 (N7833, N7832, N4364, N1840, N3446);
buf BUF1 (N7834, N7833);
nand NAND2 (N7835, N7822, N6396);
nor NOR4 (N7836, N7830, N6099, N4884, N4942);
not NOT1 (N7837, N7828);
or OR2 (N7838, N7831, N7659);
or OR2 (N7839, N7816, N4651);
or OR3 (N7840, N7835, N626, N3000);
not NOT1 (N7841, N7838);
xor XOR2 (N7842, N7808, N6653);
nor NOR2 (N7843, N7839, N690);
buf BUF1 (N7844, N7840);
and AND2 (N7845, N7823, N977);
xor XOR2 (N7846, N7827, N2948);
buf BUF1 (N7847, N7819);
not NOT1 (N7848, N7845);
or OR2 (N7849, N7848, N4171);
xor XOR2 (N7850, N7844, N2253);
xor XOR2 (N7851, N7836, N6398);
xor XOR2 (N7852, N7842, N6401);
not NOT1 (N7853, N7852);
not NOT1 (N7854, N7849);
buf BUF1 (N7855, N7846);
buf BUF1 (N7856, N7851);
not NOT1 (N7857, N7834);
buf BUF1 (N7858, N7855);
nand NAND4 (N7859, N7856, N1936, N1830, N4221);
nor NOR3 (N7860, N7858, N2124, N3989);
not NOT1 (N7861, N7859);
or OR4 (N7862, N7847, N4014, N635, N3154);
or OR4 (N7863, N7853, N7788, N7767, N3201);
xor XOR2 (N7864, N7863, N4189);
not NOT1 (N7865, N7861);
xor XOR2 (N7866, N7841, N6362);
buf BUF1 (N7867, N7854);
xor XOR2 (N7868, N7843, N847);
xor XOR2 (N7869, N7857, N2729);
or OR3 (N7870, N7868, N627, N7367);
not NOT1 (N7871, N7867);
xor XOR2 (N7872, N7860, N4301);
and AND3 (N7873, N7869, N974, N1772);
and AND3 (N7874, N7872, N7424, N6266);
xor XOR2 (N7875, N7870, N6064);
xor XOR2 (N7876, N7850, N5613);
or OR4 (N7877, N7875, N7608, N7486, N2725);
buf BUF1 (N7878, N7837);
buf BUF1 (N7879, N7876);
not NOT1 (N7880, N7874);
not NOT1 (N7881, N7871);
buf BUF1 (N7882, N7878);
or OR4 (N7883, N7864, N7594, N1556, N2096);
xor XOR2 (N7884, N7879, N7370);
and AND4 (N7885, N7862, N2619, N7707, N7423);
buf BUF1 (N7886, N7881);
or OR2 (N7887, N7880, N3616);
nand NAND3 (N7888, N7886, N6471, N3258);
nand NAND4 (N7889, N7884, N6758, N1420, N186);
nor NOR2 (N7890, N7877, N4717);
xor XOR2 (N7891, N7866, N6042);
and AND4 (N7892, N7885, N1339, N6580, N4503);
buf BUF1 (N7893, N7890);
buf BUF1 (N7894, N7892);
nor NOR4 (N7895, N7873, N3105, N5575, N3649);
not NOT1 (N7896, N7889);
xor XOR2 (N7897, N7882, N6081);
nand NAND3 (N7898, N7897, N2549, N4763);
or OR2 (N7899, N7895, N1962);
nand NAND3 (N7900, N7883, N946, N1713);
xor XOR2 (N7901, N7896, N921);
or OR3 (N7902, N7894, N7397, N4846);
and AND3 (N7903, N7888, N1409, N6030);
nand NAND3 (N7904, N7887, N3699, N1444);
nand NAND3 (N7905, N7891, N7156, N5699);
or OR4 (N7906, N7905, N33, N2110, N1001);
nand NAND4 (N7907, N7904, N2789, N3128, N4092);
nand NAND3 (N7908, N7865, N1237, N2074);
xor XOR2 (N7909, N7902, N4356);
buf BUF1 (N7910, N7903);
xor XOR2 (N7911, N7893, N1577);
nand NAND3 (N7912, N7910, N754, N6713);
nor NOR2 (N7913, N7898, N5730);
nor NOR3 (N7914, N7913, N2257, N4444);
or OR4 (N7915, N7906, N7888, N2988, N377);
nor NOR2 (N7916, N7900, N2619);
and AND2 (N7917, N7901, N2009);
not NOT1 (N7918, N7916);
nor NOR2 (N7919, N7908, N4724);
or OR3 (N7920, N7919, N845, N3075);
and AND4 (N7921, N7920, N6296, N1906, N6949);
not NOT1 (N7922, N7912);
not NOT1 (N7923, N7909);
nor NOR2 (N7924, N7914, N3417);
nand NAND3 (N7925, N7911, N1855, N4263);
and AND3 (N7926, N7917, N7645, N267);
and AND3 (N7927, N7925, N6852, N2941);
xor XOR2 (N7928, N7927, N3163);
and AND2 (N7929, N7899, N3765);
nor NOR3 (N7930, N7923, N2377, N7763);
or OR2 (N7931, N7915, N4370);
xor XOR2 (N7932, N7918, N6540);
nand NAND4 (N7933, N7921, N4310, N7918, N3682);
not NOT1 (N7934, N7929);
or OR4 (N7935, N7907, N4554, N7016, N7887);
nand NAND2 (N7936, N7931, N845);
buf BUF1 (N7937, N7936);
or OR3 (N7938, N7924, N6055, N4654);
or OR2 (N7939, N7933, N255);
and AND2 (N7940, N7922, N11);
xor XOR2 (N7941, N7934, N4119);
nor NOR2 (N7942, N7926, N2945);
or OR3 (N7943, N7930, N6437, N3425);
nand NAND2 (N7944, N7935, N2422);
buf BUF1 (N7945, N7939);
not NOT1 (N7946, N7943);
not NOT1 (N7947, N7938);
xor XOR2 (N7948, N7942, N7773);
nand NAND3 (N7949, N7928, N903, N1189);
not NOT1 (N7950, N7946);
nor NOR3 (N7951, N7948, N6237, N4846);
not NOT1 (N7952, N7937);
nor NOR2 (N7953, N7945, N813);
xor XOR2 (N7954, N7947, N245);
or OR2 (N7955, N7949, N4065);
not NOT1 (N7956, N7932);
nor NOR2 (N7957, N7953, N3673);
and AND2 (N7958, N7954, N4379);
nor NOR3 (N7959, N7940, N6999, N7202);
buf BUF1 (N7960, N7951);
xor XOR2 (N7961, N7950, N1094);
or OR4 (N7962, N7956, N952, N537, N1642);
or OR2 (N7963, N7962, N3909);
not NOT1 (N7964, N7961);
nand NAND2 (N7965, N7959, N7698);
and AND4 (N7966, N7941, N1788, N513, N2490);
buf BUF1 (N7967, N7952);
xor XOR2 (N7968, N7966, N5937);
and AND4 (N7969, N7955, N7284, N5141, N1753);
nand NAND2 (N7970, N7963, N2936);
nand NAND2 (N7971, N7969, N5256);
xor XOR2 (N7972, N7970, N1432);
or OR3 (N7973, N7967, N581, N1781);
xor XOR2 (N7974, N7944, N6004);
xor XOR2 (N7975, N7965, N2747);
nand NAND4 (N7976, N7958, N6882, N1360, N1911);
and AND3 (N7977, N7971, N326, N2961);
or OR2 (N7978, N7973, N5315);
buf BUF1 (N7979, N7960);
not NOT1 (N7980, N7975);
and AND2 (N7981, N7964, N2228);
nand NAND3 (N7982, N7976, N942, N365);
xor XOR2 (N7983, N7972, N2679);
or OR2 (N7984, N7968, N2069);
and AND4 (N7985, N7978, N4730, N6700, N1468);
not NOT1 (N7986, N7957);
buf BUF1 (N7987, N7974);
nand NAND2 (N7988, N7979, N284);
or OR4 (N7989, N7986, N1282, N5511, N913);
xor XOR2 (N7990, N7988, N3999);
not NOT1 (N7991, N7990);
xor XOR2 (N7992, N7987, N2163);
xor XOR2 (N7993, N7992, N5138);
or OR3 (N7994, N7991, N156, N2471);
nand NAND4 (N7995, N7982, N5268, N6512, N6467);
and AND2 (N7996, N7980, N6947);
nor NOR2 (N7997, N7984, N3767);
or OR4 (N7998, N7985, N2372, N1138, N6201);
nand NAND2 (N7999, N7997, N3546);
buf BUF1 (N8000, N7993);
nor NOR2 (N8001, N7994, N5824);
nand NAND4 (N8002, N7981, N1519, N2246, N4524);
nor NOR4 (N8003, N8001, N6873, N4447, N7295);
nand NAND4 (N8004, N7983, N1919, N1012, N6860);
not NOT1 (N8005, N7989);
or OR4 (N8006, N7999, N4330, N3990, N2946);
buf BUF1 (N8007, N7998);
or OR4 (N8008, N8003, N3774, N1136, N4364);
nor NOR3 (N8009, N8002, N4298, N2568);
or OR4 (N8010, N7977, N4315, N3186, N2828);
not NOT1 (N8011, N8000);
xor XOR2 (N8012, N8007, N1741);
not NOT1 (N8013, N8012);
nor NOR3 (N8014, N8005, N1467, N4203);
and AND3 (N8015, N7996, N2199, N1312);
and AND3 (N8016, N8014, N6949, N660);
buf BUF1 (N8017, N8011);
not NOT1 (N8018, N8006);
not NOT1 (N8019, N8013);
or OR2 (N8020, N8016, N3367);
xor XOR2 (N8021, N8018, N5530);
xor XOR2 (N8022, N7995, N2952);
nand NAND3 (N8023, N8021, N4713, N303);
not NOT1 (N8024, N8008);
and AND3 (N8025, N8010, N348, N3797);
xor XOR2 (N8026, N8015, N6703);
nand NAND4 (N8027, N8026, N2615, N2939, N7055);
and AND3 (N8028, N8025, N1693, N5630);
xor XOR2 (N8029, N8028, N5441);
nand NAND2 (N8030, N8017, N2393);
or OR2 (N8031, N8029, N6792);
nor NOR3 (N8032, N8031, N2872, N6259);
xor XOR2 (N8033, N8022, N5761);
and AND2 (N8034, N8020, N6149);
buf BUF1 (N8035, N8009);
buf BUF1 (N8036, N8035);
xor XOR2 (N8037, N8034, N5601);
xor XOR2 (N8038, N8024, N5341);
buf BUF1 (N8039, N8032);
xor XOR2 (N8040, N8033, N1784);
xor XOR2 (N8041, N8019, N107);
xor XOR2 (N8042, N8038, N3825);
nand NAND3 (N8043, N8030, N1990, N3388);
or OR4 (N8044, N8036, N7678, N3974, N4720);
not NOT1 (N8045, N8027);
not NOT1 (N8046, N8040);
nor NOR4 (N8047, N8004, N553, N6081, N1876);
buf BUF1 (N8048, N8044);
xor XOR2 (N8049, N8042, N4764);
not NOT1 (N8050, N8047);
buf BUF1 (N8051, N8049);
xor XOR2 (N8052, N8048, N5395);
or OR2 (N8053, N8045, N4712);
nor NOR2 (N8054, N8051, N903);
buf BUF1 (N8055, N8053);
or OR4 (N8056, N8055, N2880, N5033, N7024);
and AND3 (N8057, N8050, N1278, N3143);
not NOT1 (N8058, N8039);
or OR2 (N8059, N8046, N3682);
buf BUF1 (N8060, N8058);
not NOT1 (N8061, N8054);
buf BUF1 (N8062, N8041);
xor XOR2 (N8063, N8057, N1996);
buf BUF1 (N8064, N8052);
xor XOR2 (N8065, N8062, N2403);
and AND3 (N8066, N8059, N3875, N4627);
nor NOR2 (N8067, N8061, N5929);
and AND4 (N8068, N8067, N2981, N1757, N4821);
nand NAND4 (N8069, N8068, N7539, N1637, N7795);
buf BUF1 (N8070, N8064);
xor XOR2 (N8071, N8056, N3074);
nand NAND2 (N8072, N8023, N344);
buf BUF1 (N8073, N8063);
nand NAND3 (N8074, N8066, N6543, N2596);
not NOT1 (N8075, N8070);
and AND4 (N8076, N8075, N4210, N7672, N252);
xor XOR2 (N8077, N8060, N453);
xor XOR2 (N8078, N8073, N2752);
not NOT1 (N8079, N8071);
and AND4 (N8080, N8043, N4356, N7142, N5824);
xor XOR2 (N8081, N8078, N6066);
not NOT1 (N8082, N8079);
nand NAND4 (N8083, N8069, N3076, N113, N6744);
or OR3 (N8084, N8081, N5894, N4796);
xor XOR2 (N8085, N8080, N7221);
nand NAND4 (N8086, N8082, N6003, N7542, N1032);
and AND3 (N8087, N8085, N710, N4785);
or OR2 (N8088, N8074, N5870);
xor XOR2 (N8089, N8087, N3960);
or OR3 (N8090, N8077, N5090, N7100);
nand NAND2 (N8091, N8037, N267);
nand NAND3 (N8092, N8089, N7070, N2105);
nor NOR4 (N8093, N8076, N702, N5381, N4825);
buf BUF1 (N8094, N8092);
or OR4 (N8095, N8091, N1586, N2556, N4127);
or OR2 (N8096, N8090, N3038);
nand NAND2 (N8097, N8094, N6183);
and AND3 (N8098, N8095, N6824, N3215);
nor NOR3 (N8099, N8083, N2776, N2398);
or OR3 (N8100, N8098, N4879, N6537);
nor NOR2 (N8101, N8096, N6981);
not NOT1 (N8102, N8100);
nor NOR4 (N8103, N8065, N5739, N2998, N2274);
or OR4 (N8104, N8099, N6845, N6634, N1993);
not NOT1 (N8105, N8103);
or OR3 (N8106, N8093, N4948, N4598);
nand NAND4 (N8107, N8101, N7699, N7217, N7920);
or OR3 (N8108, N8104, N4000, N2023);
not NOT1 (N8109, N8105);
xor XOR2 (N8110, N8086, N5071);
nor NOR4 (N8111, N8097, N5979, N3061, N2082);
nor NOR3 (N8112, N8102, N2851, N1375);
and AND4 (N8113, N8110, N4583, N7153, N3765);
buf BUF1 (N8114, N8113);
nand NAND4 (N8115, N8108, N4634, N193, N2947);
xor XOR2 (N8116, N8109, N4274);
and AND3 (N8117, N8115, N3549, N4995);
and AND4 (N8118, N8084, N2838, N6734, N6414);
and AND4 (N8119, N8118, N7368, N3896, N4879);
or OR2 (N8120, N8112, N7242);
buf BUF1 (N8121, N8117);
or OR4 (N8122, N8072, N6036, N1037, N3546);
and AND2 (N8123, N8119, N2878);
nor NOR4 (N8124, N8121, N7051, N2831, N2275);
not NOT1 (N8125, N8111);
buf BUF1 (N8126, N8120);
xor XOR2 (N8127, N8106, N4630);
xor XOR2 (N8128, N8124, N2010);
xor XOR2 (N8129, N8116, N831);
nor NOR3 (N8130, N8107, N4254, N204);
buf BUF1 (N8131, N8128);
nand NAND4 (N8132, N8114, N7106, N5976, N1074);
not NOT1 (N8133, N8123);
and AND3 (N8134, N8126, N7508, N5979);
not NOT1 (N8135, N8132);
or OR3 (N8136, N8130, N1254, N2914);
or OR4 (N8137, N8127, N1840, N826, N6805);
nand NAND4 (N8138, N8131, N3728, N3936, N6732);
nor NOR3 (N8139, N8133, N2262, N977);
nand NAND3 (N8140, N8129, N1032, N3527);
and AND2 (N8141, N8137, N6515);
or OR4 (N8142, N8134, N1361, N6360, N6305);
or OR3 (N8143, N8141, N7459, N5188);
xor XOR2 (N8144, N8138, N7853);
xor XOR2 (N8145, N8122, N7875);
and AND4 (N8146, N8135, N3979, N1538, N2586);
xor XOR2 (N8147, N8143, N5309);
nand NAND4 (N8148, N8146, N7497, N3012, N4279);
nor NOR2 (N8149, N8125, N1538);
xor XOR2 (N8150, N8139, N4875);
buf BUF1 (N8151, N8148);
and AND4 (N8152, N8145, N1278, N4859, N234);
xor XOR2 (N8153, N8147, N2612);
nand NAND2 (N8154, N8136, N5549);
buf BUF1 (N8155, N8140);
not NOT1 (N8156, N8149);
nand NAND4 (N8157, N8155, N1335, N4405, N1335);
buf BUF1 (N8158, N8150);
or OR3 (N8159, N8156, N6363, N7989);
not NOT1 (N8160, N8151);
xor XOR2 (N8161, N8158, N7613);
nor NOR4 (N8162, N8088, N5993, N4892, N106);
buf BUF1 (N8163, N8142);
buf BUF1 (N8164, N8144);
not NOT1 (N8165, N8161);
nor NOR3 (N8166, N8157, N5384, N25);
or OR4 (N8167, N8165, N4639, N4862, N2114);
nor NOR4 (N8168, N8167, N2579, N900, N7328);
and AND3 (N8169, N8162, N5692, N3214);
nor NOR2 (N8170, N8169, N5056);
buf BUF1 (N8171, N8168);
or OR4 (N8172, N8153, N2187, N4784, N2140);
xor XOR2 (N8173, N8171, N1574);
not NOT1 (N8174, N8152);
nand NAND4 (N8175, N8173, N2349, N3176, N462);
nand NAND2 (N8176, N8166, N3620);
xor XOR2 (N8177, N8164, N7915);
nand NAND4 (N8178, N8160, N8033, N3669, N4720);
not NOT1 (N8179, N8176);
and AND2 (N8180, N8159, N4941);
xor XOR2 (N8181, N8154, N1562);
buf BUF1 (N8182, N8174);
buf BUF1 (N8183, N8180);
xor XOR2 (N8184, N8179, N2792);
nand NAND4 (N8185, N8177, N7222, N1612, N3826);
not NOT1 (N8186, N8182);
nor NOR3 (N8187, N8184, N496, N2053);
nand NAND4 (N8188, N8172, N1365, N552, N3244);
not NOT1 (N8189, N8178);
or OR2 (N8190, N8170, N2232);
buf BUF1 (N8191, N8190);
or OR2 (N8192, N8188, N7820);
xor XOR2 (N8193, N8192, N6773);
not NOT1 (N8194, N8186);
buf BUF1 (N8195, N8163);
not NOT1 (N8196, N8181);
nor NOR4 (N8197, N8185, N3241, N5591, N5974);
not NOT1 (N8198, N8195);
and AND3 (N8199, N8175, N7120, N5348);
xor XOR2 (N8200, N8197, N5799);
nor NOR4 (N8201, N8187, N3707, N5562, N3197);
buf BUF1 (N8202, N8189);
nand NAND2 (N8203, N8198, N574);
not NOT1 (N8204, N8191);
buf BUF1 (N8205, N8183);
and AND3 (N8206, N8196, N6030, N5190);
nand NAND3 (N8207, N8203, N6826, N2832);
buf BUF1 (N8208, N8206);
nor NOR3 (N8209, N8193, N321, N2844);
buf BUF1 (N8210, N8207);
or OR2 (N8211, N8200, N381);
xor XOR2 (N8212, N8202, N3518);
not NOT1 (N8213, N8201);
nand NAND2 (N8214, N8199, N2595);
buf BUF1 (N8215, N8211);
xor XOR2 (N8216, N8209, N3193);
and AND3 (N8217, N8215, N5488, N5616);
buf BUF1 (N8218, N8194);
xor XOR2 (N8219, N8205, N6766);
buf BUF1 (N8220, N8212);
nand NAND2 (N8221, N8204, N2);
not NOT1 (N8222, N8218);
xor XOR2 (N8223, N8216, N275);
and AND3 (N8224, N8221, N1756, N852);
not NOT1 (N8225, N8219);
nand NAND2 (N8226, N8213, N5108);
and AND4 (N8227, N8222, N4186, N213, N4292);
buf BUF1 (N8228, N8227);
buf BUF1 (N8229, N8225);
buf BUF1 (N8230, N8228);
nor NOR3 (N8231, N8223, N6029, N7664);
xor XOR2 (N8232, N8220, N2469);
nand NAND4 (N8233, N8224, N2455, N4774, N8156);
buf BUF1 (N8234, N8214);
xor XOR2 (N8235, N8208, N7695);
nand NAND3 (N8236, N8232, N4310, N1330);
nor NOR2 (N8237, N8234, N7141);
xor XOR2 (N8238, N8236, N1754);
nand NAND3 (N8239, N8235, N3903, N8189);
or OR3 (N8240, N8237, N3394, N2717);
nand NAND4 (N8241, N8238, N6615, N1508, N555);
not NOT1 (N8242, N8210);
not NOT1 (N8243, N8231);
not NOT1 (N8244, N8241);
xor XOR2 (N8245, N8243, N2461);
and AND2 (N8246, N8240, N5513);
and AND4 (N8247, N8242, N8200, N7447, N7002);
xor XOR2 (N8248, N8245, N4212);
nand NAND4 (N8249, N8226, N3661, N1452, N7586);
not NOT1 (N8250, N8247);
buf BUF1 (N8251, N8230);
not NOT1 (N8252, N8246);
nand NAND3 (N8253, N8251, N605, N1982);
not NOT1 (N8254, N8250);
nor NOR2 (N8255, N8233, N4417);
or OR2 (N8256, N8244, N5778);
xor XOR2 (N8257, N8249, N2993);
xor XOR2 (N8258, N8256, N751);
buf BUF1 (N8259, N8257);
xor XOR2 (N8260, N8229, N7501);
not NOT1 (N8261, N8239);
or OR2 (N8262, N8259, N4121);
nor NOR4 (N8263, N8248, N7170, N4580, N6613);
xor XOR2 (N8264, N8263, N1526);
or OR2 (N8265, N8264, N3329);
buf BUF1 (N8266, N8258);
not NOT1 (N8267, N8217);
not NOT1 (N8268, N8254);
nor NOR4 (N8269, N8255, N7156, N5743, N4590);
not NOT1 (N8270, N8261);
xor XOR2 (N8271, N8260, N2020);
nand NAND4 (N8272, N8270, N1610, N2599, N1524);
nor NOR4 (N8273, N8262, N6433, N2333, N6926);
and AND2 (N8274, N8265, N3269);
not NOT1 (N8275, N8274);
and AND3 (N8276, N8266, N5992, N521);
xor XOR2 (N8277, N8267, N4976);
buf BUF1 (N8278, N8271);
xor XOR2 (N8279, N8277, N4947);
buf BUF1 (N8280, N8272);
nand NAND2 (N8281, N8280, N8224);
not NOT1 (N8282, N8275);
xor XOR2 (N8283, N8269, N4060);
buf BUF1 (N8284, N8281);
or OR4 (N8285, N8252, N7449, N6979, N1647);
nor NOR2 (N8286, N8284, N1045);
and AND3 (N8287, N8286, N4619, N6020);
or OR2 (N8288, N8253, N5681);
buf BUF1 (N8289, N8278);
or OR2 (N8290, N8288, N638);
xor XOR2 (N8291, N8268, N3092);
nor NOR4 (N8292, N8279, N361, N2950, N7545);
buf BUF1 (N8293, N8291);
xor XOR2 (N8294, N8287, N645);
not NOT1 (N8295, N8282);
nor NOR4 (N8296, N8294, N3369, N6931, N1205);
or OR2 (N8297, N8296, N3261);
nand NAND4 (N8298, N8297, N7021, N4520, N3093);
nand NAND4 (N8299, N8290, N8061, N7883, N3411);
or OR2 (N8300, N8295, N7182);
or OR4 (N8301, N8300, N5382, N4410, N2380);
nand NAND3 (N8302, N8298, N516, N2648);
or OR4 (N8303, N8293, N1316, N1218, N2382);
not NOT1 (N8304, N8283);
buf BUF1 (N8305, N8304);
and AND4 (N8306, N8303, N8087, N4262, N1878);
and AND2 (N8307, N8306, N41);
xor XOR2 (N8308, N8292, N6924);
buf BUF1 (N8309, N8307);
xor XOR2 (N8310, N8276, N7492);
xor XOR2 (N8311, N8302, N774);
xor XOR2 (N8312, N8285, N2736);
nor NOR4 (N8313, N8299, N8156, N6479, N3285);
nand NAND2 (N8314, N8311, N5234);
and AND2 (N8315, N8313, N5893);
not NOT1 (N8316, N8314);
and AND4 (N8317, N8312, N7807, N4239, N503);
xor XOR2 (N8318, N8305, N3243);
nor NOR2 (N8319, N8301, N4596);
xor XOR2 (N8320, N8309, N2557);
nor NOR2 (N8321, N8273, N30);
xor XOR2 (N8322, N8289, N4679);
and AND3 (N8323, N8315, N6575, N695);
and AND4 (N8324, N8319, N4090, N3275, N111);
or OR4 (N8325, N8321, N5119, N7217, N6970);
not NOT1 (N8326, N8324);
or OR4 (N8327, N8325, N4524, N7008, N8086);
or OR4 (N8328, N8317, N4769, N6906, N6634);
buf BUF1 (N8329, N8318);
xor XOR2 (N8330, N8329, N3);
not NOT1 (N8331, N8326);
not NOT1 (N8332, N8308);
nand NAND4 (N8333, N8320, N6694, N5870, N2155);
not NOT1 (N8334, N8316);
not NOT1 (N8335, N8310);
buf BUF1 (N8336, N8322);
xor XOR2 (N8337, N8323, N5310);
and AND3 (N8338, N8332, N5080, N7220);
xor XOR2 (N8339, N8328, N1363);
and AND3 (N8340, N8330, N4690, N6394);
or OR4 (N8341, N8340, N3840, N4120, N2378);
buf BUF1 (N8342, N8331);
buf BUF1 (N8343, N8337);
xor XOR2 (N8344, N8336, N1251);
nor NOR3 (N8345, N8341, N2762, N5967);
nand NAND2 (N8346, N8333, N2287);
xor XOR2 (N8347, N8327, N6100);
and AND3 (N8348, N8334, N3167, N747);
not NOT1 (N8349, N8343);
buf BUF1 (N8350, N8342);
or OR2 (N8351, N8349, N7670);
and AND3 (N8352, N8345, N4011, N3157);
xor XOR2 (N8353, N8347, N1794);
buf BUF1 (N8354, N8351);
or OR4 (N8355, N8346, N7983, N7843, N5441);
and AND2 (N8356, N8335, N143);
not NOT1 (N8357, N8356);
nand NAND3 (N8358, N8353, N1849, N4545);
and AND2 (N8359, N8352, N1038);
nand NAND2 (N8360, N8355, N6234);
nand NAND3 (N8361, N8354, N4983, N1687);
or OR4 (N8362, N8360, N6899, N7178, N3120);
nor NOR4 (N8363, N8357, N4285, N822, N3189);
xor XOR2 (N8364, N8361, N409);
and AND4 (N8365, N8363, N6113, N3064, N6424);
nor NOR4 (N8366, N8348, N5995, N4788, N7026);
xor XOR2 (N8367, N8359, N2900);
or OR4 (N8368, N8344, N68, N338, N2295);
nor NOR3 (N8369, N8368, N1286, N4130);
nand NAND4 (N8370, N8339, N7823, N6200, N5875);
and AND3 (N8371, N8358, N5225, N735);
nor NOR3 (N8372, N8367, N5289, N3630);
nor NOR4 (N8373, N8369, N4985, N7474, N2187);
xor XOR2 (N8374, N8338, N7203);
xor XOR2 (N8375, N8350, N6389);
nand NAND3 (N8376, N8373, N1703, N5565);
not NOT1 (N8377, N8370);
or OR3 (N8378, N8374, N472, N3924);
and AND4 (N8379, N8377, N2700, N4630, N1606);
buf BUF1 (N8380, N8364);
not NOT1 (N8381, N8375);
and AND3 (N8382, N8366, N1575, N566);
not NOT1 (N8383, N8365);
and AND2 (N8384, N8383, N6845);
xor XOR2 (N8385, N8372, N5923);
not NOT1 (N8386, N8378);
nand NAND3 (N8387, N8384, N8168, N715);
xor XOR2 (N8388, N8387, N507);
xor XOR2 (N8389, N8382, N2686);
xor XOR2 (N8390, N8388, N848);
nand NAND3 (N8391, N8381, N5666, N4713);
or OR3 (N8392, N8371, N3821, N7026);
nand NAND2 (N8393, N8376, N2951);
nand NAND3 (N8394, N8386, N7294, N740);
buf BUF1 (N8395, N8391);
not NOT1 (N8396, N8379);
not NOT1 (N8397, N8394);
nor NOR3 (N8398, N8380, N1207, N6840);
buf BUF1 (N8399, N8392);
nor NOR4 (N8400, N8385, N834, N6721, N7322);
not NOT1 (N8401, N8396);
nand NAND3 (N8402, N8393, N7227, N2333);
nand NAND3 (N8403, N8399, N6269, N4785);
or OR2 (N8404, N8403, N1073);
xor XOR2 (N8405, N8401, N6367);
xor XOR2 (N8406, N8362, N8321);
or OR3 (N8407, N8397, N4384, N7960);
nor NOR3 (N8408, N8390, N114, N1423);
xor XOR2 (N8409, N8406, N3307);
xor XOR2 (N8410, N8398, N8248);
not NOT1 (N8411, N8400);
nor NOR4 (N8412, N8410, N6235, N6579, N2776);
not NOT1 (N8413, N8409);
and AND3 (N8414, N8408, N2171, N4067);
and AND4 (N8415, N8413, N5562, N3136, N8107);
or OR4 (N8416, N8411, N6928, N4895, N1568);
or OR3 (N8417, N8412, N288, N2094);
xor XOR2 (N8418, N8389, N942);
buf BUF1 (N8419, N8416);
nand NAND3 (N8420, N8415, N445, N4289);
nor NOR3 (N8421, N8418, N7431, N3513);
not NOT1 (N8422, N8420);
or OR2 (N8423, N8407, N542);
nor NOR3 (N8424, N8422, N4740, N7341);
not NOT1 (N8425, N8395);
not NOT1 (N8426, N8402);
nor NOR2 (N8427, N8414, N131);
and AND4 (N8428, N8424, N6821, N4063, N3302);
nand NAND4 (N8429, N8423, N548, N1227, N814);
and AND4 (N8430, N8426, N2438, N2958, N3095);
or OR3 (N8431, N8417, N4887, N2473);
and AND2 (N8432, N8425, N6055);
nor NOR4 (N8433, N8428, N60, N3239, N6864);
xor XOR2 (N8434, N8421, N3476);
buf BUF1 (N8435, N8430);
xor XOR2 (N8436, N8404, N5128);
and AND4 (N8437, N8405, N2260, N4960, N121);
nand NAND2 (N8438, N8419, N5439);
and AND4 (N8439, N8432, N199, N3853, N5145);
not NOT1 (N8440, N8434);
nand NAND4 (N8441, N8429, N4147, N3216, N8134);
buf BUF1 (N8442, N8427);
or OR2 (N8443, N8437, N4361);
or OR4 (N8444, N8438, N3166, N4095, N5940);
and AND3 (N8445, N8439, N7128, N4886);
nor NOR4 (N8446, N8445, N5248, N3178, N6791);
buf BUF1 (N8447, N8446);
nand NAND3 (N8448, N8442, N4982, N2917);
and AND2 (N8449, N8435, N4865);
or OR2 (N8450, N8436, N7286);
or OR4 (N8451, N8449, N3763, N2554, N4828);
buf BUF1 (N8452, N8431);
and AND2 (N8453, N8440, N5719);
buf BUF1 (N8454, N8448);
xor XOR2 (N8455, N8443, N5165);
nor NOR3 (N8456, N8450, N1872, N3171);
or OR2 (N8457, N8447, N8423);
nor NOR2 (N8458, N8457, N7290);
nor NOR2 (N8459, N8453, N7071);
nor NOR2 (N8460, N8459, N3727);
and AND3 (N8461, N8455, N5712, N1396);
nor NOR2 (N8462, N8456, N2797);
nor NOR3 (N8463, N8454, N6331, N5957);
xor XOR2 (N8464, N8451, N7911);
or OR3 (N8465, N8441, N4667, N8071);
not NOT1 (N8466, N8461);
not NOT1 (N8467, N8452);
xor XOR2 (N8468, N8458, N8013);
xor XOR2 (N8469, N8444, N3282);
nand NAND2 (N8470, N8468, N7850);
buf BUF1 (N8471, N8433);
nor NOR3 (N8472, N8463, N7981, N1914);
and AND3 (N8473, N8471, N5021, N4254);
nor NOR2 (N8474, N8472, N8017);
nand NAND3 (N8475, N8474, N3160, N2249);
or OR2 (N8476, N8475, N5676);
not NOT1 (N8477, N8466);
or OR2 (N8478, N8460, N3319);
and AND2 (N8479, N8473, N2440);
not NOT1 (N8480, N8476);
or OR4 (N8481, N8478, N6207, N4870, N2280);
or OR3 (N8482, N8462, N6285, N6967);
nor NOR3 (N8483, N8465, N2967, N570);
not NOT1 (N8484, N8479);
not NOT1 (N8485, N8484);
not NOT1 (N8486, N8480);
and AND4 (N8487, N8486, N4854, N5079, N7005);
buf BUF1 (N8488, N8464);
buf BUF1 (N8489, N8483);
not NOT1 (N8490, N8481);
nor NOR2 (N8491, N8477, N7406);
and AND3 (N8492, N8487, N8368, N6771);
nand NAND2 (N8493, N8488, N2542);
nor NOR2 (N8494, N8490, N6582);
xor XOR2 (N8495, N8470, N5078);
and AND4 (N8496, N8495, N6669, N8280, N8158);
nor NOR2 (N8497, N8467, N4395);
xor XOR2 (N8498, N8497, N8438);
or OR3 (N8499, N8485, N7348, N7400);
not NOT1 (N8500, N8489);
nand NAND4 (N8501, N8491, N3760, N7986, N5279);
not NOT1 (N8502, N8501);
xor XOR2 (N8503, N8482, N4164);
not NOT1 (N8504, N8499);
nor NOR2 (N8505, N8493, N6720);
xor XOR2 (N8506, N8492, N4332);
or OR3 (N8507, N8494, N4722, N4519);
buf BUF1 (N8508, N8505);
buf BUF1 (N8509, N8498);
nor NOR4 (N8510, N8509, N6447, N1128, N5684);
nand NAND2 (N8511, N8496, N7911);
not NOT1 (N8512, N8504);
xor XOR2 (N8513, N8469, N580);
nand NAND4 (N8514, N8510, N7717, N8386, N7317);
nor NOR4 (N8515, N8502, N4154, N7390, N875);
xor XOR2 (N8516, N8503, N4232);
not NOT1 (N8517, N8508);
nand NAND2 (N8518, N8516, N591);
not NOT1 (N8519, N8511);
nand NAND3 (N8520, N8514, N599, N7345);
and AND3 (N8521, N8518, N6405, N230);
nand NAND4 (N8522, N8507, N1865, N7505, N407);
nand NAND3 (N8523, N8521, N1596, N2665);
or OR3 (N8524, N8520, N991, N6157);
nand NAND4 (N8525, N8515, N8499, N1945, N3622);
buf BUF1 (N8526, N8506);
xor XOR2 (N8527, N8517, N5513);
or OR2 (N8528, N8500, N5821);
buf BUF1 (N8529, N8522);
buf BUF1 (N8530, N8529);
nand NAND2 (N8531, N8524, N8468);
nand NAND2 (N8532, N8512, N5464);
xor XOR2 (N8533, N8528, N3101);
not NOT1 (N8534, N8527);
not NOT1 (N8535, N8534);
buf BUF1 (N8536, N8531);
or OR2 (N8537, N8533, N2859);
nor NOR2 (N8538, N8532, N12);
buf BUF1 (N8539, N8535);
buf BUF1 (N8540, N8519);
xor XOR2 (N8541, N8526, N6374);
and AND2 (N8542, N8513, N1706);
and AND3 (N8543, N8536, N6702, N6703);
or OR2 (N8544, N8540, N24);
not NOT1 (N8545, N8523);
nand NAND3 (N8546, N8542, N7448, N4311);
buf BUF1 (N8547, N8544);
nor NOR3 (N8548, N8541, N434, N3955);
nor NOR3 (N8549, N8538, N4310, N1739);
xor XOR2 (N8550, N8525, N5787);
nor NOR3 (N8551, N8543, N5951, N2567);
and AND2 (N8552, N8546, N1595);
or OR2 (N8553, N8537, N8076);
buf BUF1 (N8554, N8549);
buf BUF1 (N8555, N8554);
and AND4 (N8556, N8539, N8418, N5640, N100);
not NOT1 (N8557, N8552);
or OR2 (N8558, N8550, N8327);
or OR2 (N8559, N8553, N1040);
nor NOR4 (N8560, N8558, N4826, N8445, N4911);
buf BUF1 (N8561, N8548);
nor NOR3 (N8562, N8559, N3114, N1549);
not NOT1 (N8563, N8556);
and AND2 (N8564, N8555, N1200);
nand NAND2 (N8565, N8564, N6290);
buf BUF1 (N8566, N8545);
not NOT1 (N8567, N8562);
not NOT1 (N8568, N8551);
buf BUF1 (N8569, N8565);
nand NAND2 (N8570, N8530, N4430);
not NOT1 (N8571, N8561);
or OR2 (N8572, N8547, N6500);
xor XOR2 (N8573, N8557, N5261);
xor XOR2 (N8574, N8569, N1931);
xor XOR2 (N8575, N8566, N1288);
not NOT1 (N8576, N8568);
nand NAND2 (N8577, N8573, N7918);
and AND4 (N8578, N8570, N3139, N4856, N288);
nand NAND4 (N8579, N8576, N4183, N1698, N5221);
or OR2 (N8580, N8574, N8372);
nor NOR2 (N8581, N8579, N8544);
nor NOR3 (N8582, N8577, N7571, N1583);
or OR2 (N8583, N8582, N4369);
and AND2 (N8584, N8578, N7632);
not NOT1 (N8585, N8575);
xor XOR2 (N8586, N8571, N7377);
nor NOR4 (N8587, N8581, N5994, N7201, N6698);
not NOT1 (N8588, N8585);
nand NAND2 (N8589, N8580, N5734);
not NOT1 (N8590, N8586);
xor XOR2 (N8591, N8590, N2925);
or OR2 (N8592, N8583, N1280);
nand NAND4 (N8593, N8567, N5197, N3880, N1349);
nor NOR3 (N8594, N8588, N1475, N8218);
nand NAND2 (N8595, N8589, N8067);
nand NAND4 (N8596, N8560, N7642, N7540, N3135);
nand NAND2 (N8597, N8592, N4214);
not NOT1 (N8598, N8584);
and AND3 (N8599, N8591, N2698, N5829);
or OR4 (N8600, N8587, N8264, N8269, N5984);
or OR3 (N8601, N8594, N1156, N2634);
or OR2 (N8602, N8601, N5284);
nand NAND3 (N8603, N8597, N5936, N4630);
or OR2 (N8604, N8600, N6010);
nor NOR3 (N8605, N8599, N3515, N7069);
not NOT1 (N8606, N8593);
not NOT1 (N8607, N8596);
and AND3 (N8608, N8598, N4731, N1506);
or OR4 (N8609, N8606, N852, N7460, N6359);
and AND3 (N8610, N8605, N1522, N1126);
nand NAND3 (N8611, N8602, N7320, N4333);
xor XOR2 (N8612, N8608, N3027);
and AND2 (N8613, N8604, N8005);
xor XOR2 (N8614, N8609, N3319);
or OR2 (N8615, N8610, N599);
nand NAND3 (N8616, N8614, N2883, N5395);
nand NAND4 (N8617, N8607, N6099, N8081, N841);
or OR3 (N8618, N8617, N4060, N3562);
or OR2 (N8619, N8603, N3501);
xor XOR2 (N8620, N8613, N3994);
not NOT1 (N8621, N8612);
not NOT1 (N8622, N8621);
and AND2 (N8623, N8615, N8338);
or OR4 (N8624, N8616, N8446, N4449, N7736);
or OR2 (N8625, N8611, N711);
and AND3 (N8626, N8563, N6248, N747);
nand NAND2 (N8627, N8626, N7258);
buf BUF1 (N8628, N8627);
xor XOR2 (N8629, N8622, N4388);
or OR3 (N8630, N8625, N2494, N7809);
and AND4 (N8631, N8624, N5064, N8270, N4450);
nor NOR2 (N8632, N8620, N8430);
nand NAND2 (N8633, N8631, N7152);
or OR2 (N8634, N8623, N4392);
nand NAND3 (N8635, N8619, N8428, N3484);
nand NAND2 (N8636, N8595, N4983);
xor XOR2 (N8637, N8636, N8234);
not NOT1 (N8638, N8618);
and AND2 (N8639, N8634, N3218);
and AND4 (N8640, N8638, N4670, N5565, N6866);
nor NOR3 (N8641, N8632, N4727, N8117);
buf BUF1 (N8642, N8635);
not NOT1 (N8643, N8629);
nor NOR4 (N8644, N8643, N3356, N7958, N4268);
not NOT1 (N8645, N8572);
xor XOR2 (N8646, N8630, N334);
nand NAND3 (N8647, N8637, N722, N289);
and AND3 (N8648, N8645, N858, N7501);
nand NAND2 (N8649, N8648, N4049);
not NOT1 (N8650, N8646);
not NOT1 (N8651, N8641);
nand NAND3 (N8652, N8650, N796, N3529);
and AND2 (N8653, N8649, N6234);
nor NOR2 (N8654, N8647, N6916);
buf BUF1 (N8655, N8653);
and AND4 (N8656, N8654, N7009, N5925, N6816);
nand NAND3 (N8657, N8656, N8170, N6969);
nor NOR4 (N8658, N8640, N5525, N241, N588);
not NOT1 (N8659, N8657);
not NOT1 (N8660, N8655);
or OR2 (N8661, N8633, N685);
buf BUF1 (N8662, N8658);
and AND3 (N8663, N8628, N1206, N545);
nand NAND2 (N8664, N8644, N6792);
and AND4 (N8665, N8663, N8542, N392, N8244);
not NOT1 (N8666, N8652);
nand NAND4 (N8667, N8639, N2565, N2685, N8646);
or OR3 (N8668, N8667, N7268, N1359);
or OR3 (N8669, N8666, N8471, N8287);
buf BUF1 (N8670, N8651);
nand NAND3 (N8671, N8664, N3060, N2342);
buf BUF1 (N8672, N8671);
nor NOR3 (N8673, N8660, N7041, N5766);
not NOT1 (N8674, N8670);
not NOT1 (N8675, N8673);
or OR4 (N8676, N8659, N3688, N2738, N4778);
nor NOR3 (N8677, N8642, N4528, N3020);
not NOT1 (N8678, N8676);
xor XOR2 (N8679, N8678, N3449);
or OR3 (N8680, N8668, N953, N7584);
buf BUF1 (N8681, N8672);
and AND3 (N8682, N8669, N3923, N5891);
buf BUF1 (N8683, N8665);
nand NAND3 (N8684, N8674, N3520, N3838);
xor XOR2 (N8685, N8675, N7070);
buf BUF1 (N8686, N8685);
not NOT1 (N8687, N8679);
not NOT1 (N8688, N8681);
or OR3 (N8689, N8662, N8638, N2340);
not NOT1 (N8690, N8682);
and AND2 (N8691, N8686, N6206);
nor NOR4 (N8692, N8677, N7340, N6308, N3593);
nor NOR2 (N8693, N8684, N7391);
or OR4 (N8694, N8688, N2935, N5031, N1702);
or OR3 (N8695, N8690, N7558, N4830);
or OR4 (N8696, N8695, N1454, N4533, N2949);
not NOT1 (N8697, N8693);
buf BUF1 (N8698, N8683);
and AND3 (N8699, N8687, N8546, N2692);
xor XOR2 (N8700, N8696, N8492);
nand NAND3 (N8701, N8680, N3353, N7314);
buf BUF1 (N8702, N8692);
and AND4 (N8703, N8698, N2104, N1105, N2164);
and AND4 (N8704, N8661, N2265, N1405, N1670);
buf BUF1 (N8705, N8701);
xor XOR2 (N8706, N8704, N2841);
buf BUF1 (N8707, N8689);
or OR4 (N8708, N8699, N7283, N7273, N4905);
buf BUF1 (N8709, N8697);
and AND4 (N8710, N8707, N2761, N1712, N2496);
nor NOR3 (N8711, N8705, N7847, N4082);
and AND4 (N8712, N8706, N6465, N1875, N1020);
xor XOR2 (N8713, N8711, N4303);
nor NOR4 (N8714, N8713, N4714, N7177, N6495);
and AND4 (N8715, N8714, N8183, N5339, N6527);
or OR2 (N8716, N8715, N3139);
nand NAND4 (N8717, N8703, N173, N2464, N1572);
nor NOR4 (N8718, N8712, N3698, N5356, N6255);
and AND4 (N8719, N8710, N2248, N6364, N7566);
nor NOR4 (N8720, N8694, N5235, N6663, N8316);
xor XOR2 (N8721, N8708, N2523);
nand NAND3 (N8722, N8721, N7332, N1971);
or OR4 (N8723, N8716, N7337, N6809, N4644);
xor XOR2 (N8724, N8723, N8477);
xor XOR2 (N8725, N8724, N3620);
nor NOR4 (N8726, N8717, N6159, N6551, N2067);
or OR2 (N8727, N8691, N287);
not NOT1 (N8728, N8719);
and AND2 (N8729, N8725, N8580);
xor XOR2 (N8730, N8718, N6591);
buf BUF1 (N8731, N8728);
not NOT1 (N8732, N8730);
xor XOR2 (N8733, N8726, N4859);
nor NOR4 (N8734, N8720, N144, N6864, N7111);
and AND3 (N8735, N8731, N1938, N4701);
and AND3 (N8736, N8700, N4709, N5946);
not NOT1 (N8737, N8734);
and AND4 (N8738, N8733, N5778, N4236, N5000);
nand NAND3 (N8739, N8727, N3447, N5592);
not NOT1 (N8740, N8702);
buf BUF1 (N8741, N8709);
or OR3 (N8742, N8740, N1890, N5104);
and AND4 (N8743, N8729, N152, N1540, N2816);
nor NOR4 (N8744, N8736, N5715, N8458, N2422);
nand NAND4 (N8745, N8742, N8183, N5838, N8283);
not NOT1 (N8746, N8743);
not NOT1 (N8747, N8745);
and AND2 (N8748, N8739, N3799);
or OR4 (N8749, N8732, N1536, N4166, N3752);
nand NAND2 (N8750, N8748, N2220);
xor XOR2 (N8751, N8738, N6801);
not NOT1 (N8752, N8746);
buf BUF1 (N8753, N8752);
and AND4 (N8754, N8741, N6256, N3456, N8422);
nand NAND2 (N8755, N8737, N6680);
buf BUF1 (N8756, N8751);
buf BUF1 (N8757, N8744);
nor NOR3 (N8758, N8722, N8142, N7674);
or OR2 (N8759, N8749, N6763);
xor XOR2 (N8760, N8754, N8515);
nand NAND2 (N8761, N8747, N803);
xor XOR2 (N8762, N8755, N2526);
not NOT1 (N8763, N8758);
nor NOR4 (N8764, N8753, N8023, N1091, N1435);
nand NAND2 (N8765, N8761, N4205);
nor NOR2 (N8766, N8763, N3549);
buf BUF1 (N8767, N8764);
not NOT1 (N8768, N8767);
nor NOR2 (N8769, N8735, N4929);
not NOT1 (N8770, N8750);
nor NOR4 (N8771, N8760, N7773, N1123, N3702);
nand NAND4 (N8772, N8757, N681, N1355, N533);
nand NAND3 (N8773, N8765, N5900, N1698);
xor XOR2 (N8774, N8766, N8237);
nor NOR4 (N8775, N8770, N2521, N4495, N4072);
buf BUF1 (N8776, N8769);
buf BUF1 (N8777, N8771);
or OR2 (N8778, N8762, N1585);
and AND2 (N8779, N8776, N5480);
or OR3 (N8780, N8773, N4678, N7977);
and AND3 (N8781, N8768, N1309, N2247);
not NOT1 (N8782, N8772);
xor XOR2 (N8783, N8759, N137);
nand NAND4 (N8784, N8782, N5992, N6485, N3095);
or OR2 (N8785, N8775, N1487);
xor XOR2 (N8786, N8777, N3747);
nor NOR3 (N8787, N8774, N2870, N2827);
and AND4 (N8788, N8783, N1930, N4925, N8631);
not NOT1 (N8789, N8781);
nand NAND4 (N8790, N8789, N3600, N7294, N2928);
not NOT1 (N8791, N8780);
nand NAND4 (N8792, N8787, N7305, N550, N3914);
buf BUF1 (N8793, N8790);
buf BUF1 (N8794, N8778);
nor NOR3 (N8795, N8792, N3848, N7164);
nand NAND2 (N8796, N8756, N2122);
nand NAND2 (N8797, N8779, N6660);
not NOT1 (N8798, N8797);
or OR4 (N8799, N8785, N6220, N498, N3841);
and AND2 (N8800, N8786, N4505);
nor NOR3 (N8801, N8784, N1224, N8746);
buf BUF1 (N8802, N8793);
and AND4 (N8803, N8799, N8120, N4483, N2960);
buf BUF1 (N8804, N8795);
buf BUF1 (N8805, N8803);
nand NAND2 (N8806, N8798, N8149);
nand NAND2 (N8807, N8788, N7885);
and AND4 (N8808, N8800, N976, N5602, N4412);
or OR2 (N8809, N8804, N7732);
buf BUF1 (N8810, N8802);
nand NAND3 (N8811, N8809, N1345, N979);
and AND2 (N8812, N8794, N2121);
nor NOR4 (N8813, N8812, N6974, N1372, N5144);
not NOT1 (N8814, N8791);
nor NOR2 (N8815, N8810, N6445);
not NOT1 (N8816, N8801);
or OR2 (N8817, N8796, N8423);
and AND3 (N8818, N8816, N1036, N4286);
or OR3 (N8819, N8808, N5883, N7053);
not NOT1 (N8820, N8819);
buf BUF1 (N8821, N8820);
or OR4 (N8822, N8815, N1652, N5358, N4824);
or OR3 (N8823, N8806, N4500, N3424);
nand NAND3 (N8824, N8813, N117, N1163);
buf BUF1 (N8825, N8814);
not NOT1 (N8826, N8825);
buf BUF1 (N8827, N8805);
not NOT1 (N8828, N8807);
not NOT1 (N8829, N8828);
nor NOR2 (N8830, N8822, N445);
nand NAND4 (N8831, N8811, N2195, N2291, N5920);
buf BUF1 (N8832, N8831);
xor XOR2 (N8833, N8818, N4561);
nand NAND2 (N8834, N8832, N1887);
buf BUF1 (N8835, N8823);
or OR2 (N8836, N8827, N2667);
nor NOR3 (N8837, N8836, N3438, N5315);
not NOT1 (N8838, N8817);
nor NOR2 (N8839, N8835, N5828);
nand NAND3 (N8840, N8829, N46, N4642);
not NOT1 (N8841, N8821);
xor XOR2 (N8842, N8833, N2357);
buf BUF1 (N8843, N8830);
or OR2 (N8844, N8840, N367);
nor NOR3 (N8845, N8839, N7066, N7946);
xor XOR2 (N8846, N8834, N860);
xor XOR2 (N8847, N8846, N3864);
not NOT1 (N8848, N8824);
not NOT1 (N8849, N8837);
and AND4 (N8850, N8845, N4861, N968, N2185);
and AND4 (N8851, N8826, N2399, N3227, N8096);
xor XOR2 (N8852, N8843, N8022);
and AND4 (N8853, N8844, N4359, N5973, N1233);
and AND4 (N8854, N8853, N5407, N995, N7265);
and AND4 (N8855, N8851, N7410, N1485, N5595);
and AND4 (N8856, N8847, N767, N2818, N6841);
nand NAND3 (N8857, N8841, N1150, N767);
nor NOR4 (N8858, N8857, N4419, N7318, N4456);
buf BUF1 (N8859, N8842);
not NOT1 (N8860, N8852);
nand NAND2 (N8861, N8848, N8592);
and AND3 (N8862, N8856, N6595, N5152);
nand NAND2 (N8863, N8858, N2736);
not NOT1 (N8864, N8849);
nor NOR4 (N8865, N8860, N3744, N4991, N7290);
and AND3 (N8866, N8854, N955, N1529);
or OR3 (N8867, N8855, N6677, N3841);
or OR3 (N8868, N8838, N3153, N7629);
and AND3 (N8869, N8865, N823, N8814);
buf BUF1 (N8870, N8861);
and AND2 (N8871, N8864, N4265);
nor NOR4 (N8872, N8870, N1663, N6430, N7376);
and AND4 (N8873, N8866, N2317, N7592, N6852);
not NOT1 (N8874, N8863);
xor XOR2 (N8875, N8874, N2253);
nand NAND4 (N8876, N8872, N5001, N8868, N4172);
or OR4 (N8877, N7411, N8857, N7086, N7991);
xor XOR2 (N8878, N8877, N2914);
or OR3 (N8879, N8871, N2459, N2288);
and AND2 (N8880, N8873, N4016);
xor XOR2 (N8881, N8876, N2318);
not NOT1 (N8882, N8850);
buf BUF1 (N8883, N8867);
nor NOR4 (N8884, N8881, N4002, N3117, N2122);
and AND2 (N8885, N8880, N5093);
nor NOR4 (N8886, N8878, N6310, N1585, N5286);
nor NOR4 (N8887, N8859, N5390, N4511, N3620);
nand NAND2 (N8888, N8875, N7890);
or OR2 (N8889, N8887, N8226);
buf BUF1 (N8890, N8882);
nand NAND2 (N8891, N8886, N387);
or OR3 (N8892, N8889, N210, N8801);
nor NOR4 (N8893, N8862, N400, N2946, N5171);
not NOT1 (N8894, N8888);
and AND2 (N8895, N8884, N2767);
not NOT1 (N8896, N8890);
or OR4 (N8897, N8893, N7784, N2620, N7019);
or OR3 (N8898, N8883, N5264, N3983);
and AND3 (N8899, N8895, N3191, N7589);
buf BUF1 (N8900, N8896);
nor NOR2 (N8901, N8885, N6717);
and AND4 (N8902, N8900, N7100, N7127, N1858);
or OR4 (N8903, N8879, N8096, N1997, N234);
nand NAND3 (N8904, N8891, N6900, N6732);
nand NAND3 (N8905, N8892, N2748, N4452);
nand NAND2 (N8906, N8902, N1849);
not NOT1 (N8907, N8905);
or OR3 (N8908, N8898, N2173, N7646);
or OR3 (N8909, N8908, N1820, N1661);
or OR4 (N8910, N8894, N2718, N7867, N6193);
nor NOR3 (N8911, N8899, N5545, N384);
buf BUF1 (N8912, N8901);
or OR4 (N8913, N8897, N5864, N485, N748);
not NOT1 (N8914, N8909);
nor NOR4 (N8915, N8911, N2347, N7831, N4254);
nand NAND2 (N8916, N8914, N4715);
not NOT1 (N8917, N8912);
buf BUF1 (N8918, N8910);
nand NAND3 (N8919, N8917, N1438, N8833);
nor NOR4 (N8920, N8916, N7372, N3477, N4283);
nor NOR3 (N8921, N8907, N4280, N6303);
or OR3 (N8922, N8919, N8384, N4646);
or OR4 (N8923, N8920, N2061, N4804, N5009);
nand NAND3 (N8924, N8918, N6210, N2776);
or OR4 (N8925, N8924, N2914, N7922, N3080);
xor XOR2 (N8926, N8925, N617);
nand NAND3 (N8927, N8869, N4787, N4665);
not NOT1 (N8928, N8915);
nor NOR2 (N8929, N8903, N3842);
nand NAND3 (N8930, N8921, N4874, N306);
and AND2 (N8931, N8922, N3317);
buf BUF1 (N8932, N8923);
nor NOR3 (N8933, N8929, N1534, N6402);
buf BUF1 (N8934, N8928);
xor XOR2 (N8935, N8926, N8339);
nand NAND4 (N8936, N8927, N8049, N8564, N1197);
and AND2 (N8937, N8931, N3008);
or OR4 (N8938, N8932, N6572, N7314, N8399);
xor XOR2 (N8939, N8934, N4578);
xor XOR2 (N8940, N8913, N2515);
nor NOR4 (N8941, N8939, N2822, N2980, N3007);
xor XOR2 (N8942, N8937, N7535);
nand NAND2 (N8943, N8930, N8896);
and AND4 (N8944, N8935, N7666, N8145, N2986);
nor NOR3 (N8945, N8936, N6924, N7362);
and AND4 (N8946, N8941, N1034, N775, N2511);
buf BUF1 (N8947, N8933);
not NOT1 (N8948, N8945);
or OR4 (N8949, N8948, N8295, N785, N6577);
buf BUF1 (N8950, N8906);
buf BUF1 (N8951, N8940);
buf BUF1 (N8952, N8946);
nand NAND4 (N8953, N8952, N7243, N7238, N5138);
nor NOR3 (N8954, N8947, N3064, N8502);
and AND4 (N8955, N8949, N7759, N4694, N312);
buf BUF1 (N8956, N8953);
and AND3 (N8957, N8956, N4538, N3175);
or OR2 (N8958, N8955, N5715);
xor XOR2 (N8959, N8954, N5224);
or OR2 (N8960, N8950, N7727);
not NOT1 (N8961, N8960);
not NOT1 (N8962, N8961);
or OR2 (N8963, N8958, N8686);
or OR3 (N8964, N8938, N2401, N6708);
xor XOR2 (N8965, N8943, N8105);
not NOT1 (N8966, N8904);
and AND4 (N8967, N8964, N5853, N1909, N2422);
nand NAND2 (N8968, N8962, N5812);
or OR2 (N8969, N8967, N5404);
and AND4 (N8970, N8965, N1774, N1739, N2169);
not NOT1 (N8971, N8969);
buf BUF1 (N8972, N8944);
buf BUF1 (N8973, N8963);
nand NAND4 (N8974, N8951, N3911, N6195, N5652);
nor NOR3 (N8975, N8942, N1069, N1028);
nor NOR4 (N8976, N8959, N2154, N4917, N3529);
and AND2 (N8977, N8972, N639);
or OR4 (N8978, N8971, N3082, N4344, N3039);
buf BUF1 (N8979, N8978);
not NOT1 (N8980, N8957);
not NOT1 (N8981, N8975);
nand NAND4 (N8982, N8981, N6420, N8344, N1158);
not NOT1 (N8983, N8973);
or OR4 (N8984, N8983, N1170, N6017, N714);
nand NAND4 (N8985, N8982, N1200, N3860, N19);
not NOT1 (N8986, N8985);
xor XOR2 (N8987, N8979, N5448);
xor XOR2 (N8988, N8977, N1799);
buf BUF1 (N8989, N8966);
and AND4 (N8990, N8988, N1491, N6864, N7271);
or OR2 (N8991, N8974, N7713);
or OR4 (N8992, N8976, N4856, N8324, N1846);
xor XOR2 (N8993, N8991, N1263);
not NOT1 (N8994, N8968);
or OR4 (N8995, N8984, N6718, N3189, N8062);
not NOT1 (N8996, N8994);
or OR2 (N8997, N8986, N2405);
xor XOR2 (N8998, N8993, N4664);
and AND2 (N8999, N8997, N1171);
or OR2 (N9000, N8998, N5353);
nand NAND4 (N9001, N9000, N6656, N2650, N7173);
not NOT1 (N9002, N8995);
not NOT1 (N9003, N8989);
or OR2 (N9004, N8987, N3476);
or OR2 (N9005, N8980, N2720);
nand NAND4 (N9006, N8992, N5125, N7013, N4031);
not NOT1 (N9007, N9006);
nor NOR4 (N9008, N9002, N3733, N8430, N5508);
nor NOR2 (N9009, N8999, N5837);
or OR4 (N9010, N8990, N4407, N2567, N3276);
not NOT1 (N9011, N8970);
buf BUF1 (N9012, N9001);
and AND4 (N9013, N9008, N7050, N4004, N1121);
buf BUF1 (N9014, N9013);
and AND2 (N9015, N9012, N3260);
buf BUF1 (N9016, N8996);
not NOT1 (N9017, N9007);
and AND2 (N9018, N9004, N4928);
not NOT1 (N9019, N9014);
buf BUF1 (N9020, N9011);
not NOT1 (N9021, N9017);
nor NOR3 (N9022, N9003, N953, N7516);
nand NAND2 (N9023, N9021, N4977);
nand NAND4 (N9024, N9010, N5075, N4072, N4873);
nand NAND2 (N9025, N9023, N7792);
buf BUF1 (N9026, N9018);
or OR4 (N9027, N9015, N7734, N5272, N2927);
xor XOR2 (N9028, N9026, N4599);
buf BUF1 (N9029, N9020);
buf BUF1 (N9030, N9029);
nand NAND4 (N9031, N9027, N828, N6828, N3361);
nor NOR3 (N9032, N9028, N3810, N7121);
nor NOR2 (N9033, N9009, N1913);
nand NAND3 (N9034, N9019, N2522, N5235);
buf BUF1 (N9035, N9025);
not NOT1 (N9036, N9035);
nand NAND4 (N9037, N9032, N5478, N2456, N6287);
buf BUF1 (N9038, N9031);
nand NAND4 (N9039, N9034, N7671, N5228, N8072);
buf BUF1 (N9040, N9037);
nor NOR3 (N9041, N9022, N1903, N6873);
buf BUF1 (N9042, N9016);
or OR3 (N9043, N9005, N481, N1042);
nand NAND2 (N9044, N9042, N6149);
nand NAND4 (N9045, N9030, N3140, N2177, N8107);
buf BUF1 (N9046, N9044);
xor XOR2 (N9047, N9033, N3524);
or OR2 (N9048, N9040, N6173);
and AND3 (N9049, N9039, N4978, N2631);
xor XOR2 (N9050, N9043, N6460);
or OR2 (N9051, N9050, N7390);
buf BUF1 (N9052, N9046);
nor NOR4 (N9053, N9052, N2928, N1086, N7053);
or OR2 (N9054, N9048, N3437);
nor NOR3 (N9055, N9053, N4125, N7708);
and AND4 (N9056, N9051, N575, N2405, N8325);
nand NAND2 (N9057, N9038, N8067);
buf BUF1 (N9058, N9055);
not NOT1 (N9059, N9024);
nor NOR3 (N9060, N9054, N6414, N602);
buf BUF1 (N9061, N9058);
not NOT1 (N9062, N9036);
not NOT1 (N9063, N9056);
nand NAND4 (N9064, N9041, N396, N6648, N3737);
or OR3 (N9065, N9057, N4206, N6522);
xor XOR2 (N9066, N9065, N5021);
nor NOR3 (N9067, N9064, N9042, N6946);
xor XOR2 (N9068, N9049, N245);
buf BUF1 (N9069, N9062);
and AND2 (N9070, N9047, N6736);
not NOT1 (N9071, N9063);
nand NAND3 (N9072, N9060, N2075, N8440);
or OR3 (N9073, N9069, N5492, N5649);
nand NAND4 (N9074, N9066, N2871, N90, N6713);
buf BUF1 (N9075, N9068);
or OR3 (N9076, N9074, N8501, N8916);
or OR4 (N9077, N9067, N4480, N5180, N1314);
nor NOR3 (N9078, N9073, N5276, N4333);
and AND4 (N9079, N9059, N893, N473, N8748);
nor NOR2 (N9080, N9079, N2951);
or OR4 (N9081, N9071, N636, N4246, N4828);
xor XOR2 (N9082, N9072, N3219);
nand NAND2 (N9083, N9082, N5759);
and AND4 (N9084, N9045, N3413, N9057, N4919);
xor XOR2 (N9085, N9076, N6745);
not NOT1 (N9086, N9081);
not NOT1 (N9087, N9086);
and AND3 (N9088, N9077, N1580, N3167);
nand NAND2 (N9089, N9088, N1304);
not NOT1 (N9090, N9083);
xor XOR2 (N9091, N9075, N8024);
not NOT1 (N9092, N9085);
not NOT1 (N9093, N9090);
not NOT1 (N9094, N9061);
xor XOR2 (N9095, N9078, N1686);
and AND3 (N9096, N9080, N476, N4528);
or OR2 (N9097, N9087, N6519);
xor XOR2 (N9098, N9094, N1102);
not NOT1 (N9099, N9098);
xor XOR2 (N9100, N9089, N6118);
and AND3 (N9101, N9091, N6338, N2756);
or OR3 (N9102, N9093, N5057, N2818);
xor XOR2 (N9103, N9084, N7918);
and AND4 (N9104, N9102, N8018, N511, N6232);
and AND3 (N9105, N9070, N1222, N1558);
buf BUF1 (N9106, N9100);
buf BUF1 (N9107, N9103);
nand NAND3 (N9108, N9107, N6010, N5068);
buf BUF1 (N9109, N9108);
not NOT1 (N9110, N9099);
buf BUF1 (N9111, N9095);
and AND3 (N9112, N9096, N3828, N1283);
not NOT1 (N9113, N9106);
nand NAND2 (N9114, N9109, N6453);
and AND2 (N9115, N9104, N6734);
not NOT1 (N9116, N9111);
not NOT1 (N9117, N9113);
not NOT1 (N9118, N9112);
or OR4 (N9119, N9101, N5899, N7310, N2987);
xor XOR2 (N9120, N9117, N4018);
not NOT1 (N9121, N9119);
buf BUF1 (N9122, N9110);
not NOT1 (N9123, N9122);
nand NAND2 (N9124, N9092, N7940);
or OR3 (N9125, N9105, N931, N2221);
and AND4 (N9126, N9114, N920, N8645, N6759);
or OR3 (N9127, N9115, N2274, N6906);
and AND4 (N9128, N9121, N2403, N4006, N3446);
buf BUF1 (N9129, N9125);
nor NOR3 (N9130, N9116, N2875, N2883);
xor XOR2 (N9131, N9124, N8993);
or OR3 (N9132, N9097, N5157, N4620);
buf BUF1 (N9133, N9132);
nand NAND2 (N9134, N9126, N4896);
or OR3 (N9135, N9129, N6956, N3633);
xor XOR2 (N9136, N9134, N3023);
or OR2 (N9137, N9130, N3103);
nand NAND2 (N9138, N9131, N3954);
and AND3 (N9139, N9133, N2663, N8210);
or OR4 (N9140, N9136, N8017, N3338, N6320);
or OR2 (N9141, N9118, N8793);
nand NAND2 (N9142, N9137, N5747);
or OR3 (N9143, N9140, N958, N6053);
and AND2 (N9144, N9141, N3966);
nand NAND2 (N9145, N9135, N7368);
not NOT1 (N9146, N9123);
xor XOR2 (N9147, N9128, N3788);
buf BUF1 (N9148, N9144);
and AND2 (N9149, N9127, N777);
and AND3 (N9150, N9143, N1070, N5244);
not NOT1 (N9151, N9145);
nand NAND4 (N9152, N9151, N2263, N8316, N3775);
or OR2 (N9153, N9147, N8747);
or OR3 (N9154, N9150, N4955, N8101);
or OR2 (N9155, N9142, N4403);
and AND4 (N9156, N9120, N6971, N2616, N6486);
nand NAND4 (N9157, N9153, N5888, N6335, N161);
or OR3 (N9158, N9139, N2373, N4373);
xor XOR2 (N9159, N9158, N2935);
buf BUF1 (N9160, N9148);
nand NAND2 (N9161, N9146, N6720);
and AND2 (N9162, N9161, N5126);
buf BUF1 (N9163, N9160);
xor XOR2 (N9164, N9155, N2326);
or OR4 (N9165, N9159, N390, N4704, N5299);
nor NOR2 (N9166, N9154, N5137);
xor XOR2 (N9167, N9166, N8877);
nand NAND2 (N9168, N9163, N3163);
nand NAND3 (N9169, N9149, N5425, N673);
nor NOR4 (N9170, N9162, N7530, N5076, N3176);
nand NAND3 (N9171, N9168, N5388, N1557);
nand NAND2 (N9172, N9165, N2678);
buf BUF1 (N9173, N9152);
and AND3 (N9174, N9157, N5320, N2102);
nor NOR3 (N9175, N9169, N7299, N1389);
xor XOR2 (N9176, N9170, N1157);
nand NAND4 (N9177, N9176, N7584, N7842, N4643);
nand NAND2 (N9178, N9174, N460);
or OR2 (N9179, N9173, N4688);
nor NOR4 (N9180, N9138, N2295, N6170, N8593);
and AND3 (N9181, N9175, N8641, N1105);
not NOT1 (N9182, N9181);
or OR2 (N9183, N9156, N3822);
nor NOR2 (N9184, N9182, N5652);
and AND3 (N9185, N9164, N3332, N5466);
xor XOR2 (N9186, N9177, N2132);
nor NOR3 (N9187, N9179, N6235, N3316);
or OR3 (N9188, N9178, N6122, N2568);
nand NAND3 (N9189, N9187, N8553, N1506);
nor NOR3 (N9190, N9172, N5838, N660);
xor XOR2 (N9191, N9188, N1487);
not NOT1 (N9192, N9189);
or OR3 (N9193, N9171, N4344, N3458);
buf BUF1 (N9194, N9167);
nor NOR2 (N9195, N9194, N1726);
nand NAND2 (N9196, N9191, N4447);
xor XOR2 (N9197, N9185, N6462);
or OR3 (N9198, N9186, N3336, N2458);
and AND3 (N9199, N9196, N1623, N4532);
nor NOR2 (N9200, N9180, N534);
buf BUF1 (N9201, N9183);
nor NOR2 (N9202, N9192, N5325);
and AND3 (N9203, N9184, N8760, N4325);
nand NAND2 (N9204, N9190, N8859);
nor NOR4 (N9205, N9204, N7354, N7313, N7437);
not NOT1 (N9206, N9202);
or OR3 (N9207, N9197, N4076, N6958);
and AND2 (N9208, N9193, N8640);
xor XOR2 (N9209, N9203, N1111);
buf BUF1 (N9210, N9208);
or OR4 (N9211, N9206, N7291, N6035, N8993);
not NOT1 (N9212, N9201);
xor XOR2 (N9213, N9195, N7345);
not NOT1 (N9214, N9211);
nor NOR4 (N9215, N9207, N38, N7625, N4976);
xor XOR2 (N9216, N9213, N5420);
buf BUF1 (N9217, N9205);
xor XOR2 (N9218, N9214, N4686);
or OR2 (N9219, N9217, N3281);
nor NOR3 (N9220, N9212, N8015, N8296);
nand NAND2 (N9221, N9215, N1366);
nand NAND4 (N9222, N9216, N2188, N7564, N7659);
not NOT1 (N9223, N9220);
nor NOR3 (N9224, N9221, N6654, N5417);
buf BUF1 (N9225, N9209);
buf BUF1 (N9226, N9218);
xor XOR2 (N9227, N9223, N1018);
or OR4 (N9228, N9227, N5161, N6402, N6946);
and AND3 (N9229, N9198, N8994, N8637);
nor NOR4 (N9230, N9225, N653, N5873, N8776);
nor NOR3 (N9231, N9219, N1504, N1160);
nand NAND3 (N9232, N9229, N884, N5914);
nand NAND4 (N9233, N9231, N8107, N4127, N8104);
nor NOR2 (N9234, N9233, N8350);
nor NOR2 (N9235, N9234, N2172);
buf BUF1 (N9236, N9224);
or OR4 (N9237, N9236, N7859, N7996, N6240);
buf BUF1 (N9238, N9199);
nor NOR4 (N9239, N9200, N6098, N6231, N5495);
xor XOR2 (N9240, N9232, N8819);
xor XOR2 (N9241, N9210, N5078);
and AND4 (N9242, N9235, N3314, N4661, N4595);
nand NAND3 (N9243, N9241, N2263, N1679);
buf BUF1 (N9244, N9230);
or OR3 (N9245, N9222, N6392, N8280);
and AND4 (N9246, N9243, N7346, N2085, N2696);
or OR2 (N9247, N9246, N3167);
or OR4 (N9248, N9228, N436, N4375, N3230);
nor NOR4 (N9249, N9226, N623, N7665, N5073);
and AND4 (N9250, N9244, N679, N6338, N1171);
nand NAND2 (N9251, N9250, N6359);
not NOT1 (N9252, N9242);
and AND4 (N9253, N9239, N8790, N7681, N1148);
xor XOR2 (N9254, N9252, N431);
and AND2 (N9255, N9238, N5514);
and AND2 (N9256, N9253, N3599);
xor XOR2 (N9257, N9248, N1153);
nand NAND2 (N9258, N9256, N6979);
or OR2 (N9259, N9258, N1037);
and AND3 (N9260, N9249, N7561, N7199);
or OR4 (N9261, N9240, N196, N4417, N8398);
xor XOR2 (N9262, N9259, N7923);
nand NAND3 (N9263, N9257, N5965, N1665);
and AND3 (N9264, N9261, N8447, N3773);
and AND2 (N9265, N9262, N4394);
and AND3 (N9266, N9245, N2033, N1074);
buf BUF1 (N9267, N9255);
and AND2 (N9268, N9267, N6089);
xor XOR2 (N9269, N9266, N7286);
buf BUF1 (N9270, N9264);
xor XOR2 (N9271, N9265, N2284);
nand NAND2 (N9272, N9254, N667);
nand NAND4 (N9273, N9272, N5064, N3025, N8222);
and AND4 (N9274, N9247, N3110, N6679, N6020);
and AND4 (N9275, N9268, N7622, N7511, N5536);
xor XOR2 (N9276, N9251, N4964);
xor XOR2 (N9277, N9270, N4762);
xor XOR2 (N9278, N9277, N5108);
and AND2 (N9279, N9263, N7067);
nand NAND3 (N9280, N9278, N1984, N5649);
and AND4 (N9281, N9279, N4233, N7137, N4124);
xor XOR2 (N9282, N9275, N3728);
or OR2 (N9283, N9276, N8978);
or OR3 (N9284, N9281, N7081, N2530);
xor XOR2 (N9285, N9274, N4977);
buf BUF1 (N9286, N9284);
nor NOR4 (N9287, N9280, N6093, N6661, N3303);
xor XOR2 (N9288, N9283, N5951);
not NOT1 (N9289, N9287);
xor XOR2 (N9290, N9285, N2933);
nand NAND4 (N9291, N9282, N197, N5827, N2262);
nand NAND2 (N9292, N9290, N3999);
buf BUF1 (N9293, N9237);
and AND2 (N9294, N9292, N5966);
buf BUF1 (N9295, N9293);
and AND4 (N9296, N9289, N4790, N681, N7367);
nor NOR2 (N9297, N9294, N2928);
or OR3 (N9298, N9288, N3064, N718);
nor NOR4 (N9299, N9271, N1123, N2021, N518);
nand NAND2 (N9300, N9298, N4434);
buf BUF1 (N9301, N9299);
nand NAND4 (N9302, N9301, N8529, N4930, N8289);
nor NOR3 (N9303, N9260, N1322, N8815);
or OR4 (N9304, N9297, N1295, N4892, N2313);
buf BUF1 (N9305, N9302);
not NOT1 (N9306, N9295);
buf BUF1 (N9307, N9273);
not NOT1 (N9308, N9304);
and AND3 (N9309, N9296, N4189, N1913);
nor NOR4 (N9310, N9291, N3305, N2257, N6232);
not NOT1 (N9311, N9305);
nor NOR2 (N9312, N9308, N5902);
buf BUF1 (N9313, N9306);
buf BUF1 (N9314, N9309);
buf BUF1 (N9315, N9300);
buf BUF1 (N9316, N9312);
xor XOR2 (N9317, N9303, N3583);
not NOT1 (N9318, N9315);
or OR2 (N9319, N9286, N889);
and AND3 (N9320, N9310, N1120, N102);
or OR2 (N9321, N9319, N7206);
nand NAND4 (N9322, N9311, N5455, N5482, N3780);
nand NAND2 (N9323, N9316, N2189);
and AND3 (N9324, N9323, N2010, N7355);
xor XOR2 (N9325, N9321, N7205);
xor XOR2 (N9326, N9269, N34);
nand NAND3 (N9327, N9313, N6961, N2445);
xor XOR2 (N9328, N9318, N4663);
and AND4 (N9329, N9320, N3886, N6713, N2156);
or OR3 (N9330, N9328, N7310, N7543);
or OR3 (N9331, N9317, N8240, N7673);
not NOT1 (N9332, N9331);
buf BUF1 (N9333, N9314);
buf BUF1 (N9334, N9332);
nand NAND4 (N9335, N9333, N4904, N1146, N2899);
xor XOR2 (N9336, N9330, N8565);
nor NOR2 (N9337, N9334, N1172);
and AND3 (N9338, N9337, N279, N5611);
not NOT1 (N9339, N9338);
buf BUF1 (N9340, N9326);
xor XOR2 (N9341, N9339, N720);
and AND2 (N9342, N9327, N6615);
or OR2 (N9343, N9341, N220);
xor XOR2 (N9344, N9325, N4278);
and AND2 (N9345, N9342, N6204);
nand NAND2 (N9346, N9340, N6571);
buf BUF1 (N9347, N9343);
not NOT1 (N9348, N9324);
nor NOR3 (N9349, N9345, N4633, N4354);
not NOT1 (N9350, N9347);
or OR2 (N9351, N9346, N3903);
nor NOR2 (N9352, N9322, N3034);
xor XOR2 (N9353, N9335, N3179);
nor NOR3 (N9354, N9350, N8058, N3795);
or OR2 (N9355, N9352, N8771);
buf BUF1 (N9356, N9307);
not NOT1 (N9357, N9344);
buf BUF1 (N9358, N9353);
not NOT1 (N9359, N9358);
buf BUF1 (N9360, N9348);
not NOT1 (N9361, N9336);
buf BUF1 (N9362, N9351);
xor XOR2 (N9363, N9362, N528);
or OR2 (N9364, N9363, N5233);
or OR2 (N9365, N9359, N7103);
buf BUF1 (N9366, N9355);
or OR4 (N9367, N9329, N766, N4348, N1919);
nand NAND4 (N9368, N9365, N8363, N5886, N1908);
nor NOR2 (N9369, N9356, N1483);
and AND2 (N9370, N9369, N1184);
xor XOR2 (N9371, N9370, N3168);
and AND4 (N9372, N9371, N6389, N3521, N2327);
nand NAND2 (N9373, N9360, N2181);
nor NOR4 (N9374, N9349, N315, N9336, N7658);
buf BUF1 (N9375, N9366);
xor XOR2 (N9376, N9375, N6444);
not NOT1 (N9377, N9357);
buf BUF1 (N9378, N9377);
and AND2 (N9379, N9376, N5465);
and AND3 (N9380, N9367, N8041, N5125);
nor NOR2 (N9381, N9373, N4931);
not NOT1 (N9382, N9380);
buf BUF1 (N9383, N9368);
buf BUF1 (N9384, N9379);
or OR4 (N9385, N9381, N1567, N1664, N7771);
nand NAND3 (N9386, N9378, N6747, N8186);
xor XOR2 (N9387, N9386, N6746);
not NOT1 (N9388, N9374);
nand NAND3 (N9389, N9364, N5516, N4087);
nand NAND3 (N9390, N9387, N8298, N8828);
nor NOR3 (N9391, N9372, N3223, N6225);
nor NOR3 (N9392, N9383, N5911, N4998);
not NOT1 (N9393, N9384);
nor NOR3 (N9394, N9385, N6718, N8862);
xor XOR2 (N9395, N9388, N9001);
nand NAND3 (N9396, N9382, N5254, N1387);
nor NOR3 (N9397, N9395, N6079, N6024);
nor NOR3 (N9398, N9393, N7588, N1231);
nor NOR3 (N9399, N9397, N4230, N4416);
nand NAND2 (N9400, N9394, N53);
and AND4 (N9401, N9392, N2774, N1427, N2003);
and AND4 (N9402, N9399, N4397, N1539, N2866);
nand NAND2 (N9403, N9402, N1181);
or OR2 (N9404, N9354, N6622);
not NOT1 (N9405, N9361);
not NOT1 (N9406, N9396);
xor XOR2 (N9407, N9391, N7108);
nor NOR2 (N9408, N9389, N6434);
not NOT1 (N9409, N9407);
xor XOR2 (N9410, N9408, N3464);
or OR3 (N9411, N9409, N9253, N176);
or OR2 (N9412, N9403, N4120);
not NOT1 (N9413, N9412);
nor NOR2 (N9414, N9398, N7336);
or OR3 (N9415, N9400, N8895, N2242);
not NOT1 (N9416, N9401);
nand NAND2 (N9417, N9406, N4934);
nor NOR2 (N9418, N9417, N4017);
buf BUF1 (N9419, N9416);
not NOT1 (N9420, N9414);
nor NOR2 (N9421, N9419, N6264);
and AND4 (N9422, N9410, N2028, N4321, N3877);
or OR4 (N9423, N9415, N6586, N786, N8462);
xor XOR2 (N9424, N9422, N7587);
nand NAND3 (N9425, N9421, N7395, N1411);
and AND2 (N9426, N9413, N4012);
not NOT1 (N9427, N9418);
buf BUF1 (N9428, N9404);
not NOT1 (N9429, N9405);
buf BUF1 (N9430, N9426);
buf BUF1 (N9431, N9429);
nand NAND4 (N9432, N9425, N3013, N6414, N3626);
not NOT1 (N9433, N9420);
xor XOR2 (N9434, N9430, N3703);
nor NOR2 (N9435, N9390, N1930);
buf BUF1 (N9436, N9432);
not NOT1 (N9437, N9424);
buf BUF1 (N9438, N9411);
or OR2 (N9439, N9437, N6869);
nor NOR4 (N9440, N9433, N2202, N28, N2739);
or OR4 (N9441, N9431, N3690, N336, N3871);
or OR4 (N9442, N9434, N4989, N6726, N2069);
or OR2 (N9443, N9428, N9415);
buf BUF1 (N9444, N9438);
nand NAND2 (N9445, N9436, N2295);
not NOT1 (N9446, N9445);
or OR4 (N9447, N9440, N5303, N3503, N9055);
and AND3 (N9448, N9444, N861, N1172);
xor XOR2 (N9449, N9443, N699);
and AND2 (N9450, N9441, N7829);
nand NAND3 (N9451, N9427, N754, N2708);
or OR3 (N9452, N9449, N8632, N4189);
or OR2 (N9453, N9442, N3296);
and AND3 (N9454, N9435, N7412, N5296);
or OR4 (N9455, N9454, N3615, N2123, N7988);
not NOT1 (N9456, N9453);
xor XOR2 (N9457, N9423, N7621);
or OR3 (N9458, N9446, N4260, N6278);
xor XOR2 (N9459, N9456, N390);
nor NOR2 (N9460, N9457, N4850);
and AND4 (N9461, N9439, N1692, N167, N7912);
nor NOR2 (N9462, N9452, N7220);
and AND3 (N9463, N9460, N7040, N434);
buf BUF1 (N9464, N9448);
not NOT1 (N9465, N9459);
nor NOR2 (N9466, N9458, N2235);
nand NAND2 (N9467, N9466, N8415);
not NOT1 (N9468, N9464);
buf BUF1 (N9469, N9465);
buf BUF1 (N9470, N9450);
or OR3 (N9471, N9447, N3028, N2123);
xor XOR2 (N9472, N9470, N4102);
nand NAND2 (N9473, N9455, N8491);
not NOT1 (N9474, N9471);
or OR3 (N9475, N9461, N7255, N6607);
not NOT1 (N9476, N9462);
or OR2 (N9477, N9475, N2578);
nor NOR3 (N9478, N9474, N858, N1476);
nand NAND4 (N9479, N9473, N3678, N582, N5708);
and AND2 (N9480, N9468, N8794);
or OR4 (N9481, N9472, N7628, N3583, N3493);
and AND2 (N9482, N9469, N5212);
not NOT1 (N9483, N9477);
not NOT1 (N9484, N9481);
or OR2 (N9485, N9478, N6097);
nor NOR4 (N9486, N9483, N1686, N2742, N3883);
not NOT1 (N9487, N9479);
nand NAND3 (N9488, N9485, N3464, N2151);
or OR2 (N9489, N9482, N5660);
nor NOR2 (N9490, N9488, N5095);
and AND2 (N9491, N9490, N6952);
buf BUF1 (N9492, N9486);
or OR4 (N9493, N9492, N6423, N3865, N2461);
nor NOR3 (N9494, N9487, N1756, N6290);
and AND2 (N9495, N9467, N7820);
and AND4 (N9496, N9451, N4048, N846, N5455);
buf BUF1 (N9497, N9496);
nor NOR2 (N9498, N9463, N6719);
or OR3 (N9499, N9489, N3523, N4618);
nor NOR2 (N9500, N9493, N3276);
nor NOR2 (N9501, N9494, N3499);
xor XOR2 (N9502, N9476, N3441);
xor XOR2 (N9503, N9497, N9076);
nor NOR3 (N9504, N9499, N5104, N8019);
nand NAND4 (N9505, N9500, N698, N5930, N4057);
and AND2 (N9506, N9498, N6260);
nand NAND2 (N9507, N9495, N1470);
nand NAND2 (N9508, N9505, N4076);
and AND4 (N9509, N9501, N2356, N3202, N936);
xor XOR2 (N9510, N9509, N5019);
xor XOR2 (N9511, N9510, N5657);
and AND2 (N9512, N9491, N289);
nor NOR3 (N9513, N9484, N957, N8587);
nand NAND3 (N9514, N9503, N4227, N4132);
xor XOR2 (N9515, N9512, N9019);
buf BUF1 (N9516, N9506);
and AND2 (N9517, N9508, N7962);
xor XOR2 (N9518, N9511, N1144);
buf BUF1 (N9519, N9502);
xor XOR2 (N9520, N9513, N3040);
nand NAND3 (N9521, N9517, N6228, N4707);
and AND2 (N9522, N9514, N1496);
nand NAND4 (N9523, N9520, N1070, N705, N5331);
buf BUF1 (N9524, N9523);
nand NAND4 (N9525, N9518, N6556, N1715, N5324);
and AND2 (N9526, N9516, N2315);
or OR3 (N9527, N9522, N9257, N6496);
nand NAND4 (N9528, N9519, N6301, N2994, N2033);
not NOT1 (N9529, N9526);
or OR4 (N9530, N9480, N3533, N8324, N913);
and AND3 (N9531, N9515, N5027, N2196);
buf BUF1 (N9532, N9531);
not NOT1 (N9533, N9525);
nand NAND2 (N9534, N9529, N4316);
nand NAND4 (N9535, N9524, N910, N451, N56);
nor NOR3 (N9536, N9530, N5872, N5397);
nand NAND2 (N9537, N9507, N9011);
or OR2 (N9538, N9528, N3996);
buf BUF1 (N9539, N9536);
buf BUF1 (N9540, N9537);
or OR4 (N9541, N9521, N2801, N6248, N4863);
buf BUF1 (N9542, N9532);
or OR2 (N9543, N9527, N3025);
xor XOR2 (N9544, N9540, N910);
or OR2 (N9545, N9538, N6291);
and AND3 (N9546, N9534, N1621, N110);
nor NOR2 (N9547, N9504, N6798);
and AND3 (N9548, N9539, N1292, N5197);
or OR2 (N9549, N9544, N5592);
nor NOR2 (N9550, N9549, N203);
nand NAND4 (N9551, N9546, N712, N2928, N4569);
nand NAND4 (N9552, N9547, N4114, N655, N5129);
nor NOR2 (N9553, N9548, N3797);
nor NOR3 (N9554, N9552, N8391, N2878);
buf BUF1 (N9555, N9543);
xor XOR2 (N9556, N9555, N4052);
xor XOR2 (N9557, N9550, N5005);
buf BUF1 (N9558, N9556);
nor NOR2 (N9559, N9545, N5638);
xor XOR2 (N9560, N9558, N6659);
nor NOR3 (N9561, N9559, N1324, N226);
or OR3 (N9562, N9560, N4179, N6923);
or OR3 (N9563, N9533, N9228, N3746);
buf BUF1 (N9564, N9535);
not NOT1 (N9565, N9551);
buf BUF1 (N9566, N9542);
nand NAND3 (N9567, N9563, N7153, N5039);
buf BUF1 (N9568, N9565);
and AND4 (N9569, N9562, N4614, N6348, N7725);
and AND2 (N9570, N9554, N8473);
buf BUF1 (N9571, N9568);
nand NAND4 (N9572, N9567, N896, N1273, N8798);
or OR2 (N9573, N9561, N3767);
and AND2 (N9574, N9572, N8131);
nand NAND3 (N9575, N9566, N8687, N2096);
and AND2 (N9576, N9564, N3045);
xor XOR2 (N9577, N9575, N7573);
xor XOR2 (N9578, N9553, N1971);
or OR3 (N9579, N9578, N3151, N5005);
and AND3 (N9580, N9569, N8046, N5874);
not NOT1 (N9581, N9580);
or OR4 (N9582, N9577, N4216, N3141, N3006);
or OR2 (N9583, N9570, N5227);
xor XOR2 (N9584, N9574, N1877);
nand NAND4 (N9585, N9579, N446, N8373, N3605);
not NOT1 (N9586, N9584);
buf BUF1 (N9587, N9541);
xor XOR2 (N9588, N9585, N9030);
nand NAND3 (N9589, N9571, N7734, N3044);
and AND2 (N9590, N9586, N5103);
and AND2 (N9591, N9590, N9143);
buf BUF1 (N9592, N9581);
or OR3 (N9593, N9587, N4331, N4539);
and AND2 (N9594, N9588, N4961);
nand NAND4 (N9595, N9592, N9432, N9163, N5558);
nor NOR3 (N9596, N9594, N3176, N1599);
not NOT1 (N9597, N9576);
nor NOR2 (N9598, N9591, N6338);
buf BUF1 (N9599, N9597);
and AND3 (N9600, N9596, N8440, N8316);
nor NOR2 (N9601, N9589, N5864);
nor NOR3 (N9602, N9573, N1506, N2725);
nand NAND2 (N9603, N9601, N751);
or OR3 (N9604, N9595, N5614, N205);
buf BUF1 (N9605, N9583);
and AND2 (N9606, N9602, N2180);
or OR3 (N9607, N9598, N1031, N3604);
or OR3 (N9608, N9582, N9228, N8092);
not NOT1 (N9609, N9600);
nand NAND3 (N9610, N9605, N6766, N232);
nor NOR4 (N9611, N9610, N1440, N7631, N2640);
or OR3 (N9612, N9603, N2322, N6900);
xor XOR2 (N9613, N9604, N6340);
xor XOR2 (N9614, N9613, N235);
nand NAND3 (N9615, N9607, N4384, N4083);
or OR2 (N9616, N9615, N6641);
nand NAND2 (N9617, N9616, N6982);
nor NOR2 (N9618, N9609, N9429);
not NOT1 (N9619, N9617);
nand NAND2 (N9620, N9619, N8331);
buf BUF1 (N9621, N9606);
xor XOR2 (N9622, N9611, N857);
not NOT1 (N9623, N9612);
or OR2 (N9624, N9608, N5318);
nor NOR2 (N9625, N9624, N4651);
buf BUF1 (N9626, N9593);
nand NAND3 (N9627, N9625, N4893, N4535);
nand NAND3 (N9628, N9557, N7099, N8655);
nor NOR2 (N9629, N9618, N8275);
or OR4 (N9630, N9614, N3967, N1016, N6871);
or OR2 (N9631, N9629, N7264);
buf BUF1 (N9632, N9621);
not NOT1 (N9633, N9626);
not NOT1 (N9634, N9630);
xor XOR2 (N9635, N9620, N961);
or OR4 (N9636, N9635, N5279, N8642, N7378);
not NOT1 (N9637, N9634);
nor NOR3 (N9638, N9628, N7232, N6584);
nand NAND4 (N9639, N9623, N5439, N1328, N2125);
not NOT1 (N9640, N9637);
xor XOR2 (N9641, N9627, N5954);
not NOT1 (N9642, N9631);
not NOT1 (N9643, N9632);
nand NAND4 (N9644, N9599, N759, N6325, N8127);
or OR2 (N9645, N9643, N3367);
buf BUF1 (N9646, N9642);
not NOT1 (N9647, N9641);
and AND3 (N9648, N9636, N3609, N4246);
nor NOR2 (N9649, N9647, N143);
xor XOR2 (N9650, N9639, N830);
nand NAND4 (N9651, N9640, N1735, N9431, N3944);
or OR3 (N9652, N9650, N2267, N6721);
and AND3 (N9653, N9645, N4895, N2363);
or OR2 (N9654, N9653, N7699);
nor NOR4 (N9655, N9638, N4732, N1589, N4847);
nor NOR2 (N9656, N9654, N4872);
not NOT1 (N9657, N9646);
or OR3 (N9658, N9648, N8707, N2389);
xor XOR2 (N9659, N9655, N894);
not NOT1 (N9660, N9649);
nand NAND4 (N9661, N9644, N5113, N5733, N4126);
not NOT1 (N9662, N9658);
nand NAND4 (N9663, N9652, N8194, N4213, N5547);
and AND3 (N9664, N9657, N5445, N2321);
not NOT1 (N9665, N9661);
nor NOR3 (N9666, N9665, N2038, N8815);
buf BUF1 (N9667, N9663);
or OR3 (N9668, N9664, N4982, N2392);
and AND3 (N9669, N9659, N9628, N2679);
xor XOR2 (N9670, N9662, N2894);
buf BUF1 (N9671, N9668);
not NOT1 (N9672, N9651);
or OR3 (N9673, N9672, N1101, N9027);
nor NOR2 (N9674, N9667, N813);
nor NOR4 (N9675, N9622, N8431, N3424, N7660);
xor XOR2 (N9676, N9660, N3886);
nand NAND2 (N9677, N9676, N4321);
buf BUF1 (N9678, N9673);
or OR3 (N9679, N9678, N2764, N3080);
and AND3 (N9680, N9670, N1705, N7609);
nand NAND4 (N9681, N9666, N4827, N6251, N6927);
nor NOR4 (N9682, N9679, N7220, N444, N5600);
or OR3 (N9683, N9677, N74, N6491);
nand NAND4 (N9684, N9671, N4154, N6845, N6718);
nor NOR3 (N9685, N9674, N5169, N8055);
nor NOR4 (N9686, N9684, N4985, N4709, N774);
nor NOR2 (N9687, N9633, N1597);
or OR4 (N9688, N9685, N3945, N818, N6911);
nand NAND4 (N9689, N9681, N1965, N715, N3904);
not NOT1 (N9690, N9680);
not NOT1 (N9691, N9675);
xor XOR2 (N9692, N9687, N936);
or OR2 (N9693, N9691, N7150);
or OR3 (N9694, N9669, N1296, N154);
and AND3 (N9695, N9693, N8203, N7908);
nor NOR4 (N9696, N9689, N5277, N5931, N6980);
nor NOR4 (N9697, N9694, N9601, N1542, N9516);
nor NOR4 (N9698, N9690, N6171, N6707, N6803);
xor XOR2 (N9699, N9686, N8713);
or OR3 (N9700, N9698, N2619, N7564);
not NOT1 (N9701, N9699);
or OR3 (N9702, N9683, N4653, N7665);
buf BUF1 (N9703, N9696);
nand NAND3 (N9704, N9702, N2608, N6049);
nand NAND4 (N9705, N9703, N1460, N7909, N2799);
nand NAND2 (N9706, N9688, N5636);
and AND4 (N9707, N9682, N943, N6173, N8137);
not NOT1 (N9708, N9707);
xor XOR2 (N9709, N9700, N5727);
nand NAND2 (N9710, N9704, N6838);
nor NOR4 (N9711, N9695, N9476, N6722, N4305);
and AND2 (N9712, N9701, N1217);
and AND2 (N9713, N9705, N5447);
nor NOR4 (N9714, N9708, N6617, N9546, N4694);
and AND3 (N9715, N9714, N162, N4914);
nor NOR4 (N9716, N9715, N7596, N7185, N8776);
buf BUF1 (N9717, N9710);
buf BUF1 (N9718, N9706);
not NOT1 (N9719, N9656);
not NOT1 (N9720, N9697);
and AND3 (N9721, N9713, N3853, N9049);
xor XOR2 (N9722, N9720, N4051);
xor XOR2 (N9723, N9719, N456);
not NOT1 (N9724, N9692);
nor NOR2 (N9725, N9721, N2704);
nor NOR3 (N9726, N9725, N191, N7340);
buf BUF1 (N9727, N9716);
not NOT1 (N9728, N9718);
not NOT1 (N9729, N9722);
or OR4 (N9730, N9711, N2599, N2200, N3493);
nor NOR4 (N9731, N9709, N2059, N3260, N2264);
buf BUF1 (N9732, N9727);
and AND3 (N9733, N9730, N5728, N9265);
nand NAND3 (N9734, N9732, N4000, N5832);
and AND3 (N9735, N9712, N7942, N9145);
xor XOR2 (N9736, N9726, N2366);
and AND3 (N9737, N9728, N5517, N4844);
xor XOR2 (N9738, N9737, N1842);
xor XOR2 (N9739, N9738, N9535);
nor NOR3 (N9740, N9735, N3109, N7873);
or OR2 (N9741, N9736, N6161);
nor NOR4 (N9742, N9733, N167, N6236, N5751);
xor XOR2 (N9743, N9740, N4377);
buf BUF1 (N9744, N9741);
not NOT1 (N9745, N9739);
and AND2 (N9746, N9743, N3597);
or OR4 (N9747, N9723, N699, N8189, N1523);
or OR3 (N9748, N9717, N5584, N4870);
buf BUF1 (N9749, N9724);
not NOT1 (N9750, N9731);
buf BUF1 (N9751, N9750);
nor NOR4 (N9752, N9751, N4707, N748, N4115);
not NOT1 (N9753, N9748);
nand NAND4 (N9754, N9747, N5719, N7139, N3414);
buf BUF1 (N9755, N9742);
xor XOR2 (N9756, N9752, N490);
buf BUF1 (N9757, N9746);
nor NOR4 (N9758, N9749, N3165, N8239, N2248);
buf BUF1 (N9759, N9753);
or OR3 (N9760, N9755, N3707, N4325);
not NOT1 (N9761, N9744);
and AND4 (N9762, N9729, N3405, N8071, N900);
xor XOR2 (N9763, N9757, N5117);
nand NAND3 (N9764, N9745, N8225, N1884);
buf BUF1 (N9765, N9762);
and AND4 (N9766, N9758, N2854, N2454, N6587);
or OR4 (N9767, N9766, N4928, N1976, N9675);
or OR3 (N9768, N9761, N9101, N8717);
nand NAND2 (N9769, N9734, N5019);
not NOT1 (N9770, N9767);
nand NAND3 (N9771, N9759, N2745, N8631);
nand NAND2 (N9772, N9754, N7218);
nor NOR3 (N9773, N9770, N3333, N8698);
nand NAND4 (N9774, N9756, N2672, N2797, N5550);
nand NAND2 (N9775, N9765, N3631);
not NOT1 (N9776, N9775);
or OR4 (N9777, N9776, N5616, N5043, N7144);
xor XOR2 (N9778, N9777, N4864);
xor XOR2 (N9779, N9760, N2860);
nand NAND3 (N9780, N9779, N8426, N199);
nand NAND2 (N9781, N9763, N8988);
nand NAND2 (N9782, N9774, N1534);
nand NAND3 (N9783, N9782, N6420, N6875);
buf BUF1 (N9784, N9771);
or OR2 (N9785, N9781, N6701);
buf BUF1 (N9786, N9772);
xor XOR2 (N9787, N9783, N4763);
buf BUF1 (N9788, N9784);
buf BUF1 (N9789, N9773);
nor NOR3 (N9790, N9764, N1850, N7960);
and AND2 (N9791, N9787, N3465);
or OR2 (N9792, N9768, N7357);
nor NOR4 (N9793, N9790, N700, N6776, N2199);
xor XOR2 (N9794, N9769, N8042);
nor NOR2 (N9795, N9791, N2129);
and AND4 (N9796, N9786, N3117, N5069, N5004);
or OR2 (N9797, N9792, N7273);
nand NAND4 (N9798, N9788, N8444, N3526, N4686);
not NOT1 (N9799, N9798);
buf BUF1 (N9800, N9794);
xor XOR2 (N9801, N9793, N5187);
and AND3 (N9802, N9789, N8410, N9283);
not NOT1 (N9803, N9796);
buf BUF1 (N9804, N9778);
or OR2 (N9805, N9785, N1948);
xor XOR2 (N9806, N9803, N3165);
not NOT1 (N9807, N9795);
nor NOR2 (N9808, N9804, N8215);
not NOT1 (N9809, N9800);
nor NOR3 (N9810, N9799, N761, N5424);
xor XOR2 (N9811, N9809, N4904);
nor NOR3 (N9812, N9780, N668, N3364);
and AND4 (N9813, N9801, N2947, N5941, N7995);
not NOT1 (N9814, N9805);
or OR2 (N9815, N9811, N9005);
nand NAND3 (N9816, N9807, N2745, N9418);
not NOT1 (N9817, N9797);
not NOT1 (N9818, N9810);
and AND4 (N9819, N9808, N9144, N6028, N6913);
and AND3 (N9820, N9816, N9539, N7423);
xor XOR2 (N9821, N9802, N6154);
or OR2 (N9822, N9814, N1938);
xor XOR2 (N9823, N9813, N9542);
buf BUF1 (N9824, N9823);
and AND2 (N9825, N9818, N8987);
xor XOR2 (N9826, N9817, N2387);
or OR2 (N9827, N9820, N3787);
nand NAND3 (N9828, N9826, N1385, N4135);
xor XOR2 (N9829, N9819, N7183);
xor XOR2 (N9830, N9827, N2478);
and AND3 (N9831, N9821, N2054, N8661);
nand NAND2 (N9832, N9831, N6324);
buf BUF1 (N9833, N9815);
and AND4 (N9834, N9830, N6326, N4251, N6154);
and AND4 (N9835, N9806, N3893, N9561, N2677);
xor XOR2 (N9836, N9834, N7756);
xor XOR2 (N9837, N9833, N5058);
or OR3 (N9838, N9825, N8690, N2806);
or OR3 (N9839, N9835, N4892, N9337);
nand NAND2 (N9840, N9837, N413);
not NOT1 (N9841, N9832);
and AND4 (N9842, N9829, N6276, N3792, N233);
or OR2 (N9843, N9839, N5169);
and AND4 (N9844, N9824, N3173, N4229, N9837);
not NOT1 (N9845, N9836);
or OR3 (N9846, N9842, N2494, N648);
or OR4 (N9847, N9843, N4000, N1614, N6051);
buf BUF1 (N9848, N9840);
nor NOR4 (N9849, N9846, N8293, N7277, N7240);
xor XOR2 (N9850, N9847, N7305);
nand NAND2 (N9851, N9844, N1855);
not NOT1 (N9852, N9841);
buf BUF1 (N9853, N9845);
and AND2 (N9854, N9812, N6220);
nand NAND3 (N9855, N9852, N3557, N2197);
buf BUF1 (N9856, N9850);
buf BUF1 (N9857, N9851);
nand NAND4 (N9858, N9838, N889, N4940, N5728);
nand NAND3 (N9859, N9848, N1824, N2468);
not NOT1 (N9860, N9853);
xor XOR2 (N9861, N9858, N1034);
nor NOR4 (N9862, N9861, N8329, N4474, N5290);
xor XOR2 (N9863, N9854, N5311);
buf BUF1 (N9864, N9849);
nand NAND2 (N9865, N9860, N724);
and AND2 (N9866, N9863, N7289);
or OR4 (N9867, N9859, N6312, N8354, N5771);
nor NOR2 (N9868, N9866, N4448);
and AND2 (N9869, N9867, N2761);
and AND3 (N9870, N9869, N2392, N5862);
xor XOR2 (N9871, N9857, N4930);
buf BUF1 (N9872, N9870);
and AND2 (N9873, N9865, N8923);
buf BUF1 (N9874, N9828);
not NOT1 (N9875, N9864);
not NOT1 (N9876, N9871);
xor XOR2 (N9877, N9874, N9525);
xor XOR2 (N9878, N9856, N4359);
not NOT1 (N9879, N9862);
xor XOR2 (N9880, N9822, N9728);
not NOT1 (N9881, N9873);
buf BUF1 (N9882, N9881);
xor XOR2 (N9883, N9880, N6023);
or OR3 (N9884, N9868, N1014, N6472);
buf BUF1 (N9885, N9878);
xor XOR2 (N9886, N9875, N2730);
xor XOR2 (N9887, N9879, N7525);
xor XOR2 (N9888, N9882, N1071);
xor XOR2 (N9889, N9888, N3179);
and AND2 (N9890, N9855, N1162);
nand NAND3 (N9891, N9872, N5548, N4959);
and AND3 (N9892, N9883, N5638, N1283);
or OR4 (N9893, N9885, N373, N8716, N7657);
nand NAND3 (N9894, N9877, N7353, N6326);
xor XOR2 (N9895, N9876, N2895);
xor XOR2 (N9896, N9889, N5797);
or OR2 (N9897, N9893, N6902);
xor XOR2 (N9898, N9890, N4256);
and AND3 (N9899, N9884, N3526, N4220);
nand NAND4 (N9900, N9894, N1591, N6335, N4779);
and AND4 (N9901, N9898, N1575, N8716, N5752);
nor NOR4 (N9902, N9896, N5472, N1601, N6293);
nor NOR2 (N9903, N9900, N667);
not NOT1 (N9904, N9887);
or OR3 (N9905, N9891, N2389, N9332);
nand NAND4 (N9906, N9886, N2007, N507, N8075);
or OR2 (N9907, N9897, N7268);
or OR4 (N9908, N9892, N4673, N6686, N5771);
nand NAND4 (N9909, N9908, N6846, N9413, N995);
and AND3 (N9910, N9895, N848, N7743);
xor XOR2 (N9911, N9906, N6196);
buf BUF1 (N9912, N9904);
nor NOR2 (N9913, N9903, N6310);
and AND4 (N9914, N9899, N2667, N3759, N3694);
nand NAND4 (N9915, N9912, N5989, N4445, N6722);
not NOT1 (N9916, N9907);
xor XOR2 (N9917, N9916, N5765);
and AND3 (N9918, N9901, N1689, N5600);
nand NAND4 (N9919, N9905, N2197, N3569, N2649);
or OR2 (N9920, N9914, N1506);
buf BUF1 (N9921, N9902);
buf BUF1 (N9922, N9910);
and AND4 (N9923, N9919, N2438, N7215, N968);
xor XOR2 (N9924, N9913, N6415);
or OR3 (N9925, N9924, N4262, N6030);
not NOT1 (N9926, N9917);
buf BUF1 (N9927, N9920);
nand NAND2 (N9928, N9918, N218);
nand NAND2 (N9929, N9925, N2980);
or OR3 (N9930, N9915, N5251, N4804);
or OR2 (N9931, N9922, N1380);
xor XOR2 (N9932, N9931, N8358);
not NOT1 (N9933, N9927);
and AND3 (N9934, N9928, N2418, N560);
and AND4 (N9935, N9929, N2195, N2865, N259);
or OR4 (N9936, N9926, N627, N6016, N8985);
nand NAND3 (N9937, N9936, N5887, N5364);
not NOT1 (N9938, N9935);
buf BUF1 (N9939, N9911);
or OR2 (N9940, N9933, N6528);
buf BUF1 (N9941, N9940);
and AND2 (N9942, N9909, N3398);
buf BUF1 (N9943, N9942);
nand NAND2 (N9944, N9923, N7436);
or OR3 (N9945, N9932, N2869, N6526);
nor NOR4 (N9946, N9945, N6863, N2952, N6441);
buf BUF1 (N9947, N9944);
or OR4 (N9948, N9930, N9740, N1650, N4292);
buf BUF1 (N9949, N9948);
nor NOR4 (N9950, N9939, N989, N834, N7152);
nand NAND3 (N9951, N9938, N3585, N6058);
nor NOR4 (N9952, N9950, N7545, N7114, N7631);
or OR3 (N9953, N9949, N1733, N9176);
buf BUF1 (N9954, N9937);
and AND2 (N9955, N9934, N6725);
buf BUF1 (N9956, N9943);
and AND3 (N9957, N9941, N6250, N7987);
nand NAND2 (N9958, N9953, N5640);
buf BUF1 (N9959, N9955);
xor XOR2 (N9960, N9946, N8974);
buf BUF1 (N9961, N9957);
or OR4 (N9962, N9960, N8086, N2551, N9430);
not NOT1 (N9963, N9959);
not NOT1 (N9964, N9958);
not NOT1 (N9965, N9952);
and AND3 (N9966, N9965, N928, N3228);
buf BUF1 (N9967, N9956);
not NOT1 (N9968, N9967);
nor NOR3 (N9969, N9961, N3497, N4757);
xor XOR2 (N9970, N9963, N4668);
and AND3 (N9971, N9947, N6950, N123);
buf BUF1 (N9972, N9971);
or OR2 (N9973, N9969, N1596);
not NOT1 (N9974, N9921);
nand NAND3 (N9975, N9972, N9275, N1291);
nand NAND2 (N9976, N9968, N2623);
buf BUF1 (N9977, N9970);
and AND2 (N9978, N9974, N8005);
not NOT1 (N9979, N9975);
and AND3 (N9980, N9962, N8259, N8760);
xor XOR2 (N9981, N9966, N5193);
nor NOR3 (N9982, N9976, N6289, N4612);
xor XOR2 (N9983, N9982, N278);
and AND4 (N9984, N9954, N9028, N4044, N4027);
and AND3 (N9985, N9979, N355, N1054);
xor XOR2 (N9986, N9978, N4409);
or OR3 (N9987, N9951, N6897, N2998);
and AND4 (N9988, N9977, N612, N7107, N4033);
xor XOR2 (N9989, N9983, N5004);
not NOT1 (N9990, N9987);
nand NAND2 (N9991, N9989, N7069);
or OR4 (N9992, N9973, N5376, N6573, N1316);
nand NAND2 (N9993, N9984, N7152);
and AND3 (N9994, N9993, N6609, N8051);
nand NAND2 (N9995, N9992, N9267);
buf BUF1 (N9996, N9994);
nand NAND2 (N9997, N9991, N9587);
buf BUF1 (N9998, N9997);
buf BUF1 (N9999, N9964);
nand NAND4 (N10000, N9998, N8740, N1336, N1885);
not NOT1 (N10001, N9996);
xor XOR2 (N10002, N9986, N1664);
or OR4 (N10003, N9981, N7546, N9913, N5050);
xor XOR2 (N10004, N9990, N6785);
not NOT1 (N10005, N9980);
not NOT1 (N10006, N10005);
or OR2 (N10007, N9988, N2932);
nor NOR4 (N10008, N10006, N5135, N3540, N5108);
buf BUF1 (N10009, N9995);
buf BUF1 (N10010, N10003);
or OR3 (N10011, N10004, N8481, N5880);
nor NOR3 (N10012, N10011, N3460, N1746);
buf BUF1 (N10013, N9999);
or OR4 (N10014, N10010, N6374, N4359, N9349);
or OR4 (N10015, N10001, N4529, N8682, N9798);
nor NOR4 (N10016, N10009, N2530, N1374, N3592);
buf BUF1 (N10017, N10014);
and AND4 (N10018, N10002, N5602, N6919, N1095);
buf BUF1 (N10019, N10008);
and AND4 (N10020, N10015, N3295, N7341, N994);
xor XOR2 (N10021, N10020, N9947);
and AND3 (N10022, N10000, N45, N2369);
nand NAND4 (N10023, N10018, N9089, N5653, N7905);
nand NAND4 (N10024, N10021, N4345, N1051, N5206);
and AND3 (N10025, N10024, N6438, N2825);
nand NAND4 (N10026, N10022, N1482, N1010, N2726);
nor NOR3 (N10027, N10013, N2550, N6211);
nor NOR3 (N10028, N10019, N4809, N1588);
nand NAND3 (N10029, N10028, N4495, N4452);
or OR3 (N10030, N10027, N4708, N3403);
buf BUF1 (N10031, N10016);
nand NAND4 (N10032, N10031, N9123, N6310, N6679);
buf BUF1 (N10033, N10029);
nand NAND3 (N10034, N10025, N6924, N1908);
or OR3 (N10035, N10023, N9782, N4201);
buf BUF1 (N10036, N10012);
and AND2 (N10037, N10007, N1509);
buf BUF1 (N10038, N10026);
xor XOR2 (N10039, N10035, N1370);
xor XOR2 (N10040, N10034, N1147);
and AND3 (N10041, N10033, N8942, N2856);
nand NAND2 (N10042, N10041, N2402);
nand NAND4 (N10043, N10030, N3702, N9211, N603);
xor XOR2 (N10044, N9985, N7168);
or OR4 (N10045, N10039, N8445, N9960, N7547);
buf BUF1 (N10046, N10037);
not NOT1 (N10047, N10045);
or OR3 (N10048, N10017, N4004, N9615);
xor XOR2 (N10049, N10044, N1568);
nand NAND4 (N10050, N10038, N3907, N5483, N9181);
xor XOR2 (N10051, N10036, N9967);
not NOT1 (N10052, N10043);
nor NOR3 (N10053, N10042, N4740, N4922);
buf BUF1 (N10054, N10053);
nor NOR2 (N10055, N10052, N9608);
nor NOR3 (N10056, N10046, N8280, N2265);
nand NAND2 (N10057, N10056, N1065);
xor XOR2 (N10058, N10032, N2543);
and AND3 (N10059, N10054, N9871, N6242);
or OR3 (N10060, N10047, N2533, N1756);
and AND2 (N10061, N10051, N6916);
or OR4 (N10062, N10055, N2310, N6284, N8635);
and AND2 (N10063, N10058, N5124);
and AND4 (N10064, N10063, N620, N9478, N8190);
buf BUF1 (N10065, N10050);
nor NOR3 (N10066, N10049, N3319, N1251);
buf BUF1 (N10067, N10061);
nor NOR4 (N10068, N10048, N9039, N9137, N6988);
nand NAND3 (N10069, N10065, N7489, N1075);
nor NOR3 (N10070, N10060, N1114, N9026);
or OR3 (N10071, N10070, N6110, N5900);
and AND4 (N10072, N10059, N2646, N4869, N4197);
nand NAND4 (N10073, N10057, N9905, N9011, N9493);
nor NOR4 (N10074, N10040, N7000, N7167, N6157);
nor NOR4 (N10075, N10071, N5082, N9465, N317);
nand NAND3 (N10076, N10073, N6125, N8657);
buf BUF1 (N10077, N10075);
xor XOR2 (N10078, N10066, N3014);
xor XOR2 (N10079, N10078, N7919);
or OR3 (N10080, N10067, N6261, N814);
and AND3 (N10081, N10072, N7563, N9813);
buf BUF1 (N10082, N10068);
xor XOR2 (N10083, N10062, N7537);
or OR4 (N10084, N10076, N8524, N5695, N4167);
xor XOR2 (N10085, N10074, N1091);
nand NAND3 (N10086, N10077, N2345, N1106);
xor XOR2 (N10087, N10064, N7286);
nor NOR4 (N10088, N10069, N8860, N3855, N3642);
nor NOR2 (N10089, N10085, N2063);
and AND4 (N10090, N10087, N3330, N1303, N2584);
xor XOR2 (N10091, N10083, N3034);
and AND3 (N10092, N10082, N300, N3947);
and AND4 (N10093, N10084, N4174, N7291, N100);
and AND2 (N10094, N10079, N681);
xor XOR2 (N10095, N10080, N5661);
or OR2 (N10096, N10088, N3546);
nor NOR4 (N10097, N10089, N666, N3091, N7081);
not NOT1 (N10098, N10090);
buf BUF1 (N10099, N10097);
or OR4 (N10100, N10096, N3654, N4207, N5839);
nor NOR3 (N10101, N10098, N6902, N2422);
nand NAND3 (N10102, N10091, N4678, N4812);
nor NOR3 (N10103, N10092, N4749, N2972);
xor XOR2 (N10104, N10095, N4290);
and AND2 (N10105, N10100, N6204);
buf BUF1 (N10106, N10105);
nor NOR2 (N10107, N10081, N7860);
nand NAND3 (N10108, N10102, N5645, N5658);
or OR2 (N10109, N10101, N6098);
not NOT1 (N10110, N10093);
nor NOR2 (N10111, N10104, N3585);
and AND2 (N10112, N10111, N9236);
nor NOR3 (N10113, N10099, N521, N110);
xor XOR2 (N10114, N10113, N5945);
nor NOR3 (N10115, N10108, N4430, N7895);
and AND3 (N10116, N10110, N1449, N10081);
or OR3 (N10117, N10112, N8599, N5918);
not NOT1 (N10118, N10114);
and AND2 (N10119, N10116, N9373);
nand NAND2 (N10120, N10106, N7126);
and AND3 (N10121, N10107, N6265, N8668);
xor XOR2 (N10122, N10109, N8003);
and AND2 (N10123, N10103, N3961);
and AND4 (N10124, N10094, N9426, N3599, N7655);
not NOT1 (N10125, N10117);
not NOT1 (N10126, N10120);
buf BUF1 (N10127, N10124);
nor NOR2 (N10128, N10123, N136);
nor NOR3 (N10129, N10122, N1678, N560);
xor XOR2 (N10130, N10125, N7432);
nor NOR2 (N10131, N10118, N1921);
or OR3 (N10132, N10128, N1085, N672);
nand NAND2 (N10133, N10127, N7283);
or OR2 (N10134, N10086, N318);
or OR2 (N10135, N10133, N6286);
xor XOR2 (N10136, N10119, N5135);
buf BUF1 (N10137, N10115);
not NOT1 (N10138, N10121);
nand NAND4 (N10139, N10136, N290, N1109, N9832);
or OR3 (N10140, N10138, N889, N7332);
not NOT1 (N10141, N10137);
xor XOR2 (N10142, N10131, N421);
buf BUF1 (N10143, N10141);
buf BUF1 (N10144, N10134);
nand NAND2 (N10145, N10135, N2880);
not NOT1 (N10146, N10129);
or OR4 (N10147, N10142, N5446, N2013, N7164);
buf BUF1 (N10148, N10147);
xor XOR2 (N10149, N10132, N7001);
or OR2 (N10150, N10144, N4803);
nand NAND3 (N10151, N10148, N3832, N6593);
xor XOR2 (N10152, N10146, N3109);
nor NOR2 (N10153, N10150, N8649);
not NOT1 (N10154, N10145);
not NOT1 (N10155, N10130);
or OR4 (N10156, N10126, N8643, N8671, N1691);
not NOT1 (N10157, N10155);
nand NAND3 (N10158, N10143, N2515, N7663);
or OR2 (N10159, N10158, N5823);
or OR3 (N10160, N10149, N6956, N7323);
or OR3 (N10161, N10152, N7336, N566);
not NOT1 (N10162, N10139);
nor NOR3 (N10163, N10151, N1299, N2641);
not NOT1 (N10164, N10153);
nand NAND3 (N10165, N10159, N4061, N6459);
and AND2 (N10166, N10162, N2047);
not NOT1 (N10167, N10166);
or OR3 (N10168, N10167, N3996, N6927);
nand NAND4 (N10169, N10154, N2616, N1549, N9716);
buf BUF1 (N10170, N10140);
nor NOR2 (N10171, N10164, N7013);
or OR2 (N10172, N10156, N5716);
and AND4 (N10173, N10160, N9193, N7277, N9937);
and AND2 (N10174, N10157, N4247);
and AND4 (N10175, N10173, N9531, N7299, N3035);
nor NOR3 (N10176, N10165, N7571, N6698);
buf BUF1 (N10177, N10176);
or OR4 (N10178, N10177, N8739, N6420, N3099);
not NOT1 (N10179, N10178);
not NOT1 (N10180, N10170);
or OR4 (N10181, N10172, N8845, N2735, N1402);
nand NAND4 (N10182, N10180, N4235, N8380, N4419);
not NOT1 (N10183, N10171);
or OR3 (N10184, N10179, N3795, N2218);
buf BUF1 (N10185, N10169);
or OR4 (N10186, N10181, N9275, N7617, N1560);
or OR4 (N10187, N10184, N8466, N8297, N10156);
xor XOR2 (N10188, N10161, N3314);
not NOT1 (N10189, N10183);
xor XOR2 (N10190, N10189, N7422);
or OR4 (N10191, N10190, N7510, N7215, N8705);
buf BUF1 (N10192, N10175);
xor XOR2 (N10193, N10174, N4717);
and AND3 (N10194, N10191, N1286, N9523);
not NOT1 (N10195, N10185);
xor XOR2 (N10196, N10194, N10068);
not NOT1 (N10197, N10193);
xor XOR2 (N10198, N10187, N1774);
nand NAND2 (N10199, N10163, N6763);
nand NAND4 (N10200, N10195, N6474, N4745, N3874);
nor NOR4 (N10201, N10188, N7018, N5709, N8571);
and AND2 (N10202, N10196, N4254);
nand NAND4 (N10203, N10197, N6900, N7016, N1267);
not NOT1 (N10204, N10182);
xor XOR2 (N10205, N10204, N2810);
nand NAND2 (N10206, N10203, N7390);
nor NOR3 (N10207, N10205, N7515, N3378);
nor NOR3 (N10208, N10199, N3078, N454);
not NOT1 (N10209, N10201);
not NOT1 (N10210, N10206);
nor NOR3 (N10211, N10192, N3085, N4615);
buf BUF1 (N10212, N10202);
xor XOR2 (N10213, N10198, N9223);
not NOT1 (N10214, N10208);
buf BUF1 (N10215, N10210);
xor XOR2 (N10216, N10212, N2388);
xor XOR2 (N10217, N10213, N8443);
not NOT1 (N10218, N10168);
nor NOR2 (N10219, N10186, N2450);
buf BUF1 (N10220, N10207);
and AND4 (N10221, N10200, N1916, N2818, N9676);
or OR3 (N10222, N10221, N9030, N6811);
nand NAND2 (N10223, N10209, N3730);
and AND4 (N10224, N10223, N324, N8892, N5855);
or OR2 (N10225, N10219, N1907);
nor NOR3 (N10226, N10220, N9983, N2007);
and AND4 (N10227, N10225, N3274, N9288, N3559);
not NOT1 (N10228, N10217);
not NOT1 (N10229, N10214);
nor NOR3 (N10230, N10227, N1976, N6042);
buf BUF1 (N10231, N10226);
xor XOR2 (N10232, N10222, N197);
or OR4 (N10233, N10232, N7738, N173, N6041);
or OR3 (N10234, N10215, N920, N9929);
or OR2 (N10235, N10211, N2026);
or OR3 (N10236, N10234, N5577, N9411);
xor XOR2 (N10237, N10236, N4569);
buf BUF1 (N10238, N10235);
xor XOR2 (N10239, N10231, N591);
buf BUF1 (N10240, N10238);
and AND3 (N10241, N10239, N7065, N5997);
xor XOR2 (N10242, N10241, N3139);
not NOT1 (N10243, N10237);
nand NAND2 (N10244, N10233, N6524);
and AND3 (N10245, N10229, N6845, N613);
nand NAND2 (N10246, N10245, N5667);
nand NAND3 (N10247, N10218, N7063, N8016);
xor XOR2 (N10248, N10240, N906);
nand NAND2 (N10249, N10243, N6173);
or OR2 (N10250, N10246, N140);
nor NOR4 (N10251, N10224, N163, N873, N1558);
nand NAND2 (N10252, N10244, N1647);
nand NAND3 (N10253, N10248, N9668, N7060);
xor XOR2 (N10254, N10252, N1835);
xor XOR2 (N10255, N10216, N2086);
buf BUF1 (N10256, N10247);
buf BUF1 (N10257, N10253);
and AND3 (N10258, N10254, N8370, N456);
and AND4 (N10259, N10251, N10149, N6056, N6260);
not NOT1 (N10260, N10249);
not NOT1 (N10261, N10230);
nor NOR4 (N10262, N10255, N6184, N6955, N7136);
nor NOR3 (N10263, N10262, N8092, N4551);
nand NAND4 (N10264, N10258, N5867, N2837, N1696);
xor XOR2 (N10265, N10257, N4636);
and AND2 (N10266, N10261, N9274);
buf BUF1 (N10267, N10260);
not NOT1 (N10268, N10259);
or OR2 (N10269, N10268, N1263);
nand NAND4 (N10270, N10228, N7243, N1679, N2160);
xor XOR2 (N10271, N10242, N639);
buf BUF1 (N10272, N10256);
nor NOR4 (N10273, N10264, N5004, N2415, N1859);
xor XOR2 (N10274, N10267, N345);
nor NOR2 (N10275, N10271, N3326);
nor NOR3 (N10276, N10270, N4816, N1751);
xor XOR2 (N10277, N10274, N300);
buf BUF1 (N10278, N10265);
not NOT1 (N10279, N10278);
or OR3 (N10280, N10279, N201, N8259);
nor NOR4 (N10281, N10263, N9253, N7852, N3124);
not NOT1 (N10282, N10266);
xor XOR2 (N10283, N10269, N6503);
nor NOR4 (N10284, N10282, N1353, N4016, N7012);
or OR3 (N10285, N10277, N3338, N8364);
and AND2 (N10286, N10285, N9947);
and AND3 (N10287, N10250, N9105, N5733);
not NOT1 (N10288, N10273);
nand NAND3 (N10289, N10272, N6465, N7891);
and AND3 (N10290, N10284, N6377, N666);
nor NOR2 (N10291, N10287, N5174);
buf BUF1 (N10292, N10290);
and AND4 (N10293, N10280, N8075, N3546, N6572);
xor XOR2 (N10294, N10286, N4709);
not NOT1 (N10295, N10281);
and AND3 (N10296, N10275, N1192, N1522);
not NOT1 (N10297, N10294);
nor NOR2 (N10298, N10291, N4862);
not NOT1 (N10299, N10298);
not NOT1 (N10300, N10283);
and AND4 (N10301, N10276, N4125, N6870, N1873);
not NOT1 (N10302, N10288);
and AND4 (N10303, N10295, N3426, N10239, N3904);
or OR3 (N10304, N10289, N5990, N5756);
not NOT1 (N10305, N10293);
and AND2 (N10306, N10303, N8718);
or OR2 (N10307, N10300, N10013);
xor XOR2 (N10308, N10292, N9519);
not NOT1 (N10309, N10307);
buf BUF1 (N10310, N10299);
not NOT1 (N10311, N10306);
nor NOR2 (N10312, N10302, N2402);
not NOT1 (N10313, N10311);
nor NOR3 (N10314, N10309, N9064, N1435);
and AND4 (N10315, N10310, N3605, N2732, N5984);
or OR2 (N10316, N10314, N7560);
nor NOR4 (N10317, N10304, N7307, N4883, N2794);
buf BUF1 (N10318, N10315);
nand NAND4 (N10319, N10305, N5381, N10212, N6215);
nand NAND3 (N10320, N10308, N2370, N4674);
buf BUF1 (N10321, N10318);
xor XOR2 (N10322, N10297, N6404);
or OR3 (N10323, N10319, N2713, N5970);
or OR3 (N10324, N10321, N5381, N2093);
not NOT1 (N10325, N10312);
not NOT1 (N10326, N10317);
xor XOR2 (N10327, N10320, N6996);
xor XOR2 (N10328, N10325, N9769);
nor NOR3 (N10329, N10301, N6966, N7563);
xor XOR2 (N10330, N10316, N8714);
and AND2 (N10331, N10327, N6725);
and AND2 (N10332, N10328, N845);
nor NOR2 (N10333, N10296, N7903);
and AND4 (N10334, N10313, N9800, N3761, N2610);
or OR3 (N10335, N10334, N8917, N7222);
nor NOR2 (N10336, N10335, N6916);
and AND3 (N10337, N10333, N4613, N1018);
xor XOR2 (N10338, N10324, N3857);
xor XOR2 (N10339, N10332, N46);
nand NAND2 (N10340, N10322, N1213);
nand NAND2 (N10341, N10338, N386);
or OR4 (N10342, N10326, N10336, N1344, N7094);
xor XOR2 (N10343, N9502, N5059);
or OR3 (N10344, N10323, N164, N8763);
nor NOR4 (N10345, N10339, N2790, N9982, N3968);
nand NAND2 (N10346, N10341, N1227);
nor NOR3 (N10347, N10330, N5249, N3176);
nand NAND4 (N10348, N10329, N388, N6761, N5477);
buf BUF1 (N10349, N10344);
and AND4 (N10350, N10348, N1300, N7037, N2323);
nor NOR2 (N10351, N10337, N9316);
nor NOR3 (N10352, N10343, N7621, N9508);
nand NAND3 (N10353, N10349, N5769, N411);
or OR4 (N10354, N10350, N4805, N7471, N7286);
not NOT1 (N10355, N10346);
and AND4 (N10356, N10354, N5928, N4115, N3804);
nand NAND2 (N10357, N10356, N1018);
not NOT1 (N10358, N10357);
buf BUF1 (N10359, N10345);
nor NOR4 (N10360, N10351, N7039, N2702, N1261);
and AND2 (N10361, N10353, N7011);
nand NAND2 (N10362, N10360, N6064);
nand NAND2 (N10363, N10359, N2489);
not NOT1 (N10364, N10358);
nor NOR3 (N10365, N10364, N2297, N588);
nor NOR3 (N10366, N10342, N2995, N3636);
nand NAND2 (N10367, N10352, N1728);
xor XOR2 (N10368, N10355, N7806);
nor NOR3 (N10369, N10361, N428, N2948);
not NOT1 (N10370, N10363);
nor NOR3 (N10371, N10347, N1606, N8639);
and AND4 (N10372, N10367, N9078, N146, N5760);
nor NOR2 (N10373, N10366, N9363);
buf BUF1 (N10374, N10372);
or OR2 (N10375, N10374, N8687);
xor XOR2 (N10376, N10373, N1902);
nor NOR4 (N10377, N10340, N7823, N6044, N7706);
nand NAND3 (N10378, N10375, N10007, N7350);
or OR4 (N10379, N10362, N7753, N6957, N612);
not NOT1 (N10380, N10331);
nand NAND4 (N10381, N10368, N5678, N758, N10003);
and AND3 (N10382, N10377, N2624, N160);
not NOT1 (N10383, N10371);
buf BUF1 (N10384, N10378);
and AND3 (N10385, N10380, N2366, N5633);
and AND4 (N10386, N10379, N4896, N6465, N3266);
buf BUF1 (N10387, N10385);
not NOT1 (N10388, N10384);
and AND4 (N10389, N10370, N6707, N7336, N10125);
buf BUF1 (N10390, N10383);
or OR4 (N10391, N10387, N5246, N2084, N636);
or OR4 (N10392, N10382, N5640, N1620, N980);
or OR4 (N10393, N10392, N7516, N3461, N6740);
and AND2 (N10394, N10369, N5210);
and AND2 (N10395, N10376, N1909);
xor XOR2 (N10396, N10386, N1163);
or OR4 (N10397, N10391, N10053, N3239, N7381);
nand NAND3 (N10398, N10389, N3411, N4833);
nor NOR2 (N10399, N10394, N1596);
nor NOR4 (N10400, N10388, N2855, N6859, N7058);
xor XOR2 (N10401, N10396, N7357);
xor XOR2 (N10402, N10397, N4);
nor NOR4 (N10403, N10398, N5338, N8492, N9750);
and AND2 (N10404, N10403, N3371);
buf BUF1 (N10405, N10399);
nand NAND2 (N10406, N10390, N4674);
not NOT1 (N10407, N10381);
buf BUF1 (N10408, N10402);
buf BUF1 (N10409, N10406);
and AND4 (N10410, N10401, N107, N482, N6316);
nor NOR2 (N10411, N10400, N2794);
not NOT1 (N10412, N10365);
or OR3 (N10413, N10411, N5128, N6480);
nand NAND4 (N10414, N10404, N5922, N2402, N2783);
nand NAND4 (N10415, N10413, N10313, N10144, N10249);
buf BUF1 (N10416, N10410);
buf BUF1 (N10417, N10408);
nor NOR3 (N10418, N10417, N4350, N2215);
buf BUF1 (N10419, N10407);
nand NAND3 (N10420, N10395, N5343, N1551);
and AND3 (N10421, N10414, N3887, N6141);
nand NAND2 (N10422, N10415, N2537);
and AND3 (N10423, N10393, N1327, N2346);
not NOT1 (N10424, N10412);
or OR3 (N10425, N10422, N10318, N3324);
and AND2 (N10426, N10418, N5020);
and AND2 (N10427, N10425, N4862);
nand NAND4 (N10428, N10421, N2205, N6043, N471);
not NOT1 (N10429, N10409);
not NOT1 (N10430, N10427);
xor XOR2 (N10431, N10424, N3786);
nand NAND4 (N10432, N10429, N320, N2449, N4665);
and AND4 (N10433, N10431, N4358, N6547, N5659);
nand NAND2 (N10434, N10428, N5853);
xor XOR2 (N10435, N10423, N6928);
nor NOR3 (N10436, N10433, N3475, N9749);
nor NOR3 (N10437, N10435, N549, N5005);
not NOT1 (N10438, N10432);
and AND2 (N10439, N10436, N7446);
xor XOR2 (N10440, N10439, N1391);
not NOT1 (N10441, N10437);
nand NAND3 (N10442, N10416, N1276, N6801);
and AND3 (N10443, N10405, N8882, N3473);
buf BUF1 (N10444, N10426);
not NOT1 (N10445, N10442);
xor XOR2 (N10446, N10438, N5107);
nor NOR2 (N10447, N10444, N2099);
nand NAND4 (N10448, N10420, N2702, N3973, N3906);
xor XOR2 (N10449, N10419, N7577);
and AND4 (N10450, N10445, N4380, N2133, N8477);
not NOT1 (N10451, N10449);
or OR4 (N10452, N10448, N6783, N518, N6790);
and AND2 (N10453, N10446, N7404);
buf BUF1 (N10454, N10453);
xor XOR2 (N10455, N10450, N3126);
nor NOR4 (N10456, N10451, N965, N3906, N9914);
nor NOR2 (N10457, N10443, N5150);
nand NAND4 (N10458, N10441, N6924, N628, N9927);
buf BUF1 (N10459, N10454);
xor XOR2 (N10460, N10452, N10451);
or OR2 (N10461, N10434, N5236);
or OR4 (N10462, N10456, N620, N9585, N3486);
nand NAND2 (N10463, N10430, N1518);
and AND3 (N10464, N10455, N64, N8763);
and AND3 (N10465, N10440, N4961, N8986);
buf BUF1 (N10466, N10463);
xor XOR2 (N10467, N10461, N3249);
and AND2 (N10468, N10460, N5648);
nand NAND3 (N10469, N10457, N7002, N1671);
and AND3 (N10470, N10466, N6707, N1880);
or OR4 (N10471, N10467, N5223, N1775, N1432);
xor XOR2 (N10472, N10458, N5995);
nand NAND2 (N10473, N10468, N1211);
and AND3 (N10474, N10469, N1550, N5725);
nand NAND3 (N10475, N10459, N6797, N10431);
and AND2 (N10476, N10447, N4398);
buf BUF1 (N10477, N10470);
nand NAND4 (N10478, N10477, N7467, N886, N2628);
nor NOR2 (N10479, N10476, N5806);
xor XOR2 (N10480, N10474, N5507);
and AND4 (N10481, N10465, N7856, N5161, N6203);
buf BUF1 (N10482, N10479);
and AND2 (N10483, N10482, N616);
nor NOR2 (N10484, N10483, N809);
nor NOR2 (N10485, N10472, N1776);
or OR2 (N10486, N10485, N7113);
xor XOR2 (N10487, N10475, N5439);
nor NOR3 (N10488, N10462, N3035, N4697);
or OR4 (N10489, N10484, N8098, N3876, N1442);
xor XOR2 (N10490, N10488, N4740);
nor NOR4 (N10491, N10481, N1996, N1045, N8960);
buf BUF1 (N10492, N10478);
or OR3 (N10493, N10492, N4358, N10402);
nor NOR4 (N10494, N10489, N53, N4599, N2002);
or OR4 (N10495, N10487, N10118, N9628, N6573);
xor XOR2 (N10496, N10486, N37);
nor NOR2 (N10497, N10496, N7743);
nand NAND4 (N10498, N10497, N7728, N8916, N4315);
nor NOR3 (N10499, N10471, N9048, N9633);
xor XOR2 (N10500, N10495, N3293);
not NOT1 (N10501, N10493);
buf BUF1 (N10502, N10464);
and AND3 (N10503, N10500, N4246, N1832);
nand NAND2 (N10504, N10473, N10160);
and AND3 (N10505, N10494, N9480, N7138);
nor NOR2 (N10506, N10504, N7470);
and AND3 (N10507, N10498, N2083, N2336);
nor NOR4 (N10508, N10505, N896, N10295, N5027);
or OR2 (N10509, N10491, N5060);
buf BUF1 (N10510, N10507);
and AND3 (N10511, N10509, N4309, N9976);
and AND3 (N10512, N10490, N8277, N8423);
or OR3 (N10513, N10508, N5525, N8986);
nand NAND3 (N10514, N10511, N4406, N1390);
xor XOR2 (N10515, N10510, N7896);
not NOT1 (N10516, N10499);
nand NAND3 (N10517, N10516, N9819, N4559);
xor XOR2 (N10518, N10502, N3959);
xor XOR2 (N10519, N10515, N6446);
or OR4 (N10520, N10506, N5105, N9212, N9368);
or OR3 (N10521, N10520, N10358, N7524);
nand NAND3 (N10522, N10517, N6736, N6745);
or OR2 (N10523, N10512, N1812);
or OR2 (N10524, N10480, N4445);
not NOT1 (N10525, N10518);
buf BUF1 (N10526, N10525);
or OR2 (N10527, N10524, N7618);
nand NAND3 (N10528, N10501, N1407, N6651);
xor XOR2 (N10529, N10528, N9223);
or OR3 (N10530, N10522, N6368, N8562);
nor NOR3 (N10531, N10530, N6614, N5071);
and AND2 (N10532, N10529, N8770);
nor NOR4 (N10533, N10503, N319, N9520, N7717);
nor NOR2 (N10534, N10526, N98);
xor XOR2 (N10535, N10519, N2061);
or OR3 (N10536, N10514, N2715, N1725);
nor NOR4 (N10537, N10513, N4712, N869, N7086);
buf BUF1 (N10538, N10535);
xor XOR2 (N10539, N10527, N2051);
nor NOR2 (N10540, N10534, N2514);
xor XOR2 (N10541, N10523, N8598);
buf BUF1 (N10542, N10521);
nand NAND3 (N10543, N10532, N5609, N6447);
and AND3 (N10544, N10542, N809, N10147);
not NOT1 (N10545, N10537);
xor XOR2 (N10546, N10544, N9368);
not NOT1 (N10547, N10543);
not NOT1 (N10548, N10533);
nand NAND2 (N10549, N10547, N5030);
nand NAND4 (N10550, N10538, N5872, N9318, N1772);
and AND4 (N10551, N10540, N3823, N5992, N4450);
buf BUF1 (N10552, N10548);
or OR4 (N10553, N10551, N1601, N7113, N2521);
not NOT1 (N10554, N10546);
buf BUF1 (N10555, N10549);
buf BUF1 (N10556, N10545);
not NOT1 (N10557, N10552);
xor XOR2 (N10558, N10541, N7793);
nor NOR2 (N10559, N10553, N2571);
nor NOR3 (N10560, N10559, N7421, N5560);
and AND3 (N10561, N10550, N2955, N10030);
or OR3 (N10562, N10536, N2252, N3784);
nor NOR3 (N10563, N10560, N7156, N4405);
or OR3 (N10564, N10562, N8241, N4393);
xor XOR2 (N10565, N10554, N5585);
nand NAND4 (N10566, N10558, N6701, N530, N4883);
not NOT1 (N10567, N10556);
or OR4 (N10568, N10564, N227, N8589, N7845);
or OR4 (N10569, N10565, N267, N6770, N3042);
not NOT1 (N10570, N10569);
nand NAND4 (N10571, N10555, N10546, N5709, N2462);
buf BUF1 (N10572, N10563);
nor NOR4 (N10573, N10568, N397, N155, N1199);
or OR2 (N10574, N10561, N303);
buf BUF1 (N10575, N10566);
nand NAND3 (N10576, N10531, N4136, N8237);
not NOT1 (N10577, N10576);
nand NAND3 (N10578, N10577, N7833, N8840);
nand NAND2 (N10579, N10578, N6347);
nor NOR4 (N10580, N10575, N8127, N1307, N9000);
buf BUF1 (N10581, N10574);
buf BUF1 (N10582, N10567);
nand NAND3 (N10583, N10570, N7134, N8804);
nand NAND4 (N10584, N10581, N1432, N9732, N7840);
nand NAND2 (N10585, N10571, N8608);
or OR2 (N10586, N10585, N6917);
xor XOR2 (N10587, N10582, N839);
not NOT1 (N10588, N10583);
xor XOR2 (N10589, N10557, N3184);
buf BUF1 (N10590, N10539);
nor NOR4 (N10591, N10588, N1511, N3727, N4489);
or OR4 (N10592, N10586, N4520, N8597, N8323);
or OR2 (N10593, N10580, N10435);
buf BUF1 (N10594, N10590);
xor XOR2 (N10595, N10592, N7915);
or OR3 (N10596, N10589, N2508, N1589);
and AND4 (N10597, N10584, N1832, N4118, N1348);
or OR2 (N10598, N10595, N7622);
or OR3 (N10599, N10593, N6206, N23);
nand NAND4 (N10600, N10597, N3217, N9327, N2121);
nor NOR2 (N10601, N10598, N2993);
nand NAND3 (N10602, N10587, N7609, N419);
and AND3 (N10603, N10599, N2083, N7120);
nand NAND4 (N10604, N10579, N8284, N8392, N10270);
buf BUF1 (N10605, N10594);
buf BUF1 (N10606, N10596);
or OR2 (N10607, N10602, N7943);
or OR4 (N10608, N10603, N1076, N1236, N9888);
not NOT1 (N10609, N10607);
not NOT1 (N10610, N10573);
nand NAND2 (N10611, N10609, N7360);
buf BUF1 (N10612, N10591);
nor NOR4 (N10613, N10600, N9547, N9898, N3248);
nor NOR2 (N10614, N10604, N4005);
buf BUF1 (N10615, N10612);
nand NAND2 (N10616, N10601, N5161);
buf BUF1 (N10617, N10611);
not NOT1 (N10618, N10605);
nor NOR2 (N10619, N10608, N2939);
not NOT1 (N10620, N10613);
xor XOR2 (N10621, N10614, N6120);
not NOT1 (N10622, N10618);
or OR2 (N10623, N10572, N3669);
buf BUF1 (N10624, N10615);
nand NAND3 (N10625, N10620, N7321, N10383);
buf BUF1 (N10626, N10616);
not NOT1 (N10627, N10624);
nor NOR2 (N10628, N10627, N661);
nand NAND3 (N10629, N10621, N4399, N1162);
not NOT1 (N10630, N10622);
or OR3 (N10631, N10630, N9909, N4722);
or OR2 (N10632, N10623, N6738);
nand NAND2 (N10633, N10628, N5516);
nor NOR3 (N10634, N10625, N1357, N2814);
nor NOR2 (N10635, N10606, N5094);
xor XOR2 (N10636, N10634, N1798);
xor XOR2 (N10637, N10631, N3871);
or OR3 (N10638, N10617, N9101, N2797);
xor XOR2 (N10639, N10638, N5469);
nor NOR2 (N10640, N10632, N2148);
buf BUF1 (N10641, N10636);
nand NAND2 (N10642, N10637, N10037);
buf BUF1 (N10643, N10629);
nand NAND2 (N10644, N10635, N2637);
nor NOR3 (N10645, N10641, N7146, N6342);
or OR3 (N10646, N10642, N3788, N1517);
nand NAND4 (N10647, N10639, N7958, N5905, N1753);
or OR4 (N10648, N10644, N7764, N8830, N745);
and AND2 (N10649, N10643, N6435);
nand NAND3 (N10650, N10645, N4859, N3699);
buf BUF1 (N10651, N10633);
nand NAND3 (N10652, N10647, N4910, N2892);
not NOT1 (N10653, N10651);
xor XOR2 (N10654, N10653, N1974);
nand NAND4 (N10655, N10610, N3299, N6893, N10032);
nor NOR2 (N10656, N10655, N3106);
xor XOR2 (N10657, N10619, N1009);
buf BUF1 (N10658, N10640);
and AND3 (N10659, N10650, N9691, N10066);
or OR3 (N10660, N10658, N5028, N1979);
nand NAND3 (N10661, N10660, N3684, N1911);
or OR4 (N10662, N10646, N2401, N3177, N115);
or OR3 (N10663, N10649, N3614, N2335);
xor XOR2 (N10664, N10652, N1319);
not NOT1 (N10665, N10663);
nand NAND3 (N10666, N10659, N9836, N1738);
buf BUF1 (N10667, N10648);
nand NAND4 (N10668, N10661, N474, N7048, N9138);
xor XOR2 (N10669, N10657, N1030);
nand NAND3 (N10670, N10662, N8826, N10553);
nand NAND2 (N10671, N10669, N6950);
and AND4 (N10672, N10667, N5423, N6680, N10179);
buf BUF1 (N10673, N10664);
or OR4 (N10674, N10672, N7980, N5592, N9579);
or OR3 (N10675, N10665, N909, N9852);
nand NAND2 (N10676, N10666, N2959);
nand NAND4 (N10677, N10654, N2203, N2123, N7847);
buf BUF1 (N10678, N10668);
nand NAND3 (N10679, N10678, N9415, N10128);
nor NOR3 (N10680, N10670, N466, N4976);
xor XOR2 (N10681, N10674, N1033);
and AND3 (N10682, N10677, N3060, N7360);
not NOT1 (N10683, N10656);
nand NAND2 (N10684, N10682, N3197);
buf BUF1 (N10685, N10675);
or OR2 (N10686, N10671, N8072);
not NOT1 (N10687, N10680);
xor XOR2 (N10688, N10626, N7578);
xor XOR2 (N10689, N10684, N10322);
xor XOR2 (N10690, N10688, N7357);
buf BUF1 (N10691, N10685);
nand NAND2 (N10692, N10683, N754);
and AND2 (N10693, N10681, N5236);
nand NAND4 (N10694, N10691, N6317, N9446, N8929);
nand NAND4 (N10695, N10679, N8282, N9882, N7705);
xor XOR2 (N10696, N10687, N10674);
and AND3 (N10697, N10694, N4664, N4565);
not NOT1 (N10698, N10696);
not NOT1 (N10699, N10695);
and AND3 (N10700, N10673, N2606, N5338);
nand NAND4 (N10701, N10693, N6551, N3658, N3749);
or OR4 (N10702, N10690, N1928, N7352, N5196);
and AND2 (N10703, N10702, N8390);
and AND2 (N10704, N10676, N1563);
nor NOR3 (N10705, N10703, N2976, N6355);
and AND3 (N10706, N10698, N4504, N1435);
buf BUF1 (N10707, N10701);
and AND3 (N10708, N10699, N5780, N1550);
nand NAND3 (N10709, N10697, N8453, N9053);
and AND3 (N10710, N10689, N4028, N5007);
xor XOR2 (N10711, N10709, N8985);
nor NOR2 (N10712, N10707, N999);
nand NAND3 (N10713, N10705, N276, N8071);
buf BUF1 (N10714, N10692);
buf BUF1 (N10715, N10686);
or OR4 (N10716, N10712, N5597, N3110, N8262);
buf BUF1 (N10717, N10710);
nand NAND4 (N10718, N10716, N5102, N3916, N10543);
not NOT1 (N10719, N10708);
nor NOR2 (N10720, N10718, N8388);
nor NOR4 (N10721, N10714, N7952, N8395, N3973);
not NOT1 (N10722, N10719);
not NOT1 (N10723, N10720);
or OR2 (N10724, N10721, N2397);
or OR3 (N10725, N10706, N292, N7837);
and AND3 (N10726, N10704, N6633, N8013);
nand NAND4 (N10727, N10700, N1361, N10041, N3625);
and AND3 (N10728, N10713, N4608, N6621);
and AND3 (N10729, N10724, N10611, N860);
not NOT1 (N10730, N10722);
nand NAND2 (N10731, N10727, N4221);
or OR4 (N10732, N10726, N933, N3846, N6119);
not NOT1 (N10733, N10728);
xor XOR2 (N10734, N10715, N1271);
nor NOR3 (N10735, N10733, N4121, N2829);
not NOT1 (N10736, N10732);
nor NOR3 (N10737, N10711, N8296, N5685);
nor NOR3 (N10738, N10737, N6171, N5364);
and AND2 (N10739, N10723, N8210);
buf BUF1 (N10740, N10739);
xor XOR2 (N10741, N10738, N3895);
xor XOR2 (N10742, N10735, N6508);
buf BUF1 (N10743, N10741);
xor XOR2 (N10744, N10725, N708);
xor XOR2 (N10745, N10730, N3964);
buf BUF1 (N10746, N10740);
nand NAND4 (N10747, N10744, N4596, N3395, N5700);
or OR3 (N10748, N10734, N9341, N3367);
xor XOR2 (N10749, N10717, N3395);
nor NOR3 (N10750, N10743, N7683, N4319);
not NOT1 (N10751, N10745);
buf BUF1 (N10752, N10742);
and AND3 (N10753, N10748, N9849, N3839);
or OR3 (N10754, N10749, N2718, N10138);
and AND4 (N10755, N10729, N360, N2068, N3507);
or OR2 (N10756, N10731, N2049);
or OR3 (N10757, N10752, N7044, N6408);
and AND4 (N10758, N10755, N3755, N492, N6173);
buf BUF1 (N10759, N10751);
not NOT1 (N10760, N10758);
nor NOR2 (N10761, N10747, N8903);
xor XOR2 (N10762, N10759, N125);
nor NOR3 (N10763, N10753, N9947, N4984);
not NOT1 (N10764, N10736);
xor XOR2 (N10765, N10763, N8247);
or OR4 (N10766, N10757, N2475, N7618, N8793);
nor NOR2 (N10767, N10761, N5141);
and AND3 (N10768, N10765, N3491, N1974);
buf BUF1 (N10769, N10764);
xor XOR2 (N10770, N10746, N6558);
or OR2 (N10771, N10769, N4778);
not NOT1 (N10772, N10756);
nand NAND4 (N10773, N10762, N10719, N3378, N3647);
nor NOR2 (N10774, N10771, N3312);
xor XOR2 (N10775, N10767, N4955);
and AND4 (N10776, N10766, N5435, N5705, N9003);
and AND2 (N10777, N10772, N4290);
or OR2 (N10778, N10760, N3579);
or OR3 (N10779, N10776, N3334, N2911);
or OR4 (N10780, N10768, N1815, N3411, N2706);
buf BUF1 (N10781, N10780);
xor XOR2 (N10782, N10777, N10168);
xor XOR2 (N10783, N10775, N2966);
and AND3 (N10784, N10774, N2045, N2031);
xor XOR2 (N10785, N10778, N10329);
nand NAND3 (N10786, N10783, N2563, N6725);
nor NOR2 (N10787, N10750, N7150);
not NOT1 (N10788, N10779);
nor NOR3 (N10789, N10770, N8067, N4772);
or OR3 (N10790, N10786, N8744, N10035);
not NOT1 (N10791, N10781);
xor XOR2 (N10792, N10773, N7435);
buf BUF1 (N10793, N10787);
nor NOR2 (N10794, N10790, N3721);
buf BUF1 (N10795, N10788);
nand NAND3 (N10796, N10792, N8977, N1824);
buf BUF1 (N10797, N10754);
xor XOR2 (N10798, N10785, N3645);
not NOT1 (N10799, N10797);
not NOT1 (N10800, N10798);
or OR3 (N10801, N10789, N9887, N2704);
xor XOR2 (N10802, N10796, N9225);
and AND4 (N10803, N10793, N2352, N8781, N3319);
nand NAND3 (N10804, N10784, N8475, N9120);
or OR4 (N10805, N10800, N2066, N662, N9646);
or OR3 (N10806, N10804, N8480, N5560);
xor XOR2 (N10807, N10795, N9266);
not NOT1 (N10808, N10791);
xor XOR2 (N10809, N10806, N8656);
and AND3 (N10810, N10805, N767, N4985);
nor NOR3 (N10811, N10808, N9076, N9367);
not NOT1 (N10812, N10810);
not NOT1 (N10813, N10802);
xor XOR2 (N10814, N10813, N3440);
and AND2 (N10815, N10811, N8618);
nor NOR4 (N10816, N10809, N4677, N6813, N7568);
and AND4 (N10817, N10803, N6981, N3083, N1278);
buf BUF1 (N10818, N10815);
not NOT1 (N10819, N10807);
xor XOR2 (N10820, N10816, N6437);
and AND2 (N10821, N10799, N3310);
and AND4 (N10822, N10819, N5419, N9776, N7321);
and AND2 (N10823, N10820, N936);
not NOT1 (N10824, N10821);
buf BUF1 (N10825, N10823);
or OR3 (N10826, N10782, N5115, N10378);
buf BUF1 (N10827, N10822);
buf BUF1 (N10828, N10812);
buf BUF1 (N10829, N10801);
and AND3 (N10830, N10825, N10094, N5060);
and AND3 (N10831, N10814, N3180, N4896);
nor NOR4 (N10832, N10826, N7090, N6018, N7531);
or OR4 (N10833, N10829, N123, N8316, N4969);
nand NAND3 (N10834, N10830, N8981, N9701);
or OR4 (N10835, N10818, N10102, N1456, N1051);
nand NAND2 (N10836, N10835, N1483);
and AND2 (N10837, N10834, N5128);
or OR3 (N10838, N10837, N10643, N8940);
xor XOR2 (N10839, N10836, N2234);
nor NOR4 (N10840, N10828, N7291, N3697, N5740);
and AND4 (N10841, N10831, N1769, N3955, N6816);
or OR2 (N10842, N10839, N10504);
xor XOR2 (N10843, N10838, N8447);
and AND3 (N10844, N10842, N6830, N9765);
xor XOR2 (N10845, N10832, N4733);
and AND2 (N10846, N10794, N5876);
or OR2 (N10847, N10846, N4965);
xor XOR2 (N10848, N10845, N7623);
or OR3 (N10849, N10827, N3539, N10566);
or OR3 (N10850, N10844, N7105, N990);
and AND4 (N10851, N10843, N3916, N6214, N4864);
buf BUF1 (N10852, N10817);
or OR2 (N10853, N10852, N3787);
and AND3 (N10854, N10840, N8982, N4428);
or OR4 (N10855, N10854, N3560, N1437, N1641);
xor XOR2 (N10856, N10848, N7996);
or OR4 (N10857, N10853, N5022, N4762, N1805);
not NOT1 (N10858, N10856);
nor NOR2 (N10859, N10841, N795);
nor NOR4 (N10860, N10824, N2493, N10476, N6536);
and AND2 (N10861, N10849, N7014);
buf BUF1 (N10862, N10855);
xor XOR2 (N10863, N10851, N7778);
xor XOR2 (N10864, N10857, N5247);
buf BUF1 (N10865, N10862);
and AND4 (N10866, N10861, N5860, N5524, N5903);
xor XOR2 (N10867, N10863, N360);
buf BUF1 (N10868, N10867);
buf BUF1 (N10869, N10859);
and AND3 (N10870, N10865, N3026, N7776);
nand NAND2 (N10871, N10850, N6284);
and AND2 (N10872, N10833, N1578);
and AND4 (N10873, N10870, N6483, N7295, N10575);
or OR2 (N10874, N10868, N3806);
nor NOR2 (N10875, N10873, N2378);
nor NOR3 (N10876, N10869, N3893, N5522);
not NOT1 (N10877, N10864);
and AND3 (N10878, N10875, N2533, N5197);
not NOT1 (N10879, N10872);
buf BUF1 (N10880, N10879);
buf BUF1 (N10881, N10858);
and AND2 (N10882, N10871, N241);
nand NAND4 (N10883, N10877, N1276, N6406, N10654);
or OR4 (N10884, N10881, N1043, N5338, N6720);
buf BUF1 (N10885, N10880);
buf BUF1 (N10886, N10885);
xor XOR2 (N10887, N10866, N6727);
buf BUF1 (N10888, N10878);
buf BUF1 (N10889, N10886);
nor NOR4 (N10890, N10888, N8904, N917, N2420);
and AND2 (N10891, N10874, N8210);
or OR3 (N10892, N10883, N1497, N4975);
and AND3 (N10893, N10860, N3518, N9671);
buf BUF1 (N10894, N10891);
and AND4 (N10895, N10890, N2944, N9461, N10392);
nand NAND2 (N10896, N10884, N3114);
and AND4 (N10897, N10892, N5663, N2626, N9634);
nand NAND4 (N10898, N10894, N8312, N2901, N3026);
not NOT1 (N10899, N10897);
not NOT1 (N10900, N10882);
buf BUF1 (N10901, N10899);
and AND2 (N10902, N10900, N8685);
not NOT1 (N10903, N10876);
buf BUF1 (N10904, N10887);
and AND4 (N10905, N10893, N5157, N9628, N7313);
buf BUF1 (N10906, N10902);
nor NOR2 (N10907, N10898, N8703);
not NOT1 (N10908, N10903);
nor NOR2 (N10909, N10904, N885);
or OR4 (N10910, N10901, N2844, N10732, N2172);
and AND3 (N10911, N10896, N5056, N3073);
and AND3 (N10912, N10847, N3929, N5482);
or OR3 (N10913, N10906, N1715, N1849);
buf BUF1 (N10914, N10908);
and AND2 (N10915, N10912, N10549);
not NOT1 (N10916, N10910);
and AND3 (N10917, N10916, N7696, N3928);
buf BUF1 (N10918, N10909);
not NOT1 (N10919, N10911);
buf BUF1 (N10920, N10918);
nand NAND3 (N10921, N10915, N7186, N3450);
or OR2 (N10922, N10889, N3578);
xor XOR2 (N10923, N10922, N791);
and AND3 (N10924, N10913, N5656, N5117);
nor NOR4 (N10925, N10923, N7325, N4869, N6377);
nand NAND3 (N10926, N10905, N2082, N3959);
or OR4 (N10927, N10925, N9287, N538, N6942);
nand NAND2 (N10928, N10919, N6051);
xor XOR2 (N10929, N10895, N7527);
xor XOR2 (N10930, N10907, N3586);
or OR4 (N10931, N10924, N8606, N8070, N3101);
xor XOR2 (N10932, N10927, N10153);
nor NOR3 (N10933, N10928, N1548, N5921);
not NOT1 (N10934, N10931);
nand NAND4 (N10935, N10917, N7747, N9269, N5228);
nand NAND4 (N10936, N10933, N10622, N2838, N8477);
or OR3 (N10937, N10932, N191, N1559);
and AND3 (N10938, N10937, N523, N5643);
nor NOR4 (N10939, N10921, N2304, N10578, N9110);
nand NAND3 (N10940, N10935, N2546, N2973);
xor XOR2 (N10941, N10934, N8247);
nand NAND4 (N10942, N10914, N10742, N649, N2494);
or OR4 (N10943, N10941, N2431, N10358, N3880);
buf BUF1 (N10944, N10942);
buf BUF1 (N10945, N10926);
buf BUF1 (N10946, N10936);
nor NOR2 (N10947, N10938, N490);
or OR2 (N10948, N10940, N3998);
nor NOR2 (N10949, N10929, N5044);
not NOT1 (N10950, N10946);
nor NOR2 (N10951, N10943, N7511);
or OR3 (N10952, N10944, N8080, N6177);
or OR3 (N10953, N10948, N7977, N917);
xor XOR2 (N10954, N10949, N2719);
or OR3 (N10955, N10954, N7199, N9741);
xor XOR2 (N10956, N10955, N9802);
or OR4 (N10957, N10953, N1318, N7149, N2079);
xor XOR2 (N10958, N10956, N7559);
or OR3 (N10959, N10930, N8685, N6452);
nand NAND2 (N10960, N10920, N5128);
or OR3 (N10961, N10959, N4167, N8586);
and AND2 (N10962, N10951, N9008);
or OR3 (N10963, N10961, N8053, N10431);
and AND2 (N10964, N10957, N2291);
nand NAND3 (N10965, N10964, N3795, N10766);
xor XOR2 (N10966, N10947, N6657);
buf BUF1 (N10967, N10966);
buf BUF1 (N10968, N10939);
or OR3 (N10969, N10963, N2432, N2671);
and AND3 (N10970, N10965, N8846, N9258);
nand NAND2 (N10971, N10960, N8655);
nand NAND4 (N10972, N10969, N9219, N2152, N2591);
or OR2 (N10973, N10972, N8035);
xor XOR2 (N10974, N10968, N7398);
or OR4 (N10975, N10971, N1521, N2781, N5243);
buf BUF1 (N10976, N10973);
nand NAND4 (N10977, N10952, N4849, N5473, N9378);
or OR4 (N10978, N10950, N56, N1330, N7349);
and AND2 (N10979, N10962, N8972);
not NOT1 (N10980, N10978);
buf BUF1 (N10981, N10967);
and AND2 (N10982, N10981, N10213);
xor XOR2 (N10983, N10976, N2854);
nand NAND2 (N10984, N10979, N2936);
nand NAND4 (N10985, N10983, N8366, N6796, N5815);
nand NAND2 (N10986, N10975, N5319);
not NOT1 (N10987, N10986);
nand NAND4 (N10988, N10977, N4759, N10893, N1369);
nand NAND3 (N10989, N10970, N7759, N3029);
buf BUF1 (N10990, N10984);
nor NOR3 (N10991, N10988, N5261, N4793);
nand NAND2 (N10992, N10990, N10932);
xor XOR2 (N10993, N10980, N7562);
nand NAND2 (N10994, N10945, N2396);
or OR2 (N10995, N10974, N115);
xor XOR2 (N10996, N10958, N697);
or OR2 (N10997, N10992, N10513);
buf BUF1 (N10998, N10989);
and AND4 (N10999, N10997, N1452, N6381, N10058);
nor NOR2 (N11000, N10995, N2004);
buf BUF1 (N11001, N10993);
nand NAND3 (N11002, N10985, N5905, N5981);
nor NOR3 (N11003, N10999, N4764, N3536);
buf BUF1 (N11004, N11001);
nor NOR2 (N11005, N10982, N8998);
not NOT1 (N11006, N10991);
buf BUF1 (N11007, N10996);
and AND2 (N11008, N11006, N10696);
or OR3 (N11009, N10998, N4922, N10013);
nand NAND2 (N11010, N11009, N3191);
buf BUF1 (N11011, N11008);
nand NAND2 (N11012, N11010, N9830);
buf BUF1 (N11013, N11011);
xor XOR2 (N11014, N11007, N1703);
buf BUF1 (N11015, N10994);
buf BUF1 (N11016, N11014);
nand NAND3 (N11017, N11000, N6829, N2102);
or OR4 (N11018, N11012, N8210, N7909, N7601);
and AND3 (N11019, N11018, N4359, N6761);
buf BUF1 (N11020, N11017);
not NOT1 (N11021, N11020);
nand NAND4 (N11022, N11003, N9836, N5120, N6895);
not NOT1 (N11023, N11021);
buf BUF1 (N11024, N11015);
nand NAND2 (N11025, N11004, N9789);
and AND4 (N11026, N11002, N6577, N4307, N2010);
nand NAND2 (N11027, N11019, N8946);
xor XOR2 (N11028, N11016, N1515);
buf BUF1 (N11029, N10987);
nor NOR2 (N11030, N11024, N6542);
xor XOR2 (N11031, N11030, N2366);
or OR3 (N11032, N11027, N507, N8125);
not NOT1 (N11033, N11028);
and AND2 (N11034, N11022, N1099);
not NOT1 (N11035, N11026);
nor NOR2 (N11036, N11035, N968);
xor XOR2 (N11037, N11034, N8508);
not NOT1 (N11038, N11031);
nand NAND2 (N11039, N11038, N6291);
not NOT1 (N11040, N11036);
nor NOR3 (N11041, N11032, N136, N7692);
not NOT1 (N11042, N11041);
nand NAND3 (N11043, N11039, N1204, N1932);
nor NOR2 (N11044, N11040, N1315);
buf BUF1 (N11045, N11029);
nor NOR4 (N11046, N11042, N6240, N10140, N4184);
nand NAND4 (N11047, N11033, N1941, N10834, N9888);
or OR3 (N11048, N11013, N946, N7837);
xor XOR2 (N11049, N11043, N3199);
not NOT1 (N11050, N11045);
not NOT1 (N11051, N11025);
nor NOR3 (N11052, N11046, N3491, N8202);
xor XOR2 (N11053, N11005, N5617);
and AND3 (N11054, N11023, N4896, N783);
not NOT1 (N11055, N11054);
or OR3 (N11056, N11037, N7813, N782);
not NOT1 (N11057, N11053);
nand NAND4 (N11058, N11056, N2592, N9686, N9733);
buf BUF1 (N11059, N11050);
and AND3 (N11060, N11044, N906, N7505);
nor NOR2 (N11061, N11047, N4623);
buf BUF1 (N11062, N11060);
nand NAND2 (N11063, N11061, N2416);
nor NOR2 (N11064, N11052, N10840);
not NOT1 (N11065, N11064);
buf BUF1 (N11066, N11058);
not NOT1 (N11067, N11057);
nand NAND2 (N11068, N11051, N5654);
buf BUF1 (N11069, N11055);
buf BUF1 (N11070, N11065);
not NOT1 (N11071, N11066);
nor NOR4 (N11072, N11059, N5646, N4400, N9619);
not NOT1 (N11073, N11070);
nor NOR2 (N11074, N11068, N2532);
or OR4 (N11075, N11062, N6381, N2751, N9532);
or OR2 (N11076, N11073, N4512);
nand NAND2 (N11077, N11067, N9906);
buf BUF1 (N11078, N11075);
xor XOR2 (N11079, N11072, N4821);
and AND3 (N11080, N11071, N2016, N2662);
or OR3 (N11081, N11063, N7807, N2552);
and AND4 (N11082, N11079, N7491, N9511, N2488);
and AND4 (N11083, N11076, N3254, N8379, N1405);
and AND3 (N11084, N11048, N9434, N9865);
xor XOR2 (N11085, N11069, N2951);
nand NAND4 (N11086, N11081, N7935, N10380, N2314);
xor XOR2 (N11087, N11086, N10750);
xor XOR2 (N11088, N11082, N6675);
nor NOR3 (N11089, N11077, N730, N8371);
or OR3 (N11090, N11084, N96, N3027);
and AND3 (N11091, N11090, N11087, N3426);
nor NOR3 (N11092, N4528, N4460, N10855);
and AND2 (N11093, N11092, N3190);
xor XOR2 (N11094, N11078, N6540);
xor XOR2 (N11095, N11091, N6204);
not NOT1 (N11096, N11080);
not NOT1 (N11097, N11095);
nand NAND2 (N11098, N11088, N7827);
or OR4 (N11099, N11097, N5742, N9393, N6383);
or OR2 (N11100, N11074, N9568);
buf BUF1 (N11101, N11100);
nand NAND4 (N11102, N11093, N3112, N4871, N3662);
not NOT1 (N11103, N11049);
and AND4 (N11104, N11103, N8675, N1444, N1956);
nand NAND2 (N11105, N11102, N10518);
and AND3 (N11106, N11085, N8545, N4484);
or OR4 (N11107, N11096, N5828, N10199, N9278);
nand NAND2 (N11108, N11089, N2782);
buf BUF1 (N11109, N11099);
nand NAND2 (N11110, N11094, N4513);
nand NAND3 (N11111, N11106, N2280, N3473);
nor NOR4 (N11112, N11111, N3809, N4388, N4804);
and AND3 (N11113, N11112, N2427, N6778);
or OR4 (N11114, N11109, N1874, N8852, N4538);
nand NAND2 (N11115, N11083, N3340);
xor XOR2 (N11116, N11098, N4288);
or OR4 (N11117, N11105, N7353, N4589, N6880);
buf BUF1 (N11118, N11101);
not NOT1 (N11119, N11104);
not NOT1 (N11120, N11107);
or OR4 (N11121, N11117, N5098, N2109, N750);
and AND2 (N11122, N11119, N990);
not NOT1 (N11123, N11122);
not NOT1 (N11124, N11114);
xor XOR2 (N11125, N11123, N5036);
nor NOR2 (N11126, N11113, N10771);
nand NAND4 (N11127, N11115, N1260, N5738, N2327);
buf BUF1 (N11128, N11118);
not NOT1 (N11129, N11124);
nor NOR3 (N11130, N11127, N7392, N8744);
xor XOR2 (N11131, N11110, N3781);
nor NOR2 (N11132, N11121, N6468);
buf BUF1 (N11133, N11108);
and AND4 (N11134, N11132, N6096, N6148, N10719);
xor XOR2 (N11135, N11116, N367);
buf BUF1 (N11136, N11133);
not NOT1 (N11137, N11131);
and AND3 (N11138, N11129, N8730, N7516);
nand NAND3 (N11139, N11137, N5384, N9943);
or OR2 (N11140, N11125, N8166);
not NOT1 (N11141, N11136);
xor XOR2 (N11142, N11141, N7518);
and AND2 (N11143, N11140, N3242);
not NOT1 (N11144, N11120);
nor NOR4 (N11145, N11138, N7204, N3649, N2988);
xor XOR2 (N11146, N11145, N3530);
nand NAND3 (N11147, N11144, N100, N8450);
buf BUF1 (N11148, N11126);
nor NOR3 (N11149, N11146, N2835, N2150);
nor NOR4 (N11150, N11148, N7733, N1386, N429);
nor NOR4 (N11151, N11135, N10429, N5889, N3854);
nor NOR3 (N11152, N11150, N785, N4247);
nand NAND2 (N11153, N11147, N8258);
buf BUF1 (N11154, N11134);
nor NOR4 (N11155, N11153, N10676, N8633, N3914);
nor NOR4 (N11156, N11151, N245, N6135, N799);
nand NAND2 (N11157, N11142, N4616);
not NOT1 (N11158, N11149);
xor XOR2 (N11159, N11154, N222);
and AND3 (N11160, N11158, N4452, N789);
buf BUF1 (N11161, N11143);
buf BUF1 (N11162, N11157);
buf BUF1 (N11163, N11130);
buf BUF1 (N11164, N11161);
or OR3 (N11165, N11156, N8603, N6195);
nand NAND2 (N11166, N11128, N4115);
nor NOR4 (N11167, N11159, N10276, N8595, N5075);
and AND4 (N11168, N11139, N2260, N5192, N4407);
xor XOR2 (N11169, N11164, N10441);
nor NOR4 (N11170, N11155, N8058, N5970, N5174);
nand NAND3 (N11171, N11170, N316, N9936);
buf BUF1 (N11172, N11168);
buf BUF1 (N11173, N11163);
xor XOR2 (N11174, N11172, N8822);
not NOT1 (N11175, N11173);
xor XOR2 (N11176, N11160, N263);
nand NAND2 (N11177, N11167, N10836);
or OR4 (N11178, N11174, N3262, N7810, N5453);
nor NOR3 (N11179, N11171, N4636, N5416);
xor XOR2 (N11180, N11178, N3174);
and AND2 (N11181, N11166, N10472);
buf BUF1 (N11182, N11177);
or OR4 (N11183, N11165, N7121, N10889, N4823);
xor XOR2 (N11184, N11181, N6879);
xor XOR2 (N11185, N11184, N10606);
xor XOR2 (N11186, N11175, N81);
buf BUF1 (N11187, N11183);
and AND2 (N11188, N11176, N1028);
buf BUF1 (N11189, N11185);
or OR3 (N11190, N11187, N5982, N3612);
xor XOR2 (N11191, N11162, N172);
nor NOR2 (N11192, N11179, N5271);
buf BUF1 (N11193, N11182);
not NOT1 (N11194, N11193);
xor XOR2 (N11195, N11192, N6405);
or OR4 (N11196, N11191, N9128, N799, N10678);
not NOT1 (N11197, N11189);
nor NOR3 (N11198, N11190, N9418, N6082);
xor XOR2 (N11199, N11196, N9280);
buf BUF1 (N11200, N11194);
not NOT1 (N11201, N11195);
xor XOR2 (N11202, N11188, N9418);
not NOT1 (N11203, N11198);
xor XOR2 (N11204, N11203, N6928);
buf BUF1 (N11205, N11201);
xor XOR2 (N11206, N11197, N7276);
xor XOR2 (N11207, N11180, N6636);
nand NAND4 (N11208, N11204, N637, N7162, N1898);
and AND3 (N11209, N11206, N7261, N8865);
buf BUF1 (N11210, N11208);
buf BUF1 (N11211, N11199);
xor XOR2 (N11212, N11205, N3664);
nor NOR2 (N11213, N11169, N8092);
nand NAND4 (N11214, N11212, N5380, N104, N3535);
buf BUF1 (N11215, N11186);
nand NAND3 (N11216, N11202, N2589, N627);
nor NOR4 (N11217, N11209, N8595, N8916, N3052);
and AND2 (N11218, N11214, N7977);
xor XOR2 (N11219, N11152, N3180);
nand NAND3 (N11220, N11213, N4697, N7939);
nand NAND4 (N11221, N11200, N900, N9744, N1180);
or OR4 (N11222, N11221, N8307, N11121, N6372);
not NOT1 (N11223, N11210);
or OR4 (N11224, N11223, N3742, N8143, N2340);
nand NAND2 (N11225, N11215, N2932);
nand NAND4 (N11226, N11219, N674, N4861, N2111);
not NOT1 (N11227, N11218);
xor XOR2 (N11228, N11227, N10387);
nand NAND4 (N11229, N11211, N5843, N7839, N5744);
xor XOR2 (N11230, N11224, N8495);
nand NAND2 (N11231, N11226, N10777);
or OR2 (N11232, N11229, N9053);
and AND3 (N11233, N11216, N2634, N4374);
buf BUF1 (N11234, N11232);
or OR4 (N11235, N11231, N2920, N2068, N5029);
and AND3 (N11236, N11220, N5573, N9920);
nand NAND3 (N11237, N11235, N4186, N9458);
xor XOR2 (N11238, N11228, N3657);
and AND4 (N11239, N11225, N3120, N4922, N2344);
nand NAND3 (N11240, N11234, N6083, N628);
and AND4 (N11241, N11240, N9144, N5048, N11180);
nand NAND4 (N11242, N11239, N8562, N10088, N2543);
and AND4 (N11243, N11238, N1157, N115, N9887);
and AND2 (N11244, N11222, N3244);
nor NOR3 (N11245, N11217, N8235, N10494);
not NOT1 (N11246, N11207);
not NOT1 (N11247, N11243);
nor NOR4 (N11248, N11242, N5270, N7337, N193);
nor NOR4 (N11249, N11233, N843, N9213, N8783);
and AND2 (N11250, N11230, N10903);
nor NOR2 (N11251, N11237, N5704);
and AND3 (N11252, N11251, N2065, N10846);
nand NAND2 (N11253, N11249, N322);
buf BUF1 (N11254, N11248);
nor NOR3 (N11255, N11253, N4532, N7087);
not NOT1 (N11256, N11236);
and AND3 (N11257, N11255, N9562, N10378);
buf BUF1 (N11258, N11245);
not NOT1 (N11259, N11250);
buf BUF1 (N11260, N11246);
nor NOR2 (N11261, N11244, N710);
or OR2 (N11262, N11259, N8417);
not NOT1 (N11263, N11258);
or OR3 (N11264, N11263, N2692, N8925);
nor NOR4 (N11265, N11264, N2767, N356, N11079);
nor NOR2 (N11266, N11241, N5236);
nor NOR2 (N11267, N11266, N8509);
xor XOR2 (N11268, N11265, N9095);
xor XOR2 (N11269, N11268, N10377);
nor NOR3 (N11270, N11252, N4895, N4697);
buf BUF1 (N11271, N11261);
buf BUF1 (N11272, N11267);
buf BUF1 (N11273, N11262);
nand NAND4 (N11274, N11271, N4778, N7051, N8478);
not NOT1 (N11275, N11274);
not NOT1 (N11276, N11257);
xor XOR2 (N11277, N11270, N563);
xor XOR2 (N11278, N11269, N8381);
or OR2 (N11279, N11260, N7032);
not NOT1 (N11280, N11277);
nand NAND4 (N11281, N11272, N8623, N6605, N3836);
not NOT1 (N11282, N11276);
or OR3 (N11283, N11275, N6728, N10001);
or OR3 (N11284, N11256, N2771, N6277);
buf BUF1 (N11285, N11283);
nor NOR4 (N11286, N11254, N3797, N3291, N8899);
buf BUF1 (N11287, N11282);
or OR3 (N11288, N11284, N2956, N3771);
not NOT1 (N11289, N11278);
or OR4 (N11290, N11280, N8778, N7238, N2441);
and AND3 (N11291, N11289, N319, N786);
or OR3 (N11292, N11287, N9160, N4341);
xor XOR2 (N11293, N11292, N6410);
nand NAND2 (N11294, N11273, N1354);
nor NOR3 (N11295, N11279, N7821, N10099);
or OR2 (N11296, N11291, N6607);
and AND3 (N11297, N11295, N2688, N2481);
xor XOR2 (N11298, N11281, N5874);
buf BUF1 (N11299, N11290);
nand NAND2 (N11300, N11299, N5590);
or OR3 (N11301, N11286, N3499, N3436);
not NOT1 (N11302, N11293);
buf BUF1 (N11303, N11285);
or OR4 (N11304, N11247, N6151, N4020, N8071);
buf BUF1 (N11305, N11300);
and AND2 (N11306, N11304, N9650);
and AND2 (N11307, N11297, N945);
xor XOR2 (N11308, N11306, N3898);
not NOT1 (N11309, N11298);
not NOT1 (N11310, N11308);
nor NOR3 (N11311, N11309, N6303, N3251);
not NOT1 (N11312, N11294);
and AND2 (N11313, N11312, N6682);
or OR2 (N11314, N11313, N7722);
or OR3 (N11315, N11310, N5629, N4722);
not NOT1 (N11316, N11305);
nor NOR4 (N11317, N11316, N10946, N1866, N7271);
nor NOR3 (N11318, N11302, N7092, N9158);
xor XOR2 (N11319, N11314, N10669);
and AND3 (N11320, N11307, N10148, N7428);
not NOT1 (N11321, N11317);
and AND2 (N11322, N11296, N2115);
nand NAND4 (N11323, N11321, N341, N9632, N8207);
buf BUF1 (N11324, N11319);
buf BUF1 (N11325, N11288);
nand NAND4 (N11326, N11303, N5536, N6431, N7235);
or OR2 (N11327, N11323, N4572);
nor NOR4 (N11328, N11301, N6177, N9445, N8436);
buf BUF1 (N11329, N11328);
nand NAND3 (N11330, N11325, N2250, N1946);
buf BUF1 (N11331, N11315);
and AND4 (N11332, N11320, N3599, N955, N3979);
and AND2 (N11333, N11326, N9480);
buf BUF1 (N11334, N11333);
and AND2 (N11335, N11334, N4142);
xor XOR2 (N11336, N11311, N10282);
or OR4 (N11337, N11330, N3628, N152, N6933);
xor XOR2 (N11338, N11336, N6147);
buf BUF1 (N11339, N11318);
not NOT1 (N11340, N11337);
buf BUF1 (N11341, N11322);
xor XOR2 (N11342, N11339, N7191);
and AND2 (N11343, N11341, N7588);
or OR2 (N11344, N11332, N6492);
nand NAND4 (N11345, N11331, N8062, N3508, N5396);
nand NAND3 (N11346, N11342, N6740, N3987);
and AND4 (N11347, N11335, N1005, N7064, N4684);
nor NOR4 (N11348, N11329, N3129, N9404, N3361);
or OR4 (N11349, N11324, N5851, N994, N1572);
and AND4 (N11350, N11346, N2406, N6983, N9976);
nand NAND2 (N11351, N11347, N2906);
xor XOR2 (N11352, N11338, N2962);
nand NAND4 (N11353, N11345, N9775, N6166, N6853);
xor XOR2 (N11354, N11344, N3249);
buf BUF1 (N11355, N11349);
buf BUF1 (N11356, N11351);
xor XOR2 (N11357, N11356, N5968);
buf BUF1 (N11358, N11343);
and AND2 (N11359, N11355, N10704);
nor NOR4 (N11360, N11340, N710, N2620, N1030);
and AND2 (N11361, N11357, N5866);
nand NAND4 (N11362, N11359, N4080, N1682, N7078);
xor XOR2 (N11363, N11327, N7739);
buf BUF1 (N11364, N11363);
nor NOR4 (N11365, N11354, N3496, N3268, N7235);
or OR3 (N11366, N11364, N10983, N5358);
nor NOR3 (N11367, N11362, N2103, N10916);
nand NAND3 (N11368, N11366, N10666, N11071);
xor XOR2 (N11369, N11353, N1077);
xor XOR2 (N11370, N11361, N7604);
not NOT1 (N11371, N11352);
not NOT1 (N11372, N11368);
buf BUF1 (N11373, N11358);
and AND4 (N11374, N11350, N113, N10089, N2905);
or OR4 (N11375, N11374, N11163, N273, N8700);
nor NOR2 (N11376, N11373, N2724);
and AND2 (N11377, N11375, N8217);
or OR2 (N11378, N11365, N10954);
xor XOR2 (N11379, N11376, N5291);
nand NAND3 (N11380, N11348, N875, N2161);
nor NOR2 (N11381, N11379, N10251);
not NOT1 (N11382, N11377);
and AND4 (N11383, N11369, N10118, N6776, N9291);
and AND3 (N11384, N11382, N6721, N2678);
or OR4 (N11385, N11380, N5888, N8206, N1059);
or OR2 (N11386, N11381, N10761);
buf BUF1 (N11387, N11370);
nand NAND3 (N11388, N11384, N5862, N1657);
nand NAND2 (N11389, N11385, N3766);
nor NOR3 (N11390, N11388, N3073, N10415);
not NOT1 (N11391, N11387);
xor XOR2 (N11392, N11390, N2598);
and AND3 (N11393, N11372, N4192, N6964);
nand NAND3 (N11394, N11386, N2211, N2704);
nor NOR3 (N11395, N11394, N2028, N4658);
or OR2 (N11396, N11389, N4761);
not NOT1 (N11397, N11392);
nor NOR3 (N11398, N11391, N5227, N6496);
not NOT1 (N11399, N11396);
not NOT1 (N11400, N11393);
or OR3 (N11401, N11399, N501, N10550);
or OR2 (N11402, N11367, N10882);
or OR2 (N11403, N11402, N8992);
nand NAND2 (N11404, N11400, N10306);
or OR3 (N11405, N11378, N3326, N4370);
buf BUF1 (N11406, N11371);
nand NAND4 (N11407, N11360, N1345, N1183, N1606);
nor NOR4 (N11408, N11395, N3129, N9108, N10354);
or OR3 (N11409, N11407, N6360, N230);
and AND2 (N11410, N11408, N9293);
nor NOR2 (N11411, N11403, N1137);
nand NAND3 (N11412, N11406, N7858, N10900);
nor NOR2 (N11413, N11383, N1274);
nor NOR2 (N11414, N11398, N3178);
nand NAND4 (N11415, N11410, N6500, N4532, N1859);
buf BUF1 (N11416, N11411);
or OR3 (N11417, N11415, N8082, N6254);
buf BUF1 (N11418, N11401);
nor NOR3 (N11419, N11416, N4258, N3757);
nor NOR2 (N11420, N11405, N11042);
nand NAND4 (N11421, N11404, N2456, N8000, N11307);
buf BUF1 (N11422, N11413);
nand NAND2 (N11423, N11414, N535);
and AND2 (N11424, N11421, N3539);
nand NAND4 (N11425, N11419, N7831, N1177, N2587);
buf BUF1 (N11426, N11417);
nor NOR4 (N11427, N11418, N10831, N8527, N1312);
xor XOR2 (N11428, N11412, N9138);
xor XOR2 (N11429, N11426, N239);
nand NAND4 (N11430, N11425, N10854, N504, N6180);
nor NOR3 (N11431, N11424, N9694, N6793);
nand NAND2 (N11432, N11427, N6523);
buf BUF1 (N11433, N11397);
or OR3 (N11434, N11430, N3154, N6069);
and AND2 (N11435, N11409, N7251);
xor XOR2 (N11436, N11431, N8699);
nor NOR4 (N11437, N11423, N7240, N7676, N9693);
xor XOR2 (N11438, N11429, N5172);
and AND4 (N11439, N11438, N4383, N1336, N8419);
nand NAND3 (N11440, N11422, N280, N3931);
nand NAND2 (N11441, N11437, N10510);
not NOT1 (N11442, N11432);
or OR4 (N11443, N11436, N2936, N3573, N3718);
nand NAND2 (N11444, N11428, N4818);
nor NOR3 (N11445, N11420, N2894, N8115);
not NOT1 (N11446, N11441);
not NOT1 (N11447, N11442);
xor XOR2 (N11448, N11446, N4108);
and AND2 (N11449, N11434, N1513);
not NOT1 (N11450, N11443);
buf BUF1 (N11451, N11435);
and AND2 (N11452, N11449, N3098);
nor NOR2 (N11453, N11445, N6846);
xor XOR2 (N11454, N11448, N10239);
and AND4 (N11455, N11450, N7501, N8184, N10627);
nand NAND4 (N11456, N11454, N3575, N9665, N8281);
xor XOR2 (N11457, N11440, N7002);
nor NOR2 (N11458, N11433, N3140);
and AND3 (N11459, N11453, N672, N3373);
buf BUF1 (N11460, N11451);
buf BUF1 (N11461, N11459);
or OR3 (N11462, N11458, N10236, N2396);
or OR4 (N11463, N11455, N11139, N6815, N2943);
nand NAND2 (N11464, N11457, N463);
not NOT1 (N11465, N11460);
or OR2 (N11466, N11462, N701);
or OR4 (N11467, N11439, N3327, N9534, N7076);
not NOT1 (N11468, N11466);
and AND2 (N11469, N11463, N11361);
nor NOR4 (N11470, N11452, N5310, N8078, N4781);
nor NOR2 (N11471, N11467, N9040);
xor XOR2 (N11472, N11469, N2640);
not NOT1 (N11473, N11465);
nand NAND4 (N11474, N11456, N145, N7354, N3372);
or OR2 (N11475, N11474, N2882);
not NOT1 (N11476, N11470);
nor NOR3 (N11477, N11444, N1815, N5208);
xor XOR2 (N11478, N11461, N2635);
not NOT1 (N11479, N11476);
nor NOR3 (N11480, N11468, N9182, N10670);
and AND4 (N11481, N11477, N5372, N51, N899);
buf BUF1 (N11482, N11478);
or OR4 (N11483, N11480, N4887, N2318, N8795);
buf BUF1 (N11484, N11479);
and AND4 (N11485, N11483, N1429, N1283, N2571);
not NOT1 (N11486, N11481);
nand NAND4 (N11487, N11473, N380, N5051, N3801);
or OR3 (N11488, N11487, N2187, N10513);
or OR4 (N11489, N11488, N5096, N3464, N7906);
nand NAND2 (N11490, N11475, N4127);
or OR2 (N11491, N11471, N10467);
and AND2 (N11492, N11490, N9715);
or OR2 (N11493, N11491, N5691);
xor XOR2 (N11494, N11472, N4338);
nor NOR4 (N11495, N11492, N1607, N6363, N6885);
xor XOR2 (N11496, N11495, N5997);
or OR4 (N11497, N11482, N2383, N10376, N3388);
and AND3 (N11498, N11485, N5568, N8753);
not NOT1 (N11499, N11494);
xor XOR2 (N11500, N11493, N8683);
not NOT1 (N11501, N11489);
or OR3 (N11502, N11501, N10807, N5948);
nand NAND4 (N11503, N11484, N8389, N11099, N476);
xor XOR2 (N11504, N11447, N4081);
nor NOR3 (N11505, N11464, N6428, N10855);
and AND3 (N11506, N11496, N1151, N6000);
not NOT1 (N11507, N11505);
or OR3 (N11508, N11503, N10976, N1812);
buf BUF1 (N11509, N11497);
nor NOR2 (N11510, N11502, N10367);
nand NAND2 (N11511, N11504, N10956);
nor NOR2 (N11512, N11510, N4902);
or OR4 (N11513, N11511, N7566, N9962, N9173);
and AND4 (N11514, N11508, N3946, N3452, N11251);
nor NOR2 (N11515, N11498, N4607);
nor NOR3 (N11516, N11500, N9832, N8822);
or OR2 (N11517, N11516, N156);
buf BUF1 (N11518, N11499);
or OR2 (N11519, N11509, N6279);
and AND3 (N11520, N11507, N2641, N7530);
xor XOR2 (N11521, N11486, N7420);
not NOT1 (N11522, N11506);
nor NOR3 (N11523, N11521, N1525, N9156);
xor XOR2 (N11524, N11523, N8348);
nor NOR4 (N11525, N11520, N9549, N9908, N5517);
and AND4 (N11526, N11525, N4031, N1808, N5633);
nor NOR3 (N11527, N11515, N5112, N8857);
not NOT1 (N11528, N11527);
not NOT1 (N11529, N11524);
buf BUF1 (N11530, N11512);
not NOT1 (N11531, N11529);
xor XOR2 (N11532, N11519, N2262);
buf BUF1 (N11533, N11532);
buf BUF1 (N11534, N11533);
not NOT1 (N11535, N11513);
nor NOR2 (N11536, N11517, N1915);
and AND4 (N11537, N11522, N6752, N11493, N6107);
or OR4 (N11538, N11534, N3475, N10464, N8175);
buf BUF1 (N11539, N11526);
or OR2 (N11540, N11536, N6754);
buf BUF1 (N11541, N11538);
xor XOR2 (N11542, N11535, N4373);
nand NAND2 (N11543, N11539, N10009);
nor NOR3 (N11544, N11543, N7807, N6259);
or OR4 (N11545, N11528, N5806, N870, N4492);
nor NOR4 (N11546, N11531, N8665, N9699, N8114);
buf BUF1 (N11547, N11518);
xor XOR2 (N11548, N11537, N3378);
not NOT1 (N11549, N11547);
not NOT1 (N11550, N11541);
buf BUF1 (N11551, N11549);
or OR3 (N11552, N11550, N2557, N10367);
and AND4 (N11553, N11545, N7692, N9996, N11304);
or OR3 (N11554, N11552, N11050, N3262);
and AND2 (N11555, N11553, N4679);
not NOT1 (N11556, N11530);
xor XOR2 (N11557, N11540, N8392);
xor XOR2 (N11558, N11546, N1423);
and AND3 (N11559, N11542, N9171, N255);
nand NAND2 (N11560, N11559, N7229);
buf BUF1 (N11561, N11557);
nor NOR3 (N11562, N11556, N8680, N1919);
buf BUF1 (N11563, N11551);
nand NAND4 (N11564, N11562, N1832, N472, N4417);
not NOT1 (N11565, N11560);
and AND4 (N11566, N11564, N2889, N100, N11559);
and AND3 (N11567, N11565, N3763, N3431);
nand NAND2 (N11568, N11555, N4870);
xor XOR2 (N11569, N11561, N7023);
or OR4 (N11570, N11514, N5146, N10965, N2883);
and AND2 (N11571, N11567, N8834);
or OR4 (N11572, N11569, N9321, N2916, N2381);
buf BUF1 (N11573, N11572);
xor XOR2 (N11574, N11568, N1795);
and AND3 (N11575, N11570, N1927, N7565);
xor XOR2 (N11576, N11554, N5059);
not NOT1 (N11577, N11573);
or OR2 (N11578, N11563, N6153);
buf BUF1 (N11579, N11577);
or OR2 (N11580, N11548, N8349);
buf BUF1 (N11581, N11574);
not NOT1 (N11582, N11581);
xor XOR2 (N11583, N11582, N2605);
and AND4 (N11584, N11571, N478, N3207, N7761);
xor XOR2 (N11585, N11580, N7166);
and AND4 (N11586, N11576, N10143, N59, N2892);
and AND4 (N11587, N11579, N3, N4467, N1062);
nand NAND2 (N11588, N11544, N3352);
nor NOR2 (N11589, N11586, N1236);
nor NOR3 (N11590, N11578, N4475, N4415);
nand NAND4 (N11591, N11587, N10406, N8426, N5751);
xor XOR2 (N11592, N11583, N6911);
nor NOR2 (N11593, N11588, N5857);
not NOT1 (N11594, N11585);
buf BUF1 (N11595, N11589);
and AND4 (N11596, N11593, N5298, N456, N4253);
xor XOR2 (N11597, N11594, N905);
nand NAND2 (N11598, N11558, N7316);
not NOT1 (N11599, N11596);
buf BUF1 (N11600, N11598);
buf BUF1 (N11601, N11599);
buf BUF1 (N11602, N11584);
or OR3 (N11603, N11590, N1516, N7731);
nor NOR2 (N11604, N11592, N10862);
or OR4 (N11605, N11597, N11079, N3873, N10296);
and AND4 (N11606, N11605, N5948, N11049, N1633);
not NOT1 (N11607, N11591);
nand NAND4 (N11608, N11607, N1341, N6156, N2582);
buf BUF1 (N11609, N11566);
nor NOR3 (N11610, N11595, N10209, N6877);
nand NAND3 (N11611, N11610, N7337, N214);
buf BUF1 (N11612, N11611);
buf BUF1 (N11613, N11606);
or OR4 (N11614, N11601, N7566, N10490, N4677);
nand NAND3 (N11615, N11614, N10784, N10716);
or OR3 (N11616, N11608, N10937, N8846);
or OR3 (N11617, N11616, N6821, N10411);
and AND4 (N11618, N11612, N8830, N1114, N9839);
xor XOR2 (N11619, N11600, N3400);
not NOT1 (N11620, N11615);
xor XOR2 (N11621, N11618, N6008);
xor XOR2 (N11622, N11609, N2715);
buf BUF1 (N11623, N11604);
nand NAND3 (N11624, N11623, N6346, N9270);
nor NOR4 (N11625, N11613, N6507, N302, N156);
not NOT1 (N11626, N11617);
nor NOR2 (N11627, N11603, N6803);
buf BUF1 (N11628, N11625);
and AND3 (N11629, N11622, N8186, N3134);
not NOT1 (N11630, N11627);
or OR2 (N11631, N11620, N9350);
or OR3 (N11632, N11629, N8470, N8474);
and AND3 (N11633, N11630, N11503, N11534);
not NOT1 (N11634, N11631);
xor XOR2 (N11635, N11624, N213);
not NOT1 (N11636, N11621);
not NOT1 (N11637, N11626);
buf BUF1 (N11638, N11575);
not NOT1 (N11639, N11636);
buf BUF1 (N11640, N11637);
and AND3 (N11641, N11632, N10313, N8792);
and AND2 (N11642, N11634, N4376);
nand NAND2 (N11643, N11602, N11303);
buf BUF1 (N11644, N11633);
buf BUF1 (N11645, N11640);
nand NAND3 (N11646, N11644, N6991, N4235);
nor NOR3 (N11647, N11645, N4531, N7631);
nand NAND2 (N11648, N11646, N6837);
nor NOR2 (N11649, N11639, N8929);
nand NAND3 (N11650, N11642, N11423, N4628);
buf BUF1 (N11651, N11628);
nand NAND3 (N11652, N11648, N10106, N934);
nor NOR2 (N11653, N11650, N1418);
nor NOR3 (N11654, N11641, N11265, N7976);
buf BUF1 (N11655, N11643);
not NOT1 (N11656, N11649);
nor NOR2 (N11657, N11638, N5251);
and AND2 (N11658, N11651, N7140);
and AND2 (N11659, N11635, N3225);
and AND2 (N11660, N11654, N2809);
not NOT1 (N11661, N11647);
and AND4 (N11662, N11619, N8936, N10688, N2968);
and AND2 (N11663, N11657, N412);
buf BUF1 (N11664, N11663);
not NOT1 (N11665, N11659);
not NOT1 (N11666, N11664);
or OR3 (N11667, N11661, N8337, N8026);
nand NAND2 (N11668, N11652, N1779);
nor NOR4 (N11669, N11665, N6209, N2645, N6309);
nor NOR3 (N11670, N11668, N2734, N4402);
nor NOR2 (N11671, N11658, N10613);
xor XOR2 (N11672, N11671, N7752);
not NOT1 (N11673, N11669);
xor XOR2 (N11674, N11667, N7920);
nor NOR3 (N11675, N11653, N4600, N10825);
buf BUF1 (N11676, N11670);
xor XOR2 (N11677, N11676, N5869);
nor NOR2 (N11678, N11660, N7457);
not NOT1 (N11679, N11672);
buf BUF1 (N11680, N11675);
buf BUF1 (N11681, N11662);
xor XOR2 (N11682, N11678, N3187);
not NOT1 (N11683, N11674);
nand NAND3 (N11684, N11679, N4201, N1);
nor NOR3 (N11685, N11680, N9816, N825);
and AND3 (N11686, N11666, N638, N4710);
nor NOR2 (N11687, N11681, N6925);
buf BUF1 (N11688, N11686);
nor NOR3 (N11689, N11684, N2108, N9816);
xor XOR2 (N11690, N11655, N10987);
or OR3 (N11691, N11685, N928, N5467);
xor XOR2 (N11692, N11673, N2541);
and AND3 (N11693, N11688, N8264, N648);
xor XOR2 (N11694, N11689, N6715);
xor XOR2 (N11695, N11690, N1637);
xor XOR2 (N11696, N11692, N9909);
xor XOR2 (N11697, N11696, N6029);
or OR2 (N11698, N11683, N8686);
or OR3 (N11699, N11697, N8843, N3857);
or OR2 (N11700, N11693, N1290);
or OR2 (N11701, N11691, N8881);
nor NOR2 (N11702, N11700, N7675);
not NOT1 (N11703, N11701);
nand NAND2 (N11704, N11698, N6536);
or OR3 (N11705, N11699, N11333, N11633);
and AND2 (N11706, N11656, N8454);
or OR3 (N11707, N11702, N4746, N4833);
xor XOR2 (N11708, N11677, N8718);
and AND2 (N11709, N11703, N8828);
xor XOR2 (N11710, N11706, N7256);
not NOT1 (N11711, N11710);
nand NAND2 (N11712, N11705, N10382);
or OR3 (N11713, N11712, N11673, N9981);
nor NOR3 (N11714, N11695, N10582, N10465);
buf BUF1 (N11715, N11694);
or OR2 (N11716, N11714, N5515);
nor NOR3 (N11717, N11709, N9172, N8256);
nor NOR3 (N11718, N11707, N3305, N3302);
xor XOR2 (N11719, N11715, N9696);
buf BUF1 (N11720, N11682);
and AND4 (N11721, N11717, N2249, N5135, N6194);
or OR3 (N11722, N11704, N6223, N5169);
or OR4 (N11723, N11718, N3390, N9494, N6716);
buf BUF1 (N11724, N11720);
buf BUF1 (N11725, N11716);
xor XOR2 (N11726, N11722, N10438);
not NOT1 (N11727, N11721);
buf BUF1 (N11728, N11719);
not NOT1 (N11729, N11726);
nand NAND3 (N11730, N11708, N9058, N9972);
buf BUF1 (N11731, N11725);
nor NOR4 (N11732, N11724, N8616, N4306, N10708);
xor XOR2 (N11733, N11731, N6107);
or OR2 (N11734, N11727, N1235);
or OR4 (N11735, N11728, N10311, N1915, N11189);
not NOT1 (N11736, N11729);
and AND3 (N11737, N11734, N3057, N6900);
and AND2 (N11738, N11735, N11397);
nor NOR2 (N11739, N11732, N8651);
or OR4 (N11740, N11733, N5528, N1716, N10177);
not NOT1 (N11741, N11687);
nor NOR4 (N11742, N11711, N2790, N2139, N5042);
or OR4 (N11743, N11736, N11438, N11257, N5963);
not NOT1 (N11744, N11723);
buf BUF1 (N11745, N11713);
buf BUF1 (N11746, N11739);
buf BUF1 (N11747, N11740);
nand NAND3 (N11748, N11747, N421, N11487);
or OR3 (N11749, N11744, N10795, N9080);
nand NAND3 (N11750, N11737, N7651, N7596);
and AND3 (N11751, N11738, N4362, N1700);
or OR2 (N11752, N11745, N4357);
nor NOR3 (N11753, N11741, N6374, N864);
or OR2 (N11754, N11746, N11210);
nand NAND2 (N11755, N11750, N3022);
nor NOR3 (N11756, N11730, N6177, N4790);
nor NOR2 (N11757, N11749, N3697);
nor NOR3 (N11758, N11742, N8739, N11285);
not NOT1 (N11759, N11748);
or OR4 (N11760, N11743, N7294, N2535, N4098);
not NOT1 (N11761, N11757);
and AND4 (N11762, N11752, N797, N4830, N9033);
not NOT1 (N11763, N11754);
buf BUF1 (N11764, N11753);
nand NAND2 (N11765, N11751, N3660);
and AND4 (N11766, N11760, N10839, N8950, N8385);
buf BUF1 (N11767, N11764);
nand NAND2 (N11768, N11765, N5366);
nand NAND3 (N11769, N11755, N8901, N8209);
and AND3 (N11770, N11768, N11454, N875);
or OR2 (N11771, N11759, N10735);
or OR4 (N11772, N11758, N5654, N4178, N4308);
and AND3 (N11773, N11761, N7115, N10483);
not NOT1 (N11774, N11767);
and AND2 (N11775, N11774, N625);
xor XOR2 (N11776, N11762, N9104);
nand NAND2 (N11777, N11773, N10563);
not NOT1 (N11778, N11766);
or OR4 (N11779, N11772, N6052, N6470, N5096);
and AND4 (N11780, N11779, N3227, N6359, N11082);
nor NOR2 (N11781, N11776, N9677);
and AND2 (N11782, N11756, N1865);
buf BUF1 (N11783, N11770);
xor XOR2 (N11784, N11781, N8590);
xor XOR2 (N11785, N11775, N4331);
buf BUF1 (N11786, N11782);
buf BUF1 (N11787, N11769);
and AND4 (N11788, N11787, N11215, N7411, N5709);
nand NAND4 (N11789, N11786, N3506, N653, N6835);
and AND2 (N11790, N11789, N8683);
xor XOR2 (N11791, N11780, N112);
and AND4 (N11792, N11771, N11346, N9710, N10851);
buf BUF1 (N11793, N11777);
not NOT1 (N11794, N11790);
nand NAND2 (N11795, N11785, N2902);
not NOT1 (N11796, N11792);
nand NAND4 (N11797, N11788, N5666, N7356, N1160);
not NOT1 (N11798, N11795);
xor XOR2 (N11799, N11784, N4509);
xor XOR2 (N11800, N11794, N5810);
not NOT1 (N11801, N11800);
nor NOR3 (N11802, N11796, N5741, N2040);
nor NOR3 (N11803, N11763, N9402, N4872);
not NOT1 (N11804, N11793);
nand NAND4 (N11805, N11802, N4848, N48, N7338);
and AND3 (N11806, N11799, N1982, N11556);
not NOT1 (N11807, N11791);
or OR3 (N11808, N11805, N8077, N11230);
not NOT1 (N11809, N11807);
xor XOR2 (N11810, N11798, N1332);
buf BUF1 (N11811, N11806);
nand NAND3 (N11812, N11808, N7523, N11402);
nand NAND2 (N11813, N11809, N4704);
not NOT1 (N11814, N11812);
and AND4 (N11815, N11804, N10035, N477, N5426);
nand NAND3 (N11816, N11778, N5162, N1362);
buf BUF1 (N11817, N11801);
and AND4 (N11818, N11783, N7747, N9298, N9745);
nor NOR2 (N11819, N11813, N3380);
nor NOR2 (N11820, N11816, N11099);
nor NOR4 (N11821, N11820, N10409, N4659, N5965);
nor NOR3 (N11822, N11803, N6410, N5758);
or OR2 (N11823, N11797, N10056);
or OR2 (N11824, N11814, N2598);
and AND3 (N11825, N11823, N11470, N693);
nor NOR3 (N11826, N11819, N1413, N8795);
xor XOR2 (N11827, N11818, N260);
nand NAND2 (N11828, N11827, N9307);
nand NAND4 (N11829, N11826, N6446, N6195, N6683);
not NOT1 (N11830, N11828);
not NOT1 (N11831, N11822);
nand NAND4 (N11832, N11829, N8965, N9889, N5932);
buf BUF1 (N11833, N11824);
and AND4 (N11834, N11810, N8998, N988, N5268);
xor XOR2 (N11835, N11817, N1418);
xor XOR2 (N11836, N11835, N3267);
nand NAND4 (N11837, N11815, N7470, N2336, N2186);
xor XOR2 (N11838, N11830, N11689);
and AND3 (N11839, N11834, N10521, N2370);
nor NOR2 (N11840, N11837, N11406);
and AND2 (N11841, N11838, N9975);
xor XOR2 (N11842, N11836, N11484);
xor XOR2 (N11843, N11841, N4730);
xor XOR2 (N11844, N11825, N11202);
or OR4 (N11845, N11839, N8504, N3172, N2540);
buf BUF1 (N11846, N11821);
or OR3 (N11847, N11833, N8306, N7746);
nand NAND3 (N11848, N11811, N4199, N9793);
buf BUF1 (N11849, N11832);
and AND2 (N11850, N11847, N598);
nor NOR4 (N11851, N11846, N9702, N7050, N5820);
xor XOR2 (N11852, N11849, N4344);
buf BUF1 (N11853, N11851);
nor NOR4 (N11854, N11840, N7746, N7751, N8501);
nand NAND2 (N11855, N11842, N11404);
and AND2 (N11856, N11852, N6210);
and AND3 (N11857, N11855, N4904, N7202);
nand NAND2 (N11858, N11843, N11003);
nor NOR4 (N11859, N11857, N5004, N11450, N7187);
xor XOR2 (N11860, N11844, N1899);
or OR3 (N11861, N11853, N1452, N4998);
xor XOR2 (N11862, N11860, N8939);
and AND2 (N11863, N11861, N7049);
or OR4 (N11864, N11854, N7705, N11276, N4634);
buf BUF1 (N11865, N11856);
not NOT1 (N11866, N11831);
nor NOR2 (N11867, N11862, N10596);
xor XOR2 (N11868, N11865, N9982);
not NOT1 (N11869, N11859);
or OR3 (N11870, N11863, N10638, N6267);
not NOT1 (N11871, N11850);
buf BUF1 (N11872, N11868);
not NOT1 (N11873, N11866);
nor NOR2 (N11874, N11858, N8779);
not NOT1 (N11875, N11873);
or OR3 (N11876, N11870, N10490, N2653);
nand NAND3 (N11877, N11867, N10796, N10883);
buf BUF1 (N11878, N11877);
nand NAND2 (N11879, N11869, N828);
or OR2 (N11880, N11872, N8404);
buf BUF1 (N11881, N11864);
nor NOR4 (N11882, N11875, N3994, N2035, N8052);
and AND3 (N11883, N11880, N2788, N1470);
nand NAND4 (N11884, N11848, N6171, N11279, N3093);
xor XOR2 (N11885, N11878, N817);
xor XOR2 (N11886, N11845, N5256);
nand NAND2 (N11887, N11886, N2422);
or OR2 (N11888, N11887, N415);
nor NOR4 (N11889, N11879, N10421, N6803, N2718);
buf BUF1 (N11890, N11882);
xor XOR2 (N11891, N11888, N10328);
xor XOR2 (N11892, N11871, N11245);
xor XOR2 (N11893, N11881, N4888);
and AND2 (N11894, N11883, N2353);
nand NAND2 (N11895, N11890, N1458);
nor NOR3 (N11896, N11891, N5288, N8398);
not NOT1 (N11897, N11896);
or OR3 (N11898, N11893, N7369, N11595);
or OR2 (N11899, N11892, N5315);
or OR2 (N11900, N11895, N10117);
and AND4 (N11901, N11884, N769, N10715, N1331);
not NOT1 (N11902, N11885);
buf BUF1 (N11903, N11898);
nor NOR4 (N11904, N11876, N11018, N11791, N11087);
not NOT1 (N11905, N11901);
and AND3 (N11906, N11900, N7975, N8023);
or OR4 (N11907, N11894, N6172, N2293, N4862);
nand NAND2 (N11908, N11897, N6365);
not NOT1 (N11909, N11906);
nand NAND3 (N11910, N11899, N1777, N5839);
nand NAND3 (N11911, N11907, N11413, N354);
xor XOR2 (N11912, N11905, N3209);
nor NOR3 (N11913, N11911, N2711, N7948);
buf BUF1 (N11914, N11889);
not NOT1 (N11915, N11909);
not NOT1 (N11916, N11904);
not NOT1 (N11917, N11908);
xor XOR2 (N11918, N11913, N3057);
xor XOR2 (N11919, N11902, N6695);
xor XOR2 (N11920, N11919, N3752);
xor XOR2 (N11921, N11910, N1193);
and AND4 (N11922, N11914, N666, N530, N7447);
buf BUF1 (N11923, N11903);
nor NOR4 (N11924, N11923, N5756, N3411, N8998);
nor NOR2 (N11925, N11921, N10417);
or OR2 (N11926, N11920, N4154);
buf BUF1 (N11927, N11924);
nand NAND2 (N11928, N11926, N9009);
buf BUF1 (N11929, N11917);
xor XOR2 (N11930, N11929, N5248);
nand NAND3 (N11931, N11925, N994, N9381);
xor XOR2 (N11932, N11922, N2153);
and AND3 (N11933, N11918, N5039, N4025);
nor NOR2 (N11934, N11915, N4577);
nor NOR3 (N11935, N11933, N7, N5054);
xor XOR2 (N11936, N11932, N954);
not NOT1 (N11937, N11935);
and AND2 (N11938, N11937, N10820);
nor NOR3 (N11939, N11874, N2636, N8365);
or OR2 (N11940, N11934, N600);
xor XOR2 (N11941, N11940, N4397);
xor XOR2 (N11942, N11938, N4781);
not NOT1 (N11943, N11936);
not NOT1 (N11944, N11942);
and AND2 (N11945, N11939, N2235);
buf BUF1 (N11946, N11931);
buf BUF1 (N11947, N11945);
nor NOR3 (N11948, N11912, N8208, N770);
xor XOR2 (N11949, N11930, N2713);
not NOT1 (N11950, N11946);
buf BUF1 (N11951, N11927);
and AND4 (N11952, N11928, N11476, N3091, N229);
or OR2 (N11953, N11947, N6929);
nand NAND2 (N11954, N11949, N11136);
nor NOR2 (N11955, N11951, N5316);
xor XOR2 (N11956, N11943, N2291);
or OR3 (N11957, N11950, N573, N2148);
nand NAND3 (N11958, N11952, N8335, N7478);
nor NOR2 (N11959, N11948, N11650);
nand NAND4 (N11960, N11958, N1806, N1152, N6573);
nand NAND3 (N11961, N11956, N8248, N6329);
nand NAND2 (N11962, N11954, N4079);
and AND3 (N11963, N11953, N857, N3711);
buf BUF1 (N11964, N11941);
nor NOR4 (N11965, N11961, N11337, N6516, N10758);
buf BUF1 (N11966, N11965);
buf BUF1 (N11967, N11916);
xor XOR2 (N11968, N11959, N7658);
buf BUF1 (N11969, N11964);
or OR2 (N11970, N11967, N2781);
xor XOR2 (N11971, N11963, N294);
nand NAND3 (N11972, N11969, N8647, N11227);
nor NOR4 (N11973, N11966, N5468, N3826, N11163);
and AND4 (N11974, N11957, N11123, N8102, N7859);
not NOT1 (N11975, N11973);
and AND2 (N11976, N11968, N7658);
nand NAND3 (N11977, N11970, N8428, N5775);
xor XOR2 (N11978, N11955, N5483);
and AND2 (N11979, N11972, N4381);
nor NOR3 (N11980, N11979, N7214, N10151);
nand NAND3 (N11981, N11980, N8118, N7409);
buf BUF1 (N11982, N11960);
and AND3 (N11983, N11962, N4494, N4405);
nand NAND2 (N11984, N11983, N2762);
nor NOR2 (N11985, N11982, N1935);
xor XOR2 (N11986, N11977, N10324);
xor XOR2 (N11987, N11985, N2759);
or OR4 (N11988, N11975, N2204, N767, N6068);
xor XOR2 (N11989, N11986, N3038);
buf BUF1 (N11990, N11944);
nor NOR2 (N11991, N11990, N11507);
nor NOR4 (N11992, N11987, N2650, N10996, N5892);
nand NAND4 (N11993, N11989, N1271, N3787, N6897);
or OR3 (N11994, N11974, N2932, N6851);
or OR3 (N11995, N11978, N6360, N5732);
not NOT1 (N11996, N11995);
xor XOR2 (N11997, N11971, N5952);
and AND3 (N11998, N11988, N5761, N2578);
buf BUF1 (N11999, N11976);
or OR3 (N12000, N11994, N1012, N3971);
buf BUF1 (N12001, N11999);
nand NAND4 (N12002, N11996, N3507, N6701, N1845);
or OR4 (N12003, N11992, N5952, N6631, N43);
nand NAND3 (N12004, N11993, N10229, N4213);
or OR3 (N12005, N11991, N4248, N3970);
nor NOR3 (N12006, N12000, N4735, N500);
not NOT1 (N12007, N11981);
nor NOR4 (N12008, N12007, N1223, N10236, N7339);
buf BUF1 (N12009, N12001);
nor NOR4 (N12010, N11997, N6116, N5001, N518);
nor NOR4 (N12011, N12010, N1287, N2032, N10178);
nor NOR2 (N12012, N12003, N4256);
xor XOR2 (N12013, N12012, N2089);
nor NOR4 (N12014, N12006, N476, N10325, N10511);
or OR3 (N12015, N12005, N10886, N10902);
or OR4 (N12016, N11998, N3352, N2851, N10538);
buf BUF1 (N12017, N12009);
and AND3 (N12018, N12011, N1994, N4908);
buf BUF1 (N12019, N12016);
nor NOR2 (N12020, N12013, N1425);
buf BUF1 (N12021, N12002);
buf BUF1 (N12022, N12019);
or OR3 (N12023, N12014, N1365, N11741);
or OR4 (N12024, N12008, N9087, N7979, N2928);
or OR3 (N12025, N12018, N7024, N2775);
and AND3 (N12026, N12020, N8486, N9256);
and AND4 (N12027, N12022, N5690, N1070, N9604);
buf BUF1 (N12028, N12023);
nor NOR3 (N12029, N12004, N801, N5964);
nand NAND4 (N12030, N12021, N8371, N6441, N10681);
nand NAND3 (N12031, N12030, N8591, N8918);
or OR4 (N12032, N12028, N2918, N8089, N1324);
buf BUF1 (N12033, N12026);
xor XOR2 (N12034, N12024, N4267);
nand NAND2 (N12035, N12027, N4152);
nand NAND4 (N12036, N12025, N10202, N4225, N3482);
and AND3 (N12037, N12033, N2092, N2600);
nor NOR3 (N12038, N12015, N5134, N1517);
nor NOR3 (N12039, N12038, N9047, N7402);
or OR2 (N12040, N12036, N8360);
and AND3 (N12041, N12035, N9208, N5535);
and AND4 (N12042, N12032, N9607, N72, N10820);
nand NAND2 (N12043, N12037, N10962);
not NOT1 (N12044, N11984);
and AND3 (N12045, N12029, N11041, N9342);
nand NAND2 (N12046, N12039, N2209);
buf BUF1 (N12047, N12041);
xor XOR2 (N12048, N12046, N7141);
nand NAND3 (N12049, N12047, N11808, N4390);
nand NAND3 (N12050, N12031, N8680, N1037);
and AND2 (N12051, N12040, N8242);
nand NAND2 (N12052, N12017, N4352);
and AND3 (N12053, N12045, N9189, N5608);
buf BUF1 (N12054, N12053);
buf BUF1 (N12055, N12049);
not NOT1 (N12056, N12051);
not NOT1 (N12057, N12050);
xor XOR2 (N12058, N12034, N7951);
nand NAND3 (N12059, N12048, N7984, N5018);
buf BUF1 (N12060, N12055);
buf BUF1 (N12061, N12056);
not NOT1 (N12062, N12044);
nor NOR3 (N12063, N12043, N8207, N9636);
nor NOR4 (N12064, N12052, N6891, N10553, N405);
or OR4 (N12065, N12064, N10766, N3349, N8478);
and AND2 (N12066, N12059, N5467);
not NOT1 (N12067, N12061);
or OR3 (N12068, N12062, N7411, N6563);
nand NAND2 (N12069, N12068, N9209);
nand NAND4 (N12070, N12067, N9121, N3402, N2466);
nand NAND3 (N12071, N12066, N22, N1481);
buf BUF1 (N12072, N12071);
not NOT1 (N12073, N12060);
not NOT1 (N12074, N12063);
and AND2 (N12075, N12054, N1944);
not NOT1 (N12076, N12058);
and AND4 (N12077, N12075, N9330, N11725, N3657);
or OR2 (N12078, N12057, N6571);
not NOT1 (N12079, N12072);
or OR2 (N12080, N12073, N10031);
nand NAND2 (N12081, N12069, N855);
xor XOR2 (N12082, N12070, N4881);
not NOT1 (N12083, N12076);
nor NOR3 (N12084, N12042, N10944, N10130);
or OR4 (N12085, N12078, N12073, N812, N10963);
xor XOR2 (N12086, N12080, N12069);
nand NAND4 (N12087, N12085, N8131, N6601, N8176);
or OR3 (N12088, N12081, N1958, N7248);
and AND2 (N12089, N12079, N8935);
xor XOR2 (N12090, N12086, N9297);
and AND4 (N12091, N12082, N122, N6705, N88);
or OR4 (N12092, N12074, N10732, N4289, N5717);
not NOT1 (N12093, N12087);
and AND4 (N12094, N12091, N10984, N1362, N7337);
and AND3 (N12095, N12065, N1026, N9736);
xor XOR2 (N12096, N12093, N83);
nor NOR4 (N12097, N12089, N1608, N190, N3477);
xor XOR2 (N12098, N12094, N11758);
buf BUF1 (N12099, N12090);
not NOT1 (N12100, N12097);
nor NOR2 (N12101, N12077, N5012);
nor NOR3 (N12102, N12100, N5355, N11568);
or OR3 (N12103, N12083, N5382, N10151);
nor NOR3 (N12104, N12092, N1990, N9640);
nor NOR2 (N12105, N12099, N8163);
nor NOR2 (N12106, N12104, N4872);
or OR2 (N12107, N12095, N2553);
or OR3 (N12108, N12103, N8642, N3386);
and AND2 (N12109, N12098, N5883);
and AND4 (N12110, N12105, N10095, N7589, N7461);
buf BUF1 (N12111, N12109);
xor XOR2 (N12112, N12096, N5001);
or OR4 (N12113, N12110, N11849, N5329, N2814);
buf BUF1 (N12114, N12111);
buf BUF1 (N12115, N12106);
not NOT1 (N12116, N12084);
or OR2 (N12117, N12115, N5045);
nor NOR3 (N12118, N12113, N6077, N9846);
nor NOR3 (N12119, N12118, N10347, N2943);
nor NOR2 (N12120, N12116, N4411);
nand NAND4 (N12121, N12120, N3334, N9671, N3628);
or OR2 (N12122, N12101, N4130);
nand NAND4 (N12123, N12108, N4854, N5021, N2417);
nor NOR4 (N12124, N12122, N7641, N8910, N2948);
buf BUF1 (N12125, N12117);
xor XOR2 (N12126, N12125, N1377);
nand NAND2 (N12127, N12119, N11046);
nand NAND2 (N12128, N12112, N3858);
and AND2 (N12129, N12107, N4666);
nor NOR3 (N12130, N12088, N5312, N8483);
not NOT1 (N12131, N12130);
buf BUF1 (N12132, N12126);
nand NAND3 (N12133, N12123, N4023, N524);
not NOT1 (N12134, N12131);
buf BUF1 (N12135, N12114);
or OR2 (N12136, N12121, N6248);
xor XOR2 (N12137, N12133, N3419);
xor XOR2 (N12138, N12129, N2164);
buf BUF1 (N12139, N12132);
nor NOR3 (N12140, N12124, N6948, N5082);
not NOT1 (N12141, N12102);
and AND4 (N12142, N12141, N3332, N6396, N3384);
nor NOR3 (N12143, N12136, N4814, N3340);
not NOT1 (N12144, N12134);
or OR3 (N12145, N12139, N3099, N1248);
and AND4 (N12146, N12145, N2733, N11282, N1633);
and AND2 (N12147, N12135, N2631);
nor NOR2 (N12148, N12128, N9662);
buf BUF1 (N12149, N12138);
nor NOR4 (N12150, N12142, N4427, N7988, N9823);
and AND3 (N12151, N12144, N3780, N9464);
buf BUF1 (N12152, N12148);
and AND3 (N12153, N12140, N8699, N8484);
xor XOR2 (N12154, N12147, N10256);
xor XOR2 (N12155, N12151, N11576);
nor NOR3 (N12156, N12137, N7110, N5445);
buf BUF1 (N12157, N12155);
and AND2 (N12158, N12152, N813);
or OR3 (N12159, N12146, N2541, N5844);
xor XOR2 (N12160, N12150, N186);
nor NOR4 (N12161, N12156, N10271, N10411, N3205);
nor NOR2 (N12162, N12160, N9832);
nor NOR2 (N12163, N12162, N9673);
nand NAND2 (N12164, N12149, N9986);
nand NAND2 (N12165, N12157, N8757);
and AND4 (N12166, N12159, N7300, N5916, N4310);
and AND2 (N12167, N12166, N9137);
and AND3 (N12168, N12167, N4049, N5317);
not NOT1 (N12169, N12154);
not NOT1 (N12170, N12169);
nor NOR3 (N12171, N12170, N9892, N1698);
buf BUF1 (N12172, N12163);
xor XOR2 (N12173, N12158, N11874);
or OR4 (N12174, N12153, N5760, N8973, N9750);
buf BUF1 (N12175, N12165);
xor XOR2 (N12176, N12127, N6950);
or OR2 (N12177, N12175, N449);
or OR3 (N12178, N12174, N9400, N11663);
nand NAND3 (N12179, N12143, N4103, N7496);
not NOT1 (N12180, N12173);
nand NAND2 (N12181, N12176, N8725);
not NOT1 (N12182, N12177);
nor NOR2 (N12183, N12171, N933);
or OR2 (N12184, N12178, N3487);
nor NOR4 (N12185, N12183, N4916, N3573, N10976);
not NOT1 (N12186, N12164);
or OR3 (N12187, N12161, N351, N7483);
nand NAND4 (N12188, N12182, N8478, N3136, N9631);
not NOT1 (N12189, N12172);
buf BUF1 (N12190, N12189);
buf BUF1 (N12191, N12181);
or OR3 (N12192, N12188, N7579, N101);
nor NOR2 (N12193, N12190, N7287);
not NOT1 (N12194, N12185);
and AND4 (N12195, N12192, N2769, N2556, N4538);
xor XOR2 (N12196, N12180, N7630);
nor NOR2 (N12197, N12194, N850);
xor XOR2 (N12198, N12191, N1746);
buf BUF1 (N12199, N12196);
nand NAND2 (N12200, N12193, N10926);
xor XOR2 (N12201, N12184, N2200);
and AND3 (N12202, N12197, N6456, N422);
nor NOR2 (N12203, N12187, N10740);
buf BUF1 (N12204, N12199);
or OR2 (N12205, N12179, N4567);
xor XOR2 (N12206, N12186, N10182);
buf BUF1 (N12207, N12201);
nor NOR2 (N12208, N12207, N11078);
xor XOR2 (N12209, N12206, N2419);
xor XOR2 (N12210, N12209, N2853);
nor NOR2 (N12211, N12205, N7920);
nor NOR2 (N12212, N12203, N10678);
xor XOR2 (N12213, N12200, N8478);
and AND4 (N12214, N12202, N4309, N2291, N6072);
buf BUF1 (N12215, N12210);
nand NAND4 (N12216, N12212, N4874, N3617, N1969);
nand NAND3 (N12217, N12168, N8363, N3222);
nand NAND2 (N12218, N12216, N11979);
or OR2 (N12219, N12211, N8018);
and AND3 (N12220, N12204, N5640, N3079);
xor XOR2 (N12221, N12208, N187);
buf BUF1 (N12222, N12217);
buf BUF1 (N12223, N12220);
not NOT1 (N12224, N12195);
not NOT1 (N12225, N12218);
or OR3 (N12226, N12219, N2794, N5535);
not NOT1 (N12227, N12222);
not NOT1 (N12228, N12198);
xor XOR2 (N12229, N12226, N2857);
not NOT1 (N12230, N12215);
nand NAND3 (N12231, N12224, N5436, N34);
not NOT1 (N12232, N12223);
or OR3 (N12233, N12214, N7718, N1413);
or OR4 (N12234, N12233, N11748, N1259, N10542);
buf BUF1 (N12235, N12230);
and AND2 (N12236, N12213, N2897);
not NOT1 (N12237, N12227);
xor XOR2 (N12238, N12232, N1338);
nor NOR3 (N12239, N12237, N2680, N12137);
and AND2 (N12240, N12221, N1752);
and AND4 (N12241, N12229, N1524, N9159, N1240);
nand NAND2 (N12242, N12239, N1055);
nand NAND3 (N12243, N12238, N9505, N12029);
xor XOR2 (N12244, N12231, N9325);
nor NOR4 (N12245, N12241, N4475, N6688, N319);
xor XOR2 (N12246, N12236, N2635);
buf BUF1 (N12247, N12245);
and AND4 (N12248, N12235, N325, N11214, N6089);
buf BUF1 (N12249, N12246);
nor NOR4 (N12250, N12240, N4247, N2445, N6760);
xor XOR2 (N12251, N12250, N5784);
and AND2 (N12252, N12234, N11864);
xor XOR2 (N12253, N12252, N4840);
xor XOR2 (N12254, N12244, N1590);
xor XOR2 (N12255, N12253, N2153);
not NOT1 (N12256, N12248);
nor NOR2 (N12257, N12242, N2386);
and AND3 (N12258, N12249, N2209, N606);
nor NOR4 (N12259, N12228, N3131, N553, N11210);
not NOT1 (N12260, N12259);
buf BUF1 (N12261, N12260);
nor NOR3 (N12262, N12247, N5374, N4314);
nand NAND2 (N12263, N12255, N10202);
nor NOR3 (N12264, N12225, N11393, N44);
xor XOR2 (N12265, N12262, N7104);
or OR4 (N12266, N12264, N5205, N214, N11491);
and AND2 (N12267, N12256, N7523);
and AND3 (N12268, N12266, N146, N9265);
nand NAND3 (N12269, N12251, N2044, N6417);
buf BUF1 (N12270, N12269);
or OR2 (N12271, N12268, N11789);
xor XOR2 (N12272, N12261, N10262);
xor XOR2 (N12273, N12263, N5968);
or OR4 (N12274, N12267, N7198, N10591, N1483);
not NOT1 (N12275, N12243);
or OR4 (N12276, N12272, N3790, N1261, N8342);
nand NAND4 (N12277, N12270, N8011, N1602, N6460);
not NOT1 (N12278, N12254);
nand NAND3 (N12279, N12276, N7270, N2997);
xor XOR2 (N12280, N12279, N3345);
nor NOR4 (N12281, N12277, N11647, N7427, N2436);
nor NOR4 (N12282, N12257, N9778, N3158, N9221);
xor XOR2 (N12283, N12265, N4557);
nor NOR3 (N12284, N12278, N12158, N1910);
xor XOR2 (N12285, N12281, N7885);
nor NOR3 (N12286, N12282, N1158, N2008);
or OR4 (N12287, N12274, N5724, N3447, N11772);
not NOT1 (N12288, N12275);
nand NAND4 (N12289, N12273, N8046, N6976, N6819);
or OR2 (N12290, N12283, N11257);
and AND4 (N12291, N12289, N4938, N11050, N12019);
or OR3 (N12292, N12291, N6130, N409);
nor NOR4 (N12293, N12271, N6841, N1504, N5427);
buf BUF1 (N12294, N12258);
nor NOR4 (N12295, N12287, N1335, N8538, N429);
buf BUF1 (N12296, N12286);
or OR4 (N12297, N12292, N11100, N7264, N12271);
or OR3 (N12298, N12297, N5810, N7533);
or OR3 (N12299, N12294, N8936, N4215);
nand NAND3 (N12300, N12295, N11504, N8015);
nand NAND3 (N12301, N12296, N845, N2164);
xor XOR2 (N12302, N12285, N2061);
or OR2 (N12303, N12288, N529);
nand NAND2 (N12304, N12299, N12196);
not NOT1 (N12305, N12301);
or OR4 (N12306, N12293, N7725, N8950, N5018);
buf BUF1 (N12307, N12303);
buf BUF1 (N12308, N12298);
or OR4 (N12309, N12284, N8189, N3438, N3022);
not NOT1 (N12310, N12304);
xor XOR2 (N12311, N12307, N4302);
and AND3 (N12312, N12311, N5309, N6483);
and AND4 (N12313, N12300, N9802, N1585, N2129);
buf BUF1 (N12314, N12290);
nand NAND3 (N12315, N12310, N4795, N10067);
nor NOR2 (N12316, N12314, N10524);
buf BUF1 (N12317, N12306);
nor NOR4 (N12318, N12308, N3984, N8068, N4645);
nor NOR2 (N12319, N12302, N5099);
and AND4 (N12320, N12312, N4540, N4092, N7599);
buf BUF1 (N12321, N12315);
xor XOR2 (N12322, N12309, N3758);
xor XOR2 (N12323, N12316, N12083);
xor XOR2 (N12324, N12322, N11488);
or OR2 (N12325, N12318, N7414);
nand NAND2 (N12326, N12280, N8527);
and AND2 (N12327, N12326, N5121);
nand NAND2 (N12328, N12319, N4394);
or OR3 (N12329, N12328, N7153, N8226);
or OR2 (N12330, N12320, N10139);
or OR4 (N12331, N12329, N1775, N10885, N9269);
nand NAND3 (N12332, N12305, N3800, N5793);
nand NAND2 (N12333, N12323, N10228);
not NOT1 (N12334, N12325);
and AND3 (N12335, N12331, N9766, N9181);
and AND4 (N12336, N12327, N7651, N1687, N3604);
not NOT1 (N12337, N12321);
nor NOR3 (N12338, N12333, N3057, N6733);
or OR4 (N12339, N12336, N10576, N1581, N6857);
not NOT1 (N12340, N12332);
nand NAND2 (N12341, N12330, N3229);
xor XOR2 (N12342, N12324, N10525);
not NOT1 (N12343, N12334);
not NOT1 (N12344, N12340);
and AND4 (N12345, N12335, N604, N1938, N9947);
not NOT1 (N12346, N12341);
buf BUF1 (N12347, N12317);
xor XOR2 (N12348, N12346, N5781);
not NOT1 (N12349, N12347);
or OR4 (N12350, N12348, N12117, N995, N2460);
or OR3 (N12351, N12339, N12270, N9752);
nor NOR3 (N12352, N12351, N7718, N1395);
not NOT1 (N12353, N12350);
nor NOR3 (N12354, N12353, N6605, N8729);
or OR2 (N12355, N12344, N8241);
or OR3 (N12356, N12349, N3751, N6987);
and AND2 (N12357, N12342, N5674);
nand NAND2 (N12358, N12313, N4285);
or OR4 (N12359, N12358, N1296, N1127, N7055);
not NOT1 (N12360, N12359);
not NOT1 (N12361, N12360);
not NOT1 (N12362, N12352);
nand NAND3 (N12363, N12345, N2295, N8509);
nand NAND4 (N12364, N12354, N8485, N1591, N5490);
not NOT1 (N12365, N12361);
not NOT1 (N12366, N12362);
not NOT1 (N12367, N12337);
nand NAND4 (N12368, N12366, N9772, N11930, N877);
buf BUF1 (N12369, N12363);
and AND3 (N12370, N12364, N5876, N1626);
or OR3 (N12371, N12365, N2655, N440);
and AND2 (N12372, N12370, N9405);
and AND4 (N12373, N12368, N126, N454, N851);
xor XOR2 (N12374, N12372, N8623);
nor NOR3 (N12375, N12374, N12028, N11279);
nor NOR3 (N12376, N12369, N4592, N3918);
or OR3 (N12377, N12373, N3097, N8152);
nor NOR4 (N12378, N12357, N2485, N658, N5816);
nand NAND4 (N12379, N12343, N4448, N8063, N6177);
xor XOR2 (N12380, N12338, N8509);
not NOT1 (N12381, N12378);
and AND4 (N12382, N12371, N6051, N11722, N10663);
not NOT1 (N12383, N12355);
xor XOR2 (N12384, N12367, N5473);
not NOT1 (N12385, N12356);
nor NOR2 (N12386, N12379, N8113);
nor NOR2 (N12387, N12386, N7767);
not NOT1 (N12388, N12382);
and AND3 (N12389, N12381, N8417, N7822);
not NOT1 (N12390, N12376);
not NOT1 (N12391, N12387);
xor XOR2 (N12392, N12375, N5694);
xor XOR2 (N12393, N12389, N8045);
xor XOR2 (N12394, N12390, N2348);
not NOT1 (N12395, N12384);
not NOT1 (N12396, N12391);
and AND2 (N12397, N12392, N5843);
buf BUF1 (N12398, N12383);
not NOT1 (N12399, N12388);
and AND2 (N12400, N12380, N6374);
and AND4 (N12401, N12377, N7414, N12322, N5616);
and AND3 (N12402, N12396, N9767, N8144);
and AND2 (N12403, N12394, N85);
buf BUF1 (N12404, N12402);
nand NAND4 (N12405, N12395, N4099, N7712, N505);
nor NOR2 (N12406, N12398, N435);
and AND4 (N12407, N12401, N765, N10132, N7926);
xor XOR2 (N12408, N12397, N5082);
and AND3 (N12409, N12400, N6713, N9013);
nor NOR3 (N12410, N12404, N9026, N6020);
and AND2 (N12411, N12406, N10042);
and AND3 (N12412, N12399, N11750, N1557);
or OR2 (N12413, N12403, N12394);
and AND3 (N12414, N12393, N3980, N11329);
and AND2 (N12415, N12409, N9919);
not NOT1 (N12416, N12410);
or OR2 (N12417, N12405, N6674);
xor XOR2 (N12418, N12411, N8668);
nor NOR2 (N12419, N12408, N12064);
or OR2 (N12420, N12415, N7222);
not NOT1 (N12421, N12385);
nor NOR2 (N12422, N12416, N3250);
not NOT1 (N12423, N12412);
nor NOR2 (N12424, N12422, N1017);
xor XOR2 (N12425, N12414, N7152);
nor NOR4 (N12426, N12417, N7227, N9753, N6974);
not NOT1 (N12427, N12421);
nand NAND4 (N12428, N12423, N8143, N8929, N3990);
and AND4 (N12429, N12424, N1134, N10294, N7270);
and AND4 (N12430, N12418, N1191, N9713, N9284);
not NOT1 (N12431, N12420);
xor XOR2 (N12432, N12430, N11067);
nor NOR2 (N12433, N12413, N9351);
nand NAND3 (N12434, N12426, N12358, N10338);
xor XOR2 (N12435, N12428, N916);
nand NAND3 (N12436, N12419, N9062, N11626);
nand NAND3 (N12437, N12433, N939, N1584);
not NOT1 (N12438, N12432);
and AND4 (N12439, N12425, N8460, N4758, N480);
nand NAND2 (N12440, N12407, N8493);
nor NOR3 (N12441, N12435, N10744, N11371);
or OR3 (N12442, N12438, N6953, N3414);
nand NAND4 (N12443, N12439, N11138, N2884, N949);
and AND2 (N12444, N12443, N4674);
nor NOR4 (N12445, N12431, N1471, N9156, N7027);
nand NAND2 (N12446, N12442, N10940);
xor XOR2 (N12447, N12436, N3416);
and AND3 (N12448, N12446, N10308, N5440);
and AND2 (N12449, N12440, N767);
buf BUF1 (N12450, N12448);
nand NAND3 (N12451, N12437, N4689, N8996);
buf BUF1 (N12452, N12447);
and AND3 (N12453, N12449, N11110, N7012);
or OR2 (N12454, N12434, N2073);
nor NOR3 (N12455, N12427, N7500, N3808);
not NOT1 (N12456, N12451);
buf BUF1 (N12457, N12429);
buf BUF1 (N12458, N12444);
nand NAND3 (N12459, N12441, N9234, N1973);
or OR2 (N12460, N12445, N8170);
xor XOR2 (N12461, N12459, N8335);
or OR4 (N12462, N12460, N10989, N9457, N3485);
xor XOR2 (N12463, N12453, N1923);
nand NAND3 (N12464, N12463, N2501, N8911);
or OR2 (N12465, N12450, N2347);
nand NAND2 (N12466, N12464, N5939);
buf BUF1 (N12467, N12452);
or OR3 (N12468, N12455, N9182, N11012);
nand NAND3 (N12469, N12458, N3527, N8283);
nor NOR2 (N12470, N12469, N12048);
nand NAND3 (N12471, N12466, N6317, N663);
nand NAND2 (N12472, N12465, N9593);
not NOT1 (N12473, N12462);
or OR2 (N12474, N12467, N3522);
nand NAND4 (N12475, N12474, N4087, N252, N10215);
or OR4 (N12476, N12461, N7783, N2268, N11297);
xor XOR2 (N12477, N12475, N11848);
nor NOR2 (N12478, N12471, N11824);
and AND2 (N12479, N12476, N12079);
and AND4 (N12480, N12477, N234, N6986, N7916);
nor NOR2 (N12481, N12473, N2021);
and AND2 (N12482, N12481, N1525);
and AND2 (N12483, N12454, N6139);
buf BUF1 (N12484, N12482);
nor NOR2 (N12485, N12478, N8547);
or OR4 (N12486, N12472, N9248, N7546, N9870);
buf BUF1 (N12487, N12485);
and AND4 (N12488, N12457, N5743, N10526, N7940);
xor XOR2 (N12489, N12484, N9261);
not NOT1 (N12490, N12470);
nor NOR4 (N12491, N12486, N11794, N409, N3345);
and AND4 (N12492, N12479, N11361, N1558, N10694);
buf BUF1 (N12493, N12489);
or OR2 (N12494, N12493, N8004);
xor XOR2 (N12495, N12487, N11857);
not NOT1 (N12496, N12492);
nand NAND4 (N12497, N12483, N349, N3751, N9497);
nand NAND4 (N12498, N12491, N6994, N8614, N2973);
nand NAND3 (N12499, N12495, N5789, N8600);
nand NAND3 (N12500, N12496, N1797, N1669);
and AND4 (N12501, N12468, N11622, N12152, N4816);
nor NOR2 (N12502, N12499, N7039);
and AND3 (N12503, N12480, N7064, N5903);
nor NOR4 (N12504, N12498, N8804, N5794, N6628);
not NOT1 (N12505, N12504);
buf BUF1 (N12506, N12494);
not NOT1 (N12507, N12490);
buf BUF1 (N12508, N12501);
xor XOR2 (N12509, N12497, N2588);
not NOT1 (N12510, N12503);
not NOT1 (N12511, N12502);
or OR3 (N12512, N12507, N3309, N866);
nor NOR4 (N12513, N12511, N11400, N6266, N875);
xor XOR2 (N12514, N12510, N7677);
nor NOR2 (N12515, N12512, N5490);
nor NOR2 (N12516, N12508, N5826);
and AND2 (N12517, N12515, N7185);
not NOT1 (N12518, N12513);
nand NAND3 (N12519, N12500, N5936, N3174);
not NOT1 (N12520, N12514);
or OR3 (N12521, N12506, N10552, N8171);
nand NAND2 (N12522, N12509, N10805);
xor XOR2 (N12523, N12519, N8407);
nand NAND3 (N12524, N12516, N4796, N8887);
xor XOR2 (N12525, N12505, N5217);
or OR4 (N12526, N12517, N2916, N10275, N12019);
nand NAND2 (N12527, N12488, N9914);
nand NAND2 (N12528, N12523, N7269);
xor XOR2 (N12529, N12528, N3492);
buf BUF1 (N12530, N12527);
nand NAND2 (N12531, N12518, N2286);
xor XOR2 (N12532, N12526, N6787);
not NOT1 (N12533, N12522);
nor NOR4 (N12534, N12530, N1972, N3567, N4986);
or OR4 (N12535, N12531, N6530, N11072, N10970);
or OR2 (N12536, N12521, N9619);
buf BUF1 (N12537, N12535);
buf BUF1 (N12538, N12537);
nor NOR3 (N12539, N12456, N9544, N7028);
or OR3 (N12540, N12525, N7916, N7346);
or OR3 (N12541, N12533, N3158, N9756);
nand NAND4 (N12542, N12534, N2440, N5800, N1403);
buf BUF1 (N12543, N12542);
nor NOR3 (N12544, N12524, N646, N3894);
nor NOR2 (N12545, N12543, N8641);
not NOT1 (N12546, N12538);
buf BUF1 (N12547, N12539);
buf BUF1 (N12548, N12520);
nand NAND3 (N12549, N12546, N12116, N5134);
or OR4 (N12550, N12536, N6070, N9208, N5238);
nand NAND2 (N12551, N12529, N2974);
or OR3 (N12552, N12550, N3228, N4987);
or OR4 (N12553, N12547, N1627, N7354, N1236);
nand NAND4 (N12554, N12551, N5512, N6294, N8999);
buf BUF1 (N12555, N12554);
buf BUF1 (N12556, N12553);
nor NOR4 (N12557, N12556, N11558, N9925, N11701);
or OR4 (N12558, N12541, N11774, N8196, N10150);
nor NOR4 (N12559, N12552, N2969, N9747, N3813);
nor NOR2 (N12560, N12544, N8437);
nor NOR3 (N12561, N12549, N10836, N6967);
and AND4 (N12562, N12532, N2962, N11922, N3643);
buf BUF1 (N12563, N12562);
nand NAND2 (N12564, N12557, N8042);
buf BUF1 (N12565, N12540);
or OR4 (N12566, N12559, N5761, N12247, N7437);
or OR3 (N12567, N12558, N7918, N8672);
nand NAND2 (N12568, N12555, N4403);
xor XOR2 (N12569, N12567, N10936);
buf BUF1 (N12570, N12568);
nor NOR4 (N12571, N12561, N1808, N9597, N1519);
not NOT1 (N12572, N12565);
nor NOR3 (N12573, N12571, N11238, N12141);
not NOT1 (N12574, N12572);
xor XOR2 (N12575, N12564, N10526);
nor NOR3 (N12576, N12566, N11732, N1649);
and AND3 (N12577, N12574, N812, N1882);
buf BUF1 (N12578, N12560);
nor NOR2 (N12579, N12575, N3623);
not NOT1 (N12580, N12569);
not NOT1 (N12581, N12579);
nand NAND2 (N12582, N12580, N5333);
or OR3 (N12583, N12545, N5148, N10196);
xor XOR2 (N12584, N12548, N2118);
or OR4 (N12585, N12573, N5322, N11645, N10542);
not NOT1 (N12586, N12578);
nor NOR3 (N12587, N12584, N3548, N2064);
xor XOR2 (N12588, N12576, N4322);
buf BUF1 (N12589, N12581);
buf BUF1 (N12590, N12589);
or OR3 (N12591, N12577, N11970, N8870);
nor NOR4 (N12592, N12588, N2044, N7963, N5549);
or OR2 (N12593, N12585, N9538);
and AND2 (N12594, N12587, N7173);
buf BUF1 (N12595, N12594);
nor NOR2 (N12596, N12586, N10415);
buf BUF1 (N12597, N12582);
nand NAND4 (N12598, N12593, N4331, N12595, N1514);
and AND2 (N12599, N379, N7353);
buf BUF1 (N12600, N12570);
nor NOR2 (N12601, N12598, N12007);
and AND3 (N12602, N12599, N4244, N3977);
not NOT1 (N12603, N12590);
and AND4 (N12604, N12592, N2814, N5317, N10601);
nand NAND3 (N12605, N12601, N2766, N8934);
nand NAND2 (N12606, N12605, N2169);
and AND4 (N12607, N12563, N8358, N506, N5032);
not NOT1 (N12608, N12597);
nand NAND2 (N12609, N12591, N11599);
nand NAND4 (N12610, N12603, N10395, N6339, N4969);
and AND2 (N12611, N12604, N12127);
xor XOR2 (N12612, N12583, N4847);
xor XOR2 (N12613, N12608, N3285);
not NOT1 (N12614, N12611);
and AND3 (N12615, N12602, N4662, N11547);
nor NOR2 (N12616, N12614, N8079);
not NOT1 (N12617, N12615);
not NOT1 (N12618, N12612);
xor XOR2 (N12619, N12610, N5307);
nor NOR3 (N12620, N12609, N11376, N9389);
nand NAND3 (N12621, N12618, N9093, N9214);
xor XOR2 (N12622, N12621, N2433);
nor NOR4 (N12623, N12600, N7492, N6941, N5526);
buf BUF1 (N12624, N12607);
and AND2 (N12625, N12606, N7980);
or OR4 (N12626, N12616, N5719, N5798, N24);
nor NOR2 (N12627, N12617, N6672);
nand NAND3 (N12628, N12613, N3161, N10609);
nor NOR4 (N12629, N12619, N8352, N4992, N5376);
xor XOR2 (N12630, N12625, N2929);
not NOT1 (N12631, N12624);
and AND4 (N12632, N12628, N3362, N11198, N9145);
or OR3 (N12633, N12631, N11929, N8696);
xor XOR2 (N12634, N12630, N12450);
not NOT1 (N12635, N12596);
buf BUF1 (N12636, N12634);
or OR2 (N12637, N12632, N2900);
and AND3 (N12638, N12636, N7438, N11558);
or OR4 (N12639, N12629, N6518, N2596, N5883);
buf BUF1 (N12640, N12638);
and AND3 (N12641, N12623, N2772, N2958);
buf BUF1 (N12642, N12627);
and AND4 (N12643, N12620, N1634, N2031, N2102);
buf BUF1 (N12644, N12639);
and AND4 (N12645, N12643, N238, N7541, N1680);
buf BUF1 (N12646, N12633);
nand NAND2 (N12647, N12637, N2265);
xor XOR2 (N12648, N12647, N103);
nor NOR3 (N12649, N12640, N6154, N3681);
xor XOR2 (N12650, N12635, N9365);
and AND4 (N12651, N12644, N6683, N10806, N5481);
and AND3 (N12652, N12649, N2051, N141);
or OR2 (N12653, N12651, N4595);
nand NAND2 (N12654, N12645, N3573);
xor XOR2 (N12655, N12642, N3016);
nand NAND4 (N12656, N12641, N4332, N4344, N6389);
xor XOR2 (N12657, N12653, N6874);
xor XOR2 (N12658, N12656, N8583);
or OR3 (N12659, N12652, N12240, N10175);
buf BUF1 (N12660, N12648);
not NOT1 (N12661, N12626);
buf BUF1 (N12662, N12622);
or OR3 (N12663, N12657, N12012, N7430);
nor NOR4 (N12664, N12650, N6081, N5709, N8555);
and AND3 (N12665, N12662, N10711, N8634);
not NOT1 (N12666, N12665);
buf BUF1 (N12667, N12646);
xor XOR2 (N12668, N12664, N10074);
nor NOR2 (N12669, N12668, N11979);
not NOT1 (N12670, N12655);
nand NAND2 (N12671, N12663, N3411);
xor XOR2 (N12672, N12671, N11422);
nand NAND2 (N12673, N12658, N10259);
nand NAND2 (N12674, N12669, N10188);
buf BUF1 (N12675, N12660);
or OR3 (N12676, N12666, N1194, N7881);
not NOT1 (N12677, N12675);
xor XOR2 (N12678, N12677, N10167);
nand NAND2 (N12679, N12674, N4228);
or OR2 (N12680, N12661, N5883);
not NOT1 (N12681, N12659);
and AND4 (N12682, N12654, N9295, N2163, N2430);
nor NOR2 (N12683, N12682, N3943);
buf BUF1 (N12684, N12676);
or OR3 (N12685, N12683, N6362, N1343);
nor NOR4 (N12686, N12678, N7835, N10606, N221);
or OR3 (N12687, N12667, N9941, N11693);
nor NOR2 (N12688, N12679, N365);
nand NAND3 (N12689, N12680, N1010, N9946);
xor XOR2 (N12690, N12681, N8110);
buf BUF1 (N12691, N12673);
nand NAND2 (N12692, N12690, N5629);
nor NOR2 (N12693, N12686, N2120);
and AND2 (N12694, N12689, N8387);
and AND4 (N12695, N12685, N4487, N1951, N11296);
nor NOR3 (N12696, N12672, N9850, N10987);
or OR4 (N12697, N12687, N951, N12505, N11363);
nand NAND3 (N12698, N12695, N11719, N12430);
not NOT1 (N12699, N12693);
nor NOR2 (N12700, N12694, N2526);
nor NOR4 (N12701, N12691, N8294, N2004, N3103);
nand NAND2 (N12702, N12692, N4238);
xor XOR2 (N12703, N12688, N5544);
buf BUF1 (N12704, N12684);
xor XOR2 (N12705, N12704, N5313);
buf BUF1 (N12706, N12701);
xor XOR2 (N12707, N12670, N802);
nand NAND4 (N12708, N12707, N1255, N6645, N7100);
not NOT1 (N12709, N12696);
and AND2 (N12710, N12697, N12523);
buf BUF1 (N12711, N12706);
and AND2 (N12712, N12700, N218);
and AND4 (N12713, N12705, N9150, N4136, N11707);
buf BUF1 (N12714, N12709);
not NOT1 (N12715, N12708);
nor NOR3 (N12716, N12714, N204, N10650);
or OR4 (N12717, N12711, N4966, N5750, N2804);
buf BUF1 (N12718, N12713);
buf BUF1 (N12719, N12698);
xor XOR2 (N12720, N12715, N1483);
not NOT1 (N12721, N12720);
xor XOR2 (N12722, N12712, N10552);
or OR2 (N12723, N12719, N9705);
not NOT1 (N12724, N12722);
nor NOR2 (N12725, N12703, N1115);
or OR4 (N12726, N12723, N5363, N2451, N5667);
or OR2 (N12727, N12721, N7492);
and AND3 (N12728, N12718, N10069, N5263);
nor NOR2 (N12729, N12727, N9109);
xor XOR2 (N12730, N12699, N4121);
not NOT1 (N12731, N12710);
nor NOR3 (N12732, N12717, N8622, N4593);
nor NOR3 (N12733, N12726, N3093, N9395);
nand NAND3 (N12734, N12730, N6889, N5783);
not NOT1 (N12735, N12733);
not NOT1 (N12736, N12728);
xor XOR2 (N12737, N12734, N4694);
and AND3 (N12738, N12737, N788, N4497);
nor NOR4 (N12739, N12736, N5588, N6463, N9911);
xor XOR2 (N12740, N12729, N6874);
not NOT1 (N12741, N12740);
nor NOR4 (N12742, N12702, N9837, N4624, N9445);
buf BUF1 (N12743, N12732);
not NOT1 (N12744, N12742);
xor XOR2 (N12745, N12743, N4882);
buf BUF1 (N12746, N12731);
nand NAND3 (N12747, N12741, N11335, N10644);
not NOT1 (N12748, N12725);
xor XOR2 (N12749, N12744, N4054);
nor NOR4 (N12750, N12738, N2195, N10600, N10688);
buf BUF1 (N12751, N12735);
or OR4 (N12752, N12716, N9654, N8993, N10713);
and AND3 (N12753, N12748, N4895, N1370);
nor NOR4 (N12754, N12724, N7076, N12370, N3479);
buf BUF1 (N12755, N12751);
and AND2 (N12756, N12752, N11284);
not NOT1 (N12757, N12739);
or OR4 (N12758, N12745, N12436, N8537, N138);
or OR2 (N12759, N12757, N3039);
not NOT1 (N12760, N12759);
nor NOR4 (N12761, N12756, N8393, N12424, N3044);
xor XOR2 (N12762, N12750, N10363);
nand NAND4 (N12763, N12747, N2077, N2698, N10976);
not NOT1 (N12764, N12746);
buf BUF1 (N12765, N12749);
nor NOR2 (N12766, N12758, N12287);
nor NOR4 (N12767, N12766, N8355, N11452, N1272);
buf BUF1 (N12768, N12765);
nor NOR4 (N12769, N12768, N11207, N6116, N6189);
and AND3 (N12770, N12754, N10879, N339);
xor XOR2 (N12771, N12769, N3042);
nor NOR4 (N12772, N12761, N12364, N3162, N4228);
xor XOR2 (N12773, N12760, N5724);
or OR4 (N12774, N12771, N878, N11956, N4583);
and AND2 (N12775, N12772, N7326);
nor NOR4 (N12776, N12774, N1352, N831, N8468);
buf BUF1 (N12777, N12770);
nor NOR4 (N12778, N12755, N399, N1528, N4893);
nor NOR3 (N12779, N12764, N1763, N1376);
not NOT1 (N12780, N12773);
buf BUF1 (N12781, N12763);
xor XOR2 (N12782, N12762, N2891);
buf BUF1 (N12783, N12777);
and AND4 (N12784, N12780, N5907, N12653, N6648);
nand NAND4 (N12785, N12776, N1780, N6803, N7907);
buf BUF1 (N12786, N12779);
and AND2 (N12787, N12784, N4859);
not NOT1 (N12788, N12767);
buf BUF1 (N12789, N12787);
buf BUF1 (N12790, N12778);
and AND4 (N12791, N12781, N10670, N9156, N11748);
or OR4 (N12792, N12790, N8447, N9449, N5675);
nor NOR4 (N12793, N12775, N2746, N6201, N7748);
and AND3 (N12794, N12792, N6162, N10611);
xor XOR2 (N12795, N12789, N1435);
or OR3 (N12796, N12785, N7291, N6138);
xor XOR2 (N12797, N12791, N8937);
nand NAND2 (N12798, N12786, N9656);
not NOT1 (N12799, N12796);
nor NOR2 (N12800, N12794, N11940);
nor NOR3 (N12801, N12797, N10679, N359);
nor NOR4 (N12802, N12782, N3221, N606, N10253);
xor XOR2 (N12803, N12795, N8038);
buf BUF1 (N12804, N12783);
or OR4 (N12805, N12793, N8742, N4084, N12387);
nand NAND3 (N12806, N12800, N3228, N8146);
not NOT1 (N12807, N12802);
nor NOR2 (N12808, N12801, N10399);
buf BUF1 (N12809, N12753);
not NOT1 (N12810, N12804);
buf BUF1 (N12811, N12805);
buf BUF1 (N12812, N12807);
xor XOR2 (N12813, N12799, N2931);
or OR4 (N12814, N12811, N5655, N7030, N3160);
not NOT1 (N12815, N12806);
buf BUF1 (N12816, N12803);
nor NOR3 (N12817, N12809, N4846, N11087);
nand NAND3 (N12818, N12815, N12232, N8013);
endmodule