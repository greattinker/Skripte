// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N1512,N1483,N1511,N1506,N1502,N1505,N1510,N1508,N1495,N1513;

buf BUF1 (N14, N5);
and AND2 (N15, N14, N13);
not NOT1 (N16, N13);
nand NAND4 (N17, N5, N6, N13, N13);
buf BUF1 (N18, N16);
nor NOR4 (N19, N18, N6, N16, N8);
xor XOR2 (N20, N8, N17);
xor XOR2 (N21, N12, N19);
and AND2 (N22, N12, N16);
buf BUF1 (N23, N5);
nand NAND4 (N24, N8, N8, N8, N19);
and AND3 (N25, N7, N13, N6);
nand NAND4 (N26, N20, N2, N24, N19);
or OR2 (N27, N7, N24);
or OR2 (N28, N6, N24);
nand NAND4 (N29, N22, N28, N4, N2);
buf BUF1 (N30, N29);
or OR2 (N31, N21, N28);
and AND3 (N32, N16, N27, N18);
nand NAND3 (N33, N21, N26, N26);
not NOT1 (N34, N1);
nor NOR3 (N35, N6, N28, N4);
xor XOR2 (N36, N17, N31);
or OR2 (N37, N35, N22);
nand NAND4 (N38, N9, N37, N17, N4);
nor NOR2 (N39, N31, N12);
nor NOR3 (N40, N23, N12, N11);
not NOT1 (N41, N39);
or OR4 (N42, N34, N5, N5, N29);
or OR4 (N43, N41, N8, N31, N10);
buf BUF1 (N44, N36);
and AND2 (N45, N30, N28);
nand NAND2 (N46, N43, N6);
or OR3 (N47, N15, N22, N7);
xor XOR2 (N48, N40, N6);
nor NOR4 (N49, N25, N39, N35, N33);
not NOT1 (N50, N38);
xor XOR2 (N51, N25, N47);
nor NOR2 (N52, N12, N29);
xor XOR2 (N53, N45, N39);
and AND4 (N54, N52, N33, N17, N46);
nor NOR3 (N55, N4, N26, N42);
or OR2 (N56, N36, N2);
nand NAND3 (N57, N44, N15, N22);
or OR3 (N58, N50, N18, N53);
buf BUF1 (N59, N57);
nor NOR2 (N60, N29, N23);
nor NOR2 (N61, N49, N21);
xor XOR2 (N62, N55, N6);
and AND2 (N63, N32, N47);
and AND3 (N64, N59, N39, N14);
nor NOR2 (N65, N63, N7);
nand NAND3 (N66, N54, N3, N21);
nor NOR4 (N67, N65, N22, N14, N24);
nor NOR2 (N68, N58, N35);
not NOT1 (N69, N66);
or OR2 (N70, N56, N66);
nor NOR2 (N71, N64, N4);
not NOT1 (N72, N70);
nand NAND4 (N73, N69, N63, N19, N21);
nand NAND4 (N74, N61, N37, N24, N62);
not NOT1 (N75, N47);
not NOT1 (N76, N68);
nand NAND3 (N77, N74, N41, N57);
and AND3 (N78, N72, N19, N17);
and AND3 (N79, N71, N48, N7);
nand NAND4 (N80, N7, N58, N19, N58);
or OR2 (N81, N60, N23);
buf BUF1 (N82, N81);
nand NAND4 (N83, N80, N46, N54, N8);
not NOT1 (N84, N73);
not NOT1 (N85, N83);
not NOT1 (N86, N67);
nand NAND2 (N87, N86, N55);
nor NOR4 (N88, N75, N44, N61, N72);
nor NOR2 (N89, N78, N18);
xor XOR2 (N90, N85, N60);
nor NOR2 (N91, N90, N58);
buf BUF1 (N92, N77);
nand NAND3 (N93, N89, N24, N81);
buf BUF1 (N94, N91);
or OR3 (N95, N87, N64, N92);
buf BUF1 (N96, N35);
or OR2 (N97, N51, N41);
buf BUF1 (N98, N96);
nand NAND4 (N99, N82, N94, N81, N60);
xor XOR2 (N100, N86, N24);
nand NAND2 (N101, N99, N72);
xor XOR2 (N102, N88, N69);
nand NAND3 (N103, N95, N69, N74);
not NOT1 (N104, N97);
xor XOR2 (N105, N98, N15);
nand NAND4 (N106, N100, N101, N88, N38);
and AND2 (N107, N60, N97);
xor XOR2 (N108, N102, N69);
and AND4 (N109, N107, N59, N79, N49);
not NOT1 (N110, N18);
nor NOR4 (N111, N76, N107, N110, N48);
not NOT1 (N112, N92);
xor XOR2 (N113, N111, N50);
nor NOR2 (N114, N112, N16);
nand NAND2 (N115, N84, N84);
nor NOR3 (N116, N105, N68, N35);
not NOT1 (N117, N116);
buf BUF1 (N118, N106);
buf BUF1 (N119, N93);
nand NAND3 (N120, N113, N83, N70);
and AND2 (N121, N103, N15);
or OR3 (N122, N121, N31, N85);
nand NAND3 (N123, N109, N81, N71);
nand NAND4 (N124, N123, N87, N35, N91);
nand NAND2 (N125, N118, N59);
not NOT1 (N126, N117);
or OR2 (N127, N126, N49);
nand NAND4 (N128, N125, N126, N111, N94);
xor XOR2 (N129, N115, N76);
xor XOR2 (N130, N108, N44);
buf BUF1 (N131, N128);
or OR3 (N132, N114, N34, N12);
nand NAND4 (N133, N120, N104, N3, N37);
nand NAND4 (N134, N109, N82, N42, N73);
and AND3 (N135, N134, N121, N9);
or OR2 (N136, N131, N20);
buf BUF1 (N137, N136);
nor NOR2 (N138, N130, N92);
and AND2 (N139, N135, N31);
xor XOR2 (N140, N122, N59);
nor NOR4 (N141, N133, N103, N16, N8);
nor NOR4 (N142, N119, N113, N21, N56);
nor NOR3 (N143, N132, N107, N86);
and AND2 (N144, N129, N52);
nor NOR3 (N145, N142, N47, N32);
xor XOR2 (N146, N143, N12);
not NOT1 (N147, N145);
and AND4 (N148, N147, N98, N134, N88);
and AND3 (N149, N127, N12, N99);
and AND4 (N150, N138, N123, N132, N11);
not NOT1 (N151, N149);
nor NOR2 (N152, N144, N111);
nand NAND3 (N153, N141, N50, N47);
nand NAND4 (N154, N153, N105, N73, N25);
xor XOR2 (N155, N140, N134);
xor XOR2 (N156, N155, N61);
xor XOR2 (N157, N146, N1);
nor NOR3 (N158, N152, N123, N114);
or OR4 (N159, N157, N81, N33, N46);
xor XOR2 (N160, N156, N123);
nor NOR2 (N161, N158, N41);
buf BUF1 (N162, N137);
or OR4 (N163, N148, N152, N35, N108);
nand NAND3 (N164, N160, N34, N64);
not NOT1 (N165, N159);
and AND3 (N166, N139, N146, N64);
nor NOR4 (N167, N150, N37, N142, N155);
nor NOR4 (N168, N163, N97, N57, N140);
not NOT1 (N169, N161);
nor NOR2 (N170, N154, N84);
xor XOR2 (N171, N162, N9);
and AND3 (N172, N168, N117, N135);
buf BUF1 (N173, N169);
xor XOR2 (N174, N170, N76);
and AND2 (N175, N164, N149);
xor XOR2 (N176, N151, N79);
not NOT1 (N177, N167);
xor XOR2 (N178, N176, N147);
or OR3 (N179, N172, N85, N72);
buf BUF1 (N180, N166);
nor NOR2 (N181, N179, N75);
buf BUF1 (N182, N180);
nand NAND3 (N183, N171, N45, N15);
or OR2 (N184, N183, N115);
buf BUF1 (N185, N165);
buf BUF1 (N186, N185);
xor XOR2 (N187, N175, N143);
and AND3 (N188, N174, N170, N43);
nand NAND3 (N189, N177, N155, N159);
nor NOR3 (N190, N173, N71, N118);
not NOT1 (N191, N182);
buf BUF1 (N192, N178);
nor NOR4 (N193, N190, N127, N8, N147);
nand NAND2 (N194, N184, N87);
and AND3 (N195, N188, N136, N174);
or OR2 (N196, N186, N113);
not NOT1 (N197, N192);
buf BUF1 (N198, N191);
xor XOR2 (N199, N194, N88);
and AND4 (N200, N198, N102, N30, N60);
not NOT1 (N201, N195);
nor NOR3 (N202, N193, N64, N96);
nor NOR4 (N203, N189, N186, N148, N101);
xor XOR2 (N204, N202, N100);
nand NAND3 (N205, N181, N160, N199);
nor NOR2 (N206, N15, N119);
and AND2 (N207, N187, N70);
nand NAND4 (N208, N201, N19, N167, N159);
buf BUF1 (N209, N205);
not NOT1 (N210, N124);
buf BUF1 (N211, N203);
and AND3 (N212, N196, N167, N29);
or OR2 (N213, N209, N59);
xor XOR2 (N214, N212, N115);
buf BUF1 (N215, N214);
xor XOR2 (N216, N207, N56);
buf BUF1 (N217, N200);
or OR4 (N218, N208, N112, N170, N32);
not NOT1 (N219, N216);
buf BUF1 (N220, N219);
and AND4 (N221, N210, N19, N164, N139);
xor XOR2 (N222, N197, N104);
and AND4 (N223, N221, N99, N103, N94);
not NOT1 (N224, N222);
buf BUF1 (N225, N211);
or OR3 (N226, N217, N184, N103);
nand NAND4 (N227, N226, N52, N7, N18);
nand NAND4 (N228, N220, N86, N174, N139);
and AND4 (N229, N223, N216, N100, N169);
nor NOR4 (N230, N215, N4, N139, N124);
nand NAND4 (N231, N218, N56, N71, N220);
not NOT1 (N232, N224);
nand NAND2 (N233, N232, N203);
and AND4 (N234, N213, N114, N110, N170);
xor XOR2 (N235, N204, N58);
not NOT1 (N236, N227);
nand NAND3 (N237, N206, N3, N127);
and AND2 (N238, N234, N69);
xor XOR2 (N239, N229, N220);
xor XOR2 (N240, N225, N47);
buf BUF1 (N241, N238);
xor XOR2 (N242, N241, N147);
buf BUF1 (N243, N235);
buf BUF1 (N244, N228);
or OR3 (N245, N236, N65, N32);
or OR2 (N246, N239, N22);
xor XOR2 (N247, N246, N236);
and AND4 (N248, N233, N169, N42, N126);
xor XOR2 (N249, N230, N133);
xor XOR2 (N250, N231, N190);
not NOT1 (N251, N237);
and AND4 (N252, N240, N98, N124, N85);
nor NOR2 (N253, N244, N97);
or OR2 (N254, N249, N44);
nand NAND2 (N255, N250, N22);
not NOT1 (N256, N243);
or OR3 (N257, N253, N90, N116);
nand NAND2 (N258, N257, N26);
nand NAND4 (N259, N258, N127, N220, N157);
or OR2 (N260, N245, N105);
not NOT1 (N261, N252);
buf BUF1 (N262, N259);
xor XOR2 (N263, N262, N235);
or OR4 (N264, N260, N255, N75, N95);
xor XOR2 (N265, N213, N100);
or OR2 (N266, N256, N2);
nand NAND2 (N267, N266, N30);
xor XOR2 (N268, N247, N241);
buf BUF1 (N269, N251);
nand NAND2 (N270, N269, N226);
or OR2 (N271, N270, N157);
and AND2 (N272, N267, N86);
nor NOR3 (N273, N263, N178, N57);
or OR4 (N274, N242, N203, N130, N152);
xor XOR2 (N275, N268, N54);
or OR2 (N276, N275, N181);
xor XOR2 (N277, N273, N91);
not NOT1 (N278, N265);
buf BUF1 (N279, N278);
xor XOR2 (N280, N277, N45);
not NOT1 (N281, N261);
buf BUF1 (N282, N271);
nand NAND3 (N283, N280, N123, N20);
and AND2 (N284, N264, N176);
not NOT1 (N285, N276);
nand NAND3 (N286, N284, N174, N191);
not NOT1 (N287, N281);
nand NAND3 (N288, N248, N278, N90);
buf BUF1 (N289, N288);
buf BUF1 (N290, N286);
nor NOR2 (N291, N283, N279);
not NOT1 (N292, N7);
and AND4 (N293, N290, N14, N123, N86);
nor NOR3 (N294, N285, N84, N67);
xor XOR2 (N295, N294, N132);
buf BUF1 (N296, N292);
and AND4 (N297, N296, N87, N2, N195);
or OR3 (N298, N291, N4, N38);
or OR2 (N299, N272, N223);
nor NOR2 (N300, N274, N199);
nor NOR3 (N301, N300, N225, N61);
and AND3 (N302, N254, N294, N230);
or OR4 (N303, N297, N263, N73, N276);
and AND2 (N304, N287, N172);
not NOT1 (N305, N295);
nor NOR4 (N306, N289, N152, N215, N166);
not NOT1 (N307, N306);
nor NOR3 (N308, N303, N27, N236);
not NOT1 (N309, N308);
buf BUF1 (N310, N309);
nand NAND4 (N311, N310, N278, N279, N209);
not NOT1 (N312, N304);
xor XOR2 (N313, N307, N73);
nand NAND3 (N314, N312, N115, N116);
nor NOR3 (N315, N299, N52, N170);
xor XOR2 (N316, N282, N69);
or OR4 (N317, N301, N117, N37, N307);
buf BUF1 (N318, N305);
and AND3 (N319, N314, N174, N272);
and AND4 (N320, N302, N82, N214, N184);
nand NAND2 (N321, N298, N248);
buf BUF1 (N322, N293);
buf BUF1 (N323, N313);
or OR4 (N324, N315, N277, N32, N269);
nand NAND4 (N325, N321, N228, N199, N40);
nor NOR4 (N326, N323, N234, N6, N3);
and AND3 (N327, N317, N293, N67);
buf BUF1 (N328, N326);
nor NOR4 (N329, N319, N187, N2, N42);
xor XOR2 (N330, N328, N319);
xor XOR2 (N331, N311, N67);
xor XOR2 (N332, N320, N285);
buf BUF1 (N333, N331);
nor NOR4 (N334, N322, N189, N202, N21);
and AND4 (N335, N324, N48, N143, N7);
and AND2 (N336, N325, N160);
not NOT1 (N337, N329);
nor NOR2 (N338, N337, N97);
buf BUF1 (N339, N330);
or OR3 (N340, N338, N101, N65);
nand NAND3 (N341, N339, N176, N306);
nand NAND4 (N342, N333, N282, N97, N140);
xor XOR2 (N343, N316, N39);
and AND4 (N344, N327, N230, N20, N177);
nor NOR2 (N345, N332, N106);
not NOT1 (N346, N318);
nor NOR3 (N347, N346, N62, N346);
nand NAND4 (N348, N347, N340, N117, N117);
nand NAND2 (N349, N300, N316);
buf BUF1 (N350, N343);
or OR2 (N351, N341, N314);
buf BUF1 (N352, N348);
buf BUF1 (N353, N335);
not NOT1 (N354, N352);
and AND3 (N355, N334, N195, N283);
buf BUF1 (N356, N344);
or OR2 (N357, N336, N136);
and AND3 (N358, N354, N293, N233);
xor XOR2 (N359, N350, N104);
not NOT1 (N360, N353);
and AND2 (N361, N345, N324);
xor XOR2 (N362, N357, N215);
nor NOR3 (N363, N356, N172, N176);
not NOT1 (N364, N359);
nor NOR4 (N365, N342, N291, N281, N113);
nor NOR2 (N366, N362, N360);
and AND4 (N367, N118, N162, N307, N133);
and AND3 (N368, N364, N97, N183);
or OR2 (N369, N351, N45);
and AND2 (N370, N367, N309);
xor XOR2 (N371, N355, N349);
not NOT1 (N372, N16);
or OR4 (N373, N371, N347, N154, N262);
buf BUF1 (N374, N369);
buf BUF1 (N375, N361);
not NOT1 (N376, N370);
buf BUF1 (N377, N375);
not NOT1 (N378, N372);
nor NOR4 (N379, N368, N257, N162, N81);
or OR3 (N380, N358, N132, N95);
xor XOR2 (N381, N373, N100);
and AND2 (N382, N380, N361);
and AND4 (N383, N381, N148, N56, N79);
or OR2 (N384, N376, N118);
or OR2 (N385, N379, N231);
buf BUF1 (N386, N383);
or OR4 (N387, N365, N359, N212, N287);
not NOT1 (N388, N366);
and AND3 (N389, N377, N101, N265);
not NOT1 (N390, N387);
and AND2 (N391, N390, N111);
or OR2 (N392, N378, N285);
xor XOR2 (N393, N392, N48);
and AND4 (N394, N393, N266, N338, N267);
xor XOR2 (N395, N363, N127);
or OR2 (N396, N384, N66);
xor XOR2 (N397, N374, N72);
buf BUF1 (N398, N396);
and AND4 (N399, N391, N312, N241, N332);
nor NOR3 (N400, N398, N59, N25);
not NOT1 (N401, N399);
nand NAND2 (N402, N386, N233);
nand NAND3 (N403, N389, N123, N368);
buf BUF1 (N404, N403);
or OR2 (N405, N394, N32);
buf BUF1 (N406, N402);
and AND2 (N407, N400, N7);
or OR2 (N408, N405, N69);
nand NAND4 (N409, N408, N81, N23, N85);
nor NOR2 (N410, N401, N110);
xor XOR2 (N411, N388, N217);
nand NAND4 (N412, N406, N16, N18, N58);
buf BUF1 (N413, N382);
or OR2 (N414, N410, N342);
not NOT1 (N415, N411);
buf BUF1 (N416, N404);
and AND3 (N417, N412, N124, N400);
nand NAND4 (N418, N397, N90, N331, N156);
and AND4 (N419, N416, N113, N34, N377);
nor NOR3 (N420, N407, N263, N132);
or OR2 (N421, N414, N81);
nor NOR4 (N422, N395, N98, N270, N121);
xor XOR2 (N423, N420, N208);
nor NOR4 (N424, N421, N163, N109, N122);
buf BUF1 (N425, N415);
buf BUF1 (N426, N413);
or OR4 (N427, N423, N380, N279, N148);
buf BUF1 (N428, N424);
and AND3 (N429, N422, N225, N343);
xor XOR2 (N430, N427, N354);
buf BUF1 (N431, N385);
and AND2 (N432, N425, N85);
and AND2 (N433, N419, N30);
nand NAND3 (N434, N430, N169, N201);
nor NOR3 (N435, N434, N247, N254);
nand NAND4 (N436, N417, N282, N326, N44);
xor XOR2 (N437, N409, N79);
nand NAND4 (N438, N418, N133, N46, N185);
not NOT1 (N439, N431);
nand NAND2 (N440, N435, N290);
buf BUF1 (N441, N428);
nor NOR4 (N442, N439, N118, N400, N62);
nor NOR2 (N443, N436, N145);
buf BUF1 (N444, N441);
and AND4 (N445, N429, N78, N348, N422);
nor NOR3 (N446, N444, N399, N148);
nor NOR4 (N447, N432, N228, N61, N204);
not NOT1 (N448, N440);
buf BUF1 (N449, N443);
nand NAND4 (N450, N448, N345, N34, N38);
buf BUF1 (N451, N438);
xor XOR2 (N452, N449, N103);
not NOT1 (N453, N450);
nor NOR3 (N454, N445, N399, N414);
buf BUF1 (N455, N447);
nand NAND2 (N456, N452, N236);
xor XOR2 (N457, N442, N221);
xor XOR2 (N458, N456, N251);
or OR3 (N459, N453, N169, N84);
xor XOR2 (N460, N451, N72);
not NOT1 (N461, N455);
buf BUF1 (N462, N454);
nor NOR2 (N463, N459, N383);
nand NAND2 (N464, N463, N317);
and AND3 (N465, N464, N28, N413);
buf BUF1 (N466, N446);
or OR3 (N467, N458, N226, N373);
and AND2 (N468, N437, N286);
nor NOR4 (N469, N468, N98, N228, N435);
xor XOR2 (N470, N460, N1);
or OR4 (N471, N465, N187, N212, N62);
buf BUF1 (N472, N462);
nor NOR2 (N473, N457, N333);
not NOT1 (N474, N461);
nor NOR4 (N475, N466, N173, N290, N204);
buf BUF1 (N476, N474);
or OR4 (N477, N476, N383, N468, N453);
or OR3 (N478, N469, N443, N458);
xor XOR2 (N479, N473, N284);
not NOT1 (N480, N479);
nor NOR2 (N481, N478, N459);
nor NOR4 (N482, N481, N27, N36, N122);
nor NOR3 (N483, N470, N139, N252);
not NOT1 (N484, N477);
and AND2 (N485, N426, N95);
nor NOR2 (N486, N467, N361);
or OR3 (N487, N472, N160, N200);
not NOT1 (N488, N486);
nand NAND4 (N489, N483, N385, N344, N138);
not NOT1 (N490, N482);
buf BUF1 (N491, N489);
buf BUF1 (N492, N433);
xor XOR2 (N493, N490, N342);
nand NAND4 (N494, N493, N239, N253, N341);
or OR2 (N495, N492, N8);
and AND3 (N496, N480, N168, N83);
nor NOR3 (N497, N495, N103, N388);
nand NAND4 (N498, N484, N431, N279, N21);
nand NAND3 (N499, N494, N224, N64);
xor XOR2 (N500, N487, N93);
nor NOR3 (N501, N488, N106, N276);
nand NAND3 (N502, N475, N287, N491);
buf BUF1 (N503, N293);
not NOT1 (N504, N498);
nor NOR4 (N505, N500, N139, N197, N5);
xor XOR2 (N506, N499, N70);
buf BUF1 (N507, N505);
xor XOR2 (N508, N503, N421);
or OR4 (N509, N501, N254, N123, N500);
or OR3 (N510, N497, N391, N478);
and AND2 (N511, N507, N447);
and AND4 (N512, N496, N86, N128, N486);
not NOT1 (N513, N485);
buf BUF1 (N514, N504);
nand NAND3 (N515, N506, N400, N444);
xor XOR2 (N516, N508, N288);
nand NAND2 (N517, N509, N88);
xor XOR2 (N518, N516, N55);
not NOT1 (N519, N517);
nand NAND3 (N520, N511, N506, N354);
buf BUF1 (N521, N520);
xor XOR2 (N522, N513, N488);
buf BUF1 (N523, N514);
xor XOR2 (N524, N510, N323);
or OR2 (N525, N519, N335);
nand NAND4 (N526, N522, N14, N304, N310);
nor NOR4 (N527, N502, N46, N165, N325);
nor NOR3 (N528, N515, N460, N274);
or OR3 (N529, N471, N14, N54);
buf BUF1 (N530, N527);
or OR4 (N531, N530, N242, N245, N501);
nor NOR2 (N532, N521, N163);
nand NAND2 (N533, N518, N445);
nand NAND3 (N534, N529, N147, N324);
nand NAND4 (N535, N512, N458, N74, N270);
nor NOR4 (N536, N532, N349, N12, N171);
not NOT1 (N537, N524);
buf BUF1 (N538, N523);
and AND4 (N539, N528, N419, N351, N212);
xor XOR2 (N540, N538, N169);
or OR3 (N541, N533, N344, N229);
or OR4 (N542, N531, N22, N524, N215);
or OR2 (N543, N536, N442);
xor XOR2 (N544, N539, N188);
nor NOR3 (N545, N542, N487, N67);
xor XOR2 (N546, N526, N3);
nand NAND2 (N547, N544, N422);
not NOT1 (N548, N537);
buf BUF1 (N549, N543);
not NOT1 (N550, N525);
nor NOR2 (N551, N548, N466);
and AND2 (N552, N535, N96);
not NOT1 (N553, N549);
or OR4 (N554, N552, N133, N166, N44);
xor XOR2 (N555, N547, N86);
nor NOR4 (N556, N546, N393, N108, N292);
nor NOR3 (N557, N551, N114, N199);
not NOT1 (N558, N556);
nand NAND4 (N559, N534, N390, N200, N523);
xor XOR2 (N560, N553, N427);
or OR2 (N561, N557, N27);
nand NAND2 (N562, N561, N47);
nand NAND4 (N563, N562, N437, N150, N407);
nand NAND2 (N564, N540, N261);
and AND3 (N565, N560, N110, N284);
or OR4 (N566, N555, N134, N278, N86);
not NOT1 (N567, N564);
and AND3 (N568, N559, N378, N90);
not NOT1 (N569, N550);
xor XOR2 (N570, N545, N256);
xor XOR2 (N571, N569, N465);
and AND3 (N572, N568, N78, N247);
and AND3 (N573, N570, N127, N128);
xor XOR2 (N574, N565, N388);
nand NAND4 (N575, N574, N137, N511, N222);
buf BUF1 (N576, N573);
buf BUF1 (N577, N567);
or OR2 (N578, N575, N421);
buf BUF1 (N579, N572);
nor NOR2 (N580, N571, N73);
nor NOR4 (N581, N577, N433, N256, N325);
nand NAND3 (N582, N579, N137, N349);
buf BUF1 (N583, N581);
nor NOR4 (N584, N558, N356, N254, N514);
buf BUF1 (N585, N578);
nand NAND4 (N586, N584, N79, N126, N147);
nor NOR4 (N587, N580, N470, N413, N259);
not NOT1 (N588, N587);
nor NOR4 (N589, N583, N511, N458, N448);
and AND3 (N590, N563, N502, N148);
or OR2 (N591, N590, N590);
not NOT1 (N592, N589);
nand NAND3 (N593, N541, N262, N47);
xor XOR2 (N594, N586, N280);
and AND3 (N595, N592, N5, N342);
nand NAND2 (N596, N591, N548);
or OR3 (N597, N593, N572, N17);
or OR4 (N598, N566, N494, N499, N301);
xor XOR2 (N599, N598, N488);
buf BUF1 (N600, N588);
and AND4 (N601, N594, N332, N359, N293);
and AND2 (N602, N554, N495);
buf BUF1 (N603, N599);
xor XOR2 (N604, N585, N14);
or OR3 (N605, N603, N541, N91);
and AND3 (N606, N601, N196, N517);
xor XOR2 (N607, N597, N1);
nor NOR2 (N608, N595, N104);
or OR3 (N609, N608, N213, N497);
buf BUF1 (N610, N600);
and AND3 (N611, N602, N359, N311);
or OR2 (N612, N609, N276);
buf BUF1 (N613, N611);
buf BUF1 (N614, N610);
nor NOR4 (N615, N582, N481, N112, N212);
buf BUF1 (N616, N615);
and AND3 (N617, N616, N56, N38);
nor NOR3 (N618, N604, N100, N333);
nand NAND3 (N619, N614, N502, N332);
nor NOR2 (N620, N619, N590);
nand NAND3 (N621, N618, N366, N528);
xor XOR2 (N622, N605, N191);
nor NOR3 (N623, N617, N486, N145);
nor NOR2 (N624, N576, N337);
not NOT1 (N625, N612);
or OR3 (N626, N596, N54, N614);
xor XOR2 (N627, N621, N558);
not NOT1 (N628, N626);
buf BUF1 (N629, N628);
nor NOR3 (N630, N607, N124, N155);
nand NAND3 (N631, N620, N218, N79);
not NOT1 (N632, N625);
and AND3 (N633, N613, N104, N432);
xor XOR2 (N634, N606, N496);
nor NOR3 (N635, N631, N365, N629);
not NOT1 (N636, N27);
buf BUF1 (N637, N627);
nand NAND4 (N638, N634, N179, N363, N624);
xor XOR2 (N639, N225, N71);
and AND4 (N640, N636, N369, N173, N193);
nor NOR3 (N641, N632, N398, N220);
or OR2 (N642, N638, N1);
not NOT1 (N643, N640);
xor XOR2 (N644, N633, N516);
and AND4 (N645, N630, N234, N364, N152);
or OR4 (N646, N644, N585, N431, N522);
and AND4 (N647, N637, N568, N286, N563);
not NOT1 (N648, N645);
or OR3 (N649, N623, N36, N607);
and AND4 (N650, N646, N634, N13, N25);
nand NAND3 (N651, N650, N129, N530);
and AND4 (N652, N641, N16, N390, N553);
not NOT1 (N653, N622);
xor XOR2 (N654, N647, N142);
and AND2 (N655, N642, N462);
nor NOR2 (N656, N652, N26);
or OR4 (N657, N643, N595, N416, N204);
or OR4 (N658, N657, N265, N255, N401);
buf BUF1 (N659, N656);
nor NOR3 (N660, N649, N374, N142);
nor NOR3 (N661, N648, N535, N393);
nand NAND3 (N662, N655, N591, N415);
xor XOR2 (N663, N635, N105);
or OR4 (N664, N662, N430, N206, N174);
not NOT1 (N665, N651);
buf BUF1 (N666, N653);
nor NOR3 (N667, N666, N634, N179);
not NOT1 (N668, N667);
xor XOR2 (N669, N639, N560);
and AND2 (N670, N663, N370);
or OR4 (N671, N654, N145, N621, N251);
not NOT1 (N672, N669);
nand NAND3 (N673, N672, N230, N634);
or OR3 (N674, N668, N207, N158);
or OR3 (N675, N674, N331, N543);
nor NOR2 (N676, N675, N294);
or OR4 (N677, N661, N324, N179, N342);
nor NOR3 (N678, N670, N13, N42);
not NOT1 (N679, N677);
and AND4 (N680, N676, N92, N261, N163);
nand NAND2 (N681, N664, N200);
not NOT1 (N682, N671);
or OR4 (N683, N682, N643, N226, N606);
buf BUF1 (N684, N680);
or OR2 (N685, N678, N239);
nand NAND2 (N686, N658, N523);
not NOT1 (N687, N686);
or OR2 (N688, N660, N271);
or OR4 (N689, N688, N192, N296, N455);
not NOT1 (N690, N659);
or OR3 (N691, N665, N646, N131);
or OR4 (N692, N690, N29, N174, N450);
or OR3 (N693, N679, N612, N307);
buf BUF1 (N694, N691);
xor XOR2 (N695, N683, N653);
nand NAND4 (N696, N692, N420, N210, N285);
xor XOR2 (N697, N687, N377);
and AND3 (N698, N695, N142, N537);
nor NOR4 (N699, N684, N287, N74, N104);
nor NOR4 (N700, N698, N99, N225, N26);
nor NOR3 (N701, N699, N700, N350);
nor NOR3 (N702, N46, N529, N52);
not NOT1 (N703, N701);
and AND2 (N704, N685, N167);
buf BUF1 (N705, N693);
nor NOR2 (N706, N704, N140);
or OR2 (N707, N705, N297);
buf BUF1 (N708, N703);
not NOT1 (N709, N706);
buf BUF1 (N710, N681);
or OR4 (N711, N709, N293, N560, N89);
not NOT1 (N712, N694);
or OR3 (N713, N711, N540, N404);
nand NAND3 (N714, N689, N113, N147);
xor XOR2 (N715, N713, N500);
buf BUF1 (N716, N702);
buf BUF1 (N717, N716);
or OR3 (N718, N697, N617, N258);
xor XOR2 (N719, N718, N65);
nor NOR3 (N720, N710, N509, N188);
or OR4 (N721, N714, N21, N235, N134);
not NOT1 (N722, N720);
nand NAND2 (N723, N696, N5);
not NOT1 (N724, N719);
or OR2 (N725, N724, N720);
and AND3 (N726, N715, N327, N529);
nand NAND4 (N727, N712, N657, N276, N41);
buf BUF1 (N728, N717);
buf BUF1 (N729, N725);
not NOT1 (N730, N729);
nand NAND4 (N731, N721, N60, N249, N358);
and AND4 (N732, N707, N714, N499, N581);
not NOT1 (N733, N731);
and AND2 (N734, N733, N514);
and AND2 (N735, N708, N453);
and AND4 (N736, N727, N389, N152, N598);
buf BUF1 (N737, N726);
nor NOR4 (N738, N734, N640, N216, N524);
not NOT1 (N739, N673);
xor XOR2 (N740, N722, N703);
buf BUF1 (N741, N730);
or OR3 (N742, N741, N113, N301);
xor XOR2 (N743, N740, N629);
or OR3 (N744, N737, N515, N588);
and AND4 (N745, N736, N260, N453, N50);
or OR2 (N746, N745, N551);
xor XOR2 (N747, N739, N447);
or OR4 (N748, N747, N642, N181, N41);
and AND3 (N749, N728, N184, N485);
or OR4 (N750, N732, N597, N622, N339);
xor XOR2 (N751, N750, N511);
or OR2 (N752, N751, N384);
buf BUF1 (N753, N723);
and AND3 (N754, N735, N552, N699);
and AND2 (N755, N749, N103);
and AND3 (N756, N746, N100, N468);
xor XOR2 (N757, N755, N390);
or OR3 (N758, N743, N39, N568);
nor NOR3 (N759, N756, N333, N385);
not NOT1 (N760, N753);
nand NAND4 (N761, N758, N643, N428, N575);
not NOT1 (N762, N759);
or OR4 (N763, N754, N19, N239, N518);
nand NAND4 (N764, N757, N206, N439, N343);
nand NAND2 (N765, N748, N627);
nand NAND4 (N766, N742, N455, N25, N652);
or OR4 (N767, N744, N716, N377, N750);
not NOT1 (N768, N761);
not NOT1 (N769, N760);
buf BUF1 (N770, N762);
or OR3 (N771, N764, N661, N361);
nor NOR3 (N772, N770, N514, N668);
nand NAND2 (N773, N768, N13);
xor XOR2 (N774, N765, N155);
or OR3 (N775, N766, N414, N22);
xor XOR2 (N776, N775, N388);
buf BUF1 (N777, N776);
buf BUF1 (N778, N738);
and AND4 (N779, N767, N256, N199, N137);
nor NOR4 (N780, N772, N644, N322, N490);
nor NOR2 (N781, N752, N35);
xor XOR2 (N782, N778, N513);
xor XOR2 (N783, N777, N211);
and AND4 (N784, N781, N333, N221, N345);
and AND4 (N785, N779, N594, N76, N645);
or OR4 (N786, N785, N766, N536, N628);
not NOT1 (N787, N786);
not NOT1 (N788, N771);
nor NOR4 (N789, N773, N22, N497, N349);
nand NAND2 (N790, N787, N119);
not NOT1 (N791, N763);
buf BUF1 (N792, N780);
and AND3 (N793, N789, N348, N325);
xor XOR2 (N794, N790, N616);
nand NAND3 (N795, N784, N85, N93);
buf BUF1 (N796, N794);
or OR2 (N797, N782, N178);
not NOT1 (N798, N796);
and AND4 (N799, N797, N277, N194, N51);
and AND3 (N800, N769, N482, N772);
nand NAND4 (N801, N798, N53, N560, N520);
not NOT1 (N802, N795);
nor NOR2 (N803, N774, N702);
xor XOR2 (N804, N791, N350);
not NOT1 (N805, N803);
nand NAND3 (N806, N804, N498, N160);
nor NOR4 (N807, N801, N781, N703, N680);
nand NAND3 (N808, N807, N146, N62);
and AND2 (N809, N805, N216);
and AND3 (N810, N808, N656, N505);
and AND4 (N811, N783, N222, N110, N483);
nand NAND2 (N812, N788, N99);
and AND4 (N813, N802, N44, N251, N596);
buf BUF1 (N814, N810);
and AND2 (N815, N799, N355);
nand NAND4 (N816, N809, N534, N280, N145);
buf BUF1 (N817, N815);
nor NOR2 (N818, N811, N94);
nor NOR3 (N819, N793, N427, N303);
nor NOR4 (N820, N819, N667, N331, N741);
and AND4 (N821, N792, N161, N758, N525);
and AND3 (N822, N806, N407, N84);
nand NAND2 (N823, N813, N234);
xor XOR2 (N824, N818, N60);
and AND2 (N825, N817, N218);
buf BUF1 (N826, N820);
or OR3 (N827, N816, N433, N632);
nor NOR4 (N828, N814, N259, N585, N514);
not NOT1 (N829, N812);
and AND4 (N830, N824, N478, N81, N156);
not NOT1 (N831, N821);
nand NAND3 (N832, N825, N792, N374);
and AND2 (N833, N826, N618);
not NOT1 (N834, N829);
not NOT1 (N835, N800);
or OR2 (N836, N831, N231);
or OR3 (N837, N828, N123, N249);
and AND2 (N838, N830, N558);
and AND4 (N839, N836, N233, N827, N307);
or OR2 (N840, N511, N400);
buf BUF1 (N841, N822);
nor NOR2 (N842, N840, N813);
buf BUF1 (N843, N834);
and AND2 (N844, N833, N281);
or OR4 (N845, N842, N1, N597, N389);
and AND3 (N846, N841, N505, N759);
and AND4 (N847, N846, N200, N45, N181);
not NOT1 (N848, N845);
buf BUF1 (N849, N823);
and AND3 (N850, N835, N638, N399);
nor NOR3 (N851, N848, N708, N262);
or OR3 (N852, N839, N731, N822);
and AND3 (N853, N843, N284, N524);
not NOT1 (N854, N853);
not NOT1 (N855, N851);
and AND3 (N856, N838, N61, N104);
buf BUF1 (N857, N850);
not NOT1 (N858, N856);
nor NOR2 (N859, N844, N578);
and AND3 (N860, N857, N761, N610);
xor XOR2 (N861, N854, N711);
buf BUF1 (N862, N859);
not NOT1 (N863, N855);
nand NAND3 (N864, N832, N856, N258);
xor XOR2 (N865, N837, N334);
or OR3 (N866, N849, N43, N91);
not NOT1 (N867, N852);
or OR3 (N868, N860, N68, N839);
and AND2 (N869, N847, N112);
or OR3 (N870, N866, N818, N574);
not NOT1 (N871, N865);
buf BUF1 (N872, N868);
and AND2 (N873, N863, N650);
xor XOR2 (N874, N858, N589);
xor XOR2 (N875, N861, N57);
buf BUF1 (N876, N862);
or OR2 (N877, N875, N31);
buf BUF1 (N878, N864);
xor XOR2 (N879, N874, N819);
or OR2 (N880, N873, N585);
nor NOR3 (N881, N876, N60, N180);
or OR2 (N882, N869, N562);
nand NAND2 (N883, N871, N263);
and AND3 (N884, N872, N680, N171);
xor XOR2 (N885, N879, N748);
xor XOR2 (N886, N877, N822);
buf BUF1 (N887, N884);
nand NAND2 (N888, N886, N590);
not NOT1 (N889, N882);
and AND3 (N890, N885, N338, N556);
not NOT1 (N891, N888);
buf BUF1 (N892, N890);
or OR3 (N893, N887, N633, N475);
and AND2 (N894, N891, N169);
buf BUF1 (N895, N880);
nand NAND2 (N896, N878, N484);
xor XOR2 (N897, N896, N661);
not NOT1 (N898, N870);
and AND4 (N899, N898, N522, N212, N748);
or OR2 (N900, N881, N353);
nand NAND3 (N901, N894, N405, N506);
xor XOR2 (N902, N892, N692);
and AND4 (N903, N883, N455, N135, N168);
and AND3 (N904, N895, N455, N418);
nand NAND2 (N905, N901, N426);
or OR4 (N906, N900, N488, N551, N88);
buf BUF1 (N907, N893);
and AND2 (N908, N867, N405);
xor XOR2 (N909, N902, N730);
and AND2 (N910, N909, N7);
nand NAND4 (N911, N906, N276, N60, N664);
buf BUF1 (N912, N910);
buf BUF1 (N913, N904);
nand NAND4 (N914, N911, N896, N76, N592);
nor NOR3 (N915, N903, N477, N497);
and AND2 (N916, N889, N574);
or OR4 (N917, N908, N449, N263, N93);
not NOT1 (N918, N916);
not NOT1 (N919, N917);
nand NAND3 (N920, N915, N221, N347);
and AND4 (N921, N918, N358, N25, N915);
not NOT1 (N922, N920);
nor NOR3 (N923, N914, N495, N485);
xor XOR2 (N924, N897, N693);
and AND3 (N925, N921, N494, N62);
nor NOR4 (N926, N924, N768, N590, N756);
nor NOR2 (N927, N923, N490);
not NOT1 (N928, N922);
buf BUF1 (N929, N928);
not NOT1 (N930, N926);
and AND2 (N931, N905, N394);
nand NAND3 (N932, N929, N381, N45);
xor XOR2 (N933, N927, N572);
nor NOR2 (N934, N919, N164);
xor XOR2 (N935, N930, N31);
nand NAND4 (N936, N913, N813, N160, N489);
not NOT1 (N937, N935);
nand NAND4 (N938, N937, N750, N822, N581);
nor NOR4 (N939, N932, N428, N109, N640);
buf BUF1 (N940, N907);
buf BUF1 (N941, N899);
buf BUF1 (N942, N939);
or OR4 (N943, N934, N839, N594, N110);
buf BUF1 (N944, N912);
or OR4 (N945, N943, N397, N159, N732);
not NOT1 (N946, N925);
nand NAND4 (N947, N938, N791, N443, N880);
or OR4 (N948, N946, N564, N242, N112);
nand NAND4 (N949, N947, N311, N696, N497);
and AND2 (N950, N942, N596);
or OR2 (N951, N933, N794);
xor XOR2 (N952, N940, N692);
buf BUF1 (N953, N948);
xor XOR2 (N954, N953, N798);
buf BUF1 (N955, N950);
or OR3 (N956, N941, N356, N227);
nand NAND3 (N957, N931, N96, N239);
buf BUF1 (N958, N945);
buf BUF1 (N959, N955);
xor XOR2 (N960, N952, N827);
not NOT1 (N961, N956);
xor XOR2 (N962, N957, N558);
nor NOR2 (N963, N962, N172);
nor NOR2 (N964, N954, N944);
nand NAND4 (N965, N371, N344, N616, N891);
and AND2 (N966, N961, N945);
xor XOR2 (N967, N958, N695);
nor NOR4 (N968, N965, N375, N664, N822);
xor XOR2 (N969, N949, N478);
nand NAND4 (N970, N968, N87, N448, N617);
buf BUF1 (N971, N970);
buf BUF1 (N972, N936);
xor XOR2 (N973, N969, N185);
or OR4 (N974, N966, N758, N129, N103);
buf BUF1 (N975, N960);
nor NOR3 (N976, N959, N563, N481);
xor XOR2 (N977, N975, N173);
xor XOR2 (N978, N971, N615);
xor XOR2 (N979, N976, N741);
nor NOR2 (N980, N979, N654);
xor XOR2 (N981, N963, N143);
or OR4 (N982, N972, N331, N133, N26);
and AND2 (N983, N973, N593);
nand NAND2 (N984, N951, N556);
not NOT1 (N985, N982);
or OR4 (N986, N967, N694, N737, N503);
and AND4 (N987, N983, N270, N332, N395);
not NOT1 (N988, N987);
nand NAND2 (N989, N984, N719);
not NOT1 (N990, N980);
or OR2 (N991, N989, N375);
buf BUF1 (N992, N974);
not NOT1 (N993, N981);
or OR2 (N994, N985, N361);
buf BUF1 (N995, N991);
or OR3 (N996, N990, N498, N318);
or OR2 (N997, N995, N268);
not NOT1 (N998, N978);
or OR2 (N999, N996, N455);
buf BUF1 (N1000, N964);
nor NOR4 (N1001, N986, N767, N518, N187);
xor XOR2 (N1002, N977, N13);
not NOT1 (N1003, N992);
nor NOR2 (N1004, N1002, N364);
xor XOR2 (N1005, N1000, N897);
nor NOR2 (N1006, N993, N139);
buf BUF1 (N1007, N994);
nor NOR3 (N1008, N1007, N141, N230);
nand NAND4 (N1009, N988, N107, N927, N981);
xor XOR2 (N1010, N998, N470);
xor XOR2 (N1011, N1001, N317);
and AND2 (N1012, N997, N90);
not NOT1 (N1013, N1008);
nor NOR2 (N1014, N1003, N645);
nor NOR2 (N1015, N999, N675);
nor NOR2 (N1016, N1015, N703);
nor NOR2 (N1017, N1006, N768);
buf BUF1 (N1018, N1012);
and AND3 (N1019, N1011, N391, N489);
nor NOR2 (N1020, N1004, N62);
buf BUF1 (N1021, N1017);
buf BUF1 (N1022, N1014);
nand NAND4 (N1023, N1016, N715, N778, N58);
or OR4 (N1024, N1013, N799, N1009, N365);
nor NOR3 (N1025, N35, N520, N535);
not NOT1 (N1026, N1019);
not NOT1 (N1027, N1025);
nand NAND3 (N1028, N1005, N1011, N1013);
nor NOR3 (N1029, N1021, N507, N864);
nand NAND4 (N1030, N1018, N611, N153, N840);
not NOT1 (N1031, N1024);
nor NOR4 (N1032, N1028, N288, N97, N557);
not NOT1 (N1033, N1031);
buf BUF1 (N1034, N1030);
and AND2 (N1035, N1023, N827);
nand NAND4 (N1036, N1027, N236, N941, N326);
or OR4 (N1037, N1010, N606, N623, N428);
or OR4 (N1038, N1022, N68, N697, N61);
nor NOR3 (N1039, N1038, N778, N651);
nor NOR3 (N1040, N1026, N270, N442);
nor NOR4 (N1041, N1020, N593, N253, N346);
nand NAND4 (N1042, N1037, N530, N896, N343);
xor XOR2 (N1043, N1040, N854);
xor XOR2 (N1044, N1034, N291);
nand NAND4 (N1045, N1029, N279, N559, N457);
not NOT1 (N1046, N1036);
nor NOR3 (N1047, N1032, N813, N773);
and AND2 (N1048, N1041, N659);
xor XOR2 (N1049, N1044, N174);
or OR4 (N1050, N1033, N616, N728, N412);
or OR2 (N1051, N1046, N985);
and AND4 (N1052, N1050, N839, N286, N379);
not NOT1 (N1053, N1042);
buf BUF1 (N1054, N1048);
and AND4 (N1055, N1054, N62, N814, N35);
nor NOR3 (N1056, N1055, N400, N372);
not NOT1 (N1057, N1049);
buf BUF1 (N1058, N1043);
buf BUF1 (N1059, N1045);
and AND4 (N1060, N1053, N775, N918, N310);
nand NAND4 (N1061, N1035, N187, N931, N721);
not NOT1 (N1062, N1047);
nor NOR2 (N1063, N1052, N851);
nand NAND4 (N1064, N1062, N118, N514, N706);
not NOT1 (N1065, N1057);
xor XOR2 (N1066, N1061, N747);
nand NAND2 (N1067, N1066, N626);
or OR2 (N1068, N1063, N906);
buf BUF1 (N1069, N1056);
buf BUF1 (N1070, N1059);
nand NAND2 (N1071, N1058, N30);
not NOT1 (N1072, N1065);
or OR2 (N1073, N1072, N1032);
buf BUF1 (N1074, N1070);
nor NOR2 (N1075, N1069, N165);
not NOT1 (N1076, N1074);
nand NAND2 (N1077, N1071, N180);
buf BUF1 (N1078, N1076);
and AND4 (N1079, N1067, N325, N740, N647);
nand NAND3 (N1080, N1075, N497, N140);
nor NOR4 (N1081, N1051, N677, N10, N121);
nor NOR3 (N1082, N1039, N592, N676);
and AND4 (N1083, N1064, N109, N808, N600);
or OR4 (N1084, N1080, N895, N339, N1047);
nand NAND4 (N1085, N1078, N341, N241, N1082);
xor XOR2 (N1086, N292, N275);
not NOT1 (N1087, N1077);
buf BUF1 (N1088, N1060);
xor XOR2 (N1089, N1087, N193);
and AND2 (N1090, N1086, N97);
buf BUF1 (N1091, N1085);
not NOT1 (N1092, N1090);
not NOT1 (N1093, N1068);
buf BUF1 (N1094, N1083);
nor NOR2 (N1095, N1094, N1051);
or OR3 (N1096, N1088, N248, N712);
buf BUF1 (N1097, N1091);
xor XOR2 (N1098, N1096, N276);
and AND4 (N1099, N1073, N745, N387, N514);
xor XOR2 (N1100, N1092, N38);
nor NOR4 (N1101, N1097, N133, N384, N280);
and AND2 (N1102, N1089, N741);
or OR3 (N1103, N1081, N545, N476);
buf BUF1 (N1104, N1101);
nand NAND4 (N1105, N1095, N490, N878, N340);
or OR2 (N1106, N1098, N754);
buf BUF1 (N1107, N1100);
xor XOR2 (N1108, N1084, N320);
or OR2 (N1109, N1079, N360);
xor XOR2 (N1110, N1108, N555);
nand NAND2 (N1111, N1106, N1074);
xor XOR2 (N1112, N1111, N926);
nor NOR3 (N1113, N1102, N7, N516);
and AND4 (N1114, N1113, N152, N524, N47);
and AND4 (N1115, N1093, N332, N538, N834);
not NOT1 (N1116, N1099);
nand NAND2 (N1117, N1104, N191);
and AND4 (N1118, N1107, N590, N987, N688);
xor XOR2 (N1119, N1115, N531);
not NOT1 (N1120, N1109);
nand NAND3 (N1121, N1117, N1028, N464);
xor XOR2 (N1122, N1110, N487);
nor NOR4 (N1123, N1122, N111, N930, N328);
xor XOR2 (N1124, N1114, N594);
nand NAND4 (N1125, N1120, N891, N679, N805);
and AND4 (N1126, N1103, N115, N53, N314);
xor XOR2 (N1127, N1116, N549);
and AND2 (N1128, N1127, N68);
nand NAND2 (N1129, N1118, N192);
buf BUF1 (N1130, N1112);
and AND3 (N1131, N1126, N1077, N969);
nand NAND4 (N1132, N1123, N366, N1131, N867);
not NOT1 (N1133, N1063);
buf BUF1 (N1134, N1119);
or OR4 (N1135, N1124, N390, N319, N1108);
xor XOR2 (N1136, N1135, N1073);
buf BUF1 (N1137, N1132);
nor NOR2 (N1138, N1105, N195);
xor XOR2 (N1139, N1121, N624);
buf BUF1 (N1140, N1128);
nand NAND4 (N1141, N1140, N618, N1035, N311);
buf BUF1 (N1142, N1125);
xor XOR2 (N1143, N1139, N132);
nor NOR3 (N1144, N1136, N843, N1059);
buf BUF1 (N1145, N1144);
not NOT1 (N1146, N1134);
or OR4 (N1147, N1133, N315, N821, N360);
and AND3 (N1148, N1143, N476, N762);
buf BUF1 (N1149, N1129);
nand NAND2 (N1150, N1148, N401);
not NOT1 (N1151, N1146);
or OR3 (N1152, N1130, N706, N862);
xor XOR2 (N1153, N1147, N510);
or OR3 (N1154, N1138, N195, N441);
and AND4 (N1155, N1137, N990, N1027, N235);
and AND4 (N1156, N1153, N1065, N107, N613);
nor NOR4 (N1157, N1154, N542, N68, N476);
xor XOR2 (N1158, N1152, N727);
and AND3 (N1159, N1142, N952, N374);
or OR3 (N1160, N1150, N844, N645);
xor XOR2 (N1161, N1155, N1142);
buf BUF1 (N1162, N1161);
nor NOR4 (N1163, N1160, N434, N690, N987);
xor XOR2 (N1164, N1149, N763);
xor XOR2 (N1165, N1162, N686);
nor NOR4 (N1166, N1158, N188, N50, N226);
nand NAND2 (N1167, N1145, N485);
nand NAND2 (N1168, N1163, N847);
nor NOR4 (N1169, N1157, N884, N764, N897);
xor XOR2 (N1170, N1167, N255);
nor NOR4 (N1171, N1156, N751, N641, N886);
nor NOR4 (N1172, N1151, N41, N1017, N1143);
nand NAND2 (N1173, N1159, N341);
not NOT1 (N1174, N1165);
buf BUF1 (N1175, N1166);
not NOT1 (N1176, N1170);
xor XOR2 (N1177, N1168, N947);
buf BUF1 (N1178, N1169);
or OR4 (N1179, N1174, N92, N860, N85);
nand NAND2 (N1180, N1171, N132);
and AND2 (N1181, N1180, N1178);
and AND3 (N1182, N881, N1168, N48);
or OR3 (N1183, N1172, N571, N1011);
and AND4 (N1184, N1182, N899, N1053, N139);
and AND3 (N1185, N1164, N221, N638);
not NOT1 (N1186, N1181);
and AND3 (N1187, N1177, N69, N126);
nor NOR4 (N1188, N1179, N209, N179, N75);
or OR2 (N1189, N1141, N235);
buf BUF1 (N1190, N1186);
nor NOR4 (N1191, N1187, N1144, N496, N279);
buf BUF1 (N1192, N1188);
or OR3 (N1193, N1184, N109, N627);
buf BUF1 (N1194, N1190);
buf BUF1 (N1195, N1193);
buf BUF1 (N1196, N1176);
and AND3 (N1197, N1173, N845, N151);
and AND4 (N1198, N1192, N879, N31, N793);
nand NAND3 (N1199, N1189, N1091, N629);
or OR4 (N1200, N1194, N610, N1156, N252);
xor XOR2 (N1201, N1200, N1172);
xor XOR2 (N1202, N1195, N824);
nor NOR3 (N1203, N1196, N92, N963);
or OR4 (N1204, N1191, N795, N469, N1018);
nor NOR2 (N1205, N1183, N955);
nand NAND3 (N1206, N1185, N822, N517);
nand NAND3 (N1207, N1202, N1057, N1006);
or OR3 (N1208, N1205, N100, N983);
and AND3 (N1209, N1203, N1183, N484);
and AND3 (N1210, N1206, N1089, N893);
nor NOR2 (N1211, N1209, N965);
and AND4 (N1212, N1208, N403, N558, N82);
not NOT1 (N1213, N1201);
buf BUF1 (N1214, N1199);
buf BUF1 (N1215, N1175);
nand NAND3 (N1216, N1213, N1040, N803);
buf BUF1 (N1217, N1207);
or OR4 (N1218, N1217, N106, N582, N921);
nand NAND4 (N1219, N1204, N280, N1194, N360);
not NOT1 (N1220, N1198);
and AND4 (N1221, N1215, N24, N609, N74);
or OR2 (N1222, N1210, N192);
and AND2 (N1223, N1197, N253);
nand NAND2 (N1224, N1221, N379);
buf BUF1 (N1225, N1222);
nor NOR4 (N1226, N1214, N575, N316, N891);
or OR3 (N1227, N1219, N398, N249);
nand NAND2 (N1228, N1212, N585);
buf BUF1 (N1229, N1228);
or OR3 (N1230, N1220, N558, N200);
nor NOR2 (N1231, N1225, N170);
and AND4 (N1232, N1227, N1206, N1039, N359);
and AND2 (N1233, N1231, N302);
buf BUF1 (N1234, N1229);
or OR4 (N1235, N1211, N769, N1076, N1090);
not NOT1 (N1236, N1226);
and AND2 (N1237, N1234, N941);
or OR2 (N1238, N1218, N585);
nand NAND4 (N1239, N1232, N862, N610, N895);
nor NOR4 (N1240, N1230, N529, N217, N1140);
xor XOR2 (N1241, N1236, N803);
nand NAND2 (N1242, N1240, N1217);
or OR4 (N1243, N1238, N272, N1003, N885);
and AND3 (N1244, N1224, N976, N309);
nand NAND3 (N1245, N1241, N877, N398);
or OR3 (N1246, N1216, N1153, N1065);
not NOT1 (N1247, N1223);
xor XOR2 (N1248, N1233, N1141);
nor NOR4 (N1249, N1242, N781, N991, N828);
buf BUF1 (N1250, N1235);
and AND4 (N1251, N1243, N437, N1242, N1217);
nand NAND4 (N1252, N1237, N705, N409, N901);
nor NOR3 (N1253, N1247, N140, N87);
xor XOR2 (N1254, N1252, N383);
buf BUF1 (N1255, N1248);
and AND4 (N1256, N1251, N785, N754, N810);
nand NAND2 (N1257, N1253, N143);
nand NAND3 (N1258, N1257, N660, N716);
nand NAND4 (N1259, N1256, N836, N518, N377);
nand NAND4 (N1260, N1258, N664, N1051, N972);
or OR3 (N1261, N1245, N1089, N110);
nor NOR2 (N1262, N1250, N402);
buf BUF1 (N1263, N1239);
nor NOR3 (N1264, N1261, N97, N523);
nand NAND4 (N1265, N1259, N966, N617, N320);
xor XOR2 (N1266, N1260, N897);
xor XOR2 (N1267, N1262, N768);
nor NOR2 (N1268, N1249, N802);
nand NAND2 (N1269, N1267, N122);
nor NOR3 (N1270, N1264, N151, N175);
or OR2 (N1271, N1269, N1);
not NOT1 (N1272, N1244);
xor XOR2 (N1273, N1272, N465);
not NOT1 (N1274, N1246);
not NOT1 (N1275, N1254);
nand NAND2 (N1276, N1268, N215);
not NOT1 (N1277, N1265);
nand NAND4 (N1278, N1271, N933, N1031, N218);
buf BUF1 (N1279, N1274);
or OR3 (N1280, N1273, N265, N1024);
xor XOR2 (N1281, N1279, N904);
or OR4 (N1282, N1270, N291, N406, N1069);
and AND3 (N1283, N1280, N645, N136);
not NOT1 (N1284, N1275);
xor XOR2 (N1285, N1281, N176);
buf BUF1 (N1286, N1278);
xor XOR2 (N1287, N1266, N1173);
and AND3 (N1288, N1263, N43, N863);
nand NAND2 (N1289, N1286, N165);
buf BUF1 (N1290, N1284);
buf BUF1 (N1291, N1288);
buf BUF1 (N1292, N1287);
xor XOR2 (N1293, N1283, N524);
buf BUF1 (N1294, N1255);
nand NAND2 (N1295, N1282, N383);
nand NAND3 (N1296, N1276, N474, N209);
not NOT1 (N1297, N1291);
not NOT1 (N1298, N1296);
or OR2 (N1299, N1292, N1141);
not NOT1 (N1300, N1293);
not NOT1 (N1301, N1285);
not NOT1 (N1302, N1299);
not NOT1 (N1303, N1298);
buf BUF1 (N1304, N1294);
xor XOR2 (N1305, N1290, N20);
buf BUF1 (N1306, N1297);
or OR3 (N1307, N1304, N1115, N1073);
not NOT1 (N1308, N1306);
nand NAND2 (N1309, N1277, N835);
or OR3 (N1310, N1308, N58, N1049);
not NOT1 (N1311, N1303);
nand NAND3 (N1312, N1309, N830, N838);
nand NAND4 (N1313, N1312, N827, N1078, N24);
nor NOR4 (N1314, N1289, N168, N206, N1308);
or OR3 (N1315, N1311, N480, N1123);
and AND2 (N1316, N1302, N1046);
buf BUF1 (N1317, N1295);
nor NOR3 (N1318, N1300, N52, N60);
buf BUF1 (N1319, N1301);
not NOT1 (N1320, N1319);
and AND4 (N1321, N1317, N272, N732, N749);
and AND2 (N1322, N1318, N1226);
and AND3 (N1323, N1315, N420, N372);
or OR2 (N1324, N1305, N980);
nor NOR4 (N1325, N1313, N888, N526, N1235);
nor NOR4 (N1326, N1314, N712, N1108, N699);
or OR2 (N1327, N1323, N1072);
or OR4 (N1328, N1327, N154, N483, N610);
not NOT1 (N1329, N1321);
buf BUF1 (N1330, N1310);
or OR2 (N1331, N1307, N479);
buf BUF1 (N1332, N1330);
nand NAND4 (N1333, N1316, N647, N163, N685);
buf BUF1 (N1334, N1325);
nand NAND3 (N1335, N1333, N319, N638);
xor XOR2 (N1336, N1332, N1279);
not NOT1 (N1337, N1334);
nand NAND3 (N1338, N1331, N158, N1287);
or OR2 (N1339, N1335, N258);
nor NOR3 (N1340, N1329, N1, N33);
xor XOR2 (N1341, N1336, N816);
nand NAND4 (N1342, N1328, N357, N1306, N1136);
and AND4 (N1343, N1326, N1323, N1019, N250);
not NOT1 (N1344, N1339);
and AND2 (N1345, N1338, N1020);
xor XOR2 (N1346, N1340, N37);
or OR2 (N1347, N1324, N1320);
nor NOR4 (N1348, N242, N23, N783, N342);
nand NAND2 (N1349, N1342, N601);
xor XOR2 (N1350, N1343, N1088);
not NOT1 (N1351, N1337);
not NOT1 (N1352, N1347);
not NOT1 (N1353, N1346);
nand NAND4 (N1354, N1353, N815, N795, N871);
nor NOR2 (N1355, N1349, N68);
buf BUF1 (N1356, N1354);
and AND4 (N1357, N1322, N849, N376, N534);
buf BUF1 (N1358, N1352);
or OR3 (N1359, N1357, N281, N1154);
and AND2 (N1360, N1355, N67);
buf BUF1 (N1361, N1350);
buf BUF1 (N1362, N1361);
nand NAND3 (N1363, N1359, N809, N347);
not NOT1 (N1364, N1363);
not NOT1 (N1365, N1364);
xor XOR2 (N1366, N1351, N1055);
not NOT1 (N1367, N1344);
or OR2 (N1368, N1367, N219);
not NOT1 (N1369, N1358);
nor NOR2 (N1370, N1362, N1259);
or OR4 (N1371, N1365, N37, N572, N995);
buf BUF1 (N1372, N1345);
xor XOR2 (N1373, N1371, N953);
nand NAND2 (N1374, N1370, N105);
buf BUF1 (N1375, N1373);
buf BUF1 (N1376, N1375);
buf BUF1 (N1377, N1372);
nand NAND2 (N1378, N1374, N15);
nand NAND2 (N1379, N1368, N712);
and AND2 (N1380, N1369, N281);
not NOT1 (N1381, N1377);
xor XOR2 (N1382, N1381, N1054);
or OR3 (N1383, N1341, N998, N796);
nand NAND4 (N1384, N1348, N736, N804, N473);
not NOT1 (N1385, N1360);
and AND3 (N1386, N1379, N823, N213);
not NOT1 (N1387, N1366);
not NOT1 (N1388, N1382);
nand NAND2 (N1389, N1387, N669);
nor NOR2 (N1390, N1389, N489);
or OR3 (N1391, N1383, N748, N1380);
or OR4 (N1392, N428, N968, N1079, N1159);
xor XOR2 (N1393, N1356, N947);
and AND3 (N1394, N1392, N1181, N776);
xor XOR2 (N1395, N1378, N1034);
nor NOR4 (N1396, N1376, N813, N863, N1198);
or OR4 (N1397, N1391, N278, N1290, N299);
not NOT1 (N1398, N1396);
and AND4 (N1399, N1398, N574, N24, N503);
xor XOR2 (N1400, N1385, N53);
xor XOR2 (N1401, N1395, N1224);
xor XOR2 (N1402, N1400, N638);
not NOT1 (N1403, N1394);
or OR2 (N1404, N1403, N15);
or OR4 (N1405, N1399, N739, N1335, N823);
buf BUF1 (N1406, N1384);
and AND3 (N1407, N1405, N22, N360);
not NOT1 (N1408, N1406);
and AND2 (N1409, N1397, N1390);
buf BUF1 (N1410, N1131);
xor XOR2 (N1411, N1410, N1056);
nor NOR4 (N1412, N1388, N762, N157, N190);
nand NAND4 (N1413, N1393, N204, N755, N274);
buf BUF1 (N1414, N1402);
nor NOR3 (N1415, N1411, N147, N1153);
not NOT1 (N1416, N1412);
and AND4 (N1417, N1414, N186, N879, N256);
xor XOR2 (N1418, N1413, N423);
nand NAND4 (N1419, N1409, N511, N777, N515);
buf BUF1 (N1420, N1419);
nor NOR4 (N1421, N1404, N1028, N1255, N1047);
or OR2 (N1422, N1401, N874);
not NOT1 (N1423, N1386);
nand NAND3 (N1424, N1421, N816, N954);
or OR3 (N1425, N1422, N65, N836);
buf BUF1 (N1426, N1416);
or OR4 (N1427, N1408, N391, N1158, N1136);
xor XOR2 (N1428, N1418, N1078);
nor NOR4 (N1429, N1423, N190, N50, N941);
buf BUF1 (N1430, N1428);
buf BUF1 (N1431, N1407);
or OR2 (N1432, N1415, N380);
or OR3 (N1433, N1424, N1162, N1303);
xor XOR2 (N1434, N1433, N318);
xor XOR2 (N1435, N1430, N197);
nand NAND3 (N1436, N1417, N306, N1123);
nor NOR2 (N1437, N1427, N215);
nor NOR2 (N1438, N1432, N542);
xor XOR2 (N1439, N1438, N613);
nor NOR4 (N1440, N1439, N978, N1367, N718);
or OR3 (N1441, N1429, N286, N1146);
buf BUF1 (N1442, N1425);
xor XOR2 (N1443, N1434, N872);
not NOT1 (N1444, N1426);
or OR3 (N1445, N1431, N279, N723);
or OR3 (N1446, N1441, N1117, N107);
and AND4 (N1447, N1440, N1364, N646, N1150);
nand NAND4 (N1448, N1420, N1341, N1382, N943);
xor XOR2 (N1449, N1448, N441);
xor XOR2 (N1450, N1447, N48);
not NOT1 (N1451, N1437);
or OR4 (N1452, N1449, N161, N315, N1146);
not NOT1 (N1453, N1451);
nand NAND4 (N1454, N1443, N369, N1308, N1421);
not NOT1 (N1455, N1436);
buf BUF1 (N1456, N1445);
xor XOR2 (N1457, N1442, N1214);
nand NAND2 (N1458, N1455, N980);
not NOT1 (N1459, N1458);
nor NOR3 (N1460, N1453, N254, N1376);
nor NOR2 (N1461, N1459, N830);
or OR2 (N1462, N1444, N1061);
nor NOR2 (N1463, N1454, N739);
and AND4 (N1464, N1446, N1349, N1446, N628);
or OR4 (N1465, N1457, N808, N255, N1);
or OR2 (N1466, N1463, N778);
xor XOR2 (N1467, N1435, N627);
not NOT1 (N1468, N1450);
not NOT1 (N1469, N1467);
and AND3 (N1470, N1456, N975, N967);
xor XOR2 (N1471, N1470, N1246);
nand NAND3 (N1472, N1469, N414, N759);
buf BUF1 (N1473, N1461);
buf BUF1 (N1474, N1472);
and AND2 (N1475, N1452, N354);
nand NAND4 (N1476, N1460, N819, N796, N906);
xor XOR2 (N1477, N1466, N490);
xor XOR2 (N1478, N1465, N1378);
nor NOR3 (N1479, N1473, N790, N284);
and AND4 (N1480, N1476, N249, N922, N1174);
and AND3 (N1481, N1474, N1248, N256);
or OR3 (N1482, N1468, N167, N1348);
nand NAND3 (N1483, N1475, N283, N541);
nor NOR3 (N1484, N1462, N452, N385);
xor XOR2 (N1485, N1464, N1406);
buf BUF1 (N1486, N1484);
nand NAND3 (N1487, N1480, N683, N1097);
and AND4 (N1488, N1479, N746, N1181, N1131);
nor NOR3 (N1489, N1478, N234, N616);
xor XOR2 (N1490, N1488, N1163);
or OR4 (N1491, N1489, N1173, N1062, N1163);
buf BUF1 (N1492, N1486);
buf BUF1 (N1493, N1490);
and AND2 (N1494, N1485, N561);
or OR2 (N1495, N1493, N1091);
buf BUF1 (N1496, N1492);
xor XOR2 (N1497, N1496, N560);
xor XOR2 (N1498, N1494, N800);
or OR2 (N1499, N1471, N1430);
and AND4 (N1500, N1499, N28, N186, N134);
nand NAND3 (N1501, N1482, N649, N582);
xor XOR2 (N1502, N1481, N1226);
or OR2 (N1503, N1501, N561);
xor XOR2 (N1504, N1500, N888);
or OR4 (N1505, N1487, N1050, N837, N227);
buf BUF1 (N1506, N1477);
xor XOR2 (N1507, N1503, N531);
and AND4 (N1508, N1504, N1251, N1066, N503);
nand NAND2 (N1509, N1498, N1047);
and AND4 (N1510, N1507, N711, N1368, N116);
xor XOR2 (N1511, N1509, N486);
and AND4 (N1512, N1497, N13, N672, N258);
or OR4 (N1513, N1491, N1207, N112, N154);
endmodule