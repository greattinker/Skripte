// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N16000,N16005,N16010,N15993,N16011,N16013,N16003,N16001,N15997,N16014;

and AND2 (N15, N13, N14);
xor XOR2 (N16, N1, N2);
not NOT1 (N17, N12);
and AND4 (N18, N15, N15, N16, N5);
xor XOR2 (N19, N14, N16);
buf BUF1 (N20, N1);
or OR4 (N21, N19, N3, N6, N5);
and AND2 (N22, N14, N7);
or OR4 (N23, N19, N3, N13, N13);
and AND4 (N24, N17, N13, N4, N4);
nand NAND2 (N25, N3, N13);
nor NOR3 (N26, N10, N2, N6);
and AND4 (N27, N2, N12, N21, N18);
and AND2 (N28, N1, N16);
not NOT1 (N29, N19);
and AND2 (N30, N1, N28);
nor NOR4 (N31, N11, N1, N13, N23);
buf BUF1 (N32, N1);
xor XOR2 (N33, N24, N4);
buf BUF1 (N34, N29);
nor NOR2 (N35, N32, N11);
buf BUF1 (N36, N33);
not NOT1 (N37, N26);
nand NAND4 (N38, N35, N26, N19, N33);
nor NOR2 (N39, N34, N9);
and AND4 (N40, N22, N23, N2, N10);
nand NAND2 (N41, N40, N26);
or OR2 (N42, N25, N3);
nand NAND2 (N43, N30, N7);
nand NAND2 (N44, N41, N10);
buf BUF1 (N45, N27);
and AND3 (N46, N45, N24, N23);
or OR4 (N47, N36, N39, N27, N28);
and AND4 (N48, N45, N9, N26, N38);
nand NAND2 (N49, N8, N27);
nor NOR3 (N50, N31, N2, N14);
nand NAND4 (N51, N48, N23, N28, N32);
buf BUF1 (N52, N47);
or OR4 (N53, N49, N26, N29, N48);
xor XOR2 (N54, N43, N37);
or OR3 (N55, N23, N1, N4);
xor XOR2 (N56, N50, N16);
or OR2 (N57, N46, N6);
or OR2 (N58, N44, N48);
nand NAND3 (N59, N55, N38, N55);
or OR4 (N60, N59, N40, N14, N12);
nor NOR3 (N61, N51, N3, N3);
xor XOR2 (N62, N52, N4);
nand NAND2 (N63, N60, N58);
nand NAND2 (N64, N4, N35);
not NOT1 (N65, N62);
nand NAND4 (N66, N20, N14, N4, N33);
nand NAND3 (N67, N56, N12, N65);
nand NAND3 (N68, N52, N46, N60);
nand NAND2 (N69, N64, N22);
or OR3 (N70, N68, N55, N61);
xor XOR2 (N71, N56, N19);
buf BUF1 (N72, N42);
and AND2 (N73, N67, N67);
not NOT1 (N74, N72);
nor NOR3 (N75, N66, N64, N52);
nor NOR2 (N76, N75, N42);
nor NOR4 (N77, N74, N48, N57, N73);
nor NOR2 (N78, N18, N28);
nor NOR3 (N79, N11, N7, N50);
buf BUF1 (N80, N69);
xor XOR2 (N81, N78, N66);
and AND2 (N82, N54, N72);
nor NOR2 (N83, N71, N7);
and AND3 (N84, N76, N28, N20);
nand NAND3 (N85, N80, N6, N52);
and AND2 (N86, N81, N43);
or OR4 (N87, N85, N59, N5, N58);
xor XOR2 (N88, N82, N44);
and AND2 (N89, N63, N80);
nand NAND3 (N90, N77, N51, N50);
not NOT1 (N91, N86);
or OR2 (N92, N88, N65);
nor NOR3 (N93, N90, N87, N59);
xor XOR2 (N94, N89, N12);
nand NAND2 (N95, N34, N28);
not NOT1 (N96, N92);
buf BUF1 (N97, N83);
xor XOR2 (N98, N53, N54);
buf BUF1 (N99, N98);
nand NAND2 (N100, N94, N60);
nand NAND2 (N101, N79, N13);
not NOT1 (N102, N97);
not NOT1 (N103, N96);
nand NAND3 (N104, N103, N76, N92);
buf BUF1 (N105, N99);
and AND2 (N106, N101, N10);
nand NAND3 (N107, N104, N77, N19);
and AND2 (N108, N106, N19);
and AND3 (N109, N91, N52, N101);
and AND2 (N110, N100, N43);
buf BUF1 (N111, N107);
buf BUF1 (N112, N102);
xor XOR2 (N113, N109, N111);
xor XOR2 (N114, N14, N39);
or OR4 (N115, N93, N84, N73, N28);
and AND3 (N116, N3, N16, N49);
xor XOR2 (N117, N108, N14);
nor NOR2 (N118, N95, N20);
nor NOR2 (N119, N112, N97);
or OR4 (N120, N117, N65, N84, N87);
not NOT1 (N121, N120);
nand NAND3 (N122, N113, N70, N10);
or OR3 (N123, N68, N46, N104);
nand NAND4 (N124, N119, N42, N38, N89);
nor NOR2 (N125, N116, N114);
xor XOR2 (N126, N50, N58);
nand NAND2 (N127, N126, N9);
nor NOR3 (N128, N125, N60, N24);
nand NAND4 (N129, N124, N19, N57, N90);
buf BUF1 (N130, N110);
and AND3 (N131, N130, N102, N86);
and AND3 (N132, N122, N79, N131);
buf BUF1 (N133, N130);
xor XOR2 (N134, N123, N46);
buf BUF1 (N135, N105);
nand NAND2 (N136, N129, N62);
xor XOR2 (N137, N133, N43);
not NOT1 (N138, N127);
nor NOR2 (N139, N115, N64);
buf BUF1 (N140, N137);
or OR4 (N141, N132, N120, N62, N101);
and AND2 (N142, N140, N62);
buf BUF1 (N143, N135);
nand NAND2 (N144, N138, N76);
and AND3 (N145, N136, N69, N105);
nor NOR2 (N146, N118, N77);
not NOT1 (N147, N128);
or OR4 (N148, N142, N59, N47, N21);
nand NAND2 (N149, N141, N101);
xor XOR2 (N150, N149, N115);
not NOT1 (N151, N144);
not NOT1 (N152, N121);
and AND3 (N153, N145, N21, N58);
xor XOR2 (N154, N146, N13);
nand NAND3 (N155, N143, N143, N132);
and AND3 (N156, N147, N41, N61);
nor NOR3 (N157, N155, N94, N71);
or OR3 (N158, N154, N114, N130);
nand NAND3 (N159, N151, N51, N126);
buf BUF1 (N160, N152);
not NOT1 (N161, N159);
nand NAND3 (N162, N156, N117, N27);
nor NOR3 (N163, N150, N110, N33);
xor XOR2 (N164, N157, N104);
nand NAND2 (N165, N139, N155);
nor NOR2 (N166, N160, N27);
buf BUF1 (N167, N164);
buf BUF1 (N168, N162);
not NOT1 (N169, N166);
or OR4 (N170, N165, N79, N129, N55);
buf BUF1 (N171, N148);
not NOT1 (N172, N171);
xor XOR2 (N173, N161, N6);
or OR2 (N174, N167, N4);
and AND3 (N175, N168, N3, N67);
xor XOR2 (N176, N163, N128);
and AND3 (N177, N172, N65, N119);
buf BUF1 (N178, N177);
buf BUF1 (N179, N175);
nand NAND3 (N180, N178, N158, N121);
buf BUF1 (N181, N41);
nor NOR4 (N182, N134, N18, N93, N76);
buf BUF1 (N183, N153);
and AND4 (N184, N179, N50, N10, N105);
or OR3 (N185, N169, N87, N39);
buf BUF1 (N186, N181);
not NOT1 (N187, N180);
nor NOR3 (N188, N182, N114, N43);
and AND2 (N189, N188, N114);
xor XOR2 (N190, N189, N23);
nand NAND2 (N191, N170, N11);
buf BUF1 (N192, N186);
or OR3 (N193, N190, N44, N108);
nor NOR2 (N194, N193, N20);
nor NOR4 (N195, N192, N188, N119, N171);
or OR4 (N196, N173, N14, N84, N140);
nor NOR3 (N197, N184, N48, N87);
nand NAND2 (N198, N187, N164);
not NOT1 (N199, N198);
and AND3 (N200, N199, N178, N140);
buf BUF1 (N201, N200);
and AND3 (N202, N201, N132, N191);
nand NAND4 (N203, N139, N16, N72, N23);
nor NOR3 (N204, N174, N25, N186);
nor NOR3 (N205, N204, N174, N116);
nor NOR2 (N206, N203, N36);
buf BUF1 (N207, N195);
nand NAND4 (N208, N176, N197, N195, N95);
xor XOR2 (N209, N203, N185);
and AND3 (N210, N200, N105, N109);
nand NAND3 (N211, N194, N46, N169);
and AND3 (N212, N206, N120, N84);
not NOT1 (N213, N209);
xor XOR2 (N214, N208, N127);
xor XOR2 (N215, N210, N208);
nor NOR4 (N216, N212, N213, N48, N70);
buf BUF1 (N217, N78);
xor XOR2 (N218, N183, N26);
nand NAND2 (N219, N205, N186);
nand NAND4 (N220, N215, N77, N200, N39);
buf BUF1 (N221, N218);
xor XOR2 (N222, N216, N112);
not NOT1 (N223, N207);
buf BUF1 (N224, N222);
nor NOR3 (N225, N221, N90, N116);
buf BUF1 (N226, N219);
nor NOR4 (N227, N202, N98, N138, N69);
buf BUF1 (N228, N223);
not NOT1 (N229, N227);
not NOT1 (N230, N225);
nor NOR4 (N231, N224, N152, N89, N72);
nor NOR4 (N232, N217, N35, N80, N161);
xor XOR2 (N233, N226, N175);
and AND4 (N234, N231, N206, N1, N157);
buf BUF1 (N235, N232);
not NOT1 (N236, N214);
xor XOR2 (N237, N220, N152);
buf BUF1 (N238, N211);
or OR4 (N239, N196, N107, N159, N189);
and AND4 (N240, N229, N22, N7, N70);
nand NAND2 (N241, N228, N23);
or OR3 (N242, N241, N22, N63);
nor NOR4 (N243, N240, N230, N33, N112);
not NOT1 (N244, N84);
and AND3 (N245, N233, N148, N215);
not NOT1 (N246, N243);
nor NOR2 (N247, N236, N89);
not NOT1 (N248, N247);
xor XOR2 (N249, N238, N205);
not NOT1 (N250, N249);
and AND4 (N251, N237, N85, N176, N210);
nor NOR3 (N252, N242, N206, N90);
not NOT1 (N253, N235);
or OR4 (N254, N245, N21, N135, N12);
xor XOR2 (N255, N248, N152);
not NOT1 (N256, N239);
nand NAND2 (N257, N251, N113);
and AND2 (N258, N234, N247);
nand NAND3 (N259, N254, N162, N185);
and AND4 (N260, N257, N140, N215, N245);
xor XOR2 (N261, N258, N129);
nor NOR3 (N262, N259, N183, N260);
nand NAND3 (N263, N3, N85, N27);
xor XOR2 (N264, N244, N262);
xor XOR2 (N265, N190, N157);
nor NOR4 (N266, N256, N147, N95, N226);
xor XOR2 (N267, N252, N107);
buf BUF1 (N268, N250);
nor NOR3 (N269, N266, N259, N97);
nor NOR4 (N270, N246, N154, N148, N204);
not NOT1 (N271, N267);
and AND4 (N272, N255, N73, N104, N227);
buf BUF1 (N273, N270);
not NOT1 (N274, N273);
nand NAND4 (N275, N272, N49, N239, N225);
xor XOR2 (N276, N275, N69);
xor XOR2 (N277, N265, N220);
buf BUF1 (N278, N253);
nor NOR3 (N279, N268, N89, N3);
nor NOR3 (N280, N264, N196, N148);
and AND3 (N281, N279, N260, N174);
not NOT1 (N282, N276);
and AND2 (N283, N280, N8);
or OR4 (N284, N263, N239, N209, N230);
or OR4 (N285, N284, N37, N180, N15);
xor XOR2 (N286, N277, N156);
nor NOR2 (N287, N271, N18);
buf BUF1 (N288, N269);
nand NAND3 (N289, N288, N163, N25);
not NOT1 (N290, N289);
nand NAND2 (N291, N274, N246);
or OR3 (N292, N290, N134, N248);
xor XOR2 (N293, N292, N76);
not NOT1 (N294, N281);
nand NAND4 (N295, N285, N212, N151, N278);
nand NAND3 (N296, N246, N279, N78);
nor NOR3 (N297, N291, N28, N257);
or OR4 (N298, N296, N160, N196, N228);
buf BUF1 (N299, N294);
and AND2 (N300, N297, N58);
buf BUF1 (N301, N283);
or OR3 (N302, N295, N82, N14);
and AND4 (N303, N261, N124, N136, N92);
xor XOR2 (N304, N293, N232);
buf BUF1 (N305, N282);
not NOT1 (N306, N301);
buf BUF1 (N307, N299);
nor NOR4 (N308, N303, N210, N139, N291);
buf BUF1 (N309, N286);
or OR4 (N310, N287, N74, N239, N156);
and AND2 (N311, N308, N230);
not NOT1 (N312, N310);
nor NOR2 (N313, N312, N304);
not NOT1 (N314, N193);
nand NAND4 (N315, N313, N164, N247, N74);
or OR2 (N316, N305, N315);
nand NAND2 (N317, N98, N294);
not NOT1 (N318, N298);
and AND4 (N319, N311, N196, N88, N180);
or OR4 (N320, N317, N10, N177, N317);
or OR3 (N321, N318, N302, N46);
nand NAND3 (N322, N104, N185, N13);
and AND2 (N323, N322, N107);
buf BUF1 (N324, N320);
not NOT1 (N325, N319);
xor XOR2 (N326, N323, N51);
buf BUF1 (N327, N309);
nor NOR2 (N328, N321, N240);
buf BUF1 (N329, N328);
and AND4 (N330, N326, N163, N318, N49);
or OR4 (N331, N316, N183, N138, N77);
or OR2 (N332, N300, N288);
nor NOR2 (N333, N325, N31);
nand NAND2 (N334, N327, N323);
xor XOR2 (N335, N334, N300);
not NOT1 (N336, N307);
xor XOR2 (N337, N330, N188);
or OR4 (N338, N337, N26, N45, N262);
nor NOR2 (N339, N324, N54);
nand NAND2 (N340, N332, N338);
nand NAND3 (N341, N230, N200, N270);
not NOT1 (N342, N333);
or OR2 (N343, N306, N110);
nor NOR2 (N344, N314, N331);
and AND3 (N345, N135, N314, N88);
xor XOR2 (N346, N343, N95);
nand NAND2 (N347, N346, N313);
or OR4 (N348, N335, N197, N237, N135);
and AND2 (N349, N345, N84);
or OR4 (N350, N340, N193, N244, N316);
nand NAND4 (N351, N329, N225, N162, N255);
or OR2 (N352, N339, N238);
buf BUF1 (N353, N350);
buf BUF1 (N354, N336);
buf BUF1 (N355, N342);
and AND3 (N356, N351, N112, N46);
nor NOR2 (N357, N348, N32);
xor XOR2 (N358, N355, N314);
buf BUF1 (N359, N352);
xor XOR2 (N360, N356, N246);
nor NOR4 (N361, N344, N203, N67, N351);
nor NOR3 (N362, N361, N80, N288);
xor XOR2 (N363, N349, N217);
buf BUF1 (N364, N357);
or OR2 (N365, N364, N280);
buf BUF1 (N366, N359);
buf BUF1 (N367, N347);
buf BUF1 (N368, N358);
xor XOR2 (N369, N354, N189);
nor NOR3 (N370, N368, N1, N352);
buf BUF1 (N371, N369);
buf BUF1 (N372, N360);
and AND4 (N373, N366, N267, N352, N143);
xor XOR2 (N374, N367, N225);
not NOT1 (N375, N365);
or OR2 (N376, N371, N205);
buf BUF1 (N377, N363);
xor XOR2 (N378, N377, N37);
or OR2 (N379, N375, N369);
xor XOR2 (N380, N378, N366);
nand NAND3 (N381, N372, N336, N108);
nor NOR4 (N382, N362, N378, N183, N369);
nor NOR3 (N383, N341, N258, N255);
buf BUF1 (N384, N376);
xor XOR2 (N385, N373, N308);
nand NAND2 (N386, N381, N250);
nor NOR2 (N387, N382, N96);
xor XOR2 (N388, N384, N123);
buf BUF1 (N389, N353);
and AND2 (N390, N387, N198);
buf BUF1 (N391, N388);
xor XOR2 (N392, N383, N73);
nand NAND4 (N393, N385, N76, N267, N77);
and AND3 (N394, N380, N65, N316);
and AND3 (N395, N386, N61, N171);
nor NOR4 (N396, N391, N115, N17, N101);
nand NAND3 (N397, N374, N288, N59);
nor NOR3 (N398, N396, N227, N187);
not NOT1 (N399, N398);
and AND2 (N400, N397, N234);
xor XOR2 (N401, N394, N262);
or OR2 (N402, N400, N213);
and AND2 (N403, N389, N380);
or OR4 (N404, N390, N258, N200, N31);
buf BUF1 (N405, N401);
and AND4 (N406, N405, N380, N240, N123);
buf BUF1 (N407, N402);
xor XOR2 (N408, N393, N395);
buf BUF1 (N409, N218);
buf BUF1 (N410, N379);
nand NAND4 (N411, N408, N107, N303, N258);
nand NAND4 (N412, N399, N295, N265, N270);
buf BUF1 (N413, N370);
nor NOR4 (N414, N403, N400, N247, N205);
buf BUF1 (N415, N412);
nor NOR3 (N416, N415, N133, N380);
and AND3 (N417, N413, N98, N88);
and AND3 (N418, N404, N375, N141);
nor NOR2 (N419, N392, N41);
not NOT1 (N420, N406);
not NOT1 (N421, N419);
buf BUF1 (N422, N418);
nor NOR4 (N423, N421, N165, N34, N314);
xor XOR2 (N424, N423, N367);
xor XOR2 (N425, N411, N309);
nand NAND2 (N426, N409, N182);
xor XOR2 (N427, N414, N347);
or OR2 (N428, N407, N279);
nand NAND2 (N429, N420, N243);
buf BUF1 (N430, N426);
not NOT1 (N431, N427);
nor NOR4 (N432, N425, N195, N67, N271);
xor XOR2 (N433, N432, N286);
and AND3 (N434, N424, N229, N168);
nand NAND4 (N435, N416, N231, N3, N154);
nand NAND4 (N436, N430, N69, N342, N339);
buf BUF1 (N437, N422);
and AND2 (N438, N417, N301);
xor XOR2 (N439, N428, N422);
nor NOR4 (N440, N438, N212, N417, N325);
nand NAND2 (N441, N433, N388);
nand NAND4 (N442, N434, N168, N60, N289);
nand NAND3 (N443, N440, N129, N209);
nand NAND3 (N444, N443, N15, N396);
nand NAND4 (N445, N429, N190, N274, N160);
nor NOR2 (N446, N444, N189);
buf BUF1 (N447, N441);
not NOT1 (N448, N435);
or OR3 (N449, N410, N322, N290);
not NOT1 (N450, N439);
buf BUF1 (N451, N445);
nand NAND3 (N452, N449, N231, N378);
nand NAND3 (N453, N431, N253, N98);
or OR3 (N454, N446, N101, N238);
nor NOR2 (N455, N436, N179);
not NOT1 (N456, N437);
and AND2 (N457, N454, N195);
nor NOR3 (N458, N456, N379, N421);
nor NOR3 (N459, N453, N393, N289);
and AND2 (N460, N447, N238);
nand NAND2 (N461, N451, N449);
nand NAND3 (N462, N459, N445, N164);
or OR2 (N463, N442, N126);
buf BUF1 (N464, N448);
and AND3 (N465, N464, N405, N163);
not NOT1 (N466, N461);
buf BUF1 (N467, N457);
or OR3 (N468, N455, N148, N72);
xor XOR2 (N469, N450, N85);
buf BUF1 (N470, N468);
not NOT1 (N471, N452);
nor NOR2 (N472, N466, N109);
nand NAND2 (N473, N458, N109);
or OR2 (N474, N472, N331);
xor XOR2 (N475, N474, N473);
not NOT1 (N476, N320);
buf BUF1 (N477, N476);
nand NAND2 (N478, N462, N328);
or OR4 (N479, N467, N152, N81, N196);
and AND3 (N480, N470, N469, N351);
or OR4 (N481, N18, N400, N331, N112);
nor NOR3 (N482, N478, N457, N168);
buf BUF1 (N483, N480);
buf BUF1 (N484, N460);
nor NOR3 (N485, N481, N202, N53);
and AND3 (N486, N483, N460, N318);
xor XOR2 (N487, N475, N196);
buf BUF1 (N488, N479);
not NOT1 (N489, N482);
buf BUF1 (N490, N471);
or OR4 (N491, N489, N96, N93, N9);
not NOT1 (N492, N491);
not NOT1 (N493, N486);
or OR2 (N494, N484, N362);
xor XOR2 (N495, N490, N268);
nor NOR4 (N496, N493, N46, N35, N395);
and AND3 (N497, N496, N233, N239);
nand NAND4 (N498, N487, N20, N47, N144);
not NOT1 (N499, N494);
not NOT1 (N500, N488);
or OR3 (N501, N465, N39, N125);
xor XOR2 (N502, N497, N463);
and AND2 (N503, N222, N338);
buf BUF1 (N504, N499);
and AND3 (N505, N503, N39, N444);
xor XOR2 (N506, N504, N285);
nand NAND2 (N507, N477, N108);
and AND4 (N508, N492, N101, N316, N186);
and AND4 (N509, N495, N366, N11, N52);
xor XOR2 (N510, N506, N117);
xor XOR2 (N511, N505, N396);
nor NOR2 (N512, N500, N188);
nand NAND3 (N513, N512, N102, N391);
xor XOR2 (N514, N498, N481);
xor XOR2 (N515, N485, N396);
nor NOR4 (N516, N510, N121, N35, N221);
xor XOR2 (N517, N508, N487);
buf BUF1 (N518, N502);
xor XOR2 (N519, N511, N188);
or OR3 (N520, N514, N108, N400);
or OR3 (N521, N501, N98, N20);
not NOT1 (N522, N517);
and AND2 (N523, N515, N284);
buf BUF1 (N524, N507);
and AND3 (N525, N523, N200, N502);
nor NOR4 (N526, N521, N222, N159, N415);
not NOT1 (N527, N513);
buf BUF1 (N528, N527);
not NOT1 (N529, N525);
xor XOR2 (N530, N528, N370);
nand NAND2 (N531, N529, N329);
nand NAND2 (N532, N509, N236);
not NOT1 (N533, N526);
buf BUF1 (N534, N530);
nand NAND4 (N535, N519, N455, N459, N111);
nor NOR3 (N536, N518, N528, N483);
not NOT1 (N537, N534);
not NOT1 (N538, N536);
buf BUF1 (N539, N516);
or OR2 (N540, N537, N132);
and AND2 (N541, N532, N133);
buf BUF1 (N542, N539);
nand NAND4 (N543, N535, N123, N497, N358);
or OR2 (N544, N533, N109);
and AND4 (N545, N531, N532, N196, N152);
or OR2 (N546, N538, N524);
buf BUF1 (N547, N271);
buf BUF1 (N548, N542);
nor NOR4 (N549, N548, N243, N95, N187);
xor XOR2 (N550, N522, N57);
buf BUF1 (N551, N541);
buf BUF1 (N552, N544);
xor XOR2 (N553, N550, N66);
not NOT1 (N554, N552);
xor XOR2 (N555, N540, N471);
buf BUF1 (N556, N555);
buf BUF1 (N557, N549);
xor XOR2 (N558, N520, N246);
not NOT1 (N559, N556);
nor NOR3 (N560, N553, N403, N268);
nor NOR4 (N561, N559, N221, N297, N32);
nand NAND4 (N562, N546, N469, N8, N301);
nand NAND4 (N563, N557, N243, N401, N297);
and AND2 (N564, N543, N47);
nor NOR2 (N565, N551, N370);
nor NOR3 (N566, N563, N546, N319);
not NOT1 (N567, N545);
nor NOR2 (N568, N558, N158);
buf BUF1 (N569, N566);
nor NOR2 (N570, N560, N555);
not NOT1 (N571, N568);
buf BUF1 (N572, N562);
xor XOR2 (N573, N570, N474);
not NOT1 (N574, N573);
buf BUF1 (N575, N561);
nor NOR4 (N576, N554, N574, N378, N140);
buf BUF1 (N577, N110);
buf BUF1 (N578, N567);
nor NOR4 (N579, N578, N476, N320, N132);
nand NAND2 (N580, N575, N497);
and AND4 (N581, N565, N500, N314, N29);
and AND4 (N582, N569, N407, N324, N329);
xor XOR2 (N583, N571, N332);
and AND3 (N584, N581, N96, N38);
nor NOR4 (N585, N580, N426, N550, N14);
and AND4 (N586, N576, N157, N469, N325);
buf BUF1 (N587, N585);
buf BUF1 (N588, N579);
or OR3 (N589, N584, N444, N277);
xor XOR2 (N590, N547, N55);
and AND4 (N591, N577, N415, N535, N339);
not NOT1 (N592, N590);
not NOT1 (N593, N587);
or OR3 (N594, N591, N91, N516);
nand NAND2 (N595, N594, N207);
buf BUF1 (N596, N572);
or OR4 (N597, N593, N5, N297, N121);
and AND4 (N598, N592, N118, N136, N99);
not NOT1 (N599, N586);
nand NAND2 (N600, N564, N16);
nor NOR3 (N601, N588, N54, N297);
not NOT1 (N602, N596);
not NOT1 (N603, N595);
and AND3 (N604, N597, N119, N530);
not NOT1 (N605, N604);
xor XOR2 (N606, N589, N187);
and AND3 (N607, N605, N539, N497);
buf BUF1 (N608, N583);
not NOT1 (N609, N606);
buf BUF1 (N610, N602);
and AND4 (N611, N608, N106, N404, N165);
nand NAND3 (N612, N611, N371, N256);
not NOT1 (N613, N599);
nand NAND3 (N614, N601, N103, N442);
nand NAND3 (N615, N614, N148, N411);
buf BUF1 (N616, N582);
nor NOR4 (N617, N607, N556, N332, N134);
nor NOR4 (N618, N603, N499, N104, N358);
or OR2 (N619, N615, N402);
buf BUF1 (N620, N613);
nand NAND3 (N621, N617, N580, N418);
or OR4 (N622, N600, N110, N471, N291);
xor XOR2 (N623, N609, N619);
xor XOR2 (N624, N329, N432);
or OR2 (N625, N623, N359);
buf BUF1 (N626, N598);
nor NOR2 (N627, N624, N565);
nor NOR3 (N628, N616, N125, N71);
buf BUF1 (N629, N622);
not NOT1 (N630, N610);
or OR2 (N631, N630, N6);
or OR2 (N632, N618, N599);
nor NOR2 (N633, N621, N437);
buf BUF1 (N634, N625);
and AND3 (N635, N620, N603, N440);
nand NAND2 (N636, N626, N547);
buf BUF1 (N637, N627);
not NOT1 (N638, N636);
not NOT1 (N639, N635);
and AND4 (N640, N629, N420, N181, N302);
buf BUF1 (N641, N637);
xor XOR2 (N642, N632, N376);
xor XOR2 (N643, N642, N627);
xor XOR2 (N644, N639, N258);
or OR3 (N645, N640, N318, N289);
and AND3 (N646, N631, N638, N400);
not NOT1 (N647, N65);
buf BUF1 (N648, N647);
not NOT1 (N649, N634);
xor XOR2 (N650, N648, N250);
and AND4 (N651, N612, N610, N416, N545);
or OR4 (N652, N650, N294, N274, N61);
xor XOR2 (N653, N645, N454);
not NOT1 (N654, N641);
nand NAND4 (N655, N652, N546, N582, N262);
or OR4 (N656, N633, N537, N524, N115);
not NOT1 (N657, N649);
nand NAND2 (N658, N655, N479);
or OR4 (N659, N653, N356, N618, N207);
xor XOR2 (N660, N646, N525);
buf BUF1 (N661, N654);
nor NOR2 (N662, N659, N578);
or OR3 (N663, N651, N551, N589);
not NOT1 (N664, N660);
xor XOR2 (N665, N664, N622);
not NOT1 (N666, N643);
or OR3 (N667, N661, N328, N296);
xor XOR2 (N668, N657, N566);
nor NOR4 (N669, N662, N478, N126, N411);
xor XOR2 (N670, N658, N125);
not NOT1 (N671, N656);
nor NOR2 (N672, N668, N192);
nand NAND2 (N673, N666, N76);
nor NOR2 (N674, N669, N240);
not NOT1 (N675, N672);
xor XOR2 (N676, N671, N149);
xor XOR2 (N677, N670, N65);
nand NAND3 (N678, N675, N218, N506);
xor XOR2 (N679, N673, N119);
nor NOR3 (N680, N679, N558, N301);
nand NAND2 (N681, N678, N277);
or OR2 (N682, N676, N157);
xor XOR2 (N683, N667, N213);
not NOT1 (N684, N677);
xor XOR2 (N685, N684, N485);
nor NOR4 (N686, N628, N678, N511, N239);
or OR4 (N687, N665, N523, N509, N42);
nand NAND4 (N688, N686, N19, N279, N349);
nand NAND4 (N689, N682, N526, N546, N666);
or OR4 (N690, N663, N267, N127, N246);
nor NOR4 (N691, N683, N343, N583, N77);
buf BUF1 (N692, N689);
nand NAND2 (N693, N688, N276);
xor XOR2 (N694, N690, N582);
not NOT1 (N695, N674);
nor NOR2 (N696, N644, N361);
nor NOR2 (N697, N692, N201);
not NOT1 (N698, N694);
not NOT1 (N699, N698);
nor NOR4 (N700, N695, N226, N137, N479);
nand NAND4 (N701, N680, N611, N467, N253);
nand NAND2 (N702, N681, N604);
or OR2 (N703, N697, N144);
xor XOR2 (N704, N699, N286);
nand NAND3 (N705, N700, N64, N418);
not NOT1 (N706, N703);
and AND3 (N707, N701, N397, N467);
not NOT1 (N708, N706);
and AND4 (N709, N702, N151, N344, N28);
nor NOR2 (N710, N705, N487);
and AND2 (N711, N704, N303);
xor XOR2 (N712, N710, N280);
and AND3 (N713, N685, N592, N335);
not NOT1 (N714, N709);
buf BUF1 (N715, N708);
nand NAND4 (N716, N707, N564, N94, N384);
buf BUF1 (N717, N713);
xor XOR2 (N718, N715, N578);
or OR4 (N719, N711, N107, N148, N192);
xor XOR2 (N720, N718, N692);
buf BUF1 (N721, N714);
nor NOR2 (N722, N693, N379);
buf BUF1 (N723, N720);
nor NOR4 (N724, N712, N134, N122, N266);
not NOT1 (N725, N687);
not NOT1 (N726, N725);
nand NAND4 (N727, N719, N54, N688, N24);
buf BUF1 (N728, N716);
not NOT1 (N729, N723);
xor XOR2 (N730, N726, N387);
nand NAND4 (N731, N717, N186, N526, N183);
not NOT1 (N732, N730);
nand NAND2 (N733, N729, N341);
buf BUF1 (N734, N728);
or OR2 (N735, N732, N236);
nand NAND4 (N736, N731, N477, N679, N186);
and AND2 (N737, N724, N540);
xor XOR2 (N738, N734, N717);
nand NAND2 (N739, N737, N382);
not NOT1 (N740, N739);
and AND3 (N741, N733, N661, N28);
xor XOR2 (N742, N722, N236);
and AND3 (N743, N742, N533, N448);
nor NOR2 (N744, N721, N179);
and AND4 (N745, N740, N601, N319, N166);
nor NOR3 (N746, N744, N553, N132);
buf BUF1 (N747, N696);
or OR4 (N748, N743, N722, N608, N731);
not NOT1 (N749, N745);
nand NAND3 (N750, N749, N366, N321);
and AND2 (N751, N741, N426);
or OR2 (N752, N748, N279);
xor XOR2 (N753, N735, N418);
nand NAND3 (N754, N751, N81, N251);
nor NOR2 (N755, N750, N275);
not NOT1 (N756, N727);
not NOT1 (N757, N746);
and AND3 (N758, N738, N592, N730);
and AND2 (N759, N747, N273);
buf BUF1 (N760, N756);
xor XOR2 (N761, N752, N430);
nand NAND2 (N762, N760, N30);
or OR4 (N763, N759, N281, N100, N179);
xor XOR2 (N764, N757, N341);
not NOT1 (N765, N758);
nand NAND4 (N766, N691, N559, N236, N179);
buf BUF1 (N767, N764);
nor NOR2 (N768, N762, N91);
nor NOR2 (N769, N766, N153);
buf BUF1 (N770, N754);
nand NAND4 (N771, N736, N768, N178, N759);
buf BUF1 (N772, N118);
xor XOR2 (N773, N755, N396);
xor XOR2 (N774, N773, N437);
not NOT1 (N775, N767);
xor XOR2 (N776, N769, N38);
nor NOR4 (N777, N772, N244, N335, N131);
buf BUF1 (N778, N770);
nand NAND2 (N779, N775, N372);
buf BUF1 (N780, N779);
xor XOR2 (N781, N763, N490);
nor NOR4 (N782, N765, N492, N27, N111);
buf BUF1 (N783, N780);
xor XOR2 (N784, N776, N146);
xor XOR2 (N785, N753, N146);
and AND2 (N786, N782, N521);
nand NAND3 (N787, N761, N571, N23);
or OR4 (N788, N774, N490, N748, N652);
and AND4 (N789, N787, N239, N601, N431);
not NOT1 (N790, N784);
or OR3 (N791, N777, N26, N306);
and AND4 (N792, N785, N330, N267, N665);
nor NOR4 (N793, N790, N642, N321, N24);
xor XOR2 (N794, N788, N198);
or OR3 (N795, N791, N434, N445);
not NOT1 (N796, N783);
or OR2 (N797, N771, N154);
nor NOR2 (N798, N778, N699);
xor XOR2 (N799, N795, N789);
or OR4 (N800, N106, N56, N615, N728);
nor NOR3 (N801, N798, N32, N440);
not NOT1 (N802, N792);
nor NOR4 (N803, N801, N764, N634, N318);
xor XOR2 (N804, N794, N397);
or OR3 (N805, N793, N152, N119);
not NOT1 (N806, N786);
xor XOR2 (N807, N803, N581);
nor NOR3 (N808, N804, N76, N568);
and AND3 (N809, N806, N81, N449);
nand NAND2 (N810, N808, N8);
or OR3 (N811, N810, N335, N438);
nand NAND4 (N812, N807, N642, N481, N533);
not NOT1 (N813, N796);
nand NAND2 (N814, N809, N96);
buf BUF1 (N815, N802);
not NOT1 (N816, N797);
not NOT1 (N817, N799);
or OR3 (N818, N815, N579, N163);
nand NAND4 (N819, N805, N798, N171, N385);
buf BUF1 (N820, N814);
buf BUF1 (N821, N811);
xor XOR2 (N822, N816, N572);
buf BUF1 (N823, N781);
xor XOR2 (N824, N823, N81);
and AND2 (N825, N818, N101);
or OR3 (N826, N820, N444, N201);
nor NOR4 (N827, N825, N156, N171, N325);
not NOT1 (N828, N822);
nor NOR2 (N829, N817, N30);
buf BUF1 (N830, N821);
nor NOR2 (N831, N824, N407);
or OR4 (N832, N827, N522, N40, N784);
or OR2 (N833, N829, N732);
and AND2 (N834, N830, N807);
and AND3 (N835, N819, N528, N650);
nand NAND3 (N836, N826, N773, N75);
nand NAND4 (N837, N832, N593, N492, N623);
buf BUF1 (N838, N836);
or OR3 (N839, N833, N803, N375);
xor XOR2 (N840, N828, N228);
nand NAND2 (N841, N835, N836);
nor NOR2 (N842, N834, N54);
or OR2 (N843, N812, N798);
nor NOR4 (N844, N840, N89, N215, N55);
nor NOR4 (N845, N813, N330, N750, N288);
xor XOR2 (N846, N800, N355);
or OR4 (N847, N842, N175, N228, N144);
and AND2 (N848, N846, N24);
buf BUF1 (N849, N831);
or OR4 (N850, N844, N558, N349, N621);
not NOT1 (N851, N849);
or OR4 (N852, N839, N371, N756, N340);
buf BUF1 (N853, N845);
xor XOR2 (N854, N848, N770);
xor XOR2 (N855, N852, N475);
xor XOR2 (N856, N838, N188);
not NOT1 (N857, N837);
nand NAND3 (N858, N843, N390, N99);
or OR3 (N859, N853, N522, N129);
or OR3 (N860, N858, N590, N578);
buf BUF1 (N861, N855);
xor XOR2 (N862, N860, N538);
not NOT1 (N863, N851);
nor NOR3 (N864, N861, N358, N528);
and AND2 (N865, N857, N819);
nor NOR3 (N866, N850, N730, N558);
xor XOR2 (N867, N859, N207);
and AND3 (N868, N864, N784, N38);
or OR4 (N869, N854, N601, N574, N414);
nand NAND2 (N870, N869, N556);
buf BUF1 (N871, N856);
not NOT1 (N872, N841);
nor NOR2 (N873, N871, N319);
xor XOR2 (N874, N863, N316);
nor NOR4 (N875, N847, N507, N678, N764);
nor NOR4 (N876, N872, N364, N586, N478);
not NOT1 (N877, N873);
nor NOR4 (N878, N865, N98, N17, N173);
xor XOR2 (N879, N870, N363);
not NOT1 (N880, N866);
or OR4 (N881, N876, N624, N852, N92);
not NOT1 (N882, N874);
buf BUF1 (N883, N875);
not NOT1 (N884, N882);
nor NOR4 (N885, N881, N43, N173, N539);
buf BUF1 (N886, N879);
buf BUF1 (N887, N886);
nand NAND3 (N888, N868, N623, N745);
not NOT1 (N889, N877);
buf BUF1 (N890, N888);
nand NAND2 (N891, N880, N310);
and AND4 (N892, N883, N645, N287, N150);
not NOT1 (N893, N890);
xor XOR2 (N894, N893, N180);
buf BUF1 (N895, N885);
not NOT1 (N896, N892);
or OR4 (N897, N862, N668, N57, N208);
or OR3 (N898, N867, N717, N271);
buf BUF1 (N899, N898);
xor XOR2 (N900, N899, N832);
xor XOR2 (N901, N887, N748);
xor XOR2 (N902, N894, N226);
nand NAND3 (N903, N902, N258, N662);
xor XOR2 (N904, N889, N359);
and AND2 (N905, N891, N184);
not NOT1 (N906, N895);
or OR2 (N907, N906, N65);
xor XOR2 (N908, N900, N704);
and AND2 (N909, N901, N311);
xor XOR2 (N910, N896, N263);
not NOT1 (N911, N907);
nand NAND3 (N912, N910, N108, N789);
nand NAND2 (N913, N878, N613);
buf BUF1 (N914, N912);
xor XOR2 (N915, N904, N252);
not NOT1 (N916, N914);
nand NAND4 (N917, N908, N512, N592, N696);
or OR4 (N918, N911, N100, N883, N375);
buf BUF1 (N919, N897);
nor NOR3 (N920, N917, N219, N326);
nor NOR2 (N921, N919, N868);
or OR4 (N922, N921, N713, N618, N38);
xor XOR2 (N923, N884, N285);
and AND4 (N924, N903, N376, N180, N418);
buf BUF1 (N925, N916);
xor XOR2 (N926, N905, N347);
buf BUF1 (N927, N925);
nor NOR4 (N928, N913, N9, N860, N169);
and AND2 (N929, N922, N135);
or OR4 (N930, N926, N549, N560, N381);
nand NAND3 (N931, N929, N536, N542);
and AND2 (N932, N931, N463);
or OR4 (N933, N932, N826, N153, N106);
and AND2 (N934, N918, N534);
and AND2 (N935, N915, N590);
nand NAND4 (N936, N928, N752, N711, N807);
xor XOR2 (N937, N927, N769);
nand NAND4 (N938, N923, N907, N844, N559);
and AND2 (N939, N934, N528);
buf BUF1 (N940, N930);
and AND3 (N941, N920, N180, N99);
nor NOR4 (N942, N938, N158, N293, N210);
xor XOR2 (N943, N924, N340);
or OR4 (N944, N936, N301, N211, N490);
xor XOR2 (N945, N933, N553);
xor XOR2 (N946, N909, N337);
buf BUF1 (N947, N945);
and AND2 (N948, N943, N143);
buf BUF1 (N949, N940);
nand NAND3 (N950, N941, N744, N150);
nor NOR3 (N951, N939, N492, N123);
nor NOR3 (N952, N937, N650, N295);
xor XOR2 (N953, N946, N872);
and AND3 (N954, N935, N620, N251);
nand NAND2 (N955, N952, N537);
nand NAND2 (N956, N947, N133);
or OR4 (N957, N949, N462, N559, N931);
nand NAND3 (N958, N942, N767, N799);
and AND2 (N959, N951, N109);
nor NOR2 (N960, N957, N417);
buf BUF1 (N961, N958);
and AND3 (N962, N956, N236, N614);
and AND4 (N963, N953, N591, N408, N209);
buf BUF1 (N964, N948);
nand NAND2 (N965, N944, N707);
not NOT1 (N966, N962);
nor NOR4 (N967, N961, N180, N302, N197);
and AND3 (N968, N960, N456, N955);
not NOT1 (N969, N597);
or OR3 (N970, N963, N888, N411);
or OR3 (N971, N966, N416, N930);
or OR2 (N972, N967, N525);
nand NAND4 (N973, N965, N427, N736, N275);
and AND2 (N974, N950, N524);
nor NOR3 (N975, N954, N805, N686);
or OR2 (N976, N969, N399);
not NOT1 (N977, N973);
and AND3 (N978, N959, N718, N211);
nor NOR4 (N979, N971, N962, N28, N363);
nand NAND4 (N980, N968, N733, N30, N300);
and AND2 (N981, N980, N737);
or OR3 (N982, N976, N151, N249);
not NOT1 (N983, N982);
not NOT1 (N984, N979);
or OR3 (N985, N983, N68, N280);
or OR2 (N986, N981, N269);
or OR4 (N987, N964, N829, N522, N520);
buf BUF1 (N988, N987);
and AND3 (N989, N986, N733, N284);
buf BUF1 (N990, N970);
not NOT1 (N991, N977);
nand NAND4 (N992, N975, N857, N682, N599);
and AND4 (N993, N989, N866, N101, N515);
nor NOR2 (N994, N988, N409);
buf BUF1 (N995, N992);
or OR3 (N996, N974, N635, N112);
and AND4 (N997, N972, N450, N130, N187);
not NOT1 (N998, N996);
nand NAND2 (N999, N990, N674);
buf BUF1 (N1000, N995);
buf BUF1 (N1001, N985);
nand NAND3 (N1002, N1000, N446, N387);
nor NOR2 (N1003, N978, N636);
xor XOR2 (N1004, N1001, N45);
buf BUF1 (N1005, N994);
or OR3 (N1006, N998, N837, N472);
nor NOR3 (N1007, N993, N452, N872);
not NOT1 (N1008, N1005);
xor XOR2 (N1009, N997, N153);
and AND2 (N1010, N1003, N668);
nand NAND4 (N1011, N1002, N908, N360, N815);
nor NOR4 (N1012, N984, N593, N878, N169);
not NOT1 (N1013, N1009);
nand NAND3 (N1014, N991, N448, N535);
xor XOR2 (N1015, N1008, N732);
nor NOR4 (N1016, N1014, N857, N92, N302);
buf BUF1 (N1017, N1015);
xor XOR2 (N1018, N1013, N236);
buf BUF1 (N1019, N1011);
nand NAND2 (N1020, N1017, N970);
nor NOR4 (N1021, N1012, N740, N710, N544);
and AND2 (N1022, N1021, N213);
nor NOR4 (N1023, N1010, N746, N815, N37);
nand NAND2 (N1024, N1016, N105);
not NOT1 (N1025, N999);
nor NOR2 (N1026, N1007, N567);
and AND4 (N1027, N1006, N792, N365, N58);
xor XOR2 (N1028, N1027, N899);
and AND3 (N1029, N1025, N658, N3);
nand NAND3 (N1030, N1019, N534, N390);
or OR4 (N1031, N1024, N465, N739, N953);
buf BUF1 (N1032, N1023);
nand NAND2 (N1033, N1004, N406);
buf BUF1 (N1034, N1022);
buf BUF1 (N1035, N1031);
nand NAND2 (N1036, N1028, N135);
and AND2 (N1037, N1032, N971);
buf BUF1 (N1038, N1018);
or OR4 (N1039, N1020, N229, N498, N529);
buf BUF1 (N1040, N1026);
or OR3 (N1041, N1037, N1026, N352);
buf BUF1 (N1042, N1033);
nor NOR3 (N1043, N1034, N324, N787);
xor XOR2 (N1044, N1038, N831);
nor NOR3 (N1045, N1042, N571, N895);
not NOT1 (N1046, N1029);
nand NAND3 (N1047, N1044, N183, N533);
xor XOR2 (N1048, N1043, N367);
and AND3 (N1049, N1035, N875, N476);
buf BUF1 (N1050, N1049);
nand NAND3 (N1051, N1040, N259, N766);
nor NOR3 (N1052, N1048, N143, N938);
buf BUF1 (N1053, N1030);
not NOT1 (N1054, N1036);
xor XOR2 (N1055, N1050, N929);
nand NAND3 (N1056, N1053, N793, N815);
nand NAND3 (N1057, N1039, N529, N827);
buf BUF1 (N1058, N1054);
nand NAND3 (N1059, N1056, N128, N263);
or OR2 (N1060, N1041, N305);
buf BUF1 (N1061, N1045);
and AND3 (N1062, N1055, N884, N73);
and AND2 (N1063, N1062, N757);
buf BUF1 (N1064, N1051);
buf BUF1 (N1065, N1052);
xor XOR2 (N1066, N1063, N698);
and AND2 (N1067, N1066, N343);
nor NOR2 (N1068, N1058, N660);
and AND4 (N1069, N1060, N562, N383, N293);
buf BUF1 (N1070, N1065);
nand NAND3 (N1071, N1070, N1058, N45);
not NOT1 (N1072, N1071);
nand NAND2 (N1073, N1072, N213);
buf BUF1 (N1074, N1064);
or OR2 (N1075, N1068, N792);
buf BUF1 (N1076, N1069);
nor NOR3 (N1077, N1057, N187, N1030);
xor XOR2 (N1078, N1074, N171);
buf BUF1 (N1079, N1078);
nand NAND2 (N1080, N1077, N3);
and AND2 (N1081, N1061, N721);
nand NAND2 (N1082, N1081, N735);
not NOT1 (N1083, N1059);
xor XOR2 (N1084, N1079, N507);
not NOT1 (N1085, N1073);
nand NAND4 (N1086, N1075, N964, N849, N277);
buf BUF1 (N1087, N1082);
or OR2 (N1088, N1080, N797);
not NOT1 (N1089, N1084);
buf BUF1 (N1090, N1046);
xor XOR2 (N1091, N1067, N463);
xor XOR2 (N1092, N1089, N788);
and AND2 (N1093, N1086, N124);
nand NAND4 (N1094, N1091, N371, N928, N956);
xor XOR2 (N1095, N1047, N230);
xor XOR2 (N1096, N1085, N782);
or OR2 (N1097, N1096, N7);
nand NAND2 (N1098, N1076, N426);
or OR2 (N1099, N1097, N653);
nand NAND4 (N1100, N1092, N226, N917, N66);
xor XOR2 (N1101, N1093, N438);
nand NAND3 (N1102, N1088, N157, N703);
nand NAND4 (N1103, N1102, N521, N300, N453);
buf BUF1 (N1104, N1098);
and AND3 (N1105, N1100, N273, N262);
xor XOR2 (N1106, N1099, N672);
nor NOR4 (N1107, N1090, N1063, N23, N33);
xor XOR2 (N1108, N1107, N464);
and AND2 (N1109, N1095, N645);
and AND3 (N1110, N1101, N598, N83);
and AND4 (N1111, N1083, N514, N601, N638);
or OR3 (N1112, N1087, N1052, N143);
nor NOR4 (N1113, N1112, N852, N901, N542);
buf BUF1 (N1114, N1110);
not NOT1 (N1115, N1094);
not NOT1 (N1116, N1104);
not NOT1 (N1117, N1103);
nand NAND2 (N1118, N1111, N172);
xor XOR2 (N1119, N1113, N47);
nor NOR2 (N1120, N1109, N819);
xor XOR2 (N1121, N1117, N368);
xor XOR2 (N1122, N1120, N727);
buf BUF1 (N1123, N1116);
or OR3 (N1124, N1123, N566, N258);
and AND2 (N1125, N1108, N719);
not NOT1 (N1126, N1124);
buf BUF1 (N1127, N1119);
nand NAND2 (N1128, N1127, N367);
xor XOR2 (N1129, N1115, N79);
xor XOR2 (N1130, N1105, N664);
or OR4 (N1131, N1114, N269, N863, N756);
not NOT1 (N1132, N1129);
nand NAND3 (N1133, N1126, N821, N832);
nor NOR3 (N1134, N1106, N781, N484);
nor NOR4 (N1135, N1130, N9, N1087, N550);
nand NAND4 (N1136, N1128, N326, N368, N803);
not NOT1 (N1137, N1121);
nand NAND3 (N1138, N1132, N36, N1117);
and AND2 (N1139, N1118, N473);
or OR4 (N1140, N1135, N313, N351, N247);
and AND4 (N1141, N1131, N897, N1031, N454);
nand NAND3 (N1142, N1136, N690, N1034);
xor XOR2 (N1143, N1137, N961);
and AND4 (N1144, N1133, N985, N318, N198);
and AND3 (N1145, N1140, N984, N326);
buf BUF1 (N1146, N1145);
and AND4 (N1147, N1125, N901, N617, N459);
not NOT1 (N1148, N1143);
xor XOR2 (N1149, N1148, N1092);
xor XOR2 (N1150, N1139, N42);
and AND3 (N1151, N1122, N218, N598);
xor XOR2 (N1152, N1151, N1023);
nor NOR2 (N1153, N1149, N846);
nand NAND3 (N1154, N1147, N675, N336);
and AND3 (N1155, N1146, N216, N855);
and AND4 (N1156, N1142, N908, N651, N132);
nand NAND2 (N1157, N1134, N1062);
buf BUF1 (N1158, N1155);
xor XOR2 (N1159, N1158, N559);
xor XOR2 (N1160, N1159, N114);
or OR2 (N1161, N1138, N8);
nor NOR2 (N1162, N1157, N482);
or OR3 (N1163, N1160, N441, N1035);
and AND3 (N1164, N1144, N331, N490);
nor NOR2 (N1165, N1161, N723);
nor NOR4 (N1166, N1141, N711, N228, N739);
or OR2 (N1167, N1156, N728);
nor NOR3 (N1168, N1166, N486, N948);
nand NAND3 (N1169, N1165, N357, N1081);
nand NAND2 (N1170, N1169, N851);
or OR4 (N1171, N1152, N764, N681, N987);
nor NOR3 (N1172, N1153, N836, N828);
and AND3 (N1173, N1162, N388, N529);
nor NOR3 (N1174, N1170, N986, N263);
nand NAND2 (N1175, N1163, N266);
nor NOR2 (N1176, N1175, N501);
nor NOR2 (N1177, N1174, N253);
or OR3 (N1178, N1168, N958, N724);
nand NAND3 (N1179, N1176, N504, N734);
nor NOR2 (N1180, N1164, N167);
nor NOR2 (N1181, N1171, N687);
buf BUF1 (N1182, N1177);
or OR4 (N1183, N1182, N245, N68, N1104);
nor NOR3 (N1184, N1167, N195, N697);
nor NOR3 (N1185, N1172, N33, N923);
nor NOR4 (N1186, N1183, N51, N773, N1052);
not NOT1 (N1187, N1179);
buf BUF1 (N1188, N1178);
nor NOR3 (N1189, N1187, N807, N276);
or OR4 (N1190, N1184, N1113, N516, N1149);
not NOT1 (N1191, N1189);
xor XOR2 (N1192, N1181, N1007);
not NOT1 (N1193, N1192);
not NOT1 (N1194, N1186);
and AND2 (N1195, N1188, N143);
or OR3 (N1196, N1194, N935, N693);
and AND3 (N1197, N1154, N641, N366);
or OR4 (N1198, N1195, N804, N207, N35);
or OR4 (N1199, N1196, N1001, N1190, N386);
buf BUF1 (N1200, N679);
not NOT1 (N1201, N1197);
xor XOR2 (N1202, N1185, N1079);
and AND4 (N1203, N1173, N885, N366, N1192);
nor NOR4 (N1204, N1198, N1203, N691, N465);
buf BUF1 (N1205, N523);
nor NOR2 (N1206, N1180, N1107);
or OR3 (N1207, N1191, N671, N760);
and AND4 (N1208, N1150, N1083, N1, N477);
xor XOR2 (N1209, N1202, N1038);
or OR3 (N1210, N1209, N992, N975);
and AND3 (N1211, N1206, N639, N1030);
or OR4 (N1212, N1201, N610, N994, N128);
not NOT1 (N1213, N1205);
not NOT1 (N1214, N1193);
not NOT1 (N1215, N1211);
buf BUF1 (N1216, N1215);
nor NOR3 (N1217, N1207, N1043, N389);
nor NOR2 (N1218, N1208, N699);
buf BUF1 (N1219, N1217);
nand NAND4 (N1220, N1218, N534, N217, N1189);
not NOT1 (N1221, N1213);
and AND4 (N1222, N1204, N73, N244, N296);
nand NAND4 (N1223, N1210, N976, N9, N650);
nor NOR3 (N1224, N1223, N928, N1109);
not NOT1 (N1225, N1212);
xor XOR2 (N1226, N1199, N520);
not NOT1 (N1227, N1214);
and AND3 (N1228, N1220, N1057, N718);
nand NAND2 (N1229, N1222, N606);
not NOT1 (N1230, N1224);
not NOT1 (N1231, N1228);
nand NAND2 (N1232, N1227, N81);
or OR2 (N1233, N1216, N671);
not NOT1 (N1234, N1231);
not NOT1 (N1235, N1229);
nor NOR3 (N1236, N1225, N571, N884);
nor NOR3 (N1237, N1219, N1037, N4);
xor XOR2 (N1238, N1237, N899);
xor XOR2 (N1239, N1234, N394);
not NOT1 (N1240, N1221);
buf BUF1 (N1241, N1238);
or OR4 (N1242, N1226, N441, N1158, N1204);
xor XOR2 (N1243, N1235, N490);
buf BUF1 (N1244, N1240);
or OR4 (N1245, N1243, N171, N1128, N507);
nor NOR2 (N1246, N1200, N784);
or OR4 (N1247, N1241, N1241, N1034, N1231);
nor NOR3 (N1248, N1236, N494, N80);
buf BUF1 (N1249, N1239);
not NOT1 (N1250, N1248);
xor XOR2 (N1251, N1230, N1191);
nand NAND4 (N1252, N1249, N1199, N358, N157);
not NOT1 (N1253, N1244);
nand NAND4 (N1254, N1253, N861, N186, N868);
nor NOR2 (N1255, N1251, N915);
and AND2 (N1256, N1247, N126);
not NOT1 (N1257, N1254);
buf BUF1 (N1258, N1255);
xor XOR2 (N1259, N1252, N279);
nor NOR3 (N1260, N1242, N311, N1209);
nor NOR2 (N1261, N1232, N929);
not NOT1 (N1262, N1258);
nor NOR2 (N1263, N1245, N972);
buf BUF1 (N1264, N1260);
xor XOR2 (N1265, N1246, N915);
not NOT1 (N1266, N1233);
nor NOR3 (N1267, N1266, N1199, N1200);
or OR4 (N1268, N1263, N1241, N883, N925);
or OR3 (N1269, N1264, N970, N603);
and AND2 (N1270, N1269, N440);
nor NOR4 (N1271, N1270, N1149, N522, N768);
or OR4 (N1272, N1256, N828, N570, N342);
or OR4 (N1273, N1272, N1045, N1090, N168);
nand NAND2 (N1274, N1262, N1251);
xor XOR2 (N1275, N1273, N1212);
and AND4 (N1276, N1265, N1170, N913, N630);
nor NOR3 (N1277, N1261, N268, N574);
or OR3 (N1278, N1250, N581, N808);
xor XOR2 (N1279, N1278, N1197);
and AND3 (N1280, N1275, N628, N397);
nand NAND3 (N1281, N1274, N385, N191);
xor XOR2 (N1282, N1280, N542);
nand NAND2 (N1283, N1282, N391);
and AND3 (N1284, N1279, N910, N98);
buf BUF1 (N1285, N1276);
and AND3 (N1286, N1284, N910, N278);
nor NOR4 (N1287, N1259, N134, N154, N78);
nand NAND3 (N1288, N1281, N268, N1183);
nand NAND2 (N1289, N1285, N866);
and AND4 (N1290, N1286, N226, N392, N512);
nor NOR2 (N1291, N1267, N528);
nor NOR2 (N1292, N1290, N13);
xor XOR2 (N1293, N1287, N756);
buf BUF1 (N1294, N1283);
xor XOR2 (N1295, N1292, N237);
not NOT1 (N1296, N1277);
nor NOR2 (N1297, N1257, N28);
or OR2 (N1298, N1289, N925);
buf BUF1 (N1299, N1298);
xor XOR2 (N1300, N1268, N1167);
or OR3 (N1301, N1291, N865, N649);
nand NAND4 (N1302, N1294, N53, N935, N863);
xor XOR2 (N1303, N1297, N307);
not NOT1 (N1304, N1293);
or OR3 (N1305, N1296, N1259, N867);
xor XOR2 (N1306, N1288, N920);
nor NOR3 (N1307, N1306, N706, N947);
xor XOR2 (N1308, N1271, N308);
or OR2 (N1309, N1295, N771);
buf BUF1 (N1310, N1304);
xor XOR2 (N1311, N1310, N910);
nor NOR3 (N1312, N1301, N1208, N950);
and AND2 (N1313, N1308, N599);
nor NOR3 (N1314, N1307, N273, N1049);
and AND2 (N1315, N1313, N216);
xor XOR2 (N1316, N1303, N892);
or OR2 (N1317, N1305, N1312);
not NOT1 (N1318, N110);
xor XOR2 (N1319, N1314, N874);
nor NOR2 (N1320, N1315, N610);
or OR4 (N1321, N1318, N287, N1160, N1198);
or OR4 (N1322, N1299, N613, N465, N1276);
xor XOR2 (N1323, N1302, N732);
and AND2 (N1324, N1300, N162);
xor XOR2 (N1325, N1323, N258);
buf BUF1 (N1326, N1309);
nor NOR3 (N1327, N1326, N9, N1132);
not NOT1 (N1328, N1325);
buf BUF1 (N1329, N1320);
not NOT1 (N1330, N1319);
not NOT1 (N1331, N1317);
buf BUF1 (N1332, N1327);
nand NAND3 (N1333, N1316, N378, N542);
buf BUF1 (N1334, N1330);
not NOT1 (N1335, N1311);
not NOT1 (N1336, N1331);
not NOT1 (N1337, N1332);
and AND2 (N1338, N1329, N1264);
nor NOR4 (N1339, N1336, N44, N347, N1315);
xor XOR2 (N1340, N1322, N637);
nor NOR4 (N1341, N1328, N851, N318, N793);
nand NAND3 (N1342, N1339, N643, N1163);
not NOT1 (N1343, N1337);
or OR4 (N1344, N1333, N749, N121, N1197);
nor NOR2 (N1345, N1344, N1014);
or OR2 (N1346, N1334, N412);
or OR4 (N1347, N1345, N1278, N394, N1325);
or OR4 (N1348, N1343, N1108, N928, N642);
xor XOR2 (N1349, N1338, N1164);
nand NAND3 (N1350, N1341, N1304, N688);
xor XOR2 (N1351, N1324, N1011);
nand NAND2 (N1352, N1349, N690);
nand NAND2 (N1353, N1346, N1275);
nand NAND4 (N1354, N1348, N174, N906, N193);
not NOT1 (N1355, N1350);
xor XOR2 (N1356, N1354, N37);
and AND2 (N1357, N1321, N452);
or OR3 (N1358, N1342, N820, N1356);
buf BUF1 (N1359, N24);
nor NOR3 (N1360, N1359, N1282, N1263);
xor XOR2 (N1361, N1360, N844);
nor NOR3 (N1362, N1347, N962, N207);
buf BUF1 (N1363, N1362);
buf BUF1 (N1364, N1351);
xor XOR2 (N1365, N1353, N216);
and AND4 (N1366, N1340, N509, N1279, N942);
nand NAND2 (N1367, N1357, N446);
nor NOR2 (N1368, N1355, N891);
xor XOR2 (N1369, N1367, N379);
nand NAND3 (N1370, N1365, N955, N426);
nor NOR2 (N1371, N1352, N223);
buf BUF1 (N1372, N1371);
or OR2 (N1373, N1369, N537);
or OR2 (N1374, N1363, N265);
xor XOR2 (N1375, N1364, N201);
and AND4 (N1376, N1374, N1083, N337, N907);
xor XOR2 (N1377, N1366, N716);
nand NAND2 (N1378, N1375, N516);
not NOT1 (N1379, N1361);
buf BUF1 (N1380, N1376);
nor NOR2 (N1381, N1370, N353);
xor XOR2 (N1382, N1368, N1064);
nor NOR3 (N1383, N1372, N55, N135);
nand NAND4 (N1384, N1377, N530, N354, N1262);
and AND4 (N1385, N1335, N1046, N17, N275);
buf BUF1 (N1386, N1379);
or OR2 (N1387, N1382, N1108);
nor NOR2 (N1388, N1378, N681);
or OR4 (N1389, N1373, N551, N923, N1204);
or OR2 (N1390, N1386, N1361);
buf BUF1 (N1391, N1388);
not NOT1 (N1392, N1380);
and AND3 (N1393, N1383, N307, N809);
and AND2 (N1394, N1389, N784);
buf BUF1 (N1395, N1394);
nand NAND3 (N1396, N1358, N540, N1247);
xor XOR2 (N1397, N1381, N648);
xor XOR2 (N1398, N1397, N945);
and AND4 (N1399, N1396, N208, N611, N522);
or OR3 (N1400, N1395, N496, N7);
or OR4 (N1401, N1398, N1339, N183, N764);
or OR3 (N1402, N1399, N1344, N695);
nand NAND3 (N1403, N1400, N1251, N818);
xor XOR2 (N1404, N1403, N415);
xor XOR2 (N1405, N1385, N501);
not NOT1 (N1406, N1392);
or OR2 (N1407, N1405, N485);
and AND4 (N1408, N1387, N1332, N48, N603);
nand NAND2 (N1409, N1390, N263);
buf BUF1 (N1410, N1401);
xor XOR2 (N1411, N1384, N868);
not NOT1 (N1412, N1408);
not NOT1 (N1413, N1409);
nor NOR4 (N1414, N1412, N1382, N266, N491);
and AND2 (N1415, N1414, N146);
xor XOR2 (N1416, N1407, N1338);
nand NAND4 (N1417, N1391, N1378, N842, N1179);
nand NAND4 (N1418, N1406, N748, N618, N128);
buf BUF1 (N1419, N1393);
xor XOR2 (N1420, N1415, N1331);
and AND3 (N1421, N1416, N324, N448);
nand NAND2 (N1422, N1419, N276);
nand NAND4 (N1423, N1420, N112, N1379, N302);
not NOT1 (N1424, N1410);
and AND4 (N1425, N1423, N601, N25, N1334);
or OR4 (N1426, N1411, N708, N772, N204);
xor XOR2 (N1427, N1402, N1002);
nor NOR3 (N1428, N1418, N844, N1288);
nor NOR4 (N1429, N1427, N336, N584, N311);
not NOT1 (N1430, N1428);
buf BUF1 (N1431, N1424);
buf BUF1 (N1432, N1413);
xor XOR2 (N1433, N1425, N1081);
xor XOR2 (N1434, N1430, N818);
buf BUF1 (N1435, N1434);
xor XOR2 (N1436, N1435, N131);
nand NAND2 (N1437, N1422, N367);
or OR4 (N1438, N1429, N1228, N503, N921);
or OR4 (N1439, N1417, N33, N438, N1225);
nand NAND2 (N1440, N1439, N1436);
buf BUF1 (N1441, N350);
or OR4 (N1442, N1431, N175, N956, N419);
nand NAND3 (N1443, N1421, N868, N1266);
buf BUF1 (N1444, N1432);
xor XOR2 (N1445, N1440, N1393);
nor NOR3 (N1446, N1433, N18, N503);
buf BUF1 (N1447, N1441);
not NOT1 (N1448, N1444);
or OR4 (N1449, N1442, N1180, N1312, N272);
nor NOR4 (N1450, N1437, N885, N1050, N740);
or OR2 (N1451, N1446, N1430);
and AND2 (N1452, N1426, N110);
not NOT1 (N1453, N1438);
xor XOR2 (N1454, N1451, N1276);
buf BUF1 (N1455, N1450);
and AND3 (N1456, N1453, N1084, N1159);
not NOT1 (N1457, N1445);
not NOT1 (N1458, N1449);
and AND4 (N1459, N1458, N405, N498, N1008);
not NOT1 (N1460, N1459);
buf BUF1 (N1461, N1460);
nand NAND2 (N1462, N1452, N733);
or OR4 (N1463, N1447, N321, N508, N1040);
and AND3 (N1464, N1454, N1375, N744);
xor XOR2 (N1465, N1456, N639);
buf BUF1 (N1466, N1455);
buf BUF1 (N1467, N1466);
or OR4 (N1468, N1443, N832, N898, N1257);
or OR4 (N1469, N1448, N1418, N917, N408);
or OR4 (N1470, N1469, N781, N1131, N974);
or OR4 (N1471, N1467, N247, N181, N233);
and AND2 (N1472, N1465, N619);
and AND4 (N1473, N1462, N1448, N1424, N1278);
nor NOR3 (N1474, N1468, N866, N1095);
not NOT1 (N1475, N1474);
or OR2 (N1476, N1470, N506);
not NOT1 (N1477, N1473);
xor XOR2 (N1478, N1463, N277);
nor NOR2 (N1479, N1475, N395);
buf BUF1 (N1480, N1477);
and AND3 (N1481, N1478, N1173, N329);
nor NOR3 (N1482, N1404, N443, N1077);
nand NAND2 (N1483, N1461, N167);
nand NAND4 (N1484, N1476, N1437, N664, N960);
buf BUF1 (N1485, N1464);
not NOT1 (N1486, N1457);
and AND4 (N1487, N1482, N1408, N932, N963);
and AND4 (N1488, N1480, N1132, N1445, N579);
not NOT1 (N1489, N1481);
xor XOR2 (N1490, N1486, N381);
xor XOR2 (N1491, N1471, N794);
nand NAND2 (N1492, N1489, N669);
and AND2 (N1493, N1492, N598);
nand NAND4 (N1494, N1483, N1127, N311, N26);
buf BUF1 (N1495, N1472);
not NOT1 (N1496, N1495);
and AND4 (N1497, N1494, N228, N761, N372);
xor XOR2 (N1498, N1488, N103);
xor XOR2 (N1499, N1484, N1042);
not NOT1 (N1500, N1487);
not NOT1 (N1501, N1497);
nor NOR2 (N1502, N1498, N1047);
not NOT1 (N1503, N1499);
nand NAND2 (N1504, N1501, N689);
xor XOR2 (N1505, N1504, N1188);
nor NOR3 (N1506, N1479, N384, N1459);
buf BUF1 (N1507, N1500);
buf BUF1 (N1508, N1490);
nor NOR3 (N1509, N1507, N1185, N895);
xor XOR2 (N1510, N1503, N799);
buf BUF1 (N1511, N1485);
buf BUF1 (N1512, N1510);
nand NAND2 (N1513, N1508, N36);
xor XOR2 (N1514, N1506, N1146);
buf BUF1 (N1515, N1502);
buf BUF1 (N1516, N1511);
nand NAND3 (N1517, N1491, N544, N285);
xor XOR2 (N1518, N1517, N884);
buf BUF1 (N1519, N1516);
nor NOR2 (N1520, N1519, N982);
nor NOR4 (N1521, N1513, N123, N870, N492);
buf BUF1 (N1522, N1496);
buf BUF1 (N1523, N1521);
xor XOR2 (N1524, N1505, N917);
not NOT1 (N1525, N1515);
not NOT1 (N1526, N1523);
and AND3 (N1527, N1525, N197, N260);
or OR4 (N1528, N1518, N1167, N536, N1007);
nor NOR4 (N1529, N1524, N225, N707, N462);
or OR3 (N1530, N1529, N1452, N121);
nand NAND4 (N1531, N1514, N317, N127, N390);
nand NAND2 (N1532, N1520, N633);
buf BUF1 (N1533, N1532);
and AND2 (N1534, N1526, N148);
nand NAND3 (N1535, N1533, N449, N1404);
nand NAND2 (N1536, N1534, N76);
or OR4 (N1537, N1535, N1465, N219, N681);
and AND3 (N1538, N1509, N1456, N243);
or OR2 (N1539, N1512, N1345);
nand NAND3 (N1540, N1522, N1514, N1263);
buf BUF1 (N1541, N1527);
or OR2 (N1542, N1539, N829);
not NOT1 (N1543, N1537);
nand NAND3 (N1544, N1542, N481, N322);
xor XOR2 (N1545, N1530, N1295);
nor NOR3 (N1546, N1493, N697, N991);
nand NAND3 (N1547, N1538, N625, N956);
nand NAND2 (N1548, N1540, N920);
xor XOR2 (N1549, N1548, N884);
nor NOR2 (N1550, N1544, N782);
not NOT1 (N1551, N1549);
and AND2 (N1552, N1547, N659);
or OR3 (N1553, N1531, N893, N490);
nand NAND3 (N1554, N1551, N1450, N355);
and AND4 (N1555, N1554, N501, N927, N433);
nor NOR4 (N1556, N1553, N393, N558, N795);
nor NOR4 (N1557, N1550, N1106, N1290, N885);
nand NAND3 (N1558, N1541, N698, N62);
or OR2 (N1559, N1556, N217);
and AND3 (N1560, N1557, N1536, N76);
not NOT1 (N1561, N749);
nand NAND2 (N1562, N1558, N215);
xor XOR2 (N1563, N1528, N336);
nor NOR2 (N1564, N1561, N1352);
nor NOR2 (N1565, N1560, N1095);
buf BUF1 (N1566, N1559);
not NOT1 (N1567, N1543);
buf BUF1 (N1568, N1564);
xor XOR2 (N1569, N1568, N548);
or OR2 (N1570, N1569, N1525);
xor XOR2 (N1571, N1567, N221);
nand NAND4 (N1572, N1562, N1346, N1489, N1267);
or OR2 (N1573, N1572, N1074);
xor XOR2 (N1574, N1573, N409);
not NOT1 (N1575, N1563);
nand NAND2 (N1576, N1566, N190);
buf BUF1 (N1577, N1576);
or OR2 (N1578, N1545, N598);
nor NOR2 (N1579, N1571, N976);
xor XOR2 (N1580, N1555, N1509);
or OR4 (N1581, N1546, N1031, N395, N1020);
not NOT1 (N1582, N1580);
and AND4 (N1583, N1552, N1147, N161, N1569);
or OR2 (N1584, N1575, N771);
nand NAND2 (N1585, N1574, N186);
or OR4 (N1586, N1582, N474, N787, N285);
buf BUF1 (N1587, N1578);
nor NOR3 (N1588, N1581, N155, N638);
nand NAND4 (N1589, N1579, N81, N527, N1028);
or OR3 (N1590, N1588, N29, N309);
xor XOR2 (N1591, N1590, N1360);
nand NAND3 (N1592, N1583, N1303, N246);
buf BUF1 (N1593, N1577);
and AND3 (N1594, N1592, N950, N479);
and AND3 (N1595, N1565, N664, N520);
and AND4 (N1596, N1591, N1088, N677, N717);
nor NOR2 (N1597, N1593, N1029);
not NOT1 (N1598, N1589);
buf BUF1 (N1599, N1586);
or OR3 (N1600, N1570, N183, N768);
not NOT1 (N1601, N1598);
or OR2 (N1602, N1597, N1298);
buf BUF1 (N1603, N1595);
xor XOR2 (N1604, N1601, N1398);
nor NOR2 (N1605, N1585, N1329);
buf BUF1 (N1606, N1596);
buf BUF1 (N1607, N1594);
nor NOR2 (N1608, N1607, N1025);
and AND2 (N1609, N1608, N870);
and AND4 (N1610, N1609, N833, N1224, N10);
buf BUF1 (N1611, N1603);
nand NAND2 (N1612, N1599, N843);
xor XOR2 (N1613, N1602, N1100);
or OR2 (N1614, N1611, N723);
or OR2 (N1615, N1614, N1408);
buf BUF1 (N1616, N1606);
or OR4 (N1617, N1584, N706, N1519, N708);
xor XOR2 (N1618, N1612, N299);
or OR3 (N1619, N1617, N650, N339);
nand NAND4 (N1620, N1605, N566, N632, N779);
buf BUF1 (N1621, N1613);
not NOT1 (N1622, N1620);
not NOT1 (N1623, N1621);
not NOT1 (N1624, N1616);
or OR4 (N1625, N1623, N830, N1371, N1172);
and AND3 (N1626, N1619, N1536, N385);
xor XOR2 (N1627, N1618, N544);
or OR4 (N1628, N1610, N1455, N1004, N60);
and AND4 (N1629, N1625, N79, N483, N1500);
xor XOR2 (N1630, N1600, N1530);
or OR3 (N1631, N1604, N406, N601);
xor XOR2 (N1632, N1624, N555);
nor NOR2 (N1633, N1587, N71);
or OR3 (N1634, N1629, N381, N14);
or OR4 (N1635, N1615, N20, N1500, N372);
and AND4 (N1636, N1626, N434, N1324, N477);
buf BUF1 (N1637, N1622);
nor NOR3 (N1638, N1637, N633, N201);
or OR2 (N1639, N1631, N1324);
or OR2 (N1640, N1634, N1142);
xor XOR2 (N1641, N1639, N429);
and AND2 (N1642, N1630, N1620);
nand NAND2 (N1643, N1632, N1359);
or OR4 (N1644, N1633, N1065, N803, N1057);
nor NOR3 (N1645, N1628, N636, N101);
nand NAND4 (N1646, N1627, N540, N1441, N293);
or OR2 (N1647, N1643, N667);
nand NAND2 (N1648, N1642, N300);
not NOT1 (N1649, N1635);
buf BUF1 (N1650, N1646);
not NOT1 (N1651, N1641);
and AND3 (N1652, N1636, N99, N1034);
or OR4 (N1653, N1645, N655, N1123, N122);
nand NAND4 (N1654, N1640, N823, N316, N1634);
nor NOR2 (N1655, N1649, N667);
nor NOR4 (N1656, N1647, N458, N327, N1186);
and AND2 (N1657, N1651, N607);
not NOT1 (N1658, N1655);
not NOT1 (N1659, N1652);
and AND3 (N1660, N1650, N534, N133);
xor XOR2 (N1661, N1654, N1133);
or OR3 (N1662, N1660, N1109, N1318);
xor XOR2 (N1663, N1653, N1225);
buf BUF1 (N1664, N1662);
not NOT1 (N1665, N1663);
or OR4 (N1666, N1656, N635, N168, N799);
or OR4 (N1667, N1661, N1156, N824, N1282);
not NOT1 (N1668, N1664);
xor XOR2 (N1669, N1657, N1243);
xor XOR2 (N1670, N1648, N526);
not NOT1 (N1671, N1658);
nand NAND2 (N1672, N1670, N391);
and AND4 (N1673, N1644, N367, N272, N893);
nor NOR3 (N1674, N1669, N1093, N123);
buf BUF1 (N1675, N1638);
and AND2 (N1676, N1665, N933);
and AND2 (N1677, N1671, N1442);
xor XOR2 (N1678, N1673, N340);
and AND2 (N1679, N1666, N998);
nand NAND4 (N1680, N1675, N1242, N905, N1048);
or OR4 (N1681, N1667, N1642, N1050, N1240);
buf BUF1 (N1682, N1668);
xor XOR2 (N1683, N1679, N1345);
nor NOR2 (N1684, N1672, N140);
or OR4 (N1685, N1680, N172, N574, N1014);
nor NOR3 (N1686, N1676, N444, N1492);
nor NOR4 (N1687, N1677, N1267, N301, N699);
buf BUF1 (N1688, N1687);
nand NAND4 (N1689, N1686, N1326, N682, N844);
or OR2 (N1690, N1683, N1677);
nor NOR4 (N1691, N1688, N186, N1095, N727);
not NOT1 (N1692, N1659);
nand NAND3 (N1693, N1674, N1297, N267);
not NOT1 (N1694, N1681);
buf BUF1 (N1695, N1690);
xor XOR2 (N1696, N1692, N1540);
nor NOR2 (N1697, N1693, N1459);
nor NOR2 (N1698, N1695, N174);
and AND4 (N1699, N1694, N742, N337, N1058);
xor XOR2 (N1700, N1684, N1235);
buf BUF1 (N1701, N1697);
nor NOR2 (N1702, N1691, N1357);
or OR3 (N1703, N1702, N263, N291);
nor NOR4 (N1704, N1701, N1575, N697, N1692);
nand NAND2 (N1705, N1678, N112);
buf BUF1 (N1706, N1698);
nor NOR3 (N1707, N1703, N517, N355);
or OR4 (N1708, N1685, N1062, N1094, N1517);
buf BUF1 (N1709, N1699);
nand NAND3 (N1710, N1689, N552, N933);
and AND2 (N1711, N1709, N1254);
nor NOR4 (N1712, N1700, N360, N283, N1198);
nand NAND4 (N1713, N1708, N1654, N1516, N1613);
buf BUF1 (N1714, N1696);
or OR4 (N1715, N1704, N944, N130, N868);
nor NOR4 (N1716, N1713, N1483, N24, N555);
xor XOR2 (N1717, N1712, N1113);
buf BUF1 (N1718, N1710);
buf BUF1 (N1719, N1716);
or OR2 (N1720, N1715, N118);
or OR3 (N1721, N1719, N418, N814);
or OR2 (N1722, N1718, N1052);
buf BUF1 (N1723, N1706);
buf BUF1 (N1724, N1714);
buf BUF1 (N1725, N1724);
nor NOR4 (N1726, N1723, N351, N99, N1247);
not NOT1 (N1727, N1707);
nand NAND4 (N1728, N1721, N887, N570, N422);
nand NAND2 (N1729, N1682, N567);
nand NAND3 (N1730, N1729, N421, N1476);
xor XOR2 (N1731, N1727, N1395);
or OR2 (N1732, N1711, N1074);
nand NAND2 (N1733, N1731, N1581);
or OR2 (N1734, N1720, N679);
nand NAND4 (N1735, N1734, N113, N1578, N1651);
not NOT1 (N1736, N1728);
xor XOR2 (N1737, N1725, N1700);
nand NAND2 (N1738, N1737, N297);
not NOT1 (N1739, N1717);
xor XOR2 (N1740, N1738, N1646);
buf BUF1 (N1741, N1735);
nand NAND4 (N1742, N1740, N1736, N682, N126);
and AND3 (N1743, N58, N253, N1566);
not NOT1 (N1744, N1742);
buf BUF1 (N1745, N1739);
buf BUF1 (N1746, N1743);
buf BUF1 (N1747, N1733);
or OR2 (N1748, N1744, N1535);
not NOT1 (N1749, N1746);
and AND3 (N1750, N1726, N135, N886);
not NOT1 (N1751, N1730);
nand NAND4 (N1752, N1722, N1220, N167, N1661);
or OR3 (N1753, N1732, N1738, N1019);
xor XOR2 (N1754, N1741, N494);
xor XOR2 (N1755, N1752, N566);
xor XOR2 (N1756, N1753, N279);
or OR4 (N1757, N1747, N236, N1199, N1462);
nor NOR3 (N1758, N1750, N1568, N826);
nor NOR3 (N1759, N1754, N1118, N219);
buf BUF1 (N1760, N1759);
and AND3 (N1761, N1751, N459, N1006);
nand NAND4 (N1762, N1745, N1379, N1051, N1120);
not NOT1 (N1763, N1755);
xor XOR2 (N1764, N1756, N1461);
nor NOR4 (N1765, N1749, N1642, N123, N1451);
and AND3 (N1766, N1761, N116, N1431);
and AND4 (N1767, N1757, N1413, N1263, N831);
xor XOR2 (N1768, N1765, N290);
or OR3 (N1769, N1758, N704, N851);
buf BUF1 (N1770, N1768);
not NOT1 (N1771, N1762);
xor XOR2 (N1772, N1767, N540);
nand NAND3 (N1773, N1770, N960, N1276);
and AND2 (N1774, N1748, N1290);
not NOT1 (N1775, N1705);
nand NAND3 (N1776, N1774, N972, N1317);
nand NAND2 (N1777, N1775, N995);
or OR3 (N1778, N1773, N1160, N787);
or OR3 (N1779, N1777, N1342, N1072);
nor NOR3 (N1780, N1764, N879, N1142);
nor NOR4 (N1781, N1771, N670, N613, N482);
nand NAND3 (N1782, N1763, N732, N31);
not NOT1 (N1783, N1780);
buf BUF1 (N1784, N1782);
buf BUF1 (N1785, N1769);
xor XOR2 (N1786, N1784, N1456);
and AND2 (N1787, N1783, N1354);
not NOT1 (N1788, N1776);
not NOT1 (N1789, N1786);
nand NAND2 (N1790, N1772, N332);
buf BUF1 (N1791, N1788);
nand NAND3 (N1792, N1789, N1450, N1755);
nand NAND3 (N1793, N1779, N860, N526);
nand NAND4 (N1794, N1778, N35, N1497, N1155);
and AND4 (N1795, N1781, N1430, N1302, N1091);
nor NOR4 (N1796, N1795, N569, N485, N1190);
or OR2 (N1797, N1793, N257);
nor NOR4 (N1798, N1790, N1133, N352, N811);
not NOT1 (N1799, N1792);
nor NOR3 (N1800, N1794, N827, N1733);
nor NOR4 (N1801, N1800, N313, N1590, N393);
xor XOR2 (N1802, N1787, N64);
nand NAND2 (N1803, N1766, N849);
and AND2 (N1804, N1797, N1194);
nand NAND2 (N1805, N1791, N364);
and AND2 (N1806, N1760, N22);
xor XOR2 (N1807, N1798, N1552);
and AND3 (N1808, N1804, N106, N1414);
and AND2 (N1809, N1803, N675);
nand NAND4 (N1810, N1802, N959, N1427, N757);
not NOT1 (N1811, N1807);
and AND2 (N1812, N1801, N267);
buf BUF1 (N1813, N1805);
nor NOR3 (N1814, N1813, N607, N1791);
nor NOR2 (N1815, N1812, N749);
nor NOR4 (N1816, N1808, N253, N855, N588);
buf BUF1 (N1817, N1814);
not NOT1 (N1818, N1810);
or OR2 (N1819, N1799, N511);
xor XOR2 (N1820, N1811, N1230);
buf BUF1 (N1821, N1817);
not NOT1 (N1822, N1820);
nor NOR3 (N1823, N1818, N827, N1093);
or OR4 (N1824, N1823, N534, N786, N921);
buf BUF1 (N1825, N1816);
and AND2 (N1826, N1815, N782);
xor XOR2 (N1827, N1822, N1535);
buf BUF1 (N1828, N1825);
buf BUF1 (N1829, N1806);
nand NAND2 (N1830, N1824, N1337);
or OR4 (N1831, N1809, N343, N367, N472);
or OR2 (N1832, N1826, N1354);
and AND4 (N1833, N1785, N277, N950, N677);
or OR4 (N1834, N1830, N90, N1114, N950);
nor NOR3 (N1835, N1829, N1600, N1394);
not NOT1 (N1836, N1828);
nand NAND4 (N1837, N1833, N1623, N1565, N1142);
nand NAND4 (N1838, N1819, N1408, N1470, N1239);
buf BUF1 (N1839, N1831);
buf BUF1 (N1840, N1827);
not NOT1 (N1841, N1837);
xor XOR2 (N1842, N1832, N34);
nor NOR2 (N1843, N1796, N1637);
nor NOR3 (N1844, N1839, N1372, N969);
nor NOR4 (N1845, N1821, N1773, N201, N3);
not NOT1 (N1846, N1842);
nor NOR4 (N1847, N1843, N55, N256, N220);
nor NOR2 (N1848, N1835, N43);
and AND2 (N1849, N1834, N667);
and AND3 (N1850, N1848, N488, N1212);
xor XOR2 (N1851, N1844, N1506);
xor XOR2 (N1852, N1841, N972);
or OR4 (N1853, N1838, N475, N298, N1657);
not NOT1 (N1854, N1850);
nand NAND4 (N1855, N1847, N863, N629, N1402);
or OR2 (N1856, N1836, N1545);
buf BUF1 (N1857, N1855);
and AND3 (N1858, N1857, N1172, N1358);
not NOT1 (N1859, N1854);
xor XOR2 (N1860, N1856, N243);
not NOT1 (N1861, N1853);
nand NAND3 (N1862, N1846, N422, N418);
nor NOR4 (N1863, N1852, N81, N1170, N1204);
xor XOR2 (N1864, N1862, N503);
xor XOR2 (N1865, N1863, N149);
not NOT1 (N1866, N1858);
nor NOR4 (N1867, N1851, N1641, N909, N1628);
or OR2 (N1868, N1860, N1634);
or OR4 (N1869, N1865, N1674, N476, N230);
xor XOR2 (N1870, N1869, N1099);
and AND4 (N1871, N1870, N968, N304, N1504);
xor XOR2 (N1872, N1871, N1242);
and AND4 (N1873, N1849, N1430, N1007, N1771);
and AND4 (N1874, N1864, N1414, N1850, N1147);
or OR4 (N1875, N1845, N1102, N1310, N1044);
and AND3 (N1876, N1867, N1010, N1515);
nor NOR4 (N1877, N1840, N826, N1487, N1695);
nor NOR2 (N1878, N1874, N1769);
xor XOR2 (N1879, N1866, N1249);
nor NOR4 (N1880, N1875, N5, N622, N1009);
buf BUF1 (N1881, N1868);
buf BUF1 (N1882, N1876);
or OR3 (N1883, N1877, N1858, N1882);
nor NOR3 (N1884, N694, N1042, N1264);
nor NOR4 (N1885, N1884, N1487, N1211, N1724);
not NOT1 (N1886, N1881);
buf BUF1 (N1887, N1859);
nor NOR4 (N1888, N1878, N266, N1110, N501);
buf BUF1 (N1889, N1888);
not NOT1 (N1890, N1879);
and AND2 (N1891, N1890, N603);
nand NAND4 (N1892, N1889, N978, N871, N919);
xor XOR2 (N1893, N1885, N1706);
and AND4 (N1894, N1873, N140, N588, N1389);
not NOT1 (N1895, N1886);
nand NAND2 (N1896, N1872, N1777);
or OR4 (N1897, N1880, N423, N429, N265);
nor NOR4 (N1898, N1861, N1608, N1659, N672);
or OR3 (N1899, N1892, N801, N244);
buf BUF1 (N1900, N1898);
and AND4 (N1901, N1896, N1043, N1005, N199);
nor NOR3 (N1902, N1895, N1748, N1365);
and AND4 (N1903, N1900, N226, N808, N1292);
nand NAND3 (N1904, N1894, N94, N1246);
nand NAND3 (N1905, N1901, N290, N383);
nand NAND3 (N1906, N1883, N1088, N524);
nor NOR3 (N1907, N1897, N1125, N1160);
and AND4 (N1908, N1893, N612, N1066, N1797);
or OR3 (N1909, N1887, N52, N323);
and AND2 (N1910, N1891, N6);
not NOT1 (N1911, N1910);
and AND2 (N1912, N1899, N25);
and AND2 (N1913, N1912, N1477);
xor XOR2 (N1914, N1907, N928);
and AND3 (N1915, N1909, N1701, N862);
nor NOR4 (N1916, N1913, N1663, N1728, N123);
or OR4 (N1917, N1905, N622, N1353, N1831);
buf BUF1 (N1918, N1908);
and AND4 (N1919, N1903, N729, N1468, N309);
and AND4 (N1920, N1902, N1288, N871, N239);
not NOT1 (N1921, N1916);
buf BUF1 (N1922, N1921);
and AND3 (N1923, N1906, N1580, N594);
nor NOR2 (N1924, N1923, N1413);
and AND3 (N1925, N1917, N942, N1673);
nand NAND2 (N1926, N1925, N1378);
xor XOR2 (N1927, N1911, N366);
nand NAND2 (N1928, N1927, N748);
or OR3 (N1929, N1919, N1474, N1347);
xor XOR2 (N1930, N1918, N652);
and AND3 (N1931, N1928, N964, N1296);
xor XOR2 (N1932, N1931, N1542);
buf BUF1 (N1933, N1932);
nand NAND4 (N1934, N1920, N1152, N1771, N1784);
not NOT1 (N1935, N1930);
buf BUF1 (N1936, N1933);
not NOT1 (N1937, N1924);
or OR2 (N1938, N1922, N1390);
buf BUF1 (N1939, N1934);
not NOT1 (N1940, N1936);
buf BUF1 (N1941, N1929);
xor XOR2 (N1942, N1939, N646);
nand NAND3 (N1943, N1938, N1919, N252);
xor XOR2 (N1944, N1926, N1243);
xor XOR2 (N1945, N1940, N1739);
not NOT1 (N1946, N1942);
xor XOR2 (N1947, N1943, N1172);
nand NAND2 (N1948, N1945, N448);
nand NAND2 (N1949, N1915, N337);
nand NAND3 (N1950, N1947, N1131, N589);
nor NOR2 (N1951, N1904, N1552);
xor XOR2 (N1952, N1937, N1776);
buf BUF1 (N1953, N1944);
and AND4 (N1954, N1941, N1161, N1498, N1371);
nand NAND2 (N1955, N1951, N991);
nor NOR2 (N1956, N1953, N508);
nor NOR4 (N1957, N1935, N1521, N221, N908);
and AND4 (N1958, N1955, N71, N555, N1160);
and AND2 (N1959, N1946, N1068);
nand NAND4 (N1960, N1948, N675, N1151, N1307);
nand NAND3 (N1961, N1960, N970, N1434);
not NOT1 (N1962, N1956);
and AND4 (N1963, N1949, N1800, N1109, N1597);
or OR2 (N1964, N1952, N875);
nor NOR2 (N1965, N1957, N27);
buf BUF1 (N1966, N1961);
and AND4 (N1967, N1914, N537, N1822, N970);
not NOT1 (N1968, N1962);
and AND3 (N1969, N1959, N156, N1625);
or OR2 (N1970, N1969, N1696);
or OR3 (N1971, N1958, N804, N1090);
xor XOR2 (N1972, N1954, N1734);
buf BUF1 (N1973, N1968);
not NOT1 (N1974, N1950);
xor XOR2 (N1975, N1973, N944);
nor NOR2 (N1976, N1963, N937);
not NOT1 (N1977, N1970);
nand NAND2 (N1978, N1964, N1441);
nor NOR4 (N1979, N1965, N1643, N1772, N1947);
or OR2 (N1980, N1977, N1662);
nor NOR3 (N1981, N1974, N978, N95);
not NOT1 (N1982, N1967);
nor NOR2 (N1983, N1976, N536);
nor NOR4 (N1984, N1975, N103, N803, N83);
and AND2 (N1985, N1980, N130);
nor NOR4 (N1986, N1978, N1733, N474, N746);
xor XOR2 (N1987, N1979, N286);
nor NOR3 (N1988, N1987, N1016, N1978);
and AND3 (N1989, N1982, N1732, N355);
xor XOR2 (N1990, N1988, N1778);
nor NOR4 (N1991, N1989, N44, N586, N1043);
not NOT1 (N1992, N1984);
or OR4 (N1993, N1992, N372, N769, N28);
xor XOR2 (N1994, N1971, N886);
nand NAND4 (N1995, N1966, N1244, N1394, N1414);
not NOT1 (N1996, N1993);
or OR4 (N1997, N1985, N1375, N438, N923);
not NOT1 (N1998, N1981);
nand NAND2 (N1999, N1990, N862);
nand NAND4 (N2000, N1972, N1547, N81, N953);
buf BUF1 (N2001, N1986);
buf BUF1 (N2002, N1997);
and AND4 (N2003, N2002, N498, N1877, N707);
buf BUF1 (N2004, N1983);
nand NAND3 (N2005, N1999, N422, N2000);
xor XOR2 (N2006, N1731, N72);
or OR2 (N2007, N1996, N1045);
and AND3 (N2008, N1998, N84, N1981);
and AND2 (N2009, N1995, N1738);
nand NAND2 (N2010, N2006, N1890);
not NOT1 (N2011, N1994);
xor XOR2 (N2012, N2009, N1299);
and AND4 (N2013, N2008, N762, N1520, N1037);
and AND2 (N2014, N2004, N1607);
or OR3 (N2015, N2003, N1039, N1825);
nand NAND4 (N2016, N1991, N1842, N1394, N242);
or OR2 (N2017, N2011, N454);
nor NOR2 (N2018, N2001, N1646);
or OR4 (N2019, N2010, N987, N1192, N1469);
and AND4 (N2020, N2005, N1018, N1427, N1577);
not NOT1 (N2021, N2012);
or OR4 (N2022, N2013, N1137, N1751, N1928);
or OR3 (N2023, N2022, N1057, N1182);
nand NAND3 (N2024, N2020, N1917, N14);
nand NAND2 (N2025, N2015, N248);
not NOT1 (N2026, N2018);
buf BUF1 (N2027, N2024);
or OR3 (N2028, N2014, N775, N1984);
not NOT1 (N2029, N2019);
buf BUF1 (N2030, N2026);
or OR2 (N2031, N2023, N1784);
nand NAND2 (N2032, N2027, N715);
not NOT1 (N2033, N2025);
nand NAND3 (N2034, N2030, N481, N1643);
or OR3 (N2035, N2017, N2014, N993);
not NOT1 (N2036, N2007);
or OR3 (N2037, N2035, N1766, N1123);
buf BUF1 (N2038, N2016);
and AND4 (N2039, N2028, N87, N394, N1656);
buf BUF1 (N2040, N2037);
or OR4 (N2041, N2033, N1828, N962, N521);
xor XOR2 (N2042, N2021, N662);
or OR4 (N2043, N2031, N10, N257, N1376);
buf BUF1 (N2044, N2041);
xor XOR2 (N2045, N2039, N1729);
xor XOR2 (N2046, N2040, N857);
buf BUF1 (N2047, N2046);
nand NAND3 (N2048, N2045, N1516, N1286);
and AND4 (N2049, N2032, N1837, N1668, N1349);
and AND3 (N2050, N2036, N396, N525);
or OR4 (N2051, N2047, N527, N1695, N175);
or OR2 (N2052, N2029, N1092);
xor XOR2 (N2053, N2044, N1091);
or OR2 (N2054, N2051, N1703);
nand NAND4 (N2055, N2054, N1200, N1309, N579);
xor XOR2 (N2056, N2042, N666);
nor NOR4 (N2057, N2038, N1581, N1123, N1525);
nand NAND3 (N2058, N2053, N1844, N2031);
buf BUF1 (N2059, N2050);
not NOT1 (N2060, N2043);
not NOT1 (N2061, N2052);
and AND4 (N2062, N2059, N517, N167, N1813);
not NOT1 (N2063, N2034);
nand NAND2 (N2064, N2058, N384);
buf BUF1 (N2065, N2048);
buf BUF1 (N2066, N2063);
not NOT1 (N2067, N2049);
buf BUF1 (N2068, N2064);
and AND4 (N2069, N2055, N1078, N1066, N425);
nor NOR2 (N2070, N2065, N1047);
not NOT1 (N2071, N2060);
nand NAND3 (N2072, N2070, N501, N712);
and AND3 (N2073, N2057, N1253, N358);
not NOT1 (N2074, N2061);
nand NAND4 (N2075, N2074, N2034, N229, N1272);
nand NAND2 (N2076, N2075, N2069);
or OR4 (N2077, N944, N342, N1804, N192);
not NOT1 (N2078, N2073);
or OR3 (N2079, N2068, N185, N947);
nand NAND2 (N2080, N2062, N1821);
or OR4 (N2081, N2071, N1356, N2048, N1489);
nand NAND4 (N2082, N2080, N179, N306, N1172);
not NOT1 (N2083, N2082);
or OR3 (N2084, N2083, N1070, N1055);
buf BUF1 (N2085, N2078);
nand NAND3 (N2086, N2085, N2040, N438);
and AND3 (N2087, N2072, N1713, N1817);
or OR3 (N2088, N2056, N658, N1201);
nand NAND3 (N2089, N2086, N935, N531);
nand NAND3 (N2090, N2089, N325, N1512);
not NOT1 (N2091, N2081);
buf BUF1 (N2092, N2077);
buf BUF1 (N2093, N2088);
not NOT1 (N2094, N2087);
nor NOR4 (N2095, N2092, N32, N295, N1717);
buf BUF1 (N2096, N2066);
and AND2 (N2097, N2093, N431);
and AND3 (N2098, N2079, N498, N129);
nand NAND4 (N2099, N2091, N865, N16, N247);
xor XOR2 (N2100, N2094, N1670);
xor XOR2 (N2101, N2095, N581);
nand NAND2 (N2102, N2076, N1747);
buf BUF1 (N2103, N2090);
xor XOR2 (N2104, N2084, N1880);
and AND3 (N2105, N2104, N346, N1432);
xor XOR2 (N2106, N2067, N1148);
nor NOR2 (N2107, N2100, N1250);
and AND2 (N2108, N2102, N710);
and AND2 (N2109, N2103, N722);
not NOT1 (N2110, N2101);
nor NOR4 (N2111, N2096, N240, N259, N797);
nor NOR4 (N2112, N2106, N120, N502, N1835);
xor XOR2 (N2113, N2097, N927);
nand NAND2 (N2114, N2099, N926);
nor NOR3 (N2115, N2107, N1409, N158);
not NOT1 (N2116, N2105);
nor NOR2 (N2117, N2098, N1897);
xor XOR2 (N2118, N2117, N463);
buf BUF1 (N2119, N2115);
nand NAND4 (N2120, N2108, N1972, N566, N1398);
xor XOR2 (N2121, N2111, N1159);
nand NAND4 (N2122, N2116, N363, N921, N246);
nand NAND2 (N2123, N2109, N1338);
and AND2 (N2124, N2114, N593);
and AND3 (N2125, N2118, N1257, N682);
not NOT1 (N2126, N2119);
nor NOR2 (N2127, N2112, N1127);
buf BUF1 (N2128, N2121);
or OR2 (N2129, N2120, N1967);
xor XOR2 (N2130, N2129, N907);
buf BUF1 (N2131, N2122);
not NOT1 (N2132, N2123);
nand NAND4 (N2133, N2113, N1775, N1205, N80);
nor NOR4 (N2134, N2110, N624, N1542, N499);
nand NAND2 (N2135, N2127, N1487);
and AND3 (N2136, N2132, N966, N1732);
and AND3 (N2137, N2124, N2013, N2087);
nor NOR3 (N2138, N2131, N1825, N1183);
xor XOR2 (N2139, N2133, N1345);
nor NOR2 (N2140, N2136, N1067);
nand NAND3 (N2141, N2130, N1342, N1188);
nand NAND4 (N2142, N2135, N406, N1683, N340);
not NOT1 (N2143, N2139);
not NOT1 (N2144, N2134);
not NOT1 (N2145, N2143);
nor NOR2 (N2146, N2142, N1869);
nand NAND2 (N2147, N2146, N1416);
buf BUF1 (N2148, N2138);
nand NAND2 (N2149, N2147, N557);
or OR4 (N2150, N2126, N1910, N1189, N194);
or OR4 (N2151, N2137, N1681, N1659, N943);
xor XOR2 (N2152, N2149, N1566);
nand NAND2 (N2153, N2150, N1093);
not NOT1 (N2154, N2152);
nor NOR4 (N2155, N2145, N559, N316, N611);
nor NOR2 (N2156, N2148, N140);
not NOT1 (N2157, N2151);
nor NOR4 (N2158, N2156, N549, N649, N1178);
or OR4 (N2159, N2125, N1625, N1119, N1389);
xor XOR2 (N2160, N2159, N861);
xor XOR2 (N2161, N2158, N1307);
xor XOR2 (N2162, N2140, N541);
nor NOR2 (N2163, N2128, N657);
or OR4 (N2164, N2153, N370, N1958, N359);
buf BUF1 (N2165, N2160);
buf BUF1 (N2166, N2165);
nor NOR4 (N2167, N2164, N1794, N972, N382);
buf BUF1 (N2168, N2157);
xor XOR2 (N2169, N2166, N253);
xor XOR2 (N2170, N2163, N699);
buf BUF1 (N2171, N2155);
xor XOR2 (N2172, N2167, N980);
nand NAND4 (N2173, N2144, N860, N441, N253);
buf BUF1 (N2174, N2172);
nand NAND2 (N2175, N2161, N2153);
xor XOR2 (N2176, N2141, N970);
xor XOR2 (N2177, N2174, N323);
xor XOR2 (N2178, N2168, N1251);
xor XOR2 (N2179, N2175, N997);
xor XOR2 (N2180, N2178, N146);
and AND3 (N2181, N2180, N945, N1595);
or OR2 (N2182, N2162, N44);
and AND2 (N2183, N2173, N739);
buf BUF1 (N2184, N2154);
not NOT1 (N2185, N2171);
xor XOR2 (N2186, N2185, N339);
xor XOR2 (N2187, N2186, N2092);
xor XOR2 (N2188, N2183, N617);
buf BUF1 (N2189, N2170);
buf BUF1 (N2190, N2181);
xor XOR2 (N2191, N2190, N1131);
nor NOR2 (N2192, N2182, N386);
xor XOR2 (N2193, N2192, N1125);
or OR4 (N2194, N2193, N1626, N640, N537);
xor XOR2 (N2195, N2169, N1205);
nand NAND3 (N2196, N2191, N825, N188);
nand NAND4 (N2197, N2187, N1416, N1855, N591);
not NOT1 (N2198, N2176);
nand NAND4 (N2199, N2184, N930, N1472, N1616);
not NOT1 (N2200, N2197);
buf BUF1 (N2201, N2177);
nor NOR3 (N2202, N2200, N1672, N51);
xor XOR2 (N2203, N2199, N988);
buf BUF1 (N2204, N2194);
and AND2 (N2205, N2201, N1178);
xor XOR2 (N2206, N2203, N527);
or OR2 (N2207, N2179, N2158);
buf BUF1 (N2208, N2202);
not NOT1 (N2209, N2196);
nor NOR2 (N2210, N2207, N2126);
nand NAND2 (N2211, N2206, N1424);
or OR2 (N2212, N2195, N1758);
not NOT1 (N2213, N2211);
or OR4 (N2214, N2212, N1254, N495, N734);
or OR3 (N2215, N2205, N1077, N708);
not NOT1 (N2216, N2215);
and AND4 (N2217, N2204, N1176, N865, N1889);
nor NOR4 (N2218, N2188, N1852, N13, N682);
not NOT1 (N2219, N2218);
or OR2 (N2220, N2219, N262);
buf BUF1 (N2221, N2213);
nand NAND2 (N2222, N2210, N1406);
and AND4 (N2223, N2189, N1384, N2197, N89);
buf BUF1 (N2224, N2216);
not NOT1 (N2225, N2208);
buf BUF1 (N2226, N2221);
buf BUF1 (N2227, N2226);
nand NAND4 (N2228, N2214, N198, N1075, N1920);
and AND4 (N2229, N2228, N1825, N818, N763);
xor XOR2 (N2230, N2229, N1501);
and AND3 (N2231, N2222, N19, N1474);
not NOT1 (N2232, N2230);
nor NOR4 (N2233, N2217, N1625, N2179, N1305);
and AND3 (N2234, N2225, N796, N1293);
or OR2 (N2235, N2227, N336);
or OR2 (N2236, N2231, N428);
xor XOR2 (N2237, N2224, N1235);
and AND2 (N2238, N2209, N598);
nor NOR2 (N2239, N2235, N894);
xor XOR2 (N2240, N2234, N1488);
not NOT1 (N2241, N2239);
nand NAND2 (N2242, N2220, N1954);
or OR4 (N2243, N2238, N711, N1703, N1530);
nand NAND2 (N2244, N2233, N197);
or OR2 (N2245, N2236, N938);
and AND4 (N2246, N2223, N525, N1894, N68);
nand NAND3 (N2247, N2232, N2072, N431);
buf BUF1 (N2248, N2198);
xor XOR2 (N2249, N2241, N967);
nor NOR2 (N2250, N2242, N195);
nor NOR4 (N2251, N2245, N1920, N1392, N2083);
xor XOR2 (N2252, N2237, N1505);
nor NOR4 (N2253, N2240, N1860, N2003, N544);
and AND3 (N2254, N2244, N28, N504);
buf BUF1 (N2255, N2252);
buf BUF1 (N2256, N2247);
nor NOR3 (N2257, N2251, N1015, N1395);
xor XOR2 (N2258, N2246, N1440);
and AND4 (N2259, N2258, N2156, N1164, N1866);
xor XOR2 (N2260, N2250, N75);
xor XOR2 (N2261, N2243, N1511);
nor NOR3 (N2262, N2255, N62, N2061);
not NOT1 (N2263, N2261);
xor XOR2 (N2264, N2256, N1478);
xor XOR2 (N2265, N2259, N1385);
and AND2 (N2266, N2263, N1203);
and AND2 (N2267, N2260, N1724);
and AND2 (N2268, N2249, N613);
not NOT1 (N2269, N2265);
nand NAND2 (N2270, N2253, N769);
buf BUF1 (N2271, N2268);
buf BUF1 (N2272, N2267);
xor XOR2 (N2273, N2264, N1289);
xor XOR2 (N2274, N2257, N2128);
not NOT1 (N2275, N2266);
and AND3 (N2276, N2271, N1051, N1705);
buf BUF1 (N2277, N2262);
buf BUF1 (N2278, N2275);
and AND2 (N2279, N2277, N1549);
xor XOR2 (N2280, N2278, N1694);
nor NOR4 (N2281, N2248, N807, N551, N1415);
or OR4 (N2282, N2280, N1858, N2220, N2209);
and AND2 (N2283, N2276, N1335);
or OR4 (N2284, N2254, N2261, N791, N555);
nand NAND4 (N2285, N2270, N1178, N1008, N581);
or OR4 (N2286, N2269, N734, N1129, N109);
not NOT1 (N2287, N2283);
nor NOR4 (N2288, N2279, N250, N439, N636);
buf BUF1 (N2289, N2273);
nor NOR2 (N2290, N2286, N1249);
or OR2 (N2291, N2287, N910);
and AND2 (N2292, N2285, N89);
buf BUF1 (N2293, N2289);
xor XOR2 (N2294, N2284, N2235);
nor NOR2 (N2295, N2274, N14);
and AND4 (N2296, N2288, N438, N636, N1310);
or OR4 (N2297, N2292, N980, N470, N1029);
buf BUF1 (N2298, N2297);
or OR2 (N2299, N2296, N11);
not NOT1 (N2300, N2272);
buf BUF1 (N2301, N2281);
not NOT1 (N2302, N2298);
nand NAND4 (N2303, N2290, N2012, N795, N150);
xor XOR2 (N2304, N2294, N2096);
buf BUF1 (N2305, N2302);
or OR3 (N2306, N2300, N1286, N1557);
buf BUF1 (N2307, N2291);
nor NOR3 (N2308, N2282, N1828, N1188);
or OR2 (N2309, N2295, N2196);
not NOT1 (N2310, N2306);
xor XOR2 (N2311, N2309, N1458);
or OR2 (N2312, N2299, N1240);
buf BUF1 (N2313, N2304);
nor NOR4 (N2314, N2301, N345, N744, N1719);
xor XOR2 (N2315, N2303, N908);
and AND4 (N2316, N2293, N1872, N39, N1729);
nor NOR4 (N2317, N2312, N866, N2287, N2224);
and AND3 (N2318, N2305, N962, N302);
buf BUF1 (N2319, N2317);
buf BUF1 (N2320, N2315);
nor NOR4 (N2321, N2311, N1686, N1957, N1182);
or OR2 (N2322, N2319, N1030);
not NOT1 (N2323, N2308);
buf BUF1 (N2324, N2322);
or OR2 (N2325, N2318, N364);
buf BUF1 (N2326, N2313);
or OR4 (N2327, N2321, N556, N1220, N1706);
nand NAND2 (N2328, N2310, N796);
or OR4 (N2329, N2316, N975, N2254, N2291);
not NOT1 (N2330, N2323);
nand NAND3 (N2331, N2326, N262, N1453);
and AND3 (N2332, N2330, N1784, N1275);
xor XOR2 (N2333, N2320, N1045);
xor XOR2 (N2334, N2314, N2228);
nand NAND4 (N2335, N2325, N1885, N316, N298);
buf BUF1 (N2336, N2333);
xor XOR2 (N2337, N2332, N278);
nor NOR2 (N2338, N2307, N539);
not NOT1 (N2339, N2331);
xor XOR2 (N2340, N2327, N117);
nand NAND2 (N2341, N2337, N1668);
xor XOR2 (N2342, N2339, N392);
nand NAND2 (N2343, N2342, N375);
xor XOR2 (N2344, N2341, N255);
and AND2 (N2345, N2329, N186);
or OR4 (N2346, N2345, N597, N2288, N1368);
and AND2 (N2347, N2334, N156);
buf BUF1 (N2348, N2346);
xor XOR2 (N2349, N2344, N977);
nor NOR3 (N2350, N2328, N447, N1257);
xor XOR2 (N2351, N2349, N1817);
or OR3 (N2352, N2340, N2246, N1608);
nor NOR4 (N2353, N2352, N1944, N642, N1040);
not NOT1 (N2354, N2338);
or OR2 (N2355, N2324, N749);
or OR2 (N2356, N2355, N535);
buf BUF1 (N2357, N2350);
nand NAND2 (N2358, N2343, N1821);
xor XOR2 (N2359, N2358, N693);
not NOT1 (N2360, N2348);
not NOT1 (N2361, N2354);
and AND2 (N2362, N2353, N1324);
buf BUF1 (N2363, N2356);
not NOT1 (N2364, N2335);
and AND3 (N2365, N2364, N2094, N1820);
not NOT1 (N2366, N2362);
nor NOR2 (N2367, N2351, N1572);
nor NOR2 (N2368, N2357, N171);
and AND4 (N2369, N2365, N1765, N961, N938);
nor NOR4 (N2370, N2336, N230, N246, N40);
or OR3 (N2371, N2359, N1690, N894);
xor XOR2 (N2372, N2366, N987);
buf BUF1 (N2373, N2372);
buf BUF1 (N2374, N2370);
xor XOR2 (N2375, N2361, N794);
and AND2 (N2376, N2374, N1575);
xor XOR2 (N2377, N2376, N621);
or OR2 (N2378, N2377, N1714);
xor XOR2 (N2379, N2378, N225);
and AND4 (N2380, N2368, N667, N368, N1051);
or OR4 (N2381, N2347, N1340, N1361, N405);
buf BUF1 (N2382, N2360);
nand NAND4 (N2383, N2381, N662, N41, N729);
and AND3 (N2384, N2382, N1600, N1772);
buf BUF1 (N2385, N2369);
nand NAND3 (N2386, N2367, N723, N805);
not NOT1 (N2387, N2379);
or OR3 (N2388, N2384, N196, N837);
nor NOR2 (N2389, N2371, N1185);
buf BUF1 (N2390, N2375);
or OR3 (N2391, N2363, N2181, N1505);
buf BUF1 (N2392, N2388);
or OR3 (N2393, N2391, N28, N1290);
nand NAND2 (N2394, N2380, N1536);
nand NAND2 (N2395, N2394, N867);
xor XOR2 (N2396, N2383, N1597);
not NOT1 (N2397, N2395);
buf BUF1 (N2398, N2385);
nor NOR4 (N2399, N2373, N511, N2255, N1699);
or OR3 (N2400, N2387, N2242, N1360);
nor NOR3 (N2401, N2400, N1380, N569);
xor XOR2 (N2402, N2396, N1978);
and AND4 (N2403, N2392, N789, N432, N2226);
and AND4 (N2404, N2402, N313, N686, N1319);
and AND4 (N2405, N2401, N1882, N1637, N143);
not NOT1 (N2406, N2390);
nor NOR2 (N2407, N2405, N1057);
not NOT1 (N2408, N2397);
nand NAND2 (N2409, N2386, N1001);
xor XOR2 (N2410, N2407, N229);
buf BUF1 (N2411, N2408);
buf BUF1 (N2412, N2389);
or OR3 (N2413, N2404, N947, N1321);
xor XOR2 (N2414, N2393, N1134);
nor NOR4 (N2415, N2403, N927, N126, N105);
buf BUF1 (N2416, N2414);
xor XOR2 (N2417, N2406, N8);
not NOT1 (N2418, N2398);
nand NAND2 (N2419, N2415, N848);
nand NAND3 (N2420, N2399, N882, N1540);
xor XOR2 (N2421, N2419, N2143);
or OR2 (N2422, N2410, N84);
buf BUF1 (N2423, N2420);
and AND3 (N2424, N2411, N1634, N852);
and AND2 (N2425, N2422, N623);
or OR2 (N2426, N2413, N725);
and AND4 (N2427, N2425, N384, N2035, N1166);
not NOT1 (N2428, N2416);
and AND2 (N2429, N2428, N861);
nand NAND4 (N2430, N2426, N2248, N1679, N1685);
and AND2 (N2431, N2429, N2354);
buf BUF1 (N2432, N2421);
not NOT1 (N2433, N2424);
and AND4 (N2434, N2409, N478, N1531, N617);
not NOT1 (N2435, N2431);
or OR3 (N2436, N2435, N1631, N1882);
nor NOR4 (N2437, N2427, N2061, N1150, N1708);
buf BUF1 (N2438, N2423);
and AND3 (N2439, N2437, N2319, N121);
nand NAND4 (N2440, N2412, N351, N2106, N1187);
nor NOR2 (N2441, N2418, N97);
and AND4 (N2442, N2432, N92, N767, N1398);
nor NOR2 (N2443, N2440, N1387);
or OR3 (N2444, N2443, N1646, N1160);
nor NOR3 (N2445, N2434, N1033, N2018);
buf BUF1 (N2446, N2444);
buf BUF1 (N2447, N2433);
or OR4 (N2448, N2436, N555, N1855, N1182);
or OR2 (N2449, N2442, N1290);
buf BUF1 (N2450, N2430);
buf BUF1 (N2451, N2449);
buf BUF1 (N2452, N2417);
not NOT1 (N2453, N2450);
nand NAND2 (N2454, N2447, N88);
nor NOR3 (N2455, N2441, N1006, N1556);
nor NOR2 (N2456, N2452, N205);
nor NOR3 (N2457, N2453, N969, N1061);
not NOT1 (N2458, N2446);
xor XOR2 (N2459, N2458, N1866);
and AND4 (N2460, N2448, N2199, N939, N1717);
nor NOR3 (N2461, N2438, N583, N1953);
not NOT1 (N2462, N2451);
and AND3 (N2463, N2461, N510, N326);
and AND3 (N2464, N2439, N2199, N2071);
nor NOR3 (N2465, N2460, N213, N1257);
xor XOR2 (N2466, N2463, N1176);
buf BUF1 (N2467, N2464);
xor XOR2 (N2468, N2462, N686);
nand NAND3 (N2469, N2468, N255, N2070);
buf BUF1 (N2470, N2465);
not NOT1 (N2471, N2467);
or OR2 (N2472, N2466, N1760);
nand NAND2 (N2473, N2471, N1537);
nor NOR2 (N2474, N2457, N519);
nand NAND4 (N2475, N2472, N1982, N128, N831);
buf BUF1 (N2476, N2456);
nor NOR2 (N2477, N2455, N1279);
or OR4 (N2478, N2445, N2022, N890, N2000);
xor XOR2 (N2479, N2473, N712);
and AND3 (N2480, N2454, N1280, N1422);
buf BUF1 (N2481, N2459);
xor XOR2 (N2482, N2477, N2161);
nand NAND3 (N2483, N2476, N1262, N211);
not NOT1 (N2484, N2481);
or OR2 (N2485, N2484, N1412);
nand NAND2 (N2486, N2478, N2231);
xor XOR2 (N2487, N2482, N2274);
xor XOR2 (N2488, N2475, N2375);
and AND2 (N2489, N2479, N1099);
buf BUF1 (N2490, N2489);
not NOT1 (N2491, N2480);
not NOT1 (N2492, N2474);
nor NOR4 (N2493, N2483, N376, N1470, N1483);
not NOT1 (N2494, N2492);
and AND4 (N2495, N2493, N1077, N2288, N877);
not NOT1 (N2496, N2488);
not NOT1 (N2497, N2490);
nand NAND4 (N2498, N2469, N832, N422, N1637);
xor XOR2 (N2499, N2491, N13);
not NOT1 (N2500, N2494);
nor NOR4 (N2501, N2496, N1518, N367, N1338);
buf BUF1 (N2502, N2485);
not NOT1 (N2503, N2495);
xor XOR2 (N2504, N2503, N1114);
or OR3 (N2505, N2487, N615, N81);
and AND3 (N2506, N2504, N2043, N2434);
not NOT1 (N2507, N2498);
and AND3 (N2508, N2502, N2245, N878);
buf BUF1 (N2509, N2499);
buf BUF1 (N2510, N2506);
nor NOR3 (N2511, N2500, N2349, N474);
and AND4 (N2512, N2511, N1525, N336, N1315);
nor NOR4 (N2513, N2470, N755, N1738, N78);
not NOT1 (N2514, N2505);
xor XOR2 (N2515, N2514, N2337);
nand NAND2 (N2516, N2512, N2338);
nand NAND2 (N2517, N2509, N1435);
not NOT1 (N2518, N2508);
and AND3 (N2519, N2516, N510, N1806);
and AND2 (N2520, N2507, N828);
nor NOR4 (N2521, N2501, N2286, N1124, N2159);
nand NAND3 (N2522, N2486, N2351, N930);
nand NAND2 (N2523, N2521, N1599);
or OR4 (N2524, N2517, N1373, N1402, N1067);
not NOT1 (N2525, N2497);
or OR2 (N2526, N2525, N1649);
not NOT1 (N2527, N2520);
buf BUF1 (N2528, N2515);
not NOT1 (N2529, N2526);
not NOT1 (N2530, N2510);
or OR4 (N2531, N2519, N1660, N1812, N150);
nor NOR2 (N2532, N2513, N1535);
buf BUF1 (N2533, N2527);
buf BUF1 (N2534, N2533);
nor NOR3 (N2535, N2530, N1800, N1996);
buf BUF1 (N2536, N2524);
not NOT1 (N2537, N2536);
not NOT1 (N2538, N2523);
or OR4 (N2539, N2528, N2243, N2032, N1522);
buf BUF1 (N2540, N2531);
not NOT1 (N2541, N2529);
nand NAND2 (N2542, N2538, N994);
nor NOR4 (N2543, N2534, N1682, N555, N1227);
nand NAND2 (N2544, N2522, N1043);
not NOT1 (N2545, N2539);
xor XOR2 (N2546, N2543, N1633);
xor XOR2 (N2547, N2537, N836);
and AND4 (N2548, N2535, N307, N92, N2230);
buf BUF1 (N2549, N2548);
and AND3 (N2550, N2545, N1452, N49);
nor NOR4 (N2551, N2532, N147, N1637, N1107);
xor XOR2 (N2552, N2549, N902);
or OR4 (N2553, N2552, N1778, N1156, N1632);
nor NOR3 (N2554, N2540, N1736, N2322);
buf BUF1 (N2555, N2544);
or OR2 (N2556, N2555, N1000);
not NOT1 (N2557, N2518);
and AND4 (N2558, N2553, N1331, N1452, N627);
nor NOR2 (N2559, N2550, N2229);
nand NAND3 (N2560, N2557, N986, N2465);
and AND3 (N2561, N2560, N843, N1975);
nor NOR2 (N2562, N2558, N1561);
xor XOR2 (N2563, N2541, N2076);
and AND2 (N2564, N2562, N278);
xor XOR2 (N2565, N2563, N714);
nor NOR2 (N2566, N2547, N2355);
nor NOR4 (N2567, N2566, N1541, N603, N2466);
xor XOR2 (N2568, N2561, N1740);
nand NAND2 (N2569, N2564, N842);
not NOT1 (N2570, N2565);
or OR2 (N2571, N2551, N1244);
nand NAND3 (N2572, N2569, N1143, N599);
nor NOR4 (N2573, N2559, N65, N13, N957);
xor XOR2 (N2574, N2542, N116);
nand NAND2 (N2575, N2572, N1734);
not NOT1 (N2576, N2570);
or OR2 (N2577, N2554, N741);
or OR2 (N2578, N2571, N2047);
nor NOR4 (N2579, N2575, N1666, N1002, N776);
xor XOR2 (N2580, N2567, N1499);
buf BUF1 (N2581, N2546);
or OR4 (N2582, N2574, N327, N2180, N834);
xor XOR2 (N2583, N2581, N226);
and AND4 (N2584, N2579, N1974, N350, N449);
nor NOR4 (N2585, N2580, N2218, N1646, N76);
xor XOR2 (N2586, N2573, N2488);
xor XOR2 (N2587, N2577, N16);
or OR2 (N2588, N2587, N2400);
buf BUF1 (N2589, N2585);
xor XOR2 (N2590, N2582, N440);
xor XOR2 (N2591, N2588, N797);
and AND4 (N2592, N2556, N779, N485, N1601);
xor XOR2 (N2593, N2586, N337);
and AND3 (N2594, N2590, N356, N972);
not NOT1 (N2595, N2591);
not NOT1 (N2596, N2568);
xor XOR2 (N2597, N2578, N2122);
or OR3 (N2598, N2593, N2443, N972);
and AND4 (N2599, N2589, N1605, N1573, N727);
and AND2 (N2600, N2592, N2212);
not NOT1 (N2601, N2598);
and AND4 (N2602, N2601, N2292, N142, N2154);
xor XOR2 (N2603, N2584, N1475);
nand NAND3 (N2604, N2594, N1806, N466);
xor XOR2 (N2605, N2602, N428);
nor NOR3 (N2606, N2597, N1014, N1206);
nand NAND2 (N2607, N2583, N2270);
buf BUF1 (N2608, N2605);
not NOT1 (N2609, N2595);
nor NOR3 (N2610, N2603, N1239, N1377);
nand NAND3 (N2611, N2599, N1074, N882);
not NOT1 (N2612, N2609);
buf BUF1 (N2613, N2610);
and AND4 (N2614, N2606, N2092, N2152, N1123);
nor NOR4 (N2615, N2576, N2090, N1833, N1368);
and AND3 (N2616, N2613, N1266, N1781);
or OR4 (N2617, N2611, N1060, N267, N216);
or OR4 (N2618, N2607, N865, N1081, N2415);
xor XOR2 (N2619, N2612, N1498);
and AND4 (N2620, N2615, N1346, N1469, N116);
and AND4 (N2621, N2600, N1130, N52, N643);
buf BUF1 (N2622, N2608);
and AND3 (N2623, N2619, N1620, N1464);
not NOT1 (N2624, N2604);
or OR3 (N2625, N2621, N2077, N2175);
nor NOR2 (N2626, N2614, N1653);
or OR2 (N2627, N2616, N1187);
nor NOR4 (N2628, N2623, N1974, N1416, N1607);
nand NAND3 (N2629, N2620, N266, N1736);
and AND2 (N2630, N2617, N1639);
nand NAND2 (N2631, N2627, N589);
nor NOR2 (N2632, N2628, N944);
and AND4 (N2633, N2624, N2163, N2030, N687);
nand NAND2 (N2634, N2622, N1481);
not NOT1 (N2635, N2596);
and AND2 (N2636, N2629, N1134);
buf BUF1 (N2637, N2630);
and AND4 (N2638, N2626, N1265, N662, N726);
and AND2 (N2639, N2634, N2168);
or OR2 (N2640, N2637, N2627);
nand NAND4 (N2641, N2638, N2546, N2318, N1622);
or OR4 (N2642, N2636, N1855, N862, N329);
xor XOR2 (N2643, N2639, N1019);
or OR4 (N2644, N2633, N863, N1920, N498);
nor NOR2 (N2645, N2644, N1664);
or OR2 (N2646, N2635, N2382);
nand NAND3 (N2647, N2618, N1664, N2501);
xor XOR2 (N2648, N2642, N1731);
and AND4 (N2649, N2631, N345, N871, N1354);
not NOT1 (N2650, N2643);
not NOT1 (N2651, N2640);
xor XOR2 (N2652, N2646, N1754);
nand NAND4 (N2653, N2625, N769, N1249, N702);
xor XOR2 (N2654, N2647, N526);
not NOT1 (N2655, N2654);
nor NOR2 (N2656, N2641, N1347);
or OR4 (N2657, N2645, N129, N1314, N1198);
xor XOR2 (N2658, N2657, N1120);
buf BUF1 (N2659, N2655);
buf BUF1 (N2660, N2658);
nand NAND4 (N2661, N2649, N1759, N2456, N2623);
nor NOR4 (N2662, N2661, N886, N1522, N2225);
not NOT1 (N2663, N2650);
not NOT1 (N2664, N2652);
nand NAND3 (N2665, N2648, N50, N2273);
buf BUF1 (N2666, N2651);
nor NOR4 (N2667, N2663, N513, N1010, N648);
not NOT1 (N2668, N2667);
not NOT1 (N2669, N2662);
buf BUF1 (N2670, N2660);
not NOT1 (N2671, N2670);
or OR4 (N2672, N2664, N778, N1509, N331);
or OR4 (N2673, N2665, N1602, N1460, N1494);
and AND2 (N2674, N2659, N1747);
xor XOR2 (N2675, N2666, N2481);
and AND2 (N2676, N2675, N32);
nand NAND3 (N2677, N2669, N1523, N2598);
buf BUF1 (N2678, N2676);
not NOT1 (N2679, N2673);
nor NOR3 (N2680, N2656, N870, N1405);
buf BUF1 (N2681, N2632);
and AND3 (N2682, N2677, N1345, N2670);
and AND3 (N2683, N2674, N891, N334);
or OR3 (N2684, N2668, N689, N1453);
nand NAND2 (N2685, N2653, N1963);
xor XOR2 (N2686, N2678, N1593);
nand NAND4 (N2687, N2683, N2076, N1632, N575);
or OR3 (N2688, N2672, N378, N2284);
nand NAND4 (N2689, N2685, N1718, N14, N786);
xor XOR2 (N2690, N2686, N2188);
buf BUF1 (N2691, N2682);
or OR2 (N2692, N2671, N2652);
not NOT1 (N2693, N2692);
and AND4 (N2694, N2693, N2193, N433, N407);
and AND4 (N2695, N2689, N1279, N1315, N1542);
nand NAND4 (N2696, N2684, N2, N1127, N634);
nor NOR4 (N2697, N2696, N1949, N168, N2491);
nand NAND4 (N2698, N2690, N2194, N1495, N1548);
and AND3 (N2699, N2695, N7, N1595);
and AND3 (N2700, N2698, N1040, N2229);
nand NAND2 (N2701, N2680, N932);
not NOT1 (N2702, N2699);
or OR2 (N2703, N2691, N1194);
not NOT1 (N2704, N2697);
or OR2 (N2705, N2703, N92);
not NOT1 (N2706, N2681);
nand NAND4 (N2707, N2687, N445, N1603, N1471);
not NOT1 (N2708, N2688);
nand NAND2 (N2709, N2700, N1654);
not NOT1 (N2710, N2706);
or OR4 (N2711, N2709, N605, N2559, N1290);
buf BUF1 (N2712, N2707);
or OR2 (N2713, N2694, N1996);
and AND2 (N2714, N2704, N1348);
nand NAND4 (N2715, N2712, N1649, N2196, N1013);
nor NOR2 (N2716, N2708, N129);
and AND2 (N2717, N2679, N2484);
not NOT1 (N2718, N2717);
or OR3 (N2719, N2705, N1583, N927);
nand NAND3 (N2720, N2713, N2127, N2270);
nand NAND2 (N2721, N2711, N998);
buf BUF1 (N2722, N2718);
not NOT1 (N2723, N2701);
and AND2 (N2724, N2721, N2185);
and AND4 (N2725, N2702, N1063, N2428, N741);
or OR2 (N2726, N2720, N1830);
nand NAND2 (N2727, N2724, N10);
and AND3 (N2728, N2714, N2029, N1813);
buf BUF1 (N2729, N2728);
nand NAND2 (N2730, N2729, N883);
not NOT1 (N2731, N2716);
or OR2 (N2732, N2715, N676);
nor NOR3 (N2733, N2710, N1806, N2356);
xor XOR2 (N2734, N2725, N899);
xor XOR2 (N2735, N2734, N2125);
xor XOR2 (N2736, N2727, N2529);
and AND2 (N2737, N2733, N2001);
and AND4 (N2738, N2736, N1344, N2546, N1253);
nand NAND2 (N2739, N2737, N1062);
or OR2 (N2740, N2722, N2607);
and AND4 (N2741, N2726, N2619, N1387, N1300);
buf BUF1 (N2742, N2730);
nor NOR2 (N2743, N2735, N1797);
xor XOR2 (N2744, N2740, N1001);
and AND3 (N2745, N2731, N2072, N1013);
nand NAND3 (N2746, N2742, N2494, N1519);
nor NOR3 (N2747, N2744, N2123, N642);
or OR2 (N2748, N2746, N390);
nand NAND2 (N2749, N2738, N1127);
or OR2 (N2750, N2749, N2181);
not NOT1 (N2751, N2732);
or OR4 (N2752, N2743, N2288, N2687, N2463);
not NOT1 (N2753, N2748);
or OR2 (N2754, N2751, N1200);
and AND2 (N2755, N2752, N1414);
nand NAND3 (N2756, N2741, N2145, N1813);
and AND4 (N2757, N2756, N2485, N1571, N718);
and AND3 (N2758, N2757, N2462, N1101);
not NOT1 (N2759, N2754);
and AND2 (N2760, N2739, N739);
not NOT1 (N2761, N2745);
nor NOR4 (N2762, N2758, N1925, N457, N1339);
or OR2 (N2763, N2760, N2541);
nor NOR2 (N2764, N2719, N370);
nand NAND3 (N2765, N2753, N2035, N1477);
buf BUF1 (N2766, N2723);
nor NOR3 (N2767, N2750, N1687, N2145);
buf BUF1 (N2768, N2747);
or OR4 (N2769, N2761, N899, N1784, N88);
xor XOR2 (N2770, N2764, N328);
xor XOR2 (N2771, N2769, N671);
and AND4 (N2772, N2771, N1668, N1333, N173);
not NOT1 (N2773, N2770);
buf BUF1 (N2774, N2773);
nand NAND3 (N2775, N2767, N1529, N91);
or OR2 (N2776, N2763, N2380);
buf BUF1 (N2777, N2776);
buf BUF1 (N2778, N2775);
or OR2 (N2779, N2755, N2702);
nor NOR4 (N2780, N2766, N162, N2664, N668);
xor XOR2 (N2781, N2777, N492);
and AND3 (N2782, N2765, N1287, N134);
and AND3 (N2783, N2778, N69, N212);
or OR3 (N2784, N2780, N1371, N144);
and AND3 (N2785, N2782, N2530, N1894);
xor XOR2 (N2786, N2785, N89);
or OR2 (N2787, N2781, N1595);
not NOT1 (N2788, N2779);
not NOT1 (N2789, N2762);
and AND2 (N2790, N2787, N445);
nand NAND2 (N2791, N2784, N1408);
and AND4 (N2792, N2789, N1841, N795, N1440);
not NOT1 (N2793, N2791);
buf BUF1 (N2794, N2759);
and AND2 (N2795, N2774, N2598);
not NOT1 (N2796, N2783);
buf BUF1 (N2797, N2795);
xor XOR2 (N2798, N2793, N1227);
buf BUF1 (N2799, N2797);
or OR4 (N2800, N2799, N1369, N1434, N2257);
buf BUF1 (N2801, N2796);
or OR4 (N2802, N2790, N1584, N973, N1202);
nor NOR2 (N2803, N2786, N1334);
buf BUF1 (N2804, N2798);
not NOT1 (N2805, N2794);
buf BUF1 (N2806, N2768);
or OR3 (N2807, N2802, N1746, N225);
buf BUF1 (N2808, N2805);
nand NAND2 (N2809, N2807, N1624);
buf BUF1 (N2810, N2803);
nor NOR4 (N2811, N2810, N370, N736, N1451);
or OR3 (N2812, N2811, N1672, N359);
buf BUF1 (N2813, N2804);
nor NOR2 (N2814, N2808, N1694);
nand NAND3 (N2815, N2800, N2130, N1590);
nand NAND2 (N2816, N2812, N567);
not NOT1 (N2817, N2815);
nand NAND2 (N2818, N2792, N2595);
or OR3 (N2819, N2817, N1292, N1299);
nor NOR3 (N2820, N2801, N2170, N980);
nand NAND4 (N2821, N2820, N2791, N1580, N632);
nor NOR3 (N2822, N2821, N585, N159);
nor NOR3 (N2823, N2822, N2627, N504);
buf BUF1 (N2824, N2772);
or OR2 (N2825, N2814, N902);
nand NAND3 (N2826, N2818, N1688, N2422);
nand NAND3 (N2827, N2806, N2027, N2320);
buf BUF1 (N2828, N2816);
buf BUF1 (N2829, N2819);
not NOT1 (N2830, N2813);
not NOT1 (N2831, N2824);
not NOT1 (N2832, N2823);
not NOT1 (N2833, N2830);
buf BUF1 (N2834, N2833);
or OR3 (N2835, N2829, N213, N643);
xor XOR2 (N2836, N2835, N276);
nor NOR3 (N2837, N2836, N748, N1118);
not NOT1 (N2838, N2809);
not NOT1 (N2839, N2826);
xor XOR2 (N2840, N2828, N2425);
xor XOR2 (N2841, N2788, N2246);
and AND3 (N2842, N2841, N71, N2538);
or OR4 (N2843, N2827, N352, N1770, N1386);
and AND3 (N2844, N2825, N1662, N1095);
nand NAND4 (N2845, N2837, N606, N1661, N1295);
nor NOR2 (N2846, N2831, N1258);
buf BUF1 (N2847, N2846);
xor XOR2 (N2848, N2832, N1361);
and AND2 (N2849, N2840, N226);
or OR2 (N2850, N2844, N754);
not NOT1 (N2851, N2839);
not NOT1 (N2852, N2834);
buf BUF1 (N2853, N2848);
nor NOR4 (N2854, N2847, N929, N2717, N210);
xor XOR2 (N2855, N2853, N956);
buf BUF1 (N2856, N2850);
and AND2 (N2857, N2854, N2341);
and AND3 (N2858, N2849, N1321, N2408);
or OR2 (N2859, N2842, N1899);
nor NOR4 (N2860, N2856, N1274, N2169, N331);
buf BUF1 (N2861, N2857);
buf BUF1 (N2862, N2855);
nand NAND2 (N2863, N2843, N1679);
not NOT1 (N2864, N2851);
and AND2 (N2865, N2860, N801);
xor XOR2 (N2866, N2858, N2165);
nor NOR3 (N2867, N2861, N717, N942);
or OR2 (N2868, N2859, N946);
or OR3 (N2869, N2868, N2542, N2053);
or OR4 (N2870, N2838, N341, N1936, N1286);
xor XOR2 (N2871, N2867, N233);
or OR2 (N2872, N2870, N1047);
nand NAND2 (N2873, N2852, N2212);
buf BUF1 (N2874, N2869);
and AND3 (N2875, N2872, N2810, N484);
buf BUF1 (N2876, N2875);
and AND2 (N2877, N2863, N674);
xor XOR2 (N2878, N2874, N1870);
buf BUF1 (N2879, N2876);
or OR4 (N2880, N2877, N779, N1462, N1528);
and AND3 (N2881, N2864, N1557, N2599);
nand NAND4 (N2882, N2880, N2685, N1073, N2174);
buf BUF1 (N2883, N2879);
and AND2 (N2884, N2883, N1881);
and AND4 (N2885, N2882, N2416, N597, N2378);
xor XOR2 (N2886, N2873, N1370);
not NOT1 (N2887, N2884);
nor NOR4 (N2888, N2878, N1022, N1529, N805);
or OR2 (N2889, N2888, N896);
buf BUF1 (N2890, N2886);
nand NAND3 (N2891, N2865, N2513, N1091);
not NOT1 (N2892, N2881);
buf BUF1 (N2893, N2891);
xor XOR2 (N2894, N2845, N1176);
buf BUF1 (N2895, N2890);
buf BUF1 (N2896, N2894);
nor NOR3 (N2897, N2887, N2355, N1721);
nand NAND2 (N2898, N2895, N73);
or OR3 (N2899, N2893, N1609, N1465);
buf BUF1 (N2900, N2899);
or OR4 (N2901, N2889, N1958, N1668, N517);
nand NAND2 (N2902, N2897, N1002);
or OR4 (N2903, N2902, N2678, N1940, N2489);
nor NOR2 (N2904, N2862, N1345);
not NOT1 (N2905, N2896);
xor XOR2 (N2906, N2904, N2656);
nand NAND3 (N2907, N2898, N2264, N244);
nor NOR4 (N2908, N2866, N2245, N2691, N1631);
and AND3 (N2909, N2903, N2074, N214);
xor XOR2 (N2910, N2905, N566);
xor XOR2 (N2911, N2892, N2302);
nor NOR3 (N2912, N2900, N2289, N605);
and AND3 (N2913, N2906, N382, N1092);
xor XOR2 (N2914, N2885, N1662);
or OR3 (N2915, N2908, N1515, N153);
nor NOR2 (N2916, N2915, N1248);
and AND4 (N2917, N2871, N755, N161, N2320);
not NOT1 (N2918, N2913);
nor NOR4 (N2919, N2911, N2022, N622, N1748);
xor XOR2 (N2920, N2914, N2841);
nor NOR4 (N2921, N2907, N1813, N126, N1080);
nand NAND4 (N2922, N2920, N2283, N1548, N1632);
and AND3 (N2923, N2919, N2599, N1786);
buf BUF1 (N2924, N2922);
and AND4 (N2925, N2918, N484, N560, N2188);
or OR4 (N2926, N2923, N765, N2031, N301);
or OR4 (N2927, N2910, N2720, N2444, N429);
or OR3 (N2928, N2921, N1489, N2743);
not NOT1 (N2929, N2924);
nand NAND3 (N2930, N2909, N1029, N440);
buf BUF1 (N2931, N2901);
nand NAND2 (N2932, N2912, N1853);
buf BUF1 (N2933, N2931);
buf BUF1 (N2934, N2926);
xor XOR2 (N2935, N2930, N2288);
nor NOR4 (N2936, N2935, N45, N1902, N566);
not NOT1 (N2937, N2917);
nor NOR3 (N2938, N2929, N1024, N672);
and AND4 (N2939, N2932, N1756, N2109, N168);
or OR3 (N2940, N2916, N2042, N1423);
or OR4 (N2941, N2928, N2929, N1007, N1536);
not NOT1 (N2942, N2936);
and AND3 (N2943, N2927, N1491, N1048);
or OR3 (N2944, N2941, N1685, N2344);
and AND3 (N2945, N2938, N1108, N841);
xor XOR2 (N2946, N2934, N2811);
not NOT1 (N2947, N2933);
nor NOR2 (N2948, N2925, N2798);
nand NAND3 (N2949, N2940, N1086, N770);
nand NAND4 (N2950, N2944, N507, N1943, N2388);
xor XOR2 (N2951, N2947, N2451);
nor NOR3 (N2952, N2943, N2107, N1766);
nor NOR2 (N2953, N2937, N2262);
not NOT1 (N2954, N2951);
and AND2 (N2955, N2942, N1599);
nor NOR3 (N2956, N2949, N2738, N1858);
nand NAND2 (N2957, N2956, N2053);
nand NAND3 (N2958, N2945, N890, N1830);
nor NOR4 (N2959, N2950, N1518, N528, N1888);
not NOT1 (N2960, N2946);
buf BUF1 (N2961, N2955);
nor NOR2 (N2962, N2959, N1047);
or OR2 (N2963, N2954, N2496);
or OR2 (N2964, N2958, N983);
or OR2 (N2965, N2961, N1310);
or OR3 (N2966, N2953, N2708, N778);
and AND3 (N2967, N2939, N1734, N2350);
or OR2 (N2968, N2963, N1410);
or OR2 (N2969, N2948, N974);
and AND4 (N2970, N2969, N2768, N702, N328);
or OR4 (N2971, N2968, N1666, N1342, N2540);
or OR2 (N2972, N2960, N1346);
xor XOR2 (N2973, N2965, N526);
buf BUF1 (N2974, N2962);
and AND2 (N2975, N2967, N277);
not NOT1 (N2976, N2957);
xor XOR2 (N2977, N2973, N1132);
or OR4 (N2978, N2966, N2168, N2354, N2366);
buf BUF1 (N2979, N2964);
xor XOR2 (N2980, N2972, N372);
not NOT1 (N2981, N2980);
or OR4 (N2982, N2981, N143, N2596, N1952);
nor NOR4 (N2983, N2975, N1263, N2529, N2579);
or OR2 (N2984, N2971, N1583);
not NOT1 (N2985, N2982);
xor XOR2 (N2986, N2974, N683);
not NOT1 (N2987, N2970);
xor XOR2 (N2988, N2983, N2628);
nor NOR3 (N2989, N2987, N2928, N2412);
xor XOR2 (N2990, N2988, N1843);
nand NAND3 (N2991, N2985, N208, N2110);
and AND4 (N2992, N2991, N2090, N685, N945);
and AND4 (N2993, N2976, N2704, N2750, N631);
and AND4 (N2994, N2990, N1181, N1604, N896);
xor XOR2 (N2995, N2993, N2243);
and AND4 (N2996, N2984, N1127, N838, N2537);
xor XOR2 (N2997, N2979, N570);
or OR4 (N2998, N2997, N1294, N1124, N1668);
nand NAND2 (N2999, N2989, N429);
buf BUF1 (N3000, N2986);
xor XOR2 (N3001, N2995, N2591);
buf BUF1 (N3002, N2978);
or OR4 (N3003, N3002, N774, N1273, N974);
and AND2 (N3004, N3003, N2780);
buf BUF1 (N3005, N2992);
xor XOR2 (N3006, N2952, N1484);
xor XOR2 (N3007, N2977, N396);
nand NAND4 (N3008, N3004, N2706, N1726, N2739);
xor XOR2 (N3009, N3000, N1854);
or OR3 (N3010, N3008, N1708, N13);
buf BUF1 (N3011, N3005);
and AND4 (N3012, N2994, N1171, N402, N2236);
nor NOR4 (N3013, N2998, N1911, N186, N318);
and AND4 (N3014, N3011, N2376, N778, N238);
not NOT1 (N3015, N3012);
nor NOR4 (N3016, N2999, N1673, N1999, N2854);
or OR3 (N3017, N3001, N1471, N260);
nor NOR2 (N3018, N3010, N750);
buf BUF1 (N3019, N3017);
nor NOR2 (N3020, N3006, N2029);
nand NAND2 (N3021, N3018, N922);
buf BUF1 (N3022, N3019);
or OR3 (N3023, N3009, N2709, N454);
xor XOR2 (N3024, N3021, N1815);
or OR3 (N3025, N3016, N440, N1987);
xor XOR2 (N3026, N3024, N2147);
xor XOR2 (N3027, N3023, N1854);
nor NOR3 (N3028, N3022, N2103, N1027);
and AND3 (N3029, N3027, N1838, N2019);
not NOT1 (N3030, N3007);
nand NAND2 (N3031, N3025, N1626);
nand NAND2 (N3032, N3029, N1767);
xor XOR2 (N3033, N3014, N612);
not NOT1 (N3034, N3028);
xor XOR2 (N3035, N3015, N1556);
xor XOR2 (N3036, N3034, N1209);
nand NAND3 (N3037, N3033, N408, N1398);
nor NOR4 (N3038, N3026, N1453, N1600, N1450);
xor XOR2 (N3039, N3030, N1063);
or OR3 (N3040, N3013, N1352, N2176);
and AND4 (N3041, N3038, N933, N773, N346);
buf BUF1 (N3042, N3040);
buf BUF1 (N3043, N3020);
nor NOR4 (N3044, N3039, N138, N89, N2640);
nand NAND2 (N3045, N3031, N1514);
and AND2 (N3046, N3042, N1409);
nor NOR2 (N3047, N3032, N2431);
buf BUF1 (N3048, N3036);
nor NOR3 (N3049, N3045, N383, N1887);
not NOT1 (N3050, N3048);
not NOT1 (N3051, N3041);
nand NAND3 (N3052, N3049, N382, N1756);
or OR4 (N3053, N3047, N3050, N273, N1069);
nor NOR4 (N3054, N2405, N1990, N2610, N1788);
not NOT1 (N3055, N3044);
or OR3 (N3056, N3054, N700, N2082);
not NOT1 (N3057, N3052);
not NOT1 (N3058, N3046);
nand NAND3 (N3059, N3055, N163, N347);
or OR4 (N3060, N3053, N1171, N2383, N563);
xor XOR2 (N3061, N3058, N1083);
xor XOR2 (N3062, N3037, N613);
or OR3 (N3063, N2996, N785, N1954);
xor XOR2 (N3064, N3060, N2276);
xor XOR2 (N3065, N3051, N2232);
nand NAND2 (N3066, N3057, N405);
xor XOR2 (N3067, N3061, N729);
not NOT1 (N3068, N3067);
xor XOR2 (N3069, N3065, N129);
buf BUF1 (N3070, N3056);
buf BUF1 (N3071, N3068);
not NOT1 (N3072, N3071);
nor NOR4 (N3073, N3064, N107, N3069, N2130);
buf BUF1 (N3074, N1073);
nor NOR3 (N3075, N3063, N35, N969);
not NOT1 (N3076, N3059);
buf BUF1 (N3077, N3066);
nor NOR4 (N3078, N3076, N392, N2279, N2918);
xor XOR2 (N3079, N3072, N12);
or OR3 (N3080, N3074, N851, N1534);
and AND4 (N3081, N3035, N263, N186, N2633);
xor XOR2 (N3082, N3080, N2418);
or OR4 (N3083, N3082, N512, N1703, N1272);
or OR3 (N3084, N3062, N1213, N2240);
and AND2 (N3085, N3070, N1190);
buf BUF1 (N3086, N3073);
or OR3 (N3087, N3085, N1625, N1650);
buf BUF1 (N3088, N3084);
not NOT1 (N3089, N3088);
and AND3 (N3090, N3089, N1646, N2778);
nand NAND4 (N3091, N3081, N2729, N2818, N314);
nand NAND4 (N3092, N3091, N2668, N58, N2095);
or OR3 (N3093, N3090, N775, N1854);
nand NAND4 (N3094, N3092, N2614, N228, N631);
and AND2 (N3095, N3075, N2848);
nand NAND3 (N3096, N3093, N1038, N382);
buf BUF1 (N3097, N3077);
or OR4 (N3098, N3096, N3074, N2515, N2043);
buf BUF1 (N3099, N3078);
nor NOR2 (N3100, N3079, N2452);
buf BUF1 (N3101, N3043);
nor NOR4 (N3102, N3098, N1540, N875, N2293);
not NOT1 (N3103, N3100);
not NOT1 (N3104, N3083);
nand NAND2 (N3105, N3102, N2168);
xor XOR2 (N3106, N3087, N1296);
nand NAND4 (N3107, N3106, N1922, N1460, N3093);
and AND2 (N3108, N3095, N2210);
nor NOR3 (N3109, N3101, N2698, N1802);
nor NOR2 (N3110, N3104, N2799);
xor XOR2 (N3111, N3107, N766);
nand NAND3 (N3112, N3099, N665, N764);
nor NOR2 (N3113, N3110, N277);
nand NAND3 (N3114, N3103, N471, N1303);
buf BUF1 (N3115, N3114);
nand NAND3 (N3116, N3086, N237, N1210);
or OR4 (N3117, N3108, N2937, N3109, N2742);
not NOT1 (N3118, N897);
nor NOR4 (N3119, N3105, N1401, N873, N1758);
nand NAND4 (N3120, N3113, N867, N360, N433);
and AND2 (N3121, N3116, N1274);
and AND2 (N3122, N3119, N261);
buf BUF1 (N3123, N3122);
or OR2 (N3124, N3094, N1124);
not NOT1 (N3125, N3123);
nor NOR2 (N3126, N3097, N2451);
xor XOR2 (N3127, N3120, N836);
buf BUF1 (N3128, N3121);
buf BUF1 (N3129, N3118);
or OR2 (N3130, N3115, N689);
nor NOR4 (N3131, N3124, N1588, N3119, N1454);
buf BUF1 (N3132, N3126);
not NOT1 (N3133, N3112);
not NOT1 (N3134, N3133);
buf BUF1 (N3135, N3131);
or OR3 (N3136, N3129, N346, N1745);
buf BUF1 (N3137, N3132);
nand NAND2 (N3138, N3136, N986);
nand NAND2 (N3139, N3138, N144);
nand NAND3 (N3140, N3130, N350, N24);
or OR2 (N3141, N3139, N2176);
xor XOR2 (N3142, N3117, N1903);
xor XOR2 (N3143, N3128, N768);
and AND3 (N3144, N3142, N315, N1788);
xor XOR2 (N3145, N3140, N2162);
buf BUF1 (N3146, N3141);
nand NAND2 (N3147, N3134, N1441);
nor NOR2 (N3148, N3147, N2328);
not NOT1 (N3149, N3137);
buf BUF1 (N3150, N3144);
or OR2 (N3151, N3146, N909);
not NOT1 (N3152, N3149);
not NOT1 (N3153, N3150);
nand NAND4 (N3154, N3151, N2455, N2711, N544);
nand NAND2 (N3155, N3111, N1039);
nor NOR4 (N3156, N3125, N1178, N1923, N3144);
xor XOR2 (N3157, N3153, N2076);
not NOT1 (N3158, N3127);
buf BUF1 (N3159, N3158);
and AND2 (N3160, N3156, N678);
xor XOR2 (N3161, N3148, N971);
or OR4 (N3162, N3145, N440, N2199, N611);
or OR2 (N3163, N3154, N3021);
xor XOR2 (N3164, N3161, N2132);
and AND3 (N3165, N3159, N2669, N565);
nand NAND3 (N3166, N3162, N1194, N994);
nor NOR2 (N3167, N3135, N1566);
xor XOR2 (N3168, N3157, N2411);
or OR2 (N3169, N3152, N15);
xor XOR2 (N3170, N3163, N691);
or OR3 (N3171, N3165, N980, N91);
buf BUF1 (N3172, N3155);
or OR2 (N3173, N3167, N521);
xor XOR2 (N3174, N3171, N875);
buf BUF1 (N3175, N3173);
nand NAND2 (N3176, N3168, N2336);
buf BUF1 (N3177, N3170);
nor NOR2 (N3178, N3160, N82);
or OR3 (N3179, N3172, N2160, N2103);
nor NOR4 (N3180, N3179, N1388, N1859, N2527);
or OR2 (N3181, N3169, N1784);
not NOT1 (N3182, N3143);
or OR3 (N3183, N3174, N9, N760);
nand NAND2 (N3184, N3181, N541);
nand NAND3 (N3185, N3164, N602, N1014);
not NOT1 (N3186, N3180);
and AND4 (N3187, N3166, N22, N165, N2235);
and AND4 (N3188, N3175, N1892, N2619, N1780);
xor XOR2 (N3189, N3184, N1086);
not NOT1 (N3190, N3185);
nand NAND2 (N3191, N3186, N1170);
or OR3 (N3192, N3191, N1329, N487);
not NOT1 (N3193, N3188);
nor NOR4 (N3194, N3183, N2899, N1142, N482);
buf BUF1 (N3195, N3178);
or OR2 (N3196, N3177, N1559);
xor XOR2 (N3197, N3189, N1527);
or OR2 (N3198, N3192, N1665);
buf BUF1 (N3199, N3197);
nor NOR4 (N3200, N3196, N1531, N381, N1969);
nand NAND2 (N3201, N3193, N2166);
buf BUF1 (N3202, N3194);
buf BUF1 (N3203, N3200);
or OR2 (N3204, N3182, N1709);
nor NOR4 (N3205, N3195, N1563, N2340, N552);
nor NOR3 (N3206, N3204, N1187, N1264);
buf BUF1 (N3207, N3203);
buf BUF1 (N3208, N3190);
nand NAND4 (N3209, N3199, N1563, N2581, N2266);
and AND3 (N3210, N3206, N1887, N1066);
not NOT1 (N3211, N3198);
and AND4 (N3212, N3187, N2119, N466, N518);
xor XOR2 (N3213, N3209, N1932);
buf BUF1 (N3214, N3201);
nand NAND3 (N3215, N3176, N2521, N1356);
or OR3 (N3216, N3208, N448, N566);
and AND3 (N3217, N3207, N2372, N2554);
buf BUF1 (N3218, N3205);
nor NOR2 (N3219, N3216, N2869);
buf BUF1 (N3220, N3218);
not NOT1 (N3221, N3202);
or OR3 (N3222, N3217, N344, N2603);
buf BUF1 (N3223, N3214);
nand NAND3 (N3224, N3215, N1705, N2818);
and AND2 (N3225, N3224, N1658);
xor XOR2 (N3226, N3223, N1448);
buf BUF1 (N3227, N3213);
not NOT1 (N3228, N3221);
xor XOR2 (N3229, N3226, N2918);
nor NOR4 (N3230, N3227, N1127, N2375, N1738);
buf BUF1 (N3231, N3211);
buf BUF1 (N3232, N3212);
nand NAND4 (N3233, N3219, N2411, N2627, N1361);
xor XOR2 (N3234, N3228, N677);
nor NOR4 (N3235, N3231, N772, N1125, N2964);
or OR4 (N3236, N3222, N2739, N1911, N1018);
buf BUF1 (N3237, N3236);
nand NAND2 (N3238, N3229, N2526);
or OR2 (N3239, N3233, N2848);
buf BUF1 (N3240, N3225);
and AND4 (N3241, N3234, N766, N630, N296);
buf BUF1 (N3242, N3235);
xor XOR2 (N3243, N3232, N314);
nor NOR2 (N3244, N3230, N632);
and AND4 (N3245, N3241, N304, N198, N2997);
and AND2 (N3246, N3243, N440);
xor XOR2 (N3247, N3244, N1807);
nor NOR4 (N3248, N3240, N2784, N2603, N2640);
nand NAND2 (N3249, N3238, N242);
and AND4 (N3250, N3248, N1317, N3126, N370);
and AND4 (N3251, N3250, N2999, N17, N1799);
buf BUF1 (N3252, N3239);
nor NOR4 (N3253, N3242, N1478, N687, N1471);
and AND3 (N3254, N3220, N2958, N1679);
nor NOR3 (N3255, N3249, N2135, N542);
buf BUF1 (N3256, N3253);
buf BUF1 (N3257, N3237);
and AND3 (N3258, N3257, N1604, N1175);
nand NAND4 (N3259, N3247, N959, N3184, N1070);
buf BUF1 (N3260, N3256);
not NOT1 (N3261, N3260);
nand NAND3 (N3262, N3245, N438, N2196);
and AND4 (N3263, N3259, N632, N2766, N877);
not NOT1 (N3264, N3252);
or OR4 (N3265, N3210, N1185, N1378, N2340);
and AND2 (N3266, N3258, N754);
xor XOR2 (N3267, N3261, N2183);
not NOT1 (N3268, N3263);
not NOT1 (N3269, N3266);
or OR4 (N3270, N3254, N2467, N791, N2136);
and AND3 (N3271, N3255, N2392, N1204);
xor XOR2 (N3272, N3264, N1701);
nor NOR2 (N3273, N3251, N2655);
or OR2 (N3274, N3269, N750);
nand NAND2 (N3275, N3265, N2754);
or OR3 (N3276, N3273, N489, N766);
nand NAND3 (N3277, N3272, N1425, N693);
nor NOR2 (N3278, N3246, N2112);
not NOT1 (N3279, N3267);
nor NOR4 (N3280, N3279, N845, N2100, N2665);
nand NAND2 (N3281, N3274, N120);
not NOT1 (N3282, N3271);
not NOT1 (N3283, N3282);
or OR4 (N3284, N3283, N154, N1805, N1633);
not NOT1 (N3285, N3280);
buf BUF1 (N3286, N3276);
and AND2 (N3287, N3262, N1908);
not NOT1 (N3288, N3275);
nor NOR4 (N3289, N3278, N2043, N3034, N227);
or OR3 (N3290, N3285, N1023, N1712);
or OR2 (N3291, N3288, N2399);
nand NAND2 (N3292, N3284, N1859);
xor XOR2 (N3293, N3291, N2947);
xor XOR2 (N3294, N3293, N2337);
nand NAND4 (N3295, N3287, N3164, N1881, N2052);
or OR4 (N3296, N3286, N3069, N1372, N1467);
buf BUF1 (N3297, N3289);
nor NOR4 (N3298, N3294, N494, N1458, N2803);
or OR4 (N3299, N3297, N2070, N2708, N879);
buf BUF1 (N3300, N3268);
nand NAND3 (N3301, N3292, N224, N342);
nand NAND2 (N3302, N3296, N186);
buf BUF1 (N3303, N3290);
or OR2 (N3304, N3270, N972);
buf BUF1 (N3305, N3300);
not NOT1 (N3306, N3298);
nand NAND3 (N3307, N3277, N2430, N1935);
xor XOR2 (N3308, N3306, N1085);
nand NAND2 (N3309, N3299, N51);
buf BUF1 (N3310, N3281);
buf BUF1 (N3311, N3305);
xor XOR2 (N3312, N3301, N3172);
buf BUF1 (N3313, N3295);
xor XOR2 (N3314, N3308, N2370);
and AND3 (N3315, N3311, N2439, N1970);
buf BUF1 (N3316, N3307);
not NOT1 (N3317, N3302);
xor XOR2 (N3318, N3303, N2060);
not NOT1 (N3319, N3317);
buf BUF1 (N3320, N3310);
nor NOR2 (N3321, N3320, N1022);
nor NOR2 (N3322, N3319, N2339);
or OR2 (N3323, N3313, N3089);
xor XOR2 (N3324, N3304, N2982);
nor NOR2 (N3325, N3314, N621);
xor XOR2 (N3326, N3315, N838);
buf BUF1 (N3327, N3321);
xor XOR2 (N3328, N3312, N599);
buf BUF1 (N3329, N3324);
xor XOR2 (N3330, N3323, N774);
not NOT1 (N3331, N3327);
not NOT1 (N3332, N3330);
buf BUF1 (N3333, N3316);
nand NAND3 (N3334, N3326, N559, N3063);
xor XOR2 (N3335, N3334, N2901);
xor XOR2 (N3336, N3332, N2326);
nor NOR4 (N3337, N3333, N1972, N1386, N871);
xor XOR2 (N3338, N3322, N527);
not NOT1 (N3339, N3325);
xor XOR2 (N3340, N3335, N786);
buf BUF1 (N3341, N3338);
or OR3 (N3342, N3336, N3309, N2528);
nor NOR3 (N3343, N3089, N455, N562);
buf BUF1 (N3344, N3343);
or OR2 (N3345, N3342, N3064);
and AND2 (N3346, N3328, N1904);
and AND4 (N3347, N3344, N235, N2499, N1941);
or OR4 (N3348, N3347, N1795, N3142, N1581);
or OR4 (N3349, N3341, N2688, N1327, N1012);
and AND3 (N3350, N3331, N2003, N967);
nor NOR3 (N3351, N3345, N1215, N2287);
and AND4 (N3352, N3318, N2958, N781, N1196);
nor NOR4 (N3353, N3351, N554, N1072, N1193);
buf BUF1 (N3354, N3329);
nand NAND4 (N3355, N3353, N2245, N1578, N2559);
buf BUF1 (N3356, N3352);
nand NAND2 (N3357, N3340, N1203);
nor NOR2 (N3358, N3349, N1804);
and AND3 (N3359, N3348, N2590, N2005);
buf BUF1 (N3360, N3355);
and AND3 (N3361, N3350, N3104, N1105);
nor NOR3 (N3362, N3337, N649, N3118);
buf BUF1 (N3363, N3358);
or OR4 (N3364, N3354, N2999, N1864, N164);
nor NOR2 (N3365, N3357, N431);
and AND2 (N3366, N3361, N3147);
and AND4 (N3367, N3356, N3327, N2180, N150);
nor NOR3 (N3368, N3339, N2790, N2296);
nand NAND4 (N3369, N3362, N785, N2764, N3073);
nor NOR3 (N3370, N3366, N2505, N851);
nand NAND4 (N3371, N3363, N2500, N3130, N523);
buf BUF1 (N3372, N3364);
nand NAND4 (N3373, N3360, N2906, N1934, N1515);
and AND3 (N3374, N3367, N3082, N2548);
buf BUF1 (N3375, N3359);
xor XOR2 (N3376, N3373, N183);
nand NAND3 (N3377, N3369, N661, N2789);
buf BUF1 (N3378, N3368);
or OR4 (N3379, N3372, N468, N608, N2553);
not NOT1 (N3380, N3365);
nor NOR3 (N3381, N3370, N2997, N1227);
nand NAND3 (N3382, N3371, N2104, N2883);
xor XOR2 (N3383, N3374, N634);
buf BUF1 (N3384, N3383);
and AND2 (N3385, N3376, N3278);
nand NAND4 (N3386, N3375, N2880, N1499, N2642);
nor NOR4 (N3387, N3381, N511, N2610, N2811);
or OR3 (N3388, N3385, N2458, N848);
nor NOR4 (N3389, N3386, N1516, N2838, N2077);
xor XOR2 (N3390, N3379, N63);
nor NOR2 (N3391, N3384, N2639);
nor NOR2 (N3392, N3382, N1064);
nand NAND2 (N3393, N3387, N668);
not NOT1 (N3394, N3390);
buf BUF1 (N3395, N3377);
nor NOR2 (N3396, N3380, N1770);
or OR3 (N3397, N3395, N3189, N2342);
not NOT1 (N3398, N3397);
nor NOR3 (N3399, N3392, N2054, N695);
xor XOR2 (N3400, N3391, N747);
xor XOR2 (N3401, N3346, N616);
and AND3 (N3402, N3393, N922, N2442);
and AND4 (N3403, N3388, N1141, N122, N2979);
nand NAND2 (N3404, N3403, N2487);
nor NOR3 (N3405, N3402, N255, N898);
nand NAND4 (N3406, N3396, N461, N1260, N1918);
nor NOR2 (N3407, N3394, N1807);
nor NOR4 (N3408, N3378, N2401, N923, N1621);
nand NAND3 (N3409, N3399, N1539, N762);
and AND4 (N3410, N3409, N2962, N2771, N2863);
nand NAND2 (N3411, N3401, N2319);
xor XOR2 (N3412, N3411, N568);
xor XOR2 (N3413, N3412, N3383);
and AND2 (N3414, N3406, N1069);
not NOT1 (N3415, N3398);
xor XOR2 (N3416, N3413, N1907);
not NOT1 (N3417, N3414);
xor XOR2 (N3418, N3405, N3322);
and AND2 (N3419, N3410, N3263);
buf BUF1 (N3420, N3416);
or OR3 (N3421, N3408, N1026, N1730);
xor XOR2 (N3422, N3389, N687);
nand NAND2 (N3423, N3404, N858);
xor XOR2 (N3424, N3422, N1502);
nand NAND3 (N3425, N3419, N3063, N277);
buf BUF1 (N3426, N3417);
buf BUF1 (N3427, N3426);
and AND3 (N3428, N3423, N3050, N2814);
buf BUF1 (N3429, N3425);
or OR3 (N3430, N3424, N1180, N349);
nand NAND3 (N3431, N3418, N312, N3023);
and AND4 (N3432, N3400, N2470, N70, N2908);
not NOT1 (N3433, N3432);
nand NAND2 (N3434, N3427, N1501);
nor NOR3 (N3435, N3420, N2107, N301);
not NOT1 (N3436, N3407);
nand NAND2 (N3437, N3434, N3317);
or OR4 (N3438, N3430, N1690, N718, N2253);
xor XOR2 (N3439, N3429, N1071);
xor XOR2 (N3440, N3415, N1740);
or OR3 (N3441, N3440, N746, N653);
nand NAND2 (N3442, N3435, N1850);
or OR2 (N3443, N3436, N2666);
buf BUF1 (N3444, N3421);
not NOT1 (N3445, N3443);
buf BUF1 (N3446, N3428);
xor XOR2 (N3447, N3438, N733);
or OR3 (N3448, N3441, N2333, N3332);
and AND3 (N3449, N3444, N1727, N606);
nor NOR4 (N3450, N3446, N2090, N2401, N2512);
or OR3 (N3451, N3437, N719, N1026);
and AND2 (N3452, N3451, N2969);
and AND4 (N3453, N3433, N1456, N920, N1185);
buf BUF1 (N3454, N3445);
and AND4 (N3455, N3448, N2080, N418, N1800);
xor XOR2 (N3456, N3452, N163);
xor XOR2 (N3457, N3456, N2361);
or OR4 (N3458, N3450, N315, N1908, N3190);
buf BUF1 (N3459, N3447);
buf BUF1 (N3460, N3449);
not NOT1 (N3461, N3455);
nand NAND3 (N3462, N3431, N1377, N2150);
or OR3 (N3463, N3457, N3389, N887);
and AND3 (N3464, N3461, N1108, N2690);
and AND2 (N3465, N3459, N980);
buf BUF1 (N3466, N3463);
nand NAND3 (N3467, N3453, N1482, N1200);
nor NOR3 (N3468, N3467, N2235, N369);
buf BUF1 (N3469, N3468);
and AND4 (N3470, N3469, N1276, N2885, N2361);
buf BUF1 (N3471, N3462);
nand NAND4 (N3472, N3442, N2330, N2717, N2181);
xor XOR2 (N3473, N3471, N2470);
buf BUF1 (N3474, N3458);
nor NOR4 (N3475, N3470, N2013, N1696, N2000);
not NOT1 (N3476, N3473);
not NOT1 (N3477, N3464);
and AND2 (N3478, N3474, N3463);
not NOT1 (N3479, N3477);
nor NOR4 (N3480, N3439, N1763, N748, N1627);
buf BUF1 (N3481, N3454);
or OR2 (N3482, N3472, N180);
buf BUF1 (N3483, N3475);
nor NOR3 (N3484, N3465, N1730, N2070);
nor NOR3 (N3485, N3480, N1347, N2274);
xor XOR2 (N3486, N3476, N2972);
or OR3 (N3487, N3460, N3427, N917);
nand NAND4 (N3488, N3479, N1009, N2271, N2261);
xor XOR2 (N3489, N3486, N630);
and AND3 (N3490, N3478, N104, N203);
or OR4 (N3491, N3485, N1312, N2856, N2770);
nor NOR4 (N3492, N3491, N3423, N2438, N1164);
xor XOR2 (N3493, N3481, N1312);
not NOT1 (N3494, N3492);
not NOT1 (N3495, N3489);
and AND4 (N3496, N3483, N2967, N143, N931);
buf BUF1 (N3497, N3493);
not NOT1 (N3498, N3488);
xor XOR2 (N3499, N3497, N2586);
nor NOR3 (N3500, N3484, N2311, N3182);
and AND4 (N3501, N3466, N1770, N3351, N1448);
nor NOR4 (N3502, N3487, N2648, N2397, N286);
nand NAND3 (N3503, N3494, N1558, N1719);
not NOT1 (N3504, N3502);
nor NOR2 (N3505, N3496, N2551);
xor XOR2 (N3506, N3482, N1668);
and AND3 (N3507, N3506, N237, N2237);
nand NAND4 (N3508, N3507, N1317, N553, N2184);
xor XOR2 (N3509, N3505, N2164);
nand NAND3 (N3510, N3500, N1214, N2498);
and AND4 (N3511, N3510, N2732, N3288, N266);
nor NOR3 (N3512, N3490, N602, N292);
nand NAND4 (N3513, N3498, N3049, N2077, N109);
nor NOR2 (N3514, N3512, N782);
buf BUF1 (N3515, N3508);
buf BUF1 (N3516, N3509);
not NOT1 (N3517, N3515);
or OR4 (N3518, N3517, N3366, N267, N1347);
not NOT1 (N3519, N3514);
not NOT1 (N3520, N3504);
or OR3 (N3521, N3499, N3264, N3453);
xor XOR2 (N3522, N3520, N3084);
nand NAND2 (N3523, N3495, N1624);
and AND3 (N3524, N3513, N2853, N2504);
and AND4 (N3525, N3518, N1773, N1275, N606);
nand NAND3 (N3526, N3521, N2822, N2223);
or OR2 (N3527, N3524, N1129);
buf BUF1 (N3528, N3516);
or OR4 (N3529, N3503, N1817, N821, N1564);
nand NAND2 (N3530, N3526, N3368);
and AND3 (N3531, N3523, N2047, N1295);
and AND4 (N3532, N3501, N2354, N3030, N2693);
buf BUF1 (N3533, N3530);
nand NAND3 (N3534, N3528, N1485, N2210);
buf BUF1 (N3535, N3533);
nand NAND2 (N3536, N3525, N1983);
not NOT1 (N3537, N3527);
or OR4 (N3538, N3519, N2253, N1637, N3410);
nand NAND2 (N3539, N3537, N573);
or OR4 (N3540, N3538, N1898, N64, N1946);
nor NOR2 (N3541, N3531, N3303);
and AND4 (N3542, N3540, N656, N3215, N3019);
or OR3 (N3543, N3522, N1291, N2079);
and AND2 (N3544, N3532, N1758);
or OR4 (N3545, N3534, N3192, N642, N1651);
or OR2 (N3546, N3544, N1488);
or OR3 (N3547, N3545, N883, N1056);
xor XOR2 (N3548, N3536, N724);
not NOT1 (N3549, N3542);
nand NAND2 (N3550, N3535, N312);
and AND3 (N3551, N3547, N3491, N549);
nand NAND3 (N3552, N3511, N1495, N1880);
xor XOR2 (N3553, N3550, N1306);
nor NOR2 (N3554, N3539, N1096);
buf BUF1 (N3555, N3551);
nor NOR3 (N3556, N3555, N3097, N568);
not NOT1 (N3557, N3549);
nor NOR4 (N3558, N3554, N351, N1062, N3193);
and AND3 (N3559, N3543, N3310, N296);
or OR3 (N3560, N3541, N1746, N424);
not NOT1 (N3561, N3552);
xor XOR2 (N3562, N3560, N1459);
nand NAND2 (N3563, N3559, N329);
not NOT1 (N3564, N3558);
not NOT1 (N3565, N3557);
and AND3 (N3566, N3548, N2543, N3193);
and AND4 (N3567, N3566, N3289, N1646, N917);
and AND2 (N3568, N3556, N806);
nor NOR4 (N3569, N3553, N1528, N1895, N3191);
not NOT1 (N3570, N3563);
and AND3 (N3571, N3561, N1530, N1591);
not NOT1 (N3572, N3564);
nand NAND3 (N3573, N3567, N1351, N2960);
or OR4 (N3574, N3570, N2729, N1847, N64);
and AND4 (N3575, N3574, N2791, N3187, N2702);
xor XOR2 (N3576, N3573, N2840);
nor NOR4 (N3577, N3572, N1090, N371, N2535);
xor XOR2 (N3578, N3577, N2441);
not NOT1 (N3579, N3565);
xor XOR2 (N3580, N3579, N1574);
xor XOR2 (N3581, N3569, N834);
buf BUF1 (N3582, N3581);
nor NOR4 (N3583, N3568, N1377, N436, N2015);
and AND3 (N3584, N3582, N212, N2415);
nor NOR2 (N3585, N3562, N1033);
or OR4 (N3586, N3571, N174, N962, N2232);
nor NOR4 (N3587, N3578, N2446, N1070, N1631);
nand NAND4 (N3588, N3575, N2416, N3054, N36);
or OR4 (N3589, N3588, N1297, N260, N3136);
nand NAND2 (N3590, N3529, N736);
nand NAND2 (N3591, N3586, N2762);
nand NAND3 (N3592, N3583, N3054, N2188);
buf BUF1 (N3593, N3546);
xor XOR2 (N3594, N3587, N1906);
not NOT1 (N3595, N3592);
xor XOR2 (N3596, N3584, N3379);
nor NOR2 (N3597, N3589, N460);
nor NOR3 (N3598, N3596, N389, N3558);
xor XOR2 (N3599, N3585, N1451);
nand NAND4 (N3600, N3598, N880, N2366, N2028);
xor XOR2 (N3601, N3597, N629);
or OR4 (N3602, N3600, N296, N754, N534);
nand NAND4 (N3603, N3602, N1165, N25, N574);
buf BUF1 (N3604, N3590);
or OR2 (N3605, N3593, N202);
nor NOR4 (N3606, N3603, N876, N1651, N230);
nor NOR2 (N3607, N3580, N1230);
nor NOR4 (N3608, N3607, N292, N2790, N875);
or OR4 (N3609, N3606, N164, N227, N3486);
or OR3 (N3610, N3599, N2237, N2261);
nor NOR4 (N3611, N3594, N1236, N3428, N1416);
nor NOR4 (N3612, N3595, N2266, N1848, N135);
buf BUF1 (N3613, N3605);
not NOT1 (N3614, N3604);
and AND3 (N3615, N3613, N56, N2157);
not NOT1 (N3616, N3576);
not NOT1 (N3617, N3616);
nand NAND2 (N3618, N3614, N1263);
xor XOR2 (N3619, N3611, N2025);
buf BUF1 (N3620, N3601);
nor NOR3 (N3621, N3608, N2810, N1106);
nand NAND2 (N3622, N3615, N932);
nor NOR3 (N3623, N3619, N1023, N1994);
and AND2 (N3624, N3621, N1537);
nor NOR3 (N3625, N3610, N1919, N1217);
or OR2 (N3626, N3624, N979);
buf BUF1 (N3627, N3618);
nor NOR2 (N3628, N3609, N164);
nand NAND3 (N3629, N3622, N1029, N605);
nand NAND3 (N3630, N3625, N2821, N2933);
nor NOR3 (N3631, N3627, N2112, N1429);
not NOT1 (N3632, N3628);
not NOT1 (N3633, N3630);
not NOT1 (N3634, N3617);
xor XOR2 (N3635, N3626, N3004);
nor NOR3 (N3636, N3591, N2669, N966);
nand NAND4 (N3637, N3633, N610, N408, N1525);
xor XOR2 (N3638, N3620, N392);
or OR4 (N3639, N3636, N1588, N2197, N2260);
xor XOR2 (N3640, N3612, N826);
nand NAND4 (N3641, N3631, N2984, N2785, N2655);
and AND4 (N3642, N3639, N676, N3469, N1791);
or OR4 (N3643, N3623, N817, N2319, N161);
and AND3 (N3644, N3642, N2108, N412);
or OR2 (N3645, N3635, N2805);
buf BUF1 (N3646, N3643);
or OR4 (N3647, N3634, N817, N2650, N3547);
nor NOR4 (N3648, N3638, N302, N3212, N1762);
and AND3 (N3649, N3646, N1233, N2691);
or OR2 (N3650, N3641, N1550);
xor XOR2 (N3651, N3637, N3524);
and AND2 (N3652, N3644, N451);
not NOT1 (N3653, N3629);
and AND3 (N3654, N3651, N1322, N1088);
nor NOR3 (N3655, N3653, N562, N527);
buf BUF1 (N3656, N3655);
or OR3 (N3657, N3640, N3222, N1132);
nor NOR4 (N3658, N3648, N2496, N3446, N2792);
or OR3 (N3659, N3657, N3420, N659);
xor XOR2 (N3660, N3647, N2942);
and AND2 (N3661, N3659, N960);
or OR2 (N3662, N3645, N2638);
nor NOR4 (N3663, N3650, N2456, N2017, N2525);
nand NAND3 (N3664, N3656, N1934, N694);
not NOT1 (N3665, N3649);
buf BUF1 (N3666, N3664);
or OR3 (N3667, N3666, N598, N3164);
and AND2 (N3668, N3661, N2949);
nand NAND2 (N3669, N3652, N2317);
nand NAND2 (N3670, N3654, N107);
xor XOR2 (N3671, N3665, N3185);
not NOT1 (N3672, N3660);
nand NAND3 (N3673, N3658, N2715, N1005);
nand NAND4 (N3674, N3632, N1361, N2257, N2301);
or OR3 (N3675, N3670, N1571, N1203);
xor XOR2 (N3676, N3672, N3160);
xor XOR2 (N3677, N3675, N2410);
buf BUF1 (N3678, N3668);
nand NAND3 (N3679, N3673, N1445, N2043);
xor XOR2 (N3680, N3678, N314);
and AND4 (N3681, N3677, N577, N2730, N97);
and AND3 (N3682, N3680, N1329, N2933);
nand NAND2 (N3683, N3669, N2783);
buf BUF1 (N3684, N3676);
nand NAND2 (N3685, N3667, N55);
and AND2 (N3686, N3679, N966);
or OR4 (N3687, N3684, N2770, N2807, N3098);
or OR3 (N3688, N3671, N2752, N2554);
not NOT1 (N3689, N3663);
nand NAND2 (N3690, N3662, N2417);
nor NOR4 (N3691, N3689, N1774, N2244, N1205);
nor NOR2 (N3692, N3685, N3272);
nand NAND3 (N3693, N3682, N2011, N110);
or OR3 (N3694, N3688, N1353, N796);
xor XOR2 (N3695, N3693, N3602);
or OR4 (N3696, N3687, N1574, N63, N3165);
xor XOR2 (N3697, N3686, N1927);
nand NAND4 (N3698, N3681, N339, N1899, N1377);
or OR2 (N3699, N3692, N1462);
buf BUF1 (N3700, N3695);
nand NAND3 (N3701, N3691, N1198, N1595);
or OR3 (N3702, N3696, N1827, N1688);
or OR4 (N3703, N3701, N578, N2355, N116);
and AND3 (N3704, N3698, N2343, N1850);
xor XOR2 (N3705, N3690, N1913);
not NOT1 (N3706, N3699);
buf BUF1 (N3707, N3700);
nand NAND2 (N3708, N3707, N1386);
buf BUF1 (N3709, N3705);
and AND2 (N3710, N3704, N2208);
not NOT1 (N3711, N3694);
xor XOR2 (N3712, N3697, N1835);
or OR2 (N3713, N3674, N2441);
and AND2 (N3714, N3703, N3515);
or OR2 (N3715, N3711, N1193);
and AND3 (N3716, N3713, N1465, N2153);
and AND4 (N3717, N3702, N2109, N925, N1673);
or OR3 (N3718, N3715, N1329, N1966);
not NOT1 (N3719, N3709);
xor XOR2 (N3720, N3712, N2956);
nand NAND2 (N3721, N3714, N1441);
not NOT1 (N3722, N3708);
not NOT1 (N3723, N3719);
buf BUF1 (N3724, N3683);
nand NAND3 (N3725, N3721, N1099, N1097);
and AND4 (N3726, N3722, N3621, N3152, N1671);
or OR3 (N3727, N3710, N43, N3669);
or OR2 (N3728, N3726, N395);
or OR3 (N3729, N3720, N1850, N307);
xor XOR2 (N3730, N3723, N2268);
or OR4 (N3731, N3729, N1192, N820, N1366);
not NOT1 (N3732, N3728);
nand NAND2 (N3733, N3706, N2008);
buf BUF1 (N3734, N3732);
buf BUF1 (N3735, N3727);
xor XOR2 (N3736, N3730, N2684);
buf BUF1 (N3737, N3718);
buf BUF1 (N3738, N3736);
nand NAND3 (N3739, N3738, N3044, N933);
nand NAND2 (N3740, N3735, N1879);
or OR3 (N3741, N3740, N1657, N1900);
and AND4 (N3742, N3739, N1372, N3433, N83);
nand NAND4 (N3743, N3734, N3702, N3724, N2885);
buf BUF1 (N3744, N412);
buf BUF1 (N3745, N3741);
or OR3 (N3746, N3725, N2788, N3223);
or OR2 (N3747, N3746, N3065);
nand NAND3 (N3748, N3743, N1478, N1411);
buf BUF1 (N3749, N3731);
xor XOR2 (N3750, N3747, N817);
xor XOR2 (N3751, N3742, N1269);
nor NOR4 (N3752, N3749, N2397, N1794, N2577);
not NOT1 (N3753, N3737);
not NOT1 (N3754, N3751);
xor XOR2 (N3755, N3716, N3413);
and AND2 (N3756, N3748, N1155);
nand NAND2 (N3757, N3754, N1671);
not NOT1 (N3758, N3717);
nor NOR2 (N3759, N3757, N3425);
and AND2 (N3760, N3755, N2036);
nand NAND4 (N3761, N3759, N177, N2874, N1466);
not NOT1 (N3762, N3744);
and AND4 (N3763, N3750, N396, N2703, N334);
nor NOR2 (N3764, N3763, N1588);
nor NOR2 (N3765, N3762, N2267);
nand NAND2 (N3766, N3765, N1392);
and AND4 (N3767, N3761, N2331, N3122, N109);
xor XOR2 (N3768, N3764, N2273);
and AND3 (N3769, N3758, N3026, N3254);
nor NOR4 (N3770, N3768, N1982, N221, N1537);
buf BUF1 (N3771, N3752);
buf BUF1 (N3772, N3769);
nor NOR2 (N3773, N3771, N1017);
buf BUF1 (N3774, N3770);
nor NOR3 (N3775, N3733, N3628, N2570);
not NOT1 (N3776, N3745);
nand NAND4 (N3777, N3760, N218, N2549, N770);
buf BUF1 (N3778, N3776);
xor XOR2 (N3779, N3774, N1913);
not NOT1 (N3780, N3779);
and AND4 (N3781, N3778, N1026, N848, N1574);
nand NAND3 (N3782, N3775, N1317, N1002);
or OR4 (N3783, N3753, N1577, N109, N2089);
and AND3 (N3784, N3766, N2191, N1327);
nand NAND4 (N3785, N3780, N2524, N472, N236);
nand NAND4 (N3786, N3772, N5, N209, N150);
nand NAND4 (N3787, N3777, N3207, N3324, N49);
or OR2 (N3788, N3783, N13);
not NOT1 (N3789, N3767);
nand NAND4 (N3790, N3786, N162, N445, N3038);
xor XOR2 (N3791, N3784, N1806);
not NOT1 (N3792, N3773);
and AND3 (N3793, N3788, N461, N1397);
or OR2 (N3794, N3782, N855);
and AND4 (N3795, N3789, N3384, N2892, N3043);
not NOT1 (N3796, N3795);
xor XOR2 (N3797, N3781, N3708);
nand NAND4 (N3798, N3791, N3261, N68, N3618);
and AND3 (N3799, N3793, N2745, N3517);
buf BUF1 (N3800, N3794);
and AND3 (N3801, N3785, N1638, N1279);
xor XOR2 (N3802, N3797, N2783);
or OR4 (N3803, N3790, N77, N653, N323);
xor XOR2 (N3804, N3802, N963);
not NOT1 (N3805, N3756);
nand NAND3 (N3806, N3801, N1111, N2194);
nor NOR3 (N3807, N3796, N1780, N2979);
nor NOR4 (N3808, N3804, N3265, N2594, N2980);
and AND3 (N3809, N3808, N1717, N2904);
and AND4 (N3810, N3787, N1045, N2869, N3793);
xor XOR2 (N3811, N3807, N384);
nor NOR4 (N3812, N3803, N2730, N182, N1724);
not NOT1 (N3813, N3805);
not NOT1 (N3814, N3810);
not NOT1 (N3815, N3798);
nand NAND4 (N3816, N3806, N1506, N2154, N873);
or OR4 (N3817, N3799, N48, N114, N2267);
not NOT1 (N3818, N3817);
nor NOR4 (N3819, N3812, N1805, N2909, N2303);
buf BUF1 (N3820, N3813);
nor NOR2 (N3821, N3809, N851);
or OR3 (N3822, N3792, N2028, N2847);
nor NOR3 (N3823, N3800, N3046, N3571);
nand NAND3 (N3824, N3822, N3636, N2987);
or OR4 (N3825, N3820, N429, N1482, N3361);
nand NAND4 (N3826, N3824, N509, N1700, N3242);
buf BUF1 (N3827, N3819);
not NOT1 (N3828, N3826);
nor NOR3 (N3829, N3827, N1347, N565);
xor XOR2 (N3830, N3814, N2062);
nor NOR2 (N3831, N3830, N300);
nor NOR4 (N3832, N3811, N1723, N1657, N1098);
nand NAND3 (N3833, N3818, N1557, N892);
not NOT1 (N3834, N3832);
or OR3 (N3835, N3833, N1610, N812);
xor XOR2 (N3836, N3823, N2508);
nor NOR3 (N3837, N3835, N3530, N3317);
and AND4 (N3838, N3815, N1190, N2117, N3103);
nor NOR4 (N3839, N3836, N2661, N2738, N8);
or OR2 (N3840, N3839, N1322);
nand NAND3 (N3841, N3831, N1845, N1214);
and AND4 (N3842, N3841, N2273, N1227, N2769);
not NOT1 (N3843, N3842);
and AND2 (N3844, N3837, N1512);
or OR2 (N3845, N3843, N1690);
xor XOR2 (N3846, N3844, N1734);
and AND3 (N3847, N3816, N438, N786);
and AND4 (N3848, N3840, N2120, N3633, N1474);
not NOT1 (N3849, N3847);
buf BUF1 (N3850, N3846);
xor XOR2 (N3851, N3850, N1206);
xor XOR2 (N3852, N3845, N2126);
and AND4 (N3853, N3851, N2828, N3497, N2612);
buf BUF1 (N3854, N3852);
buf BUF1 (N3855, N3853);
nor NOR3 (N3856, N3855, N3409, N3461);
nand NAND4 (N3857, N3854, N2813, N3505, N959);
xor XOR2 (N3858, N3849, N3237);
and AND4 (N3859, N3857, N3095, N3215, N1219);
xor XOR2 (N3860, N3856, N3131);
or OR2 (N3861, N3859, N1663);
buf BUF1 (N3862, N3838);
or OR2 (N3863, N3834, N1206);
or OR3 (N3864, N3860, N1026, N2490);
or OR2 (N3865, N3863, N3856);
buf BUF1 (N3866, N3864);
nor NOR4 (N3867, N3862, N1047, N578, N908);
and AND4 (N3868, N3867, N867, N248, N501);
not NOT1 (N3869, N3828);
nand NAND2 (N3870, N3829, N2224);
and AND3 (N3871, N3866, N2357, N2501);
buf BUF1 (N3872, N3848);
not NOT1 (N3873, N3821);
xor XOR2 (N3874, N3858, N3658);
nor NOR3 (N3875, N3861, N1421, N3624);
nand NAND4 (N3876, N3872, N3560, N1232, N2885);
and AND4 (N3877, N3825, N128, N2819, N582);
nor NOR4 (N3878, N3876, N298, N88, N3169);
and AND2 (N3879, N3869, N3080);
buf BUF1 (N3880, N3874);
or OR4 (N3881, N3865, N2039, N823, N735);
buf BUF1 (N3882, N3871);
buf BUF1 (N3883, N3881);
xor XOR2 (N3884, N3877, N1920);
xor XOR2 (N3885, N3882, N3739);
nor NOR3 (N3886, N3884, N3124, N1469);
nand NAND3 (N3887, N3870, N3575, N843);
nand NAND4 (N3888, N3868, N743, N2146, N1210);
and AND2 (N3889, N3887, N3335);
nor NOR4 (N3890, N3888, N3086, N1077, N2448);
nand NAND3 (N3891, N3873, N330, N1121);
buf BUF1 (N3892, N3875);
xor XOR2 (N3893, N3883, N3367);
xor XOR2 (N3894, N3885, N2959);
xor XOR2 (N3895, N3879, N1455);
or OR4 (N3896, N3880, N930, N1647, N1613);
buf BUF1 (N3897, N3895);
not NOT1 (N3898, N3878);
nand NAND3 (N3899, N3889, N563, N1124);
nor NOR3 (N3900, N3886, N2838, N3171);
or OR2 (N3901, N3899, N1819);
or OR2 (N3902, N3891, N587);
not NOT1 (N3903, N3890);
not NOT1 (N3904, N3902);
nand NAND3 (N3905, N3898, N3346, N1261);
buf BUF1 (N3906, N3903);
or OR3 (N3907, N3896, N35, N331);
xor XOR2 (N3908, N3904, N1421);
or OR2 (N3909, N3892, N2686);
xor XOR2 (N3910, N3908, N2024);
and AND2 (N3911, N3905, N350);
buf BUF1 (N3912, N3900);
not NOT1 (N3913, N3907);
buf BUF1 (N3914, N3912);
or OR2 (N3915, N3897, N3895);
or OR2 (N3916, N3915, N701);
and AND2 (N3917, N3909, N1432);
or OR3 (N3918, N3916, N2213, N96);
or OR4 (N3919, N3911, N357, N2729, N226);
and AND3 (N3920, N3919, N2636, N2940);
or OR4 (N3921, N3920, N1391, N957, N420);
nor NOR4 (N3922, N3914, N1174, N229, N1368);
not NOT1 (N3923, N3922);
nor NOR4 (N3924, N3901, N3749, N2573, N805);
buf BUF1 (N3925, N3913);
nand NAND4 (N3926, N3924, N2928, N2507, N910);
xor XOR2 (N3927, N3917, N825);
or OR4 (N3928, N3927, N3378, N3318, N1741);
and AND2 (N3929, N3893, N787);
nor NOR3 (N3930, N3894, N1988, N2062);
buf BUF1 (N3931, N3923);
nand NAND4 (N3932, N3930, N2257, N2063, N2542);
not NOT1 (N3933, N3925);
buf BUF1 (N3934, N3910);
or OR4 (N3935, N3933, N1468, N1045, N3920);
xor XOR2 (N3936, N3934, N3905);
buf BUF1 (N3937, N3932);
and AND2 (N3938, N3928, N1512);
nand NAND2 (N3939, N3937, N791);
not NOT1 (N3940, N3921);
xor XOR2 (N3941, N3929, N2967);
or OR3 (N3942, N3935, N1611, N3471);
buf BUF1 (N3943, N3926);
nand NAND2 (N3944, N3936, N161);
nand NAND4 (N3945, N3940, N731, N115, N859);
and AND3 (N3946, N3942, N2613, N729);
or OR2 (N3947, N3946, N98);
xor XOR2 (N3948, N3918, N1569);
not NOT1 (N3949, N3939);
nor NOR2 (N3950, N3941, N3797);
not NOT1 (N3951, N3931);
or OR3 (N3952, N3943, N2619, N709);
and AND3 (N3953, N3947, N3638, N485);
xor XOR2 (N3954, N3950, N2972);
buf BUF1 (N3955, N3906);
xor XOR2 (N3956, N3952, N3513);
nand NAND4 (N3957, N3956, N1606, N2521, N1099);
or OR2 (N3958, N3951, N425);
buf BUF1 (N3959, N3948);
or OR4 (N3960, N3958, N910, N2601, N3518);
buf BUF1 (N3961, N3944);
buf BUF1 (N3962, N3959);
xor XOR2 (N3963, N3957, N369);
buf BUF1 (N3964, N3960);
xor XOR2 (N3965, N3964, N604);
nor NOR4 (N3966, N3961, N637, N3545, N1780);
nand NAND4 (N3967, N3949, N1540, N10, N1220);
not NOT1 (N3968, N3965);
buf BUF1 (N3969, N3945);
xor XOR2 (N3970, N3968, N116);
nor NOR2 (N3971, N3966, N2262);
nor NOR3 (N3972, N3971, N858, N2787);
nand NAND2 (N3973, N3938, N3194);
not NOT1 (N3974, N3967);
nor NOR4 (N3975, N3954, N1248, N1548, N2581);
buf BUF1 (N3976, N3955);
and AND2 (N3977, N3963, N3555);
or OR3 (N3978, N3972, N3308, N3721);
nand NAND4 (N3979, N3962, N548, N2432, N3264);
not NOT1 (N3980, N3977);
buf BUF1 (N3981, N3978);
nand NAND2 (N3982, N3969, N3190);
not NOT1 (N3983, N3979);
or OR3 (N3984, N3974, N2105, N677);
nor NOR4 (N3985, N3970, N1952, N744, N3017);
or OR4 (N3986, N3981, N1095, N2488, N684);
or OR4 (N3987, N3986, N1334, N20, N2832);
buf BUF1 (N3988, N3985);
not NOT1 (N3989, N3983);
not NOT1 (N3990, N3980);
nand NAND2 (N3991, N3973, N1787);
and AND2 (N3992, N3975, N201);
not NOT1 (N3993, N3987);
nor NOR2 (N3994, N3990, N2535);
nand NAND2 (N3995, N3994, N3615);
nor NOR3 (N3996, N3988, N57, N2313);
nor NOR2 (N3997, N3984, N359);
and AND2 (N3998, N3991, N3550);
or OR2 (N3999, N3997, N3093);
buf BUF1 (N4000, N3953);
not NOT1 (N4001, N3996);
buf BUF1 (N4002, N3999);
and AND4 (N4003, N3993, N286, N2665, N1806);
and AND2 (N4004, N3995, N2611);
or OR3 (N4005, N3976, N695, N2839);
or OR2 (N4006, N3989, N3750);
and AND2 (N4007, N3982, N767);
xor XOR2 (N4008, N4000, N1749);
nor NOR3 (N4009, N4004, N2758, N2104);
nand NAND4 (N4010, N4001, N1366, N2784, N3084);
not NOT1 (N4011, N4010);
xor XOR2 (N4012, N3998, N2057);
nor NOR2 (N4013, N4005, N2822);
nand NAND3 (N4014, N4003, N716, N3094);
xor XOR2 (N4015, N4011, N1199);
nor NOR2 (N4016, N4015, N3507);
xor XOR2 (N4017, N3992, N2309);
xor XOR2 (N4018, N4014, N1763);
nor NOR2 (N4019, N4007, N2644);
nand NAND2 (N4020, N4013, N2188);
nor NOR4 (N4021, N4019, N3227, N1501, N2545);
nor NOR3 (N4022, N4008, N3347, N1007);
xor XOR2 (N4023, N4016, N171);
nor NOR3 (N4024, N4018, N1453, N4013);
and AND4 (N4025, N4021, N3739, N196, N699);
and AND2 (N4026, N4006, N882);
xor XOR2 (N4027, N4026, N3156);
nand NAND3 (N4028, N4023, N3629, N3656);
nor NOR2 (N4029, N4024, N3355);
xor XOR2 (N4030, N4025, N658);
and AND3 (N4031, N4002, N2209, N1085);
nor NOR2 (N4032, N4031, N3182);
or OR3 (N4033, N4020, N1783, N2961);
not NOT1 (N4034, N4030);
buf BUF1 (N4035, N4032);
nor NOR2 (N4036, N4034, N2181);
or OR3 (N4037, N4012, N1703, N3703);
buf BUF1 (N4038, N4028);
nor NOR3 (N4039, N4022, N1886, N2974);
nand NAND2 (N4040, N4009, N94);
buf BUF1 (N4041, N4036);
xor XOR2 (N4042, N4035, N1659);
xor XOR2 (N4043, N4027, N148);
buf BUF1 (N4044, N4017);
not NOT1 (N4045, N4039);
nor NOR2 (N4046, N4043, N1657);
buf BUF1 (N4047, N4041);
not NOT1 (N4048, N4046);
and AND3 (N4049, N4044, N2318, N2305);
or OR2 (N4050, N4038, N3178);
xor XOR2 (N4051, N4040, N2401);
buf BUF1 (N4052, N4029);
nand NAND3 (N4053, N4045, N1786, N2239);
nor NOR3 (N4054, N4052, N260, N3756);
nor NOR2 (N4055, N4037, N3579);
or OR3 (N4056, N4042, N347, N602);
nand NAND2 (N4057, N4055, N2318);
nor NOR2 (N4058, N4049, N2237);
nand NAND4 (N4059, N4056, N1150, N3409, N1859);
or OR3 (N4060, N4057, N1538, N1885);
buf BUF1 (N4061, N4060);
nand NAND3 (N4062, N4054, N1860, N2433);
and AND3 (N4063, N4047, N523, N3400);
nor NOR3 (N4064, N4059, N3499, N634);
or OR4 (N4065, N4053, N4050, N719, N2510);
or OR3 (N4066, N3617, N1590, N2933);
and AND3 (N4067, N4064, N2353, N27);
xor XOR2 (N4068, N4062, N1654);
or OR3 (N4069, N4061, N2121, N1436);
xor XOR2 (N4070, N4033, N993);
nor NOR4 (N4071, N4068, N3933, N2239, N324);
buf BUF1 (N4072, N4070);
nor NOR4 (N4073, N4072, N2502, N741, N2872);
buf BUF1 (N4074, N4066);
buf BUF1 (N4075, N4069);
nand NAND3 (N4076, N4048, N1199, N3847);
buf BUF1 (N4077, N4065);
buf BUF1 (N4078, N4051);
nor NOR2 (N4079, N4076, N390);
not NOT1 (N4080, N4063);
not NOT1 (N4081, N4077);
xor XOR2 (N4082, N4071, N2917);
not NOT1 (N4083, N4082);
not NOT1 (N4084, N4073);
and AND4 (N4085, N4080, N419, N1683, N361);
not NOT1 (N4086, N4067);
and AND2 (N4087, N4084, N781);
not NOT1 (N4088, N4085);
nand NAND3 (N4089, N4087, N3371, N3664);
buf BUF1 (N4090, N4089);
or OR3 (N4091, N4081, N1103, N3929);
buf BUF1 (N4092, N4090);
not NOT1 (N4093, N4083);
or OR3 (N4094, N4093, N777, N1150);
buf BUF1 (N4095, N4058);
xor XOR2 (N4096, N4078, N2769);
or OR4 (N4097, N4079, N3120, N727, N499);
or OR3 (N4098, N4094, N1016, N544);
nand NAND4 (N4099, N4091, N2721, N1512, N2565);
or OR3 (N4100, N4098, N1630, N2339);
xor XOR2 (N4101, N4074, N235);
xor XOR2 (N4102, N4099, N2345);
not NOT1 (N4103, N4095);
nor NOR4 (N4104, N4100, N2240, N1855, N1970);
not NOT1 (N4105, N4075);
nand NAND3 (N4106, N4097, N1423, N3716);
buf BUF1 (N4107, N4105);
xor XOR2 (N4108, N4102, N1350);
buf BUF1 (N4109, N4086);
and AND3 (N4110, N4104, N1911, N3574);
xor XOR2 (N4111, N4109, N746);
buf BUF1 (N4112, N4092);
nor NOR4 (N4113, N4110, N3301, N3435, N3749);
xor XOR2 (N4114, N4113, N759);
or OR4 (N4115, N4111, N2485, N948, N3122);
nand NAND4 (N4116, N4101, N1493, N2234, N3217);
nand NAND4 (N4117, N4107, N2762, N549, N785);
not NOT1 (N4118, N4112);
nor NOR2 (N4119, N4106, N835);
and AND2 (N4120, N4117, N2309);
nor NOR3 (N4121, N4088, N4106, N2938);
nand NAND3 (N4122, N4119, N1747, N3825);
xor XOR2 (N4123, N4108, N3114);
nor NOR2 (N4124, N4122, N1871);
nor NOR2 (N4125, N4121, N2266);
xor XOR2 (N4126, N4114, N1844);
nor NOR4 (N4127, N4124, N2834, N558, N2801);
and AND3 (N4128, N4096, N1250, N730);
nand NAND3 (N4129, N4125, N3792, N1680);
nand NAND3 (N4130, N4127, N2740, N3704);
nand NAND3 (N4131, N4129, N1028, N2301);
or OR3 (N4132, N4115, N2752, N2553);
buf BUF1 (N4133, N4131);
nand NAND2 (N4134, N4123, N3279);
and AND4 (N4135, N4128, N2603, N4053, N407);
nand NAND4 (N4136, N4126, N1420, N2957, N2005);
not NOT1 (N4137, N4135);
buf BUF1 (N4138, N4130);
buf BUF1 (N4139, N4134);
not NOT1 (N4140, N4137);
not NOT1 (N4141, N4116);
not NOT1 (N4142, N4133);
and AND3 (N4143, N4140, N279, N1965);
xor XOR2 (N4144, N4141, N1218);
or OR3 (N4145, N4143, N3044, N3686);
and AND4 (N4146, N4142, N1989, N203, N3278);
and AND4 (N4147, N4103, N584, N1009, N960);
and AND2 (N4148, N4138, N414);
nand NAND3 (N4149, N4146, N3226, N959);
and AND2 (N4150, N4120, N1440);
xor XOR2 (N4151, N4150, N2969);
or OR3 (N4152, N4139, N4119, N609);
buf BUF1 (N4153, N4118);
nand NAND3 (N4154, N4132, N894, N916);
buf BUF1 (N4155, N4153);
buf BUF1 (N4156, N4149);
xor XOR2 (N4157, N4156, N3442);
not NOT1 (N4158, N4154);
xor XOR2 (N4159, N4152, N2328);
not NOT1 (N4160, N4148);
not NOT1 (N4161, N4157);
or OR3 (N4162, N4161, N2701, N3929);
buf BUF1 (N4163, N4151);
not NOT1 (N4164, N4158);
nor NOR2 (N4165, N4162, N2304);
nand NAND3 (N4166, N4145, N865, N889);
buf BUF1 (N4167, N4136);
and AND2 (N4168, N4164, N226);
and AND3 (N4169, N4165, N1805, N3257);
buf BUF1 (N4170, N4159);
nor NOR2 (N4171, N4163, N2466);
xor XOR2 (N4172, N4160, N2765);
nor NOR4 (N4173, N4167, N2810, N925, N1479);
nor NOR4 (N4174, N4171, N457, N2952, N2459);
and AND3 (N4175, N4173, N1089, N948);
and AND2 (N4176, N4168, N2443);
not NOT1 (N4177, N4155);
and AND2 (N4178, N4144, N3786);
and AND2 (N4179, N4177, N4078);
or OR2 (N4180, N4170, N2720);
or OR4 (N4181, N4172, N3834, N720, N37);
or OR2 (N4182, N4180, N3410);
xor XOR2 (N4183, N4169, N2878);
xor XOR2 (N4184, N4176, N3287);
buf BUF1 (N4185, N4166);
nand NAND4 (N4186, N4175, N919, N3611, N2643);
or OR4 (N4187, N4186, N612, N1223, N1395);
nor NOR3 (N4188, N4185, N3358, N2564);
nand NAND4 (N4189, N4182, N3796, N1981, N1095);
xor XOR2 (N4190, N4174, N608);
buf BUF1 (N4191, N4189);
buf BUF1 (N4192, N4191);
buf BUF1 (N4193, N4179);
buf BUF1 (N4194, N4187);
buf BUF1 (N4195, N4183);
nor NOR3 (N4196, N4188, N1257, N3652);
not NOT1 (N4197, N4193);
nor NOR3 (N4198, N4147, N856, N1411);
buf BUF1 (N4199, N4178);
xor XOR2 (N4200, N4194, N1377);
nor NOR2 (N4201, N4195, N3026);
xor XOR2 (N4202, N4199, N1949);
nor NOR2 (N4203, N4181, N1863);
buf BUF1 (N4204, N4196);
nor NOR4 (N4205, N4190, N279, N250, N374);
nor NOR4 (N4206, N4198, N3035, N1369, N2338);
and AND2 (N4207, N4205, N2353);
not NOT1 (N4208, N4201);
xor XOR2 (N4209, N4208, N2885);
xor XOR2 (N4210, N4202, N1973);
buf BUF1 (N4211, N4203);
xor XOR2 (N4212, N4210, N923);
buf BUF1 (N4213, N4197);
or OR2 (N4214, N4200, N380);
nor NOR2 (N4215, N4184, N731);
and AND4 (N4216, N4207, N783, N1705, N3630);
nand NAND3 (N4217, N4206, N1280, N1362);
or OR3 (N4218, N4214, N2026, N3248);
buf BUF1 (N4219, N4217);
buf BUF1 (N4220, N4192);
xor XOR2 (N4221, N4204, N4134);
or OR4 (N4222, N4220, N3672, N3308, N2888);
buf BUF1 (N4223, N4215);
nor NOR2 (N4224, N4212, N2039);
and AND3 (N4225, N4222, N3530, N1822);
not NOT1 (N4226, N4211);
xor XOR2 (N4227, N4226, N2322);
and AND3 (N4228, N4225, N1752, N1122);
buf BUF1 (N4229, N4224);
xor XOR2 (N4230, N4219, N1668);
nand NAND4 (N4231, N4227, N1986, N2331, N4164);
nor NOR4 (N4232, N4223, N3012, N800, N250);
not NOT1 (N4233, N4213);
buf BUF1 (N4234, N4228);
or OR3 (N4235, N4229, N1628, N727);
not NOT1 (N4236, N4221);
and AND4 (N4237, N4235, N380, N499, N2105);
not NOT1 (N4238, N4233);
nor NOR2 (N4239, N4236, N2444);
xor XOR2 (N4240, N4232, N3728);
xor XOR2 (N4241, N4240, N1795);
or OR4 (N4242, N4209, N3182, N2273, N1115);
and AND4 (N4243, N4218, N766, N761, N2590);
and AND3 (N4244, N4234, N660, N817);
xor XOR2 (N4245, N4242, N4084);
and AND2 (N4246, N4237, N3695);
buf BUF1 (N4247, N4230);
nand NAND2 (N4248, N4246, N1248);
nor NOR4 (N4249, N4241, N2056, N3442, N1870);
buf BUF1 (N4250, N4239);
and AND2 (N4251, N4243, N885);
nor NOR4 (N4252, N4249, N563, N1404, N1542);
buf BUF1 (N4253, N4247);
nand NAND3 (N4254, N4248, N2771, N1592);
and AND4 (N4255, N4250, N784, N2148, N3938);
xor XOR2 (N4256, N4238, N1545);
and AND3 (N4257, N4251, N2720, N997);
not NOT1 (N4258, N4255);
or OR2 (N4259, N4244, N3331);
or OR2 (N4260, N4252, N310);
and AND3 (N4261, N4254, N684, N2687);
buf BUF1 (N4262, N4260);
xor XOR2 (N4263, N4245, N1451);
xor XOR2 (N4264, N4262, N3602);
nand NAND4 (N4265, N4256, N990, N3000, N1405);
nand NAND2 (N4266, N4263, N1485);
buf BUF1 (N4267, N4265);
nand NAND4 (N4268, N4258, N2280, N57, N689);
not NOT1 (N4269, N4216);
and AND4 (N4270, N4253, N2015, N3186, N3796);
and AND4 (N4271, N4266, N3686, N1183, N3571);
buf BUF1 (N4272, N4271);
xor XOR2 (N4273, N4261, N407);
not NOT1 (N4274, N4270);
buf BUF1 (N4275, N4272);
nand NAND2 (N4276, N4264, N179);
buf BUF1 (N4277, N4273);
xor XOR2 (N4278, N4259, N939);
xor XOR2 (N4279, N4274, N4046);
xor XOR2 (N4280, N4257, N726);
nor NOR2 (N4281, N4267, N2455);
not NOT1 (N4282, N4279);
buf BUF1 (N4283, N4268);
nand NAND3 (N4284, N4277, N2547, N3333);
buf BUF1 (N4285, N4231);
or OR2 (N4286, N4283, N1434);
buf BUF1 (N4287, N4286);
buf BUF1 (N4288, N4275);
or OR3 (N4289, N4285, N2089, N2906);
not NOT1 (N4290, N4288);
or OR3 (N4291, N4280, N2202, N461);
xor XOR2 (N4292, N4291, N1072);
and AND2 (N4293, N4287, N3988);
not NOT1 (N4294, N4290);
nor NOR4 (N4295, N4278, N2970, N4212, N1836);
buf BUF1 (N4296, N4293);
nand NAND4 (N4297, N4281, N1987, N2376, N4065);
nand NAND3 (N4298, N4292, N3788, N2777);
not NOT1 (N4299, N4289);
and AND2 (N4300, N4297, N1271);
and AND2 (N4301, N4294, N876);
and AND3 (N4302, N4301, N2776, N1785);
nor NOR2 (N4303, N4298, N3185);
buf BUF1 (N4304, N4300);
xor XOR2 (N4305, N4299, N398);
nand NAND2 (N4306, N4276, N694);
buf BUF1 (N4307, N4282);
xor XOR2 (N4308, N4307, N1501);
buf BUF1 (N4309, N4306);
nor NOR2 (N4310, N4284, N3185);
nand NAND2 (N4311, N4296, N3126);
not NOT1 (N4312, N4269);
or OR4 (N4313, N4310, N2057, N3145, N965);
nor NOR3 (N4314, N4305, N149, N2526);
xor XOR2 (N4315, N4303, N1886);
buf BUF1 (N4316, N4309);
nand NAND4 (N4317, N4313, N372, N664, N3579);
and AND2 (N4318, N4312, N393);
and AND2 (N4319, N4302, N1155);
not NOT1 (N4320, N4317);
not NOT1 (N4321, N4316);
nor NOR4 (N4322, N4314, N3957, N388, N2015);
xor XOR2 (N4323, N4321, N2900);
and AND2 (N4324, N4320, N2506);
not NOT1 (N4325, N4323);
buf BUF1 (N4326, N4322);
and AND4 (N4327, N4311, N3665, N2474, N1955);
not NOT1 (N4328, N4308);
and AND3 (N4329, N4326, N250, N2363);
not NOT1 (N4330, N4319);
nor NOR4 (N4331, N4304, N3970, N2047, N3480);
nand NAND2 (N4332, N4324, N1302);
and AND4 (N4333, N4295, N3507, N4226, N3555);
or OR2 (N4334, N4325, N2626);
buf BUF1 (N4335, N4333);
xor XOR2 (N4336, N4332, N3049);
xor XOR2 (N4337, N4318, N2147);
nor NOR4 (N4338, N4330, N3800, N3800, N703);
or OR3 (N4339, N4328, N1246, N3165);
or OR3 (N4340, N4334, N2011, N694);
not NOT1 (N4341, N4335);
or OR2 (N4342, N4339, N2013);
nor NOR4 (N4343, N4331, N1117, N714, N2414);
or OR4 (N4344, N4315, N1766, N3328, N2126);
nand NAND4 (N4345, N4336, N226, N2407, N3137);
buf BUF1 (N4346, N4344);
nand NAND2 (N4347, N4341, N3648);
xor XOR2 (N4348, N4347, N4276);
xor XOR2 (N4349, N4340, N1643);
not NOT1 (N4350, N4346);
buf BUF1 (N4351, N4350);
buf BUF1 (N4352, N4337);
nor NOR3 (N4353, N4345, N3381, N1858);
xor XOR2 (N4354, N4349, N239);
xor XOR2 (N4355, N4338, N2583);
and AND2 (N4356, N4355, N2130);
nand NAND4 (N4357, N4348, N3076, N2970, N1498);
not NOT1 (N4358, N4352);
xor XOR2 (N4359, N4351, N1050);
buf BUF1 (N4360, N4353);
nor NOR3 (N4361, N4360, N564, N1605);
and AND3 (N4362, N4358, N1166, N940);
or OR4 (N4363, N4342, N3688, N2119, N4157);
xor XOR2 (N4364, N4343, N608);
or OR2 (N4365, N4357, N4217);
or OR4 (N4366, N4363, N423, N82, N1109);
xor XOR2 (N4367, N4356, N1604);
and AND4 (N4368, N4327, N3776, N1971, N3599);
or OR4 (N4369, N4329, N1622, N464, N3916);
buf BUF1 (N4370, N4362);
nor NOR3 (N4371, N4369, N2975, N2878);
nand NAND2 (N4372, N4367, N2133);
nand NAND3 (N4373, N4359, N2741, N3395);
or OR2 (N4374, N4368, N2285);
buf BUF1 (N4375, N4365);
and AND3 (N4376, N4364, N250, N1577);
and AND3 (N4377, N4374, N1739, N1252);
not NOT1 (N4378, N4370);
not NOT1 (N4379, N4378);
nor NOR3 (N4380, N4372, N2024, N933);
nand NAND3 (N4381, N4380, N3847, N3978);
buf BUF1 (N4382, N4381);
or OR2 (N4383, N4354, N407);
and AND4 (N4384, N4383, N274, N4268, N1885);
nor NOR3 (N4385, N4366, N2788, N3808);
or OR3 (N4386, N4384, N3469, N4157);
buf BUF1 (N4387, N4382);
not NOT1 (N4388, N4379);
nor NOR3 (N4389, N4375, N591, N775);
not NOT1 (N4390, N4376);
and AND4 (N4391, N4361, N1471, N343, N756);
buf BUF1 (N4392, N4389);
nand NAND3 (N4393, N4392, N1818, N2585);
or OR4 (N4394, N4371, N4112, N3284, N170);
not NOT1 (N4395, N4377);
or OR4 (N4396, N4387, N2959, N349, N3459);
buf BUF1 (N4397, N4394);
nor NOR4 (N4398, N4395, N1929, N180, N367);
and AND3 (N4399, N4391, N1002, N2398);
and AND4 (N4400, N4396, N979, N3463, N3261);
xor XOR2 (N4401, N4397, N60);
and AND2 (N4402, N4393, N4357);
not NOT1 (N4403, N4401);
nor NOR4 (N4404, N4399, N3572, N4108, N183);
nor NOR3 (N4405, N4385, N4041, N2957);
buf BUF1 (N4406, N4373);
not NOT1 (N4407, N4406);
buf BUF1 (N4408, N4390);
or OR2 (N4409, N4405, N3726);
or OR3 (N4410, N4403, N696, N4147);
or OR2 (N4411, N4408, N3347);
nand NAND4 (N4412, N4409, N4316, N1578, N828);
or OR3 (N4413, N4410, N3615, N1233);
and AND2 (N4414, N4402, N3739);
not NOT1 (N4415, N4388);
not NOT1 (N4416, N4411);
buf BUF1 (N4417, N4413);
not NOT1 (N4418, N4407);
buf BUF1 (N4419, N4417);
buf BUF1 (N4420, N4400);
or OR4 (N4421, N4412, N2851, N3275, N4189);
not NOT1 (N4422, N4386);
and AND4 (N4423, N4421, N4138, N1430, N2308);
xor XOR2 (N4424, N4404, N3828);
not NOT1 (N4425, N4416);
or OR3 (N4426, N4420, N1125, N227);
not NOT1 (N4427, N4398);
nand NAND2 (N4428, N4424, N3228);
or OR2 (N4429, N4414, N2252);
nor NOR4 (N4430, N4429, N1318, N188, N3205);
xor XOR2 (N4431, N4418, N3851);
and AND3 (N4432, N4430, N561, N2023);
nor NOR2 (N4433, N4428, N1384);
xor XOR2 (N4434, N4427, N758);
buf BUF1 (N4435, N4426);
nand NAND4 (N4436, N4433, N2750, N3766, N3075);
and AND2 (N4437, N4425, N791);
xor XOR2 (N4438, N4437, N1916);
buf BUF1 (N4439, N4435);
nor NOR4 (N4440, N4419, N819, N3445, N2258);
buf BUF1 (N4441, N4439);
and AND3 (N4442, N4415, N1740, N3701);
or OR3 (N4443, N4434, N1146, N3178);
nand NAND2 (N4444, N4442, N1708);
nor NOR2 (N4445, N4422, N1176);
not NOT1 (N4446, N4441);
and AND3 (N4447, N4443, N646, N575);
nor NOR2 (N4448, N4423, N602);
not NOT1 (N4449, N4444);
nand NAND2 (N4450, N4440, N3007);
nand NAND3 (N4451, N4448, N4343, N4011);
xor XOR2 (N4452, N4446, N2855);
and AND3 (N4453, N4447, N2095, N925);
xor XOR2 (N4454, N4449, N1525);
not NOT1 (N4455, N4431);
xor XOR2 (N4456, N4454, N2449);
xor XOR2 (N4457, N4455, N365);
nand NAND4 (N4458, N4450, N1714, N3196, N4428);
buf BUF1 (N4459, N4458);
not NOT1 (N4460, N4445);
or OR3 (N4461, N4438, N195, N1345);
nor NOR3 (N4462, N4456, N3062, N2570);
nor NOR2 (N4463, N4457, N1361);
buf BUF1 (N4464, N4452);
not NOT1 (N4465, N4462);
not NOT1 (N4466, N4465);
nor NOR2 (N4467, N4451, N1529);
nor NOR4 (N4468, N4464, N84, N161, N3019);
not NOT1 (N4469, N4453);
or OR4 (N4470, N4460, N8, N1485, N766);
xor XOR2 (N4471, N4467, N2036);
xor XOR2 (N4472, N4436, N2751);
xor XOR2 (N4473, N4470, N40);
and AND3 (N4474, N4459, N3805, N3152);
buf BUF1 (N4475, N4468);
xor XOR2 (N4476, N4461, N2732);
xor XOR2 (N4477, N4475, N763);
xor XOR2 (N4478, N4469, N467);
buf BUF1 (N4479, N4471);
nand NAND4 (N4480, N4476, N2403, N1433, N2161);
not NOT1 (N4481, N4463);
or OR3 (N4482, N4473, N2018, N4380);
nor NOR3 (N4483, N4480, N631, N1779);
buf BUF1 (N4484, N4477);
and AND3 (N4485, N4483, N2605, N1333);
nand NAND4 (N4486, N4478, N3884, N2543, N3145);
or OR4 (N4487, N4486, N655, N2341, N3505);
and AND3 (N4488, N4485, N3505, N1715);
and AND2 (N4489, N4482, N927);
buf BUF1 (N4490, N4432);
or OR4 (N4491, N4472, N3649, N695, N3491);
nand NAND3 (N4492, N4490, N1746, N4109);
or OR3 (N4493, N4487, N1886, N395);
not NOT1 (N4494, N4491);
or OR3 (N4495, N4466, N551, N2019);
not NOT1 (N4496, N4479);
or OR4 (N4497, N4493, N3806, N306, N4256);
xor XOR2 (N4498, N4489, N2887);
or OR3 (N4499, N4488, N122, N2130);
or OR3 (N4500, N4499, N3248, N389);
and AND4 (N4501, N4494, N116, N964, N3452);
not NOT1 (N4502, N4498);
not NOT1 (N4503, N4501);
xor XOR2 (N4504, N4481, N71);
and AND3 (N4505, N4503, N1333, N2587);
nand NAND3 (N4506, N4502, N1044, N2093);
xor XOR2 (N4507, N4497, N2517);
and AND2 (N4508, N4505, N1365);
nand NAND4 (N4509, N4500, N2914, N3336, N3776);
nand NAND3 (N4510, N4509, N3467, N3606);
xor XOR2 (N4511, N4506, N4303);
and AND4 (N4512, N4507, N471, N1776, N2684);
not NOT1 (N4513, N4511);
xor XOR2 (N4514, N4474, N1587);
xor XOR2 (N4515, N4504, N2499);
buf BUF1 (N4516, N4510);
not NOT1 (N4517, N4515);
buf BUF1 (N4518, N4516);
nand NAND3 (N4519, N4508, N3507, N1007);
nor NOR2 (N4520, N4492, N2300);
not NOT1 (N4521, N4517);
not NOT1 (N4522, N4521);
xor XOR2 (N4523, N4513, N2777);
buf BUF1 (N4524, N4519);
xor XOR2 (N4525, N4495, N557);
or OR4 (N4526, N4524, N742, N3801, N665);
nor NOR2 (N4527, N4523, N3634);
buf BUF1 (N4528, N4526);
xor XOR2 (N4529, N4512, N3929);
xor XOR2 (N4530, N4514, N3313);
not NOT1 (N4531, N4522);
or OR3 (N4532, N4528, N781, N702);
and AND4 (N4533, N4531, N1738, N4096, N3922);
not NOT1 (N4534, N4520);
and AND2 (N4535, N4496, N4044);
buf BUF1 (N4536, N4535);
not NOT1 (N4537, N4532);
nand NAND2 (N4538, N4536, N2760);
or OR3 (N4539, N4518, N3729, N4398);
buf BUF1 (N4540, N4537);
or OR3 (N4541, N4533, N3001, N3282);
xor XOR2 (N4542, N4530, N2779);
or OR2 (N4543, N4484, N4102);
not NOT1 (N4544, N4525);
buf BUF1 (N4545, N4542);
nand NAND4 (N4546, N4534, N3770, N4492, N3874);
buf BUF1 (N4547, N4540);
xor XOR2 (N4548, N4546, N514);
and AND4 (N4549, N4541, N608, N4444, N2655);
nor NOR3 (N4550, N4543, N2226, N1120);
or OR3 (N4551, N4550, N1918, N2733);
nand NAND3 (N4552, N4551, N379, N3470);
not NOT1 (N4553, N4539);
not NOT1 (N4554, N4538);
xor XOR2 (N4555, N4549, N836);
xor XOR2 (N4556, N4527, N2523);
buf BUF1 (N4557, N4552);
or OR3 (N4558, N4548, N260, N1431);
and AND4 (N4559, N4544, N2416, N3265, N3420);
buf BUF1 (N4560, N4555);
xor XOR2 (N4561, N4554, N3953);
nand NAND2 (N4562, N4556, N2101);
nor NOR4 (N4563, N4557, N2370, N3979, N552);
and AND2 (N4564, N4561, N2090);
and AND3 (N4565, N4563, N3642, N4048);
and AND2 (N4566, N4547, N359);
xor XOR2 (N4567, N4558, N2718);
xor XOR2 (N4568, N4553, N1236);
buf BUF1 (N4569, N4559);
nor NOR2 (N4570, N4567, N1290);
not NOT1 (N4571, N4568);
not NOT1 (N4572, N4565);
not NOT1 (N4573, N4545);
buf BUF1 (N4574, N4573);
xor XOR2 (N4575, N4562, N4356);
buf BUF1 (N4576, N4529);
nand NAND3 (N4577, N4576, N2946, N3944);
buf BUF1 (N4578, N4566);
nand NAND3 (N4579, N4560, N3104, N2919);
and AND3 (N4580, N4571, N1312, N2972);
nor NOR2 (N4581, N4579, N3688);
and AND4 (N4582, N4581, N359, N3833, N2040);
xor XOR2 (N4583, N4575, N4579);
or OR3 (N4584, N4574, N3248, N4014);
and AND2 (N4585, N4577, N3233);
or OR2 (N4586, N4585, N3874);
nand NAND2 (N4587, N4564, N4025);
or OR2 (N4588, N4583, N1495);
or OR2 (N4589, N4587, N2607);
not NOT1 (N4590, N4570);
nor NOR4 (N4591, N4582, N2622, N1483, N3105);
xor XOR2 (N4592, N4591, N4500);
buf BUF1 (N4593, N4580);
nand NAND4 (N4594, N4586, N795, N1860, N2634);
and AND4 (N4595, N4593, N1276, N204, N2498);
nand NAND4 (N4596, N4594, N1229, N2430, N4276);
or OR4 (N4597, N4572, N1594, N184, N2170);
xor XOR2 (N4598, N4584, N4091);
and AND2 (N4599, N4588, N385);
nor NOR3 (N4600, N4569, N269, N395);
nor NOR4 (N4601, N4578, N4364, N3957, N1850);
or OR3 (N4602, N4590, N4458, N1880);
and AND3 (N4603, N4596, N1698, N3949);
xor XOR2 (N4604, N4599, N320);
buf BUF1 (N4605, N4597);
buf BUF1 (N4606, N4598);
and AND2 (N4607, N4600, N703);
xor XOR2 (N4608, N4607, N3035);
not NOT1 (N4609, N4589);
and AND4 (N4610, N4609, N1659, N2361, N1605);
or OR2 (N4611, N4610, N3290);
xor XOR2 (N4612, N4611, N4054);
nor NOR2 (N4613, N4604, N2810);
nor NOR3 (N4614, N4606, N2418, N1770);
and AND4 (N4615, N4613, N1309, N3885, N2576);
not NOT1 (N4616, N4602);
nor NOR2 (N4617, N4595, N2742);
and AND2 (N4618, N4592, N3959);
or OR4 (N4619, N4617, N2043, N1380, N513);
and AND4 (N4620, N4608, N2368, N3048, N3061);
buf BUF1 (N4621, N4601);
or OR3 (N4622, N4618, N1956, N3894);
or OR2 (N4623, N4614, N3196);
nor NOR3 (N4624, N4605, N3199, N547);
nor NOR3 (N4625, N4603, N3623, N826);
nand NAND2 (N4626, N4612, N4564);
or OR3 (N4627, N4623, N3926, N2398);
xor XOR2 (N4628, N4620, N1574);
nand NAND3 (N4629, N4615, N3003, N4041);
buf BUF1 (N4630, N4629);
nor NOR3 (N4631, N4626, N1933, N1859);
not NOT1 (N4632, N4616);
nand NAND3 (N4633, N4619, N3758, N796);
nand NAND4 (N4634, N4630, N581, N2760, N4102);
not NOT1 (N4635, N4627);
or OR4 (N4636, N4635, N3370, N14, N2527);
and AND4 (N4637, N4625, N4368, N1562, N4602);
or OR4 (N4638, N4633, N2625, N447, N190);
buf BUF1 (N4639, N4622);
or OR3 (N4640, N4631, N274, N3297);
or OR4 (N4641, N4621, N1061, N4356, N552);
nand NAND4 (N4642, N4638, N3981, N4489, N4160);
nand NAND3 (N4643, N4637, N4391, N180);
buf BUF1 (N4644, N4641);
not NOT1 (N4645, N4628);
not NOT1 (N4646, N4640);
and AND2 (N4647, N4645, N403);
or OR4 (N4648, N4644, N3801, N1046, N4316);
buf BUF1 (N4649, N4646);
or OR4 (N4650, N4634, N3896, N339, N4238);
buf BUF1 (N4651, N4650);
nand NAND4 (N4652, N4632, N638, N1891, N2121);
not NOT1 (N4653, N4642);
buf BUF1 (N4654, N4643);
or OR4 (N4655, N4651, N4095, N4287, N2461);
nor NOR3 (N4656, N4654, N3207, N1391);
nor NOR4 (N4657, N4639, N1311, N1264, N4497);
nor NOR3 (N4658, N4624, N1021, N1047);
nor NOR3 (N4659, N4636, N3200, N4331);
buf BUF1 (N4660, N4649);
nor NOR3 (N4661, N4647, N3293, N2934);
not NOT1 (N4662, N4661);
nand NAND3 (N4663, N4655, N2323, N4084);
and AND3 (N4664, N4652, N3706, N242);
nor NOR4 (N4665, N4653, N3677, N176, N782);
or OR4 (N4666, N4664, N2490, N2190, N4157);
nor NOR4 (N4667, N4659, N448, N2879, N2527);
not NOT1 (N4668, N4663);
and AND3 (N4669, N4658, N2462, N722);
not NOT1 (N4670, N4667);
and AND3 (N4671, N4656, N1861, N2117);
nor NOR2 (N4672, N4648, N2200);
buf BUF1 (N4673, N4672);
and AND3 (N4674, N4657, N4368, N583);
nor NOR3 (N4675, N4674, N3973, N4348);
xor XOR2 (N4676, N4662, N2753);
nor NOR2 (N4677, N4671, N1570);
not NOT1 (N4678, N4665);
not NOT1 (N4679, N4675);
xor XOR2 (N4680, N4670, N1821);
nand NAND2 (N4681, N4668, N916);
and AND3 (N4682, N4679, N3946, N3887);
not NOT1 (N4683, N4660);
and AND4 (N4684, N4681, N2958, N4171, N1056);
buf BUF1 (N4685, N4678);
and AND3 (N4686, N4685, N3960, N788);
nand NAND2 (N4687, N4673, N2882);
buf BUF1 (N4688, N4684);
and AND4 (N4689, N4682, N4381, N4246, N3511);
and AND2 (N4690, N4689, N1976);
buf BUF1 (N4691, N4680);
not NOT1 (N4692, N4686);
nand NAND3 (N4693, N4687, N3287, N1519);
and AND4 (N4694, N4669, N1803, N4574, N530);
xor XOR2 (N4695, N4688, N2380);
nor NOR2 (N4696, N4677, N2711);
and AND4 (N4697, N4683, N2777, N3226, N2538);
or OR2 (N4698, N4697, N4420);
nor NOR4 (N4699, N4666, N2232, N3257, N955);
and AND3 (N4700, N4676, N2005, N2032);
buf BUF1 (N4701, N4699);
nand NAND3 (N4702, N4696, N3963, N2468);
buf BUF1 (N4703, N4698);
buf BUF1 (N4704, N4691);
xor XOR2 (N4705, N4694, N2301);
xor XOR2 (N4706, N4702, N4197);
xor XOR2 (N4707, N4690, N559);
nor NOR4 (N4708, N4706, N2989, N1084, N3059);
nor NOR4 (N4709, N4708, N541, N1963, N2604);
not NOT1 (N4710, N4703);
nor NOR4 (N4711, N4700, N3812, N1932, N4398);
xor XOR2 (N4712, N4701, N4458);
and AND3 (N4713, N4707, N1025, N4398);
or OR3 (N4714, N4709, N2767, N4692);
and AND2 (N4715, N2165, N4508);
and AND4 (N4716, N4695, N2303, N2459, N2224);
xor XOR2 (N4717, N4715, N2917);
nand NAND4 (N4718, N4704, N3149, N4436, N3761);
not NOT1 (N4719, N4711);
or OR4 (N4720, N4693, N3263, N3800, N3068);
nor NOR4 (N4721, N4713, N1490, N3759, N1919);
not NOT1 (N4722, N4705);
nand NAND3 (N4723, N4716, N2755, N1799);
buf BUF1 (N4724, N4719);
buf BUF1 (N4725, N4720);
xor XOR2 (N4726, N4724, N1351);
nand NAND3 (N4727, N4726, N3922, N247);
nand NAND2 (N4728, N4717, N3418);
xor XOR2 (N4729, N4714, N3568);
xor XOR2 (N4730, N4712, N1943);
nand NAND2 (N4731, N4721, N1414);
nor NOR4 (N4732, N4728, N4662, N1832, N3598);
nor NOR2 (N4733, N4723, N3456);
nor NOR3 (N4734, N4718, N4567, N4098);
nor NOR2 (N4735, N4722, N656);
or OR4 (N4736, N4734, N1430, N2648, N3910);
nor NOR4 (N4737, N4725, N4613, N4170, N1260);
xor XOR2 (N4738, N4710, N645);
not NOT1 (N4739, N4737);
and AND4 (N4740, N4730, N253, N2425, N4701);
or OR4 (N4741, N4733, N208, N3904, N3602);
and AND2 (N4742, N4732, N2770);
xor XOR2 (N4743, N4739, N904);
xor XOR2 (N4744, N4740, N2962);
nand NAND2 (N4745, N4741, N4264);
xor XOR2 (N4746, N4742, N3885);
nand NAND3 (N4747, N4738, N3288, N138);
nand NAND3 (N4748, N4745, N1470, N2241);
nand NAND4 (N4749, N4731, N2434, N3595, N3012);
nor NOR2 (N4750, N4735, N4155);
buf BUF1 (N4751, N4747);
not NOT1 (N4752, N4746);
xor XOR2 (N4753, N4748, N1941);
and AND4 (N4754, N4751, N1795, N613, N3861);
xor XOR2 (N4755, N4752, N45);
and AND4 (N4756, N4753, N219, N19, N3034);
buf BUF1 (N4757, N4736);
and AND3 (N4758, N4743, N3221, N3858);
and AND3 (N4759, N4750, N2907, N992);
or OR3 (N4760, N4727, N3091, N1742);
xor XOR2 (N4761, N4744, N1419);
nand NAND2 (N4762, N4754, N1575);
and AND4 (N4763, N4760, N3828, N1449, N1034);
nor NOR3 (N4764, N4759, N1937, N13);
and AND4 (N4765, N4758, N4540, N4432, N903);
and AND2 (N4766, N4756, N1584);
xor XOR2 (N4767, N4749, N3425);
not NOT1 (N4768, N4764);
buf BUF1 (N4769, N4766);
nor NOR3 (N4770, N4768, N3163, N2377);
not NOT1 (N4771, N4757);
or OR4 (N4772, N4769, N1505, N134, N1921);
xor XOR2 (N4773, N4761, N4555);
xor XOR2 (N4774, N4755, N3939);
and AND2 (N4775, N4773, N3333);
not NOT1 (N4776, N4770);
not NOT1 (N4777, N4763);
nor NOR4 (N4778, N4772, N2625, N2959, N4279);
not NOT1 (N4779, N4777);
not NOT1 (N4780, N4765);
buf BUF1 (N4781, N4780);
nand NAND3 (N4782, N4771, N1425, N4197);
nand NAND2 (N4783, N4776, N2384);
buf BUF1 (N4784, N4783);
nand NAND2 (N4785, N4782, N232);
nand NAND3 (N4786, N4774, N462, N4464);
and AND4 (N4787, N4767, N632, N3918, N1192);
nor NOR3 (N4788, N4785, N2582, N2266);
nand NAND2 (N4789, N4788, N2427);
nand NAND3 (N4790, N4787, N4329, N2401);
not NOT1 (N4791, N4781);
and AND4 (N4792, N4790, N127, N2088, N3267);
or OR3 (N4793, N4784, N3702, N4070);
nand NAND4 (N4794, N4791, N3867, N1655, N2196);
not NOT1 (N4795, N4793);
or OR3 (N4796, N4729, N3953, N3938);
nor NOR4 (N4797, N4795, N4334, N1268, N229);
and AND4 (N4798, N4779, N2924, N4712, N1156);
nand NAND4 (N4799, N4798, N4310, N2345, N3501);
nand NAND4 (N4800, N4778, N958, N3638, N3561);
xor XOR2 (N4801, N4786, N454);
nand NAND3 (N4802, N4796, N550, N3440);
nand NAND3 (N4803, N4789, N4506, N2322);
nor NOR4 (N4804, N4797, N2737, N3850, N1753);
or OR3 (N4805, N4803, N2342, N568);
and AND3 (N4806, N4804, N4528, N2863);
and AND4 (N4807, N4792, N4292, N2121, N2622);
or OR2 (N4808, N4794, N4234);
xor XOR2 (N4809, N4808, N1198);
and AND3 (N4810, N4809, N1254, N672);
xor XOR2 (N4811, N4810, N2307);
not NOT1 (N4812, N4799);
xor XOR2 (N4813, N4812, N4654);
or OR3 (N4814, N4807, N3130, N352);
xor XOR2 (N4815, N4805, N30);
and AND2 (N4816, N4801, N904);
nand NAND4 (N4817, N4814, N1230, N403, N4127);
or OR2 (N4818, N4775, N4009);
nor NOR4 (N4819, N4762, N3650, N1289, N110);
nand NAND3 (N4820, N4818, N3444, N2826);
or OR2 (N4821, N4813, N3954);
or OR3 (N4822, N4820, N1387, N3717);
nand NAND4 (N4823, N4816, N4799, N3342, N3118);
and AND3 (N4824, N4823, N136, N4349);
nand NAND2 (N4825, N4822, N1541);
and AND2 (N4826, N4806, N2714);
or OR3 (N4827, N4821, N2866, N3621);
not NOT1 (N4828, N4824);
nand NAND2 (N4829, N4826, N3271);
and AND2 (N4830, N4811, N442);
buf BUF1 (N4831, N4829);
or OR3 (N4832, N4802, N1568, N1636);
or OR4 (N4833, N4832, N764, N966, N4094);
not NOT1 (N4834, N4800);
xor XOR2 (N4835, N4834, N4585);
nand NAND4 (N4836, N4831, N4278, N3348, N2782);
nand NAND3 (N4837, N4817, N3544, N3122);
and AND3 (N4838, N4827, N556, N3844);
nand NAND3 (N4839, N4815, N2763, N4039);
nand NAND2 (N4840, N4819, N2131);
xor XOR2 (N4841, N4828, N3357);
buf BUF1 (N4842, N4835);
or OR4 (N4843, N4830, N3276, N74, N3693);
not NOT1 (N4844, N4837);
nand NAND3 (N4845, N4840, N1194, N3305);
xor XOR2 (N4846, N4844, N3827);
buf BUF1 (N4847, N4845);
and AND2 (N4848, N4825, N3771);
buf BUF1 (N4849, N4842);
xor XOR2 (N4850, N4848, N1094);
or OR3 (N4851, N4841, N356, N4113);
buf BUF1 (N4852, N4838);
buf BUF1 (N4853, N4851);
not NOT1 (N4854, N4846);
or OR2 (N4855, N4849, N3027);
xor XOR2 (N4856, N4836, N2486);
nand NAND4 (N4857, N4853, N2354, N1443, N3262);
not NOT1 (N4858, N4847);
or OR4 (N4859, N4843, N1305, N640, N4158);
not NOT1 (N4860, N4833);
and AND2 (N4861, N4854, N2105);
and AND2 (N4862, N4857, N4842);
nor NOR3 (N4863, N4860, N4375, N4460);
not NOT1 (N4864, N4850);
xor XOR2 (N4865, N4856, N1211);
and AND2 (N4866, N4852, N4322);
or OR4 (N4867, N4863, N730, N2546, N1785);
buf BUF1 (N4868, N4855);
nor NOR3 (N4869, N4858, N2766, N3422);
not NOT1 (N4870, N4865);
buf BUF1 (N4871, N4839);
nor NOR2 (N4872, N4870, N3495);
nand NAND4 (N4873, N4862, N3806, N3323, N2504);
nand NAND2 (N4874, N4869, N1894);
and AND3 (N4875, N4866, N4874, N1637);
nand NAND4 (N4876, N767, N1285, N942, N1669);
nor NOR4 (N4877, N4871, N2128, N3336, N4802);
nand NAND4 (N4878, N4861, N458, N4006, N4256);
buf BUF1 (N4879, N4873);
and AND4 (N4880, N4867, N2472, N2115, N2454);
not NOT1 (N4881, N4880);
buf BUF1 (N4882, N4868);
and AND4 (N4883, N4882, N2067, N2187, N1470);
xor XOR2 (N4884, N4859, N3730);
nor NOR4 (N4885, N4875, N635, N477, N4163);
not NOT1 (N4886, N4877);
xor XOR2 (N4887, N4881, N1121);
and AND2 (N4888, N4887, N3550);
or OR2 (N4889, N4872, N2167);
not NOT1 (N4890, N4888);
nor NOR2 (N4891, N4883, N3014);
buf BUF1 (N4892, N4889);
nand NAND2 (N4893, N4890, N4363);
or OR3 (N4894, N4864, N1736, N4326);
or OR3 (N4895, N4876, N3513, N4587);
nand NAND4 (N4896, N4895, N2411, N3563, N2654);
xor XOR2 (N4897, N4884, N3751);
xor XOR2 (N4898, N4891, N2002);
nor NOR4 (N4899, N4886, N1019, N4809, N1662);
or OR2 (N4900, N4878, N4301);
buf BUF1 (N4901, N4899);
nand NAND2 (N4902, N4897, N1747);
nand NAND3 (N4903, N4892, N509, N1996);
nor NOR4 (N4904, N4896, N98, N4785, N2787);
and AND2 (N4905, N4885, N3050);
and AND2 (N4906, N4903, N3511);
not NOT1 (N4907, N4906);
xor XOR2 (N4908, N4905, N565);
and AND4 (N4909, N4894, N4422, N2387, N1910);
not NOT1 (N4910, N4909);
nor NOR3 (N4911, N4902, N190, N3335);
nand NAND3 (N4912, N4893, N3616, N3958);
or OR3 (N4913, N4911, N4522, N3803);
nor NOR4 (N4914, N4901, N4862, N1253, N1222);
buf BUF1 (N4915, N4910);
and AND2 (N4916, N4908, N3225);
not NOT1 (N4917, N4913);
buf BUF1 (N4918, N4914);
nand NAND4 (N4919, N4918, N4914, N4628, N2906);
buf BUF1 (N4920, N4919);
nor NOR2 (N4921, N4879, N2612);
nor NOR2 (N4922, N4920, N4389);
nor NOR4 (N4923, N4907, N2047, N253, N2231);
or OR3 (N4924, N4900, N2986, N2793);
buf BUF1 (N4925, N4898);
and AND4 (N4926, N4915, N3803, N1634, N2602);
not NOT1 (N4927, N4923);
and AND4 (N4928, N4925, N657, N1242, N1334);
nand NAND4 (N4929, N4904, N1887, N3297, N3243);
buf BUF1 (N4930, N4927);
nor NOR3 (N4931, N4912, N161, N2491);
or OR3 (N4932, N4924, N2404, N3512);
or OR3 (N4933, N4931, N3762, N714);
nor NOR4 (N4934, N4922, N3647, N2805, N274);
and AND2 (N4935, N4928, N1025);
nor NOR2 (N4936, N4916, N4323);
or OR2 (N4937, N4934, N259);
xor XOR2 (N4938, N4929, N531);
and AND3 (N4939, N4933, N2370, N1204);
nor NOR3 (N4940, N4930, N1233, N1679);
xor XOR2 (N4941, N4926, N3427);
and AND3 (N4942, N4932, N387, N1780);
nor NOR4 (N4943, N4935, N365, N4755, N544);
nand NAND3 (N4944, N4940, N2524, N4452);
or OR4 (N4945, N4941, N4912, N1753, N116);
nand NAND2 (N4946, N4944, N4834);
nor NOR4 (N4947, N4942, N2834, N292, N2499);
xor XOR2 (N4948, N4946, N644);
or OR2 (N4949, N4943, N1807);
not NOT1 (N4950, N4938);
not NOT1 (N4951, N4945);
buf BUF1 (N4952, N4936);
or OR2 (N4953, N4948, N4852);
or OR3 (N4954, N4949, N1901, N3117);
and AND4 (N4955, N4951, N2263, N545, N3238);
buf BUF1 (N4956, N4921);
not NOT1 (N4957, N4956);
buf BUF1 (N4958, N4957);
nand NAND4 (N4959, N4958, N3458, N2392, N2421);
not NOT1 (N4960, N4954);
xor XOR2 (N4961, N4950, N2760);
nand NAND4 (N4962, N4959, N3323, N3867, N2471);
xor XOR2 (N4963, N4937, N2255);
not NOT1 (N4964, N4962);
nor NOR3 (N4965, N4963, N3834, N1340);
and AND4 (N4966, N4955, N167, N1238, N3485);
nand NAND4 (N4967, N4953, N3897, N2027, N1516);
xor XOR2 (N4968, N4939, N723);
or OR4 (N4969, N4960, N655, N4756, N2304);
nor NOR2 (N4970, N4968, N2673);
and AND2 (N4971, N4947, N2579);
nand NAND4 (N4972, N4966, N3659, N3184, N4012);
or OR2 (N4973, N4952, N1069);
not NOT1 (N4974, N4967);
xor XOR2 (N4975, N4917, N3041);
xor XOR2 (N4976, N4964, N526);
and AND2 (N4977, N4969, N130);
and AND2 (N4978, N4975, N3531);
and AND4 (N4979, N4971, N2113, N1003, N151);
and AND2 (N4980, N4970, N3983);
nor NOR3 (N4981, N4973, N2350, N596);
and AND3 (N4982, N4979, N1032, N4281);
xor XOR2 (N4983, N4961, N63);
not NOT1 (N4984, N4974);
and AND4 (N4985, N4978, N3187, N585, N3190);
and AND3 (N4986, N4984, N4276, N3004);
xor XOR2 (N4987, N4980, N583);
or OR2 (N4988, N4983, N4128);
or OR4 (N4989, N4977, N1439, N2685, N3103);
nand NAND3 (N4990, N4972, N3692, N1710);
not NOT1 (N4991, N4965);
nor NOR3 (N4992, N4982, N1058, N1865);
not NOT1 (N4993, N4985);
xor XOR2 (N4994, N4988, N123);
not NOT1 (N4995, N4989);
nand NAND3 (N4996, N4976, N3794, N254);
nor NOR3 (N4997, N4990, N6, N1696);
not NOT1 (N4998, N4986);
or OR2 (N4999, N4992, N2227);
and AND3 (N5000, N4993, N1276, N4646);
buf BUF1 (N5001, N4981);
nor NOR3 (N5002, N4998, N1947, N204);
buf BUF1 (N5003, N4994);
nor NOR2 (N5004, N4995, N1585);
or OR2 (N5005, N5000, N3929);
buf BUF1 (N5006, N5004);
nand NAND2 (N5007, N4987, N640);
buf BUF1 (N5008, N5003);
and AND2 (N5009, N5005, N3071);
and AND2 (N5010, N4997, N2556);
not NOT1 (N5011, N5006);
nor NOR3 (N5012, N4991, N39, N1464);
not NOT1 (N5013, N5007);
or OR4 (N5014, N5010, N1818, N2234, N4136);
buf BUF1 (N5015, N4996);
xor XOR2 (N5016, N4999, N2153);
and AND4 (N5017, N5001, N4343, N583, N2124);
nor NOR2 (N5018, N5011, N1149);
buf BUF1 (N5019, N5017);
and AND3 (N5020, N5008, N306, N4289);
nand NAND2 (N5021, N5014, N4825);
not NOT1 (N5022, N5021);
nor NOR2 (N5023, N5013, N90);
nand NAND4 (N5024, N5020, N4052, N270, N4259);
and AND4 (N5025, N5012, N2204, N1628, N3099);
nand NAND3 (N5026, N5016, N1952, N3718);
not NOT1 (N5027, N5018);
buf BUF1 (N5028, N5026);
not NOT1 (N5029, N5024);
buf BUF1 (N5030, N5025);
or OR3 (N5031, N5022, N3605, N3);
and AND2 (N5032, N5031, N4264);
or OR4 (N5033, N5029, N2663, N4229, N3118);
nand NAND2 (N5034, N5019, N1768);
xor XOR2 (N5035, N5033, N4758);
buf BUF1 (N5036, N5009);
not NOT1 (N5037, N5032);
buf BUF1 (N5038, N5036);
nand NAND3 (N5039, N5002, N1203, N4667);
nor NOR3 (N5040, N5035, N577, N3658);
nand NAND4 (N5041, N5030, N3782, N685, N3753);
nand NAND2 (N5042, N5037, N2935);
or OR4 (N5043, N5023, N3730, N2317, N2166);
and AND2 (N5044, N5027, N4867);
buf BUF1 (N5045, N5042);
nor NOR4 (N5046, N5041, N2349, N3250, N4514);
not NOT1 (N5047, N5040);
not NOT1 (N5048, N5038);
nand NAND2 (N5049, N5039, N4290);
nor NOR3 (N5050, N5015, N2424, N3334);
nand NAND2 (N5051, N5044, N4271);
xor XOR2 (N5052, N5043, N1114);
not NOT1 (N5053, N5049);
nand NAND4 (N5054, N5052, N25, N4689, N5014);
or OR3 (N5055, N5028, N2163, N2134);
xor XOR2 (N5056, N5045, N3188);
nand NAND3 (N5057, N5047, N330, N1807);
xor XOR2 (N5058, N5046, N2679);
nand NAND3 (N5059, N5056, N1645, N850);
not NOT1 (N5060, N5054);
nand NAND4 (N5061, N5050, N1335, N3298, N921);
and AND4 (N5062, N5051, N1887, N1418, N2831);
not NOT1 (N5063, N5057);
xor XOR2 (N5064, N5062, N379);
or OR2 (N5065, N5048, N2181);
nor NOR4 (N5066, N5055, N427, N4136, N2604);
buf BUF1 (N5067, N5053);
not NOT1 (N5068, N5061);
not NOT1 (N5069, N5058);
xor XOR2 (N5070, N5059, N2203);
xor XOR2 (N5071, N5060, N845);
nand NAND4 (N5072, N5034, N475, N2605, N527);
nand NAND4 (N5073, N5067, N1240, N1567, N3623);
and AND2 (N5074, N5065, N4294);
xor XOR2 (N5075, N5069, N3894);
and AND4 (N5076, N5064, N1422, N851, N869);
nor NOR3 (N5077, N5075, N2216, N4189);
not NOT1 (N5078, N5073);
xor XOR2 (N5079, N5063, N3986);
or OR2 (N5080, N5079, N3159);
not NOT1 (N5081, N5070);
or OR3 (N5082, N5071, N2552, N2831);
nor NOR2 (N5083, N5078, N2054);
nand NAND2 (N5084, N5068, N1533);
nor NOR2 (N5085, N5076, N2096);
not NOT1 (N5086, N5074);
or OR2 (N5087, N5072, N2648);
not NOT1 (N5088, N5081);
nand NAND4 (N5089, N5087, N2239, N2236, N1844);
buf BUF1 (N5090, N5077);
and AND2 (N5091, N5089, N1167);
or OR2 (N5092, N5082, N3122);
and AND4 (N5093, N5066, N3733, N3808, N4930);
and AND4 (N5094, N5088, N2982, N4302, N897);
buf BUF1 (N5095, N5093);
buf BUF1 (N5096, N5085);
nand NAND2 (N5097, N5091, N1533);
or OR3 (N5098, N5083, N847, N1804);
xor XOR2 (N5099, N5092, N2734);
xor XOR2 (N5100, N5096, N177);
buf BUF1 (N5101, N5100);
xor XOR2 (N5102, N5084, N1734);
and AND3 (N5103, N5097, N3476, N3707);
buf BUF1 (N5104, N5080);
nor NOR3 (N5105, N5101, N2795, N4004);
or OR3 (N5106, N5099, N4891, N3183);
or OR3 (N5107, N5104, N4918, N943);
not NOT1 (N5108, N5106);
xor XOR2 (N5109, N5095, N1989);
buf BUF1 (N5110, N5109);
not NOT1 (N5111, N5102);
or OR2 (N5112, N5110, N1039);
nor NOR4 (N5113, N5086, N1429, N3336, N3918);
xor XOR2 (N5114, N5105, N3217);
buf BUF1 (N5115, N5090);
nand NAND2 (N5116, N5115, N3195);
not NOT1 (N5117, N5113);
buf BUF1 (N5118, N5098);
nor NOR4 (N5119, N5108, N926, N4920, N541);
nand NAND4 (N5120, N5103, N1977, N2857, N4071);
buf BUF1 (N5121, N5111);
and AND4 (N5122, N5120, N4287, N4748, N2418);
xor XOR2 (N5123, N5094, N705);
and AND3 (N5124, N5107, N3293, N14);
not NOT1 (N5125, N5121);
or OR4 (N5126, N5122, N2411, N4827, N3810);
xor XOR2 (N5127, N5123, N1658);
not NOT1 (N5128, N5116);
xor XOR2 (N5129, N5127, N4841);
nor NOR2 (N5130, N5126, N1313);
nand NAND3 (N5131, N5117, N4205, N4850);
nand NAND2 (N5132, N5114, N4037);
buf BUF1 (N5133, N5129);
nor NOR2 (N5134, N5132, N3386);
buf BUF1 (N5135, N5112);
and AND2 (N5136, N5133, N4654);
xor XOR2 (N5137, N5119, N1033);
buf BUF1 (N5138, N5134);
not NOT1 (N5139, N5137);
nor NOR3 (N5140, N5124, N2851, N350);
xor XOR2 (N5141, N5131, N1210);
xor XOR2 (N5142, N5140, N51);
not NOT1 (N5143, N5128);
and AND4 (N5144, N5136, N4893, N4427, N3433);
not NOT1 (N5145, N5142);
buf BUF1 (N5146, N5118);
xor XOR2 (N5147, N5145, N3490);
not NOT1 (N5148, N5125);
buf BUF1 (N5149, N5147);
nor NOR3 (N5150, N5138, N1089, N126);
xor XOR2 (N5151, N5148, N253);
buf BUF1 (N5152, N5149);
nor NOR2 (N5153, N5135, N2034);
nand NAND4 (N5154, N5153, N4962, N3637, N1099);
nor NOR2 (N5155, N5143, N3353);
not NOT1 (N5156, N5155);
or OR4 (N5157, N5130, N4760, N3178, N3028);
and AND3 (N5158, N5150, N1911, N4038);
nand NAND2 (N5159, N5144, N940);
nand NAND3 (N5160, N5146, N453, N2009);
buf BUF1 (N5161, N5156);
xor XOR2 (N5162, N5161, N2750);
nand NAND4 (N5163, N5160, N326, N1096, N209);
nor NOR3 (N5164, N5139, N1354, N4653);
buf BUF1 (N5165, N5164);
buf BUF1 (N5166, N5162);
buf BUF1 (N5167, N5151);
or OR4 (N5168, N5166, N4481, N1896, N3810);
nor NOR3 (N5169, N5168, N3377, N3497);
not NOT1 (N5170, N5158);
nand NAND2 (N5171, N5141, N1081);
xor XOR2 (N5172, N5163, N3414);
buf BUF1 (N5173, N5157);
nor NOR3 (N5174, N5167, N516, N122);
xor XOR2 (N5175, N5165, N3797);
buf BUF1 (N5176, N5171);
and AND3 (N5177, N5174, N2629, N1717);
and AND3 (N5178, N5170, N3127, N16);
or OR2 (N5179, N5178, N3228);
nand NAND4 (N5180, N5159, N3525, N497, N5143);
nand NAND4 (N5181, N5152, N3433, N2817, N4103);
buf BUF1 (N5182, N5169);
or OR3 (N5183, N5182, N677, N588);
xor XOR2 (N5184, N5180, N197);
nand NAND3 (N5185, N5172, N3558, N3777);
nor NOR2 (N5186, N5175, N3868);
or OR4 (N5187, N5177, N4533, N4122, N3242);
nor NOR4 (N5188, N5173, N2210, N1184, N4495);
xor XOR2 (N5189, N5154, N3646);
not NOT1 (N5190, N5189);
nand NAND3 (N5191, N5184, N2254, N3191);
nor NOR3 (N5192, N5188, N2402, N677);
not NOT1 (N5193, N5185);
and AND3 (N5194, N5187, N4235, N852);
buf BUF1 (N5195, N5176);
and AND2 (N5196, N5186, N1198);
nor NOR4 (N5197, N5192, N4946, N385, N975);
nor NOR4 (N5198, N5196, N2040, N306, N1259);
or OR4 (N5199, N5195, N4477, N4866, N4279);
nor NOR2 (N5200, N5181, N2204);
buf BUF1 (N5201, N5200);
nand NAND4 (N5202, N5194, N442, N736, N4963);
or OR4 (N5203, N5191, N3882, N883, N4826);
nor NOR3 (N5204, N5190, N3181, N4586);
nor NOR2 (N5205, N5203, N3704);
xor XOR2 (N5206, N5205, N3633);
or OR4 (N5207, N5201, N415, N170, N4422);
not NOT1 (N5208, N5197);
xor XOR2 (N5209, N5199, N5000);
nand NAND2 (N5210, N5202, N793);
buf BUF1 (N5211, N5204);
buf BUF1 (N5212, N5208);
xor XOR2 (N5213, N5206, N211);
buf BUF1 (N5214, N5193);
nor NOR2 (N5215, N5213, N2397);
nor NOR2 (N5216, N5210, N509);
nand NAND2 (N5217, N5212, N3241);
not NOT1 (N5218, N5215);
nor NOR2 (N5219, N5211, N3520);
and AND4 (N5220, N5217, N2248, N4851, N484);
not NOT1 (N5221, N5179);
nor NOR2 (N5222, N5207, N941);
xor XOR2 (N5223, N5218, N2288);
nand NAND4 (N5224, N5183, N1715, N4183, N2918);
nor NOR3 (N5225, N5220, N4788, N3054);
xor XOR2 (N5226, N5216, N2221);
not NOT1 (N5227, N5223);
nand NAND2 (N5228, N5226, N3356);
buf BUF1 (N5229, N5224);
nand NAND4 (N5230, N5227, N559, N3377, N377);
xor XOR2 (N5231, N5219, N1700);
nor NOR4 (N5232, N5222, N645, N1697, N1101);
nand NAND3 (N5233, N5232, N1199, N3594);
nand NAND3 (N5234, N5198, N2109, N2191);
and AND4 (N5235, N5225, N4327, N5035, N2648);
xor XOR2 (N5236, N5228, N3786);
not NOT1 (N5237, N5214);
xor XOR2 (N5238, N5235, N2492);
nor NOR2 (N5239, N5234, N389);
and AND3 (N5240, N5233, N1569, N3161);
and AND2 (N5241, N5229, N4066);
and AND4 (N5242, N5231, N3467, N2153, N4663);
or OR4 (N5243, N5236, N1066, N1633, N2501);
nand NAND4 (N5244, N5240, N206, N508, N1329);
or OR3 (N5245, N5238, N1935, N3895);
nand NAND2 (N5246, N5242, N700);
nand NAND2 (N5247, N5237, N5229);
and AND2 (N5248, N5241, N2073);
not NOT1 (N5249, N5247);
nor NOR2 (N5250, N5244, N2256);
not NOT1 (N5251, N5246);
and AND2 (N5252, N5249, N3395);
buf BUF1 (N5253, N5248);
xor XOR2 (N5254, N5230, N2296);
nand NAND4 (N5255, N5250, N3908, N4976, N5043);
buf BUF1 (N5256, N5239);
nor NOR2 (N5257, N5245, N230);
xor XOR2 (N5258, N5221, N232);
nor NOR2 (N5259, N5255, N2134);
or OR2 (N5260, N5254, N2006);
and AND3 (N5261, N5256, N3081, N3074);
and AND4 (N5262, N5259, N3245, N4681, N1614);
and AND4 (N5263, N5261, N4570, N1893, N49);
not NOT1 (N5264, N5263);
nand NAND4 (N5265, N5260, N3920, N3831, N802);
not NOT1 (N5266, N5264);
nand NAND3 (N5267, N5253, N2655, N5151);
and AND3 (N5268, N5266, N3137, N1214);
or OR2 (N5269, N5268, N558);
or OR3 (N5270, N5257, N110, N1981);
nor NOR3 (N5271, N5267, N3966, N4820);
xor XOR2 (N5272, N5251, N1931);
buf BUF1 (N5273, N5258);
not NOT1 (N5274, N5262);
xor XOR2 (N5275, N5273, N905);
or OR3 (N5276, N5274, N4515, N208);
nor NOR2 (N5277, N5271, N3398);
or OR4 (N5278, N5209, N5020, N3074, N3636);
nand NAND3 (N5279, N5243, N3092, N4476);
or OR2 (N5280, N5277, N1792);
buf BUF1 (N5281, N5272);
or OR3 (N5282, N5275, N4547, N3469);
nor NOR2 (N5283, N5280, N3424);
and AND4 (N5284, N5282, N4398, N1517, N5255);
not NOT1 (N5285, N5283);
not NOT1 (N5286, N5252);
buf BUF1 (N5287, N5286);
nand NAND2 (N5288, N5278, N2469);
xor XOR2 (N5289, N5287, N4492);
nand NAND4 (N5290, N5270, N5177, N4982, N3241);
nand NAND3 (N5291, N5265, N2739, N1623);
or OR3 (N5292, N5285, N4183, N1444);
xor XOR2 (N5293, N5281, N4778);
nor NOR3 (N5294, N5288, N3647, N4763);
nor NOR2 (N5295, N5291, N670);
not NOT1 (N5296, N5276);
or OR2 (N5297, N5293, N2067);
buf BUF1 (N5298, N5294);
nor NOR2 (N5299, N5279, N1240);
nand NAND4 (N5300, N5289, N2456, N4102, N4100);
or OR4 (N5301, N5297, N4536, N1103, N4868);
buf BUF1 (N5302, N5300);
or OR3 (N5303, N5284, N4653, N810);
xor XOR2 (N5304, N5302, N3492);
nor NOR2 (N5305, N5304, N3373);
xor XOR2 (N5306, N5295, N3128);
not NOT1 (N5307, N5306);
or OR4 (N5308, N5298, N4523, N2420, N769);
nand NAND4 (N5309, N5305, N1275, N4476, N3039);
buf BUF1 (N5310, N5301);
or OR4 (N5311, N5290, N4400, N346, N3889);
buf BUF1 (N5312, N5311);
not NOT1 (N5313, N5269);
xor XOR2 (N5314, N5307, N3958);
not NOT1 (N5315, N5308);
not NOT1 (N5316, N5310);
nand NAND2 (N5317, N5316, N4324);
xor XOR2 (N5318, N5315, N2907);
not NOT1 (N5319, N5303);
nand NAND4 (N5320, N5319, N3461, N1460, N4861);
nor NOR4 (N5321, N5312, N2129, N1748, N69);
not NOT1 (N5322, N5321);
nand NAND4 (N5323, N5299, N4672, N2265, N548);
not NOT1 (N5324, N5317);
nor NOR4 (N5325, N5296, N2933, N2575, N1660);
xor XOR2 (N5326, N5323, N4669);
nor NOR2 (N5327, N5324, N3092);
nand NAND2 (N5328, N5325, N4139);
and AND3 (N5329, N5313, N324, N4173);
not NOT1 (N5330, N5322);
nor NOR2 (N5331, N5309, N4662);
not NOT1 (N5332, N5314);
nor NOR4 (N5333, N5326, N386, N1733, N2200);
buf BUF1 (N5334, N5292);
not NOT1 (N5335, N5327);
buf BUF1 (N5336, N5330);
or OR2 (N5337, N5335, N314);
and AND2 (N5338, N5333, N1420);
nand NAND2 (N5339, N5320, N3579);
and AND4 (N5340, N5331, N4422, N600, N916);
nor NOR4 (N5341, N5340, N1216, N1222, N5001);
nor NOR2 (N5342, N5339, N2370);
xor XOR2 (N5343, N5329, N172);
not NOT1 (N5344, N5332);
and AND4 (N5345, N5336, N1827, N1583, N4417);
or OR2 (N5346, N5343, N2752);
not NOT1 (N5347, N5337);
not NOT1 (N5348, N5347);
not NOT1 (N5349, N5341);
or OR4 (N5350, N5338, N1484, N325, N4833);
nor NOR3 (N5351, N5334, N3366, N1039);
not NOT1 (N5352, N5344);
xor XOR2 (N5353, N5342, N3733);
buf BUF1 (N5354, N5349);
not NOT1 (N5355, N5345);
and AND2 (N5356, N5351, N1791);
or OR4 (N5357, N5318, N3212, N2334, N1531);
or OR4 (N5358, N5348, N694, N4163, N3644);
xor XOR2 (N5359, N5357, N4182);
nand NAND2 (N5360, N5353, N3412);
or OR2 (N5361, N5360, N3881);
buf BUF1 (N5362, N5328);
not NOT1 (N5363, N5352);
not NOT1 (N5364, N5359);
buf BUF1 (N5365, N5355);
xor XOR2 (N5366, N5346, N439);
nor NOR2 (N5367, N5350, N765);
xor XOR2 (N5368, N5366, N1288);
xor XOR2 (N5369, N5368, N930);
nor NOR3 (N5370, N5361, N3192, N4314);
nand NAND4 (N5371, N5370, N4221, N1467, N2600);
nor NOR2 (N5372, N5363, N4350);
nor NOR3 (N5373, N5354, N4775, N4703);
not NOT1 (N5374, N5362);
nand NAND2 (N5375, N5372, N2966);
not NOT1 (N5376, N5373);
buf BUF1 (N5377, N5365);
buf BUF1 (N5378, N5358);
not NOT1 (N5379, N5369);
not NOT1 (N5380, N5367);
nand NAND2 (N5381, N5371, N4361);
xor XOR2 (N5382, N5356, N891);
buf BUF1 (N5383, N5381);
nor NOR2 (N5384, N5377, N2586);
nor NOR2 (N5385, N5378, N1314);
or OR4 (N5386, N5382, N2790, N4728, N2674);
xor XOR2 (N5387, N5364, N2672);
and AND3 (N5388, N5374, N1675, N141);
or OR2 (N5389, N5383, N5284);
nand NAND3 (N5390, N5385, N2131, N758);
xor XOR2 (N5391, N5384, N649);
nor NOR4 (N5392, N5387, N622, N3712, N3650);
nor NOR3 (N5393, N5390, N2334, N4203);
nand NAND4 (N5394, N5375, N3045, N1119, N1726);
not NOT1 (N5395, N5388);
nand NAND3 (N5396, N5386, N986, N559);
or OR4 (N5397, N5396, N1611, N5244, N1631);
nor NOR2 (N5398, N5392, N1037);
nand NAND4 (N5399, N5394, N2064, N5208, N213);
xor XOR2 (N5400, N5393, N3601);
or OR4 (N5401, N5389, N3348, N2176, N1606);
or OR2 (N5402, N5399, N3350);
buf BUF1 (N5403, N5395);
buf BUF1 (N5404, N5397);
xor XOR2 (N5405, N5398, N1242);
nor NOR3 (N5406, N5405, N2512, N3705);
nand NAND2 (N5407, N5379, N3652);
not NOT1 (N5408, N5404);
or OR4 (N5409, N5380, N2244, N5154, N5202);
nand NAND2 (N5410, N5408, N2406);
nor NOR4 (N5411, N5402, N3442, N1042, N2742);
buf BUF1 (N5412, N5411);
or OR4 (N5413, N5391, N4599, N4194, N1212);
buf BUF1 (N5414, N5413);
xor XOR2 (N5415, N5403, N342);
nand NAND2 (N5416, N5415, N633);
nor NOR2 (N5417, N5400, N2515);
buf BUF1 (N5418, N5410);
not NOT1 (N5419, N5407);
not NOT1 (N5420, N5412);
or OR4 (N5421, N5376, N2204, N2613, N926);
nor NOR3 (N5422, N5419, N1018, N1187);
and AND3 (N5423, N5416, N1723, N1537);
nand NAND3 (N5424, N5414, N3242, N4535);
not NOT1 (N5425, N5423);
xor XOR2 (N5426, N5421, N4883);
buf BUF1 (N5427, N5406);
or OR4 (N5428, N5418, N287, N3839, N383);
nor NOR4 (N5429, N5426, N4734, N5333, N730);
buf BUF1 (N5430, N5424);
nand NAND3 (N5431, N5417, N823, N4754);
xor XOR2 (N5432, N5420, N3600);
buf BUF1 (N5433, N5409);
nor NOR2 (N5434, N5428, N2063);
not NOT1 (N5435, N5434);
buf BUF1 (N5436, N5433);
not NOT1 (N5437, N5401);
and AND4 (N5438, N5437, N1068, N894, N1719);
not NOT1 (N5439, N5436);
xor XOR2 (N5440, N5422, N1632);
nand NAND2 (N5441, N5438, N196);
buf BUF1 (N5442, N5441);
not NOT1 (N5443, N5439);
nand NAND3 (N5444, N5430, N1499, N323);
nand NAND4 (N5445, N5432, N2385, N5281, N2950);
nor NOR2 (N5446, N5442, N3411);
and AND3 (N5447, N5425, N108, N2274);
nand NAND2 (N5448, N5446, N4940);
buf BUF1 (N5449, N5444);
xor XOR2 (N5450, N5427, N1630);
buf BUF1 (N5451, N5450);
buf BUF1 (N5452, N5435);
and AND3 (N5453, N5440, N3215, N3028);
and AND2 (N5454, N5452, N5224);
nor NOR3 (N5455, N5454, N3106, N2707);
not NOT1 (N5456, N5429);
nand NAND3 (N5457, N5447, N246, N4085);
nand NAND2 (N5458, N5431, N3150);
nor NOR2 (N5459, N5449, N2175);
buf BUF1 (N5460, N5451);
or OR3 (N5461, N5453, N1128, N2469);
and AND3 (N5462, N5460, N1704, N4456);
not NOT1 (N5463, N5458);
xor XOR2 (N5464, N5445, N431);
xor XOR2 (N5465, N5459, N2563);
buf BUF1 (N5466, N5457);
nand NAND3 (N5467, N5455, N4754, N161);
nand NAND2 (N5468, N5465, N3743);
nand NAND4 (N5469, N5467, N3876, N5462, N2063);
xor XOR2 (N5470, N693, N2227);
or OR3 (N5471, N5463, N1510, N1195);
nand NAND3 (N5472, N5468, N3773, N798);
nor NOR3 (N5473, N5448, N2704, N1076);
nand NAND4 (N5474, N5461, N5231, N5034, N1309);
and AND4 (N5475, N5471, N3008, N1434, N3261);
nor NOR3 (N5476, N5473, N1649, N4629);
not NOT1 (N5477, N5474);
not NOT1 (N5478, N5443);
and AND4 (N5479, N5476, N4072, N5228, N4141);
nand NAND2 (N5480, N5475, N1031);
buf BUF1 (N5481, N5477);
nor NOR4 (N5482, N5470, N3234, N3643, N3349);
or OR3 (N5483, N5469, N4173, N1610);
buf BUF1 (N5484, N5482);
buf BUF1 (N5485, N5481);
buf BUF1 (N5486, N5485);
or OR2 (N5487, N5472, N5335);
nand NAND3 (N5488, N5487, N682, N3090);
xor XOR2 (N5489, N5479, N527);
nor NOR3 (N5490, N5486, N2158, N4231);
nor NOR2 (N5491, N5464, N2057);
nor NOR3 (N5492, N5478, N4324, N2290);
or OR4 (N5493, N5488, N1363, N4058, N3980);
and AND2 (N5494, N5489, N1438);
nand NAND2 (N5495, N5494, N4466);
nand NAND3 (N5496, N5490, N3364, N4981);
nand NAND4 (N5497, N5492, N5027, N4125, N3704);
nand NAND4 (N5498, N5456, N1612, N2755, N1911);
not NOT1 (N5499, N5484);
xor XOR2 (N5500, N5491, N3877);
not NOT1 (N5501, N5493);
not NOT1 (N5502, N5480);
or OR2 (N5503, N5499, N3933);
nand NAND4 (N5504, N5501, N4641, N2496, N1438);
nor NOR3 (N5505, N5496, N3122, N3732);
not NOT1 (N5506, N5504);
nor NOR3 (N5507, N5497, N1341, N3403);
not NOT1 (N5508, N5503);
nor NOR2 (N5509, N5505, N1773);
buf BUF1 (N5510, N5508);
not NOT1 (N5511, N5495);
nor NOR3 (N5512, N5498, N2901, N86);
nand NAND2 (N5513, N5512, N2226);
or OR3 (N5514, N5507, N191, N3849);
nor NOR2 (N5515, N5510, N4227);
or OR3 (N5516, N5502, N3015, N3191);
xor XOR2 (N5517, N5511, N3253);
and AND2 (N5518, N5515, N177);
xor XOR2 (N5519, N5513, N4500);
nor NOR3 (N5520, N5466, N1212, N1367);
not NOT1 (N5521, N5483);
xor XOR2 (N5522, N5518, N691);
xor XOR2 (N5523, N5517, N5495);
not NOT1 (N5524, N5520);
nor NOR3 (N5525, N5524, N4253, N4327);
buf BUF1 (N5526, N5523);
xor XOR2 (N5527, N5521, N13);
and AND4 (N5528, N5500, N268, N4206, N1999);
nor NOR2 (N5529, N5514, N134);
or OR3 (N5530, N5527, N5341, N3144);
and AND2 (N5531, N5509, N188);
or OR3 (N5532, N5528, N3618, N2532);
xor XOR2 (N5533, N5530, N2784);
or OR4 (N5534, N5532, N3539, N5151, N2990);
buf BUF1 (N5535, N5533);
not NOT1 (N5536, N5525);
and AND4 (N5537, N5536, N223, N4816, N3584);
buf BUF1 (N5538, N5519);
and AND2 (N5539, N5531, N209);
and AND4 (N5540, N5526, N1209, N772, N2482);
xor XOR2 (N5541, N5535, N4398);
nor NOR4 (N5542, N5522, N3966, N5427, N2818);
nand NAND4 (N5543, N5541, N1735, N299, N916);
nand NAND2 (N5544, N5537, N5428);
not NOT1 (N5545, N5544);
xor XOR2 (N5546, N5539, N1598);
not NOT1 (N5547, N5534);
buf BUF1 (N5548, N5506);
nor NOR4 (N5549, N5543, N5226, N3962, N3046);
and AND3 (N5550, N5542, N1299, N1280);
not NOT1 (N5551, N5545);
not NOT1 (N5552, N5540);
buf BUF1 (N5553, N5548);
xor XOR2 (N5554, N5516, N458);
nor NOR3 (N5555, N5551, N1167, N1269);
xor XOR2 (N5556, N5529, N738);
buf BUF1 (N5557, N5555);
or OR3 (N5558, N5547, N450, N2740);
xor XOR2 (N5559, N5552, N3971);
xor XOR2 (N5560, N5557, N5328);
buf BUF1 (N5561, N5554);
nor NOR2 (N5562, N5538, N1943);
and AND4 (N5563, N5558, N2807, N1696, N2690);
nor NOR2 (N5564, N5559, N5342);
buf BUF1 (N5565, N5562);
nor NOR2 (N5566, N5560, N453);
nor NOR4 (N5567, N5550, N2237, N2997, N1533);
nor NOR2 (N5568, N5556, N652);
and AND4 (N5569, N5568, N1335, N4683, N5427);
nor NOR2 (N5570, N5553, N2082);
and AND3 (N5571, N5565, N840, N1003);
xor XOR2 (N5572, N5566, N1812);
buf BUF1 (N5573, N5569);
not NOT1 (N5574, N5573);
and AND4 (N5575, N5549, N4441, N4967, N4977);
nand NAND3 (N5576, N5563, N1115, N947);
and AND3 (N5577, N5571, N1597, N2192);
nor NOR3 (N5578, N5561, N4179, N4284);
not NOT1 (N5579, N5572);
or OR3 (N5580, N5546, N5556, N3654);
or OR4 (N5581, N5579, N3787, N5175, N1586);
not NOT1 (N5582, N5567);
and AND2 (N5583, N5570, N3024);
nor NOR2 (N5584, N5582, N1935);
or OR3 (N5585, N5564, N1475, N1919);
nand NAND3 (N5586, N5575, N2060, N942);
buf BUF1 (N5587, N5577);
buf BUF1 (N5588, N5581);
not NOT1 (N5589, N5585);
buf BUF1 (N5590, N5574);
and AND4 (N5591, N5580, N4421, N30, N4190);
or OR3 (N5592, N5586, N4982, N1102);
xor XOR2 (N5593, N5590, N2171);
xor XOR2 (N5594, N5593, N3414);
nand NAND2 (N5595, N5587, N396);
or OR3 (N5596, N5591, N3468, N1090);
or OR4 (N5597, N5595, N2897, N2254, N2190);
xor XOR2 (N5598, N5588, N1923);
buf BUF1 (N5599, N5583);
nand NAND2 (N5600, N5578, N5278);
or OR4 (N5601, N5594, N3297, N3161, N2897);
nand NAND2 (N5602, N5584, N1836);
nand NAND3 (N5603, N5601, N4539, N2021);
nor NOR4 (N5604, N5600, N171, N697, N4555);
nor NOR4 (N5605, N5603, N1777, N1635, N4751);
xor XOR2 (N5606, N5592, N5501);
not NOT1 (N5607, N5604);
not NOT1 (N5608, N5589);
nand NAND4 (N5609, N5596, N1004, N4627, N5483);
nor NOR3 (N5610, N5597, N1198, N1466);
nor NOR3 (N5611, N5608, N2530, N3570);
not NOT1 (N5612, N5605);
xor XOR2 (N5613, N5598, N2508);
xor XOR2 (N5614, N5609, N3007);
nand NAND3 (N5615, N5602, N4723, N2693);
not NOT1 (N5616, N5606);
not NOT1 (N5617, N5607);
xor XOR2 (N5618, N5599, N1278);
not NOT1 (N5619, N5611);
buf BUF1 (N5620, N5617);
not NOT1 (N5621, N5616);
nor NOR3 (N5622, N5618, N139, N4833);
nand NAND2 (N5623, N5612, N1869);
not NOT1 (N5624, N5576);
nor NOR2 (N5625, N5621, N3932);
or OR2 (N5626, N5623, N4757);
not NOT1 (N5627, N5626);
or OR3 (N5628, N5619, N3119, N1692);
nor NOR2 (N5629, N5620, N1764);
nor NOR2 (N5630, N5629, N5453);
buf BUF1 (N5631, N5613);
or OR3 (N5632, N5628, N5065, N59);
xor XOR2 (N5633, N5625, N4656);
or OR4 (N5634, N5614, N2177, N3693, N2668);
or OR3 (N5635, N5634, N1797, N2279);
nor NOR2 (N5636, N5615, N2081);
xor XOR2 (N5637, N5610, N4127);
not NOT1 (N5638, N5632);
nand NAND3 (N5639, N5636, N3273, N1888);
xor XOR2 (N5640, N5624, N2047);
buf BUF1 (N5641, N5638);
xor XOR2 (N5642, N5637, N1930);
nor NOR4 (N5643, N5633, N3132, N5287, N679);
xor XOR2 (N5644, N5643, N4810);
xor XOR2 (N5645, N5627, N1094);
xor XOR2 (N5646, N5635, N2693);
and AND4 (N5647, N5639, N5187, N21, N4432);
or OR2 (N5648, N5647, N1588);
nand NAND4 (N5649, N5631, N3772, N2964, N1697);
nor NOR4 (N5650, N5646, N4840, N723, N2390);
buf BUF1 (N5651, N5642);
or OR3 (N5652, N5650, N1949, N1953);
or OR2 (N5653, N5645, N2746);
and AND4 (N5654, N5653, N2091, N2824, N754);
and AND3 (N5655, N5640, N376, N4008);
xor XOR2 (N5656, N5655, N5227);
buf BUF1 (N5657, N5652);
and AND2 (N5658, N5648, N4293);
or OR3 (N5659, N5654, N2404, N5310);
xor XOR2 (N5660, N5659, N3486);
nor NOR4 (N5661, N5644, N855, N1051, N4033);
and AND4 (N5662, N5656, N1747, N1166, N681);
and AND2 (N5663, N5641, N1700);
buf BUF1 (N5664, N5651);
nor NOR3 (N5665, N5663, N305, N560);
not NOT1 (N5666, N5630);
nor NOR3 (N5667, N5662, N3421, N665);
not NOT1 (N5668, N5664);
xor XOR2 (N5669, N5658, N4971);
nor NOR2 (N5670, N5668, N3292);
and AND4 (N5671, N5670, N5411, N4139, N4868);
nor NOR3 (N5672, N5622, N5533, N779);
or OR3 (N5673, N5657, N3692, N1445);
buf BUF1 (N5674, N5669);
buf BUF1 (N5675, N5661);
nand NAND4 (N5676, N5660, N2070, N3687, N2870);
or OR2 (N5677, N5671, N659);
nor NOR4 (N5678, N5675, N2584, N4529, N216);
buf BUF1 (N5679, N5665);
nor NOR3 (N5680, N5679, N5337, N5356);
xor XOR2 (N5681, N5649, N2392);
buf BUF1 (N5682, N5676);
xor XOR2 (N5683, N5678, N491);
buf BUF1 (N5684, N5674);
not NOT1 (N5685, N5681);
nor NOR3 (N5686, N5672, N1119, N1567);
xor XOR2 (N5687, N5666, N3414);
nor NOR4 (N5688, N5673, N2642, N511, N1285);
not NOT1 (N5689, N5667);
nor NOR4 (N5690, N5688, N1384, N2378, N5136);
and AND2 (N5691, N5680, N5458);
nand NAND2 (N5692, N5687, N3900);
nand NAND2 (N5693, N5677, N3965);
and AND2 (N5694, N5691, N1368);
nand NAND4 (N5695, N5692, N433, N2524, N12);
not NOT1 (N5696, N5682);
or OR2 (N5697, N5684, N5550);
xor XOR2 (N5698, N5696, N4288);
buf BUF1 (N5699, N5698);
not NOT1 (N5700, N5699);
xor XOR2 (N5701, N5683, N3018);
and AND2 (N5702, N5690, N4507);
or OR3 (N5703, N5697, N3590, N3624);
nor NOR3 (N5704, N5689, N3660, N155);
xor XOR2 (N5705, N5694, N2184);
nor NOR3 (N5706, N5700, N1724, N3707);
and AND2 (N5707, N5705, N975);
xor XOR2 (N5708, N5695, N648);
not NOT1 (N5709, N5706);
nand NAND2 (N5710, N5701, N2640);
or OR3 (N5711, N5686, N4486, N3721);
and AND3 (N5712, N5707, N4377, N2246);
and AND4 (N5713, N5703, N3838, N1218, N615);
nand NAND2 (N5714, N5713, N4112);
or OR3 (N5715, N5693, N4828, N4521);
and AND3 (N5716, N5704, N2743, N5010);
xor XOR2 (N5717, N5685, N4254);
not NOT1 (N5718, N5710);
nor NOR2 (N5719, N5712, N3357);
nor NOR4 (N5720, N5714, N3487, N1020, N55);
buf BUF1 (N5721, N5718);
nor NOR3 (N5722, N5702, N2401, N1529);
and AND3 (N5723, N5708, N2087, N1377);
and AND3 (N5724, N5709, N439, N3279);
and AND4 (N5725, N5724, N4169, N2563, N2075);
buf BUF1 (N5726, N5721);
and AND3 (N5727, N5725, N1695, N3329);
xor XOR2 (N5728, N5715, N394);
or OR4 (N5729, N5727, N2546, N945, N2130);
nor NOR2 (N5730, N5728, N3061);
xor XOR2 (N5731, N5726, N3120);
nand NAND4 (N5732, N5717, N3390, N897, N539);
nor NOR3 (N5733, N5730, N1137, N4189);
not NOT1 (N5734, N5711);
buf BUF1 (N5735, N5716);
nor NOR3 (N5736, N5734, N3629, N5597);
not NOT1 (N5737, N5732);
not NOT1 (N5738, N5729);
nor NOR2 (N5739, N5735, N5472);
xor XOR2 (N5740, N5720, N3054);
xor XOR2 (N5741, N5733, N1375);
not NOT1 (N5742, N5741);
nand NAND2 (N5743, N5719, N2814);
nand NAND4 (N5744, N5738, N473, N512, N4774);
nor NOR3 (N5745, N5736, N4327, N5407);
or OR4 (N5746, N5740, N3660, N1109, N623);
buf BUF1 (N5747, N5723);
xor XOR2 (N5748, N5737, N1856);
nor NOR4 (N5749, N5747, N3588, N347, N528);
nand NAND2 (N5750, N5739, N4313);
xor XOR2 (N5751, N5750, N4634);
not NOT1 (N5752, N5748);
buf BUF1 (N5753, N5731);
nor NOR2 (N5754, N5746, N5226);
not NOT1 (N5755, N5742);
buf BUF1 (N5756, N5751);
and AND4 (N5757, N5752, N2882, N3381, N5226);
xor XOR2 (N5758, N5749, N3685);
and AND2 (N5759, N5757, N3438);
nand NAND3 (N5760, N5756, N1092, N2522);
buf BUF1 (N5761, N5722);
nand NAND3 (N5762, N5754, N358, N4478);
nor NOR4 (N5763, N5762, N4139, N876, N1034);
not NOT1 (N5764, N5744);
nand NAND4 (N5765, N5745, N2195, N4266, N3732);
nor NOR3 (N5766, N5753, N4232, N4759);
xor XOR2 (N5767, N5765, N1240);
not NOT1 (N5768, N5743);
and AND2 (N5769, N5767, N4492);
and AND2 (N5770, N5760, N1608);
or OR4 (N5771, N5764, N4535, N2177, N713);
not NOT1 (N5772, N5755);
not NOT1 (N5773, N5771);
buf BUF1 (N5774, N5772);
or OR3 (N5775, N5763, N714, N4524);
nand NAND4 (N5776, N5761, N5274, N2357, N4845);
not NOT1 (N5777, N5774);
or OR3 (N5778, N5759, N821, N1099);
or OR4 (N5779, N5770, N1514, N3556, N3503);
and AND3 (N5780, N5773, N5280, N1510);
buf BUF1 (N5781, N5775);
xor XOR2 (N5782, N5769, N753);
buf BUF1 (N5783, N5780);
nand NAND2 (N5784, N5779, N3060);
xor XOR2 (N5785, N5778, N5443);
not NOT1 (N5786, N5782);
buf BUF1 (N5787, N5781);
or OR3 (N5788, N5776, N737, N1939);
xor XOR2 (N5789, N5758, N3551);
nand NAND2 (N5790, N5777, N4698);
and AND3 (N5791, N5788, N144, N4413);
buf BUF1 (N5792, N5790);
buf BUF1 (N5793, N5783);
nor NOR2 (N5794, N5784, N3783);
nor NOR3 (N5795, N5768, N1335, N171);
and AND4 (N5796, N5791, N1831, N1417, N5726);
not NOT1 (N5797, N5785);
not NOT1 (N5798, N5794);
nand NAND2 (N5799, N5792, N800);
not NOT1 (N5800, N5795);
xor XOR2 (N5801, N5799, N3180);
nand NAND3 (N5802, N5796, N404, N5786);
not NOT1 (N5803, N2906);
xor XOR2 (N5804, N5793, N1033);
xor XOR2 (N5805, N5789, N407);
and AND3 (N5806, N5804, N4212, N3327);
not NOT1 (N5807, N5797);
or OR2 (N5808, N5800, N3936);
nor NOR2 (N5809, N5806, N1215);
xor XOR2 (N5810, N5803, N4578);
nand NAND4 (N5811, N5766, N1324, N1943, N1996);
nand NAND2 (N5812, N5807, N4943);
or OR4 (N5813, N5810, N3040, N5154, N1299);
buf BUF1 (N5814, N5802);
nand NAND2 (N5815, N5808, N1453);
not NOT1 (N5816, N5814);
buf BUF1 (N5817, N5809);
not NOT1 (N5818, N5817);
or OR3 (N5819, N5787, N5325, N2000);
xor XOR2 (N5820, N5812, N4380);
nor NOR2 (N5821, N5815, N2118);
buf BUF1 (N5822, N5820);
buf BUF1 (N5823, N5798);
nand NAND2 (N5824, N5818, N5465);
buf BUF1 (N5825, N5823);
buf BUF1 (N5826, N5816);
buf BUF1 (N5827, N5801);
buf BUF1 (N5828, N5811);
not NOT1 (N5829, N5819);
not NOT1 (N5830, N5827);
nand NAND4 (N5831, N5813, N1841, N3905, N3057);
nor NOR4 (N5832, N5829, N5214, N2582, N1045);
or OR4 (N5833, N5830, N2093, N1999, N333);
nand NAND3 (N5834, N5826, N686, N727);
xor XOR2 (N5835, N5834, N438);
nand NAND4 (N5836, N5825, N1704, N5071, N1186);
or OR3 (N5837, N5835, N3772, N630);
or OR4 (N5838, N5822, N220, N5661, N870);
buf BUF1 (N5839, N5821);
or OR2 (N5840, N5838, N408);
nand NAND3 (N5841, N5805, N4801, N2413);
buf BUF1 (N5842, N5831);
nand NAND3 (N5843, N5824, N4676, N1242);
or OR3 (N5844, N5832, N1631, N5012);
and AND2 (N5845, N5841, N819);
xor XOR2 (N5846, N5836, N4768);
nand NAND2 (N5847, N5833, N3998);
buf BUF1 (N5848, N5844);
and AND2 (N5849, N5828, N4313);
nand NAND2 (N5850, N5848, N3254);
buf BUF1 (N5851, N5842);
or OR4 (N5852, N5849, N879, N4500, N2064);
nand NAND2 (N5853, N5852, N905);
buf BUF1 (N5854, N5846);
xor XOR2 (N5855, N5853, N670);
or OR2 (N5856, N5855, N2498);
not NOT1 (N5857, N5840);
not NOT1 (N5858, N5837);
buf BUF1 (N5859, N5854);
nor NOR2 (N5860, N5851, N4952);
buf BUF1 (N5861, N5847);
and AND2 (N5862, N5857, N1267);
and AND3 (N5863, N5850, N4502, N724);
xor XOR2 (N5864, N5861, N796);
buf BUF1 (N5865, N5858);
xor XOR2 (N5866, N5845, N4089);
nand NAND2 (N5867, N5839, N4913);
or OR3 (N5868, N5860, N1925, N1834);
or OR4 (N5869, N5863, N2740, N2721, N5340);
and AND4 (N5870, N5867, N3375, N1404, N1217);
or OR4 (N5871, N5862, N4039, N2716, N5794);
nand NAND2 (N5872, N5871, N26);
xor XOR2 (N5873, N5859, N945);
or OR4 (N5874, N5843, N2848, N937, N2311);
not NOT1 (N5875, N5870);
or OR3 (N5876, N5868, N3759, N1835);
buf BUF1 (N5877, N5872);
xor XOR2 (N5878, N5869, N4935);
xor XOR2 (N5879, N5877, N1842);
nand NAND2 (N5880, N5864, N4634);
xor XOR2 (N5881, N5873, N3527);
nand NAND4 (N5882, N5874, N2250, N5717, N452);
or OR4 (N5883, N5865, N1208, N2865, N701);
or OR4 (N5884, N5866, N953, N5073, N2875);
nor NOR4 (N5885, N5882, N5465, N2220, N2963);
xor XOR2 (N5886, N5875, N4169);
and AND2 (N5887, N5876, N3051);
not NOT1 (N5888, N5879);
xor XOR2 (N5889, N5887, N1833);
nand NAND2 (N5890, N5886, N832);
nor NOR3 (N5891, N5888, N2393, N1601);
or OR3 (N5892, N5881, N2426, N548);
nor NOR4 (N5893, N5891, N1376, N1959, N1095);
nor NOR3 (N5894, N5856, N507, N838);
buf BUF1 (N5895, N5878);
not NOT1 (N5896, N5880);
or OR4 (N5897, N5890, N2608, N3715, N3939);
buf BUF1 (N5898, N5892);
and AND3 (N5899, N5889, N3114, N2982);
nand NAND3 (N5900, N5899, N4904, N918);
xor XOR2 (N5901, N5883, N5425);
nand NAND2 (N5902, N5898, N38);
or OR3 (N5903, N5894, N2762, N122);
nor NOR2 (N5904, N5893, N2545);
not NOT1 (N5905, N5895);
xor XOR2 (N5906, N5902, N5658);
or OR4 (N5907, N5901, N924, N339, N116);
not NOT1 (N5908, N5904);
buf BUF1 (N5909, N5884);
xor XOR2 (N5910, N5903, N4044);
xor XOR2 (N5911, N5908, N5722);
and AND2 (N5912, N5885, N673);
and AND2 (N5913, N5905, N3232);
nand NAND4 (N5914, N5900, N4325, N5340, N1124);
nand NAND2 (N5915, N5910, N3436);
and AND4 (N5916, N5907, N2924, N2640, N3636);
or OR4 (N5917, N5915, N1059, N350, N2774);
xor XOR2 (N5918, N5909, N4702);
nor NOR2 (N5919, N5906, N4494);
buf BUF1 (N5920, N5913);
and AND4 (N5921, N5916, N5528, N1499, N2850);
not NOT1 (N5922, N5917);
not NOT1 (N5923, N5919);
nand NAND2 (N5924, N5920, N337);
xor XOR2 (N5925, N5896, N5385);
xor XOR2 (N5926, N5925, N1269);
nand NAND4 (N5927, N5912, N2198, N1514, N5595);
nor NOR3 (N5928, N5921, N5203, N1877);
buf BUF1 (N5929, N5927);
and AND2 (N5930, N5929, N5137);
buf BUF1 (N5931, N5923);
xor XOR2 (N5932, N5924, N1662);
xor XOR2 (N5933, N5932, N689);
buf BUF1 (N5934, N5933);
and AND4 (N5935, N5897, N4551, N4521, N3108);
not NOT1 (N5936, N5930);
nand NAND4 (N5937, N5928, N1380, N2244, N3158);
and AND2 (N5938, N5936, N5680);
buf BUF1 (N5939, N5914);
not NOT1 (N5940, N5939);
and AND4 (N5941, N5918, N4735, N5497, N4298);
nor NOR3 (N5942, N5911, N5305, N2047);
and AND2 (N5943, N5922, N5090);
xor XOR2 (N5944, N5941, N4329);
not NOT1 (N5945, N5937);
buf BUF1 (N5946, N5931);
buf BUF1 (N5947, N5938);
nand NAND3 (N5948, N5945, N5241, N3711);
buf BUF1 (N5949, N5935);
and AND4 (N5950, N5946, N2472, N199, N1724);
nand NAND2 (N5951, N5947, N2712);
nand NAND2 (N5952, N5926, N1489);
nand NAND4 (N5953, N5950, N4912, N2245, N4977);
buf BUF1 (N5954, N5940);
buf BUF1 (N5955, N5954);
nor NOR4 (N5956, N5942, N2221, N5797, N797);
nand NAND2 (N5957, N5949, N2793);
buf BUF1 (N5958, N5953);
xor XOR2 (N5959, N5934, N2241);
and AND4 (N5960, N5943, N5217, N1132, N1409);
nor NOR4 (N5961, N5958, N509, N2304, N5761);
nor NOR4 (N5962, N5960, N2864, N4259, N3678);
xor XOR2 (N5963, N5948, N857);
not NOT1 (N5964, N5957);
nand NAND4 (N5965, N5951, N3131, N825, N4527);
nand NAND2 (N5966, N5962, N4196);
buf BUF1 (N5967, N5955);
or OR3 (N5968, N5967, N2765, N1712);
xor XOR2 (N5969, N5966, N4594);
nand NAND3 (N5970, N5965, N5376, N4847);
not NOT1 (N5971, N5970);
not NOT1 (N5972, N5968);
and AND3 (N5973, N5956, N1328, N507);
nand NAND3 (N5974, N5969, N5174, N5016);
not NOT1 (N5975, N5952);
not NOT1 (N5976, N5971);
nand NAND2 (N5977, N5975, N4393);
not NOT1 (N5978, N5964);
nor NOR3 (N5979, N5959, N2237, N397);
not NOT1 (N5980, N5944);
not NOT1 (N5981, N5977);
nand NAND2 (N5982, N5963, N1218);
nand NAND2 (N5983, N5979, N949);
or OR3 (N5984, N5972, N5947, N1950);
nand NAND4 (N5985, N5976, N1135, N4486, N4886);
xor XOR2 (N5986, N5981, N656);
and AND3 (N5987, N5980, N434, N5272);
nor NOR3 (N5988, N5961, N1309, N4370);
xor XOR2 (N5989, N5986, N1883);
not NOT1 (N5990, N5989);
or OR3 (N5991, N5988, N357, N2969);
not NOT1 (N5992, N5984);
not NOT1 (N5993, N5985);
and AND4 (N5994, N5973, N1279, N5348, N2623);
buf BUF1 (N5995, N5982);
nor NOR2 (N5996, N5993, N2366);
and AND4 (N5997, N5994, N3056, N5874, N5166);
or OR4 (N5998, N5974, N689, N4381, N3043);
not NOT1 (N5999, N5998);
buf BUF1 (N6000, N5995);
not NOT1 (N6001, N5983);
nand NAND4 (N6002, N5987, N5787, N5483, N1855);
xor XOR2 (N6003, N5996, N1028);
or OR2 (N6004, N5991, N3892);
xor XOR2 (N6005, N5992, N3515);
or OR3 (N6006, N6001, N3031, N1743);
and AND2 (N6007, N5990, N1606);
or OR4 (N6008, N6007, N2010, N4963, N4318);
buf BUF1 (N6009, N6005);
or OR3 (N6010, N5999, N4388, N2767);
buf BUF1 (N6011, N6004);
buf BUF1 (N6012, N6011);
buf BUF1 (N6013, N6000);
nand NAND2 (N6014, N6013, N5503);
not NOT1 (N6015, N6009);
and AND2 (N6016, N6006, N5667);
not NOT1 (N6017, N6014);
buf BUF1 (N6018, N6012);
and AND4 (N6019, N6003, N4703, N76, N5942);
not NOT1 (N6020, N6002);
nand NAND4 (N6021, N6018, N5567, N4331, N647);
nand NAND3 (N6022, N6010, N1757, N1658);
buf BUF1 (N6023, N6008);
not NOT1 (N6024, N6021);
not NOT1 (N6025, N6022);
xor XOR2 (N6026, N6025, N3894);
buf BUF1 (N6027, N6026);
nand NAND2 (N6028, N5997, N5857);
nor NOR4 (N6029, N6020, N140, N5254, N1695);
or OR4 (N6030, N6016, N1826, N277, N5376);
xor XOR2 (N6031, N6017, N1315);
xor XOR2 (N6032, N5978, N476);
not NOT1 (N6033, N6031);
buf BUF1 (N6034, N6015);
nor NOR3 (N6035, N6027, N5073, N3992);
nand NAND4 (N6036, N6035, N3419, N4663, N3632);
nor NOR2 (N6037, N6028, N1375);
nor NOR2 (N6038, N6034, N119);
buf BUF1 (N6039, N6029);
xor XOR2 (N6040, N6037, N3284);
buf BUF1 (N6041, N6032);
nand NAND2 (N6042, N6019, N4357);
nand NAND3 (N6043, N6033, N1320, N1223);
buf BUF1 (N6044, N6023);
xor XOR2 (N6045, N6042, N4952);
nor NOR4 (N6046, N6030, N5914, N4556, N5439);
nor NOR3 (N6047, N6036, N5206, N479);
or OR4 (N6048, N6039, N1593, N4511, N3819);
nand NAND3 (N6049, N6038, N5584, N997);
buf BUF1 (N6050, N6041);
or OR2 (N6051, N6043, N4094);
or OR3 (N6052, N6048, N3363, N779);
not NOT1 (N6053, N6052);
buf BUF1 (N6054, N6045);
and AND2 (N6055, N6040, N1007);
xor XOR2 (N6056, N6046, N4403);
and AND2 (N6057, N6056, N393);
nor NOR4 (N6058, N6024, N1893, N5488, N2023);
or OR4 (N6059, N6053, N382, N4000, N1055);
nand NAND3 (N6060, N6047, N5356, N3535);
and AND3 (N6061, N6058, N1479, N2557);
nand NAND3 (N6062, N6054, N5379, N5973);
nor NOR2 (N6063, N6062, N3631);
xor XOR2 (N6064, N6055, N4663);
or OR2 (N6065, N6063, N743);
nor NOR2 (N6066, N6065, N4066);
and AND2 (N6067, N6051, N4648);
and AND2 (N6068, N6066, N3988);
and AND4 (N6069, N6050, N3534, N1802, N4246);
buf BUF1 (N6070, N6049);
and AND4 (N6071, N6060, N4669, N3631, N4539);
and AND3 (N6072, N6044, N5938, N3147);
not NOT1 (N6073, N6068);
nor NOR2 (N6074, N6069, N5373);
nor NOR4 (N6075, N6070, N3760, N5193, N4663);
nand NAND4 (N6076, N6071, N4893, N326, N1650);
xor XOR2 (N6077, N6076, N770);
and AND3 (N6078, N6075, N4047, N3454);
or OR4 (N6079, N6057, N3056, N2449, N1422);
nand NAND2 (N6080, N6078, N1990);
buf BUF1 (N6081, N6061);
or OR4 (N6082, N6059, N1203, N1001, N3136);
and AND4 (N6083, N6077, N5769, N4495, N404);
buf BUF1 (N6084, N6067);
buf BUF1 (N6085, N6074);
xor XOR2 (N6086, N6073, N5285);
nor NOR4 (N6087, N6081, N3416, N5666, N1570);
and AND3 (N6088, N6086, N3331, N1147);
buf BUF1 (N6089, N6082);
not NOT1 (N6090, N6079);
nand NAND2 (N6091, N6080, N1962);
nand NAND3 (N6092, N6088, N1630, N3132);
and AND4 (N6093, N6064, N1621, N687, N1394);
or OR3 (N6094, N6085, N5398, N2216);
or OR3 (N6095, N6087, N356, N2817);
nor NOR3 (N6096, N6084, N3304, N1617);
not NOT1 (N6097, N6072);
not NOT1 (N6098, N6092);
and AND4 (N6099, N6093, N2018, N5903, N5456);
and AND4 (N6100, N6099, N5514, N4679, N5269);
buf BUF1 (N6101, N6089);
buf BUF1 (N6102, N6100);
xor XOR2 (N6103, N6090, N3795);
nor NOR2 (N6104, N6098, N2986);
buf BUF1 (N6105, N6103);
nor NOR4 (N6106, N6091, N3050, N5895, N265);
or OR2 (N6107, N6102, N965);
nand NAND4 (N6108, N6083, N266, N5525, N4351);
nand NAND2 (N6109, N6108, N1480);
and AND4 (N6110, N6094, N2165, N2026, N2699);
xor XOR2 (N6111, N6107, N249);
nand NAND3 (N6112, N6096, N1340, N766);
and AND4 (N6113, N6101, N2062, N2946, N5533);
xor XOR2 (N6114, N6110, N2237);
and AND3 (N6115, N6114, N3526, N3881);
buf BUF1 (N6116, N6105);
nor NOR2 (N6117, N6115, N4380);
buf BUF1 (N6118, N6097);
and AND2 (N6119, N6112, N3862);
xor XOR2 (N6120, N6106, N5738);
and AND3 (N6121, N6119, N5959, N430);
buf BUF1 (N6122, N6109);
nor NOR4 (N6123, N6117, N3593, N1693, N4225);
xor XOR2 (N6124, N6118, N4989);
xor XOR2 (N6125, N6095, N367);
nor NOR3 (N6126, N6121, N256, N4574);
xor XOR2 (N6127, N6120, N4182);
and AND3 (N6128, N6113, N5171, N4561);
nand NAND4 (N6129, N6126, N6123, N4201, N2471);
nor NOR4 (N6130, N448, N496, N2842, N3197);
buf BUF1 (N6131, N6104);
or OR2 (N6132, N6116, N796);
or OR2 (N6133, N6127, N2648);
buf BUF1 (N6134, N6124);
not NOT1 (N6135, N6132);
not NOT1 (N6136, N6131);
nand NAND2 (N6137, N6130, N3453);
xor XOR2 (N6138, N6133, N4011);
buf BUF1 (N6139, N6135);
nand NAND4 (N6140, N6138, N1495, N4560, N713);
and AND4 (N6141, N6111, N3227, N1475, N1003);
not NOT1 (N6142, N6122);
buf BUF1 (N6143, N6134);
buf BUF1 (N6144, N6143);
and AND3 (N6145, N6139, N3760, N5142);
or OR2 (N6146, N6145, N5588);
xor XOR2 (N6147, N6142, N4242);
nor NOR4 (N6148, N6125, N749, N2873, N5431);
xor XOR2 (N6149, N6148, N2196);
nor NOR4 (N6150, N6144, N5581, N1007, N1598);
not NOT1 (N6151, N6150);
nand NAND3 (N6152, N6151, N798, N392);
not NOT1 (N6153, N6149);
or OR3 (N6154, N6129, N878, N1615);
xor XOR2 (N6155, N6141, N1188);
nand NAND4 (N6156, N6146, N452, N2323, N4128);
xor XOR2 (N6157, N6140, N2703);
nor NOR2 (N6158, N6156, N6048);
not NOT1 (N6159, N6158);
nor NOR2 (N6160, N6153, N1637);
and AND3 (N6161, N6152, N3835, N2182);
or OR4 (N6162, N6137, N2813, N373, N3028);
and AND4 (N6163, N6155, N131, N93, N1516);
or OR3 (N6164, N6147, N2828, N5076);
or OR3 (N6165, N6160, N1937, N5573);
buf BUF1 (N6166, N6159);
or OR2 (N6167, N6164, N5083);
nor NOR4 (N6168, N6128, N4672, N2256, N3449);
or OR2 (N6169, N6154, N3497);
or OR2 (N6170, N6157, N4995);
or OR2 (N6171, N6161, N1659);
or OR3 (N6172, N6163, N3263, N1738);
buf BUF1 (N6173, N6166);
buf BUF1 (N6174, N6169);
nor NOR2 (N6175, N6165, N110);
nor NOR3 (N6176, N6175, N4078, N2126);
and AND4 (N6177, N6172, N1746, N2199, N2175);
nand NAND2 (N6178, N6170, N5476);
nor NOR4 (N6179, N6168, N440, N3054, N1044);
nor NOR2 (N6180, N6178, N4669);
xor XOR2 (N6181, N6174, N4839);
or OR4 (N6182, N6136, N2300, N2064, N4219);
nor NOR4 (N6183, N6171, N3608, N1542, N5651);
nand NAND3 (N6184, N6183, N5995, N494);
nand NAND3 (N6185, N6184, N2455, N5980);
buf BUF1 (N6186, N6185);
nand NAND3 (N6187, N6179, N3655, N1840);
nand NAND3 (N6188, N6186, N4474, N1111);
nand NAND4 (N6189, N6177, N4234, N5769, N5816);
not NOT1 (N6190, N6176);
buf BUF1 (N6191, N6188);
xor XOR2 (N6192, N6167, N5317);
buf BUF1 (N6193, N6173);
or OR2 (N6194, N6190, N4669);
nor NOR2 (N6195, N6182, N488);
nand NAND3 (N6196, N6191, N5324, N2034);
or OR2 (N6197, N6162, N4197);
xor XOR2 (N6198, N6193, N2187);
and AND3 (N6199, N6194, N985, N167);
xor XOR2 (N6200, N6189, N442);
nor NOR4 (N6201, N6200, N544, N1630, N4230);
and AND3 (N6202, N6187, N5091, N4176);
and AND2 (N6203, N6197, N1528);
not NOT1 (N6204, N6203);
or OR4 (N6205, N6192, N5801, N5385, N2433);
nor NOR4 (N6206, N6201, N2332, N602, N5659);
nand NAND4 (N6207, N6180, N720, N406, N1716);
not NOT1 (N6208, N6199);
and AND4 (N6209, N6198, N302, N1302, N4070);
xor XOR2 (N6210, N6181, N4468);
or OR2 (N6211, N6206, N1654);
nor NOR4 (N6212, N6210, N35, N126, N1559);
nand NAND2 (N6213, N6212, N6033);
nor NOR4 (N6214, N6205, N412, N3450, N5962);
not NOT1 (N6215, N6195);
or OR2 (N6216, N6202, N5555);
not NOT1 (N6217, N6204);
xor XOR2 (N6218, N6214, N986);
and AND4 (N6219, N6218, N3374, N1039, N5670);
nand NAND2 (N6220, N6215, N5869);
not NOT1 (N6221, N6213);
or OR4 (N6222, N6208, N3837, N3724, N3483);
xor XOR2 (N6223, N6211, N174);
xor XOR2 (N6224, N6219, N4024);
xor XOR2 (N6225, N6216, N4367);
not NOT1 (N6226, N6224);
xor XOR2 (N6227, N6225, N1748);
xor XOR2 (N6228, N6220, N1340);
not NOT1 (N6229, N6222);
not NOT1 (N6230, N6227);
xor XOR2 (N6231, N6209, N1667);
nor NOR4 (N6232, N6196, N4113, N2120, N1982);
not NOT1 (N6233, N6221);
not NOT1 (N6234, N6228);
nand NAND2 (N6235, N6217, N4007);
and AND4 (N6236, N6233, N3137, N3498, N1228);
nor NOR3 (N6237, N6234, N2807, N506);
buf BUF1 (N6238, N6223);
nor NOR3 (N6239, N6235, N2255, N4541);
xor XOR2 (N6240, N6238, N3727);
or OR3 (N6241, N6231, N5317, N488);
not NOT1 (N6242, N6232);
buf BUF1 (N6243, N6240);
xor XOR2 (N6244, N6207, N5278);
and AND3 (N6245, N6244, N2660, N3925);
xor XOR2 (N6246, N6226, N1734);
nor NOR4 (N6247, N6236, N3414, N5385, N4016);
nor NOR4 (N6248, N6230, N3681, N715, N3150);
nor NOR3 (N6249, N6237, N4165, N839);
nand NAND4 (N6250, N6243, N3230, N3975, N933);
xor XOR2 (N6251, N6249, N3691);
xor XOR2 (N6252, N6246, N6113);
buf BUF1 (N6253, N6248);
and AND3 (N6254, N6229, N5758, N3976);
not NOT1 (N6255, N6247);
not NOT1 (N6256, N6254);
xor XOR2 (N6257, N6253, N253);
or OR4 (N6258, N6256, N2900, N4268, N2004);
nand NAND4 (N6259, N6245, N3422, N1160, N6235);
buf BUF1 (N6260, N6255);
xor XOR2 (N6261, N6250, N2928);
nand NAND3 (N6262, N6261, N2004, N4856);
nor NOR2 (N6263, N6251, N3378);
and AND2 (N6264, N6260, N3728);
nor NOR2 (N6265, N6262, N2162);
or OR2 (N6266, N6263, N4204);
nor NOR4 (N6267, N6266, N2263, N2043, N3394);
and AND4 (N6268, N6267, N130, N3435, N1726);
and AND3 (N6269, N6241, N1158, N2668);
buf BUF1 (N6270, N6264);
nor NOR4 (N6271, N6242, N5811, N2619, N3053);
nor NOR2 (N6272, N6270, N1892);
nor NOR4 (N6273, N6268, N1828, N981, N3909);
buf BUF1 (N6274, N6272);
nand NAND4 (N6275, N6252, N783, N1015, N5463);
buf BUF1 (N6276, N6275);
and AND3 (N6277, N6258, N1252, N3972);
buf BUF1 (N6278, N6239);
nand NAND4 (N6279, N6257, N229, N4690, N861);
not NOT1 (N6280, N6277);
or OR4 (N6281, N6269, N4000, N5748, N1944);
and AND4 (N6282, N6278, N4668, N4571, N4699);
nand NAND3 (N6283, N6280, N3141, N713);
buf BUF1 (N6284, N6274);
or OR4 (N6285, N6265, N2002, N1668, N3370);
buf BUF1 (N6286, N6271);
nand NAND3 (N6287, N6282, N2216, N3781);
or OR2 (N6288, N6284, N1236);
nand NAND4 (N6289, N6273, N1178, N5872, N1240);
or OR3 (N6290, N6289, N356, N1670);
nand NAND4 (N6291, N6259, N2439, N492, N4460);
nand NAND2 (N6292, N6290, N4807);
nor NOR3 (N6293, N6286, N3550, N730);
buf BUF1 (N6294, N6283);
buf BUF1 (N6295, N6293);
xor XOR2 (N6296, N6279, N5657);
nor NOR4 (N6297, N6276, N4406, N6038, N1336);
not NOT1 (N6298, N6292);
not NOT1 (N6299, N6287);
nand NAND2 (N6300, N6297, N2932);
nor NOR3 (N6301, N6298, N5019, N1976);
buf BUF1 (N6302, N6301);
xor XOR2 (N6303, N6302, N210);
nor NOR2 (N6304, N6281, N4690);
or OR4 (N6305, N6304, N92, N659, N1742);
nor NOR3 (N6306, N6303, N3482, N6114);
nor NOR3 (N6307, N6288, N3679, N6248);
not NOT1 (N6308, N6305);
not NOT1 (N6309, N6294);
buf BUF1 (N6310, N6309);
nor NOR4 (N6311, N6291, N1613, N1195, N5372);
not NOT1 (N6312, N6308);
nor NOR4 (N6313, N6306, N1989, N1751, N4819);
or OR4 (N6314, N6300, N2167, N6025, N1753);
or OR2 (N6315, N6299, N1351);
nor NOR3 (N6316, N6313, N2604, N1367);
not NOT1 (N6317, N6315);
not NOT1 (N6318, N6310);
nor NOR4 (N6319, N6285, N1889, N1623, N1319);
nor NOR4 (N6320, N6312, N1409, N3313, N4255);
xor XOR2 (N6321, N6316, N4);
not NOT1 (N6322, N6311);
not NOT1 (N6323, N6322);
and AND2 (N6324, N6319, N4938);
not NOT1 (N6325, N6295);
not NOT1 (N6326, N6318);
xor XOR2 (N6327, N6317, N738);
not NOT1 (N6328, N6314);
nand NAND3 (N6329, N6323, N6125, N2715);
or OR2 (N6330, N6325, N5405);
nand NAND2 (N6331, N6307, N6183);
nor NOR3 (N6332, N6327, N1477, N4538);
nand NAND4 (N6333, N6330, N2287, N322, N1410);
nor NOR2 (N6334, N6332, N133);
and AND4 (N6335, N6331, N1419, N1140, N1851);
xor XOR2 (N6336, N6333, N17);
not NOT1 (N6337, N6336);
or OR4 (N6338, N6328, N4604, N1065, N758);
nand NAND2 (N6339, N6338, N5419);
nor NOR4 (N6340, N6334, N5990, N5601, N2188);
nand NAND3 (N6341, N6324, N5703, N298);
and AND3 (N6342, N6341, N2771, N1398);
xor XOR2 (N6343, N6321, N2681);
xor XOR2 (N6344, N6343, N3206);
xor XOR2 (N6345, N6339, N4737);
xor XOR2 (N6346, N6329, N5943);
buf BUF1 (N6347, N6344);
and AND2 (N6348, N6337, N1664);
or OR3 (N6349, N6335, N5899, N347);
buf BUF1 (N6350, N6326);
or OR4 (N6351, N6350, N3656, N674, N4751);
nor NOR2 (N6352, N6346, N554);
and AND3 (N6353, N6345, N3323, N2365);
and AND2 (N6354, N6340, N451);
not NOT1 (N6355, N6353);
xor XOR2 (N6356, N6354, N1791);
buf BUF1 (N6357, N6352);
nor NOR3 (N6358, N6349, N5822, N5392);
buf BUF1 (N6359, N6358);
or OR2 (N6360, N6348, N2208);
not NOT1 (N6361, N6360);
buf BUF1 (N6362, N6347);
or OR2 (N6363, N6320, N5600);
nor NOR3 (N6364, N6359, N5005, N433);
and AND3 (N6365, N6362, N5412, N5990);
and AND4 (N6366, N6296, N5085, N2460, N4283);
nor NOR4 (N6367, N6357, N5100, N2461, N3894);
and AND3 (N6368, N6351, N2193, N3018);
not NOT1 (N6369, N6367);
xor XOR2 (N6370, N6356, N2164);
xor XOR2 (N6371, N6342, N2589);
or OR2 (N6372, N6368, N1024);
nor NOR2 (N6373, N6370, N4220);
nor NOR3 (N6374, N6373, N5207, N2678);
or OR3 (N6375, N6363, N4124, N4552);
xor XOR2 (N6376, N6372, N3788);
and AND3 (N6377, N6371, N3195, N3110);
or OR2 (N6378, N6365, N4273);
nand NAND4 (N6379, N6374, N4330, N3013, N3322);
or OR4 (N6380, N6369, N262, N2964, N1151);
buf BUF1 (N6381, N6375);
or OR4 (N6382, N6380, N610, N2832, N6066);
xor XOR2 (N6383, N6378, N4845);
not NOT1 (N6384, N6366);
nand NAND4 (N6385, N6382, N3110, N552, N1650);
and AND4 (N6386, N6385, N785, N1733, N267);
nand NAND3 (N6387, N6386, N3169, N251);
and AND3 (N6388, N6387, N2913, N5327);
nand NAND2 (N6389, N6384, N2202);
or OR3 (N6390, N6381, N2068, N2808);
xor XOR2 (N6391, N6388, N2023);
nor NOR4 (N6392, N6379, N1920, N875, N1072);
or OR4 (N6393, N6391, N4628, N513, N4190);
xor XOR2 (N6394, N6393, N2417);
nand NAND2 (N6395, N6361, N867);
nand NAND2 (N6396, N6395, N3923);
buf BUF1 (N6397, N6355);
not NOT1 (N6398, N6364);
or OR2 (N6399, N6376, N4900);
buf BUF1 (N6400, N6398);
or OR2 (N6401, N6394, N4025);
xor XOR2 (N6402, N6396, N5800);
nor NOR3 (N6403, N6377, N543, N4790);
and AND4 (N6404, N6399, N5390, N2815, N724);
and AND4 (N6405, N6403, N5956, N680, N4228);
nor NOR2 (N6406, N6397, N4352);
or OR2 (N6407, N6404, N1106);
nand NAND3 (N6408, N6406, N1470, N761);
buf BUF1 (N6409, N6401);
and AND2 (N6410, N6392, N44);
nand NAND2 (N6411, N6408, N3962);
not NOT1 (N6412, N6410);
buf BUF1 (N6413, N6405);
or OR4 (N6414, N6383, N561, N6159, N5631);
not NOT1 (N6415, N6411);
nor NOR2 (N6416, N6409, N328);
not NOT1 (N6417, N6412);
or OR3 (N6418, N6417, N3458, N1548);
not NOT1 (N6419, N6416);
not NOT1 (N6420, N6390);
and AND2 (N6421, N6414, N4932);
or OR3 (N6422, N6389, N6306, N4559);
xor XOR2 (N6423, N6415, N5202);
nor NOR3 (N6424, N6423, N3186, N3204);
and AND2 (N6425, N6402, N3054);
xor XOR2 (N6426, N6420, N2276);
or OR3 (N6427, N6426, N4376, N464);
not NOT1 (N6428, N6400);
buf BUF1 (N6429, N6418);
xor XOR2 (N6430, N6419, N3081);
not NOT1 (N6431, N6422);
xor XOR2 (N6432, N6421, N3458);
or OR4 (N6433, N6424, N1514, N552, N261);
and AND4 (N6434, N6432, N4407, N6386, N5391);
xor XOR2 (N6435, N6425, N339);
not NOT1 (N6436, N6413);
nor NOR4 (N6437, N6427, N3746, N2405, N4053);
nor NOR4 (N6438, N6433, N4926, N1028, N2819);
and AND2 (N6439, N6430, N6374);
nor NOR4 (N6440, N6436, N3275, N854, N3315);
buf BUF1 (N6441, N6435);
and AND2 (N6442, N6439, N6014);
xor XOR2 (N6443, N6441, N353);
or OR4 (N6444, N6431, N137, N1559, N144);
not NOT1 (N6445, N6443);
buf BUF1 (N6446, N6437);
and AND4 (N6447, N6438, N1881, N5440, N5705);
or OR2 (N6448, N6407, N2775);
and AND2 (N6449, N6444, N4838);
or OR4 (N6450, N6446, N2177, N1244, N2374);
or OR3 (N6451, N6442, N5891, N6197);
not NOT1 (N6452, N6448);
or OR3 (N6453, N6434, N1345, N622);
or OR4 (N6454, N6453, N2979, N5700, N5927);
xor XOR2 (N6455, N6440, N4347);
and AND3 (N6456, N6452, N2523, N3997);
not NOT1 (N6457, N6449);
buf BUF1 (N6458, N6451);
and AND4 (N6459, N6456, N4655, N1728, N1811);
nand NAND2 (N6460, N6457, N1802);
not NOT1 (N6461, N6445);
buf BUF1 (N6462, N6447);
or OR4 (N6463, N6450, N5427, N5329, N4475);
or OR2 (N6464, N6461, N143);
nand NAND2 (N6465, N6460, N5012);
not NOT1 (N6466, N6429);
nand NAND3 (N6467, N6454, N5082, N1644);
not NOT1 (N6468, N6467);
xor XOR2 (N6469, N6428, N5493);
buf BUF1 (N6470, N6465);
buf BUF1 (N6471, N6463);
or OR2 (N6472, N6455, N6150);
xor XOR2 (N6473, N6469, N981);
nand NAND2 (N6474, N6458, N1902);
or OR4 (N6475, N6472, N2533, N1644, N2185);
and AND2 (N6476, N6470, N5143);
or OR3 (N6477, N6471, N3031, N2232);
or OR3 (N6478, N6468, N2917, N6014);
xor XOR2 (N6479, N6477, N5784);
buf BUF1 (N6480, N6479);
and AND2 (N6481, N6462, N3441);
buf BUF1 (N6482, N6476);
or OR4 (N6483, N6480, N4218, N2506, N2630);
nor NOR2 (N6484, N6482, N5129);
not NOT1 (N6485, N6481);
nand NAND3 (N6486, N6464, N3136, N3419);
not NOT1 (N6487, N6475);
and AND4 (N6488, N6487, N914, N4632, N4362);
not NOT1 (N6489, N6474);
or OR4 (N6490, N6484, N4890, N75, N5058);
xor XOR2 (N6491, N6488, N2178);
not NOT1 (N6492, N6491);
or OR4 (N6493, N6459, N5542, N1881, N3818);
not NOT1 (N6494, N6478);
not NOT1 (N6495, N6466);
nor NOR2 (N6496, N6483, N430);
xor XOR2 (N6497, N6485, N464);
buf BUF1 (N6498, N6495);
or OR2 (N6499, N6486, N5607);
not NOT1 (N6500, N6494);
buf BUF1 (N6501, N6500);
or OR3 (N6502, N6499, N3242, N6335);
nand NAND2 (N6503, N6490, N6341);
xor XOR2 (N6504, N6502, N921);
not NOT1 (N6505, N6504);
nor NOR4 (N6506, N6498, N3680, N2571, N1079);
not NOT1 (N6507, N6473);
buf BUF1 (N6508, N6497);
nor NOR4 (N6509, N6493, N1301, N5693, N948);
xor XOR2 (N6510, N6501, N5120);
nor NOR2 (N6511, N6509, N854);
nand NAND3 (N6512, N6507, N6127, N1373);
not NOT1 (N6513, N6511);
or OR3 (N6514, N6510, N4154, N854);
nor NOR3 (N6515, N6506, N3170, N567);
nor NOR3 (N6516, N6513, N3329, N1887);
buf BUF1 (N6517, N6508);
and AND4 (N6518, N6489, N2033, N5406, N4925);
nor NOR2 (N6519, N6512, N2038);
nor NOR4 (N6520, N6505, N4023, N4943, N5366);
nor NOR4 (N6521, N6496, N2404, N2219, N3387);
nand NAND3 (N6522, N6521, N4139, N4726);
nand NAND2 (N6523, N6522, N1192);
and AND4 (N6524, N6514, N4180, N4724, N1814);
buf BUF1 (N6525, N6515);
nor NOR2 (N6526, N6525, N1399);
nand NAND2 (N6527, N6526, N3292);
nor NOR4 (N6528, N6492, N2965, N2149, N6149);
xor XOR2 (N6529, N6516, N1702);
or OR3 (N6530, N6528, N816, N2389);
buf BUF1 (N6531, N6518);
and AND4 (N6532, N6520, N772, N6490, N4741);
xor XOR2 (N6533, N6527, N3014);
nand NAND3 (N6534, N6517, N833, N6203);
buf BUF1 (N6535, N6523);
xor XOR2 (N6536, N6534, N4111);
or OR4 (N6537, N6531, N6052, N4982, N1351);
and AND2 (N6538, N6530, N4044);
buf BUF1 (N6539, N6532);
nand NAND3 (N6540, N6503, N1571, N4641);
nand NAND4 (N6541, N6537, N6526, N4008, N5868);
nor NOR2 (N6542, N6535, N475);
nand NAND3 (N6543, N6539, N4265, N68);
and AND2 (N6544, N6542, N3965);
not NOT1 (N6545, N6543);
and AND3 (N6546, N6533, N3822, N5720);
nor NOR4 (N6547, N6538, N1156, N459, N5008);
not NOT1 (N6548, N6524);
and AND4 (N6549, N6548, N3443, N3980, N4853);
nand NAND4 (N6550, N6547, N2170, N1298, N1327);
nor NOR2 (N6551, N6540, N6092);
xor XOR2 (N6552, N6550, N5630);
buf BUF1 (N6553, N6544);
or OR3 (N6554, N6552, N499, N350);
and AND2 (N6555, N6541, N4924);
nand NAND3 (N6556, N6519, N5142, N780);
nor NOR2 (N6557, N6529, N5070);
buf BUF1 (N6558, N6536);
nor NOR2 (N6559, N6554, N6137);
nand NAND3 (N6560, N6551, N3028, N824);
or OR4 (N6561, N6555, N5869, N3143, N4695);
not NOT1 (N6562, N6558);
nand NAND2 (N6563, N6562, N3316);
nand NAND4 (N6564, N6549, N945, N5642, N3454);
xor XOR2 (N6565, N6553, N6233);
xor XOR2 (N6566, N6556, N2665);
or OR4 (N6567, N6559, N5789, N5701, N6169);
nor NOR2 (N6568, N6561, N5307);
or OR4 (N6569, N6565, N4389, N1185, N1026);
and AND2 (N6570, N6563, N829);
xor XOR2 (N6571, N6564, N5757);
and AND3 (N6572, N6560, N5843, N2416);
or OR3 (N6573, N6545, N5635, N2168);
and AND4 (N6574, N6557, N677, N3222, N2377);
or OR3 (N6575, N6566, N6043, N4246);
buf BUF1 (N6576, N6573);
nor NOR3 (N6577, N6575, N2332, N3403);
or OR3 (N6578, N6569, N3753, N5432);
xor XOR2 (N6579, N6567, N441);
or OR4 (N6580, N6577, N3658, N6243, N4715);
and AND4 (N6581, N6570, N2917, N6203, N4792);
not NOT1 (N6582, N6546);
or OR3 (N6583, N6576, N67, N1846);
and AND4 (N6584, N6579, N6426, N3709, N710);
nor NOR3 (N6585, N6568, N3169, N5327);
nand NAND3 (N6586, N6583, N2858, N2728);
not NOT1 (N6587, N6572);
nor NOR3 (N6588, N6578, N5971, N4079);
not NOT1 (N6589, N6587);
nand NAND2 (N6590, N6580, N2613);
buf BUF1 (N6591, N6581);
or OR3 (N6592, N6589, N6471, N5129);
and AND2 (N6593, N6590, N3538);
xor XOR2 (N6594, N6582, N299);
nand NAND4 (N6595, N6586, N6203, N4658, N3206);
or OR4 (N6596, N6595, N3118, N490, N3135);
not NOT1 (N6597, N6571);
nor NOR3 (N6598, N6597, N3422, N2222);
buf BUF1 (N6599, N6596);
buf BUF1 (N6600, N6584);
not NOT1 (N6601, N6591);
nor NOR4 (N6602, N6599, N3098, N6480, N2492);
or OR4 (N6603, N6574, N4305, N1023, N1766);
or OR3 (N6604, N6600, N6527, N989);
nand NAND3 (N6605, N6604, N547, N4193);
not NOT1 (N6606, N6605);
nand NAND4 (N6607, N6606, N6076, N5784, N3224);
not NOT1 (N6608, N6588);
nor NOR4 (N6609, N6598, N1229, N280, N5472);
or OR4 (N6610, N6593, N2047, N4853, N4677);
xor XOR2 (N6611, N6592, N1616);
nor NOR4 (N6612, N6609, N5061, N3503, N3065);
buf BUF1 (N6613, N6585);
nand NAND3 (N6614, N6611, N3068, N6155);
buf BUF1 (N6615, N6603);
nor NOR2 (N6616, N6594, N2778);
nor NOR2 (N6617, N6601, N604);
or OR2 (N6618, N6608, N5916);
and AND2 (N6619, N6616, N2116);
buf BUF1 (N6620, N6612);
buf BUF1 (N6621, N6620);
and AND3 (N6622, N6610, N3398, N1478);
not NOT1 (N6623, N6618);
or OR4 (N6624, N6613, N3116, N849, N5477);
or OR3 (N6625, N6607, N4847, N3911);
buf BUF1 (N6626, N6615);
and AND2 (N6627, N6626, N3724);
or OR3 (N6628, N6614, N1113, N903);
nand NAND3 (N6629, N6602, N3893, N46);
buf BUF1 (N6630, N6627);
buf BUF1 (N6631, N6624);
not NOT1 (N6632, N6625);
or OR2 (N6633, N6622, N1281);
nor NOR4 (N6634, N6630, N2259, N1083, N4701);
xor XOR2 (N6635, N6629, N1223);
buf BUF1 (N6636, N6633);
or OR4 (N6637, N6636, N5265, N2654, N4016);
nand NAND3 (N6638, N6637, N4550, N4177);
buf BUF1 (N6639, N6631);
xor XOR2 (N6640, N6621, N317);
and AND3 (N6641, N6640, N1954, N1406);
nand NAND4 (N6642, N6638, N5006, N2324, N2133);
buf BUF1 (N6643, N6641);
nor NOR2 (N6644, N6623, N5889);
nor NOR4 (N6645, N6642, N6524, N753, N2612);
buf BUF1 (N6646, N6619);
nor NOR3 (N6647, N6632, N27, N5024);
or OR4 (N6648, N6646, N3661, N2169, N544);
or OR2 (N6649, N6644, N189);
nor NOR2 (N6650, N6649, N3509);
buf BUF1 (N6651, N6634);
not NOT1 (N6652, N6635);
and AND3 (N6653, N6645, N6415, N6254);
or OR3 (N6654, N6639, N4633, N6051);
and AND3 (N6655, N6647, N4602, N6251);
buf BUF1 (N6656, N6648);
not NOT1 (N6657, N6650);
nand NAND3 (N6658, N6654, N5151, N5548);
nor NOR3 (N6659, N6643, N4946, N3554);
and AND4 (N6660, N6658, N283, N5568, N114);
buf BUF1 (N6661, N6656);
buf BUF1 (N6662, N6617);
nand NAND3 (N6663, N6628, N6073, N4765);
nand NAND3 (N6664, N6653, N6101, N1042);
and AND3 (N6665, N6651, N5454, N1087);
and AND4 (N6666, N6659, N6031, N365, N4515);
and AND2 (N6667, N6655, N663);
buf BUF1 (N6668, N6663);
buf BUF1 (N6669, N6668);
nand NAND3 (N6670, N6662, N726, N1233);
buf BUF1 (N6671, N6657);
nand NAND2 (N6672, N6652, N2835);
not NOT1 (N6673, N6666);
nand NAND2 (N6674, N6667, N3793);
and AND3 (N6675, N6673, N5590, N959);
buf BUF1 (N6676, N6661);
nand NAND2 (N6677, N6670, N685);
xor XOR2 (N6678, N6671, N4407);
and AND2 (N6679, N6677, N1544);
nand NAND2 (N6680, N6665, N284);
and AND2 (N6681, N6675, N6556);
nor NOR4 (N6682, N6676, N5393, N4075, N1948);
or OR4 (N6683, N6678, N5117, N3737, N6220);
and AND3 (N6684, N6672, N379, N2240);
nand NAND2 (N6685, N6684, N1492);
xor XOR2 (N6686, N6683, N6639);
or OR2 (N6687, N6669, N2027);
or OR3 (N6688, N6680, N3159, N6598);
buf BUF1 (N6689, N6674);
nor NOR4 (N6690, N6664, N4207, N3818, N2832);
or OR3 (N6691, N6685, N5430, N3750);
nand NAND3 (N6692, N6681, N275, N3316);
nor NOR4 (N6693, N6660, N1660, N6052, N1664);
nand NAND2 (N6694, N6690, N2337);
and AND3 (N6695, N6679, N1941, N6031);
not NOT1 (N6696, N6686);
and AND3 (N6697, N6689, N6487, N2109);
nand NAND3 (N6698, N6682, N2164, N5467);
and AND4 (N6699, N6687, N992, N4697, N2576);
or OR4 (N6700, N6696, N5457, N2394, N2992);
and AND3 (N6701, N6691, N5802, N6324);
not NOT1 (N6702, N6693);
nor NOR4 (N6703, N6695, N1727, N4410, N3761);
buf BUF1 (N6704, N6702);
nor NOR2 (N6705, N6697, N6366);
nor NOR2 (N6706, N6701, N631);
and AND2 (N6707, N6699, N3465);
xor XOR2 (N6708, N6703, N1533);
not NOT1 (N6709, N6705);
and AND4 (N6710, N6688, N3994, N3625, N2195);
nor NOR2 (N6711, N6704, N2900);
buf BUF1 (N6712, N6710);
not NOT1 (N6713, N6707);
xor XOR2 (N6714, N6692, N2058);
nor NOR2 (N6715, N6712, N3986);
buf BUF1 (N6716, N6698);
or OR2 (N6717, N6714, N2288);
and AND3 (N6718, N6694, N3564, N6075);
xor XOR2 (N6719, N6709, N1621);
not NOT1 (N6720, N6711);
buf BUF1 (N6721, N6715);
or OR3 (N6722, N6716, N6620, N3116);
buf BUF1 (N6723, N6722);
not NOT1 (N6724, N6720);
nand NAND3 (N6725, N6718, N4253, N4491);
and AND4 (N6726, N6724, N4456, N6375, N2685);
not NOT1 (N6727, N6723);
xor XOR2 (N6728, N6727, N2888);
not NOT1 (N6729, N6717);
xor XOR2 (N6730, N6729, N419);
or OR4 (N6731, N6725, N168, N1507, N6501);
xor XOR2 (N6732, N6708, N1272);
nand NAND2 (N6733, N6732, N3438);
nor NOR3 (N6734, N6726, N6184, N4721);
and AND3 (N6735, N6730, N4180, N1297);
nor NOR4 (N6736, N6734, N4975, N5257, N2231);
xor XOR2 (N6737, N6733, N6643);
and AND4 (N6738, N6713, N4167, N357, N2954);
and AND3 (N6739, N6706, N1233, N6283);
or OR4 (N6740, N6719, N5901, N646, N2844);
or OR4 (N6741, N6721, N1050, N4630, N2281);
or OR3 (N6742, N6740, N4602, N1499);
not NOT1 (N6743, N6735);
buf BUF1 (N6744, N6728);
nor NOR2 (N6745, N6743, N5824);
nand NAND2 (N6746, N6745, N1967);
not NOT1 (N6747, N6731);
nor NOR2 (N6748, N6742, N1216);
or OR3 (N6749, N6737, N436, N6673);
nand NAND3 (N6750, N6746, N508, N5107);
or OR2 (N6751, N6741, N2862);
nand NAND3 (N6752, N6739, N3149, N4844);
buf BUF1 (N6753, N6751);
and AND3 (N6754, N6750, N1847, N613);
xor XOR2 (N6755, N6748, N4098);
and AND3 (N6756, N6747, N4663, N3273);
and AND2 (N6757, N6744, N3874);
or OR2 (N6758, N6749, N3095);
or OR3 (N6759, N6755, N1978, N471);
or OR4 (N6760, N6756, N3887, N6272, N6222);
or OR2 (N6761, N6757, N5292);
nor NOR2 (N6762, N6752, N3308);
nand NAND4 (N6763, N6736, N3257, N1798, N2806);
and AND4 (N6764, N6760, N3250, N1068, N1285);
xor XOR2 (N6765, N6761, N301);
nand NAND2 (N6766, N6753, N661);
nand NAND3 (N6767, N6758, N3058, N1070);
nor NOR2 (N6768, N6765, N2852);
xor XOR2 (N6769, N6738, N95);
xor XOR2 (N6770, N6767, N26);
not NOT1 (N6771, N6766);
nor NOR3 (N6772, N6771, N163, N351);
and AND3 (N6773, N6763, N2239, N3434);
buf BUF1 (N6774, N6769);
not NOT1 (N6775, N6773);
buf BUF1 (N6776, N6700);
not NOT1 (N6777, N6774);
nor NOR3 (N6778, N6762, N2665, N763);
buf BUF1 (N6779, N6778);
nor NOR2 (N6780, N6754, N461);
nor NOR4 (N6781, N6759, N6680, N1999, N6091);
or OR2 (N6782, N6768, N1306);
and AND3 (N6783, N6779, N4653, N5841);
nand NAND3 (N6784, N6783, N3196, N6562);
nand NAND3 (N6785, N6784, N873, N1265);
and AND2 (N6786, N6777, N2572);
or OR2 (N6787, N6775, N4977);
and AND2 (N6788, N6781, N2835);
buf BUF1 (N6789, N6786);
not NOT1 (N6790, N6788);
xor XOR2 (N6791, N6782, N2207);
or OR3 (N6792, N6764, N671, N4919);
or OR2 (N6793, N6791, N3048);
or OR2 (N6794, N6776, N450);
xor XOR2 (N6795, N6789, N4779);
xor XOR2 (N6796, N6793, N3944);
buf BUF1 (N6797, N6790);
nand NAND3 (N6798, N6796, N1577, N4731);
nand NAND4 (N6799, N6772, N484, N2638, N3797);
xor XOR2 (N6800, N6787, N6715);
nor NOR3 (N6801, N6799, N3245, N2649);
nor NOR2 (N6802, N6785, N4503);
xor XOR2 (N6803, N6770, N2682);
buf BUF1 (N6804, N6803);
nand NAND3 (N6805, N6800, N6348, N1830);
buf BUF1 (N6806, N6780);
or OR4 (N6807, N6794, N1887, N1624, N5685);
and AND3 (N6808, N6804, N1838, N4844);
nand NAND2 (N6809, N6795, N786);
nor NOR4 (N6810, N6809, N6071, N5698, N1067);
not NOT1 (N6811, N6802);
not NOT1 (N6812, N6810);
and AND3 (N6813, N6792, N2746, N3133);
not NOT1 (N6814, N6806);
and AND4 (N6815, N6801, N3768, N4606, N3774);
and AND3 (N6816, N6814, N3510, N1604);
xor XOR2 (N6817, N6813, N1782);
nor NOR3 (N6818, N6807, N4883, N1079);
or OR4 (N6819, N6808, N2332, N5538, N4446);
nand NAND4 (N6820, N6811, N1960, N6097, N2817);
and AND2 (N6821, N6819, N4855);
xor XOR2 (N6822, N6816, N396);
xor XOR2 (N6823, N6821, N1973);
not NOT1 (N6824, N6798);
and AND3 (N6825, N6817, N5987, N1646);
or OR2 (N6826, N6824, N4829);
not NOT1 (N6827, N6826);
or OR2 (N6828, N6827, N98);
buf BUF1 (N6829, N6820);
buf BUF1 (N6830, N6805);
nor NOR3 (N6831, N6830, N5940, N4118);
nand NAND3 (N6832, N6828, N143, N4215);
nor NOR2 (N6833, N6825, N5974);
nor NOR3 (N6834, N6831, N746, N1863);
and AND4 (N6835, N6822, N2697, N6029, N6359);
not NOT1 (N6836, N6818);
nand NAND2 (N6837, N6812, N5460);
and AND2 (N6838, N6836, N4154);
or OR4 (N6839, N6823, N6567, N1565, N5167);
or OR2 (N6840, N6839, N460);
or OR2 (N6841, N6832, N6075);
not NOT1 (N6842, N6834);
xor XOR2 (N6843, N6797, N6829);
xor XOR2 (N6844, N6133, N3836);
not NOT1 (N6845, N6841);
nor NOR2 (N6846, N6843, N6523);
nand NAND4 (N6847, N6842, N1663, N3228, N987);
xor XOR2 (N6848, N6815, N6298);
and AND4 (N6849, N6847, N1136, N3550, N771);
nor NOR4 (N6850, N6848, N4075, N2838, N477);
buf BUF1 (N6851, N6845);
xor XOR2 (N6852, N6844, N2048);
nor NOR3 (N6853, N6838, N2277, N4444);
xor XOR2 (N6854, N6846, N4126);
nor NOR3 (N6855, N6849, N2029, N4554);
not NOT1 (N6856, N6850);
nand NAND2 (N6857, N6855, N769);
xor XOR2 (N6858, N6854, N5838);
or OR4 (N6859, N6853, N219, N1807, N1628);
xor XOR2 (N6860, N6856, N2155);
or OR3 (N6861, N6833, N2277, N384);
or OR3 (N6862, N6857, N6245, N6533);
nor NOR4 (N6863, N6851, N5686, N3229, N5647);
nand NAND4 (N6864, N6840, N338, N5147, N2541);
not NOT1 (N6865, N6864);
or OR2 (N6866, N6852, N4814);
buf BUF1 (N6867, N6865);
and AND4 (N6868, N6866, N569, N202, N1930);
xor XOR2 (N6869, N6837, N754);
nor NOR3 (N6870, N6861, N2289, N3112);
or OR2 (N6871, N6835, N2573);
xor XOR2 (N6872, N6859, N1460);
nand NAND3 (N6873, N6870, N550, N2581);
xor XOR2 (N6874, N6869, N6149);
buf BUF1 (N6875, N6868);
and AND3 (N6876, N6862, N5139, N3108);
buf BUF1 (N6877, N6873);
buf BUF1 (N6878, N6877);
not NOT1 (N6879, N6860);
buf BUF1 (N6880, N6876);
nor NOR3 (N6881, N6858, N1482, N3270);
xor XOR2 (N6882, N6879, N1470);
nor NOR3 (N6883, N6880, N2535, N4665);
not NOT1 (N6884, N6883);
and AND2 (N6885, N6878, N1573);
and AND2 (N6886, N6874, N278);
nand NAND4 (N6887, N6867, N215, N1343, N1976);
xor XOR2 (N6888, N6872, N2694);
nor NOR3 (N6889, N6875, N6725, N6392);
nand NAND4 (N6890, N6871, N4151, N440, N6467);
nand NAND2 (N6891, N6889, N4665);
and AND3 (N6892, N6886, N5711, N1250);
nor NOR2 (N6893, N6885, N3869);
nor NOR4 (N6894, N6882, N5971, N3576, N2942);
buf BUF1 (N6895, N6891);
xor XOR2 (N6896, N6890, N5619);
xor XOR2 (N6897, N6888, N5169);
not NOT1 (N6898, N6892);
nor NOR3 (N6899, N6887, N6372, N2124);
buf BUF1 (N6900, N6897);
nand NAND4 (N6901, N6899, N536, N1557, N5336);
buf BUF1 (N6902, N6901);
or OR3 (N6903, N6895, N4460, N2334);
buf BUF1 (N6904, N6903);
nor NOR4 (N6905, N6902, N947, N3978, N551);
or OR2 (N6906, N6893, N2396);
nor NOR4 (N6907, N6863, N2750, N2388, N3914);
and AND3 (N6908, N6896, N2737, N3991);
or OR4 (N6909, N6884, N1500, N938, N3197);
buf BUF1 (N6910, N6909);
xor XOR2 (N6911, N6908, N2973);
buf BUF1 (N6912, N6910);
nand NAND4 (N6913, N6912, N3247, N478, N2608);
or OR4 (N6914, N6906, N6116, N5695, N627);
nand NAND3 (N6915, N6894, N3508, N4964);
nor NOR4 (N6916, N6914, N1720, N5548, N4086);
not NOT1 (N6917, N6913);
nor NOR2 (N6918, N6905, N2529);
and AND2 (N6919, N6898, N708);
xor XOR2 (N6920, N6900, N1798);
buf BUF1 (N6921, N6881);
buf BUF1 (N6922, N6917);
and AND3 (N6923, N6922, N1942, N5876);
buf BUF1 (N6924, N6921);
nand NAND4 (N6925, N6916, N6160, N3935, N3756);
or OR3 (N6926, N6920, N1337, N6722);
not NOT1 (N6927, N6925);
and AND2 (N6928, N6919, N5734);
not NOT1 (N6929, N6904);
buf BUF1 (N6930, N6924);
nand NAND4 (N6931, N6928, N5716, N6013, N1184);
nor NOR4 (N6932, N6918, N263, N1354, N5449);
or OR3 (N6933, N6923, N4573, N18);
nor NOR2 (N6934, N6911, N6579);
and AND4 (N6935, N6934, N6450, N2887, N2907);
buf BUF1 (N6936, N6927);
not NOT1 (N6937, N6930);
not NOT1 (N6938, N6907);
buf BUF1 (N6939, N6933);
xor XOR2 (N6940, N6915, N1179);
and AND2 (N6941, N6926, N4673);
not NOT1 (N6942, N6941);
not NOT1 (N6943, N6939);
and AND4 (N6944, N6932, N5331, N4013, N4084);
nor NOR2 (N6945, N6940, N2653);
xor XOR2 (N6946, N6943, N2914);
and AND4 (N6947, N6931, N4458, N2489, N5296);
nor NOR4 (N6948, N6937, N6028, N2637, N6224);
xor XOR2 (N6949, N6942, N3355);
buf BUF1 (N6950, N6948);
nor NOR3 (N6951, N6938, N3536, N6566);
and AND3 (N6952, N6945, N3876, N4972);
xor XOR2 (N6953, N6950, N5960);
buf BUF1 (N6954, N6953);
nand NAND4 (N6955, N6944, N553, N6404, N1948);
nor NOR2 (N6956, N6947, N5058);
nor NOR3 (N6957, N6956, N4188, N2029);
nand NAND2 (N6958, N6935, N2609);
or OR4 (N6959, N6946, N4338, N4038, N5806);
nand NAND4 (N6960, N6936, N3654, N5481, N1787);
or OR3 (N6961, N6929, N553, N5539);
xor XOR2 (N6962, N6955, N3293);
nor NOR3 (N6963, N6960, N3409, N2509);
nor NOR3 (N6964, N6959, N6076, N6417);
or OR2 (N6965, N6952, N1117);
not NOT1 (N6966, N6949);
or OR2 (N6967, N6957, N4822);
and AND3 (N6968, N6967, N6946, N3893);
and AND4 (N6969, N6964, N1686, N989, N3726);
nor NOR4 (N6970, N6963, N109, N1988, N516);
buf BUF1 (N6971, N6965);
xor XOR2 (N6972, N6966, N2278);
buf BUF1 (N6973, N6961);
and AND3 (N6974, N6958, N1067, N1702);
nor NOR3 (N6975, N6974, N365, N424);
and AND4 (N6976, N6969, N3981, N5465, N1661);
or OR4 (N6977, N6962, N279, N6433, N5693);
not NOT1 (N6978, N6972);
or OR2 (N6979, N6978, N3025);
xor XOR2 (N6980, N6954, N3987);
nand NAND2 (N6981, N6977, N3025);
nand NAND2 (N6982, N6968, N1689);
or OR3 (N6983, N6970, N4622, N4390);
and AND2 (N6984, N6981, N4381);
xor XOR2 (N6985, N6984, N3533);
nor NOR2 (N6986, N6982, N6973);
nor NOR2 (N6987, N6226, N3583);
nand NAND2 (N6988, N6987, N3194);
nand NAND4 (N6989, N6988, N1750, N862, N4134);
nor NOR3 (N6990, N6989, N2935, N6275);
and AND3 (N6991, N6980, N4403, N3088);
xor XOR2 (N6992, N6975, N677);
and AND4 (N6993, N6990, N4692, N6524, N4782);
nor NOR2 (N6994, N6993, N2326);
xor XOR2 (N6995, N6976, N929);
nand NAND2 (N6996, N6971, N3227);
not NOT1 (N6997, N6983);
or OR3 (N6998, N6951, N6489, N5149);
not NOT1 (N6999, N6995);
buf BUF1 (N7000, N6999);
nor NOR2 (N7001, N6992, N6410);
nand NAND3 (N7002, N6997, N471, N2168);
not NOT1 (N7003, N6994);
or OR2 (N7004, N7000, N2726);
or OR2 (N7005, N7003, N1390);
nor NOR4 (N7006, N6998, N6051, N97, N2124);
or OR2 (N7007, N6979, N3910);
nand NAND4 (N7008, N6986, N734, N5636, N3607);
nand NAND3 (N7009, N7004, N5472, N29);
buf BUF1 (N7010, N6985);
or OR4 (N7011, N7007, N3419, N3852, N2181);
xor XOR2 (N7012, N6991, N757);
xor XOR2 (N7013, N7009, N5374);
nor NOR4 (N7014, N7005, N1047, N1984, N6050);
nor NOR2 (N7015, N7013, N833);
and AND4 (N7016, N7012, N222, N1434, N3699);
and AND4 (N7017, N7014, N2160, N5468, N4147);
and AND4 (N7018, N7010, N5300, N5731, N2040);
and AND4 (N7019, N7006, N6325, N5923, N3163);
and AND4 (N7020, N7008, N3670, N2310, N561);
and AND4 (N7021, N6996, N289, N1755, N5668);
not NOT1 (N7022, N7017);
and AND2 (N7023, N7002, N4857);
and AND4 (N7024, N7011, N1064, N3870, N7010);
nor NOR3 (N7025, N7016, N6819, N6809);
nand NAND3 (N7026, N7021, N2189, N5782);
or OR2 (N7027, N7019, N6335);
buf BUF1 (N7028, N7015);
nor NOR2 (N7029, N7018, N3231);
or OR3 (N7030, N7020, N3263, N2730);
not NOT1 (N7031, N7022);
nand NAND4 (N7032, N7001, N1236, N1617, N2542);
or OR3 (N7033, N7030, N6712, N2253);
nand NAND2 (N7034, N7025, N4858);
not NOT1 (N7035, N7033);
xor XOR2 (N7036, N7024, N4885);
not NOT1 (N7037, N7031);
and AND3 (N7038, N7023, N2600, N3016);
buf BUF1 (N7039, N7038);
nor NOR4 (N7040, N7037, N3850, N6365, N5152);
nand NAND2 (N7041, N7026, N4188);
buf BUF1 (N7042, N7034);
xor XOR2 (N7043, N7039, N239);
nor NOR4 (N7044, N7035, N6104, N2381, N2102);
not NOT1 (N7045, N7041);
nand NAND2 (N7046, N7027, N1918);
or OR2 (N7047, N7029, N4128);
buf BUF1 (N7048, N7040);
and AND4 (N7049, N7046, N491, N3450, N462);
not NOT1 (N7050, N7047);
nand NAND3 (N7051, N7032, N5424, N6203);
nor NOR4 (N7052, N7048, N4379, N1074, N4472);
not NOT1 (N7053, N7028);
or OR2 (N7054, N7042, N1423);
not NOT1 (N7055, N7051);
or OR4 (N7056, N7045, N3764, N3231, N6632);
buf BUF1 (N7057, N7056);
not NOT1 (N7058, N7043);
or OR4 (N7059, N7036, N4285, N1796, N6825);
nor NOR2 (N7060, N7057, N5855);
or OR3 (N7061, N7044, N2015, N3854);
not NOT1 (N7062, N7052);
buf BUF1 (N7063, N7062);
nor NOR3 (N7064, N7058, N152, N6999);
or OR4 (N7065, N7063, N5611, N3455, N1461);
xor XOR2 (N7066, N7065, N1177);
and AND2 (N7067, N7059, N4510);
xor XOR2 (N7068, N7067, N5415);
nand NAND2 (N7069, N7068, N689);
nor NOR3 (N7070, N7064, N4360, N3830);
xor XOR2 (N7071, N7061, N6207);
not NOT1 (N7072, N7069);
buf BUF1 (N7073, N7071);
or OR4 (N7074, N7066, N5963, N2268, N4376);
not NOT1 (N7075, N7050);
nand NAND3 (N7076, N7060, N167, N4110);
not NOT1 (N7077, N7076);
buf BUF1 (N7078, N7054);
or OR3 (N7079, N7074, N1009, N875);
or OR3 (N7080, N7053, N6164, N2866);
and AND3 (N7081, N7072, N4749, N3375);
nor NOR3 (N7082, N7070, N668, N1024);
and AND4 (N7083, N7079, N4436, N2829, N3704);
and AND2 (N7084, N7081, N2967);
nand NAND2 (N7085, N7073, N2563);
or OR3 (N7086, N7049, N3049, N6974);
nor NOR4 (N7087, N7078, N2889, N3705, N2446);
nor NOR3 (N7088, N7082, N3030, N3905);
xor XOR2 (N7089, N7080, N3370);
and AND2 (N7090, N7083, N5398);
xor XOR2 (N7091, N7085, N530);
not NOT1 (N7092, N7090);
xor XOR2 (N7093, N7089, N3931);
nand NAND4 (N7094, N7088, N4201, N1720, N6145);
and AND4 (N7095, N7094, N2008, N5603, N5421);
or OR3 (N7096, N7092, N5387, N1274);
or OR3 (N7097, N7086, N5336, N1295);
nand NAND3 (N7098, N7084, N1482, N992);
and AND2 (N7099, N7098, N2247);
not NOT1 (N7100, N7075);
xor XOR2 (N7101, N7099, N670);
nand NAND3 (N7102, N7077, N270, N5494);
and AND2 (N7103, N7101, N6755);
xor XOR2 (N7104, N7091, N4683);
xor XOR2 (N7105, N7103, N519);
xor XOR2 (N7106, N7095, N894);
buf BUF1 (N7107, N7106);
and AND4 (N7108, N7096, N6940, N3543, N2037);
xor XOR2 (N7109, N7105, N1785);
or OR3 (N7110, N7087, N372, N2160);
nor NOR3 (N7111, N7093, N3056, N2114);
and AND3 (N7112, N7100, N813, N6363);
or OR2 (N7113, N7112, N6115);
buf BUF1 (N7114, N7111);
nand NAND4 (N7115, N7109, N2113, N1094, N359);
not NOT1 (N7116, N7113);
nand NAND2 (N7117, N7115, N2618);
nor NOR2 (N7118, N7107, N2801);
nand NAND4 (N7119, N7116, N3900, N3390, N3354);
nor NOR4 (N7120, N7055, N5212, N4134, N880);
or OR2 (N7121, N7102, N6922);
not NOT1 (N7122, N7117);
xor XOR2 (N7123, N7104, N5411);
not NOT1 (N7124, N7118);
not NOT1 (N7125, N7122);
nand NAND2 (N7126, N7097, N3938);
xor XOR2 (N7127, N7119, N1966);
nand NAND2 (N7128, N7123, N5476);
not NOT1 (N7129, N7124);
nand NAND2 (N7130, N7127, N4298);
nand NAND2 (N7131, N7126, N2240);
xor XOR2 (N7132, N7131, N3853);
and AND2 (N7133, N7120, N4310);
xor XOR2 (N7134, N7133, N2204);
xor XOR2 (N7135, N7128, N1996);
xor XOR2 (N7136, N7121, N2147);
or OR3 (N7137, N7136, N172, N6630);
or OR3 (N7138, N7134, N2122, N3461);
or OR4 (N7139, N7137, N1606, N4530, N1023);
nor NOR2 (N7140, N7108, N2287);
nand NAND3 (N7141, N7132, N911, N5476);
or OR4 (N7142, N7138, N572, N174, N5794);
nand NAND2 (N7143, N7129, N4831);
buf BUF1 (N7144, N7140);
xor XOR2 (N7145, N7114, N3222);
nand NAND3 (N7146, N7145, N6646, N4494);
nor NOR3 (N7147, N7135, N326, N788);
and AND2 (N7148, N7142, N1549);
nand NAND3 (N7149, N7141, N3560, N5484);
or OR3 (N7150, N7125, N468, N5995);
xor XOR2 (N7151, N7149, N1748);
or OR4 (N7152, N7148, N2076, N2455, N4110);
nor NOR4 (N7153, N7110, N3605, N481, N4821);
nor NOR3 (N7154, N7147, N6522, N4534);
nor NOR3 (N7155, N7154, N4549, N4863);
or OR3 (N7156, N7151, N2465, N2589);
and AND2 (N7157, N7150, N5278);
or OR3 (N7158, N7144, N6558, N3374);
buf BUF1 (N7159, N7143);
or OR3 (N7160, N7130, N5923, N6133);
buf BUF1 (N7161, N7139);
nand NAND4 (N7162, N7152, N2374, N1635, N6381);
not NOT1 (N7163, N7146);
xor XOR2 (N7164, N7153, N4667);
nor NOR2 (N7165, N7157, N5365);
buf BUF1 (N7166, N7156);
and AND3 (N7167, N7155, N388, N6185);
or OR2 (N7168, N7158, N3480);
nor NOR4 (N7169, N7168, N4531, N112, N6183);
buf BUF1 (N7170, N7165);
and AND4 (N7171, N7170, N932, N398, N197);
and AND4 (N7172, N7159, N2780, N5162, N4008);
xor XOR2 (N7173, N7171, N3514);
and AND3 (N7174, N7161, N4411, N1825);
buf BUF1 (N7175, N7174);
not NOT1 (N7176, N7162);
nor NOR2 (N7177, N7167, N5232);
buf BUF1 (N7178, N7177);
buf BUF1 (N7179, N7160);
or OR4 (N7180, N7179, N2317, N6123, N6748);
or OR3 (N7181, N7173, N2626, N3579);
not NOT1 (N7182, N7176);
and AND3 (N7183, N7164, N3082, N2529);
nor NOR4 (N7184, N7172, N3869, N4987, N3609);
not NOT1 (N7185, N7182);
not NOT1 (N7186, N7183);
or OR2 (N7187, N7180, N428);
buf BUF1 (N7188, N7166);
nand NAND4 (N7189, N7184, N2475, N2373, N2729);
nand NAND3 (N7190, N7188, N1475, N3824);
or OR4 (N7191, N7189, N3051, N1559, N6456);
and AND2 (N7192, N7175, N3727);
not NOT1 (N7193, N7186);
or OR3 (N7194, N7187, N5627, N2462);
nand NAND4 (N7195, N7163, N2202, N6957, N6400);
buf BUF1 (N7196, N7181);
buf BUF1 (N7197, N7194);
nor NOR3 (N7198, N7178, N1306, N1083);
nand NAND3 (N7199, N7190, N6433, N2829);
xor XOR2 (N7200, N7185, N5730);
nor NOR4 (N7201, N7192, N2273, N3110, N6248);
not NOT1 (N7202, N7191);
nand NAND2 (N7203, N7199, N3459);
and AND3 (N7204, N7195, N2556, N4778);
xor XOR2 (N7205, N7203, N1425);
and AND3 (N7206, N7200, N3015, N3387);
xor XOR2 (N7207, N7205, N4645);
or OR3 (N7208, N7198, N1325, N6370);
and AND4 (N7209, N7204, N6163, N5232, N1517);
nand NAND3 (N7210, N7202, N6100, N6980);
nor NOR4 (N7211, N7193, N1846, N5749, N4307);
xor XOR2 (N7212, N7169, N6182);
or OR3 (N7213, N7207, N3331, N6562);
and AND3 (N7214, N7208, N1450, N4313);
and AND2 (N7215, N7210, N5858);
not NOT1 (N7216, N7196);
nor NOR2 (N7217, N7211, N2470);
nand NAND4 (N7218, N7214, N3356, N1690, N2292);
nor NOR3 (N7219, N7216, N919, N2126);
and AND2 (N7220, N7217, N328);
xor XOR2 (N7221, N7219, N3220);
xor XOR2 (N7222, N7220, N4152);
not NOT1 (N7223, N7218);
and AND3 (N7224, N7212, N1949, N5341);
or OR3 (N7225, N7223, N3385, N7219);
not NOT1 (N7226, N7213);
nand NAND2 (N7227, N7206, N7163);
buf BUF1 (N7228, N7197);
nand NAND2 (N7229, N7222, N3433);
nor NOR4 (N7230, N7226, N3709, N4381, N2015);
buf BUF1 (N7231, N7215);
xor XOR2 (N7232, N7231, N6368);
xor XOR2 (N7233, N7230, N6842);
or OR4 (N7234, N7224, N682, N3346, N4625);
buf BUF1 (N7235, N7234);
or OR4 (N7236, N7225, N2317, N4088, N2140);
and AND2 (N7237, N7221, N5475);
not NOT1 (N7238, N7232);
not NOT1 (N7239, N7227);
nand NAND2 (N7240, N7201, N6830);
or OR4 (N7241, N7236, N5338, N3185, N1427);
and AND3 (N7242, N7240, N6036, N4173);
nand NAND4 (N7243, N7241, N3339, N2183, N3259);
xor XOR2 (N7244, N7229, N281);
not NOT1 (N7245, N7228);
not NOT1 (N7246, N7245);
nor NOR2 (N7247, N7242, N6801);
nand NAND4 (N7248, N7244, N6611, N3063, N4671);
buf BUF1 (N7249, N7237);
nand NAND4 (N7250, N7238, N6187, N6760, N2233);
not NOT1 (N7251, N7243);
buf BUF1 (N7252, N7209);
and AND4 (N7253, N7249, N2794, N5777, N2837);
nor NOR2 (N7254, N7252, N1717);
and AND3 (N7255, N7254, N149, N3314);
and AND4 (N7256, N7247, N2379, N222, N3980);
xor XOR2 (N7257, N7239, N5769);
or OR4 (N7258, N7256, N5167, N5536, N2311);
xor XOR2 (N7259, N7251, N2982);
or OR3 (N7260, N7253, N4080, N5031);
nand NAND2 (N7261, N7257, N3269);
or OR4 (N7262, N7250, N3882, N6209, N4289);
not NOT1 (N7263, N7255);
nand NAND3 (N7264, N7263, N6551, N3774);
not NOT1 (N7265, N7235);
buf BUF1 (N7266, N7264);
nand NAND2 (N7267, N7233, N2541);
not NOT1 (N7268, N7265);
and AND3 (N7269, N7262, N6330, N6258);
or OR4 (N7270, N7259, N4050, N176, N6269);
nand NAND2 (N7271, N7258, N6234);
and AND3 (N7272, N7246, N910, N5610);
nor NOR4 (N7273, N7267, N5508, N1387, N6423);
nand NAND4 (N7274, N7268, N2120, N2128, N4861);
nand NAND4 (N7275, N7266, N7257, N2416, N2871);
buf BUF1 (N7276, N7270);
buf BUF1 (N7277, N7272);
nand NAND4 (N7278, N7260, N1685, N2092, N7083);
not NOT1 (N7279, N7273);
nor NOR2 (N7280, N7261, N5366);
and AND2 (N7281, N7248, N4801);
buf BUF1 (N7282, N7280);
and AND2 (N7283, N7271, N2047);
and AND4 (N7284, N7275, N4893, N2060, N3722);
nand NAND4 (N7285, N7281, N3362, N6828, N3457);
not NOT1 (N7286, N7276);
and AND3 (N7287, N7286, N5963, N3109);
buf BUF1 (N7288, N7279);
and AND2 (N7289, N7288, N3952);
nand NAND3 (N7290, N7282, N3691, N7078);
xor XOR2 (N7291, N7285, N3265);
nand NAND3 (N7292, N7269, N4483, N1112);
xor XOR2 (N7293, N7290, N5853);
nor NOR4 (N7294, N7287, N7264, N7109, N1063);
not NOT1 (N7295, N7277);
or OR2 (N7296, N7274, N2898);
or OR4 (N7297, N7294, N6567, N6369, N5073);
buf BUF1 (N7298, N7292);
or OR3 (N7299, N7298, N245, N1523);
not NOT1 (N7300, N7284);
xor XOR2 (N7301, N7296, N294);
xor XOR2 (N7302, N7300, N6940);
or OR4 (N7303, N7291, N5640, N6425, N5213);
not NOT1 (N7304, N7278);
or OR2 (N7305, N7299, N6684);
xor XOR2 (N7306, N7297, N1187);
xor XOR2 (N7307, N7305, N2007);
buf BUF1 (N7308, N7283);
or OR2 (N7309, N7302, N6535);
not NOT1 (N7310, N7289);
nor NOR3 (N7311, N7306, N4901, N4467);
xor XOR2 (N7312, N7304, N4279);
xor XOR2 (N7313, N7308, N5600);
nor NOR4 (N7314, N7313, N2963, N4212, N3540);
or OR3 (N7315, N7312, N5985, N2991);
and AND2 (N7316, N7293, N5370);
and AND3 (N7317, N7303, N3312, N4219);
not NOT1 (N7318, N7314);
buf BUF1 (N7319, N7309);
nor NOR3 (N7320, N7316, N2813, N1281);
nor NOR3 (N7321, N7295, N323, N1472);
or OR3 (N7322, N7315, N5746, N723);
buf BUF1 (N7323, N7317);
or OR3 (N7324, N7320, N3265, N7149);
buf BUF1 (N7325, N7301);
or OR2 (N7326, N7322, N5287);
nor NOR3 (N7327, N7324, N4762, N2716);
or OR3 (N7328, N7321, N253, N4138);
xor XOR2 (N7329, N7323, N6678);
xor XOR2 (N7330, N7328, N4997);
nand NAND3 (N7331, N7329, N1929, N5618);
buf BUF1 (N7332, N7326);
not NOT1 (N7333, N7327);
nand NAND4 (N7334, N7307, N6662, N3244, N3692);
nand NAND2 (N7335, N7330, N7253);
not NOT1 (N7336, N7333);
nor NOR3 (N7337, N7318, N5026, N1718);
nand NAND4 (N7338, N7332, N6342, N3044, N2232);
nor NOR4 (N7339, N7325, N2941, N1737, N5632);
nor NOR2 (N7340, N7339, N4949);
or OR3 (N7341, N7310, N5110, N4942);
nand NAND3 (N7342, N7340, N4066, N2038);
not NOT1 (N7343, N7341);
not NOT1 (N7344, N7337);
nand NAND4 (N7345, N7311, N3734, N3021, N5285);
nand NAND4 (N7346, N7334, N5710, N1181, N4228);
or OR4 (N7347, N7343, N7047, N4714, N4957);
not NOT1 (N7348, N7346);
xor XOR2 (N7349, N7348, N1502);
or OR2 (N7350, N7347, N2626);
and AND2 (N7351, N7331, N4830);
or OR3 (N7352, N7336, N5291, N3322);
or OR3 (N7353, N7352, N6112, N295);
not NOT1 (N7354, N7319);
not NOT1 (N7355, N7353);
or OR2 (N7356, N7342, N3217);
not NOT1 (N7357, N7344);
buf BUF1 (N7358, N7356);
and AND3 (N7359, N7338, N1672, N3256);
nand NAND3 (N7360, N7354, N4104, N2720);
or OR3 (N7361, N7345, N3142, N1799);
not NOT1 (N7362, N7359);
nor NOR2 (N7363, N7350, N5991);
and AND2 (N7364, N7335, N7355);
buf BUF1 (N7365, N4286);
or OR4 (N7366, N7364, N4453, N5912, N1200);
nor NOR3 (N7367, N7357, N3213, N2491);
nand NAND2 (N7368, N7366, N327);
nor NOR4 (N7369, N7368, N6850, N3802, N5675);
not NOT1 (N7370, N7365);
and AND4 (N7371, N7367, N5980, N2654, N3541);
or OR4 (N7372, N7370, N4371, N4187, N3727);
not NOT1 (N7373, N7361);
buf BUF1 (N7374, N7371);
not NOT1 (N7375, N7363);
buf BUF1 (N7376, N7349);
and AND2 (N7377, N7358, N740);
or OR2 (N7378, N7362, N4139);
or OR4 (N7379, N7375, N1346, N5335, N2060);
nand NAND2 (N7380, N7369, N2975);
and AND2 (N7381, N7379, N778);
buf BUF1 (N7382, N7372);
nor NOR3 (N7383, N7380, N5489, N590);
xor XOR2 (N7384, N7383, N3769);
nand NAND2 (N7385, N7376, N1319);
nand NAND2 (N7386, N7381, N5986);
xor XOR2 (N7387, N7384, N588);
or OR4 (N7388, N7374, N866, N7140, N435);
and AND2 (N7389, N7377, N1601);
nand NAND2 (N7390, N7388, N1490);
buf BUF1 (N7391, N7360);
not NOT1 (N7392, N7385);
nor NOR3 (N7393, N7351, N473, N2358);
xor XOR2 (N7394, N7386, N4180);
buf BUF1 (N7395, N7394);
buf BUF1 (N7396, N7378);
buf BUF1 (N7397, N7387);
nor NOR2 (N7398, N7392, N6387);
nor NOR4 (N7399, N7391, N1343, N1043, N2822);
or OR4 (N7400, N7398, N3325, N1734, N1106);
not NOT1 (N7401, N7396);
nand NAND2 (N7402, N7397, N5689);
nor NOR3 (N7403, N7402, N1707, N5344);
and AND4 (N7404, N7403, N3462, N4752, N6057);
nor NOR3 (N7405, N7401, N4938, N6656);
nand NAND2 (N7406, N7400, N5758);
buf BUF1 (N7407, N7373);
not NOT1 (N7408, N7399);
xor XOR2 (N7409, N7393, N6386);
nor NOR4 (N7410, N7390, N1234, N1010, N2462);
buf BUF1 (N7411, N7406);
and AND3 (N7412, N7409, N2386, N6859);
nand NAND3 (N7413, N7405, N541, N3616);
buf BUF1 (N7414, N7395);
xor XOR2 (N7415, N7408, N73);
buf BUF1 (N7416, N7415);
not NOT1 (N7417, N7407);
and AND2 (N7418, N7413, N2297);
nand NAND2 (N7419, N7416, N4212);
nor NOR3 (N7420, N7404, N1769, N1951);
or OR4 (N7421, N7410, N6504, N70, N2880);
nand NAND2 (N7422, N7382, N728);
or OR4 (N7423, N7418, N1711, N6170, N5697);
or OR3 (N7424, N7423, N6166, N6800);
and AND4 (N7425, N7421, N5271, N1468, N4631);
not NOT1 (N7426, N7412);
nand NAND2 (N7427, N7389, N5683);
nor NOR3 (N7428, N7417, N6807, N1659);
and AND3 (N7429, N7425, N5898, N6178);
and AND3 (N7430, N7414, N2554, N5196);
not NOT1 (N7431, N7428);
and AND3 (N7432, N7426, N717, N6755);
nor NOR2 (N7433, N7420, N5820);
or OR2 (N7434, N7430, N4271);
nor NOR2 (N7435, N7429, N1163);
and AND4 (N7436, N7433, N5612, N2283, N557);
nand NAND2 (N7437, N7419, N1976);
nand NAND4 (N7438, N7422, N4322, N7120, N3854);
not NOT1 (N7439, N7427);
xor XOR2 (N7440, N7437, N1318);
and AND4 (N7441, N7424, N6942, N2642, N2988);
nand NAND4 (N7442, N7436, N6932, N3119, N2413);
not NOT1 (N7443, N7439);
not NOT1 (N7444, N7442);
nand NAND2 (N7445, N7440, N7031);
buf BUF1 (N7446, N7431);
not NOT1 (N7447, N7444);
not NOT1 (N7448, N7446);
buf BUF1 (N7449, N7447);
nor NOR3 (N7450, N7432, N1366, N4099);
nand NAND4 (N7451, N7443, N2578, N3613, N1585);
and AND3 (N7452, N7438, N5636, N4852);
nand NAND2 (N7453, N7445, N6765);
and AND3 (N7454, N7448, N4313, N1);
nor NOR4 (N7455, N7411, N6215, N7026, N2809);
nand NAND3 (N7456, N7453, N1014, N5042);
nor NOR2 (N7457, N7455, N831);
xor XOR2 (N7458, N7457, N73);
buf BUF1 (N7459, N7434);
nand NAND2 (N7460, N7454, N4078);
nor NOR3 (N7461, N7456, N447, N234);
buf BUF1 (N7462, N7450);
xor XOR2 (N7463, N7458, N5451);
or OR4 (N7464, N7449, N6244, N2935, N3341);
nand NAND4 (N7465, N7462, N2893, N6030, N4390);
xor XOR2 (N7466, N7459, N4742);
or OR3 (N7467, N7451, N5829, N5438);
or OR4 (N7468, N7465, N7416, N5648, N108);
not NOT1 (N7469, N7441);
nand NAND3 (N7470, N7460, N405, N7165);
and AND4 (N7471, N7461, N2978, N4224, N2374);
not NOT1 (N7472, N7435);
xor XOR2 (N7473, N7469, N2267);
nor NOR3 (N7474, N7464, N3374, N6461);
xor XOR2 (N7475, N7468, N1078);
not NOT1 (N7476, N7472);
and AND4 (N7477, N7467, N5366, N5525, N6428);
nand NAND2 (N7478, N7477, N6645);
buf BUF1 (N7479, N7463);
xor XOR2 (N7480, N7471, N3727);
nand NAND2 (N7481, N7452, N5952);
or OR4 (N7482, N7481, N6086, N1251, N6165);
nand NAND4 (N7483, N7480, N1016, N5794, N3059);
xor XOR2 (N7484, N7466, N571);
nand NAND2 (N7485, N7483, N3245);
buf BUF1 (N7486, N7474);
xor XOR2 (N7487, N7475, N6934);
and AND4 (N7488, N7482, N4468, N4720, N1000);
nand NAND2 (N7489, N7484, N1988);
or OR3 (N7490, N7489, N4305, N4879);
nor NOR4 (N7491, N7476, N5052, N2573, N3431);
nor NOR3 (N7492, N7486, N5973, N2165);
or OR4 (N7493, N7470, N1317, N1643, N916);
buf BUF1 (N7494, N7473);
buf BUF1 (N7495, N7492);
nor NOR4 (N7496, N7495, N2295, N3810, N5517);
or OR4 (N7497, N7494, N4512, N2666, N4428);
xor XOR2 (N7498, N7497, N383);
not NOT1 (N7499, N7479);
nor NOR2 (N7500, N7485, N382);
buf BUF1 (N7501, N7500);
nand NAND3 (N7502, N7487, N5721, N4033);
not NOT1 (N7503, N7478);
nand NAND3 (N7504, N7491, N5049, N5878);
buf BUF1 (N7505, N7498);
or OR3 (N7506, N7490, N6528, N7098);
nor NOR2 (N7507, N7502, N6413);
nand NAND2 (N7508, N7501, N2328);
buf BUF1 (N7509, N7508);
nand NAND3 (N7510, N7506, N5151, N1817);
or OR3 (N7511, N7505, N2364, N4534);
or OR3 (N7512, N7511, N5789, N6823);
nand NAND3 (N7513, N7504, N5093, N1134);
nand NAND4 (N7514, N7513, N130, N5744, N5665);
not NOT1 (N7515, N7493);
nand NAND3 (N7516, N7499, N4680, N3805);
buf BUF1 (N7517, N7516);
and AND2 (N7518, N7509, N1576);
not NOT1 (N7519, N7496);
nor NOR4 (N7520, N7515, N2958, N3554, N7192);
and AND3 (N7521, N7510, N1494, N3031);
xor XOR2 (N7522, N7512, N3200);
not NOT1 (N7523, N7520);
buf BUF1 (N7524, N7521);
and AND2 (N7525, N7488, N605);
nand NAND4 (N7526, N7519, N1028, N5274, N3917);
and AND3 (N7527, N7525, N2323, N6424);
not NOT1 (N7528, N7518);
buf BUF1 (N7529, N7527);
not NOT1 (N7530, N7529);
nor NOR4 (N7531, N7528, N466, N3478, N5477);
and AND4 (N7532, N7507, N3600, N402, N3813);
not NOT1 (N7533, N7523);
nand NAND3 (N7534, N7533, N242, N4203);
and AND4 (N7535, N7517, N5937, N2238, N1702);
nand NAND2 (N7536, N7526, N1745);
buf BUF1 (N7537, N7530);
not NOT1 (N7538, N7522);
buf BUF1 (N7539, N7514);
or OR4 (N7540, N7539, N1467, N5815, N4035);
or OR4 (N7541, N7531, N3099, N2509, N6817);
nand NAND3 (N7542, N7534, N6265, N1523);
not NOT1 (N7543, N7540);
not NOT1 (N7544, N7535);
buf BUF1 (N7545, N7524);
and AND4 (N7546, N7536, N655, N4710, N5233);
or OR2 (N7547, N7546, N560);
and AND2 (N7548, N7541, N2049);
and AND4 (N7549, N7542, N535, N4098, N7197);
nor NOR2 (N7550, N7548, N5779);
buf BUF1 (N7551, N7547);
or OR2 (N7552, N7538, N2804);
not NOT1 (N7553, N7544);
and AND4 (N7554, N7553, N3413, N1163, N2711);
or OR3 (N7555, N7549, N3109, N6594);
or OR2 (N7556, N7545, N2391);
nand NAND2 (N7557, N7550, N3219);
xor XOR2 (N7558, N7503, N7142);
not NOT1 (N7559, N7554);
xor XOR2 (N7560, N7556, N4444);
nor NOR4 (N7561, N7552, N6536, N6442, N2216);
nand NAND4 (N7562, N7561, N6627, N6178, N3340);
or OR4 (N7563, N7537, N889, N5688, N7343);
and AND4 (N7564, N7562, N3323, N3380, N1300);
or OR3 (N7565, N7543, N5304, N6884);
nor NOR3 (N7566, N7559, N1011, N7420);
not NOT1 (N7567, N7560);
or OR4 (N7568, N7565, N6035, N360, N5558);
and AND4 (N7569, N7558, N5883, N5771, N7350);
xor XOR2 (N7570, N7532, N3638);
buf BUF1 (N7571, N7563);
buf BUF1 (N7572, N7551);
xor XOR2 (N7573, N7568, N1249);
and AND2 (N7574, N7570, N4181);
nor NOR2 (N7575, N7564, N388);
nor NOR4 (N7576, N7566, N2211, N2780, N284);
buf BUF1 (N7577, N7575);
not NOT1 (N7578, N7567);
or OR3 (N7579, N7576, N7326, N7227);
and AND4 (N7580, N7572, N1780, N3179, N2136);
and AND3 (N7581, N7569, N2894, N1234);
nand NAND4 (N7582, N7581, N5691, N7355, N3328);
nor NOR4 (N7583, N7580, N3863, N3392, N453);
or OR2 (N7584, N7579, N1321);
not NOT1 (N7585, N7582);
buf BUF1 (N7586, N7555);
nand NAND2 (N7587, N7584, N2312);
buf BUF1 (N7588, N7574);
nand NAND3 (N7589, N7585, N4185, N6605);
xor XOR2 (N7590, N7583, N7227);
nor NOR2 (N7591, N7589, N593);
or OR3 (N7592, N7571, N3304, N2877);
not NOT1 (N7593, N7573);
buf BUF1 (N7594, N7592);
nor NOR3 (N7595, N7594, N4596, N479);
or OR4 (N7596, N7593, N1636, N1021, N7509);
buf BUF1 (N7597, N7586);
and AND4 (N7598, N7596, N7199, N3999, N1887);
or OR4 (N7599, N7557, N3439, N1931, N3366);
nand NAND4 (N7600, N7591, N19, N2786, N2211);
or OR2 (N7601, N7597, N1607);
xor XOR2 (N7602, N7577, N3909);
nor NOR4 (N7603, N7595, N659, N535, N674);
nor NOR2 (N7604, N7601, N2852);
nor NOR4 (N7605, N7604, N2758, N1263, N4579);
not NOT1 (N7606, N7599);
nor NOR3 (N7607, N7602, N2180, N456);
not NOT1 (N7608, N7590);
and AND2 (N7609, N7607, N553);
not NOT1 (N7610, N7598);
buf BUF1 (N7611, N7603);
and AND4 (N7612, N7588, N2264, N140, N2982);
nand NAND3 (N7613, N7610, N3062, N5580);
nand NAND4 (N7614, N7612, N5036, N6679, N7091);
nor NOR4 (N7615, N7605, N6206, N2860, N1700);
nor NOR2 (N7616, N7578, N4093);
or OR2 (N7617, N7611, N5905);
xor XOR2 (N7618, N7613, N1631);
xor XOR2 (N7619, N7618, N464);
not NOT1 (N7620, N7600);
buf BUF1 (N7621, N7616);
nand NAND2 (N7622, N7609, N7478);
nand NAND4 (N7623, N7614, N4091, N6155, N1136);
nand NAND3 (N7624, N7608, N3264, N2766);
or OR4 (N7625, N7587, N1687, N2327, N6793);
or OR2 (N7626, N7617, N1260);
nor NOR2 (N7627, N7619, N1110);
or OR3 (N7628, N7624, N3570, N4264);
nand NAND3 (N7629, N7615, N1367, N6901);
nor NOR2 (N7630, N7621, N2310);
nand NAND3 (N7631, N7626, N387, N1110);
nor NOR2 (N7632, N7622, N6522);
and AND3 (N7633, N7632, N316, N4334);
buf BUF1 (N7634, N7625);
and AND2 (N7635, N7620, N1740);
xor XOR2 (N7636, N7627, N5045);
xor XOR2 (N7637, N7633, N1199);
and AND4 (N7638, N7635, N5410, N4633, N6557);
xor XOR2 (N7639, N7628, N6193);
nand NAND4 (N7640, N7629, N3294, N6707, N398);
buf BUF1 (N7641, N7638);
nor NOR3 (N7642, N7606, N5266, N2855);
nand NAND3 (N7643, N7623, N2341, N5534);
xor XOR2 (N7644, N7642, N4328);
or OR2 (N7645, N7644, N6278);
not NOT1 (N7646, N7631);
xor XOR2 (N7647, N7637, N494);
nand NAND3 (N7648, N7646, N3957, N4092);
xor XOR2 (N7649, N7640, N6721);
and AND2 (N7650, N7649, N3999);
nor NOR4 (N7651, N7648, N2095, N404, N3226);
buf BUF1 (N7652, N7645);
nand NAND3 (N7653, N7639, N645, N2869);
and AND3 (N7654, N7641, N3538, N4896);
or OR4 (N7655, N7636, N5019, N1348, N4089);
or OR3 (N7656, N7653, N7246, N4378);
and AND2 (N7657, N7652, N6113);
nor NOR2 (N7658, N7654, N6735);
nor NOR2 (N7659, N7657, N7251);
not NOT1 (N7660, N7656);
and AND3 (N7661, N7659, N6938, N4252);
buf BUF1 (N7662, N7660);
not NOT1 (N7663, N7650);
or OR4 (N7664, N7661, N7640, N4775, N5768);
buf BUF1 (N7665, N7664);
nor NOR4 (N7666, N7655, N2568, N3730, N5424);
not NOT1 (N7667, N7663);
buf BUF1 (N7668, N7630);
and AND3 (N7669, N7668, N92, N793);
xor XOR2 (N7670, N7634, N5033);
not NOT1 (N7671, N7669);
not NOT1 (N7672, N7647);
nand NAND3 (N7673, N7670, N4912, N3896);
and AND3 (N7674, N7658, N1907, N4764);
or OR4 (N7675, N7651, N5800, N4259, N6335);
and AND2 (N7676, N7675, N656);
buf BUF1 (N7677, N7676);
buf BUF1 (N7678, N7671);
not NOT1 (N7679, N7674);
not NOT1 (N7680, N7672);
nand NAND3 (N7681, N7677, N2137, N2424);
and AND4 (N7682, N7681, N1381, N1261, N5067);
buf BUF1 (N7683, N7666);
not NOT1 (N7684, N7643);
and AND3 (N7685, N7684, N4654, N1698);
buf BUF1 (N7686, N7679);
or OR3 (N7687, N7667, N1956, N6810);
nand NAND2 (N7688, N7686, N6230);
not NOT1 (N7689, N7665);
and AND4 (N7690, N7678, N1300, N6622, N3586);
not NOT1 (N7691, N7662);
not NOT1 (N7692, N7689);
xor XOR2 (N7693, N7680, N3600);
or OR4 (N7694, N7673, N753, N270, N3847);
xor XOR2 (N7695, N7690, N9);
and AND2 (N7696, N7682, N6723);
nand NAND2 (N7697, N7687, N5764);
nor NOR4 (N7698, N7693, N2235, N7089, N6225);
nand NAND2 (N7699, N7691, N3048);
or OR3 (N7700, N7692, N6670, N1801);
and AND3 (N7701, N7697, N271, N867);
nor NOR4 (N7702, N7688, N2902, N5914, N6553);
buf BUF1 (N7703, N7696);
nand NAND3 (N7704, N7683, N3546, N1749);
nor NOR4 (N7705, N7704, N5010, N7477, N6759);
and AND3 (N7706, N7702, N6446, N6291);
nor NOR4 (N7707, N7695, N5115, N7665, N3088);
not NOT1 (N7708, N7698);
and AND4 (N7709, N7706, N24, N2500, N4994);
xor XOR2 (N7710, N7701, N574);
or OR3 (N7711, N7685, N7355, N1588);
not NOT1 (N7712, N7709);
buf BUF1 (N7713, N7712);
nor NOR3 (N7714, N7700, N5691, N7014);
buf BUF1 (N7715, N7707);
nor NOR2 (N7716, N7705, N4509);
or OR3 (N7717, N7714, N429, N6365);
xor XOR2 (N7718, N7703, N2869);
buf BUF1 (N7719, N7718);
nor NOR3 (N7720, N7719, N3820, N4640);
not NOT1 (N7721, N7720);
xor XOR2 (N7722, N7721, N6251);
nor NOR2 (N7723, N7711, N3197);
or OR4 (N7724, N7699, N4741, N85, N2927);
buf BUF1 (N7725, N7724);
nand NAND2 (N7726, N7725, N2599);
nand NAND3 (N7727, N7723, N2279, N3426);
nor NOR3 (N7728, N7717, N3084, N6339);
or OR4 (N7729, N7713, N4798, N1645, N3338);
nand NAND3 (N7730, N7726, N301, N3521);
or OR4 (N7731, N7716, N1600, N2218, N3965);
not NOT1 (N7732, N7727);
or OR3 (N7733, N7708, N4289, N1110);
or OR2 (N7734, N7730, N4407);
not NOT1 (N7735, N7733);
not NOT1 (N7736, N7734);
nand NAND3 (N7737, N7732, N2171, N2463);
and AND3 (N7738, N7731, N5488, N1160);
nor NOR4 (N7739, N7735, N3803, N3746, N5384);
or OR4 (N7740, N7738, N4313, N3996, N3146);
xor XOR2 (N7741, N7736, N4622);
buf BUF1 (N7742, N7740);
nor NOR3 (N7743, N7742, N1133, N706);
and AND3 (N7744, N7739, N17, N7243);
nand NAND3 (N7745, N7729, N4303, N3544);
xor XOR2 (N7746, N7715, N2742);
buf BUF1 (N7747, N7745);
xor XOR2 (N7748, N7728, N5870);
nand NAND3 (N7749, N7737, N5868, N922);
or OR3 (N7750, N7746, N3385, N7412);
nor NOR3 (N7751, N7744, N1558, N5574);
nor NOR2 (N7752, N7741, N4085);
and AND3 (N7753, N7748, N5453, N1764);
xor XOR2 (N7754, N7722, N1191);
not NOT1 (N7755, N7749);
nand NAND3 (N7756, N7747, N2267, N3575);
and AND4 (N7757, N7755, N4116, N5088, N786);
nand NAND2 (N7758, N7743, N1827);
buf BUF1 (N7759, N7752);
xor XOR2 (N7760, N7756, N3074);
xor XOR2 (N7761, N7757, N2099);
xor XOR2 (N7762, N7753, N1544);
and AND3 (N7763, N7694, N1802, N397);
nand NAND4 (N7764, N7762, N1119, N151, N2816);
xor XOR2 (N7765, N7759, N5254);
buf BUF1 (N7766, N7763);
nand NAND2 (N7767, N7760, N4894);
nand NAND3 (N7768, N7750, N3524, N3252);
not NOT1 (N7769, N7758);
and AND2 (N7770, N7768, N3668);
nor NOR3 (N7771, N7761, N2121, N4558);
not NOT1 (N7772, N7765);
nand NAND3 (N7773, N7764, N6539, N4144);
or OR4 (N7774, N7767, N2119, N5223, N1443);
buf BUF1 (N7775, N7751);
xor XOR2 (N7776, N7774, N7720);
buf BUF1 (N7777, N7770);
nand NAND4 (N7778, N7777, N5360, N5375, N5139);
or OR3 (N7779, N7775, N3953, N1751);
nand NAND2 (N7780, N7754, N3366);
and AND2 (N7781, N7780, N5234);
or OR3 (N7782, N7776, N831, N6913);
nand NAND3 (N7783, N7773, N1152, N5056);
buf BUF1 (N7784, N7783);
and AND4 (N7785, N7784, N6497, N7651, N3072);
and AND3 (N7786, N7785, N3503, N7712);
nor NOR4 (N7787, N7786, N4959, N268, N2600);
and AND3 (N7788, N7782, N1782, N2295);
or OR4 (N7789, N7771, N3799, N6327, N5851);
buf BUF1 (N7790, N7769);
not NOT1 (N7791, N7710);
nand NAND2 (N7792, N7787, N5168);
and AND3 (N7793, N7766, N1815, N2138);
xor XOR2 (N7794, N7790, N5653);
nand NAND2 (N7795, N7792, N3370);
not NOT1 (N7796, N7779);
nor NOR2 (N7797, N7772, N2618);
not NOT1 (N7798, N7793);
not NOT1 (N7799, N7791);
not NOT1 (N7800, N7797);
nand NAND4 (N7801, N7796, N4060, N4009, N4721);
nor NOR3 (N7802, N7799, N1051, N4571);
not NOT1 (N7803, N7801);
xor XOR2 (N7804, N7802, N4481);
xor XOR2 (N7805, N7795, N4849);
nand NAND2 (N7806, N7798, N1757);
not NOT1 (N7807, N7805);
not NOT1 (N7808, N7789);
xor XOR2 (N7809, N7806, N428);
xor XOR2 (N7810, N7800, N817);
and AND3 (N7811, N7794, N1889, N3566);
not NOT1 (N7812, N7810);
or OR2 (N7813, N7812, N7428);
not NOT1 (N7814, N7781);
or OR3 (N7815, N7804, N3479, N6087);
nor NOR3 (N7816, N7778, N3126, N7645);
buf BUF1 (N7817, N7808);
or OR3 (N7818, N7813, N6277, N5827);
or OR2 (N7819, N7807, N6365);
or OR2 (N7820, N7811, N5163);
buf BUF1 (N7821, N7819);
not NOT1 (N7822, N7815);
xor XOR2 (N7823, N7788, N771);
or OR3 (N7824, N7814, N1285, N7463);
and AND2 (N7825, N7818, N7254);
nor NOR2 (N7826, N7816, N1842);
not NOT1 (N7827, N7822);
buf BUF1 (N7828, N7820);
or OR2 (N7829, N7828, N1101);
or OR3 (N7830, N7827, N7371, N107);
nand NAND3 (N7831, N7830, N2318, N878);
buf BUF1 (N7832, N7829);
nor NOR2 (N7833, N7817, N3494);
xor XOR2 (N7834, N7824, N1132);
nor NOR3 (N7835, N7834, N7203, N1455);
buf BUF1 (N7836, N7826);
nand NAND2 (N7837, N7836, N4336);
nand NAND4 (N7838, N7831, N4897, N3807, N5411);
nor NOR3 (N7839, N7837, N6743, N1860);
and AND3 (N7840, N7838, N2181, N7350);
not NOT1 (N7841, N7840);
and AND4 (N7842, N7841, N608, N5982, N5045);
buf BUF1 (N7843, N7825);
and AND4 (N7844, N7823, N3295, N3801, N2156);
buf BUF1 (N7845, N7833);
and AND2 (N7846, N7803, N5890);
xor XOR2 (N7847, N7821, N341);
buf BUF1 (N7848, N7809);
or OR3 (N7849, N7835, N2368, N1488);
nand NAND2 (N7850, N7844, N6642);
and AND2 (N7851, N7850, N4547);
nor NOR3 (N7852, N7845, N5442, N5684);
nand NAND2 (N7853, N7849, N2940);
buf BUF1 (N7854, N7847);
nor NOR4 (N7855, N7851, N1379, N448, N5839);
nand NAND4 (N7856, N7853, N2274, N1723, N3245);
nor NOR4 (N7857, N7846, N1994, N367, N7478);
or OR3 (N7858, N7852, N3468, N3567);
or OR4 (N7859, N7843, N7654, N5480, N7347);
xor XOR2 (N7860, N7858, N3132);
buf BUF1 (N7861, N7855);
not NOT1 (N7862, N7859);
buf BUF1 (N7863, N7861);
xor XOR2 (N7864, N7863, N4931);
xor XOR2 (N7865, N7842, N6033);
nand NAND2 (N7866, N7839, N3959);
nand NAND3 (N7867, N7864, N3757, N3733);
or OR2 (N7868, N7862, N458);
or OR3 (N7869, N7856, N6488, N702);
and AND2 (N7870, N7868, N7426);
not NOT1 (N7871, N7848);
buf BUF1 (N7872, N7857);
or OR2 (N7873, N7871, N6065);
or OR3 (N7874, N7870, N7129, N94);
buf BUF1 (N7875, N7866);
xor XOR2 (N7876, N7872, N2902);
or OR3 (N7877, N7860, N2, N3573);
xor XOR2 (N7878, N7867, N7470);
not NOT1 (N7879, N7876);
xor XOR2 (N7880, N7874, N2475);
and AND4 (N7881, N7869, N1359, N2066, N7519);
not NOT1 (N7882, N7879);
not NOT1 (N7883, N7865);
not NOT1 (N7884, N7878);
or OR3 (N7885, N7875, N6945, N3363);
nor NOR4 (N7886, N7877, N1541, N1840, N3565);
buf BUF1 (N7887, N7880);
buf BUF1 (N7888, N7886);
nor NOR3 (N7889, N7883, N5756, N6071);
or OR4 (N7890, N7888, N6396, N2842, N2336);
not NOT1 (N7891, N7884);
buf BUF1 (N7892, N7891);
nor NOR3 (N7893, N7873, N68, N7559);
not NOT1 (N7894, N7885);
xor XOR2 (N7895, N7854, N5865);
or OR3 (N7896, N7890, N6991, N5605);
buf BUF1 (N7897, N7881);
and AND4 (N7898, N7896, N7765, N7081, N7750);
buf BUF1 (N7899, N7889);
xor XOR2 (N7900, N7893, N5078);
nor NOR2 (N7901, N7895, N4842);
and AND4 (N7902, N7899, N4672, N6253, N4283);
nor NOR4 (N7903, N7894, N432, N778, N7276);
and AND2 (N7904, N7902, N7032);
nand NAND4 (N7905, N7882, N7766, N3983, N1653);
not NOT1 (N7906, N7887);
nor NOR4 (N7907, N7906, N6190, N392, N2694);
nand NAND2 (N7908, N7892, N906);
not NOT1 (N7909, N7904);
not NOT1 (N7910, N7898);
and AND4 (N7911, N7905, N3419, N3551, N2663);
not NOT1 (N7912, N7900);
xor XOR2 (N7913, N7911, N673);
xor XOR2 (N7914, N7907, N7754);
nand NAND4 (N7915, N7910, N4863, N3138, N7253);
nand NAND4 (N7916, N7909, N6934, N3631, N5006);
not NOT1 (N7917, N7897);
and AND4 (N7918, N7914, N1518, N1545, N3979);
and AND3 (N7919, N7908, N3736, N4016);
and AND3 (N7920, N7919, N6244, N5944);
and AND4 (N7921, N7916, N6838, N5562, N5425);
not NOT1 (N7922, N7912);
not NOT1 (N7923, N7922);
or OR3 (N7924, N7921, N6595, N1979);
not NOT1 (N7925, N7917);
nor NOR2 (N7926, N7832, N7754);
nand NAND4 (N7927, N7918, N2866, N6917, N6374);
and AND3 (N7928, N7901, N6090, N7322);
xor XOR2 (N7929, N7920, N2855);
and AND3 (N7930, N7925, N3544, N2107);
nor NOR2 (N7931, N7924, N5434);
nor NOR2 (N7932, N7931, N7018);
nand NAND4 (N7933, N7930, N5818, N2529, N7132);
nor NOR2 (N7934, N7913, N3033);
nand NAND3 (N7935, N7928, N1044, N3365);
xor XOR2 (N7936, N7926, N2388);
xor XOR2 (N7937, N7929, N932);
nor NOR3 (N7938, N7934, N5495, N1784);
not NOT1 (N7939, N7935);
and AND4 (N7940, N7903, N1554, N5491, N1499);
xor XOR2 (N7941, N7932, N4385);
buf BUF1 (N7942, N7936);
or OR4 (N7943, N7940, N7916, N2136, N3576);
not NOT1 (N7944, N7938);
nand NAND2 (N7945, N7939, N6050);
nor NOR3 (N7946, N7945, N4083, N6789);
or OR4 (N7947, N7923, N4010, N5576, N1201);
and AND3 (N7948, N7927, N6056, N3840);
nor NOR3 (N7949, N7946, N1923, N4810);
or OR4 (N7950, N7937, N3663, N1359, N2904);
not NOT1 (N7951, N7947);
nor NOR3 (N7952, N7942, N1049, N803);
nand NAND4 (N7953, N7949, N7476, N6257, N37);
nor NOR3 (N7954, N7948, N6585, N322);
and AND4 (N7955, N7954, N6659, N7170, N4310);
and AND2 (N7956, N7941, N3059);
xor XOR2 (N7957, N7952, N6783);
nand NAND2 (N7958, N7950, N581);
not NOT1 (N7959, N7955);
and AND3 (N7960, N7958, N3570, N255);
or OR3 (N7961, N7957, N3215, N2844);
xor XOR2 (N7962, N7944, N5505);
nor NOR3 (N7963, N7962, N4024, N3401);
nor NOR2 (N7964, N7960, N7624);
or OR4 (N7965, N7961, N4729, N7215, N5954);
nor NOR3 (N7966, N7956, N3634, N5125);
not NOT1 (N7967, N7953);
not NOT1 (N7968, N7943);
not NOT1 (N7969, N7915);
xor XOR2 (N7970, N7951, N4596);
buf BUF1 (N7971, N7933);
and AND4 (N7972, N7966, N7002, N2297, N6411);
xor XOR2 (N7973, N7969, N774);
nand NAND3 (N7974, N7959, N2032, N7649);
nor NOR4 (N7975, N7965, N4791, N2750, N3498);
nand NAND4 (N7976, N7971, N2591, N1179, N7404);
xor XOR2 (N7977, N7964, N1505);
not NOT1 (N7978, N7976);
not NOT1 (N7979, N7963);
not NOT1 (N7980, N7978);
xor XOR2 (N7981, N7980, N5600);
nand NAND2 (N7982, N7973, N7186);
buf BUF1 (N7983, N7982);
xor XOR2 (N7984, N7975, N7420);
nor NOR3 (N7985, N7977, N4070, N223);
xor XOR2 (N7986, N7974, N2787);
nand NAND2 (N7987, N7972, N4919);
nor NOR3 (N7988, N7985, N6955, N6014);
buf BUF1 (N7989, N7988);
nor NOR2 (N7990, N7986, N7053);
nand NAND3 (N7991, N7981, N4986, N1282);
buf BUF1 (N7992, N7968);
nor NOR2 (N7993, N7991, N5285);
or OR4 (N7994, N7984, N4858, N1919, N4068);
xor XOR2 (N7995, N7987, N3072);
not NOT1 (N7996, N7989);
buf BUF1 (N7997, N7992);
nand NAND2 (N7998, N7990, N1459);
nand NAND2 (N7999, N7967, N227);
buf BUF1 (N8000, N7979);
and AND3 (N8001, N7999, N2547, N1564);
nor NOR3 (N8002, N7995, N3026, N7687);
nand NAND4 (N8003, N8001, N6028, N1968, N7154);
buf BUF1 (N8004, N8002);
not NOT1 (N8005, N7970);
and AND2 (N8006, N7983, N6969);
not NOT1 (N8007, N7994);
nor NOR4 (N8008, N8003, N3787, N1459, N7024);
xor XOR2 (N8009, N7993, N6710);
nor NOR2 (N8010, N8009, N67);
nor NOR4 (N8011, N7997, N1279, N5495, N6835);
buf BUF1 (N8012, N8000);
buf BUF1 (N8013, N8008);
and AND4 (N8014, N8004, N3178, N6445, N6440);
nand NAND3 (N8015, N8010, N3693, N2698);
not NOT1 (N8016, N8007);
nor NOR4 (N8017, N8016, N3672, N5267, N7617);
and AND2 (N8018, N7998, N3681);
xor XOR2 (N8019, N7996, N4885);
nor NOR3 (N8020, N8014, N2859, N1192);
buf BUF1 (N8021, N8020);
not NOT1 (N8022, N8011);
not NOT1 (N8023, N8013);
xor XOR2 (N8024, N8023, N7017);
not NOT1 (N8025, N8017);
or OR3 (N8026, N8018, N6056, N7403);
xor XOR2 (N8027, N8024, N2715);
and AND4 (N8028, N8021, N5459, N7338, N5557);
not NOT1 (N8029, N8005);
nor NOR4 (N8030, N8027, N6775, N6409, N3083);
nand NAND4 (N8031, N8026, N1526, N4319, N6184);
buf BUF1 (N8032, N8019);
xor XOR2 (N8033, N8032, N6099);
buf BUF1 (N8034, N8006);
or OR3 (N8035, N8029, N5482, N7202);
and AND2 (N8036, N8035, N1767);
or OR4 (N8037, N8034, N5476, N5140, N382);
xor XOR2 (N8038, N8012, N5620);
or OR3 (N8039, N8025, N5641, N2227);
or OR4 (N8040, N8031, N3434, N2319, N4539);
nand NAND2 (N8041, N8039, N3396);
nor NOR3 (N8042, N8030, N3779, N3524);
and AND4 (N8043, N8028, N2268, N4423, N7063);
and AND3 (N8044, N8042, N7026, N7421);
nand NAND2 (N8045, N8033, N7023);
nor NOR3 (N8046, N8044, N1062, N5791);
nor NOR2 (N8047, N8036, N7660);
buf BUF1 (N8048, N8038);
and AND2 (N8049, N8015, N7935);
not NOT1 (N8050, N8047);
and AND4 (N8051, N8045, N5903, N976, N2932);
xor XOR2 (N8052, N8043, N3929);
not NOT1 (N8053, N8048);
nand NAND3 (N8054, N8022, N5730, N3530);
not NOT1 (N8055, N8053);
xor XOR2 (N8056, N8050, N2130);
and AND4 (N8057, N8052, N4991, N1596, N6557);
nor NOR3 (N8058, N8041, N410, N606);
and AND4 (N8059, N8049, N7981, N7544, N963);
not NOT1 (N8060, N8040);
and AND3 (N8061, N8060, N3825, N1356);
not NOT1 (N8062, N8057);
and AND3 (N8063, N8055, N1543, N6284);
nand NAND3 (N8064, N8062, N3120, N5103);
and AND3 (N8065, N8059, N7514, N5110);
nor NOR4 (N8066, N8061, N2076, N1264, N5406);
nor NOR3 (N8067, N8066, N8000, N3271);
xor XOR2 (N8068, N8067, N1837);
and AND4 (N8069, N8046, N2649, N6437, N1393);
buf BUF1 (N8070, N8058);
xor XOR2 (N8071, N8063, N5323);
nor NOR4 (N8072, N8037, N3528, N3756, N7809);
xor XOR2 (N8073, N8069, N2774);
and AND2 (N8074, N8064, N7619);
and AND4 (N8075, N8071, N4541, N5351, N3363);
and AND2 (N8076, N8054, N7473);
nor NOR3 (N8077, N8076, N6109, N2513);
xor XOR2 (N8078, N8051, N1839);
nor NOR3 (N8079, N8070, N2132, N6961);
xor XOR2 (N8080, N8075, N7745);
not NOT1 (N8081, N8068);
not NOT1 (N8082, N8077);
not NOT1 (N8083, N8081);
buf BUF1 (N8084, N8078);
or OR2 (N8085, N8080, N2278);
or OR2 (N8086, N8085, N5797);
or OR2 (N8087, N8083, N1320);
nand NAND3 (N8088, N8073, N4765, N206);
nand NAND2 (N8089, N8082, N5);
nor NOR4 (N8090, N8086, N7663, N6598, N6963);
buf BUF1 (N8091, N8089);
not NOT1 (N8092, N8079);
nor NOR4 (N8093, N8072, N6185, N7557, N1848);
buf BUF1 (N8094, N8092);
or OR2 (N8095, N8090, N7831);
or OR3 (N8096, N8084, N4660, N2511);
or OR3 (N8097, N8065, N2028, N2644);
buf BUF1 (N8098, N8095);
nor NOR2 (N8099, N8096, N1646);
nand NAND2 (N8100, N8091, N7143);
nor NOR4 (N8101, N8100, N2470, N3085, N1750);
xor XOR2 (N8102, N8074, N8055);
not NOT1 (N8103, N8101);
nand NAND2 (N8104, N8056, N1207);
nor NOR2 (N8105, N8102, N2048);
and AND2 (N8106, N8104, N1153);
nor NOR3 (N8107, N8094, N193, N7280);
buf BUF1 (N8108, N8097);
xor XOR2 (N8109, N8093, N2016);
buf BUF1 (N8110, N8098);
not NOT1 (N8111, N8107);
not NOT1 (N8112, N8105);
nand NAND4 (N8113, N8087, N1307, N5822, N6919);
xor XOR2 (N8114, N8099, N7339);
xor XOR2 (N8115, N8110, N1960);
and AND4 (N8116, N8112, N2403, N5120, N3134);
not NOT1 (N8117, N8115);
nor NOR2 (N8118, N8114, N5003);
xor XOR2 (N8119, N8108, N4070);
nand NAND3 (N8120, N8109, N5461, N6312);
not NOT1 (N8121, N8088);
nand NAND3 (N8122, N8111, N6293, N8040);
and AND4 (N8123, N8116, N2699, N3608, N311);
buf BUF1 (N8124, N8118);
nand NAND2 (N8125, N8121, N2173);
xor XOR2 (N8126, N8125, N1985);
not NOT1 (N8127, N8124);
nor NOR2 (N8128, N8106, N5860);
and AND4 (N8129, N8120, N3886, N2899, N2553);
and AND2 (N8130, N8103, N127);
xor XOR2 (N8131, N8117, N5417);
and AND4 (N8132, N8123, N3071, N3373, N2887);
xor XOR2 (N8133, N8132, N321);
or OR4 (N8134, N8119, N987, N6853, N6924);
and AND2 (N8135, N8126, N4150);
not NOT1 (N8136, N8129);
nor NOR3 (N8137, N8135, N2811, N1767);
not NOT1 (N8138, N8137);
buf BUF1 (N8139, N8113);
nor NOR2 (N8140, N8128, N4302);
not NOT1 (N8141, N8136);
or OR4 (N8142, N8130, N6463, N1781, N1623);
nand NAND3 (N8143, N8133, N2789, N7325);
buf BUF1 (N8144, N8140);
or OR2 (N8145, N8127, N2829);
xor XOR2 (N8146, N8134, N5132);
nor NOR2 (N8147, N8144, N2547);
nand NAND2 (N8148, N8141, N2374);
not NOT1 (N8149, N8146);
xor XOR2 (N8150, N8139, N7512);
nor NOR4 (N8151, N8149, N4946, N3686, N6780);
and AND4 (N8152, N8148, N5939, N3289, N7795);
xor XOR2 (N8153, N8131, N5209);
nand NAND3 (N8154, N8150, N3745, N30);
or OR4 (N8155, N8142, N481, N270, N5947);
not NOT1 (N8156, N8145);
nor NOR3 (N8157, N8138, N3007, N1294);
nand NAND4 (N8158, N8147, N4596, N7902, N1711);
buf BUF1 (N8159, N8153);
nand NAND4 (N8160, N8157, N2773, N7638, N730);
nand NAND4 (N8161, N8143, N6, N7905, N4775);
or OR3 (N8162, N8122, N3211, N3111);
nand NAND3 (N8163, N8152, N7461, N1511);
nor NOR4 (N8164, N8158, N1112, N181, N6238);
nand NAND4 (N8165, N8163, N7958, N1087, N7894);
nand NAND2 (N8166, N8164, N1375);
xor XOR2 (N8167, N8166, N5394);
buf BUF1 (N8168, N8160);
buf BUF1 (N8169, N8168);
buf BUF1 (N8170, N8162);
buf BUF1 (N8171, N8161);
or OR3 (N8172, N8155, N5256, N1176);
nor NOR4 (N8173, N8167, N555, N1116, N4049);
nor NOR4 (N8174, N8170, N7259, N6025, N2452);
not NOT1 (N8175, N8151);
and AND4 (N8176, N8174, N2977, N4766, N7528);
nor NOR3 (N8177, N8172, N5254, N3674);
not NOT1 (N8178, N8165);
buf BUF1 (N8179, N8177);
nor NOR2 (N8180, N8156, N5925);
nand NAND4 (N8181, N8154, N5075, N3302, N426);
not NOT1 (N8182, N8173);
not NOT1 (N8183, N8176);
nand NAND3 (N8184, N8175, N7720, N6944);
or OR4 (N8185, N8179, N5540, N4424, N6942);
nand NAND2 (N8186, N8171, N6820);
nand NAND3 (N8187, N8183, N6694, N321);
nor NOR4 (N8188, N8180, N301, N6348, N7808);
nand NAND4 (N8189, N8187, N2457, N4195, N1371);
and AND2 (N8190, N8178, N185);
not NOT1 (N8191, N8182);
xor XOR2 (N8192, N8185, N409);
nor NOR3 (N8193, N8191, N4222, N4857);
nor NOR2 (N8194, N8169, N6725);
or OR3 (N8195, N8193, N4747, N7265);
buf BUF1 (N8196, N8190);
nand NAND2 (N8197, N8186, N4356);
and AND3 (N8198, N8189, N6924, N2603);
not NOT1 (N8199, N8188);
not NOT1 (N8200, N8194);
or OR4 (N8201, N8181, N2947, N1532, N3357);
nand NAND3 (N8202, N8199, N5095, N3982);
or OR2 (N8203, N8159, N5225);
buf BUF1 (N8204, N8184);
buf BUF1 (N8205, N8204);
not NOT1 (N8206, N8197);
or OR3 (N8207, N8195, N1228, N2543);
xor XOR2 (N8208, N8201, N360);
or OR2 (N8209, N8206, N2592);
nor NOR3 (N8210, N8205, N2256, N2486);
or OR4 (N8211, N8207, N5447, N4425, N859);
nor NOR4 (N8212, N8192, N4156, N6095, N1081);
nor NOR4 (N8213, N8209, N2526, N4891, N7426);
not NOT1 (N8214, N8202);
not NOT1 (N8215, N8196);
buf BUF1 (N8216, N8211);
or OR2 (N8217, N8215, N5714);
and AND2 (N8218, N8208, N4550);
buf BUF1 (N8219, N8214);
not NOT1 (N8220, N8212);
xor XOR2 (N8221, N8198, N1261);
nand NAND3 (N8222, N8218, N7574, N963);
nor NOR2 (N8223, N8200, N7137);
and AND4 (N8224, N8219, N3290, N6400, N4007);
xor XOR2 (N8225, N8216, N2747);
nor NOR4 (N8226, N8203, N869, N1236, N2246);
buf BUF1 (N8227, N8221);
not NOT1 (N8228, N8227);
nand NAND4 (N8229, N8223, N5325, N3114, N3787);
nand NAND2 (N8230, N8220, N938);
and AND2 (N8231, N8226, N5204);
buf BUF1 (N8232, N8224);
xor XOR2 (N8233, N8228, N7352);
or OR2 (N8234, N8210, N3140);
xor XOR2 (N8235, N8233, N7099);
xor XOR2 (N8236, N8231, N8047);
or OR3 (N8237, N8217, N3395, N2412);
not NOT1 (N8238, N8230);
buf BUF1 (N8239, N8235);
not NOT1 (N8240, N8237);
nor NOR3 (N8241, N8229, N6977, N6607);
or OR2 (N8242, N8213, N2927);
nand NAND3 (N8243, N8239, N5771, N2190);
not NOT1 (N8244, N8222);
buf BUF1 (N8245, N8241);
or OR3 (N8246, N8240, N6176, N2432);
or OR3 (N8247, N8246, N232, N4137);
not NOT1 (N8248, N8238);
or OR4 (N8249, N8243, N8202, N8013, N7896);
xor XOR2 (N8250, N8247, N1172);
and AND3 (N8251, N8250, N4877, N7911);
buf BUF1 (N8252, N8245);
or OR3 (N8253, N8248, N3164, N4396);
not NOT1 (N8254, N8234);
nand NAND4 (N8255, N8242, N2449, N5691, N1236);
nand NAND4 (N8256, N8251, N6090, N3792, N6797);
nand NAND2 (N8257, N8256, N2217);
nand NAND4 (N8258, N8252, N1971, N8082, N4686);
and AND2 (N8259, N8225, N1628);
buf BUF1 (N8260, N8236);
and AND3 (N8261, N8254, N2945, N7402);
nor NOR3 (N8262, N8257, N2954, N1651);
xor XOR2 (N8263, N8261, N1808);
xor XOR2 (N8264, N8255, N6781);
and AND4 (N8265, N8232, N683, N7131, N681);
and AND2 (N8266, N8258, N2263);
and AND4 (N8267, N8265, N2544, N2554, N4572);
xor XOR2 (N8268, N8244, N6489);
nor NOR3 (N8269, N8263, N8026, N7380);
nand NAND3 (N8270, N8249, N6384, N1367);
and AND3 (N8271, N8253, N271, N1916);
not NOT1 (N8272, N8262);
nor NOR3 (N8273, N8271, N4413, N5755);
and AND4 (N8274, N8270, N828, N3252, N7625);
xor XOR2 (N8275, N8264, N4712);
nand NAND4 (N8276, N8266, N3502, N4699, N2818);
nor NOR4 (N8277, N8272, N4736, N1007, N959);
and AND4 (N8278, N8269, N1665, N686, N8116);
not NOT1 (N8279, N8260);
buf BUF1 (N8280, N8267);
or OR2 (N8281, N8268, N6439);
or OR2 (N8282, N8273, N2573);
not NOT1 (N8283, N8282);
or OR2 (N8284, N8274, N137);
not NOT1 (N8285, N8284);
xor XOR2 (N8286, N8280, N2326);
or OR2 (N8287, N8279, N1158);
or OR2 (N8288, N8283, N4050);
nand NAND4 (N8289, N8276, N5339, N736, N1594);
not NOT1 (N8290, N8289);
nor NOR4 (N8291, N8290, N6737, N1422, N4882);
or OR2 (N8292, N8288, N7984);
or OR4 (N8293, N8277, N6749, N7891, N4031);
xor XOR2 (N8294, N8291, N2980);
nand NAND3 (N8295, N8259, N4886, N7697);
buf BUF1 (N8296, N8275);
buf BUF1 (N8297, N8293);
nor NOR3 (N8298, N8281, N2371, N6719);
nor NOR4 (N8299, N8297, N361, N1659, N2986);
nor NOR2 (N8300, N8294, N94);
and AND3 (N8301, N8285, N6974, N1728);
or OR3 (N8302, N8300, N1588, N1403);
buf BUF1 (N8303, N8301);
or OR2 (N8304, N8278, N569);
or OR3 (N8305, N8287, N5674, N4903);
nor NOR3 (N8306, N8305, N1164, N5121);
not NOT1 (N8307, N8286);
nand NAND2 (N8308, N8299, N668);
nor NOR2 (N8309, N8307, N6679);
or OR2 (N8310, N8292, N1648);
and AND4 (N8311, N8306, N4637, N3145, N4861);
and AND3 (N8312, N8298, N4791, N192);
or OR4 (N8313, N8311, N1725, N699, N228);
nor NOR4 (N8314, N8296, N4852, N589, N560);
buf BUF1 (N8315, N8303);
buf BUF1 (N8316, N8315);
and AND2 (N8317, N8295, N6049);
xor XOR2 (N8318, N8313, N3807);
or OR4 (N8319, N8316, N7981, N3605, N1384);
xor XOR2 (N8320, N8302, N6419);
and AND4 (N8321, N8320, N3392, N6284, N4815);
nand NAND3 (N8322, N8318, N2593, N5080);
xor XOR2 (N8323, N8310, N2638);
xor XOR2 (N8324, N8323, N3036);
nand NAND2 (N8325, N8319, N3632);
nor NOR2 (N8326, N8321, N164);
or OR4 (N8327, N8326, N2925, N6600, N2222);
xor XOR2 (N8328, N8325, N4956);
or OR2 (N8329, N8304, N7953);
nor NOR3 (N8330, N8328, N3656, N4010);
not NOT1 (N8331, N8329);
not NOT1 (N8332, N8317);
buf BUF1 (N8333, N8312);
not NOT1 (N8334, N8327);
nor NOR3 (N8335, N8330, N1855, N6600);
not NOT1 (N8336, N8333);
xor XOR2 (N8337, N8334, N6198);
and AND4 (N8338, N8324, N3665, N1334, N1311);
or OR4 (N8339, N8308, N3689, N2729, N7527);
nand NAND3 (N8340, N8314, N2178, N8201);
nor NOR3 (N8341, N8339, N5089, N2421);
nand NAND2 (N8342, N8322, N7079);
nand NAND3 (N8343, N8331, N4227, N8000);
not NOT1 (N8344, N8335);
not NOT1 (N8345, N8341);
nor NOR2 (N8346, N8332, N2674);
xor XOR2 (N8347, N8342, N3850);
xor XOR2 (N8348, N8347, N8036);
xor XOR2 (N8349, N8343, N7884);
buf BUF1 (N8350, N8336);
buf BUF1 (N8351, N8309);
nand NAND3 (N8352, N8350, N3508, N7737);
and AND3 (N8353, N8337, N4154, N8214);
and AND2 (N8354, N8352, N8103);
nand NAND2 (N8355, N8340, N7430);
not NOT1 (N8356, N8355);
nand NAND2 (N8357, N8349, N253);
not NOT1 (N8358, N8357);
or OR2 (N8359, N8345, N8001);
and AND4 (N8360, N8354, N6738, N7169, N1489);
nor NOR2 (N8361, N8359, N6200);
buf BUF1 (N8362, N8348);
and AND2 (N8363, N8338, N7071);
buf BUF1 (N8364, N8351);
nand NAND3 (N8365, N8364, N4031, N6640);
and AND3 (N8366, N8362, N38, N1247);
or OR3 (N8367, N8366, N7718, N1695);
nand NAND3 (N8368, N8356, N6855, N3031);
and AND4 (N8369, N8361, N6661, N2310, N4543);
nor NOR4 (N8370, N8367, N5517, N6772, N407);
nand NAND4 (N8371, N8358, N3236, N7514, N4989);
xor XOR2 (N8372, N8370, N7642);
buf BUF1 (N8373, N8368);
xor XOR2 (N8374, N8371, N653);
nand NAND3 (N8375, N8365, N4974, N5078);
xor XOR2 (N8376, N8353, N7956);
nor NOR2 (N8377, N8373, N3638);
or OR2 (N8378, N8363, N5495);
not NOT1 (N8379, N8372);
or OR2 (N8380, N8377, N7179);
buf BUF1 (N8381, N8344);
nor NOR3 (N8382, N8369, N7076, N372);
buf BUF1 (N8383, N8379);
buf BUF1 (N8384, N8375);
buf BUF1 (N8385, N8374);
nor NOR2 (N8386, N8380, N3160);
xor XOR2 (N8387, N8386, N4821);
nor NOR2 (N8388, N8384, N1540);
xor XOR2 (N8389, N8385, N6379);
nand NAND3 (N8390, N8383, N8019, N1102);
and AND2 (N8391, N8360, N3165);
nor NOR3 (N8392, N8387, N6092, N7536);
or OR3 (N8393, N8389, N2257, N4189);
xor XOR2 (N8394, N8381, N2368);
nand NAND2 (N8395, N8391, N8075);
nor NOR2 (N8396, N8388, N2983);
not NOT1 (N8397, N8376);
buf BUF1 (N8398, N8395);
buf BUF1 (N8399, N8394);
nor NOR2 (N8400, N8399, N7288);
or OR4 (N8401, N8397, N7306, N2776, N1294);
nor NOR2 (N8402, N8396, N4314);
nor NOR3 (N8403, N8378, N1597, N5585);
xor XOR2 (N8404, N8390, N2984);
nor NOR3 (N8405, N8382, N7321, N2308);
nand NAND4 (N8406, N8400, N3977, N511, N7953);
not NOT1 (N8407, N8346);
nor NOR4 (N8408, N8403, N6224, N4448, N4604);
or OR4 (N8409, N8401, N3176, N7308, N7429);
buf BUF1 (N8410, N8405);
xor XOR2 (N8411, N8408, N8092);
or OR3 (N8412, N8393, N3863, N680);
xor XOR2 (N8413, N8409, N4528);
nand NAND4 (N8414, N8407, N5329, N1127, N589);
not NOT1 (N8415, N8398);
not NOT1 (N8416, N8410);
buf BUF1 (N8417, N8413);
nor NOR3 (N8418, N8412, N6745, N7551);
or OR4 (N8419, N8416, N5877, N7832, N7466);
not NOT1 (N8420, N8392);
buf BUF1 (N8421, N8404);
and AND3 (N8422, N8402, N2905, N3016);
not NOT1 (N8423, N8422);
nor NOR3 (N8424, N8411, N5875, N5140);
nor NOR3 (N8425, N8414, N4709, N1617);
xor XOR2 (N8426, N8421, N7922);
and AND3 (N8427, N8406, N4316, N6906);
not NOT1 (N8428, N8418);
nand NAND2 (N8429, N8428, N2051);
and AND3 (N8430, N8417, N6802, N7313);
nor NOR4 (N8431, N8420, N1643, N6635, N6619);
xor XOR2 (N8432, N8426, N2464);
nor NOR4 (N8433, N8429, N1099, N7694, N2928);
or OR2 (N8434, N8419, N1842);
nand NAND2 (N8435, N8425, N1645);
nor NOR2 (N8436, N8415, N2258);
nor NOR2 (N8437, N8424, N7838);
not NOT1 (N8438, N8430);
nand NAND4 (N8439, N8435, N7229, N6577, N6866);
or OR3 (N8440, N8427, N3935, N4011);
xor XOR2 (N8441, N8439, N4184);
nor NOR2 (N8442, N8423, N2010);
and AND2 (N8443, N8431, N2616);
nand NAND2 (N8444, N8443, N3872);
and AND4 (N8445, N8441, N2083, N440, N1925);
xor XOR2 (N8446, N8433, N290);
nand NAND4 (N8447, N8442, N4277, N7406, N7890);
xor XOR2 (N8448, N8434, N2150);
nand NAND2 (N8449, N8432, N7855);
buf BUF1 (N8450, N8448);
buf BUF1 (N8451, N8447);
xor XOR2 (N8452, N8451, N119);
xor XOR2 (N8453, N8445, N3655);
nor NOR4 (N8454, N8450, N6282, N2772, N627);
and AND2 (N8455, N8436, N7451);
xor XOR2 (N8456, N8438, N8187);
nand NAND2 (N8457, N8456, N3869);
or OR3 (N8458, N8440, N8234, N2002);
not NOT1 (N8459, N8452);
nand NAND4 (N8460, N8454, N7314, N5609, N6862);
or OR3 (N8461, N8437, N4570, N1704);
xor XOR2 (N8462, N8461, N967);
nand NAND3 (N8463, N8455, N8408, N1492);
and AND2 (N8464, N8460, N7244);
nand NAND2 (N8465, N8458, N2880);
not NOT1 (N8466, N8464);
buf BUF1 (N8467, N8459);
and AND2 (N8468, N8444, N3154);
xor XOR2 (N8469, N8453, N4323);
not NOT1 (N8470, N8469);
buf BUF1 (N8471, N8470);
and AND4 (N8472, N8462, N3440, N223, N5884);
and AND3 (N8473, N8465, N6617, N7054);
or OR3 (N8474, N8472, N4511, N7504);
buf BUF1 (N8475, N8467);
nor NOR3 (N8476, N8474, N1297, N1346);
buf BUF1 (N8477, N8475);
buf BUF1 (N8478, N8449);
and AND3 (N8479, N8466, N336, N7511);
xor XOR2 (N8480, N8446, N4591);
or OR3 (N8481, N8477, N2752, N3510);
not NOT1 (N8482, N8471);
buf BUF1 (N8483, N8476);
not NOT1 (N8484, N8473);
or OR4 (N8485, N8484, N3652, N949, N862);
xor XOR2 (N8486, N8468, N3481);
buf BUF1 (N8487, N8457);
buf BUF1 (N8488, N8479);
not NOT1 (N8489, N8488);
nor NOR3 (N8490, N8481, N3268, N1206);
not NOT1 (N8491, N8489);
or OR3 (N8492, N8486, N5445, N4964);
buf BUF1 (N8493, N8463);
xor XOR2 (N8494, N8492, N3650);
nor NOR3 (N8495, N8482, N5007, N5469);
xor XOR2 (N8496, N8493, N2071);
xor XOR2 (N8497, N8487, N4168);
and AND4 (N8498, N8494, N4193, N1872, N6857);
nor NOR2 (N8499, N8478, N5593);
nand NAND4 (N8500, N8491, N3013, N956, N504);
and AND3 (N8501, N8497, N896, N5776);
xor XOR2 (N8502, N8500, N7039);
or OR2 (N8503, N8496, N5158);
xor XOR2 (N8504, N8501, N496);
not NOT1 (N8505, N8480);
not NOT1 (N8506, N8499);
or OR2 (N8507, N8495, N1427);
or OR2 (N8508, N8498, N176);
and AND3 (N8509, N8508, N6544, N1059);
xor XOR2 (N8510, N8506, N4663);
and AND2 (N8511, N8507, N2435);
not NOT1 (N8512, N8504);
nand NAND2 (N8513, N8502, N3473);
xor XOR2 (N8514, N8511, N3567);
nor NOR4 (N8515, N8485, N5227, N3279, N3400);
xor XOR2 (N8516, N8503, N4726);
nor NOR3 (N8517, N8505, N4178, N4514);
nor NOR2 (N8518, N8512, N8121);
buf BUF1 (N8519, N8515);
buf BUF1 (N8520, N8518);
buf BUF1 (N8521, N8520);
not NOT1 (N8522, N8519);
not NOT1 (N8523, N8521);
nor NOR2 (N8524, N8509, N8092);
xor XOR2 (N8525, N8514, N437);
and AND2 (N8526, N8490, N4746);
nor NOR2 (N8527, N8517, N7432);
nand NAND3 (N8528, N8525, N4995, N930);
nand NAND4 (N8529, N8524, N4309, N4915, N1364);
nor NOR3 (N8530, N8513, N4840, N278);
nor NOR4 (N8531, N8522, N6943, N5393, N5318);
and AND4 (N8532, N8528, N6863, N4852, N7690);
nor NOR2 (N8533, N8532, N2911);
buf BUF1 (N8534, N8526);
xor XOR2 (N8535, N8527, N2198);
not NOT1 (N8536, N8510);
buf BUF1 (N8537, N8523);
nand NAND2 (N8538, N8516, N2100);
and AND3 (N8539, N8530, N5813, N7941);
buf BUF1 (N8540, N8538);
buf BUF1 (N8541, N8537);
and AND2 (N8542, N8529, N6073);
buf BUF1 (N8543, N8541);
or OR4 (N8544, N8531, N2331, N1480, N556);
xor XOR2 (N8545, N8540, N2752);
nor NOR4 (N8546, N8543, N7742, N4422, N1675);
not NOT1 (N8547, N8542);
xor XOR2 (N8548, N8533, N5670);
and AND3 (N8549, N8539, N7881, N5916);
and AND2 (N8550, N8544, N6877);
buf BUF1 (N8551, N8534);
buf BUF1 (N8552, N8550);
nor NOR4 (N8553, N8546, N2101, N5693, N967);
nand NAND4 (N8554, N8548, N7332, N6847, N5770);
and AND2 (N8555, N8554, N5543);
nor NOR4 (N8556, N8547, N1384, N7931, N2059);
buf BUF1 (N8557, N8553);
and AND2 (N8558, N8555, N247);
and AND2 (N8559, N8536, N8258);
nor NOR3 (N8560, N8559, N6597, N1482);
not NOT1 (N8561, N8535);
not NOT1 (N8562, N8558);
not NOT1 (N8563, N8560);
nand NAND4 (N8564, N8562, N757, N3415, N4302);
xor XOR2 (N8565, N8564, N2809);
nor NOR2 (N8566, N8483, N994);
and AND3 (N8567, N8552, N6654, N7400);
nor NOR4 (N8568, N8561, N2848, N5439, N1010);
nor NOR4 (N8569, N8556, N3053, N5389, N7807);
nand NAND4 (N8570, N8565, N449, N8225, N7236);
or OR3 (N8571, N8567, N2285, N7636);
or OR2 (N8572, N8568, N4586);
nor NOR3 (N8573, N8571, N3427, N5322);
not NOT1 (N8574, N8551);
nand NAND2 (N8575, N8569, N978);
not NOT1 (N8576, N8545);
xor XOR2 (N8577, N8563, N2809);
xor XOR2 (N8578, N8575, N3735);
and AND2 (N8579, N8549, N81);
not NOT1 (N8580, N8566);
xor XOR2 (N8581, N8574, N333);
buf BUF1 (N8582, N8557);
buf BUF1 (N8583, N8576);
xor XOR2 (N8584, N8580, N5610);
nand NAND3 (N8585, N8572, N8453, N6927);
not NOT1 (N8586, N8577);
xor XOR2 (N8587, N8579, N2870);
not NOT1 (N8588, N8570);
nand NAND2 (N8589, N8573, N7915);
xor XOR2 (N8590, N8578, N1205);
nand NAND3 (N8591, N8589, N3041, N1417);
buf BUF1 (N8592, N8584);
or OR3 (N8593, N8590, N1941, N7617);
nand NAND3 (N8594, N8588, N3268, N7332);
nand NAND2 (N8595, N8587, N1112);
nand NAND4 (N8596, N8582, N4861, N7763, N6278);
nand NAND4 (N8597, N8583, N3360, N3441, N7878);
nand NAND2 (N8598, N8586, N5263);
buf BUF1 (N8599, N8594);
or OR3 (N8600, N8599, N5430, N1648);
nor NOR4 (N8601, N8585, N7350, N6738, N1093);
and AND2 (N8602, N8600, N3392);
nor NOR4 (N8603, N8601, N5745, N465, N5);
or OR3 (N8604, N8597, N4254, N90);
and AND4 (N8605, N8581, N1273, N1447, N1809);
or OR4 (N8606, N8598, N2321, N4003, N8112);
not NOT1 (N8607, N8603);
nand NAND3 (N8608, N8602, N4112, N6537);
nand NAND3 (N8609, N8595, N1806, N4070);
or OR2 (N8610, N8609, N6858);
xor XOR2 (N8611, N8592, N4741);
nand NAND3 (N8612, N8606, N4094, N121);
buf BUF1 (N8613, N8611);
nand NAND4 (N8614, N8604, N6661, N4993, N8030);
buf BUF1 (N8615, N8613);
nand NAND4 (N8616, N8614, N1285, N1209, N90);
nor NOR2 (N8617, N8607, N3393);
nor NOR3 (N8618, N8612, N1168, N5314);
nand NAND4 (N8619, N8616, N1373, N3679, N5856);
nand NAND2 (N8620, N8596, N7995);
not NOT1 (N8621, N8619);
buf BUF1 (N8622, N8605);
nor NOR4 (N8623, N8621, N7925, N5691, N3493);
not NOT1 (N8624, N8620);
nor NOR2 (N8625, N8623, N420);
or OR4 (N8626, N8625, N6040, N4232, N588);
xor XOR2 (N8627, N8615, N2236);
nand NAND2 (N8628, N8593, N2561);
or OR2 (N8629, N8610, N6578);
and AND3 (N8630, N8617, N7390, N7737);
nor NOR4 (N8631, N8591, N499, N249, N2788);
not NOT1 (N8632, N8618);
xor XOR2 (N8633, N8627, N4614);
nand NAND2 (N8634, N8631, N6713);
xor XOR2 (N8635, N8626, N329);
xor XOR2 (N8636, N8633, N4235);
buf BUF1 (N8637, N8636);
nand NAND4 (N8638, N8608, N1661, N880, N6197);
buf BUF1 (N8639, N8628);
or OR4 (N8640, N8634, N6895, N2502, N3684);
buf BUF1 (N8641, N8624);
and AND3 (N8642, N8640, N7946, N5004);
or OR3 (N8643, N8637, N3034, N6831);
or OR4 (N8644, N8638, N7552, N5491, N1393);
and AND4 (N8645, N8629, N1288, N4746, N8182);
nand NAND3 (N8646, N8645, N174, N4578);
or OR4 (N8647, N8641, N2363, N7416, N3280);
nand NAND4 (N8648, N8642, N6124, N6031, N5949);
nand NAND2 (N8649, N8630, N8115);
nand NAND4 (N8650, N8644, N5306, N434, N5854);
buf BUF1 (N8651, N8632);
buf BUF1 (N8652, N8647);
buf BUF1 (N8653, N8648);
and AND3 (N8654, N8653, N1009, N7255);
nor NOR4 (N8655, N8649, N5128, N4452, N5275);
xor XOR2 (N8656, N8643, N4593);
nand NAND3 (N8657, N8652, N7959, N5566);
nand NAND3 (N8658, N8622, N8166, N5429);
buf BUF1 (N8659, N8646);
and AND3 (N8660, N8639, N8168, N2432);
nor NOR2 (N8661, N8651, N5373);
xor XOR2 (N8662, N8650, N7904);
not NOT1 (N8663, N8635);
nand NAND4 (N8664, N8660, N578, N2629, N5244);
or OR3 (N8665, N8662, N7888, N7765);
or OR4 (N8666, N8655, N5919, N7250, N7067);
and AND4 (N8667, N8657, N5049, N2758, N3171);
not NOT1 (N8668, N8665);
buf BUF1 (N8669, N8658);
or OR3 (N8670, N8664, N7351, N7580);
nand NAND2 (N8671, N8656, N7466);
or OR3 (N8672, N8668, N2240, N204);
or OR3 (N8673, N8659, N5355, N1968);
or OR2 (N8674, N8670, N1790);
and AND4 (N8675, N8673, N7580, N4877, N7976);
not NOT1 (N8676, N8666);
nand NAND4 (N8677, N8675, N3807, N7627, N7164);
nor NOR4 (N8678, N8663, N8228, N151, N4108);
or OR2 (N8679, N8676, N2245);
xor XOR2 (N8680, N8661, N277);
or OR2 (N8681, N8679, N2617);
and AND2 (N8682, N8654, N3268);
buf BUF1 (N8683, N8678);
xor XOR2 (N8684, N8669, N6117);
not NOT1 (N8685, N8683);
not NOT1 (N8686, N8681);
nand NAND2 (N8687, N8685, N3829);
and AND3 (N8688, N8680, N2655, N8642);
nor NOR3 (N8689, N8674, N2973, N5223);
or OR2 (N8690, N8687, N6986);
nand NAND4 (N8691, N8684, N2491, N6516, N1162);
buf BUF1 (N8692, N8672);
or OR4 (N8693, N8689, N5564, N1434, N8283);
or OR2 (N8694, N8691, N2846);
xor XOR2 (N8695, N8692, N151);
or OR4 (N8696, N8667, N2874, N6784, N744);
and AND3 (N8697, N8688, N4163, N7023);
or OR4 (N8698, N8696, N3686, N7465, N1093);
or OR4 (N8699, N8698, N2155, N7214, N6576);
xor XOR2 (N8700, N8695, N148);
not NOT1 (N8701, N8686);
not NOT1 (N8702, N8694);
and AND2 (N8703, N8697, N6327);
nor NOR4 (N8704, N8682, N7232, N2623, N612);
nand NAND4 (N8705, N8704, N1357, N8062, N3472);
nand NAND4 (N8706, N8693, N1719, N4961, N6366);
xor XOR2 (N8707, N8702, N8568);
and AND2 (N8708, N8701, N300);
xor XOR2 (N8709, N8707, N7832);
and AND2 (N8710, N8706, N834);
nor NOR4 (N8711, N8677, N627, N7325, N7674);
nor NOR3 (N8712, N8699, N4132, N48);
and AND2 (N8713, N8690, N3387);
nor NOR2 (N8714, N8708, N4995);
or OR4 (N8715, N8710, N6324, N1627, N49);
nand NAND2 (N8716, N8711, N6337);
not NOT1 (N8717, N8712);
or OR4 (N8718, N8703, N4243, N3303, N93);
buf BUF1 (N8719, N8716);
and AND4 (N8720, N8709, N4779, N5832, N8447);
not NOT1 (N8721, N8715);
nor NOR4 (N8722, N8671, N8174, N652, N4286);
buf BUF1 (N8723, N8718);
nor NOR2 (N8724, N8700, N6460);
not NOT1 (N8725, N8717);
and AND2 (N8726, N8714, N562);
nor NOR4 (N8727, N8720, N2468, N8483, N3915);
nor NOR3 (N8728, N8723, N7233, N4618);
or OR2 (N8729, N8722, N3876);
nor NOR2 (N8730, N8726, N6784);
xor XOR2 (N8731, N8719, N913);
not NOT1 (N8732, N8713);
not NOT1 (N8733, N8727);
buf BUF1 (N8734, N8729);
not NOT1 (N8735, N8728);
nor NOR2 (N8736, N8730, N1721);
nand NAND3 (N8737, N8725, N409, N6645);
and AND2 (N8738, N8705, N2252);
buf BUF1 (N8739, N8724);
not NOT1 (N8740, N8731);
not NOT1 (N8741, N8739);
not NOT1 (N8742, N8721);
and AND3 (N8743, N8741, N44, N1165);
xor XOR2 (N8744, N8735, N2662);
xor XOR2 (N8745, N8738, N885);
nor NOR3 (N8746, N8732, N3454, N7431);
nand NAND3 (N8747, N8744, N4510, N5115);
buf BUF1 (N8748, N8747);
nand NAND4 (N8749, N8740, N4854, N1442, N5393);
or OR4 (N8750, N8749, N3854, N8117, N8636);
nand NAND4 (N8751, N8734, N7027, N3355, N6421);
not NOT1 (N8752, N8746);
buf BUF1 (N8753, N8750);
nor NOR3 (N8754, N8733, N2022, N8300);
not NOT1 (N8755, N8753);
or OR4 (N8756, N8737, N1494, N1029, N1899);
nor NOR3 (N8757, N8743, N6893, N3626);
not NOT1 (N8758, N8751);
nand NAND2 (N8759, N8757, N3127);
and AND2 (N8760, N8745, N7994);
buf BUF1 (N8761, N8736);
not NOT1 (N8762, N8756);
xor XOR2 (N8763, N8758, N5986);
buf BUF1 (N8764, N8759);
or OR3 (N8765, N8763, N1363, N3421);
xor XOR2 (N8766, N8755, N5158);
nand NAND2 (N8767, N8748, N5282);
nand NAND3 (N8768, N8765, N381, N6217);
nand NAND4 (N8769, N8767, N3735, N8433, N1463);
not NOT1 (N8770, N8754);
xor XOR2 (N8771, N8768, N7082);
buf BUF1 (N8772, N8752);
nor NOR4 (N8773, N8742, N2283, N695, N1274);
or OR4 (N8774, N8772, N6903, N4310, N4227);
xor XOR2 (N8775, N8766, N4228);
and AND2 (N8776, N8769, N7729);
or OR4 (N8777, N8774, N202, N6038, N8735);
xor XOR2 (N8778, N8775, N6001);
and AND3 (N8779, N8776, N1638, N2520);
nor NOR2 (N8780, N8773, N7822);
nand NAND4 (N8781, N8760, N7731, N7252, N8183);
or OR4 (N8782, N8764, N6634, N745, N177);
buf BUF1 (N8783, N8781);
not NOT1 (N8784, N8780);
xor XOR2 (N8785, N8762, N6079);
xor XOR2 (N8786, N8777, N7003);
nor NOR2 (N8787, N8761, N434);
nand NAND3 (N8788, N8784, N8048, N7025);
and AND2 (N8789, N8779, N7319);
not NOT1 (N8790, N8787);
nand NAND4 (N8791, N8770, N6565, N6468, N3917);
and AND2 (N8792, N8786, N2137);
or OR4 (N8793, N8792, N6509, N8073, N62);
nand NAND4 (N8794, N8771, N6693, N5361, N3348);
buf BUF1 (N8795, N8794);
and AND3 (N8796, N8785, N4051, N174);
nor NOR4 (N8797, N8778, N6677, N5562, N5111);
nand NAND4 (N8798, N8789, N2538, N4833, N1575);
or OR3 (N8799, N8783, N3361, N4193);
buf BUF1 (N8800, N8788);
nand NAND2 (N8801, N8790, N6735);
nor NOR2 (N8802, N8795, N2107);
buf BUF1 (N8803, N8799);
nor NOR4 (N8804, N8798, N5545, N5995, N6324);
nand NAND3 (N8805, N8796, N6693, N2397);
or OR3 (N8806, N8803, N5239, N1223);
or OR3 (N8807, N8800, N6977, N1692);
buf BUF1 (N8808, N8802);
nor NOR4 (N8809, N8805, N810, N2348, N4989);
nor NOR4 (N8810, N8793, N7409, N1857, N3226);
nor NOR4 (N8811, N8806, N1778, N7439, N3272);
not NOT1 (N8812, N8808);
and AND4 (N8813, N8782, N6935, N227, N5589);
not NOT1 (N8814, N8804);
or OR2 (N8815, N8797, N5218);
not NOT1 (N8816, N8814);
xor XOR2 (N8817, N8816, N1201);
nand NAND2 (N8818, N8811, N3644);
nor NOR4 (N8819, N8791, N7373, N7176, N5781);
buf BUF1 (N8820, N8817);
nor NOR4 (N8821, N8820, N5433, N5734, N8784);
and AND3 (N8822, N8818, N4740, N240);
nor NOR4 (N8823, N8810, N6037, N4341, N3427);
xor XOR2 (N8824, N8815, N2074);
xor XOR2 (N8825, N8807, N3211);
xor XOR2 (N8826, N8801, N7335);
or OR3 (N8827, N8824, N4348, N3393);
or OR3 (N8828, N8822, N7125, N4166);
buf BUF1 (N8829, N8821);
or OR4 (N8830, N8829, N848, N8002, N1781);
and AND4 (N8831, N8830, N852, N7864, N5405);
nor NOR4 (N8832, N8828, N4374, N6200, N3618);
and AND3 (N8833, N8826, N8041, N4799);
nor NOR2 (N8834, N8825, N5619);
nor NOR2 (N8835, N8812, N7261);
not NOT1 (N8836, N8813);
or OR2 (N8837, N8836, N1153);
or OR4 (N8838, N8835, N4756, N5908, N5567);
buf BUF1 (N8839, N8823);
buf BUF1 (N8840, N8819);
buf BUF1 (N8841, N8839);
nand NAND4 (N8842, N8840, N4613, N1675, N6441);
buf BUF1 (N8843, N8841);
xor XOR2 (N8844, N8842, N6795);
buf BUF1 (N8845, N8843);
not NOT1 (N8846, N8837);
not NOT1 (N8847, N8809);
or OR2 (N8848, N8831, N5258);
or OR3 (N8849, N8845, N7402, N3839);
nor NOR3 (N8850, N8847, N3062, N2209);
buf BUF1 (N8851, N8848);
buf BUF1 (N8852, N8838);
nor NOR4 (N8853, N8851, N7762, N6374, N1136);
xor XOR2 (N8854, N8844, N7991);
or OR3 (N8855, N8834, N1308, N4808);
or OR3 (N8856, N8849, N7477, N4047);
buf BUF1 (N8857, N8855);
nand NAND2 (N8858, N8852, N6516);
or OR3 (N8859, N8832, N107, N8338);
xor XOR2 (N8860, N8854, N8043);
and AND4 (N8861, N8846, N6002, N6447, N7385);
not NOT1 (N8862, N8860);
buf BUF1 (N8863, N8850);
not NOT1 (N8864, N8858);
xor XOR2 (N8865, N8857, N5505);
or OR2 (N8866, N8853, N3618);
nor NOR3 (N8867, N8863, N2061, N4975);
or OR2 (N8868, N8856, N8861);
not NOT1 (N8869, N7921);
nand NAND3 (N8870, N8862, N8503, N1756);
xor XOR2 (N8871, N8865, N6094);
xor XOR2 (N8872, N8864, N722);
or OR3 (N8873, N8833, N4246, N3073);
and AND2 (N8874, N8859, N7571);
nor NOR4 (N8875, N8866, N1650, N648, N4532);
buf BUF1 (N8876, N8869);
not NOT1 (N8877, N8867);
xor XOR2 (N8878, N8877, N3751);
not NOT1 (N8879, N8878);
nor NOR2 (N8880, N8873, N6443);
or OR3 (N8881, N8870, N2931, N459);
xor XOR2 (N8882, N8875, N4884);
xor XOR2 (N8883, N8871, N1502);
buf BUF1 (N8884, N8876);
nand NAND3 (N8885, N8881, N6283, N2805);
nand NAND3 (N8886, N8880, N428, N4545);
xor XOR2 (N8887, N8882, N6337);
nand NAND3 (N8888, N8874, N1620, N1793);
buf BUF1 (N8889, N8883);
buf BUF1 (N8890, N8827);
nor NOR4 (N8891, N8889, N8241, N8539, N4334);
nand NAND3 (N8892, N8891, N3849, N2691);
or OR4 (N8893, N8888, N256, N1778, N4263);
and AND3 (N8894, N8890, N6261, N6344);
xor XOR2 (N8895, N8868, N348);
and AND2 (N8896, N8893, N6671);
nand NAND2 (N8897, N8885, N3401);
and AND4 (N8898, N8884, N5406, N1786, N2862);
xor XOR2 (N8899, N8892, N6735);
nand NAND2 (N8900, N8886, N5551);
buf BUF1 (N8901, N8900);
nor NOR3 (N8902, N8872, N4256, N4135);
or OR4 (N8903, N8899, N2212, N3200, N4130);
and AND2 (N8904, N8901, N3675);
nand NAND4 (N8905, N8894, N4119, N6122, N2483);
nor NOR2 (N8906, N8904, N3987);
xor XOR2 (N8907, N8903, N5995);
and AND2 (N8908, N8887, N2943);
nor NOR2 (N8909, N8897, N4179);
and AND2 (N8910, N8908, N6372);
buf BUF1 (N8911, N8905);
nand NAND3 (N8912, N8911, N937, N2890);
nor NOR3 (N8913, N8879, N255, N6758);
or OR4 (N8914, N8913, N825, N43, N6868);
and AND3 (N8915, N8910, N607, N6827);
nand NAND3 (N8916, N8898, N4368, N8803);
or OR4 (N8917, N8909, N1720, N7724, N3839);
and AND4 (N8918, N8902, N5587, N7052, N131);
not NOT1 (N8919, N8914);
and AND2 (N8920, N8907, N7476);
buf BUF1 (N8921, N8906);
not NOT1 (N8922, N8895);
xor XOR2 (N8923, N8920, N8200);
xor XOR2 (N8924, N8915, N3625);
nand NAND2 (N8925, N8919, N1459);
and AND4 (N8926, N8924, N1535, N2038, N8715);
not NOT1 (N8927, N8896);
buf BUF1 (N8928, N8923);
xor XOR2 (N8929, N8917, N1115);
buf BUF1 (N8930, N8918);
and AND2 (N8931, N8929, N5861);
or OR4 (N8932, N8922, N272, N8763, N8523);
nor NOR2 (N8933, N8927, N461);
buf BUF1 (N8934, N8926);
buf BUF1 (N8935, N8934);
nand NAND2 (N8936, N8930, N3209);
not NOT1 (N8937, N8933);
or OR4 (N8938, N8921, N2608, N8201, N8375);
not NOT1 (N8939, N8932);
or OR2 (N8940, N8931, N2073);
or OR3 (N8941, N8940, N7062, N2589);
buf BUF1 (N8942, N8941);
nor NOR3 (N8943, N8912, N7523, N3112);
and AND2 (N8944, N8942, N7632);
not NOT1 (N8945, N8936);
nand NAND2 (N8946, N8916, N7137);
buf BUF1 (N8947, N8928);
or OR4 (N8948, N8939, N6702, N8734, N7806);
or OR2 (N8949, N8944, N7843);
not NOT1 (N8950, N8935);
not NOT1 (N8951, N8946);
nand NAND2 (N8952, N8949, N1595);
nand NAND3 (N8953, N8943, N7232, N3167);
nand NAND4 (N8954, N8945, N5370, N90, N7502);
nor NOR4 (N8955, N8951, N4643, N4186, N6646);
xor XOR2 (N8956, N8947, N6084);
nand NAND4 (N8957, N8937, N4892, N7732, N8812);
nor NOR2 (N8958, N8925, N8549);
and AND4 (N8959, N8958, N1035, N7129, N2638);
nand NAND2 (N8960, N8959, N5301);
or OR3 (N8961, N8950, N2566, N4506);
xor XOR2 (N8962, N8948, N5800);
not NOT1 (N8963, N8954);
buf BUF1 (N8964, N8962);
nor NOR2 (N8965, N8963, N1689);
or OR3 (N8966, N8961, N540, N1497);
buf BUF1 (N8967, N8957);
nor NOR3 (N8968, N8956, N2579, N4660);
nand NAND4 (N8969, N8952, N8363, N5921, N8745);
nand NAND3 (N8970, N8965, N4044, N7705);
nand NAND4 (N8971, N8960, N2847, N2342, N6078);
not NOT1 (N8972, N8969);
xor XOR2 (N8973, N8953, N3162);
not NOT1 (N8974, N8970);
or OR3 (N8975, N8955, N5203, N7733);
not NOT1 (N8976, N8971);
xor XOR2 (N8977, N8966, N7060);
not NOT1 (N8978, N8977);
nand NAND3 (N8979, N8938, N8072, N6384);
nand NAND4 (N8980, N8974, N1971, N297, N5594);
and AND4 (N8981, N8978, N2072, N7837, N1011);
or OR4 (N8982, N8976, N3378, N3524, N1639);
or OR2 (N8983, N8975, N5232);
or OR3 (N8984, N8981, N5861, N2736);
not NOT1 (N8985, N8982);
not NOT1 (N8986, N8967);
buf BUF1 (N8987, N8964);
not NOT1 (N8988, N8980);
nor NOR3 (N8989, N8984, N4508, N5158);
not NOT1 (N8990, N8989);
or OR4 (N8991, N8985, N3733, N5044, N4196);
and AND2 (N8992, N8973, N7350);
and AND2 (N8993, N8988, N439);
or OR2 (N8994, N8987, N1789);
nand NAND2 (N8995, N8992, N4369);
buf BUF1 (N8996, N8983);
nor NOR4 (N8997, N8979, N5583, N4351, N4555);
nand NAND2 (N8998, N8968, N8688);
nand NAND3 (N8999, N8972, N5232, N5850);
nand NAND2 (N9000, N8999, N6003);
nor NOR2 (N9001, N8997, N886);
nand NAND3 (N9002, N8995, N7934, N72);
xor XOR2 (N9003, N8993, N4307);
not NOT1 (N9004, N9000);
nand NAND2 (N9005, N8990, N6909);
nor NOR3 (N9006, N8994, N5991, N8438);
nand NAND3 (N9007, N9004, N752, N658);
nor NOR2 (N9008, N9005, N6004);
and AND3 (N9009, N8996, N1893, N522);
not NOT1 (N9010, N9006);
or OR4 (N9011, N9008, N3971, N2730, N278);
nor NOR3 (N9012, N9001, N3620, N3171);
or OR4 (N9013, N9002, N6902, N4510, N8500);
xor XOR2 (N9014, N8998, N3114);
or OR4 (N9015, N8986, N2185, N2080, N5547);
xor XOR2 (N9016, N9015, N3619);
or OR2 (N9017, N9012, N1578);
not NOT1 (N9018, N9007);
nor NOR2 (N9019, N9016, N6060);
and AND4 (N9020, N9013, N2977, N969, N5049);
nor NOR4 (N9021, N9019, N960, N8918, N4645);
xor XOR2 (N9022, N9018, N3029);
buf BUF1 (N9023, N9011);
nor NOR4 (N9024, N9014, N4112, N3263, N7720);
nand NAND3 (N9025, N9024, N7651, N5688);
and AND2 (N9026, N9009, N6411);
and AND3 (N9027, N9010, N3093, N8176);
nor NOR2 (N9028, N9027, N5884);
nand NAND2 (N9029, N9025, N4625);
not NOT1 (N9030, N9023);
xor XOR2 (N9031, N9029, N2746);
nor NOR3 (N9032, N9026, N3485, N250);
not NOT1 (N9033, N9017);
not NOT1 (N9034, N9003);
not NOT1 (N9035, N9033);
nand NAND3 (N9036, N9031, N5974, N8719);
and AND3 (N9037, N9032, N3791, N3706);
buf BUF1 (N9038, N9022);
or OR3 (N9039, N8991, N4112, N5005);
not NOT1 (N9040, N9030);
nand NAND3 (N9041, N9039, N887, N204);
nor NOR2 (N9042, N9040, N7735);
nor NOR4 (N9043, N9021, N2567, N3775, N7799);
and AND3 (N9044, N9034, N4075, N6796);
nor NOR2 (N9045, N9037, N1039);
and AND4 (N9046, N9038, N5685, N288, N4644);
and AND2 (N9047, N9044, N5904);
buf BUF1 (N9048, N9028);
nand NAND3 (N9049, N9042, N7004, N5177);
xor XOR2 (N9050, N9043, N4753);
nor NOR2 (N9051, N9046, N2961);
nand NAND4 (N9052, N9020, N6360, N2481, N3457);
buf BUF1 (N9053, N9049);
or OR3 (N9054, N9041, N5030, N5811);
and AND4 (N9055, N9052, N7600, N5980, N339);
or OR3 (N9056, N9035, N3812, N4069);
and AND2 (N9057, N9050, N7367);
nor NOR3 (N9058, N9055, N654, N4219);
nor NOR4 (N9059, N9045, N5932, N2550, N5260);
xor XOR2 (N9060, N9057, N2114);
or OR4 (N9061, N9048, N1792, N6760, N625);
not NOT1 (N9062, N9036);
xor XOR2 (N9063, N9051, N1942);
nand NAND2 (N9064, N9060, N8509);
or OR3 (N9065, N9054, N3594, N4151);
not NOT1 (N9066, N9058);
buf BUF1 (N9067, N9053);
buf BUF1 (N9068, N9064);
nand NAND3 (N9069, N9059, N8178, N6837);
xor XOR2 (N9070, N9056, N6978);
xor XOR2 (N9071, N9067, N7091);
buf BUF1 (N9072, N9068);
or OR3 (N9073, N9072, N301, N8464);
or OR4 (N9074, N9062, N9024, N6162, N2105);
or OR2 (N9075, N9073, N6113);
nor NOR4 (N9076, N9066, N1928, N2261, N3648);
xor XOR2 (N9077, N9076, N4813);
not NOT1 (N9078, N9065);
buf BUF1 (N9079, N9071);
nor NOR2 (N9080, N9063, N3808);
xor XOR2 (N9081, N9074, N161);
buf BUF1 (N9082, N9081);
xor XOR2 (N9083, N9075, N4681);
buf BUF1 (N9084, N9083);
or OR3 (N9085, N9061, N7731, N7732);
nor NOR3 (N9086, N9084, N2939, N3419);
nor NOR4 (N9087, N9077, N4489, N2200, N7743);
buf BUF1 (N9088, N9087);
and AND2 (N9089, N9078, N4899);
and AND4 (N9090, N9047, N2853, N4592, N3658);
buf BUF1 (N9091, N9082);
or OR4 (N9092, N9070, N2686, N8650, N1538);
xor XOR2 (N9093, N9080, N8690);
and AND4 (N9094, N9086, N2691, N6287, N7019);
buf BUF1 (N9095, N9090);
and AND2 (N9096, N9088, N2555);
nor NOR3 (N9097, N9095, N4313, N6664);
and AND4 (N9098, N9094, N8179, N5346, N454);
and AND3 (N9099, N9096, N1723, N4273);
or OR4 (N9100, N9099, N7341, N4168, N6772);
xor XOR2 (N9101, N9092, N6374);
buf BUF1 (N9102, N9100);
xor XOR2 (N9103, N9085, N5029);
or OR2 (N9104, N9098, N8402);
nand NAND3 (N9105, N9101, N6702, N8296);
buf BUF1 (N9106, N9102);
or OR2 (N9107, N9091, N6316);
not NOT1 (N9108, N9107);
nor NOR4 (N9109, N9104, N7872, N8083, N6794);
buf BUF1 (N9110, N9069);
or OR3 (N9111, N9089, N1324, N8904);
and AND2 (N9112, N9093, N890);
not NOT1 (N9113, N9105);
nor NOR4 (N9114, N9110, N8661, N4637, N5479);
nor NOR3 (N9115, N9079, N6673, N3526);
or OR4 (N9116, N9111, N7747, N2084, N5071);
or OR3 (N9117, N9114, N2929, N2947);
nor NOR2 (N9118, N9116, N7769);
nand NAND3 (N9119, N9115, N4054, N5202);
xor XOR2 (N9120, N9097, N4120);
xor XOR2 (N9121, N9120, N7232);
xor XOR2 (N9122, N9117, N6362);
xor XOR2 (N9123, N9106, N2122);
and AND2 (N9124, N9123, N2140);
xor XOR2 (N9125, N9121, N1668);
nor NOR2 (N9126, N9119, N8510);
nand NAND4 (N9127, N9118, N2724, N6898, N185);
or OR4 (N9128, N9109, N6087, N8561, N5749);
xor XOR2 (N9129, N9112, N304);
and AND2 (N9130, N9125, N4910);
and AND3 (N9131, N9128, N2642, N4000);
xor XOR2 (N9132, N9130, N4813);
buf BUF1 (N9133, N9132);
or OR2 (N9134, N9113, N2191);
nor NOR2 (N9135, N9126, N2351);
or OR2 (N9136, N9124, N560);
nand NAND2 (N9137, N9135, N1673);
xor XOR2 (N9138, N9108, N6738);
or OR4 (N9139, N9129, N5373, N6980, N5992);
nand NAND3 (N9140, N9133, N181, N7910);
not NOT1 (N9141, N9136);
or OR4 (N9142, N9141, N7969, N8173, N4563);
not NOT1 (N9143, N9140);
nor NOR2 (N9144, N9134, N3560);
xor XOR2 (N9145, N9127, N4897);
xor XOR2 (N9146, N9144, N8809);
xor XOR2 (N9147, N9143, N5004);
and AND3 (N9148, N9131, N3303, N3329);
nor NOR3 (N9149, N9103, N5532, N6094);
xor XOR2 (N9150, N9149, N1303);
or OR4 (N9151, N9148, N3106, N6740, N3875);
nand NAND2 (N9152, N9142, N301);
nor NOR2 (N9153, N9138, N4986);
not NOT1 (N9154, N9150);
not NOT1 (N9155, N9145);
nor NOR4 (N9156, N9147, N3620, N6892, N7097);
nor NOR2 (N9157, N9154, N8947);
buf BUF1 (N9158, N9139);
and AND4 (N9159, N9137, N7239, N410, N5421);
buf BUF1 (N9160, N9155);
not NOT1 (N9161, N9156);
xor XOR2 (N9162, N9160, N4567);
nand NAND2 (N9163, N9152, N1361);
or OR2 (N9164, N9163, N1877);
or OR2 (N9165, N9162, N2841);
nor NOR2 (N9166, N9161, N6962);
xor XOR2 (N9167, N9164, N2435);
xor XOR2 (N9168, N9122, N648);
nor NOR4 (N9169, N9167, N1141, N6669, N1019);
xor XOR2 (N9170, N9157, N8645);
buf BUF1 (N9171, N9165);
not NOT1 (N9172, N9158);
buf BUF1 (N9173, N9146);
nor NOR4 (N9174, N9168, N1936, N3431, N3040);
not NOT1 (N9175, N9173);
nor NOR3 (N9176, N9174, N6642, N1003);
nand NAND2 (N9177, N9171, N3088);
not NOT1 (N9178, N9176);
nor NOR4 (N9179, N9178, N2012, N1248, N9132);
buf BUF1 (N9180, N9177);
xor XOR2 (N9181, N9175, N7341);
nor NOR2 (N9182, N9151, N5845);
not NOT1 (N9183, N9180);
and AND4 (N9184, N9179, N4028, N5395, N8751);
nand NAND2 (N9185, N9170, N117);
nor NOR2 (N9186, N9169, N3182);
and AND2 (N9187, N9153, N8963);
buf BUF1 (N9188, N9181);
nand NAND3 (N9189, N9183, N3860, N4992);
not NOT1 (N9190, N9159);
or OR4 (N9191, N9187, N3036, N8994, N7434);
or OR4 (N9192, N9166, N6663, N6121, N5203);
and AND4 (N9193, N9186, N3233, N5703, N2092);
buf BUF1 (N9194, N9192);
nand NAND4 (N9195, N9190, N6032, N5417, N2788);
nand NAND2 (N9196, N9195, N7316);
and AND4 (N9197, N9184, N6735, N2405, N6417);
and AND2 (N9198, N9189, N6233);
buf BUF1 (N9199, N9196);
not NOT1 (N9200, N9198);
buf BUF1 (N9201, N9188);
nor NOR4 (N9202, N9191, N8493, N5325, N1079);
xor XOR2 (N9203, N9194, N7855);
nor NOR4 (N9204, N9200, N6043, N8750, N7136);
nand NAND2 (N9205, N9199, N5176);
or OR3 (N9206, N9172, N4913, N6374);
not NOT1 (N9207, N9197);
and AND4 (N9208, N9193, N3829, N3536, N880);
or OR3 (N9209, N9202, N1386, N5387);
buf BUF1 (N9210, N9201);
nand NAND2 (N9211, N9206, N655);
or OR4 (N9212, N9205, N5901, N3658, N7477);
and AND4 (N9213, N9182, N7327, N494, N7805);
not NOT1 (N9214, N9212);
not NOT1 (N9215, N9204);
buf BUF1 (N9216, N9208);
buf BUF1 (N9217, N9216);
or OR3 (N9218, N9207, N1802, N1028);
xor XOR2 (N9219, N9209, N5201);
nor NOR3 (N9220, N9213, N8725, N5781);
nor NOR3 (N9221, N9218, N1384, N5185);
xor XOR2 (N9222, N9220, N7933);
or OR4 (N9223, N9217, N3912, N5171, N5052);
xor XOR2 (N9224, N9210, N4936);
or OR4 (N9225, N9203, N5160, N640, N306);
nor NOR4 (N9226, N9222, N8993, N2114, N3597);
not NOT1 (N9227, N9221);
or OR4 (N9228, N9225, N5660, N5869, N7586);
nor NOR4 (N9229, N9211, N4272, N6383, N1575);
not NOT1 (N9230, N9224);
nor NOR4 (N9231, N9215, N8462, N4466, N953);
and AND4 (N9232, N9229, N6165, N3583, N6644);
or OR3 (N9233, N9232, N9002, N8477);
not NOT1 (N9234, N9214);
not NOT1 (N9235, N9231);
buf BUF1 (N9236, N9219);
and AND4 (N9237, N9236, N2980, N5111, N7970);
and AND3 (N9238, N9234, N8089, N1775);
and AND4 (N9239, N9230, N605, N2999, N6342);
or OR4 (N9240, N9228, N725, N3654, N2594);
xor XOR2 (N9241, N9235, N5630);
nor NOR4 (N9242, N9226, N3487, N6958, N6349);
not NOT1 (N9243, N9233);
and AND2 (N9244, N9241, N5640);
nand NAND2 (N9245, N9243, N665);
or OR3 (N9246, N9244, N1438, N7515);
nor NOR2 (N9247, N9246, N1469);
nand NAND2 (N9248, N9185, N7720);
not NOT1 (N9249, N9238);
buf BUF1 (N9250, N9248);
and AND4 (N9251, N9247, N300, N5112, N3184);
xor XOR2 (N9252, N9239, N4572);
or OR4 (N9253, N9242, N725, N7065, N6645);
nand NAND4 (N9254, N9250, N3687, N4539, N3843);
not NOT1 (N9255, N9240);
and AND4 (N9256, N9254, N8826, N3213, N5754);
or OR3 (N9257, N9253, N1192, N6970);
xor XOR2 (N9258, N9245, N6279);
nor NOR3 (N9259, N9237, N8768, N4682);
not NOT1 (N9260, N9252);
and AND2 (N9261, N9256, N7298);
or OR4 (N9262, N9255, N7448, N8440, N6253);
buf BUF1 (N9263, N9262);
buf BUF1 (N9264, N9263);
not NOT1 (N9265, N9223);
and AND2 (N9266, N9260, N4396);
buf BUF1 (N9267, N9259);
and AND3 (N9268, N9267, N4765, N5965);
buf BUF1 (N9269, N9227);
nand NAND3 (N9270, N9258, N7463, N7148);
nor NOR2 (N9271, N9257, N6026);
xor XOR2 (N9272, N9261, N4152);
or OR2 (N9273, N9268, N1731);
nor NOR2 (N9274, N9251, N6281);
nor NOR4 (N9275, N9265, N7960, N3222, N2539);
or OR2 (N9276, N9275, N7316);
nor NOR2 (N9277, N9270, N2290);
nor NOR3 (N9278, N9269, N6700, N8791);
buf BUF1 (N9279, N9278);
or OR3 (N9280, N9276, N2896, N4460);
and AND3 (N9281, N9271, N8991, N5444);
and AND4 (N9282, N9264, N3887, N8476, N3904);
not NOT1 (N9283, N9272);
and AND3 (N9284, N9283, N5588, N5882);
nor NOR4 (N9285, N9266, N7826, N8644, N8669);
buf BUF1 (N9286, N9284);
not NOT1 (N9287, N9280);
nand NAND3 (N9288, N9281, N2412, N7286);
nor NOR3 (N9289, N9286, N7512, N3441);
buf BUF1 (N9290, N9287);
xor XOR2 (N9291, N9285, N7886);
not NOT1 (N9292, N9289);
xor XOR2 (N9293, N9277, N1072);
xor XOR2 (N9294, N9274, N2603);
buf BUF1 (N9295, N9292);
not NOT1 (N9296, N9290);
or OR2 (N9297, N9288, N6435);
buf BUF1 (N9298, N9295);
xor XOR2 (N9299, N9291, N9209);
and AND2 (N9300, N9294, N769);
nand NAND3 (N9301, N9298, N6122, N7425);
or OR4 (N9302, N9249, N5861, N3772, N5730);
not NOT1 (N9303, N9279);
xor XOR2 (N9304, N9296, N894);
xor XOR2 (N9305, N9302, N5681);
and AND2 (N9306, N9299, N5375);
and AND3 (N9307, N9301, N3622, N8961);
not NOT1 (N9308, N9307);
nand NAND2 (N9309, N9293, N7829);
xor XOR2 (N9310, N9303, N1991);
xor XOR2 (N9311, N9305, N7757);
nand NAND2 (N9312, N9273, N3725);
xor XOR2 (N9313, N9309, N1543);
nand NAND2 (N9314, N9306, N1900);
or OR4 (N9315, N9297, N7889, N5088, N5492);
or OR4 (N9316, N9300, N6632, N7507, N1054);
not NOT1 (N9317, N9310);
and AND2 (N9318, N9304, N34);
nor NOR3 (N9319, N9312, N7998, N714);
not NOT1 (N9320, N9317);
xor XOR2 (N9321, N9311, N279);
nand NAND4 (N9322, N9318, N884, N3711, N735);
and AND4 (N9323, N9308, N4860, N1106, N6516);
nand NAND4 (N9324, N9282, N8234, N1052, N6042);
buf BUF1 (N9325, N9316);
and AND4 (N9326, N9313, N11, N1578, N7307);
buf BUF1 (N9327, N9315);
nor NOR2 (N9328, N9314, N963);
xor XOR2 (N9329, N9323, N2663);
nor NOR3 (N9330, N9322, N7300, N1752);
xor XOR2 (N9331, N9326, N1502);
and AND3 (N9332, N9328, N5665, N2424);
xor XOR2 (N9333, N9325, N2928);
and AND2 (N9334, N9332, N4633);
not NOT1 (N9335, N9320);
and AND4 (N9336, N9321, N3199, N2360, N5922);
xor XOR2 (N9337, N9331, N4696);
and AND2 (N9338, N9333, N7285);
and AND3 (N9339, N9330, N2397, N3597);
nor NOR3 (N9340, N9338, N918, N4521);
nand NAND3 (N9341, N9324, N7046, N6415);
buf BUF1 (N9342, N9329);
nand NAND4 (N9343, N9336, N2418, N5217, N727);
nand NAND4 (N9344, N9335, N6158, N9094, N6856);
not NOT1 (N9345, N9327);
not NOT1 (N9346, N9340);
xor XOR2 (N9347, N9344, N4379);
or OR4 (N9348, N9319, N8748, N7313, N739);
buf BUF1 (N9349, N9342);
nand NAND2 (N9350, N9337, N5713);
nor NOR2 (N9351, N9334, N5720);
nand NAND2 (N9352, N9341, N1146);
and AND4 (N9353, N9348, N2930, N47, N5528);
and AND3 (N9354, N9343, N2966, N1094);
nor NOR2 (N9355, N9350, N2813);
buf BUF1 (N9356, N9353);
buf BUF1 (N9357, N9345);
buf BUF1 (N9358, N9351);
xor XOR2 (N9359, N9358, N8269);
nand NAND4 (N9360, N9346, N7910, N8818, N5096);
buf BUF1 (N9361, N9355);
nor NOR3 (N9362, N9339, N8332, N8318);
nor NOR3 (N9363, N9356, N2989, N9237);
buf BUF1 (N9364, N9361);
and AND2 (N9365, N9347, N2694);
and AND2 (N9366, N9357, N4866);
xor XOR2 (N9367, N9354, N4466);
or OR3 (N9368, N9367, N8278, N2498);
nor NOR4 (N9369, N9362, N3884, N4851, N4808);
not NOT1 (N9370, N9363);
or OR3 (N9371, N9365, N7900, N4187);
or OR4 (N9372, N9368, N6041, N8990, N1791);
nor NOR3 (N9373, N9360, N1370, N4497);
or OR2 (N9374, N9369, N2832);
buf BUF1 (N9375, N9366);
and AND2 (N9376, N9373, N4306);
or OR4 (N9377, N9370, N3168, N2446, N2913);
nand NAND2 (N9378, N9349, N4444);
buf BUF1 (N9379, N9364);
nand NAND3 (N9380, N9371, N1090, N821);
not NOT1 (N9381, N9372);
xor XOR2 (N9382, N9359, N98);
not NOT1 (N9383, N9381);
buf BUF1 (N9384, N9375);
nor NOR3 (N9385, N9352, N8419, N474);
buf BUF1 (N9386, N9380);
not NOT1 (N9387, N9376);
and AND3 (N9388, N9387, N4933, N3723);
or OR4 (N9389, N9385, N3196, N7938, N2934);
xor XOR2 (N9390, N9386, N7098);
buf BUF1 (N9391, N9383);
not NOT1 (N9392, N9378);
and AND2 (N9393, N9384, N5081);
xor XOR2 (N9394, N9377, N5898);
not NOT1 (N9395, N9389);
and AND3 (N9396, N9394, N5254, N1142);
xor XOR2 (N9397, N9392, N3824);
or OR4 (N9398, N9393, N6147, N7832, N9329);
or OR2 (N9399, N9391, N989);
nor NOR3 (N9400, N9374, N6152, N5150);
xor XOR2 (N9401, N9390, N5433);
xor XOR2 (N9402, N9396, N2384);
xor XOR2 (N9403, N9382, N4047);
buf BUF1 (N9404, N9397);
xor XOR2 (N9405, N9388, N1969);
xor XOR2 (N9406, N9401, N285);
or OR4 (N9407, N9395, N6546, N2766, N7215);
not NOT1 (N9408, N9379);
not NOT1 (N9409, N9398);
or OR4 (N9410, N9402, N7784, N4105, N8332);
nor NOR2 (N9411, N9407, N8492);
or OR3 (N9412, N9411, N5757, N3088);
or OR4 (N9413, N9409, N4425, N3971, N479);
buf BUF1 (N9414, N9406);
nor NOR4 (N9415, N9404, N3985, N9228, N920);
nand NAND4 (N9416, N9399, N934, N1004, N3540);
nor NOR2 (N9417, N9400, N5785);
and AND4 (N9418, N9417, N6234, N380, N929);
nor NOR2 (N9419, N9403, N4213);
not NOT1 (N9420, N9408);
not NOT1 (N9421, N9413);
or OR3 (N9422, N9412, N5748, N7879);
not NOT1 (N9423, N9414);
buf BUF1 (N9424, N9421);
nand NAND2 (N9425, N9420, N6345);
not NOT1 (N9426, N9418);
and AND3 (N9427, N9405, N321, N2461);
buf BUF1 (N9428, N9410);
or OR4 (N9429, N9424, N1505, N603, N747);
or OR2 (N9430, N9425, N8133);
buf BUF1 (N9431, N9430);
nor NOR4 (N9432, N9423, N420, N4265, N6087);
nand NAND4 (N9433, N9429, N4397, N7635, N4785);
not NOT1 (N9434, N9433);
xor XOR2 (N9435, N9415, N831);
xor XOR2 (N9436, N9416, N7219);
buf BUF1 (N9437, N9422);
not NOT1 (N9438, N9428);
nor NOR4 (N9439, N9419, N5496, N802, N7266);
not NOT1 (N9440, N9434);
nand NAND2 (N9441, N9437, N6857);
or OR4 (N9442, N9426, N3510, N2915, N980);
nor NOR3 (N9443, N9440, N1049, N3926);
nand NAND3 (N9444, N9439, N2059, N9425);
nor NOR4 (N9445, N9435, N5267, N6182, N5148);
nor NOR3 (N9446, N9431, N7340, N1535);
xor XOR2 (N9447, N9427, N3753);
and AND2 (N9448, N9432, N4000);
nand NAND4 (N9449, N9447, N841, N1581, N3504);
nor NOR2 (N9450, N9441, N4430);
and AND4 (N9451, N9450, N1371, N9329, N1651);
or OR4 (N9452, N9449, N618, N7402, N5493);
buf BUF1 (N9453, N9438);
nand NAND4 (N9454, N9445, N5749, N3409, N8608);
not NOT1 (N9455, N9444);
nor NOR2 (N9456, N9455, N4708);
not NOT1 (N9457, N9456);
and AND3 (N9458, N9453, N8548, N7532);
and AND2 (N9459, N9443, N4828);
xor XOR2 (N9460, N9459, N8829);
nor NOR3 (N9461, N9454, N6931, N6540);
xor XOR2 (N9462, N9436, N3437);
xor XOR2 (N9463, N9458, N1886);
not NOT1 (N9464, N9462);
nand NAND2 (N9465, N9442, N9037);
buf BUF1 (N9466, N9446);
nand NAND3 (N9467, N9464, N9078, N9113);
or OR2 (N9468, N9448, N5155);
buf BUF1 (N9469, N9465);
and AND4 (N9470, N9457, N6408, N7684, N4229);
buf BUF1 (N9471, N9470);
not NOT1 (N9472, N9469);
nand NAND4 (N9473, N9451, N6824, N1864, N488);
nand NAND2 (N9474, N9467, N9319);
nand NAND2 (N9475, N9460, N7533);
not NOT1 (N9476, N9452);
and AND2 (N9477, N9472, N6677);
and AND2 (N9478, N9475, N5312);
nand NAND3 (N9479, N9474, N2885, N4411);
and AND2 (N9480, N9479, N6487);
nor NOR4 (N9481, N9476, N3730, N318, N558);
or OR4 (N9482, N9478, N4545, N9034, N275);
nand NAND3 (N9483, N9482, N1096, N7946);
not NOT1 (N9484, N9463);
nor NOR4 (N9485, N9483, N4616, N1266, N1651);
or OR4 (N9486, N9477, N493, N8792, N6962);
nand NAND2 (N9487, N9473, N9052);
buf BUF1 (N9488, N9461);
not NOT1 (N9489, N9486);
xor XOR2 (N9490, N9468, N8259);
and AND4 (N9491, N9490, N5747, N7184, N8144);
xor XOR2 (N9492, N9491, N301);
nand NAND3 (N9493, N9471, N3551, N1484);
xor XOR2 (N9494, N9489, N8657);
or OR3 (N9495, N9480, N7215, N6215);
and AND2 (N9496, N9466, N110);
not NOT1 (N9497, N9484);
xor XOR2 (N9498, N9492, N8912);
or OR2 (N9499, N9494, N5469);
nand NAND4 (N9500, N9495, N5160, N6809, N5048);
xor XOR2 (N9501, N9481, N1810);
nand NAND2 (N9502, N9500, N1786);
not NOT1 (N9503, N9497);
or OR4 (N9504, N9502, N3677, N8927, N9460);
and AND2 (N9505, N9504, N69);
not NOT1 (N9506, N9487);
nor NOR4 (N9507, N9488, N7623, N6807, N9151);
and AND3 (N9508, N9498, N7745, N7634);
or OR2 (N9509, N9508, N4443);
not NOT1 (N9510, N9485);
xor XOR2 (N9511, N9499, N7051);
not NOT1 (N9512, N9506);
and AND3 (N9513, N9503, N3909, N4176);
nand NAND2 (N9514, N9496, N595);
and AND3 (N9515, N9511, N4885, N3024);
and AND4 (N9516, N9493, N7004, N7016, N3762);
and AND4 (N9517, N9512, N8650, N8830, N8644);
and AND3 (N9518, N9515, N6133, N2475);
or OR2 (N9519, N9517, N6372);
and AND3 (N9520, N9510, N5039, N4114);
nand NAND4 (N9521, N9519, N4240, N8724, N390);
xor XOR2 (N9522, N9501, N1884);
nand NAND4 (N9523, N9513, N7022, N6258, N4430);
nor NOR2 (N9524, N9514, N4273);
or OR3 (N9525, N9505, N735, N7259);
or OR2 (N9526, N9522, N362);
or OR2 (N9527, N9523, N6204);
xor XOR2 (N9528, N9527, N4151);
and AND4 (N9529, N9516, N2411, N4913, N3158);
nand NAND3 (N9530, N9525, N7544, N6046);
nor NOR4 (N9531, N9524, N7676, N1784, N991);
buf BUF1 (N9532, N9518);
not NOT1 (N9533, N9507);
and AND3 (N9534, N9520, N8173, N2868);
and AND2 (N9535, N9530, N5611);
nor NOR3 (N9536, N9533, N2905, N895);
and AND3 (N9537, N9521, N2522, N359);
xor XOR2 (N9538, N9526, N6623);
nor NOR3 (N9539, N9534, N5187, N2272);
buf BUF1 (N9540, N9529);
nand NAND4 (N9541, N9509, N6358, N5853, N6325);
nand NAND4 (N9542, N9538, N8819, N9426, N243);
buf BUF1 (N9543, N9541);
not NOT1 (N9544, N9537);
or OR4 (N9545, N9544, N8221, N8459, N8051);
nor NOR4 (N9546, N9531, N5078, N810, N6413);
nand NAND2 (N9547, N9539, N5663);
and AND3 (N9548, N9545, N709, N4536);
not NOT1 (N9549, N9532);
buf BUF1 (N9550, N9540);
or OR2 (N9551, N9536, N4375);
nand NAND4 (N9552, N9546, N6713, N7523, N8890);
nor NOR4 (N9553, N9548, N3182, N4923, N9085);
not NOT1 (N9554, N9528);
and AND2 (N9555, N9553, N6040);
and AND2 (N9556, N9543, N2792);
nand NAND3 (N9557, N9555, N3994, N4972);
buf BUF1 (N9558, N9542);
not NOT1 (N9559, N9547);
nand NAND3 (N9560, N9551, N5198, N5203);
or OR3 (N9561, N9554, N331, N2895);
not NOT1 (N9562, N9552);
nor NOR4 (N9563, N9535, N6760, N385, N6625);
buf BUF1 (N9564, N9559);
or OR4 (N9565, N9558, N4805, N5074, N6214);
not NOT1 (N9566, N9549);
nor NOR3 (N9567, N9556, N3747, N7420);
and AND3 (N9568, N9567, N599, N204);
nand NAND4 (N9569, N9564, N6131, N5945, N1922);
xor XOR2 (N9570, N9568, N6916);
or OR2 (N9571, N9563, N4630);
nand NAND3 (N9572, N9566, N6877, N57);
and AND4 (N9573, N9557, N5416, N5302, N6720);
buf BUF1 (N9574, N9569);
nor NOR3 (N9575, N9570, N9038, N6420);
nand NAND4 (N9576, N9561, N1867, N5274, N5046);
nor NOR2 (N9577, N9574, N4818);
xor XOR2 (N9578, N9562, N4822);
nor NOR2 (N9579, N9572, N3790);
nor NOR3 (N9580, N9550, N6171, N7987);
nor NOR3 (N9581, N9578, N1572, N215);
nand NAND4 (N9582, N9581, N976, N9053, N8588);
not NOT1 (N9583, N9576);
and AND4 (N9584, N9580, N9565, N2723, N2015);
xor XOR2 (N9585, N1996, N1747);
buf BUF1 (N9586, N9575);
or OR3 (N9587, N9584, N2880, N7521);
nand NAND2 (N9588, N9585, N1521);
and AND3 (N9589, N9560, N9497, N3399);
nand NAND4 (N9590, N9571, N1784, N4598, N201);
not NOT1 (N9591, N9587);
nor NOR4 (N9592, N9586, N121, N2036, N8140);
and AND3 (N9593, N9590, N4327, N8691);
and AND4 (N9594, N9577, N4930, N6929, N4077);
nor NOR4 (N9595, N9594, N8894, N4079, N6589);
xor XOR2 (N9596, N9573, N9009);
xor XOR2 (N9597, N9588, N4517);
buf BUF1 (N9598, N9591);
nor NOR4 (N9599, N9583, N2534, N1148, N7579);
nand NAND4 (N9600, N9589, N3177, N5557, N899);
or OR2 (N9601, N9598, N5239);
nand NAND2 (N9602, N9592, N7739);
xor XOR2 (N9603, N9601, N5194);
buf BUF1 (N9604, N9593);
xor XOR2 (N9605, N9599, N1547);
xor XOR2 (N9606, N9582, N1964);
buf BUF1 (N9607, N9596);
and AND2 (N9608, N9604, N1337);
not NOT1 (N9609, N9595);
and AND3 (N9610, N9600, N3552, N2988);
or OR3 (N9611, N9597, N9569, N7123);
not NOT1 (N9612, N9611);
xor XOR2 (N9613, N9603, N5171);
and AND2 (N9614, N9605, N8755);
buf BUF1 (N9615, N9612);
buf BUF1 (N9616, N9602);
xor XOR2 (N9617, N9615, N2463);
buf BUF1 (N9618, N9616);
or OR4 (N9619, N9606, N8176, N698, N2527);
xor XOR2 (N9620, N9618, N9553);
or OR4 (N9621, N9619, N3908, N7585, N4409);
buf BUF1 (N9622, N9621);
buf BUF1 (N9623, N9607);
or OR4 (N9624, N9617, N2196, N3022, N31);
xor XOR2 (N9625, N9614, N3881);
buf BUF1 (N9626, N9620);
buf BUF1 (N9627, N9625);
nor NOR2 (N9628, N9613, N5810);
xor XOR2 (N9629, N9579, N4180);
or OR2 (N9630, N9628, N3650);
nand NAND3 (N9631, N9622, N4877, N4980);
and AND2 (N9632, N9624, N1704);
buf BUF1 (N9633, N9609);
not NOT1 (N9634, N9630);
and AND3 (N9635, N9627, N3544, N8348);
xor XOR2 (N9636, N9629, N8606);
not NOT1 (N9637, N9632);
and AND2 (N9638, N9631, N1957);
xor XOR2 (N9639, N9635, N5566);
xor XOR2 (N9640, N9626, N6726);
nand NAND3 (N9641, N9638, N9565, N8659);
not NOT1 (N9642, N9640);
xor XOR2 (N9643, N9633, N1584);
nand NAND4 (N9644, N9634, N6959, N7637, N2515);
or OR2 (N9645, N9637, N1504);
or OR2 (N9646, N9639, N49);
or OR2 (N9647, N9642, N8276);
or OR2 (N9648, N9644, N5351);
not NOT1 (N9649, N9646);
nand NAND2 (N9650, N9641, N4309);
buf BUF1 (N9651, N9648);
xor XOR2 (N9652, N9645, N9523);
not NOT1 (N9653, N9636);
xor XOR2 (N9654, N9649, N2059);
nand NAND2 (N9655, N9654, N3219);
buf BUF1 (N9656, N9623);
or OR2 (N9657, N9647, N6376);
nand NAND4 (N9658, N9652, N2579, N1835, N8603);
or OR3 (N9659, N9610, N8274, N6904);
and AND2 (N9660, N9643, N1775);
xor XOR2 (N9661, N9650, N4158);
and AND3 (N9662, N9656, N6686, N850);
or OR4 (N9663, N9658, N7093, N3719, N5642);
nor NOR3 (N9664, N9660, N549, N6542);
xor XOR2 (N9665, N9662, N4064);
and AND4 (N9666, N9651, N3706, N3042, N4157);
and AND3 (N9667, N9659, N8006, N8653);
xor XOR2 (N9668, N9655, N5748);
and AND3 (N9669, N9657, N8475, N6719);
nor NOR3 (N9670, N9668, N4744, N8638);
xor XOR2 (N9671, N9666, N8281);
not NOT1 (N9672, N9671);
buf BUF1 (N9673, N9661);
nor NOR3 (N9674, N9663, N5825, N9187);
and AND4 (N9675, N9673, N5232, N3635, N1144);
not NOT1 (N9676, N9608);
buf BUF1 (N9677, N9665);
nor NOR2 (N9678, N9677, N5701);
and AND4 (N9679, N9674, N3196, N4183, N1187);
buf BUF1 (N9680, N9664);
or OR2 (N9681, N9676, N1341);
nand NAND4 (N9682, N9670, N7550, N3957, N7591);
and AND2 (N9683, N9679, N8835);
xor XOR2 (N9684, N9681, N2448);
nor NOR4 (N9685, N9672, N7647, N8262, N8345);
buf BUF1 (N9686, N9653);
xor XOR2 (N9687, N9669, N927);
nand NAND2 (N9688, N9685, N2774);
nand NAND3 (N9689, N9675, N5142, N7332);
not NOT1 (N9690, N9683);
and AND4 (N9691, N9688, N6741, N5608, N6198);
buf BUF1 (N9692, N9678);
xor XOR2 (N9693, N9692, N3521);
and AND4 (N9694, N9684, N3738, N4324, N4132);
or OR4 (N9695, N9680, N7903, N9000, N4600);
nor NOR2 (N9696, N9687, N7894);
and AND4 (N9697, N9696, N754, N2874, N2637);
nand NAND4 (N9698, N9694, N4492, N7052, N4385);
and AND4 (N9699, N9690, N1137, N4424, N1326);
nor NOR4 (N9700, N9699, N8346, N2356, N5531);
not NOT1 (N9701, N9700);
not NOT1 (N9702, N9693);
nand NAND2 (N9703, N9682, N6308);
not NOT1 (N9704, N9695);
and AND2 (N9705, N9667, N6272);
xor XOR2 (N9706, N9691, N4775);
xor XOR2 (N9707, N9686, N4655);
buf BUF1 (N9708, N9697);
nand NAND3 (N9709, N9689, N1557, N655);
xor XOR2 (N9710, N9702, N1891);
nor NOR2 (N9711, N9704, N3671);
buf BUF1 (N9712, N9703);
xor XOR2 (N9713, N9710, N2015);
nor NOR2 (N9714, N9709, N1314);
buf BUF1 (N9715, N9698);
nand NAND2 (N9716, N9707, N8774);
nand NAND4 (N9717, N9701, N1218, N6504, N1526);
buf BUF1 (N9718, N9713);
nand NAND2 (N9719, N9718, N5001);
or OR2 (N9720, N9706, N4594);
buf BUF1 (N9721, N9708);
buf BUF1 (N9722, N9714);
xor XOR2 (N9723, N9720, N5769);
nor NOR3 (N9724, N9705, N8409, N6625);
nand NAND3 (N9725, N9719, N1524, N812);
xor XOR2 (N9726, N9723, N4584);
or OR3 (N9727, N9721, N382, N6746);
buf BUF1 (N9728, N9717);
nand NAND3 (N9729, N9726, N3259, N1319);
nand NAND4 (N9730, N9724, N2341, N7720, N6133);
buf BUF1 (N9731, N9715);
nand NAND4 (N9732, N9725, N8594, N4993, N3893);
buf BUF1 (N9733, N9732);
or OR2 (N9734, N9711, N4737);
or OR4 (N9735, N9730, N9707, N1919, N8232);
xor XOR2 (N9736, N9729, N4083);
not NOT1 (N9737, N9722);
nand NAND3 (N9738, N9737, N1981, N3098);
xor XOR2 (N9739, N9736, N8977);
nand NAND3 (N9740, N9735, N1365, N5289);
nor NOR3 (N9741, N9740, N5095, N3864);
and AND4 (N9742, N9728, N2799, N1728, N2992);
nand NAND3 (N9743, N9716, N9612, N3435);
not NOT1 (N9744, N9742);
not NOT1 (N9745, N9727);
buf BUF1 (N9746, N9733);
buf BUF1 (N9747, N9745);
buf BUF1 (N9748, N9747);
nand NAND2 (N9749, N9743, N1173);
nand NAND3 (N9750, N9744, N2909, N5753);
xor XOR2 (N9751, N9750, N940);
xor XOR2 (N9752, N9739, N9008);
nor NOR4 (N9753, N9741, N7491, N307, N5435);
and AND3 (N9754, N9731, N5737, N6756);
and AND2 (N9755, N9746, N4278);
nor NOR2 (N9756, N9749, N5804);
buf BUF1 (N9757, N9755);
nand NAND4 (N9758, N9751, N7961, N527, N3690);
xor XOR2 (N9759, N9748, N2898);
or OR3 (N9760, N9738, N8174, N1850);
buf BUF1 (N9761, N9758);
and AND2 (N9762, N9752, N8166);
or OR3 (N9763, N9757, N8587, N8615);
not NOT1 (N9764, N9763);
buf BUF1 (N9765, N9760);
and AND3 (N9766, N9712, N5553, N1786);
not NOT1 (N9767, N9756);
nand NAND3 (N9768, N9762, N6303, N6457);
nand NAND4 (N9769, N9767, N7590, N7474, N211);
buf BUF1 (N9770, N9768);
nor NOR3 (N9771, N9766, N680, N1280);
nor NOR3 (N9772, N9759, N1552, N4626);
buf BUF1 (N9773, N9772);
nand NAND4 (N9774, N9770, N532, N5133, N5046);
not NOT1 (N9775, N9761);
buf BUF1 (N9776, N9775);
xor XOR2 (N9777, N9773, N2846);
and AND3 (N9778, N9764, N5400, N5272);
or OR4 (N9779, N9753, N2292, N6025, N7151);
buf BUF1 (N9780, N9778);
buf BUF1 (N9781, N9780);
buf BUF1 (N9782, N9781);
buf BUF1 (N9783, N9734);
buf BUF1 (N9784, N9779);
nand NAND2 (N9785, N9765, N6920);
and AND4 (N9786, N9784, N5115, N4884, N8629);
nor NOR3 (N9787, N9754, N2916, N2276);
nand NAND2 (N9788, N9771, N4198);
or OR2 (N9789, N9783, N9788);
nand NAND4 (N9790, N7625, N4392, N1733, N5325);
or OR3 (N9791, N9790, N2491, N1081);
xor XOR2 (N9792, N9774, N6801);
not NOT1 (N9793, N9769);
not NOT1 (N9794, N9777);
nor NOR4 (N9795, N9776, N4099, N6915, N7709);
not NOT1 (N9796, N9792);
nand NAND2 (N9797, N9795, N9124);
nand NAND3 (N9798, N9785, N3777, N649);
not NOT1 (N9799, N9797);
not NOT1 (N9800, N9789);
nand NAND3 (N9801, N9796, N5467, N4521);
or OR4 (N9802, N9791, N8600, N7693, N2500);
xor XOR2 (N9803, N9802, N6603);
nor NOR3 (N9804, N9787, N238, N607);
or OR3 (N9805, N9786, N6125, N7240);
and AND2 (N9806, N9799, N4269);
or OR2 (N9807, N9801, N7738);
nor NOR3 (N9808, N9793, N3637, N7534);
nor NOR2 (N9809, N9806, N7378);
or OR2 (N9810, N9809, N9380);
or OR3 (N9811, N9804, N945, N9805);
nand NAND4 (N9812, N5911, N4338, N3492, N8456);
nor NOR2 (N9813, N9807, N393);
not NOT1 (N9814, N9810);
buf BUF1 (N9815, N9808);
xor XOR2 (N9816, N9813, N7851);
or OR3 (N9817, N9814, N3127, N7546);
xor XOR2 (N9818, N9803, N5078);
or OR4 (N9819, N9794, N1238, N5332, N7608);
and AND3 (N9820, N9782, N932, N1022);
nor NOR2 (N9821, N9800, N3728);
or OR4 (N9822, N9820, N9125, N7464, N7700);
nor NOR2 (N9823, N9818, N2366);
and AND4 (N9824, N9815, N5119, N1528, N4819);
not NOT1 (N9825, N9823);
nor NOR3 (N9826, N9812, N3185, N5008);
nor NOR3 (N9827, N9819, N3622, N4231);
and AND4 (N9828, N9827, N7866, N7642, N4101);
not NOT1 (N9829, N9811);
buf BUF1 (N9830, N9826);
nor NOR4 (N9831, N9829, N3554, N8222, N2629);
or OR3 (N9832, N9817, N72, N5700);
nand NAND4 (N9833, N9798, N6886, N5566, N1229);
nor NOR2 (N9834, N9828, N4260);
nor NOR3 (N9835, N9821, N1517, N4165);
nand NAND3 (N9836, N9833, N3343, N8786);
or OR3 (N9837, N9816, N492, N4062);
xor XOR2 (N9838, N9834, N6179);
or OR3 (N9839, N9831, N9524, N9469);
xor XOR2 (N9840, N9822, N1245);
nor NOR3 (N9841, N9825, N3433, N9409);
xor XOR2 (N9842, N9838, N6406);
not NOT1 (N9843, N9839);
buf BUF1 (N9844, N9824);
not NOT1 (N9845, N9832);
buf BUF1 (N9846, N9844);
or OR2 (N9847, N9845, N1737);
nand NAND4 (N9848, N9835, N4294, N6317, N7266);
not NOT1 (N9849, N9847);
nand NAND4 (N9850, N9842, N4621, N3306, N4430);
not NOT1 (N9851, N9841);
and AND4 (N9852, N9837, N4049, N1097, N4790);
and AND3 (N9853, N9851, N9220, N8892);
not NOT1 (N9854, N9843);
or OR2 (N9855, N9853, N4792);
xor XOR2 (N9856, N9840, N8669);
nor NOR3 (N9857, N9849, N5805, N4306);
not NOT1 (N9858, N9854);
nor NOR3 (N9859, N9836, N2096, N4890);
nand NAND4 (N9860, N9850, N4157, N5445, N973);
nand NAND4 (N9861, N9856, N1858, N6881, N5462);
buf BUF1 (N9862, N9859);
or OR3 (N9863, N9861, N4882, N1318);
buf BUF1 (N9864, N9858);
nor NOR2 (N9865, N9846, N5261);
not NOT1 (N9866, N9863);
nand NAND4 (N9867, N9866, N8875, N9253, N4839);
nor NOR4 (N9868, N9865, N3675, N2442, N8409);
nor NOR4 (N9869, N9848, N5470, N6960, N4385);
nand NAND4 (N9870, N9852, N6149, N5528, N4561);
or OR2 (N9871, N9864, N2041);
nor NOR4 (N9872, N9869, N6858, N3586, N4001);
not NOT1 (N9873, N9871);
nand NAND2 (N9874, N9830, N7192);
xor XOR2 (N9875, N9874, N9418);
nor NOR4 (N9876, N9872, N6414, N6535, N5281);
or OR3 (N9877, N9868, N614, N3076);
nand NAND2 (N9878, N9875, N813);
xor XOR2 (N9879, N9862, N577);
and AND4 (N9880, N9857, N8263, N45, N6567);
nor NOR2 (N9881, N9876, N8614);
nor NOR4 (N9882, N9855, N9838, N8429, N8572);
and AND3 (N9883, N9860, N8621, N372);
buf BUF1 (N9884, N9879);
not NOT1 (N9885, N9881);
and AND4 (N9886, N9882, N2757, N6415, N8936);
and AND4 (N9887, N9885, N3075, N764, N3424);
and AND2 (N9888, N9873, N1654);
nor NOR3 (N9889, N9880, N6888, N7874);
and AND4 (N9890, N9887, N4207, N9594, N6120);
nor NOR3 (N9891, N9889, N3661, N7690);
buf BUF1 (N9892, N9878);
xor XOR2 (N9893, N9888, N9408);
xor XOR2 (N9894, N9867, N1366);
buf BUF1 (N9895, N9891);
nand NAND4 (N9896, N9890, N5920, N2319, N1929);
nor NOR2 (N9897, N9886, N8131);
and AND4 (N9898, N9870, N5857, N9892, N3888);
buf BUF1 (N9899, N5455);
not NOT1 (N9900, N9895);
and AND3 (N9901, N9896, N3277, N561);
nor NOR3 (N9902, N9884, N9031, N9359);
and AND2 (N9903, N9900, N4922);
buf BUF1 (N9904, N9877);
buf BUF1 (N9905, N9902);
xor XOR2 (N9906, N9904, N4689);
or OR4 (N9907, N9903, N3745, N3778, N9381);
or OR3 (N9908, N9894, N911, N930);
buf BUF1 (N9909, N9893);
nand NAND4 (N9910, N9898, N1364, N3230, N5873);
or OR2 (N9911, N9899, N6983);
xor XOR2 (N9912, N9910, N160);
not NOT1 (N9913, N9911);
and AND3 (N9914, N9905, N4465, N24);
and AND3 (N9915, N9897, N6684, N5251);
xor XOR2 (N9916, N9906, N7903);
or OR4 (N9917, N9901, N5850, N4525, N916);
nand NAND2 (N9918, N9883, N7465);
not NOT1 (N9919, N9907);
or OR3 (N9920, N9917, N2221, N7711);
or OR3 (N9921, N9919, N7141, N7394);
or OR2 (N9922, N9916, N3779);
nand NAND2 (N9923, N9912, N5147);
nand NAND3 (N9924, N9921, N4847, N8556);
not NOT1 (N9925, N9909);
nor NOR4 (N9926, N9918, N6844, N5097, N5385);
or OR2 (N9927, N9913, N6396);
or OR4 (N9928, N9914, N4652, N5263, N3762);
nor NOR2 (N9929, N9928, N3416);
and AND2 (N9930, N9922, N8667);
xor XOR2 (N9931, N9925, N3764);
or OR3 (N9932, N9929, N521, N6252);
nor NOR4 (N9933, N9926, N6493, N7207, N8764);
not NOT1 (N9934, N9920);
buf BUF1 (N9935, N9932);
nor NOR4 (N9936, N9935, N3770, N1664, N9556);
or OR4 (N9937, N9908, N8220, N715, N3739);
and AND4 (N9938, N9933, N7219, N6459, N5301);
and AND3 (N9939, N9915, N9469, N8414);
not NOT1 (N9940, N9936);
and AND2 (N9941, N9934, N8333);
buf BUF1 (N9942, N9923);
nor NOR3 (N9943, N9938, N3909, N460);
buf BUF1 (N9944, N9937);
nand NAND4 (N9945, N9924, N1698, N2344, N3028);
xor XOR2 (N9946, N9927, N4440);
or OR2 (N9947, N9939, N3084);
nor NOR2 (N9948, N9945, N4375);
and AND3 (N9949, N9941, N5057, N8383);
buf BUF1 (N9950, N9940);
nor NOR2 (N9951, N9930, N9155);
xor XOR2 (N9952, N9947, N6814);
or OR2 (N9953, N9943, N371);
not NOT1 (N9954, N9949);
nand NAND3 (N9955, N9942, N4178, N2639);
not NOT1 (N9956, N9931);
xor XOR2 (N9957, N9944, N6803);
or OR2 (N9958, N9953, N1365);
or OR3 (N9959, N9958, N5400, N1649);
or OR3 (N9960, N9946, N7467, N465);
nand NAND3 (N9961, N9952, N5776, N5342);
nand NAND2 (N9962, N9955, N6859);
and AND2 (N9963, N9961, N5256);
not NOT1 (N9964, N9954);
nor NOR3 (N9965, N9964, N2511, N3742);
and AND4 (N9966, N9965, N6790, N1579, N1158);
nor NOR2 (N9967, N9966, N1935);
xor XOR2 (N9968, N9956, N1619);
and AND3 (N9969, N9959, N8160, N3765);
buf BUF1 (N9970, N9967);
or OR2 (N9971, N9960, N3573);
nand NAND3 (N9972, N9957, N885, N134);
xor XOR2 (N9973, N9962, N7335);
xor XOR2 (N9974, N9950, N4134);
nand NAND3 (N9975, N9970, N8136, N5917);
xor XOR2 (N9976, N9971, N2871);
nand NAND4 (N9977, N9976, N3822, N1482, N5894);
and AND3 (N9978, N9974, N6359, N6956);
and AND3 (N9979, N9973, N9821, N9263);
xor XOR2 (N9980, N9977, N3046);
xor XOR2 (N9981, N9963, N6693);
and AND3 (N9982, N9969, N7554, N205);
nand NAND2 (N9983, N9948, N3661);
nor NOR2 (N9984, N9951, N1438);
nor NOR4 (N9985, N9981, N4695, N7900, N3792);
buf BUF1 (N9986, N9968);
nand NAND4 (N9987, N9978, N8939, N564, N69);
buf BUF1 (N9988, N9983);
nor NOR4 (N9989, N9982, N5540, N8654, N7454);
buf BUF1 (N9990, N9985);
nand NAND3 (N9991, N9972, N6065, N8207);
or OR4 (N9992, N9989, N7942, N1390, N6732);
or OR3 (N9993, N9987, N6288, N274);
not NOT1 (N9994, N9990);
nand NAND4 (N9995, N9975, N9389, N460, N2591);
xor XOR2 (N9996, N9979, N4973);
nor NOR3 (N9997, N9992, N5027, N1406);
or OR3 (N9998, N9988, N1212, N1251);
and AND4 (N9999, N9991, N7727, N9868, N8516);
nor NOR4 (N10000, N9997, N1297, N762, N7855);
buf BUF1 (N10001, N9998);
buf BUF1 (N10002, N9984);
not NOT1 (N10003, N10002);
nor NOR4 (N10004, N9999, N4459, N2800, N5468);
xor XOR2 (N10005, N9996, N4137);
or OR4 (N10006, N9993, N5536, N7586, N4106);
xor XOR2 (N10007, N10001, N5099);
buf BUF1 (N10008, N10003);
nor NOR4 (N10009, N10007, N2949, N8328, N9904);
buf BUF1 (N10010, N10005);
and AND4 (N10011, N9986, N8607, N7852, N7956);
nor NOR4 (N10012, N9995, N8168, N8445, N4577);
and AND2 (N10013, N10009, N5582);
and AND4 (N10014, N10004, N3193, N3483, N8084);
xor XOR2 (N10015, N10014, N4734);
buf BUF1 (N10016, N10010);
or OR3 (N10017, N10008, N4651, N4459);
not NOT1 (N10018, N10012);
xor XOR2 (N10019, N10018, N1111);
not NOT1 (N10020, N10000);
not NOT1 (N10021, N9980);
buf BUF1 (N10022, N9994);
not NOT1 (N10023, N10013);
nor NOR3 (N10024, N10017, N6609, N6425);
xor XOR2 (N10025, N10015, N7523);
or OR3 (N10026, N10020, N3596, N8601);
not NOT1 (N10027, N10021);
not NOT1 (N10028, N10025);
nand NAND2 (N10029, N10026, N5751);
nand NAND2 (N10030, N10027, N5622);
or OR2 (N10031, N10029, N1861);
xor XOR2 (N10032, N10023, N1658);
not NOT1 (N10033, N10022);
xor XOR2 (N10034, N10030, N4417);
nand NAND4 (N10035, N10016, N6219, N965, N9511);
nor NOR4 (N10036, N10035, N7540, N3690, N271);
nand NAND4 (N10037, N10034, N4615, N7548, N699);
and AND4 (N10038, N10024, N9036, N646, N1965);
and AND2 (N10039, N10032, N4975);
not NOT1 (N10040, N10033);
and AND2 (N10041, N10031, N7281);
or OR2 (N10042, N10019, N8291);
buf BUF1 (N10043, N10038);
nand NAND4 (N10044, N10040, N4296, N6647, N4773);
not NOT1 (N10045, N10044);
nor NOR3 (N10046, N10037, N7761, N7071);
buf BUF1 (N10047, N10046);
nand NAND3 (N10048, N10011, N6394, N7178);
nand NAND4 (N10049, N10045, N82, N409, N8856);
xor XOR2 (N10050, N10042, N7314);
nor NOR4 (N10051, N10049, N917, N908, N4133);
not NOT1 (N10052, N10043);
xor XOR2 (N10053, N10036, N5543);
not NOT1 (N10054, N10006);
not NOT1 (N10055, N10053);
or OR2 (N10056, N10039, N8570);
not NOT1 (N10057, N10052);
or OR3 (N10058, N10055, N2653, N4613);
not NOT1 (N10059, N10054);
xor XOR2 (N10060, N10028, N7638);
nor NOR3 (N10061, N10058, N4541, N6947);
xor XOR2 (N10062, N10041, N5340);
or OR3 (N10063, N10047, N1334, N622);
or OR3 (N10064, N10056, N4021, N6323);
nor NOR4 (N10065, N10048, N3989, N2753, N117);
xor XOR2 (N10066, N10060, N2914);
not NOT1 (N10067, N10057);
and AND4 (N10068, N10061, N8533, N5292, N4356);
and AND4 (N10069, N10067, N3628, N1414, N2198);
nand NAND2 (N10070, N10064, N5868);
or OR4 (N10071, N10065, N6676, N7069, N5565);
buf BUF1 (N10072, N10063);
or OR4 (N10073, N10069, N4877, N3587, N3766);
or OR3 (N10074, N10068, N6339, N6963);
buf BUF1 (N10075, N10070);
buf BUF1 (N10076, N10066);
buf BUF1 (N10077, N10075);
nand NAND3 (N10078, N10050, N462, N3365);
not NOT1 (N10079, N10059);
nand NAND2 (N10080, N10071, N2886);
buf BUF1 (N10081, N10076);
and AND4 (N10082, N10051, N2719, N754, N8286);
not NOT1 (N10083, N10074);
or OR2 (N10084, N10077, N4012);
and AND2 (N10085, N10079, N7365);
or OR3 (N10086, N10083, N6661, N9590);
or OR3 (N10087, N10081, N7429, N2680);
or OR4 (N10088, N10085, N3216, N5766, N10058);
nor NOR2 (N10089, N10072, N6994);
or OR4 (N10090, N10086, N3017, N2704, N8457);
or OR2 (N10091, N10080, N5943);
buf BUF1 (N10092, N10090);
not NOT1 (N10093, N10091);
not NOT1 (N10094, N10093);
nand NAND3 (N10095, N10084, N796, N9864);
xor XOR2 (N10096, N10095, N2728);
not NOT1 (N10097, N10073);
not NOT1 (N10098, N10088);
buf BUF1 (N10099, N10097);
and AND4 (N10100, N10062, N6478, N9730, N2073);
or OR3 (N10101, N10082, N6167, N8845);
nand NAND3 (N10102, N10100, N8199, N9484);
or OR4 (N10103, N10094, N3733, N6271, N9660);
and AND2 (N10104, N10078, N4155);
and AND2 (N10105, N10092, N4237);
and AND2 (N10106, N10087, N314);
xor XOR2 (N10107, N10102, N8653);
buf BUF1 (N10108, N10107);
or OR4 (N10109, N10089, N9532, N8775, N4957);
xor XOR2 (N10110, N10109, N9202);
nor NOR4 (N10111, N10096, N8855, N5718, N7590);
and AND3 (N10112, N10101, N1350, N4876);
not NOT1 (N10113, N10108);
not NOT1 (N10114, N10111);
buf BUF1 (N10115, N10103);
not NOT1 (N10116, N10113);
xor XOR2 (N10117, N10106, N4692);
buf BUF1 (N10118, N10099);
buf BUF1 (N10119, N10104);
xor XOR2 (N10120, N10115, N2987);
not NOT1 (N10121, N10112);
buf BUF1 (N10122, N10118);
or OR2 (N10123, N10122, N7489);
not NOT1 (N10124, N10123);
nor NOR2 (N10125, N10105, N2686);
xor XOR2 (N10126, N10120, N1891);
not NOT1 (N10127, N10110);
nor NOR3 (N10128, N10116, N4217, N1394);
buf BUF1 (N10129, N10128);
xor XOR2 (N10130, N10129, N1128);
and AND3 (N10131, N10130, N6680, N4505);
nor NOR3 (N10132, N10127, N4871, N9887);
nand NAND3 (N10133, N10132, N5310, N3100);
nor NOR3 (N10134, N10114, N132, N4081);
nor NOR2 (N10135, N10117, N2429);
buf BUF1 (N10136, N10126);
nand NAND2 (N10137, N10124, N3570);
and AND2 (N10138, N10137, N513);
not NOT1 (N10139, N10119);
nand NAND2 (N10140, N10135, N9451);
xor XOR2 (N10141, N10125, N7359);
or OR2 (N10142, N10140, N4598);
not NOT1 (N10143, N10136);
buf BUF1 (N10144, N10121);
and AND2 (N10145, N10139, N8666);
not NOT1 (N10146, N10142);
not NOT1 (N10147, N10146);
nand NAND3 (N10148, N10145, N496, N8777);
and AND3 (N10149, N10131, N4469, N9633);
nand NAND2 (N10150, N10144, N9364);
buf BUF1 (N10151, N10143);
and AND3 (N10152, N10151, N1834, N9781);
and AND2 (N10153, N10138, N3321);
buf BUF1 (N10154, N10152);
xor XOR2 (N10155, N10147, N8709);
not NOT1 (N10156, N10141);
xor XOR2 (N10157, N10148, N4385);
and AND3 (N10158, N10098, N6387, N1925);
nor NOR3 (N10159, N10150, N3115, N8047);
and AND2 (N10160, N10133, N8294);
buf BUF1 (N10161, N10160);
not NOT1 (N10162, N10149);
nand NAND4 (N10163, N10153, N7664, N2104, N868);
buf BUF1 (N10164, N10158);
buf BUF1 (N10165, N10154);
buf BUF1 (N10166, N10165);
and AND3 (N10167, N10155, N803, N10067);
and AND2 (N10168, N10161, N5188);
or OR4 (N10169, N10162, N1658, N1659, N3013);
buf BUF1 (N10170, N10166);
and AND3 (N10171, N10164, N3251, N9388);
nor NOR2 (N10172, N10167, N2683);
buf BUF1 (N10173, N10157);
not NOT1 (N10174, N10173);
nor NOR3 (N10175, N10168, N8774, N3139);
not NOT1 (N10176, N10171);
nand NAND4 (N10177, N10174, N7911, N7014, N7403);
buf BUF1 (N10178, N10169);
xor XOR2 (N10179, N10177, N2601);
nor NOR4 (N10180, N10178, N4267, N3052, N8604);
nand NAND4 (N10181, N10159, N1823, N2000, N4177);
and AND3 (N10182, N10175, N2553, N435);
xor XOR2 (N10183, N10182, N2843);
xor XOR2 (N10184, N10181, N1376);
not NOT1 (N10185, N10180);
nand NAND2 (N10186, N10134, N3485);
not NOT1 (N10187, N10185);
or OR2 (N10188, N10170, N4303);
xor XOR2 (N10189, N10183, N1164);
xor XOR2 (N10190, N10163, N7742);
nor NOR3 (N10191, N10189, N4416, N3107);
xor XOR2 (N10192, N10186, N9206);
buf BUF1 (N10193, N10184);
nand NAND2 (N10194, N10188, N9414);
not NOT1 (N10195, N10179);
not NOT1 (N10196, N10187);
or OR4 (N10197, N10172, N8336, N1547, N7543);
nor NOR4 (N10198, N10195, N4545, N9878, N6207);
not NOT1 (N10199, N10196);
or OR4 (N10200, N10190, N6309, N58, N226);
nor NOR3 (N10201, N10199, N7915, N2374);
nand NAND4 (N10202, N10156, N417, N7995, N6601);
not NOT1 (N10203, N10197);
nand NAND3 (N10204, N10192, N7757, N4606);
or OR2 (N10205, N10191, N4448);
nor NOR4 (N10206, N10176, N3104, N8749, N4453);
or OR2 (N10207, N10203, N6288);
not NOT1 (N10208, N10202);
xor XOR2 (N10209, N10194, N3776);
buf BUF1 (N10210, N10204);
nand NAND2 (N10211, N10206, N2515);
or OR4 (N10212, N10201, N9976, N2431, N227);
or OR4 (N10213, N10193, N1768, N3908, N7638);
nand NAND3 (N10214, N10198, N3631, N302);
buf BUF1 (N10215, N10211);
not NOT1 (N10216, N10212);
and AND2 (N10217, N10216, N9860);
or OR2 (N10218, N10217, N7409);
nor NOR2 (N10219, N10205, N10155);
buf BUF1 (N10220, N10219);
and AND2 (N10221, N10215, N1851);
nor NOR2 (N10222, N10213, N7544);
nor NOR3 (N10223, N10222, N5692, N5006);
and AND4 (N10224, N10214, N3307, N1784, N4925);
and AND2 (N10225, N10221, N3933);
nor NOR2 (N10226, N10218, N1490);
xor XOR2 (N10227, N10224, N9999);
nand NAND3 (N10228, N10225, N5836, N5647);
nand NAND4 (N10229, N10209, N813, N8900, N6181);
not NOT1 (N10230, N10228);
xor XOR2 (N10231, N10227, N1891);
xor XOR2 (N10232, N10223, N733);
not NOT1 (N10233, N10207);
nand NAND2 (N10234, N10220, N6911);
xor XOR2 (N10235, N10200, N302);
nand NAND3 (N10236, N10229, N8983, N2570);
nand NAND3 (N10237, N10235, N4551, N7007);
nand NAND4 (N10238, N10208, N4864, N9829, N2349);
xor XOR2 (N10239, N10210, N1743);
xor XOR2 (N10240, N10234, N8360);
and AND4 (N10241, N10233, N8110, N10057, N3530);
and AND3 (N10242, N10237, N9561, N10032);
or OR2 (N10243, N10230, N8426);
or OR4 (N10244, N10243, N9552, N171, N10186);
or OR2 (N10245, N10236, N6360);
nor NOR2 (N10246, N10241, N5475);
or OR3 (N10247, N10240, N5954, N161);
nand NAND2 (N10248, N10231, N6487);
buf BUF1 (N10249, N10246);
xor XOR2 (N10250, N10244, N6584);
xor XOR2 (N10251, N10242, N4639);
not NOT1 (N10252, N10249);
not NOT1 (N10253, N10247);
xor XOR2 (N10254, N10239, N5701);
nor NOR3 (N10255, N10226, N7461, N7762);
and AND4 (N10256, N10245, N6484, N8462, N3849);
buf BUF1 (N10257, N10238);
nand NAND2 (N10258, N10255, N1017);
xor XOR2 (N10259, N10251, N206);
nand NAND2 (N10260, N10258, N796);
xor XOR2 (N10261, N10232, N3632);
nand NAND3 (N10262, N10254, N9884, N3850);
not NOT1 (N10263, N10256);
or OR3 (N10264, N10261, N8030, N9499);
nor NOR4 (N10265, N10252, N6179, N2370, N9593);
not NOT1 (N10266, N10263);
or OR4 (N10267, N10259, N5397, N9639, N1231);
nor NOR3 (N10268, N10264, N3525, N10164);
and AND3 (N10269, N10267, N4778, N6060);
not NOT1 (N10270, N10260);
not NOT1 (N10271, N10268);
not NOT1 (N10272, N10257);
nor NOR3 (N10273, N10248, N3693, N1107);
nor NOR4 (N10274, N10270, N8121, N3020, N636);
buf BUF1 (N10275, N10253);
not NOT1 (N10276, N10273);
nand NAND4 (N10277, N10274, N920, N8235, N5974);
nand NAND4 (N10278, N10277, N2905, N8300, N7185);
buf BUF1 (N10279, N10262);
nand NAND3 (N10280, N10272, N4077, N4755);
not NOT1 (N10281, N10280);
not NOT1 (N10282, N10281);
nand NAND4 (N10283, N10269, N1157, N7536, N987);
not NOT1 (N10284, N10283);
buf BUF1 (N10285, N10271);
or OR2 (N10286, N10276, N6828);
buf BUF1 (N10287, N10285);
not NOT1 (N10288, N10275);
buf BUF1 (N10289, N10284);
buf BUF1 (N10290, N10278);
nor NOR4 (N10291, N10279, N9658, N2112, N5357);
nand NAND3 (N10292, N10282, N159, N4453);
nand NAND3 (N10293, N10250, N3377, N3552);
and AND2 (N10294, N10291, N3729);
not NOT1 (N10295, N10290);
xor XOR2 (N10296, N10289, N9100);
and AND2 (N10297, N10292, N590);
or OR4 (N10298, N10286, N9929, N9063, N6931);
xor XOR2 (N10299, N10287, N3219);
buf BUF1 (N10300, N10294);
not NOT1 (N10301, N10297);
nand NAND2 (N10302, N10288, N3284);
xor XOR2 (N10303, N10295, N9689);
buf BUF1 (N10304, N10302);
xor XOR2 (N10305, N10293, N1447);
or OR3 (N10306, N10305, N6494, N8022);
nor NOR2 (N10307, N10296, N3308);
and AND4 (N10308, N10303, N6940, N2339, N3219);
or OR3 (N10309, N10299, N3888, N462);
nand NAND4 (N10310, N10309, N586, N6922, N8425);
nand NAND2 (N10311, N10304, N1589);
not NOT1 (N10312, N10300);
nor NOR4 (N10313, N10308, N8458, N5724, N9362);
not NOT1 (N10314, N10311);
buf BUF1 (N10315, N10312);
or OR2 (N10316, N10315, N1826);
xor XOR2 (N10317, N10266, N7008);
or OR3 (N10318, N10265, N6079, N5641);
nand NAND3 (N10319, N10301, N7199, N5500);
not NOT1 (N10320, N10314);
xor XOR2 (N10321, N10298, N4149);
or OR3 (N10322, N10319, N9036, N6900);
nand NAND4 (N10323, N10317, N9403, N5173, N5426);
and AND3 (N10324, N10306, N1820, N3761);
and AND2 (N10325, N10307, N4781);
nor NOR3 (N10326, N10316, N9341, N290);
or OR2 (N10327, N10325, N2008);
or OR3 (N10328, N10326, N9652, N1379);
nor NOR3 (N10329, N10324, N7146, N7094);
not NOT1 (N10330, N10329);
not NOT1 (N10331, N10322);
nand NAND3 (N10332, N10330, N3989, N4163);
buf BUF1 (N10333, N10313);
xor XOR2 (N10334, N10321, N8160);
or OR2 (N10335, N10310, N2100);
buf BUF1 (N10336, N10335);
nand NAND3 (N10337, N10320, N7195, N5205);
and AND2 (N10338, N10331, N2014);
xor XOR2 (N10339, N10338, N3200);
and AND2 (N10340, N10318, N6736);
nand NAND3 (N10341, N10340, N9358, N6012);
nand NAND2 (N10342, N10328, N6012);
not NOT1 (N10343, N10341);
nor NOR4 (N10344, N10336, N1779, N6918, N2852);
buf BUF1 (N10345, N10332);
or OR2 (N10346, N10323, N7252);
nor NOR2 (N10347, N10327, N8401);
nand NAND2 (N10348, N10344, N967);
xor XOR2 (N10349, N10345, N8387);
not NOT1 (N10350, N10347);
xor XOR2 (N10351, N10339, N570);
nand NAND4 (N10352, N10337, N977, N3589, N4956);
and AND2 (N10353, N10333, N113);
buf BUF1 (N10354, N10352);
or OR3 (N10355, N10350, N606, N5498);
or OR3 (N10356, N10342, N7231, N6108);
buf BUF1 (N10357, N10343);
buf BUF1 (N10358, N10351);
and AND4 (N10359, N10348, N4076, N4528, N36);
xor XOR2 (N10360, N10357, N2696);
xor XOR2 (N10361, N10355, N3605);
or OR4 (N10362, N10360, N2536, N3790, N6405);
buf BUF1 (N10363, N10346);
or OR2 (N10364, N10334, N5609);
and AND4 (N10365, N10361, N4022, N3948, N824);
nand NAND2 (N10366, N10353, N1180);
nand NAND4 (N10367, N10365, N7741, N1825, N3457);
or OR4 (N10368, N10349, N7881, N5112, N2361);
or OR4 (N10369, N10363, N7184, N612, N5857);
xor XOR2 (N10370, N10358, N7799);
nor NOR4 (N10371, N10359, N5241, N2065, N5794);
buf BUF1 (N10372, N10354);
not NOT1 (N10373, N10356);
xor XOR2 (N10374, N10367, N678);
xor XOR2 (N10375, N10372, N8998);
xor XOR2 (N10376, N10364, N2055);
nand NAND2 (N10377, N10371, N7985);
and AND3 (N10378, N10376, N6612, N5661);
nand NAND3 (N10379, N10368, N9350, N1182);
nor NOR2 (N10380, N10377, N2336);
buf BUF1 (N10381, N10375);
or OR3 (N10382, N10381, N6299, N3336);
and AND4 (N10383, N10374, N5671, N3507, N4923);
nand NAND2 (N10384, N10362, N4079);
xor XOR2 (N10385, N10383, N1730);
not NOT1 (N10386, N10378);
or OR2 (N10387, N10370, N3689);
nand NAND4 (N10388, N10366, N3779, N1941, N8054);
xor XOR2 (N10389, N10373, N5618);
nand NAND3 (N10390, N10369, N4560, N10328);
not NOT1 (N10391, N10380);
and AND3 (N10392, N10387, N5890, N9542);
or OR3 (N10393, N10392, N82, N3258);
nand NAND2 (N10394, N10389, N10258);
buf BUF1 (N10395, N10385);
xor XOR2 (N10396, N10388, N6385);
and AND2 (N10397, N10394, N3859);
not NOT1 (N10398, N10379);
nand NAND4 (N10399, N10390, N1420, N2800, N9824);
not NOT1 (N10400, N10382);
buf BUF1 (N10401, N10399);
and AND3 (N10402, N10391, N2401, N8142);
and AND3 (N10403, N10400, N2490, N2899);
xor XOR2 (N10404, N10398, N3272);
buf BUF1 (N10405, N10393);
or OR4 (N10406, N10384, N425, N5938, N7232);
not NOT1 (N10407, N10401);
and AND4 (N10408, N10407, N8635, N1906, N3665);
buf BUF1 (N10409, N10408);
nor NOR3 (N10410, N10386, N6178, N9172);
buf BUF1 (N10411, N10405);
nor NOR4 (N10412, N10397, N993, N591, N8371);
and AND2 (N10413, N10403, N8257);
buf BUF1 (N10414, N10412);
or OR3 (N10415, N10413, N10080, N1166);
xor XOR2 (N10416, N10410, N8275);
and AND3 (N10417, N10409, N5890, N1774);
xor XOR2 (N10418, N10406, N9661);
nor NOR3 (N10419, N10414, N7176, N9791);
or OR2 (N10420, N10404, N2762);
and AND4 (N10421, N10415, N3590, N2379, N2881);
xor XOR2 (N10422, N10418, N6701);
nor NOR2 (N10423, N10396, N5596);
nor NOR4 (N10424, N10402, N1069, N9935, N7539);
nor NOR2 (N10425, N10423, N134);
buf BUF1 (N10426, N10421);
xor XOR2 (N10427, N10422, N8630);
buf BUF1 (N10428, N10411);
not NOT1 (N10429, N10417);
xor XOR2 (N10430, N10395, N6896);
and AND4 (N10431, N10419, N2979, N4103, N1593);
and AND3 (N10432, N10430, N5034, N6244);
buf BUF1 (N10433, N10416);
buf BUF1 (N10434, N10425);
nor NOR4 (N10435, N10433, N1281, N8767, N2724);
nor NOR4 (N10436, N10420, N4866, N2133, N1353);
buf BUF1 (N10437, N10426);
not NOT1 (N10438, N10435);
not NOT1 (N10439, N10429);
or OR3 (N10440, N10436, N8563, N4060);
and AND4 (N10441, N10427, N5427, N230, N8844);
xor XOR2 (N10442, N10439, N5303);
nor NOR3 (N10443, N10432, N10242, N9118);
buf BUF1 (N10444, N10442);
and AND2 (N10445, N10438, N5464);
not NOT1 (N10446, N10441);
nand NAND3 (N10447, N10437, N6598, N3392);
nor NOR3 (N10448, N10444, N940, N87);
nand NAND4 (N10449, N10443, N4840, N59, N1527);
nor NOR2 (N10450, N10431, N8085);
xor XOR2 (N10451, N10446, N7850);
xor XOR2 (N10452, N10445, N880);
nand NAND4 (N10453, N10450, N5392, N302, N4894);
nand NAND3 (N10454, N10428, N3239, N8769);
and AND3 (N10455, N10449, N2132, N6661);
or OR3 (N10456, N10448, N6429, N7626);
or OR2 (N10457, N10424, N1926);
buf BUF1 (N10458, N10447);
buf BUF1 (N10459, N10452);
nand NAND2 (N10460, N10455, N2198);
xor XOR2 (N10461, N10458, N8823);
or OR3 (N10462, N10461, N7786, N6432);
not NOT1 (N10463, N10454);
buf BUF1 (N10464, N10460);
and AND4 (N10465, N10456, N8271, N4283, N4950);
not NOT1 (N10466, N10465);
nor NOR3 (N10467, N10434, N4085, N2207);
buf BUF1 (N10468, N10463);
nor NOR4 (N10469, N10453, N1488, N1590, N7834);
buf BUF1 (N10470, N10469);
or OR2 (N10471, N10462, N9522);
xor XOR2 (N10472, N10451, N6740);
nand NAND4 (N10473, N10457, N2610, N8115, N9663);
nand NAND3 (N10474, N10471, N5, N5174);
not NOT1 (N10475, N10464);
buf BUF1 (N10476, N10459);
nand NAND4 (N10477, N10476, N2967, N8235, N3189);
nor NOR3 (N10478, N10477, N6019, N7793);
xor XOR2 (N10479, N10470, N4788);
and AND3 (N10480, N10478, N5512, N6497);
nand NAND4 (N10481, N10472, N7299, N4836, N1595);
nand NAND4 (N10482, N10475, N10385, N10163, N9916);
nand NAND2 (N10483, N10466, N1861);
not NOT1 (N10484, N10474);
and AND4 (N10485, N10468, N813, N3473, N1334);
and AND3 (N10486, N10484, N7196, N5946);
not NOT1 (N10487, N10480);
nor NOR3 (N10488, N10479, N7284, N10153);
not NOT1 (N10489, N10467);
xor XOR2 (N10490, N10440, N8304);
and AND3 (N10491, N10486, N2149, N3683);
not NOT1 (N10492, N10491);
xor XOR2 (N10493, N10488, N6880);
xor XOR2 (N10494, N10487, N2388);
not NOT1 (N10495, N10482);
nor NOR2 (N10496, N10493, N5255);
xor XOR2 (N10497, N10494, N326);
xor XOR2 (N10498, N10473, N3372);
and AND3 (N10499, N10485, N328, N2234);
and AND2 (N10500, N10496, N7822);
and AND4 (N10501, N10500, N8511, N10491, N548);
nand NAND2 (N10502, N10489, N8370);
nand NAND4 (N10503, N10497, N2538, N4954, N3867);
buf BUF1 (N10504, N10498);
or OR4 (N10505, N10501, N4885, N4892, N8686);
xor XOR2 (N10506, N10483, N8203);
not NOT1 (N10507, N10503);
or OR4 (N10508, N10506, N7959, N10218, N424);
buf BUF1 (N10509, N10504);
not NOT1 (N10510, N10505);
nand NAND2 (N10511, N10481, N5662);
xor XOR2 (N10512, N10508, N5976);
and AND3 (N10513, N10490, N7601, N7400);
buf BUF1 (N10514, N10512);
xor XOR2 (N10515, N10499, N3449);
and AND4 (N10516, N10511, N4201, N7653, N1107);
not NOT1 (N10517, N10516);
or OR4 (N10518, N10513, N2857, N1514, N6619);
nor NOR3 (N10519, N10517, N1437, N6048);
buf BUF1 (N10520, N10519);
or OR3 (N10521, N10515, N3662, N4013);
xor XOR2 (N10522, N10518, N5801);
or OR3 (N10523, N10495, N543, N3372);
buf BUF1 (N10524, N10514);
nor NOR4 (N10525, N10509, N4310, N2308, N3666);
nor NOR2 (N10526, N10522, N1016);
and AND3 (N10527, N10510, N3046, N321);
not NOT1 (N10528, N10527);
and AND2 (N10529, N10523, N357);
or OR4 (N10530, N10492, N754, N581, N3877);
xor XOR2 (N10531, N10530, N745);
buf BUF1 (N10532, N10507);
not NOT1 (N10533, N10502);
or OR2 (N10534, N10526, N934);
nor NOR3 (N10535, N10524, N7159, N6308);
nand NAND4 (N10536, N10534, N923, N9716, N10454);
xor XOR2 (N10537, N10520, N8876);
and AND3 (N10538, N10521, N439, N2362);
and AND2 (N10539, N10536, N10192);
not NOT1 (N10540, N10531);
nand NAND4 (N10541, N10525, N2914, N6178, N4215);
buf BUF1 (N10542, N10540);
nand NAND3 (N10543, N10535, N8231, N3664);
not NOT1 (N10544, N10532);
not NOT1 (N10545, N10533);
nor NOR3 (N10546, N10542, N5955, N5131);
or OR2 (N10547, N10544, N4718);
not NOT1 (N10548, N10529);
nor NOR4 (N10549, N10539, N1668, N5811, N7226);
nand NAND2 (N10550, N10541, N2732);
nor NOR2 (N10551, N10543, N9485);
buf BUF1 (N10552, N10550);
and AND2 (N10553, N10538, N7428);
xor XOR2 (N10554, N10537, N6987);
nor NOR3 (N10555, N10547, N8920, N7672);
or OR3 (N10556, N10555, N6486, N10460);
and AND2 (N10557, N10549, N2701);
not NOT1 (N10558, N10545);
or OR2 (N10559, N10558, N2633);
buf BUF1 (N10560, N10559);
or OR2 (N10561, N10553, N3878);
nand NAND4 (N10562, N10556, N673, N5612, N2542);
nor NOR2 (N10563, N10557, N3493);
and AND4 (N10564, N10546, N2347, N10359, N2315);
or OR3 (N10565, N10561, N9454, N889);
nor NOR4 (N10566, N10528, N4028, N8107, N7876);
xor XOR2 (N10567, N10566, N1571);
xor XOR2 (N10568, N10565, N5648);
and AND2 (N10569, N10568, N10468);
buf BUF1 (N10570, N10567);
and AND3 (N10571, N10562, N6103, N5468);
and AND4 (N10572, N10564, N8651, N8272, N8323);
or OR3 (N10573, N10563, N7470, N60);
nand NAND2 (N10574, N10572, N2750);
xor XOR2 (N10575, N10554, N5853);
nand NAND4 (N10576, N10569, N2038, N10045, N7276);
not NOT1 (N10577, N10571);
nor NOR2 (N10578, N10551, N7340);
or OR2 (N10579, N10574, N2295);
nand NAND4 (N10580, N10579, N9804, N4253, N6722);
xor XOR2 (N10581, N10577, N2600);
not NOT1 (N10582, N10560);
not NOT1 (N10583, N10573);
or OR2 (N10584, N10582, N4637);
nor NOR2 (N10585, N10581, N6363);
not NOT1 (N10586, N10580);
nand NAND2 (N10587, N10575, N5429);
xor XOR2 (N10588, N10585, N440);
and AND3 (N10589, N10576, N9878, N7502);
nor NOR2 (N10590, N10570, N9894);
nor NOR4 (N10591, N10586, N8356, N4459, N3247);
buf BUF1 (N10592, N10591);
nor NOR2 (N10593, N10583, N7667);
and AND4 (N10594, N10593, N463, N953, N526);
nor NOR2 (N10595, N10552, N6478);
not NOT1 (N10596, N10589);
or OR2 (N10597, N10595, N444);
or OR3 (N10598, N10587, N4157, N5721);
and AND3 (N10599, N10594, N7611, N5871);
nand NAND3 (N10600, N10592, N9605, N1205);
and AND2 (N10601, N10599, N6414);
xor XOR2 (N10602, N10590, N8907);
and AND2 (N10603, N10597, N5731);
xor XOR2 (N10604, N10596, N6181);
xor XOR2 (N10605, N10578, N9624);
xor XOR2 (N10606, N10600, N7560);
and AND3 (N10607, N10584, N2810, N2906);
and AND4 (N10608, N10601, N7266, N9262, N5515);
or OR4 (N10609, N10598, N5709, N7148, N8708);
nand NAND4 (N10610, N10607, N717, N6335, N551);
nand NAND2 (N10611, N10548, N1044);
or OR3 (N10612, N10588, N2576, N9470);
and AND2 (N10613, N10612, N5195);
or OR4 (N10614, N10604, N9868, N4144, N3767);
or OR4 (N10615, N10614, N4856, N4614, N9617);
nor NOR3 (N10616, N10615, N3166, N9810);
not NOT1 (N10617, N10616);
xor XOR2 (N10618, N10610, N3839);
xor XOR2 (N10619, N10609, N7069);
nand NAND3 (N10620, N10611, N3437, N4748);
or OR3 (N10621, N10603, N3946, N1354);
xor XOR2 (N10622, N10613, N1790);
buf BUF1 (N10623, N10606);
or OR3 (N10624, N10621, N1739, N3582);
buf BUF1 (N10625, N10605);
not NOT1 (N10626, N10619);
and AND4 (N10627, N10620, N6043, N9462, N7173);
nand NAND3 (N10628, N10626, N622, N6142);
nor NOR4 (N10629, N10623, N2520, N9304, N4917);
nor NOR2 (N10630, N10618, N1833);
buf BUF1 (N10631, N10608);
not NOT1 (N10632, N10630);
buf BUF1 (N10633, N10632);
buf BUF1 (N10634, N10617);
or OR2 (N10635, N10622, N10553);
and AND4 (N10636, N10628, N2422, N9877, N8546);
or OR4 (N10637, N10631, N4469, N7302, N6468);
and AND3 (N10638, N10633, N575, N2164);
or OR3 (N10639, N10634, N5846, N6253);
not NOT1 (N10640, N10637);
buf BUF1 (N10641, N10638);
nand NAND4 (N10642, N10602, N6178, N2113, N6527);
xor XOR2 (N10643, N10625, N1561);
xor XOR2 (N10644, N10636, N609);
nand NAND4 (N10645, N10635, N10578, N5441, N6991);
not NOT1 (N10646, N10639);
and AND4 (N10647, N10624, N247, N1712, N5908);
not NOT1 (N10648, N10642);
or OR4 (N10649, N10629, N4239, N2634, N4073);
buf BUF1 (N10650, N10649);
xor XOR2 (N10651, N10650, N1383);
buf BUF1 (N10652, N10644);
buf BUF1 (N10653, N10647);
or OR2 (N10654, N10640, N1474);
nand NAND4 (N10655, N10648, N1406, N2193, N10473);
or OR2 (N10656, N10652, N41);
xor XOR2 (N10657, N10643, N9766);
and AND2 (N10658, N10646, N6117);
xor XOR2 (N10659, N10657, N6351);
and AND3 (N10660, N10627, N10651, N4318);
not NOT1 (N10661, N7948);
buf BUF1 (N10662, N10659);
or OR3 (N10663, N10653, N9597, N7802);
buf BUF1 (N10664, N10655);
or OR4 (N10665, N10656, N2683, N2577, N4454);
and AND3 (N10666, N10664, N8453, N3175);
buf BUF1 (N10667, N10654);
not NOT1 (N10668, N10645);
nand NAND2 (N10669, N10660, N1363);
buf BUF1 (N10670, N10663);
or OR3 (N10671, N10666, N9873, N7958);
buf BUF1 (N10672, N10665);
buf BUF1 (N10673, N10658);
nand NAND4 (N10674, N10673, N504, N3196, N8300);
and AND3 (N10675, N10662, N3843, N6306);
xor XOR2 (N10676, N10671, N8303);
nor NOR4 (N10677, N10641, N8582, N277, N5932);
nand NAND4 (N10678, N10670, N3004, N3223, N6027);
or OR4 (N10679, N10678, N1234, N1975, N5786);
nand NAND2 (N10680, N10668, N9666);
buf BUF1 (N10681, N10674);
not NOT1 (N10682, N10672);
nor NOR4 (N10683, N10679, N2219, N567, N8058);
not NOT1 (N10684, N10669);
xor XOR2 (N10685, N10684, N10619);
nor NOR3 (N10686, N10675, N8564, N6546);
buf BUF1 (N10687, N10681);
not NOT1 (N10688, N10677);
buf BUF1 (N10689, N10685);
and AND4 (N10690, N10667, N1304, N4066, N7152);
nor NOR2 (N10691, N10690, N8604);
xor XOR2 (N10692, N10687, N2640);
or OR2 (N10693, N10692, N1883);
buf BUF1 (N10694, N10676);
and AND2 (N10695, N10693, N9518);
and AND2 (N10696, N10695, N1068);
not NOT1 (N10697, N10689);
nor NOR2 (N10698, N10682, N10345);
or OR2 (N10699, N10694, N8273);
buf BUF1 (N10700, N10661);
not NOT1 (N10701, N10696);
nor NOR3 (N10702, N10680, N10467, N9454);
nor NOR4 (N10703, N10697, N3407, N2829, N3422);
nand NAND2 (N10704, N10699, N3673);
nor NOR2 (N10705, N10701, N1702);
nand NAND3 (N10706, N10704, N6062, N9360);
buf BUF1 (N10707, N10698);
buf BUF1 (N10708, N10707);
nor NOR2 (N10709, N10708, N3011);
buf BUF1 (N10710, N10691);
and AND3 (N10711, N10683, N6554, N8727);
and AND3 (N10712, N10711, N1849, N1585);
buf BUF1 (N10713, N10686);
nor NOR2 (N10714, N10700, N8217);
nor NOR2 (N10715, N10710, N7741);
or OR2 (N10716, N10703, N7582);
buf BUF1 (N10717, N10706);
nand NAND3 (N10718, N10714, N10561, N9322);
buf BUF1 (N10719, N10712);
xor XOR2 (N10720, N10705, N1371);
and AND3 (N10721, N10688, N7238, N4453);
not NOT1 (N10722, N10719);
or OR4 (N10723, N10720, N1317, N8937, N2733);
not NOT1 (N10724, N10723);
xor XOR2 (N10725, N10721, N4537);
nor NOR3 (N10726, N10709, N752, N5242);
and AND2 (N10727, N10717, N7396);
not NOT1 (N10728, N10702);
or OR2 (N10729, N10715, N3877);
not NOT1 (N10730, N10722);
or OR4 (N10731, N10727, N6238, N2339, N6771);
and AND4 (N10732, N10716, N10526, N6052, N3139);
or OR3 (N10733, N10729, N1190, N10466);
and AND3 (N10734, N10713, N4308, N4543);
or OR2 (N10735, N10725, N7948);
and AND2 (N10736, N10728, N1090);
not NOT1 (N10737, N10733);
not NOT1 (N10738, N10726);
and AND3 (N10739, N10730, N9697, N8164);
and AND4 (N10740, N10737, N7778, N4393, N5644);
nand NAND2 (N10741, N10734, N10628);
xor XOR2 (N10742, N10731, N1956);
or OR2 (N10743, N10736, N8254);
xor XOR2 (N10744, N10740, N808);
nor NOR3 (N10745, N10718, N2324, N2587);
xor XOR2 (N10746, N10744, N10572);
not NOT1 (N10747, N10732);
and AND2 (N10748, N10743, N10506);
not NOT1 (N10749, N10746);
xor XOR2 (N10750, N10735, N5001);
and AND3 (N10751, N10745, N8772, N9676);
nand NAND3 (N10752, N10750, N4869, N110);
nor NOR2 (N10753, N10747, N2907);
not NOT1 (N10754, N10751);
or OR4 (N10755, N10752, N5637, N9888, N3539);
not NOT1 (N10756, N10754);
and AND4 (N10757, N10739, N4962, N301, N7147);
xor XOR2 (N10758, N10756, N2257);
xor XOR2 (N10759, N10741, N5985);
not NOT1 (N10760, N10758);
xor XOR2 (N10761, N10748, N9617);
xor XOR2 (N10762, N10757, N5651);
and AND2 (N10763, N10759, N3417);
xor XOR2 (N10764, N10742, N2177);
xor XOR2 (N10765, N10763, N8038);
buf BUF1 (N10766, N10765);
xor XOR2 (N10767, N10764, N5053);
and AND2 (N10768, N10766, N3439);
buf BUF1 (N10769, N10761);
not NOT1 (N10770, N10762);
and AND2 (N10771, N10749, N1949);
and AND2 (N10772, N10760, N308);
nor NOR2 (N10773, N10769, N6212);
and AND2 (N10774, N10738, N8651);
and AND3 (N10775, N10772, N6822, N6285);
xor XOR2 (N10776, N10755, N3393);
or OR3 (N10777, N10770, N1692, N4038);
xor XOR2 (N10778, N10767, N4614);
xor XOR2 (N10779, N10776, N7332);
xor XOR2 (N10780, N10724, N8271);
and AND2 (N10781, N10775, N8103);
and AND2 (N10782, N10753, N9545);
and AND3 (N10783, N10780, N3124, N7993);
not NOT1 (N10784, N10771);
nor NOR3 (N10785, N10774, N9370, N7953);
not NOT1 (N10786, N10768);
or OR2 (N10787, N10779, N10068);
buf BUF1 (N10788, N10778);
xor XOR2 (N10789, N10781, N4789);
nand NAND4 (N10790, N10784, N6037, N8787, N10588);
nand NAND4 (N10791, N10773, N3804, N1336, N4191);
or OR3 (N10792, N10783, N7508, N4466);
and AND3 (N10793, N10782, N1437, N5704);
xor XOR2 (N10794, N10792, N6328);
nor NOR4 (N10795, N10785, N6795, N6527, N7284);
buf BUF1 (N10796, N10777);
not NOT1 (N10797, N10794);
xor XOR2 (N10798, N10789, N9970);
not NOT1 (N10799, N10798);
buf BUF1 (N10800, N10796);
not NOT1 (N10801, N10793);
nand NAND4 (N10802, N10790, N6725, N688, N4880);
nor NOR2 (N10803, N10797, N1875);
buf BUF1 (N10804, N10802);
xor XOR2 (N10805, N10803, N4643);
nor NOR4 (N10806, N10795, N10157, N7285, N1412);
nor NOR3 (N10807, N10801, N6603, N3527);
or OR4 (N10808, N10787, N4926, N5749, N10353);
and AND3 (N10809, N10786, N4931, N3144);
nor NOR4 (N10810, N10791, N9589, N4562, N7771);
nand NAND3 (N10811, N10810, N8270, N9986);
not NOT1 (N10812, N10800);
buf BUF1 (N10813, N10808);
and AND2 (N10814, N10806, N8104);
not NOT1 (N10815, N10807);
and AND2 (N10816, N10805, N6265);
not NOT1 (N10817, N10812);
buf BUF1 (N10818, N10813);
or OR4 (N10819, N10818, N3185, N7110, N9221);
not NOT1 (N10820, N10804);
or OR2 (N10821, N10811, N724);
nor NOR3 (N10822, N10815, N1214, N1422);
buf BUF1 (N10823, N10819);
and AND2 (N10824, N10817, N4751);
xor XOR2 (N10825, N10822, N7429);
nand NAND3 (N10826, N10814, N34, N8688);
not NOT1 (N10827, N10816);
nand NAND2 (N10828, N10824, N9519);
nand NAND2 (N10829, N10827, N4540);
and AND3 (N10830, N10823, N2013, N7250);
and AND4 (N10831, N10821, N159, N4693, N8580);
and AND3 (N10832, N10788, N7535, N2365);
or OR4 (N10833, N10799, N9722, N6942, N4188);
not NOT1 (N10834, N10830);
and AND3 (N10835, N10829, N1838, N7625);
nand NAND3 (N10836, N10835, N7886, N3071);
buf BUF1 (N10837, N10826);
or OR2 (N10838, N10825, N7220);
nand NAND4 (N10839, N10836, N8027, N3733, N8313);
nand NAND4 (N10840, N10837, N9261, N7953, N4239);
and AND2 (N10841, N10838, N5901);
xor XOR2 (N10842, N10831, N6651);
buf BUF1 (N10843, N10833);
nor NOR3 (N10844, N10834, N10824, N3361);
xor XOR2 (N10845, N10820, N509);
xor XOR2 (N10846, N10809, N1356);
xor XOR2 (N10847, N10845, N5816);
or OR4 (N10848, N10839, N5654, N1240, N7595);
not NOT1 (N10849, N10844);
or OR4 (N10850, N10841, N5907, N10577, N1796);
not NOT1 (N10851, N10840);
nor NOR4 (N10852, N10847, N3722, N3870, N2424);
or OR2 (N10853, N10849, N387);
buf BUF1 (N10854, N10828);
or OR4 (N10855, N10851, N7989, N4179, N7125);
buf BUF1 (N10856, N10832);
and AND2 (N10857, N10856, N8649);
not NOT1 (N10858, N10854);
nand NAND4 (N10859, N10857, N1185, N2815, N1508);
not NOT1 (N10860, N10850);
not NOT1 (N10861, N10855);
xor XOR2 (N10862, N10846, N3435);
or OR4 (N10863, N10852, N8017, N2138, N8460);
not NOT1 (N10864, N10848);
buf BUF1 (N10865, N10863);
buf BUF1 (N10866, N10865);
nor NOR3 (N10867, N10866, N5230, N3088);
or OR2 (N10868, N10862, N3953);
not NOT1 (N10869, N10867);
or OR3 (N10870, N10858, N5534, N4755);
nand NAND4 (N10871, N10861, N10265, N1025, N5995);
buf BUF1 (N10872, N10871);
and AND3 (N10873, N10870, N2267, N8309);
nor NOR4 (N10874, N10869, N4432, N8009, N1560);
buf BUF1 (N10875, N10873);
and AND4 (N10876, N10842, N189, N2657, N9112);
or OR2 (N10877, N10859, N6956);
nor NOR4 (N10878, N10843, N1782, N6652, N7276);
not NOT1 (N10879, N10864);
nor NOR4 (N10880, N10875, N6905, N7369, N8458);
not NOT1 (N10881, N10880);
xor XOR2 (N10882, N10879, N8747);
or OR2 (N10883, N10868, N2313);
buf BUF1 (N10884, N10860);
not NOT1 (N10885, N10872);
nor NOR3 (N10886, N10884, N5850, N723);
not NOT1 (N10887, N10885);
not NOT1 (N10888, N10876);
nand NAND2 (N10889, N10878, N6810);
buf BUF1 (N10890, N10883);
not NOT1 (N10891, N10887);
buf BUF1 (N10892, N10888);
nand NAND2 (N10893, N10891, N3817);
buf BUF1 (N10894, N10877);
xor XOR2 (N10895, N10892, N10321);
not NOT1 (N10896, N10889);
nand NAND2 (N10897, N10896, N10698);
nor NOR2 (N10898, N10894, N6557);
nor NOR2 (N10899, N10886, N9534);
xor XOR2 (N10900, N10874, N5725);
not NOT1 (N10901, N10893);
or OR4 (N10902, N10853, N10854, N5825, N10679);
not NOT1 (N10903, N10895);
and AND2 (N10904, N10901, N503);
nand NAND3 (N10905, N10899, N9094, N9912);
nor NOR4 (N10906, N10881, N687, N3574, N2900);
nand NAND2 (N10907, N10903, N3758);
and AND2 (N10908, N10902, N1095);
buf BUF1 (N10909, N10897);
not NOT1 (N10910, N10906);
nand NAND3 (N10911, N10905, N162, N971);
nor NOR2 (N10912, N10911, N10709);
and AND4 (N10913, N10909, N10589, N1944, N688);
xor XOR2 (N10914, N10898, N9423);
and AND3 (N10915, N10882, N7980, N4451);
nand NAND3 (N10916, N10914, N134, N1617);
buf BUF1 (N10917, N10907);
nor NOR4 (N10918, N10917, N10639, N10777, N4552);
xor XOR2 (N10919, N10916, N3443);
and AND4 (N10920, N10890, N7842, N10051, N5743);
or OR4 (N10921, N10913, N239, N1765, N8933);
not NOT1 (N10922, N10904);
not NOT1 (N10923, N10920);
not NOT1 (N10924, N10910);
and AND3 (N10925, N10900, N7863, N3603);
buf BUF1 (N10926, N10923);
buf BUF1 (N10927, N10924);
buf BUF1 (N10928, N10908);
and AND2 (N10929, N10915, N10314);
xor XOR2 (N10930, N10927, N5004);
or OR2 (N10931, N10919, N33);
nor NOR2 (N10932, N10912, N615);
not NOT1 (N10933, N10921);
buf BUF1 (N10934, N10922);
or OR2 (N10935, N10933, N925);
xor XOR2 (N10936, N10934, N5084);
or OR2 (N10937, N10930, N3131);
and AND2 (N10938, N10935, N6434);
buf BUF1 (N10939, N10929);
nand NAND4 (N10940, N10939, N3570, N4760, N300);
or OR3 (N10941, N10932, N8473, N211);
nor NOR4 (N10942, N10925, N3069, N7307, N2215);
xor XOR2 (N10943, N10942, N4245);
nand NAND2 (N10944, N10931, N5819);
xor XOR2 (N10945, N10936, N5990);
nor NOR3 (N10946, N10943, N4605, N797);
nor NOR2 (N10947, N10938, N6130);
buf BUF1 (N10948, N10926);
buf BUF1 (N10949, N10918);
buf BUF1 (N10950, N10941);
or OR2 (N10951, N10948, N10641);
and AND3 (N10952, N10947, N5798, N7084);
nor NOR4 (N10953, N10944, N2923, N8956, N3263);
nand NAND3 (N10954, N10945, N10158, N8449);
nand NAND3 (N10955, N10950, N608, N2379);
or OR3 (N10956, N10954, N6297, N7454);
or OR2 (N10957, N10937, N10616);
not NOT1 (N10958, N10951);
not NOT1 (N10959, N10957);
buf BUF1 (N10960, N10959);
nand NAND2 (N10961, N10928, N8284);
nor NOR2 (N10962, N10940, N7564);
nand NAND4 (N10963, N10958, N7094, N6409, N9436);
xor XOR2 (N10964, N10962, N1994);
buf BUF1 (N10965, N10953);
and AND2 (N10966, N10960, N10367);
and AND2 (N10967, N10949, N105);
buf BUF1 (N10968, N10966);
not NOT1 (N10969, N10952);
or OR3 (N10970, N10963, N6911, N4322);
buf BUF1 (N10971, N10946);
or OR3 (N10972, N10970, N6781, N9716);
nand NAND2 (N10973, N10964, N8191);
nand NAND4 (N10974, N10955, N10610, N4141, N8098);
buf BUF1 (N10975, N10974);
not NOT1 (N10976, N10975);
nor NOR3 (N10977, N10972, N4170, N2241);
or OR3 (N10978, N10961, N727, N5989);
and AND4 (N10979, N10973, N7330, N3889, N7056);
and AND4 (N10980, N10965, N2912, N24, N1798);
not NOT1 (N10981, N10967);
buf BUF1 (N10982, N10969);
xor XOR2 (N10983, N10968, N2270);
buf BUF1 (N10984, N10983);
nand NAND3 (N10985, N10979, N907, N10541);
nand NAND4 (N10986, N10956, N3874, N3268, N5987);
xor XOR2 (N10987, N10981, N9011);
xor XOR2 (N10988, N10987, N1004);
nand NAND4 (N10989, N10971, N3603, N9109, N5811);
nand NAND2 (N10990, N10988, N75);
buf BUF1 (N10991, N10985);
not NOT1 (N10992, N10986);
and AND2 (N10993, N10976, N6662);
and AND3 (N10994, N10984, N6119, N7870);
nand NAND2 (N10995, N10994, N2053);
nand NAND2 (N10996, N10990, N90);
or OR2 (N10997, N10991, N10006);
nor NOR3 (N10998, N10992, N8909, N5469);
or OR2 (N10999, N10993, N9901);
xor XOR2 (N11000, N10997, N3645);
xor XOR2 (N11001, N10989, N1211);
buf BUF1 (N11002, N10996);
buf BUF1 (N11003, N11001);
xor XOR2 (N11004, N10982, N383);
or OR2 (N11005, N10977, N10510);
nor NOR4 (N11006, N10999, N8490, N1839, N6470);
nand NAND2 (N11007, N11002, N3431);
nor NOR3 (N11008, N11007, N198, N6666);
not NOT1 (N11009, N11000);
buf BUF1 (N11010, N10978);
nor NOR2 (N11011, N11006, N4713);
nand NAND4 (N11012, N11004, N10790, N10411, N8349);
or OR2 (N11013, N11005, N3457);
nor NOR3 (N11014, N10980, N4237, N5132);
and AND2 (N11015, N11012, N9079);
nand NAND3 (N11016, N11009, N3842, N1363);
xor XOR2 (N11017, N11011, N184);
buf BUF1 (N11018, N11015);
xor XOR2 (N11019, N11017, N4515);
buf BUF1 (N11020, N11008);
nand NAND3 (N11021, N11020, N4722, N9438);
and AND4 (N11022, N11018, N1738, N5488, N10382);
and AND4 (N11023, N11016, N4723, N1174, N7151);
not NOT1 (N11024, N11022);
nand NAND2 (N11025, N10998, N1339);
nand NAND4 (N11026, N11010, N8775, N4953, N51);
not NOT1 (N11027, N11019);
or OR3 (N11028, N10995, N9065, N4468);
and AND3 (N11029, N11023, N4786, N1865);
or OR3 (N11030, N11026, N7912, N5685);
nand NAND2 (N11031, N11027, N7259);
nor NOR4 (N11032, N11030, N6035, N10582, N53);
and AND3 (N11033, N11029, N707, N6141);
not NOT1 (N11034, N11032);
and AND4 (N11035, N11028, N7230, N1899, N8121);
buf BUF1 (N11036, N11025);
nor NOR2 (N11037, N11033, N5076);
and AND4 (N11038, N11034, N3659, N684, N817);
buf BUF1 (N11039, N11003);
or OR3 (N11040, N11013, N4020, N9693);
nand NAND2 (N11041, N11021, N8336);
nor NOR2 (N11042, N11038, N1728);
and AND2 (N11043, N11040, N265);
and AND4 (N11044, N11036, N6397, N2639, N7418);
nor NOR4 (N11045, N11031, N9910, N8855, N4644);
buf BUF1 (N11046, N11045);
nand NAND3 (N11047, N11042, N10481, N1846);
or OR3 (N11048, N11024, N9768, N994);
and AND4 (N11049, N11044, N723, N5038, N9801);
nor NOR2 (N11050, N11043, N886);
and AND4 (N11051, N11048, N4447, N5310, N7151);
and AND2 (N11052, N11014, N7);
buf BUF1 (N11053, N11039);
and AND4 (N11054, N11052, N1994, N546, N8301);
buf BUF1 (N11055, N11047);
xor XOR2 (N11056, N11050, N3086);
and AND2 (N11057, N11037, N5676);
not NOT1 (N11058, N11055);
or OR4 (N11059, N11056, N7117, N4109, N9168);
or OR3 (N11060, N11051, N1901, N411);
not NOT1 (N11061, N11059);
or OR2 (N11062, N11061, N1864);
buf BUF1 (N11063, N11058);
buf BUF1 (N11064, N11049);
buf BUF1 (N11065, N11062);
and AND3 (N11066, N11041, N9631, N10965);
or OR3 (N11067, N11064, N1496, N9750);
xor XOR2 (N11068, N11067, N9489);
nor NOR2 (N11069, N11054, N596);
or OR2 (N11070, N11035, N275);
not NOT1 (N11071, N11066);
buf BUF1 (N11072, N11071);
nand NAND2 (N11073, N11070, N6247);
not NOT1 (N11074, N11072);
or OR2 (N11075, N11073, N10102);
or OR2 (N11076, N11060, N4775);
nor NOR2 (N11077, N11046, N1270);
or OR4 (N11078, N11077, N3959, N595, N10024);
or OR2 (N11079, N11065, N10702);
or OR2 (N11080, N11079, N7333);
or OR2 (N11081, N11078, N4836);
nor NOR3 (N11082, N11074, N3618, N4752);
nor NOR4 (N11083, N11081, N3320, N93, N7734);
or OR2 (N11084, N11069, N4098);
xor XOR2 (N11085, N11080, N2755);
nand NAND3 (N11086, N11082, N3436, N7230);
nor NOR4 (N11087, N11076, N10857, N967, N8549);
and AND2 (N11088, N11085, N1381);
nand NAND3 (N11089, N11075, N3982, N1531);
buf BUF1 (N11090, N11068);
nor NOR4 (N11091, N11057, N1353, N7941, N1186);
xor XOR2 (N11092, N11086, N494);
xor XOR2 (N11093, N11053, N10336);
or OR3 (N11094, N11087, N7173, N2728);
xor XOR2 (N11095, N11091, N10769);
or OR4 (N11096, N11083, N5540, N5030, N2794);
buf BUF1 (N11097, N11084);
and AND3 (N11098, N11063, N7220, N3681);
not NOT1 (N11099, N11094);
nor NOR4 (N11100, N11099, N3889, N6104, N400);
not NOT1 (N11101, N11096);
not NOT1 (N11102, N11088);
buf BUF1 (N11103, N11092);
not NOT1 (N11104, N11090);
and AND2 (N11105, N11104, N3973);
not NOT1 (N11106, N11101);
nand NAND4 (N11107, N11106, N384, N639, N9728);
not NOT1 (N11108, N11100);
xor XOR2 (N11109, N11103, N3434);
and AND4 (N11110, N11105, N1703, N4539, N996);
and AND3 (N11111, N11098, N9177, N1743);
not NOT1 (N11112, N11097);
and AND3 (N11113, N11112, N5164, N3777);
not NOT1 (N11114, N11107);
not NOT1 (N11115, N11110);
nand NAND4 (N11116, N11115, N500, N6661, N3963);
and AND3 (N11117, N11114, N11107, N3825);
and AND3 (N11118, N11109, N2857, N3391);
buf BUF1 (N11119, N11117);
and AND4 (N11120, N11108, N10261, N2155, N1914);
buf BUF1 (N11121, N11113);
nor NOR2 (N11122, N11121, N1272);
nand NAND3 (N11123, N11102, N6867, N385);
and AND3 (N11124, N11123, N6536, N8203);
nor NOR4 (N11125, N11119, N786, N7362, N1164);
not NOT1 (N11126, N11116);
xor XOR2 (N11127, N11095, N3090);
nand NAND4 (N11128, N11093, N947, N2832, N2135);
nor NOR3 (N11129, N11120, N8135, N9415);
buf BUF1 (N11130, N11089);
not NOT1 (N11131, N11130);
or OR4 (N11132, N11122, N715, N7496, N979);
not NOT1 (N11133, N11129);
or OR3 (N11134, N11132, N4334, N9734);
buf BUF1 (N11135, N11128);
or OR4 (N11136, N11131, N4911, N4189, N10580);
and AND3 (N11137, N11136, N3583, N1439);
or OR4 (N11138, N11118, N2789, N8522, N8516);
not NOT1 (N11139, N11111);
nand NAND3 (N11140, N11127, N5535, N5079);
buf BUF1 (N11141, N11135);
not NOT1 (N11142, N11138);
nor NOR3 (N11143, N11137, N3407, N8192);
buf BUF1 (N11144, N11126);
and AND2 (N11145, N11124, N3749);
or OR2 (N11146, N11141, N5446);
nand NAND2 (N11147, N11146, N604);
not NOT1 (N11148, N11144);
nor NOR2 (N11149, N11148, N19);
not NOT1 (N11150, N11143);
buf BUF1 (N11151, N11134);
and AND2 (N11152, N11140, N1339);
nor NOR4 (N11153, N11133, N1591, N5538, N11087);
xor XOR2 (N11154, N11147, N8952);
or OR4 (N11155, N11150, N4570, N8458, N5571);
xor XOR2 (N11156, N11152, N7467);
nand NAND4 (N11157, N11149, N592, N9679, N10023);
buf BUF1 (N11158, N11154);
and AND2 (N11159, N11145, N4234);
nor NOR2 (N11160, N11151, N9702);
or OR4 (N11161, N11142, N4174, N1046, N1051);
nand NAND4 (N11162, N11160, N3299, N6192, N10742);
buf BUF1 (N11163, N11153);
nor NOR3 (N11164, N11139, N6887, N8174);
nor NOR2 (N11165, N11156, N15);
nor NOR3 (N11166, N11155, N7397, N7168);
nand NAND2 (N11167, N11163, N1163);
xor XOR2 (N11168, N11159, N4893);
nor NOR4 (N11169, N11157, N8073, N6263, N3227);
not NOT1 (N11170, N11158);
buf BUF1 (N11171, N11166);
buf BUF1 (N11172, N11171);
or OR4 (N11173, N11125, N9288, N6582, N1738);
and AND4 (N11174, N11161, N11102, N9427, N5209);
buf BUF1 (N11175, N11167);
nor NOR3 (N11176, N11169, N5909, N6576);
xor XOR2 (N11177, N11162, N1159);
nor NOR2 (N11178, N11170, N4427);
nor NOR2 (N11179, N11177, N4150);
xor XOR2 (N11180, N11165, N5887);
nand NAND3 (N11181, N11175, N7978, N4156);
and AND3 (N11182, N11174, N3051, N3755);
nand NAND3 (N11183, N11178, N7979, N5936);
nor NOR4 (N11184, N11173, N2822, N8158, N3798);
not NOT1 (N11185, N11184);
xor XOR2 (N11186, N11179, N8190);
nor NOR2 (N11187, N11172, N8072);
and AND4 (N11188, N11176, N9858, N7824, N2198);
nand NAND2 (N11189, N11185, N3324);
or OR2 (N11190, N11181, N5777);
and AND2 (N11191, N11190, N5850);
or OR4 (N11192, N11188, N5342, N2625, N7467);
buf BUF1 (N11193, N11164);
nand NAND4 (N11194, N11183, N4165, N8589, N1569);
and AND4 (N11195, N11193, N6484, N1491, N9626);
buf BUF1 (N11196, N11168);
not NOT1 (N11197, N11191);
nand NAND3 (N11198, N11196, N8743, N1925);
or OR4 (N11199, N11198, N4103, N4770, N2282);
not NOT1 (N11200, N11189);
nor NOR2 (N11201, N11194, N3856);
nor NOR2 (N11202, N11186, N4741);
buf BUF1 (N11203, N11195);
nor NOR2 (N11204, N11203, N1059);
nand NAND4 (N11205, N11199, N6865, N5261, N6278);
xor XOR2 (N11206, N11204, N5157);
and AND3 (N11207, N11192, N1163, N2260);
and AND4 (N11208, N11202, N5478, N7724, N621);
buf BUF1 (N11209, N11207);
xor XOR2 (N11210, N11187, N313);
or OR4 (N11211, N11208, N4350, N8905, N7642);
xor XOR2 (N11212, N11209, N213);
and AND2 (N11213, N11210, N2625);
xor XOR2 (N11214, N11182, N5333);
nand NAND4 (N11215, N11197, N3957, N628, N9804);
xor XOR2 (N11216, N11215, N5385);
buf BUF1 (N11217, N11214);
buf BUF1 (N11218, N11213);
buf BUF1 (N11219, N11211);
and AND2 (N11220, N11206, N5919);
buf BUF1 (N11221, N11201);
and AND3 (N11222, N11216, N6752, N5993);
or OR4 (N11223, N11217, N5600, N6656, N6322);
xor XOR2 (N11224, N11180, N4136);
nand NAND3 (N11225, N11220, N10248, N4994);
xor XOR2 (N11226, N11222, N10201);
and AND2 (N11227, N11200, N8765);
not NOT1 (N11228, N11225);
not NOT1 (N11229, N11219);
nor NOR3 (N11230, N11223, N3871, N7558);
not NOT1 (N11231, N11227);
or OR2 (N11232, N11212, N7785);
not NOT1 (N11233, N11230);
buf BUF1 (N11234, N11229);
not NOT1 (N11235, N11228);
buf BUF1 (N11236, N11234);
not NOT1 (N11237, N11232);
xor XOR2 (N11238, N11218, N424);
buf BUF1 (N11239, N11233);
not NOT1 (N11240, N11224);
nand NAND4 (N11241, N11239, N3020, N2572, N1333);
not NOT1 (N11242, N11237);
not NOT1 (N11243, N11241);
buf BUF1 (N11244, N11205);
nor NOR3 (N11245, N11226, N9189, N5221);
nand NAND4 (N11246, N11231, N2226, N6061, N9055);
nor NOR4 (N11247, N11246, N7139, N9683, N9910);
or OR4 (N11248, N11247, N3059, N10665, N10950);
nand NAND3 (N11249, N11238, N3222, N2571);
not NOT1 (N11250, N11244);
or OR3 (N11251, N11248, N3423, N10068);
or OR4 (N11252, N11251, N6397, N6800, N9781);
buf BUF1 (N11253, N11252);
and AND3 (N11254, N11236, N2369, N1109);
and AND3 (N11255, N11243, N5051, N10643);
not NOT1 (N11256, N11250);
not NOT1 (N11257, N11235);
nand NAND4 (N11258, N11257, N10627, N2062, N1511);
xor XOR2 (N11259, N11253, N6493);
nand NAND2 (N11260, N11254, N2357);
xor XOR2 (N11261, N11255, N10370);
nand NAND2 (N11262, N11221, N9713);
nor NOR3 (N11263, N11261, N1240, N170);
or OR2 (N11264, N11245, N8832);
or OR4 (N11265, N11264, N2215, N7640, N4922);
or OR4 (N11266, N11258, N10732, N1710, N6777);
nor NOR4 (N11267, N11260, N6015, N392, N9072);
and AND4 (N11268, N11267, N4198, N9192, N3777);
or OR3 (N11269, N11265, N4604, N6337);
nand NAND4 (N11270, N11242, N6252, N7092, N1963);
xor XOR2 (N11271, N11249, N2431);
not NOT1 (N11272, N11266);
not NOT1 (N11273, N11271);
nor NOR3 (N11274, N11270, N6408, N5428);
nand NAND4 (N11275, N11262, N2586, N9987, N7688);
or OR2 (N11276, N11240, N10909);
and AND3 (N11277, N11272, N10687, N3688);
nand NAND3 (N11278, N11275, N992, N1340);
nor NOR3 (N11279, N11276, N7078, N1334);
nor NOR2 (N11280, N11259, N7916);
or OR2 (N11281, N11263, N10464);
xor XOR2 (N11282, N11269, N857);
and AND4 (N11283, N11278, N9234, N10719, N6460);
not NOT1 (N11284, N11279);
or OR4 (N11285, N11256, N3145, N2329, N7714);
xor XOR2 (N11286, N11281, N2332);
nand NAND4 (N11287, N11285, N8954, N3171, N7713);
xor XOR2 (N11288, N11280, N889);
buf BUF1 (N11289, N11287);
not NOT1 (N11290, N11268);
nor NOR2 (N11291, N11282, N10566);
buf BUF1 (N11292, N11273);
nor NOR4 (N11293, N11291, N4073, N4320, N1298);
nand NAND3 (N11294, N11277, N1502, N2721);
nand NAND2 (N11295, N11289, N7355);
not NOT1 (N11296, N11286);
not NOT1 (N11297, N11284);
and AND2 (N11298, N11296, N4067);
buf BUF1 (N11299, N11290);
and AND3 (N11300, N11294, N9239, N10675);
buf BUF1 (N11301, N11299);
not NOT1 (N11302, N11298);
and AND3 (N11303, N11301, N1079, N1984);
not NOT1 (N11304, N11283);
and AND3 (N11305, N11304, N7285, N6223);
buf BUF1 (N11306, N11297);
nor NOR2 (N11307, N11274, N11000);
or OR2 (N11308, N11293, N175);
xor XOR2 (N11309, N11307, N7474);
xor XOR2 (N11310, N11302, N10479);
and AND4 (N11311, N11306, N3605, N4108, N3501);
buf BUF1 (N11312, N11305);
xor XOR2 (N11313, N11310, N6015);
and AND3 (N11314, N11312, N7890, N3026);
nand NAND4 (N11315, N11309, N9255, N3115, N6248);
nor NOR2 (N11316, N11303, N5543);
not NOT1 (N11317, N11314);
nor NOR2 (N11318, N11313, N5240);
buf BUF1 (N11319, N11315);
and AND2 (N11320, N11295, N10154);
nand NAND2 (N11321, N11316, N10320);
not NOT1 (N11322, N11320);
nor NOR3 (N11323, N11311, N9944, N3915);
and AND4 (N11324, N11317, N11171, N10019, N10717);
or OR2 (N11325, N11323, N3337);
nand NAND3 (N11326, N11322, N5192, N7714);
not NOT1 (N11327, N11288);
not NOT1 (N11328, N11327);
and AND3 (N11329, N11319, N1228, N4402);
buf BUF1 (N11330, N11318);
nor NOR4 (N11331, N11292, N10906, N11191, N5042);
and AND4 (N11332, N11324, N8348, N6872, N8618);
xor XOR2 (N11333, N11321, N2155);
xor XOR2 (N11334, N11300, N8654);
not NOT1 (N11335, N11326);
and AND3 (N11336, N11335, N10865, N1048);
nor NOR2 (N11337, N11325, N5389);
or OR4 (N11338, N11329, N5331, N7585, N9308);
xor XOR2 (N11339, N11330, N601);
buf BUF1 (N11340, N11339);
xor XOR2 (N11341, N11308, N5502);
nor NOR3 (N11342, N11338, N1251, N3625);
buf BUF1 (N11343, N11341);
not NOT1 (N11344, N11331);
xor XOR2 (N11345, N11343, N10123);
not NOT1 (N11346, N11336);
or OR3 (N11347, N11337, N8391, N1876);
not NOT1 (N11348, N11340);
buf BUF1 (N11349, N11342);
or OR3 (N11350, N11345, N6404, N4025);
and AND3 (N11351, N11328, N8806, N6983);
buf BUF1 (N11352, N11350);
and AND3 (N11353, N11334, N5535, N5393);
xor XOR2 (N11354, N11332, N2279);
nand NAND3 (N11355, N11346, N4141, N9737);
not NOT1 (N11356, N11349);
and AND3 (N11357, N11356, N8937, N9716);
buf BUF1 (N11358, N11355);
nand NAND2 (N11359, N11352, N10567);
buf BUF1 (N11360, N11347);
and AND3 (N11361, N11333, N9005, N4901);
buf BUF1 (N11362, N11354);
not NOT1 (N11363, N11344);
or OR4 (N11364, N11348, N2461, N4598, N10592);
not NOT1 (N11365, N11362);
or OR2 (N11366, N11364, N11249);
nand NAND3 (N11367, N11365, N8257, N730);
buf BUF1 (N11368, N11358);
nand NAND4 (N11369, N11353, N2381, N10016, N4472);
not NOT1 (N11370, N11357);
or OR2 (N11371, N11369, N269);
nor NOR3 (N11372, N11351, N9647, N9464);
xor XOR2 (N11373, N11371, N3058);
and AND4 (N11374, N11366, N1264, N5178, N1570);
buf BUF1 (N11375, N11373);
not NOT1 (N11376, N11360);
xor XOR2 (N11377, N11361, N9988);
and AND2 (N11378, N11359, N6771);
nor NOR2 (N11379, N11377, N4900);
xor XOR2 (N11380, N11379, N2554);
xor XOR2 (N11381, N11372, N3802);
and AND4 (N11382, N11374, N7189, N8511, N8631);
or OR2 (N11383, N11376, N98);
buf BUF1 (N11384, N11378);
xor XOR2 (N11385, N11382, N3476);
or OR2 (N11386, N11383, N5926);
xor XOR2 (N11387, N11380, N9007);
nand NAND2 (N11388, N11370, N6058);
or OR4 (N11389, N11384, N8129, N6731, N8224);
and AND2 (N11390, N11375, N10441);
and AND4 (N11391, N11386, N3632, N5487, N8207);
xor XOR2 (N11392, N11385, N7838);
buf BUF1 (N11393, N11388);
and AND3 (N11394, N11389, N10361, N7080);
or OR2 (N11395, N11391, N8106);
and AND2 (N11396, N11393, N4842);
or OR4 (N11397, N11392, N2928, N3273, N9147);
nor NOR3 (N11398, N11395, N10937, N9889);
nand NAND2 (N11399, N11398, N958);
nor NOR2 (N11400, N11368, N10520);
or OR4 (N11401, N11367, N5605, N3876, N9740);
or OR2 (N11402, N11387, N2565);
buf BUF1 (N11403, N11397);
nand NAND2 (N11404, N11396, N2975);
xor XOR2 (N11405, N11402, N7673);
buf BUF1 (N11406, N11363);
not NOT1 (N11407, N11403);
or OR3 (N11408, N11407, N10356, N5700);
and AND3 (N11409, N11405, N7194, N159);
buf BUF1 (N11410, N11408);
nor NOR4 (N11411, N11406, N1353, N8699, N3972);
or OR4 (N11412, N11381, N8811, N6836, N2087);
nor NOR3 (N11413, N11390, N5473, N9462);
buf BUF1 (N11414, N11410);
and AND2 (N11415, N11412, N1097);
nor NOR2 (N11416, N11399, N11048);
or OR3 (N11417, N11401, N2072, N9326);
buf BUF1 (N11418, N11400);
xor XOR2 (N11419, N11416, N11343);
nor NOR4 (N11420, N11413, N6211, N3315, N2732);
buf BUF1 (N11421, N11411);
or OR3 (N11422, N11404, N9043, N5377);
nand NAND3 (N11423, N11417, N365, N11);
not NOT1 (N11424, N11419);
or OR3 (N11425, N11424, N5648, N4551);
nand NAND4 (N11426, N11420, N2186, N3879, N7248);
and AND2 (N11427, N11415, N2731);
buf BUF1 (N11428, N11423);
buf BUF1 (N11429, N11426);
nor NOR3 (N11430, N11394, N4378, N1375);
nor NOR2 (N11431, N11427, N7125);
and AND3 (N11432, N11431, N5186, N1405);
or OR2 (N11433, N11414, N1009);
buf BUF1 (N11434, N11422);
nand NAND4 (N11435, N11425, N2756, N10346, N5466);
nand NAND2 (N11436, N11434, N11066);
or OR2 (N11437, N11435, N11230);
not NOT1 (N11438, N11433);
nand NAND4 (N11439, N11418, N2402, N3166, N7840);
nor NOR3 (N11440, N11436, N10086, N6315);
nor NOR4 (N11441, N11440, N2596, N6378, N10169);
buf BUF1 (N11442, N11439);
nor NOR2 (N11443, N11438, N7775);
and AND4 (N11444, N11441, N10605, N5390, N2144);
buf BUF1 (N11445, N11442);
xor XOR2 (N11446, N11444, N3684);
nand NAND4 (N11447, N11437, N9353, N404, N2058);
xor XOR2 (N11448, N11443, N1817);
and AND2 (N11449, N11445, N890);
nor NOR4 (N11450, N11447, N10509, N3258, N1501);
not NOT1 (N11451, N11446);
and AND4 (N11452, N11409, N4852, N8501, N4647);
nor NOR4 (N11453, N11429, N3235, N4462, N2157);
buf BUF1 (N11454, N11453);
nand NAND4 (N11455, N11421, N5949, N5036, N10887);
nand NAND2 (N11456, N11449, N1164);
nor NOR3 (N11457, N11432, N28, N2853);
xor XOR2 (N11458, N11450, N5077);
nand NAND2 (N11459, N11428, N8872);
not NOT1 (N11460, N11430);
buf BUF1 (N11461, N11454);
buf BUF1 (N11462, N11460);
not NOT1 (N11463, N11456);
nor NOR4 (N11464, N11461, N11451, N3475, N5833);
nand NAND4 (N11465, N1143, N2842, N8860, N1333);
nand NAND2 (N11466, N11455, N3612);
xor XOR2 (N11467, N11466, N3643);
or OR3 (N11468, N11452, N9151, N10881);
xor XOR2 (N11469, N11457, N6872);
xor XOR2 (N11470, N11463, N6415);
nor NOR2 (N11471, N11468, N255);
buf BUF1 (N11472, N11462);
buf BUF1 (N11473, N11464);
xor XOR2 (N11474, N11448, N2309);
and AND2 (N11475, N11472, N3202);
nand NAND4 (N11476, N11473, N9365, N10851, N2941);
nand NAND4 (N11477, N11476, N1369, N10736, N4932);
nor NOR3 (N11478, N11459, N79, N9954);
nand NAND3 (N11479, N11469, N9393, N10053);
and AND4 (N11480, N11458, N1095, N7951, N10852);
and AND4 (N11481, N11465, N4919, N2175, N1834);
nor NOR3 (N11482, N11475, N3424, N5829);
nand NAND2 (N11483, N11471, N1712);
nor NOR2 (N11484, N11483, N9019);
nand NAND2 (N11485, N11470, N7922);
nand NAND3 (N11486, N11481, N7711, N8020);
or OR2 (N11487, N11486, N5285);
nand NAND2 (N11488, N11482, N2909);
not NOT1 (N11489, N11488);
buf BUF1 (N11490, N11484);
or OR4 (N11491, N11477, N7291, N6607, N1860);
and AND2 (N11492, N11479, N10629);
or OR3 (N11493, N11490, N4387, N10127);
not NOT1 (N11494, N11487);
nand NAND2 (N11495, N11480, N8639);
and AND4 (N11496, N11485, N5304, N518, N1159);
nand NAND2 (N11497, N11495, N8348);
or OR3 (N11498, N11493, N10159, N8895);
xor XOR2 (N11499, N11491, N7172);
and AND3 (N11500, N11496, N10930, N2422);
not NOT1 (N11501, N11497);
nand NAND2 (N11502, N11498, N6595);
nand NAND2 (N11503, N11501, N3444);
buf BUF1 (N11504, N11500);
xor XOR2 (N11505, N11478, N2092);
buf BUF1 (N11506, N11467);
nand NAND3 (N11507, N11494, N2573, N2883);
xor XOR2 (N11508, N11504, N93);
or OR4 (N11509, N11489, N9415, N1690, N5848);
nand NAND4 (N11510, N11505, N11345, N5656, N8667);
and AND4 (N11511, N11492, N10825, N855, N9925);
or OR2 (N11512, N11474, N9211);
buf BUF1 (N11513, N11509);
xor XOR2 (N11514, N11508, N9758);
buf BUF1 (N11515, N11502);
and AND4 (N11516, N11510, N939, N2265, N564);
or OR4 (N11517, N11514, N8482, N10529, N6040);
xor XOR2 (N11518, N11503, N5560);
buf BUF1 (N11519, N11513);
buf BUF1 (N11520, N11518);
xor XOR2 (N11521, N11517, N904);
nand NAND3 (N11522, N11506, N11273, N9734);
and AND4 (N11523, N11522, N4674, N1392, N10032);
buf BUF1 (N11524, N11519);
nor NOR2 (N11525, N11507, N1435);
and AND4 (N11526, N11512, N7962, N8202, N4909);
not NOT1 (N11527, N11515);
or OR2 (N11528, N11526, N9033);
not NOT1 (N11529, N11516);
buf BUF1 (N11530, N11529);
buf BUF1 (N11531, N11528);
nand NAND3 (N11532, N11523, N2813, N11404);
nand NAND3 (N11533, N11511, N3414, N29);
buf BUF1 (N11534, N11531);
nand NAND4 (N11535, N11520, N9458, N5617, N3855);
nor NOR2 (N11536, N11532, N3092);
nand NAND4 (N11537, N11527, N7948, N7728, N2982);
nor NOR4 (N11538, N11521, N4215, N10497, N1840);
xor XOR2 (N11539, N11538, N5928);
nor NOR2 (N11540, N11499, N10275);
xor XOR2 (N11541, N11535, N1400);
xor XOR2 (N11542, N11540, N4199);
nand NAND2 (N11543, N11539, N9141);
nor NOR4 (N11544, N11534, N2300, N5940, N4052);
and AND2 (N11545, N11542, N1620);
not NOT1 (N11546, N11533);
not NOT1 (N11547, N11536);
not NOT1 (N11548, N11545);
buf BUF1 (N11549, N11524);
not NOT1 (N11550, N11530);
not NOT1 (N11551, N11548);
xor XOR2 (N11552, N11550, N4159);
buf BUF1 (N11553, N11549);
buf BUF1 (N11554, N11537);
nor NOR3 (N11555, N11551, N4245, N10999);
xor XOR2 (N11556, N11553, N4165);
nor NOR4 (N11557, N11541, N8084, N9217, N4282);
not NOT1 (N11558, N11525);
and AND4 (N11559, N11555, N10631, N10923, N8771);
xor XOR2 (N11560, N11543, N4355);
nor NOR2 (N11561, N11554, N10973);
and AND2 (N11562, N11557, N11131);
xor XOR2 (N11563, N11560, N295);
and AND3 (N11564, N11552, N2598, N2964);
buf BUF1 (N11565, N11544);
xor XOR2 (N11566, N11559, N3454);
buf BUF1 (N11567, N11558);
nor NOR4 (N11568, N11564, N10244, N4940, N11214);
nand NAND2 (N11569, N11568, N3885);
or OR2 (N11570, N11546, N7020);
nand NAND3 (N11571, N11562, N2758, N4012);
and AND2 (N11572, N11565, N6368);
or OR2 (N11573, N11563, N4177);
nor NOR2 (N11574, N11571, N9537);
xor XOR2 (N11575, N11566, N8822);
nand NAND3 (N11576, N11570, N8715, N3283);
buf BUF1 (N11577, N11576);
not NOT1 (N11578, N11574);
nor NOR4 (N11579, N11572, N8283, N9010, N8532);
xor XOR2 (N11580, N11569, N11168);
nor NOR3 (N11581, N11575, N5058, N7697);
buf BUF1 (N11582, N11579);
not NOT1 (N11583, N11556);
xor XOR2 (N11584, N11581, N6688);
nand NAND2 (N11585, N11567, N4355);
buf BUF1 (N11586, N11584);
and AND4 (N11587, N11586, N6855, N6312, N3197);
nor NOR3 (N11588, N11547, N10944, N4048);
nand NAND4 (N11589, N11587, N8509, N8641, N8342);
nor NOR3 (N11590, N11577, N4260, N7407);
and AND2 (N11591, N11580, N2000);
and AND2 (N11592, N11589, N4533);
buf BUF1 (N11593, N11588);
or OR4 (N11594, N11561, N8854, N7122, N6332);
nor NOR3 (N11595, N11592, N9053, N8894);
buf BUF1 (N11596, N11578);
nand NAND3 (N11597, N11573, N2437, N10654);
xor XOR2 (N11598, N11597, N4748);
and AND2 (N11599, N11582, N322);
or OR4 (N11600, N11583, N10977, N3417, N191);
nand NAND2 (N11601, N11590, N8118);
nor NOR2 (N11602, N11591, N10201);
nand NAND3 (N11603, N11596, N773, N4251);
nand NAND2 (N11604, N11602, N5686);
and AND4 (N11605, N11603, N269, N10402, N1253);
or OR3 (N11606, N11605, N7293, N7136);
or OR4 (N11607, N11598, N1768, N1032, N9543);
nor NOR2 (N11608, N11585, N6760);
nor NOR4 (N11609, N11600, N8159, N9517, N7788);
nand NAND4 (N11610, N11608, N7806, N713, N8084);
nand NAND3 (N11611, N11593, N4701, N6948);
xor XOR2 (N11612, N11607, N5210);
and AND3 (N11613, N11595, N1940, N10479);
nor NOR4 (N11614, N11599, N5146, N11015, N537);
or OR3 (N11615, N11609, N2185, N248);
xor XOR2 (N11616, N11613, N11598);
nand NAND3 (N11617, N11606, N6193, N8007);
and AND3 (N11618, N11617, N2090, N6684);
nand NAND4 (N11619, N11610, N1244, N2411, N9994);
xor XOR2 (N11620, N11619, N6032);
and AND4 (N11621, N11618, N3936, N4849, N4859);
or OR3 (N11622, N11621, N8358, N2181);
not NOT1 (N11623, N11615);
nand NAND3 (N11624, N11594, N3671, N2109);
nand NAND4 (N11625, N11622, N2225, N541, N11274);
and AND2 (N11626, N11601, N11484);
nand NAND2 (N11627, N11604, N183);
nor NOR4 (N11628, N11611, N2974, N5945, N10279);
xor XOR2 (N11629, N11628, N4927);
xor XOR2 (N11630, N11629, N1247);
buf BUF1 (N11631, N11624);
and AND3 (N11632, N11625, N10019, N7347);
xor XOR2 (N11633, N11616, N10101);
buf BUF1 (N11634, N11623);
and AND4 (N11635, N11632, N6142, N11595, N11195);
buf BUF1 (N11636, N11626);
not NOT1 (N11637, N11634);
nand NAND4 (N11638, N11637, N1674, N6825, N9589);
and AND2 (N11639, N11630, N8048);
and AND2 (N11640, N11612, N839);
nand NAND3 (N11641, N11627, N1691, N589);
or OR4 (N11642, N11640, N439, N9665, N6792);
or OR3 (N11643, N11636, N10443, N9860);
or OR3 (N11644, N11641, N793, N5041);
nor NOR4 (N11645, N11635, N7080, N8507, N536);
nand NAND3 (N11646, N11639, N1177, N8416);
buf BUF1 (N11647, N11620);
and AND3 (N11648, N11645, N1447, N84);
not NOT1 (N11649, N11648);
buf BUF1 (N11650, N11647);
or OR4 (N11651, N11646, N2019, N2290, N3108);
not NOT1 (N11652, N11644);
nand NAND2 (N11653, N11649, N10101);
or OR3 (N11654, N11650, N8115, N9690);
buf BUF1 (N11655, N11653);
nand NAND3 (N11656, N11643, N3875, N4339);
nand NAND4 (N11657, N11631, N4866, N10860, N10572);
not NOT1 (N11658, N11654);
buf BUF1 (N11659, N11651);
nor NOR3 (N11660, N11657, N8368, N1903);
not NOT1 (N11661, N11642);
buf BUF1 (N11662, N11655);
buf BUF1 (N11663, N11658);
or OR2 (N11664, N11659, N8599);
or OR4 (N11665, N11663, N3581, N1085, N9826);
not NOT1 (N11666, N11656);
nand NAND4 (N11667, N11638, N516, N9878, N2645);
xor XOR2 (N11668, N11665, N2989);
not NOT1 (N11669, N11660);
not NOT1 (N11670, N11669);
or OR2 (N11671, N11668, N3631);
nand NAND4 (N11672, N11633, N3106, N1461, N204);
xor XOR2 (N11673, N11614, N6959);
xor XOR2 (N11674, N11671, N7452);
or OR2 (N11675, N11673, N11139);
xor XOR2 (N11676, N11667, N8969);
or OR4 (N11677, N11662, N1348, N11516, N10929);
xor XOR2 (N11678, N11675, N9473);
nand NAND2 (N11679, N11674, N7306);
and AND2 (N11680, N11677, N3149);
and AND3 (N11681, N11664, N5738, N7414);
buf BUF1 (N11682, N11676);
buf BUF1 (N11683, N11661);
not NOT1 (N11684, N11678);
xor XOR2 (N11685, N11682, N2284);
not NOT1 (N11686, N11680);
not NOT1 (N11687, N11666);
buf BUF1 (N11688, N11685);
buf BUF1 (N11689, N11672);
or OR2 (N11690, N11683, N785);
buf BUF1 (N11691, N11681);
and AND2 (N11692, N11652, N2142);
and AND4 (N11693, N11691, N10320, N1317, N782);
or OR2 (N11694, N11692, N9768);
nand NAND2 (N11695, N11693, N11287);
not NOT1 (N11696, N11670);
or OR3 (N11697, N11679, N9680, N10773);
not NOT1 (N11698, N11688);
xor XOR2 (N11699, N11684, N6801);
buf BUF1 (N11700, N11694);
nand NAND2 (N11701, N11697, N438);
xor XOR2 (N11702, N11698, N6429);
and AND3 (N11703, N11690, N3837, N7156);
or OR2 (N11704, N11703, N1269);
not NOT1 (N11705, N11704);
xor XOR2 (N11706, N11700, N9445);
nor NOR2 (N11707, N11701, N11473);
buf BUF1 (N11708, N11696);
xor XOR2 (N11709, N11689, N9306);
buf BUF1 (N11710, N11706);
buf BUF1 (N11711, N11705);
not NOT1 (N11712, N11695);
or OR2 (N11713, N11708, N7503);
nand NAND3 (N11714, N11687, N2908, N8396);
buf BUF1 (N11715, N11710);
nand NAND2 (N11716, N11715, N2006);
nand NAND3 (N11717, N11712, N7979, N9670);
or OR4 (N11718, N11714, N7548, N4662, N652);
nand NAND2 (N11719, N11707, N2915);
not NOT1 (N11720, N11713);
nand NAND4 (N11721, N11718, N4404, N5579, N4921);
nor NOR2 (N11722, N11719, N10385);
buf BUF1 (N11723, N11686);
or OR4 (N11724, N11722, N6848, N8831, N1478);
nor NOR3 (N11725, N11721, N7831, N8569);
and AND2 (N11726, N11717, N4585);
nand NAND4 (N11727, N11726, N9684, N10204, N5881);
xor XOR2 (N11728, N11727, N10634);
or OR4 (N11729, N11728, N3986, N6731, N8258);
or OR4 (N11730, N11724, N10, N3614, N433);
or OR4 (N11731, N11711, N9618, N1350, N7665);
or OR4 (N11732, N11723, N10743, N2662, N9526);
nor NOR4 (N11733, N11732, N7078, N7798, N626);
not NOT1 (N11734, N11730);
or OR3 (N11735, N11716, N7365, N10079);
not NOT1 (N11736, N11735);
or OR2 (N11737, N11702, N148);
nand NAND4 (N11738, N11709, N1205, N6444, N4222);
nor NOR2 (N11739, N11729, N3343);
nor NOR4 (N11740, N11739, N6816, N7386, N7098);
not NOT1 (N11741, N11733);
nor NOR4 (N11742, N11731, N6298, N6183, N9780);
nand NAND4 (N11743, N11720, N4945, N8636, N10841);
not NOT1 (N11744, N11741);
not NOT1 (N11745, N11734);
buf BUF1 (N11746, N11738);
or OR3 (N11747, N11743, N2281, N10716);
not NOT1 (N11748, N11740);
and AND2 (N11749, N11737, N802);
xor XOR2 (N11750, N11744, N10851);
nor NOR3 (N11751, N11699, N9028, N3217);
not NOT1 (N11752, N11745);
nor NOR3 (N11753, N11736, N8524, N6712);
and AND4 (N11754, N11748, N13, N6393, N3250);
and AND3 (N11755, N11746, N10163, N9465);
not NOT1 (N11756, N11747);
xor XOR2 (N11757, N11725, N9322);
and AND4 (N11758, N11750, N1608, N11311, N1731);
buf BUF1 (N11759, N11755);
nor NOR3 (N11760, N11756, N3945, N9964);
nor NOR4 (N11761, N11759, N4362, N5707, N7202);
xor XOR2 (N11762, N11761, N7231);
nor NOR2 (N11763, N11751, N8531);
and AND4 (N11764, N11760, N8147, N2289, N6643);
buf BUF1 (N11765, N11762);
not NOT1 (N11766, N11757);
xor XOR2 (N11767, N11758, N11137);
nor NOR2 (N11768, N11767, N255);
and AND3 (N11769, N11764, N8565, N1734);
buf BUF1 (N11770, N11769);
not NOT1 (N11771, N11763);
or OR3 (N11772, N11749, N10079, N8028);
nor NOR2 (N11773, N11771, N8406);
nand NAND2 (N11774, N11768, N8977);
buf BUF1 (N11775, N11773);
xor XOR2 (N11776, N11752, N1615);
buf BUF1 (N11777, N11772);
nor NOR4 (N11778, N11777, N2609, N846, N4191);
buf BUF1 (N11779, N11774);
xor XOR2 (N11780, N11775, N10457);
or OR3 (N11781, N11765, N6457, N6109);
nand NAND2 (N11782, N11770, N3049);
or OR4 (N11783, N11779, N3870, N585, N1498);
buf BUF1 (N11784, N11783);
and AND4 (N11785, N11776, N10484, N10401, N10461);
nor NOR2 (N11786, N11766, N2418);
xor XOR2 (N11787, N11742, N11682);
or OR3 (N11788, N11754, N6866, N11399);
nand NAND4 (N11789, N11786, N6952, N8343, N4840);
and AND3 (N11790, N11781, N4160, N11106);
xor XOR2 (N11791, N11788, N10510);
nor NOR4 (N11792, N11791, N11254, N5750, N4827);
xor XOR2 (N11793, N11780, N4332);
nand NAND3 (N11794, N11793, N8832, N25);
or OR2 (N11795, N11790, N9932);
and AND3 (N11796, N11782, N11580, N9511);
nor NOR4 (N11797, N11778, N5677, N979, N3882);
buf BUF1 (N11798, N11785);
nand NAND3 (N11799, N11784, N8323, N1810);
nand NAND4 (N11800, N11798, N10114, N10972, N5299);
buf BUF1 (N11801, N11789);
not NOT1 (N11802, N11753);
nor NOR3 (N11803, N11795, N9319, N10947);
nand NAND4 (N11804, N11803, N3676, N11572, N5181);
and AND2 (N11805, N11796, N6415);
xor XOR2 (N11806, N11801, N1832);
nor NOR4 (N11807, N11797, N5567, N10996, N7622);
nand NAND2 (N11808, N11787, N10003);
buf BUF1 (N11809, N11807);
nand NAND2 (N11810, N11799, N182);
or OR2 (N11811, N11794, N11002);
buf BUF1 (N11812, N11804);
not NOT1 (N11813, N11811);
nand NAND2 (N11814, N11802, N3383);
nand NAND4 (N11815, N11800, N1107, N9924, N5446);
nand NAND4 (N11816, N11813, N6628, N9688, N8078);
and AND4 (N11817, N11810, N2552, N10056, N4524);
nand NAND3 (N11818, N11814, N10905, N5824);
not NOT1 (N11819, N11806);
xor XOR2 (N11820, N11792, N4030);
nand NAND2 (N11821, N11809, N5673);
nor NOR3 (N11822, N11821, N11001, N3011);
xor XOR2 (N11823, N11815, N1060);
and AND2 (N11824, N11812, N7278);
xor XOR2 (N11825, N11824, N11270);
buf BUF1 (N11826, N11805);
or OR4 (N11827, N11823, N3909, N2487, N11406);
nand NAND2 (N11828, N11820, N1066);
nor NOR2 (N11829, N11828, N5526);
xor XOR2 (N11830, N11822, N1664);
nand NAND2 (N11831, N11825, N8327);
not NOT1 (N11832, N11830);
or OR2 (N11833, N11817, N4605);
nor NOR4 (N11834, N11829, N6741, N9640, N1717);
nor NOR2 (N11835, N11826, N4600);
not NOT1 (N11836, N11831);
nand NAND3 (N11837, N11816, N904, N4163);
not NOT1 (N11838, N11833);
xor XOR2 (N11839, N11827, N8017);
xor XOR2 (N11840, N11839, N9058);
nor NOR2 (N11841, N11819, N9673);
nor NOR4 (N11842, N11837, N7650, N5204, N1340);
nand NAND4 (N11843, N11834, N8434, N6600, N4418);
not NOT1 (N11844, N11835);
nand NAND3 (N11845, N11808, N2762, N6254);
nand NAND4 (N11846, N11844, N1663, N4474, N10462);
and AND4 (N11847, N11838, N6395, N8083, N269);
buf BUF1 (N11848, N11845);
and AND3 (N11849, N11848, N10030, N7102);
buf BUF1 (N11850, N11843);
or OR4 (N11851, N11836, N8715, N1423, N4706);
or OR2 (N11852, N11847, N5365);
buf BUF1 (N11853, N11832);
xor XOR2 (N11854, N11850, N3645);
xor XOR2 (N11855, N11851, N9664);
or OR4 (N11856, N11840, N9386, N5755, N10814);
not NOT1 (N11857, N11854);
buf BUF1 (N11858, N11846);
buf BUF1 (N11859, N11849);
nor NOR2 (N11860, N11856, N1958);
buf BUF1 (N11861, N11842);
buf BUF1 (N11862, N11858);
not NOT1 (N11863, N11861);
nand NAND2 (N11864, N11859, N820);
or OR2 (N11865, N11818, N8233);
nand NAND3 (N11866, N11863, N1313, N124);
xor XOR2 (N11867, N11862, N4500);
or OR4 (N11868, N11852, N9429, N11866, N2028);
not NOT1 (N11869, N8206);
buf BUF1 (N11870, N11868);
or OR4 (N11871, N11857, N4967, N10436, N2444);
xor XOR2 (N11872, N11853, N11727);
xor XOR2 (N11873, N11864, N4663);
nor NOR2 (N11874, N11871, N8983);
nand NAND4 (N11875, N11874, N1966, N4744, N2789);
or OR4 (N11876, N11860, N6422, N1761, N10148);
or OR2 (N11877, N11873, N6968);
and AND4 (N11878, N11855, N9171, N9624, N9642);
nand NAND4 (N11879, N11872, N4916, N8066, N7337);
xor XOR2 (N11880, N11870, N10520);
nor NOR3 (N11881, N11867, N1720, N10567);
not NOT1 (N11882, N11878);
not NOT1 (N11883, N11879);
nor NOR4 (N11884, N11869, N4832, N7890, N9851);
buf BUF1 (N11885, N11882);
buf BUF1 (N11886, N11884);
nand NAND2 (N11887, N11883, N10672);
or OR4 (N11888, N11880, N1237, N3786, N5777);
not NOT1 (N11889, N11877);
or OR2 (N11890, N11887, N10721);
not NOT1 (N11891, N11881);
or OR2 (N11892, N11841, N10936);
xor XOR2 (N11893, N11891, N1594);
nor NOR2 (N11894, N11876, N3523);
nor NOR4 (N11895, N11892, N10992, N4078, N6398);
and AND2 (N11896, N11893, N3931);
not NOT1 (N11897, N11886);
nand NAND3 (N11898, N11875, N649, N8971);
nor NOR2 (N11899, N11898, N7980);
or OR2 (N11900, N11896, N3041);
buf BUF1 (N11901, N11888);
and AND3 (N11902, N11899, N3884, N8394);
not NOT1 (N11903, N11889);
nor NOR4 (N11904, N11885, N2189, N1819, N2115);
or OR3 (N11905, N11900, N9221, N972);
nor NOR2 (N11906, N11903, N5866);
nor NOR3 (N11907, N11897, N1505, N6213);
xor XOR2 (N11908, N11865, N820);
and AND4 (N11909, N11894, N2061, N4691, N11170);
nor NOR2 (N11910, N11895, N10734);
and AND4 (N11911, N11910, N3093, N10011, N10692);
or OR2 (N11912, N11890, N7358);
and AND3 (N11913, N11906, N9576, N797);
and AND4 (N11914, N11902, N7865, N1765, N9555);
not NOT1 (N11915, N11907);
or OR4 (N11916, N11912, N8767, N7961, N1304);
buf BUF1 (N11917, N11913);
buf BUF1 (N11918, N11916);
or OR2 (N11919, N11901, N4982);
buf BUF1 (N11920, N11918);
buf BUF1 (N11921, N11909);
or OR4 (N11922, N11911, N441, N6966, N7263);
buf BUF1 (N11923, N11922);
xor XOR2 (N11924, N11923, N2071);
or OR3 (N11925, N11921, N816, N2341);
nand NAND4 (N11926, N11905, N4722, N10973, N4860);
or OR2 (N11927, N11920, N1176);
nand NAND4 (N11928, N11908, N11572, N2293, N3070);
buf BUF1 (N11929, N11904);
not NOT1 (N11930, N11928);
xor XOR2 (N11931, N11915, N7350);
nor NOR2 (N11932, N11927, N4551);
nor NOR4 (N11933, N11931, N7656, N2616, N9525);
or OR3 (N11934, N11919, N2358, N1372);
and AND2 (N11935, N11925, N7656);
xor XOR2 (N11936, N11924, N2219);
nor NOR2 (N11937, N11930, N6470);
xor XOR2 (N11938, N11937, N2914);
nor NOR3 (N11939, N11936, N5118, N1236);
or OR3 (N11940, N11939, N2329, N6265);
nand NAND3 (N11941, N11932, N1954, N11391);
and AND2 (N11942, N11938, N1335);
nor NOR2 (N11943, N11940, N3433);
or OR4 (N11944, N11941, N2340, N11885, N1459);
nor NOR2 (N11945, N11914, N2839);
buf BUF1 (N11946, N11944);
nor NOR2 (N11947, N11945, N5131);
or OR3 (N11948, N11926, N3984, N5148);
not NOT1 (N11949, N11933);
xor XOR2 (N11950, N11948, N4065);
xor XOR2 (N11951, N11950, N1700);
or OR2 (N11952, N11929, N8319);
xor XOR2 (N11953, N11934, N1056);
nor NOR2 (N11954, N11949, N8115);
buf BUF1 (N11955, N11953);
xor XOR2 (N11956, N11942, N9422);
and AND4 (N11957, N11956, N4690, N10115, N6806);
xor XOR2 (N11958, N11954, N4194);
xor XOR2 (N11959, N11943, N4808);
and AND3 (N11960, N11958, N7674, N1572);
or OR2 (N11961, N11955, N994);
xor XOR2 (N11962, N11957, N2014);
nand NAND3 (N11963, N11935, N3969, N11717);
nand NAND3 (N11964, N11960, N3658, N2916);
or OR2 (N11965, N11951, N11920);
nand NAND2 (N11966, N11947, N7010);
and AND4 (N11967, N11963, N8404, N8117, N3848);
xor XOR2 (N11968, N11946, N5714);
buf BUF1 (N11969, N11965);
nand NAND4 (N11970, N11964, N3399, N8714, N7120);
nand NAND3 (N11971, N11966, N3599, N2578);
nand NAND2 (N11972, N11959, N7845);
nor NOR3 (N11973, N11972, N2518, N2368);
nand NAND3 (N11974, N11917, N778, N11880);
and AND2 (N11975, N11961, N8102);
and AND4 (N11976, N11971, N11630, N5087, N1950);
or OR3 (N11977, N11969, N7631, N8231);
not NOT1 (N11978, N11973);
not NOT1 (N11979, N11968);
and AND2 (N11980, N11977, N11499);
not NOT1 (N11981, N11979);
not NOT1 (N11982, N11976);
and AND2 (N11983, N11974, N9365);
nor NOR4 (N11984, N11952, N7387, N4225, N396);
nand NAND2 (N11985, N11962, N8755);
or OR4 (N11986, N11981, N11060, N981, N9553);
and AND4 (N11987, N11984, N11140, N10919, N4837);
not NOT1 (N11988, N11986);
buf BUF1 (N11989, N11978);
or OR4 (N11990, N11985, N3947, N3541, N8752);
nand NAND3 (N11991, N11988, N6784, N3504);
xor XOR2 (N11992, N11970, N6560);
nand NAND4 (N11993, N11989, N4676, N3084, N4254);
or OR4 (N11994, N11983, N6221, N1242, N4898);
buf BUF1 (N11995, N11982);
not NOT1 (N11996, N11992);
and AND2 (N11997, N11987, N6576);
or OR4 (N11998, N11967, N7491, N1069, N4389);
nand NAND2 (N11999, N11994, N8555);
and AND3 (N12000, N11996, N6330, N9397);
xor XOR2 (N12001, N11997, N1615);
buf BUF1 (N12002, N12001);
or OR3 (N12003, N11999, N4020, N178);
or OR3 (N12004, N11993, N8368, N2979);
or OR2 (N12005, N11975, N7617);
not NOT1 (N12006, N11995);
nand NAND2 (N12007, N11998, N826);
buf BUF1 (N12008, N12007);
not NOT1 (N12009, N11980);
nand NAND3 (N12010, N12009, N9180, N11386);
nand NAND4 (N12011, N12003, N7565, N4146, N10708);
buf BUF1 (N12012, N12010);
buf BUF1 (N12013, N11991);
nor NOR3 (N12014, N12006, N11838, N5932);
nor NOR4 (N12015, N12013, N5552, N971, N4481);
or OR3 (N12016, N12008, N5383, N3681);
not NOT1 (N12017, N12016);
not NOT1 (N12018, N12012);
xor XOR2 (N12019, N12005, N9449);
or OR4 (N12020, N12002, N1957, N4832, N9951);
and AND2 (N12021, N12011, N6825);
or OR4 (N12022, N12021, N10870, N6774, N1977);
buf BUF1 (N12023, N12000);
or OR4 (N12024, N12020, N7759, N2170, N3081);
not NOT1 (N12025, N12023);
and AND3 (N12026, N12014, N2399, N1688);
and AND4 (N12027, N12025, N3000, N10689, N171);
xor XOR2 (N12028, N12024, N7976);
buf BUF1 (N12029, N11990);
not NOT1 (N12030, N12022);
xor XOR2 (N12031, N12030, N4007);
nand NAND3 (N12032, N12004, N9755, N7512);
and AND3 (N12033, N12028, N9843, N6950);
nor NOR4 (N12034, N12019, N460, N4627, N1663);
and AND4 (N12035, N12031, N3328, N4423, N9553);
not NOT1 (N12036, N12017);
nor NOR4 (N12037, N12036, N6474, N2123, N10934);
nor NOR3 (N12038, N12015, N1712, N3858);
xor XOR2 (N12039, N12029, N603);
buf BUF1 (N12040, N12027);
not NOT1 (N12041, N12039);
nand NAND3 (N12042, N12035, N3276, N1811);
xor XOR2 (N12043, N12018, N6915);
buf BUF1 (N12044, N12038);
and AND3 (N12045, N12040, N6216, N3737);
nor NOR2 (N12046, N12041, N6144);
xor XOR2 (N12047, N12045, N6472);
buf BUF1 (N12048, N12046);
and AND3 (N12049, N12047, N7566, N1305);
nor NOR4 (N12050, N12032, N11340, N1016, N4065);
and AND4 (N12051, N12033, N3873, N10450, N3312);
xor XOR2 (N12052, N12051, N292);
or OR3 (N12053, N12044, N7380, N1022);
or OR4 (N12054, N12049, N5559, N8322, N6056);
nor NOR4 (N12055, N12054, N10182, N11610, N10264);
not NOT1 (N12056, N12042);
not NOT1 (N12057, N12056);
buf BUF1 (N12058, N12037);
xor XOR2 (N12059, N12034, N7917);
nor NOR2 (N12060, N12059, N8208);
nor NOR2 (N12061, N12057, N3877);
or OR3 (N12062, N12055, N1010, N10891);
not NOT1 (N12063, N12052);
or OR3 (N12064, N12060, N7739, N6042);
nand NAND3 (N12065, N12053, N3940, N1563);
and AND2 (N12066, N12050, N2596);
not NOT1 (N12067, N12043);
xor XOR2 (N12068, N12026, N7288);
nand NAND3 (N12069, N12064, N7802, N2246);
xor XOR2 (N12070, N12063, N173);
buf BUF1 (N12071, N12048);
buf BUF1 (N12072, N12062);
nand NAND4 (N12073, N12070, N6153, N9876, N7129);
or OR4 (N12074, N12071, N1479, N6039, N11804);
or OR2 (N12075, N12073, N2100);
buf BUF1 (N12076, N12067);
and AND3 (N12077, N12074, N10312, N7321);
and AND2 (N12078, N12069, N9402);
nor NOR2 (N12079, N12077, N10186);
or OR3 (N12080, N12079, N2606, N8318);
nand NAND3 (N12081, N12072, N3358, N6236);
buf BUF1 (N12082, N12080);
nand NAND4 (N12083, N12082, N9759, N11749, N4383);
xor XOR2 (N12084, N12083, N10955);
not NOT1 (N12085, N12078);
xor XOR2 (N12086, N12075, N1709);
and AND4 (N12087, N12085, N1097, N11577, N9890);
and AND3 (N12088, N12086, N6343, N9763);
or OR2 (N12089, N12065, N9981);
xor XOR2 (N12090, N12066, N1151);
nand NAND3 (N12091, N12089, N8012, N2245);
not NOT1 (N12092, N12088);
xor XOR2 (N12093, N12081, N2077);
buf BUF1 (N12094, N12084);
nand NAND4 (N12095, N12093, N4479, N6570, N6301);
nand NAND3 (N12096, N12061, N11507, N3262);
buf BUF1 (N12097, N12091);
nand NAND4 (N12098, N12087, N4767, N7400, N7724);
xor XOR2 (N12099, N12096, N5825);
or OR2 (N12100, N12092, N8782);
buf BUF1 (N12101, N12098);
not NOT1 (N12102, N12095);
not NOT1 (N12103, N12058);
and AND4 (N12104, N12094, N3150, N10887, N867);
xor XOR2 (N12105, N12100, N6722);
not NOT1 (N12106, N12103);
xor XOR2 (N12107, N12090, N4711);
and AND4 (N12108, N12097, N6568, N2887, N9145);
not NOT1 (N12109, N12104);
or OR2 (N12110, N12101, N3852);
buf BUF1 (N12111, N12099);
not NOT1 (N12112, N12110);
nor NOR2 (N12113, N12106, N5947);
not NOT1 (N12114, N12109);
buf BUF1 (N12115, N12068);
nand NAND3 (N12116, N12076, N3435, N1323);
or OR4 (N12117, N12111, N5166, N4943, N2388);
xor XOR2 (N12118, N12116, N7848);
nand NAND2 (N12119, N12115, N1608);
nand NAND4 (N12120, N12102, N4187, N6571, N11856);
nand NAND3 (N12121, N12108, N1187, N11097);
nand NAND3 (N12122, N12113, N3556, N7220);
not NOT1 (N12123, N12107);
or OR3 (N12124, N12117, N6875, N8949);
not NOT1 (N12125, N12114);
buf BUF1 (N12126, N12120);
nand NAND3 (N12127, N12124, N11885, N1175);
nor NOR2 (N12128, N12127, N4720);
buf BUF1 (N12129, N12123);
or OR2 (N12130, N12119, N2998);
or OR3 (N12131, N12129, N6712, N5382);
not NOT1 (N12132, N12131);
nand NAND2 (N12133, N12118, N8399);
not NOT1 (N12134, N12112);
nor NOR4 (N12135, N12130, N8408, N5523, N6710);
or OR3 (N12136, N12126, N51, N9065);
buf BUF1 (N12137, N12132);
nor NOR2 (N12138, N12128, N7474);
nand NAND2 (N12139, N12105, N4741);
not NOT1 (N12140, N12139);
or OR4 (N12141, N12125, N10194, N7303, N7447);
and AND3 (N12142, N12122, N8471, N6459);
nand NAND2 (N12143, N12137, N148);
not NOT1 (N12144, N12134);
nor NOR2 (N12145, N12121, N5718);
not NOT1 (N12146, N12141);
or OR4 (N12147, N12145, N5794, N5907, N7201);
nand NAND3 (N12148, N12136, N5094, N1276);
buf BUF1 (N12149, N12147);
and AND4 (N12150, N12146, N9101, N426, N3507);
nor NOR4 (N12151, N12144, N6335, N2591, N10075);
or OR4 (N12152, N12149, N8155, N5397, N2558);
nor NOR3 (N12153, N12151, N3930, N11477);
nand NAND3 (N12154, N12138, N7135, N1382);
buf BUF1 (N12155, N12153);
or OR2 (N12156, N12154, N4674);
or OR3 (N12157, N12140, N342, N4256);
nor NOR3 (N12158, N12156, N352, N9068);
not NOT1 (N12159, N12158);
xor XOR2 (N12160, N12135, N1032);
not NOT1 (N12161, N12142);
xor XOR2 (N12162, N12160, N11601);
nor NOR3 (N12163, N12162, N3222, N3181);
not NOT1 (N12164, N12163);
and AND4 (N12165, N12143, N1471, N2385, N2356);
or OR2 (N12166, N12150, N355);
and AND2 (N12167, N12133, N5522);
buf BUF1 (N12168, N12167);
buf BUF1 (N12169, N12155);
xor XOR2 (N12170, N12169, N3635);
nand NAND2 (N12171, N12165, N9734);
nand NAND2 (N12172, N12148, N2172);
or OR3 (N12173, N12166, N2840, N9927);
or OR2 (N12174, N12172, N7862);
nor NOR4 (N12175, N12161, N858, N5604, N5032);
nor NOR4 (N12176, N12159, N4038, N5345, N9407);
or OR2 (N12177, N12168, N4817);
buf BUF1 (N12178, N12177);
nor NOR4 (N12179, N12175, N498, N905, N7641);
or OR2 (N12180, N12164, N8832);
nor NOR4 (N12181, N12174, N7009, N11653, N11421);
buf BUF1 (N12182, N12152);
and AND3 (N12183, N12157, N6755, N3554);
xor XOR2 (N12184, N12183, N1149);
not NOT1 (N12185, N12173);
and AND3 (N12186, N12182, N11281, N10982);
not NOT1 (N12187, N12176);
and AND3 (N12188, N12171, N7530, N10922);
or OR2 (N12189, N12185, N6964);
nand NAND2 (N12190, N12189, N3482);
xor XOR2 (N12191, N12181, N8014);
or OR3 (N12192, N12191, N913, N5815);
nand NAND4 (N12193, N12184, N7336, N9856, N7125);
nor NOR2 (N12194, N12180, N2904);
not NOT1 (N12195, N12186);
xor XOR2 (N12196, N12188, N1485);
and AND3 (N12197, N12196, N7477, N7150);
nor NOR3 (N12198, N12194, N800, N9816);
buf BUF1 (N12199, N12179);
not NOT1 (N12200, N12198);
nand NAND3 (N12201, N12170, N1990, N1109);
and AND2 (N12202, N12192, N1719);
buf BUF1 (N12203, N12200);
and AND3 (N12204, N12178, N3147, N3761);
nor NOR4 (N12205, N12190, N10665, N6444, N9124);
xor XOR2 (N12206, N12201, N5744);
buf BUF1 (N12207, N12204);
xor XOR2 (N12208, N12203, N406);
or OR3 (N12209, N12202, N10642, N4823);
xor XOR2 (N12210, N12205, N4325);
xor XOR2 (N12211, N12195, N10457);
buf BUF1 (N12212, N12210);
xor XOR2 (N12213, N12209, N4100);
buf BUF1 (N12214, N12213);
xor XOR2 (N12215, N12197, N9334);
or OR2 (N12216, N12193, N1838);
not NOT1 (N12217, N12207);
xor XOR2 (N12218, N12208, N12163);
or OR2 (N12219, N12212, N11374);
nor NOR3 (N12220, N12211, N3939, N5027);
xor XOR2 (N12221, N12217, N11311);
xor XOR2 (N12222, N12199, N9442);
nor NOR4 (N12223, N12220, N8607, N720, N8705);
nand NAND2 (N12224, N12216, N9360);
xor XOR2 (N12225, N12206, N867);
or OR4 (N12226, N12214, N1563, N5709, N1132);
xor XOR2 (N12227, N12215, N10937);
not NOT1 (N12228, N12224);
nand NAND2 (N12229, N12226, N8041);
nor NOR2 (N12230, N12187, N10768);
nand NAND2 (N12231, N12218, N1776);
not NOT1 (N12232, N12222);
not NOT1 (N12233, N12231);
not NOT1 (N12234, N12225);
buf BUF1 (N12235, N12229);
nor NOR4 (N12236, N12230, N4322, N8364, N9006);
or OR2 (N12237, N12227, N4617);
and AND4 (N12238, N12237, N8668, N11879, N4101);
or OR3 (N12239, N12238, N10992, N4623);
buf BUF1 (N12240, N12219);
buf BUF1 (N12241, N12233);
or OR4 (N12242, N12223, N3368, N3088, N2895);
buf BUF1 (N12243, N12236);
nor NOR2 (N12244, N12242, N7646);
and AND4 (N12245, N12244, N10432, N492, N3480);
or OR4 (N12246, N12243, N1221, N3745, N703);
nor NOR3 (N12247, N12235, N5147, N12140);
and AND2 (N12248, N12245, N9552);
xor XOR2 (N12249, N12241, N1207);
xor XOR2 (N12250, N12232, N1547);
or OR4 (N12251, N12240, N3738, N1372, N2473);
xor XOR2 (N12252, N12239, N826);
or OR3 (N12253, N12252, N9158, N5440);
nor NOR4 (N12254, N12221, N5758, N2061, N2633);
buf BUF1 (N12255, N12246);
or OR4 (N12256, N12253, N3074, N5748, N11710);
not NOT1 (N12257, N12247);
nand NAND3 (N12258, N12249, N1863, N9297);
not NOT1 (N12259, N12250);
buf BUF1 (N12260, N12259);
nor NOR2 (N12261, N12260, N7256);
xor XOR2 (N12262, N12255, N1325);
or OR2 (N12263, N12254, N2141);
xor XOR2 (N12264, N12263, N9502);
nor NOR3 (N12265, N12256, N2204, N5993);
buf BUF1 (N12266, N12264);
nand NAND3 (N12267, N12261, N6237, N5225);
xor XOR2 (N12268, N12266, N4466);
or OR3 (N12269, N12265, N5801, N6901);
buf BUF1 (N12270, N12258);
and AND3 (N12271, N12251, N3580, N1178);
xor XOR2 (N12272, N12228, N10662);
buf BUF1 (N12273, N12270);
xor XOR2 (N12274, N12234, N6379);
not NOT1 (N12275, N12269);
and AND4 (N12276, N12272, N3629, N3842, N8829);
or OR3 (N12277, N12262, N3871, N12112);
xor XOR2 (N12278, N12271, N10480);
and AND3 (N12279, N12267, N6246, N5504);
xor XOR2 (N12280, N12274, N3660);
buf BUF1 (N12281, N12268);
buf BUF1 (N12282, N12257);
xor XOR2 (N12283, N12276, N11745);
buf BUF1 (N12284, N12283);
xor XOR2 (N12285, N12278, N3426);
nand NAND2 (N12286, N12248, N2746);
nor NOR2 (N12287, N12275, N5450);
xor XOR2 (N12288, N12279, N1004);
not NOT1 (N12289, N12280);
xor XOR2 (N12290, N12282, N8527);
xor XOR2 (N12291, N12288, N636);
not NOT1 (N12292, N12284);
not NOT1 (N12293, N12290);
nor NOR4 (N12294, N12289, N7968, N12067, N8891);
and AND2 (N12295, N12292, N6997);
xor XOR2 (N12296, N12295, N206);
and AND4 (N12297, N12273, N5008, N4750, N2992);
or OR4 (N12298, N12281, N10842, N636, N7521);
and AND4 (N12299, N12298, N4722, N8520, N3127);
not NOT1 (N12300, N12286);
buf BUF1 (N12301, N12285);
buf BUF1 (N12302, N12277);
nand NAND2 (N12303, N12294, N6491);
nand NAND4 (N12304, N12299, N5266, N5483, N6741);
nand NAND4 (N12305, N12297, N11222, N3090, N9905);
not NOT1 (N12306, N12293);
and AND4 (N12307, N12301, N10329, N6541, N6114);
or OR3 (N12308, N12306, N93, N9173);
and AND3 (N12309, N12308, N10273, N3475);
xor XOR2 (N12310, N12309, N5727);
or OR3 (N12311, N12287, N7656, N1574);
xor XOR2 (N12312, N12307, N2372);
buf BUF1 (N12313, N12311);
nor NOR3 (N12314, N12300, N3205, N1755);
nor NOR2 (N12315, N12304, N9768);
and AND2 (N12316, N12310, N7955);
xor XOR2 (N12317, N12305, N4210);
nand NAND3 (N12318, N12291, N12007, N10665);
buf BUF1 (N12319, N12317);
nor NOR2 (N12320, N12315, N6315);
nor NOR2 (N12321, N12318, N2336);
not NOT1 (N12322, N12313);
or OR4 (N12323, N12322, N4081, N2803, N5265);
nor NOR4 (N12324, N12312, N2574, N4830, N6433);
xor XOR2 (N12325, N12302, N11475);
xor XOR2 (N12326, N12323, N10537);
nor NOR3 (N12327, N12314, N4361, N2977);
and AND3 (N12328, N12320, N8236, N11511);
or OR4 (N12329, N12303, N9866, N1165, N9430);
xor XOR2 (N12330, N12319, N5286);
nand NAND4 (N12331, N12326, N4752, N12257, N4411);
nor NOR2 (N12332, N12316, N516);
buf BUF1 (N12333, N12329);
and AND4 (N12334, N12325, N10196, N4227, N12150);
nand NAND2 (N12335, N12328, N4523);
or OR2 (N12336, N12324, N8482);
or OR2 (N12337, N12327, N6583);
nor NOR4 (N12338, N12333, N10682, N2210, N1660);
nor NOR4 (N12339, N12338, N6468, N8798, N9644);
and AND4 (N12340, N12335, N7245, N7749, N8397);
buf BUF1 (N12341, N12296);
xor XOR2 (N12342, N12339, N10203);
nand NAND3 (N12343, N12334, N3005, N2386);
xor XOR2 (N12344, N12341, N9669);
nor NOR2 (N12345, N12331, N8914);
xor XOR2 (N12346, N12336, N4085);
and AND4 (N12347, N12343, N6661, N2734, N6301);
and AND2 (N12348, N12347, N202);
not NOT1 (N12349, N12346);
nand NAND2 (N12350, N12321, N7114);
xor XOR2 (N12351, N12344, N7924);
nand NAND3 (N12352, N12348, N9647, N3156);
not NOT1 (N12353, N12345);
and AND3 (N12354, N12350, N3397, N7029);
not NOT1 (N12355, N12342);
nand NAND2 (N12356, N12340, N5115);
not NOT1 (N12357, N12356);
and AND2 (N12358, N12357, N1733);
not NOT1 (N12359, N12330);
or OR4 (N12360, N12351, N8072, N10627, N4020);
not NOT1 (N12361, N12337);
buf BUF1 (N12362, N12360);
buf BUF1 (N12363, N12349);
xor XOR2 (N12364, N12355, N995);
or OR2 (N12365, N12358, N1162);
and AND4 (N12366, N12359, N5949, N7798, N7215);
nor NOR3 (N12367, N12363, N9173, N1812);
nor NOR3 (N12368, N12353, N11096, N6466);
or OR4 (N12369, N12364, N10869, N11183, N5400);
or OR3 (N12370, N12352, N7284, N3786);
xor XOR2 (N12371, N12367, N12262);
nor NOR4 (N12372, N12365, N2172, N647, N202);
xor XOR2 (N12373, N12362, N5176);
not NOT1 (N12374, N12373);
or OR3 (N12375, N12368, N4606, N662);
nor NOR3 (N12376, N12370, N2130, N9096);
not NOT1 (N12377, N12366);
xor XOR2 (N12378, N12375, N112);
xor XOR2 (N12379, N12371, N8803);
not NOT1 (N12380, N12372);
and AND2 (N12381, N12379, N6073);
nand NAND3 (N12382, N12381, N751, N1613);
buf BUF1 (N12383, N12382);
or OR2 (N12384, N12376, N3383);
buf BUF1 (N12385, N12332);
xor XOR2 (N12386, N12384, N9996);
or OR2 (N12387, N12385, N10493);
xor XOR2 (N12388, N12386, N1580);
and AND4 (N12389, N12369, N4929, N9765, N8632);
not NOT1 (N12390, N12383);
xor XOR2 (N12391, N12377, N2782);
xor XOR2 (N12392, N12391, N4404);
xor XOR2 (N12393, N12390, N9377);
xor XOR2 (N12394, N12354, N10150);
nor NOR2 (N12395, N12374, N2342);
nand NAND4 (N12396, N12394, N8038, N7773, N1507);
buf BUF1 (N12397, N12395);
and AND3 (N12398, N12388, N4828, N3723);
xor XOR2 (N12399, N12396, N1429);
xor XOR2 (N12400, N12392, N2363);
not NOT1 (N12401, N12389);
buf BUF1 (N12402, N12387);
nand NAND3 (N12403, N12399, N8699, N3140);
buf BUF1 (N12404, N12397);
xor XOR2 (N12405, N12404, N9559);
xor XOR2 (N12406, N12361, N9166);
nor NOR3 (N12407, N12405, N1269, N7684);
or OR2 (N12408, N12378, N4534);
xor XOR2 (N12409, N12393, N1336);
and AND3 (N12410, N12407, N4619, N5241);
not NOT1 (N12411, N12406);
not NOT1 (N12412, N12380);
and AND2 (N12413, N12409, N892);
nand NAND3 (N12414, N12408, N3216, N12237);
or OR2 (N12415, N12410, N7643);
and AND3 (N12416, N12411, N10172, N6580);
or OR3 (N12417, N12401, N11410, N10806);
not NOT1 (N12418, N12413);
xor XOR2 (N12419, N12418, N7512);
nor NOR3 (N12420, N12415, N2169, N9496);
or OR4 (N12421, N12398, N5754, N11754, N10214);
not NOT1 (N12422, N12414);
or OR2 (N12423, N12400, N193);
and AND3 (N12424, N12416, N11367, N10856);
buf BUF1 (N12425, N12424);
buf BUF1 (N12426, N12422);
buf BUF1 (N12427, N12425);
or OR3 (N12428, N12417, N10815, N8637);
or OR3 (N12429, N12419, N9711, N10561);
nor NOR4 (N12430, N12429, N11742, N935, N2968);
or OR3 (N12431, N12402, N4439, N5837);
buf BUF1 (N12432, N12421);
nand NAND4 (N12433, N12423, N8155, N7775, N10872);
nand NAND4 (N12434, N12431, N10260, N12217, N5038);
or OR4 (N12435, N12427, N2681, N11294, N11049);
nand NAND4 (N12436, N12426, N11999, N7837, N2051);
nand NAND3 (N12437, N12430, N7118, N539);
and AND3 (N12438, N12434, N4517, N10570);
xor XOR2 (N12439, N12432, N10375);
xor XOR2 (N12440, N12438, N3432);
xor XOR2 (N12441, N12433, N8007);
xor XOR2 (N12442, N12435, N10267);
not NOT1 (N12443, N12437);
buf BUF1 (N12444, N12441);
and AND3 (N12445, N12442, N9099, N2821);
nand NAND3 (N12446, N12443, N5276, N6102);
buf BUF1 (N12447, N12439);
and AND3 (N12448, N12440, N1344, N6930);
not NOT1 (N12449, N12446);
or OR3 (N12450, N12436, N3122, N537);
nor NOR2 (N12451, N12428, N4190);
buf BUF1 (N12452, N12448);
or OR2 (N12453, N12450, N1338);
nor NOR2 (N12454, N12412, N7090);
xor XOR2 (N12455, N12445, N4178);
and AND4 (N12456, N12452, N11813, N9006, N3638);
nor NOR4 (N12457, N12451, N10335, N7786, N8016);
nor NOR4 (N12458, N12457, N2013, N1998, N1275);
xor XOR2 (N12459, N12454, N12339);
nand NAND2 (N12460, N12458, N6653);
nor NOR2 (N12461, N12455, N9292);
xor XOR2 (N12462, N12447, N10467);
and AND2 (N12463, N12403, N3232);
nor NOR2 (N12464, N12462, N1889);
or OR3 (N12465, N12464, N1548, N11122);
or OR3 (N12466, N12449, N2614, N9077);
and AND2 (N12467, N12461, N9284);
not NOT1 (N12468, N12466);
and AND3 (N12469, N12463, N8498, N2829);
buf BUF1 (N12470, N12453);
nand NAND3 (N12471, N12460, N4055, N11551);
xor XOR2 (N12472, N12444, N483);
buf BUF1 (N12473, N12456);
and AND4 (N12474, N12420, N9847, N7164, N9510);
and AND3 (N12475, N12465, N7113, N3939);
nor NOR3 (N12476, N12472, N5769, N9121);
xor XOR2 (N12477, N12469, N8648);
xor XOR2 (N12478, N12470, N6519);
not NOT1 (N12479, N12459);
not NOT1 (N12480, N12473);
nand NAND2 (N12481, N12468, N789);
nor NOR4 (N12482, N12477, N10298, N1518, N10895);
and AND4 (N12483, N12475, N981, N1927, N10247);
nor NOR3 (N12484, N12481, N9297, N7531);
or OR2 (N12485, N12476, N3989);
nor NOR4 (N12486, N12474, N1224, N4365, N8231);
nor NOR2 (N12487, N12482, N8036);
nor NOR2 (N12488, N12486, N9915);
buf BUF1 (N12489, N12485);
nand NAND2 (N12490, N12471, N9800);
and AND2 (N12491, N12489, N5413);
and AND2 (N12492, N12484, N2387);
or OR3 (N12493, N12490, N880, N194);
and AND2 (N12494, N12479, N7160);
xor XOR2 (N12495, N12480, N10382);
and AND4 (N12496, N12494, N6615, N8523, N10827);
and AND2 (N12497, N12478, N6535);
buf BUF1 (N12498, N12492);
nor NOR2 (N12499, N12495, N4019);
nor NOR4 (N12500, N12496, N2984, N10275, N8714);
nor NOR4 (N12501, N12499, N517, N11711, N9946);
or OR2 (N12502, N12500, N9464);
nor NOR3 (N12503, N12491, N4821, N11884);
not NOT1 (N12504, N12502);
not NOT1 (N12505, N12497);
and AND4 (N12506, N12498, N1659, N9294, N2138);
xor XOR2 (N12507, N12488, N5110);
not NOT1 (N12508, N12483);
buf BUF1 (N12509, N12503);
not NOT1 (N12510, N12509);
or OR3 (N12511, N12504, N1929, N4763);
not NOT1 (N12512, N12505);
or OR4 (N12513, N12501, N7324, N6337, N9583);
nor NOR4 (N12514, N12511, N1737, N5934, N9067);
not NOT1 (N12515, N12508);
and AND2 (N12516, N12514, N37);
nand NAND4 (N12517, N12493, N9162, N8052, N4043);
buf BUF1 (N12518, N12515);
nor NOR3 (N12519, N12487, N1510, N1324);
or OR4 (N12520, N12517, N3085, N2779, N3939);
xor XOR2 (N12521, N12467, N6113);
nor NOR2 (N12522, N12507, N1675);
xor XOR2 (N12523, N12513, N1649);
nand NAND3 (N12524, N12512, N466, N4391);
not NOT1 (N12525, N12524);
buf BUF1 (N12526, N12506);
xor XOR2 (N12527, N12516, N4661);
not NOT1 (N12528, N12526);
xor XOR2 (N12529, N12519, N1873);
and AND3 (N12530, N12529, N10774, N7567);
nand NAND2 (N12531, N12510, N7538);
not NOT1 (N12532, N12518);
not NOT1 (N12533, N12525);
xor XOR2 (N12534, N12522, N9232);
xor XOR2 (N12535, N12531, N6333);
buf BUF1 (N12536, N12528);
and AND3 (N12537, N12535, N7944, N7557);
or OR3 (N12538, N12533, N5095, N10102);
xor XOR2 (N12539, N12536, N1379);
and AND3 (N12540, N12537, N11415, N8121);
xor XOR2 (N12541, N12521, N7180);
nor NOR2 (N12542, N12532, N8198);
or OR2 (N12543, N12534, N6065);
or OR2 (N12544, N12543, N11144);
xor XOR2 (N12545, N12527, N6923);
xor XOR2 (N12546, N12544, N5673);
or OR4 (N12547, N12540, N10299, N3212, N6213);
buf BUF1 (N12548, N12541);
buf BUF1 (N12549, N12530);
buf BUF1 (N12550, N12539);
and AND2 (N12551, N12520, N537);
xor XOR2 (N12552, N12551, N3486);
nand NAND4 (N12553, N12550, N11812, N12432, N12289);
or OR3 (N12554, N12547, N12289, N12489);
xor XOR2 (N12555, N12545, N981);
xor XOR2 (N12556, N12546, N4201);
nor NOR3 (N12557, N12556, N5731, N12121);
buf BUF1 (N12558, N12548);
buf BUF1 (N12559, N12549);
nand NAND4 (N12560, N12559, N215, N7320, N6491);
nand NAND3 (N12561, N12553, N6557, N2033);
not NOT1 (N12562, N12523);
and AND4 (N12563, N12558, N11306, N7792, N6631);
not NOT1 (N12564, N12563);
and AND3 (N12565, N12552, N7672, N2534);
xor XOR2 (N12566, N12538, N5355);
nor NOR4 (N12567, N12565, N3329, N8763, N11552);
not NOT1 (N12568, N12561);
and AND2 (N12569, N12557, N4728);
xor XOR2 (N12570, N12566, N3730);
and AND3 (N12571, N12570, N1503, N3302);
or OR4 (N12572, N12555, N5026, N3376, N9887);
and AND3 (N12573, N12569, N10804, N3428);
xor XOR2 (N12574, N12568, N9617);
and AND2 (N12575, N12572, N6179);
nand NAND3 (N12576, N12567, N3577, N2607);
nand NAND3 (N12577, N12575, N724, N10594);
xor XOR2 (N12578, N12577, N5230);
nor NOR4 (N12579, N12562, N3893, N1030, N6333);
buf BUF1 (N12580, N12573);
nand NAND2 (N12581, N12554, N11467);
nand NAND4 (N12582, N12581, N1094, N2157, N4433);
not NOT1 (N12583, N12564);
not NOT1 (N12584, N12583);
and AND3 (N12585, N12571, N3588, N10844);
buf BUF1 (N12586, N12578);
nor NOR4 (N12587, N12584, N2312, N9626, N10586);
not NOT1 (N12588, N12542);
or OR2 (N12589, N12560, N11541);
nand NAND3 (N12590, N12574, N11802, N2992);
or OR2 (N12591, N12579, N10889);
and AND3 (N12592, N12591, N9815, N8402);
xor XOR2 (N12593, N12586, N12096);
nand NAND2 (N12594, N12593, N11588);
or OR3 (N12595, N12585, N2305, N632);
nor NOR2 (N12596, N12582, N8863);
nor NOR2 (N12597, N12590, N9705);
nor NOR3 (N12598, N12592, N455, N12325);
nor NOR4 (N12599, N12576, N3717, N6265, N9216);
xor XOR2 (N12600, N12580, N11421);
not NOT1 (N12601, N12596);
nand NAND4 (N12602, N12594, N3413, N1889, N10436);
or OR2 (N12603, N12588, N4220);
buf BUF1 (N12604, N12595);
or OR3 (N12605, N12587, N3352, N4335);
xor XOR2 (N12606, N12589, N11790);
buf BUF1 (N12607, N12598);
nand NAND3 (N12608, N12600, N974, N3396);
and AND2 (N12609, N12607, N10008);
not NOT1 (N12610, N12599);
not NOT1 (N12611, N12608);
or OR3 (N12612, N12604, N4431, N4974);
buf BUF1 (N12613, N12601);
and AND4 (N12614, N12605, N10654, N3733, N3877);
nand NAND4 (N12615, N12611, N5080, N1299, N8868);
nor NOR2 (N12616, N12614, N8568);
or OR2 (N12617, N12603, N891);
or OR2 (N12618, N12613, N2966);
buf BUF1 (N12619, N12618);
xor XOR2 (N12620, N12616, N3937);
xor XOR2 (N12621, N12612, N10990);
nor NOR4 (N12622, N12606, N9011, N5034, N5178);
xor XOR2 (N12623, N12597, N11422);
not NOT1 (N12624, N12602);
not NOT1 (N12625, N12620);
buf BUF1 (N12626, N12623);
not NOT1 (N12627, N12617);
nor NOR3 (N12628, N12627, N12167, N6917);
nor NOR2 (N12629, N12625, N379);
xor XOR2 (N12630, N12626, N2680);
nor NOR4 (N12631, N12630, N7343, N12565, N6392);
not NOT1 (N12632, N12622);
and AND4 (N12633, N12631, N10821, N9860, N4088);
or OR4 (N12634, N12610, N9037, N10310, N4014);
not NOT1 (N12635, N12624);
nor NOR4 (N12636, N12609, N2008, N8175, N9086);
buf BUF1 (N12637, N12633);
not NOT1 (N12638, N12634);
or OR2 (N12639, N12628, N7622);
xor XOR2 (N12640, N12632, N10648);
buf BUF1 (N12641, N12640);
nand NAND4 (N12642, N12635, N5974, N2356, N639);
not NOT1 (N12643, N12615);
nor NOR4 (N12644, N12639, N12374, N8911, N4896);
xor XOR2 (N12645, N12643, N11129);
not NOT1 (N12646, N12619);
buf BUF1 (N12647, N12621);
nor NOR2 (N12648, N12646, N3948);
buf BUF1 (N12649, N12648);
and AND2 (N12650, N12638, N11292);
buf BUF1 (N12651, N12647);
not NOT1 (N12652, N12629);
or OR2 (N12653, N12651, N3384);
or OR4 (N12654, N12644, N6927, N11263, N1948);
not NOT1 (N12655, N12645);
or OR3 (N12656, N12652, N3588, N6332);
nand NAND4 (N12657, N12650, N2375, N10500, N5839);
nand NAND4 (N12658, N12654, N498, N6266, N11113);
and AND2 (N12659, N12653, N8217);
buf BUF1 (N12660, N12656);
not NOT1 (N12661, N12636);
nor NOR2 (N12662, N12649, N12456);
and AND4 (N12663, N12658, N8326, N1764, N646);
buf BUF1 (N12664, N12659);
nand NAND2 (N12665, N12657, N11706);
xor XOR2 (N12666, N12641, N10577);
buf BUF1 (N12667, N12663);
nand NAND4 (N12668, N12660, N9911, N1668, N2562);
nand NAND3 (N12669, N12668, N4271, N11307);
xor XOR2 (N12670, N12664, N10819);
nor NOR4 (N12671, N12655, N9615, N2178, N1414);
nor NOR4 (N12672, N12637, N4044, N3362, N5661);
buf BUF1 (N12673, N12667);
nor NOR4 (N12674, N12673, N5349, N7261, N7019);
nand NAND3 (N12675, N12671, N3051, N12191);
nor NOR2 (N12676, N12670, N3875);
or OR4 (N12677, N12674, N8533, N12213, N6493);
buf BUF1 (N12678, N12642);
or OR3 (N12679, N12676, N3658, N8595);
nor NOR3 (N12680, N12679, N7238, N4678);
and AND3 (N12681, N12665, N7473, N468);
or OR2 (N12682, N12677, N10802);
nand NAND4 (N12683, N12680, N11643, N4678, N5837);
nand NAND4 (N12684, N12675, N11060, N5867, N11668);
buf BUF1 (N12685, N12662);
or OR4 (N12686, N12669, N10939, N11075, N11532);
xor XOR2 (N12687, N12683, N8690);
nor NOR4 (N12688, N12681, N2699, N7594, N3861);
buf BUF1 (N12689, N12682);
nor NOR2 (N12690, N12689, N6108);
nand NAND3 (N12691, N12686, N8885, N3198);
buf BUF1 (N12692, N12672);
nor NOR4 (N12693, N12678, N7848, N3220, N6635);
nor NOR4 (N12694, N12661, N1477, N2134, N1302);
nand NAND4 (N12695, N12694, N5013, N9960, N11384);
not NOT1 (N12696, N12688);
nand NAND4 (N12697, N12687, N12348, N30, N5969);
nor NOR3 (N12698, N12684, N10176, N12509);
xor XOR2 (N12699, N12685, N8044);
nor NOR4 (N12700, N12692, N3552, N10306, N5612);
nor NOR3 (N12701, N12693, N6127, N1928);
or OR2 (N12702, N12700, N7338);
or OR2 (N12703, N12691, N4155);
not NOT1 (N12704, N12690);
not NOT1 (N12705, N12703);
buf BUF1 (N12706, N12702);
and AND3 (N12707, N12698, N1482, N5030);
nor NOR4 (N12708, N12701, N4162, N7006, N12659);
or OR2 (N12709, N12706, N4479);
not NOT1 (N12710, N12699);
buf BUF1 (N12711, N12697);
and AND4 (N12712, N12705, N9737, N1350, N2513);
xor XOR2 (N12713, N12708, N11952);
nand NAND4 (N12714, N12707, N3187, N3172, N5728);
nor NOR4 (N12715, N12710, N1072, N9028, N8618);
nand NAND2 (N12716, N12695, N6236);
nor NOR4 (N12717, N12714, N740, N5471, N9133);
xor XOR2 (N12718, N12716, N4221);
xor XOR2 (N12719, N12713, N3849);
or OR2 (N12720, N12719, N5334);
and AND2 (N12721, N12717, N3730);
nand NAND2 (N12722, N12666, N11220);
nor NOR3 (N12723, N12704, N2700, N8512);
and AND4 (N12724, N12712, N76, N9093, N8433);
or OR3 (N12725, N12709, N8197, N5523);
or OR2 (N12726, N12725, N7502);
xor XOR2 (N12727, N12723, N2583);
buf BUF1 (N12728, N12724);
or OR4 (N12729, N12720, N4261, N12278, N5571);
nand NAND4 (N12730, N12726, N1838, N8463, N4832);
not NOT1 (N12731, N12696);
not NOT1 (N12732, N12721);
nor NOR2 (N12733, N12711, N10766);
buf BUF1 (N12734, N12729);
and AND4 (N12735, N12732, N12488, N2319, N4017);
nor NOR3 (N12736, N12718, N10419, N197);
nand NAND2 (N12737, N12734, N8375);
buf BUF1 (N12738, N12728);
nand NAND3 (N12739, N12736, N11620, N10003);
not NOT1 (N12740, N12730);
nand NAND2 (N12741, N12715, N3824);
or OR4 (N12742, N12727, N8326, N12527, N5498);
nand NAND3 (N12743, N12731, N7387, N4080);
buf BUF1 (N12744, N12741);
or OR2 (N12745, N12722, N10741);
nor NOR4 (N12746, N12743, N2281, N12006, N7985);
nor NOR3 (N12747, N12744, N3303, N11383);
nand NAND4 (N12748, N12740, N10966, N10248, N5169);
nand NAND3 (N12749, N12737, N10639, N6728);
and AND3 (N12750, N12747, N7432, N11523);
not NOT1 (N12751, N12739);
nand NAND2 (N12752, N12738, N4075);
xor XOR2 (N12753, N12746, N9763);
nand NAND3 (N12754, N12742, N5504, N1026);
or OR4 (N12755, N12752, N7438, N8175, N8527);
not NOT1 (N12756, N12735);
nor NOR4 (N12757, N12733, N9788, N298, N1231);
xor XOR2 (N12758, N12753, N481);
not NOT1 (N12759, N12754);
nand NAND4 (N12760, N12758, N1054, N7880, N5961);
not NOT1 (N12761, N12755);
and AND3 (N12762, N12750, N4161, N20);
buf BUF1 (N12763, N12762);
xor XOR2 (N12764, N12761, N10929);
nand NAND3 (N12765, N12751, N7720, N6311);
or OR3 (N12766, N12760, N11985, N10049);
nand NAND4 (N12767, N12764, N3277, N5503, N10560);
and AND3 (N12768, N12766, N1395, N11078);
and AND2 (N12769, N12745, N2242);
nor NOR3 (N12770, N12756, N10349, N9512);
not NOT1 (N12771, N12748);
and AND3 (N12772, N12749, N8122, N1066);
nand NAND3 (N12773, N12768, N11814, N12274);
and AND3 (N12774, N12767, N7040, N2619);
nor NOR4 (N12775, N12772, N1858, N3827, N5504);
nor NOR3 (N12776, N12765, N489, N1076);
nand NAND4 (N12777, N12769, N5154, N7274, N4906);
xor XOR2 (N12778, N12776, N6099);
nor NOR2 (N12779, N12763, N3673);
nand NAND2 (N12780, N12770, N5451);
nand NAND3 (N12781, N12773, N11835, N10655);
and AND2 (N12782, N12759, N11470);
or OR2 (N12783, N12771, N8062);
or OR2 (N12784, N12782, N1307);
or OR4 (N12785, N12781, N7297, N3125, N8984);
buf BUF1 (N12786, N12775);
not NOT1 (N12787, N12783);
nor NOR2 (N12788, N12787, N3280);
nand NAND2 (N12789, N12780, N1647);
buf BUF1 (N12790, N12789);
buf BUF1 (N12791, N12774);
nor NOR3 (N12792, N12790, N11174, N6232);
nand NAND2 (N12793, N12791, N1389);
nor NOR2 (N12794, N12757, N7069);
nand NAND4 (N12795, N12785, N8534, N10459, N4588);
not NOT1 (N12796, N12788);
buf BUF1 (N12797, N12793);
buf BUF1 (N12798, N12794);
buf BUF1 (N12799, N12798);
and AND4 (N12800, N12779, N1317, N1435, N6249);
not NOT1 (N12801, N12786);
and AND3 (N12802, N12799, N1124, N10198);
xor XOR2 (N12803, N12800, N11997);
buf BUF1 (N12804, N12797);
nor NOR4 (N12805, N12792, N2983, N7303, N8287);
not NOT1 (N12806, N12796);
nor NOR3 (N12807, N12795, N2277, N11671);
or OR2 (N12808, N12802, N2080);
not NOT1 (N12809, N12784);
buf BUF1 (N12810, N12807);
nor NOR2 (N12811, N12803, N1166);
not NOT1 (N12812, N12777);
not NOT1 (N12813, N12809);
nor NOR4 (N12814, N12811, N8740, N11482, N6568);
nand NAND2 (N12815, N12813, N10163);
or OR2 (N12816, N12815, N1637);
and AND2 (N12817, N12806, N3682);
and AND4 (N12818, N12810, N11703, N11618, N9701);
and AND3 (N12819, N12805, N2448, N10898);
not NOT1 (N12820, N12814);
buf BUF1 (N12821, N12804);
xor XOR2 (N12822, N12820, N2859);
nand NAND2 (N12823, N12812, N8449);
not NOT1 (N12824, N12816);
nor NOR4 (N12825, N12778, N249, N7533, N7629);
nor NOR3 (N12826, N12824, N12124, N1060);
buf BUF1 (N12827, N12822);
not NOT1 (N12828, N12819);
nand NAND4 (N12829, N12827, N3692, N12453, N6175);
and AND4 (N12830, N12825, N5625, N5838, N10350);
nor NOR2 (N12831, N12801, N3659);
nor NOR3 (N12832, N12821, N2295, N12724);
nor NOR2 (N12833, N12830, N9086);
nor NOR2 (N12834, N12833, N11237);
or OR2 (N12835, N12834, N6412);
and AND2 (N12836, N12831, N11775);
xor XOR2 (N12837, N12808, N6317);
xor XOR2 (N12838, N12837, N4958);
and AND3 (N12839, N12828, N4573, N5579);
nor NOR4 (N12840, N12832, N358, N6097, N9307);
or OR3 (N12841, N12823, N4538, N309);
nor NOR2 (N12842, N12838, N9045);
nor NOR2 (N12843, N12829, N6875);
nand NAND2 (N12844, N12826, N3491);
not NOT1 (N12845, N12818);
nor NOR3 (N12846, N12843, N3142, N12473);
nand NAND4 (N12847, N12835, N12050, N4447, N3998);
nand NAND3 (N12848, N12845, N11857, N6);
and AND4 (N12849, N12841, N10480, N4975, N11902);
buf BUF1 (N12850, N12840);
or OR3 (N12851, N12846, N1635, N2023);
nand NAND3 (N12852, N12849, N9657, N9944);
xor XOR2 (N12853, N12850, N6733);
not NOT1 (N12854, N12842);
buf BUF1 (N12855, N12851);
and AND4 (N12856, N12844, N5832, N11474, N12400);
not NOT1 (N12857, N12836);
or OR2 (N12858, N12853, N11923);
nor NOR2 (N12859, N12855, N76);
nor NOR3 (N12860, N12847, N1743, N2101);
and AND2 (N12861, N12854, N817);
not NOT1 (N12862, N12817);
buf BUF1 (N12863, N12839);
not NOT1 (N12864, N12857);
buf BUF1 (N12865, N12862);
not NOT1 (N12866, N12861);
or OR2 (N12867, N12848, N7858);
xor XOR2 (N12868, N12863, N12235);
or OR3 (N12869, N12864, N1500, N9020);
not NOT1 (N12870, N12852);
nand NAND2 (N12871, N12870, N8512);
buf BUF1 (N12872, N12869);
nand NAND3 (N12873, N12871, N12716, N1138);
and AND3 (N12874, N12873, N1278, N8432);
nand NAND2 (N12875, N12859, N7488);
nor NOR4 (N12876, N12866, N3331, N4457, N1650);
and AND4 (N12877, N12868, N8083, N2348, N609);
nor NOR3 (N12878, N12875, N6264, N10303);
and AND2 (N12879, N12865, N6955);
or OR3 (N12880, N12878, N1477, N7209);
xor XOR2 (N12881, N12856, N8940);
or OR4 (N12882, N12880, N4463, N8713, N7197);
xor XOR2 (N12883, N12858, N8960);
buf BUF1 (N12884, N12876);
nor NOR3 (N12885, N12883, N4232, N2394);
or OR4 (N12886, N12877, N2225, N8248, N10669);
xor XOR2 (N12887, N12884, N12760);
or OR2 (N12888, N12887, N3549);
nor NOR3 (N12889, N12888, N4113, N5794);
and AND3 (N12890, N12885, N9954, N8843);
nor NOR4 (N12891, N12886, N11957, N8765, N1712);
nor NOR2 (N12892, N12872, N7335);
nand NAND3 (N12893, N12889, N202, N7402);
nor NOR4 (N12894, N12882, N9984, N862, N5071);
and AND2 (N12895, N12893, N2737);
buf BUF1 (N12896, N12895);
xor XOR2 (N12897, N12892, N12189);
and AND2 (N12898, N12874, N919);
or OR3 (N12899, N12896, N6917, N2878);
and AND4 (N12900, N12860, N12382, N468, N5624);
nand NAND3 (N12901, N12891, N12719, N3722);
nand NAND4 (N12902, N12894, N7045, N8389, N10223);
not NOT1 (N12903, N12879);
not NOT1 (N12904, N12901);
buf BUF1 (N12905, N12867);
and AND4 (N12906, N12905, N3434, N699, N2551);
xor XOR2 (N12907, N12881, N5386);
or OR4 (N12908, N12906, N8888, N11332, N7986);
nand NAND4 (N12909, N12903, N6689, N130, N10049);
and AND4 (N12910, N12909, N5230, N8566, N3567);
nor NOR4 (N12911, N12902, N10844, N6781, N2132);
nand NAND2 (N12912, N12900, N2788);
nand NAND3 (N12913, N12890, N4901, N3403);
xor XOR2 (N12914, N12897, N2616);
or OR3 (N12915, N12898, N2440, N11915);
buf BUF1 (N12916, N12908);
and AND4 (N12917, N12913, N7149, N5439, N12801);
nand NAND3 (N12918, N12904, N8625, N12699);
and AND3 (N12919, N12916, N10295, N12870);
nor NOR2 (N12920, N12914, N11615);
and AND2 (N12921, N12910, N39);
nand NAND4 (N12922, N12918, N3001, N11398, N9666);
and AND4 (N12923, N12915, N11461, N1930, N1843);
or OR3 (N12924, N12911, N11615, N12808);
or OR2 (N12925, N12917, N10549);
nand NAND3 (N12926, N12919, N5376, N10350);
and AND2 (N12927, N12923, N7774);
buf BUF1 (N12928, N12926);
xor XOR2 (N12929, N12922, N6809);
xor XOR2 (N12930, N12907, N8301);
nor NOR2 (N12931, N12928, N7746);
buf BUF1 (N12932, N12899);
nand NAND3 (N12933, N12925, N6945, N7824);
and AND3 (N12934, N12931, N10942, N5790);
xor XOR2 (N12935, N12927, N11813);
or OR3 (N12936, N12933, N1277, N7243);
not NOT1 (N12937, N12932);
or OR3 (N12938, N12934, N9199, N787);
and AND4 (N12939, N12937, N2172, N4652, N7081);
buf BUF1 (N12940, N12921);
not NOT1 (N12941, N12924);
not NOT1 (N12942, N12940);
nor NOR3 (N12943, N12939, N881, N3630);
nand NAND4 (N12944, N12942, N11046, N4069, N2014);
not NOT1 (N12945, N12941);
buf BUF1 (N12946, N12935);
buf BUF1 (N12947, N12946);
nor NOR2 (N12948, N12930, N8825);
and AND2 (N12949, N12912, N9460);
buf BUF1 (N12950, N12929);
not NOT1 (N12951, N12938);
or OR3 (N12952, N12936, N6945, N2486);
nand NAND3 (N12953, N12943, N12915, N11033);
nor NOR2 (N12954, N12948, N4105);
or OR3 (N12955, N12944, N6198, N2235);
buf BUF1 (N12956, N12950);
and AND3 (N12957, N12947, N7673, N4889);
buf BUF1 (N12958, N12957);
nand NAND4 (N12959, N12949, N12431, N6399, N9339);
not NOT1 (N12960, N12959);
xor XOR2 (N12961, N12954, N7168);
nand NAND3 (N12962, N12952, N3691, N9653);
xor XOR2 (N12963, N12945, N9309);
not NOT1 (N12964, N12953);
nand NAND3 (N12965, N12960, N6275, N4851);
nor NOR4 (N12966, N12965, N1263, N6447, N9170);
not NOT1 (N12967, N12951);
and AND4 (N12968, N12963, N3671, N10417, N9723);
not NOT1 (N12969, N12958);
buf BUF1 (N12970, N12962);
or OR2 (N12971, N12967, N3985);
and AND2 (N12972, N12964, N11501);
or OR2 (N12973, N12972, N4474);
buf BUF1 (N12974, N12956);
and AND4 (N12975, N12961, N1655, N4021, N4087);
and AND2 (N12976, N12975, N5509);
nor NOR4 (N12977, N12974, N8218, N4306, N516);
nor NOR2 (N12978, N12970, N11565);
buf BUF1 (N12979, N12920);
buf BUF1 (N12980, N12969);
or OR3 (N12981, N12977, N6157, N156);
not NOT1 (N12982, N12978);
xor XOR2 (N12983, N12980, N8112);
not NOT1 (N12984, N12971);
buf BUF1 (N12985, N12973);
buf BUF1 (N12986, N12976);
nand NAND4 (N12987, N12966, N6481, N5332, N9099);
or OR4 (N12988, N12985, N1489, N11439, N5624);
nand NAND4 (N12989, N12983, N11513, N11529, N4147);
nand NAND3 (N12990, N12986, N7028, N4706);
nand NAND4 (N12991, N12981, N5774, N1358, N2653);
buf BUF1 (N12992, N12990);
nor NOR4 (N12993, N12982, N2139, N4149, N6640);
not NOT1 (N12994, N12968);
nand NAND3 (N12995, N12979, N1905, N2531);
not NOT1 (N12996, N12987);
nor NOR2 (N12997, N12991, N7561);
buf BUF1 (N12998, N12955);
not NOT1 (N12999, N12997);
buf BUF1 (N13000, N12998);
nor NOR2 (N13001, N12988, N5507);
and AND2 (N13002, N12994, N4403);
xor XOR2 (N13003, N13002, N12045);
buf BUF1 (N13004, N13001);
or OR4 (N13005, N12992, N12456, N11712, N9947);
nand NAND4 (N13006, N13003, N9268, N4479, N7847);
buf BUF1 (N13007, N13004);
nor NOR2 (N13008, N12996, N1067);
buf BUF1 (N13009, N12993);
buf BUF1 (N13010, N13009);
not NOT1 (N13011, N12984);
not NOT1 (N13012, N12999);
and AND2 (N13013, N13012, N7759);
nor NOR3 (N13014, N12989, N80, N5723);
and AND2 (N13015, N12995, N7323);
and AND4 (N13016, N13014, N6064, N4781, N9084);
buf BUF1 (N13017, N13007);
xor XOR2 (N13018, N13006, N42);
not NOT1 (N13019, N13018);
nor NOR2 (N13020, N13008, N7962);
nand NAND4 (N13021, N13017, N9576, N5513, N4788);
not NOT1 (N13022, N13013);
or OR2 (N13023, N13019, N9295);
nor NOR3 (N13024, N13020, N11358, N12297);
xor XOR2 (N13025, N13023, N1614);
nor NOR4 (N13026, N13025, N2667, N11818, N346);
or OR3 (N13027, N13011, N6085, N9740);
buf BUF1 (N13028, N13026);
nor NOR4 (N13029, N13028, N3834, N1942, N12088);
nand NAND4 (N13030, N13016, N7036, N8765, N3978);
nor NOR4 (N13031, N13027, N3555, N6082, N1693);
buf BUF1 (N13032, N13010);
xor XOR2 (N13033, N13024, N10193);
or OR2 (N13034, N13021, N5073);
and AND4 (N13035, N13022, N6046, N1084, N3581);
not NOT1 (N13036, N13034);
nor NOR3 (N13037, N13035, N12133, N10130);
not NOT1 (N13038, N13005);
buf BUF1 (N13039, N13000);
xor XOR2 (N13040, N13038, N3848);
not NOT1 (N13041, N13030);
and AND4 (N13042, N13039, N3408, N12856, N11256);
xor XOR2 (N13043, N13031, N10515);
buf BUF1 (N13044, N13029);
nand NAND4 (N13045, N13037, N8148, N4040, N192);
xor XOR2 (N13046, N13045, N645);
not NOT1 (N13047, N13044);
nor NOR3 (N13048, N13032, N2244, N1566);
and AND3 (N13049, N13040, N10512, N9201);
nand NAND3 (N13050, N13015, N5574, N8435);
and AND4 (N13051, N13033, N3135, N10866, N8680);
not NOT1 (N13052, N13041);
xor XOR2 (N13053, N13050, N9685);
or OR4 (N13054, N13052, N4135, N11235, N12041);
buf BUF1 (N13055, N13048);
buf BUF1 (N13056, N13042);
not NOT1 (N13057, N13055);
xor XOR2 (N13058, N13056, N4194);
nand NAND4 (N13059, N13053, N4820, N241, N5223);
buf BUF1 (N13060, N13058);
nor NOR3 (N13061, N13047, N11041, N180);
and AND4 (N13062, N13046, N2317, N4781, N11770);
nand NAND4 (N13063, N13054, N1827, N5518, N12544);
nor NOR2 (N13064, N13062, N9697);
not NOT1 (N13065, N13063);
buf BUF1 (N13066, N13051);
nor NOR2 (N13067, N13066, N6587);
and AND2 (N13068, N13064, N10729);
not NOT1 (N13069, N13049);
and AND2 (N13070, N13060, N4351);
nand NAND4 (N13071, N13067, N3655, N7662, N2698);
buf BUF1 (N13072, N13070);
xor XOR2 (N13073, N13059, N11026);
nor NOR4 (N13074, N13043, N7713, N5040, N12451);
and AND3 (N13075, N13074, N3833, N2049);
nand NAND4 (N13076, N13073, N356, N2335, N10713);
nor NOR4 (N13077, N13036, N338, N10936, N3623);
not NOT1 (N13078, N13076);
nand NAND3 (N13079, N13071, N37, N6091);
not NOT1 (N13080, N13077);
nand NAND2 (N13081, N13075, N1444);
and AND3 (N13082, N13057, N7330, N1079);
nand NAND4 (N13083, N13065, N12306, N8976, N8762);
buf BUF1 (N13084, N13082);
and AND3 (N13085, N13068, N2099, N1700);
buf BUF1 (N13086, N13079);
buf BUF1 (N13087, N13085);
not NOT1 (N13088, N13080);
nand NAND3 (N13089, N13086, N2165, N4698);
nor NOR3 (N13090, N13089, N9890, N4001);
not NOT1 (N13091, N13069);
not NOT1 (N13092, N13061);
nand NAND4 (N13093, N13088, N6329, N8419, N12496);
nor NOR4 (N13094, N13084, N11160, N2535, N6811);
buf BUF1 (N13095, N13081);
nor NOR4 (N13096, N13095, N7160, N11601, N7123);
nand NAND3 (N13097, N13072, N5257, N5891);
or OR3 (N13098, N13092, N4168, N10936);
not NOT1 (N13099, N13083);
nor NOR2 (N13100, N13093, N2772);
buf BUF1 (N13101, N13078);
buf BUF1 (N13102, N13096);
buf BUF1 (N13103, N13097);
and AND4 (N13104, N13103, N10889, N11830, N3524);
buf BUF1 (N13105, N13101);
not NOT1 (N13106, N13099);
nand NAND3 (N13107, N13090, N3295, N535);
buf BUF1 (N13108, N13106);
or OR4 (N13109, N13087, N11543, N4214, N8743);
not NOT1 (N13110, N13098);
buf BUF1 (N13111, N13091);
and AND4 (N13112, N13109, N11162, N5173, N19);
nor NOR3 (N13113, N13100, N10639, N12004);
nor NOR4 (N13114, N13111, N10916, N7002, N12616);
xor XOR2 (N13115, N13107, N7316);
nor NOR4 (N13116, N13115, N8222, N1911, N8796);
buf BUF1 (N13117, N13094);
nor NOR2 (N13118, N13108, N10269);
or OR3 (N13119, N13117, N3742, N6755);
buf BUF1 (N13120, N13105);
nor NOR4 (N13121, N13110, N3539, N6928, N7867);
nand NAND3 (N13122, N13114, N9780, N2604);
or OR4 (N13123, N13112, N5382, N6660, N1570);
and AND3 (N13124, N13121, N5141, N9159);
not NOT1 (N13125, N13104);
buf BUF1 (N13126, N13118);
not NOT1 (N13127, N13102);
xor XOR2 (N13128, N13127, N8445);
nand NAND4 (N13129, N13126, N8043, N1283, N10997);
nor NOR4 (N13130, N13113, N5478, N7838, N10914);
not NOT1 (N13131, N13123);
and AND2 (N13132, N13131, N9680);
xor XOR2 (N13133, N13124, N10848);
nor NOR3 (N13134, N13129, N8264, N7856);
not NOT1 (N13135, N13116);
and AND4 (N13136, N13135, N1479, N10887, N6261);
nand NAND2 (N13137, N13128, N7594);
nor NOR4 (N13138, N13137, N11938, N7523, N2266);
buf BUF1 (N13139, N13125);
xor XOR2 (N13140, N13132, N6951);
buf BUF1 (N13141, N13133);
buf BUF1 (N13142, N13136);
nor NOR2 (N13143, N13120, N5543);
nand NAND4 (N13144, N13142, N3209, N7149, N1310);
buf BUF1 (N13145, N13140);
not NOT1 (N13146, N13139);
nor NOR3 (N13147, N13146, N2153, N2974);
buf BUF1 (N13148, N13145);
and AND3 (N13149, N13144, N13058, N4142);
buf BUF1 (N13150, N13130);
nor NOR4 (N13151, N13147, N5915, N3749, N12080);
or OR3 (N13152, N13141, N13016, N11260);
or OR4 (N13153, N13119, N1027, N7093, N3502);
not NOT1 (N13154, N13153);
buf BUF1 (N13155, N13134);
not NOT1 (N13156, N13143);
buf BUF1 (N13157, N13149);
not NOT1 (N13158, N13150);
not NOT1 (N13159, N13155);
not NOT1 (N13160, N13152);
xor XOR2 (N13161, N13122, N11171);
xor XOR2 (N13162, N13156, N2893);
nand NAND2 (N13163, N13148, N1973);
xor XOR2 (N13164, N13151, N5743);
buf BUF1 (N13165, N13161);
and AND2 (N13166, N13157, N2322);
and AND3 (N13167, N13166, N11054, N5661);
not NOT1 (N13168, N13154);
and AND2 (N13169, N13167, N91);
buf BUF1 (N13170, N13165);
xor XOR2 (N13171, N13159, N3614);
or OR3 (N13172, N13162, N4216, N11468);
buf BUF1 (N13173, N13170);
or OR4 (N13174, N13163, N7752, N3611, N5244);
and AND2 (N13175, N13172, N3693);
or OR4 (N13176, N13169, N8714, N8022, N8491);
and AND3 (N13177, N13164, N8855, N1436);
and AND4 (N13178, N13176, N6923, N10125, N6006);
and AND4 (N13179, N13175, N4788, N4615, N184);
and AND3 (N13180, N13168, N5741, N12449);
nand NAND2 (N13181, N13177, N2077);
nor NOR3 (N13182, N13138, N387, N2749);
buf BUF1 (N13183, N13158);
or OR2 (N13184, N13181, N11597);
buf BUF1 (N13185, N13178);
nand NAND4 (N13186, N13185, N5550, N1199, N2079);
buf BUF1 (N13187, N13180);
and AND3 (N13188, N13186, N4603, N1503);
xor XOR2 (N13189, N13171, N1283);
nand NAND2 (N13190, N13187, N12506);
nor NOR3 (N13191, N13190, N705, N4846);
and AND4 (N13192, N13179, N7711, N131, N4124);
or OR2 (N13193, N13173, N1993);
not NOT1 (N13194, N13191);
nand NAND3 (N13195, N13189, N5729, N12941);
nand NAND4 (N13196, N13188, N5456, N8926, N11952);
nand NAND2 (N13197, N13160, N4532);
buf BUF1 (N13198, N13195);
buf BUF1 (N13199, N13194);
nor NOR3 (N13200, N13198, N478, N7275);
and AND3 (N13201, N13174, N617, N4993);
and AND4 (N13202, N13183, N2224, N1194, N1503);
xor XOR2 (N13203, N13197, N8999);
buf BUF1 (N13204, N13196);
and AND2 (N13205, N13200, N2483);
xor XOR2 (N13206, N13203, N7504);
and AND2 (N13207, N13182, N7661);
nand NAND2 (N13208, N13201, N11866);
or OR2 (N13209, N13184, N4634);
nand NAND2 (N13210, N13209, N13016);
or OR4 (N13211, N13204, N4582, N4213, N5604);
xor XOR2 (N13212, N13206, N2636);
or OR4 (N13213, N13211, N4565, N12590, N2871);
nor NOR2 (N13214, N13210, N6413);
not NOT1 (N13215, N13207);
nor NOR3 (N13216, N13199, N12343, N13054);
nand NAND2 (N13217, N13208, N3706);
or OR3 (N13218, N13202, N7439, N6071);
or OR4 (N13219, N13215, N6567, N12870, N5080);
nor NOR3 (N13220, N13192, N12490, N9226);
buf BUF1 (N13221, N13212);
buf BUF1 (N13222, N13221);
not NOT1 (N13223, N13214);
nand NAND4 (N13224, N13218, N4102, N7059, N2009);
buf BUF1 (N13225, N13205);
and AND2 (N13226, N13222, N4481);
nor NOR4 (N13227, N13226, N6674, N3075, N9789);
nand NAND3 (N13228, N13193, N2934, N9356);
buf BUF1 (N13229, N13216);
not NOT1 (N13230, N13219);
nor NOR4 (N13231, N13223, N5595, N12659, N55);
buf BUF1 (N13232, N13224);
buf BUF1 (N13233, N13217);
and AND4 (N13234, N13230, N5616, N7073, N6968);
nand NAND2 (N13235, N13233, N4761);
buf BUF1 (N13236, N13228);
not NOT1 (N13237, N13213);
xor XOR2 (N13238, N13220, N8523);
xor XOR2 (N13239, N13229, N8616);
nor NOR3 (N13240, N13239, N5403, N11999);
buf BUF1 (N13241, N13237);
buf BUF1 (N13242, N13225);
nor NOR4 (N13243, N13234, N439, N483, N9263);
xor XOR2 (N13244, N13231, N7343);
and AND4 (N13245, N13240, N10013, N8738, N6427);
not NOT1 (N13246, N13232);
nor NOR4 (N13247, N13227, N11169, N4132, N8979);
nor NOR4 (N13248, N13245, N12740, N2615, N6672);
nand NAND3 (N13249, N13243, N11030, N4554);
xor XOR2 (N13250, N13235, N7030);
xor XOR2 (N13251, N13241, N5025);
buf BUF1 (N13252, N13249);
buf BUF1 (N13253, N13247);
nand NAND4 (N13254, N13251, N535, N8635, N5272);
not NOT1 (N13255, N13246);
and AND3 (N13256, N13236, N11342, N6310);
not NOT1 (N13257, N13248);
buf BUF1 (N13258, N13252);
nor NOR2 (N13259, N13250, N691);
xor XOR2 (N13260, N13259, N7659);
and AND4 (N13261, N13256, N2718, N10860, N13128);
buf BUF1 (N13262, N13238);
buf BUF1 (N13263, N13242);
xor XOR2 (N13264, N13253, N1909);
nand NAND2 (N13265, N13254, N944);
buf BUF1 (N13266, N13264);
not NOT1 (N13267, N13262);
or OR4 (N13268, N13263, N8467, N11089, N12516);
nor NOR4 (N13269, N13266, N10817, N11547, N2264);
nand NAND2 (N13270, N13257, N10308);
or OR3 (N13271, N13258, N6982, N13093);
and AND3 (N13272, N13268, N1617, N10315);
and AND2 (N13273, N13269, N2167);
buf BUF1 (N13274, N13261);
xor XOR2 (N13275, N13244, N3921);
xor XOR2 (N13276, N13274, N10622);
buf BUF1 (N13277, N13276);
or OR2 (N13278, N13267, N6890);
xor XOR2 (N13279, N13265, N2095);
buf BUF1 (N13280, N13273);
nand NAND2 (N13281, N13260, N6057);
nor NOR3 (N13282, N13275, N11227, N1676);
buf BUF1 (N13283, N13279);
and AND4 (N13284, N13283, N11099, N3903, N3058);
not NOT1 (N13285, N13271);
nor NOR4 (N13286, N13255, N7718, N2071, N1239);
nand NAND4 (N13287, N13280, N11504, N1767, N2562);
nand NAND3 (N13288, N13278, N8836, N11477);
nor NOR4 (N13289, N13281, N10585, N5311, N1011);
xor XOR2 (N13290, N13277, N7503);
nor NOR3 (N13291, N13286, N1179, N4862);
and AND3 (N13292, N13282, N10305, N342);
not NOT1 (N13293, N13287);
nor NOR3 (N13294, N13272, N9841, N10823);
and AND4 (N13295, N13290, N25, N8362, N5883);
xor XOR2 (N13296, N13295, N8520);
not NOT1 (N13297, N13293);
nand NAND3 (N13298, N13296, N11420, N10130);
buf BUF1 (N13299, N13298);
and AND3 (N13300, N13285, N7935, N12115);
not NOT1 (N13301, N13284);
nor NOR4 (N13302, N13294, N2012, N8585, N11568);
not NOT1 (N13303, N13292);
nor NOR4 (N13304, N13270, N6577, N5095, N3887);
or OR4 (N13305, N13301, N9103, N5284, N10525);
xor XOR2 (N13306, N13305, N3107);
or OR4 (N13307, N13289, N3662, N8466, N10592);
xor XOR2 (N13308, N13288, N2296);
and AND2 (N13309, N13304, N3315);
or OR4 (N13310, N13306, N3686, N3043, N4588);
buf BUF1 (N13311, N13302);
or OR2 (N13312, N13291, N4299);
buf BUF1 (N13313, N13297);
nand NAND4 (N13314, N13312, N10064, N7992, N7552);
and AND3 (N13315, N13300, N7274, N4747);
xor XOR2 (N13316, N13303, N3577);
xor XOR2 (N13317, N13316, N4250);
and AND4 (N13318, N13309, N3425, N1165, N11015);
xor XOR2 (N13319, N13317, N7504);
not NOT1 (N13320, N13315);
nor NOR3 (N13321, N13307, N11265, N5955);
nand NAND4 (N13322, N13318, N852, N11979, N4734);
nand NAND2 (N13323, N13319, N5008);
nor NOR3 (N13324, N13320, N4953, N1363);
buf BUF1 (N13325, N13314);
nand NAND4 (N13326, N13308, N4527, N8604, N3347);
not NOT1 (N13327, N13323);
nand NAND2 (N13328, N13310, N7876);
buf BUF1 (N13329, N13326);
and AND2 (N13330, N13324, N8858);
nor NOR4 (N13331, N13321, N11177, N4226, N8398);
nor NOR3 (N13332, N13322, N4314, N11727);
nor NOR2 (N13333, N13331, N10530);
buf BUF1 (N13334, N13332);
nor NOR2 (N13335, N13334, N3933);
or OR3 (N13336, N13325, N12742, N10360);
and AND2 (N13337, N13329, N2071);
nor NOR4 (N13338, N13333, N4085, N7816, N5192);
and AND2 (N13339, N13338, N1918);
buf BUF1 (N13340, N13330);
buf BUF1 (N13341, N13299);
nand NAND3 (N13342, N13336, N6384, N1993);
not NOT1 (N13343, N13339);
nor NOR4 (N13344, N13327, N9193, N8249, N12000);
nand NAND2 (N13345, N13343, N11146);
not NOT1 (N13346, N13341);
and AND3 (N13347, N13335, N8727, N961);
not NOT1 (N13348, N13346);
xor XOR2 (N13349, N13348, N1059);
buf BUF1 (N13350, N13347);
nand NAND4 (N13351, N13345, N4720, N900, N4835);
buf BUF1 (N13352, N13313);
and AND4 (N13353, N13340, N3732, N423, N9289);
and AND3 (N13354, N13349, N7834, N7539);
buf BUF1 (N13355, N13352);
nor NOR4 (N13356, N13354, N4322, N344, N11223);
or OR4 (N13357, N13328, N12435, N4459, N3906);
or OR3 (N13358, N13344, N8445, N8338);
nand NAND2 (N13359, N13355, N11671);
or OR3 (N13360, N13358, N13227, N7439);
nor NOR2 (N13361, N13350, N6202);
nand NAND2 (N13362, N13337, N1975);
nor NOR2 (N13363, N13311, N2408);
or OR4 (N13364, N13361, N2998, N2754, N2221);
nor NOR3 (N13365, N13363, N1929, N9033);
xor XOR2 (N13366, N13353, N2158);
xor XOR2 (N13367, N13362, N216);
nand NAND3 (N13368, N13359, N11616, N4586);
or OR3 (N13369, N13342, N9423, N349);
xor XOR2 (N13370, N13364, N2600);
nor NOR4 (N13371, N13367, N1662, N9208, N10041);
nand NAND4 (N13372, N13360, N67, N11169, N7638);
not NOT1 (N13373, N13365);
not NOT1 (N13374, N13372);
not NOT1 (N13375, N13366);
nor NOR4 (N13376, N13351, N9355, N672, N9992);
and AND2 (N13377, N13376, N31);
nand NAND3 (N13378, N13370, N851, N9319);
or OR4 (N13379, N13378, N2064, N12652, N3162);
nor NOR2 (N13380, N13371, N3716);
xor XOR2 (N13381, N13369, N7598);
or OR4 (N13382, N13356, N12588, N486, N10220);
buf BUF1 (N13383, N13379);
xor XOR2 (N13384, N13374, N10441);
nor NOR4 (N13385, N13384, N9808, N4778, N1224);
not NOT1 (N13386, N13385);
buf BUF1 (N13387, N13383);
nand NAND2 (N13388, N13375, N9998);
not NOT1 (N13389, N13381);
or OR4 (N13390, N13357, N4358, N12292, N9745);
buf BUF1 (N13391, N13389);
nand NAND2 (N13392, N13386, N4281);
buf BUF1 (N13393, N13391);
and AND2 (N13394, N13368, N3278);
xor XOR2 (N13395, N13390, N1679);
nand NAND3 (N13396, N13380, N13363, N12525);
or OR2 (N13397, N13388, N7121);
and AND3 (N13398, N13377, N12678, N3555);
buf BUF1 (N13399, N13393);
and AND3 (N13400, N13387, N1819, N1919);
buf BUF1 (N13401, N13382);
nor NOR2 (N13402, N13373, N12928);
buf BUF1 (N13403, N13395);
nor NOR2 (N13404, N13402, N4155);
nand NAND2 (N13405, N13394, N4259);
nand NAND2 (N13406, N13401, N14);
nor NOR4 (N13407, N13397, N10108, N9095, N3339);
and AND4 (N13408, N13407, N11115, N5648, N11065);
nor NOR2 (N13409, N13399, N9810);
buf BUF1 (N13410, N13404);
not NOT1 (N13411, N13409);
and AND4 (N13412, N13392, N13120, N4792, N1872);
nand NAND2 (N13413, N13408, N237);
xor XOR2 (N13414, N13403, N7466);
and AND3 (N13415, N13400, N4233, N9981);
not NOT1 (N13416, N13405);
and AND2 (N13417, N13411, N524);
and AND4 (N13418, N13396, N1548, N6431, N255);
not NOT1 (N13419, N13416);
or OR3 (N13420, N13419, N11731, N12467);
and AND4 (N13421, N13412, N2303, N13318, N10969);
and AND3 (N13422, N13398, N7693, N9491);
nand NAND3 (N13423, N13421, N6333, N8886);
not NOT1 (N13424, N13423);
or OR2 (N13425, N13418, N2812);
or OR2 (N13426, N13422, N12578);
nor NOR2 (N13427, N13415, N8690);
nand NAND2 (N13428, N13420, N7700);
and AND4 (N13429, N13426, N7202, N10050, N403);
xor XOR2 (N13430, N13428, N2557);
xor XOR2 (N13431, N13410, N2254);
xor XOR2 (N13432, N13427, N11957);
buf BUF1 (N13433, N13414);
xor XOR2 (N13434, N13425, N13220);
and AND2 (N13435, N13413, N11041);
or OR4 (N13436, N13435, N9596, N8011, N799);
nand NAND3 (N13437, N13432, N6465, N7956);
nand NAND4 (N13438, N13429, N2558, N6595, N3305);
nand NAND3 (N13439, N13424, N734, N1182);
not NOT1 (N13440, N13417);
nand NAND3 (N13441, N13439, N11911, N4379);
not NOT1 (N13442, N13438);
nand NAND3 (N13443, N13441, N10298, N12226);
nand NAND2 (N13444, N13430, N2430);
nor NOR2 (N13445, N13443, N12428);
buf BUF1 (N13446, N13406);
nor NOR3 (N13447, N13442, N7241, N10);
nor NOR4 (N13448, N13437, N2290, N9242, N13127);
or OR2 (N13449, N13431, N8911);
buf BUF1 (N13450, N13446);
or OR3 (N13451, N13448, N10153, N7640);
and AND4 (N13452, N13433, N9758, N9998, N4242);
not NOT1 (N13453, N13450);
nor NOR4 (N13454, N13434, N1029, N2420, N10146);
nand NAND4 (N13455, N13436, N6793, N4661, N6379);
nor NOR3 (N13456, N13445, N1424, N10295);
nand NAND2 (N13457, N13444, N2775);
not NOT1 (N13458, N13452);
buf BUF1 (N13459, N13455);
nand NAND4 (N13460, N13457, N6356, N69, N1805);
nand NAND3 (N13461, N13459, N10475, N6976);
xor XOR2 (N13462, N13461, N8849);
and AND2 (N13463, N13453, N6822);
nand NAND2 (N13464, N13460, N12574);
not NOT1 (N13465, N13440);
nand NAND2 (N13466, N13456, N6961);
not NOT1 (N13467, N13464);
not NOT1 (N13468, N13454);
xor XOR2 (N13469, N13451, N7956);
nand NAND4 (N13470, N13463, N9798, N1511, N4562);
buf BUF1 (N13471, N13447);
nor NOR3 (N13472, N13470, N12954, N2521);
nor NOR4 (N13473, N13462, N3989, N11827, N13004);
and AND4 (N13474, N13465, N7753, N1710, N3760);
nor NOR2 (N13475, N13467, N11705);
buf BUF1 (N13476, N13473);
not NOT1 (N13477, N13476);
not NOT1 (N13478, N13469);
not NOT1 (N13479, N13477);
not NOT1 (N13480, N13466);
or OR3 (N13481, N13449, N1149, N10140);
nand NAND3 (N13482, N13458, N11543, N2900);
xor XOR2 (N13483, N13475, N10433);
nand NAND3 (N13484, N13472, N2035, N8514);
xor XOR2 (N13485, N13482, N2738);
not NOT1 (N13486, N13468);
nand NAND3 (N13487, N13478, N12524, N6492);
buf BUF1 (N13488, N13485);
not NOT1 (N13489, N13481);
or OR2 (N13490, N13484, N8814);
or OR4 (N13491, N13474, N6194, N931, N488);
nor NOR4 (N13492, N13471, N2129, N1234, N8088);
nor NOR4 (N13493, N13489, N10520, N1322, N12058);
and AND3 (N13494, N13491, N12416, N589);
xor XOR2 (N13495, N13493, N3708);
or OR2 (N13496, N13479, N5990);
buf BUF1 (N13497, N13488);
nand NAND4 (N13498, N13486, N11068, N2877, N3403);
nor NOR2 (N13499, N13480, N4914);
nor NOR4 (N13500, N13487, N4910, N2741, N9890);
nor NOR3 (N13501, N13496, N7432, N12086);
not NOT1 (N13502, N13483);
xor XOR2 (N13503, N13494, N6601);
not NOT1 (N13504, N13499);
or OR3 (N13505, N13502, N851, N8935);
buf BUF1 (N13506, N13490);
not NOT1 (N13507, N13497);
not NOT1 (N13508, N13500);
buf BUF1 (N13509, N13492);
buf BUF1 (N13510, N13504);
nand NAND2 (N13511, N13503, N7626);
nor NOR3 (N13512, N13501, N1904, N1721);
not NOT1 (N13513, N13505);
not NOT1 (N13514, N13508);
nand NAND3 (N13515, N13509, N12883, N2786);
buf BUF1 (N13516, N13513);
nor NOR2 (N13517, N13514, N9560);
or OR4 (N13518, N13506, N10735, N12936, N2626);
buf BUF1 (N13519, N13518);
buf BUF1 (N13520, N13517);
and AND2 (N13521, N13511, N6287);
not NOT1 (N13522, N13515);
nand NAND3 (N13523, N13498, N9217, N6750);
nor NOR2 (N13524, N13507, N7176);
buf BUF1 (N13525, N13495);
nor NOR2 (N13526, N13510, N10998);
and AND3 (N13527, N13512, N2145, N1353);
nor NOR4 (N13528, N13522, N10062, N5279, N10712);
and AND4 (N13529, N13523, N10155, N8497, N13460);
not NOT1 (N13530, N13529);
not NOT1 (N13531, N13520);
not NOT1 (N13532, N13519);
and AND4 (N13533, N13528, N3815, N4446, N245);
buf BUF1 (N13534, N13527);
buf BUF1 (N13535, N13526);
or OR4 (N13536, N13533, N5239, N7427, N7123);
nor NOR3 (N13537, N13524, N4805, N6169);
not NOT1 (N13538, N13531);
buf BUF1 (N13539, N13537);
xor XOR2 (N13540, N13532, N11760);
nor NOR3 (N13541, N13539, N40, N11451);
nor NOR3 (N13542, N13535, N1778, N5426);
xor XOR2 (N13543, N13541, N3525);
xor XOR2 (N13544, N13540, N6595);
not NOT1 (N13545, N13543);
nand NAND2 (N13546, N13536, N10993);
and AND3 (N13547, N13521, N9036, N2060);
nand NAND4 (N13548, N13547, N825, N3589, N2073);
not NOT1 (N13549, N13538);
nand NAND3 (N13550, N13534, N77, N4549);
and AND3 (N13551, N13546, N12389, N5764);
nand NAND2 (N13552, N13530, N11953);
nand NAND2 (N13553, N13516, N5824);
nand NAND2 (N13554, N13553, N10874);
nor NOR4 (N13555, N13549, N4349, N862, N13426);
buf BUF1 (N13556, N13552);
nor NOR4 (N13557, N13525, N11502, N8207, N8164);
nor NOR3 (N13558, N13548, N375, N11476);
not NOT1 (N13559, N13544);
and AND4 (N13560, N13554, N5965, N4035, N11547);
buf BUF1 (N13561, N13559);
and AND3 (N13562, N13542, N11317, N11188);
or OR2 (N13563, N13557, N6154);
nand NAND3 (N13564, N13560, N4139, N8415);
nor NOR4 (N13565, N13562, N4522, N6745, N7527);
and AND3 (N13566, N13550, N5484, N1175);
and AND2 (N13567, N13563, N3564);
not NOT1 (N13568, N13556);
and AND2 (N13569, N13551, N977);
and AND2 (N13570, N13565, N5114);
xor XOR2 (N13571, N13545, N437);
and AND3 (N13572, N13566, N2151, N1423);
buf BUF1 (N13573, N13561);
nand NAND4 (N13574, N13555, N6861, N8113, N10917);
xor XOR2 (N13575, N13567, N1479);
or OR4 (N13576, N13569, N2485, N8789, N9031);
buf BUF1 (N13577, N13572);
not NOT1 (N13578, N13574);
and AND4 (N13579, N13564, N4973, N6888, N6986);
not NOT1 (N13580, N13576);
buf BUF1 (N13581, N13577);
xor XOR2 (N13582, N13578, N6747);
buf BUF1 (N13583, N13575);
xor XOR2 (N13584, N13558, N5021);
xor XOR2 (N13585, N13579, N9113);
and AND3 (N13586, N13582, N4357, N1076);
not NOT1 (N13587, N13570);
buf BUF1 (N13588, N13585);
or OR3 (N13589, N13573, N9015, N969);
not NOT1 (N13590, N13588);
and AND4 (N13591, N13586, N12063, N12458, N6866);
or OR4 (N13592, N13581, N1634, N10144, N3297);
nand NAND2 (N13593, N13584, N5377);
nor NOR2 (N13594, N13587, N4887);
nor NOR2 (N13595, N13590, N9056);
nand NAND4 (N13596, N13593, N10967, N8482, N5952);
not NOT1 (N13597, N13589);
xor XOR2 (N13598, N13583, N1174);
and AND4 (N13599, N13592, N323, N4124, N4800);
and AND3 (N13600, N13571, N56, N12272);
not NOT1 (N13601, N13596);
nor NOR3 (N13602, N13591, N1322, N7551);
nand NAND4 (N13603, N13568, N363, N4857, N11839);
xor XOR2 (N13604, N13594, N9918);
xor XOR2 (N13605, N13604, N8922);
nand NAND4 (N13606, N13602, N7449, N5946, N10672);
nand NAND3 (N13607, N13605, N769, N289);
and AND2 (N13608, N13601, N2451);
buf BUF1 (N13609, N13607);
buf BUF1 (N13610, N13599);
and AND3 (N13611, N13603, N3242, N7685);
not NOT1 (N13612, N13595);
not NOT1 (N13613, N13612);
nand NAND3 (N13614, N13611, N11409, N1411);
nor NOR4 (N13615, N13606, N8502, N6990, N5429);
nand NAND3 (N13616, N13580, N80, N9259);
nor NOR4 (N13617, N13613, N11599, N10390, N190);
nor NOR3 (N13618, N13597, N11411, N1082);
xor XOR2 (N13619, N13616, N10747);
buf BUF1 (N13620, N13608);
and AND3 (N13621, N13615, N12857, N5079);
buf BUF1 (N13622, N13610);
nand NAND4 (N13623, N13621, N11936, N9690, N7404);
and AND4 (N13624, N13619, N10385, N2814, N5486);
nor NOR2 (N13625, N13614, N1757);
buf BUF1 (N13626, N13598);
or OR4 (N13627, N13624, N7982, N5078, N10369);
xor XOR2 (N13628, N13627, N1048);
and AND2 (N13629, N13609, N1489);
nand NAND4 (N13630, N13622, N6417, N3624, N12772);
not NOT1 (N13631, N13600);
or OR4 (N13632, N13617, N715, N6189, N6273);
nor NOR3 (N13633, N13631, N11994, N13004);
or OR2 (N13634, N13630, N11250);
buf BUF1 (N13635, N13620);
nor NOR3 (N13636, N13629, N8312, N7436);
and AND4 (N13637, N13618, N3878, N10595, N8441);
nand NAND3 (N13638, N13632, N9536, N5762);
not NOT1 (N13639, N13637);
not NOT1 (N13640, N13626);
nor NOR2 (N13641, N13635, N1451);
or OR4 (N13642, N13634, N8791, N5443, N3684);
and AND3 (N13643, N13628, N417, N8266);
and AND4 (N13644, N13633, N1831, N5230, N13170);
not NOT1 (N13645, N13643);
not NOT1 (N13646, N13640);
and AND2 (N13647, N13642, N12112);
or OR3 (N13648, N13647, N5328, N3036);
or OR2 (N13649, N13645, N4683);
and AND3 (N13650, N13623, N12041, N7312);
xor XOR2 (N13651, N13646, N11441);
nor NOR2 (N13652, N13644, N2053);
and AND3 (N13653, N13639, N4383, N13248);
nand NAND4 (N13654, N13625, N7546, N12859, N12515);
nand NAND2 (N13655, N13654, N4287);
not NOT1 (N13656, N13641);
xor XOR2 (N13657, N13656, N4725);
or OR3 (N13658, N13648, N8937, N9660);
or OR3 (N13659, N13653, N6017, N8725);
and AND3 (N13660, N13650, N3468, N4848);
or OR4 (N13661, N13658, N12491, N1250, N6836);
xor XOR2 (N13662, N13636, N1936);
buf BUF1 (N13663, N13661);
xor XOR2 (N13664, N13659, N10061);
or OR3 (N13665, N13657, N1445, N7356);
not NOT1 (N13666, N13655);
nor NOR4 (N13667, N13638, N9178, N12370, N3501);
buf BUF1 (N13668, N13651);
or OR2 (N13669, N13660, N10231);
buf BUF1 (N13670, N13667);
or OR3 (N13671, N13670, N1346, N2669);
xor XOR2 (N13672, N13666, N13180);
nand NAND3 (N13673, N13649, N11818, N11026);
nor NOR4 (N13674, N13672, N11371, N11064, N11551);
xor XOR2 (N13675, N13669, N9985);
buf BUF1 (N13676, N13671);
buf BUF1 (N13677, N13663);
xor XOR2 (N13678, N13674, N3627);
buf BUF1 (N13679, N13675);
and AND4 (N13680, N13678, N484, N5202, N3149);
nand NAND2 (N13681, N13676, N4930);
not NOT1 (N13682, N13652);
nand NAND2 (N13683, N13664, N5693);
buf BUF1 (N13684, N13682);
not NOT1 (N13685, N13668);
nor NOR2 (N13686, N13677, N10941);
nand NAND4 (N13687, N13685, N3648, N2887, N5318);
xor XOR2 (N13688, N13665, N6075);
buf BUF1 (N13689, N13686);
and AND4 (N13690, N13687, N12373, N13489, N6999);
nor NOR2 (N13691, N13681, N9487);
xor XOR2 (N13692, N13680, N10803);
nand NAND3 (N13693, N13691, N587, N6153);
buf BUF1 (N13694, N13679);
or OR2 (N13695, N13693, N9471);
or OR3 (N13696, N13689, N12737, N3011);
and AND2 (N13697, N13688, N6480);
or OR2 (N13698, N13684, N12075);
or OR3 (N13699, N13695, N2182, N1955);
and AND4 (N13700, N13696, N10763, N9492, N5633);
and AND2 (N13701, N13699, N67);
xor XOR2 (N13702, N13694, N11388);
buf BUF1 (N13703, N13673);
or OR4 (N13704, N13703, N8718, N3101, N13042);
nand NAND3 (N13705, N13690, N3276, N1777);
not NOT1 (N13706, N13701);
or OR2 (N13707, N13705, N10349);
buf BUF1 (N13708, N13707);
nor NOR3 (N13709, N13697, N7410, N8376);
nor NOR4 (N13710, N13683, N7407, N9438, N9849);
and AND3 (N13711, N13662, N288, N13387);
nand NAND4 (N13712, N13706, N3422, N7030, N12933);
and AND2 (N13713, N13702, N1895);
and AND3 (N13714, N13700, N5644, N5549);
nor NOR2 (N13715, N13692, N2918);
not NOT1 (N13716, N13713);
buf BUF1 (N13717, N13709);
not NOT1 (N13718, N13698);
buf BUF1 (N13719, N13704);
nand NAND4 (N13720, N13708, N8488, N7299, N5279);
and AND2 (N13721, N13716, N8989);
nor NOR3 (N13722, N13717, N3595, N6585);
xor XOR2 (N13723, N13711, N2199);
nor NOR2 (N13724, N13710, N5575);
nor NOR4 (N13725, N13722, N9032, N6105, N1957);
or OR3 (N13726, N13723, N4599, N986);
nor NOR4 (N13727, N13719, N11118, N12319, N5356);
nor NOR3 (N13728, N13718, N1154, N5214);
or OR2 (N13729, N13721, N3163);
and AND4 (N13730, N13729, N8471, N6774, N4277);
or OR4 (N13731, N13730, N8028, N11895, N12558);
or OR4 (N13732, N13731, N4408, N5533, N1315);
and AND2 (N13733, N13720, N13229);
buf BUF1 (N13734, N13725);
not NOT1 (N13735, N13733);
or OR4 (N13736, N13728, N9753, N3062, N6816);
or OR3 (N13737, N13714, N1226, N4739);
nand NAND3 (N13738, N13734, N12991, N12708);
not NOT1 (N13739, N13737);
and AND4 (N13740, N13739, N7234, N9570, N10923);
nor NOR3 (N13741, N13736, N2701, N3164);
xor XOR2 (N13742, N13741, N9271);
nand NAND4 (N13743, N13735, N13666, N9353, N2935);
nand NAND4 (N13744, N13743, N5448, N2339, N11022);
not NOT1 (N13745, N13727);
or OR4 (N13746, N13745, N13411, N1582, N5108);
nor NOR2 (N13747, N13715, N13333);
buf BUF1 (N13748, N13738);
nand NAND4 (N13749, N13724, N10580, N5713, N8395);
nand NAND4 (N13750, N13742, N7890, N12447, N2263);
or OR4 (N13751, N13748, N10545, N7244, N10032);
nand NAND2 (N13752, N13740, N9536);
buf BUF1 (N13753, N13712);
buf BUF1 (N13754, N13747);
and AND4 (N13755, N13749, N11712, N12861, N1397);
not NOT1 (N13756, N13755);
xor XOR2 (N13757, N13744, N3299);
buf BUF1 (N13758, N13754);
or OR3 (N13759, N13751, N862, N7474);
nor NOR4 (N13760, N13732, N8841, N7759, N10294);
nor NOR4 (N13761, N13752, N2759, N12502, N3161);
nand NAND3 (N13762, N13761, N3273, N5463);
xor XOR2 (N13763, N13746, N7520);
or OR3 (N13764, N13757, N5826, N3875);
nor NOR2 (N13765, N13756, N12249);
nor NOR4 (N13766, N13763, N9253, N536, N7318);
not NOT1 (N13767, N13753);
not NOT1 (N13768, N13760);
not NOT1 (N13769, N13726);
or OR3 (N13770, N13759, N6688, N5796);
nand NAND3 (N13771, N13769, N9062, N2302);
or OR2 (N13772, N13767, N10464);
nor NOR4 (N13773, N13768, N10368, N3518, N10668);
nand NAND4 (N13774, N13765, N1843, N9053, N347);
nor NOR2 (N13775, N13764, N4144);
or OR3 (N13776, N13774, N5755, N4775);
nor NOR4 (N13777, N13772, N11387, N6510, N6934);
or OR3 (N13778, N13777, N9259, N9209);
nand NAND4 (N13779, N13750, N3134, N2613, N8179);
nand NAND2 (N13780, N13775, N7447);
xor XOR2 (N13781, N13758, N10430);
nor NOR3 (N13782, N13773, N3567, N2612);
buf BUF1 (N13783, N13770);
not NOT1 (N13784, N13762);
and AND2 (N13785, N13766, N7792);
not NOT1 (N13786, N13784);
nor NOR3 (N13787, N13779, N5715, N1783);
and AND3 (N13788, N13787, N254, N130);
not NOT1 (N13789, N13781);
or OR2 (N13790, N13771, N3996);
not NOT1 (N13791, N13785);
buf BUF1 (N13792, N13789);
and AND2 (N13793, N13791, N6998);
nor NOR2 (N13794, N13778, N13137);
or OR4 (N13795, N13788, N4330, N13487, N8844);
xor XOR2 (N13796, N13776, N11338);
buf BUF1 (N13797, N13795);
xor XOR2 (N13798, N13792, N10864);
buf BUF1 (N13799, N13796);
buf BUF1 (N13800, N13790);
nor NOR3 (N13801, N13798, N10763, N9119);
nor NOR4 (N13802, N13800, N11636, N3250, N5543);
xor XOR2 (N13803, N13786, N3278);
not NOT1 (N13804, N13780);
and AND2 (N13805, N13793, N12548);
or OR2 (N13806, N13804, N2226);
xor XOR2 (N13807, N13801, N12561);
or OR4 (N13808, N13783, N3073, N10878, N7415);
not NOT1 (N13809, N13803);
nand NAND3 (N13810, N13809, N1755, N6443);
and AND3 (N13811, N13807, N6240, N1564);
and AND4 (N13812, N13806, N6866, N13680, N4814);
xor XOR2 (N13813, N13812, N6443);
xor XOR2 (N13814, N13802, N755);
and AND3 (N13815, N13794, N8659, N3005);
nor NOR2 (N13816, N13811, N6656);
and AND3 (N13817, N13805, N11997, N536);
nor NOR4 (N13818, N13782, N4199, N6597, N10246);
nor NOR4 (N13819, N13808, N1913, N7030, N12995);
nor NOR3 (N13820, N13819, N1750, N1767);
buf BUF1 (N13821, N13799);
nor NOR4 (N13822, N13820, N4058, N3142, N4249);
buf BUF1 (N13823, N13810);
nand NAND2 (N13824, N13821, N8418);
or OR2 (N13825, N13815, N1930);
nor NOR2 (N13826, N13813, N4588);
not NOT1 (N13827, N13817);
buf BUF1 (N13828, N13816);
and AND2 (N13829, N13826, N7148);
not NOT1 (N13830, N13797);
nor NOR4 (N13831, N13822, N6581, N10312, N12779);
and AND2 (N13832, N13818, N4982);
xor XOR2 (N13833, N13814, N10171);
xor XOR2 (N13834, N13829, N5404);
buf BUF1 (N13835, N13833);
and AND4 (N13836, N13830, N8526, N12995, N4749);
and AND3 (N13837, N13835, N4518, N12591);
not NOT1 (N13838, N13831);
nand NAND2 (N13839, N13825, N830);
or OR2 (N13840, N13837, N4869);
or OR4 (N13841, N13838, N13233, N7441, N3957);
not NOT1 (N13842, N13840);
xor XOR2 (N13843, N13842, N11367);
xor XOR2 (N13844, N13827, N3385);
xor XOR2 (N13845, N13843, N1456);
buf BUF1 (N13846, N13844);
or OR3 (N13847, N13832, N8879, N11321);
not NOT1 (N13848, N13828);
nand NAND2 (N13849, N13845, N8645);
nor NOR2 (N13850, N13841, N10568);
xor XOR2 (N13851, N13839, N1563);
and AND2 (N13852, N13834, N12001);
nor NOR4 (N13853, N13847, N10385, N6064, N2690);
and AND2 (N13854, N13824, N7146);
nand NAND4 (N13855, N13849, N1828, N12716, N1035);
nor NOR3 (N13856, N13846, N4029, N1379);
buf BUF1 (N13857, N13848);
or OR3 (N13858, N13852, N9357, N3514);
nor NOR4 (N13859, N13851, N5410, N351, N3895);
nand NAND3 (N13860, N13823, N4902, N13158);
and AND4 (N13861, N13856, N4817, N8703, N11476);
and AND3 (N13862, N13853, N12039, N8022);
buf BUF1 (N13863, N13860);
buf BUF1 (N13864, N13850);
or OR4 (N13865, N13861, N1492, N9562, N5247);
xor XOR2 (N13866, N13836, N11168);
nand NAND4 (N13867, N13866, N3207, N9655, N1073);
xor XOR2 (N13868, N13867, N4255);
xor XOR2 (N13869, N13862, N777);
or OR3 (N13870, N13869, N13544, N6211);
or OR2 (N13871, N13864, N8329);
buf BUF1 (N13872, N13870);
nand NAND2 (N13873, N13865, N10621);
not NOT1 (N13874, N13868);
buf BUF1 (N13875, N13873);
and AND4 (N13876, N13863, N10140, N3438, N5192);
not NOT1 (N13877, N13855);
nor NOR3 (N13878, N13857, N8646, N2071);
nand NAND4 (N13879, N13877, N11278, N8160, N6196);
not NOT1 (N13880, N13872);
nand NAND4 (N13881, N13875, N9603, N7527, N6617);
buf BUF1 (N13882, N13858);
or OR2 (N13883, N13859, N6735);
nand NAND4 (N13884, N13879, N11936, N974, N10114);
or OR4 (N13885, N13871, N1728, N1541, N1861);
nor NOR4 (N13886, N13885, N4041, N6688, N10230);
xor XOR2 (N13887, N13882, N2335);
or OR3 (N13888, N13884, N7962, N6016);
buf BUF1 (N13889, N13886);
nand NAND3 (N13890, N13889, N13102, N9619);
xor XOR2 (N13891, N13887, N7134);
not NOT1 (N13892, N13854);
nand NAND2 (N13893, N13883, N212);
not NOT1 (N13894, N13892);
buf BUF1 (N13895, N13881);
nor NOR2 (N13896, N13891, N13060);
not NOT1 (N13897, N13895);
not NOT1 (N13898, N13878);
nand NAND2 (N13899, N13897, N4070);
xor XOR2 (N13900, N13893, N604);
nor NOR3 (N13901, N13894, N10031, N10154);
nor NOR3 (N13902, N13898, N4552, N9904);
buf BUF1 (N13903, N13902);
xor XOR2 (N13904, N13901, N10637);
and AND4 (N13905, N13896, N4074, N8730, N13501);
not NOT1 (N13906, N13890);
or OR2 (N13907, N13900, N11938);
xor XOR2 (N13908, N13904, N7270);
nand NAND4 (N13909, N13906, N2225, N9007, N7101);
or OR4 (N13910, N13909, N3466, N8925, N1384);
buf BUF1 (N13911, N13910);
nor NOR2 (N13912, N13903, N13842);
not NOT1 (N13913, N13907);
buf BUF1 (N13914, N13880);
nor NOR3 (N13915, N13908, N10027, N1129);
and AND3 (N13916, N13911, N20, N13203);
not NOT1 (N13917, N13912);
and AND3 (N13918, N13874, N12161, N6652);
nand NAND3 (N13919, N13905, N79, N10810);
nor NOR2 (N13920, N13876, N4011);
nor NOR3 (N13921, N13918, N3257, N5028);
or OR2 (N13922, N13920, N3438);
not NOT1 (N13923, N13888);
nand NAND2 (N13924, N13921, N9783);
buf BUF1 (N13925, N13922);
xor XOR2 (N13926, N13925, N1611);
nand NAND2 (N13927, N13914, N5854);
not NOT1 (N13928, N13923);
nor NOR2 (N13929, N13899, N352);
buf BUF1 (N13930, N13928);
xor XOR2 (N13931, N13916, N4650);
xor XOR2 (N13932, N13926, N7077);
and AND2 (N13933, N13929, N75);
buf BUF1 (N13934, N13927);
xor XOR2 (N13935, N13915, N6676);
or OR2 (N13936, N13924, N12040);
or OR2 (N13937, N13930, N13807);
xor XOR2 (N13938, N13919, N9184);
and AND3 (N13939, N13934, N6181, N6108);
buf BUF1 (N13940, N13939);
buf BUF1 (N13941, N13913);
nand NAND4 (N13942, N13938, N5117, N9082, N8025);
not NOT1 (N13943, N13936);
nand NAND4 (N13944, N13935, N6145, N12942, N11868);
not NOT1 (N13945, N13933);
nor NOR4 (N13946, N13931, N10381, N11782, N7351);
nor NOR2 (N13947, N13945, N7437);
nor NOR2 (N13948, N13940, N2110);
or OR4 (N13949, N13917, N7457, N13831, N6370);
and AND4 (N13950, N13941, N13931, N5020, N4304);
not NOT1 (N13951, N13942);
buf BUF1 (N13952, N13949);
nor NOR4 (N13953, N13932, N11344, N12739, N13584);
nor NOR4 (N13954, N13950, N12000, N13128, N7924);
and AND3 (N13955, N13954, N2161, N1481);
nor NOR3 (N13956, N13948, N10053, N11997);
or OR4 (N13957, N13955, N13134, N7076, N2837);
buf BUF1 (N13958, N13947);
and AND4 (N13959, N13957, N9672, N6207, N4481);
or OR3 (N13960, N13937, N7523, N7133);
xor XOR2 (N13961, N13952, N3642);
nor NOR2 (N13962, N13960, N3556);
nor NOR4 (N13963, N13961, N13720, N5257, N5817);
xor XOR2 (N13964, N13943, N664);
buf BUF1 (N13965, N13944);
buf BUF1 (N13966, N13946);
not NOT1 (N13967, N13966);
or OR4 (N13968, N13967, N5836, N7620, N8438);
buf BUF1 (N13969, N13951);
xor XOR2 (N13970, N13956, N2067);
xor XOR2 (N13971, N13970, N12632);
not NOT1 (N13972, N13958);
buf BUF1 (N13973, N13965);
not NOT1 (N13974, N13972);
buf BUF1 (N13975, N13953);
xor XOR2 (N13976, N13959, N13457);
nand NAND2 (N13977, N13968, N9);
or OR4 (N13978, N13962, N8217, N3073, N13794);
nand NAND3 (N13979, N13974, N8584, N10771);
nor NOR3 (N13980, N13963, N6006, N1406);
and AND2 (N13981, N13971, N9948);
nand NAND2 (N13982, N13975, N4424);
nor NOR3 (N13983, N13979, N13640, N13227);
or OR3 (N13984, N13983, N10924, N4432);
and AND4 (N13985, N13980, N1944, N4973, N5761);
xor XOR2 (N13986, N13984, N6605);
nand NAND2 (N13987, N13964, N12871);
nand NAND3 (N13988, N13986, N3088, N3315);
nor NOR3 (N13989, N13987, N8862, N275);
not NOT1 (N13990, N13988);
nand NAND3 (N13991, N13977, N13157, N4926);
xor XOR2 (N13992, N13973, N10573);
xor XOR2 (N13993, N13992, N10226);
or OR4 (N13994, N13982, N8988, N8627, N637);
and AND3 (N13995, N13991, N4422, N2537);
buf BUF1 (N13996, N13976);
buf BUF1 (N13997, N13993);
nor NOR2 (N13998, N13990, N1470);
not NOT1 (N13999, N13985);
buf BUF1 (N14000, N13989);
buf BUF1 (N14001, N14000);
xor XOR2 (N14002, N13978, N3352);
or OR3 (N14003, N13997, N13672, N3677);
nor NOR4 (N14004, N13996, N4971, N8805, N3208);
nor NOR4 (N14005, N14001, N12748, N7534, N13128);
buf BUF1 (N14006, N13995);
not NOT1 (N14007, N14002);
and AND4 (N14008, N13999, N508, N6925, N6535);
nor NOR2 (N14009, N14006, N8143);
xor XOR2 (N14010, N13969, N6856);
and AND3 (N14011, N13981, N2180, N12695);
not NOT1 (N14012, N13994);
not NOT1 (N14013, N14008);
and AND3 (N14014, N14011, N7047, N7605);
nor NOR2 (N14015, N14007, N7924);
and AND3 (N14016, N14009, N9693, N1421);
nand NAND3 (N14017, N14015, N4134, N8635);
xor XOR2 (N14018, N14003, N7136);
nor NOR3 (N14019, N14016, N12032, N7407);
or OR4 (N14020, N14012, N9401, N1337, N7638);
buf BUF1 (N14021, N14020);
nor NOR4 (N14022, N14019, N4093, N3270, N12910);
nand NAND2 (N14023, N14014, N2993);
not NOT1 (N14024, N14005);
buf BUF1 (N14025, N14018);
or OR2 (N14026, N14025, N6277);
and AND2 (N14027, N14021, N13784);
buf BUF1 (N14028, N14026);
xor XOR2 (N14029, N14013, N11669);
or OR4 (N14030, N14028, N6031, N4447, N5985);
or OR3 (N14031, N14029, N6124, N1274);
or OR3 (N14032, N14027, N1851, N1363);
nand NAND3 (N14033, N14017, N1157, N9130);
nand NAND2 (N14034, N14004, N13745);
nand NAND3 (N14035, N14023, N5267, N9769);
or OR3 (N14036, N14022, N2735, N4517);
xor XOR2 (N14037, N14034, N594);
xor XOR2 (N14038, N14024, N5957);
xor XOR2 (N14039, N14036, N11804);
not NOT1 (N14040, N14030);
nor NOR3 (N14041, N14035, N9882, N13125);
buf BUF1 (N14042, N14041);
nand NAND3 (N14043, N14010, N10787, N3351);
not NOT1 (N14044, N14039);
buf BUF1 (N14045, N14038);
buf BUF1 (N14046, N14037);
nor NOR2 (N14047, N14046, N9490);
and AND3 (N14048, N14044, N13795, N11139);
xor XOR2 (N14049, N14047, N3794);
buf BUF1 (N14050, N14033);
and AND2 (N14051, N14031, N13183);
nand NAND4 (N14052, N14049, N3751, N8124, N2078);
buf BUF1 (N14053, N14045);
buf BUF1 (N14054, N14032);
nor NOR3 (N14055, N14053, N7527, N13345);
and AND2 (N14056, N14043, N4748);
nand NAND3 (N14057, N14051, N12596, N8642);
nor NOR3 (N14058, N14057, N4635, N3917);
and AND3 (N14059, N14040, N9797, N12187);
xor XOR2 (N14060, N14050, N5214);
not NOT1 (N14061, N14060);
nor NOR4 (N14062, N14056, N11995, N9042, N10949);
buf BUF1 (N14063, N14048);
and AND2 (N14064, N14054, N5311);
buf BUF1 (N14065, N14063);
nand NAND4 (N14066, N14058, N12791, N5207, N8319);
or OR2 (N14067, N14065, N11247);
not NOT1 (N14068, N14055);
nor NOR3 (N14069, N14067, N8566, N2455);
nand NAND3 (N14070, N14062, N12231, N1433);
nor NOR3 (N14071, N14064, N13777, N8314);
nor NOR2 (N14072, N14071, N10605);
and AND2 (N14073, N14066, N7284);
or OR2 (N14074, N14061, N4184);
and AND2 (N14075, N14042, N12300);
nor NOR3 (N14076, N14059, N1877, N2354);
nand NAND2 (N14077, N14072, N9934);
nor NOR2 (N14078, N14076, N3415);
not NOT1 (N14079, N14075);
nor NOR3 (N14080, N14079, N5909, N8447);
nor NOR3 (N14081, N14069, N11560, N7296);
not NOT1 (N14082, N14070);
buf BUF1 (N14083, N13998);
buf BUF1 (N14084, N14052);
nor NOR4 (N14085, N14082, N11574, N9329, N9660);
or OR2 (N14086, N14081, N12741);
and AND3 (N14087, N14083, N13940, N5985);
and AND4 (N14088, N14087, N13190, N3385, N6511);
nand NAND2 (N14089, N14085, N4540);
not NOT1 (N14090, N14088);
not NOT1 (N14091, N14086);
or OR2 (N14092, N14078, N3308);
nand NAND4 (N14093, N14090, N5364, N7775, N4645);
and AND4 (N14094, N14080, N1016, N13017, N7265);
not NOT1 (N14095, N14074);
xor XOR2 (N14096, N14089, N10309);
nand NAND4 (N14097, N14073, N8015, N5182, N2098);
nand NAND3 (N14098, N14094, N11883, N10003);
and AND3 (N14099, N14098, N4245, N997);
or OR2 (N14100, N14096, N12348);
nand NAND4 (N14101, N14093, N176, N11761, N4961);
and AND4 (N14102, N14101, N5437, N6032, N11519);
nor NOR4 (N14103, N14077, N12258, N6824, N10713);
or OR3 (N14104, N14099, N924, N4511);
not NOT1 (N14105, N14103);
xor XOR2 (N14106, N14095, N3359);
not NOT1 (N14107, N14106);
or OR4 (N14108, N14100, N4151, N3102, N2838);
not NOT1 (N14109, N14097);
nand NAND2 (N14110, N14091, N6841);
and AND4 (N14111, N14068, N10333, N5890, N12152);
not NOT1 (N14112, N14092);
nand NAND2 (N14113, N14102, N3320);
and AND2 (N14114, N14109, N7951);
and AND4 (N14115, N14113, N13392, N5085, N4828);
and AND2 (N14116, N14112, N10390);
nand NAND2 (N14117, N14115, N12315);
buf BUF1 (N14118, N14104);
xor XOR2 (N14119, N14110, N1372);
nand NAND2 (N14120, N14084, N2727);
or OR3 (N14121, N14120, N9913, N2005);
or OR2 (N14122, N14108, N9142);
xor XOR2 (N14123, N14122, N9632);
nor NOR3 (N14124, N14116, N7922, N2396);
buf BUF1 (N14125, N14117);
nor NOR2 (N14126, N14118, N7778);
buf BUF1 (N14127, N14107);
nand NAND2 (N14128, N14119, N5032);
nor NOR2 (N14129, N14128, N1299);
and AND3 (N14130, N14129, N7606, N12229);
or OR2 (N14131, N14114, N9426);
and AND2 (N14132, N14124, N12697);
nand NAND3 (N14133, N14125, N3712, N10326);
and AND3 (N14134, N14123, N1498, N10143);
and AND4 (N14135, N14105, N4169, N11399, N7750);
buf BUF1 (N14136, N14127);
nor NOR4 (N14137, N14135, N8912, N6357, N3486);
buf BUF1 (N14138, N14121);
nand NAND2 (N14139, N14111, N8605);
xor XOR2 (N14140, N14137, N6146);
xor XOR2 (N14141, N14132, N5692);
nor NOR4 (N14142, N14140, N4765, N13588, N13691);
or OR3 (N14143, N14139, N6906, N10452);
nand NAND2 (N14144, N14126, N6280);
and AND4 (N14145, N14142, N6289, N4903, N5235);
buf BUF1 (N14146, N14143);
and AND2 (N14147, N14138, N3392);
or OR2 (N14148, N14145, N1068);
buf BUF1 (N14149, N14134);
or OR4 (N14150, N14149, N9646, N493, N3877);
and AND2 (N14151, N14147, N11968);
nor NOR2 (N14152, N14146, N2574);
nor NOR4 (N14153, N14148, N5990, N9773, N4979);
buf BUF1 (N14154, N14136);
xor XOR2 (N14155, N14144, N1115);
nand NAND4 (N14156, N14153, N6326, N45, N9864);
xor XOR2 (N14157, N14155, N9847);
nand NAND3 (N14158, N14151, N2133, N2301);
nor NOR2 (N14159, N14141, N10300);
not NOT1 (N14160, N14159);
xor XOR2 (N14161, N14160, N10390);
not NOT1 (N14162, N14130);
buf BUF1 (N14163, N14131);
nor NOR3 (N14164, N14157, N7134, N11641);
and AND2 (N14165, N14158, N9968);
nor NOR4 (N14166, N14150, N11166, N657, N1776);
nor NOR2 (N14167, N14166, N13950);
or OR3 (N14168, N14161, N7050, N7063);
nor NOR4 (N14169, N14154, N12255, N5253, N2926);
or OR2 (N14170, N14162, N9064);
nor NOR4 (N14171, N14167, N5635, N212, N7879);
nand NAND4 (N14172, N14152, N601, N6984, N10234);
xor XOR2 (N14173, N14165, N12571);
buf BUF1 (N14174, N14163);
nand NAND2 (N14175, N14156, N2622);
xor XOR2 (N14176, N14173, N13989);
nor NOR2 (N14177, N14175, N12897);
xor XOR2 (N14178, N14176, N3013);
not NOT1 (N14179, N14133);
or OR4 (N14180, N14174, N3715, N9163, N4945);
or OR3 (N14181, N14177, N3959, N11771);
not NOT1 (N14182, N14178);
nor NOR2 (N14183, N14180, N13234);
or OR3 (N14184, N14179, N12235, N6539);
not NOT1 (N14185, N14171);
xor XOR2 (N14186, N14172, N8603);
xor XOR2 (N14187, N14164, N1753);
nand NAND2 (N14188, N14182, N500);
not NOT1 (N14189, N14183);
xor XOR2 (N14190, N14169, N888);
not NOT1 (N14191, N14181);
or OR4 (N14192, N14185, N7750, N2408, N3477);
or OR3 (N14193, N14188, N10756, N12522);
not NOT1 (N14194, N14170);
buf BUF1 (N14195, N14192);
or OR3 (N14196, N14190, N7533, N12898);
and AND3 (N14197, N14195, N1560, N3203);
xor XOR2 (N14198, N14184, N10190);
and AND3 (N14199, N14194, N6414, N386);
not NOT1 (N14200, N14187);
or OR3 (N14201, N14197, N1843, N11218);
and AND3 (N14202, N14201, N13556, N11428);
nor NOR2 (N14203, N14200, N10038);
and AND3 (N14204, N14186, N9607, N8824);
nor NOR3 (N14205, N14202, N13724, N498);
nor NOR4 (N14206, N14198, N10858, N1456, N2198);
buf BUF1 (N14207, N14206);
nand NAND4 (N14208, N14203, N5349, N12676, N5962);
nor NOR3 (N14209, N14205, N4924, N4000);
xor XOR2 (N14210, N14189, N12856);
and AND4 (N14211, N14209, N3123, N8474, N13742);
xor XOR2 (N14212, N14208, N11931);
or OR4 (N14213, N14193, N6115, N13805, N13817);
buf BUF1 (N14214, N14199);
xor XOR2 (N14215, N14196, N1602);
not NOT1 (N14216, N14191);
buf BUF1 (N14217, N14210);
buf BUF1 (N14218, N14211);
buf BUF1 (N14219, N14217);
and AND2 (N14220, N14212, N8368);
buf BUF1 (N14221, N14219);
xor XOR2 (N14222, N14220, N4811);
nand NAND3 (N14223, N14218, N12365, N8533);
and AND3 (N14224, N14214, N8968, N2392);
buf BUF1 (N14225, N14222);
and AND2 (N14226, N14223, N7329);
xor XOR2 (N14227, N14168, N4285);
nor NOR2 (N14228, N14204, N5476);
xor XOR2 (N14229, N14228, N13000);
xor XOR2 (N14230, N14215, N11233);
buf BUF1 (N14231, N14224);
nand NAND3 (N14232, N14213, N6698, N1068);
not NOT1 (N14233, N14221);
and AND3 (N14234, N14233, N7760, N13633);
nor NOR4 (N14235, N14232, N8070, N1757, N8856);
and AND3 (N14236, N14225, N13114, N6570);
nor NOR4 (N14237, N14226, N3171, N2639, N13097);
or OR3 (N14238, N14207, N8446, N1118);
nor NOR3 (N14239, N14238, N4982, N13248);
nand NAND2 (N14240, N14236, N574);
xor XOR2 (N14241, N14227, N11390);
nor NOR4 (N14242, N14237, N5865, N6392, N13324);
nor NOR2 (N14243, N14241, N11573);
xor XOR2 (N14244, N14242, N5230);
buf BUF1 (N14245, N14235);
nand NAND3 (N14246, N14216, N7921, N14175);
or OR3 (N14247, N14239, N2089, N9852);
or OR3 (N14248, N14246, N3826, N5341);
nand NAND3 (N14249, N14229, N10827, N1625);
xor XOR2 (N14250, N14248, N7655);
not NOT1 (N14251, N14245);
nor NOR2 (N14252, N14243, N13849);
nor NOR4 (N14253, N14249, N3146, N6389, N5294);
xor XOR2 (N14254, N14252, N2812);
nand NAND3 (N14255, N14234, N13068, N5010);
nand NAND2 (N14256, N14240, N3045);
or OR2 (N14257, N14251, N13313);
buf BUF1 (N14258, N14250);
or OR3 (N14259, N14253, N3841, N11139);
xor XOR2 (N14260, N14247, N2644);
or OR2 (N14261, N14230, N11174);
and AND3 (N14262, N14256, N3429, N2966);
nand NAND4 (N14263, N14231, N2301, N11723, N6697);
or OR2 (N14264, N14259, N11205);
nand NAND4 (N14265, N14260, N2803, N9733, N9538);
buf BUF1 (N14266, N14257);
or OR4 (N14267, N14265, N12129, N13308, N6583);
xor XOR2 (N14268, N14255, N7260);
xor XOR2 (N14269, N14264, N646);
and AND2 (N14270, N14269, N1216);
xor XOR2 (N14271, N14258, N12199);
or OR4 (N14272, N14266, N8328, N44, N7993);
not NOT1 (N14273, N14263);
nor NOR2 (N14274, N14270, N10708);
nand NAND4 (N14275, N14271, N6272, N13877, N4449);
buf BUF1 (N14276, N14272);
nand NAND2 (N14277, N14261, N7568);
buf BUF1 (N14278, N14274);
xor XOR2 (N14279, N14268, N2441);
and AND3 (N14280, N14244, N10114, N244);
buf BUF1 (N14281, N14280);
and AND3 (N14282, N14254, N4180, N323);
and AND4 (N14283, N14273, N10593, N12183, N2273);
nor NOR4 (N14284, N14282, N2611, N13680, N7177);
xor XOR2 (N14285, N14267, N7924);
nor NOR4 (N14286, N14275, N7213, N1968, N12811);
or OR2 (N14287, N14277, N8954);
nor NOR4 (N14288, N14286, N5010, N6590, N9206);
or OR4 (N14289, N14287, N637, N6648, N11145);
not NOT1 (N14290, N14276);
xor XOR2 (N14291, N14262, N1589);
buf BUF1 (N14292, N14285);
not NOT1 (N14293, N14278);
nor NOR4 (N14294, N14281, N9769, N14006, N10463);
xor XOR2 (N14295, N14294, N5822);
and AND3 (N14296, N14292, N7084, N9660);
nor NOR3 (N14297, N14279, N8644, N5325);
buf BUF1 (N14298, N14288);
and AND3 (N14299, N14291, N11934, N13570);
nor NOR2 (N14300, N14298, N9282);
nand NAND4 (N14301, N14290, N12294, N6798, N4115);
or OR2 (N14302, N14300, N12445);
and AND3 (N14303, N14283, N5075, N5142);
nor NOR4 (N14304, N14296, N5690, N11612, N2977);
and AND2 (N14305, N14301, N3639);
buf BUF1 (N14306, N14284);
xor XOR2 (N14307, N14304, N7227);
nor NOR4 (N14308, N14303, N9872, N4765, N13631);
or OR4 (N14309, N14293, N3742, N4318, N9952);
not NOT1 (N14310, N14295);
and AND2 (N14311, N14297, N14190);
xor XOR2 (N14312, N14302, N5249);
not NOT1 (N14313, N14312);
xor XOR2 (N14314, N14289, N13826);
xor XOR2 (N14315, N14310, N11244);
and AND4 (N14316, N14309, N6065, N7832, N8589);
nor NOR4 (N14317, N14313, N7983, N9078, N1187);
or OR2 (N14318, N14314, N13651);
nand NAND3 (N14319, N14299, N9933, N9026);
buf BUF1 (N14320, N14308);
or OR4 (N14321, N14311, N6585, N4800, N2588);
not NOT1 (N14322, N14305);
or OR4 (N14323, N14316, N3110, N4915, N13544);
nand NAND3 (N14324, N14321, N12344, N4960);
and AND4 (N14325, N14307, N466, N7867, N12960);
nand NAND3 (N14326, N14317, N5319, N356);
not NOT1 (N14327, N14306);
nand NAND2 (N14328, N14319, N11502);
nor NOR4 (N14329, N14327, N11172, N11204, N7583);
nand NAND4 (N14330, N14324, N1893, N5827, N6359);
or OR2 (N14331, N14328, N2141);
buf BUF1 (N14332, N14325);
nand NAND3 (N14333, N14326, N7129, N1001);
or OR2 (N14334, N14318, N10514);
buf BUF1 (N14335, N14333);
buf BUF1 (N14336, N14335);
buf BUF1 (N14337, N14336);
buf BUF1 (N14338, N14330);
buf BUF1 (N14339, N14332);
and AND2 (N14340, N14334, N13964);
buf BUF1 (N14341, N14340);
and AND4 (N14342, N14322, N6581, N9566, N2415);
nor NOR4 (N14343, N14331, N7801, N9308, N4088);
nand NAND2 (N14344, N14339, N12153);
not NOT1 (N14345, N14343);
buf BUF1 (N14346, N14337);
not NOT1 (N14347, N14341);
not NOT1 (N14348, N14347);
nand NAND3 (N14349, N14338, N11113, N8775);
buf BUF1 (N14350, N14349);
and AND2 (N14351, N14342, N12184);
xor XOR2 (N14352, N14351, N6830);
and AND2 (N14353, N14346, N6360);
xor XOR2 (N14354, N14315, N1234);
buf BUF1 (N14355, N14354);
not NOT1 (N14356, N14348);
and AND4 (N14357, N14345, N12293, N1472, N8022);
and AND4 (N14358, N14357, N7149, N1605, N12967);
xor XOR2 (N14359, N14353, N11005);
nand NAND3 (N14360, N14356, N4482, N7308);
or OR2 (N14361, N14344, N834);
xor XOR2 (N14362, N14358, N11521);
and AND4 (N14363, N14323, N671, N4747, N10695);
nand NAND2 (N14364, N14355, N4702);
and AND2 (N14365, N14363, N6679);
nor NOR3 (N14366, N14350, N13804, N12347);
buf BUF1 (N14367, N14320);
not NOT1 (N14368, N14367);
buf BUF1 (N14369, N14329);
buf BUF1 (N14370, N14359);
nand NAND4 (N14371, N14352, N2742, N373, N4996);
nand NAND2 (N14372, N14369, N3826);
or OR3 (N14373, N14366, N13969, N2782);
buf BUF1 (N14374, N14360);
and AND3 (N14375, N14362, N381, N4792);
and AND3 (N14376, N14373, N6353, N9572);
buf BUF1 (N14377, N14376);
not NOT1 (N14378, N14361);
nand NAND3 (N14379, N14378, N5752, N182);
not NOT1 (N14380, N14368);
nand NAND2 (N14381, N14379, N5279);
and AND2 (N14382, N14374, N10742);
xor XOR2 (N14383, N14377, N9158);
buf BUF1 (N14384, N14375);
xor XOR2 (N14385, N14371, N12979);
or OR4 (N14386, N14383, N9112, N12379, N3180);
and AND2 (N14387, N14364, N11575);
xor XOR2 (N14388, N14387, N556);
xor XOR2 (N14389, N14372, N7069);
buf BUF1 (N14390, N14389);
and AND2 (N14391, N14384, N12021);
buf BUF1 (N14392, N14385);
not NOT1 (N14393, N14391);
not NOT1 (N14394, N14386);
not NOT1 (N14395, N14365);
and AND3 (N14396, N14393, N9448, N13257);
nand NAND2 (N14397, N14370, N1577);
not NOT1 (N14398, N14392);
not NOT1 (N14399, N14390);
or OR2 (N14400, N14388, N10872);
nand NAND4 (N14401, N14399, N11872, N13509, N5994);
or OR3 (N14402, N14395, N11708, N11229);
or OR2 (N14403, N14394, N11618);
nor NOR3 (N14404, N14401, N1261, N10399);
or OR4 (N14405, N14380, N7607, N13591, N1405);
not NOT1 (N14406, N14382);
nand NAND3 (N14407, N14396, N6559, N11155);
nand NAND3 (N14408, N14397, N1498, N12588);
xor XOR2 (N14409, N14400, N7512);
nand NAND3 (N14410, N14407, N8703, N7192);
nand NAND3 (N14411, N14402, N7322, N9228);
not NOT1 (N14412, N14410);
buf BUF1 (N14413, N14409);
nor NOR3 (N14414, N14412, N8513, N13180);
nor NOR3 (N14415, N14413, N8263, N1857);
buf BUF1 (N14416, N14398);
or OR3 (N14417, N14411, N853, N2291);
nor NOR4 (N14418, N14405, N11734, N3989, N7589);
xor XOR2 (N14419, N14414, N5184);
xor XOR2 (N14420, N14419, N5849);
and AND3 (N14421, N14416, N6538, N8591);
buf BUF1 (N14422, N14420);
buf BUF1 (N14423, N14403);
xor XOR2 (N14424, N14406, N6594);
or OR4 (N14425, N14381, N12857, N3307, N3078);
or OR4 (N14426, N14424, N6734, N1924, N2464);
and AND4 (N14427, N14425, N1963, N13597, N5606);
xor XOR2 (N14428, N14426, N109);
not NOT1 (N14429, N14422);
not NOT1 (N14430, N14421);
and AND4 (N14431, N14415, N9648, N1329, N8843);
xor XOR2 (N14432, N14423, N14317);
nor NOR4 (N14433, N14404, N8714, N13693, N1709);
nor NOR3 (N14434, N14431, N12183, N2860);
or OR3 (N14435, N14408, N9402, N13579);
buf BUF1 (N14436, N14428);
nand NAND3 (N14437, N14430, N9966, N10896);
xor XOR2 (N14438, N14435, N2344);
nor NOR3 (N14439, N14437, N5322, N12);
or OR4 (N14440, N14427, N3638, N12792, N7962);
nor NOR3 (N14441, N14440, N8544, N7464);
and AND4 (N14442, N14432, N5178, N6653, N3489);
and AND3 (N14443, N14441, N6306, N2041);
and AND2 (N14444, N14433, N2116);
nand NAND2 (N14445, N14443, N5472);
and AND4 (N14446, N14417, N4730, N8411, N7319);
xor XOR2 (N14447, N14442, N6206);
and AND3 (N14448, N14446, N2914, N6743);
nand NAND3 (N14449, N14445, N9167, N3835);
nand NAND2 (N14450, N14439, N11554);
nor NOR2 (N14451, N14438, N7512);
not NOT1 (N14452, N14449);
xor XOR2 (N14453, N14429, N2714);
nand NAND4 (N14454, N14452, N11314, N9869, N13523);
or OR2 (N14455, N14447, N648);
not NOT1 (N14456, N14418);
not NOT1 (N14457, N14448);
xor XOR2 (N14458, N14444, N2811);
and AND3 (N14459, N14451, N11061, N1024);
nor NOR2 (N14460, N14434, N2478);
xor XOR2 (N14461, N14436, N130);
xor XOR2 (N14462, N14457, N3320);
and AND4 (N14463, N14454, N7019, N3055, N12750);
nor NOR2 (N14464, N14450, N2312);
buf BUF1 (N14465, N14462);
nand NAND2 (N14466, N14465, N12881);
xor XOR2 (N14467, N14461, N161);
nand NAND3 (N14468, N14459, N12823, N11869);
nand NAND4 (N14469, N14463, N8853, N5564, N4293);
or OR2 (N14470, N14467, N1811);
buf BUF1 (N14471, N14453);
buf BUF1 (N14472, N14466);
xor XOR2 (N14473, N14455, N4543);
xor XOR2 (N14474, N14469, N13882);
and AND4 (N14475, N14456, N12623, N14313, N10855);
and AND4 (N14476, N14475, N3659, N12570, N10135);
buf BUF1 (N14477, N14472);
or OR4 (N14478, N14464, N641, N558, N459);
not NOT1 (N14479, N14477);
or OR4 (N14480, N14458, N363, N11064, N13692);
not NOT1 (N14481, N14476);
nor NOR4 (N14482, N14480, N14420, N8940, N9657);
buf BUF1 (N14483, N14482);
and AND4 (N14484, N14478, N13572, N3200, N13893);
and AND2 (N14485, N14471, N11990);
xor XOR2 (N14486, N14468, N7329);
xor XOR2 (N14487, N14483, N8148);
not NOT1 (N14488, N14485);
or OR4 (N14489, N14479, N390, N1849, N7420);
and AND3 (N14490, N14487, N3831, N4936);
nand NAND3 (N14491, N14484, N13591, N3692);
or OR4 (N14492, N14490, N27, N4877, N1644);
not NOT1 (N14493, N14473);
nand NAND3 (N14494, N14486, N11795, N2367);
nor NOR3 (N14495, N14460, N7830, N6974);
nor NOR3 (N14496, N14491, N3973, N2062);
xor XOR2 (N14497, N14495, N3823);
or OR2 (N14498, N14493, N10366);
not NOT1 (N14499, N14497);
or OR2 (N14500, N14489, N8987);
not NOT1 (N14501, N14500);
not NOT1 (N14502, N14494);
or OR2 (N14503, N14499, N11145);
xor XOR2 (N14504, N14474, N3630);
not NOT1 (N14505, N14488);
xor XOR2 (N14506, N14503, N7382);
and AND3 (N14507, N14470, N14350, N12165);
nor NOR2 (N14508, N14505, N13957);
xor XOR2 (N14509, N14496, N2554);
nand NAND4 (N14510, N14509, N13446, N4958, N4653);
or OR3 (N14511, N14508, N1376, N2744);
buf BUF1 (N14512, N14510);
and AND3 (N14513, N14481, N5266, N2738);
nand NAND4 (N14514, N14506, N7689, N2733, N12499);
or OR2 (N14515, N14504, N11658);
and AND2 (N14516, N14515, N14276);
xor XOR2 (N14517, N14498, N12862);
buf BUF1 (N14518, N14502);
or OR3 (N14519, N14514, N10516, N11706);
and AND3 (N14520, N14519, N4565, N13218);
nand NAND4 (N14521, N14507, N14125, N8191, N2552);
not NOT1 (N14522, N14520);
or OR3 (N14523, N14512, N13813, N11759);
nor NOR2 (N14524, N14521, N2221);
or OR2 (N14525, N14524, N8486);
nor NOR4 (N14526, N14518, N4472, N5401, N10421);
buf BUF1 (N14527, N14526);
nor NOR4 (N14528, N14511, N10532, N9772, N6258);
or OR4 (N14529, N14513, N9832, N10264, N9284);
nor NOR3 (N14530, N14527, N510, N2483);
buf BUF1 (N14531, N14522);
nand NAND2 (N14532, N14516, N6700);
nand NAND4 (N14533, N14492, N5776, N13100, N2296);
not NOT1 (N14534, N14529);
xor XOR2 (N14535, N14528, N8903);
nor NOR4 (N14536, N14501, N2326, N10487, N322);
nand NAND2 (N14537, N14532, N5506);
nand NAND3 (N14538, N14534, N6713, N8696);
not NOT1 (N14539, N14536);
and AND4 (N14540, N14535, N3590, N13176, N11799);
or OR3 (N14541, N14540, N915, N2510);
or OR4 (N14542, N14541, N11585, N8785, N1627);
or OR2 (N14543, N14517, N6091);
xor XOR2 (N14544, N14531, N13568);
nor NOR3 (N14545, N14530, N13960, N8246);
or OR4 (N14546, N14545, N6383, N8183, N10263);
or OR3 (N14547, N14537, N8473, N13730);
and AND4 (N14548, N14525, N8731, N1580, N12209);
nand NAND2 (N14549, N14533, N9815);
or OR3 (N14550, N14538, N6349, N559);
and AND3 (N14551, N14539, N1152, N9971);
or OR4 (N14552, N14551, N2559, N868, N11871);
nand NAND2 (N14553, N14547, N7887);
not NOT1 (N14554, N14553);
and AND2 (N14555, N14552, N4469);
nand NAND2 (N14556, N14542, N9131);
not NOT1 (N14557, N14544);
nor NOR2 (N14558, N14556, N119);
buf BUF1 (N14559, N14550);
not NOT1 (N14560, N14549);
xor XOR2 (N14561, N14546, N2017);
and AND2 (N14562, N14561, N6518);
nand NAND3 (N14563, N14548, N4300, N9174);
nor NOR2 (N14564, N14554, N3635);
nand NAND3 (N14565, N14559, N6138, N4921);
buf BUF1 (N14566, N14557);
and AND3 (N14567, N14558, N7533, N2752);
buf BUF1 (N14568, N14523);
or OR3 (N14569, N14543, N4931, N7282);
nor NOR3 (N14570, N14555, N3243, N1009);
or OR3 (N14571, N14567, N1556, N2632);
xor XOR2 (N14572, N14566, N14403);
not NOT1 (N14573, N14568);
not NOT1 (N14574, N14565);
not NOT1 (N14575, N14569);
nor NOR4 (N14576, N14563, N1171, N9391, N4115);
and AND3 (N14577, N14560, N1504, N12570);
buf BUF1 (N14578, N14562);
xor XOR2 (N14579, N14564, N11063);
or OR2 (N14580, N14574, N6552);
and AND3 (N14581, N14570, N2895, N6361);
and AND2 (N14582, N14571, N2002);
nor NOR4 (N14583, N14575, N13733, N3472, N1975);
not NOT1 (N14584, N14580);
or OR2 (N14585, N14576, N11370);
nor NOR2 (N14586, N14579, N14442);
and AND2 (N14587, N14583, N6394);
buf BUF1 (N14588, N14587);
nor NOR2 (N14589, N14582, N10078);
not NOT1 (N14590, N14573);
xor XOR2 (N14591, N14584, N1226);
nand NAND2 (N14592, N14590, N13306);
and AND2 (N14593, N14591, N8623);
or OR4 (N14594, N14593, N14265, N6577, N14462);
xor XOR2 (N14595, N14588, N9227);
or OR3 (N14596, N14585, N9440, N754);
and AND4 (N14597, N14577, N7735, N6293, N11802);
not NOT1 (N14598, N14586);
or OR4 (N14599, N14572, N819, N5182, N3712);
not NOT1 (N14600, N14598);
buf BUF1 (N14601, N14600);
or OR4 (N14602, N14592, N8529, N3131, N9455);
nand NAND4 (N14603, N14578, N1088, N10812, N4983);
not NOT1 (N14604, N14595);
not NOT1 (N14605, N14602);
buf BUF1 (N14606, N14604);
nand NAND2 (N14607, N14597, N4940);
or OR4 (N14608, N14594, N20, N11603, N2059);
xor XOR2 (N14609, N14603, N8262);
and AND3 (N14610, N14589, N9088, N3884);
or OR3 (N14611, N14605, N5676, N14321);
nor NOR3 (N14612, N14596, N7383, N456);
nand NAND4 (N14613, N14609, N4548, N9022, N9232);
xor XOR2 (N14614, N14606, N8939);
not NOT1 (N14615, N14613);
buf BUF1 (N14616, N14608);
and AND4 (N14617, N14615, N8738, N6478, N4130);
buf BUF1 (N14618, N14607);
not NOT1 (N14619, N14618);
not NOT1 (N14620, N14581);
not NOT1 (N14621, N14610);
buf BUF1 (N14622, N14617);
and AND4 (N14623, N14611, N12325, N9803, N771);
or OR2 (N14624, N14599, N9740);
buf BUF1 (N14625, N14623);
buf BUF1 (N14626, N14612);
or OR2 (N14627, N14625, N8791);
buf BUF1 (N14628, N14620);
xor XOR2 (N14629, N14622, N9902);
nor NOR3 (N14630, N14629, N6300, N531);
nor NOR3 (N14631, N14630, N14505, N6120);
nor NOR4 (N14632, N14616, N9248, N1308, N1374);
xor XOR2 (N14633, N14628, N9352);
and AND4 (N14634, N14632, N14547, N2621, N9514);
not NOT1 (N14635, N14633);
and AND4 (N14636, N14624, N6086, N4126, N1122);
or OR2 (N14637, N14635, N8191);
or OR4 (N14638, N14619, N4494, N4111, N9018);
buf BUF1 (N14639, N14626);
buf BUF1 (N14640, N14631);
buf BUF1 (N14641, N14638);
buf BUF1 (N14642, N14634);
and AND3 (N14643, N14642, N13603, N11344);
not NOT1 (N14644, N14637);
xor XOR2 (N14645, N14601, N12824);
nor NOR2 (N14646, N14639, N7679);
xor XOR2 (N14647, N14641, N1701);
buf BUF1 (N14648, N14621);
and AND4 (N14649, N14640, N3361, N2272, N3349);
and AND4 (N14650, N14643, N7310, N5577, N4247);
xor XOR2 (N14651, N14648, N11210);
and AND2 (N14652, N14650, N12949);
or OR4 (N14653, N14652, N6325, N12181, N12756);
buf BUF1 (N14654, N14653);
buf BUF1 (N14655, N14645);
xor XOR2 (N14656, N14644, N3036);
buf BUF1 (N14657, N14655);
nand NAND4 (N14658, N14649, N6426, N4380, N13692);
nor NOR3 (N14659, N14627, N14261, N6646);
nand NAND4 (N14660, N14636, N9584, N8777, N2251);
xor XOR2 (N14661, N14658, N7689);
not NOT1 (N14662, N14656);
not NOT1 (N14663, N14651);
nand NAND3 (N14664, N14661, N7489, N11215);
nand NAND4 (N14665, N14614, N12458, N1826, N13373);
not NOT1 (N14666, N14654);
not NOT1 (N14667, N14646);
or OR4 (N14668, N14667, N213, N7834, N5508);
buf BUF1 (N14669, N14660);
not NOT1 (N14670, N14659);
nor NOR4 (N14671, N14668, N14597, N9753, N13754);
nand NAND2 (N14672, N14671, N11417);
buf BUF1 (N14673, N14647);
and AND2 (N14674, N14657, N365);
xor XOR2 (N14675, N14665, N10793);
or OR4 (N14676, N14664, N10240, N4857, N9988);
not NOT1 (N14677, N14675);
not NOT1 (N14678, N14674);
not NOT1 (N14679, N14662);
nand NAND2 (N14680, N14679, N5165);
nor NOR2 (N14681, N14672, N6358);
nand NAND2 (N14682, N14676, N9898);
buf BUF1 (N14683, N14677);
nor NOR4 (N14684, N14682, N3695, N1798, N11501);
or OR4 (N14685, N14670, N14226, N7920, N2803);
and AND4 (N14686, N14680, N10493, N14311, N11379);
nand NAND3 (N14687, N14666, N12770, N11305);
not NOT1 (N14688, N14669);
xor XOR2 (N14689, N14678, N2828);
or OR2 (N14690, N14663, N8033);
or OR2 (N14691, N14689, N10819);
nor NOR2 (N14692, N14687, N14612);
nor NOR2 (N14693, N14685, N6644);
not NOT1 (N14694, N14688);
and AND2 (N14695, N14694, N7745);
nor NOR4 (N14696, N14686, N1131, N4679, N14008);
or OR2 (N14697, N14683, N9454);
and AND4 (N14698, N14697, N1270, N516, N3691);
or OR4 (N14699, N14698, N9676, N9202, N60);
nand NAND3 (N14700, N14692, N7185, N13562);
or OR2 (N14701, N14691, N915);
nor NOR3 (N14702, N14673, N6235, N2520);
not NOT1 (N14703, N14693);
nor NOR4 (N14704, N14702, N9454, N8371, N3273);
not NOT1 (N14705, N14704);
buf BUF1 (N14706, N14696);
or OR2 (N14707, N14705, N7756);
nand NAND4 (N14708, N14701, N13939, N11184, N12329);
nand NAND3 (N14709, N14707, N384, N10245);
and AND4 (N14710, N14690, N9037, N11427, N5621);
not NOT1 (N14711, N14709);
nor NOR4 (N14712, N14706, N2717, N1951, N2967);
not NOT1 (N14713, N14711);
or OR2 (N14714, N14708, N578);
or OR2 (N14715, N14684, N10109);
and AND4 (N14716, N14700, N578, N14476, N11802);
not NOT1 (N14717, N14716);
or OR4 (N14718, N14710, N12200, N13641, N5085);
buf BUF1 (N14719, N14712);
not NOT1 (N14720, N14713);
and AND3 (N14721, N14719, N10307, N727);
and AND2 (N14722, N14720, N11576);
or OR4 (N14723, N14714, N4297, N9452, N5586);
xor XOR2 (N14724, N14723, N5146);
not NOT1 (N14725, N14722);
or OR3 (N14726, N14725, N12178, N13987);
nand NAND3 (N14727, N14721, N13133, N5580);
not NOT1 (N14728, N14699);
nor NOR3 (N14729, N14681, N9720, N4534);
not NOT1 (N14730, N14726);
nand NAND4 (N14731, N14728, N5483, N13652, N4090);
nor NOR2 (N14732, N14717, N6995);
xor XOR2 (N14733, N14703, N9822);
nand NAND3 (N14734, N14733, N8378, N1226);
nor NOR4 (N14735, N14695, N5735, N8009, N1431);
not NOT1 (N14736, N14718);
nor NOR2 (N14737, N14734, N10035);
and AND4 (N14738, N14715, N13499, N12599, N14271);
and AND3 (N14739, N14730, N4713, N14408);
and AND3 (N14740, N14731, N14187, N8571);
xor XOR2 (N14741, N14732, N8801);
and AND2 (N14742, N14736, N14398);
or OR3 (N14743, N14737, N10393, N13533);
buf BUF1 (N14744, N14724);
nand NAND3 (N14745, N14735, N3216, N1006);
or OR2 (N14746, N14744, N3761);
buf BUF1 (N14747, N14727);
nand NAND2 (N14748, N14747, N7766);
or OR2 (N14749, N14729, N5919);
buf BUF1 (N14750, N14745);
xor XOR2 (N14751, N14750, N14588);
not NOT1 (N14752, N14739);
xor XOR2 (N14753, N14740, N10721);
nor NOR4 (N14754, N14742, N3913, N6875, N10577);
buf BUF1 (N14755, N14743);
nand NAND3 (N14756, N14738, N4295, N10437);
xor XOR2 (N14757, N14755, N9021);
nor NOR4 (N14758, N14752, N6824, N11664, N8027);
or OR4 (N14759, N14746, N11809, N4197, N5080);
nor NOR2 (N14760, N14741, N4697);
nor NOR3 (N14761, N14760, N4226, N11422);
xor XOR2 (N14762, N14758, N11550);
buf BUF1 (N14763, N14751);
not NOT1 (N14764, N14754);
buf BUF1 (N14765, N14753);
nor NOR3 (N14766, N14762, N7237, N9536);
nor NOR2 (N14767, N14759, N9820);
nand NAND2 (N14768, N14761, N4313);
not NOT1 (N14769, N14748);
not NOT1 (N14770, N14764);
xor XOR2 (N14771, N14768, N8458);
or OR3 (N14772, N14767, N2867, N7529);
nand NAND4 (N14773, N14771, N8850, N9459, N12633);
nor NOR2 (N14774, N14773, N518);
and AND3 (N14775, N14770, N8099, N13780);
buf BUF1 (N14776, N14765);
nand NAND3 (N14777, N14766, N6081, N13326);
xor XOR2 (N14778, N14772, N11640);
or OR2 (N14779, N14757, N11775);
nor NOR2 (N14780, N14777, N3069);
xor XOR2 (N14781, N14756, N5429);
xor XOR2 (N14782, N14778, N534);
buf BUF1 (N14783, N14780);
not NOT1 (N14784, N14775);
or OR4 (N14785, N14784, N11580, N1398, N10239);
and AND2 (N14786, N14774, N7132);
not NOT1 (N14787, N14781);
xor XOR2 (N14788, N14769, N4448);
not NOT1 (N14789, N14787);
or OR2 (N14790, N14789, N3491);
nand NAND3 (N14791, N14788, N2256, N12797);
nor NOR4 (N14792, N14763, N13055, N2127, N5502);
nand NAND3 (N14793, N14776, N11524, N593);
or OR2 (N14794, N14792, N1478);
xor XOR2 (N14795, N14794, N11256);
and AND2 (N14796, N14785, N1848);
buf BUF1 (N14797, N14795);
nor NOR4 (N14798, N14782, N4894, N7576, N4149);
xor XOR2 (N14799, N14783, N9536);
and AND3 (N14800, N14791, N13896, N2645);
not NOT1 (N14801, N14793);
buf BUF1 (N14802, N14779);
nand NAND4 (N14803, N14797, N7638, N9946, N12161);
xor XOR2 (N14804, N14796, N190);
nor NOR3 (N14805, N14801, N8444, N9705);
nand NAND4 (N14806, N14786, N8423, N7108, N7748);
not NOT1 (N14807, N14803);
buf BUF1 (N14808, N14798);
or OR4 (N14809, N14805, N7277, N9, N6403);
xor XOR2 (N14810, N14802, N4308);
buf BUF1 (N14811, N14807);
nor NOR2 (N14812, N14806, N10995);
nand NAND3 (N14813, N14804, N12840, N14809);
xor XOR2 (N14814, N2053, N3302);
nor NOR4 (N14815, N14814, N1652, N3566, N12438);
and AND4 (N14816, N14810, N203, N2638, N1760);
not NOT1 (N14817, N14813);
and AND3 (N14818, N14815, N13309, N1699);
nand NAND4 (N14819, N14790, N10101, N8053, N4758);
nor NOR4 (N14820, N14811, N2033, N5838, N1976);
buf BUF1 (N14821, N14817);
xor XOR2 (N14822, N14819, N8150);
buf BUF1 (N14823, N14818);
xor XOR2 (N14824, N14808, N726);
and AND3 (N14825, N14822, N12355, N2455);
not NOT1 (N14826, N14823);
nor NOR2 (N14827, N14820, N4382);
nand NAND4 (N14828, N14825, N8865, N5112, N11231);
xor XOR2 (N14829, N14826, N10580);
nor NOR4 (N14830, N14799, N14174, N11352, N9383);
or OR2 (N14831, N14800, N13365);
and AND2 (N14832, N14828, N10572);
and AND4 (N14833, N14827, N8828, N4098, N598);
nand NAND3 (N14834, N14832, N2203, N814);
not NOT1 (N14835, N14824);
xor XOR2 (N14836, N14821, N6925);
buf BUF1 (N14837, N14831);
buf BUF1 (N14838, N14812);
or OR3 (N14839, N14838, N6588, N4109);
and AND4 (N14840, N14834, N12389, N571, N10027);
xor XOR2 (N14841, N14840, N524);
and AND3 (N14842, N14835, N3574, N3430);
not NOT1 (N14843, N14837);
not NOT1 (N14844, N14829);
or OR3 (N14845, N14843, N12028, N9397);
xor XOR2 (N14846, N14836, N13879);
not NOT1 (N14847, N14841);
not NOT1 (N14848, N14816);
and AND4 (N14849, N14749, N1965, N10605, N11680);
nand NAND2 (N14850, N14846, N5133);
not NOT1 (N14851, N14842);
nand NAND4 (N14852, N14839, N10555, N5526, N2498);
nand NAND2 (N14853, N14851, N10386);
nor NOR2 (N14854, N14853, N3793);
buf BUF1 (N14855, N14844);
or OR4 (N14856, N14847, N3569, N2462, N2749);
nor NOR4 (N14857, N14830, N4657, N2985, N10876);
nor NOR2 (N14858, N14852, N4522);
buf BUF1 (N14859, N14858);
or OR2 (N14860, N14855, N14619);
nor NOR2 (N14861, N14859, N6048);
nand NAND2 (N14862, N14850, N4333);
nor NOR4 (N14863, N14849, N155, N3943, N385);
nor NOR2 (N14864, N14863, N9329);
or OR2 (N14865, N14864, N11946);
nor NOR4 (N14866, N14845, N7847, N8519, N10870);
and AND4 (N14867, N14833, N5584, N889, N8125);
buf BUF1 (N14868, N14865);
nor NOR3 (N14869, N14867, N472, N2578);
xor XOR2 (N14870, N14854, N6397);
or OR3 (N14871, N14868, N12136, N11388);
nor NOR4 (N14872, N14870, N4461, N2912, N2384);
xor XOR2 (N14873, N14860, N7384);
nand NAND3 (N14874, N14848, N1706, N11513);
buf BUF1 (N14875, N14874);
not NOT1 (N14876, N14862);
or OR2 (N14877, N14871, N710);
nor NOR2 (N14878, N14872, N10807);
and AND3 (N14879, N14877, N10873, N9071);
nor NOR4 (N14880, N14866, N12353, N10311, N6909);
nor NOR3 (N14881, N14879, N1224, N10029);
buf BUF1 (N14882, N14881);
or OR3 (N14883, N14869, N5017, N4940);
and AND3 (N14884, N14875, N10, N136);
buf BUF1 (N14885, N14857);
and AND4 (N14886, N14882, N4300, N14486, N1073);
xor XOR2 (N14887, N14884, N1997);
not NOT1 (N14888, N14856);
nand NAND4 (N14889, N14885, N4211, N2057, N6830);
and AND4 (N14890, N14888, N7944, N10545, N5251);
and AND3 (N14891, N14873, N13842, N3243);
nor NOR4 (N14892, N14861, N4283, N2669, N873);
and AND2 (N14893, N14892, N4086);
or OR3 (N14894, N14890, N6447, N12142);
and AND2 (N14895, N14891, N7320);
and AND2 (N14896, N14886, N285);
and AND3 (N14897, N14887, N7572, N6836);
not NOT1 (N14898, N14878);
buf BUF1 (N14899, N14895);
not NOT1 (N14900, N14894);
xor XOR2 (N14901, N14899, N11374);
xor XOR2 (N14902, N14883, N4494);
not NOT1 (N14903, N14896);
or OR2 (N14904, N14880, N9772);
buf BUF1 (N14905, N14897);
not NOT1 (N14906, N14901);
nand NAND2 (N14907, N14903, N9517);
nor NOR4 (N14908, N14905, N4291, N8271, N8855);
and AND3 (N14909, N14906, N10539, N7045);
xor XOR2 (N14910, N14876, N6882);
and AND2 (N14911, N14900, N6465);
or OR2 (N14912, N14907, N12275);
and AND3 (N14913, N14912, N14629, N8226);
xor XOR2 (N14914, N14893, N2635);
nand NAND4 (N14915, N14911, N520, N5106, N2581);
nor NOR2 (N14916, N14909, N8543);
nor NOR2 (N14917, N14902, N13093);
xor XOR2 (N14918, N14910, N1280);
and AND2 (N14919, N14917, N858);
not NOT1 (N14920, N14914);
buf BUF1 (N14921, N14919);
buf BUF1 (N14922, N14898);
nand NAND4 (N14923, N14916, N11236, N4037, N3347);
nor NOR3 (N14924, N14889, N6091, N12274);
or OR3 (N14925, N14924, N11004, N10052);
xor XOR2 (N14926, N14921, N4483);
nor NOR2 (N14927, N14918, N12767);
and AND3 (N14928, N14926, N6480, N1131);
not NOT1 (N14929, N14927);
xor XOR2 (N14930, N14928, N11501);
nand NAND2 (N14931, N14929, N13398);
or OR3 (N14932, N14920, N10768, N455);
not NOT1 (N14933, N14923);
nor NOR2 (N14934, N14931, N12512);
not NOT1 (N14935, N14933);
nand NAND4 (N14936, N14922, N13838, N13252, N13438);
or OR4 (N14937, N14935, N1531, N10286, N12694);
buf BUF1 (N14938, N14936);
buf BUF1 (N14939, N14913);
or OR4 (N14940, N14915, N13161, N10292, N11870);
buf BUF1 (N14941, N14934);
nor NOR2 (N14942, N14940, N10312);
nor NOR2 (N14943, N14938, N13021);
nand NAND4 (N14944, N14930, N3068, N8148, N12613);
and AND2 (N14945, N14908, N9271);
buf BUF1 (N14946, N14939);
nor NOR3 (N14947, N14946, N12110, N4168);
not NOT1 (N14948, N14925);
buf BUF1 (N14949, N14942);
not NOT1 (N14950, N14948);
not NOT1 (N14951, N14932);
buf BUF1 (N14952, N14937);
xor XOR2 (N14953, N14945, N7353);
xor XOR2 (N14954, N14944, N8813);
not NOT1 (N14955, N14953);
nor NOR2 (N14956, N14949, N189);
buf BUF1 (N14957, N14952);
nand NAND2 (N14958, N14951, N7049);
not NOT1 (N14959, N14955);
nand NAND3 (N14960, N14958, N13920, N2463);
nand NAND3 (N14961, N14960, N10476, N4162);
nand NAND4 (N14962, N14941, N5306, N8621, N14586);
nor NOR2 (N14963, N14904, N9683);
buf BUF1 (N14964, N14957);
buf BUF1 (N14965, N14961);
or OR2 (N14966, N14954, N315);
or OR4 (N14967, N14962, N442, N1937, N13622);
and AND4 (N14968, N14943, N10586, N4420, N8071);
buf BUF1 (N14969, N14964);
or OR4 (N14970, N14950, N4465, N13355, N4339);
not NOT1 (N14971, N14956);
or OR4 (N14972, N14967, N6363, N1004, N2514);
not NOT1 (N14973, N14966);
nor NOR2 (N14974, N14947, N2968);
nand NAND2 (N14975, N14965, N1363);
nand NAND2 (N14976, N14972, N13154);
nor NOR3 (N14977, N14973, N8142, N10793);
or OR2 (N14978, N14976, N10062);
or OR2 (N14979, N14975, N10811);
nand NAND2 (N14980, N14968, N12229);
not NOT1 (N14981, N14979);
not NOT1 (N14982, N14970);
buf BUF1 (N14983, N14974);
xor XOR2 (N14984, N14971, N1925);
nand NAND4 (N14985, N14982, N6726, N12511, N6190);
and AND3 (N14986, N14978, N10650, N10794);
or OR4 (N14987, N14959, N2027, N3219, N11776);
and AND3 (N14988, N14985, N5756, N10384);
nand NAND4 (N14989, N14988, N11815, N5785, N3986);
and AND3 (N14990, N14984, N12968, N10130);
or OR4 (N14991, N14987, N11614, N9131, N8106);
not NOT1 (N14992, N14981);
buf BUF1 (N14993, N14990);
or OR2 (N14994, N14992, N1351);
or OR2 (N14995, N14977, N10760);
or OR3 (N14996, N14989, N12877, N6071);
not NOT1 (N14997, N14995);
nand NAND4 (N14998, N14980, N13402, N4413, N12820);
or OR2 (N14999, N14986, N14360);
or OR4 (N15000, N14969, N6350, N11872, N14186);
buf BUF1 (N15001, N14963);
nor NOR3 (N15002, N14983, N9758, N592);
xor XOR2 (N15003, N14998, N12885);
nor NOR2 (N15004, N15000, N8331);
or OR3 (N15005, N15002, N6767, N11527);
buf BUF1 (N15006, N15004);
buf BUF1 (N15007, N15001);
xor XOR2 (N15008, N14991, N9340);
not NOT1 (N15009, N14993);
nand NAND3 (N15010, N14996, N7730, N1214);
and AND4 (N15011, N15010, N12588, N6749, N8556);
and AND3 (N15012, N15003, N1274, N10247);
nor NOR4 (N15013, N14994, N6782, N3888, N4688);
nand NAND2 (N15014, N14999, N5153);
or OR3 (N15015, N15012, N3525, N1586);
nor NOR4 (N15016, N15006, N4910, N5208, N7926);
buf BUF1 (N15017, N15009);
and AND4 (N15018, N15015, N13225, N7410, N804);
xor XOR2 (N15019, N15018, N2619);
nand NAND3 (N15020, N15011, N11845, N12421);
or OR2 (N15021, N15016, N10528);
nand NAND2 (N15022, N14997, N9632);
and AND3 (N15023, N15007, N3463, N314);
nor NOR2 (N15024, N15021, N13673);
nor NOR4 (N15025, N15022, N405, N1513, N2062);
xor XOR2 (N15026, N15023, N6865);
buf BUF1 (N15027, N15020);
nand NAND4 (N15028, N15026, N8174, N412, N13851);
not NOT1 (N15029, N15025);
buf BUF1 (N15030, N15024);
buf BUF1 (N15031, N15008);
nand NAND4 (N15032, N15029, N4228, N12737, N9828);
nand NAND2 (N15033, N15027, N10653);
nor NOR2 (N15034, N15031, N10006);
xor XOR2 (N15035, N15033, N6316);
and AND4 (N15036, N15034, N12879, N5888, N7379);
nand NAND2 (N15037, N15030, N7101);
xor XOR2 (N15038, N15017, N4171);
buf BUF1 (N15039, N15019);
not NOT1 (N15040, N15032);
buf BUF1 (N15041, N15036);
nand NAND3 (N15042, N15037, N14983, N10091);
buf BUF1 (N15043, N15028);
nor NOR4 (N15044, N15040, N811, N2052, N12982);
buf BUF1 (N15045, N15035);
or OR2 (N15046, N15044, N1617);
nor NOR2 (N15047, N15005, N9008);
xor XOR2 (N15048, N15045, N3416);
and AND4 (N15049, N15038, N8694, N3550, N1507);
and AND4 (N15050, N15047, N453, N7923, N14242);
buf BUF1 (N15051, N15048);
not NOT1 (N15052, N15041);
not NOT1 (N15053, N15050);
nor NOR3 (N15054, N15049, N12520, N2625);
not NOT1 (N15055, N15051);
nor NOR3 (N15056, N15014, N6718, N10491);
xor XOR2 (N15057, N15039, N12946);
buf BUF1 (N15058, N15046);
or OR3 (N15059, N15055, N12851, N13386);
or OR3 (N15060, N15054, N8863, N9478);
or OR3 (N15061, N15056, N4067, N8008);
nand NAND3 (N15062, N15060, N4740, N9159);
and AND2 (N15063, N15013, N1495);
nor NOR4 (N15064, N15059, N4812, N11639, N2511);
buf BUF1 (N15065, N15062);
and AND4 (N15066, N15061, N11341, N1371, N970);
not NOT1 (N15067, N15064);
and AND2 (N15068, N15066, N7725);
buf BUF1 (N15069, N15053);
or OR3 (N15070, N15052, N12204, N8276);
nand NAND2 (N15071, N15070, N13417);
xor XOR2 (N15072, N15071, N12351);
or OR3 (N15073, N15069, N11524, N10130);
or OR2 (N15074, N15065, N1958);
and AND2 (N15075, N15074, N4828);
or OR3 (N15076, N15057, N1909, N10894);
nor NOR3 (N15077, N15068, N10743, N3714);
buf BUF1 (N15078, N15058);
nand NAND2 (N15079, N15077, N6065);
not NOT1 (N15080, N15073);
and AND2 (N15081, N15067, N1755);
xor XOR2 (N15082, N15076, N2164);
and AND3 (N15083, N15082, N253, N149);
not NOT1 (N15084, N15042);
xor XOR2 (N15085, N15063, N9665);
not NOT1 (N15086, N15085);
buf BUF1 (N15087, N15075);
not NOT1 (N15088, N15086);
xor XOR2 (N15089, N15087, N4468);
xor XOR2 (N15090, N15079, N1538);
and AND2 (N15091, N15072, N14687);
not NOT1 (N15092, N15088);
xor XOR2 (N15093, N15084, N6661);
nor NOR4 (N15094, N15091, N9447, N1645, N11720);
nand NAND4 (N15095, N15090, N7310, N13949, N842);
nor NOR2 (N15096, N15093, N1745);
or OR4 (N15097, N15078, N2852, N4591, N12130);
nor NOR2 (N15098, N15095, N2894);
and AND4 (N15099, N15098, N12052, N8596, N7046);
not NOT1 (N15100, N15096);
or OR4 (N15101, N15100, N2822, N5831, N2443);
buf BUF1 (N15102, N15101);
nor NOR2 (N15103, N15043, N14018);
or OR2 (N15104, N15103, N10954);
xor XOR2 (N15105, N15097, N1397);
nand NAND3 (N15106, N15105, N5349, N6011);
xor XOR2 (N15107, N15092, N5551);
nand NAND4 (N15108, N15104, N14524, N7190, N321);
nand NAND3 (N15109, N15081, N2672, N6038);
nand NAND3 (N15110, N15099, N1958, N3053);
or OR3 (N15111, N15106, N3343, N13430);
xor XOR2 (N15112, N15109, N14657);
buf BUF1 (N15113, N15110);
buf BUF1 (N15114, N15094);
and AND2 (N15115, N15111, N741);
nor NOR3 (N15116, N15102, N4522, N5874);
or OR4 (N15117, N15108, N8014, N10258, N3310);
or OR4 (N15118, N15113, N11778, N10825, N9892);
and AND3 (N15119, N15116, N9605, N11761);
nand NAND2 (N15120, N15119, N6944);
nor NOR3 (N15121, N15107, N10924, N124);
buf BUF1 (N15122, N15112);
and AND4 (N15123, N15114, N827, N10137, N94);
not NOT1 (N15124, N15089);
nor NOR4 (N15125, N15122, N3673, N7653, N1571);
or OR3 (N15126, N15080, N1614, N14972);
or OR4 (N15127, N15123, N6800, N12457, N12589);
nor NOR2 (N15128, N15117, N5482);
xor XOR2 (N15129, N15127, N9304);
or OR3 (N15130, N15125, N6449, N13283);
buf BUF1 (N15131, N15115);
or OR2 (N15132, N15130, N6856);
xor XOR2 (N15133, N15131, N2812);
nor NOR2 (N15134, N15128, N5985);
not NOT1 (N15135, N15133);
nand NAND4 (N15136, N15121, N8650, N2895, N11187);
nor NOR2 (N15137, N15134, N6348);
nor NOR4 (N15138, N15129, N1316, N3036, N3722);
buf BUF1 (N15139, N15132);
nand NAND3 (N15140, N15138, N14013, N11301);
buf BUF1 (N15141, N15136);
not NOT1 (N15142, N15139);
nand NAND2 (N15143, N15135, N13469);
and AND3 (N15144, N15126, N1265, N306);
and AND2 (N15145, N15120, N11827);
not NOT1 (N15146, N15118);
and AND3 (N15147, N15144, N1000, N4688);
not NOT1 (N15148, N15137);
and AND2 (N15149, N15146, N10701);
not NOT1 (N15150, N15149);
buf BUF1 (N15151, N15147);
nand NAND3 (N15152, N15151, N9945, N12786);
nand NAND3 (N15153, N15152, N14103, N217);
buf BUF1 (N15154, N15142);
nand NAND4 (N15155, N15141, N4935, N7764, N4357);
and AND2 (N15156, N15140, N2104);
or OR4 (N15157, N15153, N11489, N4544, N13234);
and AND3 (N15158, N15143, N5827, N12363);
not NOT1 (N15159, N15083);
xor XOR2 (N15160, N15159, N2539);
and AND3 (N15161, N15160, N3980, N5576);
and AND4 (N15162, N15157, N14898, N10148, N11463);
nand NAND3 (N15163, N15148, N8575, N9997);
xor XOR2 (N15164, N15163, N5047);
and AND4 (N15165, N15156, N8637, N8817, N4150);
nor NOR2 (N15166, N15154, N3090);
or OR4 (N15167, N15162, N7472, N430, N5280);
xor XOR2 (N15168, N15150, N13266);
nand NAND3 (N15169, N15145, N10889, N12745);
buf BUF1 (N15170, N15155);
xor XOR2 (N15171, N15167, N12318);
or OR2 (N15172, N15164, N4811);
and AND2 (N15173, N15165, N7955);
or OR3 (N15174, N15161, N13790, N14075);
nor NOR2 (N15175, N15174, N6854);
or OR4 (N15176, N15175, N9339, N4915, N6700);
buf BUF1 (N15177, N15172);
nor NOR4 (N15178, N15171, N14839, N7614, N13844);
or OR3 (N15179, N15178, N498, N102);
xor XOR2 (N15180, N15124, N3281);
xor XOR2 (N15181, N15173, N8447);
nand NAND2 (N15182, N15170, N12438);
xor XOR2 (N15183, N15158, N5471);
nand NAND2 (N15184, N15179, N13766);
not NOT1 (N15185, N15181);
not NOT1 (N15186, N15177);
xor XOR2 (N15187, N15169, N12748);
or OR4 (N15188, N15185, N6511, N6530, N2264);
nor NOR3 (N15189, N15176, N113, N2587);
nand NAND3 (N15190, N15189, N2917, N14650);
and AND4 (N15191, N15168, N12081, N5644, N3102);
buf BUF1 (N15192, N15187);
xor XOR2 (N15193, N15190, N10820);
nand NAND4 (N15194, N15180, N13027, N1254, N4613);
or OR4 (N15195, N15183, N14903, N3809, N7675);
nor NOR4 (N15196, N15193, N12227, N3686, N950);
and AND2 (N15197, N15184, N9653);
and AND3 (N15198, N15166, N8387, N8918);
nor NOR4 (N15199, N15182, N4578, N7099, N1939);
and AND4 (N15200, N15194, N5478, N11609, N1781);
nor NOR3 (N15201, N15197, N2670, N5156);
or OR2 (N15202, N15201, N3727);
buf BUF1 (N15203, N15191);
nand NAND4 (N15204, N15199, N7938, N13729, N12097);
or OR3 (N15205, N15186, N8256, N6541);
not NOT1 (N15206, N15203);
not NOT1 (N15207, N15206);
nor NOR3 (N15208, N15200, N3152, N6549);
not NOT1 (N15209, N15205);
or OR2 (N15210, N15204, N12665);
and AND4 (N15211, N15207, N1585, N1554, N4720);
not NOT1 (N15212, N15195);
buf BUF1 (N15213, N15196);
nor NOR3 (N15214, N15198, N12714, N10732);
not NOT1 (N15215, N15192);
buf BUF1 (N15216, N15208);
xor XOR2 (N15217, N15202, N1206);
not NOT1 (N15218, N15212);
not NOT1 (N15219, N15211);
nor NOR3 (N15220, N15219, N8195, N6234);
not NOT1 (N15221, N15188);
nor NOR3 (N15222, N15214, N13502, N13225);
not NOT1 (N15223, N15215);
and AND2 (N15224, N15220, N1194);
not NOT1 (N15225, N15218);
nor NOR4 (N15226, N15222, N3516, N5317, N1820);
xor XOR2 (N15227, N15225, N8373);
and AND2 (N15228, N15217, N5774);
and AND3 (N15229, N15227, N8967, N13637);
or OR2 (N15230, N15213, N14815);
not NOT1 (N15231, N15230);
and AND3 (N15232, N15223, N8053, N10379);
not NOT1 (N15233, N15229);
buf BUF1 (N15234, N15226);
not NOT1 (N15235, N15233);
or OR3 (N15236, N15232, N3557, N4021);
xor XOR2 (N15237, N15216, N11793);
buf BUF1 (N15238, N15224);
and AND2 (N15239, N15237, N7955);
buf BUF1 (N15240, N15235);
and AND2 (N15241, N15238, N527);
nand NAND2 (N15242, N15210, N8303);
buf BUF1 (N15243, N15209);
buf BUF1 (N15244, N15242);
or OR2 (N15245, N15228, N14345);
nor NOR3 (N15246, N15221, N4477, N8953);
and AND2 (N15247, N15244, N12335);
xor XOR2 (N15248, N15247, N12411);
xor XOR2 (N15249, N15243, N7876);
xor XOR2 (N15250, N15231, N15212);
nor NOR4 (N15251, N15248, N14869, N10077, N2660);
or OR3 (N15252, N15234, N5745, N6814);
buf BUF1 (N15253, N15250);
buf BUF1 (N15254, N15240);
buf BUF1 (N15255, N15253);
xor XOR2 (N15256, N15249, N783);
nor NOR3 (N15257, N15239, N11501, N2652);
and AND4 (N15258, N15236, N2411, N9084, N3549);
buf BUF1 (N15259, N15251);
buf BUF1 (N15260, N15254);
or OR4 (N15261, N15260, N7849, N10240, N12481);
not NOT1 (N15262, N15261);
xor XOR2 (N15263, N15255, N14095);
not NOT1 (N15264, N15256);
nand NAND3 (N15265, N15246, N4476, N6037);
and AND2 (N15266, N15263, N12044);
buf BUF1 (N15267, N15241);
nor NOR4 (N15268, N15264, N11855, N11099, N12120);
nand NAND3 (N15269, N15268, N559, N13297);
not NOT1 (N15270, N15266);
buf BUF1 (N15271, N15270);
or OR2 (N15272, N15258, N8962);
not NOT1 (N15273, N15245);
and AND2 (N15274, N15259, N4976);
and AND4 (N15275, N15267, N3582, N11762, N4837);
not NOT1 (N15276, N15265);
nand NAND2 (N15277, N15252, N12524);
buf BUF1 (N15278, N15262);
not NOT1 (N15279, N15257);
xor XOR2 (N15280, N15279, N2150);
nand NAND2 (N15281, N15276, N7561);
buf BUF1 (N15282, N15278);
nor NOR3 (N15283, N15282, N5422, N4925);
not NOT1 (N15284, N15273);
xor XOR2 (N15285, N15281, N2622);
or OR3 (N15286, N15277, N14590, N3694);
xor XOR2 (N15287, N15286, N4310);
buf BUF1 (N15288, N15275);
nor NOR4 (N15289, N15271, N3482, N5974, N8938);
xor XOR2 (N15290, N15284, N10784);
and AND3 (N15291, N15274, N2938, N8391);
nor NOR2 (N15292, N15269, N14473);
nor NOR3 (N15293, N15288, N1327, N3631);
and AND2 (N15294, N15289, N8019);
xor XOR2 (N15295, N15294, N14242);
buf BUF1 (N15296, N15280);
and AND2 (N15297, N15295, N6825);
xor XOR2 (N15298, N15293, N9935);
not NOT1 (N15299, N15283);
and AND3 (N15300, N15299, N14950, N10623);
and AND2 (N15301, N15300, N11333);
or OR2 (N15302, N15285, N7711);
buf BUF1 (N15303, N15272);
nand NAND2 (N15304, N15296, N5956);
or OR2 (N15305, N15292, N9212);
not NOT1 (N15306, N15303);
xor XOR2 (N15307, N15305, N1110);
not NOT1 (N15308, N15290);
xor XOR2 (N15309, N15308, N11890);
buf BUF1 (N15310, N15291);
or OR2 (N15311, N15309, N12364);
nor NOR4 (N15312, N15310, N4853, N2644, N9035);
xor XOR2 (N15313, N15304, N8420);
buf BUF1 (N15314, N15302);
and AND3 (N15315, N15313, N3491, N15112);
xor XOR2 (N15316, N15315, N5317);
xor XOR2 (N15317, N15312, N4663);
buf BUF1 (N15318, N15317);
nand NAND2 (N15319, N15314, N14007);
not NOT1 (N15320, N15297);
xor XOR2 (N15321, N15287, N14292);
or OR2 (N15322, N15321, N9994);
nand NAND3 (N15323, N15306, N8329, N14943);
not NOT1 (N15324, N15320);
xor XOR2 (N15325, N15311, N14035);
or OR4 (N15326, N15324, N2870, N8998, N6333);
xor XOR2 (N15327, N15326, N5142);
or OR2 (N15328, N15318, N15082);
buf BUF1 (N15329, N15298);
or OR3 (N15330, N15323, N5966, N1464);
xor XOR2 (N15331, N15319, N11402);
and AND2 (N15332, N15325, N4602);
not NOT1 (N15333, N15329);
not NOT1 (N15334, N15316);
buf BUF1 (N15335, N15301);
and AND3 (N15336, N15330, N13611, N1656);
and AND2 (N15337, N15332, N744);
xor XOR2 (N15338, N15327, N2556);
xor XOR2 (N15339, N15333, N12452);
and AND4 (N15340, N15331, N1165, N5576, N5253);
xor XOR2 (N15341, N15334, N13331);
or OR3 (N15342, N15338, N2553, N14058);
or OR3 (N15343, N15340, N13765, N5661);
and AND2 (N15344, N15337, N12311);
and AND2 (N15345, N15341, N2866);
nand NAND3 (N15346, N15344, N5341, N14314);
nor NOR2 (N15347, N15342, N3956);
not NOT1 (N15348, N15345);
buf BUF1 (N15349, N15343);
not NOT1 (N15350, N15339);
buf BUF1 (N15351, N15349);
not NOT1 (N15352, N15307);
xor XOR2 (N15353, N15348, N1160);
xor XOR2 (N15354, N15328, N1562);
buf BUF1 (N15355, N15352);
buf BUF1 (N15356, N15335);
and AND2 (N15357, N15355, N936);
xor XOR2 (N15358, N15347, N8909);
nor NOR3 (N15359, N15356, N14788, N967);
or OR2 (N15360, N15358, N2481);
buf BUF1 (N15361, N15357);
nand NAND3 (N15362, N15336, N6090, N11208);
xor XOR2 (N15363, N15351, N2995);
nor NOR3 (N15364, N15353, N12437, N9907);
buf BUF1 (N15365, N15364);
xor XOR2 (N15366, N15350, N3593);
xor XOR2 (N15367, N15346, N9372);
or OR4 (N15368, N15362, N2429, N6932, N12774);
buf BUF1 (N15369, N15368);
nand NAND4 (N15370, N15365, N9844, N13977, N1999);
not NOT1 (N15371, N15322);
buf BUF1 (N15372, N15363);
nand NAND2 (N15373, N15360, N1530);
nor NOR4 (N15374, N15370, N956, N7024, N263);
xor XOR2 (N15375, N15369, N5747);
xor XOR2 (N15376, N15361, N15336);
or OR3 (N15377, N15366, N10799, N6732);
nor NOR4 (N15378, N15374, N880, N7457, N3310);
buf BUF1 (N15379, N15376);
nor NOR3 (N15380, N15371, N2436, N6493);
nand NAND4 (N15381, N15379, N10492, N11185, N12975);
buf BUF1 (N15382, N15359);
or OR4 (N15383, N15367, N13653, N8833, N1836);
nor NOR4 (N15384, N15372, N12324, N9604, N7281);
or OR4 (N15385, N15384, N4302, N95, N2629);
nor NOR4 (N15386, N15378, N8208, N9958, N2796);
not NOT1 (N15387, N15377);
xor XOR2 (N15388, N15373, N494);
not NOT1 (N15389, N15388);
nor NOR3 (N15390, N15375, N11827, N4127);
and AND2 (N15391, N15385, N5187);
or OR4 (N15392, N15354, N8530, N6231, N413);
buf BUF1 (N15393, N15386);
or OR3 (N15394, N15389, N15366, N6552);
or OR2 (N15395, N15394, N330);
and AND2 (N15396, N15387, N11788);
not NOT1 (N15397, N15395);
nand NAND3 (N15398, N15397, N7205, N6766);
nand NAND2 (N15399, N15396, N9423);
not NOT1 (N15400, N15380);
or OR3 (N15401, N15400, N6656, N5513);
or OR3 (N15402, N15401, N14218, N11494);
or OR2 (N15403, N15392, N5829);
nand NAND3 (N15404, N15383, N11532, N13685);
buf BUF1 (N15405, N15398);
not NOT1 (N15406, N15402);
not NOT1 (N15407, N15403);
nand NAND4 (N15408, N15404, N3566, N8667, N8003);
and AND3 (N15409, N15391, N5800, N3507);
not NOT1 (N15410, N15399);
not NOT1 (N15411, N15406);
xor XOR2 (N15412, N15393, N14543);
nor NOR2 (N15413, N15381, N3541);
or OR2 (N15414, N15409, N1430);
nor NOR4 (N15415, N15413, N7723, N6741, N6343);
xor XOR2 (N15416, N15412, N11935);
or OR3 (N15417, N15410, N2380, N6099);
or OR4 (N15418, N15390, N15342, N14857, N14102);
not NOT1 (N15419, N15408);
buf BUF1 (N15420, N15415);
buf BUF1 (N15421, N15418);
and AND4 (N15422, N15421, N153, N10892, N3592);
xor XOR2 (N15423, N15382, N9069);
not NOT1 (N15424, N15422);
nand NAND3 (N15425, N15405, N1610, N3397);
not NOT1 (N15426, N15419);
xor XOR2 (N15427, N15407, N12326);
or OR4 (N15428, N15426, N26, N574, N2492);
nand NAND4 (N15429, N15416, N10545, N176, N9307);
nor NOR2 (N15430, N15411, N6210);
nand NAND2 (N15431, N15417, N15336);
buf BUF1 (N15432, N15429);
and AND4 (N15433, N15431, N10587, N1942, N14719);
and AND3 (N15434, N15427, N5338, N10413);
not NOT1 (N15435, N15433);
xor XOR2 (N15436, N15434, N4700);
not NOT1 (N15437, N15436);
and AND4 (N15438, N15428, N3357, N11745, N8352);
nor NOR3 (N15439, N15424, N12113, N601);
buf BUF1 (N15440, N15435);
xor XOR2 (N15441, N15440, N106);
buf BUF1 (N15442, N15441);
nor NOR2 (N15443, N15437, N2533);
buf BUF1 (N15444, N15414);
nand NAND4 (N15445, N15443, N4182, N15055, N10865);
nor NOR4 (N15446, N15432, N99, N2851, N9159);
buf BUF1 (N15447, N15425);
and AND2 (N15448, N15420, N9830);
buf BUF1 (N15449, N15442);
xor XOR2 (N15450, N15445, N1193);
nor NOR3 (N15451, N15446, N6815, N14517);
or OR2 (N15452, N15447, N12019);
or OR3 (N15453, N15451, N7603, N7386);
nand NAND2 (N15454, N15452, N9623);
nor NOR4 (N15455, N15454, N7985, N14570, N5189);
nor NOR4 (N15456, N15453, N14712, N492, N14646);
buf BUF1 (N15457, N15450);
nand NAND3 (N15458, N15439, N6948, N9571);
buf BUF1 (N15459, N15456);
nand NAND3 (N15460, N15459, N5623, N13323);
xor XOR2 (N15461, N15449, N13833);
or OR4 (N15462, N15458, N13285, N11224, N8734);
or OR4 (N15463, N15430, N1588, N9984, N7556);
not NOT1 (N15464, N15460);
buf BUF1 (N15465, N15463);
nor NOR2 (N15466, N15448, N3252);
not NOT1 (N15467, N15466);
not NOT1 (N15468, N15438);
and AND2 (N15469, N15468, N8017);
not NOT1 (N15470, N15461);
nand NAND3 (N15471, N15455, N2578, N10037);
and AND2 (N15472, N15465, N5013);
or OR2 (N15473, N15469, N507);
and AND2 (N15474, N15473, N4515);
not NOT1 (N15475, N15464);
not NOT1 (N15476, N15475);
or OR2 (N15477, N15423, N14282);
not NOT1 (N15478, N15476);
buf BUF1 (N15479, N15471);
xor XOR2 (N15480, N15470, N10406);
and AND3 (N15481, N15477, N14787, N14340);
buf BUF1 (N15482, N15462);
not NOT1 (N15483, N15457);
buf BUF1 (N15484, N15479);
xor XOR2 (N15485, N15467, N9512);
and AND2 (N15486, N15444, N10492);
nand NAND2 (N15487, N15480, N9788);
not NOT1 (N15488, N15474);
or OR4 (N15489, N15484, N12085, N355, N11831);
nor NOR3 (N15490, N15489, N1607, N11182);
xor XOR2 (N15491, N15486, N8710);
not NOT1 (N15492, N15491);
and AND4 (N15493, N15478, N7912, N12260, N1404);
nor NOR3 (N15494, N15488, N6267, N15110);
or OR2 (N15495, N15493, N5479);
or OR2 (N15496, N15494, N10763);
and AND4 (N15497, N15482, N385, N845, N652);
or OR4 (N15498, N15483, N9645, N8389, N5426);
or OR4 (N15499, N15490, N5033, N12485, N1323);
or OR3 (N15500, N15485, N1815, N13944);
buf BUF1 (N15501, N15481);
buf BUF1 (N15502, N15499);
nand NAND2 (N15503, N15487, N636);
buf BUF1 (N15504, N15501);
nand NAND3 (N15505, N15504, N11467, N1263);
nand NAND4 (N15506, N15503, N12614, N12700, N4618);
nand NAND4 (N15507, N15497, N4985, N14302, N4678);
nor NOR2 (N15508, N15502, N15321);
nor NOR3 (N15509, N15492, N5689, N13775);
buf BUF1 (N15510, N15498);
xor XOR2 (N15511, N15507, N3821);
nor NOR2 (N15512, N15500, N14554);
nor NOR2 (N15513, N15512, N11789);
nand NAND3 (N15514, N15510, N2421, N15457);
nand NAND2 (N15515, N15495, N2915);
not NOT1 (N15516, N15511);
nor NOR2 (N15517, N15472, N11206);
or OR3 (N15518, N15516, N287, N14616);
nand NAND4 (N15519, N15517, N369, N11562, N7343);
and AND2 (N15520, N15506, N1785);
and AND4 (N15521, N15513, N11718, N479, N6771);
buf BUF1 (N15522, N15515);
not NOT1 (N15523, N15520);
nand NAND4 (N15524, N15514, N14497, N1662, N3731);
buf BUF1 (N15525, N15521);
xor XOR2 (N15526, N15509, N5362);
nor NOR2 (N15527, N15508, N7560);
buf BUF1 (N15528, N15527);
buf BUF1 (N15529, N15518);
or OR3 (N15530, N15524, N10524, N9906);
and AND4 (N15531, N15522, N8002, N13898, N11638);
not NOT1 (N15532, N15505);
nand NAND2 (N15533, N15526, N1009);
not NOT1 (N15534, N15530);
xor XOR2 (N15535, N15532, N4307);
nor NOR4 (N15536, N15531, N6502, N7784, N5986);
xor XOR2 (N15537, N15519, N1777);
or OR2 (N15538, N15535, N11706);
or OR4 (N15539, N15528, N2878, N2440, N2916);
buf BUF1 (N15540, N15533);
or OR3 (N15541, N15538, N11432, N12655);
and AND2 (N15542, N15523, N6175);
nand NAND2 (N15543, N15496, N2486);
buf BUF1 (N15544, N15540);
nor NOR4 (N15545, N15542, N3093, N4613, N1152);
buf BUF1 (N15546, N15545);
buf BUF1 (N15547, N15537);
nor NOR2 (N15548, N15534, N1376);
and AND2 (N15549, N15541, N12597);
nand NAND3 (N15550, N15549, N14337, N11999);
nor NOR4 (N15551, N15529, N2297, N4158, N6315);
buf BUF1 (N15552, N15536);
nand NAND3 (N15553, N15525, N12384, N2626);
not NOT1 (N15554, N15552);
and AND3 (N15555, N15553, N13386, N11794);
xor XOR2 (N15556, N15555, N7787);
nand NAND3 (N15557, N15539, N914, N3680);
not NOT1 (N15558, N15556);
or OR3 (N15559, N15547, N5741, N11990);
or OR2 (N15560, N15551, N1519);
or OR4 (N15561, N15557, N4395, N12748, N2866);
xor XOR2 (N15562, N15561, N7598);
or OR4 (N15563, N15543, N9493, N7402, N8682);
nand NAND2 (N15564, N15546, N14186);
xor XOR2 (N15565, N15554, N7369);
nand NAND2 (N15566, N15563, N12332);
or OR4 (N15567, N15559, N13420, N1927, N10804);
xor XOR2 (N15568, N15544, N10278);
xor XOR2 (N15569, N15562, N6288);
nand NAND3 (N15570, N15568, N13612, N12033);
and AND3 (N15571, N15565, N11617, N14207);
buf BUF1 (N15572, N15569);
not NOT1 (N15573, N15572);
buf BUF1 (N15574, N15558);
nor NOR2 (N15575, N15548, N8388);
nor NOR4 (N15576, N15564, N4417, N15203, N1994);
not NOT1 (N15577, N15567);
not NOT1 (N15578, N15576);
not NOT1 (N15579, N15577);
nor NOR4 (N15580, N15560, N5825, N5096, N2692);
nand NAND2 (N15581, N15580, N8973);
nor NOR4 (N15582, N15578, N6452, N1378, N515);
or OR3 (N15583, N15575, N4265, N7010);
nand NAND4 (N15584, N15570, N207, N9934, N13872);
nand NAND3 (N15585, N15571, N14246, N712);
xor XOR2 (N15586, N15581, N74);
nand NAND4 (N15587, N15583, N15297, N1101, N9510);
and AND3 (N15588, N15579, N3936, N5498);
nor NOR4 (N15589, N15582, N65, N10983, N5470);
and AND4 (N15590, N15586, N8637, N11564, N4855);
not NOT1 (N15591, N15588);
nand NAND3 (N15592, N15566, N3514, N6759);
nand NAND4 (N15593, N15574, N340, N7714, N11530);
nor NOR3 (N15594, N15592, N575, N13977);
buf BUF1 (N15595, N15591);
nand NAND3 (N15596, N15584, N685, N13400);
nand NAND2 (N15597, N15593, N14579);
nor NOR3 (N15598, N15590, N4971, N550);
buf BUF1 (N15599, N15573);
or OR4 (N15600, N15599, N7857, N1007, N7197);
and AND3 (N15601, N15594, N8946, N13270);
buf BUF1 (N15602, N15598);
nand NAND4 (N15603, N15597, N854, N8139, N2023);
buf BUF1 (N15604, N15550);
nand NAND3 (N15605, N15595, N2181, N8196);
xor XOR2 (N15606, N15605, N8224);
nand NAND3 (N15607, N15589, N1505, N7280);
nand NAND4 (N15608, N15587, N5882, N11651, N7541);
buf BUF1 (N15609, N15596);
and AND2 (N15610, N15601, N1400);
or OR3 (N15611, N15608, N1924, N5881);
nand NAND2 (N15612, N15602, N14091);
or OR3 (N15613, N15607, N6516, N4508);
or OR2 (N15614, N15610, N10076);
nand NAND2 (N15615, N15604, N4428);
nand NAND3 (N15616, N15609, N7703, N4705);
nand NAND4 (N15617, N15585, N2037, N9075, N12320);
buf BUF1 (N15618, N15614);
nand NAND3 (N15619, N15611, N334, N11307);
xor XOR2 (N15620, N15613, N7542);
and AND2 (N15621, N15618, N4171);
nand NAND4 (N15622, N15612, N8033, N12073, N732);
nor NOR3 (N15623, N15621, N11551, N938);
xor XOR2 (N15624, N15617, N987);
nor NOR2 (N15625, N15606, N2514);
and AND4 (N15626, N15625, N858, N14657, N13500);
not NOT1 (N15627, N15620);
buf BUF1 (N15628, N15622);
or OR4 (N15629, N15627, N1119, N12105, N5160);
nand NAND2 (N15630, N15619, N2379);
xor XOR2 (N15631, N15629, N10583);
or OR3 (N15632, N15603, N909, N7621);
xor XOR2 (N15633, N15615, N1859);
xor XOR2 (N15634, N15624, N6826);
nand NAND4 (N15635, N15626, N9606, N3826, N6074);
not NOT1 (N15636, N15630);
nor NOR2 (N15637, N15628, N6355);
nand NAND4 (N15638, N15634, N6211, N3579, N160);
nand NAND2 (N15639, N15636, N11680);
and AND2 (N15640, N15631, N4574);
nor NOR4 (N15641, N15635, N8535, N9389, N5393);
or OR4 (N15642, N15639, N13856, N4232, N69);
not NOT1 (N15643, N15633);
nand NAND3 (N15644, N15600, N3538, N9633);
or OR3 (N15645, N15637, N11693, N14512);
not NOT1 (N15646, N15643);
nand NAND2 (N15647, N15642, N14927);
and AND2 (N15648, N15623, N4925);
buf BUF1 (N15649, N15645);
not NOT1 (N15650, N15644);
or OR2 (N15651, N15647, N7014);
nor NOR4 (N15652, N15640, N9787, N10031, N3789);
xor XOR2 (N15653, N15652, N12933);
xor XOR2 (N15654, N15638, N7922);
nand NAND3 (N15655, N15651, N10741, N13375);
xor XOR2 (N15656, N15616, N7613);
nand NAND4 (N15657, N15632, N5517, N6512, N11087);
nand NAND2 (N15658, N15657, N2467);
xor XOR2 (N15659, N15655, N13745);
and AND4 (N15660, N15646, N4405, N3159, N1022);
or OR2 (N15661, N15659, N2925);
buf BUF1 (N15662, N15641);
xor XOR2 (N15663, N15653, N246);
or OR2 (N15664, N15650, N4753);
nor NOR3 (N15665, N15664, N15169, N10854);
and AND2 (N15666, N15649, N15637);
buf BUF1 (N15667, N15663);
xor XOR2 (N15668, N15660, N15455);
or OR4 (N15669, N15661, N722, N6659, N3367);
and AND2 (N15670, N15665, N3422);
xor XOR2 (N15671, N15658, N53);
nor NOR4 (N15672, N15648, N4422, N5985, N9039);
xor XOR2 (N15673, N15666, N13855);
and AND4 (N15674, N15673, N2864, N4574, N6398);
nand NAND3 (N15675, N15654, N706, N200);
not NOT1 (N15676, N15670);
and AND4 (N15677, N15669, N15564, N5888, N8695);
xor XOR2 (N15678, N15671, N5186);
or OR4 (N15679, N15667, N10978, N14060, N12703);
buf BUF1 (N15680, N15662);
not NOT1 (N15681, N15656);
nand NAND2 (N15682, N15676, N12989);
buf BUF1 (N15683, N15681);
and AND3 (N15684, N15678, N8563, N10890);
nor NOR4 (N15685, N15674, N9608, N15298, N255);
nand NAND4 (N15686, N15668, N8452, N7664, N3906);
buf BUF1 (N15687, N15680);
buf BUF1 (N15688, N15684);
nor NOR4 (N15689, N15688, N7376, N12790, N10360);
not NOT1 (N15690, N15686);
xor XOR2 (N15691, N15683, N9037);
xor XOR2 (N15692, N15690, N15662);
or OR3 (N15693, N15691, N14804, N7149);
nand NAND2 (N15694, N15689, N9245);
or OR2 (N15695, N15675, N4367);
nand NAND4 (N15696, N15687, N15482, N15484, N10543);
or OR3 (N15697, N15693, N8845, N12232);
xor XOR2 (N15698, N15695, N8151);
not NOT1 (N15699, N15685);
xor XOR2 (N15700, N15672, N9312);
nand NAND2 (N15701, N15694, N10762);
buf BUF1 (N15702, N15677);
nand NAND4 (N15703, N15698, N6782, N6762, N2850);
xor XOR2 (N15704, N15697, N2344);
and AND2 (N15705, N15700, N3037);
nor NOR2 (N15706, N15699, N10250);
nor NOR3 (N15707, N15682, N1090, N6216);
not NOT1 (N15708, N15696);
or OR2 (N15709, N15706, N101);
and AND3 (N15710, N15707, N1154, N13689);
and AND2 (N15711, N15701, N11027);
nor NOR3 (N15712, N15704, N12148, N8268);
and AND4 (N15713, N15709, N14143, N1175, N15269);
not NOT1 (N15714, N15713);
nand NAND2 (N15715, N15705, N4618);
buf BUF1 (N15716, N15710);
not NOT1 (N15717, N15708);
buf BUF1 (N15718, N15679);
xor XOR2 (N15719, N15712, N4934);
buf BUF1 (N15720, N15711);
nand NAND2 (N15721, N15718, N4115);
and AND4 (N15722, N15692, N9982, N14662, N10999);
nand NAND2 (N15723, N15716, N5001);
not NOT1 (N15724, N15717);
xor XOR2 (N15725, N15723, N14465);
nand NAND3 (N15726, N15725, N12202, N8746);
nor NOR3 (N15727, N15703, N3695, N911);
nand NAND3 (N15728, N15726, N13694, N8733);
and AND4 (N15729, N15727, N9055, N15711, N4661);
buf BUF1 (N15730, N15714);
or OR2 (N15731, N15722, N4043);
buf BUF1 (N15732, N15702);
nor NOR4 (N15733, N15724, N12310, N6000, N2813);
not NOT1 (N15734, N15719);
not NOT1 (N15735, N15721);
not NOT1 (N15736, N15733);
xor XOR2 (N15737, N15731, N3571);
not NOT1 (N15738, N15732);
not NOT1 (N15739, N15720);
and AND4 (N15740, N15737, N14591, N15371, N3464);
not NOT1 (N15741, N15738);
xor XOR2 (N15742, N15729, N11272);
and AND4 (N15743, N15736, N6225, N13956, N5767);
xor XOR2 (N15744, N15739, N2052);
or OR2 (N15745, N15728, N10672);
and AND4 (N15746, N15735, N7072, N8782, N10000);
nand NAND2 (N15747, N15741, N7155);
nor NOR3 (N15748, N15747, N11726, N10584);
or OR3 (N15749, N15740, N12400, N7780);
or OR2 (N15750, N15743, N15066);
not NOT1 (N15751, N15730);
or OR3 (N15752, N15749, N1792, N4194);
nand NAND3 (N15753, N15742, N3494, N7299);
and AND4 (N15754, N15752, N10386, N3657, N11739);
or OR3 (N15755, N15734, N2760, N6315);
buf BUF1 (N15756, N15753);
nor NOR4 (N15757, N15754, N10378, N3118, N917);
and AND4 (N15758, N15750, N583, N9458, N5340);
xor XOR2 (N15759, N15746, N15511);
and AND2 (N15760, N15745, N4415);
or OR3 (N15761, N15756, N9108, N12233);
and AND3 (N15762, N15757, N4210, N15618);
xor XOR2 (N15763, N15755, N3075);
not NOT1 (N15764, N15763);
and AND2 (N15765, N15764, N5091);
or OR4 (N15766, N15761, N11110, N3211, N13542);
nand NAND4 (N15767, N15766, N2643, N2313, N14257);
and AND4 (N15768, N15765, N6970, N6368, N13306);
buf BUF1 (N15769, N15758);
buf BUF1 (N15770, N15748);
buf BUF1 (N15771, N15768);
buf BUF1 (N15772, N15767);
not NOT1 (N15773, N15762);
or OR4 (N15774, N15744, N5080, N8228, N3992);
or OR3 (N15775, N15715, N14390, N12329);
not NOT1 (N15776, N15774);
nor NOR2 (N15777, N15771, N14098);
not NOT1 (N15778, N15777);
nor NOR2 (N15779, N15778, N9553);
nand NAND4 (N15780, N15759, N10667, N14093, N11031);
xor XOR2 (N15781, N15751, N8935);
not NOT1 (N15782, N15776);
buf BUF1 (N15783, N15782);
not NOT1 (N15784, N15773);
nor NOR2 (N15785, N15784, N1551);
buf BUF1 (N15786, N15780);
or OR3 (N15787, N15781, N8846, N13505);
or OR4 (N15788, N15785, N3799, N6259, N6671);
nand NAND3 (N15789, N15770, N9672, N14099);
not NOT1 (N15790, N15788);
and AND4 (N15791, N15789, N718, N6900, N4773);
nand NAND2 (N15792, N15775, N9918);
nand NAND3 (N15793, N15791, N5764, N7623);
nor NOR4 (N15794, N15783, N14845, N10913, N5788);
nand NAND4 (N15795, N15786, N11949, N10161, N7900);
and AND3 (N15796, N15795, N7521, N2711);
xor XOR2 (N15797, N15794, N13988);
nor NOR3 (N15798, N15779, N6450, N12537);
nor NOR4 (N15799, N15793, N4669, N33, N7547);
or OR4 (N15800, N15787, N7537, N11435, N8009);
nor NOR4 (N15801, N15798, N3984, N11250, N15543);
not NOT1 (N15802, N15797);
xor XOR2 (N15803, N15790, N2952);
buf BUF1 (N15804, N15799);
xor XOR2 (N15805, N15796, N10796);
nor NOR3 (N15806, N15802, N5868, N1162);
buf BUF1 (N15807, N15806);
not NOT1 (N15808, N15807);
nand NAND4 (N15809, N15760, N1256, N9567, N13639);
and AND2 (N15810, N15804, N3347);
buf BUF1 (N15811, N15801);
and AND3 (N15812, N15792, N15614, N15784);
xor XOR2 (N15813, N15772, N8129);
not NOT1 (N15814, N15809);
buf BUF1 (N15815, N15803);
nand NAND4 (N15816, N15812, N1449, N5175, N11116);
nand NAND2 (N15817, N15815, N13563);
nor NOR2 (N15818, N15810, N14065);
not NOT1 (N15819, N15818);
nor NOR2 (N15820, N15808, N12775);
not NOT1 (N15821, N15805);
nor NOR3 (N15822, N15816, N15686, N10707);
buf BUF1 (N15823, N15811);
and AND4 (N15824, N15819, N2206, N8181, N797);
or OR3 (N15825, N15800, N12622, N2237);
buf BUF1 (N15826, N15820);
and AND2 (N15827, N15769, N7026);
or OR4 (N15828, N15823, N14, N706, N15288);
xor XOR2 (N15829, N15827, N812);
or OR3 (N15830, N15828, N2136, N3368);
and AND3 (N15831, N15822, N6681, N11524);
nand NAND2 (N15832, N15821, N15213);
nand NAND4 (N15833, N15813, N7612, N10490, N5397);
or OR2 (N15834, N15824, N10709);
buf BUF1 (N15835, N15825);
or OR4 (N15836, N15830, N10794, N5292, N14670);
and AND3 (N15837, N15817, N11476, N9650);
xor XOR2 (N15838, N15829, N4089);
nand NAND2 (N15839, N15814, N3938);
xor XOR2 (N15840, N15839, N4602);
xor XOR2 (N15841, N15836, N8196);
nor NOR3 (N15842, N15833, N8719, N2454);
nand NAND4 (N15843, N15838, N826, N14582, N5389);
buf BUF1 (N15844, N15835);
not NOT1 (N15845, N15844);
nand NAND2 (N15846, N15832, N581);
xor XOR2 (N15847, N15837, N143);
nand NAND3 (N15848, N15841, N638, N15116);
nor NOR4 (N15849, N15845, N11231, N6345, N11540);
nand NAND4 (N15850, N15831, N12408, N9080, N5957);
not NOT1 (N15851, N15848);
xor XOR2 (N15852, N15843, N4280);
and AND2 (N15853, N15849, N15699);
and AND4 (N15854, N15842, N9593, N11881, N14575);
not NOT1 (N15855, N15826);
not NOT1 (N15856, N15840);
nor NOR2 (N15857, N15853, N15146);
or OR4 (N15858, N15834, N3577, N6351, N11140);
buf BUF1 (N15859, N15850);
xor XOR2 (N15860, N15854, N6941);
nor NOR2 (N15861, N15851, N8972);
not NOT1 (N15862, N15857);
not NOT1 (N15863, N15858);
nand NAND2 (N15864, N15861, N10979);
and AND2 (N15865, N15863, N6102);
xor XOR2 (N15866, N15865, N10859);
nand NAND3 (N15867, N15859, N15222, N12630);
xor XOR2 (N15868, N15866, N1018);
nor NOR2 (N15869, N15852, N4519);
not NOT1 (N15870, N15867);
not NOT1 (N15871, N15862);
buf BUF1 (N15872, N15870);
not NOT1 (N15873, N15855);
and AND3 (N15874, N15860, N6027, N15648);
xor XOR2 (N15875, N15856, N3471);
or OR3 (N15876, N15869, N14556, N12952);
buf BUF1 (N15877, N15875);
nor NOR4 (N15878, N15847, N7325, N10505, N6084);
xor XOR2 (N15879, N15874, N3936);
and AND3 (N15880, N15872, N9474, N4622);
or OR4 (N15881, N15846, N13181, N4837, N14597);
not NOT1 (N15882, N15881);
buf BUF1 (N15883, N15873);
buf BUF1 (N15884, N15871);
xor XOR2 (N15885, N15877, N10034);
xor XOR2 (N15886, N15868, N7091);
nand NAND3 (N15887, N15884, N8804, N7134);
xor XOR2 (N15888, N15886, N7151);
buf BUF1 (N15889, N15876);
nor NOR4 (N15890, N15883, N7716, N287, N9397);
buf BUF1 (N15891, N15879);
or OR2 (N15892, N15885, N6558);
xor XOR2 (N15893, N15878, N8982);
or OR4 (N15894, N15893, N3935, N1057, N2507);
nand NAND2 (N15895, N15890, N430);
or OR2 (N15896, N15864, N12834);
and AND2 (N15897, N15891, N12608);
nand NAND2 (N15898, N15888, N3402);
not NOT1 (N15899, N15895);
or OR3 (N15900, N15899, N11276, N1343);
xor XOR2 (N15901, N15894, N7411);
xor XOR2 (N15902, N15900, N8675);
not NOT1 (N15903, N15902);
or OR3 (N15904, N15882, N14730, N3140);
xor XOR2 (N15905, N15889, N11953);
not NOT1 (N15906, N15898);
nor NOR3 (N15907, N15896, N9957, N9249);
buf BUF1 (N15908, N15907);
nand NAND4 (N15909, N15901, N15475, N12967, N4247);
nor NOR2 (N15910, N15906, N10569);
xor XOR2 (N15911, N15908, N3133);
and AND2 (N15912, N15892, N12722);
and AND2 (N15913, N15897, N3625);
or OR3 (N15914, N15905, N5868, N618);
xor XOR2 (N15915, N15911, N2913);
xor XOR2 (N15916, N15880, N8055);
and AND4 (N15917, N15887, N13373, N11019, N7721);
or OR2 (N15918, N15903, N3445);
xor XOR2 (N15919, N15904, N13887);
nand NAND3 (N15920, N15914, N7865, N8856);
or OR2 (N15921, N15916, N9085);
nor NOR3 (N15922, N15910, N5724, N9862);
xor XOR2 (N15923, N15912, N11561);
nor NOR3 (N15924, N15920, N10281, N9679);
xor XOR2 (N15925, N15921, N5174);
xor XOR2 (N15926, N15915, N2724);
and AND2 (N15927, N15909, N12257);
or OR3 (N15928, N15923, N12081, N2653);
buf BUF1 (N15929, N15919);
or OR3 (N15930, N15924, N7482, N9888);
and AND3 (N15931, N15922, N11814, N6060);
or OR3 (N15932, N15918, N3770, N4694);
nor NOR2 (N15933, N15928, N15240);
and AND3 (N15934, N15925, N10774, N13418);
not NOT1 (N15935, N15917);
nand NAND2 (N15936, N15927, N11280);
nor NOR2 (N15937, N15935, N13351);
nand NAND3 (N15938, N15937, N5188, N3602);
or OR2 (N15939, N15934, N5355);
nand NAND3 (N15940, N15913, N5122, N5476);
buf BUF1 (N15941, N15930);
and AND2 (N15942, N15929, N11629);
and AND4 (N15943, N15932, N10546, N7124, N10906);
nor NOR3 (N15944, N15943, N2551, N8515);
not NOT1 (N15945, N15936);
nor NOR3 (N15946, N15944, N8366, N1949);
buf BUF1 (N15947, N15939);
xor XOR2 (N15948, N15938, N7490);
nor NOR2 (N15949, N15941, N1981);
nor NOR3 (N15950, N15933, N14211, N14725);
nor NOR4 (N15951, N15945, N12856, N9327, N14940);
nor NOR4 (N15952, N15949, N5830, N6213, N4715);
and AND3 (N15953, N15940, N2419, N10246);
buf BUF1 (N15954, N15942);
not NOT1 (N15955, N15952);
nand NAND3 (N15956, N15951, N7146, N3271);
nor NOR3 (N15957, N15956, N5927, N14579);
xor XOR2 (N15958, N15950, N2426);
or OR2 (N15959, N15953, N8581);
buf BUF1 (N15960, N15954);
nand NAND4 (N15961, N15958, N14422, N7137, N7966);
xor XOR2 (N15962, N15947, N6859);
buf BUF1 (N15963, N15957);
nor NOR4 (N15964, N15960, N10459, N11644, N7781);
nand NAND4 (N15965, N15963, N9097, N11597, N7685);
nand NAND3 (N15966, N15962, N15033, N6275);
and AND4 (N15967, N15948, N11534, N4648, N13500);
not NOT1 (N15968, N15931);
nand NAND2 (N15969, N15968, N6485);
nand NAND4 (N15970, N15969, N637, N1783, N11662);
and AND2 (N15971, N15965, N13636);
xor XOR2 (N15972, N15967, N14385);
xor XOR2 (N15973, N15966, N5347);
or OR3 (N15974, N15946, N8984, N9438);
nor NOR3 (N15975, N15959, N4775, N5376);
or OR3 (N15976, N15975, N7556, N7867);
xor XOR2 (N15977, N15974, N1602);
buf BUF1 (N15978, N15976);
or OR2 (N15979, N15978, N1613);
buf BUF1 (N15980, N15955);
not NOT1 (N15981, N15971);
buf BUF1 (N15982, N15973);
xor XOR2 (N15983, N15961, N10290);
not NOT1 (N15984, N15982);
buf BUF1 (N15985, N15984);
not NOT1 (N15986, N15979);
or OR4 (N15987, N15980, N5141, N1504, N8532);
nand NAND3 (N15988, N15926, N13902, N13010);
nor NOR3 (N15989, N15964, N8789, N13739);
nor NOR4 (N15990, N15988, N1245, N8363, N15179);
not NOT1 (N15991, N15977);
nor NOR4 (N15992, N15990, N5226, N4980, N7202);
xor XOR2 (N15993, N15986, N7973);
buf BUF1 (N15994, N15992);
nor NOR2 (N15995, N15983, N12713);
xor XOR2 (N15996, N15987, N14345);
and AND3 (N15997, N15985, N13017, N9829);
nor NOR4 (N15998, N15995, N12814, N12273, N8272);
and AND3 (N15999, N15994, N2105, N8723);
buf BUF1 (N16000, N15989);
or OR2 (N16001, N15996, N5315);
xor XOR2 (N16002, N15998, N14880);
xor XOR2 (N16003, N15991, N10854);
nand NAND3 (N16004, N15999, N7065, N9645);
buf BUF1 (N16005, N16004);
xor XOR2 (N16006, N15981, N3231);
xor XOR2 (N16007, N16002, N11888);
nand NAND3 (N16008, N15972, N15761, N12638);
or OR2 (N16009, N16008, N2336);
or OR2 (N16010, N16006, N14150);
or OR2 (N16011, N16007, N874);
xor XOR2 (N16012, N15970, N684);
and AND2 (N16013, N16009, N6373);
and AND2 (N16014, N16012, N9463);
endmodule