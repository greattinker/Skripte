// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N806,N801,N809,N808,N804,N795,N794,N789,N807,N810;

nand NAND2 (N11, N4, N2);
buf BUF1 (N12, N11);
and AND3 (N13, N11, N6, N4);
nand NAND4 (N14, N5, N4, N4, N1);
buf BUF1 (N15, N6);
xor XOR2 (N16, N5, N3);
nand NAND4 (N17, N14, N1, N9, N10);
nor NOR2 (N18, N12, N11);
or OR3 (N19, N16, N13, N3);
or OR4 (N20, N4, N13, N12, N17);
xor XOR2 (N21, N3, N19);
buf BUF1 (N22, N14);
not NOT1 (N23, N18);
xor XOR2 (N24, N22, N18);
not NOT1 (N25, N14);
xor XOR2 (N26, N15, N8);
or OR4 (N27, N5, N25, N25, N20);
and AND3 (N28, N12, N21, N27);
buf BUF1 (N29, N24);
xor XOR2 (N30, N20, N1);
or OR4 (N31, N30, N9, N27, N28);
nor NOR3 (N32, N25, N28, N18);
nor NOR3 (N33, N28, N28, N14);
or OR2 (N34, N23, N24);
nor NOR3 (N35, N34, N4, N16);
xor XOR2 (N36, N10, N19);
buf BUF1 (N37, N34);
and AND4 (N38, N9, N26, N37, N13);
xor XOR2 (N39, N7, N36);
nor NOR4 (N40, N39, N32, N7, N23);
and AND3 (N41, N15, N2, N9);
and AND2 (N42, N35, N2);
nor NOR2 (N43, N10, N6);
nor NOR2 (N44, N13, N32);
not NOT1 (N45, N2);
nand NAND2 (N46, N45, N6);
not NOT1 (N47, N38);
xor XOR2 (N48, N44, N32);
xor XOR2 (N49, N40, N34);
nand NAND3 (N50, N43, N2, N32);
nand NAND2 (N51, N50, N49);
nor NOR3 (N52, N46, N24, N31);
buf BUF1 (N53, N27);
buf BUF1 (N54, N37);
buf BUF1 (N55, N42);
nand NAND4 (N56, N33, N35, N18, N30);
buf BUF1 (N57, N55);
nor NOR2 (N58, N54, N45);
or OR2 (N59, N48, N54);
or OR4 (N60, N41, N22, N27, N13);
nand NAND3 (N61, N56, N15, N25);
not NOT1 (N62, N53);
nand NAND3 (N63, N51, N35, N26);
nor NOR3 (N64, N29, N11, N37);
and AND2 (N65, N62, N8);
xor XOR2 (N66, N60, N21);
and AND3 (N67, N63, N25, N58);
or OR4 (N68, N31, N54, N52, N19);
not NOT1 (N69, N22);
not NOT1 (N70, N66);
nor NOR2 (N71, N69, N36);
buf BUF1 (N72, N59);
not NOT1 (N73, N64);
nand NAND3 (N74, N73, N67, N19);
nor NOR2 (N75, N5, N50);
and AND3 (N76, N74, N8, N15);
and AND2 (N77, N71, N14);
and AND3 (N78, N65, N53, N15);
nor NOR4 (N79, N77, N71, N45, N73);
not NOT1 (N80, N70);
and AND2 (N81, N75, N48);
or OR4 (N82, N78, N3, N41, N70);
not NOT1 (N83, N81);
and AND3 (N84, N57, N15, N56);
and AND3 (N85, N68, N60, N5);
not NOT1 (N86, N84);
or OR2 (N87, N47, N85);
or OR2 (N88, N63, N10);
and AND3 (N89, N87, N37, N83);
or OR2 (N90, N86, N60);
and AND3 (N91, N79, N88, N62);
buf BUF1 (N92, N43);
nor NOR2 (N93, N81, N11);
nand NAND2 (N94, N89, N81);
and AND4 (N95, N90, N49, N19, N93);
and AND2 (N96, N28, N78);
and AND4 (N97, N91, N35, N13, N70);
or OR2 (N98, N92, N63);
not NOT1 (N99, N61);
nor NOR4 (N100, N72, N77, N52, N31);
nand NAND2 (N101, N82, N85);
nand NAND2 (N102, N100, N70);
nand NAND2 (N103, N99, N18);
and AND3 (N104, N96, N81, N28);
xor XOR2 (N105, N102, N74);
buf BUF1 (N106, N105);
xor XOR2 (N107, N97, N2);
or OR3 (N108, N80, N72, N49);
nor NOR3 (N109, N108, N46, N90);
and AND4 (N110, N76, N24, N6, N8);
buf BUF1 (N111, N107);
xor XOR2 (N112, N94, N50);
buf BUF1 (N113, N112);
not NOT1 (N114, N113);
not NOT1 (N115, N106);
not NOT1 (N116, N115);
buf BUF1 (N117, N104);
and AND2 (N118, N110, N35);
or OR4 (N119, N95, N96, N71, N96);
nand NAND4 (N120, N119, N54, N41, N68);
buf BUF1 (N121, N101);
and AND3 (N122, N116, N23, N25);
xor XOR2 (N123, N114, N80);
or OR3 (N124, N121, N44, N30);
and AND3 (N125, N117, N13, N118);
not NOT1 (N126, N63);
buf BUF1 (N127, N109);
buf BUF1 (N128, N125);
nand NAND2 (N129, N98, N64);
not NOT1 (N130, N124);
buf BUF1 (N131, N103);
or OR2 (N132, N128, N77);
and AND2 (N133, N129, N103);
and AND2 (N134, N132, N53);
not NOT1 (N135, N126);
nand NAND2 (N136, N111, N89);
not NOT1 (N137, N127);
and AND2 (N138, N120, N77);
or OR4 (N139, N133, N58, N135, N124);
xor XOR2 (N140, N138, N69);
and AND4 (N141, N133, N103, N50, N46);
and AND3 (N142, N141, N2, N82);
buf BUF1 (N143, N136);
nand NAND4 (N144, N131, N68, N66, N141);
and AND3 (N145, N142, N29, N73);
or OR4 (N146, N143, N90, N88, N71);
nor NOR2 (N147, N140, N50);
or OR2 (N148, N122, N93);
xor XOR2 (N149, N148, N81);
or OR2 (N150, N149, N63);
nand NAND3 (N151, N144, N142, N113);
and AND3 (N152, N146, N81, N130);
nor NOR4 (N153, N116, N121, N81, N63);
and AND3 (N154, N150, N125, N24);
or OR2 (N155, N152, N104);
xor XOR2 (N156, N151, N15);
not NOT1 (N157, N145);
or OR4 (N158, N123, N30, N3, N136);
buf BUF1 (N159, N137);
buf BUF1 (N160, N154);
buf BUF1 (N161, N153);
xor XOR2 (N162, N160, N8);
and AND3 (N163, N158, N28, N64);
buf BUF1 (N164, N155);
xor XOR2 (N165, N164, N154);
nand NAND3 (N166, N139, N99, N118);
nor NOR4 (N167, N165, N139, N123, N117);
or OR3 (N168, N161, N69, N55);
nor NOR4 (N169, N156, N47, N125, N107);
not NOT1 (N170, N159);
not NOT1 (N171, N168);
not NOT1 (N172, N162);
not NOT1 (N173, N134);
buf BUF1 (N174, N147);
and AND3 (N175, N171, N93, N130);
nand NAND3 (N176, N173, N168, N38);
not NOT1 (N177, N170);
nand NAND4 (N178, N175, N28, N4, N21);
nand NAND3 (N179, N176, N144, N86);
and AND4 (N180, N179, N56, N123, N138);
xor XOR2 (N181, N180, N127);
buf BUF1 (N182, N172);
and AND3 (N183, N169, N96, N31);
xor XOR2 (N184, N178, N88);
nor NOR4 (N185, N182, N52, N31, N67);
not NOT1 (N186, N183);
nand NAND4 (N187, N163, N77, N176, N46);
not NOT1 (N188, N157);
nor NOR4 (N189, N166, N43, N101, N51);
nor NOR3 (N190, N174, N106, N111);
buf BUF1 (N191, N188);
nand NAND3 (N192, N189, N69, N75);
or OR4 (N193, N186, N23, N147, N86);
xor XOR2 (N194, N177, N4);
nand NAND3 (N195, N194, N99, N121);
xor XOR2 (N196, N193, N137);
not NOT1 (N197, N192);
and AND3 (N198, N181, N3, N24);
and AND2 (N199, N167, N67);
and AND3 (N200, N190, N37, N181);
buf BUF1 (N201, N185);
nor NOR4 (N202, N197, N87, N22, N89);
not NOT1 (N203, N201);
nor NOR3 (N204, N195, N182, N14);
buf BUF1 (N205, N191);
nor NOR3 (N206, N204, N147, N76);
and AND4 (N207, N198, N27, N110, N199);
or OR3 (N208, N152, N160, N120);
buf BUF1 (N209, N202);
not NOT1 (N210, N203);
or OR2 (N211, N210, N134);
nor NOR2 (N212, N207, N205);
and AND4 (N213, N84, N17, N134, N73);
not NOT1 (N214, N209);
xor XOR2 (N215, N208, N196);
xor XOR2 (N216, N174, N12);
or OR3 (N217, N184, N197, N100);
xor XOR2 (N218, N211, N65);
xor XOR2 (N219, N212, N176);
buf BUF1 (N220, N206);
xor XOR2 (N221, N216, N209);
xor XOR2 (N222, N218, N109);
buf BUF1 (N223, N220);
not NOT1 (N224, N223);
or OR2 (N225, N213, N203);
xor XOR2 (N226, N217, N216);
buf BUF1 (N227, N226);
and AND3 (N228, N214, N220, N120);
or OR3 (N229, N221, N198, N105);
buf BUF1 (N230, N200);
not NOT1 (N231, N228);
not NOT1 (N232, N187);
and AND4 (N233, N224, N64, N23, N205);
not NOT1 (N234, N225);
and AND3 (N235, N234, N51, N4);
not NOT1 (N236, N231);
nand NAND4 (N237, N229, N203, N63, N57);
buf BUF1 (N238, N233);
buf BUF1 (N239, N237);
and AND3 (N240, N236, N27, N42);
nand NAND2 (N241, N227, N153);
nor NOR2 (N242, N235, N195);
buf BUF1 (N243, N215);
buf BUF1 (N244, N241);
xor XOR2 (N245, N239, N64);
xor XOR2 (N246, N243, N77);
not NOT1 (N247, N222);
xor XOR2 (N248, N245, N235);
and AND4 (N249, N248, N91, N177, N79);
nand NAND2 (N250, N238, N29);
xor XOR2 (N251, N232, N86);
xor XOR2 (N252, N242, N70);
buf BUF1 (N253, N251);
nand NAND2 (N254, N244, N123);
not NOT1 (N255, N230);
nand NAND3 (N256, N255, N71, N75);
nand NAND4 (N257, N240, N181, N241, N89);
not NOT1 (N258, N257);
xor XOR2 (N259, N256, N6);
nor NOR2 (N260, N219, N147);
and AND4 (N261, N260, N74, N134, N181);
nand NAND4 (N262, N254, N109, N186, N252);
not NOT1 (N263, N13);
buf BUF1 (N264, N247);
nor NOR2 (N265, N258, N231);
or OR3 (N266, N250, N31, N22);
buf BUF1 (N267, N262);
not NOT1 (N268, N259);
nand NAND4 (N269, N267, N139, N187, N247);
and AND2 (N270, N265, N91);
nor NOR2 (N271, N253, N131);
nor NOR2 (N272, N270, N231);
not NOT1 (N273, N268);
nand NAND3 (N274, N269, N21, N78);
not NOT1 (N275, N266);
and AND2 (N276, N264, N171);
not NOT1 (N277, N263);
nand NAND3 (N278, N273, N11, N85);
xor XOR2 (N279, N261, N167);
nand NAND2 (N280, N278, N21);
not NOT1 (N281, N271);
or OR3 (N282, N274, N211, N264);
or OR4 (N283, N249, N98, N117, N104);
buf BUF1 (N284, N280);
xor XOR2 (N285, N277, N210);
not NOT1 (N286, N284);
buf BUF1 (N287, N279);
not NOT1 (N288, N285);
buf BUF1 (N289, N276);
not NOT1 (N290, N288);
and AND4 (N291, N246, N235, N155, N261);
not NOT1 (N292, N287);
buf BUF1 (N293, N282);
xor XOR2 (N294, N281, N183);
not NOT1 (N295, N286);
nand NAND4 (N296, N275, N276, N32, N22);
xor XOR2 (N297, N272, N232);
or OR2 (N298, N292, N105);
nand NAND2 (N299, N283, N42);
nand NAND3 (N300, N294, N279, N171);
not NOT1 (N301, N297);
buf BUF1 (N302, N300);
buf BUF1 (N303, N293);
xor XOR2 (N304, N295, N78);
nand NAND2 (N305, N304, N59);
nor NOR3 (N306, N305, N193, N121);
not NOT1 (N307, N303);
or OR3 (N308, N302, N212, N274);
xor XOR2 (N309, N296, N292);
xor XOR2 (N310, N306, N85);
or OR3 (N311, N299, N59, N170);
nor NOR3 (N312, N298, N21, N67);
buf BUF1 (N313, N289);
buf BUF1 (N314, N291);
not NOT1 (N315, N309);
not NOT1 (N316, N308);
nor NOR2 (N317, N315, N178);
nor NOR4 (N318, N317, N202, N166, N311);
and AND3 (N319, N137, N78, N273);
nor NOR2 (N320, N301, N236);
and AND3 (N321, N310, N45, N191);
nor NOR4 (N322, N307, N196, N227, N50);
or OR4 (N323, N316, N42, N43, N160);
nor NOR2 (N324, N290, N305);
xor XOR2 (N325, N314, N116);
buf BUF1 (N326, N324);
and AND2 (N327, N312, N237);
xor XOR2 (N328, N325, N277);
buf BUF1 (N329, N326);
and AND3 (N330, N327, N102, N235);
and AND3 (N331, N321, N244, N157);
or OR2 (N332, N320, N258);
buf BUF1 (N333, N329);
buf BUF1 (N334, N330);
and AND3 (N335, N323, N162, N1);
or OR3 (N336, N331, N268, N286);
nand NAND4 (N337, N313, N95, N239, N155);
or OR4 (N338, N333, N218, N297, N298);
not NOT1 (N339, N334);
and AND3 (N340, N332, N278, N274);
not NOT1 (N341, N328);
xor XOR2 (N342, N340, N325);
xor XOR2 (N343, N338, N324);
or OR2 (N344, N339, N234);
not NOT1 (N345, N342);
and AND2 (N346, N344, N78);
not NOT1 (N347, N319);
nor NOR4 (N348, N343, N319, N130, N84);
xor XOR2 (N349, N348, N101);
nor NOR3 (N350, N336, N137, N175);
xor XOR2 (N351, N337, N49);
or OR2 (N352, N322, N24);
nand NAND2 (N353, N350, N317);
nor NOR2 (N354, N349, N293);
buf BUF1 (N355, N341);
or OR3 (N356, N345, N76, N120);
buf BUF1 (N357, N335);
xor XOR2 (N358, N353, N303);
xor XOR2 (N359, N357, N105);
nand NAND3 (N360, N346, N6, N6);
xor XOR2 (N361, N360, N326);
and AND4 (N362, N351, N52, N290, N329);
not NOT1 (N363, N359);
not NOT1 (N364, N354);
buf BUF1 (N365, N318);
nor NOR4 (N366, N356, N200, N273, N121);
buf BUF1 (N367, N365);
or OR3 (N368, N352, N115, N198);
not NOT1 (N369, N366);
nand NAND2 (N370, N361, N340);
and AND4 (N371, N368, N196, N356, N57);
nor NOR2 (N372, N347, N274);
or OR4 (N373, N362, N58, N6, N176);
and AND3 (N374, N367, N95, N278);
nand NAND4 (N375, N369, N161, N4, N353);
and AND4 (N376, N374, N14, N247, N28);
xor XOR2 (N377, N373, N15);
nand NAND2 (N378, N375, N366);
buf BUF1 (N379, N378);
xor XOR2 (N380, N370, N324);
or OR4 (N381, N372, N85, N97, N135);
not NOT1 (N382, N371);
and AND4 (N383, N380, N279, N194, N71);
nand NAND3 (N384, N355, N162, N96);
or OR3 (N385, N376, N106, N381);
buf BUF1 (N386, N358);
buf BUF1 (N387, N99);
buf BUF1 (N388, N377);
buf BUF1 (N389, N387);
xor XOR2 (N390, N363, N243);
or OR2 (N391, N379, N29);
not NOT1 (N392, N386);
nor NOR4 (N393, N391, N40, N385, N278);
xor XOR2 (N394, N34, N50);
or OR2 (N395, N388, N215);
xor XOR2 (N396, N395, N202);
not NOT1 (N397, N393);
xor XOR2 (N398, N382, N193);
or OR2 (N399, N390, N142);
not NOT1 (N400, N384);
or OR4 (N401, N383, N335, N19, N37);
not NOT1 (N402, N401);
nand NAND3 (N403, N396, N313, N6);
nand NAND2 (N404, N402, N315);
xor XOR2 (N405, N400, N148);
xor XOR2 (N406, N394, N163);
or OR2 (N407, N392, N183);
buf BUF1 (N408, N399);
not NOT1 (N409, N364);
and AND2 (N410, N406, N195);
or OR2 (N411, N398, N155);
buf BUF1 (N412, N405);
and AND2 (N413, N404, N66);
xor XOR2 (N414, N389, N198);
or OR3 (N415, N412, N16, N378);
buf BUF1 (N416, N413);
xor XOR2 (N417, N407, N172);
nor NOR2 (N418, N409, N297);
nor NOR3 (N419, N417, N330, N69);
and AND2 (N420, N408, N239);
or OR3 (N421, N410, N213, N126);
not NOT1 (N422, N420);
nand NAND3 (N423, N416, N287, N220);
nor NOR2 (N424, N422, N235);
not NOT1 (N425, N411);
and AND4 (N426, N403, N367, N69, N294);
and AND4 (N427, N414, N46, N80, N41);
nand NAND4 (N428, N415, N185, N53, N133);
xor XOR2 (N429, N427, N13);
nor NOR2 (N430, N418, N41);
or OR3 (N431, N421, N216, N144);
xor XOR2 (N432, N428, N215);
buf BUF1 (N433, N426);
buf BUF1 (N434, N433);
not NOT1 (N435, N425);
or OR2 (N436, N430, N2);
xor XOR2 (N437, N423, N247);
or OR4 (N438, N436, N203, N261, N423);
nor NOR2 (N439, N397, N322);
nand NAND2 (N440, N435, N158);
or OR3 (N441, N429, N5, N398);
nand NAND3 (N442, N431, N367, N82);
not NOT1 (N443, N441);
or OR2 (N444, N440, N405);
nand NAND2 (N445, N444, N343);
xor XOR2 (N446, N443, N316);
xor XOR2 (N447, N437, N19);
buf BUF1 (N448, N419);
not NOT1 (N449, N448);
buf BUF1 (N450, N434);
not NOT1 (N451, N445);
nand NAND2 (N452, N447, N213);
nand NAND2 (N453, N439, N447);
xor XOR2 (N454, N451, N73);
and AND4 (N455, N438, N141, N420, N232);
and AND2 (N456, N454, N102);
not NOT1 (N457, N450);
xor XOR2 (N458, N455, N102);
and AND3 (N459, N449, N405, N136);
or OR3 (N460, N459, N373, N390);
nand NAND3 (N461, N460, N336, N244);
xor XOR2 (N462, N457, N134);
not NOT1 (N463, N446);
xor XOR2 (N464, N456, N130);
nor NOR2 (N465, N442, N72);
nor NOR4 (N466, N453, N226, N15, N51);
nor NOR4 (N467, N458, N278, N172, N102);
nand NAND4 (N468, N467, N224, N110, N49);
xor XOR2 (N469, N432, N4);
or OR3 (N470, N466, N214, N201);
and AND2 (N471, N464, N413);
and AND2 (N472, N465, N217);
not NOT1 (N473, N463);
xor XOR2 (N474, N471, N170);
or OR3 (N475, N462, N281, N47);
nand NAND2 (N476, N470, N305);
buf BUF1 (N477, N452);
xor XOR2 (N478, N472, N374);
or OR3 (N479, N477, N154, N36);
buf BUF1 (N480, N478);
or OR3 (N481, N475, N100, N288);
nor NOR3 (N482, N476, N432, N316);
or OR2 (N483, N480, N456);
or OR3 (N484, N479, N81, N55);
or OR2 (N485, N469, N252);
not NOT1 (N486, N473);
or OR4 (N487, N482, N111, N82, N216);
nand NAND2 (N488, N486, N268);
and AND4 (N489, N474, N165, N392, N84);
nand NAND2 (N490, N461, N401);
buf BUF1 (N491, N488);
buf BUF1 (N492, N485);
nand NAND3 (N493, N491, N340, N249);
or OR2 (N494, N481, N240);
nor NOR2 (N495, N489, N44);
and AND4 (N496, N490, N25, N178, N341);
and AND4 (N497, N496, N278, N465, N173);
and AND3 (N498, N483, N487, N140);
nor NOR2 (N499, N415, N97);
nor NOR4 (N500, N495, N488, N298, N484);
not NOT1 (N501, N291);
nand NAND2 (N502, N501, N312);
nand NAND3 (N503, N493, N226, N372);
xor XOR2 (N504, N499, N221);
and AND4 (N505, N424, N277, N440, N354);
or OR3 (N506, N497, N70, N274);
xor XOR2 (N507, N492, N424);
xor XOR2 (N508, N506, N199);
xor XOR2 (N509, N502, N173);
buf BUF1 (N510, N509);
buf BUF1 (N511, N505);
not NOT1 (N512, N494);
buf BUF1 (N513, N500);
buf BUF1 (N514, N510);
or OR2 (N515, N508, N346);
nand NAND4 (N516, N512, N273, N371, N218);
xor XOR2 (N517, N507, N165);
and AND3 (N518, N517, N11, N148);
nand NAND4 (N519, N504, N348, N350, N508);
buf BUF1 (N520, N519);
buf BUF1 (N521, N516);
and AND2 (N522, N514, N206);
nor NOR3 (N523, N503, N327, N27);
not NOT1 (N524, N520);
nand NAND2 (N525, N521, N176);
nor NOR3 (N526, N513, N170, N100);
not NOT1 (N527, N526);
and AND3 (N528, N511, N314, N508);
and AND2 (N529, N522, N312);
and AND2 (N530, N468, N242);
xor XOR2 (N531, N518, N511);
nor NOR3 (N532, N523, N61, N187);
nor NOR4 (N533, N525, N303, N344, N285);
nor NOR2 (N534, N515, N70);
nand NAND4 (N535, N533, N429, N354, N44);
nor NOR3 (N536, N529, N304, N310);
buf BUF1 (N537, N536);
nor NOR2 (N538, N535, N308);
nor NOR3 (N539, N538, N375, N146);
nand NAND3 (N540, N532, N393, N294);
buf BUF1 (N541, N537);
xor XOR2 (N542, N498, N138);
and AND3 (N543, N534, N114, N129);
buf BUF1 (N544, N528);
or OR3 (N545, N544, N523, N371);
buf BUF1 (N546, N545);
nor NOR2 (N547, N541, N224);
nor NOR4 (N548, N530, N403, N167, N344);
not NOT1 (N549, N543);
not NOT1 (N550, N542);
or OR2 (N551, N549, N300);
and AND3 (N552, N547, N164, N499);
and AND2 (N553, N550, N455);
or OR2 (N554, N546, N205);
or OR3 (N555, N531, N533, N378);
nand NAND3 (N556, N553, N542, N379);
not NOT1 (N557, N554);
xor XOR2 (N558, N556, N226);
xor XOR2 (N559, N557, N460);
nand NAND2 (N560, N558, N114);
buf BUF1 (N561, N524);
nand NAND2 (N562, N551, N170);
or OR3 (N563, N540, N36, N494);
xor XOR2 (N564, N563, N29);
or OR4 (N565, N559, N46, N188, N432);
nand NAND4 (N566, N539, N304, N210, N469);
not NOT1 (N567, N548);
not NOT1 (N568, N527);
not NOT1 (N569, N561);
or OR4 (N570, N564, N558, N461, N74);
xor XOR2 (N571, N569, N416);
or OR2 (N572, N571, N101);
and AND2 (N573, N555, N11);
nor NOR3 (N574, N562, N105, N3);
nand NAND4 (N575, N552, N116, N123, N172);
buf BUF1 (N576, N572);
not NOT1 (N577, N573);
or OR2 (N578, N565, N122);
xor XOR2 (N579, N574, N73);
xor XOR2 (N580, N576, N226);
xor XOR2 (N581, N570, N158);
nand NAND2 (N582, N581, N103);
not NOT1 (N583, N577);
nand NAND4 (N584, N575, N559, N191, N293);
xor XOR2 (N585, N583, N234);
nor NOR4 (N586, N584, N156, N568, N139);
or OR2 (N587, N246, N528);
not NOT1 (N588, N585);
not NOT1 (N589, N586);
or OR3 (N590, N578, N416, N434);
nor NOR3 (N591, N588, N550, N538);
nand NAND3 (N592, N579, N101, N370);
nand NAND3 (N593, N567, N337, N585);
nand NAND2 (N594, N591, N526);
buf BUF1 (N595, N560);
nand NAND4 (N596, N593, N111, N445, N480);
and AND4 (N597, N590, N394, N146, N235);
buf BUF1 (N598, N597);
buf BUF1 (N599, N582);
or OR3 (N600, N599, N305, N328);
or OR3 (N601, N600, N36, N483);
xor XOR2 (N602, N595, N335);
buf BUF1 (N603, N601);
xor XOR2 (N604, N580, N83);
nor NOR2 (N605, N566, N445);
buf BUF1 (N606, N589);
xor XOR2 (N607, N606, N175);
not NOT1 (N608, N594);
not NOT1 (N609, N592);
buf BUF1 (N610, N605);
or OR4 (N611, N610, N246, N59, N415);
buf BUF1 (N612, N603);
xor XOR2 (N613, N611, N357);
and AND3 (N614, N604, N49, N395);
and AND3 (N615, N602, N282, N436);
buf BUF1 (N616, N615);
nand NAND3 (N617, N613, N203, N441);
not NOT1 (N618, N608);
and AND3 (N619, N617, N612, N457);
or OR3 (N620, N182, N149, N185);
or OR3 (N621, N616, N17, N197);
and AND3 (N622, N607, N346, N413);
xor XOR2 (N623, N587, N591);
and AND3 (N624, N614, N408, N217);
and AND4 (N625, N622, N472, N217, N350);
not NOT1 (N626, N623);
buf BUF1 (N627, N596);
buf BUF1 (N628, N625);
not NOT1 (N629, N609);
and AND2 (N630, N626, N410);
nor NOR4 (N631, N620, N12, N566, N153);
and AND2 (N632, N630, N471);
and AND4 (N633, N627, N247, N531, N24);
nand NAND2 (N634, N619, N298);
and AND2 (N635, N618, N49);
nand NAND2 (N636, N621, N383);
not NOT1 (N637, N634);
xor XOR2 (N638, N635, N318);
nor NOR3 (N639, N632, N256, N505);
nand NAND3 (N640, N629, N373, N55);
xor XOR2 (N641, N628, N120);
or OR2 (N642, N637, N511);
xor XOR2 (N643, N624, N110);
nor NOR3 (N644, N640, N234, N268);
nand NAND2 (N645, N641, N12);
xor XOR2 (N646, N644, N211);
buf BUF1 (N647, N636);
not NOT1 (N648, N645);
nand NAND3 (N649, N648, N363, N130);
and AND4 (N650, N598, N91, N200, N462);
not NOT1 (N651, N643);
xor XOR2 (N652, N647, N391);
nor NOR4 (N653, N651, N423, N357, N507);
xor XOR2 (N654, N631, N613);
nand NAND3 (N655, N653, N465, N206);
nor NOR3 (N656, N649, N162, N446);
nand NAND4 (N657, N638, N465, N602, N285);
xor XOR2 (N658, N656, N435);
and AND4 (N659, N652, N622, N33, N335);
or OR2 (N660, N639, N64);
xor XOR2 (N661, N650, N194);
or OR4 (N662, N646, N212, N8, N638);
and AND4 (N663, N642, N626, N44, N7);
xor XOR2 (N664, N663, N206);
nand NAND2 (N665, N655, N553);
not NOT1 (N666, N660);
nand NAND4 (N667, N662, N129, N74, N200);
nand NAND2 (N668, N667, N396);
not NOT1 (N669, N665);
or OR4 (N670, N657, N405, N255, N162);
nor NOR4 (N671, N670, N360, N211, N282);
or OR3 (N672, N664, N418, N118);
not NOT1 (N673, N669);
not NOT1 (N674, N672);
xor XOR2 (N675, N661, N392);
not NOT1 (N676, N666);
nor NOR3 (N677, N676, N115, N540);
buf BUF1 (N678, N654);
buf BUF1 (N679, N668);
or OR3 (N680, N673, N397, N527);
nand NAND3 (N681, N633, N200, N22);
and AND3 (N682, N658, N487, N409);
or OR3 (N683, N680, N251, N354);
nand NAND3 (N684, N681, N573, N307);
nand NAND2 (N685, N682, N104);
xor XOR2 (N686, N684, N680);
or OR2 (N687, N675, N169);
or OR4 (N688, N677, N178, N84, N486);
nand NAND3 (N689, N671, N591, N181);
or OR2 (N690, N674, N396);
xor XOR2 (N691, N687, N159);
or OR2 (N692, N659, N617);
nor NOR2 (N693, N683, N528);
xor XOR2 (N694, N686, N225);
xor XOR2 (N695, N693, N115);
or OR2 (N696, N678, N521);
xor XOR2 (N697, N689, N458);
buf BUF1 (N698, N688);
nand NAND2 (N699, N698, N71);
xor XOR2 (N700, N690, N393);
nor NOR4 (N701, N697, N51, N394, N72);
or OR4 (N702, N696, N20, N576, N665);
buf BUF1 (N703, N695);
nor NOR4 (N704, N702, N224, N107, N463);
xor XOR2 (N705, N700, N191);
not NOT1 (N706, N701);
nor NOR3 (N707, N704, N466, N16);
nand NAND3 (N708, N685, N696, N349);
not NOT1 (N709, N705);
nor NOR3 (N710, N679, N124, N268);
or OR2 (N711, N699, N332);
or OR4 (N712, N709, N4, N158, N42);
or OR4 (N713, N706, N588, N430, N641);
nor NOR4 (N714, N713, N559, N450, N151);
nand NAND2 (N715, N707, N58);
nand NAND2 (N716, N692, N578);
and AND4 (N717, N691, N218, N236, N458);
nor NOR2 (N718, N694, N536);
or OR2 (N719, N712, N331);
xor XOR2 (N720, N716, N526);
nor NOR3 (N721, N711, N706, N620);
nor NOR3 (N722, N718, N119, N466);
buf BUF1 (N723, N717);
nand NAND2 (N724, N715, N277);
or OR2 (N725, N710, N5);
nand NAND2 (N726, N724, N436);
xor XOR2 (N727, N719, N297);
nand NAND3 (N728, N723, N39, N724);
and AND3 (N729, N714, N233, N607);
nand NAND3 (N730, N708, N521, N48);
nor NOR3 (N731, N703, N620, N325);
nand NAND4 (N732, N729, N211, N543, N641);
and AND4 (N733, N720, N263, N696, N399);
or OR4 (N734, N727, N519, N676, N396);
nand NAND4 (N735, N722, N490, N682, N74);
xor XOR2 (N736, N731, N78);
and AND2 (N737, N730, N683);
nor NOR3 (N738, N721, N655, N267);
not NOT1 (N739, N728);
or OR2 (N740, N739, N378);
or OR2 (N741, N738, N493);
or OR2 (N742, N740, N303);
nand NAND2 (N743, N737, N60);
xor XOR2 (N744, N743, N169);
buf BUF1 (N745, N732);
xor XOR2 (N746, N745, N536);
buf BUF1 (N747, N735);
not NOT1 (N748, N733);
and AND4 (N749, N747, N585, N516, N208);
and AND4 (N750, N741, N707, N345, N609);
nand NAND3 (N751, N734, N164, N85);
buf BUF1 (N752, N746);
xor XOR2 (N753, N749, N109);
or OR4 (N754, N752, N80, N522, N493);
or OR2 (N755, N753, N553);
or OR3 (N756, N742, N34, N219);
xor XOR2 (N757, N736, N653);
and AND3 (N758, N726, N612, N119);
xor XOR2 (N759, N758, N436);
xor XOR2 (N760, N725, N51);
and AND3 (N761, N757, N211, N508);
nor NOR4 (N762, N750, N390, N354, N755);
nand NAND3 (N763, N394, N318, N673);
and AND3 (N764, N748, N182, N326);
not NOT1 (N765, N759);
or OR2 (N766, N751, N587);
xor XOR2 (N767, N754, N598);
not NOT1 (N768, N744);
buf BUF1 (N769, N762);
nor NOR2 (N770, N756, N190);
buf BUF1 (N771, N769);
or OR4 (N772, N766, N396, N34, N75);
xor XOR2 (N773, N767, N128);
xor XOR2 (N774, N763, N161);
or OR4 (N775, N768, N556, N581, N436);
or OR4 (N776, N775, N192, N375, N423);
nand NAND3 (N777, N772, N146, N589);
xor XOR2 (N778, N771, N762);
and AND4 (N779, N770, N113, N712, N778);
or OR4 (N780, N91, N94, N191, N449);
and AND4 (N781, N773, N735, N750, N519);
buf BUF1 (N782, N780);
buf BUF1 (N783, N764);
buf BUF1 (N784, N761);
buf BUF1 (N785, N777);
and AND4 (N786, N760, N14, N146, N668);
nand NAND2 (N787, N785, N129);
not NOT1 (N788, N765);
buf BUF1 (N789, N782);
and AND3 (N790, N781, N72, N254);
nor NOR4 (N791, N779, N15, N724, N677);
or OR4 (N792, N783, N321, N484, N697);
not NOT1 (N793, N786);
or OR2 (N794, N776, N216);
not NOT1 (N795, N788);
and AND2 (N796, N793, N21);
not NOT1 (N797, N774);
nor NOR2 (N798, N787, N567);
buf BUF1 (N799, N797);
or OR3 (N800, N798, N762, N757);
nor NOR3 (N801, N796, N178, N505);
buf BUF1 (N802, N792);
xor XOR2 (N803, N790, N542);
nor NOR2 (N804, N784, N405);
or OR3 (N805, N803, N422, N764);
nand NAND3 (N806, N791, N246, N8);
nand NAND3 (N807, N799, N602, N231);
not NOT1 (N808, N800);
nor NOR2 (N809, N805, N703);
xor XOR2 (N810, N802, N785);
endmodule