// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N2521,N2485,N2516,N2517,N2518,N2523,N2514,N2473,N2522,N2524;

buf BUF1 (N25, N7);
or OR4 (N26, N23, N24, N16, N10);
nor NOR3 (N27, N25, N22, N11);
and AND3 (N28, N5, N20, N1);
buf BUF1 (N29, N9);
nor NOR4 (N30, N16, N15, N7, N21);
buf BUF1 (N31, N19);
not NOT1 (N32, N1);
nor NOR4 (N33, N2, N2, N27, N10);
xor XOR2 (N34, N32, N6);
and AND2 (N35, N33, N18);
not NOT1 (N36, N29);
or OR2 (N37, N35, N36);
buf BUF1 (N38, N17);
nor NOR4 (N39, N18, N12, N6, N26);
xor XOR2 (N40, N21, N23);
not NOT1 (N41, N4);
nor NOR4 (N42, N39, N8, N31, N34);
buf BUF1 (N43, N21);
buf BUF1 (N44, N30);
and AND3 (N45, N7, N43, N32);
and AND4 (N46, N37, N36, N30, N14);
and AND3 (N47, N20, N19, N46);
xor XOR2 (N48, N27, N36);
not NOT1 (N49, N17);
xor XOR2 (N50, N41, N36);
buf BUF1 (N51, N47);
buf BUF1 (N52, N40);
not NOT1 (N53, N42);
nor NOR2 (N54, N44, N26);
nand NAND3 (N55, N50, N34, N29);
nand NAND4 (N56, N52, N22, N16, N11);
buf BUF1 (N57, N54);
or OR3 (N58, N56, N32, N46);
or OR3 (N59, N45, N36, N31);
and AND4 (N60, N48, N42, N46, N18);
not NOT1 (N61, N60);
not NOT1 (N62, N58);
or OR4 (N63, N38, N8, N27, N58);
or OR3 (N64, N57, N4, N42);
or OR4 (N65, N64, N30, N50, N44);
not NOT1 (N66, N49);
buf BUF1 (N67, N28);
nand NAND4 (N68, N61, N26, N21, N29);
not NOT1 (N69, N68);
xor XOR2 (N70, N66, N15);
nor NOR4 (N71, N51, N18, N27, N10);
or OR3 (N72, N69, N7, N10);
xor XOR2 (N73, N63, N63);
and AND4 (N74, N72, N68, N14, N68);
buf BUF1 (N75, N73);
and AND4 (N76, N74, N49, N5, N50);
nor NOR4 (N77, N70, N38, N29, N71);
xor XOR2 (N78, N50, N68);
not NOT1 (N79, N76);
nor NOR2 (N80, N67, N37);
and AND3 (N81, N77, N57, N80);
nand NAND3 (N82, N45, N55, N51);
not NOT1 (N83, N5);
nor NOR4 (N84, N78, N81, N18, N56);
nor NOR3 (N85, N69, N6, N72);
not NOT1 (N86, N84);
nor NOR3 (N87, N86, N31, N51);
not NOT1 (N88, N79);
nor NOR3 (N89, N75, N42, N1);
nor NOR3 (N90, N83, N62, N73);
or OR2 (N91, N27, N12);
nor NOR2 (N92, N87, N71);
buf BUF1 (N93, N82);
nand NAND3 (N94, N92, N24, N40);
nand NAND3 (N95, N85, N39, N78);
or OR3 (N96, N53, N76, N12);
not NOT1 (N97, N90);
not NOT1 (N98, N95);
buf BUF1 (N99, N65);
nor NOR4 (N100, N97, N10, N30, N9);
buf BUF1 (N101, N88);
nand NAND4 (N102, N94, N7, N26, N68);
xor XOR2 (N103, N100, N51);
nor NOR3 (N104, N96, N63, N14);
nand NAND2 (N105, N91, N49);
buf BUF1 (N106, N101);
xor XOR2 (N107, N103, N100);
and AND4 (N108, N106, N20, N107, N67);
not NOT1 (N109, N24);
buf BUF1 (N110, N98);
nand NAND4 (N111, N108, N1, N87, N76);
and AND3 (N112, N89, N82, N34);
not NOT1 (N113, N111);
not NOT1 (N114, N112);
nor NOR3 (N115, N102, N32, N107);
buf BUF1 (N116, N113);
nand NAND4 (N117, N59, N114, N12, N84);
and AND2 (N118, N11, N108);
nand NAND4 (N119, N116, N86, N19, N105);
buf BUF1 (N120, N55);
or OR2 (N121, N117, N95);
xor XOR2 (N122, N120, N67);
not NOT1 (N123, N121);
nor NOR4 (N124, N110, N49, N57, N12);
nand NAND4 (N125, N123, N92, N59, N20);
or OR3 (N126, N93, N120, N43);
xor XOR2 (N127, N126, N109);
buf BUF1 (N128, N113);
and AND2 (N129, N115, N28);
nor NOR3 (N130, N119, N20, N101);
or OR2 (N131, N130, N78);
nor NOR3 (N132, N122, N130, N11);
nor NOR4 (N133, N124, N36, N66, N48);
xor XOR2 (N134, N127, N22);
not NOT1 (N135, N129);
and AND3 (N136, N99, N27, N109);
buf BUF1 (N137, N125);
or OR3 (N138, N136, N128, N15);
buf BUF1 (N139, N127);
buf BUF1 (N140, N134);
and AND4 (N141, N135, N104, N55, N138);
not NOT1 (N142, N10);
buf BUF1 (N143, N100);
buf BUF1 (N144, N118);
or OR3 (N145, N131, N67, N77);
or OR4 (N146, N141, N34, N141, N140);
nand NAND3 (N147, N52, N65, N5);
nand NAND2 (N148, N145, N140);
or OR4 (N149, N144, N108, N58, N38);
nand NAND2 (N150, N146, N70);
not NOT1 (N151, N143);
and AND2 (N152, N148, N73);
nand NAND3 (N153, N137, N74, N133);
and AND2 (N154, N63, N40);
or OR2 (N155, N147, N97);
not NOT1 (N156, N132);
nand NAND4 (N157, N139, N32, N90, N57);
not NOT1 (N158, N149);
not NOT1 (N159, N153);
xor XOR2 (N160, N157, N140);
xor XOR2 (N161, N155, N127);
xor XOR2 (N162, N142, N48);
or OR3 (N163, N158, N94, N38);
nor NOR2 (N164, N162, N99);
or OR2 (N165, N152, N24);
xor XOR2 (N166, N159, N22);
buf BUF1 (N167, N150);
xor XOR2 (N168, N164, N155);
xor XOR2 (N169, N156, N17);
buf BUF1 (N170, N167);
or OR4 (N171, N151, N33, N39, N60);
nand NAND4 (N172, N160, N12, N37, N50);
not NOT1 (N173, N165);
buf BUF1 (N174, N166);
nand NAND3 (N175, N173, N165, N107);
not NOT1 (N176, N175);
buf BUF1 (N177, N154);
nand NAND2 (N178, N161, N3);
or OR4 (N179, N169, N13, N37, N81);
not NOT1 (N180, N176);
not NOT1 (N181, N177);
nand NAND4 (N182, N163, N99, N101, N131);
or OR3 (N183, N181, N132, N82);
xor XOR2 (N184, N172, N87);
xor XOR2 (N185, N179, N151);
nand NAND4 (N186, N180, N172, N35, N60);
or OR3 (N187, N183, N36, N68);
nand NAND2 (N188, N170, N17);
or OR4 (N189, N168, N4, N186, N35);
nor NOR3 (N190, N152, N103, N74);
buf BUF1 (N191, N189);
not NOT1 (N192, N190);
nand NAND3 (N193, N182, N14, N184);
or OR4 (N194, N9, N167, N7, N9);
and AND4 (N195, N191, N41, N96, N116);
not NOT1 (N196, N171);
xor XOR2 (N197, N185, N112);
or OR4 (N198, N187, N149, N194, N189);
buf BUF1 (N199, N60);
or OR2 (N200, N196, N54);
and AND3 (N201, N192, N54, N190);
nand NAND2 (N202, N178, N182);
and AND2 (N203, N193, N71);
and AND4 (N204, N195, N90, N68, N50);
nor NOR4 (N205, N200, N18, N202, N20);
or OR3 (N206, N8, N184, N133);
buf BUF1 (N207, N188);
xor XOR2 (N208, N174, N157);
buf BUF1 (N209, N198);
buf BUF1 (N210, N208);
not NOT1 (N211, N209);
not NOT1 (N212, N205);
buf BUF1 (N213, N201);
not NOT1 (N214, N211);
not NOT1 (N215, N212);
not NOT1 (N216, N213);
nor NOR4 (N217, N206, N199, N25, N175);
buf BUF1 (N218, N172);
nor NOR2 (N219, N203, N146);
nand NAND4 (N220, N210, N96, N218, N138);
and AND3 (N221, N136, N163, N188);
nor NOR2 (N222, N197, N130);
xor XOR2 (N223, N219, N91);
xor XOR2 (N224, N223, N25);
nand NAND4 (N225, N204, N118, N123, N95);
or OR2 (N226, N224, N184);
nor NOR3 (N227, N207, N144, N12);
or OR4 (N228, N220, N9, N82, N54);
buf BUF1 (N229, N215);
xor XOR2 (N230, N222, N84);
xor XOR2 (N231, N229, N228);
or OR2 (N232, N38, N218);
xor XOR2 (N233, N214, N184);
nand NAND4 (N234, N217, N67, N19, N164);
xor XOR2 (N235, N227, N78);
nand NAND4 (N236, N232, N60, N85, N15);
nand NAND4 (N237, N216, N185, N107, N3);
buf BUF1 (N238, N230);
nor NOR3 (N239, N234, N203, N207);
nand NAND3 (N240, N226, N93, N167);
nand NAND3 (N241, N237, N194, N211);
nor NOR4 (N242, N240, N139, N134, N50);
and AND3 (N243, N221, N34, N80);
nand NAND2 (N244, N243, N7);
buf BUF1 (N245, N239);
xor XOR2 (N246, N225, N32);
not NOT1 (N247, N241);
and AND2 (N248, N246, N111);
buf BUF1 (N249, N231);
nand NAND3 (N250, N249, N128, N195);
nand NAND4 (N251, N244, N41, N23, N107);
nor NOR4 (N252, N235, N202, N93, N25);
and AND2 (N253, N248, N63);
nor NOR3 (N254, N242, N177, N151);
not NOT1 (N255, N233);
nand NAND3 (N256, N255, N6, N30);
and AND4 (N257, N251, N189, N141, N215);
or OR2 (N258, N257, N227);
xor XOR2 (N259, N238, N71);
buf BUF1 (N260, N252);
nor NOR3 (N261, N247, N34, N199);
not NOT1 (N262, N245);
xor XOR2 (N263, N260, N158);
xor XOR2 (N264, N258, N41);
xor XOR2 (N265, N256, N206);
nor NOR4 (N266, N263, N40, N51, N260);
and AND4 (N267, N265, N116, N235, N4);
or OR4 (N268, N264, N226, N11, N74);
nor NOR4 (N269, N267, N50, N73, N4);
xor XOR2 (N270, N253, N183);
buf BUF1 (N271, N268);
or OR3 (N272, N259, N135, N258);
not NOT1 (N273, N271);
or OR2 (N274, N254, N177);
or OR3 (N275, N266, N61, N14);
or OR4 (N276, N270, N80, N189, N195);
nor NOR4 (N277, N236, N136, N10, N194);
nand NAND4 (N278, N276, N61, N247, N225);
or OR3 (N279, N275, N22, N29);
and AND2 (N280, N250, N226);
xor XOR2 (N281, N280, N272);
or OR3 (N282, N94, N278, N214);
buf BUF1 (N283, N23);
not NOT1 (N284, N277);
nand NAND2 (N285, N262, N270);
xor XOR2 (N286, N282, N182);
or OR2 (N287, N285, N108);
buf BUF1 (N288, N269);
nand NAND4 (N289, N284, N80, N166, N236);
not NOT1 (N290, N261);
not NOT1 (N291, N287);
nand NAND3 (N292, N283, N194, N4);
and AND3 (N293, N274, N53, N68);
and AND2 (N294, N288, N43);
xor XOR2 (N295, N279, N172);
buf BUF1 (N296, N294);
and AND2 (N297, N296, N231);
not NOT1 (N298, N290);
and AND3 (N299, N286, N183, N197);
xor XOR2 (N300, N298, N35);
nor NOR2 (N301, N281, N110);
and AND4 (N302, N299, N36, N297, N131);
xor XOR2 (N303, N117, N46);
nor NOR4 (N304, N289, N279, N93, N151);
xor XOR2 (N305, N302, N236);
xor XOR2 (N306, N291, N231);
not NOT1 (N307, N301);
not NOT1 (N308, N303);
or OR3 (N309, N308, N163, N199);
xor XOR2 (N310, N300, N235);
and AND2 (N311, N307, N68);
nand NAND3 (N312, N293, N142, N251);
nor NOR4 (N313, N306, N312, N199, N255);
or OR2 (N314, N192, N268);
and AND2 (N315, N309, N167);
xor XOR2 (N316, N311, N280);
nor NOR3 (N317, N316, N31, N61);
and AND3 (N318, N292, N256, N129);
not NOT1 (N319, N315);
or OR2 (N320, N318, N183);
nor NOR2 (N321, N310, N283);
xor XOR2 (N322, N320, N221);
xor XOR2 (N323, N322, N147);
nand NAND3 (N324, N304, N179, N160);
and AND3 (N325, N305, N107, N170);
not NOT1 (N326, N323);
buf BUF1 (N327, N321);
xor XOR2 (N328, N295, N265);
xor XOR2 (N329, N314, N161);
or OR4 (N330, N324, N325, N117, N177);
not NOT1 (N331, N308);
not NOT1 (N332, N326);
nor NOR3 (N333, N331, N276, N257);
nand NAND3 (N334, N330, N73, N165);
xor XOR2 (N335, N329, N255);
nand NAND2 (N336, N313, N156);
nand NAND4 (N337, N333, N13, N287, N116);
or OR4 (N338, N335, N333, N166, N198);
nor NOR4 (N339, N273, N253, N51, N242);
nor NOR3 (N340, N338, N219, N256);
nor NOR2 (N341, N339, N337);
not NOT1 (N342, N186);
not NOT1 (N343, N319);
nor NOR2 (N344, N336, N54);
not NOT1 (N345, N340);
or OR3 (N346, N345, N240, N201);
or OR3 (N347, N332, N190, N280);
or OR2 (N348, N347, N278);
not NOT1 (N349, N348);
xor XOR2 (N350, N342, N110);
and AND4 (N351, N334, N207, N304, N71);
nor NOR4 (N352, N343, N7, N306, N196);
nor NOR2 (N353, N341, N231);
nand NAND4 (N354, N327, N156, N176, N168);
and AND4 (N355, N328, N16, N115, N30);
and AND4 (N356, N350, N344, N93, N171);
and AND3 (N357, N57, N55, N205);
xor XOR2 (N358, N356, N8);
buf BUF1 (N359, N354);
xor XOR2 (N360, N317, N20);
not NOT1 (N361, N351);
or OR3 (N362, N361, N90, N106);
and AND4 (N363, N349, N76, N163, N110);
buf BUF1 (N364, N358);
nand NAND3 (N365, N357, N241, N302);
nand NAND2 (N366, N346, N304);
not NOT1 (N367, N359);
nand NAND2 (N368, N364, N216);
not NOT1 (N369, N363);
nor NOR2 (N370, N362, N196);
xor XOR2 (N371, N355, N104);
not NOT1 (N372, N368);
not NOT1 (N373, N365);
nand NAND2 (N374, N367, N325);
xor XOR2 (N375, N372, N166);
buf BUF1 (N376, N375);
xor XOR2 (N377, N360, N362);
not NOT1 (N378, N369);
buf BUF1 (N379, N377);
buf BUF1 (N380, N378);
xor XOR2 (N381, N376, N129);
nand NAND4 (N382, N352, N347, N205, N244);
and AND2 (N383, N379, N201);
buf BUF1 (N384, N383);
and AND2 (N385, N374, N324);
buf BUF1 (N386, N380);
xor XOR2 (N387, N373, N107);
and AND2 (N388, N366, N313);
and AND3 (N389, N382, N12, N2);
nor NOR3 (N390, N371, N2, N286);
nor NOR2 (N391, N384, N114);
or OR2 (N392, N391, N143);
buf BUF1 (N393, N353);
nand NAND4 (N394, N393, N352, N316, N2);
or OR3 (N395, N392, N49, N247);
nor NOR2 (N396, N389, N300);
nor NOR2 (N397, N388, N258);
nor NOR4 (N398, N397, N203, N315, N358);
xor XOR2 (N399, N396, N295);
xor XOR2 (N400, N385, N383);
buf BUF1 (N401, N399);
xor XOR2 (N402, N400, N109);
buf BUF1 (N403, N381);
and AND3 (N404, N390, N322, N38);
xor XOR2 (N405, N386, N144);
xor XOR2 (N406, N394, N29);
buf BUF1 (N407, N403);
and AND4 (N408, N401, N8, N270, N308);
or OR2 (N409, N406, N365);
buf BUF1 (N410, N402);
or OR2 (N411, N409, N384);
and AND2 (N412, N407, N263);
not NOT1 (N413, N405);
not NOT1 (N414, N404);
buf BUF1 (N415, N387);
or OR2 (N416, N413, N399);
or OR2 (N417, N398, N237);
xor XOR2 (N418, N370, N155);
buf BUF1 (N419, N410);
nor NOR2 (N420, N417, N14);
nor NOR2 (N421, N418, N257);
and AND3 (N422, N411, N297, N177);
xor XOR2 (N423, N420, N306);
and AND4 (N424, N419, N276, N76, N308);
not NOT1 (N425, N416);
not NOT1 (N426, N415);
or OR4 (N427, N425, N150, N68, N210);
not NOT1 (N428, N423);
xor XOR2 (N429, N412, N266);
not NOT1 (N430, N421);
or OR2 (N431, N395, N85);
nand NAND2 (N432, N431, N123);
nand NAND4 (N433, N430, N158, N39, N318);
not NOT1 (N434, N433);
xor XOR2 (N435, N434, N145);
not NOT1 (N436, N428);
and AND2 (N437, N427, N295);
nand NAND4 (N438, N424, N418, N324, N65);
or OR3 (N439, N435, N432, N436);
not NOT1 (N440, N123);
not NOT1 (N441, N324);
xor XOR2 (N442, N441, N344);
or OR2 (N443, N429, N7);
buf BUF1 (N444, N437);
xor XOR2 (N445, N440, N26);
xor XOR2 (N446, N442, N68);
not NOT1 (N447, N443);
not NOT1 (N448, N445);
nor NOR3 (N449, N439, N29, N170);
or OR3 (N450, N447, N239, N398);
or OR3 (N451, N446, N189, N37);
buf BUF1 (N452, N451);
xor XOR2 (N453, N448, N303);
or OR3 (N454, N453, N438, N203);
buf BUF1 (N455, N397);
nand NAND2 (N456, N454, N255);
and AND4 (N457, N444, N72, N404, N452);
or OR3 (N458, N393, N291, N382);
nand NAND3 (N459, N422, N411, N203);
or OR4 (N460, N459, N83, N319, N206);
and AND2 (N461, N460, N146);
not NOT1 (N462, N414);
or OR3 (N463, N461, N205, N248);
nand NAND3 (N464, N450, N243, N245);
and AND4 (N465, N457, N148, N348, N390);
xor XOR2 (N466, N458, N416);
buf BUF1 (N467, N465);
nor NOR2 (N468, N456, N298);
buf BUF1 (N469, N463);
or OR2 (N470, N408, N1);
not NOT1 (N471, N470);
not NOT1 (N472, N426);
or OR3 (N473, N466, N268, N407);
not NOT1 (N474, N449);
not NOT1 (N475, N467);
nand NAND2 (N476, N464, N271);
or OR4 (N477, N474, N146, N282, N281);
and AND2 (N478, N473, N455);
not NOT1 (N479, N44);
buf BUF1 (N480, N469);
xor XOR2 (N481, N478, N153);
or OR4 (N482, N479, N139, N388, N86);
xor XOR2 (N483, N482, N186);
nand NAND3 (N484, N477, N233, N235);
and AND2 (N485, N475, N455);
not NOT1 (N486, N476);
nand NAND4 (N487, N472, N405, N187, N1);
or OR4 (N488, N485, N406, N432, N244);
buf BUF1 (N489, N462);
xor XOR2 (N490, N486, N121);
xor XOR2 (N491, N484, N90);
nor NOR4 (N492, N488, N157, N450, N360);
nand NAND2 (N493, N487, N36);
nor NOR3 (N494, N493, N79, N129);
nand NAND3 (N495, N489, N427, N450);
or OR3 (N496, N483, N16, N332);
nor NOR2 (N497, N481, N158);
buf BUF1 (N498, N492);
nand NAND2 (N499, N471, N157);
buf BUF1 (N500, N497);
and AND2 (N501, N490, N177);
nor NOR2 (N502, N499, N34);
buf BUF1 (N503, N491);
or OR2 (N504, N501, N252);
nand NAND4 (N505, N502, N477, N145, N167);
nand NAND2 (N506, N496, N79);
or OR4 (N507, N503, N373, N185, N126);
and AND3 (N508, N505, N359, N367);
not NOT1 (N509, N468);
or OR4 (N510, N506, N199, N416, N51);
nor NOR2 (N511, N494, N363);
and AND3 (N512, N498, N366, N310);
xor XOR2 (N513, N495, N451);
xor XOR2 (N514, N480, N434);
nand NAND3 (N515, N509, N347, N447);
not NOT1 (N516, N515);
or OR4 (N517, N500, N401, N175, N145);
or OR3 (N518, N517, N94, N350);
buf BUF1 (N519, N513);
nand NAND3 (N520, N512, N156, N369);
nand NAND2 (N521, N520, N46);
not NOT1 (N522, N521);
xor XOR2 (N523, N504, N483);
xor XOR2 (N524, N508, N342);
buf BUF1 (N525, N511);
or OR4 (N526, N510, N402, N225, N417);
xor XOR2 (N527, N526, N464);
nand NAND4 (N528, N524, N401, N208, N3);
xor XOR2 (N529, N518, N124);
or OR4 (N530, N529, N368, N10, N134);
not NOT1 (N531, N528);
nor NOR2 (N532, N507, N97);
buf BUF1 (N533, N527);
xor XOR2 (N534, N519, N391);
nand NAND2 (N535, N531, N522);
and AND4 (N536, N522, N391, N392, N101);
nor NOR4 (N537, N532, N444, N348, N405);
xor XOR2 (N538, N534, N101);
nand NAND2 (N539, N536, N192);
nor NOR3 (N540, N538, N532, N27);
buf BUF1 (N541, N533);
nor NOR3 (N542, N514, N287, N96);
buf BUF1 (N543, N541);
and AND2 (N544, N523, N537);
and AND4 (N545, N234, N148, N224, N473);
not NOT1 (N546, N516);
xor XOR2 (N547, N540, N181);
and AND4 (N548, N539, N82, N434, N50);
and AND3 (N549, N548, N170, N404);
buf BUF1 (N550, N549);
nand NAND2 (N551, N545, N347);
nand NAND4 (N552, N530, N515, N131, N473);
xor XOR2 (N553, N547, N505);
xor XOR2 (N554, N542, N513);
buf BUF1 (N555, N546);
nor NOR4 (N556, N535, N544, N64, N378);
nand NAND2 (N557, N9, N398);
nand NAND2 (N558, N554, N199);
and AND2 (N559, N543, N554);
nor NOR3 (N560, N553, N80, N460);
and AND2 (N561, N556, N414);
not NOT1 (N562, N552);
not NOT1 (N563, N557);
nor NOR4 (N564, N555, N317, N296, N213);
xor XOR2 (N565, N562, N343);
nand NAND2 (N566, N565, N214);
xor XOR2 (N567, N564, N496);
and AND2 (N568, N550, N170);
buf BUF1 (N569, N563);
and AND2 (N570, N558, N505);
nor NOR4 (N571, N560, N447, N251, N516);
or OR3 (N572, N569, N404, N150);
or OR4 (N573, N561, N351, N436, N568);
or OR3 (N574, N24, N204, N555);
buf BUF1 (N575, N567);
or OR2 (N576, N572, N449);
xor XOR2 (N577, N559, N555);
xor XOR2 (N578, N551, N79);
nor NOR2 (N579, N577, N198);
not NOT1 (N580, N525);
buf BUF1 (N581, N573);
and AND4 (N582, N566, N491, N327, N200);
nand NAND4 (N583, N582, N493, N144, N258);
or OR3 (N584, N570, N221, N190);
xor XOR2 (N585, N578, N380);
not NOT1 (N586, N576);
or OR4 (N587, N571, N423, N487, N52);
nand NAND3 (N588, N587, N224, N357);
or OR2 (N589, N584, N406);
nor NOR4 (N590, N588, N155, N322, N396);
or OR2 (N591, N575, N547);
and AND2 (N592, N586, N248);
or OR4 (N593, N579, N103, N78, N159);
nor NOR2 (N594, N591, N421);
xor XOR2 (N595, N594, N95);
buf BUF1 (N596, N595);
and AND4 (N597, N593, N202, N266, N268);
nand NAND2 (N598, N597, N208);
xor XOR2 (N599, N574, N501);
or OR4 (N600, N583, N78, N478, N56);
and AND2 (N601, N599, N296);
nand NAND4 (N602, N589, N347, N158, N531);
nand NAND4 (N603, N590, N423, N78, N595);
nand NAND3 (N604, N580, N103, N595);
not NOT1 (N605, N592);
buf BUF1 (N606, N605);
xor XOR2 (N607, N600, N283);
xor XOR2 (N608, N602, N266);
buf BUF1 (N609, N606);
buf BUF1 (N610, N603);
nand NAND2 (N611, N585, N19);
and AND2 (N612, N608, N119);
and AND2 (N613, N609, N488);
nand NAND4 (N614, N598, N337, N585, N25);
buf BUF1 (N615, N607);
and AND2 (N616, N601, N190);
and AND2 (N617, N581, N451);
nand NAND2 (N618, N613, N7);
or OR4 (N619, N615, N471, N356, N228);
or OR3 (N620, N614, N228, N43);
and AND2 (N621, N604, N309);
and AND3 (N622, N621, N512, N482);
not NOT1 (N623, N619);
or OR4 (N624, N596, N453, N158, N107);
not NOT1 (N625, N616);
not NOT1 (N626, N622);
buf BUF1 (N627, N618);
buf BUF1 (N628, N611);
nor NOR3 (N629, N628, N609, N139);
nor NOR4 (N630, N620, N369, N248, N118);
and AND2 (N631, N612, N80);
buf BUF1 (N632, N610);
and AND2 (N633, N627, N573);
not NOT1 (N634, N629);
buf BUF1 (N635, N626);
buf BUF1 (N636, N633);
and AND4 (N637, N623, N28, N285, N584);
nor NOR3 (N638, N630, N254, N130);
not NOT1 (N639, N624);
nor NOR3 (N640, N631, N526, N441);
nor NOR4 (N641, N640, N148, N510, N17);
buf BUF1 (N642, N634);
buf BUF1 (N643, N637);
and AND2 (N644, N639, N611);
xor XOR2 (N645, N617, N502);
nand NAND4 (N646, N645, N386, N213, N134);
buf BUF1 (N647, N625);
xor XOR2 (N648, N647, N603);
nor NOR2 (N649, N646, N97);
or OR3 (N650, N636, N619, N370);
nor NOR3 (N651, N650, N560, N204);
or OR3 (N652, N643, N178, N126);
xor XOR2 (N653, N651, N401);
buf BUF1 (N654, N638);
nor NOR2 (N655, N635, N276);
nor NOR2 (N656, N642, N546);
or OR4 (N657, N648, N586, N239, N508);
buf BUF1 (N658, N655);
nand NAND2 (N659, N652, N574);
nor NOR4 (N660, N649, N353, N656, N41);
xor XOR2 (N661, N618, N355);
and AND3 (N662, N659, N175, N607);
not NOT1 (N663, N644);
not NOT1 (N664, N653);
not NOT1 (N665, N632);
not NOT1 (N666, N663);
xor XOR2 (N667, N666, N608);
buf BUF1 (N668, N661);
nor NOR4 (N669, N657, N393, N552, N15);
nor NOR4 (N670, N667, N37, N299, N194);
buf BUF1 (N671, N662);
xor XOR2 (N672, N671, N246);
xor XOR2 (N673, N654, N297);
or OR3 (N674, N658, N430, N543);
or OR4 (N675, N673, N101, N397, N5);
xor XOR2 (N676, N664, N298);
buf BUF1 (N677, N675);
and AND2 (N678, N669, N90);
and AND3 (N679, N676, N397, N459);
or OR3 (N680, N641, N427, N291);
or OR2 (N681, N674, N57);
nand NAND3 (N682, N679, N111, N485);
nand NAND2 (N683, N672, N32);
buf BUF1 (N684, N681);
and AND4 (N685, N678, N652, N131, N174);
nor NOR2 (N686, N683, N440);
xor XOR2 (N687, N677, N487);
or OR2 (N688, N668, N208);
or OR2 (N689, N687, N431);
xor XOR2 (N690, N686, N87);
and AND4 (N691, N688, N437, N216, N329);
buf BUF1 (N692, N670);
buf BUF1 (N693, N682);
xor XOR2 (N694, N693, N107);
not NOT1 (N695, N684);
not NOT1 (N696, N690);
and AND2 (N697, N680, N123);
nand NAND2 (N698, N695, N399);
buf BUF1 (N699, N691);
buf BUF1 (N700, N665);
not NOT1 (N701, N698);
nor NOR2 (N702, N685, N66);
nand NAND2 (N703, N701, N405);
or OR2 (N704, N700, N408);
nor NOR4 (N705, N696, N325, N44, N350);
nor NOR4 (N706, N702, N698, N218, N16);
nand NAND3 (N707, N704, N437, N166);
buf BUF1 (N708, N703);
not NOT1 (N709, N707);
nand NAND4 (N710, N660, N636, N281, N664);
xor XOR2 (N711, N709, N701);
buf BUF1 (N712, N706);
or OR2 (N713, N689, N155);
buf BUF1 (N714, N713);
nand NAND2 (N715, N710, N111);
not NOT1 (N716, N711);
nand NAND4 (N717, N699, N151, N659, N578);
not NOT1 (N718, N697);
or OR2 (N719, N717, N128);
or OR4 (N720, N716, N561, N520, N615);
and AND2 (N721, N715, N28);
nor NOR3 (N722, N721, N332, N335);
nand NAND3 (N723, N718, N696, N158);
or OR2 (N724, N720, N615);
buf BUF1 (N725, N714);
nand NAND3 (N726, N723, N277, N314);
and AND4 (N727, N694, N421, N294, N571);
buf BUF1 (N728, N705);
buf BUF1 (N729, N724);
xor XOR2 (N730, N712, N658);
xor XOR2 (N731, N722, N687);
not NOT1 (N732, N727);
and AND3 (N733, N708, N252, N503);
and AND2 (N734, N726, N467);
or OR4 (N735, N732, N130, N434, N163);
or OR3 (N736, N728, N415, N205);
nor NOR2 (N737, N736, N686);
nand NAND4 (N738, N730, N589, N517, N148);
buf BUF1 (N739, N734);
not NOT1 (N740, N729);
xor XOR2 (N741, N740, N255);
nand NAND4 (N742, N739, N99, N327, N223);
xor XOR2 (N743, N742, N344);
or OR2 (N744, N733, N460);
or OR2 (N745, N741, N148);
nand NAND3 (N746, N744, N443, N146);
buf BUF1 (N747, N731);
and AND2 (N748, N737, N362);
buf BUF1 (N749, N725);
buf BUF1 (N750, N748);
or OR4 (N751, N749, N2, N387, N390);
and AND2 (N752, N746, N56);
buf BUF1 (N753, N692);
nor NOR4 (N754, N750, N174, N149, N458);
xor XOR2 (N755, N738, N424);
not NOT1 (N756, N754);
buf BUF1 (N757, N755);
xor XOR2 (N758, N747, N658);
not NOT1 (N759, N719);
and AND3 (N760, N758, N470, N521);
not NOT1 (N761, N759);
or OR2 (N762, N745, N246);
xor XOR2 (N763, N743, N582);
nand NAND2 (N764, N751, N581);
nand NAND3 (N765, N763, N251, N236);
xor XOR2 (N766, N753, N603);
xor XOR2 (N767, N761, N270);
not NOT1 (N768, N764);
buf BUF1 (N769, N756);
nor NOR3 (N770, N760, N650, N728);
nand NAND2 (N771, N735, N569);
buf BUF1 (N772, N767);
not NOT1 (N773, N752);
or OR3 (N774, N770, N493, N54);
not NOT1 (N775, N765);
nor NOR4 (N776, N773, N738, N484, N696);
nor NOR2 (N777, N774, N138);
and AND3 (N778, N776, N304, N496);
and AND2 (N779, N772, N143);
xor XOR2 (N780, N766, N735);
xor XOR2 (N781, N777, N638);
nor NOR4 (N782, N771, N468, N124, N488);
and AND2 (N783, N775, N401);
buf BUF1 (N784, N778);
buf BUF1 (N785, N784);
and AND3 (N786, N780, N586, N618);
and AND2 (N787, N757, N568);
nand NAND3 (N788, N769, N428, N700);
xor XOR2 (N789, N762, N54);
buf BUF1 (N790, N785);
xor XOR2 (N791, N782, N192);
buf BUF1 (N792, N790);
or OR2 (N793, N791, N694);
and AND4 (N794, N768, N10, N95, N431);
buf BUF1 (N795, N787);
not NOT1 (N796, N792);
or OR3 (N797, N789, N470, N516);
or OR2 (N798, N786, N377);
not NOT1 (N799, N779);
or OR2 (N800, N799, N315);
nand NAND3 (N801, N793, N622, N191);
or OR3 (N802, N794, N551, N153);
xor XOR2 (N803, N801, N284);
and AND2 (N804, N802, N465);
or OR2 (N805, N804, N533);
xor XOR2 (N806, N781, N246);
buf BUF1 (N807, N800);
or OR3 (N808, N805, N336, N437);
nor NOR3 (N809, N808, N622, N205);
buf BUF1 (N810, N798);
not NOT1 (N811, N783);
and AND4 (N812, N806, N233, N709, N458);
buf BUF1 (N813, N797);
xor XOR2 (N814, N807, N114);
not NOT1 (N815, N812);
nand NAND3 (N816, N810, N182, N195);
xor XOR2 (N817, N813, N492);
buf BUF1 (N818, N811);
buf BUF1 (N819, N818);
buf BUF1 (N820, N819);
or OR3 (N821, N815, N37, N388);
nand NAND2 (N822, N809, N680);
nand NAND2 (N823, N795, N563);
xor XOR2 (N824, N788, N304);
xor XOR2 (N825, N822, N262);
nand NAND4 (N826, N823, N347, N89, N793);
buf BUF1 (N827, N824);
xor XOR2 (N828, N796, N600);
nand NAND2 (N829, N803, N430);
not NOT1 (N830, N825);
or OR3 (N831, N814, N145, N700);
xor XOR2 (N832, N826, N230);
xor XOR2 (N833, N817, N57);
xor XOR2 (N834, N827, N189);
nor NOR4 (N835, N833, N379, N635, N714);
or OR4 (N836, N816, N78, N64, N416);
and AND3 (N837, N834, N186, N778);
xor XOR2 (N838, N832, N671);
nor NOR4 (N839, N829, N670, N658, N423);
or OR3 (N840, N839, N59, N692);
nor NOR4 (N841, N837, N647, N467, N711);
xor XOR2 (N842, N836, N456);
nand NAND4 (N843, N828, N50, N175, N592);
and AND3 (N844, N835, N726, N843);
and AND4 (N845, N604, N286, N241, N169);
or OR4 (N846, N820, N598, N179, N193);
xor XOR2 (N847, N821, N649);
xor XOR2 (N848, N831, N357);
nor NOR2 (N849, N840, N841);
xor XOR2 (N850, N314, N163);
buf BUF1 (N851, N830);
and AND4 (N852, N850, N137, N192, N255);
buf BUF1 (N853, N848);
nor NOR2 (N854, N845, N172);
nor NOR4 (N855, N851, N410, N559, N247);
and AND2 (N856, N854, N209);
xor XOR2 (N857, N849, N148);
nand NAND2 (N858, N842, N115);
buf BUF1 (N859, N856);
and AND2 (N860, N859, N482);
or OR3 (N861, N855, N633, N648);
nand NAND3 (N862, N838, N580, N735);
buf BUF1 (N863, N846);
or OR2 (N864, N863, N150);
nand NAND2 (N865, N864, N695);
nand NAND2 (N866, N844, N736);
buf BUF1 (N867, N847);
not NOT1 (N868, N867);
not NOT1 (N869, N861);
nand NAND4 (N870, N852, N331, N862, N564);
buf BUF1 (N871, N125);
and AND4 (N872, N870, N496, N320, N401);
or OR3 (N873, N860, N736, N165);
nor NOR3 (N874, N873, N752, N721);
nor NOR2 (N875, N872, N319);
xor XOR2 (N876, N875, N256);
xor XOR2 (N877, N857, N383);
nand NAND3 (N878, N858, N420, N345);
and AND3 (N879, N878, N175, N629);
nor NOR3 (N880, N869, N183, N800);
and AND2 (N881, N865, N206);
nor NOR3 (N882, N853, N224, N455);
nor NOR2 (N883, N874, N110);
nor NOR3 (N884, N883, N328, N510);
buf BUF1 (N885, N876);
nand NAND4 (N886, N879, N231, N258, N775);
buf BUF1 (N887, N884);
xor XOR2 (N888, N880, N111);
xor XOR2 (N889, N871, N292);
buf BUF1 (N890, N886);
xor XOR2 (N891, N890, N167);
not NOT1 (N892, N882);
buf BUF1 (N893, N892);
xor XOR2 (N894, N877, N494);
nor NOR4 (N895, N893, N268, N429, N833);
xor XOR2 (N896, N866, N18);
or OR2 (N897, N894, N535);
and AND2 (N898, N888, N553);
nand NAND2 (N899, N887, N355);
or OR2 (N900, N898, N727);
nand NAND2 (N901, N897, N827);
nand NAND2 (N902, N900, N572);
nand NAND3 (N903, N881, N532, N141);
not NOT1 (N904, N889);
not NOT1 (N905, N904);
nor NOR4 (N906, N902, N415, N673, N115);
or OR2 (N907, N895, N59);
not NOT1 (N908, N907);
xor XOR2 (N909, N896, N264);
not NOT1 (N910, N899);
nor NOR4 (N911, N910, N162, N623, N839);
buf BUF1 (N912, N911);
and AND4 (N913, N905, N108, N284, N722);
nand NAND3 (N914, N913, N835, N158);
xor XOR2 (N915, N909, N164);
buf BUF1 (N916, N868);
xor XOR2 (N917, N916, N530);
and AND4 (N918, N908, N66, N909, N515);
or OR4 (N919, N903, N823, N291, N314);
xor XOR2 (N920, N912, N700);
nor NOR4 (N921, N885, N395, N156, N258);
buf BUF1 (N922, N891);
xor XOR2 (N923, N919, N394);
xor XOR2 (N924, N918, N560);
not NOT1 (N925, N920);
buf BUF1 (N926, N921);
and AND3 (N927, N922, N112, N478);
nand NAND2 (N928, N917, N349);
nor NOR2 (N929, N914, N680);
nand NAND4 (N930, N924, N404, N585, N244);
not NOT1 (N931, N929);
and AND3 (N932, N930, N646, N163);
or OR2 (N933, N931, N719);
nor NOR3 (N934, N928, N171, N106);
and AND4 (N935, N925, N250, N592, N541);
not NOT1 (N936, N906);
nand NAND3 (N937, N932, N796, N29);
or OR2 (N938, N901, N517);
xor XOR2 (N939, N933, N656);
xor XOR2 (N940, N939, N739);
not NOT1 (N941, N926);
or OR4 (N942, N927, N32, N170, N511);
xor XOR2 (N943, N923, N936);
nor NOR2 (N944, N830, N423);
or OR2 (N945, N915, N521);
and AND3 (N946, N938, N523, N135);
and AND2 (N947, N943, N16);
buf BUF1 (N948, N940);
not NOT1 (N949, N947);
not NOT1 (N950, N934);
nor NOR4 (N951, N944, N712, N380, N411);
nor NOR4 (N952, N946, N464, N833, N932);
not NOT1 (N953, N950);
buf BUF1 (N954, N937);
buf BUF1 (N955, N935);
nand NAND3 (N956, N954, N427, N518);
and AND3 (N957, N941, N363, N678);
xor XOR2 (N958, N953, N350);
nor NOR3 (N959, N958, N412, N847);
and AND4 (N960, N942, N84, N650, N946);
or OR4 (N961, N957, N387, N161, N68);
and AND4 (N962, N959, N347, N799, N32);
buf BUF1 (N963, N952);
nor NOR3 (N964, N963, N553, N823);
nand NAND2 (N965, N955, N84);
not NOT1 (N966, N964);
buf BUF1 (N967, N951);
or OR3 (N968, N956, N281, N532);
nand NAND4 (N969, N948, N932, N4, N12);
or OR3 (N970, N962, N885, N777);
not NOT1 (N971, N945);
nor NOR3 (N972, N965, N235, N853);
or OR4 (N973, N969, N101, N668, N325);
xor XOR2 (N974, N967, N303);
nand NAND3 (N975, N949, N699, N834);
buf BUF1 (N976, N971);
or OR4 (N977, N974, N311, N67, N968);
nand NAND4 (N978, N301, N677, N524, N589);
nor NOR4 (N979, N977, N321, N644, N676);
nand NAND3 (N980, N961, N368, N902);
buf BUF1 (N981, N975);
or OR4 (N982, N973, N560, N654, N800);
not NOT1 (N983, N976);
nor NOR4 (N984, N970, N794, N392, N745);
or OR2 (N985, N983, N103);
nor NOR2 (N986, N966, N466);
nand NAND2 (N987, N984, N200);
nor NOR4 (N988, N982, N648, N515, N418);
not NOT1 (N989, N979);
nor NOR2 (N990, N987, N121);
xor XOR2 (N991, N972, N423);
nor NOR4 (N992, N988, N104, N750, N447);
not NOT1 (N993, N960);
nand NAND2 (N994, N993, N881);
buf BUF1 (N995, N991);
and AND3 (N996, N980, N29, N238);
nand NAND4 (N997, N981, N199, N287, N150);
nand NAND4 (N998, N995, N186, N483, N179);
or OR3 (N999, N986, N91, N549);
nand NAND4 (N1000, N978, N398, N63, N753);
or OR3 (N1001, N994, N371, N527);
or OR4 (N1002, N1001, N403, N143, N240);
nand NAND3 (N1003, N1000, N101, N968);
nor NOR4 (N1004, N997, N927, N984, N21);
nor NOR2 (N1005, N999, N724);
xor XOR2 (N1006, N1003, N161);
buf BUF1 (N1007, N1006);
xor XOR2 (N1008, N989, N836);
nand NAND4 (N1009, N1004, N375, N973, N271);
nor NOR2 (N1010, N992, N670);
xor XOR2 (N1011, N996, N391);
nand NAND2 (N1012, N1002, N991);
nand NAND4 (N1013, N990, N77, N730, N501);
or OR3 (N1014, N1012, N710, N284);
nor NOR4 (N1015, N1010, N307, N562, N926);
nor NOR2 (N1016, N1013, N919);
xor XOR2 (N1017, N998, N344);
nand NAND2 (N1018, N1014, N841);
buf BUF1 (N1019, N1018);
buf BUF1 (N1020, N1019);
and AND4 (N1021, N1020, N353, N783, N501);
or OR3 (N1022, N1011, N724, N13);
or OR4 (N1023, N1008, N368, N489, N985);
xor XOR2 (N1024, N240, N943);
or OR3 (N1025, N1024, N766, N1016);
not NOT1 (N1026, N427);
nor NOR3 (N1027, N1023, N167, N680);
xor XOR2 (N1028, N1015, N998);
xor XOR2 (N1029, N1021, N33);
xor XOR2 (N1030, N1025, N224);
xor XOR2 (N1031, N1030, N784);
nor NOR3 (N1032, N1017, N854, N510);
buf BUF1 (N1033, N1009);
and AND4 (N1034, N1033, N442, N586, N318);
not NOT1 (N1035, N1005);
or OR3 (N1036, N1027, N335, N762);
nor NOR4 (N1037, N1029, N682, N92, N271);
buf BUF1 (N1038, N1035);
nor NOR2 (N1039, N1034, N811);
and AND3 (N1040, N1039, N599, N722);
and AND4 (N1041, N1007, N748, N202, N275);
buf BUF1 (N1042, N1037);
xor XOR2 (N1043, N1032, N578);
xor XOR2 (N1044, N1043, N730);
not NOT1 (N1045, N1040);
nand NAND3 (N1046, N1031, N888, N823);
buf BUF1 (N1047, N1022);
nor NOR2 (N1048, N1041, N344);
xor XOR2 (N1049, N1028, N93);
not NOT1 (N1050, N1026);
or OR3 (N1051, N1049, N87, N52);
xor XOR2 (N1052, N1047, N862);
xor XOR2 (N1053, N1048, N654);
not NOT1 (N1054, N1046);
nor NOR3 (N1055, N1054, N511, N894);
buf BUF1 (N1056, N1055);
nand NAND4 (N1057, N1056, N3, N492, N113);
nor NOR2 (N1058, N1051, N838);
not NOT1 (N1059, N1045);
not NOT1 (N1060, N1052);
and AND4 (N1061, N1050, N105, N959, N881);
nand NAND2 (N1062, N1057, N566);
xor XOR2 (N1063, N1042, N114);
xor XOR2 (N1064, N1044, N534);
nor NOR4 (N1065, N1059, N890, N110, N295);
nand NAND3 (N1066, N1063, N223, N652);
nand NAND4 (N1067, N1062, N241, N558, N433);
nor NOR4 (N1068, N1060, N1031, N254, N139);
buf BUF1 (N1069, N1053);
not NOT1 (N1070, N1068);
not NOT1 (N1071, N1066);
nor NOR3 (N1072, N1065, N900, N29);
and AND2 (N1073, N1061, N902);
buf BUF1 (N1074, N1064);
xor XOR2 (N1075, N1036, N451);
nand NAND2 (N1076, N1075, N338);
nand NAND4 (N1077, N1071, N186, N488, N181);
or OR3 (N1078, N1067, N552, N719);
nor NOR3 (N1079, N1038, N674, N480);
nand NAND3 (N1080, N1078, N501, N82);
buf BUF1 (N1081, N1070);
nor NOR2 (N1082, N1072, N1063);
xor XOR2 (N1083, N1069, N203);
nand NAND2 (N1084, N1076, N1014);
or OR3 (N1085, N1081, N457, N111);
buf BUF1 (N1086, N1083);
and AND2 (N1087, N1085, N649);
nand NAND4 (N1088, N1079, N202, N525, N455);
nor NOR4 (N1089, N1082, N189, N1052, N727);
or OR4 (N1090, N1088, N225, N560, N646);
and AND3 (N1091, N1058, N566, N496);
xor XOR2 (N1092, N1087, N1085);
and AND4 (N1093, N1077, N563, N964, N271);
and AND4 (N1094, N1092, N964, N1062, N774);
not NOT1 (N1095, N1090);
nor NOR2 (N1096, N1089, N654);
or OR2 (N1097, N1093, N587);
or OR2 (N1098, N1095, N797);
not NOT1 (N1099, N1084);
nor NOR4 (N1100, N1074, N188, N392, N582);
or OR2 (N1101, N1094, N339);
not NOT1 (N1102, N1098);
xor XOR2 (N1103, N1097, N698);
xor XOR2 (N1104, N1091, N365);
nand NAND4 (N1105, N1103, N951, N1044, N918);
nand NAND3 (N1106, N1102, N131, N729);
nand NAND4 (N1107, N1099, N780, N231, N811);
nor NOR3 (N1108, N1073, N275, N673);
not NOT1 (N1109, N1107);
not NOT1 (N1110, N1104);
buf BUF1 (N1111, N1105);
buf BUF1 (N1112, N1111);
not NOT1 (N1113, N1106);
not NOT1 (N1114, N1109);
not NOT1 (N1115, N1113);
nand NAND2 (N1116, N1096, N1022);
nand NAND2 (N1117, N1114, N214);
or OR3 (N1118, N1086, N864, N984);
or OR4 (N1119, N1110, N876, N745, N33);
buf BUF1 (N1120, N1112);
xor XOR2 (N1121, N1116, N146);
nor NOR2 (N1122, N1100, N1121);
and AND3 (N1123, N338, N979, N983);
nand NAND3 (N1124, N1080, N1022, N399);
and AND3 (N1125, N1122, N136, N123);
buf BUF1 (N1126, N1123);
or OR4 (N1127, N1124, N1003, N338, N1057);
and AND3 (N1128, N1120, N446, N193);
or OR2 (N1129, N1101, N155);
buf BUF1 (N1130, N1119);
or OR4 (N1131, N1127, N121, N960, N86);
and AND3 (N1132, N1131, N201, N577);
or OR4 (N1133, N1125, N802, N21, N817);
or OR2 (N1134, N1118, N631);
buf BUF1 (N1135, N1134);
and AND3 (N1136, N1115, N913, N986);
xor XOR2 (N1137, N1135, N797);
not NOT1 (N1138, N1128);
not NOT1 (N1139, N1137);
buf BUF1 (N1140, N1130);
and AND4 (N1141, N1108, N713, N429, N802);
or OR3 (N1142, N1132, N896, N528);
buf BUF1 (N1143, N1129);
buf BUF1 (N1144, N1117);
buf BUF1 (N1145, N1133);
and AND4 (N1146, N1126, N485, N339, N391);
or OR4 (N1147, N1139, N1089, N913, N185);
nor NOR3 (N1148, N1143, N132, N275);
nand NAND2 (N1149, N1140, N1119);
buf BUF1 (N1150, N1145);
nand NAND2 (N1151, N1149, N1086);
or OR2 (N1152, N1150, N106);
and AND4 (N1153, N1146, N704, N324, N102);
nand NAND3 (N1154, N1138, N1059, N1128);
nand NAND2 (N1155, N1152, N486);
not NOT1 (N1156, N1147);
buf BUF1 (N1157, N1156);
buf BUF1 (N1158, N1144);
xor XOR2 (N1159, N1157, N600);
xor XOR2 (N1160, N1159, N765);
nand NAND2 (N1161, N1141, N482);
nand NAND4 (N1162, N1153, N728, N763, N354);
buf BUF1 (N1163, N1142);
nand NAND2 (N1164, N1161, N1151);
xor XOR2 (N1165, N910, N928);
nand NAND4 (N1166, N1163, N537, N770, N1042);
and AND3 (N1167, N1165, N824, N372);
and AND4 (N1168, N1136, N243, N323, N1043);
or OR3 (N1169, N1154, N720, N262);
or OR3 (N1170, N1155, N83, N1017);
nand NAND3 (N1171, N1162, N1127, N539);
not NOT1 (N1172, N1167);
xor XOR2 (N1173, N1148, N451);
nand NAND3 (N1174, N1172, N692, N659);
nand NAND4 (N1175, N1160, N585, N624, N1158);
nor NOR2 (N1176, N919, N610);
buf BUF1 (N1177, N1168);
nor NOR3 (N1178, N1169, N163, N196);
nand NAND4 (N1179, N1174, N517, N337, N414);
nor NOR2 (N1180, N1170, N445);
or OR4 (N1181, N1180, N341, N1161, N330);
not NOT1 (N1182, N1176);
nand NAND3 (N1183, N1178, N846, N190);
nor NOR3 (N1184, N1182, N775, N153);
nor NOR3 (N1185, N1183, N826, N828);
not NOT1 (N1186, N1175);
buf BUF1 (N1187, N1166);
and AND4 (N1188, N1187, N798, N101, N922);
buf BUF1 (N1189, N1179);
or OR3 (N1190, N1177, N938, N161);
buf BUF1 (N1191, N1184);
xor XOR2 (N1192, N1171, N786);
and AND3 (N1193, N1181, N529, N831);
nand NAND2 (N1194, N1189, N203);
buf BUF1 (N1195, N1188);
buf BUF1 (N1196, N1194);
and AND4 (N1197, N1190, N638, N1085, N1011);
xor XOR2 (N1198, N1196, N926);
not NOT1 (N1199, N1191);
buf BUF1 (N1200, N1197);
not NOT1 (N1201, N1198);
xor XOR2 (N1202, N1185, N1040);
nor NOR2 (N1203, N1201, N959);
xor XOR2 (N1204, N1193, N1124);
not NOT1 (N1205, N1164);
xor XOR2 (N1206, N1202, N542);
nand NAND4 (N1207, N1173, N1107, N718, N45);
xor XOR2 (N1208, N1192, N86);
nor NOR3 (N1209, N1186, N567, N695);
nand NAND2 (N1210, N1200, N79);
and AND4 (N1211, N1207, N44, N675, N964);
buf BUF1 (N1212, N1204);
nor NOR3 (N1213, N1209, N1030, N1074);
xor XOR2 (N1214, N1213, N343);
xor XOR2 (N1215, N1203, N118);
or OR4 (N1216, N1215, N1161, N913, N1162);
nand NAND2 (N1217, N1214, N238);
and AND4 (N1218, N1206, N889, N191, N1018);
not NOT1 (N1219, N1212);
nand NAND4 (N1220, N1210, N51, N80, N794);
and AND3 (N1221, N1205, N1062, N720);
nor NOR4 (N1222, N1216, N993, N94, N515);
nor NOR2 (N1223, N1222, N459);
nand NAND3 (N1224, N1221, N256, N144);
and AND2 (N1225, N1211, N44);
or OR4 (N1226, N1208, N621, N164, N561);
nor NOR3 (N1227, N1217, N571, N962);
and AND4 (N1228, N1195, N1064, N693, N961);
xor XOR2 (N1229, N1223, N831);
buf BUF1 (N1230, N1199);
buf BUF1 (N1231, N1227);
nor NOR2 (N1232, N1229, N656);
or OR2 (N1233, N1230, N964);
nor NOR2 (N1234, N1233, N416);
or OR4 (N1235, N1218, N242, N995, N1010);
or OR2 (N1236, N1235, N255);
and AND4 (N1237, N1226, N305, N319, N20);
xor XOR2 (N1238, N1224, N1136);
or OR4 (N1239, N1219, N251, N1087, N704);
or OR4 (N1240, N1231, N117, N159, N953);
nand NAND4 (N1241, N1232, N73, N323, N441);
buf BUF1 (N1242, N1228);
or OR3 (N1243, N1220, N872, N273);
xor XOR2 (N1244, N1236, N748);
buf BUF1 (N1245, N1244);
and AND4 (N1246, N1238, N572, N410, N1236);
xor XOR2 (N1247, N1245, N336);
and AND3 (N1248, N1225, N1135, N359);
nand NAND4 (N1249, N1248, N1158, N991, N613);
xor XOR2 (N1250, N1247, N1073);
nand NAND3 (N1251, N1246, N1174, N224);
xor XOR2 (N1252, N1239, N721);
nor NOR4 (N1253, N1241, N896, N660, N668);
nor NOR2 (N1254, N1253, N514);
xor XOR2 (N1255, N1252, N1201);
or OR4 (N1256, N1243, N500, N934, N619);
and AND4 (N1257, N1251, N204, N744, N129);
nor NOR3 (N1258, N1256, N666, N577);
nand NAND2 (N1259, N1257, N1163);
nand NAND2 (N1260, N1258, N972);
and AND3 (N1261, N1259, N456, N165);
xor XOR2 (N1262, N1260, N39);
and AND2 (N1263, N1249, N263);
nor NOR4 (N1264, N1234, N352, N930, N140);
and AND2 (N1265, N1237, N808);
buf BUF1 (N1266, N1255);
nand NAND4 (N1267, N1240, N122, N727, N693);
not NOT1 (N1268, N1242);
not NOT1 (N1269, N1266);
buf BUF1 (N1270, N1254);
buf BUF1 (N1271, N1270);
and AND4 (N1272, N1264, N1220, N1008, N563);
and AND2 (N1273, N1263, N1245);
nand NAND4 (N1274, N1267, N99, N72, N414);
xor XOR2 (N1275, N1269, N317);
xor XOR2 (N1276, N1250, N459);
nor NOR3 (N1277, N1272, N1071, N1022);
nor NOR2 (N1278, N1262, N1200);
not NOT1 (N1279, N1273);
or OR2 (N1280, N1265, N302);
nor NOR2 (N1281, N1274, N786);
and AND3 (N1282, N1275, N748, N498);
nor NOR2 (N1283, N1271, N712);
nor NOR2 (N1284, N1280, N226);
and AND2 (N1285, N1261, N833);
xor XOR2 (N1286, N1281, N1067);
nand NAND3 (N1287, N1276, N1147, N734);
or OR2 (N1288, N1277, N622);
or OR4 (N1289, N1268, N810, N319, N697);
xor XOR2 (N1290, N1285, N44);
nand NAND4 (N1291, N1283, N1143, N240, N570);
not NOT1 (N1292, N1288);
buf BUF1 (N1293, N1279);
not NOT1 (N1294, N1287);
and AND3 (N1295, N1292, N552, N325);
xor XOR2 (N1296, N1291, N259);
nor NOR3 (N1297, N1282, N720, N1079);
nor NOR3 (N1298, N1278, N895, N596);
not NOT1 (N1299, N1297);
buf BUF1 (N1300, N1299);
nor NOR3 (N1301, N1289, N277, N1095);
or OR4 (N1302, N1298, N952, N933, N885);
nand NAND4 (N1303, N1296, N1196, N928, N445);
xor XOR2 (N1304, N1303, N1072);
and AND2 (N1305, N1286, N456);
or OR2 (N1306, N1305, N1179);
not NOT1 (N1307, N1294);
nor NOR3 (N1308, N1306, N650, N823);
nand NAND3 (N1309, N1304, N731, N202);
nand NAND3 (N1310, N1301, N737, N1);
buf BUF1 (N1311, N1300);
buf BUF1 (N1312, N1311);
and AND3 (N1313, N1307, N754, N260);
xor XOR2 (N1314, N1309, N64);
xor XOR2 (N1315, N1312, N1102);
buf BUF1 (N1316, N1313);
or OR4 (N1317, N1310, N877, N1251, N24);
nand NAND3 (N1318, N1314, N93, N164);
nand NAND4 (N1319, N1316, N1026, N912, N660);
not NOT1 (N1320, N1284);
buf BUF1 (N1321, N1295);
or OR2 (N1322, N1319, N472);
nor NOR3 (N1323, N1320, N207, N195);
and AND2 (N1324, N1321, N261);
xor XOR2 (N1325, N1302, N1290);
and AND4 (N1326, N428, N1022, N261, N926);
nor NOR4 (N1327, N1293, N588, N1259, N814);
xor XOR2 (N1328, N1327, N636);
buf BUF1 (N1329, N1325);
nand NAND2 (N1330, N1323, N807);
not NOT1 (N1331, N1315);
and AND3 (N1332, N1318, N238, N789);
buf BUF1 (N1333, N1331);
nand NAND4 (N1334, N1328, N1051, N48, N450);
not NOT1 (N1335, N1333);
or OR2 (N1336, N1308, N101);
nand NAND4 (N1337, N1334, N680, N958, N444);
xor XOR2 (N1338, N1332, N1230);
or OR4 (N1339, N1329, N255, N829, N107);
and AND2 (N1340, N1336, N734);
buf BUF1 (N1341, N1317);
xor XOR2 (N1342, N1326, N906);
not NOT1 (N1343, N1342);
buf BUF1 (N1344, N1335);
buf BUF1 (N1345, N1339);
xor XOR2 (N1346, N1341, N117);
and AND2 (N1347, N1324, N1212);
nand NAND2 (N1348, N1322, N1229);
not NOT1 (N1349, N1348);
nand NAND3 (N1350, N1337, N997, N277);
xor XOR2 (N1351, N1340, N705);
and AND3 (N1352, N1330, N1150, N1146);
and AND2 (N1353, N1343, N458);
buf BUF1 (N1354, N1351);
xor XOR2 (N1355, N1349, N860);
and AND2 (N1356, N1354, N636);
nand NAND4 (N1357, N1356, N387, N831, N770);
or OR4 (N1358, N1350, N251, N235, N949);
or OR3 (N1359, N1353, N1270, N492);
or OR2 (N1360, N1352, N225);
nor NOR4 (N1361, N1360, N1214, N1129, N127);
xor XOR2 (N1362, N1361, N1151);
nand NAND3 (N1363, N1345, N1327, N894);
and AND2 (N1364, N1355, N1178);
not NOT1 (N1365, N1362);
xor XOR2 (N1366, N1338, N1223);
not NOT1 (N1367, N1357);
xor XOR2 (N1368, N1363, N267);
not NOT1 (N1369, N1368);
buf BUF1 (N1370, N1347);
not NOT1 (N1371, N1370);
xor XOR2 (N1372, N1367, N44);
and AND3 (N1373, N1359, N238, N665);
not NOT1 (N1374, N1344);
or OR3 (N1375, N1364, N260, N711);
buf BUF1 (N1376, N1358);
or OR3 (N1377, N1375, N1051, N1265);
xor XOR2 (N1378, N1366, N565);
and AND3 (N1379, N1376, N565, N1209);
xor XOR2 (N1380, N1346, N547);
nand NAND4 (N1381, N1365, N1330, N1010, N674);
buf BUF1 (N1382, N1369);
buf BUF1 (N1383, N1371);
xor XOR2 (N1384, N1382, N343);
not NOT1 (N1385, N1372);
or OR2 (N1386, N1381, N441);
nor NOR2 (N1387, N1377, N12);
and AND4 (N1388, N1386, N1037, N1253, N20);
not NOT1 (N1389, N1380);
not NOT1 (N1390, N1387);
and AND2 (N1391, N1374, N70);
nand NAND4 (N1392, N1385, N1114, N1163, N420);
buf BUF1 (N1393, N1384);
or OR3 (N1394, N1373, N102, N1170);
or OR3 (N1395, N1393, N631, N999);
nand NAND2 (N1396, N1390, N260);
xor XOR2 (N1397, N1379, N365);
nor NOR3 (N1398, N1394, N1181, N878);
buf BUF1 (N1399, N1392);
xor XOR2 (N1400, N1378, N978);
nand NAND3 (N1401, N1397, N1145, N131);
nor NOR3 (N1402, N1400, N1098, N745);
or OR3 (N1403, N1398, N701, N1396);
buf BUF1 (N1404, N1296);
nand NAND4 (N1405, N1391, N968, N44, N1357);
xor XOR2 (N1406, N1403, N690);
nand NAND2 (N1407, N1388, N919);
buf BUF1 (N1408, N1402);
xor XOR2 (N1409, N1401, N1047);
or OR2 (N1410, N1409, N1367);
xor XOR2 (N1411, N1404, N43);
nand NAND2 (N1412, N1406, N1092);
or OR3 (N1413, N1408, N504, N680);
nor NOR2 (N1414, N1399, N979);
and AND2 (N1415, N1407, N1068);
nor NOR3 (N1416, N1383, N650, N178);
and AND4 (N1417, N1414, N517, N102, N708);
or OR4 (N1418, N1415, N641, N526, N168);
nor NOR4 (N1419, N1417, N683, N1146, N302);
not NOT1 (N1420, N1418);
not NOT1 (N1421, N1405);
buf BUF1 (N1422, N1410);
nand NAND2 (N1423, N1419, N216);
not NOT1 (N1424, N1420);
nand NAND2 (N1425, N1423, N1005);
not NOT1 (N1426, N1421);
or OR2 (N1427, N1416, N401);
buf BUF1 (N1428, N1395);
or OR2 (N1429, N1389, N945);
not NOT1 (N1430, N1429);
nand NAND3 (N1431, N1430, N18, N221);
and AND3 (N1432, N1412, N229, N1035);
nand NAND2 (N1433, N1422, N1366);
nor NOR2 (N1434, N1426, N1224);
not NOT1 (N1435, N1428);
nand NAND3 (N1436, N1427, N939, N1288);
nand NAND2 (N1437, N1434, N1436);
or OR4 (N1438, N1258, N719, N1010, N1242);
and AND4 (N1439, N1424, N438, N1264, N125);
buf BUF1 (N1440, N1432);
xor XOR2 (N1441, N1437, N1243);
xor XOR2 (N1442, N1425, N1289);
buf BUF1 (N1443, N1438);
buf BUF1 (N1444, N1431);
xor XOR2 (N1445, N1442, N1252);
nand NAND4 (N1446, N1441, N213, N318, N46);
not NOT1 (N1447, N1446);
nor NOR4 (N1448, N1433, N205, N565, N1147);
not NOT1 (N1449, N1445);
or OR2 (N1450, N1439, N844);
and AND3 (N1451, N1413, N640, N831);
nor NOR2 (N1452, N1444, N724);
or OR4 (N1453, N1450, N885, N716, N838);
buf BUF1 (N1454, N1435);
nand NAND4 (N1455, N1449, N510, N1336, N363);
not NOT1 (N1456, N1448);
nor NOR4 (N1457, N1440, N942, N31, N1286);
buf BUF1 (N1458, N1452);
or OR3 (N1459, N1454, N96, N1000);
nand NAND3 (N1460, N1443, N244, N819);
nor NOR2 (N1461, N1453, N534);
and AND2 (N1462, N1461, N489);
not NOT1 (N1463, N1458);
nand NAND2 (N1464, N1451, N1296);
and AND3 (N1465, N1455, N1454, N1085);
xor XOR2 (N1466, N1456, N99);
nand NAND2 (N1467, N1464, N502);
xor XOR2 (N1468, N1466, N1445);
or OR3 (N1469, N1467, N1213, N649);
or OR2 (N1470, N1447, N299);
and AND4 (N1471, N1468, N1051, N393, N356);
or OR3 (N1472, N1463, N1072, N757);
and AND2 (N1473, N1457, N1187);
nor NOR4 (N1474, N1411, N1375, N92, N1028);
nand NAND4 (N1475, N1465, N685, N874, N151);
or OR3 (N1476, N1474, N765, N222);
not NOT1 (N1477, N1460);
nand NAND3 (N1478, N1462, N465, N625);
buf BUF1 (N1479, N1473);
or OR3 (N1480, N1479, N1192, N1015);
buf BUF1 (N1481, N1477);
or OR4 (N1482, N1472, N1419, N830, N387);
not NOT1 (N1483, N1471);
nor NOR4 (N1484, N1469, N932, N216, N707);
not NOT1 (N1485, N1480);
and AND4 (N1486, N1481, N1131, N1443, N737);
and AND4 (N1487, N1484, N712, N297, N1395);
not NOT1 (N1488, N1485);
not NOT1 (N1489, N1478);
or OR3 (N1490, N1482, N1089, N179);
nor NOR4 (N1491, N1483, N819, N533, N1092);
buf BUF1 (N1492, N1488);
or OR3 (N1493, N1459, N58, N1095);
xor XOR2 (N1494, N1470, N121);
buf BUF1 (N1495, N1487);
and AND3 (N1496, N1486, N1075, N1382);
xor XOR2 (N1497, N1495, N527);
not NOT1 (N1498, N1494);
not NOT1 (N1499, N1493);
or OR2 (N1500, N1498, N124);
not NOT1 (N1501, N1496);
buf BUF1 (N1502, N1501);
nor NOR4 (N1503, N1500, N767, N24, N417);
nor NOR3 (N1504, N1489, N1112, N397);
nor NOR2 (N1505, N1490, N1449);
buf BUF1 (N1506, N1504);
and AND3 (N1507, N1475, N504, N1446);
nor NOR4 (N1508, N1503, N305, N399, N417);
not NOT1 (N1509, N1492);
or OR4 (N1510, N1491, N393, N1424, N1484);
nand NAND4 (N1511, N1508, N357, N783, N1015);
not NOT1 (N1512, N1497);
nand NAND4 (N1513, N1506, N1468, N1072, N531);
buf BUF1 (N1514, N1505);
nor NOR2 (N1515, N1509, N441);
nor NOR2 (N1516, N1512, N410);
and AND2 (N1517, N1499, N477);
nand NAND4 (N1518, N1515, N1244, N1331, N1297);
or OR2 (N1519, N1518, N444);
nor NOR3 (N1520, N1516, N247, N871);
buf BUF1 (N1521, N1519);
not NOT1 (N1522, N1514);
nand NAND3 (N1523, N1507, N981, N374);
or OR3 (N1524, N1510, N296, N1376);
not NOT1 (N1525, N1524);
not NOT1 (N1526, N1511);
or OR2 (N1527, N1521, N1431);
buf BUF1 (N1528, N1520);
and AND2 (N1529, N1522, N1403);
xor XOR2 (N1530, N1529, N1486);
buf BUF1 (N1531, N1502);
xor XOR2 (N1532, N1525, N1345);
or OR4 (N1533, N1523, N173, N847, N1400);
buf BUF1 (N1534, N1531);
not NOT1 (N1535, N1476);
not NOT1 (N1536, N1526);
nor NOR4 (N1537, N1517, N287, N585, N819);
and AND2 (N1538, N1534, N951);
or OR4 (N1539, N1537, N309, N30, N707);
and AND3 (N1540, N1532, N1392, N1441);
nand NAND3 (N1541, N1540, N902, N428);
xor XOR2 (N1542, N1538, N65);
nor NOR2 (N1543, N1542, N415);
not NOT1 (N1544, N1543);
buf BUF1 (N1545, N1533);
not NOT1 (N1546, N1530);
or OR4 (N1547, N1541, N1534, N1221, N469);
and AND3 (N1548, N1547, N776, N170);
buf BUF1 (N1549, N1548);
xor XOR2 (N1550, N1528, N556);
nor NOR4 (N1551, N1536, N1457, N702, N730);
nand NAND3 (N1552, N1544, N399, N685);
xor XOR2 (N1553, N1546, N466);
xor XOR2 (N1554, N1539, N808);
buf BUF1 (N1555, N1545);
and AND3 (N1556, N1527, N1172, N865);
buf BUF1 (N1557, N1552);
buf BUF1 (N1558, N1554);
or OR3 (N1559, N1550, N616, N377);
and AND3 (N1560, N1551, N427, N454);
or OR3 (N1561, N1556, N775, N528);
nor NOR2 (N1562, N1559, N794);
not NOT1 (N1563, N1557);
xor XOR2 (N1564, N1558, N251);
and AND3 (N1565, N1555, N1499, N159);
or OR2 (N1566, N1513, N451);
not NOT1 (N1567, N1560);
and AND2 (N1568, N1549, N431);
buf BUF1 (N1569, N1553);
nand NAND4 (N1570, N1569, N1238, N1434, N1300);
not NOT1 (N1571, N1566);
not NOT1 (N1572, N1562);
not NOT1 (N1573, N1563);
nand NAND4 (N1574, N1570, N495, N494, N656);
xor XOR2 (N1575, N1572, N15);
buf BUF1 (N1576, N1565);
or OR4 (N1577, N1576, N1210, N737, N1237);
xor XOR2 (N1578, N1577, N1258);
buf BUF1 (N1579, N1564);
xor XOR2 (N1580, N1535, N221);
or OR4 (N1581, N1580, N579, N596, N306);
or OR4 (N1582, N1579, N884, N1039, N1476);
nor NOR4 (N1583, N1561, N622, N108, N728);
not NOT1 (N1584, N1582);
nor NOR3 (N1585, N1567, N1561, N983);
and AND3 (N1586, N1571, N1057, N1439);
buf BUF1 (N1587, N1584);
not NOT1 (N1588, N1568);
buf BUF1 (N1589, N1575);
xor XOR2 (N1590, N1583, N1144);
or OR4 (N1591, N1574, N289, N21, N485);
and AND3 (N1592, N1581, N1477, N997);
buf BUF1 (N1593, N1588);
buf BUF1 (N1594, N1573);
xor XOR2 (N1595, N1594, N1063);
nand NAND2 (N1596, N1593, N221);
nor NOR2 (N1597, N1592, N705);
not NOT1 (N1598, N1596);
nor NOR2 (N1599, N1595, N1409);
and AND2 (N1600, N1597, N46);
or OR2 (N1601, N1589, N1328);
nor NOR2 (N1602, N1578, N494);
nand NAND3 (N1603, N1602, N256, N1399);
not NOT1 (N1604, N1586);
or OR2 (N1605, N1585, N860);
xor XOR2 (N1606, N1591, N316);
buf BUF1 (N1607, N1603);
buf BUF1 (N1608, N1600);
xor XOR2 (N1609, N1606, N637);
and AND3 (N1610, N1587, N1282, N408);
and AND3 (N1611, N1607, N763, N980);
buf BUF1 (N1612, N1608);
nor NOR3 (N1613, N1611, N278, N1245);
buf BUF1 (N1614, N1604);
nor NOR3 (N1615, N1601, N1234, N509);
or OR2 (N1616, N1599, N1570);
xor XOR2 (N1617, N1612, N1074);
nor NOR4 (N1618, N1613, N103, N1109, N682);
nand NAND3 (N1619, N1598, N1387, N317);
xor XOR2 (N1620, N1590, N204);
and AND3 (N1621, N1615, N19, N1351);
xor XOR2 (N1622, N1617, N767);
buf BUF1 (N1623, N1614);
xor XOR2 (N1624, N1605, N805);
buf BUF1 (N1625, N1610);
xor XOR2 (N1626, N1619, N428);
nor NOR2 (N1627, N1624, N927);
and AND2 (N1628, N1622, N4);
nand NAND3 (N1629, N1609, N248, N460);
nand NAND4 (N1630, N1626, N607, N1098, N41);
and AND3 (N1631, N1620, N172, N201);
nor NOR2 (N1632, N1618, N558);
buf BUF1 (N1633, N1627);
xor XOR2 (N1634, N1623, N794);
nor NOR2 (N1635, N1631, N188);
nand NAND2 (N1636, N1635, N528);
not NOT1 (N1637, N1636);
nand NAND2 (N1638, N1629, N943);
not NOT1 (N1639, N1632);
buf BUF1 (N1640, N1637);
nand NAND2 (N1641, N1634, N1205);
and AND2 (N1642, N1641, N972);
xor XOR2 (N1643, N1625, N551);
nor NOR3 (N1644, N1628, N98, N711);
nor NOR3 (N1645, N1630, N856, N1398);
nor NOR2 (N1646, N1633, N183);
or OR3 (N1647, N1643, N869, N627);
xor XOR2 (N1648, N1621, N1429);
nor NOR4 (N1649, N1644, N911, N540, N101);
and AND3 (N1650, N1639, N1150, N1073);
and AND3 (N1651, N1616, N1615, N1503);
or OR2 (N1652, N1647, N868);
xor XOR2 (N1653, N1651, N380);
nand NAND2 (N1654, N1653, N1503);
or OR4 (N1655, N1652, N823, N1601, N842);
nor NOR4 (N1656, N1649, N185, N541, N1471);
buf BUF1 (N1657, N1638);
nand NAND2 (N1658, N1645, N181);
xor XOR2 (N1659, N1657, N872);
or OR2 (N1660, N1654, N905);
nor NOR3 (N1661, N1660, N1463, N1358);
nand NAND3 (N1662, N1640, N1389, N1228);
nand NAND3 (N1663, N1646, N798, N357);
and AND2 (N1664, N1661, N340);
nand NAND3 (N1665, N1648, N1483, N1516);
nand NAND3 (N1666, N1665, N1326, N1610);
not NOT1 (N1667, N1659);
buf BUF1 (N1668, N1662);
not NOT1 (N1669, N1664);
not NOT1 (N1670, N1658);
buf BUF1 (N1671, N1656);
or OR4 (N1672, N1670, N710, N1482, N1569);
and AND3 (N1673, N1663, N988, N115);
not NOT1 (N1674, N1655);
or OR4 (N1675, N1672, N1060, N687, N53);
or OR2 (N1676, N1642, N1018);
or OR3 (N1677, N1671, N188, N424);
and AND4 (N1678, N1676, N168, N262, N1380);
or OR2 (N1679, N1677, N1000);
xor XOR2 (N1680, N1650, N799);
and AND4 (N1681, N1675, N58, N1463, N328);
nor NOR3 (N1682, N1678, N1426, N24);
buf BUF1 (N1683, N1681);
xor XOR2 (N1684, N1669, N1208);
nand NAND2 (N1685, N1667, N301);
and AND2 (N1686, N1666, N23);
not NOT1 (N1687, N1680);
nor NOR4 (N1688, N1668, N959, N1588, N1103);
nor NOR4 (N1689, N1682, N920, N624, N1143);
nand NAND4 (N1690, N1673, N1415, N69, N1569);
buf BUF1 (N1691, N1689);
buf BUF1 (N1692, N1683);
nand NAND2 (N1693, N1684, N743);
or OR2 (N1694, N1679, N1143);
and AND2 (N1695, N1685, N1247);
or OR2 (N1696, N1693, N900);
and AND3 (N1697, N1694, N215, N520);
nand NAND4 (N1698, N1695, N1527, N1360, N25);
nand NAND3 (N1699, N1698, N320, N36);
buf BUF1 (N1700, N1688);
or OR4 (N1701, N1700, N817, N401, N94);
or OR4 (N1702, N1687, N456, N1127, N1631);
and AND4 (N1703, N1690, N1511, N1033, N1580);
and AND4 (N1704, N1699, N884, N1100, N1631);
nand NAND4 (N1705, N1703, N682, N1627, N1544);
not NOT1 (N1706, N1674);
not NOT1 (N1707, N1686);
or OR4 (N1708, N1697, N705, N1105, N365);
and AND2 (N1709, N1691, N1044);
or OR3 (N1710, N1709, N466, N419);
buf BUF1 (N1711, N1705);
xor XOR2 (N1712, N1696, N769);
xor XOR2 (N1713, N1706, N1236);
nand NAND3 (N1714, N1701, N304, N149);
not NOT1 (N1715, N1702);
xor XOR2 (N1716, N1714, N298);
buf BUF1 (N1717, N1704);
not NOT1 (N1718, N1708);
xor XOR2 (N1719, N1716, N234);
not NOT1 (N1720, N1715);
not NOT1 (N1721, N1720);
and AND3 (N1722, N1712, N887, N1669);
and AND4 (N1723, N1717, N873, N1622, N217);
not NOT1 (N1724, N1723);
xor XOR2 (N1725, N1724, N695);
or OR3 (N1726, N1692, N1658, N1185);
nor NOR3 (N1727, N1726, N629, N1258);
not NOT1 (N1728, N1725);
nor NOR3 (N1729, N1713, N681, N570);
nand NAND2 (N1730, N1711, N1518);
not NOT1 (N1731, N1719);
xor XOR2 (N1732, N1707, N392);
or OR3 (N1733, N1718, N1554, N132);
not NOT1 (N1734, N1731);
buf BUF1 (N1735, N1722);
nor NOR2 (N1736, N1721, N781);
not NOT1 (N1737, N1734);
xor XOR2 (N1738, N1727, N758);
and AND2 (N1739, N1736, N191);
or OR2 (N1740, N1730, N1526);
not NOT1 (N1741, N1728);
xor XOR2 (N1742, N1710, N226);
buf BUF1 (N1743, N1732);
xor XOR2 (N1744, N1729, N4);
nor NOR2 (N1745, N1740, N1714);
xor XOR2 (N1746, N1744, N816);
or OR4 (N1747, N1737, N868, N1455, N911);
buf BUF1 (N1748, N1746);
xor XOR2 (N1749, N1748, N1026);
xor XOR2 (N1750, N1735, N1648);
and AND3 (N1751, N1742, N44, N210);
not NOT1 (N1752, N1745);
not NOT1 (N1753, N1747);
or OR4 (N1754, N1751, N311, N1483, N1229);
not NOT1 (N1755, N1752);
nor NOR2 (N1756, N1750, N358);
buf BUF1 (N1757, N1754);
nand NAND2 (N1758, N1733, N937);
nor NOR4 (N1759, N1743, N320, N1220, N353);
not NOT1 (N1760, N1756);
nor NOR4 (N1761, N1759, N1096, N1136, N1219);
xor XOR2 (N1762, N1757, N1324);
not NOT1 (N1763, N1760);
and AND3 (N1764, N1763, N1353, N1626);
and AND2 (N1765, N1739, N460);
buf BUF1 (N1766, N1764);
xor XOR2 (N1767, N1741, N87);
or OR4 (N1768, N1761, N728, N929, N972);
nor NOR3 (N1769, N1762, N247, N1187);
xor XOR2 (N1770, N1738, N1235);
nand NAND2 (N1771, N1758, N1439);
nand NAND3 (N1772, N1766, N824, N183);
and AND2 (N1773, N1770, N679);
or OR4 (N1774, N1771, N731, N1622, N1628);
xor XOR2 (N1775, N1773, N1096);
and AND3 (N1776, N1753, N381, N1712);
nand NAND3 (N1777, N1776, N875, N840);
xor XOR2 (N1778, N1777, N1517);
nand NAND4 (N1779, N1772, N542, N1537, N310);
or OR4 (N1780, N1775, N1749, N1630, N1773);
not NOT1 (N1781, N1236);
nor NOR3 (N1782, N1778, N550, N1750);
xor XOR2 (N1783, N1769, N734);
nor NOR2 (N1784, N1783, N1125);
not NOT1 (N1785, N1780);
or OR2 (N1786, N1768, N1353);
xor XOR2 (N1787, N1785, N77);
xor XOR2 (N1788, N1779, N344);
not NOT1 (N1789, N1788);
not NOT1 (N1790, N1786);
buf BUF1 (N1791, N1765);
not NOT1 (N1792, N1781);
not NOT1 (N1793, N1787);
buf BUF1 (N1794, N1782);
buf BUF1 (N1795, N1790);
xor XOR2 (N1796, N1789, N995);
xor XOR2 (N1797, N1767, N795);
nand NAND3 (N1798, N1793, N57, N662);
buf BUF1 (N1799, N1794);
buf BUF1 (N1800, N1797);
or OR4 (N1801, N1799, N1181, N802, N181);
not NOT1 (N1802, N1755);
nand NAND3 (N1803, N1784, N1133, N1209);
and AND2 (N1804, N1774, N1772);
nor NOR2 (N1805, N1796, N4);
buf BUF1 (N1806, N1798);
and AND2 (N1807, N1804, N1522);
xor XOR2 (N1808, N1800, N970);
not NOT1 (N1809, N1801);
or OR3 (N1810, N1803, N1500, N1702);
not NOT1 (N1811, N1795);
not NOT1 (N1812, N1811);
or OR4 (N1813, N1806, N1044, N174, N901);
buf BUF1 (N1814, N1813);
buf BUF1 (N1815, N1792);
nand NAND2 (N1816, N1815, N556);
nand NAND3 (N1817, N1805, N1538, N137);
xor XOR2 (N1818, N1817, N564);
and AND3 (N1819, N1814, N1199, N1322);
or OR4 (N1820, N1818, N1634, N1375, N1628);
nand NAND3 (N1821, N1809, N1475, N1482);
or OR4 (N1822, N1819, N1704, N1765, N816);
not NOT1 (N1823, N1822);
or OR4 (N1824, N1812, N1627, N1571, N379);
buf BUF1 (N1825, N1816);
xor XOR2 (N1826, N1802, N268);
buf BUF1 (N1827, N1810);
and AND3 (N1828, N1807, N407, N1015);
xor XOR2 (N1829, N1791, N1809);
or OR4 (N1830, N1821, N1070, N590, N57);
and AND3 (N1831, N1826, N1313, N308);
and AND3 (N1832, N1831, N1614, N686);
nand NAND3 (N1833, N1829, N351, N1817);
and AND3 (N1834, N1827, N618, N1030);
or OR4 (N1835, N1832, N31, N714, N926);
xor XOR2 (N1836, N1820, N299);
nand NAND4 (N1837, N1824, N31, N1068, N1042);
not NOT1 (N1838, N1828);
nor NOR2 (N1839, N1834, N1513);
not NOT1 (N1840, N1808);
and AND2 (N1841, N1823, N203);
buf BUF1 (N1842, N1837);
or OR4 (N1843, N1840, N1406, N501, N315);
not NOT1 (N1844, N1841);
and AND2 (N1845, N1844, N1094);
nor NOR3 (N1846, N1842, N1109, N399);
nor NOR4 (N1847, N1839, N1516, N109, N1140);
nor NOR4 (N1848, N1833, N673, N663, N521);
xor XOR2 (N1849, N1843, N786);
or OR3 (N1850, N1846, N741, N345);
buf BUF1 (N1851, N1849);
nand NAND3 (N1852, N1850, N26, N1376);
and AND2 (N1853, N1835, N144);
and AND2 (N1854, N1848, N1302);
nand NAND2 (N1855, N1847, N595);
not NOT1 (N1856, N1838);
nor NOR2 (N1857, N1830, N785);
not NOT1 (N1858, N1855);
not NOT1 (N1859, N1852);
and AND3 (N1860, N1845, N174, N477);
or OR2 (N1861, N1856, N32);
buf BUF1 (N1862, N1861);
not NOT1 (N1863, N1858);
nand NAND3 (N1864, N1862, N1851, N668);
or OR3 (N1865, N765, N18, N1126);
and AND2 (N1866, N1825, N143);
xor XOR2 (N1867, N1853, N1729);
xor XOR2 (N1868, N1864, N685);
and AND3 (N1869, N1859, N1228, N869);
buf BUF1 (N1870, N1863);
buf BUF1 (N1871, N1854);
not NOT1 (N1872, N1857);
not NOT1 (N1873, N1860);
and AND3 (N1874, N1868, N449, N706);
xor XOR2 (N1875, N1873, N314);
and AND3 (N1876, N1867, N1733, N663);
not NOT1 (N1877, N1875);
nor NOR2 (N1878, N1866, N1400);
buf BUF1 (N1879, N1870);
nor NOR3 (N1880, N1874, N1225, N1449);
nand NAND4 (N1881, N1880, N269, N951, N1691);
nor NOR2 (N1882, N1871, N648);
nand NAND4 (N1883, N1882, N283, N1697, N429);
and AND4 (N1884, N1876, N108, N511, N1098);
xor XOR2 (N1885, N1878, N254);
xor XOR2 (N1886, N1885, N601);
or OR2 (N1887, N1865, N1405);
nor NOR4 (N1888, N1869, N291, N1449, N1345);
buf BUF1 (N1889, N1884);
nor NOR2 (N1890, N1877, N1235);
and AND2 (N1891, N1872, N1062);
not NOT1 (N1892, N1836);
nand NAND3 (N1893, N1890, N81, N1084);
not NOT1 (N1894, N1879);
xor XOR2 (N1895, N1892, N94);
or OR3 (N1896, N1883, N33, N631);
not NOT1 (N1897, N1889);
buf BUF1 (N1898, N1886);
nor NOR4 (N1899, N1891, N1877, N1107, N824);
buf BUF1 (N1900, N1896);
not NOT1 (N1901, N1893);
xor XOR2 (N1902, N1900, N1294);
and AND2 (N1903, N1902, N422);
nand NAND4 (N1904, N1894, N1525, N328, N998);
and AND3 (N1905, N1897, N1070, N557);
and AND2 (N1906, N1898, N1510);
nor NOR3 (N1907, N1887, N1363, N26);
buf BUF1 (N1908, N1907);
buf BUF1 (N1909, N1881);
or OR4 (N1910, N1905, N1358, N650, N681);
xor XOR2 (N1911, N1895, N258);
nor NOR2 (N1912, N1901, N696);
nand NAND4 (N1913, N1903, N1771, N382, N1794);
xor XOR2 (N1914, N1913, N1792);
buf BUF1 (N1915, N1910);
or OR3 (N1916, N1912, N1442, N1386);
nor NOR4 (N1917, N1908, N527, N1497, N1625);
nand NAND4 (N1918, N1914, N59, N1686, N1572);
not NOT1 (N1919, N1916);
nor NOR4 (N1920, N1919, N751, N515, N184);
or OR3 (N1921, N1909, N1730, N863);
and AND4 (N1922, N1911, N1544, N1547, N1502);
and AND4 (N1923, N1899, N93, N1921, N1174);
nand NAND2 (N1924, N626, N999);
nand NAND4 (N1925, N1888, N44, N1609, N1357);
or OR3 (N1926, N1917, N694, N33);
or OR3 (N1927, N1906, N1708, N531);
and AND3 (N1928, N1904, N558, N1703);
nor NOR2 (N1929, N1920, N1754);
and AND2 (N1930, N1923, N557);
and AND3 (N1931, N1918, N1819, N358);
buf BUF1 (N1932, N1924);
xor XOR2 (N1933, N1927, N524);
nand NAND3 (N1934, N1933, N705, N1326);
nand NAND3 (N1935, N1932, N1826, N1073);
nand NAND2 (N1936, N1926, N142);
not NOT1 (N1937, N1930);
and AND4 (N1938, N1936, N576, N1205, N1135);
nand NAND4 (N1939, N1938, N1509, N1883, N1865);
nor NOR2 (N1940, N1915, N957);
nor NOR3 (N1941, N1935, N1692, N829);
buf BUF1 (N1942, N1929);
nor NOR2 (N1943, N1925, N718);
or OR4 (N1944, N1939, N470, N1914, N1292);
nand NAND4 (N1945, N1934, N166, N1689, N80);
or OR3 (N1946, N1931, N1504, N117);
nor NOR3 (N1947, N1941, N1049, N1438);
buf BUF1 (N1948, N1940);
xor XOR2 (N1949, N1922, N378);
nor NOR4 (N1950, N1928, N818, N389, N176);
xor XOR2 (N1951, N1949, N1053);
and AND2 (N1952, N1942, N47);
xor XOR2 (N1953, N1948, N999);
not NOT1 (N1954, N1945);
nor NOR2 (N1955, N1954, N685);
buf BUF1 (N1956, N1943);
or OR4 (N1957, N1946, N546, N1539, N725);
xor XOR2 (N1958, N1944, N1708);
nor NOR2 (N1959, N1952, N1404);
or OR2 (N1960, N1957, N1847);
buf BUF1 (N1961, N1960);
or OR4 (N1962, N1951, N765, N256, N393);
xor XOR2 (N1963, N1958, N225);
nor NOR3 (N1964, N1953, N1852, N1888);
or OR3 (N1965, N1961, N515, N783);
and AND4 (N1966, N1950, N1551, N264, N883);
and AND2 (N1967, N1964, N1938);
xor XOR2 (N1968, N1956, N990);
not NOT1 (N1969, N1937);
xor XOR2 (N1970, N1966, N49);
and AND2 (N1971, N1968, N925);
xor XOR2 (N1972, N1947, N953);
and AND3 (N1973, N1971, N800, N828);
not NOT1 (N1974, N1955);
nor NOR3 (N1975, N1967, N1828, N1183);
not NOT1 (N1976, N1963);
nor NOR2 (N1977, N1959, N1015);
nand NAND3 (N1978, N1976, N262, N1567);
or OR4 (N1979, N1974, N1905, N628, N479);
xor XOR2 (N1980, N1978, N124);
buf BUF1 (N1981, N1979);
or OR2 (N1982, N1972, N1976);
and AND3 (N1983, N1982, N1734, N956);
buf BUF1 (N1984, N1969);
buf BUF1 (N1985, N1981);
xor XOR2 (N1986, N1980, N1537);
xor XOR2 (N1987, N1965, N273);
not NOT1 (N1988, N1984);
nor NOR2 (N1989, N1987, N1786);
nand NAND2 (N1990, N1975, N1068);
xor XOR2 (N1991, N1983, N1192);
or OR2 (N1992, N1973, N1902);
and AND4 (N1993, N1985, N426, N178, N861);
xor XOR2 (N1994, N1962, N1185);
nand NAND3 (N1995, N1993, N1983, N770);
and AND2 (N1996, N1970, N763);
xor XOR2 (N1997, N1992, N1701);
nor NOR2 (N1998, N1991, N1370);
or OR3 (N1999, N1994, N1984, N1769);
and AND2 (N2000, N1986, N577);
nor NOR2 (N2001, N2000, N1077);
buf BUF1 (N2002, N1996);
not NOT1 (N2003, N1988);
nor NOR2 (N2004, N1998, N177);
nand NAND4 (N2005, N1995, N1628, N1428, N769);
or OR4 (N2006, N1977, N748, N1349, N527);
not NOT1 (N2007, N2002);
xor XOR2 (N2008, N2007, N1589);
buf BUF1 (N2009, N2008);
buf BUF1 (N2010, N1997);
nand NAND2 (N2011, N2010, N1047);
and AND3 (N2012, N2003, N1353, N1817);
and AND4 (N2013, N2005, N1005, N1310, N911);
nand NAND3 (N2014, N1999, N922, N1733);
or OR4 (N2015, N2012, N1845, N1761, N1148);
or OR3 (N2016, N1989, N946, N524);
not NOT1 (N2017, N2011);
xor XOR2 (N2018, N2017, N816);
xor XOR2 (N2019, N2016, N1428);
xor XOR2 (N2020, N2006, N1063);
or OR3 (N2021, N2018, N1515, N2009);
not NOT1 (N2022, N457);
nor NOR4 (N2023, N2014, N2019, N755, N1197);
buf BUF1 (N2024, N1019);
nand NAND4 (N2025, N2004, N24, N1474, N1770);
nor NOR3 (N2026, N2024, N1779, N377);
and AND3 (N2027, N2025, N1061, N527);
or OR2 (N2028, N2026, N1574);
xor XOR2 (N2029, N2001, N1786);
not NOT1 (N2030, N2022);
nand NAND4 (N2031, N2030, N1463, N1254, N1605);
xor XOR2 (N2032, N2031, N1772);
buf BUF1 (N2033, N2021);
xor XOR2 (N2034, N2033, N1670);
or OR4 (N2035, N2028, N916, N661, N1568);
or OR3 (N2036, N2020, N467, N1337);
nand NAND3 (N2037, N2032, N1480, N1715);
or OR3 (N2038, N2035, N744, N902);
nor NOR2 (N2039, N1990, N1653);
or OR2 (N2040, N2037, N134);
buf BUF1 (N2041, N2040);
xor XOR2 (N2042, N2027, N224);
or OR4 (N2043, N2038, N387, N1270, N5);
not NOT1 (N2044, N2036);
or OR3 (N2045, N2042, N498, N1286);
and AND3 (N2046, N2034, N1613, N267);
xor XOR2 (N2047, N2015, N411);
nor NOR2 (N2048, N2039, N398);
or OR2 (N2049, N2048, N130);
buf BUF1 (N2050, N2047);
not NOT1 (N2051, N2041);
xor XOR2 (N2052, N2051, N378);
buf BUF1 (N2053, N2013);
or OR3 (N2054, N2046, N146, N1833);
or OR4 (N2055, N2045, N2003, N596, N917);
buf BUF1 (N2056, N2049);
nor NOR3 (N2057, N2029, N46, N802);
and AND4 (N2058, N2050, N1706, N147, N2049);
buf BUF1 (N2059, N2053);
not NOT1 (N2060, N2044);
nand NAND4 (N2061, N2058, N1953, N1256, N470);
or OR4 (N2062, N2052, N1214, N1312, N1429);
not NOT1 (N2063, N2059);
not NOT1 (N2064, N2056);
xor XOR2 (N2065, N2043, N307);
nand NAND4 (N2066, N2060, N83, N1990, N329);
not NOT1 (N2067, N2054);
and AND4 (N2068, N2055, N469, N1217, N1069);
or OR2 (N2069, N2068, N1386);
or OR2 (N2070, N2061, N413);
nor NOR2 (N2071, N2064, N1139);
and AND3 (N2072, N2063, N1579, N610);
xor XOR2 (N2073, N2071, N1907);
and AND3 (N2074, N2065, N1305, N78);
not NOT1 (N2075, N2070);
or OR2 (N2076, N2075, N637);
nor NOR3 (N2077, N2057, N824, N2074);
nand NAND3 (N2078, N2066, N2007, N422);
or OR3 (N2079, N444, N207, N1150);
nand NAND3 (N2080, N2077, N247, N1543);
and AND3 (N2081, N2072, N1925, N1761);
and AND3 (N2082, N2023, N1525, N1749);
nand NAND3 (N2083, N2067, N725, N790);
not NOT1 (N2084, N2080);
nand NAND3 (N2085, N2084, N1155, N272);
buf BUF1 (N2086, N2062);
xor XOR2 (N2087, N2081, N555);
buf BUF1 (N2088, N2082);
nor NOR3 (N2089, N2076, N535, N1524);
nand NAND4 (N2090, N2073, N891, N237, N1708);
or OR3 (N2091, N2087, N1351, N566);
nor NOR4 (N2092, N2088, N391, N44, N2003);
nor NOR2 (N2093, N2092, N2088);
nand NAND2 (N2094, N2091, N1151);
and AND4 (N2095, N2079, N2007, N1866, N1131);
nor NOR3 (N2096, N2094, N803, N383);
not NOT1 (N2097, N2083);
nand NAND3 (N2098, N2085, N475, N1771);
and AND3 (N2099, N2093, N1575, N462);
nor NOR4 (N2100, N2099, N1850, N1623, N669);
and AND2 (N2101, N2096, N911);
nand NAND4 (N2102, N2086, N324, N1546, N1749);
buf BUF1 (N2103, N2102);
not NOT1 (N2104, N2089);
nor NOR2 (N2105, N2090, N1261);
buf BUF1 (N2106, N2103);
nor NOR3 (N2107, N2078, N505, N1228);
nor NOR2 (N2108, N2069, N282);
buf BUF1 (N2109, N2108);
nand NAND2 (N2110, N2104, N383);
nor NOR3 (N2111, N2098, N1168, N467);
or OR2 (N2112, N2111, N98);
nor NOR3 (N2113, N2101, N1572, N1745);
or OR2 (N2114, N2109, N1440);
or OR2 (N2115, N2095, N263);
and AND4 (N2116, N2115, N1486, N1686, N774);
nor NOR2 (N2117, N2100, N1604);
nand NAND4 (N2118, N2116, N1891, N1094, N1947);
or OR3 (N2119, N2118, N1316, N1033);
not NOT1 (N2120, N2113);
and AND4 (N2121, N2114, N1787, N1196, N2101);
xor XOR2 (N2122, N2112, N979);
and AND2 (N2123, N2107, N71);
and AND4 (N2124, N2123, N1629, N206, N1938);
or OR2 (N2125, N2106, N1200);
or OR2 (N2126, N2121, N1202);
and AND4 (N2127, N2119, N1082, N1751, N1491);
buf BUF1 (N2128, N2127);
buf BUF1 (N2129, N2128);
buf BUF1 (N2130, N2129);
nand NAND4 (N2131, N2117, N1940, N94, N1742);
not NOT1 (N2132, N2110);
and AND3 (N2133, N2097, N584, N770);
and AND4 (N2134, N2105, N2013, N185, N677);
buf BUF1 (N2135, N2126);
buf BUF1 (N2136, N2135);
or OR4 (N2137, N2134, N729, N234, N635);
or OR4 (N2138, N2133, N688, N1388, N1056);
xor XOR2 (N2139, N2124, N420);
nand NAND3 (N2140, N2139, N253, N396);
and AND3 (N2141, N2138, N935, N266);
not NOT1 (N2142, N2141);
xor XOR2 (N2143, N2132, N16);
nor NOR2 (N2144, N2122, N1598);
nand NAND2 (N2145, N2140, N807);
nand NAND2 (N2146, N2144, N745);
and AND2 (N2147, N2125, N413);
xor XOR2 (N2148, N2142, N1890);
xor XOR2 (N2149, N2146, N1139);
or OR2 (N2150, N2149, N1628);
nand NAND4 (N2151, N2143, N529, N1464, N1099);
xor XOR2 (N2152, N2130, N1558);
and AND4 (N2153, N2150, N1738, N934, N1980);
or OR2 (N2154, N2151, N1613);
xor XOR2 (N2155, N2136, N770);
or OR3 (N2156, N2131, N2095, N1547);
buf BUF1 (N2157, N2155);
or OR4 (N2158, N2120, N1986, N548, N216);
and AND3 (N2159, N2152, N317, N1147);
xor XOR2 (N2160, N2154, N611);
nand NAND2 (N2161, N2145, N135);
nand NAND2 (N2162, N2157, N1704);
xor XOR2 (N2163, N2159, N1228);
or OR4 (N2164, N2162, N1092, N1233, N1508);
nand NAND3 (N2165, N2164, N2101, N925);
not NOT1 (N2166, N2156);
buf BUF1 (N2167, N2166);
and AND3 (N2168, N2147, N2144, N817);
xor XOR2 (N2169, N2160, N617);
or OR2 (N2170, N2137, N1316);
not NOT1 (N2171, N2158);
and AND4 (N2172, N2171, N1878, N797, N967);
nor NOR4 (N2173, N2169, N1722, N1554, N900);
or OR2 (N2174, N2172, N1457);
not NOT1 (N2175, N2167);
or OR3 (N2176, N2153, N1226, N1657);
nand NAND2 (N2177, N2168, N1163);
buf BUF1 (N2178, N2173);
nor NOR2 (N2179, N2178, N284);
nor NOR2 (N2180, N2163, N1696);
nor NOR2 (N2181, N2170, N335);
buf BUF1 (N2182, N2165);
nor NOR3 (N2183, N2180, N325, N1642);
and AND3 (N2184, N2174, N1736, N1451);
nand NAND2 (N2185, N2182, N2062);
buf BUF1 (N2186, N2184);
nand NAND4 (N2187, N2183, N403, N251, N1111);
not NOT1 (N2188, N2185);
nor NOR4 (N2189, N2161, N2094, N1118, N727);
buf BUF1 (N2190, N2177);
not NOT1 (N2191, N2187);
xor XOR2 (N2192, N2176, N370);
xor XOR2 (N2193, N2192, N296);
buf BUF1 (N2194, N2186);
nand NAND4 (N2195, N2179, N354, N296, N198);
nand NAND4 (N2196, N2181, N1432, N912, N1983);
not NOT1 (N2197, N2195);
xor XOR2 (N2198, N2148, N2009);
nor NOR3 (N2199, N2191, N819, N1195);
and AND2 (N2200, N2199, N947);
xor XOR2 (N2201, N2175, N1462);
buf BUF1 (N2202, N2197);
nor NOR4 (N2203, N2188, N546, N684, N425);
buf BUF1 (N2204, N2193);
and AND2 (N2205, N2190, N650);
nor NOR2 (N2206, N2196, N765);
not NOT1 (N2207, N2206);
or OR3 (N2208, N2200, N1568, N1345);
buf BUF1 (N2209, N2201);
and AND4 (N2210, N2198, N141, N1464, N1035);
nor NOR4 (N2211, N2207, N1546, N1786, N139);
and AND3 (N2212, N2204, N606, N1638);
nand NAND4 (N2213, N2203, N547, N160, N1419);
not NOT1 (N2214, N2208);
buf BUF1 (N2215, N2211);
or OR3 (N2216, N2214, N2108, N180);
and AND2 (N2217, N2212, N1637);
buf BUF1 (N2218, N2205);
xor XOR2 (N2219, N2217, N704);
nor NOR4 (N2220, N2216, N929, N514, N1338);
and AND3 (N2221, N2213, N2043, N1035);
and AND3 (N2222, N2221, N557, N202);
nor NOR3 (N2223, N2209, N952, N1509);
nand NAND4 (N2224, N2202, N1649, N1904, N1341);
not NOT1 (N2225, N2224);
nor NOR4 (N2226, N2218, N2010, N1900, N1178);
not NOT1 (N2227, N2220);
xor XOR2 (N2228, N2227, N2198);
nand NAND4 (N2229, N2194, N2063, N1584, N729);
xor XOR2 (N2230, N2189, N977);
and AND3 (N2231, N2210, N338, N1433);
not NOT1 (N2232, N2223);
and AND4 (N2233, N2222, N613, N2156, N1339);
xor XOR2 (N2234, N2231, N1740);
nor NOR3 (N2235, N2234, N1156, N2228);
not NOT1 (N2236, N1102);
buf BUF1 (N2237, N2232);
buf BUF1 (N2238, N2233);
buf BUF1 (N2239, N2219);
nand NAND4 (N2240, N2238, N4, N528, N1745);
and AND3 (N2241, N2235, N473, N1398);
xor XOR2 (N2242, N2240, N740);
buf BUF1 (N2243, N2239);
xor XOR2 (N2244, N2229, N513);
nor NOR2 (N2245, N2225, N201);
or OR2 (N2246, N2236, N1219);
and AND4 (N2247, N2245, N405, N1935, N1171);
and AND3 (N2248, N2243, N2241, N2242);
xor XOR2 (N2249, N955, N1874);
and AND2 (N2250, N1019, N1072);
or OR2 (N2251, N2250, N254);
not NOT1 (N2252, N2248);
and AND2 (N2253, N2226, N684);
not NOT1 (N2254, N2249);
or OR2 (N2255, N2244, N2115);
not NOT1 (N2256, N2230);
nor NOR2 (N2257, N2237, N2011);
xor XOR2 (N2258, N2251, N2062);
not NOT1 (N2259, N2247);
and AND3 (N2260, N2259, N1941, N311);
nand NAND2 (N2261, N2215, N1249);
nor NOR2 (N2262, N2258, N610);
xor XOR2 (N2263, N2253, N1556);
buf BUF1 (N2264, N2262);
and AND3 (N2265, N2261, N1566, N1556);
nor NOR3 (N2266, N2246, N1042, N318);
and AND4 (N2267, N2254, N501, N1801, N1725);
buf BUF1 (N2268, N2267);
nor NOR2 (N2269, N2265, N1005);
xor XOR2 (N2270, N2266, N112);
buf BUF1 (N2271, N2264);
buf BUF1 (N2272, N2256);
xor XOR2 (N2273, N2255, N700);
and AND4 (N2274, N2269, N1326, N1349, N601);
and AND2 (N2275, N2257, N2140);
nand NAND4 (N2276, N2272, N1782, N487, N1371);
not NOT1 (N2277, N2273);
not NOT1 (N2278, N2252);
not NOT1 (N2279, N2276);
nand NAND4 (N2280, N2268, N1726, N1587, N12);
nor NOR3 (N2281, N2277, N1298, N366);
and AND4 (N2282, N2274, N1917, N24, N512);
xor XOR2 (N2283, N2271, N854);
not NOT1 (N2284, N2270);
buf BUF1 (N2285, N2284);
xor XOR2 (N2286, N2285, N1824);
not NOT1 (N2287, N2281);
and AND3 (N2288, N2280, N778, N790);
and AND2 (N2289, N2283, N178);
xor XOR2 (N2290, N2288, N475);
buf BUF1 (N2291, N2263);
and AND2 (N2292, N2282, N660);
not NOT1 (N2293, N2287);
xor XOR2 (N2294, N2279, N52);
xor XOR2 (N2295, N2278, N1086);
buf BUF1 (N2296, N2289);
and AND3 (N2297, N2292, N79, N1904);
or OR4 (N2298, N2291, N1065, N1170, N2105);
nor NOR2 (N2299, N2296, N1110);
or OR3 (N2300, N2295, N1010, N1880);
buf BUF1 (N2301, N2294);
xor XOR2 (N2302, N2286, N1785);
nand NAND2 (N2303, N2301, N1350);
nor NOR4 (N2304, N2275, N2215, N194, N1052);
xor XOR2 (N2305, N2298, N38);
nand NAND3 (N2306, N2302, N1719, N431);
or OR2 (N2307, N2300, N2021);
xor XOR2 (N2308, N2290, N868);
not NOT1 (N2309, N2304);
xor XOR2 (N2310, N2308, N88);
nor NOR3 (N2311, N2307, N1936, N402);
or OR3 (N2312, N2306, N946, N2302);
nor NOR3 (N2313, N2297, N676, N1324);
and AND2 (N2314, N2303, N2032);
and AND4 (N2315, N2293, N2216, N532, N1490);
nand NAND3 (N2316, N2313, N1218, N261);
and AND3 (N2317, N2260, N498, N1176);
not NOT1 (N2318, N2309);
or OR3 (N2319, N2312, N919, N1567);
buf BUF1 (N2320, N2299);
nor NOR2 (N2321, N2305, N1446);
and AND4 (N2322, N2311, N1222, N542, N114);
not NOT1 (N2323, N2317);
and AND2 (N2324, N2310, N559);
or OR2 (N2325, N2315, N965);
or OR2 (N2326, N2320, N1343);
and AND2 (N2327, N2318, N1218);
nor NOR4 (N2328, N2319, N1414, N429, N1720);
and AND3 (N2329, N2316, N1670, N883);
not NOT1 (N2330, N2323);
and AND4 (N2331, N2328, N458, N1149, N769);
xor XOR2 (N2332, N2322, N1765);
or OR3 (N2333, N2314, N871, N925);
not NOT1 (N2334, N2327);
nor NOR3 (N2335, N2329, N327, N1605);
not NOT1 (N2336, N2331);
xor XOR2 (N2337, N2321, N1577);
xor XOR2 (N2338, N2330, N1501);
not NOT1 (N2339, N2337);
xor XOR2 (N2340, N2336, N1062);
nor NOR2 (N2341, N2339, N632);
nor NOR4 (N2342, N2326, N859, N704, N973);
xor XOR2 (N2343, N2335, N1814);
or OR2 (N2344, N2340, N927);
not NOT1 (N2345, N2334);
nor NOR2 (N2346, N2344, N1527);
xor XOR2 (N2347, N2343, N166);
or OR2 (N2348, N2338, N2210);
nor NOR2 (N2349, N2342, N2337);
xor XOR2 (N2350, N2333, N1103);
or OR2 (N2351, N2341, N1316);
and AND4 (N2352, N2345, N1898, N1463, N581);
nand NAND4 (N2353, N2349, N1922, N125, N2210);
buf BUF1 (N2354, N2348);
and AND2 (N2355, N2351, N467);
nand NAND2 (N2356, N2324, N1760);
not NOT1 (N2357, N2350);
or OR3 (N2358, N2325, N1201, N2283);
buf BUF1 (N2359, N2353);
and AND3 (N2360, N2347, N866, N563);
nor NOR3 (N2361, N2354, N1230, N1181);
nor NOR2 (N2362, N2352, N823);
nor NOR4 (N2363, N2346, N938, N1998, N1241);
buf BUF1 (N2364, N2361);
xor XOR2 (N2365, N2355, N1400);
xor XOR2 (N2366, N2362, N465);
not NOT1 (N2367, N2332);
buf BUF1 (N2368, N2357);
nor NOR3 (N2369, N2364, N2340, N1736);
nor NOR4 (N2370, N2365, N1644, N742, N1430);
xor XOR2 (N2371, N2363, N702);
xor XOR2 (N2372, N2371, N1842);
not NOT1 (N2373, N2359);
not NOT1 (N2374, N2370);
nor NOR2 (N2375, N2374, N1264);
or OR2 (N2376, N2356, N2352);
nand NAND2 (N2377, N2368, N1942);
not NOT1 (N2378, N2377);
xor XOR2 (N2379, N2378, N2202);
or OR2 (N2380, N2379, N1337);
nor NOR2 (N2381, N2380, N1113);
xor XOR2 (N2382, N2367, N1116);
buf BUF1 (N2383, N2376);
xor XOR2 (N2384, N2382, N2311);
not NOT1 (N2385, N2366);
nand NAND4 (N2386, N2360, N541, N2350, N864);
and AND3 (N2387, N2358, N1684, N872);
xor XOR2 (N2388, N2373, N1006);
or OR4 (N2389, N2381, N1111, N2288, N2272);
xor XOR2 (N2390, N2383, N2143);
buf BUF1 (N2391, N2390);
not NOT1 (N2392, N2375);
nor NOR2 (N2393, N2392, N1130);
and AND4 (N2394, N2388, N2291, N700, N92);
nand NAND4 (N2395, N2391, N1980, N1280, N631);
not NOT1 (N2396, N2386);
xor XOR2 (N2397, N2387, N1614);
xor XOR2 (N2398, N2394, N1425);
xor XOR2 (N2399, N2369, N1495);
nand NAND2 (N2400, N2396, N1103);
nor NOR3 (N2401, N2399, N1731, N1570);
and AND4 (N2402, N2389, N1636, N683, N746);
not NOT1 (N2403, N2402);
or OR3 (N2404, N2397, N1393, N28);
nor NOR4 (N2405, N2384, N629, N526, N158);
not NOT1 (N2406, N2400);
nor NOR2 (N2407, N2403, N2033);
not NOT1 (N2408, N2385);
buf BUF1 (N2409, N2407);
buf BUF1 (N2410, N2395);
nand NAND4 (N2411, N2372, N2362, N995, N307);
buf BUF1 (N2412, N2405);
or OR2 (N2413, N2404, N2288);
buf BUF1 (N2414, N2411);
nand NAND2 (N2415, N2412, N2019);
or OR3 (N2416, N2410, N1089, N2134);
nand NAND2 (N2417, N2401, N242);
nor NOR4 (N2418, N2417, N954, N2085, N167);
nor NOR4 (N2419, N2393, N692, N61, N2054);
nand NAND2 (N2420, N2409, N763);
or OR2 (N2421, N2415, N1022);
not NOT1 (N2422, N2420);
nor NOR3 (N2423, N2398, N531, N674);
not NOT1 (N2424, N2408);
buf BUF1 (N2425, N2421);
xor XOR2 (N2426, N2406, N1849);
or OR4 (N2427, N2418, N1654, N1083, N2338);
or OR2 (N2428, N2425, N1093);
nand NAND3 (N2429, N2422, N287, N1558);
nor NOR3 (N2430, N2429, N2214, N1106);
nand NAND2 (N2431, N2426, N242);
nand NAND3 (N2432, N2428, N523, N168);
nand NAND2 (N2433, N2424, N1738);
or OR2 (N2434, N2416, N1421);
nor NOR2 (N2435, N2414, N1668);
or OR2 (N2436, N2431, N992);
buf BUF1 (N2437, N2432);
xor XOR2 (N2438, N2436, N11);
or OR3 (N2439, N2433, N2010, N756);
nor NOR2 (N2440, N2430, N1461);
nor NOR3 (N2441, N2440, N542, N762);
or OR4 (N2442, N2435, N2304, N2205, N785);
and AND2 (N2443, N2438, N2205);
xor XOR2 (N2444, N2434, N734);
nand NAND4 (N2445, N2444, N346, N2125, N550);
nand NAND3 (N2446, N2423, N155, N1583);
or OR2 (N2447, N2439, N670);
not NOT1 (N2448, N2443);
nand NAND3 (N2449, N2413, N736, N2119);
not NOT1 (N2450, N2445);
not NOT1 (N2451, N2446);
nand NAND2 (N2452, N2449, N1590);
or OR3 (N2453, N2419, N603, N153);
or OR4 (N2454, N2448, N1132, N2344, N798);
xor XOR2 (N2455, N2451, N1862);
xor XOR2 (N2456, N2441, N437);
xor XOR2 (N2457, N2442, N2456);
and AND3 (N2458, N1912, N92, N2166);
buf BUF1 (N2459, N2454);
xor XOR2 (N2460, N2437, N1463);
and AND4 (N2461, N2447, N2388, N1163, N308);
or OR4 (N2462, N2459, N1950, N2228, N2278);
not NOT1 (N2463, N2452);
nor NOR4 (N2464, N2450, N2387, N1461, N1203);
buf BUF1 (N2465, N2462);
buf BUF1 (N2466, N2458);
nor NOR3 (N2467, N2460, N1945, N629);
nand NAND3 (N2468, N2467, N507, N666);
not NOT1 (N2469, N2465);
buf BUF1 (N2470, N2463);
nor NOR4 (N2471, N2461, N2443, N159, N878);
nor NOR3 (N2472, N2471, N1809, N1754);
nand NAND3 (N2473, N2466, N585, N1151);
not NOT1 (N2474, N2464);
buf BUF1 (N2475, N2472);
not NOT1 (N2476, N2468);
not NOT1 (N2477, N2457);
buf BUF1 (N2478, N2477);
nor NOR4 (N2479, N2478, N1104, N2239, N1576);
and AND3 (N2480, N2455, N640, N805);
nand NAND2 (N2481, N2470, N1511);
buf BUF1 (N2482, N2427);
nor NOR2 (N2483, N2482, N360);
xor XOR2 (N2484, N2469, N1021);
buf BUF1 (N2485, N2476);
xor XOR2 (N2486, N2474, N803);
nor NOR3 (N2487, N2480, N1173, N984);
nand NAND3 (N2488, N2486, N681, N1140);
or OR3 (N2489, N2481, N1043, N89);
not NOT1 (N2490, N2483);
nor NOR3 (N2491, N2487, N649, N265);
nor NOR3 (N2492, N2490, N910, N396);
nand NAND2 (N2493, N2479, N720);
xor XOR2 (N2494, N2493, N2241);
nor NOR4 (N2495, N2494, N826, N614, N1106);
and AND3 (N2496, N2495, N117, N569);
nand NAND3 (N2497, N2484, N785, N382);
and AND3 (N2498, N2488, N170, N41);
nor NOR3 (N2499, N2491, N1803, N680);
and AND2 (N2500, N2492, N1624);
nor NOR2 (N2501, N2500, N1976);
xor XOR2 (N2502, N2499, N11);
or OR3 (N2503, N2498, N2335, N283);
xor XOR2 (N2504, N2489, N186);
or OR4 (N2505, N2502, N1705, N1630, N839);
nand NAND3 (N2506, N2501, N2290, N2323);
and AND4 (N2507, N2506, N1423, N2379, N158);
nand NAND4 (N2508, N2497, N108, N627, N782);
and AND2 (N2509, N2475, N1151);
or OR2 (N2510, N2505, N970);
or OR4 (N2511, N2503, N2449, N285, N742);
and AND3 (N2512, N2496, N1640, N1751);
buf BUF1 (N2513, N2512);
not NOT1 (N2514, N2508);
nand NAND4 (N2515, N2507, N2486, N342, N2495);
and AND4 (N2516, N2504, N1700, N848, N2073);
or OR3 (N2517, N2513, N1573, N1039);
and AND2 (N2518, N2453, N1447);
xor XOR2 (N2519, N2509, N303);
or OR4 (N2520, N2511, N2467, N1381, N546);
and AND3 (N2521, N2519, N776, N1673);
not NOT1 (N2522, N2520);
nor NOR3 (N2523, N2515, N2336, N318);
nor NOR3 (N2524, N2510, N2127, N1707);
endmodule