// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N306,N314,N300,N302,N317,N298,N315,N309,N308,N318;

and AND4 (N19, N12, N1, N11, N17);
not NOT1 (N20, N17);
nor NOR2 (N21, N5, N20);
buf BUF1 (N22, N12);
and AND4 (N23, N10, N3, N21, N3);
buf BUF1 (N24, N9);
nor NOR2 (N25, N14, N2);
and AND3 (N26, N3, N9, N11);
or OR4 (N27, N10, N17, N21, N25);
not NOT1 (N28, N17);
buf BUF1 (N29, N9);
and AND2 (N30, N22, N9);
and AND2 (N31, N14, N17);
xor XOR2 (N32, N31, N2);
not NOT1 (N33, N19);
and AND3 (N34, N5, N24, N6);
nor NOR4 (N35, N26, N4, N3, N6);
or OR3 (N36, N32, N21, N27);
or OR3 (N37, N3, N31, N9);
and AND2 (N38, N35, N34);
not NOT1 (N39, N5);
xor XOR2 (N40, N5, N34);
or OR4 (N41, N38, N38, N16, N17);
buf BUF1 (N42, N23);
and AND3 (N43, N40, N37, N38);
nand NAND4 (N44, N26, N22, N6, N1);
nor NOR4 (N45, N42, N28, N18, N17);
buf BUF1 (N46, N12);
xor XOR2 (N47, N43, N37);
nor NOR4 (N48, N29, N17, N16, N28);
nand NAND2 (N49, N48, N4);
or OR3 (N50, N39, N24, N36);
xor XOR2 (N51, N36, N43);
nand NAND3 (N52, N44, N6, N7);
buf BUF1 (N53, N51);
and AND2 (N54, N33, N24);
nand NAND2 (N55, N46, N11);
not NOT1 (N56, N50);
nor NOR4 (N57, N56, N34, N16, N31);
buf BUF1 (N58, N57);
nand NAND2 (N59, N52, N54);
not NOT1 (N60, N15);
nand NAND4 (N61, N47, N4, N6, N31);
buf BUF1 (N62, N58);
not NOT1 (N63, N55);
or OR4 (N64, N41, N9, N24, N51);
and AND3 (N65, N63, N53, N61);
nand NAND2 (N66, N34, N38);
and AND4 (N67, N45, N18, N34, N3);
nand NAND4 (N68, N44, N3, N66, N4);
buf BUF1 (N69, N19);
not NOT1 (N70, N59);
xor XOR2 (N71, N62, N43);
nor NOR2 (N72, N70, N25);
or OR4 (N73, N72, N68, N35, N28);
xor XOR2 (N74, N14, N25);
or OR4 (N75, N73, N71, N32, N53);
not NOT1 (N76, N40);
xor XOR2 (N77, N76, N19);
xor XOR2 (N78, N77, N42);
xor XOR2 (N79, N74, N49);
nand NAND3 (N80, N45, N66, N39);
buf BUF1 (N81, N79);
nor NOR2 (N82, N80, N35);
nor NOR3 (N83, N64, N17, N19);
not NOT1 (N84, N75);
nand NAND4 (N85, N67, N63, N70, N80);
nand NAND2 (N86, N65, N69);
nor NOR2 (N87, N2, N54);
buf BUF1 (N88, N86);
nor NOR4 (N89, N30, N77, N20, N27);
nand NAND2 (N90, N84, N45);
or OR4 (N91, N89, N15, N57, N29);
not NOT1 (N92, N91);
xor XOR2 (N93, N92, N58);
not NOT1 (N94, N88);
nor NOR4 (N95, N85, N76, N46, N13);
and AND2 (N96, N60, N6);
buf BUF1 (N97, N81);
and AND2 (N98, N95, N24);
nor NOR3 (N99, N94, N47, N75);
nand NAND2 (N100, N97, N88);
not NOT1 (N101, N87);
xor XOR2 (N102, N90, N43);
not NOT1 (N103, N98);
not NOT1 (N104, N102);
xor XOR2 (N105, N101, N17);
nor NOR3 (N106, N83, N27, N52);
xor XOR2 (N107, N78, N24);
xor XOR2 (N108, N99, N101);
or OR2 (N109, N103, N81);
nor NOR4 (N110, N96, N42, N55, N75);
nand NAND2 (N111, N108, N90);
or OR4 (N112, N110, N99, N82, N34);
or OR2 (N113, N96, N10);
or OR3 (N114, N107, N104, N21);
nor NOR4 (N115, N31, N20, N88, N31);
nand NAND4 (N116, N105, N90, N67, N83);
nor NOR4 (N117, N112, N47, N87, N33);
not NOT1 (N118, N115);
not NOT1 (N119, N111);
nand NAND3 (N120, N93, N33, N38);
not NOT1 (N121, N117);
and AND3 (N122, N121, N34, N56);
buf BUF1 (N123, N109);
or OR4 (N124, N122, N121, N86, N65);
xor XOR2 (N125, N116, N35);
or OR4 (N126, N120, N111, N1, N35);
and AND4 (N127, N106, N99, N64, N13);
xor XOR2 (N128, N127, N90);
buf BUF1 (N129, N100);
and AND2 (N130, N129, N88);
nor NOR4 (N131, N123, N19, N19, N69);
nor NOR2 (N132, N125, N16);
buf BUF1 (N133, N113);
nor NOR4 (N134, N133, N90, N4, N57);
buf BUF1 (N135, N119);
not NOT1 (N136, N131);
or OR3 (N137, N136, N62, N35);
and AND4 (N138, N135, N110, N69, N23);
buf BUF1 (N139, N118);
nand NAND2 (N140, N134, N132);
buf BUF1 (N141, N108);
not NOT1 (N142, N130);
not NOT1 (N143, N126);
or OR2 (N144, N142, N73);
not NOT1 (N145, N144);
and AND3 (N146, N128, N27, N60);
buf BUF1 (N147, N124);
buf BUF1 (N148, N143);
nor NOR4 (N149, N139, N115, N3, N77);
xor XOR2 (N150, N140, N28);
or OR2 (N151, N141, N49);
or OR2 (N152, N146, N138);
or OR4 (N153, N68, N89, N148, N127);
or OR3 (N154, N27, N32, N146);
buf BUF1 (N155, N154);
nand NAND3 (N156, N152, N5, N105);
not NOT1 (N157, N114);
buf BUF1 (N158, N147);
or OR4 (N159, N137, N58, N88, N11);
or OR4 (N160, N155, N98, N80, N120);
nor NOR3 (N161, N158, N68, N47);
nand NAND2 (N162, N151, N77);
or OR2 (N163, N145, N158);
nor NOR2 (N164, N153, N128);
xor XOR2 (N165, N156, N17);
nor NOR3 (N166, N160, N20, N47);
xor XOR2 (N167, N165, N58);
nor NOR2 (N168, N164, N161);
or OR2 (N169, N18, N11);
buf BUF1 (N170, N168);
and AND4 (N171, N149, N52, N104, N90);
and AND2 (N172, N169, N70);
and AND4 (N173, N150, N76, N30, N130);
buf BUF1 (N174, N167);
or OR4 (N175, N173, N9, N38, N57);
nor NOR4 (N176, N174, N145, N135, N30);
and AND3 (N177, N170, N115, N124);
nand NAND2 (N178, N162, N118);
nor NOR4 (N179, N177, N42, N76, N23);
and AND3 (N180, N172, N93, N127);
not NOT1 (N181, N175);
buf BUF1 (N182, N179);
and AND2 (N183, N159, N149);
not NOT1 (N184, N182);
not NOT1 (N185, N157);
nand NAND4 (N186, N181, N48, N67, N56);
buf BUF1 (N187, N183);
or OR4 (N188, N186, N175, N48, N57);
and AND4 (N189, N166, N57, N134, N7);
nand NAND2 (N190, N180, N107);
or OR4 (N191, N189, N69, N1, N100);
buf BUF1 (N192, N163);
and AND3 (N193, N171, N139, N66);
buf BUF1 (N194, N176);
xor XOR2 (N195, N192, N3);
xor XOR2 (N196, N190, N13);
buf BUF1 (N197, N191);
and AND2 (N198, N187, N162);
nor NOR2 (N199, N193, N43);
nand NAND4 (N200, N198, N199, N161, N12);
or OR2 (N201, N101, N134);
xor XOR2 (N202, N197, N132);
and AND4 (N203, N178, N161, N126, N11);
and AND3 (N204, N196, N191, N169);
not NOT1 (N205, N200);
nor NOR2 (N206, N184, N33);
and AND4 (N207, N202, N76, N70, N75);
and AND3 (N208, N195, N187, N139);
nor NOR2 (N209, N201, N29);
buf BUF1 (N210, N209);
nand NAND3 (N211, N206, N66, N90);
xor XOR2 (N212, N211, N97);
or OR2 (N213, N212, N28);
not NOT1 (N214, N213);
buf BUF1 (N215, N207);
buf BUF1 (N216, N204);
buf BUF1 (N217, N188);
not NOT1 (N218, N203);
xor XOR2 (N219, N215, N169);
buf BUF1 (N220, N216);
buf BUF1 (N221, N210);
not NOT1 (N222, N221);
nor NOR2 (N223, N214, N85);
buf BUF1 (N224, N205);
buf BUF1 (N225, N185);
buf BUF1 (N226, N217);
not NOT1 (N227, N208);
or OR4 (N228, N225, N108, N76, N88);
not NOT1 (N229, N224);
nand NAND4 (N230, N229, N67, N111, N45);
nand NAND2 (N231, N228, N205);
buf BUF1 (N232, N223);
not NOT1 (N233, N226);
xor XOR2 (N234, N233, N156);
nand NAND3 (N235, N227, N104, N165);
nor NOR4 (N236, N218, N232, N197, N161);
buf BUF1 (N237, N196);
buf BUF1 (N238, N235);
buf BUF1 (N239, N222);
not NOT1 (N240, N220);
buf BUF1 (N241, N237);
nor NOR2 (N242, N219, N120);
nor NOR3 (N243, N239, N187, N119);
buf BUF1 (N244, N194);
nand NAND4 (N245, N230, N97, N14, N11);
and AND2 (N246, N231, N224);
buf BUF1 (N247, N245);
buf BUF1 (N248, N246);
buf BUF1 (N249, N243);
buf BUF1 (N250, N247);
nor NOR3 (N251, N238, N207, N22);
buf BUF1 (N252, N236);
and AND3 (N253, N250, N126, N14);
buf BUF1 (N254, N244);
nor NOR4 (N255, N251, N39, N195, N190);
and AND3 (N256, N242, N20, N174);
and AND2 (N257, N234, N6);
or OR3 (N258, N252, N236, N181);
or OR4 (N259, N258, N94, N102, N151);
buf BUF1 (N260, N259);
not NOT1 (N261, N249);
nand NAND2 (N262, N241, N233);
buf BUF1 (N263, N257);
not NOT1 (N264, N260);
or OR3 (N265, N263, N131, N93);
buf BUF1 (N266, N254);
not NOT1 (N267, N261);
xor XOR2 (N268, N265, N142);
or OR4 (N269, N268, N245, N209, N41);
xor XOR2 (N270, N256, N148);
buf BUF1 (N271, N269);
not NOT1 (N272, N240);
xor XOR2 (N273, N255, N231);
and AND2 (N274, N266, N8);
not NOT1 (N275, N272);
xor XOR2 (N276, N273, N221);
xor XOR2 (N277, N264, N54);
xor XOR2 (N278, N270, N156);
not NOT1 (N279, N275);
buf BUF1 (N280, N253);
xor XOR2 (N281, N277, N96);
nand NAND2 (N282, N278, N97);
not NOT1 (N283, N262);
not NOT1 (N284, N282);
and AND2 (N285, N280, N135);
nor NOR2 (N286, N285, N233);
or OR4 (N287, N284, N132, N59, N163);
not NOT1 (N288, N274);
nor NOR4 (N289, N283, N4, N187, N43);
buf BUF1 (N290, N267);
nand NAND3 (N291, N276, N251, N100);
xor XOR2 (N292, N291, N254);
nand NAND4 (N293, N286, N85, N286, N248);
nand NAND2 (N294, N214, N46);
buf BUF1 (N295, N289);
xor XOR2 (N296, N292, N264);
not NOT1 (N297, N288);
not NOT1 (N298, N281);
and AND4 (N299, N297, N34, N106, N284);
not NOT1 (N300, N296);
xor XOR2 (N301, N271, N100);
nand NAND4 (N302, N299, N283, N89, N211);
and AND4 (N303, N279, N186, N132, N264);
buf BUF1 (N304, N295);
nand NAND4 (N305, N287, N134, N182, N221);
or OR3 (N306, N305, N136, N85);
nand NAND3 (N307, N290, N184, N159);
nor NOR4 (N308, N304, N232, N289, N125);
nor NOR3 (N309, N303, N39, N213);
or OR4 (N310, N293, N197, N87, N95);
and AND4 (N311, N294, N105, N27, N224);
buf BUF1 (N312, N307);
xor XOR2 (N313, N301, N167);
nand NAND4 (N314, N312, N70, N3, N110);
or OR4 (N315, N313, N143, N57, N105);
or OR3 (N316, N311, N29, N226);
xor XOR2 (N317, N316, N259);
nand NAND4 (N318, N310, N111, N126, N245);
endmodule