// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N519,N521,N522,N516,N520,N517,N515,N523,N507,N524;

or OR2 (N25, N5, N14);
nand NAND3 (N26, N13, N20, N7);
xor XOR2 (N27, N16, N2);
or OR3 (N28, N6, N14, N1);
nand NAND2 (N29, N9, N4);
nand NAND3 (N30, N19, N5, N22);
or OR4 (N31, N2, N28, N10, N23);
buf BUF1 (N32, N21);
nor NOR3 (N33, N32, N31, N14);
nor NOR2 (N34, N13, N32);
and AND3 (N35, N27, N33, N14);
and AND2 (N36, N20, N24);
or OR2 (N37, N11, N10);
and AND4 (N38, N8, N28, N3, N12);
and AND2 (N39, N15, N4);
buf BUF1 (N40, N35);
nor NOR3 (N41, N39, N36, N2);
not NOT1 (N42, N7);
or OR4 (N43, N30, N37, N11, N22);
xor XOR2 (N44, N37, N11);
not NOT1 (N45, N44);
and AND3 (N46, N34, N15, N25);
xor XOR2 (N47, N23, N41);
and AND4 (N48, N45, N32, N25, N43);
nand NAND2 (N49, N15, N15);
nor NOR4 (N50, N38, N44, N28, N35);
and AND3 (N51, N6, N39, N31);
nand NAND4 (N52, N50, N33, N3, N51);
buf BUF1 (N53, N20);
or OR4 (N54, N29, N44, N37, N10);
not NOT1 (N55, N54);
nand NAND4 (N56, N47, N35, N1, N4);
or OR4 (N57, N26, N30, N40, N4);
or OR2 (N58, N4, N36);
not NOT1 (N59, N56);
not NOT1 (N60, N42);
xor XOR2 (N61, N48, N49);
and AND3 (N62, N55, N27, N59);
not NOT1 (N63, N19);
xor XOR2 (N64, N60, N18);
xor XOR2 (N65, N19, N11);
and AND3 (N66, N46, N9, N50);
buf BUF1 (N67, N58);
xor XOR2 (N68, N53, N63);
and AND2 (N69, N26, N65);
and AND3 (N70, N49, N12, N22);
not NOT1 (N71, N52);
nand NAND3 (N72, N71, N69, N33);
and AND4 (N73, N38, N21, N67, N6);
buf BUF1 (N74, N34);
nor NOR3 (N75, N70, N35, N22);
nor NOR3 (N76, N62, N41, N71);
nor NOR2 (N77, N57, N23);
not NOT1 (N78, N61);
or OR2 (N79, N72, N61);
or OR2 (N80, N64, N62);
not NOT1 (N81, N66);
and AND3 (N82, N78, N64, N73);
xor XOR2 (N83, N29, N35);
buf BUF1 (N84, N82);
buf BUF1 (N85, N79);
not NOT1 (N86, N75);
buf BUF1 (N87, N84);
or OR4 (N88, N86, N75, N64, N31);
xor XOR2 (N89, N74, N81);
buf BUF1 (N90, N27);
nor NOR2 (N91, N76, N87);
buf BUF1 (N92, N13);
nand NAND2 (N93, N83, N77);
nand NAND2 (N94, N31, N43);
buf BUF1 (N95, N90);
nor NOR2 (N96, N95, N89);
nor NOR3 (N97, N37, N75, N46);
nand NAND3 (N98, N92, N76, N19);
or OR2 (N99, N97, N90);
or OR2 (N100, N93, N44);
not NOT1 (N101, N96);
buf BUF1 (N102, N100);
nand NAND4 (N103, N80, N53, N24, N41);
and AND4 (N104, N94, N67, N77, N64);
or OR2 (N105, N99, N23);
nand NAND2 (N106, N105, N54);
xor XOR2 (N107, N85, N13);
not NOT1 (N108, N103);
nand NAND4 (N109, N108, N60, N4, N62);
xor XOR2 (N110, N91, N58);
not NOT1 (N111, N110);
xor XOR2 (N112, N107, N63);
or OR3 (N113, N111, N112, N61);
or OR3 (N114, N112, N46, N49);
buf BUF1 (N115, N88);
nand NAND4 (N116, N109, N58, N48, N40);
and AND3 (N117, N104, N48, N49);
buf BUF1 (N118, N101);
nor NOR3 (N119, N115, N46, N41);
xor XOR2 (N120, N116, N109);
nand NAND2 (N121, N68, N36);
nand NAND3 (N122, N102, N30, N43);
xor XOR2 (N123, N114, N95);
xor XOR2 (N124, N123, N56);
nor NOR2 (N125, N121, N73);
and AND4 (N126, N117, N54, N119, N7);
or OR4 (N127, N111, N44, N25, N4);
not NOT1 (N128, N106);
nor NOR3 (N129, N118, N62, N47);
not NOT1 (N130, N126);
nor NOR2 (N131, N122, N81);
xor XOR2 (N132, N120, N86);
buf BUF1 (N133, N132);
and AND3 (N134, N127, N13, N77);
nor NOR4 (N135, N125, N32, N115, N2);
or OR4 (N136, N134, N32, N32, N25);
or OR4 (N137, N124, N87, N75, N53);
not NOT1 (N138, N136);
xor XOR2 (N139, N98, N38);
buf BUF1 (N140, N129);
or OR2 (N141, N131, N89);
not NOT1 (N142, N141);
nor NOR2 (N143, N135, N34);
and AND2 (N144, N143, N82);
or OR3 (N145, N113, N105, N34);
or OR4 (N146, N140, N62, N67, N107);
or OR4 (N147, N128, N110, N140, N84);
nand NAND3 (N148, N133, N78, N41);
nor NOR3 (N149, N139, N101, N108);
buf BUF1 (N150, N138);
or OR4 (N151, N146, N133, N125, N62);
not NOT1 (N152, N145);
or OR3 (N153, N144, N130, N20);
not NOT1 (N154, N121);
buf BUF1 (N155, N142);
nor NOR4 (N156, N152, N145, N123, N58);
nor NOR3 (N157, N154, N148, N83);
buf BUF1 (N158, N67);
and AND4 (N159, N151, N104, N35, N136);
not NOT1 (N160, N158);
buf BUF1 (N161, N149);
or OR3 (N162, N161, N65, N156);
or OR4 (N163, N157, N81, N107, N59);
buf BUF1 (N164, N123);
xor XOR2 (N165, N137, N34);
nand NAND3 (N166, N159, N127, N112);
not NOT1 (N167, N155);
buf BUF1 (N168, N163);
not NOT1 (N169, N160);
or OR2 (N170, N164, N53);
nor NOR3 (N171, N165, N132, N144);
xor XOR2 (N172, N162, N126);
not NOT1 (N173, N170);
nor NOR4 (N174, N150, N42, N137, N127);
and AND4 (N175, N167, N5, N144, N76);
nand NAND4 (N176, N147, N97, N23, N154);
and AND4 (N177, N173, N59, N143, N144);
and AND4 (N178, N175, N115, N52, N147);
buf BUF1 (N179, N168);
not NOT1 (N180, N178);
buf BUF1 (N181, N171);
xor XOR2 (N182, N180, N176);
nand NAND3 (N183, N24, N46, N171);
nand NAND2 (N184, N153, N111);
and AND4 (N185, N183, N95, N70, N2);
nand NAND2 (N186, N169, N138);
and AND2 (N187, N177, N131);
xor XOR2 (N188, N181, N18);
or OR2 (N189, N188, N100);
buf BUF1 (N190, N184);
and AND2 (N191, N186, N97);
xor XOR2 (N192, N182, N167);
or OR3 (N193, N174, N41, N47);
not NOT1 (N194, N172);
buf BUF1 (N195, N179);
and AND4 (N196, N187, N99, N45, N32);
nor NOR4 (N197, N190, N140, N46, N145);
not NOT1 (N198, N192);
and AND3 (N199, N189, N174, N14);
xor XOR2 (N200, N199, N5);
or OR2 (N201, N198, N139);
nand NAND3 (N202, N197, N94, N115);
nand NAND2 (N203, N185, N125);
xor XOR2 (N204, N196, N201);
or OR2 (N205, N200, N101);
nand NAND2 (N206, N141, N97);
or OR4 (N207, N195, N66, N83, N7);
and AND3 (N208, N193, N156, N116);
buf BUF1 (N209, N206);
buf BUF1 (N210, N208);
nor NOR2 (N211, N205, N81);
xor XOR2 (N212, N211, N179);
buf BUF1 (N213, N210);
or OR4 (N214, N204, N71, N13, N152);
buf BUF1 (N215, N212);
buf BUF1 (N216, N207);
and AND4 (N217, N203, N19, N62, N6);
or OR4 (N218, N194, N164, N99, N176);
buf BUF1 (N219, N202);
xor XOR2 (N220, N218, N210);
and AND2 (N221, N215, N99);
not NOT1 (N222, N166);
nand NAND2 (N223, N221, N147);
nand NAND4 (N224, N209, N97, N85, N218);
buf BUF1 (N225, N214);
or OR4 (N226, N223, N35, N110, N40);
nand NAND2 (N227, N213, N63);
nand NAND3 (N228, N225, N180, N115);
xor XOR2 (N229, N227, N13);
or OR4 (N230, N224, N116, N224, N74);
nor NOR2 (N231, N219, N6);
nand NAND4 (N232, N217, N177, N45, N172);
buf BUF1 (N233, N226);
nor NOR3 (N234, N216, N169, N14);
buf BUF1 (N235, N222);
nand NAND2 (N236, N230, N84);
nor NOR3 (N237, N191, N133, N33);
not NOT1 (N238, N235);
or OR4 (N239, N234, N234, N137, N24);
nor NOR2 (N240, N220, N39);
or OR2 (N241, N229, N184);
or OR4 (N242, N236, N120, N58, N70);
xor XOR2 (N243, N239, N201);
xor XOR2 (N244, N243, N17);
not NOT1 (N245, N240);
and AND2 (N246, N233, N138);
nand NAND2 (N247, N244, N222);
nand NAND4 (N248, N246, N62, N178, N185);
and AND2 (N249, N231, N174);
xor XOR2 (N250, N237, N179);
nand NAND3 (N251, N241, N87, N166);
nor NOR4 (N252, N228, N214, N193, N82);
not NOT1 (N253, N247);
nor NOR3 (N254, N253, N1, N124);
xor XOR2 (N255, N245, N79);
xor XOR2 (N256, N248, N175);
nand NAND2 (N257, N251, N5);
not NOT1 (N258, N250);
not NOT1 (N259, N254);
and AND3 (N260, N257, N161, N58);
buf BUF1 (N261, N258);
xor XOR2 (N262, N259, N188);
xor XOR2 (N263, N260, N75);
not NOT1 (N264, N256);
nand NAND4 (N265, N263, N26, N2, N242);
nor NOR3 (N266, N243, N183, N94);
not NOT1 (N267, N232);
nand NAND3 (N268, N238, N62, N43);
nand NAND2 (N269, N262, N256);
nor NOR4 (N270, N265, N245, N228, N120);
xor XOR2 (N271, N249, N253);
nand NAND4 (N272, N267, N108, N231, N33);
or OR3 (N273, N261, N71, N222);
not NOT1 (N274, N268);
and AND3 (N275, N274, N157, N225);
nand NAND4 (N276, N269, N109, N81, N60);
not NOT1 (N277, N266);
buf BUF1 (N278, N272);
nor NOR2 (N279, N271, N184);
or OR2 (N280, N252, N109);
not NOT1 (N281, N270);
nand NAND4 (N282, N277, N265, N86, N58);
or OR2 (N283, N273, N92);
buf BUF1 (N284, N283);
and AND3 (N285, N281, N167, N21);
not NOT1 (N286, N264);
nand NAND3 (N287, N280, N136, N229);
nor NOR4 (N288, N286, N224, N164, N127);
xor XOR2 (N289, N284, N95);
nand NAND3 (N290, N275, N135, N49);
nand NAND4 (N291, N285, N80, N102, N95);
xor XOR2 (N292, N289, N240);
xor XOR2 (N293, N255, N144);
nand NAND4 (N294, N291, N203, N257, N243);
or OR3 (N295, N292, N212, N98);
nor NOR2 (N296, N278, N253);
nand NAND2 (N297, N290, N109);
xor XOR2 (N298, N279, N210);
nand NAND2 (N299, N297, N295);
not NOT1 (N300, N255);
xor XOR2 (N301, N298, N100);
buf BUF1 (N302, N276);
and AND4 (N303, N287, N61, N35, N44);
xor XOR2 (N304, N303, N60);
nand NAND2 (N305, N304, N87);
nor NOR4 (N306, N293, N9, N21, N26);
nor NOR2 (N307, N306, N300);
nor NOR4 (N308, N61, N24, N139, N272);
buf BUF1 (N309, N305);
nand NAND3 (N310, N301, N1, N229);
buf BUF1 (N311, N308);
nor NOR4 (N312, N296, N257, N192, N125);
not NOT1 (N313, N307);
xor XOR2 (N314, N288, N50);
not NOT1 (N315, N311);
or OR4 (N316, N309, N28, N24, N217);
not NOT1 (N317, N312);
not NOT1 (N318, N314);
and AND2 (N319, N313, N67);
xor XOR2 (N320, N317, N224);
not NOT1 (N321, N318);
nor NOR3 (N322, N294, N120, N138);
or OR4 (N323, N310, N210, N116, N152);
xor XOR2 (N324, N302, N111);
xor XOR2 (N325, N323, N52);
and AND3 (N326, N320, N47, N101);
or OR2 (N327, N326, N34);
nor NOR4 (N328, N322, N179, N218, N84);
and AND2 (N329, N325, N88);
and AND4 (N330, N316, N275, N112, N246);
buf BUF1 (N331, N319);
buf BUF1 (N332, N315);
and AND4 (N333, N331, N186, N266, N121);
and AND4 (N334, N330, N187, N125, N175);
not NOT1 (N335, N324);
not NOT1 (N336, N321);
buf BUF1 (N337, N332);
xor XOR2 (N338, N299, N327);
buf BUF1 (N339, N134);
not NOT1 (N340, N338);
nor NOR4 (N341, N340, N289, N57, N260);
nor NOR2 (N342, N334, N141);
not NOT1 (N343, N333);
xor XOR2 (N344, N329, N50);
nor NOR3 (N345, N336, N268, N50);
nor NOR2 (N346, N328, N309);
or OR2 (N347, N343, N149);
nor NOR2 (N348, N341, N94);
or OR2 (N349, N282, N168);
and AND2 (N350, N346, N78);
nand NAND4 (N351, N349, N182, N29, N165);
xor XOR2 (N352, N350, N1);
and AND2 (N353, N351, N86);
xor XOR2 (N354, N337, N272);
xor XOR2 (N355, N348, N339);
nand NAND4 (N356, N159, N60, N5, N120);
and AND3 (N357, N354, N247, N116);
or OR2 (N358, N335, N130);
nor NOR3 (N359, N353, N144, N123);
nor NOR3 (N360, N359, N25, N22);
xor XOR2 (N361, N344, N301);
nor NOR4 (N362, N355, N257, N294, N23);
not NOT1 (N363, N345);
and AND2 (N364, N352, N239);
buf BUF1 (N365, N358);
or OR2 (N366, N365, N4);
nor NOR4 (N367, N361, N57, N66, N319);
buf BUF1 (N368, N362);
buf BUF1 (N369, N357);
or OR3 (N370, N369, N309, N211);
buf BUF1 (N371, N347);
buf BUF1 (N372, N370);
buf BUF1 (N373, N371);
nand NAND2 (N374, N368, N180);
nor NOR2 (N375, N342, N143);
not NOT1 (N376, N360);
xor XOR2 (N377, N367, N231);
not NOT1 (N378, N374);
and AND3 (N379, N373, N8, N179);
buf BUF1 (N380, N377);
and AND2 (N381, N372, N46);
nor NOR3 (N382, N380, N197, N77);
and AND2 (N383, N375, N232);
nand NAND3 (N384, N383, N306, N377);
nand NAND2 (N385, N379, N244);
xor XOR2 (N386, N382, N82);
not NOT1 (N387, N356);
or OR3 (N388, N385, N298, N275);
xor XOR2 (N389, N388, N364);
nor NOR3 (N390, N134, N211, N160);
and AND4 (N391, N387, N263, N153, N109);
nor NOR4 (N392, N381, N335, N91, N140);
buf BUF1 (N393, N378);
not NOT1 (N394, N376);
buf BUF1 (N395, N394);
or OR2 (N396, N393, N315);
nand NAND3 (N397, N392, N195, N256);
or OR4 (N398, N366, N137, N226, N282);
and AND2 (N399, N397, N231);
nor NOR2 (N400, N398, N114);
and AND2 (N401, N400, N66);
xor XOR2 (N402, N386, N157);
buf BUF1 (N403, N395);
nor NOR2 (N404, N403, N228);
nor NOR4 (N405, N391, N154, N68, N202);
xor XOR2 (N406, N402, N197);
nor NOR3 (N407, N389, N392, N306);
or OR4 (N408, N363, N233, N111, N88);
not NOT1 (N409, N396);
buf BUF1 (N410, N401);
buf BUF1 (N411, N406);
buf BUF1 (N412, N384);
and AND3 (N413, N409, N272, N176);
not NOT1 (N414, N390);
nand NAND3 (N415, N407, N368, N8);
nor NOR2 (N416, N405, N281);
xor XOR2 (N417, N413, N136);
nor NOR4 (N418, N414, N169, N185, N100);
nand NAND4 (N419, N410, N412, N91, N246);
xor XOR2 (N420, N16, N151);
nand NAND3 (N421, N415, N301, N190);
and AND4 (N422, N418, N2, N382, N287);
nor NOR4 (N423, N408, N327, N357, N260);
not NOT1 (N424, N420);
or OR4 (N425, N421, N223, N345, N329);
nor NOR4 (N426, N404, N338, N133, N414);
not NOT1 (N427, N423);
buf BUF1 (N428, N427);
and AND4 (N429, N416, N27, N411, N354);
buf BUF1 (N430, N70);
buf BUF1 (N431, N399);
or OR4 (N432, N425, N381, N167, N81);
nand NAND4 (N433, N431, N206, N209, N146);
or OR2 (N434, N417, N384);
nor NOR3 (N435, N419, N374, N254);
nand NAND4 (N436, N426, N50, N192, N242);
nand NAND2 (N437, N433, N160);
xor XOR2 (N438, N434, N338);
xor XOR2 (N439, N436, N289);
buf BUF1 (N440, N438);
nand NAND2 (N441, N432, N166);
not NOT1 (N442, N428);
and AND2 (N443, N429, N328);
nor NOR3 (N444, N442, N419, N79);
buf BUF1 (N445, N439);
not NOT1 (N446, N422);
not NOT1 (N447, N440);
nor NOR3 (N448, N437, N262, N59);
or OR3 (N449, N443, N333, N233);
nand NAND4 (N450, N444, N300, N78, N7);
or OR4 (N451, N435, N95, N67, N396);
nor NOR3 (N452, N445, N324, N165);
buf BUF1 (N453, N449);
buf BUF1 (N454, N451);
not NOT1 (N455, N446);
not NOT1 (N456, N450);
nor NOR4 (N457, N447, N69, N264, N69);
buf BUF1 (N458, N456);
nand NAND2 (N459, N458, N386);
not NOT1 (N460, N454);
xor XOR2 (N461, N441, N275);
buf BUF1 (N462, N453);
buf BUF1 (N463, N459);
buf BUF1 (N464, N424);
or OR3 (N465, N461, N191, N387);
nor NOR2 (N466, N465, N105);
and AND4 (N467, N464, N259, N441, N188);
and AND2 (N468, N466, N212);
xor XOR2 (N469, N457, N353);
buf BUF1 (N470, N460);
nor NOR4 (N471, N463, N126, N110, N344);
nand NAND2 (N472, N470, N257);
nand NAND3 (N473, N455, N294, N182);
or OR4 (N474, N473, N339, N373, N40);
buf BUF1 (N475, N468);
buf BUF1 (N476, N467);
and AND3 (N477, N448, N110, N254);
not NOT1 (N478, N476);
or OR3 (N479, N477, N410, N65);
not NOT1 (N480, N474);
xor XOR2 (N481, N480, N457);
nor NOR4 (N482, N462, N163, N128, N201);
xor XOR2 (N483, N481, N39);
xor XOR2 (N484, N452, N190);
xor XOR2 (N485, N430, N401);
not NOT1 (N486, N475);
or OR2 (N487, N485, N59);
nor NOR2 (N488, N482, N189);
xor XOR2 (N489, N479, N399);
xor XOR2 (N490, N471, N358);
xor XOR2 (N491, N489, N208);
xor XOR2 (N492, N488, N330);
nor NOR3 (N493, N492, N320, N278);
xor XOR2 (N494, N491, N338);
buf BUF1 (N495, N486);
not NOT1 (N496, N478);
or OR4 (N497, N490, N264, N207, N177);
or OR3 (N498, N487, N26, N112);
or OR2 (N499, N472, N119);
or OR2 (N500, N498, N377);
or OR3 (N501, N499, N259, N57);
not NOT1 (N502, N497);
or OR4 (N503, N494, N169, N87, N211);
nor NOR2 (N504, N501, N316);
xor XOR2 (N505, N495, N492);
not NOT1 (N506, N496);
not NOT1 (N507, N502);
nand NAND2 (N508, N483, N301);
xor XOR2 (N509, N505, N167);
not NOT1 (N510, N469);
and AND2 (N511, N510, N488);
or OR2 (N512, N511, N394);
and AND2 (N513, N504, N134);
xor XOR2 (N514, N508, N16);
xor XOR2 (N515, N484, N209);
not NOT1 (N516, N514);
not NOT1 (N517, N509);
buf BUF1 (N518, N503);
not NOT1 (N519, N513);
xor XOR2 (N520, N506, N340);
not NOT1 (N521, N512);
buf BUF1 (N522, N500);
buf BUF1 (N523, N518);
and AND3 (N524, N493, N399, N51);
endmodule