// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16;

output N7993,N8003,N8008,N8015,N8014,N8011,N8005,N8013,N8009,N8016;

or OR4 (N17, N12, N8, N16, N2);
or OR4 (N18, N5, N11, N2, N14);
or OR2 (N19, N18, N6);
xor XOR2 (N20, N4, N10);
xor XOR2 (N21, N2, N20);
buf BUF1 (N22, N18);
xor XOR2 (N23, N15, N2);
buf BUF1 (N24, N7);
and AND2 (N25, N5, N16);
xor XOR2 (N26, N8, N4);
nor NOR4 (N27, N10, N6, N21, N3);
buf BUF1 (N28, N18);
and AND2 (N29, N10, N27);
or OR4 (N30, N10, N23, N25, N5);
or OR4 (N31, N24, N1, N4, N12);
or OR2 (N32, N24, N5);
nor NOR4 (N33, N26, N21, N20, N14);
or OR2 (N34, N5, N2);
or OR3 (N35, N28, N34, N22);
buf BUF1 (N36, N18);
or OR2 (N37, N23, N29);
nor NOR3 (N38, N5, N25, N26);
or OR4 (N39, N38, N27, N34, N10);
nor NOR3 (N40, N36, N27, N11);
not NOT1 (N41, N17);
nand NAND4 (N42, N32, N39, N16, N36);
nand NAND4 (N43, N15, N35, N39, N39);
xor XOR2 (N44, N33, N9);
or OR3 (N45, N18, N21, N8);
nand NAND3 (N46, N45, N10, N5);
nor NOR2 (N47, N41, N8);
and AND3 (N48, N40, N34, N3);
buf BUF1 (N49, N43);
nand NAND2 (N50, N48, N45);
xor XOR2 (N51, N31, N28);
not NOT1 (N52, N19);
and AND2 (N53, N47, N47);
nand NAND4 (N54, N42, N17, N33, N34);
or OR4 (N55, N46, N53, N10, N42);
not NOT1 (N56, N54);
and AND3 (N57, N19, N7, N40);
xor XOR2 (N58, N49, N38);
not NOT1 (N59, N50);
and AND3 (N60, N57, N2, N59);
and AND2 (N61, N17, N19);
xor XOR2 (N62, N51, N15);
or OR2 (N63, N37, N56);
or OR2 (N64, N53, N5);
or OR3 (N65, N62, N19, N25);
not NOT1 (N66, N60);
nor NOR4 (N67, N44, N51, N23, N40);
or OR4 (N68, N61, N13, N49, N2);
buf BUF1 (N69, N52);
not NOT1 (N70, N64);
or OR3 (N71, N70, N20, N9);
not NOT1 (N72, N58);
nand NAND3 (N73, N30, N49, N27);
xor XOR2 (N74, N71, N24);
not NOT1 (N75, N72);
nor NOR3 (N76, N66, N52, N32);
nor NOR2 (N77, N75, N36);
nand NAND2 (N78, N65, N32);
buf BUF1 (N79, N76);
nand NAND3 (N80, N68, N55, N41);
nand NAND4 (N81, N4, N47, N55, N80);
not NOT1 (N82, N30);
nand NAND4 (N83, N82, N54, N33, N48);
and AND4 (N84, N63, N19, N21, N50);
and AND3 (N85, N84, N30, N63);
nand NAND3 (N86, N79, N52, N61);
nor NOR2 (N87, N81, N9);
not NOT1 (N88, N87);
xor XOR2 (N89, N73, N46);
or OR4 (N90, N89, N50, N21, N50);
and AND2 (N91, N86, N66);
buf BUF1 (N92, N85);
not NOT1 (N93, N78);
and AND3 (N94, N90, N93, N39);
nand NAND2 (N95, N86, N44);
or OR4 (N96, N94, N94, N90, N17);
and AND3 (N97, N91, N9, N82);
buf BUF1 (N98, N97);
or OR2 (N99, N67, N17);
nor NOR2 (N100, N74, N70);
xor XOR2 (N101, N98, N68);
or OR3 (N102, N95, N58, N51);
buf BUF1 (N103, N77);
not NOT1 (N104, N96);
not NOT1 (N105, N69);
nand NAND3 (N106, N104, N1, N70);
buf BUF1 (N107, N105);
nand NAND3 (N108, N88, N54, N21);
and AND4 (N109, N101, N54, N81, N51);
nor NOR4 (N110, N99, N85, N52, N1);
buf BUF1 (N111, N109);
and AND3 (N112, N110, N74, N36);
and AND4 (N113, N108, N7, N17, N29);
nand NAND3 (N114, N83, N105, N81);
not NOT1 (N115, N111);
nand NAND2 (N116, N103, N66);
xor XOR2 (N117, N102, N5);
buf BUF1 (N118, N106);
nor NOR3 (N119, N114, N27, N32);
and AND2 (N120, N113, N28);
and AND3 (N121, N107, N79, N98);
nand NAND4 (N122, N121, N26, N77, N91);
nand NAND4 (N123, N117, N106, N98, N23);
buf BUF1 (N124, N92);
and AND2 (N125, N120, N79);
nor NOR4 (N126, N124, N16, N95, N24);
buf BUF1 (N127, N126);
xor XOR2 (N128, N119, N100);
not NOT1 (N129, N97);
xor XOR2 (N130, N118, N71);
not NOT1 (N131, N122);
xor XOR2 (N132, N112, N59);
xor XOR2 (N133, N130, N40);
not NOT1 (N134, N132);
not NOT1 (N135, N128);
and AND3 (N136, N115, N95, N64);
and AND4 (N137, N135, N123, N13, N65);
buf BUF1 (N138, N68);
not NOT1 (N139, N127);
buf BUF1 (N140, N139);
nor NOR4 (N141, N137, N7, N107, N62);
not NOT1 (N142, N138);
and AND3 (N143, N116, N101, N111);
nor NOR3 (N144, N141, N14, N107);
xor XOR2 (N145, N131, N36);
buf BUF1 (N146, N125);
nand NAND4 (N147, N145, N135, N37, N124);
nand NAND3 (N148, N140, N125, N113);
nor NOR4 (N149, N148, N97, N85, N18);
nand NAND2 (N150, N136, N82);
buf BUF1 (N151, N147);
buf BUF1 (N152, N143);
or OR3 (N153, N146, N32, N91);
or OR4 (N154, N151, N8, N114, N148);
xor XOR2 (N155, N129, N137);
buf BUF1 (N156, N155);
not NOT1 (N157, N150);
xor XOR2 (N158, N144, N74);
nand NAND4 (N159, N133, N102, N135, N114);
xor XOR2 (N160, N157, N95);
not NOT1 (N161, N152);
and AND4 (N162, N160, N63, N50, N140);
or OR3 (N163, N142, N6, N82);
not NOT1 (N164, N134);
nand NAND3 (N165, N154, N111, N141);
xor XOR2 (N166, N158, N83);
nor NOR4 (N167, N166, N50, N89, N75);
xor XOR2 (N168, N163, N119);
buf BUF1 (N169, N149);
nor NOR3 (N170, N153, N90, N46);
or OR4 (N171, N170, N149, N51, N19);
not NOT1 (N172, N167);
and AND2 (N173, N156, N13);
not NOT1 (N174, N161);
and AND2 (N175, N168, N142);
and AND4 (N176, N172, N115, N170, N89);
nand NAND3 (N177, N169, N48, N143);
nand NAND2 (N178, N177, N59);
nor NOR3 (N179, N178, N94, N31);
nand NAND4 (N180, N175, N68, N173, N155);
or OR3 (N181, N40, N25, N102);
nand NAND4 (N182, N181, N92, N48, N138);
buf BUF1 (N183, N159);
and AND4 (N184, N165, N28, N6, N49);
and AND3 (N185, N183, N182, N130);
nor NOR2 (N186, N88, N12);
buf BUF1 (N187, N180);
nand NAND4 (N188, N162, N91, N153, N32);
nor NOR4 (N189, N184, N25, N111, N182);
or OR2 (N190, N188, N61);
not NOT1 (N191, N186);
buf BUF1 (N192, N176);
or OR4 (N193, N171, N88, N110, N160);
or OR2 (N194, N174, N83);
xor XOR2 (N195, N187, N99);
and AND4 (N196, N179, N43, N74, N97);
or OR2 (N197, N196, N143);
buf BUF1 (N198, N164);
nand NAND3 (N199, N185, N195, N114);
or OR3 (N200, N75, N64, N21);
or OR3 (N201, N194, N92, N84);
nand NAND3 (N202, N200, N83, N62);
not NOT1 (N203, N192);
nand NAND2 (N204, N190, N20);
nand NAND3 (N205, N189, N24, N144);
xor XOR2 (N206, N191, N182);
xor XOR2 (N207, N204, N89);
buf BUF1 (N208, N197);
or OR2 (N209, N202, N33);
and AND2 (N210, N208, N90);
and AND3 (N211, N206, N47, N65);
or OR2 (N212, N199, N52);
nand NAND3 (N213, N209, N1, N63);
buf BUF1 (N214, N203);
nor NOR2 (N215, N207, N173);
not NOT1 (N216, N213);
and AND4 (N217, N215, N38, N186, N151);
xor XOR2 (N218, N216, N53);
not NOT1 (N219, N198);
nor NOR2 (N220, N214, N195);
or OR2 (N221, N220, N59);
buf BUF1 (N222, N201);
and AND2 (N223, N222, N82);
nand NAND2 (N224, N221, N39);
or OR2 (N225, N218, N216);
xor XOR2 (N226, N223, N32);
not NOT1 (N227, N226);
nor NOR4 (N228, N210, N95, N43, N67);
and AND2 (N229, N228, N153);
and AND4 (N230, N225, N110, N183, N75);
and AND4 (N231, N227, N25, N207, N140);
and AND4 (N232, N211, N59, N90, N31);
buf BUF1 (N233, N212);
and AND2 (N234, N229, N16);
nor NOR4 (N235, N230, N146, N49, N191);
nand NAND2 (N236, N235, N208);
nor NOR3 (N237, N233, N197, N73);
and AND4 (N238, N237, N124, N170, N122);
nor NOR3 (N239, N217, N68, N192);
or OR4 (N240, N232, N64, N18, N50);
not NOT1 (N241, N193);
xor XOR2 (N242, N231, N63);
nand NAND2 (N243, N224, N218);
not NOT1 (N244, N238);
nor NOR2 (N245, N240, N213);
and AND2 (N246, N244, N145);
or OR3 (N247, N241, N162, N111);
nor NOR2 (N248, N234, N164);
not NOT1 (N249, N243);
buf BUF1 (N250, N249);
not NOT1 (N251, N250);
nand NAND3 (N252, N236, N207, N57);
nand NAND4 (N253, N252, N184, N227, N92);
nor NOR4 (N254, N246, N81, N158, N242);
buf BUF1 (N255, N158);
and AND4 (N256, N247, N59, N86, N227);
nor NOR3 (N257, N205, N249, N179);
nor NOR3 (N258, N219, N216, N120);
nor NOR3 (N259, N251, N178, N67);
not NOT1 (N260, N258);
not NOT1 (N261, N253);
nor NOR3 (N262, N260, N228, N235);
xor XOR2 (N263, N256, N95);
nor NOR4 (N264, N254, N61, N178, N88);
nand NAND3 (N265, N264, N126, N199);
not NOT1 (N266, N261);
xor XOR2 (N267, N255, N38);
and AND4 (N268, N262, N135, N157, N132);
nand NAND3 (N269, N268, N143, N124);
nor NOR3 (N270, N257, N65, N138);
nand NAND2 (N271, N263, N2);
or OR3 (N272, N267, N207, N13);
or OR2 (N273, N271, N14);
buf BUF1 (N274, N265);
xor XOR2 (N275, N259, N125);
nor NOR4 (N276, N245, N225, N211, N1);
nand NAND2 (N277, N266, N84);
nand NAND2 (N278, N239, N124);
and AND3 (N279, N275, N118, N209);
nand NAND3 (N280, N270, N217, N12);
or OR4 (N281, N278, N202, N136, N51);
nand NAND2 (N282, N281, N166);
and AND2 (N283, N248, N119);
and AND4 (N284, N273, N26, N172, N173);
nor NOR3 (N285, N283, N95, N180);
nand NAND2 (N286, N279, N88);
or OR4 (N287, N282, N14, N59, N256);
not NOT1 (N288, N276);
buf BUF1 (N289, N286);
xor XOR2 (N290, N288, N34);
buf BUF1 (N291, N269);
and AND2 (N292, N284, N126);
nor NOR4 (N293, N291, N161, N145, N55);
and AND2 (N294, N272, N63);
buf BUF1 (N295, N280);
or OR3 (N296, N295, N104, N171);
and AND2 (N297, N277, N44);
not NOT1 (N298, N296);
or OR3 (N299, N287, N66, N286);
buf BUF1 (N300, N292);
nor NOR4 (N301, N289, N222, N173, N1);
not NOT1 (N302, N293);
buf BUF1 (N303, N285);
not NOT1 (N304, N299);
nand NAND2 (N305, N294, N293);
buf BUF1 (N306, N290);
and AND4 (N307, N300, N194, N24, N151);
xor XOR2 (N308, N274, N84);
nor NOR4 (N309, N304, N115, N9, N263);
or OR4 (N310, N301, N106, N2, N76);
xor XOR2 (N311, N303, N172);
or OR4 (N312, N307, N180, N102, N190);
or OR2 (N313, N297, N192);
and AND4 (N314, N310, N14, N137, N94);
nand NAND2 (N315, N313, N247);
buf BUF1 (N316, N305);
not NOT1 (N317, N312);
not NOT1 (N318, N298);
nor NOR2 (N319, N302, N44);
buf BUF1 (N320, N309);
or OR2 (N321, N306, N295);
nand NAND2 (N322, N315, N14);
nor NOR2 (N323, N318, N165);
and AND4 (N324, N321, N216, N166, N262);
not NOT1 (N325, N319);
nand NAND3 (N326, N325, N245, N241);
nand NAND2 (N327, N317, N300);
buf BUF1 (N328, N324);
not NOT1 (N329, N327);
buf BUF1 (N330, N323);
nand NAND3 (N331, N314, N110, N216);
or OR4 (N332, N328, N78, N80, N109);
and AND3 (N333, N331, N2, N171);
nor NOR4 (N334, N326, N26, N147, N152);
or OR3 (N335, N320, N107, N232);
not NOT1 (N336, N330);
or OR3 (N337, N322, N323, N170);
buf BUF1 (N338, N329);
buf BUF1 (N339, N335);
and AND2 (N340, N339, N36);
nand NAND4 (N341, N338, N103, N285, N3);
or OR4 (N342, N332, N214, N108, N258);
nand NAND2 (N343, N337, N178);
buf BUF1 (N344, N343);
or OR2 (N345, N344, N13);
nand NAND4 (N346, N311, N5, N343, N42);
and AND3 (N347, N342, N117, N189);
nor NOR4 (N348, N340, N32, N215, N255);
buf BUF1 (N349, N308);
not NOT1 (N350, N348);
and AND3 (N351, N346, N315, N163);
not NOT1 (N352, N341);
not NOT1 (N353, N333);
not NOT1 (N354, N347);
or OR2 (N355, N350, N23);
or OR3 (N356, N345, N193, N316);
buf BUF1 (N357, N32);
not NOT1 (N358, N356);
or OR2 (N359, N353, N307);
or OR2 (N360, N352, N77);
nor NOR2 (N361, N355, N339);
and AND4 (N362, N359, N245, N297, N60);
buf BUF1 (N363, N360);
xor XOR2 (N364, N334, N83);
or OR4 (N365, N364, N306, N107, N194);
nand NAND4 (N366, N362, N114, N23, N3);
not NOT1 (N367, N361);
and AND4 (N368, N366, N78, N92, N33);
xor XOR2 (N369, N368, N6);
and AND2 (N370, N354, N239);
buf BUF1 (N371, N336);
xor XOR2 (N372, N363, N105);
or OR3 (N373, N371, N79, N242);
nor NOR2 (N374, N369, N92);
not NOT1 (N375, N370);
buf BUF1 (N376, N367);
or OR2 (N377, N374, N235);
and AND4 (N378, N377, N137, N144, N181);
or OR2 (N379, N373, N146);
and AND2 (N380, N349, N60);
nor NOR3 (N381, N375, N44, N207);
buf BUF1 (N382, N365);
nand NAND2 (N383, N351, N147);
not NOT1 (N384, N378);
xor XOR2 (N385, N384, N183);
not NOT1 (N386, N379);
nor NOR4 (N387, N358, N306, N257, N130);
nand NAND2 (N388, N357, N145);
xor XOR2 (N389, N381, N7);
nand NAND2 (N390, N382, N19);
xor XOR2 (N391, N376, N268);
or OR3 (N392, N391, N274, N196);
not NOT1 (N393, N387);
or OR3 (N394, N393, N145, N258);
buf BUF1 (N395, N380);
and AND3 (N396, N388, N202, N346);
and AND2 (N397, N385, N77);
xor XOR2 (N398, N386, N305);
and AND2 (N399, N389, N1);
and AND3 (N400, N395, N347, N62);
xor XOR2 (N401, N396, N16);
buf BUF1 (N402, N398);
xor XOR2 (N403, N400, N41);
buf BUF1 (N404, N392);
nand NAND2 (N405, N390, N51);
xor XOR2 (N406, N404, N289);
nor NOR3 (N407, N402, N264, N308);
not NOT1 (N408, N394);
xor XOR2 (N409, N397, N16);
not NOT1 (N410, N383);
nor NOR4 (N411, N406, N286, N28, N130);
and AND2 (N412, N405, N277);
and AND4 (N413, N409, N370, N126, N142);
buf BUF1 (N414, N413);
nor NOR3 (N415, N372, N394, N357);
or OR4 (N416, N399, N78, N227, N160);
not NOT1 (N417, N415);
or OR4 (N418, N401, N227, N232, N168);
nor NOR4 (N419, N418, N57, N107, N113);
and AND3 (N420, N414, N200, N99);
buf BUF1 (N421, N417);
xor XOR2 (N422, N419, N83);
nand NAND4 (N423, N403, N246, N183, N103);
and AND4 (N424, N412, N260, N212, N259);
nor NOR4 (N425, N420, N251, N159, N239);
buf BUF1 (N426, N424);
nand NAND4 (N427, N423, N199, N222, N209);
or OR3 (N428, N425, N102, N248);
or OR2 (N429, N416, N217);
buf BUF1 (N430, N411);
nand NAND3 (N431, N422, N296, N97);
nand NAND2 (N432, N421, N85);
and AND4 (N433, N427, N322, N394, N68);
xor XOR2 (N434, N432, N340);
nor NOR4 (N435, N408, N143, N123, N406);
nor NOR2 (N436, N426, N221);
and AND2 (N437, N433, N227);
not NOT1 (N438, N437);
and AND3 (N439, N431, N311, N428);
nor NOR4 (N440, N396, N2, N424, N59);
nand NAND4 (N441, N430, N112, N297, N365);
and AND4 (N442, N410, N138, N125, N165);
or OR3 (N443, N440, N411, N239);
buf BUF1 (N444, N439);
and AND2 (N445, N436, N210);
or OR3 (N446, N435, N259, N101);
or OR4 (N447, N443, N51, N46, N316);
nor NOR4 (N448, N444, N209, N431, N278);
nand NAND2 (N449, N441, N374);
nand NAND3 (N450, N445, N298, N253);
buf BUF1 (N451, N434);
buf BUF1 (N452, N407);
nand NAND2 (N453, N448, N219);
or OR4 (N454, N450, N157, N163, N68);
not NOT1 (N455, N454);
and AND2 (N456, N447, N419);
nor NOR2 (N457, N442, N9);
or OR2 (N458, N449, N456);
xor XOR2 (N459, N184, N8);
not NOT1 (N460, N457);
xor XOR2 (N461, N460, N217);
nor NOR4 (N462, N429, N385, N295, N138);
nor NOR4 (N463, N453, N359, N2, N201);
not NOT1 (N464, N446);
and AND2 (N465, N451, N70);
and AND2 (N466, N462, N147);
or OR2 (N467, N466, N394);
nand NAND3 (N468, N459, N119, N68);
and AND4 (N469, N452, N433, N430, N18);
nand NAND3 (N470, N461, N332, N155);
xor XOR2 (N471, N438, N176);
nand NAND4 (N472, N468, N96, N270, N301);
or OR4 (N473, N458, N102, N363, N347);
and AND4 (N474, N469, N176, N74, N74);
nand NAND3 (N475, N473, N446, N461);
nand NAND4 (N476, N470, N195, N227, N180);
nor NOR2 (N477, N476, N209);
buf BUF1 (N478, N467);
buf BUF1 (N479, N475);
and AND4 (N480, N478, N293, N131, N434);
not NOT1 (N481, N455);
nand NAND4 (N482, N471, N308, N19, N116);
xor XOR2 (N483, N472, N358);
nor NOR2 (N484, N482, N347);
nand NAND4 (N485, N480, N411, N477, N100);
nor NOR4 (N486, N29, N280, N479, N241);
xor XOR2 (N487, N19, N470);
and AND2 (N488, N465, N61);
and AND3 (N489, N485, N78, N21);
nor NOR3 (N490, N489, N268, N173);
and AND4 (N491, N488, N450, N19, N195);
nand NAND4 (N492, N481, N228, N367, N160);
nor NOR4 (N493, N474, N45, N84, N332);
xor XOR2 (N494, N486, N208);
and AND4 (N495, N487, N85, N268, N214);
xor XOR2 (N496, N494, N40);
xor XOR2 (N497, N491, N300);
xor XOR2 (N498, N493, N420);
xor XOR2 (N499, N490, N166);
buf BUF1 (N500, N497);
or OR4 (N501, N495, N491, N310, N21);
and AND2 (N502, N496, N161);
nand NAND3 (N503, N484, N38, N127);
nor NOR2 (N504, N501, N100);
and AND2 (N505, N499, N133);
nand NAND4 (N506, N502, N162, N270, N23);
and AND3 (N507, N492, N124, N125);
buf BUF1 (N508, N463);
nand NAND2 (N509, N464, N286);
or OR4 (N510, N504, N457, N133, N44);
nor NOR4 (N511, N506, N443, N260, N9);
nand NAND4 (N512, N508, N286, N74, N316);
nand NAND4 (N513, N511, N104, N279, N497);
xor XOR2 (N514, N505, N244);
and AND4 (N515, N510, N315, N478, N147);
or OR2 (N516, N503, N92);
xor XOR2 (N517, N507, N473);
or OR3 (N518, N509, N155, N431);
not NOT1 (N519, N516);
xor XOR2 (N520, N514, N464);
nand NAND2 (N521, N513, N41);
buf BUF1 (N522, N512);
xor XOR2 (N523, N483, N58);
buf BUF1 (N524, N500);
xor XOR2 (N525, N518, N143);
or OR2 (N526, N520, N145);
nor NOR2 (N527, N525, N518);
not NOT1 (N528, N517);
or OR4 (N529, N524, N186, N8, N193);
nor NOR2 (N530, N527, N49);
nor NOR3 (N531, N526, N315, N335);
xor XOR2 (N532, N528, N204);
buf BUF1 (N533, N529);
not NOT1 (N534, N523);
and AND3 (N535, N521, N23, N184);
buf BUF1 (N536, N498);
buf BUF1 (N537, N531);
nand NAND3 (N538, N537, N517, N173);
nand NAND4 (N539, N515, N180, N372, N382);
nor NOR4 (N540, N539, N464, N184, N273);
buf BUF1 (N541, N535);
or OR2 (N542, N541, N96);
nor NOR4 (N543, N532, N206, N356, N431);
buf BUF1 (N544, N536);
nor NOR2 (N545, N538, N537);
buf BUF1 (N546, N534);
and AND4 (N547, N533, N160, N349, N273);
nand NAND2 (N548, N540, N401);
not NOT1 (N549, N548);
or OR4 (N550, N543, N440, N490, N391);
or OR4 (N551, N549, N430, N86, N430);
and AND3 (N552, N519, N105, N80);
nor NOR2 (N553, N545, N512);
buf BUF1 (N554, N522);
nand NAND3 (N555, N544, N460, N82);
xor XOR2 (N556, N551, N33);
nor NOR3 (N557, N530, N302, N273);
buf BUF1 (N558, N542);
not NOT1 (N559, N546);
xor XOR2 (N560, N552, N521);
not NOT1 (N561, N554);
nand NAND2 (N562, N550, N538);
xor XOR2 (N563, N547, N386);
or OR3 (N564, N560, N257, N437);
and AND2 (N565, N557, N309);
buf BUF1 (N566, N562);
buf BUF1 (N567, N559);
or OR3 (N568, N558, N459, N48);
xor XOR2 (N569, N565, N77);
or OR3 (N570, N555, N384, N355);
xor XOR2 (N571, N553, N44);
nand NAND2 (N572, N563, N506);
buf BUF1 (N573, N564);
nor NOR3 (N574, N571, N248, N254);
buf BUF1 (N575, N569);
nor NOR2 (N576, N573, N264);
buf BUF1 (N577, N572);
xor XOR2 (N578, N556, N472);
buf BUF1 (N579, N568);
xor XOR2 (N580, N576, N200);
and AND2 (N581, N578, N506);
and AND2 (N582, N575, N574);
and AND2 (N583, N287, N340);
buf BUF1 (N584, N567);
not NOT1 (N585, N581);
and AND4 (N586, N561, N265, N550, N545);
or OR4 (N587, N586, N106, N373, N103);
nor NOR3 (N588, N577, N133, N313);
xor XOR2 (N589, N582, N224);
buf BUF1 (N590, N570);
not NOT1 (N591, N589);
xor XOR2 (N592, N566, N325);
nand NAND4 (N593, N583, N117, N11, N25);
nor NOR4 (N594, N587, N9, N498, N321);
nor NOR2 (N595, N579, N342);
or OR3 (N596, N592, N461, N585);
buf BUF1 (N597, N55);
xor XOR2 (N598, N597, N350);
nand NAND4 (N599, N598, N169, N82, N443);
nand NAND4 (N600, N594, N148, N199, N56);
or OR4 (N601, N593, N134, N540, N399);
nor NOR4 (N602, N595, N582, N13, N534);
buf BUF1 (N603, N599);
or OR3 (N604, N584, N57, N146);
nand NAND3 (N605, N591, N110, N306);
xor XOR2 (N606, N605, N293);
nand NAND2 (N607, N604, N441);
xor XOR2 (N608, N606, N32);
nor NOR4 (N609, N588, N330, N378, N429);
and AND2 (N610, N596, N187);
and AND2 (N611, N601, N310);
nor NOR2 (N612, N608, N459);
nand NAND2 (N613, N611, N69);
or OR2 (N614, N610, N554);
buf BUF1 (N615, N602);
or OR2 (N616, N590, N111);
xor XOR2 (N617, N607, N151);
buf BUF1 (N618, N580);
not NOT1 (N619, N618);
not NOT1 (N620, N603);
not NOT1 (N621, N612);
nor NOR2 (N622, N609, N258);
nand NAND2 (N623, N621, N104);
xor XOR2 (N624, N623, N282);
and AND4 (N625, N600, N197, N340, N386);
buf BUF1 (N626, N613);
nor NOR2 (N627, N616, N522);
buf BUF1 (N628, N622);
nand NAND4 (N629, N620, N179, N86, N198);
buf BUF1 (N630, N628);
xor XOR2 (N631, N630, N550);
buf BUF1 (N632, N631);
nand NAND3 (N633, N625, N332, N371);
nand NAND4 (N634, N615, N598, N425, N198);
buf BUF1 (N635, N633);
nor NOR2 (N636, N627, N397);
nand NAND3 (N637, N629, N207, N332);
nor NOR4 (N638, N619, N399, N597, N555);
or OR2 (N639, N635, N45);
buf BUF1 (N640, N624);
nand NAND3 (N641, N632, N367, N379);
xor XOR2 (N642, N636, N236);
buf BUF1 (N643, N641);
not NOT1 (N644, N637);
not NOT1 (N645, N642);
not NOT1 (N646, N644);
not NOT1 (N647, N643);
and AND4 (N648, N638, N295, N99, N626);
not NOT1 (N649, N414);
and AND2 (N650, N647, N264);
not NOT1 (N651, N649);
nor NOR4 (N652, N639, N125, N55, N627);
or OR2 (N653, N614, N194);
nand NAND3 (N654, N645, N649, N20);
not NOT1 (N655, N648);
or OR2 (N656, N617, N47);
nand NAND2 (N657, N640, N285);
not NOT1 (N658, N656);
and AND4 (N659, N652, N161, N640, N100);
not NOT1 (N660, N654);
nor NOR2 (N661, N655, N312);
buf BUF1 (N662, N660);
nand NAND3 (N663, N646, N297, N660);
buf BUF1 (N664, N662);
not NOT1 (N665, N658);
nor NOR4 (N666, N650, N11, N92, N409);
buf BUF1 (N667, N664);
not NOT1 (N668, N653);
xor XOR2 (N669, N665, N221);
xor XOR2 (N670, N666, N279);
nand NAND2 (N671, N670, N95);
nor NOR2 (N672, N659, N553);
not NOT1 (N673, N668);
nor NOR4 (N674, N671, N634, N65, N41);
buf BUF1 (N675, N664);
xor XOR2 (N676, N651, N92);
and AND2 (N677, N657, N276);
buf BUF1 (N678, N674);
and AND3 (N679, N667, N434, N656);
buf BUF1 (N680, N673);
not NOT1 (N681, N680);
buf BUF1 (N682, N676);
xor XOR2 (N683, N681, N360);
not NOT1 (N684, N682);
or OR2 (N685, N678, N621);
buf BUF1 (N686, N679);
not NOT1 (N687, N684);
nand NAND2 (N688, N687, N566);
nand NAND4 (N689, N669, N179, N405, N89);
nor NOR3 (N690, N661, N668, N505);
buf BUF1 (N691, N690);
and AND2 (N692, N663, N46);
xor XOR2 (N693, N672, N422);
buf BUF1 (N694, N685);
or OR4 (N695, N691, N72, N278, N84);
xor XOR2 (N696, N689, N481);
nand NAND2 (N697, N688, N71);
not NOT1 (N698, N695);
xor XOR2 (N699, N692, N238);
not NOT1 (N700, N675);
or OR4 (N701, N697, N671, N210, N640);
not NOT1 (N702, N694);
or OR4 (N703, N702, N94, N379, N56);
buf BUF1 (N704, N683);
and AND4 (N705, N686, N397, N127, N299);
nor NOR4 (N706, N696, N174, N34, N610);
buf BUF1 (N707, N701);
and AND3 (N708, N703, N114, N20);
xor XOR2 (N709, N706, N109);
nor NOR2 (N710, N707, N198);
buf BUF1 (N711, N698);
nand NAND4 (N712, N693, N68, N439, N188);
nand NAND2 (N713, N710, N500);
buf BUF1 (N714, N711);
nor NOR3 (N715, N714, N653, N321);
xor XOR2 (N716, N708, N313);
buf BUF1 (N717, N712);
nand NAND2 (N718, N716, N184);
not NOT1 (N719, N717);
or OR4 (N720, N704, N359, N186, N336);
and AND4 (N721, N719, N444, N414, N116);
or OR3 (N722, N720, N174, N451);
nor NOR3 (N723, N677, N148, N701);
not NOT1 (N724, N718);
xor XOR2 (N725, N724, N176);
nor NOR3 (N726, N715, N20, N102);
xor XOR2 (N727, N705, N346);
or OR3 (N728, N699, N655, N385);
not NOT1 (N729, N726);
not NOT1 (N730, N709);
not NOT1 (N731, N729);
xor XOR2 (N732, N713, N139);
buf BUF1 (N733, N725);
nor NOR4 (N734, N700, N61, N189, N287);
nor NOR4 (N735, N731, N373, N644, N237);
nor NOR2 (N736, N732, N401);
xor XOR2 (N737, N734, N648);
buf BUF1 (N738, N722);
or OR3 (N739, N738, N679, N459);
or OR2 (N740, N727, N227);
and AND3 (N741, N735, N317, N355);
xor XOR2 (N742, N733, N401);
xor XOR2 (N743, N737, N266);
not NOT1 (N744, N723);
buf BUF1 (N745, N736);
xor XOR2 (N746, N739, N588);
buf BUF1 (N747, N744);
buf BUF1 (N748, N745);
not NOT1 (N749, N743);
buf BUF1 (N750, N748);
or OR2 (N751, N749, N245);
nor NOR4 (N752, N728, N462, N365, N433);
nor NOR4 (N753, N730, N72, N7, N303);
nand NAND3 (N754, N746, N130, N241);
and AND3 (N755, N751, N85, N286);
nor NOR4 (N756, N752, N114, N318, N536);
and AND4 (N757, N753, N118, N385, N304);
nor NOR3 (N758, N755, N497, N85);
or OR4 (N759, N747, N32, N423, N92);
or OR2 (N760, N759, N326);
and AND2 (N761, N750, N739);
and AND3 (N762, N760, N577, N517);
not NOT1 (N763, N740);
nand NAND2 (N764, N762, N576);
xor XOR2 (N765, N721, N561);
not NOT1 (N766, N758);
not NOT1 (N767, N766);
and AND4 (N768, N742, N74, N171, N224);
nor NOR4 (N769, N767, N741, N733, N248);
and AND3 (N770, N444, N300, N645);
or OR4 (N771, N754, N691, N708, N542);
not NOT1 (N772, N764);
nor NOR4 (N773, N763, N513, N48, N678);
nor NOR3 (N774, N770, N77, N572);
not NOT1 (N775, N771);
or OR3 (N776, N775, N739, N564);
and AND4 (N777, N757, N265, N459, N539);
xor XOR2 (N778, N774, N277);
and AND3 (N779, N765, N248, N771);
and AND3 (N780, N756, N493, N204);
xor XOR2 (N781, N761, N642);
xor XOR2 (N782, N772, N402);
not NOT1 (N783, N776);
and AND2 (N784, N781, N783);
nand NAND3 (N785, N683, N288, N765);
nor NOR4 (N786, N780, N718, N652, N373);
nor NOR4 (N787, N778, N30, N118, N275);
nor NOR2 (N788, N787, N577);
buf BUF1 (N789, N786);
and AND3 (N790, N789, N691, N346);
buf BUF1 (N791, N768);
xor XOR2 (N792, N784, N716);
xor XOR2 (N793, N769, N764);
not NOT1 (N794, N779);
and AND3 (N795, N792, N428, N77);
nor NOR3 (N796, N791, N473, N283);
and AND2 (N797, N773, N82);
buf BUF1 (N798, N796);
nand NAND2 (N799, N795, N757);
and AND3 (N800, N794, N728, N327);
buf BUF1 (N801, N790);
buf BUF1 (N802, N785);
not NOT1 (N803, N797);
nand NAND2 (N804, N788, N462);
or OR3 (N805, N799, N603, N485);
buf BUF1 (N806, N802);
buf BUF1 (N807, N803);
nor NOR4 (N808, N804, N661, N336, N342);
xor XOR2 (N809, N782, N288);
buf BUF1 (N810, N800);
nor NOR3 (N811, N807, N457, N571);
xor XOR2 (N812, N806, N29);
and AND2 (N813, N793, N280);
not NOT1 (N814, N811);
not NOT1 (N815, N814);
nand NAND4 (N816, N809, N787, N217, N684);
xor XOR2 (N817, N816, N182);
xor XOR2 (N818, N801, N453);
nor NOR3 (N819, N817, N733, N565);
or OR2 (N820, N798, N61);
xor XOR2 (N821, N819, N242);
and AND3 (N822, N821, N475, N429);
nor NOR4 (N823, N812, N727, N41, N33);
or OR2 (N824, N805, N446);
buf BUF1 (N825, N818);
or OR4 (N826, N825, N427, N611, N317);
and AND3 (N827, N826, N325, N17);
and AND4 (N828, N823, N162, N597, N79);
nor NOR2 (N829, N808, N694);
and AND2 (N830, N828, N813);
nand NAND2 (N831, N484, N619);
nor NOR2 (N832, N829, N791);
nand NAND2 (N833, N827, N756);
nor NOR2 (N834, N815, N689);
xor XOR2 (N835, N832, N510);
or OR3 (N836, N830, N7, N33);
buf BUF1 (N837, N834);
xor XOR2 (N838, N820, N3);
and AND3 (N839, N838, N517, N83);
nor NOR3 (N840, N835, N563, N394);
nor NOR4 (N841, N824, N136, N145, N39);
nor NOR4 (N842, N831, N557, N270, N502);
and AND4 (N843, N837, N639, N332, N559);
nor NOR2 (N844, N843, N752);
buf BUF1 (N845, N833);
xor XOR2 (N846, N839, N119);
nand NAND4 (N847, N842, N89, N367, N276);
and AND2 (N848, N847, N38);
or OR4 (N849, N836, N94, N137, N687);
nor NOR3 (N850, N810, N120, N637);
nor NOR3 (N851, N840, N740, N455);
nor NOR2 (N852, N844, N337);
nor NOR3 (N853, N822, N404, N433);
xor XOR2 (N854, N777, N98);
not NOT1 (N855, N852);
and AND3 (N856, N851, N598, N56);
nor NOR4 (N857, N855, N33, N40, N58);
not NOT1 (N858, N857);
nor NOR3 (N859, N841, N406, N822);
buf BUF1 (N860, N850);
xor XOR2 (N861, N856, N631);
or OR4 (N862, N859, N661, N85, N571);
nor NOR2 (N863, N858, N282);
not NOT1 (N864, N860);
or OR2 (N865, N862, N654);
not NOT1 (N866, N845);
or OR4 (N867, N864, N41, N85, N823);
and AND2 (N868, N854, N62);
not NOT1 (N869, N846);
buf BUF1 (N870, N869);
not NOT1 (N871, N861);
not NOT1 (N872, N867);
xor XOR2 (N873, N872, N710);
not NOT1 (N874, N868);
not NOT1 (N875, N866);
or OR2 (N876, N875, N639);
and AND4 (N877, N853, N777, N652, N637);
not NOT1 (N878, N863);
xor XOR2 (N879, N874, N760);
xor XOR2 (N880, N849, N294);
buf BUF1 (N881, N879);
buf BUF1 (N882, N871);
nand NAND4 (N883, N881, N850, N722, N507);
nand NAND3 (N884, N876, N752, N584);
not NOT1 (N885, N848);
xor XOR2 (N886, N865, N244);
and AND3 (N887, N885, N765, N714);
and AND3 (N888, N878, N412, N671);
buf BUF1 (N889, N877);
nor NOR2 (N890, N886, N800);
xor XOR2 (N891, N883, N733);
or OR2 (N892, N880, N117);
buf BUF1 (N893, N892);
or OR2 (N894, N889, N692);
or OR3 (N895, N893, N158, N210);
nor NOR3 (N896, N890, N717, N347);
or OR3 (N897, N887, N97, N588);
or OR2 (N898, N870, N638);
nor NOR4 (N899, N898, N439, N887, N225);
xor XOR2 (N900, N896, N185);
nor NOR4 (N901, N884, N427, N730, N83);
nor NOR3 (N902, N873, N279, N431);
and AND3 (N903, N888, N224, N786);
not NOT1 (N904, N901);
or OR2 (N905, N899, N68);
or OR2 (N906, N891, N460);
nand NAND3 (N907, N906, N865, N648);
or OR4 (N908, N904, N795, N501, N484);
or OR2 (N909, N897, N850);
not NOT1 (N910, N909);
xor XOR2 (N911, N907, N157);
nor NOR4 (N912, N905, N363, N358, N440);
nand NAND4 (N913, N900, N278, N706, N598);
nand NAND4 (N914, N908, N123, N320, N129);
and AND3 (N915, N882, N263, N601);
or OR3 (N916, N894, N453, N812);
nand NAND2 (N917, N916, N254);
buf BUF1 (N918, N917);
buf BUF1 (N919, N911);
or OR2 (N920, N902, N660);
or OR2 (N921, N918, N261);
buf BUF1 (N922, N913);
xor XOR2 (N923, N912, N538);
nor NOR2 (N924, N922, N809);
or OR4 (N925, N919, N574, N281, N661);
buf BUF1 (N926, N903);
nor NOR2 (N927, N895, N893);
buf BUF1 (N928, N923);
nor NOR2 (N929, N924, N411);
and AND2 (N930, N928, N678);
and AND3 (N931, N915, N508, N718);
nand NAND3 (N932, N925, N109, N303);
nor NOR4 (N933, N910, N401, N254, N575);
buf BUF1 (N934, N921);
nor NOR4 (N935, N926, N615, N212, N379);
and AND3 (N936, N931, N532, N206);
or OR3 (N937, N933, N917, N339);
buf BUF1 (N938, N934);
buf BUF1 (N939, N930);
xor XOR2 (N940, N935, N518);
nor NOR4 (N941, N937, N118, N728, N500);
buf BUF1 (N942, N932);
or OR4 (N943, N942, N449, N291, N414);
nand NAND4 (N944, N939, N703, N524, N809);
not NOT1 (N945, N920);
buf BUF1 (N946, N943);
not NOT1 (N947, N946);
nand NAND4 (N948, N944, N792, N409, N569);
and AND4 (N949, N940, N932, N245, N758);
and AND3 (N950, N948, N783, N227);
nand NAND2 (N951, N938, N317);
nand NAND2 (N952, N949, N285);
nor NOR4 (N953, N914, N52, N523, N645);
and AND3 (N954, N952, N618, N900);
and AND4 (N955, N927, N6, N867, N138);
and AND2 (N956, N954, N692);
xor XOR2 (N957, N956, N164);
buf BUF1 (N958, N929);
buf BUF1 (N959, N951);
or OR4 (N960, N955, N937, N80, N355);
nor NOR4 (N961, N959, N71, N740, N770);
buf BUF1 (N962, N936);
nand NAND3 (N963, N941, N869, N207);
or OR4 (N964, N947, N231, N551, N303);
buf BUF1 (N965, N958);
nor NOR4 (N966, N945, N766, N854, N73);
buf BUF1 (N967, N961);
not NOT1 (N968, N957);
or OR2 (N969, N953, N512);
or OR4 (N970, N968, N671, N469, N18);
xor XOR2 (N971, N950, N308);
and AND3 (N972, N964, N705, N53);
nand NAND2 (N973, N969, N50);
not NOT1 (N974, N963);
buf BUF1 (N975, N966);
or OR4 (N976, N973, N370, N906, N253);
nor NOR4 (N977, N967, N448, N428, N553);
not NOT1 (N978, N965);
xor XOR2 (N979, N970, N447);
nor NOR4 (N980, N976, N461, N228, N742);
and AND4 (N981, N962, N954, N284, N362);
or OR4 (N982, N960, N850, N163, N814);
and AND2 (N983, N974, N613);
nand NAND3 (N984, N981, N68, N539);
nor NOR4 (N985, N978, N439, N408, N924);
or OR4 (N986, N984, N661, N894, N26);
buf BUF1 (N987, N972);
not NOT1 (N988, N975);
xor XOR2 (N989, N980, N393);
buf BUF1 (N990, N979);
and AND3 (N991, N989, N409, N664);
and AND3 (N992, N977, N350, N7);
nor NOR4 (N993, N971, N425, N621, N710);
and AND3 (N994, N985, N234, N616);
nor NOR4 (N995, N983, N898, N246, N631);
nor NOR2 (N996, N991, N57);
and AND4 (N997, N982, N835, N476, N134);
not NOT1 (N998, N993);
xor XOR2 (N999, N988, N310);
nor NOR2 (N1000, N990, N988);
nand NAND2 (N1001, N987, N763);
buf BUF1 (N1002, N986);
and AND4 (N1003, N1001, N60, N486, N827);
xor XOR2 (N1004, N1003, N685);
not NOT1 (N1005, N998);
or OR2 (N1006, N994, N815);
or OR3 (N1007, N999, N759, N381);
and AND2 (N1008, N1002, N518);
buf BUF1 (N1009, N1004);
and AND4 (N1010, N997, N669, N236, N600);
or OR4 (N1011, N996, N803, N6, N607);
buf BUF1 (N1012, N1010);
or OR3 (N1013, N1007, N182, N339);
and AND2 (N1014, N992, N692);
and AND4 (N1015, N1012, N438, N30, N913);
nor NOR2 (N1016, N1015, N83);
and AND4 (N1017, N1000, N644, N359, N210);
nor NOR2 (N1018, N995, N538);
buf BUF1 (N1019, N1011);
and AND3 (N1020, N1013, N772, N860);
or OR4 (N1021, N1018, N218, N489, N40);
nor NOR3 (N1022, N1017, N555, N429);
xor XOR2 (N1023, N1019, N806);
and AND4 (N1024, N1009, N15, N614, N636);
or OR2 (N1025, N1014, N107);
or OR3 (N1026, N1008, N119, N105);
nor NOR4 (N1027, N1006, N677, N1024, N348);
nor NOR3 (N1028, N663, N540, N760);
or OR2 (N1029, N1016, N706);
xor XOR2 (N1030, N1020, N773);
or OR3 (N1031, N1021, N1021, N150);
buf BUF1 (N1032, N1005);
nor NOR3 (N1033, N1027, N293, N1032);
nor NOR2 (N1034, N838, N66);
or OR3 (N1035, N1030, N95, N164);
nor NOR4 (N1036, N1022, N509, N71, N189);
nand NAND2 (N1037, N1028, N657);
xor XOR2 (N1038, N1029, N1000);
and AND3 (N1039, N1033, N436, N856);
buf BUF1 (N1040, N1039);
buf BUF1 (N1041, N1037);
xor XOR2 (N1042, N1040, N620);
nand NAND2 (N1043, N1035, N448);
nor NOR3 (N1044, N1034, N80, N555);
and AND3 (N1045, N1023, N34, N431);
xor XOR2 (N1046, N1043, N128);
or OR3 (N1047, N1045, N120, N513);
nand NAND4 (N1048, N1041, N637, N535, N527);
nor NOR3 (N1049, N1044, N527, N57);
nand NAND3 (N1050, N1046, N405, N407);
not NOT1 (N1051, N1036);
not NOT1 (N1052, N1026);
xor XOR2 (N1053, N1047, N402);
not NOT1 (N1054, N1048);
not NOT1 (N1055, N1050);
nor NOR2 (N1056, N1053, N704);
or OR3 (N1057, N1025, N605, N922);
or OR2 (N1058, N1052, N271);
or OR2 (N1059, N1057, N360);
or OR3 (N1060, N1054, N764, N613);
buf BUF1 (N1061, N1058);
buf BUF1 (N1062, N1060);
and AND3 (N1063, N1062, N102, N624);
not NOT1 (N1064, N1031);
nand NAND4 (N1065, N1049, N490, N930, N300);
or OR3 (N1066, N1059, N661, N200);
and AND2 (N1067, N1055, N755);
or OR2 (N1068, N1038, N570);
xor XOR2 (N1069, N1067, N300);
and AND3 (N1070, N1064, N8, N774);
xor XOR2 (N1071, N1066, N716);
and AND2 (N1072, N1056, N541);
or OR4 (N1073, N1061, N883, N869, N119);
nor NOR4 (N1074, N1068, N892, N712, N464);
xor XOR2 (N1075, N1065, N301);
buf BUF1 (N1076, N1074);
and AND4 (N1077, N1076, N1017, N229, N991);
not NOT1 (N1078, N1077);
buf BUF1 (N1079, N1071);
or OR2 (N1080, N1075, N1059);
or OR2 (N1081, N1078, N695);
nand NAND4 (N1082, N1069, N178, N718, N214);
nand NAND2 (N1083, N1080, N507);
nor NOR4 (N1084, N1042, N673, N203, N645);
nor NOR3 (N1085, N1082, N1049, N311);
or OR4 (N1086, N1063, N882, N264, N977);
and AND3 (N1087, N1051, N51, N778);
nor NOR4 (N1088, N1072, N99, N176, N429);
nor NOR4 (N1089, N1088, N744, N1050, N999);
nand NAND3 (N1090, N1085, N362, N602);
xor XOR2 (N1091, N1084, N340);
or OR3 (N1092, N1073, N235, N1013);
xor XOR2 (N1093, N1083, N301);
nand NAND4 (N1094, N1090, N517, N131, N428);
and AND2 (N1095, N1091, N531);
nand NAND3 (N1096, N1081, N354, N939);
buf BUF1 (N1097, N1079);
not NOT1 (N1098, N1092);
not NOT1 (N1099, N1086);
or OR4 (N1100, N1099, N906, N920, N1006);
nor NOR2 (N1101, N1095, N932);
and AND2 (N1102, N1096, N219);
nand NAND4 (N1103, N1094, N1039, N434, N582);
not NOT1 (N1104, N1089);
buf BUF1 (N1105, N1087);
nor NOR2 (N1106, N1104, N482);
and AND2 (N1107, N1097, N31);
and AND2 (N1108, N1070, N366);
and AND2 (N1109, N1093, N242);
or OR3 (N1110, N1098, N305, N555);
not NOT1 (N1111, N1109);
buf BUF1 (N1112, N1105);
or OR4 (N1113, N1101, N192, N530, N144);
not NOT1 (N1114, N1111);
nor NOR4 (N1115, N1107, N875, N924, N394);
nor NOR2 (N1116, N1110, N1114);
xor XOR2 (N1117, N489, N747);
xor XOR2 (N1118, N1113, N27);
not NOT1 (N1119, N1106);
xor XOR2 (N1120, N1112, N685);
nand NAND3 (N1121, N1119, N537, N442);
not NOT1 (N1122, N1116);
nand NAND2 (N1123, N1117, N423);
nand NAND3 (N1124, N1100, N690, N233);
and AND3 (N1125, N1115, N387, N1003);
and AND4 (N1126, N1118, N249, N410, N624);
nand NAND4 (N1127, N1124, N95, N908, N768);
nand NAND2 (N1128, N1120, N936);
buf BUF1 (N1129, N1127);
nor NOR2 (N1130, N1122, N819);
xor XOR2 (N1131, N1102, N377);
not NOT1 (N1132, N1108);
buf BUF1 (N1133, N1125);
xor XOR2 (N1134, N1123, N448);
or OR4 (N1135, N1131, N466, N917, N984);
or OR4 (N1136, N1121, N342, N623, N428);
or OR3 (N1137, N1103, N485, N106);
not NOT1 (N1138, N1132);
nor NOR2 (N1139, N1138, N640);
and AND2 (N1140, N1136, N1040);
nor NOR3 (N1141, N1137, N922, N1134);
xor XOR2 (N1142, N1141, N1062);
nand NAND4 (N1143, N59, N266, N908, N78);
not NOT1 (N1144, N1130);
xor XOR2 (N1145, N1140, N60);
buf BUF1 (N1146, N1142);
nor NOR4 (N1147, N1135, N64, N764, N716);
or OR4 (N1148, N1145, N121, N1120, N161);
or OR2 (N1149, N1129, N217);
not NOT1 (N1150, N1148);
nor NOR2 (N1151, N1128, N128);
buf BUF1 (N1152, N1133);
and AND2 (N1153, N1143, N951);
nor NOR4 (N1154, N1146, N196, N643, N560);
not NOT1 (N1155, N1151);
not NOT1 (N1156, N1139);
xor XOR2 (N1157, N1154, N833);
or OR2 (N1158, N1157, N386);
or OR2 (N1159, N1155, N959);
not NOT1 (N1160, N1158);
not NOT1 (N1161, N1144);
xor XOR2 (N1162, N1160, N266);
and AND4 (N1163, N1126, N786, N545, N1006);
not NOT1 (N1164, N1149);
nand NAND2 (N1165, N1164, N757);
nor NOR3 (N1166, N1152, N492, N492);
buf BUF1 (N1167, N1163);
nand NAND2 (N1168, N1166, N769);
xor XOR2 (N1169, N1153, N362);
nand NAND2 (N1170, N1161, N449);
or OR4 (N1171, N1162, N1071, N498, N409);
xor XOR2 (N1172, N1169, N772);
buf BUF1 (N1173, N1171);
and AND2 (N1174, N1173, N1091);
or OR2 (N1175, N1150, N201);
not NOT1 (N1176, N1170);
nor NOR4 (N1177, N1176, N1006, N895, N11);
or OR2 (N1178, N1168, N609);
nand NAND2 (N1179, N1174, N1165);
nand NAND4 (N1180, N700, N759, N786, N621);
nor NOR3 (N1181, N1179, N1119, N782);
buf BUF1 (N1182, N1147);
buf BUF1 (N1183, N1156);
not NOT1 (N1184, N1167);
xor XOR2 (N1185, N1172, N552);
nor NOR4 (N1186, N1184, N794, N414, N14);
nand NAND2 (N1187, N1177, N1124);
and AND2 (N1188, N1186, N198);
not NOT1 (N1189, N1180);
not NOT1 (N1190, N1159);
nand NAND3 (N1191, N1188, N428, N363);
nor NOR2 (N1192, N1189, N182);
xor XOR2 (N1193, N1182, N1163);
nor NOR2 (N1194, N1193, N615);
or OR4 (N1195, N1191, N745, N813, N190);
xor XOR2 (N1196, N1181, N1195);
nand NAND4 (N1197, N193, N511, N659, N520);
nand NAND2 (N1198, N1178, N1001);
or OR2 (N1199, N1192, N58);
not NOT1 (N1200, N1175);
not NOT1 (N1201, N1187);
nor NOR4 (N1202, N1183, N471, N878, N1031);
not NOT1 (N1203, N1199);
xor XOR2 (N1204, N1201, N766);
xor XOR2 (N1205, N1190, N210);
not NOT1 (N1206, N1198);
or OR2 (N1207, N1200, N1052);
nor NOR3 (N1208, N1196, N565, N127);
not NOT1 (N1209, N1204);
buf BUF1 (N1210, N1197);
nand NAND3 (N1211, N1210, N576, N176);
nor NOR3 (N1212, N1209, N1096, N620);
and AND4 (N1213, N1206, N449, N600, N356);
or OR4 (N1214, N1194, N929, N277, N664);
not NOT1 (N1215, N1214);
nor NOR2 (N1216, N1205, N215);
or OR4 (N1217, N1203, N1061, N368, N49);
nor NOR2 (N1218, N1207, N877);
buf BUF1 (N1219, N1202);
or OR3 (N1220, N1185, N492, N851);
buf BUF1 (N1221, N1220);
xor XOR2 (N1222, N1213, N525);
nand NAND3 (N1223, N1217, N670, N154);
or OR4 (N1224, N1219, N274, N69, N1115);
or OR2 (N1225, N1212, N627);
or OR3 (N1226, N1224, N701, N726);
buf BUF1 (N1227, N1225);
buf BUF1 (N1228, N1216);
buf BUF1 (N1229, N1223);
buf BUF1 (N1230, N1228);
nand NAND2 (N1231, N1229, N433);
and AND2 (N1232, N1230, N1182);
xor XOR2 (N1233, N1227, N989);
nor NOR4 (N1234, N1232, N511, N44, N161);
buf BUF1 (N1235, N1233);
and AND2 (N1236, N1211, N731);
nor NOR4 (N1237, N1215, N880, N215, N890);
nor NOR4 (N1238, N1218, N580, N1086, N1003);
nor NOR2 (N1239, N1238, N439);
xor XOR2 (N1240, N1234, N263);
or OR3 (N1241, N1240, N1080, N477);
nor NOR4 (N1242, N1239, N1193, N89, N735);
or OR2 (N1243, N1241, N693);
nand NAND2 (N1244, N1242, N607);
and AND3 (N1245, N1235, N252, N812);
nor NOR2 (N1246, N1208, N939);
buf BUF1 (N1247, N1222);
or OR4 (N1248, N1243, N961, N77, N123);
nor NOR4 (N1249, N1231, N659, N797, N1062);
xor XOR2 (N1250, N1248, N560);
nand NAND3 (N1251, N1250, N380, N876);
buf BUF1 (N1252, N1221);
nand NAND4 (N1253, N1247, N281, N682, N464);
nand NAND3 (N1254, N1236, N1207, N1223);
or OR2 (N1255, N1245, N786);
nand NAND2 (N1256, N1226, N540);
and AND2 (N1257, N1252, N731);
and AND2 (N1258, N1246, N699);
nor NOR2 (N1259, N1244, N558);
nand NAND2 (N1260, N1259, N813);
nor NOR3 (N1261, N1251, N1203, N1089);
nand NAND3 (N1262, N1258, N136, N120);
nand NAND4 (N1263, N1253, N953, N945, N1197);
buf BUF1 (N1264, N1257);
buf BUF1 (N1265, N1249);
or OR3 (N1266, N1261, N615, N34);
xor XOR2 (N1267, N1260, N592);
and AND3 (N1268, N1265, N301, N513);
xor XOR2 (N1269, N1266, N336);
or OR2 (N1270, N1254, N279);
xor XOR2 (N1271, N1267, N666);
and AND3 (N1272, N1262, N80, N771);
nand NAND3 (N1273, N1268, N568, N1114);
or OR3 (N1274, N1256, N56, N1060);
nand NAND3 (N1275, N1274, N450, N698);
not NOT1 (N1276, N1273);
xor XOR2 (N1277, N1276, N939);
not NOT1 (N1278, N1237);
nor NOR3 (N1279, N1269, N523, N718);
and AND2 (N1280, N1263, N813);
nor NOR3 (N1281, N1278, N1012, N1040);
xor XOR2 (N1282, N1281, N809);
nor NOR4 (N1283, N1277, N725, N886, N398);
and AND3 (N1284, N1271, N1031, N585);
nor NOR3 (N1285, N1270, N265, N1081);
buf BUF1 (N1286, N1282);
not NOT1 (N1287, N1264);
not NOT1 (N1288, N1255);
nor NOR4 (N1289, N1283, N494, N790, N1240);
buf BUF1 (N1290, N1275);
not NOT1 (N1291, N1287);
nand NAND3 (N1292, N1279, N1182, N326);
xor XOR2 (N1293, N1288, N685);
or OR2 (N1294, N1280, N1166);
xor XOR2 (N1295, N1291, N424);
and AND3 (N1296, N1289, N134, N851);
nor NOR3 (N1297, N1290, N693, N411);
xor XOR2 (N1298, N1296, N93);
xor XOR2 (N1299, N1285, N705);
or OR2 (N1300, N1272, N408);
or OR3 (N1301, N1284, N689, N8);
or OR4 (N1302, N1293, N462, N674, N35);
nand NAND2 (N1303, N1301, N188);
xor XOR2 (N1304, N1300, N1254);
nor NOR3 (N1305, N1302, N1215, N427);
not NOT1 (N1306, N1299);
or OR2 (N1307, N1295, N482);
xor XOR2 (N1308, N1286, N1164);
and AND3 (N1309, N1306, N463, N26);
or OR3 (N1310, N1305, N612, N958);
buf BUF1 (N1311, N1304);
and AND3 (N1312, N1297, N304, N1104);
nor NOR4 (N1313, N1303, N863, N787, N1206);
buf BUF1 (N1314, N1310);
xor XOR2 (N1315, N1313, N286);
nor NOR4 (N1316, N1298, N892, N1014, N870);
nor NOR2 (N1317, N1307, N1151);
xor XOR2 (N1318, N1316, N293);
not NOT1 (N1319, N1309);
and AND2 (N1320, N1319, N1295);
buf BUF1 (N1321, N1292);
and AND3 (N1322, N1318, N935, N1187);
buf BUF1 (N1323, N1320);
xor XOR2 (N1324, N1294, N9);
not NOT1 (N1325, N1323);
not NOT1 (N1326, N1321);
xor XOR2 (N1327, N1311, N19);
nand NAND3 (N1328, N1324, N295, N1157);
buf BUF1 (N1329, N1326);
buf BUF1 (N1330, N1327);
xor XOR2 (N1331, N1328, N765);
xor XOR2 (N1332, N1330, N1138);
nand NAND3 (N1333, N1314, N634, N513);
not NOT1 (N1334, N1333);
nand NAND3 (N1335, N1331, N100, N1044);
not NOT1 (N1336, N1308);
not NOT1 (N1337, N1334);
not NOT1 (N1338, N1325);
not NOT1 (N1339, N1338);
and AND2 (N1340, N1329, N898);
or OR4 (N1341, N1339, N540, N1222, N1325);
nand NAND4 (N1342, N1312, N438, N1246, N1210);
or OR2 (N1343, N1315, N1105);
xor XOR2 (N1344, N1342, N523);
not NOT1 (N1345, N1344);
nor NOR4 (N1346, N1345, N1228, N1297, N1007);
xor XOR2 (N1347, N1341, N1300);
xor XOR2 (N1348, N1317, N393);
xor XOR2 (N1349, N1332, N910);
or OR2 (N1350, N1346, N828);
nand NAND4 (N1351, N1348, N900, N1103, N764);
buf BUF1 (N1352, N1336);
and AND2 (N1353, N1352, N404);
xor XOR2 (N1354, N1349, N525);
xor XOR2 (N1355, N1335, N1182);
not NOT1 (N1356, N1343);
or OR3 (N1357, N1340, N116, N305);
nor NOR2 (N1358, N1355, N975);
xor XOR2 (N1359, N1354, N1131);
xor XOR2 (N1360, N1351, N777);
nand NAND4 (N1361, N1357, N821, N705, N312);
not NOT1 (N1362, N1347);
and AND4 (N1363, N1356, N797, N94, N486);
xor XOR2 (N1364, N1362, N1020);
buf BUF1 (N1365, N1359);
or OR3 (N1366, N1365, N520, N979);
nor NOR4 (N1367, N1337, N621, N302, N224);
buf BUF1 (N1368, N1363);
buf BUF1 (N1369, N1360);
nand NAND4 (N1370, N1358, N610, N1276, N830);
not NOT1 (N1371, N1350);
not NOT1 (N1372, N1364);
xor XOR2 (N1373, N1361, N431);
nor NOR3 (N1374, N1368, N793, N1310);
xor XOR2 (N1375, N1369, N1312);
buf BUF1 (N1376, N1366);
not NOT1 (N1377, N1376);
xor XOR2 (N1378, N1377, N1062);
xor XOR2 (N1379, N1367, N1016);
nand NAND3 (N1380, N1374, N654, N851);
and AND2 (N1381, N1380, N1341);
nand NAND2 (N1382, N1375, N362);
buf BUF1 (N1383, N1378);
or OR4 (N1384, N1379, N332, N1207, N1130);
or OR2 (N1385, N1373, N883);
and AND2 (N1386, N1382, N901);
not NOT1 (N1387, N1371);
nor NOR3 (N1388, N1381, N350, N1116);
nand NAND3 (N1389, N1353, N1230, N459);
not NOT1 (N1390, N1370);
xor XOR2 (N1391, N1322, N129);
or OR3 (N1392, N1385, N231, N488);
xor XOR2 (N1393, N1389, N314);
and AND2 (N1394, N1384, N317);
nand NAND4 (N1395, N1391, N916, N828, N1325);
and AND2 (N1396, N1386, N376);
buf BUF1 (N1397, N1395);
buf BUF1 (N1398, N1390);
nand NAND4 (N1399, N1387, N8, N140, N602);
nand NAND4 (N1400, N1388, N570, N215, N128);
not NOT1 (N1401, N1383);
buf BUF1 (N1402, N1392);
nor NOR2 (N1403, N1396, N297);
or OR2 (N1404, N1398, N822);
or OR3 (N1405, N1402, N529, N577);
or OR3 (N1406, N1399, N91, N334);
nand NAND3 (N1407, N1394, N886, N1308);
buf BUF1 (N1408, N1400);
or OR4 (N1409, N1372, N1396, N1058, N825);
nand NAND3 (N1410, N1408, N1176, N1029);
nor NOR2 (N1411, N1393, N1311);
buf BUF1 (N1412, N1411);
and AND2 (N1413, N1404, N721);
nand NAND2 (N1414, N1397, N649);
nor NOR2 (N1415, N1406, N1077);
buf BUF1 (N1416, N1414);
nor NOR2 (N1417, N1407, N410);
nand NAND2 (N1418, N1401, N1308);
nor NOR2 (N1419, N1409, N839);
or OR2 (N1420, N1412, N1218);
and AND2 (N1421, N1420, N502);
xor XOR2 (N1422, N1419, N535);
nor NOR4 (N1423, N1413, N1123, N309, N164);
nand NAND4 (N1424, N1403, N764, N415, N181);
nor NOR2 (N1425, N1421, N479);
nor NOR3 (N1426, N1417, N812, N194);
buf BUF1 (N1427, N1416);
xor XOR2 (N1428, N1422, N116);
nand NAND2 (N1429, N1418, N770);
not NOT1 (N1430, N1423);
nand NAND4 (N1431, N1426, N700, N1404, N1005);
xor XOR2 (N1432, N1427, N490);
nor NOR4 (N1433, N1428, N1077, N979, N421);
xor XOR2 (N1434, N1430, N1361);
and AND4 (N1435, N1415, N358, N1189, N359);
nor NOR4 (N1436, N1433, N1053, N722, N239);
or OR3 (N1437, N1405, N1035, N501);
and AND4 (N1438, N1436, N1287, N861, N1009);
xor XOR2 (N1439, N1424, N779);
nor NOR3 (N1440, N1425, N1197, N888);
buf BUF1 (N1441, N1410);
xor XOR2 (N1442, N1434, N943);
not NOT1 (N1443, N1442);
nor NOR4 (N1444, N1431, N1029, N185, N1097);
nand NAND3 (N1445, N1432, N1063, N822);
nor NOR2 (N1446, N1440, N985);
nand NAND4 (N1447, N1429, N214, N945, N253);
xor XOR2 (N1448, N1447, N1183);
buf BUF1 (N1449, N1446);
buf BUF1 (N1450, N1439);
nand NAND3 (N1451, N1435, N1018, N592);
buf BUF1 (N1452, N1450);
not NOT1 (N1453, N1441);
nor NOR3 (N1454, N1449, N352, N487);
nor NOR3 (N1455, N1438, N1014, N629);
xor XOR2 (N1456, N1445, N17);
xor XOR2 (N1457, N1453, N918);
and AND3 (N1458, N1452, N946, N244);
nor NOR2 (N1459, N1448, N1271);
not NOT1 (N1460, N1454);
and AND3 (N1461, N1451, N1027, N828);
and AND3 (N1462, N1443, N210, N682);
xor XOR2 (N1463, N1437, N116);
buf BUF1 (N1464, N1462);
nand NAND3 (N1465, N1460, N270, N896);
and AND2 (N1466, N1465, N548);
buf BUF1 (N1467, N1464);
buf BUF1 (N1468, N1461);
not NOT1 (N1469, N1463);
not NOT1 (N1470, N1457);
and AND2 (N1471, N1456, N104);
nor NOR3 (N1472, N1467, N1049, N1458);
nor NOR3 (N1473, N627, N1238, N167);
nor NOR4 (N1474, N1444, N513, N23, N270);
nor NOR3 (N1475, N1471, N1106, N622);
nand NAND3 (N1476, N1459, N582, N1013);
buf BUF1 (N1477, N1472);
and AND2 (N1478, N1468, N942);
and AND4 (N1479, N1470, N672, N121, N591);
or OR3 (N1480, N1477, N1388, N461);
nor NOR4 (N1481, N1479, N145, N1170, N1161);
xor XOR2 (N1482, N1466, N459);
xor XOR2 (N1483, N1469, N498);
nand NAND4 (N1484, N1455, N891, N909, N70);
xor XOR2 (N1485, N1474, N1027);
buf BUF1 (N1486, N1473);
nor NOR3 (N1487, N1486, N504, N942);
or OR4 (N1488, N1476, N774, N414, N175);
nand NAND3 (N1489, N1481, N1336, N1125);
or OR3 (N1490, N1487, N970, N1399);
buf BUF1 (N1491, N1475);
not NOT1 (N1492, N1491);
and AND2 (N1493, N1490, N354);
nor NOR4 (N1494, N1478, N1331, N995, N375);
buf BUF1 (N1495, N1488);
or OR2 (N1496, N1495, N1379);
and AND4 (N1497, N1482, N1027, N1215, N1323);
or OR2 (N1498, N1480, N1369);
or OR2 (N1499, N1492, N718);
or OR4 (N1500, N1498, N372, N1471, N72);
not NOT1 (N1501, N1494);
nand NAND4 (N1502, N1493, N1124, N946, N1022);
nor NOR2 (N1503, N1499, N652);
and AND4 (N1504, N1503, N1195, N532, N795);
not NOT1 (N1505, N1485);
buf BUF1 (N1506, N1496);
xor XOR2 (N1507, N1484, N4);
buf BUF1 (N1508, N1504);
nand NAND3 (N1509, N1501, N817, N814);
nand NAND4 (N1510, N1497, N1219, N433, N768);
buf BUF1 (N1511, N1507);
nand NAND4 (N1512, N1483, N869, N434, N692);
nand NAND4 (N1513, N1506, N638, N949, N976);
nor NOR4 (N1514, N1510, N1230, N321, N1465);
or OR2 (N1515, N1505, N492);
buf BUF1 (N1516, N1508);
and AND3 (N1517, N1515, N1483, N568);
xor XOR2 (N1518, N1502, N1208);
nor NOR4 (N1519, N1511, N492, N428, N429);
nor NOR2 (N1520, N1512, N664);
xor XOR2 (N1521, N1520, N421);
not NOT1 (N1522, N1489);
nor NOR2 (N1523, N1518, N1510);
nor NOR3 (N1524, N1500, N761, N1285);
xor XOR2 (N1525, N1516, N1180);
nand NAND2 (N1526, N1525, N937);
nor NOR3 (N1527, N1517, N1039, N332);
and AND2 (N1528, N1527, N345);
nor NOR4 (N1529, N1522, N758, N445, N1208);
nand NAND3 (N1530, N1524, N902, N972);
and AND3 (N1531, N1528, N737, N563);
and AND3 (N1532, N1526, N170, N4);
nor NOR3 (N1533, N1531, N1231, N1011);
xor XOR2 (N1534, N1514, N888);
buf BUF1 (N1535, N1532);
nor NOR3 (N1536, N1529, N840, N565);
buf BUF1 (N1537, N1534);
nor NOR3 (N1538, N1537, N767, N374);
buf BUF1 (N1539, N1521);
nand NAND4 (N1540, N1536, N974, N256, N479);
nor NOR2 (N1541, N1533, N273);
or OR3 (N1542, N1530, N2, N1310);
nand NAND3 (N1543, N1509, N709, N249);
nor NOR2 (N1544, N1513, N1467);
and AND3 (N1545, N1539, N183, N6);
nand NAND4 (N1546, N1545, N1185, N1468, N1075);
nand NAND2 (N1547, N1546, N1453);
xor XOR2 (N1548, N1543, N5);
or OR4 (N1549, N1542, N1518, N24, N100);
xor XOR2 (N1550, N1548, N121);
nor NOR3 (N1551, N1547, N287, N355);
buf BUF1 (N1552, N1544);
nor NOR4 (N1553, N1551, N1121, N14, N953);
nor NOR3 (N1554, N1552, N784, N683);
buf BUF1 (N1555, N1540);
not NOT1 (N1556, N1541);
xor XOR2 (N1557, N1550, N195);
or OR3 (N1558, N1538, N616, N724);
and AND4 (N1559, N1556, N6, N362, N320);
or OR4 (N1560, N1557, N1340, N551, N718);
nand NAND2 (N1561, N1560, N1385);
xor XOR2 (N1562, N1554, N1074);
nand NAND2 (N1563, N1535, N1230);
xor XOR2 (N1564, N1559, N464);
or OR2 (N1565, N1561, N775);
nor NOR4 (N1566, N1558, N999, N1494, N785);
not NOT1 (N1567, N1523);
not NOT1 (N1568, N1564);
xor XOR2 (N1569, N1566, N1100);
buf BUF1 (N1570, N1569);
xor XOR2 (N1571, N1553, N1324);
nor NOR2 (N1572, N1555, N749);
xor XOR2 (N1573, N1563, N697);
buf BUF1 (N1574, N1572);
xor XOR2 (N1575, N1573, N1303);
nor NOR2 (N1576, N1519, N1130);
and AND3 (N1577, N1565, N14, N289);
nor NOR3 (N1578, N1574, N858, N1285);
nand NAND3 (N1579, N1549, N1187, N608);
nand NAND4 (N1580, N1568, N514, N298, N673);
or OR2 (N1581, N1579, N658);
buf BUF1 (N1582, N1567);
or OR2 (N1583, N1581, N94);
or OR3 (N1584, N1575, N914, N1354);
not NOT1 (N1585, N1578);
not NOT1 (N1586, N1583);
not NOT1 (N1587, N1580);
or OR2 (N1588, N1585, N521);
buf BUF1 (N1589, N1584);
or OR3 (N1590, N1577, N869, N1251);
and AND3 (N1591, N1588, N602, N292);
or OR3 (N1592, N1590, N1302, N639);
and AND4 (N1593, N1562, N847, N812, N796);
buf BUF1 (N1594, N1592);
buf BUF1 (N1595, N1576);
nand NAND2 (N1596, N1591, N741);
xor XOR2 (N1597, N1596, N408);
nor NOR2 (N1598, N1593, N236);
nor NOR4 (N1599, N1598, N1510, N317, N993);
and AND3 (N1600, N1595, N56, N880);
or OR2 (N1601, N1594, N202);
xor XOR2 (N1602, N1582, N1171);
xor XOR2 (N1603, N1602, N472);
and AND4 (N1604, N1600, N1364, N1081, N208);
nand NAND4 (N1605, N1589, N1067, N330, N486);
nand NAND3 (N1606, N1603, N770, N1156);
xor XOR2 (N1607, N1586, N1058);
buf BUF1 (N1608, N1606);
xor XOR2 (N1609, N1605, N970);
buf BUF1 (N1610, N1571);
not NOT1 (N1611, N1599);
not NOT1 (N1612, N1610);
and AND2 (N1613, N1587, N734);
and AND4 (N1614, N1613, N106, N1089, N1192);
nand NAND4 (N1615, N1607, N272, N815, N848);
or OR2 (N1616, N1612, N1383);
not NOT1 (N1617, N1614);
nand NAND3 (N1618, N1601, N298, N926);
nor NOR2 (N1619, N1597, N586);
not NOT1 (N1620, N1616);
xor XOR2 (N1621, N1608, N13);
and AND2 (N1622, N1604, N1250);
nand NAND3 (N1623, N1609, N1267, N1150);
xor XOR2 (N1624, N1621, N798);
not NOT1 (N1625, N1611);
and AND2 (N1626, N1618, N400);
buf BUF1 (N1627, N1620);
nand NAND2 (N1628, N1570, N1021);
nand NAND2 (N1629, N1622, N344);
nand NAND4 (N1630, N1623, N1392, N283, N103);
buf BUF1 (N1631, N1625);
and AND3 (N1632, N1630, N1366, N1431);
and AND4 (N1633, N1617, N231, N394, N1534);
nand NAND2 (N1634, N1629, N1273);
nand NAND3 (N1635, N1632, N451, N892);
or OR3 (N1636, N1627, N1315, N757);
nand NAND4 (N1637, N1633, N928, N1427, N1031);
xor XOR2 (N1638, N1634, N928);
xor XOR2 (N1639, N1637, N1145);
or OR4 (N1640, N1624, N1634, N865, N1412);
xor XOR2 (N1641, N1640, N810);
or OR3 (N1642, N1641, N410, N1357);
not NOT1 (N1643, N1638);
nor NOR4 (N1644, N1636, N341, N123, N965);
not NOT1 (N1645, N1639);
xor XOR2 (N1646, N1615, N1606);
nand NAND2 (N1647, N1626, N1088);
and AND2 (N1648, N1642, N1522);
xor XOR2 (N1649, N1643, N1337);
not NOT1 (N1650, N1647);
and AND4 (N1651, N1650, N898, N152, N237);
not NOT1 (N1652, N1635);
buf BUF1 (N1653, N1652);
or OR2 (N1654, N1651, N552);
not NOT1 (N1655, N1619);
and AND3 (N1656, N1631, N431, N1600);
or OR2 (N1657, N1655, N1094);
and AND3 (N1658, N1656, N148, N442);
and AND2 (N1659, N1628, N1065);
xor XOR2 (N1660, N1644, N581);
not NOT1 (N1661, N1649);
nand NAND2 (N1662, N1657, N578);
xor XOR2 (N1663, N1662, N43);
buf BUF1 (N1664, N1654);
nand NAND3 (N1665, N1659, N1420, N589);
not NOT1 (N1666, N1661);
buf BUF1 (N1667, N1648);
buf BUF1 (N1668, N1645);
or OR2 (N1669, N1665, N598);
nor NOR3 (N1670, N1660, N1462, N810);
nand NAND4 (N1671, N1664, N1019, N1302, N1363);
not NOT1 (N1672, N1668);
and AND2 (N1673, N1663, N746);
buf BUF1 (N1674, N1673);
nand NAND2 (N1675, N1671, N1054);
or OR3 (N1676, N1658, N303, N426);
xor XOR2 (N1677, N1674, N1174);
not NOT1 (N1678, N1666);
nor NOR4 (N1679, N1669, N813, N4, N325);
nor NOR4 (N1680, N1646, N686, N507, N805);
buf BUF1 (N1681, N1653);
not NOT1 (N1682, N1678);
xor XOR2 (N1683, N1679, N1441);
nor NOR2 (N1684, N1675, N334);
buf BUF1 (N1685, N1677);
or OR4 (N1686, N1667, N1163, N1543, N1493);
and AND2 (N1687, N1686, N1509);
and AND2 (N1688, N1683, N1379);
nor NOR4 (N1689, N1680, N587, N486, N269);
nand NAND2 (N1690, N1682, N889);
and AND4 (N1691, N1681, N1100, N242, N253);
nor NOR2 (N1692, N1691, N975);
or OR2 (N1693, N1689, N876);
nor NOR4 (N1694, N1672, N179, N1393, N1575);
and AND2 (N1695, N1693, N438);
or OR2 (N1696, N1690, N846);
or OR4 (N1697, N1670, N1581, N729, N1531);
buf BUF1 (N1698, N1696);
nand NAND3 (N1699, N1695, N947, N1489);
nand NAND4 (N1700, N1699, N230, N578, N722);
nand NAND3 (N1701, N1676, N40, N1267);
and AND4 (N1702, N1685, N705, N1120, N26);
nand NAND2 (N1703, N1688, N510);
nand NAND4 (N1704, N1702, N145, N1613, N952);
not NOT1 (N1705, N1694);
not NOT1 (N1706, N1705);
buf BUF1 (N1707, N1706);
buf BUF1 (N1708, N1703);
nor NOR4 (N1709, N1700, N1675, N253, N881);
nor NOR3 (N1710, N1708, N248, N1504);
or OR2 (N1711, N1710, N216);
buf BUF1 (N1712, N1692);
and AND3 (N1713, N1697, N1626, N1640);
and AND3 (N1714, N1713, N748, N145);
nand NAND2 (N1715, N1711, N1661);
and AND3 (N1716, N1715, N75, N705);
xor XOR2 (N1717, N1701, N89);
nand NAND4 (N1718, N1717, N1473, N347, N1247);
nor NOR4 (N1719, N1709, N699, N696, N1315);
buf BUF1 (N1720, N1687);
xor XOR2 (N1721, N1714, N1274);
and AND3 (N1722, N1718, N1694, N920);
xor XOR2 (N1723, N1698, N185);
and AND3 (N1724, N1720, N1292, N127);
not NOT1 (N1725, N1719);
nand NAND2 (N1726, N1725, N1366);
xor XOR2 (N1727, N1684, N680);
buf BUF1 (N1728, N1704);
and AND3 (N1729, N1721, N1529, N401);
nand NAND4 (N1730, N1728, N1165, N1324, N65);
buf BUF1 (N1731, N1707);
or OR3 (N1732, N1722, N1402, N1059);
or OR3 (N1733, N1729, N1651, N608);
or OR4 (N1734, N1716, N893, N371, N886);
and AND2 (N1735, N1727, N842);
nor NOR2 (N1736, N1724, N1637);
or OR3 (N1737, N1730, N150, N175);
not NOT1 (N1738, N1732);
not NOT1 (N1739, N1712);
not NOT1 (N1740, N1734);
buf BUF1 (N1741, N1739);
nand NAND3 (N1742, N1726, N1558, N549);
buf BUF1 (N1743, N1736);
buf BUF1 (N1744, N1735);
and AND3 (N1745, N1737, N1545, N1429);
xor XOR2 (N1746, N1723, N636);
not NOT1 (N1747, N1746);
nor NOR3 (N1748, N1747, N25, N914);
or OR2 (N1749, N1731, N891);
not NOT1 (N1750, N1740);
nand NAND4 (N1751, N1749, N1202, N1616, N161);
or OR2 (N1752, N1742, N1557);
nand NAND4 (N1753, N1751, N70, N1033, N532);
not NOT1 (N1754, N1752);
buf BUF1 (N1755, N1741);
buf BUF1 (N1756, N1748);
nand NAND4 (N1757, N1753, N982, N827, N1723);
nand NAND2 (N1758, N1743, N324);
nor NOR4 (N1759, N1758, N220, N686, N502);
buf BUF1 (N1760, N1744);
not NOT1 (N1761, N1750);
not NOT1 (N1762, N1759);
and AND3 (N1763, N1745, N1177, N760);
xor XOR2 (N1764, N1733, N783);
or OR3 (N1765, N1756, N1536, N19);
xor XOR2 (N1766, N1763, N830);
xor XOR2 (N1767, N1757, N381);
or OR3 (N1768, N1738, N1140, N1699);
buf BUF1 (N1769, N1760);
buf BUF1 (N1770, N1765);
or OR3 (N1771, N1769, N589, N146);
nor NOR4 (N1772, N1761, N540, N1277, N618);
xor XOR2 (N1773, N1764, N1702);
nor NOR4 (N1774, N1768, N1516, N1332, N1751);
buf BUF1 (N1775, N1754);
and AND4 (N1776, N1762, N774, N508, N1001);
nor NOR2 (N1777, N1774, N1140);
nand NAND3 (N1778, N1777, N1623, N385);
nand NAND2 (N1779, N1755, N647);
not NOT1 (N1780, N1770);
nor NOR2 (N1781, N1775, N1500);
or OR4 (N1782, N1780, N737, N1627, N127);
xor XOR2 (N1783, N1773, N908);
not NOT1 (N1784, N1771);
buf BUF1 (N1785, N1766);
nand NAND2 (N1786, N1784, N227);
buf BUF1 (N1787, N1781);
not NOT1 (N1788, N1783);
nand NAND3 (N1789, N1778, N1491, N83);
not NOT1 (N1790, N1788);
xor XOR2 (N1791, N1787, N1077);
buf BUF1 (N1792, N1772);
not NOT1 (N1793, N1779);
buf BUF1 (N1794, N1792);
not NOT1 (N1795, N1767);
nand NAND3 (N1796, N1786, N1764, N798);
not NOT1 (N1797, N1796);
buf BUF1 (N1798, N1794);
or OR2 (N1799, N1785, N1068);
nand NAND2 (N1800, N1776, N325);
or OR2 (N1801, N1789, N1152);
nor NOR3 (N1802, N1801, N321, N166);
buf BUF1 (N1803, N1797);
nor NOR3 (N1804, N1782, N934, N1401);
or OR4 (N1805, N1798, N1394, N19, N868);
nand NAND2 (N1806, N1802, N578);
nand NAND4 (N1807, N1800, N1373, N1668, N782);
nor NOR2 (N1808, N1803, N811);
nand NAND4 (N1809, N1799, N1035, N384, N847);
buf BUF1 (N1810, N1804);
and AND3 (N1811, N1806, N1140, N1770);
not NOT1 (N1812, N1809);
xor XOR2 (N1813, N1805, N1346);
or OR4 (N1814, N1813, N1365, N491, N341);
nand NAND3 (N1815, N1791, N6, N834);
not NOT1 (N1816, N1790);
or OR4 (N1817, N1814, N1136, N226, N743);
not NOT1 (N1818, N1807);
not NOT1 (N1819, N1816);
buf BUF1 (N1820, N1795);
not NOT1 (N1821, N1808);
nand NAND2 (N1822, N1811, N47);
nand NAND4 (N1823, N1810, N369, N1302, N402);
or OR3 (N1824, N1821, N871, N508);
or OR4 (N1825, N1817, N903, N660, N807);
buf BUF1 (N1826, N1819);
not NOT1 (N1827, N1818);
buf BUF1 (N1828, N1812);
or OR2 (N1829, N1825, N849);
xor XOR2 (N1830, N1823, N1557);
nor NOR2 (N1831, N1829, N763);
or OR2 (N1832, N1827, N1366);
or OR4 (N1833, N1820, N1180, N3, N778);
buf BUF1 (N1834, N1828);
and AND2 (N1835, N1832, N313);
and AND4 (N1836, N1824, N314, N1118, N1595);
xor XOR2 (N1837, N1793, N150);
nor NOR4 (N1838, N1833, N517, N1099, N1730);
or OR3 (N1839, N1822, N1575, N138);
buf BUF1 (N1840, N1835);
nor NOR2 (N1841, N1831, N1332);
not NOT1 (N1842, N1838);
buf BUF1 (N1843, N1842);
or OR2 (N1844, N1843, N1276);
buf BUF1 (N1845, N1840);
nor NOR4 (N1846, N1830, N277, N1644, N549);
or OR3 (N1847, N1845, N506, N222);
nor NOR4 (N1848, N1841, N7, N1707, N1059);
and AND2 (N1849, N1847, N311);
nor NOR2 (N1850, N1848, N1402);
not NOT1 (N1851, N1815);
and AND2 (N1852, N1826, N236);
or OR2 (N1853, N1850, N1600);
nor NOR3 (N1854, N1836, N937, N1135);
not NOT1 (N1855, N1852);
nor NOR2 (N1856, N1834, N1798);
and AND3 (N1857, N1846, N1332, N580);
not NOT1 (N1858, N1857);
buf BUF1 (N1859, N1853);
buf BUF1 (N1860, N1856);
xor XOR2 (N1861, N1844, N542);
xor XOR2 (N1862, N1855, N1115);
xor XOR2 (N1863, N1854, N1242);
and AND3 (N1864, N1839, N110, N278);
not NOT1 (N1865, N1837);
nor NOR2 (N1866, N1861, N1775);
nand NAND4 (N1867, N1860, N418, N105, N1601);
and AND4 (N1868, N1851, N124, N1639, N934);
or OR3 (N1869, N1863, N550, N393);
xor XOR2 (N1870, N1862, N787);
nand NAND3 (N1871, N1858, N506, N744);
and AND2 (N1872, N1849, N217);
buf BUF1 (N1873, N1867);
or OR2 (N1874, N1864, N1506);
xor XOR2 (N1875, N1859, N282);
or OR3 (N1876, N1869, N1705, N56);
not NOT1 (N1877, N1868);
and AND3 (N1878, N1865, N1179, N1502);
not NOT1 (N1879, N1872);
xor XOR2 (N1880, N1879, N1855);
nand NAND4 (N1881, N1866, N87, N64, N995);
xor XOR2 (N1882, N1878, N451);
buf BUF1 (N1883, N1880);
buf BUF1 (N1884, N1881);
xor XOR2 (N1885, N1884, N1133);
xor XOR2 (N1886, N1874, N853);
or OR3 (N1887, N1885, N108, N955);
buf BUF1 (N1888, N1887);
buf BUF1 (N1889, N1877);
nand NAND4 (N1890, N1882, N1127, N442, N767);
nand NAND4 (N1891, N1886, N636, N971, N550);
xor XOR2 (N1892, N1890, N103);
or OR3 (N1893, N1883, N1159, N180);
nor NOR4 (N1894, N1873, N1299, N968, N1737);
not NOT1 (N1895, N1875);
or OR2 (N1896, N1894, N225);
nand NAND2 (N1897, N1889, N1626);
not NOT1 (N1898, N1897);
or OR3 (N1899, N1888, N672, N1122);
or OR3 (N1900, N1899, N211, N127);
buf BUF1 (N1901, N1892);
nor NOR2 (N1902, N1895, N102);
nor NOR4 (N1903, N1891, N53, N1164, N878);
nand NAND4 (N1904, N1900, N1848, N1050, N354);
xor XOR2 (N1905, N1904, N1629);
xor XOR2 (N1906, N1896, N1537);
or OR4 (N1907, N1876, N104, N1176, N950);
or OR2 (N1908, N1906, N1784);
and AND3 (N1909, N1903, N897, N319);
or OR4 (N1910, N1907, N606, N263, N320);
buf BUF1 (N1911, N1871);
buf BUF1 (N1912, N1905);
xor XOR2 (N1913, N1893, N794);
not NOT1 (N1914, N1912);
nor NOR4 (N1915, N1870, N1589, N1092, N1794);
or OR2 (N1916, N1902, N1394);
not NOT1 (N1917, N1909);
xor XOR2 (N1918, N1913, N1780);
buf BUF1 (N1919, N1916);
nand NAND4 (N1920, N1898, N1803, N427, N168);
buf BUF1 (N1921, N1910);
buf BUF1 (N1922, N1917);
buf BUF1 (N1923, N1901);
and AND2 (N1924, N1918, N869);
not NOT1 (N1925, N1919);
and AND4 (N1926, N1925, N1697, N384, N453);
and AND4 (N1927, N1915, N1835, N665, N690);
and AND4 (N1928, N1924, N1369, N1366, N319);
not NOT1 (N1929, N1920);
xor XOR2 (N1930, N1911, N239);
not NOT1 (N1931, N1908);
and AND2 (N1932, N1927, N83);
not NOT1 (N1933, N1932);
nand NAND3 (N1934, N1923, N916, N1781);
and AND2 (N1935, N1921, N577);
nor NOR4 (N1936, N1935, N1707, N1580, N291);
buf BUF1 (N1937, N1922);
nand NAND2 (N1938, N1926, N1525);
or OR4 (N1939, N1914, N505, N140, N945);
and AND4 (N1940, N1933, N717, N1116, N1020);
buf BUF1 (N1941, N1936);
not NOT1 (N1942, N1929);
not NOT1 (N1943, N1938);
nand NAND4 (N1944, N1943, N1180, N1722, N1689);
and AND4 (N1945, N1934, N274, N99, N700);
or OR2 (N1946, N1930, N1736);
buf BUF1 (N1947, N1939);
nor NOR4 (N1948, N1931, N1260, N877, N964);
and AND2 (N1949, N1947, N1809);
and AND4 (N1950, N1937, N1315, N559, N1706);
and AND4 (N1951, N1944, N1654, N368, N1036);
and AND4 (N1952, N1940, N1940, N1610, N323);
nand NAND2 (N1953, N1948, N1897);
xor XOR2 (N1954, N1945, N1899);
not NOT1 (N1955, N1950);
nor NOR2 (N1956, N1949, N810);
not NOT1 (N1957, N1946);
nand NAND4 (N1958, N1941, N1679, N1230, N1253);
xor XOR2 (N1959, N1951, N377);
nor NOR3 (N1960, N1952, N107, N251);
nor NOR3 (N1961, N1955, N121, N339);
xor XOR2 (N1962, N1960, N518);
or OR2 (N1963, N1956, N1598);
xor XOR2 (N1964, N1954, N344);
not NOT1 (N1965, N1942);
not NOT1 (N1966, N1928);
xor XOR2 (N1967, N1963, N1097);
or OR3 (N1968, N1961, N1040, N679);
nand NAND3 (N1969, N1965, N1436, N1788);
nand NAND2 (N1970, N1958, N439);
and AND2 (N1971, N1969, N1825);
or OR2 (N1972, N1968, N1590);
or OR4 (N1973, N1957, N429, N1267, N1668);
nand NAND3 (N1974, N1973, N1709, N1106);
buf BUF1 (N1975, N1964);
nor NOR4 (N1976, N1970, N816, N220, N1918);
and AND3 (N1977, N1976, N765, N539);
buf BUF1 (N1978, N1967);
buf BUF1 (N1979, N1977);
or OR4 (N1980, N1974, N814, N137, N1250);
not NOT1 (N1981, N1971);
or OR4 (N1982, N1981, N914, N1351, N1972);
and AND4 (N1983, N1192, N1470, N1139, N285);
nor NOR2 (N1984, N1975, N78);
xor XOR2 (N1985, N1982, N781);
buf BUF1 (N1986, N1953);
not NOT1 (N1987, N1962);
buf BUF1 (N1988, N1985);
and AND2 (N1989, N1979, N779);
buf BUF1 (N1990, N1966);
and AND2 (N1991, N1990, N1432);
and AND3 (N1992, N1991, N1840, N123);
xor XOR2 (N1993, N1983, N1779);
nand NAND4 (N1994, N1978, N1788, N1915, N1173);
xor XOR2 (N1995, N1992, N1109);
not NOT1 (N1996, N1959);
or OR4 (N1997, N1994, N858, N1133, N1109);
or OR4 (N1998, N1980, N926, N798, N787);
not NOT1 (N1999, N1986);
and AND3 (N2000, N1987, N59, N194);
nand NAND4 (N2001, N1995, N411, N282, N1445);
nand NAND2 (N2002, N1989, N742);
nor NOR4 (N2003, N1993, N1565, N314, N1330);
nor NOR4 (N2004, N2003, N151, N974, N379);
and AND3 (N2005, N1998, N526, N1173);
buf BUF1 (N2006, N2001);
xor XOR2 (N2007, N2000, N1461);
and AND3 (N2008, N1999, N222, N836);
buf BUF1 (N2009, N1997);
and AND2 (N2010, N2005, N493);
or OR4 (N2011, N2004, N1225, N1231, N1293);
or OR4 (N2012, N1996, N26, N1611, N724);
not NOT1 (N2013, N1988);
nor NOR3 (N2014, N2007, N1440, N788);
buf BUF1 (N2015, N2012);
or OR2 (N2016, N2013, N1803);
or OR2 (N2017, N2011, N248);
buf BUF1 (N2018, N2014);
and AND2 (N2019, N2018, N1629);
not NOT1 (N2020, N2010);
not NOT1 (N2021, N2008);
nor NOR4 (N2022, N2009, N1164, N1565, N1911);
buf BUF1 (N2023, N2006);
or OR4 (N2024, N2015, N1809, N1018, N933);
xor XOR2 (N2025, N2024, N876);
nor NOR3 (N2026, N2023, N240, N38);
not NOT1 (N2027, N2017);
nor NOR2 (N2028, N2016, N387);
or OR2 (N2029, N2026, N1483);
or OR2 (N2030, N2019, N764);
or OR2 (N2031, N2028, N432);
nand NAND4 (N2032, N2020, N998, N1028, N2021);
nand NAND2 (N2033, N633, N1321);
and AND2 (N2034, N2029, N608);
buf BUF1 (N2035, N2022);
or OR2 (N2036, N2033, N953);
buf BUF1 (N2037, N2030);
or OR3 (N2038, N2031, N1691, N1642);
nand NAND3 (N2039, N2025, N1373, N954);
and AND3 (N2040, N2035, N1576, N1653);
nand NAND3 (N2041, N2027, N1932, N1576);
not NOT1 (N2042, N2037);
xor XOR2 (N2043, N1984, N1536);
not NOT1 (N2044, N2039);
buf BUF1 (N2045, N2041);
not NOT1 (N2046, N2040);
nor NOR4 (N2047, N2042, N834, N989, N1701);
xor XOR2 (N2048, N2034, N624);
xor XOR2 (N2049, N2048, N546);
nand NAND4 (N2050, N2032, N1228, N1422, N776);
buf BUF1 (N2051, N2049);
xor XOR2 (N2052, N2046, N1703);
nor NOR2 (N2053, N2038, N555);
buf BUF1 (N2054, N2052);
xor XOR2 (N2055, N2002, N1566);
nor NOR4 (N2056, N2043, N75, N1073, N943);
and AND4 (N2057, N2051, N264, N561, N2008);
not NOT1 (N2058, N2055);
nand NAND2 (N2059, N2044, N550);
or OR3 (N2060, N2050, N395, N1891);
or OR4 (N2061, N2057, N628, N1151, N1812);
nor NOR3 (N2062, N2061, N1247, N2018);
nand NAND2 (N2063, N2054, N601);
xor XOR2 (N2064, N2036, N1915);
xor XOR2 (N2065, N2045, N2036);
xor XOR2 (N2066, N2063, N1261);
or OR3 (N2067, N2059, N826, N1183);
or OR2 (N2068, N2066, N45);
and AND2 (N2069, N2067, N367);
and AND2 (N2070, N2058, N188);
buf BUF1 (N2071, N2064);
or OR4 (N2072, N2071, N1631, N1577, N461);
or OR4 (N2073, N2060, N1189, N2064, N656);
nor NOR3 (N2074, N2065, N30, N640);
xor XOR2 (N2075, N2073, N1485);
not NOT1 (N2076, N2075);
nand NAND2 (N2077, N2070, N146);
buf BUF1 (N2078, N2072);
nor NOR4 (N2079, N2074, N844, N1813, N304);
nor NOR2 (N2080, N2062, N898);
nor NOR3 (N2081, N2080, N1032, N325);
and AND3 (N2082, N2079, N1892, N1355);
and AND3 (N2083, N2078, N764, N1990);
buf BUF1 (N2084, N2081);
not NOT1 (N2085, N2083);
not NOT1 (N2086, N2053);
buf BUF1 (N2087, N2085);
xor XOR2 (N2088, N2087, N1550);
buf BUF1 (N2089, N2088);
and AND2 (N2090, N2089, N1384);
not NOT1 (N2091, N2069);
and AND4 (N2092, N2056, N2006, N727, N41);
nor NOR4 (N2093, N2068, N1600, N2047, N589);
nand NAND3 (N2094, N407, N1822, N1575);
not NOT1 (N2095, N2082);
xor XOR2 (N2096, N2090, N1178);
nor NOR4 (N2097, N2096, N1476, N352, N446);
xor XOR2 (N2098, N2093, N1945);
not NOT1 (N2099, N2086);
xor XOR2 (N2100, N2099, N1308);
buf BUF1 (N2101, N2091);
xor XOR2 (N2102, N2076, N1833);
nor NOR2 (N2103, N2094, N327);
xor XOR2 (N2104, N2084, N322);
xor XOR2 (N2105, N2102, N495);
xor XOR2 (N2106, N2100, N599);
or OR2 (N2107, N2095, N1934);
or OR2 (N2108, N2107, N720);
not NOT1 (N2109, N2092);
xor XOR2 (N2110, N2108, N2073);
nand NAND4 (N2111, N2110, N1072, N639, N2004);
nand NAND4 (N2112, N2111, N280, N1683, N962);
not NOT1 (N2113, N2101);
nor NOR4 (N2114, N2103, N2015, N551, N2070);
buf BUF1 (N2115, N2077);
xor XOR2 (N2116, N2115, N88);
nor NOR4 (N2117, N2106, N1502, N1121, N1083);
or OR2 (N2118, N2109, N662);
or OR4 (N2119, N2098, N1348, N1713, N2043);
buf BUF1 (N2120, N2104);
buf BUF1 (N2121, N2114);
or OR2 (N2122, N2119, N1202);
and AND3 (N2123, N2122, N580, N533);
buf BUF1 (N2124, N2121);
and AND3 (N2125, N2118, N1923, N751);
buf BUF1 (N2126, N2120);
nor NOR2 (N2127, N2124, N970);
buf BUF1 (N2128, N2125);
nand NAND4 (N2129, N2127, N1502, N1860, N1502);
nand NAND2 (N2130, N2123, N1459);
not NOT1 (N2131, N2113);
or OR3 (N2132, N2117, N389, N2032);
xor XOR2 (N2133, N2126, N866);
nand NAND3 (N2134, N2112, N148, N130);
xor XOR2 (N2135, N2128, N483);
nor NOR4 (N2136, N2130, N1094, N1000, N2071);
xor XOR2 (N2137, N2129, N1489);
nand NAND2 (N2138, N2134, N1869);
buf BUF1 (N2139, N2135);
nor NOR4 (N2140, N2136, N704, N1717, N525);
xor XOR2 (N2141, N2137, N570);
buf BUF1 (N2142, N2141);
xor XOR2 (N2143, N2131, N1701);
not NOT1 (N2144, N2116);
xor XOR2 (N2145, N2132, N1270);
xor XOR2 (N2146, N2105, N791);
not NOT1 (N2147, N2138);
and AND4 (N2148, N2097, N1931, N160, N1786);
or OR2 (N2149, N2146, N732);
nand NAND3 (N2150, N2147, N1456, N1005);
buf BUF1 (N2151, N2145);
xor XOR2 (N2152, N2142, N939);
buf BUF1 (N2153, N2152);
nand NAND4 (N2154, N2140, N1682, N529, N1785);
or OR4 (N2155, N2144, N678, N712, N1263);
nand NAND3 (N2156, N2154, N1606, N2153);
and AND4 (N2157, N1282, N1523, N447, N1337);
xor XOR2 (N2158, N2148, N1212);
and AND4 (N2159, N2158, N1881, N1989, N1864);
nand NAND2 (N2160, N2157, N887);
and AND3 (N2161, N2159, N1803, N268);
and AND2 (N2162, N2139, N1867);
and AND3 (N2163, N2133, N447, N957);
not NOT1 (N2164, N2156);
buf BUF1 (N2165, N2161);
or OR3 (N2166, N2143, N437, N651);
xor XOR2 (N2167, N2149, N1596);
nand NAND4 (N2168, N2167, N584, N1205, N723);
and AND2 (N2169, N2150, N1331);
nor NOR2 (N2170, N2168, N2145);
not NOT1 (N2171, N2155);
not NOT1 (N2172, N2163);
not NOT1 (N2173, N2169);
nor NOR2 (N2174, N2162, N353);
nand NAND2 (N2175, N2166, N1838);
buf BUF1 (N2176, N2164);
or OR3 (N2177, N2170, N2017, N1387);
nor NOR2 (N2178, N2173, N291);
nand NAND3 (N2179, N2177, N1379, N1515);
xor XOR2 (N2180, N2176, N666);
nor NOR3 (N2181, N2172, N785, N1447);
nand NAND2 (N2182, N2171, N1422);
or OR3 (N2183, N2181, N1275, N1609);
or OR3 (N2184, N2175, N1017, N1692);
not NOT1 (N2185, N2184);
nor NOR2 (N2186, N2180, N1506);
buf BUF1 (N2187, N2186);
buf BUF1 (N2188, N2182);
nor NOR4 (N2189, N2188, N1868, N6, N318);
xor XOR2 (N2190, N2185, N1788);
not NOT1 (N2191, N2189);
nand NAND4 (N2192, N2178, N1194, N1254, N723);
nand NAND2 (N2193, N2151, N1499);
and AND4 (N2194, N2193, N1456, N1014, N1083);
nor NOR2 (N2195, N2183, N17);
not NOT1 (N2196, N2160);
buf BUF1 (N2197, N2179);
or OR3 (N2198, N2196, N666, N94);
xor XOR2 (N2199, N2187, N257);
xor XOR2 (N2200, N2190, N644);
and AND3 (N2201, N2198, N1420, N675);
or OR3 (N2202, N2194, N1377, N1917);
or OR3 (N2203, N2165, N868, N1767);
xor XOR2 (N2204, N2200, N966);
xor XOR2 (N2205, N2192, N1810);
xor XOR2 (N2206, N2203, N1853);
and AND2 (N2207, N2191, N913);
nor NOR3 (N2208, N2202, N1321, N1195);
buf BUF1 (N2209, N2208);
or OR3 (N2210, N2207, N1361, N562);
xor XOR2 (N2211, N2195, N2107);
or OR2 (N2212, N2206, N1833);
nor NOR2 (N2213, N2174, N1994);
nor NOR3 (N2214, N2197, N1215, N1967);
or OR4 (N2215, N2199, N798, N853, N1415);
buf BUF1 (N2216, N2210);
not NOT1 (N2217, N2211);
and AND2 (N2218, N2214, N99);
nand NAND3 (N2219, N2212, N1891, N695);
buf BUF1 (N2220, N2215);
buf BUF1 (N2221, N2216);
xor XOR2 (N2222, N2221, N1937);
and AND3 (N2223, N2205, N478, N840);
xor XOR2 (N2224, N2219, N1123);
not NOT1 (N2225, N2201);
nor NOR3 (N2226, N2220, N772, N1205);
xor XOR2 (N2227, N2222, N2003);
buf BUF1 (N2228, N2209);
nor NOR3 (N2229, N2226, N596, N38);
xor XOR2 (N2230, N2225, N1967);
buf BUF1 (N2231, N2204);
and AND4 (N2232, N2217, N1157, N1738, N634);
and AND3 (N2233, N2230, N503, N327);
not NOT1 (N2234, N2228);
not NOT1 (N2235, N2231);
or OR3 (N2236, N2223, N1939, N1735);
not NOT1 (N2237, N2218);
xor XOR2 (N2238, N2232, N336);
nand NAND2 (N2239, N2236, N1081);
and AND3 (N2240, N2234, N1221, N1241);
nor NOR2 (N2241, N2213, N1757);
xor XOR2 (N2242, N2238, N2137);
or OR4 (N2243, N2239, N1948, N299, N2138);
and AND4 (N2244, N2241, N2133, N172, N1843);
not NOT1 (N2245, N2240);
xor XOR2 (N2246, N2227, N1634);
nor NOR3 (N2247, N2246, N1090, N350);
or OR2 (N2248, N2229, N757);
nor NOR2 (N2249, N2247, N1144);
or OR3 (N2250, N2235, N1443, N1903);
not NOT1 (N2251, N2248);
and AND2 (N2252, N2233, N677);
nand NAND4 (N2253, N2252, N1563, N787, N668);
xor XOR2 (N2254, N2245, N350);
xor XOR2 (N2255, N2249, N2067);
or OR2 (N2256, N2242, N243);
xor XOR2 (N2257, N2237, N197);
and AND3 (N2258, N2250, N1223, N1004);
not NOT1 (N2259, N2255);
or OR2 (N2260, N2258, N2165);
not NOT1 (N2261, N2243);
nor NOR3 (N2262, N2224, N1931, N2170);
or OR3 (N2263, N2253, N940, N1442);
not NOT1 (N2264, N2259);
not NOT1 (N2265, N2254);
buf BUF1 (N2266, N2263);
and AND2 (N2267, N2265, N866);
buf BUF1 (N2268, N2244);
nor NOR4 (N2269, N2267, N611, N2140, N1116);
or OR4 (N2270, N2266, N2043, N929, N1857);
or OR2 (N2271, N2270, N89);
and AND4 (N2272, N2251, N958, N303, N595);
buf BUF1 (N2273, N2272);
not NOT1 (N2274, N2268);
or OR3 (N2275, N2274, N2192, N142);
nand NAND2 (N2276, N2264, N186);
not NOT1 (N2277, N2261);
buf BUF1 (N2278, N2260);
or OR4 (N2279, N2257, N1375, N959, N409);
and AND2 (N2280, N2271, N223);
or OR4 (N2281, N2277, N1123, N1964, N1552);
nand NAND3 (N2282, N2279, N497, N1034);
buf BUF1 (N2283, N2262);
nor NOR3 (N2284, N2275, N1620, N898);
and AND4 (N2285, N2282, N2032, N2071, N1272);
not NOT1 (N2286, N2281);
nor NOR2 (N2287, N2280, N1735);
nor NOR3 (N2288, N2278, N1062, N2026);
or OR2 (N2289, N2284, N654);
nor NOR3 (N2290, N2256, N1058, N1653);
and AND4 (N2291, N2286, N1969, N487, N97);
nand NAND4 (N2292, N2283, N2260, N1090, N673);
buf BUF1 (N2293, N2291);
or OR2 (N2294, N2276, N438);
nor NOR4 (N2295, N2288, N1678, N703, N1967);
nor NOR2 (N2296, N2293, N459);
xor XOR2 (N2297, N2292, N464);
or OR2 (N2298, N2269, N1423);
nand NAND4 (N2299, N2295, N2063, N1969, N2216);
buf BUF1 (N2300, N2273);
nand NAND2 (N2301, N2287, N1171);
nand NAND3 (N2302, N2294, N1875, N623);
buf BUF1 (N2303, N2296);
buf BUF1 (N2304, N2297);
buf BUF1 (N2305, N2300);
nor NOR2 (N2306, N2302, N1542);
buf BUF1 (N2307, N2303);
and AND3 (N2308, N2305, N2145, N1732);
nand NAND4 (N2309, N2304, N1626, N1163, N1721);
and AND2 (N2310, N2298, N289);
and AND2 (N2311, N2285, N1004);
xor XOR2 (N2312, N2301, N1747);
not NOT1 (N2313, N2309);
and AND2 (N2314, N2289, N459);
not NOT1 (N2315, N2307);
and AND3 (N2316, N2290, N2095, N332);
or OR2 (N2317, N2306, N2109);
xor XOR2 (N2318, N2299, N2087);
nand NAND2 (N2319, N2315, N1542);
or OR2 (N2320, N2310, N735);
nor NOR2 (N2321, N2318, N1708);
not NOT1 (N2322, N2321);
xor XOR2 (N2323, N2313, N849);
and AND3 (N2324, N2311, N1061, N998);
not NOT1 (N2325, N2314);
and AND2 (N2326, N2323, N1105);
or OR4 (N2327, N2317, N707, N210, N2000);
nand NAND3 (N2328, N2319, N1098, N1651);
xor XOR2 (N2329, N2308, N827);
nand NAND2 (N2330, N2316, N913);
xor XOR2 (N2331, N2328, N1768);
xor XOR2 (N2332, N2325, N2109);
or OR4 (N2333, N2330, N1338, N2170, N1696);
or OR2 (N2334, N2332, N1569);
and AND4 (N2335, N2312, N7, N1220, N1589);
nand NAND3 (N2336, N2329, N1339, N1910);
nand NAND2 (N2337, N2336, N2044);
nand NAND3 (N2338, N2337, N1048, N559);
and AND3 (N2339, N2338, N603, N1024);
and AND4 (N2340, N2327, N2167, N40, N2031);
or OR3 (N2341, N2326, N1406, N721);
and AND2 (N2342, N2334, N1577);
buf BUF1 (N2343, N2324);
xor XOR2 (N2344, N2331, N1345);
buf BUF1 (N2345, N2335);
not NOT1 (N2346, N2343);
nand NAND3 (N2347, N2344, N1622, N1809);
and AND3 (N2348, N2346, N2101, N1970);
not NOT1 (N2349, N2347);
xor XOR2 (N2350, N2322, N593);
nand NAND3 (N2351, N2320, N2283, N2319);
xor XOR2 (N2352, N2339, N67);
nor NOR4 (N2353, N2349, N1446, N591, N1353);
nor NOR4 (N2354, N2353, N2087, N2303, N2016);
nor NOR2 (N2355, N2354, N1380);
xor XOR2 (N2356, N2333, N1534);
nor NOR4 (N2357, N2341, N254, N1793, N860);
and AND3 (N2358, N2350, N2233, N1353);
or OR4 (N2359, N2340, N674, N753, N94);
nand NAND4 (N2360, N2359, N1119, N995, N1991);
nor NOR3 (N2361, N2357, N964, N1447);
xor XOR2 (N2362, N2361, N480);
buf BUF1 (N2363, N2345);
not NOT1 (N2364, N2351);
not NOT1 (N2365, N2348);
not NOT1 (N2366, N2358);
nor NOR4 (N2367, N2356, N900, N1784, N696);
and AND4 (N2368, N2352, N2190, N601, N2186);
or OR4 (N2369, N2362, N2046, N40, N556);
xor XOR2 (N2370, N2363, N1875);
or OR4 (N2371, N2370, N847, N1930, N809);
not NOT1 (N2372, N2368);
nand NAND3 (N2373, N2342, N2332, N197);
xor XOR2 (N2374, N2355, N1401);
xor XOR2 (N2375, N2367, N185);
nand NAND4 (N2376, N2371, N2087, N1876, N762);
buf BUF1 (N2377, N2372);
nor NOR2 (N2378, N2375, N1847);
buf BUF1 (N2379, N2365);
xor XOR2 (N2380, N2366, N1854);
nor NOR2 (N2381, N2377, N734);
nand NAND2 (N2382, N2379, N1817);
nor NOR3 (N2383, N2381, N145, N505);
not NOT1 (N2384, N2383);
nor NOR3 (N2385, N2374, N1842, N1224);
nor NOR2 (N2386, N2360, N2340);
or OR3 (N2387, N2373, N93, N1845);
or OR2 (N2388, N2384, N1976);
not NOT1 (N2389, N2387);
and AND3 (N2390, N2382, N682, N1399);
and AND4 (N2391, N2376, N1978, N643, N2251);
nor NOR2 (N2392, N2389, N809);
nand NAND3 (N2393, N2380, N725, N1724);
nor NOR3 (N2394, N2390, N2188, N259);
xor XOR2 (N2395, N2386, N623);
nor NOR4 (N2396, N2378, N1575, N1315, N1327);
or OR4 (N2397, N2396, N1792, N2119, N1275);
buf BUF1 (N2398, N2392);
nor NOR2 (N2399, N2397, N141);
and AND2 (N2400, N2385, N1633);
xor XOR2 (N2401, N2399, N1549);
buf BUF1 (N2402, N2394);
buf BUF1 (N2403, N2402);
not NOT1 (N2404, N2388);
not NOT1 (N2405, N2398);
buf BUF1 (N2406, N2393);
or OR3 (N2407, N2400, N396, N755);
nand NAND3 (N2408, N2364, N378, N2027);
or OR4 (N2409, N2404, N687, N1729, N58);
not NOT1 (N2410, N2409);
buf BUF1 (N2411, N2403);
and AND3 (N2412, N2410, N708, N275);
nand NAND4 (N2413, N2405, N1253, N1514, N1930);
and AND2 (N2414, N2413, N1162);
and AND2 (N2415, N2411, N1853);
and AND2 (N2416, N2395, N1380);
not NOT1 (N2417, N2414);
or OR2 (N2418, N2369, N1119);
xor XOR2 (N2419, N2406, N1244);
and AND2 (N2420, N2416, N2006);
not NOT1 (N2421, N2415);
not NOT1 (N2422, N2412);
nor NOR3 (N2423, N2407, N416, N826);
not NOT1 (N2424, N2422);
or OR3 (N2425, N2419, N35, N68);
nor NOR3 (N2426, N2418, N78, N2404);
and AND3 (N2427, N2391, N371, N485);
nand NAND4 (N2428, N2426, N510, N1139, N2349);
nor NOR2 (N2429, N2417, N157);
xor XOR2 (N2430, N2427, N971);
nand NAND2 (N2431, N2423, N10);
xor XOR2 (N2432, N2428, N376);
buf BUF1 (N2433, N2424);
xor XOR2 (N2434, N2401, N732);
nand NAND2 (N2435, N2434, N915);
nand NAND4 (N2436, N2430, N592, N1506, N773);
xor XOR2 (N2437, N2431, N268);
nand NAND4 (N2438, N2433, N1413, N1494, N447);
nand NAND3 (N2439, N2408, N1283, N1347);
buf BUF1 (N2440, N2436);
xor XOR2 (N2441, N2429, N1653);
not NOT1 (N2442, N2439);
nand NAND3 (N2443, N2440, N2143, N1907);
nand NAND4 (N2444, N2437, N580, N849, N2094);
nand NAND3 (N2445, N2442, N1199, N2204);
not NOT1 (N2446, N2445);
not NOT1 (N2447, N2443);
xor XOR2 (N2448, N2444, N720);
nand NAND2 (N2449, N2420, N1245);
and AND3 (N2450, N2441, N1411, N1231);
buf BUF1 (N2451, N2438);
nand NAND2 (N2452, N2432, N2438);
xor XOR2 (N2453, N2447, N2161);
or OR3 (N2454, N2451, N1708, N1551);
buf BUF1 (N2455, N2453);
nor NOR2 (N2456, N2450, N2417);
nor NOR4 (N2457, N2449, N1538, N1618, N2391);
or OR3 (N2458, N2425, N550, N2115);
or OR4 (N2459, N2456, N817, N1973, N1611);
or OR4 (N2460, N2457, N2217, N925, N1638);
or OR3 (N2461, N2460, N986, N1360);
not NOT1 (N2462, N2448);
not NOT1 (N2463, N2435);
buf BUF1 (N2464, N2461);
not NOT1 (N2465, N2463);
and AND4 (N2466, N2454, N55, N1884, N52);
xor XOR2 (N2467, N2465, N145);
and AND3 (N2468, N2467, N5, N742);
and AND2 (N2469, N2464, N1556);
or OR2 (N2470, N2446, N1756);
or OR4 (N2471, N2459, N585, N707, N1797);
and AND4 (N2472, N2469, N1903, N994, N2340);
not NOT1 (N2473, N2470);
buf BUF1 (N2474, N2462);
and AND3 (N2475, N2458, N352, N2236);
not NOT1 (N2476, N2472);
xor XOR2 (N2477, N2474, N970);
and AND2 (N2478, N2466, N335);
not NOT1 (N2479, N2455);
xor XOR2 (N2480, N2452, N1799);
xor XOR2 (N2481, N2468, N784);
nand NAND2 (N2482, N2473, N1958);
and AND3 (N2483, N2481, N1726, N255);
not NOT1 (N2484, N2480);
xor XOR2 (N2485, N2421, N758);
buf BUF1 (N2486, N2484);
nor NOR3 (N2487, N2477, N1691, N2146);
buf BUF1 (N2488, N2476);
nand NAND4 (N2489, N2471, N1712, N285, N1218);
xor XOR2 (N2490, N2489, N2129);
buf BUF1 (N2491, N2490);
and AND4 (N2492, N2488, N1675, N777, N193);
or OR3 (N2493, N2482, N1524, N1255);
not NOT1 (N2494, N2475);
and AND4 (N2495, N2479, N1644, N1382, N1270);
buf BUF1 (N2496, N2485);
and AND2 (N2497, N2486, N1570);
and AND3 (N2498, N2491, N1720, N2282);
nand NAND2 (N2499, N2478, N468);
nor NOR4 (N2500, N2492, N1463, N45, N360);
buf BUF1 (N2501, N2496);
and AND2 (N2502, N2498, N210);
not NOT1 (N2503, N2502);
buf BUF1 (N2504, N2494);
or OR4 (N2505, N2500, N1889, N1261, N43);
not NOT1 (N2506, N2487);
not NOT1 (N2507, N2493);
and AND4 (N2508, N2483, N461, N1017, N1308);
and AND3 (N2509, N2503, N1268, N676);
nand NAND4 (N2510, N2497, N952, N1215, N1745);
nor NOR3 (N2511, N2505, N1966, N1476);
xor XOR2 (N2512, N2506, N2219);
xor XOR2 (N2513, N2511, N372);
and AND4 (N2514, N2504, N728, N1518, N1851);
or OR2 (N2515, N2514, N1444);
nand NAND2 (N2516, N2515, N347);
and AND2 (N2517, N2508, N475);
buf BUF1 (N2518, N2507);
nor NOR3 (N2519, N2513, N1425, N72);
and AND2 (N2520, N2518, N602);
nor NOR2 (N2521, N2495, N1873);
xor XOR2 (N2522, N2520, N1570);
or OR2 (N2523, N2522, N1669);
and AND3 (N2524, N2510, N1909, N2277);
not NOT1 (N2525, N2512);
or OR2 (N2526, N2524, N2422);
and AND3 (N2527, N2519, N612, N819);
or OR3 (N2528, N2526, N1761, N912);
not NOT1 (N2529, N2499);
and AND4 (N2530, N2528, N2359, N1224, N862);
buf BUF1 (N2531, N2521);
nand NAND3 (N2532, N2527, N2054, N1736);
not NOT1 (N2533, N2523);
and AND2 (N2534, N2517, N1723);
nor NOR4 (N2535, N2525, N1653, N330, N1390);
not NOT1 (N2536, N2501);
not NOT1 (N2537, N2516);
xor XOR2 (N2538, N2536, N625);
and AND4 (N2539, N2532, N2277, N2153, N321);
xor XOR2 (N2540, N2538, N797);
and AND3 (N2541, N2534, N2084, N2191);
or OR2 (N2542, N2530, N724);
not NOT1 (N2543, N2537);
and AND2 (N2544, N2533, N1765);
buf BUF1 (N2545, N2539);
nand NAND4 (N2546, N2544, N1440, N2444, N1217);
xor XOR2 (N2547, N2543, N803);
xor XOR2 (N2548, N2540, N112);
nand NAND3 (N2549, N2529, N1821, N1641);
or OR4 (N2550, N2547, N432, N444, N2086);
xor XOR2 (N2551, N2546, N1448);
or OR2 (N2552, N2531, N2320);
and AND3 (N2553, N2550, N1485, N1623);
and AND3 (N2554, N2541, N1624, N1051);
or OR3 (N2555, N2545, N1810, N1744);
xor XOR2 (N2556, N2548, N339);
and AND3 (N2557, N2555, N551, N2417);
and AND4 (N2558, N2554, N524, N1181, N568);
xor XOR2 (N2559, N2558, N1847);
xor XOR2 (N2560, N2557, N2357);
and AND2 (N2561, N2535, N2149);
and AND2 (N2562, N2552, N518);
and AND4 (N2563, N2560, N1711, N577, N1718);
nand NAND2 (N2564, N2553, N806);
buf BUF1 (N2565, N2509);
xor XOR2 (N2566, N2564, N602);
buf BUF1 (N2567, N2556);
buf BUF1 (N2568, N2567);
xor XOR2 (N2569, N2542, N1571);
nand NAND3 (N2570, N2563, N471, N2082);
xor XOR2 (N2571, N2570, N554);
xor XOR2 (N2572, N2565, N2540);
nor NOR2 (N2573, N2559, N2538);
nand NAND3 (N2574, N2566, N144, N1737);
nand NAND3 (N2575, N2574, N1557, N416);
or OR4 (N2576, N2569, N2197, N1933, N2046);
nand NAND4 (N2577, N2561, N1586, N797, N506);
and AND3 (N2578, N2576, N2072, N723);
not NOT1 (N2579, N2575);
buf BUF1 (N2580, N2551);
and AND2 (N2581, N2577, N859);
nand NAND2 (N2582, N2579, N704);
nor NOR2 (N2583, N2581, N472);
or OR3 (N2584, N2562, N1594, N1454);
xor XOR2 (N2585, N2572, N605);
or OR2 (N2586, N2583, N698);
nand NAND4 (N2587, N2573, N1912, N247, N2225);
not NOT1 (N2588, N2568);
nor NOR4 (N2589, N2571, N1829, N848, N150);
buf BUF1 (N2590, N2580);
xor XOR2 (N2591, N2585, N234);
xor XOR2 (N2592, N2588, N2495);
buf BUF1 (N2593, N2591);
nor NOR4 (N2594, N2586, N682, N1847, N2003);
and AND4 (N2595, N2593, N904, N52, N2171);
and AND3 (N2596, N2592, N1276, N184);
buf BUF1 (N2597, N2549);
and AND3 (N2598, N2584, N383, N1902);
not NOT1 (N2599, N2587);
nor NOR2 (N2600, N2589, N1195);
not NOT1 (N2601, N2582);
xor XOR2 (N2602, N2599, N2106);
nor NOR3 (N2603, N2601, N822, N405);
buf BUF1 (N2604, N2603);
or OR4 (N2605, N2597, N2440, N1855, N200);
xor XOR2 (N2606, N2578, N1587);
and AND2 (N2607, N2594, N1485);
or OR4 (N2608, N2605, N2371, N2292, N96);
and AND3 (N2609, N2608, N397, N1241);
or OR3 (N2610, N2606, N1115, N1773);
buf BUF1 (N2611, N2595);
buf BUF1 (N2612, N2604);
nor NOR2 (N2613, N2590, N1267);
or OR3 (N2614, N2610, N288, N1130);
nand NAND2 (N2615, N2611, N674);
xor XOR2 (N2616, N2613, N1250);
buf BUF1 (N2617, N2609);
xor XOR2 (N2618, N2607, N629);
not NOT1 (N2619, N2598);
nor NOR4 (N2620, N2616, N183, N1658, N864);
xor XOR2 (N2621, N2617, N892);
not NOT1 (N2622, N2596);
xor XOR2 (N2623, N2614, N34);
nor NOR3 (N2624, N2622, N2019, N760);
nor NOR3 (N2625, N2619, N2478, N1328);
nor NOR3 (N2626, N2621, N265, N1083);
nor NOR2 (N2627, N2620, N805);
not NOT1 (N2628, N2623);
xor XOR2 (N2629, N2602, N1678);
and AND3 (N2630, N2628, N1730, N1611);
not NOT1 (N2631, N2615);
nor NOR2 (N2632, N2627, N2231);
nand NAND4 (N2633, N2624, N2545, N2526, N154);
nand NAND4 (N2634, N2618, N2217, N1218, N2082);
or OR3 (N2635, N2630, N2614, N229);
and AND2 (N2636, N2625, N324);
buf BUF1 (N2637, N2635);
nor NOR4 (N2638, N2600, N2138, N1538, N38);
nand NAND4 (N2639, N2631, N2274, N1665, N1865);
xor XOR2 (N2640, N2633, N1175);
nand NAND2 (N2641, N2634, N1439);
nor NOR3 (N2642, N2639, N84, N1841);
not NOT1 (N2643, N2612);
and AND4 (N2644, N2626, N1872, N984, N1644);
xor XOR2 (N2645, N2632, N63);
and AND4 (N2646, N2645, N684, N1626, N1580);
buf BUF1 (N2647, N2646);
and AND2 (N2648, N2638, N1223);
nor NOR2 (N2649, N2647, N186);
xor XOR2 (N2650, N2648, N485);
or OR3 (N2651, N2636, N1047, N701);
xor XOR2 (N2652, N2629, N2528);
nand NAND3 (N2653, N2644, N1597, N147);
buf BUF1 (N2654, N2643);
nand NAND2 (N2655, N2651, N850);
or OR2 (N2656, N2637, N933);
or OR3 (N2657, N2641, N2096, N901);
and AND2 (N2658, N2657, N1101);
and AND4 (N2659, N2642, N219, N1572, N1839);
and AND2 (N2660, N2653, N1100);
xor XOR2 (N2661, N2654, N35);
xor XOR2 (N2662, N2659, N2128);
nand NAND3 (N2663, N2661, N2656, N1789);
buf BUF1 (N2664, N638);
or OR2 (N2665, N2662, N1203);
nor NOR2 (N2666, N2652, N1440);
nor NOR2 (N2667, N2655, N148);
nor NOR2 (N2668, N2658, N1316);
buf BUF1 (N2669, N2665);
nand NAND2 (N2670, N2650, N787);
and AND2 (N2671, N2669, N1486);
and AND3 (N2672, N2649, N2204, N367);
buf BUF1 (N2673, N2663);
buf BUF1 (N2674, N2668);
nor NOR2 (N2675, N2672, N870);
nor NOR4 (N2676, N2667, N2288, N1995, N1752);
buf BUF1 (N2677, N2671);
or OR2 (N2678, N2660, N616);
nor NOR3 (N2679, N2670, N1146, N1475);
or OR2 (N2680, N2666, N2401);
nor NOR3 (N2681, N2640, N2455, N1068);
buf BUF1 (N2682, N2664);
not NOT1 (N2683, N2681);
or OR4 (N2684, N2675, N1323, N2100, N771);
not NOT1 (N2685, N2676);
buf BUF1 (N2686, N2680);
nand NAND4 (N2687, N2678, N1230, N1155, N1701);
xor XOR2 (N2688, N2673, N2205);
buf BUF1 (N2689, N2687);
not NOT1 (N2690, N2685);
not NOT1 (N2691, N2677);
not NOT1 (N2692, N2679);
buf BUF1 (N2693, N2690);
buf BUF1 (N2694, N2682);
buf BUF1 (N2695, N2691);
not NOT1 (N2696, N2686);
buf BUF1 (N2697, N2695);
or OR4 (N2698, N2693, N2599, N2063, N906);
nor NOR3 (N2699, N2688, N238, N1259);
not NOT1 (N2700, N2674);
xor XOR2 (N2701, N2689, N111);
and AND2 (N2702, N2697, N1502);
or OR2 (N2703, N2683, N1773);
not NOT1 (N2704, N2699);
not NOT1 (N2705, N2696);
xor XOR2 (N2706, N2700, N1026);
not NOT1 (N2707, N2704);
nor NOR2 (N2708, N2684, N2349);
nand NAND2 (N2709, N2694, N155);
buf BUF1 (N2710, N2709);
and AND3 (N2711, N2707, N1613, N2433);
xor XOR2 (N2712, N2698, N2379);
buf BUF1 (N2713, N2692);
buf BUF1 (N2714, N2713);
and AND3 (N2715, N2703, N1812, N1393);
xor XOR2 (N2716, N2702, N1266);
nor NOR4 (N2717, N2705, N1013, N2517, N2200);
nor NOR3 (N2718, N2716, N2161, N2436);
xor XOR2 (N2719, N2718, N928);
and AND4 (N2720, N2717, N1513, N137, N2563);
and AND4 (N2721, N2706, N1219, N1202, N505);
nor NOR4 (N2722, N2701, N1468, N2543, N1430);
and AND3 (N2723, N2715, N2094, N360);
nand NAND3 (N2724, N2719, N1286, N2519);
or OR3 (N2725, N2722, N425, N1914);
or OR2 (N2726, N2710, N39);
buf BUF1 (N2727, N2726);
nor NOR4 (N2728, N2725, N2423, N2281, N1746);
not NOT1 (N2729, N2711);
nand NAND2 (N2730, N2724, N1555);
and AND3 (N2731, N2727, N2263, N515);
xor XOR2 (N2732, N2730, N142);
buf BUF1 (N2733, N2731);
buf BUF1 (N2734, N2723);
buf BUF1 (N2735, N2729);
buf BUF1 (N2736, N2721);
buf BUF1 (N2737, N2712);
or OR3 (N2738, N2734, N1549, N2634);
not NOT1 (N2739, N2720);
and AND3 (N2740, N2732, N184, N2027);
not NOT1 (N2741, N2739);
nor NOR4 (N2742, N2737, N889, N2541, N807);
not NOT1 (N2743, N2740);
not NOT1 (N2744, N2714);
not NOT1 (N2745, N2735);
and AND2 (N2746, N2728, N656);
nand NAND2 (N2747, N2746, N1626);
buf BUF1 (N2748, N2747);
and AND3 (N2749, N2745, N2662, N2062);
buf BUF1 (N2750, N2708);
nor NOR2 (N2751, N2742, N945);
buf BUF1 (N2752, N2733);
or OR4 (N2753, N2748, N822, N313, N104);
xor XOR2 (N2754, N2736, N2309);
nand NAND3 (N2755, N2741, N1789, N2192);
and AND3 (N2756, N2738, N2023, N1037);
buf BUF1 (N2757, N2752);
nor NOR4 (N2758, N2744, N2352, N2257, N2663);
not NOT1 (N2759, N2755);
buf BUF1 (N2760, N2751);
nand NAND3 (N2761, N2753, N720, N2472);
buf BUF1 (N2762, N2757);
or OR4 (N2763, N2761, N577, N1782, N2541);
or OR3 (N2764, N2758, N576, N445);
nor NOR2 (N2765, N2763, N279);
nand NAND4 (N2766, N2764, N303, N1331, N2201);
and AND4 (N2767, N2759, N1742, N2654, N2015);
or OR4 (N2768, N2754, N1380, N582, N1328);
or OR3 (N2769, N2750, N1144, N417);
xor XOR2 (N2770, N2769, N343);
nand NAND3 (N2771, N2765, N230, N2706);
nor NOR3 (N2772, N2760, N279, N1783);
nor NOR4 (N2773, N2749, N668, N1543, N1466);
and AND4 (N2774, N2743, N1190, N207, N1223);
not NOT1 (N2775, N2768);
buf BUF1 (N2776, N2756);
nor NOR2 (N2777, N2767, N827);
nand NAND4 (N2778, N2776, N230, N1825, N2760);
not NOT1 (N2779, N2766);
or OR2 (N2780, N2762, N1629);
or OR2 (N2781, N2779, N2362);
xor XOR2 (N2782, N2772, N728);
nor NOR2 (N2783, N2781, N1290);
nor NOR4 (N2784, N2775, N1040, N671, N2710);
nor NOR3 (N2785, N2783, N1617, N1410);
buf BUF1 (N2786, N2770);
xor XOR2 (N2787, N2773, N2029);
or OR3 (N2788, N2780, N436, N1901);
buf BUF1 (N2789, N2777);
nor NOR2 (N2790, N2782, N1299);
buf BUF1 (N2791, N2790);
nor NOR2 (N2792, N2778, N780);
nor NOR2 (N2793, N2784, N666);
xor XOR2 (N2794, N2793, N546);
not NOT1 (N2795, N2792);
nor NOR4 (N2796, N2794, N866, N427, N2464);
nor NOR2 (N2797, N2787, N877);
and AND4 (N2798, N2797, N403, N1170, N2752);
not NOT1 (N2799, N2789);
buf BUF1 (N2800, N2774);
and AND4 (N2801, N2785, N2402, N440, N1179);
nor NOR4 (N2802, N2798, N254, N1284, N2762);
not NOT1 (N2803, N2799);
buf BUF1 (N2804, N2795);
nand NAND4 (N2805, N2788, N1785, N2505, N1156);
nand NAND2 (N2806, N2791, N184);
nor NOR3 (N2807, N2771, N1906, N888);
not NOT1 (N2808, N2807);
nor NOR2 (N2809, N2806, N2783);
nor NOR3 (N2810, N2804, N244, N1951);
xor XOR2 (N2811, N2805, N1495);
buf BUF1 (N2812, N2786);
nor NOR2 (N2813, N2800, N1391);
nand NAND3 (N2814, N2812, N1663, N856);
nor NOR3 (N2815, N2809, N2112, N2322);
nor NOR4 (N2816, N2796, N145, N192, N1011);
buf BUF1 (N2817, N2810);
nor NOR2 (N2818, N2801, N703);
or OR2 (N2819, N2808, N448);
xor XOR2 (N2820, N2814, N815);
nor NOR3 (N2821, N2802, N507, N1340);
xor XOR2 (N2822, N2817, N411);
not NOT1 (N2823, N2819);
xor XOR2 (N2824, N2803, N1130);
and AND3 (N2825, N2823, N661, N2224);
not NOT1 (N2826, N2815);
nor NOR3 (N2827, N2811, N824, N1196);
and AND4 (N2828, N2813, N545, N1271, N2031);
xor XOR2 (N2829, N2826, N1658);
not NOT1 (N2830, N2824);
or OR2 (N2831, N2816, N1520);
buf BUF1 (N2832, N2831);
and AND2 (N2833, N2827, N1751);
or OR3 (N2834, N2822, N2087, N412);
buf BUF1 (N2835, N2832);
and AND3 (N2836, N2825, N494, N1645);
and AND4 (N2837, N2821, N323, N61, N1380);
nand NAND4 (N2838, N2835, N330, N1594, N1760);
nor NOR3 (N2839, N2836, N644, N2375);
buf BUF1 (N2840, N2830);
nand NAND4 (N2841, N2829, N2083, N1483, N422);
or OR2 (N2842, N2818, N2166);
or OR4 (N2843, N2840, N2421, N2510, N2029);
not NOT1 (N2844, N2834);
not NOT1 (N2845, N2844);
and AND3 (N2846, N2842, N74, N2348);
xor XOR2 (N2847, N2846, N395);
nand NAND4 (N2848, N2828, N2130, N2847, N2225);
xor XOR2 (N2849, N2342, N2804);
nor NOR3 (N2850, N2833, N131, N1884);
or OR3 (N2851, N2843, N2354, N1370);
xor XOR2 (N2852, N2850, N1338);
xor XOR2 (N2853, N2841, N1975);
nand NAND4 (N2854, N2820, N1551, N2565, N783);
nand NAND4 (N2855, N2849, N591, N237, N2144);
and AND4 (N2856, N2848, N529, N1708, N1407);
nand NAND2 (N2857, N2851, N1214);
or OR4 (N2858, N2845, N76, N846, N1964);
buf BUF1 (N2859, N2858);
buf BUF1 (N2860, N2839);
not NOT1 (N2861, N2856);
nor NOR3 (N2862, N2861, N1173, N2298);
xor XOR2 (N2863, N2853, N2508);
nor NOR3 (N2864, N2852, N1570, N2336);
xor XOR2 (N2865, N2837, N2511);
nand NAND3 (N2866, N2864, N1351, N1701);
nand NAND2 (N2867, N2838, N2103);
not NOT1 (N2868, N2855);
nor NOR4 (N2869, N2866, N1456, N1321, N1911);
and AND2 (N2870, N2857, N1251);
nor NOR3 (N2871, N2868, N1631, N2180);
xor XOR2 (N2872, N2870, N2291);
or OR4 (N2873, N2862, N1951, N2707, N790);
and AND3 (N2874, N2865, N2581, N286);
or OR3 (N2875, N2872, N2221, N2508);
not NOT1 (N2876, N2854);
nand NAND4 (N2877, N2860, N1854, N584, N922);
nand NAND4 (N2878, N2859, N2425, N170, N727);
nor NOR4 (N2879, N2867, N592, N384, N344);
nand NAND3 (N2880, N2871, N61, N477);
nand NAND2 (N2881, N2869, N574);
or OR2 (N2882, N2878, N1878);
buf BUF1 (N2883, N2879);
nand NAND4 (N2884, N2881, N614, N2608, N1234);
buf BUF1 (N2885, N2882);
and AND3 (N2886, N2873, N2397, N2061);
and AND4 (N2887, N2885, N120, N709, N1116);
buf BUF1 (N2888, N2876);
not NOT1 (N2889, N2877);
nand NAND4 (N2890, N2884, N599, N1800, N2886);
buf BUF1 (N2891, N2270);
buf BUF1 (N2892, N2880);
buf BUF1 (N2893, N2889);
not NOT1 (N2894, N2875);
and AND4 (N2895, N2887, N2278, N2424, N1839);
buf BUF1 (N2896, N2888);
not NOT1 (N2897, N2895);
buf BUF1 (N2898, N2863);
xor XOR2 (N2899, N2890, N2863);
nor NOR3 (N2900, N2883, N300, N2329);
nand NAND3 (N2901, N2893, N1402, N319);
or OR3 (N2902, N2901, N2439, N1004);
and AND3 (N2903, N2897, N1429, N1160);
or OR2 (N2904, N2874, N1795);
xor XOR2 (N2905, N2903, N2328);
xor XOR2 (N2906, N2905, N812);
xor XOR2 (N2907, N2902, N236);
not NOT1 (N2908, N2891);
nor NOR3 (N2909, N2904, N1940, N1584);
nor NOR2 (N2910, N2892, N2089);
nor NOR2 (N2911, N2898, N2750);
buf BUF1 (N2912, N2911);
and AND2 (N2913, N2896, N2835);
and AND2 (N2914, N2913, N1573);
and AND2 (N2915, N2910, N1311);
and AND2 (N2916, N2908, N560);
and AND2 (N2917, N2899, N2063);
buf BUF1 (N2918, N2917);
or OR3 (N2919, N2907, N2316, N383);
buf BUF1 (N2920, N2918);
buf BUF1 (N2921, N2914);
and AND2 (N2922, N2909, N613);
xor XOR2 (N2923, N2922, N1911);
not NOT1 (N2924, N2900);
xor XOR2 (N2925, N2919, N47);
buf BUF1 (N2926, N2924);
nor NOR4 (N2927, N2923, N1524, N2756, N2424);
xor XOR2 (N2928, N2920, N253);
not NOT1 (N2929, N2921);
buf BUF1 (N2930, N2927);
nand NAND2 (N2931, N2925, N1560);
or OR2 (N2932, N2916, N1404);
or OR3 (N2933, N2930, N476, N2096);
or OR2 (N2934, N2912, N408);
and AND3 (N2935, N2929, N1729, N2239);
or OR2 (N2936, N2906, N2284);
xor XOR2 (N2937, N2932, N689);
xor XOR2 (N2938, N2931, N1415);
nand NAND2 (N2939, N2936, N2487);
not NOT1 (N2940, N2938);
or OR2 (N2941, N2934, N2088);
nor NOR4 (N2942, N2940, N2420, N1816, N2895);
nand NAND3 (N2943, N2933, N2429, N1595);
nor NOR4 (N2944, N2926, N1081, N1016, N2572);
buf BUF1 (N2945, N2941);
not NOT1 (N2946, N2942);
or OR3 (N2947, N2928, N2185, N1397);
xor XOR2 (N2948, N2915, N2934);
not NOT1 (N2949, N2943);
nor NOR2 (N2950, N2937, N2161);
nor NOR2 (N2951, N2894, N547);
and AND3 (N2952, N2939, N1448, N2795);
nand NAND3 (N2953, N2952, N2404, N1859);
nand NAND4 (N2954, N2946, N2793, N164, N2811);
buf BUF1 (N2955, N2948);
buf BUF1 (N2956, N2950);
nand NAND4 (N2957, N2935, N1874, N2181, N2081);
not NOT1 (N2958, N2951);
nand NAND3 (N2959, N2945, N2245, N230);
not NOT1 (N2960, N2955);
nor NOR3 (N2961, N2949, N634, N290);
and AND2 (N2962, N2959, N2882);
xor XOR2 (N2963, N2962, N1243);
and AND4 (N2964, N2954, N730, N992, N553);
and AND2 (N2965, N2963, N2944);
buf BUF1 (N2966, N1852);
nor NOR2 (N2967, N2953, N724);
xor XOR2 (N2968, N2966, N2588);
nand NAND4 (N2969, N2947, N296, N529, N658);
nand NAND2 (N2970, N2956, N2210);
not NOT1 (N2971, N2964);
nand NAND2 (N2972, N2961, N2263);
or OR4 (N2973, N2960, N2662, N2876, N1881);
nand NAND3 (N2974, N2968, N2597, N2335);
buf BUF1 (N2975, N2957);
not NOT1 (N2976, N2975);
nor NOR4 (N2977, N2969, N2822, N2036, N1764);
xor XOR2 (N2978, N2974, N446);
nand NAND4 (N2979, N2976, N2667, N1615, N2112);
nand NAND3 (N2980, N2967, N1608, N1731);
nand NAND3 (N2981, N2973, N1843, N1561);
buf BUF1 (N2982, N2978);
not NOT1 (N2983, N2982);
buf BUF1 (N2984, N2972);
or OR2 (N2985, N2984, N1213);
not NOT1 (N2986, N2971);
and AND4 (N2987, N2980, N2723, N395, N286);
or OR2 (N2988, N2987, N2582);
or OR4 (N2989, N2979, N1453, N791, N1815);
nor NOR4 (N2990, N2965, N1986, N2413, N1041);
not NOT1 (N2991, N2983);
nor NOR3 (N2992, N2989, N1417, N1296);
or OR4 (N2993, N2990, N1646, N2179, N1973);
not NOT1 (N2994, N2981);
or OR3 (N2995, N2985, N2660, N1866);
nand NAND4 (N2996, N2970, N1489, N1322, N1403);
and AND3 (N2997, N2996, N2433, N2113);
buf BUF1 (N2998, N2991);
nor NOR2 (N2999, N2997, N989);
nor NOR4 (N3000, N2994, N2613, N2948, N2098);
buf BUF1 (N3001, N2992);
nand NAND2 (N3002, N2977, N803);
and AND2 (N3003, N2995, N2343);
and AND4 (N3004, N3003, N2395, N546, N1422);
xor XOR2 (N3005, N3004, N82);
nand NAND2 (N3006, N3002, N1616);
buf BUF1 (N3007, N2986);
nand NAND3 (N3008, N3000, N3004, N866);
nor NOR2 (N3009, N3006, N706);
or OR3 (N3010, N2993, N929, N2113);
and AND3 (N3011, N2958, N1674, N1530);
xor XOR2 (N3012, N3007, N2984);
and AND3 (N3013, N3010, N1413, N715);
xor XOR2 (N3014, N2988, N2143);
not NOT1 (N3015, N3005);
and AND3 (N3016, N3009, N684, N2614);
xor XOR2 (N3017, N3013, N239);
xor XOR2 (N3018, N2999, N820);
nor NOR4 (N3019, N3012, N1030, N476, N730);
xor XOR2 (N3020, N3011, N725);
xor XOR2 (N3021, N3019, N457);
or OR4 (N3022, N3014, N393, N2738, N1854);
nand NAND2 (N3023, N3022, N2891);
nand NAND4 (N3024, N3021, N1731, N73, N2271);
buf BUF1 (N3025, N3016);
nand NAND2 (N3026, N3015, N412);
nand NAND2 (N3027, N3018, N136);
nand NAND3 (N3028, N3023, N2272, N1802);
nand NAND4 (N3029, N3008, N1253, N1761, N1234);
or OR3 (N3030, N3001, N1230, N2255);
not NOT1 (N3031, N3017);
nor NOR3 (N3032, N3030, N2130, N1227);
or OR2 (N3033, N2998, N525);
and AND4 (N3034, N3033, N2510, N2270, N1553);
and AND3 (N3035, N3027, N1170, N760);
or OR4 (N3036, N3032, N732, N896, N2529);
buf BUF1 (N3037, N3036);
buf BUF1 (N3038, N3029);
nor NOR3 (N3039, N3025, N2266, N481);
xor XOR2 (N3040, N3039, N1162);
nand NAND3 (N3041, N3034, N1680, N1027);
and AND4 (N3042, N3035, N396, N667, N2917);
and AND2 (N3043, N3020, N2522);
buf BUF1 (N3044, N3037);
xor XOR2 (N3045, N3043, N2009);
not NOT1 (N3046, N3031);
nand NAND4 (N3047, N3038, N325, N527, N1582);
xor XOR2 (N3048, N3024, N2461);
xor XOR2 (N3049, N3042, N2142);
buf BUF1 (N3050, N3044);
buf BUF1 (N3051, N3026);
nand NAND2 (N3052, N3045, N254);
and AND2 (N3053, N3040, N232);
buf BUF1 (N3054, N3049);
or OR3 (N3055, N3050, N3054, N1968);
buf BUF1 (N3056, N2481);
and AND2 (N3057, N3055, N540);
xor XOR2 (N3058, N3051, N2209);
nand NAND2 (N3059, N3053, N967);
nor NOR2 (N3060, N3047, N2764);
buf BUF1 (N3061, N3048);
xor XOR2 (N3062, N3056, N1944);
nor NOR3 (N3063, N3057, N1003, N2766);
nand NAND3 (N3064, N3063, N2980, N1443);
buf BUF1 (N3065, N3041);
not NOT1 (N3066, N3062);
xor XOR2 (N3067, N3060, N1621);
nand NAND2 (N3068, N3066, N1078);
nand NAND4 (N3069, N3061, N763, N281, N674);
nand NAND3 (N3070, N3065, N319, N1712);
not NOT1 (N3071, N3068);
buf BUF1 (N3072, N3046);
xor XOR2 (N3073, N3058, N570);
not NOT1 (N3074, N3073);
nor NOR2 (N3075, N3071, N2595);
xor XOR2 (N3076, N3052, N1547);
nand NAND3 (N3077, N3064, N1084, N2988);
nor NOR2 (N3078, N3028, N254);
buf BUF1 (N3079, N3067);
or OR2 (N3080, N3074, N1030);
or OR4 (N3081, N3069, N202, N26, N551);
or OR4 (N3082, N3059, N36, N237, N2960);
nor NOR4 (N3083, N3080, N516, N2833, N937);
or OR4 (N3084, N3079, N2960, N369, N1527);
buf BUF1 (N3085, N3081);
buf BUF1 (N3086, N3082);
xor XOR2 (N3087, N3077, N2242);
not NOT1 (N3088, N3086);
or OR2 (N3089, N3075, N278);
nor NOR3 (N3090, N3076, N2933, N914);
xor XOR2 (N3091, N3085, N272);
nor NOR3 (N3092, N3088, N2777, N2108);
or OR3 (N3093, N3092, N2197, N2701);
nor NOR2 (N3094, N3083, N2606);
or OR2 (N3095, N3072, N1975);
nor NOR4 (N3096, N3078, N966, N615, N355);
nor NOR3 (N3097, N3089, N539, N2885);
buf BUF1 (N3098, N3096);
not NOT1 (N3099, N3070);
and AND3 (N3100, N3084, N2330, N2780);
or OR2 (N3101, N3093, N462);
nand NAND4 (N3102, N3098, N3034, N1840, N2741);
nor NOR4 (N3103, N3101, N949, N1752, N1305);
xor XOR2 (N3104, N3097, N642);
nor NOR2 (N3105, N3103, N2961);
nor NOR2 (N3106, N3105, N1166);
xor XOR2 (N3107, N3091, N408);
nand NAND2 (N3108, N3099, N1962);
nor NOR3 (N3109, N3102, N2511, N959);
and AND2 (N3110, N3095, N55);
nor NOR2 (N3111, N3106, N725);
and AND4 (N3112, N3110, N2990, N2000, N610);
and AND4 (N3113, N3094, N952, N428, N377);
buf BUF1 (N3114, N3104);
nor NOR4 (N3115, N3107, N319, N1525, N2672);
xor XOR2 (N3116, N3109, N2849);
buf BUF1 (N3117, N3111);
xor XOR2 (N3118, N3090, N2178);
xor XOR2 (N3119, N3118, N427);
or OR3 (N3120, N3114, N119, N912);
xor XOR2 (N3121, N3112, N818);
not NOT1 (N3122, N3120);
and AND3 (N3123, N3087, N2413, N2721);
xor XOR2 (N3124, N3117, N1346);
nor NOR2 (N3125, N3108, N1948);
xor XOR2 (N3126, N3123, N906);
xor XOR2 (N3127, N3121, N2241);
not NOT1 (N3128, N3113);
not NOT1 (N3129, N3116);
buf BUF1 (N3130, N3129);
xor XOR2 (N3131, N3100, N2094);
not NOT1 (N3132, N3122);
nor NOR3 (N3133, N3125, N510, N2927);
xor XOR2 (N3134, N3119, N1770);
or OR2 (N3135, N3130, N369);
xor XOR2 (N3136, N3128, N346);
xor XOR2 (N3137, N3132, N2761);
nand NAND2 (N3138, N3126, N2665);
buf BUF1 (N3139, N3127);
or OR3 (N3140, N3138, N2095, N1011);
and AND2 (N3141, N3131, N2283);
not NOT1 (N3142, N3136);
and AND3 (N3143, N3137, N2778, N2121);
nor NOR2 (N3144, N3142, N2695);
and AND4 (N3145, N3135, N2062, N2366, N711);
not NOT1 (N3146, N3133);
not NOT1 (N3147, N3146);
buf BUF1 (N3148, N3134);
or OR2 (N3149, N3115, N1505);
or OR3 (N3150, N3144, N2837, N2842);
or OR3 (N3151, N3149, N958, N1660);
or OR4 (N3152, N3147, N1289, N265, N353);
xor XOR2 (N3153, N3152, N1083);
xor XOR2 (N3154, N3141, N3148);
nand NAND4 (N3155, N2895, N396, N2347, N2016);
nor NOR3 (N3156, N3124, N701, N2494);
or OR4 (N3157, N3151, N886, N1130, N1230);
xor XOR2 (N3158, N3155, N2504);
nand NAND4 (N3159, N3156, N3065, N2244, N3147);
buf BUF1 (N3160, N3154);
nor NOR3 (N3161, N3159, N56, N514);
not NOT1 (N3162, N3150);
and AND3 (N3163, N3161, N678, N464);
xor XOR2 (N3164, N3145, N2013);
xor XOR2 (N3165, N3162, N1726);
and AND2 (N3166, N3143, N831);
xor XOR2 (N3167, N3139, N604);
or OR2 (N3168, N3157, N524);
or OR2 (N3169, N3140, N1576);
xor XOR2 (N3170, N3160, N2988);
xor XOR2 (N3171, N3170, N1878);
or OR2 (N3172, N3168, N1466);
not NOT1 (N3173, N3171);
nor NOR4 (N3174, N3172, N2590, N2488, N126);
or OR3 (N3175, N3153, N1979, N384);
nor NOR2 (N3176, N3169, N115);
not NOT1 (N3177, N3167);
nand NAND3 (N3178, N3163, N383, N1038);
not NOT1 (N3179, N3164);
not NOT1 (N3180, N3177);
not NOT1 (N3181, N3158);
and AND2 (N3182, N3166, N2095);
or OR4 (N3183, N3174, N2698, N531, N2310);
xor XOR2 (N3184, N3175, N2048);
nand NAND2 (N3185, N3180, N2545);
not NOT1 (N3186, N3179);
nand NAND2 (N3187, N3165, N1989);
nand NAND2 (N3188, N3184, N2603);
buf BUF1 (N3189, N3187);
nor NOR4 (N3190, N3173, N2247, N1767, N1335);
not NOT1 (N3191, N3178);
not NOT1 (N3192, N3176);
nand NAND2 (N3193, N3181, N141);
not NOT1 (N3194, N3191);
nand NAND2 (N3195, N3189, N2689);
buf BUF1 (N3196, N3193);
nand NAND4 (N3197, N3194, N3179, N3196, N3083);
buf BUF1 (N3198, N764);
not NOT1 (N3199, N3185);
nor NOR4 (N3200, N3190, N1921, N1847, N2105);
nand NAND2 (N3201, N3199, N88);
xor XOR2 (N3202, N3183, N2588);
buf BUF1 (N3203, N3198);
not NOT1 (N3204, N3186);
not NOT1 (N3205, N3195);
buf BUF1 (N3206, N3205);
nor NOR2 (N3207, N3203, N1926);
and AND3 (N3208, N3201, N2013, N2012);
buf BUF1 (N3209, N3208);
xor XOR2 (N3210, N3204, N2627);
buf BUF1 (N3211, N3197);
not NOT1 (N3212, N3211);
nor NOR2 (N3213, N3182, N2635);
and AND2 (N3214, N3188, N884);
buf BUF1 (N3215, N3202);
or OR4 (N3216, N3207, N1842, N924, N1612);
nand NAND3 (N3217, N3206, N973, N3147);
not NOT1 (N3218, N3217);
not NOT1 (N3219, N3213);
xor XOR2 (N3220, N3212, N639);
nor NOR2 (N3221, N3216, N1843);
xor XOR2 (N3222, N3210, N374);
buf BUF1 (N3223, N3215);
or OR2 (N3224, N3209, N1305);
and AND4 (N3225, N3222, N728, N2312, N878);
or OR2 (N3226, N3225, N2847);
buf BUF1 (N3227, N3220);
and AND3 (N3228, N3224, N2937, N2540);
buf BUF1 (N3229, N3223);
or OR2 (N3230, N3221, N1039);
not NOT1 (N3231, N3214);
not NOT1 (N3232, N3227);
and AND4 (N3233, N3226, N766, N293, N434);
and AND2 (N3234, N3218, N459);
xor XOR2 (N3235, N3234, N2010);
or OR4 (N3236, N3219, N2392, N1838, N1994);
buf BUF1 (N3237, N3228);
nor NOR2 (N3238, N3229, N1484);
not NOT1 (N3239, N3192);
nand NAND3 (N3240, N3233, N899, N1742);
nand NAND3 (N3241, N3239, N2332, N159);
nor NOR4 (N3242, N3240, N2879, N1266, N1619);
nor NOR2 (N3243, N3232, N2433);
and AND3 (N3244, N3238, N1944, N2499);
nor NOR3 (N3245, N3235, N382, N1842);
or OR2 (N3246, N3245, N766);
not NOT1 (N3247, N3236);
nand NAND4 (N3248, N3241, N3012, N688, N3043);
xor XOR2 (N3249, N3247, N3045);
buf BUF1 (N3250, N3249);
not NOT1 (N3251, N3244);
buf BUF1 (N3252, N3237);
nand NAND4 (N3253, N3252, N2837, N758, N2008);
or OR3 (N3254, N3251, N868, N2720);
or OR2 (N3255, N3253, N2545);
nand NAND4 (N3256, N3255, N3218, N1397, N75);
buf BUF1 (N3257, N3231);
nand NAND2 (N3258, N3230, N1852);
nor NOR3 (N3259, N3243, N1101, N1512);
and AND4 (N3260, N3258, N1836, N1702, N945);
nand NAND2 (N3261, N3260, N1190);
nand NAND2 (N3262, N3200, N2840);
and AND3 (N3263, N3248, N2494, N1731);
nand NAND4 (N3264, N3263, N3256, N2847, N2143);
xor XOR2 (N3265, N969, N450);
xor XOR2 (N3266, N3257, N2566);
nor NOR2 (N3267, N3262, N1216);
not NOT1 (N3268, N3246);
or OR2 (N3269, N3266, N316);
buf BUF1 (N3270, N3259);
nor NOR3 (N3271, N3261, N1770, N1361);
buf BUF1 (N3272, N3268);
xor XOR2 (N3273, N3264, N1121);
nand NAND3 (N3274, N3267, N2701, N20);
or OR4 (N3275, N3242, N2589, N2757, N29);
nand NAND3 (N3276, N3254, N1474, N842);
nor NOR3 (N3277, N3265, N560, N1602);
xor XOR2 (N3278, N3271, N1977);
nand NAND4 (N3279, N3250, N1639, N426, N1260);
nand NAND2 (N3280, N3273, N544);
or OR3 (N3281, N3275, N759, N1712);
nand NAND2 (N3282, N3276, N82);
buf BUF1 (N3283, N3274);
or OR4 (N3284, N3278, N1283, N3168, N193);
nand NAND4 (N3285, N3283, N3242, N1359, N1553);
or OR2 (N3286, N3277, N205);
nand NAND4 (N3287, N3284, N2748, N56, N915);
and AND3 (N3288, N3279, N2591, N1419);
nand NAND2 (N3289, N3269, N2480);
nand NAND2 (N3290, N3288, N2465);
not NOT1 (N3291, N3289);
nor NOR4 (N3292, N3291, N1312, N3232, N1041);
not NOT1 (N3293, N3287);
and AND4 (N3294, N3292, N1711, N811, N2920);
nand NAND3 (N3295, N3282, N1842, N2962);
or OR4 (N3296, N3294, N1086, N1542, N2759);
buf BUF1 (N3297, N3293);
nand NAND3 (N3298, N3296, N774, N498);
nor NOR2 (N3299, N3280, N3193);
nor NOR3 (N3300, N3290, N2441, N3129);
xor XOR2 (N3301, N3298, N1991);
nor NOR2 (N3302, N3297, N2417);
or OR2 (N3303, N3302, N433);
and AND3 (N3304, N3303, N2027, N380);
or OR3 (N3305, N3272, N1687, N1698);
and AND4 (N3306, N3300, N1236, N3198, N321);
and AND3 (N3307, N3285, N134, N1419);
and AND2 (N3308, N3286, N283);
or OR2 (N3309, N3308, N1199);
nand NAND4 (N3310, N3305, N1077, N1994, N160);
nor NOR3 (N3311, N3304, N178, N1776);
buf BUF1 (N3312, N3306);
nor NOR4 (N3313, N3299, N1096, N2429, N2980);
nand NAND4 (N3314, N3295, N3250, N2377, N3123);
buf BUF1 (N3315, N3307);
buf BUF1 (N3316, N3311);
not NOT1 (N3317, N3281);
xor XOR2 (N3318, N3312, N2898);
buf BUF1 (N3319, N3318);
xor XOR2 (N3320, N3317, N278);
buf BUF1 (N3321, N3320);
and AND3 (N3322, N3310, N2014, N1099);
not NOT1 (N3323, N3309);
buf BUF1 (N3324, N3321);
nand NAND3 (N3325, N3314, N2264, N1259);
and AND4 (N3326, N3313, N1672, N3088, N2937);
not NOT1 (N3327, N3323);
buf BUF1 (N3328, N3322);
not NOT1 (N3329, N3315);
buf BUF1 (N3330, N3301);
or OR3 (N3331, N3330, N581, N2586);
xor XOR2 (N3332, N3331, N2333);
nand NAND3 (N3333, N3316, N3292, N547);
not NOT1 (N3334, N3270);
or OR3 (N3335, N3332, N617, N417);
buf BUF1 (N3336, N3324);
xor XOR2 (N3337, N3334, N2281);
xor XOR2 (N3338, N3337, N1863);
nor NOR3 (N3339, N3335, N1363, N288);
nand NAND3 (N3340, N3325, N3177, N1734);
xor XOR2 (N3341, N3333, N2534);
or OR3 (N3342, N3339, N2482, N2680);
nor NOR4 (N3343, N3329, N3241, N2926, N1179);
buf BUF1 (N3344, N3336);
xor XOR2 (N3345, N3319, N3343);
buf BUF1 (N3346, N3191);
and AND3 (N3347, N3326, N2812, N1989);
nor NOR3 (N3348, N3342, N1025, N1111);
nand NAND4 (N3349, N3327, N884, N2180, N1056);
and AND2 (N3350, N3349, N356);
or OR2 (N3351, N3348, N389);
xor XOR2 (N3352, N3340, N1353);
buf BUF1 (N3353, N3350);
buf BUF1 (N3354, N3328);
xor XOR2 (N3355, N3341, N2770);
nor NOR4 (N3356, N3344, N1917, N569, N43);
nor NOR3 (N3357, N3353, N1695, N647);
not NOT1 (N3358, N3347);
xor XOR2 (N3359, N3356, N29);
not NOT1 (N3360, N3355);
not NOT1 (N3361, N3358);
xor XOR2 (N3362, N3351, N1379);
buf BUF1 (N3363, N3362);
not NOT1 (N3364, N3346);
and AND3 (N3365, N3360, N458, N588);
nor NOR2 (N3366, N3354, N2044);
buf BUF1 (N3367, N3361);
buf BUF1 (N3368, N3364);
not NOT1 (N3369, N3352);
not NOT1 (N3370, N3338);
or OR3 (N3371, N3363, N651, N1436);
buf BUF1 (N3372, N3345);
and AND4 (N3373, N3365, N2514, N1321, N2031);
nand NAND2 (N3374, N3373, N2492);
xor XOR2 (N3375, N3357, N550);
xor XOR2 (N3376, N3375, N3300);
nand NAND4 (N3377, N3370, N1466, N2328, N3234);
buf BUF1 (N3378, N3376);
or OR3 (N3379, N3366, N444, N1007);
and AND2 (N3380, N3377, N516);
buf BUF1 (N3381, N3374);
nor NOR2 (N3382, N3369, N3070);
or OR2 (N3383, N3359, N1205);
not NOT1 (N3384, N3379);
nor NOR4 (N3385, N3383, N3128, N2811, N644);
nor NOR3 (N3386, N3368, N742, N2686);
buf BUF1 (N3387, N3367);
not NOT1 (N3388, N3385);
or OR3 (N3389, N3371, N170, N2179);
and AND3 (N3390, N3388, N1263, N1129);
nor NOR2 (N3391, N3378, N135);
buf BUF1 (N3392, N3389);
and AND2 (N3393, N3390, N3208);
not NOT1 (N3394, N3393);
xor XOR2 (N3395, N3372, N1059);
xor XOR2 (N3396, N3394, N2233);
nor NOR3 (N3397, N3391, N977, N2801);
nor NOR2 (N3398, N3387, N1235);
not NOT1 (N3399, N3395);
nand NAND2 (N3400, N3392, N1061);
nand NAND3 (N3401, N3384, N3178, N3151);
nor NOR2 (N3402, N3386, N2625);
nand NAND2 (N3403, N3400, N686);
not NOT1 (N3404, N3382);
nand NAND3 (N3405, N3402, N429, N135);
nor NOR3 (N3406, N3381, N656, N1430);
or OR4 (N3407, N3401, N1962, N2966, N3224);
xor XOR2 (N3408, N3380, N805);
and AND3 (N3409, N3406, N1670, N137);
nand NAND4 (N3410, N3407, N228, N1057, N1416);
and AND3 (N3411, N3396, N845, N151);
or OR2 (N3412, N3399, N1775);
not NOT1 (N3413, N3411);
nand NAND4 (N3414, N3409, N157, N3160, N1457);
xor XOR2 (N3415, N3404, N1475);
nand NAND2 (N3416, N3403, N2942);
xor XOR2 (N3417, N3398, N841);
or OR3 (N3418, N3413, N1284, N3331);
buf BUF1 (N3419, N3410);
and AND4 (N3420, N3397, N1977, N1901, N3064);
xor XOR2 (N3421, N3420, N1915);
or OR4 (N3422, N3412, N2265, N2027, N2073);
xor XOR2 (N3423, N3421, N336);
and AND2 (N3424, N3408, N3357);
and AND4 (N3425, N3414, N3253, N2401, N947);
buf BUF1 (N3426, N3424);
nor NOR3 (N3427, N3426, N3099, N1102);
or OR3 (N3428, N3423, N2377, N1854);
nor NOR2 (N3429, N3416, N3280);
or OR3 (N3430, N3427, N1989, N3234);
nand NAND2 (N3431, N3417, N2590);
not NOT1 (N3432, N3422);
nand NAND3 (N3433, N3415, N2607, N1754);
xor XOR2 (N3434, N3428, N937);
not NOT1 (N3435, N3430);
buf BUF1 (N3436, N3418);
or OR4 (N3437, N3432, N2938, N703, N1523);
or OR2 (N3438, N3431, N785);
xor XOR2 (N3439, N3419, N2917);
nor NOR4 (N3440, N3433, N72, N1308, N910);
nor NOR2 (N3441, N3435, N764);
nand NAND3 (N3442, N3405, N3149, N1714);
or OR2 (N3443, N3429, N449);
xor XOR2 (N3444, N3442, N1870);
buf BUF1 (N3445, N3425);
and AND2 (N3446, N3440, N3069);
xor XOR2 (N3447, N3441, N602);
or OR4 (N3448, N3438, N1616, N19, N3286);
nand NAND2 (N3449, N3439, N3325);
or OR2 (N3450, N3443, N1278);
nand NAND4 (N3451, N3448, N433, N2903, N1837);
and AND4 (N3452, N3436, N1368, N84, N3108);
nand NAND3 (N3453, N3450, N917, N1645);
and AND4 (N3454, N3447, N777, N3208, N213);
or OR3 (N3455, N3454, N3334, N3203);
and AND4 (N3456, N3437, N164, N896, N1150);
xor XOR2 (N3457, N3453, N1226);
nor NOR2 (N3458, N3434, N3137);
buf BUF1 (N3459, N3446);
not NOT1 (N3460, N3445);
nand NAND3 (N3461, N3452, N1387, N2582);
buf BUF1 (N3462, N3458);
xor XOR2 (N3463, N3459, N1229);
nor NOR2 (N3464, N3444, N1924);
not NOT1 (N3465, N3464);
and AND4 (N3466, N3460, N3220, N3123, N235);
nor NOR3 (N3467, N3461, N1141, N3207);
not NOT1 (N3468, N3467);
nand NAND2 (N3469, N3466, N407);
and AND2 (N3470, N3455, N1017);
nand NAND2 (N3471, N3451, N118);
and AND3 (N3472, N3449, N1847, N2832);
buf BUF1 (N3473, N3463);
nor NOR4 (N3474, N3470, N330, N1431, N406);
not NOT1 (N3475, N3472);
and AND3 (N3476, N3462, N902, N2742);
or OR3 (N3477, N3475, N2878, N104);
and AND3 (N3478, N3468, N655, N938);
nor NOR3 (N3479, N3465, N2402, N1243);
xor XOR2 (N3480, N3473, N987);
nor NOR4 (N3481, N3469, N1979, N28, N3405);
not NOT1 (N3482, N3456);
xor XOR2 (N3483, N3477, N224);
nor NOR3 (N3484, N3481, N3225, N449);
nand NAND4 (N3485, N3483, N2124, N1736, N2432);
buf BUF1 (N3486, N3482);
nand NAND4 (N3487, N3486, N2001, N3279, N728);
xor XOR2 (N3488, N3474, N1974);
not NOT1 (N3489, N3485);
and AND4 (N3490, N3487, N465, N1909, N2081);
buf BUF1 (N3491, N3457);
or OR2 (N3492, N3491, N316);
nor NOR2 (N3493, N3476, N2823);
not NOT1 (N3494, N3490);
buf BUF1 (N3495, N3492);
buf BUF1 (N3496, N3495);
nor NOR4 (N3497, N3471, N460, N130, N2402);
not NOT1 (N3498, N3496);
or OR3 (N3499, N3498, N2009, N2898);
or OR3 (N3500, N3494, N2401, N3175);
nor NOR2 (N3501, N3478, N3277);
nand NAND2 (N3502, N3479, N370);
or OR3 (N3503, N3493, N1554, N2276);
xor XOR2 (N3504, N3484, N2752);
xor XOR2 (N3505, N3502, N1606);
not NOT1 (N3506, N3505);
buf BUF1 (N3507, N3480);
xor XOR2 (N3508, N3500, N1537);
xor XOR2 (N3509, N3503, N2540);
or OR2 (N3510, N3489, N1691);
or OR3 (N3511, N3506, N2754, N2133);
buf BUF1 (N3512, N3497);
xor XOR2 (N3513, N3510, N2657);
xor XOR2 (N3514, N3511, N1350);
xor XOR2 (N3515, N3513, N1264);
buf BUF1 (N3516, N3512);
and AND4 (N3517, N3504, N1168, N614, N492);
not NOT1 (N3518, N3488);
not NOT1 (N3519, N3501);
xor XOR2 (N3520, N3499, N1294);
and AND2 (N3521, N3508, N1197);
xor XOR2 (N3522, N3516, N2485);
xor XOR2 (N3523, N3518, N1204);
or OR3 (N3524, N3519, N3024, N3436);
buf BUF1 (N3525, N3514);
nor NOR4 (N3526, N3524, N2258, N571, N2277);
nor NOR2 (N3527, N3522, N1139);
not NOT1 (N3528, N3509);
buf BUF1 (N3529, N3520);
nor NOR4 (N3530, N3517, N1031, N2130, N3238);
and AND2 (N3531, N3528, N859);
nor NOR4 (N3532, N3521, N2079, N2506, N3342);
xor XOR2 (N3533, N3515, N89);
not NOT1 (N3534, N3530);
not NOT1 (N3535, N3527);
buf BUF1 (N3536, N3523);
xor XOR2 (N3537, N3529, N2269);
nor NOR2 (N3538, N3534, N1371);
nand NAND2 (N3539, N3531, N173);
xor XOR2 (N3540, N3538, N569);
nor NOR2 (N3541, N3507, N187);
not NOT1 (N3542, N3541);
not NOT1 (N3543, N3532);
and AND2 (N3544, N3526, N274);
not NOT1 (N3545, N3540);
buf BUF1 (N3546, N3544);
and AND3 (N3547, N3525, N2454, N1032);
not NOT1 (N3548, N3539);
buf BUF1 (N3549, N3543);
and AND4 (N3550, N3548, N3292, N856, N104);
not NOT1 (N3551, N3535);
not NOT1 (N3552, N3547);
nand NAND4 (N3553, N3552, N3317, N823, N415);
not NOT1 (N3554, N3537);
nand NAND2 (N3555, N3550, N236);
nand NAND2 (N3556, N3542, N3341);
buf BUF1 (N3557, N3533);
nor NOR4 (N3558, N3557, N2570, N43, N1878);
not NOT1 (N3559, N3549);
nand NAND3 (N3560, N3556, N1259, N3212);
not NOT1 (N3561, N3555);
and AND3 (N3562, N3561, N482, N741);
nand NAND3 (N3563, N3562, N2936, N1621);
and AND3 (N3564, N3559, N1483, N535);
buf BUF1 (N3565, N3554);
and AND2 (N3566, N3565, N2433);
xor XOR2 (N3567, N3558, N752);
nor NOR4 (N3568, N3560, N2923, N828, N803);
buf BUF1 (N3569, N3545);
not NOT1 (N3570, N3536);
buf BUF1 (N3571, N3568);
buf BUF1 (N3572, N3570);
and AND2 (N3573, N3564, N3212);
and AND2 (N3574, N3567, N1978);
and AND3 (N3575, N3572, N282, N1706);
nand NAND4 (N3576, N3571, N3440, N2197, N380);
and AND3 (N3577, N3576, N1107, N735);
buf BUF1 (N3578, N3574);
nor NOR2 (N3579, N3578, N2836);
not NOT1 (N3580, N3579);
nor NOR4 (N3581, N3569, N548, N362, N2917);
xor XOR2 (N3582, N3551, N2034);
not NOT1 (N3583, N3581);
nor NOR4 (N3584, N3583, N1327, N2399, N1721);
not NOT1 (N3585, N3584);
nor NOR2 (N3586, N3563, N1055);
buf BUF1 (N3587, N3566);
xor XOR2 (N3588, N3575, N1115);
nor NOR4 (N3589, N3573, N3182, N2962, N64);
nor NOR2 (N3590, N3580, N2595);
xor XOR2 (N3591, N3585, N3021);
xor XOR2 (N3592, N3588, N134);
nand NAND2 (N3593, N3589, N357);
nand NAND2 (N3594, N3582, N2742);
buf BUF1 (N3595, N3546);
buf BUF1 (N3596, N3587);
xor XOR2 (N3597, N3594, N2496);
nand NAND3 (N3598, N3577, N2125, N2291);
nand NAND3 (N3599, N3597, N3306, N2340);
nand NAND4 (N3600, N3598, N2340, N181, N2689);
nand NAND2 (N3601, N3595, N3032);
or OR4 (N3602, N3596, N1071, N2042, N333);
not NOT1 (N3603, N3586);
or OR2 (N3604, N3602, N144);
nor NOR2 (N3605, N3591, N1942);
nand NAND2 (N3606, N3600, N3032);
nor NOR4 (N3607, N3601, N2558, N741, N925);
xor XOR2 (N3608, N3605, N881);
not NOT1 (N3609, N3603);
or OR3 (N3610, N3590, N2550, N3575);
and AND2 (N3611, N3553, N3587);
not NOT1 (N3612, N3610);
xor XOR2 (N3613, N3593, N1623);
and AND2 (N3614, N3604, N467);
and AND3 (N3615, N3611, N3114, N3200);
not NOT1 (N3616, N3609);
and AND2 (N3617, N3614, N2642);
nor NOR4 (N3618, N3599, N3247, N1653, N2265);
xor XOR2 (N3619, N3612, N181);
buf BUF1 (N3620, N3592);
not NOT1 (N3621, N3607);
and AND2 (N3622, N3620, N1689);
nor NOR2 (N3623, N3608, N2200);
nor NOR3 (N3624, N3615, N882, N543);
nand NAND4 (N3625, N3618, N92, N3330, N965);
and AND2 (N3626, N3617, N3481);
and AND3 (N3627, N3624, N3187, N231);
nor NOR4 (N3628, N3616, N2505, N79, N1152);
xor XOR2 (N3629, N3622, N2658);
nand NAND4 (N3630, N3623, N3459, N85, N2580);
nand NAND4 (N3631, N3626, N2194, N1896, N906);
and AND2 (N3632, N3630, N282);
xor XOR2 (N3633, N3613, N1453);
nand NAND2 (N3634, N3633, N2515);
xor XOR2 (N3635, N3632, N1852);
nor NOR4 (N3636, N3606, N577, N1582, N242);
and AND2 (N3637, N3634, N3456);
not NOT1 (N3638, N3621);
nand NAND2 (N3639, N3635, N1891);
nand NAND2 (N3640, N3619, N2811);
nor NOR3 (N3641, N3625, N2635, N2464);
not NOT1 (N3642, N3637);
xor XOR2 (N3643, N3627, N210);
or OR2 (N3644, N3639, N654);
and AND3 (N3645, N3638, N924, N2588);
buf BUF1 (N3646, N3640);
and AND3 (N3647, N3643, N2324, N815);
xor XOR2 (N3648, N3646, N2731);
buf BUF1 (N3649, N3644);
not NOT1 (N3650, N3628);
or OR2 (N3651, N3650, N2515);
and AND4 (N3652, N3642, N2661, N2384, N1481);
and AND2 (N3653, N3648, N3518);
buf BUF1 (N3654, N3631);
or OR4 (N3655, N3645, N2913, N1401, N230);
and AND3 (N3656, N3652, N2520, N3393);
or OR2 (N3657, N3653, N3239);
and AND3 (N3658, N3655, N999, N343);
not NOT1 (N3659, N3647);
buf BUF1 (N3660, N3657);
or OR2 (N3661, N3654, N807);
or OR2 (N3662, N3641, N1165);
buf BUF1 (N3663, N3662);
nand NAND4 (N3664, N3656, N1903, N2507, N2976);
or OR3 (N3665, N3651, N2956, N1711);
or OR3 (N3666, N3658, N2804, N3108);
nand NAND4 (N3667, N3666, N1007, N3383, N3091);
or OR2 (N3668, N3659, N916);
and AND2 (N3669, N3664, N2778);
xor XOR2 (N3670, N3649, N912);
not NOT1 (N3671, N3665);
xor XOR2 (N3672, N3661, N3254);
or OR3 (N3673, N3672, N2109, N2576);
nor NOR4 (N3674, N3673, N2210, N3501, N1302);
or OR2 (N3675, N3629, N887);
buf BUF1 (N3676, N3660);
nand NAND2 (N3677, N3671, N622);
and AND3 (N3678, N3674, N989, N3331);
nor NOR3 (N3679, N3677, N72, N1996);
xor XOR2 (N3680, N3669, N2525);
nor NOR4 (N3681, N3675, N603, N2371, N2220);
or OR4 (N3682, N3668, N2940, N3636, N3071);
nor NOR4 (N3683, N367, N2365, N571, N2309);
and AND4 (N3684, N3682, N2860, N1899, N3231);
xor XOR2 (N3685, N3681, N1002);
nand NAND3 (N3686, N3667, N3233, N3389);
nor NOR4 (N3687, N3686, N2308, N2499, N2211);
xor XOR2 (N3688, N3684, N2174);
xor XOR2 (N3689, N3663, N1564);
nand NAND2 (N3690, N3678, N3295);
nor NOR2 (N3691, N3670, N1473);
xor XOR2 (N3692, N3683, N452);
and AND2 (N3693, N3685, N2819);
or OR3 (N3694, N3687, N122, N2153);
and AND4 (N3695, N3693, N157, N2798, N2545);
buf BUF1 (N3696, N3680);
buf BUF1 (N3697, N3679);
or OR4 (N3698, N3695, N2362, N819, N2620);
nor NOR4 (N3699, N3694, N2039, N1539, N2890);
or OR2 (N3700, N3699, N2689);
nor NOR4 (N3701, N3700, N3639, N1401, N1173);
not NOT1 (N3702, N3696);
buf BUF1 (N3703, N3691);
buf BUF1 (N3704, N3690);
not NOT1 (N3705, N3692);
nor NOR2 (N3706, N3701, N1543);
or OR4 (N3707, N3676, N195, N127, N3418);
or OR2 (N3708, N3703, N122);
buf BUF1 (N3709, N3705);
nor NOR4 (N3710, N3709, N1290, N187, N1243);
nand NAND2 (N3711, N3697, N568);
nand NAND3 (N3712, N3704, N693, N374);
xor XOR2 (N3713, N3707, N3026);
and AND3 (N3714, N3708, N3103, N2074);
xor XOR2 (N3715, N3710, N110);
or OR2 (N3716, N3713, N433);
nand NAND2 (N3717, N3716, N952);
and AND3 (N3718, N3715, N565, N2312);
nor NOR2 (N3719, N3711, N73);
not NOT1 (N3720, N3689);
buf BUF1 (N3721, N3718);
buf BUF1 (N3722, N3714);
and AND4 (N3723, N3722, N2683, N1745, N3078);
xor XOR2 (N3724, N3712, N1658);
nor NOR3 (N3725, N3723, N1591, N815);
xor XOR2 (N3726, N3702, N2532);
buf BUF1 (N3727, N3721);
nor NOR4 (N3728, N3698, N997, N2681, N188);
nor NOR2 (N3729, N3724, N1839);
and AND3 (N3730, N3727, N283, N3645);
nor NOR4 (N3731, N3717, N3647, N2912, N515);
not NOT1 (N3732, N3725);
or OR3 (N3733, N3728, N635, N2881);
buf BUF1 (N3734, N3726);
and AND2 (N3735, N3734, N1179);
nor NOR3 (N3736, N3731, N429, N983);
xor XOR2 (N3737, N3730, N866);
nand NAND4 (N3738, N3729, N1475, N2715, N136);
and AND4 (N3739, N3737, N1540, N2024, N3033);
or OR2 (N3740, N3735, N3296);
nand NAND3 (N3741, N3740, N911, N3488);
and AND3 (N3742, N3732, N920, N3030);
or OR4 (N3743, N3688, N3472, N1270, N3527);
nor NOR4 (N3744, N3741, N1112, N2850, N520);
not NOT1 (N3745, N3743);
nand NAND4 (N3746, N3745, N1767, N1659, N1915);
nand NAND2 (N3747, N3733, N2965);
or OR4 (N3748, N3747, N1181, N984, N1017);
buf BUF1 (N3749, N3742);
buf BUF1 (N3750, N3719);
or OR3 (N3751, N3736, N2381, N3041);
nand NAND3 (N3752, N3746, N1414, N1445);
nand NAND2 (N3753, N3720, N32);
and AND3 (N3754, N3739, N517, N38);
not NOT1 (N3755, N3749);
or OR2 (N3756, N3744, N3258);
and AND2 (N3757, N3753, N191);
nand NAND4 (N3758, N3755, N1463, N1738, N3266);
or OR4 (N3759, N3758, N1780, N1696, N1101);
xor XOR2 (N3760, N3757, N3593);
nand NAND2 (N3761, N3756, N2369);
and AND2 (N3762, N3754, N1068);
or OR3 (N3763, N3759, N2664, N345);
and AND3 (N3764, N3751, N2650, N3678);
nor NOR4 (N3765, N3762, N3121, N861, N1381);
nor NOR3 (N3766, N3750, N2302, N1508);
xor XOR2 (N3767, N3763, N634);
nand NAND4 (N3768, N3761, N1062, N1526, N1088);
or OR2 (N3769, N3764, N402);
nor NOR2 (N3770, N3748, N1999);
buf BUF1 (N3771, N3760);
nand NAND2 (N3772, N3738, N3745);
nor NOR3 (N3773, N3752, N2321, N1390);
xor XOR2 (N3774, N3706, N2042);
not NOT1 (N3775, N3766);
or OR2 (N3776, N3765, N281);
buf BUF1 (N3777, N3770);
not NOT1 (N3778, N3777);
nor NOR4 (N3779, N3769, N1197, N315, N2756);
or OR2 (N3780, N3775, N1633);
nand NAND2 (N3781, N3779, N2557);
buf BUF1 (N3782, N3767);
and AND3 (N3783, N3780, N991, N938);
not NOT1 (N3784, N3783);
xor XOR2 (N3785, N3778, N2519);
or OR3 (N3786, N3781, N716, N2524);
not NOT1 (N3787, N3786);
or OR4 (N3788, N3784, N490, N3228, N3376);
nor NOR4 (N3789, N3774, N210, N2909, N3720);
nor NOR2 (N3790, N3787, N940);
or OR3 (N3791, N3771, N1334, N1318);
nand NAND4 (N3792, N3776, N2108, N1773, N1177);
not NOT1 (N3793, N3788);
and AND4 (N3794, N3791, N930, N2107, N2274);
or OR2 (N3795, N3768, N989);
nor NOR3 (N3796, N3790, N2385, N2441);
or OR3 (N3797, N3785, N2183, N945);
xor XOR2 (N3798, N3773, N2068);
buf BUF1 (N3799, N3795);
and AND2 (N3800, N3797, N494);
nor NOR2 (N3801, N3792, N3238);
or OR3 (N3802, N3798, N1093, N750);
buf BUF1 (N3803, N3799);
nor NOR3 (N3804, N3789, N1691, N2482);
nor NOR3 (N3805, N3802, N2041, N1457);
xor XOR2 (N3806, N3782, N3570);
not NOT1 (N3807, N3801);
not NOT1 (N3808, N3804);
or OR2 (N3809, N3800, N3742);
xor XOR2 (N3810, N3796, N1673);
buf BUF1 (N3811, N3793);
nor NOR4 (N3812, N3805, N643, N68, N2191);
xor XOR2 (N3813, N3808, N103);
or OR4 (N3814, N3809, N2691, N1297, N1452);
or OR3 (N3815, N3794, N1898, N742);
nor NOR3 (N3816, N3810, N3113, N2311);
nor NOR4 (N3817, N3811, N3300, N3640, N612);
nand NAND2 (N3818, N3812, N2235);
nand NAND4 (N3819, N3817, N1369, N226, N2420);
buf BUF1 (N3820, N3806);
nand NAND4 (N3821, N3803, N1239, N2337, N876);
and AND4 (N3822, N3820, N3802, N3388, N3794);
not NOT1 (N3823, N3772);
nor NOR4 (N3824, N3819, N1416, N3383, N1865);
not NOT1 (N3825, N3813);
buf BUF1 (N3826, N3807);
buf BUF1 (N3827, N3825);
not NOT1 (N3828, N3818);
not NOT1 (N3829, N3823);
and AND4 (N3830, N3822, N326, N2525, N999);
xor XOR2 (N3831, N3816, N3483);
and AND2 (N3832, N3830, N1254);
and AND2 (N3833, N3824, N3037);
nor NOR3 (N3834, N3827, N3226, N2800);
and AND4 (N3835, N3814, N1167, N3578, N2754);
and AND2 (N3836, N3832, N3591);
nand NAND4 (N3837, N3821, N3082, N3261, N1850);
or OR4 (N3838, N3834, N2897, N688, N3381);
xor XOR2 (N3839, N3826, N2353);
and AND2 (N3840, N3833, N1939);
and AND2 (N3841, N3837, N3242);
or OR3 (N3842, N3841, N3368, N833);
and AND2 (N3843, N3831, N3110);
or OR2 (N3844, N3842, N1676);
xor XOR2 (N3845, N3840, N2817);
nor NOR2 (N3846, N3838, N1771);
and AND2 (N3847, N3836, N1680);
and AND3 (N3848, N3839, N223, N2571);
nor NOR4 (N3849, N3815, N2005, N1225, N3410);
buf BUF1 (N3850, N3835);
not NOT1 (N3851, N3849);
buf BUF1 (N3852, N3844);
buf BUF1 (N3853, N3845);
xor XOR2 (N3854, N3828, N1094);
or OR3 (N3855, N3847, N25, N684);
nand NAND2 (N3856, N3846, N685);
and AND3 (N3857, N3856, N2282, N2034);
nand NAND4 (N3858, N3851, N2591, N2269, N1008);
xor XOR2 (N3859, N3853, N700);
xor XOR2 (N3860, N3843, N2621);
or OR4 (N3861, N3848, N92, N2935, N3188);
nor NOR4 (N3862, N3858, N2253, N911, N3410);
nor NOR2 (N3863, N3850, N2741);
nor NOR2 (N3864, N3857, N2158);
xor XOR2 (N3865, N3860, N259);
buf BUF1 (N3866, N3865);
not NOT1 (N3867, N3859);
xor XOR2 (N3868, N3866, N985);
or OR2 (N3869, N3868, N1782);
xor XOR2 (N3870, N3855, N837);
and AND3 (N3871, N3861, N2661, N1712);
nand NAND4 (N3872, N3852, N2409, N2682, N1396);
nand NAND2 (N3873, N3829, N1744);
xor XOR2 (N3874, N3869, N3107);
nor NOR3 (N3875, N3854, N2947, N3376);
not NOT1 (N3876, N3862);
and AND2 (N3877, N3874, N3566);
nor NOR2 (N3878, N3864, N3224);
not NOT1 (N3879, N3877);
xor XOR2 (N3880, N3871, N1913);
nand NAND3 (N3881, N3875, N608, N761);
nor NOR2 (N3882, N3863, N1853);
buf BUF1 (N3883, N3870);
or OR4 (N3884, N3876, N419, N813, N1386);
or OR3 (N3885, N3878, N1507, N2664);
nand NAND4 (N3886, N3879, N2077, N824, N2853);
nand NAND2 (N3887, N3885, N3003);
nand NAND2 (N3888, N3881, N193);
not NOT1 (N3889, N3883);
not NOT1 (N3890, N3882);
or OR3 (N3891, N3873, N2750, N3352);
buf BUF1 (N3892, N3888);
buf BUF1 (N3893, N3890);
or OR4 (N3894, N3867, N1754, N2067, N2712);
nor NOR2 (N3895, N3886, N3412);
or OR3 (N3896, N3880, N2011, N3454);
xor XOR2 (N3897, N3891, N3516);
not NOT1 (N3898, N3872);
nor NOR3 (N3899, N3893, N220, N3186);
buf BUF1 (N3900, N3887);
not NOT1 (N3901, N3892);
nor NOR4 (N3902, N3894, N363, N2900, N760);
xor XOR2 (N3903, N3884, N2420);
nor NOR2 (N3904, N3896, N314);
or OR4 (N3905, N3900, N358, N3771, N1579);
xor XOR2 (N3906, N3899, N3047);
xor XOR2 (N3907, N3906, N333);
and AND2 (N3908, N3902, N2420);
not NOT1 (N3909, N3901);
nand NAND2 (N3910, N3908, N860);
buf BUF1 (N3911, N3889);
not NOT1 (N3912, N3909);
xor XOR2 (N3913, N3898, N52);
nand NAND2 (N3914, N3897, N3176);
not NOT1 (N3915, N3903);
nor NOR2 (N3916, N3915, N3390);
and AND4 (N3917, N3907, N947, N2968, N1840);
nand NAND4 (N3918, N3910, N3430, N1517, N549);
or OR4 (N3919, N3905, N3452, N756, N3121);
nor NOR3 (N3920, N3904, N388, N732);
xor XOR2 (N3921, N3914, N990);
and AND2 (N3922, N3913, N3661);
nor NOR4 (N3923, N3919, N1345, N3870, N2497);
not NOT1 (N3924, N3911);
buf BUF1 (N3925, N3912);
and AND4 (N3926, N3923, N1215, N2363, N3006);
nand NAND4 (N3927, N3918, N303, N3461, N851);
or OR2 (N3928, N3925, N1955);
and AND3 (N3929, N3926, N2387, N343);
not NOT1 (N3930, N3928);
or OR4 (N3931, N3924, N3643, N1890, N2132);
nor NOR3 (N3932, N3931, N3701, N1423);
nand NAND4 (N3933, N3921, N295, N1051, N949);
xor XOR2 (N3934, N3895, N1277);
and AND2 (N3935, N3916, N3446);
nand NAND3 (N3936, N3932, N894, N2977);
buf BUF1 (N3937, N3927);
xor XOR2 (N3938, N3933, N2084);
not NOT1 (N3939, N3920);
not NOT1 (N3940, N3938);
and AND4 (N3941, N3940, N1081, N1407, N2076);
xor XOR2 (N3942, N3935, N370);
and AND4 (N3943, N3922, N1516, N1946, N1945);
nand NAND2 (N3944, N3936, N666);
xor XOR2 (N3945, N3943, N564);
or OR2 (N3946, N3941, N3561);
or OR4 (N3947, N3944, N1544, N3762, N2130);
not NOT1 (N3948, N3930);
and AND4 (N3949, N3948, N1173, N1984, N3298);
xor XOR2 (N3950, N3934, N301);
nor NOR4 (N3951, N3949, N449, N210, N1642);
xor XOR2 (N3952, N3942, N852);
nand NAND2 (N3953, N3946, N196);
not NOT1 (N3954, N3929);
or OR2 (N3955, N3951, N691);
xor XOR2 (N3956, N3955, N1219);
nor NOR4 (N3957, N3950, N1290, N2500, N130);
or OR3 (N3958, N3952, N564, N643);
nand NAND2 (N3959, N3945, N3115);
xor XOR2 (N3960, N3954, N1386);
and AND3 (N3961, N3957, N2438, N305);
nor NOR4 (N3962, N3939, N2444, N2867, N1042);
nor NOR3 (N3963, N3962, N2330, N3639);
and AND3 (N3964, N3959, N561, N3400);
and AND2 (N3965, N3958, N1565);
xor XOR2 (N3966, N3956, N3210);
xor XOR2 (N3967, N3917, N2218);
nand NAND2 (N3968, N3937, N146);
not NOT1 (N3969, N3965);
buf BUF1 (N3970, N3966);
or OR3 (N3971, N3964, N3494, N2119);
not NOT1 (N3972, N3970);
nor NOR2 (N3973, N3972, N1522);
xor XOR2 (N3974, N3947, N3153);
or OR3 (N3975, N3953, N3885, N3668);
nand NAND2 (N3976, N3969, N1023);
or OR4 (N3977, N3975, N127, N966, N315);
buf BUF1 (N3978, N3974);
xor XOR2 (N3979, N3963, N3596);
xor XOR2 (N3980, N3973, N3347);
nor NOR3 (N3981, N3967, N2666, N518);
xor XOR2 (N3982, N3978, N1734);
xor XOR2 (N3983, N3976, N3820);
buf BUF1 (N3984, N3968);
and AND3 (N3985, N3981, N4, N3426);
or OR2 (N3986, N3977, N3227);
xor XOR2 (N3987, N3961, N2561);
not NOT1 (N3988, N3987);
or OR3 (N3989, N3984, N1056, N3819);
not NOT1 (N3990, N3971);
buf BUF1 (N3991, N3980);
and AND3 (N3992, N3990, N72, N2607);
buf BUF1 (N3993, N3991);
not NOT1 (N3994, N3979);
and AND3 (N3995, N3994, N601, N1986);
or OR4 (N3996, N3960, N2523, N1923, N2003);
buf BUF1 (N3997, N3983);
nand NAND3 (N3998, N3993, N3856, N3702);
nor NOR2 (N3999, N3998, N3701);
buf BUF1 (N4000, N3989);
xor XOR2 (N4001, N3997, N595);
not NOT1 (N4002, N3988);
or OR2 (N4003, N3995, N2133);
nand NAND4 (N4004, N3996, N952, N2144, N2221);
and AND2 (N4005, N4003, N2136);
xor XOR2 (N4006, N3992, N294);
nand NAND2 (N4007, N4004, N814);
and AND4 (N4008, N4006, N81, N3410, N321);
nand NAND3 (N4009, N4008, N2531, N2517);
xor XOR2 (N4010, N3982, N3293);
and AND4 (N4011, N3985, N844, N3304, N1636);
and AND3 (N4012, N4000, N3060, N2400);
or OR3 (N4013, N4002, N1150, N3765);
not NOT1 (N4014, N4010);
nand NAND4 (N4015, N4009, N1620, N1935, N2987);
nor NOR3 (N4016, N4007, N3530, N3031);
xor XOR2 (N4017, N4016, N2160);
buf BUF1 (N4018, N4001);
not NOT1 (N4019, N4014);
xor XOR2 (N4020, N4012, N1937);
or OR3 (N4021, N3986, N367, N912);
and AND4 (N4022, N4005, N3888, N2808, N1168);
buf BUF1 (N4023, N4017);
nor NOR4 (N4024, N4015, N1995, N1141, N1217);
xor XOR2 (N4025, N4020, N130);
nor NOR4 (N4026, N4019, N3757, N917, N1846);
not NOT1 (N4027, N4024);
nand NAND4 (N4028, N4013, N2724, N180, N520);
buf BUF1 (N4029, N4028);
and AND4 (N4030, N4021, N1433, N793, N4017);
not NOT1 (N4031, N4011);
buf BUF1 (N4032, N4030);
not NOT1 (N4033, N4029);
xor XOR2 (N4034, N4027, N633);
buf BUF1 (N4035, N4025);
not NOT1 (N4036, N4032);
nand NAND4 (N4037, N4031, N1191, N1279, N1274);
xor XOR2 (N4038, N4036, N3132);
buf BUF1 (N4039, N4037);
or OR3 (N4040, N4022, N3447, N3060);
nor NOR3 (N4041, N4039, N3335, N1341);
not NOT1 (N4042, N4033);
nand NAND2 (N4043, N4041, N1360);
or OR3 (N4044, N4042, N91, N3433);
or OR4 (N4045, N4023, N572, N4040, N3969);
not NOT1 (N4046, N516);
nand NAND4 (N4047, N3999, N298, N1745, N3712);
xor XOR2 (N4048, N4026, N2385);
nor NOR3 (N4049, N4043, N1682, N3767);
buf BUF1 (N4050, N4049);
xor XOR2 (N4051, N4047, N1223);
buf BUF1 (N4052, N4035);
xor XOR2 (N4053, N4050, N2951);
buf BUF1 (N4054, N4038);
buf BUF1 (N4055, N4018);
buf BUF1 (N4056, N4046);
nor NOR2 (N4057, N4048, N3963);
buf BUF1 (N4058, N4044);
nor NOR2 (N4059, N4056, N2768);
not NOT1 (N4060, N4059);
buf BUF1 (N4061, N4055);
buf BUF1 (N4062, N4061);
or OR3 (N4063, N4054, N436, N3315);
nor NOR2 (N4064, N4057, N2563);
or OR3 (N4065, N4060, N10, N2668);
and AND3 (N4066, N4034, N1934, N528);
and AND2 (N4067, N4063, N3799);
nor NOR2 (N4068, N4062, N453);
xor XOR2 (N4069, N4068, N3524);
nand NAND4 (N4070, N4067, N3110, N3705, N198);
buf BUF1 (N4071, N4070);
and AND3 (N4072, N4058, N2156, N2125);
or OR3 (N4073, N4071, N3528, N924);
xor XOR2 (N4074, N4069, N473);
or OR3 (N4075, N4073, N385, N1356);
not NOT1 (N4076, N4066);
buf BUF1 (N4077, N4045);
buf BUF1 (N4078, N4052);
nand NAND4 (N4079, N4051, N2047, N662, N3032);
nor NOR4 (N4080, N4078, N1745, N3504, N1094);
buf BUF1 (N4081, N4072);
xor XOR2 (N4082, N4080, N2150);
not NOT1 (N4083, N4079);
nand NAND4 (N4084, N4077, N2656, N903, N3013);
and AND2 (N4085, N4053, N2933);
or OR2 (N4086, N4081, N1973);
nand NAND4 (N4087, N4086, N773, N3371, N1088);
and AND3 (N4088, N4084, N1217, N2664);
or OR3 (N4089, N4075, N110, N417);
buf BUF1 (N4090, N4064);
and AND2 (N4091, N4083, N75);
or OR4 (N4092, N4088, N1196, N3333, N220);
nor NOR2 (N4093, N4074, N2885);
not NOT1 (N4094, N4089);
and AND3 (N4095, N4094, N1104, N3590);
and AND2 (N4096, N4082, N2330);
not NOT1 (N4097, N4076);
or OR2 (N4098, N4093, N1112);
or OR3 (N4099, N4091, N3691, N2126);
nand NAND3 (N4100, N4097, N3545, N1892);
or OR3 (N4101, N4096, N2572, N2484);
xor XOR2 (N4102, N4099, N2662);
not NOT1 (N4103, N4065);
nor NOR2 (N4104, N4090, N2821);
nor NOR4 (N4105, N4085, N931, N1592, N948);
nor NOR4 (N4106, N4100, N791, N3892, N3081);
xor XOR2 (N4107, N4106, N2447);
nand NAND4 (N4108, N4098, N351, N382, N3097);
not NOT1 (N4109, N4104);
nand NAND4 (N4110, N4103, N3523, N1556, N676);
nand NAND2 (N4111, N4087, N3798);
nand NAND4 (N4112, N4108, N1768, N609, N1898);
or OR2 (N4113, N4111, N3792);
xor XOR2 (N4114, N4102, N3627);
nor NOR4 (N4115, N4110, N3766, N3853, N1925);
nor NOR3 (N4116, N4115, N1872, N2444);
or OR4 (N4117, N4114, N1292, N3665, N2336);
and AND3 (N4118, N4113, N898, N2174);
nor NOR2 (N4119, N4095, N2439);
nand NAND3 (N4120, N4105, N3326, N3128);
nor NOR3 (N4121, N4109, N3964, N3586);
xor XOR2 (N4122, N4107, N1304);
buf BUF1 (N4123, N4118);
nand NAND4 (N4124, N4120, N3117, N3633, N2869);
and AND3 (N4125, N4123, N3255, N241);
and AND3 (N4126, N4122, N3743, N1387);
xor XOR2 (N4127, N4121, N629);
buf BUF1 (N4128, N4116);
or OR2 (N4129, N4125, N1072);
and AND2 (N4130, N4117, N3610);
and AND4 (N4131, N4129, N565, N658, N567);
xor XOR2 (N4132, N4126, N3380);
or OR3 (N4133, N4119, N88, N1412);
not NOT1 (N4134, N4124);
buf BUF1 (N4135, N4128);
nand NAND3 (N4136, N4101, N137, N1224);
or OR2 (N4137, N4092, N472);
or OR3 (N4138, N4130, N3281, N3924);
buf BUF1 (N4139, N4133);
xor XOR2 (N4140, N4112, N3884);
nor NOR4 (N4141, N4127, N2038, N574, N3252);
buf BUF1 (N4142, N4140);
nor NOR4 (N4143, N4137, N1819, N2451, N1915);
nand NAND2 (N4144, N4139, N589);
and AND2 (N4145, N4136, N2503);
not NOT1 (N4146, N4144);
not NOT1 (N4147, N4138);
nand NAND4 (N4148, N4131, N2330, N1592, N2230);
xor XOR2 (N4149, N4132, N935);
not NOT1 (N4150, N4142);
buf BUF1 (N4151, N4143);
not NOT1 (N4152, N4151);
buf BUF1 (N4153, N4135);
nand NAND4 (N4154, N4146, N2712, N3072, N2247);
nor NOR4 (N4155, N4141, N905, N419, N1069);
not NOT1 (N4156, N4149);
and AND2 (N4157, N4134, N125);
not NOT1 (N4158, N4154);
or OR4 (N4159, N4145, N539, N748, N3052);
buf BUF1 (N4160, N4156);
and AND4 (N4161, N4160, N963, N1567, N1776);
xor XOR2 (N4162, N4155, N2608);
buf BUF1 (N4163, N4153);
not NOT1 (N4164, N4152);
buf BUF1 (N4165, N4162);
and AND2 (N4166, N4164, N234);
buf BUF1 (N4167, N4150);
xor XOR2 (N4168, N4161, N2201);
not NOT1 (N4169, N4163);
nor NOR3 (N4170, N4157, N155, N3095);
not NOT1 (N4171, N4158);
buf BUF1 (N4172, N4147);
not NOT1 (N4173, N4169);
xor XOR2 (N4174, N4159, N1622);
buf BUF1 (N4175, N4165);
and AND4 (N4176, N4175, N410, N2597, N788);
nand NAND2 (N4177, N4167, N2437);
nor NOR2 (N4178, N4148, N2003);
not NOT1 (N4179, N4170);
nor NOR3 (N4180, N4176, N2425, N3217);
nand NAND4 (N4181, N4168, N2822, N2651, N2809);
not NOT1 (N4182, N4173);
not NOT1 (N4183, N4180);
not NOT1 (N4184, N4171);
not NOT1 (N4185, N4174);
not NOT1 (N4186, N4181);
nor NOR2 (N4187, N4182, N11);
buf BUF1 (N4188, N4166);
or OR2 (N4189, N4178, N713);
buf BUF1 (N4190, N4187);
xor XOR2 (N4191, N4179, N1429);
and AND3 (N4192, N4190, N3761, N443);
nor NOR2 (N4193, N4188, N2904);
not NOT1 (N4194, N4191);
and AND2 (N4195, N4192, N2036);
not NOT1 (N4196, N4172);
or OR2 (N4197, N4189, N3746);
or OR4 (N4198, N4197, N2945, N1025, N3116);
xor XOR2 (N4199, N4184, N2836);
or OR3 (N4200, N4198, N3051, N147);
nor NOR3 (N4201, N4199, N1970, N194);
nand NAND4 (N4202, N4201, N2234, N2695, N1382);
not NOT1 (N4203, N4193);
and AND4 (N4204, N4185, N642, N1979, N1141);
and AND2 (N4205, N4183, N3063);
xor XOR2 (N4206, N4195, N3189);
xor XOR2 (N4207, N4205, N1026);
nand NAND2 (N4208, N4206, N434);
buf BUF1 (N4209, N4207);
buf BUF1 (N4210, N4196);
xor XOR2 (N4211, N4177, N2866);
buf BUF1 (N4212, N4194);
and AND4 (N4213, N4204, N140, N821, N509);
and AND4 (N4214, N4202, N1283, N3716, N2336);
xor XOR2 (N4215, N4203, N356);
not NOT1 (N4216, N4208);
not NOT1 (N4217, N4186);
and AND3 (N4218, N4200, N2739, N1752);
buf BUF1 (N4219, N4209);
nand NAND2 (N4220, N4219, N3419);
or OR2 (N4221, N4218, N2411);
and AND3 (N4222, N4220, N469, N2126);
not NOT1 (N4223, N4211);
xor XOR2 (N4224, N4223, N2092);
buf BUF1 (N4225, N4216);
or OR4 (N4226, N4213, N486, N1425, N3623);
or OR3 (N4227, N4226, N739, N2911);
nand NAND4 (N4228, N4225, N1838, N1457, N3401);
not NOT1 (N4229, N4212);
and AND3 (N4230, N4210, N1972, N921);
nand NAND2 (N4231, N4228, N238);
nand NAND2 (N4232, N4227, N1058);
and AND3 (N4233, N4230, N903, N434);
and AND2 (N4234, N4224, N1212);
xor XOR2 (N4235, N4231, N4182);
nor NOR3 (N4236, N4215, N2592, N1769);
buf BUF1 (N4237, N4229);
not NOT1 (N4238, N4217);
nor NOR2 (N4239, N4237, N1454);
or OR3 (N4240, N4233, N3165, N2417);
xor XOR2 (N4241, N4234, N1346);
nor NOR2 (N4242, N4240, N2616);
xor XOR2 (N4243, N4239, N4217);
not NOT1 (N4244, N4236);
not NOT1 (N4245, N4242);
buf BUF1 (N4246, N4232);
not NOT1 (N4247, N4246);
nand NAND4 (N4248, N4238, N1858, N2874, N2285);
xor XOR2 (N4249, N4245, N3196);
buf BUF1 (N4250, N4247);
xor XOR2 (N4251, N4235, N3412);
xor XOR2 (N4252, N4221, N3835);
nand NAND4 (N4253, N4250, N211, N3057, N3691);
nor NOR3 (N4254, N4244, N1513, N359);
buf BUF1 (N4255, N4251);
buf BUF1 (N4256, N4252);
nor NOR2 (N4257, N4222, N3515);
or OR4 (N4258, N4248, N1114, N4213, N3780);
not NOT1 (N4259, N4258);
not NOT1 (N4260, N4259);
xor XOR2 (N4261, N4254, N1692);
not NOT1 (N4262, N4255);
buf BUF1 (N4263, N4243);
not NOT1 (N4264, N4261);
nand NAND3 (N4265, N4256, N2839, N778);
nor NOR2 (N4266, N4264, N424);
and AND4 (N4267, N4241, N1187, N623, N823);
and AND2 (N4268, N4266, N3001);
or OR3 (N4269, N4257, N1552, N563);
buf BUF1 (N4270, N4263);
nor NOR2 (N4271, N4269, N816);
buf BUF1 (N4272, N4249);
or OR2 (N4273, N4265, N2925);
buf BUF1 (N4274, N4253);
nand NAND4 (N4275, N4272, N4187, N4161, N1674);
and AND3 (N4276, N4271, N1393, N2248);
xor XOR2 (N4277, N4275, N2152);
nand NAND3 (N4278, N4277, N2514, N1371);
nor NOR4 (N4279, N4278, N3919, N2322, N2623);
not NOT1 (N4280, N4273);
nand NAND3 (N4281, N4214, N4030, N3465);
and AND4 (N4282, N4279, N2500, N2584, N4139);
xor XOR2 (N4283, N4274, N2985);
not NOT1 (N4284, N4282);
nor NOR4 (N4285, N4283, N2770, N3951, N3963);
buf BUF1 (N4286, N4284);
nor NOR4 (N4287, N4281, N3576, N1544, N1400);
not NOT1 (N4288, N4286);
not NOT1 (N4289, N4268);
nor NOR4 (N4290, N4280, N3960, N835, N3883);
xor XOR2 (N4291, N4262, N3179);
buf BUF1 (N4292, N4260);
xor XOR2 (N4293, N4287, N3230);
nor NOR2 (N4294, N4285, N2504);
or OR3 (N4295, N4267, N4243, N1559);
nand NAND2 (N4296, N4276, N291);
not NOT1 (N4297, N4292);
nand NAND2 (N4298, N4291, N126);
and AND3 (N4299, N4270, N3880, N530);
or OR3 (N4300, N4293, N2649, N2742);
nand NAND3 (N4301, N4299, N4047, N4246);
nand NAND2 (N4302, N4300, N3680);
xor XOR2 (N4303, N4294, N3865);
or OR4 (N4304, N4303, N891, N757, N694);
and AND2 (N4305, N4302, N3627);
xor XOR2 (N4306, N4295, N1887);
not NOT1 (N4307, N4296);
nand NAND2 (N4308, N4304, N535);
and AND2 (N4309, N4301, N2823);
nor NOR2 (N4310, N4306, N3221);
and AND2 (N4311, N4297, N2898);
buf BUF1 (N4312, N4288);
buf BUF1 (N4313, N4305);
xor XOR2 (N4314, N4310, N595);
nor NOR4 (N4315, N4312, N3479, N1549, N3741);
nor NOR3 (N4316, N4311, N2783, N97);
or OR2 (N4317, N4316, N3820);
xor XOR2 (N4318, N4289, N3093);
not NOT1 (N4319, N4317);
or OR2 (N4320, N4319, N2589);
xor XOR2 (N4321, N4308, N3307);
and AND3 (N4322, N4298, N1190, N1);
xor XOR2 (N4323, N4318, N1364);
not NOT1 (N4324, N4323);
buf BUF1 (N4325, N4290);
nand NAND4 (N4326, N4309, N1499, N3659, N2631);
not NOT1 (N4327, N4320);
and AND3 (N4328, N4321, N1604, N1748);
nor NOR3 (N4329, N4314, N1308, N690);
nand NAND2 (N4330, N4328, N1958);
not NOT1 (N4331, N4326);
buf BUF1 (N4332, N4327);
or OR2 (N4333, N4332, N1744);
or OR3 (N4334, N4322, N1370, N534);
xor XOR2 (N4335, N4307, N3683);
and AND3 (N4336, N4315, N1053, N2745);
buf BUF1 (N4337, N4331);
nor NOR3 (N4338, N4324, N194, N3145);
not NOT1 (N4339, N4330);
xor XOR2 (N4340, N4335, N2743);
not NOT1 (N4341, N4334);
buf BUF1 (N4342, N4339);
or OR2 (N4343, N4340, N4094);
or OR2 (N4344, N4341, N309);
nor NOR4 (N4345, N4329, N3351, N482, N1214);
nand NAND4 (N4346, N4333, N3463, N114, N1564);
buf BUF1 (N4347, N4337);
nand NAND4 (N4348, N4313, N1150, N2142, N3074);
and AND3 (N4349, N4344, N1231, N1976);
and AND3 (N4350, N4342, N1994, N3131);
nor NOR2 (N4351, N4348, N349);
buf BUF1 (N4352, N4351);
nand NAND4 (N4353, N4349, N2881, N200, N157);
or OR4 (N4354, N4325, N2992, N3091, N3624);
and AND3 (N4355, N4336, N4076, N3779);
and AND4 (N4356, N4355, N1166, N115, N538);
or OR4 (N4357, N4352, N1332, N1595, N692);
nand NAND3 (N4358, N4343, N4155, N4149);
nand NAND4 (N4359, N4346, N430, N2658, N734);
buf BUF1 (N4360, N4338);
buf BUF1 (N4361, N4347);
or OR2 (N4362, N4345, N3645);
or OR2 (N4363, N4360, N186);
and AND2 (N4364, N4350, N1973);
buf BUF1 (N4365, N4361);
or OR2 (N4366, N4358, N3924);
and AND4 (N4367, N4363, N2300, N3024, N332);
nand NAND2 (N4368, N4357, N2544);
not NOT1 (N4369, N4354);
or OR2 (N4370, N4364, N2229);
not NOT1 (N4371, N4370);
and AND2 (N4372, N4359, N2527);
xor XOR2 (N4373, N4362, N578);
xor XOR2 (N4374, N4353, N2973);
xor XOR2 (N4375, N4367, N3458);
not NOT1 (N4376, N4369);
not NOT1 (N4377, N4371);
buf BUF1 (N4378, N4356);
or OR3 (N4379, N4376, N1335, N737);
nor NOR3 (N4380, N4377, N3009, N3496);
and AND2 (N4381, N4375, N1812);
nor NOR3 (N4382, N4379, N4242, N1324);
nor NOR3 (N4383, N4372, N611, N3912);
nor NOR4 (N4384, N4382, N3595, N2952, N3229);
or OR2 (N4385, N4378, N672);
and AND2 (N4386, N4381, N3925);
or OR2 (N4387, N4385, N135);
xor XOR2 (N4388, N4387, N2486);
nor NOR2 (N4389, N4383, N3842);
nor NOR3 (N4390, N4384, N2413, N2141);
or OR4 (N4391, N4389, N2502, N1693, N2854);
nor NOR4 (N4392, N4391, N2517, N2247, N3414);
and AND3 (N4393, N4390, N1952, N3946);
not NOT1 (N4394, N4386);
buf BUF1 (N4395, N4365);
nand NAND2 (N4396, N4373, N2330);
nor NOR4 (N4397, N4374, N3799, N4237, N3841);
not NOT1 (N4398, N4393);
not NOT1 (N4399, N4366);
nand NAND2 (N4400, N4399, N10);
not NOT1 (N4401, N4394);
or OR3 (N4402, N4380, N745, N2078);
not NOT1 (N4403, N4401);
or OR3 (N4404, N4398, N1219, N978);
and AND2 (N4405, N4403, N1703);
and AND2 (N4406, N4368, N2519);
nand NAND3 (N4407, N4404, N4053, N3366);
nand NAND4 (N4408, N4400, N1350, N4237, N999);
and AND3 (N4409, N4397, N2948, N2740);
nand NAND3 (N4410, N4402, N867, N1271);
nor NOR2 (N4411, N4405, N1249);
buf BUF1 (N4412, N4406);
and AND3 (N4413, N4392, N1331, N2880);
and AND2 (N4414, N4409, N1602);
and AND4 (N4415, N4411, N1132, N2518, N2023);
or OR4 (N4416, N4407, N1667, N964, N3282);
buf BUF1 (N4417, N4414);
not NOT1 (N4418, N4395);
nand NAND2 (N4419, N4418, N41);
nand NAND3 (N4420, N4413, N222, N1036);
nor NOR4 (N4421, N4396, N3681, N635, N3157);
not NOT1 (N4422, N4412);
nor NOR3 (N4423, N4416, N1059, N1775);
nand NAND3 (N4424, N4417, N2238, N1645);
or OR4 (N4425, N4424, N3776, N745, N1753);
not NOT1 (N4426, N4388);
nor NOR4 (N4427, N4420, N1406, N4092, N3340);
nor NOR4 (N4428, N4422, N2367, N2286, N798);
nor NOR3 (N4429, N4408, N3849, N2239);
nand NAND2 (N4430, N4428, N3614);
nor NOR3 (N4431, N4421, N3349, N2522);
nand NAND4 (N4432, N4427, N1997, N4334, N2142);
nand NAND2 (N4433, N4425, N161);
buf BUF1 (N4434, N4433);
not NOT1 (N4435, N4415);
nor NOR2 (N4436, N4423, N1524);
nor NOR3 (N4437, N4435, N460, N820);
nor NOR3 (N4438, N4410, N4430, N4401);
buf BUF1 (N4439, N2323);
nor NOR2 (N4440, N4437, N4291);
nor NOR3 (N4441, N4434, N3033, N405);
xor XOR2 (N4442, N4438, N2528);
not NOT1 (N4443, N4441);
not NOT1 (N4444, N4443);
not NOT1 (N4445, N4439);
not NOT1 (N4446, N4444);
or OR2 (N4447, N4432, N3663);
buf BUF1 (N4448, N4436);
or OR3 (N4449, N4446, N4268, N2369);
or OR2 (N4450, N4447, N3858);
and AND3 (N4451, N4449, N4146, N2430);
xor XOR2 (N4452, N4451, N2547);
not NOT1 (N4453, N4452);
or OR2 (N4454, N4431, N2741);
buf BUF1 (N4455, N4448);
xor XOR2 (N4456, N4442, N4135);
and AND3 (N4457, N4419, N3005, N3656);
xor XOR2 (N4458, N4429, N749);
nand NAND4 (N4459, N4445, N730, N3951, N2192);
or OR2 (N4460, N4454, N3627);
xor XOR2 (N4461, N4460, N693);
not NOT1 (N4462, N4453);
xor XOR2 (N4463, N4440, N2199);
nor NOR2 (N4464, N4455, N1211);
nand NAND3 (N4465, N4426, N4044, N2210);
xor XOR2 (N4466, N4464, N2337);
xor XOR2 (N4467, N4457, N1686);
not NOT1 (N4468, N4462);
buf BUF1 (N4469, N4465);
or OR4 (N4470, N4456, N3358, N651, N2626);
nor NOR3 (N4471, N4466, N3039, N3694);
nor NOR4 (N4472, N4450, N92, N3468, N1880);
xor XOR2 (N4473, N4468, N3817);
nor NOR3 (N4474, N4472, N3407, N3448);
nor NOR2 (N4475, N4471, N4298);
or OR3 (N4476, N4470, N472, N808);
not NOT1 (N4477, N4469);
buf BUF1 (N4478, N4476);
or OR3 (N4479, N4459, N1045, N2677);
or OR3 (N4480, N4478, N1339, N3208);
xor XOR2 (N4481, N4463, N1265);
and AND3 (N4482, N4480, N2961, N336);
xor XOR2 (N4483, N4475, N1107);
nand NAND2 (N4484, N4483, N3203);
not NOT1 (N4485, N4467);
nor NOR2 (N4486, N4482, N1254);
xor XOR2 (N4487, N4484, N380);
and AND4 (N4488, N4461, N1357, N3808, N2230);
and AND4 (N4489, N4486, N2781, N3809, N3476);
or OR2 (N4490, N4474, N3320);
or OR4 (N4491, N4477, N1449, N500, N2576);
nand NAND2 (N4492, N4479, N886);
not NOT1 (N4493, N4487);
or OR2 (N4494, N4458, N1865);
or OR2 (N4495, N4490, N2444);
and AND4 (N4496, N4481, N2850, N3325, N4240);
nand NAND3 (N4497, N4494, N4161, N1160);
buf BUF1 (N4498, N4497);
or OR2 (N4499, N4496, N3386);
not NOT1 (N4500, N4495);
and AND4 (N4501, N4500, N1497, N4482, N3826);
and AND4 (N4502, N4501, N4112, N1286, N2625);
not NOT1 (N4503, N4485);
nand NAND3 (N4504, N4503, N18, N1810);
nor NOR3 (N4505, N4492, N4232, N1306);
or OR2 (N4506, N4491, N3126);
xor XOR2 (N4507, N4473, N3194);
nand NAND2 (N4508, N4504, N3886);
xor XOR2 (N4509, N4508, N382);
and AND3 (N4510, N4509, N3342, N2501);
or OR2 (N4511, N4507, N279);
or OR3 (N4512, N4488, N2583, N845);
buf BUF1 (N4513, N4510);
or OR2 (N4514, N4489, N3032);
nor NOR2 (N4515, N4499, N455);
not NOT1 (N4516, N4505);
or OR3 (N4517, N4512, N3190, N2205);
nor NOR3 (N4518, N4514, N4497, N2620);
or OR4 (N4519, N4515, N4046, N1915, N1974);
or OR4 (N4520, N4519, N4477, N767, N3728);
xor XOR2 (N4521, N4516, N3031);
and AND3 (N4522, N4520, N980, N207);
nor NOR2 (N4523, N4506, N4390);
or OR2 (N4524, N4502, N1609);
xor XOR2 (N4525, N4521, N1671);
or OR4 (N4526, N4513, N1173, N1393, N555);
buf BUF1 (N4527, N4526);
buf BUF1 (N4528, N4498);
nand NAND4 (N4529, N4525, N136, N511, N3449);
not NOT1 (N4530, N4527);
buf BUF1 (N4531, N4517);
xor XOR2 (N4532, N4530, N3712);
nand NAND4 (N4533, N4518, N1728, N1603, N2406);
or OR2 (N4534, N4511, N2358);
buf BUF1 (N4535, N4533);
xor XOR2 (N4536, N4523, N314);
nor NOR2 (N4537, N4531, N1851);
nor NOR3 (N4538, N4536, N3484, N215);
xor XOR2 (N4539, N4538, N1939);
and AND4 (N4540, N4529, N1754, N3347, N4433);
xor XOR2 (N4541, N4537, N1063);
nor NOR4 (N4542, N4524, N4520, N141, N4094);
nor NOR2 (N4543, N4541, N2442);
not NOT1 (N4544, N4493);
buf BUF1 (N4545, N4534);
and AND2 (N4546, N4535, N2122);
xor XOR2 (N4547, N4542, N2885);
buf BUF1 (N4548, N4547);
nand NAND2 (N4549, N4543, N3402);
nand NAND2 (N4550, N4539, N1366);
nand NAND4 (N4551, N4545, N2695, N2484, N3086);
xor XOR2 (N4552, N4551, N115);
or OR4 (N4553, N4552, N1756, N55, N2137);
not NOT1 (N4554, N4548);
xor XOR2 (N4555, N4544, N3882);
not NOT1 (N4556, N4549);
or OR2 (N4557, N4555, N3205);
nor NOR4 (N4558, N4557, N130, N2670, N66);
nor NOR4 (N4559, N4556, N3175, N1108, N838);
not NOT1 (N4560, N4558);
and AND4 (N4561, N4540, N1134, N2219, N1212);
xor XOR2 (N4562, N4561, N1108);
nand NAND3 (N4563, N4560, N2176, N1258);
and AND3 (N4564, N4559, N3019, N2770);
and AND2 (N4565, N4564, N461);
nor NOR3 (N4566, N4554, N3666, N1946);
nor NOR3 (N4567, N4550, N3179, N4550);
xor XOR2 (N4568, N4522, N1880);
nand NAND4 (N4569, N4566, N1589, N2444, N588);
or OR2 (N4570, N4562, N2968);
not NOT1 (N4571, N4565);
nand NAND2 (N4572, N4563, N2186);
not NOT1 (N4573, N4569);
buf BUF1 (N4574, N4573);
buf BUF1 (N4575, N4572);
nand NAND3 (N4576, N4570, N3023, N734);
or OR3 (N4577, N4571, N4012, N4248);
and AND4 (N4578, N4532, N4168, N304, N1087);
buf BUF1 (N4579, N4567);
or OR3 (N4580, N4577, N4426, N1659);
nor NOR2 (N4581, N4568, N3420);
xor XOR2 (N4582, N4580, N4494);
not NOT1 (N4583, N4581);
buf BUF1 (N4584, N4578);
or OR2 (N4585, N4576, N4345);
nand NAND2 (N4586, N4582, N1917);
or OR4 (N4587, N4553, N3374, N3900, N824);
xor XOR2 (N4588, N4587, N2658);
nand NAND4 (N4589, N4579, N3682, N3707, N2810);
not NOT1 (N4590, N4574);
nor NOR2 (N4591, N4588, N390);
buf BUF1 (N4592, N4528);
or OR4 (N4593, N4589, N2143, N1600, N3048);
buf BUF1 (N4594, N4591);
nand NAND3 (N4595, N4585, N1007, N3105);
buf BUF1 (N4596, N4546);
or OR3 (N4597, N4593, N680, N2176);
nor NOR2 (N4598, N4590, N1254);
nor NOR4 (N4599, N4597, N1181, N3458, N2873);
or OR2 (N4600, N4592, N2320);
xor XOR2 (N4601, N4599, N4395);
xor XOR2 (N4602, N4584, N3719);
xor XOR2 (N4603, N4600, N2545);
and AND4 (N4604, N4575, N1502, N1919, N2554);
nand NAND2 (N4605, N4596, N28);
xor XOR2 (N4606, N4604, N482);
buf BUF1 (N4607, N4601);
nand NAND3 (N4608, N4598, N1284, N1400);
buf BUF1 (N4609, N4583);
and AND2 (N4610, N4603, N122);
not NOT1 (N4611, N4602);
buf BUF1 (N4612, N4608);
not NOT1 (N4613, N4607);
nor NOR4 (N4614, N4606, N2889, N2335, N1512);
not NOT1 (N4615, N4610);
and AND3 (N4616, N4594, N1032, N4020);
and AND4 (N4617, N4605, N1106, N3900, N1786);
xor XOR2 (N4618, N4612, N2085);
or OR2 (N4619, N4617, N3056);
buf BUF1 (N4620, N4616);
and AND4 (N4621, N4595, N1599, N691, N3062);
xor XOR2 (N4622, N4619, N3339);
and AND4 (N4623, N4618, N2155, N1486, N2312);
xor XOR2 (N4624, N4614, N2513);
buf BUF1 (N4625, N4615);
xor XOR2 (N4626, N4622, N1206);
xor XOR2 (N4627, N4624, N3986);
or OR4 (N4628, N4620, N2935, N3700, N2424);
or OR3 (N4629, N4626, N3763, N3538);
nor NOR2 (N4630, N4621, N2633);
xor XOR2 (N4631, N4630, N4173);
not NOT1 (N4632, N4625);
nor NOR4 (N4633, N4632, N3682, N2181, N24);
buf BUF1 (N4634, N4628);
not NOT1 (N4635, N4634);
buf BUF1 (N4636, N4609);
nor NOR4 (N4637, N4629, N4515, N1646, N3440);
nand NAND3 (N4638, N4637, N633, N3279);
buf BUF1 (N4639, N4635);
buf BUF1 (N4640, N4627);
nor NOR3 (N4641, N4638, N3171, N3549);
and AND3 (N4642, N4636, N3939, N3298);
not NOT1 (N4643, N4641);
xor XOR2 (N4644, N4631, N1697);
not NOT1 (N4645, N4644);
xor XOR2 (N4646, N4623, N2883);
not NOT1 (N4647, N4639);
and AND4 (N4648, N4613, N705, N442, N4109);
nand NAND4 (N4649, N4611, N796, N4098, N1555);
and AND4 (N4650, N4648, N2736, N4301, N4475);
xor XOR2 (N4651, N4649, N1744);
xor XOR2 (N4652, N4647, N593);
not NOT1 (N4653, N4642);
nor NOR3 (N4654, N4633, N793, N2519);
nor NOR3 (N4655, N4654, N4100, N536);
not NOT1 (N4656, N4640);
xor XOR2 (N4657, N4645, N2605);
buf BUF1 (N4658, N4650);
not NOT1 (N4659, N4651);
not NOT1 (N4660, N4646);
buf BUF1 (N4661, N4660);
or OR4 (N4662, N4659, N2129, N231, N2418);
xor XOR2 (N4663, N4657, N3997);
and AND3 (N4664, N4656, N3075, N553);
buf BUF1 (N4665, N4662);
xor XOR2 (N4666, N4652, N3097);
and AND4 (N4667, N4655, N3210, N2507, N2344);
nor NOR3 (N4668, N4586, N445, N4382);
xor XOR2 (N4669, N4653, N2981);
xor XOR2 (N4670, N4664, N3950);
nor NOR2 (N4671, N4666, N2580);
nand NAND3 (N4672, N4667, N2977, N2144);
nor NOR4 (N4673, N4670, N4125, N1334, N1927);
buf BUF1 (N4674, N4661);
or OR4 (N4675, N4673, N2706, N1921, N3381);
or OR4 (N4676, N4669, N721, N1627, N110);
nand NAND3 (N4677, N4665, N4392, N1462);
nand NAND2 (N4678, N4676, N3708);
nor NOR4 (N4679, N4663, N2829, N4446, N373);
buf BUF1 (N4680, N4671);
and AND2 (N4681, N4679, N3690);
buf BUF1 (N4682, N4680);
and AND4 (N4683, N4681, N2959, N2717, N2406);
or OR4 (N4684, N4672, N3712, N469, N980);
nor NOR2 (N4685, N4683, N3232);
buf BUF1 (N4686, N4643);
nand NAND2 (N4687, N4674, N1174);
xor XOR2 (N4688, N4658, N763);
or OR4 (N4689, N4688, N3839, N3490, N2133);
and AND4 (N4690, N4684, N4186, N470, N1173);
or OR3 (N4691, N4687, N3693, N2815);
not NOT1 (N4692, N4668);
nor NOR4 (N4693, N4678, N1976, N4485, N1409);
not NOT1 (N4694, N4691);
nand NAND3 (N4695, N4693, N3093, N2156);
and AND3 (N4696, N4695, N3965, N2973);
or OR3 (N4697, N4685, N4648, N4413);
nand NAND4 (N4698, N4697, N3479, N3955, N3357);
or OR2 (N4699, N4690, N3842);
nor NOR3 (N4700, N4675, N2260, N2984);
xor XOR2 (N4701, N4698, N4003);
or OR4 (N4702, N4694, N2327, N554, N3756);
nor NOR4 (N4703, N4677, N2244, N3934, N833);
buf BUF1 (N4704, N4686);
not NOT1 (N4705, N4689);
xor XOR2 (N4706, N4702, N4132);
or OR3 (N4707, N4701, N1967, N4412);
xor XOR2 (N4708, N4699, N1197);
xor XOR2 (N4709, N4706, N3262);
not NOT1 (N4710, N4700);
or OR3 (N4711, N4709, N1869, N1927);
not NOT1 (N4712, N4707);
xor XOR2 (N4713, N4696, N1061);
and AND4 (N4714, N4703, N1519, N802, N4476);
nand NAND2 (N4715, N4714, N2219);
not NOT1 (N4716, N4704);
xor XOR2 (N4717, N4712, N3556);
nor NOR2 (N4718, N4713, N4556);
or OR2 (N4719, N4711, N4224);
nor NOR3 (N4720, N4692, N3693, N4388);
nor NOR4 (N4721, N4708, N1278, N4167, N533);
or OR2 (N4722, N4716, N4396);
buf BUF1 (N4723, N4722);
not NOT1 (N4724, N4720);
or OR2 (N4725, N4723, N3787);
or OR3 (N4726, N4718, N2438, N3580);
or OR4 (N4727, N4705, N1955, N1702, N3582);
and AND3 (N4728, N4727, N329, N4140);
or OR3 (N4729, N4726, N2879, N3026);
buf BUF1 (N4730, N4717);
or OR3 (N4731, N4724, N538, N2971);
buf BUF1 (N4732, N4728);
nor NOR2 (N4733, N4730, N1105);
nor NOR4 (N4734, N4731, N770, N2481, N1923);
xor XOR2 (N4735, N4721, N1445);
nand NAND4 (N4736, N4725, N4494, N4057, N2066);
or OR4 (N4737, N4732, N4404, N4488, N420);
nor NOR2 (N4738, N4736, N3216);
nor NOR3 (N4739, N4682, N2284, N3133);
or OR4 (N4740, N4715, N3352, N4535, N4491);
buf BUF1 (N4741, N4734);
buf BUF1 (N4742, N4741);
or OR3 (N4743, N4710, N1027, N3995);
xor XOR2 (N4744, N4737, N2911);
buf BUF1 (N4745, N4733);
and AND2 (N4746, N4744, N2831);
xor XOR2 (N4747, N4745, N4500);
not NOT1 (N4748, N4739);
nand NAND4 (N4749, N4738, N269, N3095, N2627);
and AND2 (N4750, N4742, N1392);
and AND2 (N4751, N4747, N334);
or OR3 (N4752, N4748, N1385, N1082);
nor NOR2 (N4753, N4719, N1560);
xor XOR2 (N4754, N4750, N2904);
xor XOR2 (N4755, N4735, N1112);
buf BUF1 (N4756, N4753);
nand NAND4 (N4757, N4749, N1253, N3154, N4415);
nor NOR4 (N4758, N4746, N2328, N2123, N721);
or OR4 (N4759, N4752, N1665, N4652, N501);
not NOT1 (N4760, N4754);
buf BUF1 (N4761, N4743);
and AND2 (N4762, N4760, N3383);
and AND2 (N4763, N4761, N132);
and AND2 (N4764, N4763, N2160);
not NOT1 (N4765, N4729);
or OR4 (N4766, N4764, N1589, N924, N1287);
nand NAND4 (N4767, N4751, N3340, N3978, N2383);
nor NOR2 (N4768, N4756, N4167);
nand NAND4 (N4769, N4765, N3263, N246, N3690);
nor NOR4 (N4770, N4768, N4767, N3660, N1129);
or OR2 (N4771, N3416, N1279);
not NOT1 (N4772, N4759);
xor XOR2 (N4773, N4758, N764);
not NOT1 (N4774, N4757);
not NOT1 (N4775, N4774);
not NOT1 (N4776, N4771);
and AND4 (N4777, N4769, N4672, N958, N4500);
not NOT1 (N4778, N4775);
not NOT1 (N4779, N4778);
nor NOR3 (N4780, N4772, N3722, N1049);
and AND3 (N4781, N4776, N2554, N824);
nor NOR4 (N4782, N4773, N308, N3226, N223);
xor XOR2 (N4783, N4779, N883);
nor NOR2 (N4784, N4780, N3647);
not NOT1 (N4785, N4777);
nor NOR3 (N4786, N4770, N875, N4693);
and AND2 (N4787, N4783, N3961);
nand NAND3 (N4788, N4785, N684, N2285);
and AND4 (N4789, N4788, N1465, N3472, N44);
buf BUF1 (N4790, N4789);
and AND4 (N4791, N4787, N4661, N2512, N2606);
not NOT1 (N4792, N4790);
xor XOR2 (N4793, N4755, N4399);
buf BUF1 (N4794, N4781);
nand NAND2 (N4795, N4791, N2076);
buf BUF1 (N4796, N4766);
and AND4 (N4797, N4762, N417, N2768, N975);
nor NOR3 (N4798, N4784, N2204, N86);
xor XOR2 (N4799, N4793, N3456);
or OR4 (N4800, N4786, N3307, N2548, N2607);
not NOT1 (N4801, N4797);
or OR3 (N4802, N4800, N366, N1543);
or OR4 (N4803, N4782, N1823, N4003, N121);
and AND2 (N4804, N4795, N4660);
or OR2 (N4805, N4796, N1645);
nand NAND3 (N4806, N4805, N1764, N1154);
and AND4 (N4807, N4803, N4679, N3175, N3093);
or OR2 (N4808, N4807, N4092);
or OR2 (N4809, N4798, N4092);
and AND2 (N4810, N4802, N662);
and AND2 (N4811, N4808, N3851);
nor NOR4 (N4812, N4809, N4804, N1260, N373);
or OR3 (N4813, N1658, N4018, N1335);
nor NOR2 (N4814, N4813, N2366);
xor XOR2 (N4815, N4801, N137);
and AND2 (N4816, N4806, N1788);
xor XOR2 (N4817, N4794, N4259);
buf BUF1 (N4818, N4816);
buf BUF1 (N4819, N4814);
or OR3 (N4820, N4815, N1672, N2046);
xor XOR2 (N4821, N4811, N3846);
nand NAND2 (N4822, N4817, N1010);
and AND4 (N4823, N4821, N3936, N1478, N4782);
nor NOR3 (N4824, N4820, N123, N3786);
not NOT1 (N4825, N4818);
or OR2 (N4826, N4740, N4018);
not NOT1 (N4827, N4826);
or OR4 (N4828, N4827, N1847, N3665, N575);
or OR2 (N4829, N4812, N4668);
nor NOR2 (N4830, N4824, N2794);
not NOT1 (N4831, N4799);
or OR4 (N4832, N4792, N1486, N1102, N2934);
and AND2 (N4833, N4825, N2547);
xor XOR2 (N4834, N4823, N948);
xor XOR2 (N4835, N4834, N1228);
buf BUF1 (N4836, N4822);
nand NAND4 (N4837, N4833, N1041, N3163, N4092);
not NOT1 (N4838, N4828);
nand NAND4 (N4839, N4830, N2465, N3424, N2402);
or OR2 (N4840, N4831, N2432);
not NOT1 (N4841, N4839);
nor NOR3 (N4842, N4810, N1020, N4722);
nand NAND4 (N4843, N4835, N3117, N4524, N3382);
buf BUF1 (N4844, N4842);
and AND3 (N4845, N4829, N1868, N3934);
and AND4 (N4846, N4840, N3916, N3595, N437);
not NOT1 (N4847, N4845);
not NOT1 (N4848, N4838);
buf BUF1 (N4849, N4847);
buf BUF1 (N4850, N4832);
nand NAND2 (N4851, N4844, N3229);
nand NAND3 (N4852, N4837, N1151, N4432);
not NOT1 (N4853, N4848);
nor NOR2 (N4854, N4849, N1652);
nor NOR4 (N4855, N4854, N2692, N1841, N1307);
nor NOR2 (N4856, N4852, N686);
not NOT1 (N4857, N4853);
and AND4 (N4858, N4843, N706, N2885, N1088);
or OR3 (N4859, N4851, N3801, N2278);
not NOT1 (N4860, N4859);
or OR2 (N4861, N4850, N82);
not NOT1 (N4862, N4857);
xor XOR2 (N4863, N4860, N1011);
and AND2 (N4864, N4858, N2298);
buf BUF1 (N4865, N4864);
buf BUF1 (N4866, N4841);
or OR4 (N4867, N4819, N2612, N1720, N2121);
xor XOR2 (N4868, N4861, N2907);
xor XOR2 (N4869, N4868, N1896);
not NOT1 (N4870, N4846);
or OR3 (N4871, N4863, N4011, N2427);
or OR3 (N4872, N4866, N545, N891);
xor XOR2 (N4873, N4870, N2884);
and AND2 (N4874, N4836, N3039);
nand NAND2 (N4875, N4869, N2461);
nor NOR4 (N4876, N4867, N4004, N570, N2347);
and AND3 (N4877, N4855, N4097, N1612);
buf BUF1 (N4878, N4871);
nand NAND4 (N4879, N4862, N4615, N4577, N245);
not NOT1 (N4880, N4865);
not NOT1 (N4881, N4879);
and AND2 (N4882, N4873, N2971);
nor NOR3 (N4883, N4881, N589, N4630);
not NOT1 (N4884, N4874);
and AND2 (N4885, N4880, N1846);
nand NAND2 (N4886, N4884, N83);
not NOT1 (N4887, N4877);
nand NAND4 (N4888, N4875, N1184, N592, N3775);
nor NOR3 (N4889, N4882, N2950, N1543);
buf BUF1 (N4890, N4889);
nand NAND4 (N4891, N4872, N534, N1936, N4379);
not NOT1 (N4892, N4883);
buf BUF1 (N4893, N4891);
not NOT1 (N4894, N4888);
buf BUF1 (N4895, N4878);
nor NOR4 (N4896, N4886, N2488, N159, N553);
nor NOR4 (N4897, N4893, N4329, N4304, N4885);
nor NOR4 (N4898, N860, N3061, N3597, N1097);
buf BUF1 (N4899, N4898);
xor XOR2 (N4900, N4896, N1158);
buf BUF1 (N4901, N4856);
nor NOR3 (N4902, N4895, N4777, N4670);
not NOT1 (N4903, N4892);
or OR3 (N4904, N4900, N1913, N518);
nand NAND2 (N4905, N4901, N1405);
and AND2 (N4906, N4905, N294);
or OR2 (N4907, N4899, N2970);
and AND2 (N4908, N4897, N4165);
xor XOR2 (N4909, N4902, N2683);
and AND4 (N4910, N4887, N2244, N699, N2558);
and AND4 (N4911, N4894, N2549, N3958, N101);
or OR2 (N4912, N4909, N2591);
xor XOR2 (N4913, N4890, N831);
buf BUF1 (N4914, N4910);
and AND2 (N4915, N4913, N2896);
not NOT1 (N4916, N4908);
buf BUF1 (N4917, N4914);
nor NOR2 (N4918, N4915, N237);
nor NOR4 (N4919, N4911, N4176, N453, N3479);
nor NOR3 (N4920, N4918, N268, N4368);
xor XOR2 (N4921, N4912, N1046);
nor NOR3 (N4922, N4920, N333, N29);
xor XOR2 (N4923, N4917, N1804);
nand NAND2 (N4924, N4907, N2832);
xor XOR2 (N4925, N4919, N2201);
xor XOR2 (N4926, N4921, N4425);
and AND3 (N4927, N4922, N4682, N760);
and AND4 (N4928, N4904, N4595, N4611, N1415);
buf BUF1 (N4929, N4903);
nor NOR2 (N4930, N4927, N2059);
buf BUF1 (N4931, N4928);
nor NOR3 (N4932, N4931, N4485, N4084);
buf BUF1 (N4933, N4916);
and AND4 (N4934, N4929, N4537, N3960, N1429);
or OR3 (N4935, N4923, N3163, N3247);
buf BUF1 (N4936, N4925);
nand NAND4 (N4937, N4936, N4215, N364, N553);
buf BUF1 (N4938, N4937);
nor NOR3 (N4939, N4876, N2663, N2496);
nor NOR2 (N4940, N4935, N3487);
not NOT1 (N4941, N4938);
buf BUF1 (N4942, N4941);
or OR3 (N4943, N4942, N1560, N1910);
not NOT1 (N4944, N4930);
or OR4 (N4945, N4943, N4855, N4858, N4545);
or OR2 (N4946, N4924, N3183);
and AND2 (N4947, N4946, N1065);
xor XOR2 (N4948, N4932, N44);
not NOT1 (N4949, N4939);
buf BUF1 (N4950, N4933);
xor XOR2 (N4951, N4950, N4199);
not NOT1 (N4952, N4944);
buf BUF1 (N4953, N4951);
not NOT1 (N4954, N4906);
or OR4 (N4955, N4952, N2024, N2917, N4244);
nor NOR2 (N4956, N4948, N3586);
nand NAND2 (N4957, N4953, N3098);
xor XOR2 (N4958, N4954, N3937);
not NOT1 (N4959, N4956);
and AND2 (N4960, N4926, N2317);
nand NAND3 (N4961, N4959, N4658, N2593);
nand NAND2 (N4962, N4958, N4875);
buf BUF1 (N4963, N4955);
buf BUF1 (N4964, N4934);
nand NAND3 (N4965, N4963, N3077, N3722);
nand NAND3 (N4966, N4962, N1489, N3634);
not NOT1 (N4967, N4945);
nor NOR3 (N4968, N4961, N965, N630);
xor XOR2 (N4969, N4966, N1650);
or OR2 (N4970, N4968, N2080);
or OR3 (N4971, N4969, N4739, N3353);
xor XOR2 (N4972, N4967, N1222);
nor NOR2 (N4973, N4964, N1367);
buf BUF1 (N4974, N4940);
or OR4 (N4975, N4971, N1888, N4012, N3532);
nor NOR3 (N4976, N4975, N3296, N2199);
not NOT1 (N4977, N4970);
buf BUF1 (N4978, N4949);
xor XOR2 (N4979, N4960, N1337);
nor NOR3 (N4980, N4978, N809, N3715);
buf BUF1 (N4981, N4974);
nand NAND4 (N4982, N4977, N3501, N2270, N3780);
buf BUF1 (N4983, N4957);
nand NAND2 (N4984, N4983, N4624);
not NOT1 (N4985, N4980);
buf BUF1 (N4986, N4972);
nor NOR2 (N4987, N4976, N2639);
and AND4 (N4988, N4965, N2159, N3052, N3505);
and AND2 (N4989, N4982, N3603);
nand NAND2 (N4990, N4979, N4774);
buf BUF1 (N4991, N4987);
and AND3 (N4992, N4984, N3260, N122);
buf BUF1 (N4993, N4985);
nand NAND3 (N4994, N4990, N3397, N2913);
not NOT1 (N4995, N4991);
and AND3 (N4996, N4986, N653, N242);
nand NAND3 (N4997, N4989, N2279, N258);
xor XOR2 (N4998, N4981, N1101);
buf BUF1 (N4999, N4996);
buf BUF1 (N5000, N4992);
not NOT1 (N5001, N5000);
nand NAND3 (N5002, N4988, N2508, N2288);
not NOT1 (N5003, N4993);
not NOT1 (N5004, N4998);
nor NOR4 (N5005, N5002, N369, N1986, N2455);
or OR4 (N5006, N4947, N1379, N134, N4735);
buf BUF1 (N5007, N4973);
nand NAND4 (N5008, N4995, N3661, N1114, N2187);
xor XOR2 (N5009, N5005, N919);
or OR2 (N5010, N5007, N3523);
not NOT1 (N5011, N5009);
or OR4 (N5012, N5003, N4898, N3479, N922);
or OR2 (N5013, N4999, N4884);
not NOT1 (N5014, N4994);
not NOT1 (N5015, N5006);
nor NOR3 (N5016, N5011, N4083, N1682);
nor NOR3 (N5017, N5010, N887, N4033);
xor XOR2 (N5018, N5014, N5015);
not NOT1 (N5019, N3934);
buf BUF1 (N5020, N4997);
buf BUF1 (N5021, N5001);
or OR4 (N5022, N5019, N2784, N112, N2452);
buf BUF1 (N5023, N5017);
and AND2 (N5024, N5016, N1128);
nand NAND3 (N5025, N5020, N385, N4117);
buf BUF1 (N5026, N5024);
nand NAND3 (N5027, N5013, N4654, N3251);
and AND3 (N5028, N5022, N4084, N50);
or OR3 (N5029, N5023, N3385, N432);
nand NAND4 (N5030, N5026, N4210, N31, N4995);
or OR4 (N5031, N5027, N491, N2065, N832);
and AND4 (N5032, N5018, N749, N86, N1813);
and AND3 (N5033, N5028, N353, N1940);
xor XOR2 (N5034, N5033, N829);
not NOT1 (N5035, N5004);
xor XOR2 (N5036, N5008, N2365);
buf BUF1 (N5037, N5032);
nor NOR3 (N5038, N5012, N4172, N4271);
or OR2 (N5039, N5030, N3290);
nor NOR2 (N5040, N5037, N2187);
xor XOR2 (N5041, N5035, N3959);
and AND4 (N5042, N5036, N4430, N4485, N1083);
not NOT1 (N5043, N5039);
not NOT1 (N5044, N5043);
or OR2 (N5045, N5029, N496);
xor XOR2 (N5046, N5044, N4683);
or OR2 (N5047, N5031, N1894);
nor NOR2 (N5048, N5041, N3306);
not NOT1 (N5049, N5047);
or OR4 (N5050, N5049, N1050, N1987, N4466);
or OR3 (N5051, N5048, N623, N4855);
nor NOR4 (N5052, N5034, N622, N3278, N4575);
xor XOR2 (N5053, N5051, N109);
xor XOR2 (N5054, N5025, N3601);
nor NOR4 (N5055, N5054, N4822, N3923, N2562);
or OR4 (N5056, N5053, N3508, N977, N298);
buf BUF1 (N5057, N5040);
not NOT1 (N5058, N5055);
not NOT1 (N5059, N5021);
nor NOR2 (N5060, N5052, N3282);
xor XOR2 (N5061, N5042, N2738);
nand NAND4 (N5062, N5058, N1001, N4834, N4309);
and AND3 (N5063, N5059, N3463, N2968);
and AND3 (N5064, N5057, N327, N2043);
nand NAND4 (N5065, N5045, N991, N2027, N3453);
or OR2 (N5066, N5063, N3726);
or OR3 (N5067, N5060, N2455, N891);
and AND2 (N5068, N5066, N612);
buf BUF1 (N5069, N5038);
or OR2 (N5070, N5050, N2283);
nor NOR4 (N5071, N5046, N3137, N370, N2333);
nand NAND3 (N5072, N5071, N4272, N517);
xor XOR2 (N5073, N5068, N387);
or OR3 (N5074, N5072, N4479, N2254);
nand NAND4 (N5075, N5074, N5044, N2042, N144);
not NOT1 (N5076, N5067);
nor NOR4 (N5077, N5065, N1416, N4893, N4982);
xor XOR2 (N5078, N5077, N1295);
nand NAND4 (N5079, N5056, N2038, N2989, N4945);
and AND4 (N5080, N5073, N1995, N1008, N1809);
not NOT1 (N5081, N5075);
or OR3 (N5082, N5079, N4430, N298);
not NOT1 (N5083, N5081);
nor NOR3 (N5084, N5061, N2237, N2209);
or OR2 (N5085, N5064, N859);
buf BUF1 (N5086, N5070);
and AND4 (N5087, N5069, N1517, N4147, N1066);
nand NAND3 (N5088, N5086, N466, N2331);
nand NAND4 (N5089, N5083, N1337, N3878, N838);
xor XOR2 (N5090, N5078, N1579);
not NOT1 (N5091, N5087);
not NOT1 (N5092, N5084);
and AND4 (N5093, N5080, N1854, N3046, N145);
not NOT1 (N5094, N5082);
nor NOR3 (N5095, N5094, N3393, N595);
and AND2 (N5096, N5090, N1485);
nor NOR3 (N5097, N5096, N2060, N4083);
or OR3 (N5098, N5089, N1746, N723);
and AND2 (N5099, N5088, N4872);
not NOT1 (N5100, N5099);
buf BUF1 (N5101, N5092);
nor NOR4 (N5102, N5093, N1372, N1166, N667);
or OR4 (N5103, N5101, N575, N599, N4774);
xor XOR2 (N5104, N5076, N57);
xor XOR2 (N5105, N5102, N378);
buf BUF1 (N5106, N5100);
nor NOR3 (N5107, N5095, N4534, N4300);
not NOT1 (N5108, N5105);
or OR2 (N5109, N5062, N4072);
nand NAND4 (N5110, N5085, N4346, N4839, N231);
buf BUF1 (N5111, N5110);
xor XOR2 (N5112, N5107, N4529);
buf BUF1 (N5113, N5098);
or OR2 (N5114, N5111, N1455);
nor NOR4 (N5115, N5106, N2474, N1064, N2135);
buf BUF1 (N5116, N5114);
not NOT1 (N5117, N5103);
nor NOR2 (N5118, N5117, N4194);
buf BUF1 (N5119, N5116);
nor NOR3 (N5120, N5109, N1197, N4718);
or OR2 (N5121, N5091, N1248);
nor NOR3 (N5122, N5118, N3625, N1358);
not NOT1 (N5123, N5104);
nor NOR2 (N5124, N5097, N2261);
or OR3 (N5125, N5113, N4606, N3194);
nand NAND4 (N5126, N5112, N3053, N3688, N4322);
or OR4 (N5127, N5123, N2293, N1193, N3339);
nor NOR4 (N5128, N5124, N4873, N4425, N2006);
xor XOR2 (N5129, N5127, N2165);
nand NAND3 (N5130, N5125, N1216, N2504);
not NOT1 (N5131, N5130);
nand NAND4 (N5132, N5121, N57, N1409, N2042);
nand NAND3 (N5133, N5115, N2392, N2768);
nand NAND4 (N5134, N5126, N4009, N185, N694);
and AND4 (N5135, N5131, N1136, N1, N1727);
and AND4 (N5136, N5132, N3693, N2517, N498);
xor XOR2 (N5137, N5136, N4037);
not NOT1 (N5138, N5119);
nand NAND2 (N5139, N5128, N4607);
and AND2 (N5140, N5135, N1837);
nand NAND2 (N5141, N5129, N893);
nand NAND4 (N5142, N5140, N78, N1178, N2788);
nand NAND3 (N5143, N5108, N2044, N1865);
not NOT1 (N5144, N5139);
buf BUF1 (N5145, N5142);
nand NAND2 (N5146, N5122, N3346);
nor NOR3 (N5147, N5137, N2101, N3441);
and AND3 (N5148, N5133, N2962, N1241);
xor XOR2 (N5149, N5147, N3003);
nand NAND4 (N5150, N5149, N5140, N4737, N1881);
buf BUF1 (N5151, N5143);
not NOT1 (N5152, N5120);
not NOT1 (N5153, N5145);
not NOT1 (N5154, N5151);
and AND3 (N5155, N5141, N2501, N4046);
buf BUF1 (N5156, N5148);
xor XOR2 (N5157, N5153, N4572);
nand NAND2 (N5158, N5144, N1060);
nor NOR3 (N5159, N5158, N1437, N3520);
buf BUF1 (N5160, N5155);
xor XOR2 (N5161, N5154, N4553);
xor XOR2 (N5162, N5146, N4142);
and AND2 (N5163, N5134, N3171);
xor XOR2 (N5164, N5162, N3374);
nand NAND2 (N5165, N5160, N3338);
nand NAND4 (N5166, N5164, N2949, N677, N1863);
or OR3 (N5167, N5156, N1596, N3265);
not NOT1 (N5168, N5163);
and AND2 (N5169, N5157, N1706);
or OR2 (N5170, N5165, N3914);
or OR4 (N5171, N5167, N3074, N2251, N188);
not NOT1 (N5172, N5168);
buf BUF1 (N5173, N5171);
buf BUF1 (N5174, N5150);
not NOT1 (N5175, N5174);
not NOT1 (N5176, N5138);
not NOT1 (N5177, N5170);
nand NAND3 (N5178, N5169, N452, N1841);
not NOT1 (N5179, N5161);
or OR4 (N5180, N5152, N3288, N2341, N4985);
nand NAND3 (N5181, N5172, N4383, N4784);
or OR3 (N5182, N5179, N3507, N4017);
nor NOR3 (N5183, N5181, N3414, N4669);
or OR4 (N5184, N5183, N4674, N3560, N3179);
nor NOR3 (N5185, N5176, N2808, N2715);
and AND4 (N5186, N5182, N2124, N1924, N2173);
buf BUF1 (N5187, N5173);
buf BUF1 (N5188, N5175);
nor NOR4 (N5189, N5177, N2595, N1617, N4246);
and AND4 (N5190, N5184, N920, N357, N1415);
and AND2 (N5191, N5188, N1708);
or OR4 (N5192, N5186, N1371, N4418, N3424);
or OR2 (N5193, N5189, N767);
xor XOR2 (N5194, N5178, N4669);
and AND3 (N5195, N5193, N1978, N1980);
xor XOR2 (N5196, N5166, N4962);
buf BUF1 (N5197, N5185);
and AND2 (N5198, N5159, N285);
or OR3 (N5199, N5190, N957, N892);
nor NOR2 (N5200, N5198, N3702);
not NOT1 (N5201, N5187);
nand NAND2 (N5202, N5194, N4239);
xor XOR2 (N5203, N5202, N4775);
or OR3 (N5204, N5196, N2907, N1861);
not NOT1 (N5205, N5204);
nand NAND2 (N5206, N5201, N639);
xor XOR2 (N5207, N5195, N4932);
nor NOR2 (N5208, N5207, N3942);
and AND3 (N5209, N5200, N3654, N2287);
nand NAND4 (N5210, N5199, N2320, N3883, N970);
buf BUF1 (N5211, N5197);
xor XOR2 (N5212, N5180, N4330);
nor NOR2 (N5213, N5209, N4511);
not NOT1 (N5214, N5208);
and AND2 (N5215, N5203, N2071);
or OR4 (N5216, N5211, N2451, N337, N3571);
nor NOR2 (N5217, N5214, N558);
not NOT1 (N5218, N5217);
nand NAND2 (N5219, N5191, N1469);
or OR2 (N5220, N5213, N1034);
nor NOR2 (N5221, N5215, N2647);
buf BUF1 (N5222, N5221);
xor XOR2 (N5223, N5219, N2696);
nand NAND3 (N5224, N5206, N843, N3566);
not NOT1 (N5225, N5222);
nand NAND3 (N5226, N5212, N3137, N3427);
and AND4 (N5227, N5205, N3713, N3543, N1505);
xor XOR2 (N5228, N5227, N1078);
xor XOR2 (N5229, N5228, N100);
nor NOR4 (N5230, N5210, N769, N464, N2097);
nand NAND2 (N5231, N5220, N570);
nor NOR4 (N5232, N5192, N3425, N2243, N2252);
or OR3 (N5233, N5216, N4280, N219);
not NOT1 (N5234, N5233);
nor NOR3 (N5235, N5230, N2174, N5047);
buf BUF1 (N5236, N5223);
and AND4 (N5237, N5224, N5027, N1004, N3516);
buf BUF1 (N5238, N5237);
nor NOR3 (N5239, N5238, N4270, N151);
nand NAND3 (N5240, N5234, N5183, N4314);
and AND4 (N5241, N5236, N4482, N1809, N867);
buf BUF1 (N5242, N5241);
not NOT1 (N5243, N5218);
nor NOR4 (N5244, N5240, N1320, N896, N3393);
buf BUF1 (N5245, N5243);
not NOT1 (N5246, N5244);
buf BUF1 (N5247, N5239);
nand NAND2 (N5248, N5225, N4844);
and AND3 (N5249, N5247, N4174, N3161);
xor XOR2 (N5250, N5229, N1465);
xor XOR2 (N5251, N5231, N2695);
or OR2 (N5252, N5246, N2721);
xor XOR2 (N5253, N5248, N964);
xor XOR2 (N5254, N5232, N3681);
and AND2 (N5255, N5251, N744);
xor XOR2 (N5256, N5252, N2348);
buf BUF1 (N5257, N5255);
and AND4 (N5258, N5250, N4152, N3600, N3516);
nand NAND4 (N5259, N5235, N3878, N1473, N2139);
not NOT1 (N5260, N5245);
not NOT1 (N5261, N5258);
and AND2 (N5262, N5261, N3247);
xor XOR2 (N5263, N5260, N3849);
buf BUF1 (N5264, N5256);
nor NOR3 (N5265, N5263, N1333, N3332);
buf BUF1 (N5266, N5242);
buf BUF1 (N5267, N5259);
nand NAND3 (N5268, N5226, N3757, N2223);
nor NOR3 (N5269, N5268, N3469, N385);
nor NOR4 (N5270, N5266, N4491, N2184, N3975);
nor NOR3 (N5271, N5249, N2526, N2686);
or OR3 (N5272, N5254, N2091, N3498);
xor XOR2 (N5273, N5271, N4375);
nor NOR4 (N5274, N5265, N1710, N1898, N2199);
not NOT1 (N5275, N5270);
or OR4 (N5276, N5267, N1272, N1727, N318);
and AND4 (N5277, N5257, N4504, N3101, N5201);
not NOT1 (N5278, N5275);
nor NOR3 (N5279, N5272, N763, N1649);
xor XOR2 (N5280, N5278, N3121);
nor NOR2 (N5281, N5273, N2569);
or OR2 (N5282, N5280, N1896);
xor XOR2 (N5283, N5262, N1670);
buf BUF1 (N5284, N5283);
and AND2 (N5285, N5269, N2906);
or OR4 (N5286, N5253, N3292, N1497, N3426);
not NOT1 (N5287, N5284);
or OR4 (N5288, N5287, N4825, N775, N1756);
not NOT1 (N5289, N5288);
nor NOR4 (N5290, N5276, N1120, N1330, N1872);
and AND2 (N5291, N5274, N2890);
nand NAND3 (N5292, N5286, N4589, N940);
and AND2 (N5293, N5291, N1997);
nand NAND4 (N5294, N5290, N4985, N2547, N3036);
nor NOR3 (N5295, N5281, N3995, N2248);
not NOT1 (N5296, N5295);
nor NOR4 (N5297, N5282, N3921, N3161, N4778);
nand NAND4 (N5298, N5277, N886, N1434, N4016);
not NOT1 (N5299, N5285);
and AND4 (N5300, N5293, N1597, N1559, N5161);
nand NAND4 (N5301, N5279, N532, N3613, N1879);
buf BUF1 (N5302, N5298);
xor XOR2 (N5303, N5294, N3914);
or OR3 (N5304, N5303, N501, N2839);
nand NAND4 (N5305, N5296, N5112, N2754, N4497);
nand NAND2 (N5306, N5304, N2078);
nor NOR3 (N5307, N5289, N1233, N4444);
nor NOR2 (N5308, N5264, N1250);
and AND2 (N5309, N5305, N678);
nand NAND2 (N5310, N5302, N615);
buf BUF1 (N5311, N5307);
nor NOR3 (N5312, N5309, N2311, N1380);
buf BUF1 (N5313, N5311);
buf BUF1 (N5314, N5313);
nor NOR4 (N5315, N5314, N1932, N459, N748);
nor NOR3 (N5316, N5301, N1536, N3114);
not NOT1 (N5317, N5308);
nand NAND4 (N5318, N5297, N5089, N2477, N4238);
nand NAND4 (N5319, N5317, N2288, N510, N1539);
or OR2 (N5320, N5319, N3485);
xor XOR2 (N5321, N5315, N240);
nor NOR2 (N5322, N5318, N2042);
or OR3 (N5323, N5299, N2958, N2076);
xor XOR2 (N5324, N5306, N2652);
xor XOR2 (N5325, N5292, N2222);
or OR4 (N5326, N5320, N2237, N3963, N3429);
buf BUF1 (N5327, N5323);
nand NAND2 (N5328, N5326, N295);
buf BUF1 (N5329, N5327);
buf BUF1 (N5330, N5300);
nor NOR2 (N5331, N5321, N1940);
and AND4 (N5332, N5324, N1540, N3769, N1009);
nor NOR2 (N5333, N5332, N2550);
or OR4 (N5334, N5330, N2010, N1832, N2795);
and AND3 (N5335, N5329, N1753, N490);
xor XOR2 (N5336, N5310, N1437);
buf BUF1 (N5337, N5322);
buf BUF1 (N5338, N5337);
buf BUF1 (N5339, N5312);
or OR3 (N5340, N5333, N3065, N4905);
xor XOR2 (N5341, N5316, N401);
nor NOR4 (N5342, N5328, N4476, N3237, N5283);
nor NOR3 (N5343, N5336, N4996, N2029);
buf BUF1 (N5344, N5341);
buf BUF1 (N5345, N5340);
or OR3 (N5346, N5335, N4061, N2481);
not NOT1 (N5347, N5325);
xor XOR2 (N5348, N5346, N2125);
and AND2 (N5349, N5348, N4381);
or OR4 (N5350, N5338, N4444, N2623, N4188);
not NOT1 (N5351, N5349);
xor XOR2 (N5352, N5334, N1984);
xor XOR2 (N5353, N5331, N3360);
xor XOR2 (N5354, N5339, N3869);
xor XOR2 (N5355, N5343, N4290);
and AND4 (N5356, N5351, N3981, N4616, N3779);
xor XOR2 (N5357, N5342, N5063);
xor XOR2 (N5358, N5354, N2551);
nor NOR2 (N5359, N5353, N3256);
xor XOR2 (N5360, N5357, N1185);
xor XOR2 (N5361, N5344, N1324);
xor XOR2 (N5362, N5356, N3522);
and AND2 (N5363, N5360, N1462);
nor NOR4 (N5364, N5355, N4053, N2377, N4782);
and AND4 (N5365, N5361, N2628, N3504, N2933);
nor NOR2 (N5366, N5352, N4627);
not NOT1 (N5367, N5365);
or OR3 (N5368, N5362, N1519, N1430);
xor XOR2 (N5369, N5347, N3257);
buf BUF1 (N5370, N5366);
nor NOR4 (N5371, N5358, N1539, N3321, N1840);
nor NOR2 (N5372, N5364, N296);
nand NAND3 (N5373, N5359, N2093, N2681);
buf BUF1 (N5374, N5371);
not NOT1 (N5375, N5367);
and AND4 (N5376, N5372, N1381, N4436, N263);
buf BUF1 (N5377, N5375);
xor XOR2 (N5378, N5374, N546);
not NOT1 (N5379, N5368);
or OR4 (N5380, N5377, N4512, N2723, N984);
not NOT1 (N5381, N5373);
nor NOR3 (N5382, N5378, N4998, N462);
or OR2 (N5383, N5345, N3558);
and AND3 (N5384, N5363, N716, N235);
and AND3 (N5385, N5381, N4088, N4931);
buf BUF1 (N5386, N5350);
and AND4 (N5387, N5386, N3235, N4509, N3479);
nand NAND2 (N5388, N5382, N3179);
nand NAND4 (N5389, N5385, N4822, N5233, N1630);
not NOT1 (N5390, N5383);
nand NAND2 (N5391, N5376, N4074);
nand NAND3 (N5392, N5391, N5280, N1350);
and AND4 (N5393, N5390, N2178, N804, N1613);
xor XOR2 (N5394, N5379, N3529);
nand NAND4 (N5395, N5380, N1836, N2865, N320);
nand NAND4 (N5396, N5387, N3653, N1803, N1658);
xor XOR2 (N5397, N5395, N47);
buf BUF1 (N5398, N5396);
not NOT1 (N5399, N5393);
nand NAND2 (N5400, N5370, N3679);
nor NOR3 (N5401, N5388, N2062, N1743);
buf BUF1 (N5402, N5400);
nor NOR2 (N5403, N5384, N4581);
or OR4 (N5404, N5394, N795, N2702, N4981);
or OR2 (N5405, N5369, N3083);
xor XOR2 (N5406, N5402, N5288);
buf BUF1 (N5407, N5399);
not NOT1 (N5408, N5398);
buf BUF1 (N5409, N5401);
xor XOR2 (N5410, N5408, N999);
not NOT1 (N5411, N5404);
and AND3 (N5412, N5403, N3495, N4022);
or OR3 (N5413, N5389, N1613, N4704);
not NOT1 (N5414, N5407);
nand NAND3 (N5415, N5397, N3922, N3500);
buf BUF1 (N5416, N5410);
and AND4 (N5417, N5411, N2512, N626, N4386);
not NOT1 (N5418, N5412);
nor NOR4 (N5419, N5418, N659, N3673, N5257);
buf BUF1 (N5420, N5417);
nand NAND4 (N5421, N5392, N4719, N3745, N4057);
xor XOR2 (N5422, N5419, N5239);
buf BUF1 (N5423, N5416);
nor NOR3 (N5424, N5406, N1873, N2093);
xor XOR2 (N5425, N5422, N984);
xor XOR2 (N5426, N5414, N3009);
buf BUF1 (N5427, N5425);
not NOT1 (N5428, N5426);
not NOT1 (N5429, N5423);
not NOT1 (N5430, N5424);
not NOT1 (N5431, N5430);
buf BUF1 (N5432, N5413);
xor XOR2 (N5433, N5429, N954);
buf BUF1 (N5434, N5409);
nor NOR2 (N5435, N5415, N1297);
not NOT1 (N5436, N5428);
buf BUF1 (N5437, N5432);
not NOT1 (N5438, N5434);
xor XOR2 (N5439, N5427, N1237);
buf BUF1 (N5440, N5421);
buf BUF1 (N5441, N5436);
xor XOR2 (N5442, N5441, N3286);
buf BUF1 (N5443, N5420);
and AND4 (N5444, N5439, N4403, N1408, N4046);
not NOT1 (N5445, N5433);
nand NAND3 (N5446, N5443, N5094, N4058);
or OR4 (N5447, N5444, N1968, N181, N3415);
nand NAND2 (N5448, N5431, N1363);
nand NAND3 (N5449, N5445, N4906, N3786);
nor NOR2 (N5450, N5437, N1477);
nor NOR2 (N5451, N5440, N1466);
nand NAND4 (N5452, N5442, N970, N5375, N1727);
nand NAND4 (N5453, N5446, N2578, N2038, N152);
or OR4 (N5454, N5435, N1995, N3030, N4275);
not NOT1 (N5455, N5453);
not NOT1 (N5456, N5447);
and AND4 (N5457, N5449, N698, N870, N3256);
nor NOR3 (N5458, N5452, N2505, N4620);
xor XOR2 (N5459, N5458, N2851);
or OR2 (N5460, N5454, N2336);
not NOT1 (N5461, N5448);
or OR4 (N5462, N5450, N3186, N1508, N25);
nor NOR4 (N5463, N5456, N3059, N2964, N1477);
and AND3 (N5464, N5438, N2883, N4841);
nor NOR3 (N5465, N5463, N4027, N1227);
not NOT1 (N5466, N5461);
or OR4 (N5467, N5451, N1935, N1437, N378);
nor NOR2 (N5468, N5459, N3526);
not NOT1 (N5469, N5466);
nor NOR4 (N5470, N5465, N4050, N419, N4187);
and AND4 (N5471, N5460, N1889, N4724, N2468);
nor NOR4 (N5472, N5467, N4007, N2548, N5340);
nand NAND3 (N5473, N5472, N1886, N3112);
not NOT1 (N5474, N5469);
nor NOR2 (N5475, N5468, N852);
or OR4 (N5476, N5474, N2140, N4001, N873);
and AND4 (N5477, N5473, N2386, N2127, N2414);
nand NAND4 (N5478, N5471, N1101, N4548, N1009);
and AND3 (N5479, N5405, N145, N4209);
or OR4 (N5480, N5479, N4284, N1926, N1049);
buf BUF1 (N5481, N5470);
not NOT1 (N5482, N5462);
or OR2 (N5483, N5478, N4393);
not NOT1 (N5484, N5455);
xor XOR2 (N5485, N5475, N1282);
nor NOR4 (N5486, N5482, N1185, N167, N4362);
or OR4 (N5487, N5480, N2009, N490, N5410);
or OR4 (N5488, N5484, N5156, N171, N2885);
buf BUF1 (N5489, N5476);
not NOT1 (N5490, N5464);
or OR4 (N5491, N5483, N982, N2291, N3244);
nor NOR3 (N5492, N5457, N2854, N480);
not NOT1 (N5493, N5489);
not NOT1 (N5494, N5490);
buf BUF1 (N5495, N5492);
or OR3 (N5496, N5495, N3147, N1196);
or OR2 (N5497, N5493, N2822);
buf BUF1 (N5498, N5488);
nand NAND2 (N5499, N5486, N1718);
xor XOR2 (N5500, N5487, N4232);
nand NAND3 (N5501, N5494, N796, N2923);
xor XOR2 (N5502, N5497, N4003);
not NOT1 (N5503, N5491);
and AND3 (N5504, N5485, N4279, N3510);
or OR4 (N5505, N5503, N503, N3501, N1166);
not NOT1 (N5506, N5477);
not NOT1 (N5507, N5500);
nand NAND4 (N5508, N5504, N4715, N3678, N4407);
or OR4 (N5509, N5496, N3116, N4237, N1418);
nand NAND3 (N5510, N5499, N5058, N3102);
buf BUF1 (N5511, N5506);
and AND4 (N5512, N5507, N2766, N1499, N1348);
not NOT1 (N5513, N5501);
not NOT1 (N5514, N5481);
or OR4 (N5515, N5514, N712, N1365, N4180);
nor NOR2 (N5516, N5502, N1060);
nor NOR2 (N5517, N5515, N811);
and AND3 (N5518, N5513, N1780, N1803);
and AND4 (N5519, N5509, N2402, N3983, N5007);
and AND2 (N5520, N5510, N4072);
or OR3 (N5521, N5517, N1127, N2194);
nand NAND2 (N5522, N5520, N2282);
nand NAND3 (N5523, N5522, N4705, N1111);
nand NAND2 (N5524, N5523, N2940);
not NOT1 (N5525, N5511);
nand NAND2 (N5526, N5524, N2627);
xor XOR2 (N5527, N5521, N736);
nand NAND4 (N5528, N5498, N917, N2453, N2344);
xor XOR2 (N5529, N5508, N4553);
buf BUF1 (N5530, N5516);
and AND2 (N5531, N5527, N1998);
not NOT1 (N5532, N5518);
and AND2 (N5533, N5525, N1012);
xor XOR2 (N5534, N5519, N872);
buf BUF1 (N5535, N5532);
not NOT1 (N5536, N5512);
not NOT1 (N5537, N5534);
not NOT1 (N5538, N5537);
nor NOR2 (N5539, N5526, N3064);
nor NOR4 (N5540, N5539, N439, N74, N964);
nand NAND4 (N5541, N5540, N2187, N3106, N4797);
and AND3 (N5542, N5505, N1388, N1883);
nor NOR3 (N5543, N5533, N1131, N5356);
nor NOR4 (N5544, N5528, N2618, N1971, N1951);
buf BUF1 (N5545, N5536);
and AND4 (N5546, N5538, N4138, N3119, N2336);
and AND3 (N5547, N5545, N3103, N268);
nor NOR3 (N5548, N5542, N1332, N190);
not NOT1 (N5549, N5546);
nand NAND3 (N5550, N5529, N303, N3044);
nor NOR3 (N5551, N5530, N2750, N60);
buf BUF1 (N5552, N5550);
nand NAND3 (N5553, N5543, N3533, N3680);
xor XOR2 (N5554, N5549, N1312);
nor NOR4 (N5555, N5541, N3647, N4627, N5342);
buf BUF1 (N5556, N5553);
xor XOR2 (N5557, N5552, N3115);
buf BUF1 (N5558, N5555);
or OR2 (N5559, N5558, N744);
buf BUF1 (N5560, N5531);
and AND4 (N5561, N5548, N1920, N1039, N4167);
not NOT1 (N5562, N5551);
and AND3 (N5563, N5535, N726, N3949);
not NOT1 (N5564, N5562);
nor NOR3 (N5565, N5544, N2546, N3914);
nand NAND3 (N5566, N5554, N5018, N467);
nor NOR4 (N5567, N5561, N932, N552, N5133);
or OR4 (N5568, N5564, N2682, N199, N2351);
and AND3 (N5569, N5547, N5246, N273);
buf BUF1 (N5570, N5567);
nand NAND3 (N5571, N5568, N754, N772);
nand NAND3 (N5572, N5556, N4002, N5058);
not NOT1 (N5573, N5566);
not NOT1 (N5574, N5570);
buf BUF1 (N5575, N5571);
or OR2 (N5576, N5572, N1379);
buf BUF1 (N5577, N5559);
xor XOR2 (N5578, N5560, N942);
nor NOR4 (N5579, N5565, N2645, N4658, N60);
nand NAND2 (N5580, N5576, N3177);
nand NAND2 (N5581, N5577, N66);
nand NAND2 (N5582, N5578, N4576);
nor NOR4 (N5583, N5557, N1719, N3263, N1916);
and AND2 (N5584, N5573, N4030);
buf BUF1 (N5585, N5583);
buf BUF1 (N5586, N5582);
and AND3 (N5587, N5569, N2232, N67);
and AND2 (N5588, N5587, N3485);
and AND2 (N5589, N5584, N2539);
buf BUF1 (N5590, N5586);
not NOT1 (N5591, N5581);
nand NAND4 (N5592, N5591, N2501, N4732, N4933);
nand NAND4 (N5593, N5592, N4968, N4060, N5003);
nor NOR4 (N5594, N5588, N1051, N1014, N4363);
xor XOR2 (N5595, N5593, N4429);
nand NAND3 (N5596, N5595, N1850, N3427);
nor NOR3 (N5597, N5585, N171, N70);
nand NAND4 (N5598, N5574, N1198, N5053, N5135);
not NOT1 (N5599, N5589);
nor NOR2 (N5600, N5596, N201);
nor NOR3 (N5601, N5563, N5353, N3667);
not NOT1 (N5602, N5597);
and AND3 (N5603, N5601, N1662, N2792);
nor NOR2 (N5604, N5579, N4231);
nor NOR4 (N5605, N5604, N2065, N127, N4653);
nand NAND4 (N5606, N5599, N2312, N3369, N681);
xor XOR2 (N5607, N5598, N279);
nand NAND3 (N5608, N5603, N5021, N4183);
xor XOR2 (N5609, N5607, N3640);
and AND2 (N5610, N5600, N1374);
xor XOR2 (N5611, N5580, N1048);
buf BUF1 (N5612, N5606);
buf BUF1 (N5613, N5612);
nor NOR2 (N5614, N5613, N3128);
nand NAND3 (N5615, N5590, N5474, N2070);
nand NAND2 (N5616, N5610, N5250);
or OR4 (N5617, N5575, N1078, N3157, N3658);
nor NOR4 (N5618, N5617, N4907, N4352, N4579);
xor XOR2 (N5619, N5616, N1368);
nor NOR3 (N5620, N5615, N325, N4044);
not NOT1 (N5621, N5614);
nand NAND4 (N5622, N5608, N1634, N1057, N4663);
or OR2 (N5623, N5594, N4551);
not NOT1 (N5624, N5621);
and AND2 (N5625, N5605, N3562);
not NOT1 (N5626, N5624);
not NOT1 (N5627, N5611);
and AND3 (N5628, N5602, N3851, N5158);
nor NOR4 (N5629, N5609, N3821, N2940, N1493);
nor NOR3 (N5630, N5628, N927, N2106);
not NOT1 (N5631, N5620);
not NOT1 (N5632, N5623);
nand NAND3 (N5633, N5622, N4704, N1584);
or OR4 (N5634, N5631, N5103, N1134, N4754);
not NOT1 (N5635, N5627);
and AND4 (N5636, N5634, N1829, N2558, N1935);
nor NOR3 (N5637, N5635, N458, N4230);
buf BUF1 (N5638, N5637);
xor XOR2 (N5639, N5618, N1629);
or OR2 (N5640, N5632, N3931);
xor XOR2 (N5641, N5619, N4701);
or OR4 (N5642, N5641, N2414, N5285, N296);
nand NAND2 (N5643, N5629, N2246);
nor NOR4 (N5644, N5636, N1246, N1574, N585);
xor XOR2 (N5645, N5640, N3541);
nand NAND4 (N5646, N5638, N4117, N4779, N4219);
or OR2 (N5647, N5639, N3850);
nor NOR4 (N5648, N5644, N1350, N2536, N4396);
or OR2 (N5649, N5646, N3854);
not NOT1 (N5650, N5642);
or OR4 (N5651, N5645, N1292, N817, N4682);
xor XOR2 (N5652, N5649, N4623);
or OR3 (N5653, N5651, N4404, N3575);
buf BUF1 (N5654, N5647);
not NOT1 (N5655, N5625);
nor NOR3 (N5656, N5650, N910, N324);
and AND2 (N5657, N5643, N3156);
or OR2 (N5658, N5657, N5373);
and AND3 (N5659, N5656, N4577, N1169);
and AND3 (N5660, N5655, N1954, N1636);
nand NAND4 (N5661, N5633, N4738, N880, N5364);
buf BUF1 (N5662, N5658);
or OR2 (N5663, N5660, N3986);
not NOT1 (N5664, N5626);
xor XOR2 (N5665, N5653, N4046);
xor XOR2 (N5666, N5665, N4648);
or OR3 (N5667, N5654, N3310, N2181);
nor NOR2 (N5668, N5659, N4695);
or OR3 (N5669, N5663, N3476, N778);
nor NOR2 (N5670, N5664, N1139);
buf BUF1 (N5671, N5662);
or OR3 (N5672, N5669, N869, N1032);
and AND4 (N5673, N5630, N4270, N2641, N3970);
xor XOR2 (N5674, N5672, N3647);
nand NAND2 (N5675, N5670, N2403);
buf BUF1 (N5676, N5675);
nor NOR3 (N5677, N5666, N281, N5015);
buf BUF1 (N5678, N5667);
not NOT1 (N5679, N5674);
or OR3 (N5680, N5678, N850, N2615);
or OR4 (N5681, N5661, N1800, N1789, N1799);
or OR4 (N5682, N5676, N729, N3778, N4391);
and AND2 (N5683, N5679, N2540);
xor XOR2 (N5684, N5648, N4255);
xor XOR2 (N5685, N5673, N2624);
or OR3 (N5686, N5684, N3772, N5621);
or OR3 (N5687, N5680, N399, N1221);
or OR2 (N5688, N5685, N4712);
nor NOR4 (N5689, N5671, N2298, N5263, N1404);
not NOT1 (N5690, N5688);
and AND4 (N5691, N5681, N2100, N997, N4161);
or OR2 (N5692, N5686, N4599);
buf BUF1 (N5693, N5652);
and AND4 (N5694, N5687, N1023, N1185, N5294);
xor XOR2 (N5695, N5690, N3235);
and AND3 (N5696, N5682, N5268, N3492);
nand NAND3 (N5697, N5689, N2511, N5119);
buf BUF1 (N5698, N5696);
nand NAND2 (N5699, N5693, N1929);
xor XOR2 (N5700, N5697, N3281);
not NOT1 (N5701, N5698);
not NOT1 (N5702, N5683);
not NOT1 (N5703, N5694);
and AND3 (N5704, N5702, N1881, N5068);
nor NOR3 (N5705, N5695, N5173, N3432);
not NOT1 (N5706, N5704);
buf BUF1 (N5707, N5703);
and AND4 (N5708, N5692, N3894, N18, N3596);
buf BUF1 (N5709, N5691);
xor XOR2 (N5710, N5707, N4272);
nand NAND4 (N5711, N5705, N4003, N1754, N3982);
nand NAND2 (N5712, N5710, N1013);
buf BUF1 (N5713, N5708);
nand NAND3 (N5714, N5706, N3916, N5704);
nor NOR2 (N5715, N5709, N59);
nand NAND2 (N5716, N5700, N186);
nand NAND4 (N5717, N5712, N1853, N608, N1956);
and AND4 (N5718, N5711, N3914, N2674, N4490);
nor NOR4 (N5719, N5701, N2199, N1137, N1567);
or OR2 (N5720, N5699, N3422);
not NOT1 (N5721, N5668);
buf BUF1 (N5722, N5718);
buf BUF1 (N5723, N5720);
and AND4 (N5724, N5722, N4789, N882, N1014);
nor NOR3 (N5725, N5677, N2611, N472);
and AND4 (N5726, N5719, N4771, N4857, N4155);
nor NOR3 (N5727, N5715, N403, N4078);
nor NOR3 (N5728, N5721, N1138, N1363);
nor NOR4 (N5729, N5725, N2395, N3269, N3750);
and AND4 (N5730, N5716, N2373, N3462, N4510);
or OR4 (N5731, N5717, N1123, N3937, N4551);
or OR3 (N5732, N5731, N2760, N2630);
nor NOR2 (N5733, N5727, N4300);
not NOT1 (N5734, N5733);
and AND4 (N5735, N5714, N1357, N333, N162);
nor NOR2 (N5736, N5735, N561);
xor XOR2 (N5737, N5736, N1489);
nor NOR2 (N5738, N5732, N2343);
and AND4 (N5739, N5723, N1686, N5634, N1323);
nand NAND2 (N5740, N5738, N2073);
or OR3 (N5741, N5713, N3178, N1644);
xor XOR2 (N5742, N5724, N1038);
nor NOR2 (N5743, N5729, N1808);
xor XOR2 (N5744, N5737, N1316);
or OR2 (N5745, N5739, N876);
buf BUF1 (N5746, N5743);
or OR3 (N5747, N5728, N5186, N1351);
or OR3 (N5748, N5746, N668, N3871);
nand NAND3 (N5749, N5744, N5496, N2001);
nand NAND4 (N5750, N5726, N494, N114, N3781);
and AND2 (N5751, N5747, N3997);
nand NAND2 (N5752, N5740, N1368);
not NOT1 (N5753, N5734);
nor NOR4 (N5754, N5748, N3831, N3719, N1698);
buf BUF1 (N5755, N5750);
not NOT1 (N5756, N5749);
buf BUF1 (N5757, N5745);
not NOT1 (N5758, N5741);
nand NAND2 (N5759, N5754, N5013);
not NOT1 (N5760, N5759);
nand NAND2 (N5761, N5730, N3641);
not NOT1 (N5762, N5742);
and AND4 (N5763, N5753, N5606, N3818, N598);
nand NAND3 (N5764, N5758, N1837, N3842);
nor NOR4 (N5765, N5760, N2829, N758, N5600);
buf BUF1 (N5766, N5761);
or OR4 (N5767, N5762, N319, N2048, N1159);
xor XOR2 (N5768, N5763, N131);
nand NAND4 (N5769, N5751, N2444, N3303, N5670);
nor NOR3 (N5770, N5752, N2907, N4871);
buf BUF1 (N5771, N5764);
and AND2 (N5772, N5757, N3781);
nor NOR4 (N5773, N5772, N3457, N2519, N3938);
xor XOR2 (N5774, N5768, N1731);
not NOT1 (N5775, N5774);
nor NOR4 (N5776, N5775, N1692, N5314, N3251);
not NOT1 (N5777, N5755);
xor XOR2 (N5778, N5769, N1235);
nor NOR3 (N5779, N5756, N4708, N5233);
xor XOR2 (N5780, N5777, N4168);
nand NAND4 (N5781, N5778, N2988, N1690, N4314);
xor XOR2 (N5782, N5779, N831);
or OR2 (N5783, N5766, N2654);
xor XOR2 (N5784, N5770, N5417);
nand NAND3 (N5785, N5783, N5164, N5424);
xor XOR2 (N5786, N5782, N5729);
nor NOR3 (N5787, N5786, N4882, N2187);
buf BUF1 (N5788, N5787);
nor NOR2 (N5789, N5781, N5172);
buf BUF1 (N5790, N5780);
not NOT1 (N5791, N5784);
nand NAND3 (N5792, N5771, N3726, N143);
buf BUF1 (N5793, N5776);
and AND4 (N5794, N5789, N1593, N1341, N2759);
and AND3 (N5795, N5765, N1338, N478);
xor XOR2 (N5796, N5791, N2181);
not NOT1 (N5797, N5795);
nor NOR3 (N5798, N5767, N1234, N4382);
or OR4 (N5799, N5796, N827, N2377, N4657);
or OR4 (N5800, N5797, N4035, N4869, N2594);
nand NAND3 (N5801, N5788, N4704, N118);
nand NAND2 (N5802, N5790, N2244);
not NOT1 (N5803, N5773);
not NOT1 (N5804, N5802);
nand NAND3 (N5805, N5798, N3343, N166);
not NOT1 (N5806, N5801);
nand NAND4 (N5807, N5805, N5131, N3555, N5155);
or OR4 (N5808, N5794, N2061, N4426, N1050);
nor NOR2 (N5809, N5806, N4263);
or OR3 (N5810, N5792, N469, N3424);
nand NAND3 (N5811, N5785, N1150, N3321);
xor XOR2 (N5812, N5808, N951);
nor NOR4 (N5813, N5812, N5116, N500, N1890);
and AND2 (N5814, N5809, N5706);
xor XOR2 (N5815, N5804, N381);
or OR3 (N5816, N5810, N1980, N3774);
buf BUF1 (N5817, N5816);
or OR4 (N5818, N5813, N3308, N3672, N5221);
nor NOR4 (N5819, N5815, N1130, N4570, N4856);
nor NOR4 (N5820, N5811, N3656, N5580, N4115);
nand NAND4 (N5821, N5807, N4423, N3917, N3179);
nor NOR2 (N5822, N5793, N4279);
and AND4 (N5823, N5821, N1980, N5172, N5519);
not NOT1 (N5824, N5823);
not NOT1 (N5825, N5799);
buf BUF1 (N5826, N5822);
or OR2 (N5827, N5817, N3804);
xor XOR2 (N5828, N5820, N848);
xor XOR2 (N5829, N5819, N661);
nand NAND2 (N5830, N5818, N4501);
xor XOR2 (N5831, N5830, N4708);
xor XOR2 (N5832, N5814, N5590);
not NOT1 (N5833, N5829);
xor XOR2 (N5834, N5824, N1299);
xor XOR2 (N5835, N5827, N3931);
or OR4 (N5836, N5826, N280, N3791, N896);
not NOT1 (N5837, N5832);
nor NOR4 (N5838, N5831, N2559, N3978, N3881);
and AND2 (N5839, N5837, N81);
and AND3 (N5840, N5833, N3956, N5674);
buf BUF1 (N5841, N5803);
xor XOR2 (N5842, N5828, N578);
and AND4 (N5843, N5838, N4732, N4521, N933);
xor XOR2 (N5844, N5840, N5417);
and AND4 (N5845, N5800, N1393, N4670, N4860);
or OR3 (N5846, N5835, N3003, N2561);
xor XOR2 (N5847, N5839, N1685);
and AND2 (N5848, N5825, N259);
not NOT1 (N5849, N5847);
not NOT1 (N5850, N5836);
nor NOR4 (N5851, N5850, N3657, N1586, N754);
not NOT1 (N5852, N5841);
and AND3 (N5853, N5852, N5514, N60);
nand NAND4 (N5854, N5849, N1555, N5238, N4218);
and AND2 (N5855, N5851, N521);
and AND2 (N5856, N5853, N5385);
nand NAND2 (N5857, N5842, N1121);
xor XOR2 (N5858, N5844, N4454);
and AND2 (N5859, N5845, N5764);
buf BUF1 (N5860, N5857);
buf BUF1 (N5861, N5846);
or OR3 (N5862, N5860, N2038, N4274);
buf BUF1 (N5863, N5843);
nand NAND4 (N5864, N5834, N1425, N4507, N5215);
and AND4 (N5865, N5848, N2789, N3832, N1109);
or OR2 (N5866, N5859, N3525);
nand NAND4 (N5867, N5856, N536, N3552, N3582);
not NOT1 (N5868, N5867);
nor NOR3 (N5869, N5862, N5029, N2781);
nand NAND4 (N5870, N5865, N3122, N4892, N3197);
and AND2 (N5871, N5863, N2535);
nand NAND4 (N5872, N5858, N104, N3940, N3664);
and AND2 (N5873, N5861, N3760);
and AND3 (N5874, N5870, N4988, N1425);
xor XOR2 (N5875, N5871, N5364);
and AND2 (N5876, N5864, N4256);
not NOT1 (N5877, N5874);
buf BUF1 (N5878, N5855);
or OR2 (N5879, N5872, N1624);
buf BUF1 (N5880, N5875);
not NOT1 (N5881, N5877);
and AND4 (N5882, N5878, N5818, N4423, N395);
nand NAND4 (N5883, N5868, N2973, N984, N3043);
xor XOR2 (N5884, N5854, N1121);
nor NOR3 (N5885, N5873, N886, N4462);
and AND4 (N5886, N5876, N2619, N4198, N4874);
buf BUF1 (N5887, N5880);
or OR3 (N5888, N5866, N868, N2243);
nor NOR3 (N5889, N5888, N2770, N2975);
not NOT1 (N5890, N5887);
not NOT1 (N5891, N5886);
or OR4 (N5892, N5884, N1045, N607, N2997);
xor XOR2 (N5893, N5882, N1398);
and AND2 (N5894, N5879, N4711);
or OR3 (N5895, N5891, N3013, N4937);
buf BUF1 (N5896, N5890);
xor XOR2 (N5897, N5894, N462);
xor XOR2 (N5898, N5893, N1710);
or OR4 (N5899, N5883, N3995, N2185, N4802);
or OR2 (N5900, N5889, N5823);
nor NOR2 (N5901, N5895, N3001);
xor XOR2 (N5902, N5885, N3226);
xor XOR2 (N5903, N5902, N3750);
nor NOR4 (N5904, N5892, N4990, N3686, N3289);
buf BUF1 (N5905, N5898);
or OR2 (N5906, N5903, N2696);
nand NAND2 (N5907, N5881, N5031);
or OR2 (N5908, N5904, N76);
not NOT1 (N5909, N5901);
nor NOR4 (N5910, N5869, N1360, N3264, N5439);
nor NOR3 (N5911, N5909, N4274, N2370);
not NOT1 (N5912, N5896);
or OR3 (N5913, N5906, N886, N4648);
nor NOR2 (N5914, N5911, N2376);
nand NAND2 (N5915, N5912, N1432);
xor XOR2 (N5916, N5910, N4740);
not NOT1 (N5917, N5913);
buf BUF1 (N5918, N5914);
nand NAND4 (N5919, N5918, N4830, N116, N939);
and AND4 (N5920, N5916, N1484, N5067, N3653);
nor NOR4 (N5921, N5905, N4859, N4166, N2350);
nor NOR2 (N5922, N5920, N2331);
nand NAND2 (N5923, N5907, N5386);
and AND3 (N5924, N5908, N3356, N336);
or OR2 (N5925, N5922, N5621);
not NOT1 (N5926, N5921);
and AND4 (N5927, N5926, N1271, N5754, N822);
and AND2 (N5928, N5899, N2266);
or OR2 (N5929, N5917, N3905);
xor XOR2 (N5930, N5928, N1148);
nor NOR3 (N5931, N5930, N902, N2157);
nor NOR2 (N5932, N5897, N2289);
buf BUF1 (N5933, N5923);
nand NAND4 (N5934, N5929, N980, N4938, N2668);
and AND2 (N5935, N5915, N3581);
xor XOR2 (N5936, N5919, N5263);
or OR3 (N5937, N5925, N1991, N4660);
not NOT1 (N5938, N5927);
and AND3 (N5939, N5933, N2646, N1927);
not NOT1 (N5940, N5939);
or OR4 (N5941, N5900, N159, N552, N5039);
nand NAND2 (N5942, N5940, N5136);
or OR4 (N5943, N5931, N2117, N4660, N5789);
nand NAND2 (N5944, N5938, N4220);
not NOT1 (N5945, N5934);
nand NAND4 (N5946, N5942, N5894, N5139, N3700);
and AND2 (N5947, N5943, N5145);
nor NOR3 (N5948, N5941, N1821, N1416);
buf BUF1 (N5949, N5945);
nand NAND3 (N5950, N5947, N5694, N1870);
nand NAND2 (N5951, N5932, N801);
nand NAND2 (N5952, N5951, N2166);
buf BUF1 (N5953, N5949);
and AND3 (N5954, N5936, N1306, N2614);
nor NOR4 (N5955, N5937, N5171, N4265, N2630);
nand NAND4 (N5956, N5935, N2115, N2237, N890);
buf BUF1 (N5957, N5948);
nand NAND2 (N5958, N5954, N4164);
or OR2 (N5959, N5950, N165);
buf BUF1 (N5960, N5953);
nor NOR2 (N5961, N5924, N2444);
not NOT1 (N5962, N5952);
not NOT1 (N5963, N5960);
nand NAND3 (N5964, N5955, N4964, N2966);
nor NOR2 (N5965, N5957, N1765);
xor XOR2 (N5966, N5965, N3235);
buf BUF1 (N5967, N5958);
or OR2 (N5968, N5962, N1650);
nand NAND2 (N5969, N5946, N5577);
and AND3 (N5970, N5959, N2524, N1211);
nor NOR4 (N5971, N5970, N3872, N4311, N3632);
and AND4 (N5972, N5956, N632, N3088, N3736);
or OR2 (N5973, N5972, N913);
and AND3 (N5974, N5964, N468, N4986);
nor NOR4 (N5975, N5968, N5817, N3112, N5694);
or OR2 (N5976, N5963, N3066);
and AND2 (N5977, N5971, N397);
nand NAND4 (N5978, N5974, N1127, N2691, N3171);
xor XOR2 (N5979, N5977, N2801);
xor XOR2 (N5980, N5967, N5237);
and AND4 (N5981, N5978, N5521, N5268, N5484);
nor NOR3 (N5982, N5969, N1822, N69);
xor XOR2 (N5983, N5966, N77);
nor NOR4 (N5984, N5981, N4743, N1752, N4743);
or OR3 (N5985, N5980, N820, N5195);
and AND3 (N5986, N5979, N5030, N5472);
xor XOR2 (N5987, N5986, N5815);
and AND2 (N5988, N5976, N3332);
xor XOR2 (N5989, N5988, N3105);
and AND2 (N5990, N5984, N4618);
buf BUF1 (N5991, N5982);
and AND3 (N5992, N5961, N3488, N970);
nand NAND2 (N5993, N5973, N2441);
not NOT1 (N5994, N5989);
or OR2 (N5995, N5990, N3021);
buf BUF1 (N5996, N5944);
not NOT1 (N5997, N5992);
nor NOR2 (N5998, N5991, N5766);
not NOT1 (N5999, N5994);
not NOT1 (N6000, N5985);
not NOT1 (N6001, N6000);
xor XOR2 (N6002, N5997, N4370);
not NOT1 (N6003, N6002);
buf BUF1 (N6004, N6001);
or OR3 (N6005, N5999, N3229, N5240);
nand NAND3 (N6006, N5998, N4284, N5305);
and AND3 (N6007, N6005, N802, N5746);
nor NOR4 (N6008, N6004, N5372, N1373, N5102);
or OR3 (N6009, N6003, N2815, N2390);
and AND4 (N6010, N5983, N3857, N4733, N4814);
nand NAND3 (N6011, N6008, N2456, N3666);
nor NOR2 (N6012, N5987, N3105);
xor XOR2 (N6013, N5996, N882);
not NOT1 (N6014, N6007);
nor NOR3 (N6015, N6011, N2411, N210);
and AND3 (N6016, N6006, N4033, N5131);
and AND4 (N6017, N6010, N5406, N5475, N568);
not NOT1 (N6018, N5975);
nor NOR2 (N6019, N6009, N1812);
xor XOR2 (N6020, N6013, N2707);
xor XOR2 (N6021, N6017, N5262);
or OR3 (N6022, N5993, N2329, N1308);
buf BUF1 (N6023, N6019);
and AND3 (N6024, N6014, N5128, N3144);
buf BUF1 (N6025, N5995);
xor XOR2 (N6026, N6023, N2485);
xor XOR2 (N6027, N6025, N1306);
xor XOR2 (N6028, N6012, N4426);
xor XOR2 (N6029, N6022, N5311);
xor XOR2 (N6030, N6016, N4133);
or OR4 (N6031, N6026, N3688, N2780, N3181);
nand NAND2 (N6032, N6030, N6021);
xor XOR2 (N6033, N3748, N1177);
nand NAND4 (N6034, N6032, N88, N1230, N1525);
and AND4 (N6035, N6024, N4521, N638, N2095);
buf BUF1 (N6036, N6033);
and AND2 (N6037, N6020, N4348);
buf BUF1 (N6038, N6028);
or OR2 (N6039, N6027, N2434);
buf BUF1 (N6040, N6038);
buf BUF1 (N6041, N6040);
not NOT1 (N6042, N6034);
not NOT1 (N6043, N6041);
or OR4 (N6044, N6039, N4879, N2344, N1780);
buf BUF1 (N6045, N6018);
or OR4 (N6046, N6036, N4977, N2815, N3238);
not NOT1 (N6047, N6037);
xor XOR2 (N6048, N6045, N4035);
nand NAND3 (N6049, N6048, N2003, N6005);
not NOT1 (N6050, N6031);
not NOT1 (N6051, N6050);
not NOT1 (N6052, N6043);
xor XOR2 (N6053, N6052, N3810);
buf BUF1 (N6054, N6046);
not NOT1 (N6055, N6044);
xor XOR2 (N6056, N6053, N3153);
buf BUF1 (N6057, N6056);
nor NOR3 (N6058, N6054, N1448, N3922);
nand NAND2 (N6059, N6055, N3650);
not NOT1 (N6060, N6059);
not NOT1 (N6061, N6057);
nand NAND2 (N6062, N6058, N4856);
nor NOR2 (N6063, N6061, N1258);
xor XOR2 (N6064, N6062, N4726);
not NOT1 (N6065, N6051);
nor NOR3 (N6066, N6065, N2510, N2779);
not NOT1 (N6067, N6029);
not NOT1 (N6068, N6035);
nand NAND2 (N6069, N6042, N2215);
nor NOR3 (N6070, N6015, N5304, N1797);
buf BUF1 (N6071, N6068);
buf BUF1 (N6072, N6070);
nor NOR2 (N6073, N6064, N2811);
buf BUF1 (N6074, N6072);
not NOT1 (N6075, N6049);
nor NOR3 (N6076, N6073, N4281, N112);
buf BUF1 (N6077, N6066);
and AND4 (N6078, N6075, N2014, N2206, N1604);
xor XOR2 (N6079, N6071, N511);
buf BUF1 (N6080, N6074);
and AND3 (N6081, N6079, N1088, N3613);
nor NOR4 (N6082, N6078, N4931, N4966, N491);
and AND4 (N6083, N6060, N872, N4295, N1284);
nor NOR4 (N6084, N6083, N4539, N2616, N1006);
buf BUF1 (N6085, N6082);
buf BUF1 (N6086, N6077);
nand NAND4 (N6087, N6085, N3939, N2653, N3678);
or OR2 (N6088, N6063, N4479);
and AND4 (N6089, N6047, N1892, N5795, N1792);
xor XOR2 (N6090, N6084, N2427);
not NOT1 (N6091, N6087);
not NOT1 (N6092, N6080);
and AND3 (N6093, N6091, N5521, N2390);
nand NAND3 (N6094, N6076, N4636, N5159);
buf BUF1 (N6095, N6081);
xor XOR2 (N6096, N6093, N3869);
nand NAND3 (N6097, N6090, N4537, N5622);
xor XOR2 (N6098, N6089, N1057);
nand NAND2 (N6099, N6092, N4079);
not NOT1 (N6100, N6097);
nand NAND4 (N6101, N6098, N4399, N5318, N4654);
buf BUF1 (N6102, N6094);
and AND2 (N6103, N6099, N2667);
nand NAND3 (N6104, N6103, N4957, N4893);
buf BUF1 (N6105, N6069);
and AND4 (N6106, N6105, N3082, N256, N675);
nand NAND4 (N6107, N6101, N3288, N2748, N3579);
or OR3 (N6108, N6107, N4958, N884);
or OR4 (N6109, N6086, N5944, N1004, N1900);
and AND4 (N6110, N6096, N2635, N2566, N2695);
xor XOR2 (N6111, N6109, N5488);
nand NAND3 (N6112, N6088, N3045, N4458);
or OR2 (N6113, N6106, N4554);
nor NOR3 (N6114, N6110, N721, N4585);
xor XOR2 (N6115, N6111, N3712);
xor XOR2 (N6116, N6100, N1159);
buf BUF1 (N6117, N6108);
buf BUF1 (N6118, N6112);
not NOT1 (N6119, N6114);
buf BUF1 (N6120, N6102);
nand NAND3 (N6121, N6118, N454, N200);
xor XOR2 (N6122, N6067, N1108);
nand NAND2 (N6123, N6117, N4294);
and AND2 (N6124, N6115, N1823);
nor NOR4 (N6125, N6124, N4045, N3956, N2429);
xor XOR2 (N6126, N6121, N4487);
and AND2 (N6127, N6104, N2247);
or OR4 (N6128, N6123, N173, N749, N5725);
buf BUF1 (N6129, N6126);
or OR3 (N6130, N6125, N5066, N393);
nor NOR3 (N6131, N6129, N2495, N5655);
or OR3 (N6132, N6127, N3473, N5094);
nand NAND2 (N6133, N6132, N4378);
nor NOR3 (N6134, N6119, N436, N2086);
and AND4 (N6135, N6130, N3165, N5255, N5284);
buf BUF1 (N6136, N6133);
not NOT1 (N6137, N6120);
and AND2 (N6138, N6136, N4339);
nor NOR3 (N6139, N6135, N6092, N4979);
xor XOR2 (N6140, N6131, N3410);
xor XOR2 (N6141, N6138, N3842);
xor XOR2 (N6142, N6128, N4768);
nand NAND3 (N6143, N6139, N5332, N5688);
and AND2 (N6144, N6142, N1837);
not NOT1 (N6145, N6113);
not NOT1 (N6146, N6143);
buf BUF1 (N6147, N6140);
nand NAND3 (N6148, N6095, N544, N1038);
and AND4 (N6149, N6144, N3707, N3563, N1588);
nor NOR4 (N6150, N6145, N3864, N357, N2606);
nor NOR3 (N6151, N6122, N1889, N2424);
buf BUF1 (N6152, N6147);
xor XOR2 (N6153, N6116, N5897);
nand NAND3 (N6154, N6146, N138, N1151);
or OR4 (N6155, N6141, N5905, N6041, N5604);
nor NOR4 (N6156, N6154, N301, N5948, N3206);
nor NOR4 (N6157, N6153, N1984, N4945, N1138);
not NOT1 (N6158, N6148);
nand NAND2 (N6159, N6149, N867);
buf BUF1 (N6160, N6151);
buf BUF1 (N6161, N6134);
and AND2 (N6162, N6155, N5810);
nor NOR2 (N6163, N6152, N1747);
or OR3 (N6164, N6157, N5109, N4434);
or OR4 (N6165, N6159, N5651, N1856, N3280);
nand NAND3 (N6166, N6164, N5134, N2087);
nor NOR3 (N6167, N6137, N1053, N4176);
nand NAND2 (N6168, N6162, N5945);
not NOT1 (N6169, N6158);
nor NOR4 (N6170, N6150, N4277, N1309, N700);
xor XOR2 (N6171, N6169, N826);
xor XOR2 (N6172, N6161, N3859);
and AND2 (N6173, N6170, N3376);
not NOT1 (N6174, N6160);
xor XOR2 (N6175, N6156, N3910);
xor XOR2 (N6176, N6166, N5839);
and AND3 (N6177, N6176, N5629, N5779);
or OR3 (N6178, N6174, N4490, N4311);
not NOT1 (N6179, N6177);
xor XOR2 (N6180, N6175, N934);
and AND4 (N6181, N6171, N1800, N1831, N3962);
xor XOR2 (N6182, N6179, N1995);
or OR2 (N6183, N6178, N2525);
buf BUF1 (N6184, N6180);
buf BUF1 (N6185, N6172);
nand NAND2 (N6186, N6183, N2016);
not NOT1 (N6187, N6165);
nor NOR2 (N6188, N6167, N2336);
and AND2 (N6189, N6187, N862);
nor NOR3 (N6190, N6186, N70, N509);
and AND2 (N6191, N6182, N515);
not NOT1 (N6192, N6188);
or OR2 (N6193, N6184, N5402);
not NOT1 (N6194, N6190);
not NOT1 (N6195, N6191);
nand NAND2 (N6196, N6193, N1330);
not NOT1 (N6197, N6196);
xor XOR2 (N6198, N6197, N4705);
not NOT1 (N6199, N6192);
nor NOR4 (N6200, N6168, N3545, N138, N5135);
nor NOR4 (N6201, N6163, N3426, N5693, N3233);
xor XOR2 (N6202, N6199, N2548);
xor XOR2 (N6203, N6173, N267);
and AND3 (N6204, N6200, N2869, N4524);
xor XOR2 (N6205, N6185, N889);
nand NAND3 (N6206, N6198, N5764, N235);
xor XOR2 (N6207, N6206, N1756);
or OR3 (N6208, N6189, N2462, N2466);
nand NAND4 (N6209, N6203, N2723, N985, N446);
buf BUF1 (N6210, N6194);
and AND3 (N6211, N6201, N1410, N1351);
or OR3 (N6212, N6207, N989, N1933);
nor NOR4 (N6213, N6205, N5958, N3750, N4371);
or OR2 (N6214, N6212, N34);
or OR4 (N6215, N6209, N5536, N1559, N5078);
or OR4 (N6216, N6213, N82, N4458, N6117);
nand NAND4 (N6217, N6210, N250, N216, N2956);
buf BUF1 (N6218, N6208);
buf BUF1 (N6219, N6202);
not NOT1 (N6220, N6215);
nor NOR3 (N6221, N6216, N1165, N1348);
or OR3 (N6222, N6214, N708, N4901);
and AND3 (N6223, N6220, N1967, N912);
and AND4 (N6224, N6195, N6205, N5350, N5430);
buf BUF1 (N6225, N6221);
not NOT1 (N6226, N6222);
buf BUF1 (N6227, N6219);
not NOT1 (N6228, N6218);
and AND4 (N6229, N6204, N4142, N5986, N5538);
not NOT1 (N6230, N6229);
nand NAND3 (N6231, N6228, N1529, N4227);
not NOT1 (N6232, N6231);
nor NOR4 (N6233, N6227, N4225, N165, N4038);
and AND3 (N6234, N6217, N4654, N4355);
nand NAND4 (N6235, N6232, N1116, N2586, N2956);
nand NAND3 (N6236, N6223, N1242, N5002);
nand NAND2 (N6237, N6236, N1572);
or OR2 (N6238, N6230, N1585);
nand NAND2 (N6239, N6181, N4865);
buf BUF1 (N6240, N6233);
nor NOR4 (N6241, N6211, N4309, N1041, N3650);
nand NAND3 (N6242, N6235, N3567, N1847);
and AND4 (N6243, N6237, N966, N4310, N5379);
not NOT1 (N6244, N6239);
xor XOR2 (N6245, N6241, N4710);
not NOT1 (N6246, N6240);
xor XOR2 (N6247, N6224, N1233);
and AND2 (N6248, N6247, N1488);
xor XOR2 (N6249, N6244, N2702);
nand NAND3 (N6250, N6234, N4492, N22);
nor NOR4 (N6251, N6226, N98, N1814, N4077);
or OR2 (N6252, N6249, N3297);
not NOT1 (N6253, N6251);
nor NOR3 (N6254, N6243, N2518, N2632);
nand NAND3 (N6255, N6248, N4415, N6011);
nor NOR3 (N6256, N6254, N4200, N6193);
nand NAND3 (N6257, N6252, N1308, N3512);
not NOT1 (N6258, N6256);
and AND2 (N6259, N6257, N3271);
xor XOR2 (N6260, N6250, N1310);
or OR2 (N6261, N6259, N173);
xor XOR2 (N6262, N6260, N5806);
or OR2 (N6263, N6245, N3656);
nor NOR2 (N6264, N6242, N1946);
or OR2 (N6265, N6225, N3342);
nand NAND2 (N6266, N6261, N286);
or OR4 (N6267, N6263, N3182, N2144, N2064);
nor NOR3 (N6268, N6255, N6185, N679);
xor XOR2 (N6269, N6265, N4477);
buf BUF1 (N6270, N6246);
nor NOR3 (N6271, N6267, N5122, N5391);
nor NOR3 (N6272, N6238, N3984, N2590);
buf BUF1 (N6273, N6262);
nor NOR4 (N6274, N6253, N5457, N4499, N5275);
or OR3 (N6275, N6273, N1106, N3579);
nor NOR4 (N6276, N6275, N490, N5370, N3657);
xor XOR2 (N6277, N6266, N2725);
or OR3 (N6278, N6264, N3215, N1120);
and AND4 (N6279, N6270, N1375, N6141, N3483);
nor NOR2 (N6280, N6274, N5264);
or OR3 (N6281, N6278, N3697, N1398);
or OR3 (N6282, N6271, N5462, N5678);
or OR4 (N6283, N6269, N4283, N5911, N1321);
buf BUF1 (N6284, N6276);
buf BUF1 (N6285, N6282);
or OR3 (N6286, N6284, N5468, N4158);
not NOT1 (N6287, N6283);
buf BUF1 (N6288, N6272);
or OR3 (N6289, N6288, N6167, N1291);
xor XOR2 (N6290, N6289, N5757);
nor NOR4 (N6291, N6268, N827, N5276, N4288);
or OR2 (N6292, N6281, N5155);
nand NAND4 (N6293, N6279, N3570, N5188, N2830);
not NOT1 (N6294, N6258);
nor NOR4 (N6295, N6292, N328, N3515, N4496);
and AND2 (N6296, N6293, N5462);
buf BUF1 (N6297, N6277);
or OR4 (N6298, N6296, N4674, N4571, N3772);
buf BUF1 (N6299, N6290);
nand NAND3 (N6300, N6285, N754, N1856);
xor XOR2 (N6301, N6291, N4853);
xor XOR2 (N6302, N6299, N1994);
nor NOR2 (N6303, N6298, N2317);
buf BUF1 (N6304, N6302);
nor NOR4 (N6305, N6303, N1053, N324, N3971);
not NOT1 (N6306, N6300);
buf BUF1 (N6307, N6286);
or OR3 (N6308, N6305, N2182, N1006);
and AND2 (N6309, N6287, N4871);
nor NOR2 (N6310, N6301, N4747);
and AND2 (N6311, N6294, N4475);
not NOT1 (N6312, N6309);
nand NAND2 (N6313, N6311, N1315);
buf BUF1 (N6314, N6304);
or OR3 (N6315, N6307, N1478, N1298);
xor XOR2 (N6316, N6295, N5897);
nand NAND2 (N6317, N6313, N5191);
not NOT1 (N6318, N6315);
xor XOR2 (N6319, N6310, N2896);
not NOT1 (N6320, N6280);
buf BUF1 (N6321, N6317);
nand NAND2 (N6322, N6316, N2706);
xor XOR2 (N6323, N6321, N2098);
and AND4 (N6324, N6312, N1777, N3826, N1235);
buf BUF1 (N6325, N6318);
buf BUF1 (N6326, N6297);
nor NOR4 (N6327, N6306, N1772, N5717, N4457);
or OR2 (N6328, N6308, N3598);
buf BUF1 (N6329, N6319);
not NOT1 (N6330, N6322);
not NOT1 (N6331, N6324);
nand NAND4 (N6332, N6331, N922, N4275, N3430);
buf BUF1 (N6333, N6320);
xor XOR2 (N6334, N6328, N889);
buf BUF1 (N6335, N6323);
and AND4 (N6336, N6325, N5806, N3745, N207);
or OR3 (N6337, N6332, N3781, N5332);
or OR3 (N6338, N6334, N2955, N3887);
and AND2 (N6339, N6335, N4156);
xor XOR2 (N6340, N6327, N31);
and AND2 (N6341, N6314, N2458);
or OR3 (N6342, N6329, N1765, N1809);
nand NAND3 (N6343, N6333, N4859, N4633);
nand NAND4 (N6344, N6342, N6164, N3690, N3455);
and AND4 (N6345, N6326, N5889, N6252, N5426);
nor NOR3 (N6346, N6339, N4125, N4340);
nor NOR3 (N6347, N6336, N4267, N2192);
or OR4 (N6348, N6346, N4934, N545, N1234);
nor NOR4 (N6349, N6348, N6199, N5688, N493);
and AND4 (N6350, N6338, N5179, N1256, N3225);
or OR4 (N6351, N6340, N3691, N5307, N3761);
xor XOR2 (N6352, N6350, N5677);
or OR4 (N6353, N6330, N3185, N5884, N3974);
xor XOR2 (N6354, N6341, N1428);
nor NOR4 (N6355, N6343, N3287, N2280, N6046);
or OR4 (N6356, N6351, N234, N3579, N3744);
and AND3 (N6357, N6355, N5571, N3064);
buf BUF1 (N6358, N6357);
nand NAND4 (N6359, N6337, N12, N2174, N1443);
or OR4 (N6360, N6349, N1688, N5435, N6019);
or OR2 (N6361, N6344, N2816);
xor XOR2 (N6362, N6352, N5720);
xor XOR2 (N6363, N6356, N4674);
buf BUF1 (N6364, N6347);
or OR4 (N6365, N6364, N106, N5477, N3345);
and AND4 (N6366, N6360, N3256, N2688, N5967);
and AND3 (N6367, N6359, N3185, N2583);
nor NOR4 (N6368, N6363, N3129, N6216, N6190);
nand NAND2 (N6369, N6367, N5171);
nand NAND3 (N6370, N6366, N6146, N2837);
or OR4 (N6371, N6370, N729, N4295, N5031);
or OR2 (N6372, N6371, N4069);
and AND3 (N6373, N6345, N5380, N2044);
nand NAND4 (N6374, N6372, N1655, N3951, N4548);
not NOT1 (N6375, N6361);
buf BUF1 (N6376, N6365);
nand NAND3 (N6377, N6368, N2234, N3381);
not NOT1 (N6378, N6369);
and AND4 (N6379, N6358, N5019, N5946, N1788);
or OR2 (N6380, N6378, N604);
not NOT1 (N6381, N6373);
and AND3 (N6382, N6377, N317, N1197);
nand NAND3 (N6383, N6375, N4498, N947);
nand NAND3 (N6384, N6383, N3616, N4720);
nand NAND3 (N6385, N6354, N4621, N1327);
nor NOR4 (N6386, N6384, N2731, N4272, N3228);
buf BUF1 (N6387, N6381);
and AND4 (N6388, N6353, N5126, N3794, N1309);
xor XOR2 (N6389, N6385, N2899);
and AND2 (N6390, N6376, N4570);
xor XOR2 (N6391, N6362, N4364);
xor XOR2 (N6392, N6388, N1013);
xor XOR2 (N6393, N6389, N5900);
buf BUF1 (N6394, N6390);
and AND3 (N6395, N6387, N1665, N477);
nand NAND2 (N6396, N6391, N3882);
nor NOR4 (N6397, N6379, N5622, N5943, N4241);
nand NAND3 (N6398, N6396, N2042, N733);
and AND4 (N6399, N6393, N5673, N2624, N2529);
buf BUF1 (N6400, N6386);
nand NAND2 (N6401, N6382, N170);
nand NAND4 (N6402, N6399, N332, N70, N3561);
nand NAND4 (N6403, N6394, N2359, N5512, N5467);
and AND2 (N6404, N6401, N3149);
or OR4 (N6405, N6374, N4312, N3925, N1617);
and AND4 (N6406, N6395, N893, N1856, N5227);
buf BUF1 (N6407, N6406);
and AND3 (N6408, N6400, N5555, N5986);
nand NAND3 (N6409, N6392, N5355, N2085);
not NOT1 (N6410, N6403);
and AND2 (N6411, N6407, N5704);
xor XOR2 (N6412, N6408, N1027);
or OR3 (N6413, N6411, N2961, N1815);
not NOT1 (N6414, N6397);
not NOT1 (N6415, N6410);
buf BUF1 (N6416, N6413);
nor NOR2 (N6417, N6405, N4006);
xor XOR2 (N6418, N6412, N4912);
nand NAND4 (N6419, N6417, N3443, N5447, N767);
xor XOR2 (N6420, N6415, N3964);
nor NOR2 (N6421, N6419, N3067);
nor NOR4 (N6422, N6380, N6076, N3598, N4584);
and AND3 (N6423, N6398, N3403, N4039);
nand NAND3 (N6424, N6418, N2588, N1184);
and AND2 (N6425, N6424, N5276);
xor XOR2 (N6426, N6421, N613);
and AND4 (N6427, N6409, N844, N5229, N2511);
and AND2 (N6428, N6425, N2936);
xor XOR2 (N6429, N6423, N772);
xor XOR2 (N6430, N6402, N3449);
buf BUF1 (N6431, N6427);
buf BUF1 (N6432, N6426);
nand NAND3 (N6433, N6430, N3611, N5788);
nand NAND4 (N6434, N6431, N1784, N2366, N1421);
and AND3 (N6435, N6429, N6255, N2562);
and AND4 (N6436, N6433, N3853, N5492, N3492);
or OR3 (N6437, N6422, N4508, N5960);
xor XOR2 (N6438, N6437, N5557);
nand NAND4 (N6439, N6432, N3720, N5829, N3672);
nor NOR2 (N6440, N6420, N5569);
nand NAND4 (N6441, N6440, N324, N4864, N3320);
xor XOR2 (N6442, N6435, N5780);
buf BUF1 (N6443, N6441);
xor XOR2 (N6444, N6434, N3786);
buf BUF1 (N6445, N6414);
not NOT1 (N6446, N6445);
nor NOR4 (N6447, N6428, N3101, N4668, N509);
or OR3 (N6448, N6443, N6346, N5039);
not NOT1 (N6449, N6447);
xor XOR2 (N6450, N6436, N4556);
nand NAND3 (N6451, N6439, N1701, N4083);
buf BUF1 (N6452, N6404);
buf BUF1 (N6453, N6442);
xor XOR2 (N6454, N6444, N4069);
not NOT1 (N6455, N6438);
nand NAND3 (N6456, N6452, N185, N4441);
not NOT1 (N6457, N6456);
and AND4 (N6458, N6454, N5919, N668, N3342);
not NOT1 (N6459, N6416);
xor XOR2 (N6460, N6459, N604);
and AND2 (N6461, N6448, N4568);
xor XOR2 (N6462, N6449, N3899);
buf BUF1 (N6463, N6446);
nor NOR3 (N6464, N6455, N6134, N4961);
buf BUF1 (N6465, N6464);
buf BUF1 (N6466, N6461);
buf BUF1 (N6467, N6466);
buf BUF1 (N6468, N6450);
xor XOR2 (N6469, N6467, N196);
not NOT1 (N6470, N6468);
xor XOR2 (N6471, N6469, N6371);
nand NAND2 (N6472, N6471, N2765);
nor NOR3 (N6473, N6457, N743, N3931);
and AND3 (N6474, N6473, N944, N3958);
buf BUF1 (N6475, N6474);
nand NAND2 (N6476, N6460, N4360);
or OR2 (N6477, N6476, N3269);
and AND2 (N6478, N6465, N4867);
not NOT1 (N6479, N6462);
not NOT1 (N6480, N6470);
xor XOR2 (N6481, N6451, N6240);
and AND2 (N6482, N6478, N5764);
buf BUF1 (N6483, N6458);
and AND4 (N6484, N6482, N2821, N5338, N4857);
or OR3 (N6485, N6480, N5741, N3287);
nand NAND2 (N6486, N6477, N3241);
or OR4 (N6487, N6485, N4505, N3896, N5568);
buf BUF1 (N6488, N6484);
buf BUF1 (N6489, N6475);
nor NOR3 (N6490, N6479, N2166, N4376);
and AND4 (N6491, N6481, N1520, N2841, N1733);
and AND3 (N6492, N6472, N6356, N18);
and AND4 (N6493, N6463, N548, N5454, N2182);
nor NOR2 (N6494, N6453, N6288);
nand NAND4 (N6495, N6488, N1961, N1066, N1202);
not NOT1 (N6496, N6494);
nand NAND4 (N6497, N6487, N1194, N2594, N5090);
nand NAND2 (N6498, N6491, N2956);
xor XOR2 (N6499, N6486, N4023);
nand NAND2 (N6500, N6490, N6058);
and AND2 (N6501, N6492, N3483);
buf BUF1 (N6502, N6493);
not NOT1 (N6503, N6498);
or OR4 (N6504, N6483, N4984, N5554, N1703);
buf BUF1 (N6505, N6503);
not NOT1 (N6506, N6499);
nor NOR3 (N6507, N6500, N5154, N4662);
and AND3 (N6508, N6501, N5225, N4650);
or OR3 (N6509, N6506, N2285, N2782);
nand NAND4 (N6510, N6504, N2553, N2571, N5903);
nor NOR3 (N6511, N6509, N1268, N6035);
not NOT1 (N6512, N6505);
and AND2 (N6513, N6512, N492);
and AND4 (N6514, N6495, N3230, N5010, N1864);
xor XOR2 (N6515, N6502, N5114);
not NOT1 (N6516, N6511);
buf BUF1 (N6517, N6514);
xor XOR2 (N6518, N6508, N6210);
buf BUF1 (N6519, N6510);
not NOT1 (N6520, N6515);
or OR3 (N6521, N6520, N1919, N3074);
buf BUF1 (N6522, N6507);
nor NOR4 (N6523, N6517, N5709, N1432, N6346);
buf BUF1 (N6524, N6522);
and AND4 (N6525, N6521, N4932, N6473, N1984);
or OR3 (N6526, N6489, N3750, N2728);
xor XOR2 (N6527, N6496, N4821);
or OR3 (N6528, N6518, N1648, N5402);
buf BUF1 (N6529, N6523);
or OR2 (N6530, N6525, N3732);
nor NOR2 (N6531, N6516, N693);
buf BUF1 (N6532, N6530);
and AND2 (N6533, N6529, N3539);
xor XOR2 (N6534, N6526, N3414);
buf BUF1 (N6535, N6527);
buf BUF1 (N6536, N6531);
xor XOR2 (N6537, N6524, N763);
nand NAND4 (N6538, N6513, N2624, N2024, N1434);
not NOT1 (N6539, N6538);
nand NAND2 (N6540, N6497, N635);
nand NAND4 (N6541, N6539, N4786, N3007, N1268);
nand NAND3 (N6542, N6540, N5526, N2153);
not NOT1 (N6543, N6535);
or OR3 (N6544, N6534, N5831, N5840);
nor NOR2 (N6545, N6541, N4292);
nand NAND4 (N6546, N6545, N3622, N3940, N1649);
nand NAND3 (N6547, N6536, N6442, N672);
or OR4 (N6548, N6544, N6352, N1565, N6120);
or OR2 (N6549, N6547, N4622);
nor NOR3 (N6550, N6532, N2641, N3529);
not NOT1 (N6551, N6537);
not NOT1 (N6552, N6549);
and AND2 (N6553, N6550, N5335);
buf BUF1 (N6554, N6543);
xor XOR2 (N6555, N6546, N998);
buf BUF1 (N6556, N6519);
or OR4 (N6557, N6554, N1586, N1477, N1535);
nor NOR3 (N6558, N6556, N3447, N4789);
not NOT1 (N6559, N6542);
and AND4 (N6560, N6552, N2559, N1360, N5831);
nand NAND3 (N6561, N6551, N2479, N121);
not NOT1 (N6562, N6533);
nand NAND3 (N6563, N6528, N3389, N2516);
xor XOR2 (N6564, N6555, N5374);
xor XOR2 (N6565, N6563, N3400);
and AND2 (N6566, N6548, N4879);
nor NOR4 (N6567, N6564, N1504, N5074, N4955);
xor XOR2 (N6568, N6566, N4522);
nor NOR4 (N6569, N6565, N5875, N3234, N378);
and AND3 (N6570, N6569, N1815, N4968);
xor XOR2 (N6571, N6562, N1020);
and AND3 (N6572, N6558, N4259, N6000);
nand NAND4 (N6573, N6561, N3060, N4802, N4391);
nand NAND3 (N6574, N6568, N3558, N947);
xor XOR2 (N6575, N6574, N5337);
nand NAND4 (N6576, N6557, N1179, N3261, N385);
not NOT1 (N6577, N6559);
and AND3 (N6578, N6577, N646, N5832);
nor NOR3 (N6579, N6570, N5881, N1420);
buf BUF1 (N6580, N6553);
nand NAND2 (N6581, N6575, N238);
nor NOR2 (N6582, N6571, N377);
not NOT1 (N6583, N6578);
or OR4 (N6584, N6576, N6282, N540, N4444);
not NOT1 (N6585, N6580);
not NOT1 (N6586, N6583);
or OR2 (N6587, N6572, N3365);
xor XOR2 (N6588, N6579, N1541);
or OR2 (N6589, N6585, N2469);
not NOT1 (N6590, N6587);
nor NOR3 (N6591, N6586, N230, N3310);
or OR3 (N6592, N6584, N6028, N3945);
nor NOR4 (N6593, N6567, N4858, N3457, N954);
and AND4 (N6594, N6590, N210, N691, N2805);
or OR3 (N6595, N6589, N3366, N6107);
and AND3 (N6596, N6594, N6528, N228);
and AND2 (N6597, N6595, N1428);
buf BUF1 (N6598, N6596);
and AND3 (N6599, N6592, N2910, N1550);
or OR4 (N6600, N6597, N4885, N5138, N6260);
xor XOR2 (N6601, N6600, N4164);
buf BUF1 (N6602, N6588);
xor XOR2 (N6603, N6582, N5182);
buf BUF1 (N6604, N6602);
nor NOR3 (N6605, N6591, N706, N6140);
buf BUF1 (N6606, N6560);
buf BUF1 (N6607, N6605);
and AND3 (N6608, N6606, N2290, N5407);
nand NAND4 (N6609, N6601, N956, N3892, N6270);
or OR3 (N6610, N6609, N3012, N746);
and AND4 (N6611, N6604, N1958, N6538, N3868);
nand NAND4 (N6612, N6598, N4459, N3537, N3920);
nor NOR4 (N6613, N6581, N6315, N3217, N3185);
nor NOR3 (N6614, N6593, N1259, N2700);
xor XOR2 (N6615, N6608, N1780);
nand NAND3 (N6616, N6614, N6462, N4144);
not NOT1 (N6617, N6613);
and AND2 (N6618, N6610, N2394);
xor XOR2 (N6619, N6603, N5083);
buf BUF1 (N6620, N6619);
not NOT1 (N6621, N6617);
not NOT1 (N6622, N6611);
nand NAND3 (N6623, N6618, N4216, N4249);
nand NAND2 (N6624, N6573, N2832);
and AND4 (N6625, N6624, N232, N3854, N2133);
nand NAND3 (N6626, N6615, N3364, N4516);
and AND2 (N6627, N6599, N5644);
or OR4 (N6628, N6627, N4883, N4882, N5901);
xor XOR2 (N6629, N6616, N2618);
nand NAND2 (N6630, N6612, N1150);
and AND3 (N6631, N6607, N1809, N2011);
xor XOR2 (N6632, N6628, N2906);
buf BUF1 (N6633, N6626);
or OR4 (N6634, N6631, N6365, N633, N4101);
nand NAND3 (N6635, N6625, N5166, N1739);
nand NAND4 (N6636, N6633, N101, N2981, N996);
buf BUF1 (N6637, N6622);
and AND4 (N6638, N6623, N2221, N1858, N5955);
xor XOR2 (N6639, N6629, N4585);
buf BUF1 (N6640, N6639);
buf BUF1 (N6641, N6636);
or OR4 (N6642, N6621, N2018, N2938, N1073);
not NOT1 (N6643, N6642);
or OR3 (N6644, N6643, N5436, N1155);
buf BUF1 (N6645, N6634);
or OR2 (N6646, N6637, N3482);
nor NOR3 (N6647, N6638, N1823, N5641);
and AND3 (N6648, N6632, N2246, N5821);
nor NOR3 (N6649, N6630, N3376, N10);
not NOT1 (N6650, N6635);
nand NAND3 (N6651, N6645, N2154, N1215);
buf BUF1 (N6652, N6650);
not NOT1 (N6653, N6646);
nand NAND4 (N6654, N6644, N709, N637, N3517);
nand NAND4 (N6655, N6648, N5057, N1741, N2873);
nand NAND4 (N6656, N6641, N6455, N822, N1725);
not NOT1 (N6657, N6649);
and AND3 (N6658, N6653, N4195, N3809);
xor XOR2 (N6659, N6640, N2939);
buf BUF1 (N6660, N6655);
nand NAND4 (N6661, N6651, N2147, N2717, N2388);
nor NOR4 (N6662, N6656, N2085, N3451, N1208);
not NOT1 (N6663, N6652);
nor NOR2 (N6664, N6663, N5490);
buf BUF1 (N6665, N6657);
nand NAND2 (N6666, N6654, N1994);
and AND4 (N6667, N6661, N2617, N2154, N3184);
or OR3 (N6668, N6647, N761, N4934);
and AND2 (N6669, N6662, N288);
buf BUF1 (N6670, N6664);
not NOT1 (N6671, N6670);
nand NAND3 (N6672, N6668, N201, N1547);
buf BUF1 (N6673, N6671);
or OR2 (N6674, N6659, N959);
nand NAND3 (N6675, N6665, N4629, N796);
buf BUF1 (N6676, N6669);
buf BUF1 (N6677, N6673);
or OR4 (N6678, N6620, N2622, N6175, N4739);
nand NAND2 (N6679, N6658, N4478);
xor XOR2 (N6680, N6672, N499);
and AND3 (N6681, N6675, N4943, N757);
or OR3 (N6682, N6676, N3085, N822);
xor XOR2 (N6683, N6667, N4308);
xor XOR2 (N6684, N6681, N3067);
xor XOR2 (N6685, N6660, N6605);
buf BUF1 (N6686, N6684);
nand NAND2 (N6687, N6682, N133);
or OR2 (N6688, N6666, N2505);
or OR3 (N6689, N6674, N3462, N2316);
not NOT1 (N6690, N6678);
nor NOR2 (N6691, N6689, N3549);
nand NAND2 (N6692, N6685, N361);
not NOT1 (N6693, N6677);
or OR2 (N6694, N6687, N1757);
not NOT1 (N6695, N6680);
nand NAND3 (N6696, N6695, N3295, N2901);
xor XOR2 (N6697, N6688, N3714);
or OR4 (N6698, N6696, N5875, N2650, N1581);
or OR3 (N6699, N6691, N2497, N1604);
nand NAND3 (N6700, N6692, N1433, N3446);
buf BUF1 (N6701, N6693);
not NOT1 (N6702, N6690);
buf BUF1 (N6703, N6700);
buf BUF1 (N6704, N6698);
buf BUF1 (N6705, N6694);
nand NAND2 (N6706, N6679, N1691);
nor NOR2 (N6707, N6699, N1590);
or OR4 (N6708, N6683, N3955, N3698, N1438);
xor XOR2 (N6709, N6701, N3875);
not NOT1 (N6710, N6702);
and AND3 (N6711, N6697, N1948, N4668);
or OR3 (N6712, N6706, N925, N4518);
nand NAND3 (N6713, N6686, N1756, N2346);
and AND2 (N6714, N6703, N3983);
nand NAND3 (N6715, N6708, N638, N493);
nand NAND2 (N6716, N6704, N3121);
not NOT1 (N6717, N6716);
buf BUF1 (N6718, N6717);
nor NOR2 (N6719, N6711, N6450);
and AND4 (N6720, N6709, N5253, N6717, N5409);
or OR4 (N6721, N6712, N1877, N1078, N634);
buf BUF1 (N6722, N6721);
not NOT1 (N6723, N6707);
not NOT1 (N6724, N6718);
not NOT1 (N6725, N6723);
nand NAND3 (N6726, N6714, N1503, N3442);
xor XOR2 (N6727, N6713, N715);
not NOT1 (N6728, N6719);
and AND3 (N6729, N6727, N3473, N3823);
buf BUF1 (N6730, N6710);
nand NAND4 (N6731, N6729, N5985, N3357, N2474);
xor XOR2 (N6732, N6715, N6052);
not NOT1 (N6733, N6726);
or OR3 (N6734, N6722, N3041, N5157);
nand NAND2 (N6735, N6728, N4662);
not NOT1 (N6736, N6705);
and AND4 (N6737, N6731, N825, N450, N1301);
or OR4 (N6738, N6735, N2002, N2059, N2357);
not NOT1 (N6739, N6732);
not NOT1 (N6740, N6730);
nand NAND4 (N6741, N6720, N4359, N4303, N83);
xor XOR2 (N6742, N6736, N5516);
buf BUF1 (N6743, N6741);
and AND3 (N6744, N6737, N6741, N4371);
or OR4 (N6745, N6734, N6570, N5362, N3876);
nand NAND2 (N6746, N6733, N735);
buf BUF1 (N6747, N6746);
nor NOR2 (N6748, N6745, N6543);
not NOT1 (N6749, N6744);
buf BUF1 (N6750, N6739);
buf BUF1 (N6751, N6748);
not NOT1 (N6752, N6740);
nand NAND2 (N6753, N6751, N1150);
buf BUF1 (N6754, N6742);
nor NOR3 (N6755, N6750, N807, N3470);
and AND2 (N6756, N6752, N3007);
and AND3 (N6757, N6724, N2703, N4347);
buf BUF1 (N6758, N6757);
not NOT1 (N6759, N6753);
nor NOR3 (N6760, N6749, N2609, N6406);
nand NAND3 (N6761, N6760, N5296, N2548);
or OR3 (N6762, N6758, N4268, N4858);
buf BUF1 (N6763, N6738);
nand NAND2 (N6764, N6743, N4255);
nor NOR3 (N6765, N6756, N1315, N510);
not NOT1 (N6766, N6764);
or OR2 (N6767, N6759, N2926);
or OR2 (N6768, N6763, N3567);
and AND4 (N6769, N6765, N929, N2523, N3196);
and AND3 (N6770, N6762, N3838, N2737);
nor NOR4 (N6771, N6770, N3634, N5094, N3206);
xor XOR2 (N6772, N6747, N4496);
xor XOR2 (N6773, N6772, N1086);
and AND2 (N6774, N6773, N5444);
and AND4 (N6775, N6761, N4555, N2924, N6280);
nand NAND4 (N6776, N6755, N6281, N4890, N4941);
nand NAND4 (N6777, N6766, N648, N1723, N3437);
not NOT1 (N6778, N6771);
nor NOR3 (N6779, N6774, N6321, N604);
not NOT1 (N6780, N6775);
or OR4 (N6781, N6779, N283, N5350, N566);
nor NOR2 (N6782, N6769, N2981);
not NOT1 (N6783, N6768);
buf BUF1 (N6784, N6783);
or OR4 (N6785, N6767, N2215, N648, N5143);
xor XOR2 (N6786, N6780, N1111);
not NOT1 (N6787, N6776);
nand NAND4 (N6788, N6778, N5530, N4708, N1762);
xor XOR2 (N6789, N6781, N1973);
nand NAND4 (N6790, N6785, N3473, N891, N1898);
and AND4 (N6791, N6782, N358, N4073, N4877);
nand NAND4 (N6792, N6788, N325, N4165, N6042);
nor NOR2 (N6793, N6725, N6454);
xor XOR2 (N6794, N6790, N1796);
nand NAND2 (N6795, N6777, N6410);
buf BUF1 (N6796, N6754);
or OR2 (N6797, N6786, N5965);
nand NAND3 (N6798, N6787, N213, N4817);
not NOT1 (N6799, N6796);
or OR2 (N6800, N6792, N563);
xor XOR2 (N6801, N6799, N106);
nand NAND3 (N6802, N6800, N167, N6025);
xor XOR2 (N6803, N6791, N6124);
xor XOR2 (N6804, N6794, N3053);
nor NOR3 (N6805, N6793, N2431, N4942);
not NOT1 (N6806, N6801);
nand NAND3 (N6807, N6798, N5858, N4084);
or OR2 (N6808, N6806, N2319);
buf BUF1 (N6809, N6795);
and AND2 (N6810, N6807, N3452);
nor NOR3 (N6811, N6803, N3487, N5986);
buf BUF1 (N6812, N6805);
and AND2 (N6813, N6802, N2632);
nor NOR4 (N6814, N6809, N1405, N6198, N6689);
buf BUF1 (N6815, N6814);
xor XOR2 (N6816, N6811, N680);
xor XOR2 (N6817, N6804, N577);
and AND4 (N6818, N6784, N305, N3519, N3046);
or OR2 (N6819, N6810, N2978);
not NOT1 (N6820, N6812);
not NOT1 (N6821, N6797);
buf BUF1 (N6822, N6817);
not NOT1 (N6823, N6818);
nand NAND4 (N6824, N6820, N5752, N3484, N1608);
nand NAND4 (N6825, N6822, N2545, N4431, N6494);
not NOT1 (N6826, N6821);
or OR3 (N6827, N6808, N2256, N3320);
and AND3 (N6828, N6816, N258, N5519);
nand NAND3 (N6829, N6815, N1230, N289);
nor NOR3 (N6830, N6828, N3494, N461);
buf BUF1 (N6831, N6829);
nand NAND4 (N6832, N6789, N454, N918, N1476);
buf BUF1 (N6833, N6832);
nand NAND4 (N6834, N6823, N647, N172, N51);
buf BUF1 (N6835, N6825);
or OR4 (N6836, N6835, N3328, N2523, N4928);
buf BUF1 (N6837, N6827);
nor NOR2 (N6838, N6831, N2553);
xor XOR2 (N6839, N6838, N4543);
not NOT1 (N6840, N6839);
nand NAND2 (N6841, N6813, N5348);
nand NAND3 (N6842, N6830, N2472, N2650);
and AND2 (N6843, N6834, N965);
nor NOR3 (N6844, N6840, N2698, N5947);
not NOT1 (N6845, N6844);
xor XOR2 (N6846, N6833, N1304);
xor XOR2 (N6847, N6826, N984);
and AND3 (N6848, N6819, N5716, N4930);
not NOT1 (N6849, N6841);
or OR3 (N6850, N6845, N3291, N182);
nand NAND2 (N6851, N6836, N3404);
and AND2 (N6852, N6843, N4148);
nand NAND4 (N6853, N6837, N2239, N4584, N2565);
xor XOR2 (N6854, N6849, N6103);
and AND4 (N6855, N6853, N700, N1793, N2388);
xor XOR2 (N6856, N6851, N710);
and AND3 (N6857, N6846, N5460, N5441);
and AND2 (N6858, N6852, N4851);
buf BUF1 (N6859, N6842);
xor XOR2 (N6860, N6857, N3859);
and AND4 (N6861, N6848, N4003, N4888, N4705);
not NOT1 (N6862, N6854);
and AND3 (N6863, N6860, N3009, N6294);
and AND2 (N6864, N6859, N3631);
not NOT1 (N6865, N6855);
or OR2 (N6866, N6862, N1413);
nand NAND3 (N6867, N6866, N3942, N4708);
not NOT1 (N6868, N6847);
not NOT1 (N6869, N6858);
xor XOR2 (N6870, N6861, N3303);
nor NOR3 (N6871, N6864, N2317, N6261);
and AND4 (N6872, N6865, N2149, N4317, N407);
and AND3 (N6873, N6856, N3938, N6346);
nor NOR3 (N6874, N6850, N6549, N5883);
xor XOR2 (N6875, N6874, N2737);
nor NOR4 (N6876, N6863, N2046, N6115, N4725);
buf BUF1 (N6877, N6867);
or OR4 (N6878, N6870, N2067, N175, N36);
nor NOR4 (N6879, N6878, N2727, N3886, N6601);
nor NOR2 (N6880, N6868, N5052);
xor XOR2 (N6881, N6873, N4730);
not NOT1 (N6882, N6871);
and AND3 (N6883, N6875, N679, N4686);
xor XOR2 (N6884, N6877, N5040);
not NOT1 (N6885, N6869);
buf BUF1 (N6886, N6872);
nor NOR4 (N6887, N6882, N2786, N4336, N5880);
or OR4 (N6888, N6879, N3682, N3054, N4853);
buf BUF1 (N6889, N6884);
xor XOR2 (N6890, N6887, N1422);
or OR4 (N6891, N6886, N4579, N653, N2570);
xor XOR2 (N6892, N6885, N3726);
nor NOR3 (N6893, N6889, N2526, N255);
nor NOR2 (N6894, N6893, N1232);
buf BUF1 (N6895, N6891);
not NOT1 (N6896, N6883);
and AND4 (N6897, N6894, N1065, N1849, N2215);
nand NAND3 (N6898, N6895, N2653, N4846);
not NOT1 (N6899, N6898);
and AND3 (N6900, N6896, N3466, N4500);
nand NAND2 (N6901, N6892, N1793);
nor NOR3 (N6902, N6880, N5669, N1278);
nand NAND3 (N6903, N6899, N838, N6383);
nand NAND3 (N6904, N6900, N2846, N2847);
or OR2 (N6905, N6888, N5553);
and AND3 (N6906, N6824, N4536, N2119);
and AND4 (N6907, N6890, N6724, N396, N1701);
and AND3 (N6908, N6902, N5742, N2397);
nor NOR2 (N6909, N6876, N1527);
not NOT1 (N6910, N6881);
xor XOR2 (N6911, N6897, N1045);
buf BUF1 (N6912, N6910);
buf BUF1 (N6913, N6905);
not NOT1 (N6914, N6908);
and AND2 (N6915, N6901, N4392);
and AND3 (N6916, N6911, N6031, N1954);
not NOT1 (N6917, N6912);
not NOT1 (N6918, N6903);
buf BUF1 (N6919, N6909);
or OR4 (N6920, N6914, N2754, N1774, N1);
nor NOR2 (N6921, N6916, N2471);
or OR2 (N6922, N6915, N1462);
not NOT1 (N6923, N6907);
buf BUF1 (N6924, N6921);
and AND3 (N6925, N6917, N5457, N3427);
or OR3 (N6926, N6925, N2331, N4653);
not NOT1 (N6927, N6904);
or OR3 (N6928, N6919, N3127, N4308);
nor NOR2 (N6929, N6926, N2123);
xor XOR2 (N6930, N6913, N5015);
nand NAND2 (N6931, N6930, N4013);
nand NAND4 (N6932, N6922, N3714, N3686, N5676);
and AND3 (N6933, N6932, N507, N6458);
not NOT1 (N6934, N6924);
xor XOR2 (N6935, N6931, N4675);
buf BUF1 (N6936, N6933);
buf BUF1 (N6937, N6934);
and AND4 (N6938, N6937, N6752, N119, N6697);
and AND4 (N6939, N6918, N96, N850, N24);
nand NAND2 (N6940, N6939, N4365);
not NOT1 (N6941, N6938);
nor NOR4 (N6942, N6928, N533, N5578, N2280);
nand NAND2 (N6943, N6940, N3886);
buf BUF1 (N6944, N6942);
buf BUF1 (N6945, N6929);
or OR2 (N6946, N6943, N5058);
and AND4 (N6947, N6944, N6455, N6742, N3454);
or OR2 (N6948, N6945, N1305);
or OR2 (N6949, N6936, N327);
not NOT1 (N6950, N6946);
or OR4 (N6951, N6935, N323, N3184, N2732);
or OR3 (N6952, N6948, N3863, N1904);
nand NAND4 (N6953, N6949, N3865, N1416, N3978);
nor NOR3 (N6954, N6927, N5574, N5060);
not NOT1 (N6955, N6941);
and AND2 (N6956, N6955, N3170);
nand NAND4 (N6957, N6923, N1840, N786, N1494);
nor NOR4 (N6958, N6953, N5141, N4127, N2355);
buf BUF1 (N6959, N6952);
and AND3 (N6960, N6958, N1648, N1986);
not NOT1 (N6961, N6954);
buf BUF1 (N6962, N6956);
not NOT1 (N6963, N6951);
buf BUF1 (N6964, N6959);
not NOT1 (N6965, N6950);
or OR3 (N6966, N6963, N5558, N6766);
buf BUF1 (N6967, N6947);
or OR2 (N6968, N6967, N710);
buf BUF1 (N6969, N6960);
not NOT1 (N6970, N6965);
and AND4 (N6971, N6957, N5161, N6184, N6968);
xor XOR2 (N6972, N7, N3701);
not NOT1 (N6973, N6964);
not NOT1 (N6974, N6961);
xor XOR2 (N6975, N6969, N4273);
xor XOR2 (N6976, N6970, N6544);
buf BUF1 (N6977, N6972);
not NOT1 (N6978, N6966);
or OR4 (N6979, N6962, N5325, N5954, N5234);
nor NOR3 (N6980, N6977, N1197, N6684);
xor XOR2 (N6981, N6973, N5250);
not NOT1 (N6982, N6978);
buf BUF1 (N6983, N6974);
and AND3 (N6984, N6920, N1914, N2754);
or OR4 (N6985, N6906, N1460, N2057, N782);
buf BUF1 (N6986, N6976);
nor NOR2 (N6987, N6981, N2235);
and AND3 (N6988, N6987, N3241, N6931);
or OR2 (N6989, N6982, N2595);
xor XOR2 (N6990, N6975, N4003);
nor NOR4 (N6991, N6980, N2462, N2009, N3223);
nand NAND2 (N6992, N6990, N2572);
buf BUF1 (N6993, N6971);
and AND3 (N6994, N6992, N6139, N1015);
buf BUF1 (N6995, N6983);
xor XOR2 (N6996, N6991, N3079);
and AND2 (N6997, N6996, N2942);
nand NAND3 (N6998, N6979, N6551, N6033);
nand NAND2 (N6999, N6994, N4876);
or OR4 (N7000, N6997, N5584, N1856, N6960);
nand NAND2 (N7001, N6984, N5348);
nand NAND2 (N7002, N6985, N1863);
xor XOR2 (N7003, N6986, N5759);
nor NOR3 (N7004, N6999, N2756, N2912);
xor XOR2 (N7005, N7001, N1544);
buf BUF1 (N7006, N6988);
and AND2 (N7007, N7003, N4230);
nor NOR4 (N7008, N7007, N2035, N6578, N2509);
and AND3 (N7009, N7004, N3277, N6695);
and AND3 (N7010, N7005, N2290, N2133);
nor NOR2 (N7011, N7008, N74);
not NOT1 (N7012, N7000);
nor NOR2 (N7013, N7011, N3964);
buf BUF1 (N7014, N6995);
not NOT1 (N7015, N7012);
nand NAND3 (N7016, N6998, N3207, N6947);
not NOT1 (N7017, N7006);
nor NOR4 (N7018, N7002, N5851, N6208, N5916);
buf BUF1 (N7019, N7014);
buf BUF1 (N7020, N7018);
nand NAND4 (N7021, N7015, N368, N6975, N890);
xor XOR2 (N7022, N7017, N2879);
buf BUF1 (N7023, N7013);
nand NAND4 (N7024, N7009, N1192, N2767, N1909);
xor XOR2 (N7025, N6993, N6274);
nand NAND3 (N7026, N7023, N870, N2194);
not NOT1 (N7027, N7022);
xor XOR2 (N7028, N7016, N2045);
xor XOR2 (N7029, N7020, N2117);
or OR2 (N7030, N7021, N3098);
and AND3 (N7031, N7025, N2687, N6602);
xor XOR2 (N7032, N7029, N6197);
or OR4 (N7033, N7030, N6833, N3021, N2336);
nand NAND3 (N7034, N7010, N3595, N6334);
not NOT1 (N7035, N6989);
buf BUF1 (N7036, N7033);
buf BUF1 (N7037, N7035);
nand NAND4 (N7038, N7027, N3852, N1898, N917);
xor XOR2 (N7039, N7028, N1348);
and AND3 (N7040, N7032, N2678, N725);
xor XOR2 (N7041, N7036, N1530);
nor NOR2 (N7042, N7024, N2230);
nor NOR3 (N7043, N7040, N2622, N6955);
nor NOR4 (N7044, N7019, N6636, N4657, N6745);
nor NOR2 (N7045, N7042, N5890);
nor NOR2 (N7046, N7037, N3280);
xor XOR2 (N7047, N7026, N6497);
and AND3 (N7048, N7041, N5739, N4738);
nor NOR2 (N7049, N7038, N5648);
buf BUF1 (N7050, N7049);
nor NOR2 (N7051, N7050, N4067);
buf BUF1 (N7052, N7047);
not NOT1 (N7053, N7043);
xor XOR2 (N7054, N7053, N1808);
nand NAND2 (N7055, N7034, N5744);
or OR4 (N7056, N7055, N4931, N6145, N2051);
buf BUF1 (N7057, N7048);
not NOT1 (N7058, N7031);
xor XOR2 (N7059, N7056, N3907);
and AND2 (N7060, N7044, N2873);
or OR3 (N7061, N7052, N3588, N2513);
not NOT1 (N7062, N7058);
and AND4 (N7063, N7061, N4254, N5528, N2448);
nand NAND4 (N7064, N7062, N4295, N2236, N2994);
nor NOR2 (N7065, N7054, N230);
or OR2 (N7066, N7046, N1229);
not NOT1 (N7067, N7065);
nor NOR4 (N7068, N7051, N4307, N4514, N5419);
buf BUF1 (N7069, N7066);
xor XOR2 (N7070, N7057, N1626);
not NOT1 (N7071, N7067);
xor XOR2 (N7072, N7045, N3940);
or OR3 (N7073, N7063, N237, N1441);
not NOT1 (N7074, N7071);
or OR2 (N7075, N7070, N5247);
and AND2 (N7076, N7075, N6236);
and AND4 (N7077, N7069, N5148, N1626, N2354);
nor NOR3 (N7078, N7060, N1477, N134);
nand NAND3 (N7079, N7064, N1546, N3516);
buf BUF1 (N7080, N7077);
buf BUF1 (N7081, N7074);
or OR4 (N7082, N7039, N55, N736, N759);
nand NAND2 (N7083, N7082, N2152);
not NOT1 (N7084, N7083);
not NOT1 (N7085, N7073);
not NOT1 (N7086, N7084);
buf BUF1 (N7087, N7080);
xor XOR2 (N7088, N7076, N6205);
not NOT1 (N7089, N7086);
nor NOR3 (N7090, N7089, N6769, N3817);
buf BUF1 (N7091, N7059);
buf BUF1 (N7092, N7072);
nand NAND2 (N7093, N7079, N5262);
not NOT1 (N7094, N7081);
not NOT1 (N7095, N7088);
xor XOR2 (N7096, N7094, N4324);
nand NAND3 (N7097, N7068, N311, N6137);
and AND2 (N7098, N7091, N4735);
xor XOR2 (N7099, N7097, N1102);
nand NAND2 (N7100, N7092, N5479);
or OR3 (N7101, N7093, N4492, N5773);
buf BUF1 (N7102, N7096);
nor NOR3 (N7103, N7087, N3224, N2750);
not NOT1 (N7104, N7090);
not NOT1 (N7105, N7103);
or OR3 (N7106, N7098, N5749, N206);
or OR3 (N7107, N7105, N418, N2573);
nor NOR2 (N7108, N7095, N6359);
or OR3 (N7109, N7100, N1493, N3272);
or OR2 (N7110, N7078, N1202);
nor NOR3 (N7111, N7106, N158, N2253);
buf BUF1 (N7112, N7104);
xor XOR2 (N7113, N7101, N1811);
not NOT1 (N7114, N7113);
and AND2 (N7115, N7085, N3510);
xor XOR2 (N7116, N7108, N1235);
nand NAND4 (N7117, N7112, N4694, N3088, N137);
or OR4 (N7118, N7099, N5526, N4362, N996);
xor XOR2 (N7119, N7117, N2848);
not NOT1 (N7120, N7119);
xor XOR2 (N7121, N7102, N1936);
or OR4 (N7122, N7116, N2313, N4007, N5020);
not NOT1 (N7123, N7111);
xor XOR2 (N7124, N7110, N2284);
xor XOR2 (N7125, N7107, N5798);
buf BUF1 (N7126, N7114);
and AND3 (N7127, N7121, N7083, N1332);
xor XOR2 (N7128, N7122, N4277);
not NOT1 (N7129, N7128);
xor XOR2 (N7130, N7118, N6668);
nand NAND3 (N7131, N7127, N6953, N881);
buf BUF1 (N7132, N7124);
xor XOR2 (N7133, N7126, N462);
not NOT1 (N7134, N7130);
or OR3 (N7135, N7120, N1142, N4617);
nand NAND3 (N7136, N7123, N562, N4489);
nand NAND4 (N7137, N7109, N5359, N6960, N1154);
nand NAND3 (N7138, N7115, N1227, N6666);
buf BUF1 (N7139, N7135);
or OR2 (N7140, N7132, N6960);
or OR4 (N7141, N7138, N1576, N6578, N4453);
nor NOR3 (N7142, N7129, N2844, N889);
xor XOR2 (N7143, N7142, N2807);
buf BUF1 (N7144, N7125);
or OR3 (N7145, N7133, N6988, N6480);
nor NOR3 (N7146, N7145, N2686, N4550);
nor NOR3 (N7147, N7143, N4334, N3747);
or OR3 (N7148, N7140, N3737, N2486);
not NOT1 (N7149, N7146);
xor XOR2 (N7150, N7147, N1601);
nand NAND2 (N7151, N7137, N4416);
nor NOR3 (N7152, N7131, N4376, N3122);
xor XOR2 (N7153, N7148, N4278);
buf BUF1 (N7154, N7150);
buf BUF1 (N7155, N7151);
not NOT1 (N7156, N7136);
xor XOR2 (N7157, N7139, N3805);
nand NAND4 (N7158, N7144, N3919, N3133, N2103);
buf BUF1 (N7159, N7157);
not NOT1 (N7160, N7152);
and AND3 (N7161, N7149, N5244, N1651);
nand NAND4 (N7162, N7156, N7130, N2355, N1411);
or OR4 (N7163, N7159, N2694, N5891, N1879);
or OR2 (N7164, N7158, N2388);
nor NOR3 (N7165, N7155, N3234, N1613);
nor NOR2 (N7166, N7163, N5492);
or OR3 (N7167, N7134, N7118, N683);
not NOT1 (N7168, N7160);
and AND2 (N7169, N7162, N3313);
nand NAND2 (N7170, N7161, N6682);
nand NAND3 (N7171, N7166, N4717, N5596);
not NOT1 (N7172, N7168);
buf BUF1 (N7173, N7165);
or OR3 (N7174, N7171, N7001, N3261);
or OR4 (N7175, N7153, N676, N4948, N262);
nand NAND4 (N7176, N7170, N4882, N3448, N5111);
xor XOR2 (N7177, N7172, N6680);
xor XOR2 (N7178, N7176, N6329);
or OR2 (N7179, N7154, N196);
or OR2 (N7180, N7169, N4638);
nor NOR2 (N7181, N7167, N5559);
buf BUF1 (N7182, N7141);
xor XOR2 (N7183, N7164, N1008);
buf BUF1 (N7184, N7175);
and AND2 (N7185, N7174, N1628);
not NOT1 (N7186, N7173);
not NOT1 (N7187, N7177);
or OR2 (N7188, N7179, N4083);
or OR4 (N7189, N7188, N5228, N596, N3731);
nor NOR4 (N7190, N7181, N965, N5576, N3837);
not NOT1 (N7191, N7178);
nor NOR3 (N7192, N7186, N6740, N6849);
not NOT1 (N7193, N7182);
nand NAND2 (N7194, N7185, N6499);
xor XOR2 (N7195, N7189, N5074);
or OR2 (N7196, N7190, N862);
xor XOR2 (N7197, N7191, N474);
buf BUF1 (N7198, N7184);
nand NAND4 (N7199, N7183, N3570, N2463, N532);
not NOT1 (N7200, N7196);
and AND3 (N7201, N7197, N5702, N1980);
nand NAND4 (N7202, N7187, N143, N4313, N4758);
not NOT1 (N7203, N7180);
nand NAND2 (N7204, N7194, N5952);
nor NOR2 (N7205, N7193, N3706);
or OR3 (N7206, N7205, N3958, N1668);
and AND2 (N7207, N7192, N1778);
and AND3 (N7208, N7199, N4589, N3654);
not NOT1 (N7209, N7201);
nand NAND2 (N7210, N7195, N4458);
and AND3 (N7211, N7198, N1522, N5603);
not NOT1 (N7212, N7209);
nor NOR2 (N7213, N7203, N1503);
nor NOR2 (N7214, N7208, N2644);
or OR2 (N7215, N7204, N6118);
not NOT1 (N7216, N7214);
not NOT1 (N7217, N7215);
xor XOR2 (N7218, N7213, N1950);
not NOT1 (N7219, N7202);
and AND4 (N7220, N7200, N273, N7164, N4112);
nand NAND4 (N7221, N7216, N283, N5532, N3403);
or OR4 (N7222, N7207, N6890, N6019, N5068);
or OR4 (N7223, N7206, N744, N7160, N2497);
and AND4 (N7224, N7221, N3864, N1655, N6004);
xor XOR2 (N7225, N7222, N804);
nand NAND3 (N7226, N7219, N274, N4758);
xor XOR2 (N7227, N7210, N2087);
or OR2 (N7228, N7218, N3292);
nor NOR2 (N7229, N7226, N3719);
xor XOR2 (N7230, N7228, N205);
xor XOR2 (N7231, N7220, N3086);
nand NAND2 (N7232, N7224, N738);
not NOT1 (N7233, N7229);
nor NOR3 (N7234, N7232, N1420, N2192);
nor NOR2 (N7235, N7233, N5802);
xor XOR2 (N7236, N7227, N4554);
or OR3 (N7237, N7236, N5718, N5202);
nand NAND4 (N7238, N7212, N6281, N2667, N6206);
xor XOR2 (N7239, N7231, N6940);
buf BUF1 (N7240, N7235);
xor XOR2 (N7241, N7239, N5656);
or OR4 (N7242, N7234, N2733, N1654, N3533);
buf BUF1 (N7243, N7238);
nor NOR3 (N7244, N7243, N3563, N1998);
nor NOR2 (N7245, N7211, N4659);
not NOT1 (N7246, N7225);
buf BUF1 (N7247, N7241);
not NOT1 (N7248, N7247);
and AND3 (N7249, N7230, N2552, N6011);
or OR4 (N7250, N7223, N483, N4029, N2900);
not NOT1 (N7251, N7248);
buf BUF1 (N7252, N7245);
and AND4 (N7253, N7246, N542, N856, N2703);
buf BUF1 (N7254, N7252);
nand NAND3 (N7255, N7242, N1917, N6924);
not NOT1 (N7256, N7251);
xor XOR2 (N7257, N7256, N6760);
and AND4 (N7258, N7254, N6396, N2167, N5114);
buf BUF1 (N7259, N7257);
and AND4 (N7260, N7258, N498, N271, N4241);
not NOT1 (N7261, N7255);
and AND3 (N7262, N7240, N190, N2148);
xor XOR2 (N7263, N7261, N4706);
nand NAND4 (N7264, N7253, N6795, N5087, N341);
nand NAND2 (N7265, N7244, N3481);
and AND4 (N7266, N7262, N4210, N6709, N19);
xor XOR2 (N7267, N7217, N369);
buf BUF1 (N7268, N7267);
nor NOR4 (N7269, N7265, N1795, N3897, N7192);
or OR2 (N7270, N7263, N1757);
nand NAND4 (N7271, N7266, N3982, N6360, N2354);
nor NOR2 (N7272, N7270, N6544);
buf BUF1 (N7273, N7271);
buf BUF1 (N7274, N7272);
nand NAND3 (N7275, N7273, N4481, N6376);
xor XOR2 (N7276, N7249, N486);
or OR3 (N7277, N7276, N1906, N5340);
and AND4 (N7278, N7274, N6109, N3841, N4133);
nor NOR2 (N7279, N7277, N2275);
or OR4 (N7280, N7279, N3143, N5470, N5465);
not NOT1 (N7281, N7268);
or OR2 (N7282, N7280, N13);
nor NOR3 (N7283, N7237, N968, N5655);
and AND2 (N7284, N7282, N4274);
nor NOR4 (N7285, N7260, N2946, N4976, N4446);
buf BUF1 (N7286, N7284);
not NOT1 (N7287, N7275);
xor XOR2 (N7288, N7283, N2816);
not NOT1 (N7289, N7288);
nand NAND4 (N7290, N7250, N3265, N6320, N4194);
nand NAND3 (N7291, N7289, N3020, N7146);
buf BUF1 (N7292, N7278);
not NOT1 (N7293, N7285);
nor NOR4 (N7294, N7264, N4347, N7224, N3185);
not NOT1 (N7295, N7281);
nand NAND3 (N7296, N7269, N1594, N1997);
nand NAND4 (N7297, N7292, N5054, N591, N4694);
buf BUF1 (N7298, N7291);
nor NOR4 (N7299, N7294, N1172, N5193, N1615);
nor NOR3 (N7300, N7293, N747, N4807);
not NOT1 (N7301, N7286);
and AND4 (N7302, N7299, N4758, N6394, N5746);
not NOT1 (N7303, N7290);
not NOT1 (N7304, N7298);
and AND4 (N7305, N7296, N134, N3700, N56);
nand NAND3 (N7306, N7297, N2206, N360);
or OR2 (N7307, N7302, N2204);
buf BUF1 (N7308, N7300);
nand NAND3 (N7309, N7301, N2239, N5590);
or OR2 (N7310, N7304, N4738);
nor NOR4 (N7311, N7308, N5351, N3593, N4099);
nand NAND2 (N7312, N7307, N1108);
nor NOR4 (N7313, N7311, N1066, N2535, N6551);
buf BUF1 (N7314, N7306);
and AND2 (N7315, N7305, N6791);
or OR2 (N7316, N7312, N4623);
nor NOR2 (N7317, N7316, N1604);
nand NAND4 (N7318, N7315, N6468, N3309, N5282);
nor NOR4 (N7319, N7317, N2536, N4956, N2941);
not NOT1 (N7320, N7310);
not NOT1 (N7321, N7320);
not NOT1 (N7322, N7314);
not NOT1 (N7323, N7321);
nor NOR3 (N7324, N7322, N691, N6720);
or OR3 (N7325, N7295, N4888, N5821);
not NOT1 (N7326, N7309);
nor NOR2 (N7327, N7303, N1154);
or OR4 (N7328, N7327, N6305, N5704, N1160);
buf BUF1 (N7329, N7325);
xor XOR2 (N7330, N7319, N444);
xor XOR2 (N7331, N7313, N5431);
not NOT1 (N7332, N7318);
buf BUF1 (N7333, N7259);
xor XOR2 (N7334, N7332, N5482);
not NOT1 (N7335, N7331);
nor NOR2 (N7336, N7323, N1136);
buf BUF1 (N7337, N7326);
not NOT1 (N7338, N7336);
or OR4 (N7339, N7328, N4780, N3954, N3438);
nand NAND4 (N7340, N7337, N6002, N1095, N3948);
or OR3 (N7341, N7329, N3525, N638);
xor XOR2 (N7342, N7287, N1315);
xor XOR2 (N7343, N7342, N1264);
nand NAND4 (N7344, N7340, N3353, N3004, N1728);
buf BUF1 (N7345, N7333);
nor NOR4 (N7346, N7343, N2214, N3307, N7342);
and AND4 (N7347, N7330, N398, N2704, N5680);
nor NOR4 (N7348, N7346, N713, N4974, N7225);
or OR2 (N7349, N7348, N4901);
or OR3 (N7350, N7347, N1064, N4948);
buf BUF1 (N7351, N7324);
and AND4 (N7352, N7338, N6680, N5928, N3902);
not NOT1 (N7353, N7335);
nand NAND3 (N7354, N7339, N1160, N594);
and AND3 (N7355, N7344, N2709, N4562);
buf BUF1 (N7356, N7341);
or OR2 (N7357, N7350, N5627);
or OR3 (N7358, N7349, N5174, N4599);
nor NOR2 (N7359, N7354, N6283);
nor NOR2 (N7360, N7359, N5844);
nand NAND2 (N7361, N7352, N4039);
or OR2 (N7362, N7356, N2317);
and AND2 (N7363, N7362, N2949);
xor XOR2 (N7364, N7358, N5726);
buf BUF1 (N7365, N7353);
and AND4 (N7366, N7363, N5650, N660, N901);
nand NAND2 (N7367, N7334, N809);
not NOT1 (N7368, N7361);
xor XOR2 (N7369, N7360, N6834);
nand NAND2 (N7370, N7345, N7348);
nor NOR3 (N7371, N7369, N547, N3585);
or OR2 (N7372, N7367, N5645);
and AND3 (N7373, N7355, N2702, N1269);
nand NAND2 (N7374, N7366, N7201);
xor XOR2 (N7375, N7364, N2502);
buf BUF1 (N7376, N7357);
nor NOR3 (N7377, N7371, N3843, N6807);
not NOT1 (N7378, N7365);
nand NAND2 (N7379, N7370, N3280);
buf BUF1 (N7380, N7379);
buf BUF1 (N7381, N7380);
buf BUF1 (N7382, N7377);
nor NOR4 (N7383, N7376, N6596, N5700, N7013);
nand NAND4 (N7384, N7373, N5317, N6253, N2572);
not NOT1 (N7385, N7382);
nand NAND3 (N7386, N7375, N846, N4589);
xor XOR2 (N7387, N7386, N5618);
nand NAND2 (N7388, N7368, N3454);
not NOT1 (N7389, N7385);
or OR2 (N7390, N7383, N2792);
nand NAND4 (N7391, N7372, N3382, N4940, N963);
and AND2 (N7392, N7387, N5271);
xor XOR2 (N7393, N7384, N1497);
not NOT1 (N7394, N7389);
nor NOR3 (N7395, N7388, N5288, N737);
nor NOR2 (N7396, N7392, N1564);
nand NAND2 (N7397, N7390, N5990);
nand NAND2 (N7398, N7394, N952);
nor NOR4 (N7399, N7395, N2771, N298, N7316);
nor NOR4 (N7400, N7398, N6219, N3859, N2071);
buf BUF1 (N7401, N7391);
and AND2 (N7402, N7378, N5726);
and AND2 (N7403, N7401, N2081);
xor XOR2 (N7404, N7381, N2440);
or OR2 (N7405, N7399, N1262);
nand NAND2 (N7406, N7400, N5426);
or OR3 (N7407, N7402, N5845, N313);
xor XOR2 (N7408, N7374, N4819);
nand NAND2 (N7409, N7396, N2648);
or OR3 (N7410, N7408, N5265, N2609);
not NOT1 (N7411, N7406);
nor NOR3 (N7412, N7405, N3108, N2769);
xor XOR2 (N7413, N7410, N403);
not NOT1 (N7414, N7397);
nor NOR2 (N7415, N7411, N6265);
nand NAND3 (N7416, N7407, N6680, N678);
xor XOR2 (N7417, N7413, N1137);
and AND4 (N7418, N7351, N4675, N1110, N488);
nor NOR3 (N7419, N7403, N1347, N3514);
nand NAND4 (N7420, N7416, N912, N2800, N4224);
or OR3 (N7421, N7418, N1971, N6137);
nand NAND3 (N7422, N7415, N1277, N821);
not NOT1 (N7423, N7409);
xor XOR2 (N7424, N7404, N7399);
xor XOR2 (N7425, N7393, N4452);
and AND4 (N7426, N7419, N832, N5228, N1424);
nor NOR3 (N7427, N7425, N4615, N6104);
buf BUF1 (N7428, N7423);
and AND2 (N7429, N7427, N1103);
nand NAND3 (N7430, N7424, N111, N5366);
buf BUF1 (N7431, N7417);
xor XOR2 (N7432, N7431, N3888);
xor XOR2 (N7433, N7430, N3091);
or OR3 (N7434, N7420, N4635, N4205);
xor XOR2 (N7435, N7429, N6929);
and AND4 (N7436, N7412, N6462, N1190, N1271);
nor NOR4 (N7437, N7432, N1616, N766, N3444);
or OR2 (N7438, N7433, N4708);
nand NAND3 (N7439, N7437, N1953, N5531);
nand NAND3 (N7440, N7421, N3388, N4461);
nor NOR3 (N7441, N7414, N5112, N6087);
xor XOR2 (N7442, N7439, N7410);
xor XOR2 (N7443, N7441, N4163);
xor XOR2 (N7444, N7428, N4222);
or OR2 (N7445, N7444, N7342);
xor XOR2 (N7446, N7438, N5587);
nand NAND3 (N7447, N7434, N5519, N6049);
buf BUF1 (N7448, N7442);
not NOT1 (N7449, N7443);
nor NOR4 (N7450, N7446, N2549, N2334, N3569);
or OR3 (N7451, N7448, N3355, N5987);
xor XOR2 (N7452, N7447, N2308);
buf BUF1 (N7453, N7452);
nand NAND4 (N7454, N7450, N2787, N830, N3900);
xor XOR2 (N7455, N7453, N2272);
or OR4 (N7456, N7436, N4524, N2636, N4452);
not NOT1 (N7457, N7422);
nor NOR3 (N7458, N7426, N84, N6554);
not NOT1 (N7459, N7449);
xor XOR2 (N7460, N7455, N5489);
not NOT1 (N7461, N7435);
nand NAND2 (N7462, N7460, N3171);
or OR4 (N7463, N7445, N5385, N6799, N3114);
xor XOR2 (N7464, N7440, N4925);
not NOT1 (N7465, N7454);
buf BUF1 (N7466, N7463);
and AND2 (N7467, N7459, N7456);
and AND4 (N7468, N1348, N1341, N2774, N450);
and AND4 (N7469, N7464, N3665, N3252, N3586);
xor XOR2 (N7470, N7461, N6359);
buf BUF1 (N7471, N7457);
nand NAND4 (N7472, N7468, N342, N3477, N5014);
or OR2 (N7473, N7465, N7017);
nand NAND3 (N7474, N7467, N3693, N2896);
nand NAND2 (N7475, N7471, N4454);
and AND3 (N7476, N7474, N802, N5749);
and AND4 (N7477, N7475, N7250, N3542, N1658);
not NOT1 (N7478, N7451);
not NOT1 (N7479, N7466);
and AND2 (N7480, N7478, N4025);
nor NOR4 (N7481, N7476, N4626, N5513, N5281);
nor NOR2 (N7482, N7472, N2696);
xor XOR2 (N7483, N7473, N6200);
not NOT1 (N7484, N7479);
nor NOR2 (N7485, N7482, N942);
xor XOR2 (N7486, N7484, N2171);
buf BUF1 (N7487, N7470);
nor NOR4 (N7488, N7485, N7459, N333, N2203);
xor XOR2 (N7489, N7480, N4281);
nand NAND2 (N7490, N7487, N4906);
or OR4 (N7491, N7490, N412, N4646, N3022);
or OR4 (N7492, N7481, N1357, N4240, N4593);
nor NOR3 (N7493, N7469, N3560, N4479);
nand NAND3 (N7494, N7462, N5522, N2485);
not NOT1 (N7495, N7493);
and AND2 (N7496, N7483, N73);
and AND4 (N7497, N7486, N1882, N1817, N4422);
not NOT1 (N7498, N7489);
and AND4 (N7499, N7477, N4921, N6154, N271);
nor NOR2 (N7500, N7488, N928);
nand NAND4 (N7501, N7496, N6388, N1149, N1061);
nand NAND4 (N7502, N7499, N5429, N2042, N6329);
xor XOR2 (N7503, N7498, N1366);
or OR3 (N7504, N7494, N1913, N6472);
or OR4 (N7505, N7501, N1122, N90, N3485);
or OR2 (N7506, N7495, N5771);
or OR2 (N7507, N7458, N1588);
and AND3 (N7508, N7497, N6557, N6377);
nor NOR4 (N7509, N7504, N4933, N4704, N1406);
nand NAND2 (N7510, N7500, N357);
buf BUF1 (N7511, N7507);
or OR4 (N7512, N7508, N883, N3916, N1266);
not NOT1 (N7513, N7503);
and AND4 (N7514, N7492, N5537, N3925, N5694);
nand NAND4 (N7515, N7509, N3275, N7249, N7306);
xor XOR2 (N7516, N7513, N198);
or OR4 (N7517, N7511, N2736, N7158, N5772);
not NOT1 (N7518, N7505);
nor NOR4 (N7519, N7506, N2269, N1102, N5714);
nor NOR2 (N7520, N7491, N1624);
buf BUF1 (N7521, N7514);
and AND2 (N7522, N7518, N4204);
and AND2 (N7523, N7510, N2456);
xor XOR2 (N7524, N7502, N2333);
and AND3 (N7525, N7516, N4128, N2282);
not NOT1 (N7526, N7517);
nor NOR4 (N7527, N7523, N2231, N985, N4419);
buf BUF1 (N7528, N7515);
buf BUF1 (N7529, N7512);
nand NAND2 (N7530, N7524, N6037);
nand NAND3 (N7531, N7519, N1082, N3082);
and AND2 (N7532, N7526, N3640);
xor XOR2 (N7533, N7525, N6341);
xor XOR2 (N7534, N7522, N6120);
buf BUF1 (N7535, N7533);
xor XOR2 (N7536, N7530, N3740);
not NOT1 (N7537, N7528);
nand NAND3 (N7538, N7532, N6437, N677);
nor NOR2 (N7539, N7537, N3762);
not NOT1 (N7540, N7539);
not NOT1 (N7541, N7538);
xor XOR2 (N7542, N7535, N1718);
or OR3 (N7543, N7542, N6136, N2864);
not NOT1 (N7544, N7536);
xor XOR2 (N7545, N7541, N3774);
nand NAND4 (N7546, N7521, N108, N3628, N6144);
nand NAND3 (N7547, N7543, N3115, N5017);
xor XOR2 (N7548, N7545, N5733);
and AND2 (N7549, N7547, N3629);
or OR3 (N7550, N7527, N6672, N6608);
xor XOR2 (N7551, N7546, N3076);
or OR3 (N7552, N7550, N5497, N6532);
buf BUF1 (N7553, N7544);
nor NOR2 (N7554, N7529, N4775);
not NOT1 (N7555, N7554);
xor XOR2 (N7556, N7549, N3311);
and AND3 (N7557, N7552, N7273, N3435);
and AND4 (N7558, N7555, N2285, N775, N1011);
buf BUF1 (N7559, N7556);
not NOT1 (N7560, N7531);
not NOT1 (N7561, N7540);
buf BUF1 (N7562, N7559);
nand NAND4 (N7563, N7558, N2156, N3211, N1776);
or OR3 (N7564, N7563, N5864, N5802);
nor NOR3 (N7565, N7520, N3864, N6292);
not NOT1 (N7566, N7557);
buf BUF1 (N7567, N7548);
not NOT1 (N7568, N7566);
nand NAND2 (N7569, N7551, N6679);
not NOT1 (N7570, N7564);
buf BUF1 (N7571, N7562);
and AND3 (N7572, N7553, N218, N2236);
and AND2 (N7573, N7570, N5091);
nand NAND2 (N7574, N7572, N4369);
and AND4 (N7575, N7569, N6613, N6966, N1928);
nor NOR4 (N7576, N7575, N877, N2134, N3464);
xor XOR2 (N7577, N7567, N6153);
buf BUF1 (N7578, N7571);
not NOT1 (N7579, N7568);
nand NAND4 (N7580, N7577, N2, N5860, N5337);
nand NAND3 (N7581, N7534, N1717, N7374);
buf BUF1 (N7582, N7573);
buf BUF1 (N7583, N7581);
nand NAND2 (N7584, N7583, N4584);
xor XOR2 (N7585, N7579, N5304);
or OR3 (N7586, N7584, N5633, N2483);
xor XOR2 (N7587, N7565, N6567);
buf BUF1 (N7588, N7582);
buf BUF1 (N7589, N7576);
or OR4 (N7590, N7589, N2321, N314, N2232);
buf BUF1 (N7591, N7561);
or OR3 (N7592, N7586, N2505, N3934);
xor XOR2 (N7593, N7590, N5915);
nor NOR2 (N7594, N7580, N6116);
not NOT1 (N7595, N7593);
nand NAND4 (N7596, N7592, N2778, N954, N7313);
nand NAND2 (N7597, N7585, N5702);
xor XOR2 (N7598, N7574, N1111);
not NOT1 (N7599, N7578);
nand NAND3 (N7600, N7591, N2820, N5090);
not NOT1 (N7601, N7560);
nand NAND2 (N7602, N7588, N7426);
buf BUF1 (N7603, N7596);
and AND4 (N7604, N7603, N6040, N1466, N7536);
not NOT1 (N7605, N7587);
nand NAND4 (N7606, N7598, N457, N2362, N7604);
nor NOR4 (N7607, N1740, N6348, N2292, N1588);
buf BUF1 (N7608, N7602);
nand NAND2 (N7609, N7605, N1858);
not NOT1 (N7610, N7608);
buf BUF1 (N7611, N7597);
xor XOR2 (N7612, N7609, N4234);
nor NOR3 (N7613, N7610, N497, N1622);
not NOT1 (N7614, N7599);
or OR3 (N7615, N7594, N6891, N3603);
not NOT1 (N7616, N7600);
not NOT1 (N7617, N7615);
buf BUF1 (N7618, N7614);
xor XOR2 (N7619, N7618, N5005);
not NOT1 (N7620, N7616);
nor NOR2 (N7621, N7595, N2057);
or OR4 (N7622, N7606, N6153, N4475, N3091);
and AND4 (N7623, N7620, N3959, N4323, N4184);
xor XOR2 (N7624, N7611, N4975);
nand NAND3 (N7625, N7607, N1496, N4834);
or OR2 (N7626, N7619, N545);
or OR4 (N7627, N7601, N6213, N4634, N4662);
buf BUF1 (N7628, N7613);
buf BUF1 (N7629, N7621);
and AND3 (N7630, N7627, N2886, N2843);
nor NOR3 (N7631, N7629, N3421, N4041);
or OR4 (N7632, N7628, N4349, N6799, N7325);
xor XOR2 (N7633, N7617, N2905);
buf BUF1 (N7634, N7623);
buf BUF1 (N7635, N7633);
and AND4 (N7636, N7624, N4535, N6669, N6454);
not NOT1 (N7637, N7625);
and AND3 (N7638, N7626, N6233, N3571);
not NOT1 (N7639, N7637);
nand NAND2 (N7640, N7639, N2858);
buf BUF1 (N7641, N7630);
buf BUF1 (N7642, N7632);
or OR3 (N7643, N7640, N4369, N6299);
or OR3 (N7644, N7643, N7614, N4260);
nor NOR2 (N7645, N7612, N487);
or OR4 (N7646, N7645, N7263, N4945, N4042);
nand NAND2 (N7647, N7638, N634);
nand NAND4 (N7648, N7631, N2494, N1396, N4891);
nor NOR2 (N7649, N7634, N3522);
nor NOR4 (N7650, N7644, N244, N3367, N1373);
buf BUF1 (N7651, N7649);
nor NOR3 (N7652, N7641, N2405, N640);
not NOT1 (N7653, N7635);
buf BUF1 (N7654, N7651);
nand NAND2 (N7655, N7622, N6054);
buf BUF1 (N7656, N7652);
nand NAND2 (N7657, N7653, N7593);
or OR2 (N7658, N7655, N5788);
not NOT1 (N7659, N7657);
and AND2 (N7660, N7646, N1657);
and AND2 (N7661, N7642, N2561);
nor NOR4 (N7662, N7647, N6837, N2144, N4682);
or OR4 (N7663, N7658, N4014, N2158, N1860);
xor XOR2 (N7664, N7654, N5512);
or OR3 (N7665, N7664, N3868, N395);
or OR2 (N7666, N7662, N4323);
nand NAND2 (N7667, N7656, N4621);
xor XOR2 (N7668, N7648, N2621);
not NOT1 (N7669, N7660);
buf BUF1 (N7670, N7668);
nor NOR2 (N7671, N7665, N1618);
buf BUF1 (N7672, N7650);
or OR4 (N7673, N7666, N6802, N3125, N2743);
and AND4 (N7674, N7667, N6583, N6774, N4412);
nand NAND4 (N7675, N7661, N4631, N2164, N5821);
nand NAND3 (N7676, N7663, N6175, N2237);
xor XOR2 (N7677, N7636, N2550);
nand NAND2 (N7678, N7670, N4740);
and AND3 (N7679, N7674, N3209, N4492);
xor XOR2 (N7680, N7676, N2187);
buf BUF1 (N7681, N7672);
or OR2 (N7682, N7671, N626);
or OR2 (N7683, N7673, N1056);
or OR2 (N7684, N7682, N334);
nor NOR4 (N7685, N7684, N3238, N6179, N5833);
buf BUF1 (N7686, N7681);
nand NAND4 (N7687, N7683, N1374, N6195, N6611);
buf BUF1 (N7688, N7680);
not NOT1 (N7689, N7659);
buf BUF1 (N7690, N7686);
nand NAND4 (N7691, N7688, N3651, N180, N7488);
and AND2 (N7692, N7691, N5697);
nand NAND2 (N7693, N7677, N3407);
and AND4 (N7694, N7675, N170, N4931, N2255);
or OR4 (N7695, N7693, N6439, N3033, N3536);
nand NAND4 (N7696, N7694, N2256, N3202, N2902);
and AND2 (N7697, N7669, N4062);
nor NOR3 (N7698, N7689, N963, N4011);
not NOT1 (N7699, N7679);
buf BUF1 (N7700, N7698);
xor XOR2 (N7701, N7699, N1960);
and AND4 (N7702, N7692, N3860, N6117, N6796);
or OR3 (N7703, N7685, N970, N4130);
buf BUF1 (N7704, N7703);
nor NOR4 (N7705, N7678, N5466, N6074, N5273);
nor NOR4 (N7706, N7702, N933, N6873, N2674);
nor NOR3 (N7707, N7696, N1736, N7495);
and AND3 (N7708, N7690, N1485, N502);
nand NAND2 (N7709, N7706, N1);
xor XOR2 (N7710, N7687, N5699);
buf BUF1 (N7711, N7704);
buf BUF1 (N7712, N7708);
not NOT1 (N7713, N7695);
nor NOR4 (N7714, N7705, N2717, N1961, N2156);
and AND3 (N7715, N7710, N5066, N1056);
nand NAND2 (N7716, N7713, N3768);
buf BUF1 (N7717, N7712);
nor NOR4 (N7718, N7715, N5312, N2851, N6618);
nand NAND4 (N7719, N7718, N1741, N4146, N2466);
xor XOR2 (N7720, N7714, N727);
buf BUF1 (N7721, N7717);
not NOT1 (N7722, N7719);
nand NAND4 (N7723, N7701, N7361, N6724, N4429);
not NOT1 (N7724, N7720);
or OR2 (N7725, N7723, N1640);
or OR2 (N7726, N7725, N175);
and AND4 (N7727, N7709, N2737, N1560, N2901);
not NOT1 (N7728, N7727);
and AND3 (N7729, N7722, N2773, N7061);
not NOT1 (N7730, N7700);
not NOT1 (N7731, N7707);
buf BUF1 (N7732, N7729);
nor NOR2 (N7733, N7726, N6281);
buf BUF1 (N7734, N7721);
not NOT1 (N7735, N7728);
or OR4 (N7736, N7735, N921, N3619, N401);
nand NAND2 (N7737, N7724, N933);
nor NOR4 (N7738, N7711, N60, N7649, N124);
and AND4 (N7739, N7697, N2041, N4336, N2901);
buf BUF1 (N7740, N7732);
and AND2 (N7741, N7739, N5648);
xor XOR2 (N7742, N7737, N1637);
nor NOR2 (N7743, N7738, N5409);
and AND4 (N7744, N7743, N1754, N4447, N341);
or OR3 (N7745, N7733, N6694, N186);
buf BUF1 (N7746, N7744);
and AND3 (N7747, N7736, N7650, N7135);
or OR2 (N7748, N7731, N367);
nor NOR4 (N7749, N7742, N3791, N3917, N1129);
not NOT1 (N7750, N7741);
buf BUF1 (N7751, N7730);
nor NOR4 (N7752, N7748, N776, N7092, N1277);
or OR4 (N7753, N7734, N3903, N3036, N4045);
or OR4 (N7754, N7752, N3390, N7247, N3001);
nor NOR3 (N7755, N7746, N4677, N5432);
nand NAND4 (N7756, N7740, N7501, N2997, N2236);
nand NAND3 (N7757, N7716, N6060, N6684);
nand NAND3 (N7758, N7749, N3888, N5043);
nand NAND4 (N7759, N7753, N2915, N4076, N5892);
nor NOR3 (N7760, N7756, N3286, N3124);
buf BUF1 (N7761, N7754);
and AND2 (N7762, N7747, N5024);
not NOT1 (N7763, N7759);
buf BUF1 (N7764, N7762);
nand NAND2 (N7765, N7763, N6980);
or OR4 (N7766, N7751, N6069, N4292, N3185);
and AND2 (N7767, N7755, N5223);
or OR2 (N7768, N7758, N4320);
buf BUF1 (N7769, N7750);
and AND2 (N7770, N7769, N5276);
xor XOR2 (N7771, N7765, N3585);
buf BUF1 (N7772, N7767);
not NOT1 (N7773, N7761);
nand NAND3 (N7774, N7773, N4800, N5561);
not NOT1 (N7775, N7771);
nand NAND4 (N7776, N7764, N1774, N3265, N4351);
and AND2 (N7777, N7757, N895);
nand NAND4 (N7778, N7745, N1135, N4434, N3321);
and AND3 (N7779, N7776, N3062, N6645);
or OR3 (N7780, N7777, N3649, N7298);
nor NOR4 (N7781, N7772, N2432, N7725, N603);
or OR3 (N7782, N7768, N6256, N5022);
nand NAND2 (N7783, N7782, N2727);
nor NOR2 (N7784, N7770, N3390);
nand NAND2 (N7785, N7760, N4566);
not NOT1 (N7786, N7779);
nor NOR2 (N7787, N7780, N5382);
or OR4 (N7788, N7784, N3879, N6301, N1734);
xor XOR2 (N7789, N7775, N421);
or OR3 (N7790, N7783, N2377, N702);
and AND2 (N7791, N7766, N3886);
not NOT1 (N7792, N7791);
xor XOR2 (N7793, N7781, N4347);
or OR4 (N7794, N7778, N6720, N2143, N6912);
xor XOR2 (N7795, N7788, N5476);
nor NOR4 (N7796, N7795, N3974, N6650, N6275);
xor XOR2 (N7797, N7789, N797);
and AND3 (N7798, N7790, N2067, N2199);
or OR4 (N7799, N7786, N2431, N3278, N4974);
buf BUF1 (N7800, N7792);
or OR4 (N7801, N7787, N6182, N995, N3778);
nand NAND2 (N7802, N7785, N2830);
not NOT1 (N7803, N7793);
not NOT1 (N7804, N7794);
and AND4 (N7805, N7801, N4981, N7145, N4000);
nor NOR2 (N7806, N7799, N2855);
nand NAND2 (N7807, N7774, N1246);
or OR3 (N7808, N7802, N6960, N2633);
nand NAND4 (N7809, N7796, N2291, N402, N1419);
and AND2 (N7810, N7807, N6015);
nor NOR3 (N7811, N7798, N3266, N2003);
or OR3 (N7812, N7808, N3032, N4597);
not NOT1 (N7813, N7806);
buf BUF1 (N7814, N7809);
nand NAND4 (N7815, N7813, N779, N3099, N4929);
not NOT1 (N7816, N7810);
not NOT1 (N7817, N7804);
nor NOR4 (N7818, N7817, N7615, N648, N392);
not NOT1 (N7819, N7811);
nand NAND2 (N7820, N7805, N1511);
nand NAND4 (N7821, N7812, N3139, N6623, N6068);
nor NOR2 (N7822, N7819, N5519);
not NOT1 (N7823, N7800);
nand NAND2 (N7824, N7821, N664);
nand NAND3 (N7825, N7797, N2447, N875);
xor XOR2 (N7826, N7824, N7326);
and AND3 (N7827, N7818, N6138, N3037);
xor XOR2 (N7828, N7825, N5977);
or OR4 (N7829, N7820, N5753, N986, N570);
nand NAND3 (N7830, N7816, N1502, N7390);
buf BUF1 (N7831, N7827);
or OR2 (N7832, N7828, N6360);
and AND4 (N7833, N7826, N7527, N6967, N187);
buf BUF1 (N7834, N7829);
or OR4 (N7835, N7831, N1668, N7521, N7155);
buf BUF1 (N7836, N7830);
and AND3 (N7837, N7803, N5475, N2319);
not NOT1 (N7838, N7814);
or OR3 (N7839, N7822, N5565, N2592);
not NOT1 (N7840, N7834);
or OR4 (N7841, N7836, N1368, N6256, N4097);
nand NAND2 (N7842, N7839, N1810);
xor XOR2 (N7843, N7841, N7150);
and AND4 (N7844, N7838, N5686, N5601, N22);
nor NOR2 (N7845, N7835, N807);
and AND4 (N7846, N7833, N1016, N2795, N3857);
nand NAND3 (N7847, N7846, N3293, N206);
and AND3 (N7848, N7842, N2400, N2061);
not NOT1 (N7849, N7847);
xor XOR2 (N7850, N7845, N7173);
xor XOR2 (N7851, N7823, N871);
buf BUF1 (N7852, N7837);
xor XOR2 (N7853, N7840, N845);
or OR2 (N7854, N7852, N3403);
nand NAND3 (N7855, N7832, N6668, N1399);
nor NOR4 (N7856, N7844, N5276, N429, N4312);
buf BUF1 (N7857, N7815);
and AND2 (N7858, N7848, N4891);
not NOT1 (N7859, N7843);
xor XOR2 (N7860, N7854, N6696);
nor NOR4 (N7861, N7859, N2611, N3831, N3301);
and AND4 (N7862, N7856, N4837, N447, N4476);
nand NAND2 (N7863, N7861, N7591);
and AND4 (N7864, N7858, N4166, N7792, N6863);
xor XOR2 (N7865, N7855, N2219);
xor XOR2 (N7866, N7860, N5748);
nand NAND3 (N7867, N7853, N7587, N6387);
nor NOR2 (N7868, N7864, N2301);
nor NOR2 (N7869, N7849, N1293);
buf BUF1 (N7870, N7857);
buf BUF1 (N7871, N7865);
xor XOR2 (N7872, N7866, N5338);
not NOT1 (N7873, N7867);
buf BUF1 (N7874, N7870);
or OR3 (N7875, N7850, N7704, N5034);
xor XOR2 (N7876, N7851, N5816);
xor XOR2 (N7877, N7875, N5870);
and AND2 (N7878, N7869, N3018);
and AND2 (N7879, N7876, N2802);
buf BUF1 (N7880, N7868);
nand NAND4 (N7881, N7880, N6876, N5941, N2187);
buf BUF1 (N7882, N7877);
nand NAND3 (N7883, N7872, N6989, N4316);
or OR2 (N7884, N7871, N4004);
xor XOR2 (N7885, N7884, N3930);
not NOT1 (N7886, N7881);
nor NOR2 (N7887, N7874, N3816);
buf BUF1 (N7888, N7863);
nor NOR2 (N7889, N7887, N2930);
not NOT1 (N7890, N7862);
or OR2 (N7891, N7886, N2881);
nand NAND4 (N7892, N7888, N5324, N7718, N326);
or OR3 (N7893, N7878, N6279, N1135);
or OR4 (N7894, N7892, N6283, N4728, N2827);
nor NOR4 (N7895, N7873, N6983, N5734, N440);
nor NOR3 (N7896, N7879, N5511, N7805);
nor NOR4 (N7897, N7883, N6513, N2277, N5171);
not NOT1 (N7898, N7890);
nand NAND4 (N7899, N7897, N5806, N1317, N3878);
nor NOR3 (N7900, N7889, N3174, N6738);
xor XOR2 (N7901, N7898, N874);
xor XOR2 (N7902, N7895, N4370);
buf BUF1 (N7903, N7896);
or OR2 (N7904, N7893, N7631);
xor XOR2 (N7905, N7900, N744);
xor XOR2 (N7906, N7894, N5050);
not NOT1 (N7907, N7891);
buf BUF1 (N7908, N7904);
buf BUF1 (N7909, N7908);
nand NAND3 (N7910, N7882, N7061, N2893);
not NOT1 (N7911, N7903);
buf BUF1 (N7912, N7911);
nand NAND3 (N7913, N7885, N1341, N2085);
nand NAND4 (N7914, N7901, N666, N2768, N7514);
not NOT1 (N7915, N7906);
buf BUF1 (N7916, N7915);
not NOT1 (N7917, N7914);
xor XOR2 (N7918, N7917, N2956);
nand NAND2 (N7919, N7909, N4512);
not NOT1 (N7920, N7910);
or OR3 (N7921, N7902, N1791, N4915);
or OR4 (N7922, N7905, N6758, N7806, N606);
buf BUF1 (N7923, N7913);
or OR2 (N7924, N7916, N6655);
or OR4 (N7925, N7923, N1414, N2459, N5421);
nand NAND2 (N7926, N7922, N3059);
nor NOR4 (N7927, N7920, N7407, N1824, N43);
not NOT1 (N7928, N7927);
nand NAND3 (N7929, N7925, N2181, N3625);
xor XOR2 (N7930, N7928, N3156);
or OR3 (N7931, N7899, N6770, N4972);
not NOT1 (N7932, N7919);
or OR4 (N7933, N7932, N7155, N4861, N3405);
buf BUF1 (N7934, N7931);
nor NOR2 (N7935, N7912, N5682);
and AND3 (N7936, N7933, N4, N10);
xor XOR2 (N7937, N7918, N1546);
and AND2 (N7938, N7921, N3715);
buf BUF1 (N7939, N7937);
xor XOR2 (N7940, N7907, N2840);
or OR3 (N7941, N7929, N1053, N3044);
or OR2 (N7942, N7934, N220);
not NOT1 (N7943, N7940);
or OR4 (N7944, N7943, N3804, N1499, N4058);
not NOT1 (N7945, N7939);
or OR2 (N7946, N7936, N1006);
nand NAND2 (N7947, N7938, N4880);
and AND4 (N7948, N7942, N1284, N5873, N3600);
and AND2 (N7949, N7930, N4894);
or OR3 (N7950, N7924, N4237, N4102);
not NOT1 (N7951, N7946);
not NOT1 (N7952, N7945);
nor NOR4 (N7953, N7947, N7554, N3335, N5618);
not NOT1 (N7954, N7950);
xor XOR2 (N7955, N7949, N7309);
nand NAND4 (N7956, N7935, N7083, N1488, N4485);
nand NAND2 (N7957, N7954, N6727);
buf BUF1 (N7958, N7955);
not NOT1 (N7959, N7953);
or OR4 (N7960, N7958, N1375, N461, N3520);
nand NAND4 (N7961, N7926, N3651, N4856, N4976);
nand NAND4 (N7962, N7948, N3429, N6919, N1498);
nand NAND3 (N7963, N7956, N4664, N7462);
not NOT1 (N7964, N7957);
nand NAND2 (N7965, N7951, N155);
or OR4 (N7966, N7960, N3264, N5900, N1456);
or OR2 (N7967, N7963, N6818);
or OR4 (N7968, N7962, N7457, N2060, N3709);
nand NAND3 (N7969, N7967, N946, N1242);
buf BUF1 (N7970, N7944);
not NOT1 (N7971, N7952);
buf BUF1 (N7972, N7941);
and AND4 (N7973, N7968, N2696, N5683, N2884);
or OR3 (N7974, N7971, N5490, N3238);
and AND2 (N7975, N7961, N1547);
xor XOR2 (N7976, N7959, N2069);
xor XOR2 (N7977, N7975, N4271);
not NOT1 (N7978, N7965);
nand NAND3 (N7979, N7973, N1595, N3017);
buf BUF1 (N7980, N7964);
nor NOR3 (N7981, N7978, N3414, N7779);
buf BUF1 (N7982, N7970);
buf BUF1 (N7983, N7981);
buf BUF1 (N7984, N7976);
nand NAND2 (N7985, N7984, N1744);
nor NOR4 (N7986, N7972, N4454, N3688, N838);
xor XOR2 (N7987, N7979, N2759);
nand NAND2 (N7988, N7985, N5232);
nor NOR3 (N7989, N7982, N5845, N1696);
buf BUF1 (N7990, N7977);
nand NAND3 (N7991, N7980, N526, N7124);
nand NAND2 (N7992, N7989, N354);
buf BUF1 (N7993, N7991);
not NOT1 (N7994, N7974);
buf BUF1 (N7995, N7986);
or OR4 (N7996, N7987, N1299, N5493, N2188);
buf BUF1 (N7997, N7983);
buf BUF1 (N7998, N7995);
nand NAND3 (N7999, N7994, N1744, N511);
nand NAND4 (N8000, N7992, N3291, N931, N6249);
nor NOR3 (N8001, N7988, N7979, N4694);
xor XOR2 (N8002, N7996, N6267);
and AND2 (N8003, N8001, N5997);
buf BUF1 (N8004, N7990);
nand NAND3 (N8005, N8000, N4659, N3049);
not NOT1 (N8006, N8004);
and AND4 (N8007, N7997, N5000, N4929, N3679);
nand NAND4 (N8008, N8006, N811, N1488, N6586);
nor NOR2 (N8009, N7966, N5199);
xor XOR2 (N8010, N7969, N1299);
buf BUF1 (N8011, N7998);
nand NAND4 (N8012, N8010, N2652, N4256, N6052);
xor XOR2 (N8013, N7999, N2135);
and AND4 (N8014, N8007, N3000, N2149, N4103);
xor XOR2 (N8015, N8002, N905);
buf BUF1 (N8016, N8012);
endmodule