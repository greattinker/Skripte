// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N209,N213,N203,N184,N212,N200,N206,N187,N211,N214;

nand NAND4 (N15, N2, N5, N8, N7);
buf BUF1 (N16, N2);
nand NAND2 (N17, N7, N2);
and AND4 (N18, N12, N3, N8, N1);
xor XOR2 (N19, N1, N16);
buf BUF1 (N20, N3);
buf BUF1 (N21, N11);
not NOT1 (N22, N9);
and AND2 (N23, N14, N3);
not NOT1 (N24, N17);
and AND4 (N25, N8, N4, N17, N3);
buf BUF1 (N26, N5);
nor NOR3 (N27, N15, N19, N12);
buf BUF1 (N28, N20);
xor XOR2 (N29, N4, N21);
not NOT1 (N30, N15);
nor NOR4 (N31, N24, N27, N7, N27);
or OR2 (N32, N11, N27);
nand NAND3 (N33, N29, N6, N18);
buf BUF1 (N34, N17);
nor NOR4 (N35, N31, N20, N10, N20);
not NOT1 (N36, N32);
nor NOR2 (N37, N33, N11);
nor NOR3 (N38, N37, N8, N32);
not NOT1 (N39, N28);
xor XOR2 (N40, N30, N30);
xor XOR2 (N41, N35, N40);
buf BUF1 (N42, N21);
and AND2 (N43, N22, N34);
or OR2 (N44, N28, N9);
buf BUF1 (N45, N23);
nor NOR3 (N46, N43, N44, N35);
and AND3 (N47, N9, N38, N33);
buf BUF1 (N48, N26);
not NOT1 (N49, N46);
not NOT1 (N50, N14);
and AND4 (N51, N45, N35, N47, N31);
nand NAND4 (N52, N16, N51, N26, N41);
xor XOR2 (N53, N12, N3);
not NOT1 (N54, N14);
and AND4 (N55, N53, N46, N12, N31);
nor NOR3 (N56, N52, N32, N41);
nor NOR2 (N57, N49, N23);
and AND3 (N58, N39, N57, N18);
or OR2 (N59, N31, N13);
nor NOR3 (N60, N48, N33, N20);
or OR3 (N61, N42, N42, N47);
xor XOR2 (N62, N59, N18);
nand NAND3 (N63, N60, N3, N19);
and AND4 (N64, N56, N46, N37, N61);
and AND3 (N65, N60, N48, N40);
nor NOR3 (N66, N64, N3, N53);
xor XOR2 (N67, N66, N57);
nand NAND2 (N68, N65, N10);
buf BUF1 (N69, N58);
nor NOR4 (N70, N63, N3, N22, N33);
not NOT1 (N71, N36);
nand NAND2 (N72, N68, N17);
and AND4 (N73, N62, N61, N6, N33);
or OR4 (N74, N25, N52, N21, N70);
not NOT1 (N75, N14);
and AND3 (N76, N73, N39, N6);
or OR2 (N77, N50, N9);
nand NAND2 (N78, N75, N22);
xor XOR2 (N79, N69, N5);
buf BUF1 (N80, N77);
not NOT1 (N81, N78);
and AND4 (N82, N54, N10, N38, N4);
and AND4 (N83, N76, N77, N19, N40);
buf BUF1 (N84, N79);
and AND4 (N85, N84, N20, N40, N44);
not NOT1 (N86, N71);
xor XOR2 (N87, N67, N80);
nand NAND4 (N88, N22, N72, N59, N53);
not NOT1 (N89, N23);
buf BUF1 (N90, N87);
xor XOR2 (N91, N86, N38);
not NOT1 (N92, N55);
or OR2 (N93, N81, N42);
xor XOR2 (N94, N85, N31);
or OR2 (N95, N89, N48);
not NOT1 (N96, N95);
and AND2 (N97, N94, N65);
nand NAND3 (N98, N83, N92, N55);
nor NOR2 (N99, N30, N75);
not NOT1 (N100, N90);
nand NAND4 (N101, N100, N6, N89, N84);
or OR3 (N102, N101, N96, N3);
buf BUF1 (N103, N9);
buf BUF1 (N104, N93);
nor NOR3 (N105, N74, N13, N53);
and AND4 (N106, N88, N38, N70, N104);
and AND2 (N107, N47, N43);
nor NOR2 (N108, N97, N10);
nor NOR2 (N109, N103, N53);
and AND2 (N110, N105, N13);
and AND2 (N111, N82, N7);
xor XOR2 (N112, N109, N22);
nor NOR4 (N113, N99, N101, N50, N60);
nand NAND3 (N114, N110, N110, N91);
not NOT1 (N115, N49);
and AND3 (N116, N102, N35, N58);
and AND2 (N117, N108, N74);
xor XOR2 (N118, N107, N91);
nor NOR4 (N119, N115, N45, N106, N32);
nand NAND3 (N120, N91, N36, N85);
nand NAND4 (N121, N119, N92, N106, N78);
buf BUF1 (N122, N112);
buf BUF1 (N123, N98);
buf BUF1 (N124, N117);
or OR2 (N125, N114, N7);
nor NOR3 (N126, N125, N19, N49);
or OR4 (N127, N113, N104, N98, N13);
buf BUF1 (N128, N121);
buf BUF1 (N129, N116);
buf BUF1 (N130, N126);
not NOT1 (N131, N128);
not NOT1 (N132, N127);
nand NAND3 (N133, N124, N63, N80);
nand NAND4 (N134, N120, N114, N15, N38);
not NOT1 (N135, N129);
not NOT1 (N136, N135);
or OR2 (N137, N123, N59);
nand NAND2 (N138, N131, N12);
nand NAND4 (N139, N136, N100, N133, N22);
xor XOR2 (N140, N132, N25);
nor NOR3 (N141, N91, N140, N103);
not NOT1 (N142, N77);
and AND2 (N143, N122, N85);
nor NOR4 (N144, N134, N97, N17, N68);
nand NAND4 (N145, N139, N136, N30, N2);
nand NAND2 (N146, N145, N35);
nor NOR2 (N147, N141, N89);
or OR4 (N148, N138, N3, N34, N64);
xor XOR2 (N149, N137, N93);
buf BUF1 (N150, N146);
and AND3 (N151, N149, N85, N107);
not NOT1 (N152, N111);
nor NOR3 (N153, N150, N71, N17);
xor XOR2 (N154, N143, N3);
xor XOR2 (N155, N153, N68);
or OR3 (N156, N151, N52, N17);
xor XOR2 (N157, N148, N35);
not NOT1 (N158, N147);
nand NAND2 (N159, N142, N157);
not NOT1 (N160, N84);
or OR3 (N161, N154, N85, N86);
not NOT1 (N162, N155);
buf BUF1 (N163, N158);
nor NOR4 (N164, N161, N56, N48, N99);
and AND4 (N165, N144, N52, N155, N109);
and AND3 (N166, N164, N52, N63);
not NOT1 (N167, N165);
and AND2 (N168, N167, N114);
nor NOR4 (N169, N159, N67, N1, N128);
nand NAND4 (N170, N169, N98, N49, N99);
and AND3 (N171, N160, N97, N147);
nand NAND4 (N172, N163, N77, N61, N90);
nand NAND4 (N173, N156, N110, N134, N49);
xor XOR2 (N174, N170, N95);
xor XOR2 (N175, N130, N45);
buf BUF1 (N176, N168);
buf BUF1 (N177, N175);
buf BUF1 (N178, N152);
buf BUF1 (N179, N177);
or OR2 (N180, N166, N64);
not NOT1 (N181, N171);
nor NOR3 (N182, N178, N43, N53);
and AND2 (N183, N162, N172);
xor XOR2 (N184, N95, N92);
not NOT1 (N185, N179);
nor NOR2 (N186, N176, N30);
xor XOR2 (N187, N186, N35);
nor NOR4 (N188, N118, N71, N175, N137);
nand NAND4 (N189, N188, N147, N27, N57);
or OR2 (N190, N185, N112);
not NOT1 (N191, N173);
not NOT1 (N192, N174);
xor XOR2 (N193, N189, N182);
nand NAND3 (N194, N51, N176, N153);
and AND2 (N195, N192, N46);
nor NOR3 (N196, N194, N80, N3);
nor NOR4 (N197, N183, N139, N189, N115);
and AND2 (N198, N191, N31);
buf BUF1 (N199, N196);
buf BUF1 (N200, N181);
xor XOR2 (N201, N190, N90);
and AND3 (N202, N195, N57, N32);
or OR2 (N203, N193, N199);
not NOT1 (N204, N44);
nand NAND2 (N205, N202, N16);
nor NOR2 (N206, N198, N193);
and AND3 (N207, N197, N113, N158);
not NOT1 (N208, N201);
nand NAND3 (N209, N207, N121, N2);
buf BUF1 (N210, N180);
buf BUF1 (N211, N204);
buf BUF1 (N212, N210);
and AND4 (N213, N208, N47, N83, N114);
not NOT1 (N214, N205);
endmodule