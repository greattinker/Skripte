// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N15971,N16004,N15997,N16008,N16009,N15987,N16007,N15999,N16003,N16010;

nor NOR2 (N11, N5, N5);
buf BUF1 (N12, N3);
buf BUF1 (N13, N7);
nand NAND4 (N14, N8, N9, N13, N12);
xor XOR2 (N15, N6, N14);
nor NOR4 (N16, N8, N9, N9, N10);
buf BUF1 (N17, N2);
xor XOR2 (N18, N9, N9);
nor NOR4 (N19, N11, N17, N16, N8);
buf BUF1 (N20, N10);
xor XOR2 (N21, N14, N1);
nor NOR3 (N22, N11, N17, N11);
buf BUF1 (N23, N5);
buf BUF1 (N24, N10);
nand NAND3 (N25, N9, N22, N23);
or OR4 (N26, N17, N14, N18, N22);
nor NOR3 (N27, N14, N11, N25);
xor XOR2 (N28, N9, N2);
xor XOR2 (N29, N7, N8);
nor NOR3 (N30, N3, N10, N3);
xor XOR2 (N31, N27, N23);
not NOT1 (N32, N19);
nor NOR2 (N33, N30, N24);
nor NOR2 (N34, N8, N31);
buf BUF1 (N35, N23);
buf BUF1 (N36, N34);
nor NOR4 (N37, N20, N20, N21, N10);
not NOT1 (N38, N26);
nand NAND2 (N39, N2, N7);
and AND2 (N40, N35, N22);
and AND4 (N41, N37, N23, N26, N27);
and AND3 (N42, N41, N13, N41);
and AND4 (N43, N28, N11, N21, N17);
xor XOR2 (N44, N43, N26);
or OR3 (N45, N39, N25, N29);
not NOT1 (N46, N26);
not NOT1 (N47, N32);
nand NAND3 (N48, N47, N23, N45);
nand NAND3 (N49, N41, N21, N14);
nor NOR3 (N50, N40, N2, N38);
not NOT1 (N51, N45);
and AND3 (N52, N50, N23, N14);
or OR2 (N53, N51, N12);
and AND4 (N54, N33, N35, N2, N35);
not NOT1 (N55, N49);
nand NAND3 (N56, N44, N25, N5);
not NOT1 (N57, N48);
nor NOR4 (N58, N55, N57, N24, N30);
xor XOR2 (N59, N54, N40);
not NOT1 (N60, N1);
or OR2 (N61, N53, N11);
and AND2 (N62, N59, N14);
xor XOR2 (N63, N58, N58);
nand NAND3 (N64, N56, N20, N28);
nand NAND2 (N65, N46, N16);
and AND4 (N66, N63, N34, N18, N47);
buf BUF1 (N67, N61);
and AND2 (N68, N67, N21);
or OR4 (N69, N42, N31, N33, N50);
buf BUF1 (N70, N68);
not NOT1 (N71, N52);
nor NOR2 (N72, N36, N30);
not NOT1 (N73, N71);
nor NOR4 (N74, N62, N52, N9, N73);
and AND2 (N75, N21, N44);
or OR3 (N76, N15, N70, N58);
buf BUF1 (N77, N50);
xor XOR2 (N78, N69, N57);
buf BUF1 (N79, N72);
xor XOR2 (N80, N76, N52);
nor NOR3 (N81, N78, N15, N19);
nor NOR2 (N82, N74, N18);
buf BUF1 (N83, N82);
xor XOR2 (N84, N60, N41);
nor NOR2 (N85, N75, N58);
nor NOR2 (N86, N79, N15);
xor XOR2 (N87, N80, N1);
nor NOR3 (N88, N84, N59, N46);
and AND2 (N89, N83, N7);
buf BUF1 (N90, N88);
nand NAND2 (N91, N65, N34);
and AND4 (N92, N81, N80, N68, N41);
or OR4 (N93, N86, N63, N17, N78);
buf BUF1 (N94, N77);
nor NOR3 (N95, N87, N50, N48);
nor NOR3 (N96, N90, N83, N21);
and AND4 (N97, N94, N4, N14, N47);
and AND2 (N98, N89, N50);
xor XOR2 (N99, N93, N53);
and AND2 (N100, N85, N58);
nand NAND4 (N101, N64, N46, N83, N80);
xor XOR2 (N102, N100, N84);
buf BUF1 (N103, N97);
nand NAND3 (N104, N91, N81, N35);
or OR2 (N105, N66, N95);
nand NAND2 (N106, N47, N38);
xor XOR2 (N107, N99, N63);
and AND4 (N108, N96, N18, N103, N39);
or OR4 (N109, N16, N45, N33, N80);
and AND2 (N110, N92, N25);
nor NOR4 (N111, N110, N41, N16, N87);
xor XOR2 (N112, N109, N69);
not NOT1 (N113, N98);
not NOT1 (N114, N113);
and AND3 (N115, N105, N92, N17);
or OR3 (N116, N108, N31, N68);
nand NAND2 (N117, N112, N87);
nor NOR4 (N118, N111, N12, N8, N44);
not NOT1 (N119, N115);
xor XOR2 (N120, N116, N90);
nand NAND2 (N121, N118, N46);
or OR2 (N122, N117, N32);
buf BUF1 (N123, N104);
buf BUF1 (N124, N114);
buf BUF1 (N125, N102);
not NOT1 (N126, N119);
not NOT1 (N127, N124);
buf BUF1 (N128, N125);
nand NAND2 (N129, N126, N67);
or OR4 (N130, N107, N118, N10, N90);
or OR2 (N131, N123, N28);
nand NAND3 (N132, N130, N78, N49);
xor XOR2 (N133, N121, N118);
buf BUF1 (N134, N132);
xor XOR2 (N135, N129, N27);
buf BUF1 (N136, N131);
buf BUF1 (N137, N120);
or OR4 (N138, N106, N42, N71, N83);
and AND4 (N139, N138, N58, N81, N114);
not NOT1 (N140, N122);
xor XOR2 (N141, N140, N16);
nand NAND4 (N142, N133, N113, N46, N22);
and AND3 (N143, N127, N46, N68);
xor XOR2 (N144, N139, N93);
or OR4 (N145, N137, N41, N97, N12);
xor XOR2 (N146, N136, N104);
nand NAND4 (N147, N101, N118, N133, N7);
not NOT1 (N148, N146);
nand NAND3 (N149, N135, N2, N48);
and AND2 (N150, N134, N45);
nand NAND3 (N151, N141, N140, N54);
nand NAND4 (N152, N149, N113, N76, N86);
buf BUF1 (N153, N147);
nand NAND3 (N154, N145, N21, N142);
buf BUF1 (N155, N131);
xor XOR2 (N156, N155, N43);
buf BUF1 (N157, N143);
buf BUF1 (N158, N157);
xor XOR2 (N159, N154, N58);
and AND4 (N160, N144, N75, N1, N155);
nand NAND3 (N161, N160, N86, N83);
and AND2 (N162, N159, N15);
nor NOR4 (N163, N153, N9, N34, N118);
xor XOR2 (N164, N156, N161);
nand NAND3 (N165, N133, N144, N122);
nand NAND2 (N166, N158, N1);
not NOT1 (N167, N150);
not NOT1 (N168, N128);
nor NOR2 (N169, N152, N21);
buf BUF1 (N170, N167);
not NOT1 (N171, N168);
nor NOR2 (N172, N171, N120);
xor XOR2 (N173, N162, N96);
xor XOR2 (N174, N165, N103);
or OR3 (N175, N166, N63, N174);
or OR3 (N176, N85, N35, N123);
buf BUF1 (N177, N172);
and AND3 (N178, N151, N118, N138);
nor NOR4 (N179, N176, N148, N66, N113);
and AND2 (N180, N86, N148);
not NOT1 (N181, N180);
not NOT1 (N182, N163);
nor NOR4 (N183, N178, N144, N29, N14);
nor NOR2 (N184, N169, N15);
nand NAND2 (N185, N164, N48);
buf BUF1 (N186, N177);
and AND4 (N187, N184, N98, N95, N160);
nand NAND4 (N188, N179, N124, N176, N61);
xor XOR2 (N189, N175, N103);
not NOT1 (N190, N189);
or OR4 (N191, N181, N16, N74, N72);
or OR3 (N192, N188, N84, N132);
nor NOR4 (N193, N185, N22, N152, N130);
buf BUF1 (N194, N182);
and AND2 (N195, N193, N127);
nand NAND3 (N196, N192, N10, N63);
and AND2 (N197, N196, N83);
not NOT1 (N198, N190);
nor NOR4 (N199, N186, N48, N150, N88);
and AND2 (N200, N197, N88);
not NOT1 (N201, N200);
or OR3 (N202, N195, N36, N153);
xor XOR2 (N203, N173, N134);
or OR2 (N204, N201, N45);
and AND4 (N205, N203, N9, N64, N151);
xor XOR2 (N206, N199, N58);
nor NOR3 (N207, N198, N150, N189);
or OR4 (N208, N205, N122, N111, N78);
or OR4 (N209, N207, N39, N56, N41);
and AND4 (N210, N191, N118, N45, N160);
and AND2 (N211, N210, N84);
nor NOR2 (N212, N206, N13);
or OR2 (N213, N212, N191);
nor NOR3 (N214, N211, N34, N145);
nor NOR2 (N215, N183, N73);
xor XOR2 (N216, N213, N96);
and AND3 (N217, N187, N123, N66);
or OR3 (N218, N216, N93, N95);
not NOT1 (N219, N209);
buf BUF1 (N220, N194);
or OR3 (N221, N214, N220, N191);
not NOT1 (N222, N171);
nor NOR4 (N223, N219, N173, N150, N189);
not NOT1 (N224, N218);
nor NOR2 (N225, N215, N224);
xor XOR2 (N226, N107, N8);
not NOT1 (N227, N204);
nand NAND3 (N228, N221, N130, N178);
not NOT1 (N229, N170);
xor XOR2 (N230, N229, N192);
or OR2 (N231, N228, N105);
or OR2 (N232, N223, N70);
not NOT1 (N233, N231);
xor XOR2 (N234, N232, N28);
xor XOR2 (N235, N226, N234);
or OR4 (N236, N58, N228, N154, N187);
or OR2 (N237, N235, N9);
nor NOR2 (N238, N225, N37);
nand NAND2 (N239, N222, N183);
or OR4 (N240, N238, N67, N231, N230);
nor NOR2 (N241, N64, N13);
buf BUF1 (N242, N217);
nand NAND2 (N243, N239, N97);
xor XOR2 (N244, N236, N168);
buf BUF1 (N245, N243);
nand NAND4 (N246, N244, N150, N174, N139);
nor NOR4 (N247, N241, N56, N238, N241);
nor NOR3 (N248, N245, N172, N237);
or OR4 (N249, N47, N120, N58, N231);
buf BUF1 (N250, N227);
not NOT1 (N251, N247);
buf BUF1 (N252, N251);
nand NAND4 (N253, N242, N132, N32, N19);
xor XOR2 (N254, N208, N127);
buf BUF1 (N255, N249);
or OR2 (N256, N248, N171);
and AND2 (N257, N256, N121);
nor NOR2 (N258, N257, N13);
not NOT1 (N259, N255);
or OR4 (N260, N253, N32, N72, N43);
nor NOR2 (N261, N250, N228);
and AND4 (N262, N252, N115, N240, N87);
nand NAND4 (N263, N90, N240, N121, N185);
buf BUF1 (N264, N261);
xor XOR2 (N265, N264, N152);
or OR3 (N266, N246, N88, N111);
xor XOR2 (N267, N263, N92);
nand NAND3 (N268, N233, N181, N52);
nor NOR2 (N269, N202, N153);
buf BUF1 (N270, N267);
nand NAND2 (N271, N266, N73);
nor NOR3 (N272, N254, N190, N86);
and AND3 (N273, N272, N25, N88);
nand NAND2 (N274, N270, N240);
and AND3 (N275, N269, N232, N75);
nor NOR3 (N276, N268, N27, N164);
and AND3 (N277, N276, N267, N44);
and AND3 (N278, N259, N77, N154);
xor XOR2 (N279, N271, N32);
xor XOR2 (N280, N279, N134);
buf BUF1 (N281, N278);
nor NOR4 (N282, N275, N86, N95, N85);
and AND2 (N283, N274, N210);
nand NAND4 (N284, N277, N58, N10, N224);
or OR4 (N285, N283, N176, N30, N267);
not NOT1 (N286, N273);
nor NOR4 (N287, N262, N37, N284, N38);
nor NOR2 (N288, N187, N237);
buf BUF1 (N289, N286);
and AND2 (N290, N281, N245);
nand NAND4 (N291, N258, N140, N132, N172);
and AND4 (N292, N285, N191, N288, N69);
or OR2 (N293, N211, N106);
buf BUF1 (N294, N265);
or OR3 (N295, N280, N4, N101);
nand NAND3 (N296, N291, N236, N193);
or OR2 (N297, N287, N222);
xor XOR2 (N298, N297, N108);
xor XOR2 (N299, N292, N75);
or OR2 (N300, N295, N243);
nand NAND4 (N301, N289, N208, N72, N167);
or OR4 (N302, N296, N202, N212, N43);
nand NAND4 (N303, N301, N147, N199, N165);
not NOT1 (N304, N290);
and AND2 (N305, N302, N113);
or OR3 (N306, N304, N174, N87);
not NOT1 (N307, N294);
nand NAND3 (N308, N260, N33, N153);
buf BUF1 (N309, N299);
nand NAND4 (N310, N309, N235, N304, N269);
or OR4 (N311, N282, N166, N143, N258);
buf BUF1 (N312, N310);
not NOT1 (N313, N293);
nor NOR3 (N314, N298, N107, N51);
not NOT1 (N315, N308);
xor XOR2 (N316, N305, N115);
xor XOR2 (N317, N315, N36);
xor XOR2 (N318, N316, N53);
nor NOR4 (N319, N311, N236, N274, N166);
buf BUF1 (N320, N313);
not NOT1 (N321, N300);
buf BUF1 (N322, N317);
xor XOR2 (N323, N320, N181);
and AND2 (N324, N322, N13);
and AND3 (N325, N312, N220, N99);
buf BUF1 (N326, N303);
nand NAND3 (N327, N314, N166, N210);
xor XOR2 (N328, N324, N305);
not NOT1 (N329, N307);
and AND3 (N330, N325, N283, N296);
nand NAND2 (N331, N326, N72);
or OR4 (N332, N319, N283, N249, N40);
or OR4 (N333, N327, N114, N65, N32);
not NOT1 (N334, N318);
buf BUF1 (N335, N323);
not NOT1 (N336, N335);
nand NAND3 (N337, N333, N77, N184);
nor NOR4 (N338, N329, N198, N91, N116);
and AND2 (N339, N331, N279);
and AND4 (N340, N306, N86, N158, N97);
or OR4 (N341, N339, N139, N143, N217);
buf BUF1 (N342, N341);
nand NAND3 (N343, N336, N266, N241);
xor XOR2 (N344, N321, N152);
nor NOR2 (N345, N328, N161);
nand NAND2 (N346, N345, N254);
nand NAND4 (N347, N334, N125, N90, N298);
or OR3 (N348, N342, N189, N312);
not NOT1 (N349, N337);
and AND4 (N350, N332, N43, N295, N239);
nor NOR2 (N351, N340, N262);
nor NOR4 (N352, N330, N294, N88, N161);
or OR2 (N353, N338, N247);
xor XOR2 (N354, N343, N171);
and AND3 (N355, N346, N263, N79);
nand NAND4 (N356, N344, N249, N22, N182);
xor XOR2 (N357, N347, N69);
nand NAND2 (N358, N349, N219);
or OR2 (N359, N355, N240);
xor XOR2 (N360, N350, N280);
not NOT1 (N361, N357);
nand NAND3 (N362, N353, N297, N281);
nand NAND2 (N363, N362, N172);
and AND2 (N364, N358, N189);
or OR3 (N365, N351, N359, N74);
and AND2 (N366, N87, N208);
nand NAND2 (N367, N348, N237);
and AND3 (N368, N363, N42, N144);
nand NAND3 (N369, N356, N285, N297);
and AND3 (N370, N369, N57, N270);
or OR3 (N371, N361, N207, N7);
buf BUF1 (N372, N368);
xor XOR2 (N373, N372, N64);
nand NAND3 (N374, N360, N29, N315);
and AND4 (N375, N364, N221, N367, N12);
not NOT1 (N376, N348);
nor NOR4 (N377, N371, N235, N183, N51);
not NOT1 (N378, N366);
xor XOR2 (N379, N377, N7);
xor XOR2 (N380, N370, N17);
not NOT1 (N381, N352);
or OR2 (N382, N354, N51);
not NOT1 (N383, N382);
not NOT1 (N384, N381);
or OR2 (N385, N373, N361);
and AND2 (N386, N374, N269);
buf BUF1 (N387, N378);
nand NAND2 (N388, N380, N12);
not NOT1 (N389, N388);
not NOT1 (N390, N365);
or OR3 (N391, N390, N203, N23);
nor NOR4 (N392, N386, N106, N305, N386);
nand NAND4 (N393, N392, N227, N148, N387);
xor XOR2 (N394, N225, N307);
or OR4 (N395, N376, N276, N338, N386);
xor XOR2 (N396, N379, N55);
or OR3 (N397, N393, N396, N241);
buf BUF1 (N398, N154);
xor XOR2 (N399, N394, N188);
buf BUF1 (N400, N395);
not NOT1 (N401, N384);
nor NOR2 (N402, N385, N156);
and AND2 (N403, N401, N387);
and AND3 (N404, N389, N83, N18);
not NOT1 (N405, N399);
or OR3 (N406, N398, N392, N392);
nor NOR2 (N407, N406, N45);
nand NAND4 (N408, N397, N100, N86, N80);
or OR4 (N409, N383, N167, N177, N135);
nor NOR2 (N410, N404, N340);
nand NAND2 (N411, N402, N200);
xor XOR2 (N412, N407, N297);
nand NAND3 (N413, N403, N174, N47);
nor NOR3 (N414, N411, N75, N40);
not NOT1 (N415, N412);
xor XOR2 (N416, N410, N283);
not NOT1 (N417, N375);
not NOT1 (N418, N415);
xor XOR2 (N419, N405, N411);
buf BUF1 (N420, N419);
nor NOR4 (N421, N413, N355, N80, N11);
or OR3 (N422, N420, N201, N357);
buf BUF1 (N423, N414);
and AND4 (N424, N391, N3, N78, N314);
nor NOR4 (N425, N418, N263, N168, N88);
buf BUF1 (N426, N416);
xor XOR2 (N427, N421, N173);
nand NAND3 (N428, N426, N142, N43);
buf BUF1 (N429, N428);
nor NOR2 (N430, N424, N149);
and AND3 (N431, N408, N91, N202);
buf BUF1 (N432, N431);
nor NOR2 (N433, N432, N207);
not NOT1 (N434, N409);
and AND2 (N435, N400, N91);
not NOT1 (N436, N422);
nor NOR4 (N437, N429, N294, N173, N288);
xor XOR2 (N438, N427, N107);
buf BUF1 (N439, N430);
nand NAND2 (N440, N437, N386);
nand NAND4 (N441, N439, N36, N210, N267);
nand NAND3 (N442, N440, N141, N369);
nand NAND3 (N443, N436, N355, N250);
or OR3 (N444, N438, N163, N78);
xor XOR2 (N445, N442, N10);
nor NOR2 (N446, N444, N62);
not NOT1 (N447, N445);
nand NAND4 (N448, N425, N261, N3, N247);
buf BUF1 (N449, N433);
xor XOR2 (N450, N448, N278);
or OR3 (N451, N417, N180, N244);
and AND2 (N452, N446, N224);
or OR2 (N453, N450, N169);
not NOT1 (N454, N449);
and AND2 (N455, N435, N348);
or OR2 (N456, N447, N73);
nand NAND4 (N457, N443, N387, N181, N296);
not NOT1 (N458, N423);
buf BUF1 (N459, N451);
and AND3 (N460, N441, N413, N184);
buf BUF1 (N461, N458);
nand NAND3 (N462, N460, N112, N438);
xor XOR2 (N463, N462, N435);
nor NOR2 (N464, N457, N262);
nand NAND3 (N465, N459, N158, N164);
nor NOR2 (N466, N455, N158);
xor XOR2 (N467, N463, N280);
or OR4 (N468, N452, N158, N463, N399);
nand NAND2 (N469, N466, N366);
nand NAND2 (N470, N469, N342);
nand NAND3 (N471, N468, N369, N206);
and AND2 (N472, N465, N112);
and AND2 (N473, N453, N380);
or OR4 (N474, N434, N135, N425, N166);
xor XOR2 (N475, N461, N83);
xor XOR2 (N476, N467, N240);
nand NAND2 (N477, N471, N19);
xor XOR2 (N478, N470, N41);
or OR3 (N479, N472, N428, N100);
xor XOR2 (N480, N454, N187);
not NOT1 (N481, N456);
buf BUF1 (N482, N477);
xor XOR2 (N483, N481, N341);
or OR2 (N484, N464, N113);
nand NAND3 (N485, N480, N174, N85);
nand NAND2 (N486, N482, N16);
nand NAND4 (N487, N483, N169, N66, N287);
not NOT1 (N488, N485);
or OR4 (N489, N486, N348, N163, N308);
nand NAND4 (N490, N479, N300, N387, N486);
nand NAND4 (N491, N488, N211, N272, N171);
and AND4 (N492, N474, N331, N347, N22);
buf BUF1 (N493, N473);
buf BUF1 (N494, N476);
nor NOR3 (N495, N489, N368, N389);
or OR4 (N496, N490, N409, N42, N79);
xor XOR2 (N497, N491, N319);
xor XOR2 (N498, N494, N410);
not NOT1 (N499, N492);
not NOT1 (N500, N497);
nor NOR3 (N501, N478, N251, N39);
nand NAND2 (N502, N475, N160);
or OR4 (N503, N498, N74, N469, N485);
nand NAND3 (N504, N501, N472, N387);
xor XOR2 (N505, N484, N408);
nand NAND4 (N506, N500, N437, N426, N197);
nand NAND3 (N507, N503, N102, N184);
not NOT1 (N508, N506);
nor NOR4 (N509, N507, N493, N401, N345);
nand NAND4 (N510, N377, N120, N152, N342);
nand NAND4 (N511, N487, N198, N76, N346);
and AND3 (N512, N505, N259, N34);
or OR2 (N513, N496, N467);
or OR3 (N514, N509, N443, N447);
and AND2 (N515, N495, N175);
buf BUF1 (N516, N513);
or OR2 (N517, N512, N41);
nand NAND4 (N518, N502, N45, N451, N359);
nor NOR2 (N519, N515, N153);
buf BUF1 (N520, N514);
xor XOR2 (N521, N517, N498);
nor NOR3 (N522, N516, N59, N184);
nor NOR3 (N523, N521, N90, N175);
xor XOR2 (N524, N518, N444);
or OR3 (N525, N523, N42, N150);
nand NAND2 (N526, N524, N130);
and AND2 (N527, N522, N520);
nor NOR2 (N528, N71, N119);
xor XOR2 (N529, N527, N261);
or OR3 (N530, N499, N181, N473);
and AND4 (N531, N511, N400, N200, N115);
nor NOR2 (N532, N530, N177);
nand NAND2 (N533, N525, N279);
buf BUF1 (N534, N531);
xor XOR2 (N535, N529, N200);
and AND2 (N536, N504, N212);
not NOT1 (N537, N526);
nor NOR4 (N538, N537, N496, N259, N209);
and AND2 (N539, N532, N381);
nor NOR4 (N540, N510, N69, N322, N431);
nor NOR3 (N541, N533, N271, N295);
nand NAND4 (N542, N539, N123, N68, N454);
buf BUF1 (N543, N536);
and AND2 (N544, N538, N318);
and AND4 (N545, N542, N61, N30, N119);
not NOT1 (N546, N541);
nor NOR3 (N547, N545, N370, N495);
buf BUF1 (N548, N540);
and AND2 (N549, N519, N199);
buf BUF1 (N550, N548);
or OR2 (N551, N535, N307);
and AND2 (N552, N528, N408);
buf BUF1 (N553, N550);
xor XOR2 (N554, N552, N227);
not NOT1 (N555, N551);
and AND2 (N556, N553, N262);
or OR4 (N557, N508, N358, N163, N527);
buf BUF1 (N558, N557);
not NOT1 (N559, N558);
and AND4 (N560, N543, N375, N316, N25);
buf BUF1 (N561, N560);
nor NOR3 (N562, N554, N549, N468);
nand NAND3 (N563, N274, N525, N229);
nand NAND3 (N564, N544, N93, N340);
nor NOR4 (N565, N563, N50, N144, N78);
nor NOR2 (N566, N559, N371);
and AND3 (N567, N534, N364, N230);
buf BUF1 (N568, N561);
buf BUF1 (N569, N567);
xor XOR2 (N570, N569, N268);
not NOT1 (N571, N564);
not NOT1 (N572, N562);
xor XOR2 (N573, N555, N88);
and AND3 (N574, N572, N137, N345);
nand NAND3 (N575, N566, N303, N16);
or OR4 (N576, N547, N569, N17, N44);
xor XOR2 (N577, N568, N541);
nor NOR3 (N578, N577, N142, N388);
and AND4 (N579, N578, N567, N370, N370);
buf BUF1 (N580, N574);
not NOT1 (N581, N575);
or OR3 (N582, N573, N156, N181);
and AND3 (N583, N565, N242, N566);
nand NAND2 (N584, N581, N382);
nand NAND3 (N585, N570, N479, N128);
nand NAND3 (N586, N580, N250, N413);
xor XOR2 (N587, N556, N33);
and AND3 (N588, N582, N42, N258);
not NOT1 (N589, N579);
not NOT1 (N590, N589);
buf BUF1 (N591, N583);
and AND2 (N592, N584, N209);
xor XOR2 (N593, N588, N318);
nand NAND2 (N594, N571, N210);
nor NOR2 (N595, N585, N404);
nand NAND2 (N596, N594, N439);
or OR4 (N597, N576, N454, N481, N420);
nand NAND4 (N598, N587, N57, N350, N371);
xor XOR2 (N599, N592, N503);
or OR3 (N600, N599, N485, N352);
nor NOR2 (N601, N596, N301);
buf BUF1 (N602, N593);
or OR3 (N603, N598, N370, N268);
not NOT1 (N604, N601);
and AND2 (N605, N602, N1);
not NOT1 (N606, N591);
nor NOR4 (N607, N603, N92, N477, N189);
nand NAND4 (N608, N605, N403, N229, N594);
nand NAND2 (N609, N597, N216);
xor XOR2 (N610, N595, N364);
and AND3 (N611, N586, N45, N8);
not NOT1 (N612, N611);
buf BUF1 (N613, N612);
xor XOR2 (N614, N604, N154);
not NOT1 (N615, N590);
buf BUF1 (N616, N546);
not NOT1 (N617, N609);
and AND2 (N618, N616, N536);
xor XOR2 (N619, N617, N210);
nand NAND4 (N620, N614, N134, N394, N532);
nand NAND2 (N621, N620, N546);
nand NAND2 (N622, N621, N82);
not NOT1 (N623, N615);
and AND3 (N624, N610, N376, N97);
and AND2 (N625, N618, N183);
and AND2 (N626, N623, N600);
nor NOR4 (N627, N503, N3, N123, N260);
nor NOR2 (N628, N625, N435);
buf BUF1 (N629, N628);
and AND4 (N630, N619, N80, N311, N579);
not NOT1 (N631, N626);
nand NAND4 (N632, N608, N396, N284, N144);
nor NOR3 (N633, N632, N96, N252);
xor XOR2 (N634, N629, N189);
buf BUF1 (N635, N624);
xor XOR2 (N636, N634, N379);
not NOT1 (N637, N635);
and AND2 (N638, N607, N584);
nor NOR2 (N639, N630, N465);
or OR3 (N640, N636, N263, N340);
xor XOR2 (N641, N640, N551);
xor XOR2 (N642, N633, N1);
and AND2 (N643, N627, N196);
nor NOR3 (N644, N606, N501, N391);
xor XOR2 (N645, N644, N482);
nor NOR3 (N646, N638, N329, N495);
buf BUF1 (N647, N645);
and AND2 (N648, N642, N616);
or OR3 (N649, N643, N252, N605);
nor NOR2 (N650, N613, N286);
nand NAND3 (N651, N649, N495, N460);
and AND4 (N652, N631, N368, N279, N144);
buf BUF1 (N653, N650);
or OR4 (N654, N646, N69, N331, N41);
buf BUF1 (N655, N639);
nor NOR2 (N656, N653, N264);
nor NOR2 (N657, N647, N624);
nand NAND2 (N658, N652, N295);
nand NAND3 (N659, N648, N200, N254);
nand NAND3 (N660, N651, N91, N490);
not NOT1 (N661, N655);
or OR4 (N662, N654, N504, N520, N215);
buf BUF1 (N663, N641);
nand NAND2 (N664, N637, N596);
nand NAND4 (N665, N661, N356, N432, N491);
nor NOR3 (N666, N657, N612, N278);
buf BUF1 (N667, N658);
nor NOR2 (N668, N665, N420);
nand NAND2 (N669, N660, N448);
or OR4 (N670, N662, N189, N427, N650);
or OR2 (N671, N670, N40);
and AND3 (N672, N668, N382, N154);
nor NOR4 (N673, N671, N540, N56, N339);
xor XOR2 (N674, N622, N300);
or OR4 (N675, N669, N257, N123, N345);
xor XOR2 (N676, N659, N18);
not NOT1 (N677, N676);
buf BUF1 (N678, N675);
not NOT1 (N679, N663);
not NOT1 (N680, N679);
and AND2 (N681, N680, N96);
buf BUF1 (N682, N674);
nor NOR2 (N683, N673, N533);
not NOT1 (N684, N678);
nor NOR4 (N685, N684, N189, N100, N416);
xor XOR2 (N686, N667, N186);
nand NAND4 (N687, N682, N322, N298, N107);
nor NOR2 (N688, N656, N459);
xor XOR2 (N689, N681, N439);
not NOT1 (N690, N685);
and AND2 (N691, N664, N49);
buf BUF1 (N692, N689);
buf BUF1 (N693, N691);
nor NOR2 (N694, N677, N630);
and AND3 (N695, N672, N21, N78);
buf BUF1 (N696, N666);
not NOT1 (N697, N692);
and AND4 (N698, N686, N103, N489, N426);
xor XOR2 (N699, N687, N360);
nor NOR4 (N700, N699, N200, N574, N449);
not NOT1 (N701, N697);
or OR4 (N702, N696, N653, N679, N144);
xor XOR2 (N703, N683, N255);
buf BUF1 (N704, N698);
buf BUF1 (N705, N694);
and AND3 (N706, N701, N473, N207);
or OR4 (N707, N705, N61, N579, N569);
and AND3 (N708, N706, N64, N423);
nand NAND3 (N709, N690, N579, N232);
and AND2 (N710, N704, N513);
nor NOR4 (N711, N700, N380, N205, N551);
buf BUF1 (N712, N688);
not NOT1 (N713, N710);
not NOT1 (N714, N702);
xor XOR2 (N715, N695, N430);
nand NAND4 (N716, N714, N73, N103, N132);
nand NAND4 (N717, N713, N317, N94, N130);
and AND4 (N718, N711, N360, N308, N571);
nand NAND2 (N719, N717, N598);
nand NAND2 (N720, N708, N103);
nand NAND3 (N721, N707, N212, N679);
buf BUF1 (N722, N716);
and AND2 (N723, N709, N394);
buf BUF1 (N724, N712);
xor XOR2 (N725, N724, N435);
not NOT1 (N726, N715);
buf BUF1 (N727, N693);
nand NAND3 (N728, N725, N344, N249);
nand NAND4 (N729, N722, N642, N651, N532);
buf BUF1 (N730, N703);
nor NOR4 (N731, N728, N526, N479, N691);
not NOT1 (N732, N731);
buf BUF1 (N733, N723);
xor XOR2 (N734, N719, N136);
nand NAND2 (N735, N730, N403);
not NOT1 (N736, N727);
nand NAND3 (N737, N718, N412, N458);
xor XOR2 (N738, N735, N106);
not NOT1 (N739, N721);
nor NOR4 (N740, N732, N521, N136, N178);
not NOT1 (N741, N738);
nor NOR4 (N742, N737, N352, N198, N602);
xor XOR2 (N743, N734, N165);
or OR4 (N744, N733, N691, N717, N153);
or OR4 (N745, N739, N718, N224, N181);
nor NOR4 (N746, N726, N410, N565, N635);
or OR2 (N747, N742, N697);
not NOT1 (N748, N745);
buf BUF1 (N749, N720);
nor NOR2 (N750, N744, N99);
not NOT1 (N751, N740);
buf BUF1 (N752, N736);
nand NAND3 (N753, N729, N679, N487);
buf BUF1 (N754, N752);
nand NAND4 (N755, N750, N62, N31, N248);
not NOT1 (N756, N749);
nand NAND4 (N757, N748, N299, N427, N56);
or OR2 (N758, N753, N594);
or OR3 (N759, N758, N592, N382);
and AND3 (N760, N743, N725, N669);
nand NAND3 (N761, N751, N580, N661);
xor XOR2 (N762, N755, N759);
and AND3 (N763, N439, N561, N129);
not NOT1 (N764, N741);
buf BUF1 (N765, N756);
xor XOR2 (N766, N754, N379);
not NOT1 (N767, N764);
or OR3 (N768, N767, N231, N381);
not NOT1 (N769, N765);
nand NAND2 (N770, N761, N669);
nand NAND3 (N771, N770, N260, N457);
and AND2 (N772, N766, N564);
and AND3 (N773, N769, N259, N256);
not NOT1 (N774, N757);
buf BUF1 (N775, N763);
nand NAND3 (N776, N768, N745, N282);
or OR3 (N777, N747, N207, N378);
or OR4 (N778, N771, N484, N181, N678);
buf BUF1 (N779, N776);
and AND3 (N780, N779, N317, N187);
nor NOR3 (N781, N746, N607, N754);
nand NAND4 (N782, N781, N560, N504, N366);
and AND4 (N783, N773, N35, N543, N97);
not NOT1 (N784, N762);
nand NAND3 (N785, N775, N501, N190);
or OR3 (N786, N785, N597, N757);
nand NAND3 (N787, N783, N47, N454);
nor NOR2 (N788, N778, N346);
xor XOR2 (N789, N780, N122);
or OR3 (N790, N789, N39, N536);
and AND2 (N791, N788, N762);
buf BUF1 (N792, N760);
not NOT1 (N793, N791);
nand NAND4 (N794, N774, N699, N109, N45);
nand NAND2 (N795, N782, N8);
buf BUF1 (N796, N795);
xor XOR2 (N797, N787, N668);
and AND3 (N798, N786, N11, N619);
xor XOR2 (N799, N777, N408);
nor NOR3 (N800, N798, N710, N732);
buf BUF1 (N801, N800);
or OR2 (N802, N797, N169);
xor XOR2 (N803, N801, N529);
nand NAND3 (N804, N802, N305, N455);
nand NAND3 (N805, N799, N638, N635);
not NOT1 (N806, N784);
buf BUF1 (N807, N806);
buf BUF1 (N808, N807);
buf BUF1 (N809, N808);
nand NAND3 (N810, N772, N691, N414);
or OR4 (N811, N794, N651, N416, N51);
nand NAND2 (N812, N810, N332);
nor NOR2 (N813, N804, N673);
buf BUF1 (N814, N809);
nor NOR3 (N815, N811, N615, N456);
not NOT1 (N816, N796);
nor NOR3 (N817, N814, N574, N561);
nand NAND3 (N818, N812, N620, N133);
buf BUF1 (N819, N815);
or OR2 (N820, N813, N25);
nor NOR3 (N821, N819, N302, N397);
not NOT1 (N822, N818);
nor NOR4 (N823, N820, N460, N181, N786);
nor NOR4 (N824, N793, N323, N446, N12);
not NOT1 (N825, N823);
buf BUF1 (N826, N790);
or OR3 (N827, N817, N280, N792);
not NOT1 (N828, N774);
nor NOR4 (N829, N803, N326, N112, N330);
and AND4 (N830, N816, N175, N640, N470);
and AND4 (N831, N826, N684, N28, N708);
xor XOR2 (N832, N828, N785);
xor XOR2 (N833, N830, N330);
xor XOR2 (N834, N825, N34);
not NOT1 (N835, N821);
xor XOR2 (N836, N829, N467);
or OR3 (N837, N822, N377, N533);
not NOT1 (N838, N824);
nor NOR2 (N839, N834, N738);
or OR4 (N840, N839, N815, N695, N242);
xor XOR2 (N841, N832, N636);
buf BUF1 (N842, N836);
xor XOR2 (N843, N840, N838);
nand NAND3 (N844, N262, N175, N774);
xor XOR2 (N845, N841, N283);
not NOT1 (N846, N805);
or OR3 (N847, N827, N814, N186);
buf BUF1 (N848, N843);
buf BUF1 (N849, N848);
nand NAND3 (N850, N837, N627, N283);
and AND4 (N851, N833, N572, N120, N121);
nand NAND2 (N852, N849, N846);
or OR2 (N853, N82, N571);
nand NAND3 (N854, N831, N673, N339);
buf BUF1 (N855, N852);
nand NAND2 (N856, N847, N791);
buf BUF1 (N857, N855);
xor XOR2 (N858, N845, N169);
xor XOR2 (N859, N850, N824);
buf BUF1 (N860, N851);
buf BUF1 (N861, N844);
not NOT1 (N862, N858);
nand NAND4 (N863, N854, N536, N279, N321);
and AND3 (N864, N856, N678, N643);
nand NAND3 (N865, N853, N579, N300);
xor XOR2 (N866, N835, N421);
xor XOR2 (N867, N861, N511);
nand NAND4 (N868, N863, N67, N253, N232);
xor XOR2 (N869, N842, N527);
nor NOR4 (N870, N865, N278, N436, N534);
not NOT1 (N871, N868);
not NOT1 (N872, N869);
buf BUF1 (N873, N862);
buf BUF1 (N874, N857);
buf BUF1 (N875, N860);
buf BUF1 (N876, N872);
not NOT1 (N877, N871);
or OR4 (N878, N870, N465, N71, N368);
or OR3 (N879, N859, N292, N875);
buf BUF1 (N880, N292);
nand NAND4 (N881, N876, N495, N88, N782);
nand NAND3 (N882, N881, N156, N56);
nor NOR3 (N883, N866, N715, N370);
and AND4 (N884, N878, N88, N753, N479);
not NOT1 (N885, N867);
or OR3 (N886, N880, N370, N65);
buf BUF1 (N887, N882);
xor XOR2 (N888, N883, N632);
xor XOR2 (N889, N874, N588);
not NOT1 (N890, N884);
nor NOR4 (N891, N877, N93, N201, N488);
nor NOR4 (N892, N889, N647, N573, N60);
xor XOR2 (N893, N873, N196);
buf BUF1 (N894, N891);
xor XOR2 (N895, N879, N847);
buf BUF1 (N896, N895);
xor XOR2 (N897, N896, N828);
nand NAND4 (N898, N886, N627, N211, N258);
xor XOR2 (N899, N885, N592);
nand NAND2 (N900, N864, N763);
and AND3 (N901, N900, N271, N622);
and AND4 (N902, N888, N588, N200, N743);
buf BUF1 (N903, N892);
nand NAND2 (N904, N903, N425);
buf BUF1 (N905, N894);
nor NOR4 (N906, N904, N142, N49, N6);
nor NOR3 (N907, N906, N481, N267);
not NOT1 (N908, N887);
buf BUF1 (N909, N902);
xor XOR2 (N910, N908, N414);
nand NAND2 (N911, N893, N681);
buf BUF1 (N912, N901);
nor NOR2 (N913, N899, N241);
nor NOR2 (N914, N905, N158);
nor NOR2 (N915, N914, N47);
and AND4 (N916, N910, N117, N708, N452);
or OR3 (N917, N913, N490, N724);
buf BUF1 (N918, N912);
not NOT1 (N919, N911);
nor NOR2 (N920, N909, N394);
nor NOR4 (N921, N916, N800, N42, N877);
buf BUF1 (N922, N915);
or OR2 (N923, N907, N295);
nor NOR3 (N924, N917, N843, N574);
nor NOR4 (N925, N919, N579, N250, N87);
nor NOR3 (N926, N920, N551, N82);
nor NOR3 (N927, N924, N795, N896);
buf BUF1 (N928, N898);
nor NOR3 (N929, N918, N419, N248);
nand NAND3 (N930, N928, N265, N866);
nand NAND4 (N931, N930, N126, N19, N789);
nor NOR4 (N932, N923, N804, N377, N846);
xor XOR2 (N933, N931, N621);
xor XOR2 (N934, N929, N836);
or OR2 (N935, N922, N159);
nand NAND2 (N936, N935, N323);
nand NAND2 (N937, N933, N478);
and AND3 (N938, N937, N108, N584);
buf BUF1 (N939, N897);
nor NOR2 (N940, N932, N612);
or OR3 (N941, N938, N415, N928);
and AND2 (N942, N934, N582);
buf BUF1 (N943, N936);
and AND3 (N944, N939, N747, N931);
buf BUF1 (N945, N927);
or OR3 (N946, N942, N572, N907);
not NOT1 (N947, N890);
buf BUF1 (N948, N944);
nor NOR4 (N949, N947, N704, N184, N614);
xor XOR2 (N950, N948, N583);
buf BUF1 (N951, N949);
and AND3 (N952, N950, N599, N938);
and AND2 (N953, N926, N240);
xor XOR2 (N954, N953, N749);
xor XOR2 (N955, N941, N660);
and AND2 (N956, N925, N21);
not NOT1 (N957, N946);
xor XOR2 (N958, N943, N332);
nor NOR4 (N959, N954, N373, N300, N732);
and AND3 (N960, N957, N603, N847);
and AND4 (N961, N955, N323, N692, N586);
buf BUF1 (N962, N958);
buf BUF1 (N963, N940);
xor XOR2 (N964, N961, N155);
nor NOR3 (N965, N921, N886, N274);
buf BUF1 (N966, N964);
nand NAND3 (N967, N952, N493, N702);
and AND2 (N968, N965, N796);
or OR3 (N969, N963, N668, N629);
xor XOR2 (N970, N962, N288);
buf BUF1 (N971, N968);
and AND4 (N972, N966, N289, N3, N40);
xor XOR2 (N973, N972, N776);
xor XOR2 (N974, N973, N259);
nor NOR2 (N975, N959, N598);
and AND4 (N976, N951, N666, N487, N136);
nand NAND2 (N977, N960, N857);
not NOT1 (N978, N974);
or OR2 (N979, N971, N31);
not NOT1 (N980, N970);
not NOT1 (N981, N945);
nand NAND4 (N982, N977, N921, N235, N658);
xor XOR2 (N983, N975, N16);
nor NOR4 (N984, N980, N552, N684, N186);
or OR3 (N985, N967, N782, N929);
xor XOR2 (N986, N984, N213);
and AND3 (N987, N969, N656, N376);
or OR3 (N988, N979, N330, N918);
and AND3 (N989, N982, N713, N273);
and AND2 (N990, N956, N169);
buf BUF1 (N991, N976);
nand NAND4 (N992, N978, N595, N85, N710);
buf BUF1 (N993, N992);
nand NAND2 (N994, N991, N889);
buf BUF1 (N995, N987);
xor XOR2 (N996, N995, N515);
nor NOR2 (N997, N996, N400);
nor NOR3 (N998, N997, N680, N559);
not NOT1 (N999, N989);
xor XOR2 (N1000, N999, N830);
xor XOR2 (N1001, N981, N891);
and AND3 (N1002, N998, N770, N523);
and AND2 (N1003, N983, N742);
buf BUF1 (N1004, N986);
nand NAND2 (N1005, N1000, N586);
xor XOR2 (N1006, N990, N333);
xor XOR2 (N1007, N1002, N348);
not NOT1 (N1008, N1003);
buf BUF1 (N1009, N1008);
xor XOR2 (N1010, N993, N203);
xor XOR2 (N1011, N1005, N731);
nor NOR3 (N1012, N1007, N919, N297);
nand NAND2 (N1013, N994, N104);
xor XOR2 (N1014, N985, N447);
xor XOR2 (N1015, N1011, N6);
xor XOR2 (N1016, N1014, N290);
xor XOR2 (N1017, N1009, N130);
nand NAND3 (N1018, N1016, N588, N321);
or OR4 (N1019, N988, N672, N587, N696);
and AND2 (N1020, N1001, N970);
not NOT1 (N1021, N1006);
buf BUF1 (N1022, N1020);
nor NOR4 (N1023, N1010, N228, N535, N322);
xor XOR2 (N1024, N1022, N974);
or OR2 (N1025, N1017, N776);
xor XOR2 (N1026, N1018, N400);
nand NAND2 (N1027, N1026, N491);
nor NOR2 (N1028, N1027, N284);
and AND2 (N1029, N1021, N333);
not NOT1 (N1030, N1024);
or OR4 (N1031, N1019, N310, N570, N937);
not NOT1 (N1032, N1023);
not NOT1 (N1033, N1025);
nor NOR3 (N1034, N1028, N642, N520);
or OR4 (N1035, N1013, N566, N143, N25);
xor XOR2 (N1036, N1031, N592);
and AND3 (N1037, N1033, N388, N653);
nand NAND4 (N1038, N1015, N784, N894, N80);
nor NOR3 (N1039, N1012, N658, N58);
nor NOR3 (N1040, N1029, N892, N904);
nor NOR4 (N1041, N1032, N121, N712, N943);
buf BUF1 (N1042, N1037);
nand NAND2 (N1043, N1030, N987);
nor NOR4 (N1044, N1004, N199, N224, N797);
xor XOR2 (N1045, N1040, N654);
nand NAND3 (N1046, N1039, N318, N810);
buf BUF1 (N1047, N1046);
and AND3 (N1048, N1043, N166, N772);
nor NOR2 (N1049, N1048, N1030);
buf BUF1 (N1050, N1035);
nor NOR4 (N1051, N1038, N1031, N658, N194);
nand NAND2 (N1052, N1034, N945);
nor NOR2 (N1053, N1047, N924);
xor XOR2 (N1054, N1051, N110);
not NOT1 (N1055, N1042);
not NOT1 (N1056, N1052);
not NOT1 (N1057, N1036);
and AND4 (N1058, N1056, N324, N199, N469);
xor XOR2 (N1059, N1053, N890);
and AND3 (N1060, N1055, N374, N326);
not NOT1 (N1061, N1044);
buf BUF1 (N1062, N1060);
nor NOR3 (N1063, N1041, N799, N211);
nor NOR3 (N1064, N1045, N432, N580);
nand NAND4 (N1065, N1061, N147, N159, N823);
nand NAND4 (N1066, N1054, N843, N176, N695);
buf BUF1 (N1067, N1050);
not NOT1 (N1068, N1066);
and AND2 (N1069, N1062, N628);
not NOT1 (N1070, N1058);
buf BUF1 (N1071, N1063);
nor NOR3 (N1072, N1057, N928, N826);
nor NOR4 (N1073, N1072, N132, N174, N455);
nor NOR3 (N1074, N1065, N885, N1054);
xor XOR2 (N1075, N1069, N205);
nand NAND3 (N1076, N1075, N928, N993);
and AND2 (N1077, N1070, N506);
and AND2 (N1078, N1064, N151);
or OR2 (N1079, N1076, N152);
or OR2 (N1080, N1073, N171);
xor XOR2 (N1081, N1068, N9);
or OR4 (N1082, N1081, N294, N428, N1070);
buf BUF1 (N1083, N1077);
or OR4 (N1084, N1079, N213, N1020, N841);
not NOT1 (N1085, N1082);
not NOT1 (N1086, N1059);
buf BUF1 (N1087, N1049);
xor XOR2 (N1088, N1086, N579);
buf BUF1 (N1089, N1083);
nor NOR2 (N1090, N1078, N865);
not NOT1 (N1091, N1090);
and AND2 (N1092, N1087, N328);
xor XOR2 (N1093, N1067, N166);
or OR4 (N1094, N1071, N255, N641, N673);
xor XOR2 (N1095, N1080, N682);
nor NOR4 (N1096, N1093, N874, N1038, N341);
buf BUF1 (N1097, N1084);
and AND3 (N1098, N1096, N44, N30);
or OR4 (N1099, N1089, N980, N472, N125);
nor NOR4 (N1100, N1097, N530, N512, N643);
buf BUF1 (N1101, N1098);
not NOT1 (N1102, N1091);
nor NOR2 (N1103, N1074, N33);
xor XOR2 (N1104, N1099, N206);
nor NOR3 (N1105, N1094, N391, N344);
or OR2 (N1106, N1103, N968);
buf BUF1 (N1107, N1104);
xor XOR2 (N1108, N1106, N983);
and AND3 (N1109, N1085, N864, N1105);
xor XOR2 (N1110, N439, N845);
xor XOR2 (N1111, N1100, N637);
or OR3 (N1112, N1102, N860, N115);
buf BUF1 (N1113, N1109);
or OR2 (N1114, N1113, N843);
nand NAND4 (N1115, N1095, N210, N445, N505);
buf BUF1 (N1116, N1092);
nor NOR4 (N1117, N1112, N968, N309, N65);
or OR4 (N1118, N1101, N1115, N1100, N990);
or OR2 (N1119, N78, N644);
nand NAND2 (N1120, N1088, N1074);
nor NOR2 (N1121, N1108, N1016);
or OR4 (N1122, N1119, N938, N644, N266);
not NOT1 (N1123, N1117);
nor NOR3 (N1124, N1107, N814, N345);
and AND2 (N1125, N1123, N513);
and AND4 (N1126, N1121, N922, N86, N964);
xor XOR2 (N1127, N1110, N131);
buf BUF1 (N1128, N1120);
xor XOR2 (N1129, N1114, N491);
buf BUF1 (N1130, N1118);
xor XOR2 (N1131, N1129, N893);
not NOT1 (N1132, N1111);
nor NOR2 (N1133, N1122, N88);
or OR3 (N1134, N1116, N425, N595);
xor XOR2 (N1135, N1133, N225);
and AND3 (N1136, N1127, N381, N658);
nand NAND2 (N1137, N1128, N749);
not NOT1 (N1138, N1125);
xor XOR2 (N1139, N1134, N942);
xor XOR2 (N1140, N1131, N630);
nor NOR4 (N1141, N1124, N1064, N518, N998);
and AND2 (N1142, N1141, N164);
not NOT1 (N1143, N1139);
not NOT1 (N1144, N1136);
xor XOR2 (N1145, N1137, N960);
not NOT1 (N1146, N1135);
nand NAND4 (N1147, N1126, N437, N92, N931);
nand NAND3 (N1148, N1145, N804, N927);
nand NAND4 (N1149, N1140, N41, N831, N67);
or OR3 (N1150, N1143, N541, N310);
nor NOR2 (N1151, N1146, N571);
or OR4 (N1152, N1138, N911, N280, N1044);
or OR4 (N1153, N1152, N1129, N960, N377);
nand NAND4 (N1154, N1142, N55, N200, N570);
xor XOR2 (N1155, N1144, N7);
nand NAND2 (N1156, N1132, N975);
and AND3 (N1157, N1151, N210, N734);
nand NAND2 (N1158, N1130, N508);
xor XOR2 (N1159, N1147, N857);
nand NAND3 (N1160, N1158, N105, N660);
buf BUF1 (N1161, N1159);
and AND3 (N1162, N1148, N770, N779);
and AND2 (N1163, N1157, N380);
or OR2 (N1164, N1156, N169);
and AND4 (N1165, N1161, N292, N635, N1117);
xor XOR2 (N1166, N1149, N558);
xor XOR2 (N1167, N1150, N998);
xor XOR2 (N1168, N1163, N862);
nor NOR2 (N1169, N1164, N1039);
nor NOR4 (N1170, N1166, N13, N38, N427);
not NOT1 (N1171, N1169);
xor XOR2 (N1172, N1155, N286);
nand NAND4 (N1173, N1154, N104, N875, N246);
and AND2 (N1174, N1167, N263);
or OR2 (N1175, N1173, N499);
and AND3 (N1176, N1171, N932, N923);
not NOT1 (N1177, N1168);
and AND2 (N1178, N1165, N781);
buf BUF1 (N1179, N1177);
nand NAND2 (N1180, N1170, N102);
nor NOR3 (N1181, N1178, N408, N10);
not NOT1 (N1182, N1172);
not NOT1 (N1183, N1179);
nand NAND2 (N1184, N1175, N4);
buf BUF1 (N1185, N1183);
xor XOR2 (N1186, N1162, N673);
xor XOR2 (N1187, N1180, N773);
nand NAND2 (N1188, N1176, N692);
buf BUF1 (N1189, N1186);
not NOT1 (N1190, N1160);
buf BUF1 (N1191, N1184);
not NOT1 (N1192, N1191);
and AND4 (N1193, N1187, N480, N456, N591);
xor XOR2 (N1194, N1181, N446);
nand NAND4 (N1195, N1185, N931, N602, N711);
buf BUF1 (N1196, N1194);
nand NAND2 (N1197, N1192, N194);
or OR4 (N1198, N1189, N1092, N399, N853);
or OR3 (N1199, N1190, N734, N288);
nor NOR4 (N1200, N1193, N1104, N848, N609);
nor NOR4 (N1201, N1200, N77, N231, N844);
nand NAND3 (N1202, N1182, N232, N683);
and AND4 (N1203, N1153, N10, N899, N423);
nor NOR3 (N1204, N1196, N429, N1176);
buf BUF1 (N1205, N1203);
or OR4 (N1206, N1195, N1195, N581, N664);
nand NAND2 (N1207, N1206, N769);
and AND4 (N1208, N1199, N1182, N500, N935);
buf BUF1 (N1209, N1204);
xor XOR2 (N1210, N1209, N646);
xor XOR2 (N1211, N1198, N542);
and AND4 (N1212, N1201, N1138, N565, N472);
nand NAND3 (N1213, N1188, N1035, N118);
nand NAND4 (N1214, N1174, N63, N1015, N971);
nand NAND4 (N1215, N1202, N74, N72, N899);
and AND4 (N1216, N1215, N740, N538, N1136);
nand NAND3 (N1217, N1205, N104, N1100);
xor XOR2 (N1218, N1210, N336);
nand NAND3 (N1219, N1217, N1048, N194);
xor XOR2 (N1220, N1213, N907);
buf BUF1 (N1221, N1220);
xor XOR2 (N1222, N1208, N1106);
nor NOR4 (N1223, N1212, N641, N200, N385);
not NOT1 (N1224, N1223);
nor NOR4 (N1225, N1216, N104, N107, N213);
xor XOR2 (N1226, N1214, N767);
and AND2 (N1227, N1197, N752);
and AND3 (N1228, N1211, N668, N297);
and AND4 (N1229, N1227, N643, N1043, N421);
xor XOR2 (N1230, N1226, N894);
buf BUF1 (N1231, N1221);
xor XOR2 (N1232, N1225, N721);
xor XOR2 (N1233, N1230, N1021);
nor NOR3 (N1234, N1219, N513, N587);
nor NOR4 (N1235, N1234, N1161, N302, N685);
and AND4 (N1236, N1222, N343, N631, N609);
not NOT1 (N1237, N1232);
or OR3 (N1238, N1224, N463, N887);
buf BUF1 (N1239, N1233);
xor XOR2 (N1240, N1228, N748);
nor NOR3 (N1241, N1239, N625, N72);
or OR4 (N1242, N1241, N360, N799, N262);
buf BUF1 (N1243, N1242);
nor NOR4 (N1244, N1207, N1109, N1195, N475);
nor NOR2 (N1245, N1235, N222);
buf BUF1 (N1246, N1243);
nand NAND2 (N1247, N1244, N271);
not NOT1 (N1248, N1237);
buf BUF1 (N1249, N1229);
or OR3 (N1250, N1249, N358, N385);
nand NAND4 (N1251, N1248, N199, N1144, N418);
or OR3 (N1252, N1218, N662, N1247);
nand NAND4 (N1253, N647, N227, N508, N748);
and AND3 (N1254, N1245, N271, N676);
and AND3 (N1255, N1251, N503, N683);
nor NOR3 (N1256, N1250, N1193, N1165);
xor XOR2 (N1257, N1252, N322);
buf BUF1 (N1258, N1231);
buf BUF1 (N1259, N1258);
nand NAND3 (N1260, N1259, N538, N257);
not NOT1 (N1261, N1257);
or OR2 (N1262, N1254, N123);
and AND3 (N1263, N1236, N535, N485);
or OR3 (N1264, N1262, N1234, N498);
or OR4 (N1265, N1240, N993, N1036, N311);
nand NAND2 (N1266, N1260, N93);
not NOT1 (N1267, N1256);
buf BUF1 (N1268, N1265);
nand NAND2 (N1269, N1238, N531);
and AND2 (N1270, N1246, N1206);
not NOT1 (N1271, N1264);
xor XOR2 (N1272, N1263, N384);
xor XOR2 (N1273, N1269, N260);
buf BUF1 (N1274, N1271);
or OR3 (N1275, N1273, N2, N439);
nand NAND2 (N1276, N1266, N803);
nor NOR3 (N1277, N1275, N1127, N6);
nand NAND3 (N1278, N1276, N272, N804);
nor NOR2 (N1279, N1270, N1115);
or OR4 (N1280, N1278, N84, N250, N996);
not NOT1 (N1281, N1279);
xor XOR2 (N1282, N1277, N923);
or OR2 (N1283, N1281, N166);
not NOT1 (N1284, N1253);
xor XOR2 (N1285, N1255, N725);
and AND4 (N1286, N1274, N404, N1189, N948);
xor XOR2 (N1287, N1261, N1009);
buf BUF1 (N1288, N1287);
and AND4 (N1289, N1272, N371, N559, N30);
buf BUF1 (N1290, N1267);
nor NOR4 (N1291, N1283, N369, N340, N839);
nand NAND3 (N1292, N1285, N1126, N825);
nand NAND2 (N1293, N1284, N1094);
nand NAND3 (N1294, N1282, N589, N996);
and AND4 (N1295, N1268, N282, N533, N1278);
or OR2 (N1296, N1290, N597);
and AND2 (N1297, N1294, N1058);
and AND3 (N1298, N1292, N332, N1222);
or OR2 (N1299, N1289, N783);
buf BUF1 (N1300, N1296);
nand NAND2 (N1301, N1286, N1065);
or OR3 (N1302, N1299, N43, N510);
and AND2 (N1303, N1300, N605);
and AND2 (N1304, N1302, N63);
or OR3 (N1305, N1291, N88, N418);
or OR2 (N1306, N1301, N141);
nand NAND4 (N1307, N1305, N1118, N833, N999);
nor NOR2 (N1308, N1297, N580);
nand NAND2 (N1309, N1308, N1025);
xor XOR2 (N1310, N1304, N81);
buf BUF1 (N1311, N1306);
nor NOR2 (N1312, N1280, N937);
or OR4 (N1313, N1288, N1104, N192, N301);
nor NOR2 (N1314, N1298, N513);
not NOT1 (N1315, N1307);
or OR4 (N1316, N1315, N622, N737, N450);
and AND4 (N1317, N1295, N179, N740, N964);
xor XOR2 (N1318, N1313, N1207);
xor XOR2 (N1319, N1314, N794);
xor XOR2 (N1320, N1318, N14);
nor NOR3 (N1321, N1303, N638, N912);
and AND4 (N1322, N1317, N1097, N420, N513);
xor XOR2 (N1323, N1309, N130);
xor XOR2 (N1324, N1311, N983);
not NOT1 (N1325, N1320);
nand NAND2 (N1326, N1293, N1153);
buf BUF1 (N1327, N1321);
buf BUF1 (N1328, N1316);
or OR3 (N1329, N1312, N62, N869);
not NOT1 (N1330, N1310);
nand NAND3 (N1331, N1327, N720, N723);
xor XOR2 (N1332, N1329, N205);
and AND4 (N1333, N1332, N1120, N1182, N1234);
buf BUF1 (N1334, N1330);
or OR3 (N1335, N1331, N200, N688);
buf BUF1 (N1336, N1323);
buf BUF1 (N1337, N1322);
or OR2 (N1338, N1319, N451);
xor XOR2 (N1339, N1324, N772);
not NOT1 (N1340, N1334);
nand NAND4 (N1341, N1335, N49, N17, N1338);
xor XOR2 (N1342, N1006, N296);
or OR3 (N1343, N1341, N1140, N303);
nor NOR2 (N1344, N1326, N570);
and AND4 (N1345, N1340, N146, N574, N342);
xor XOR2 (N1346, N1339, N975);
nor NOR3 (N1347, N1345, N482, N913);
xor XOR2 (N1348, N1346, N78);
or OR3 (N1349, N1333, N430, N390);
or OR4 (N1350, N1348, N103, N565, N544);
nand NAND3 (N1351, N1344, N1041, N260);
nor NOR3 (N1352, N1342, N1221, N602);
nand NAND3 (N1353, N1328, N520, N54);
xor XOR2 (N1354, N1353, N898);
and AND4 (N1355, N1337, N1234, N597, N163);
xor XOR2 (N1356, N1352, N444);
xor XOR2 (N1357, N1347, N12);
nand NAND4 (N1358, N1349, N834, N960, N487);
xor XOR2 (N1359, N1358, N644);
nor NOR3 (N1360, N1336, N1088, N381);
or OR2 (N1361, N1351, N139);
or OR2 (N1362, N1355, N1266);
and AND3 (N1363, N1325, N1291, N875);
nor NOR3 (N1364, N1357, N586, N511);
and AND2 (N1365, N1362, N1019);
nand NAND4 (N1366, N1350, N1351, N687, N517);
xor XOR2 (N1367, N1363, N508);
buf BUF1 (N1368, N1361);
not NOT1 (N1369, N1359);
or OR3 (N1370, N1369, N248, N1273);
buf BUF1 (N1371, N1360);
nand NAND3 (N1372, N1371, N283, N1121);
or OR4 (N1373, N1365, N575, N109, N453);
buf BUF1 (N1374, N1366);
and AND4 (N1375, N1356, N1015, N1008, N1097);
xor XOR2 (N1376, N1375, N1179);
not NOT1 (N1377, N1370);
not NOT1 (N1378, N1372);
nor NOR3 (N1379, N1377, N1067, N922);
or OR4 (N1380, N1373, N671, N1095, N328);
not NOT1 (N1381, N1378);
and AND4 (N1382, N1381, N458, N1184, N595);
buf BUF1 (N1383, N1354);
nand NAND2 (N1384, N1379, N376);
nand NAND4 (N1385, N1383, N650, N82, N1355);
nand NAND4 (N1386, N1367, N1288, N452, N954);
xor XOR2 (N1387, N1386, N1346);
not NOT1 (N1388, N1376);
not NOT1 (N1389, N1374);
nand NAND4 (N1390, N1343, N167, N734, N644);
nand NAND3 (N1391, N1368, N712, N968);
buf BUF1 (N1392, N1382);
or OR2 (N1393, N1389, N1111);
and AND2 (N1394, N1384, N1091);
buf BUF1 (N1395, N1387);
nand NAND3 (N1396, N1391, N1200, N1060);
nor NOR2 (N1397, N1388, N1130);
and AND4 (N1398, N1392, N1146, N1115, N1140);
xor XOR2 (N1399, N1398, N965);
nand NAND3 (N1400, N1397, N158, N1122);
nand NAND3 (N1401, N1400, N67, N797);
and AND2 (N1402, N1394, N922);
or OR3 (N1403, N1395, N580, N1283);
buf BUF1 (N1404, N1393);
or OR2 (N1405, N1399, N149);
nor NOR2 (N1406, N1364, N861);
or OR4 (N1407, N1396, N1364, N1399, N485);
buf BUF1 (N1408, N1404);
not NOT1 (N1409, N1390);
nand NAND4 (N1410, N1385, N473, N347, N198);
not NOT1 (N1411, N1409);
buf BUF1 (N1412, N1406);
not NOT1 (N1413, N1412);
or OR3 (N1414, N1407, N28, N352);
not NOT1 (N1415, N1401);
not NOT1 (N1416, N1403);
nor NOR3 (N1417, N1416, N1231, N916);
xor XOR2 (N1418, N1380, N402);
nand NAND4 (N1419, N1418, N1409, N972, N235);
nand NAND3 (N1420, N1408, N254, N841);
buf BUF1 (N1421, N1402);
nor NOR2 (N1422, N1415, N623);
nor NOR4 (N1423, N1419, N350, N947, N1094);
xor XOR2 (N1424, N1413, N329);
and AND4 (N1425, N1414, N1228, N752, N345);
or OR2 (N1426, N1420, N1174);
or OR3 (N1427, N1425, N955, N441);
xor XOR2 (N1428, N1421, N808);
xor XOR2 (N1429, N1411, N122);
or OR3 (N1430, N1423, N386, N25);
nand NAND3 (N1431, N1422, N1233, N776);
not NOT1 (N1432, N1417);
nor NOR4 (N1433, N1428, N207, N851, N503);
or OR2 (N1434, N1429, N407);
and AND4 (N1435, N1433, N988, N396, N422);
or OR4 (N1436, N1426, N636, N1269, N66);
nor NOR2 (N1437, N1432, N59);
and AND2 (N1438, N1405, N801);
or OR3 (N1439, N1410, N1300, N532);
buf BUF1 (N1440, N1431);
nor NOR2 (N1441, N1439, N76);
not NOT1 (N1442, N1436);
xor XOR2 (N1443, N1430, N380);
not NOT1 (N1444, N1437);
not NOT1 (N1445, N1441);
nor NOR3 (N1446, N1434, N624, N716);
not NOT1 (N1447, N1444);
not NOT1 (N1448, N1427);
or OR4 (N1449, N1446, N240, N645, N81);
not NOT1 (N1450, N1438);
nand NAND3 (N1451, N1440, N570, N641);
xor XOR2 (N1452, N1445, N1083);
nor NOR4 (N1453, N1452, N90, N872, N125);
and AND4 (N1454, N1448, N332, N716, N909);
nor NOR3 (N1455, N1443, N772, N1240);
or OR3 (N1456, N1424, N1382, N419);
xor XOR2 (N1457, N1435, N413);
and AND2 (N1458, N1447, N498);
and AND3 (N1459, N1450, N276, N698);
or OR2 (N1460, N1451, N1455);
nor NOR2 (N1461, N322, N239);
or OR3 (N1462, N1454, N128, N1268);
and AND3 (N1463, N1449, N1260, N1321);
or OR4 (N1464, N1463, N650, N940, N353);
or OR4 (N1465, N1462, N49, N1389, N450);
and AND3 (N1466, N1461, N1355, N176);
nor NOR2 (N1467, N1456, N385);
xor XOR2 (N1468, N1442, N1271);
or OR2 (N1469, N1457, N317);
nor NOR3 (N1470, N1464, N635, N1458);
or OR4 (N1471, N403, N855, N60, N1429);
xor XOR2 (N1472, N1470, N540);
xor XOR2 (N1473, N1453, N270);
xor XOR2 (N1474, N1473, N1090);
buf BUF1 (N1475, N1469);
nor NOR4 (N1476, N1474, N754, N986, N788);
xor XOR2 (N1477, N1465, N362);
xor XOR2 (N1478, N1466, N1256);
not NOT1 (N1479, N1476);
and AND4 (N1480, N1459, N466, N611, N460);
nor NOR2 (N1481, N1467, N871);
and AND2 (N1482, N1475, N342);
or OR4 (N1483, N1471, N355, N174, N934);
or OR2 (N1484, N1482, N1059);
nor NOR3 (N1485, N1479, N701, N998);
and AND4 (N1486, N1481, N389, N937, N22);
nand NAND4 (N1487, N1477, N1405, N765, N929);
buf BUF1 (N1488, N1472);
nor NOR4 (N1489, N1487, N946, N909, N563);
nor NOR3 (N1490, N1483, N1211, N598);
and AND4 (N1491, N1490, N84, N670, N1038);
not NOT1 (N1492, N1484);
xor XOR2 (N1493, N1485, N1061);
or OR3 (N1494, N1486, N1122, N1149);
nor NOR2 (N1495, N1488, N513);
xor XOR2 (N1496, N1493, N972);
xor XOR2 (N1497, N1468, N774);
not NOT1 (N1498, N1491);
or OR4 (N1499, N1495, N92, N1414, N889);
xor XOR2 (N1500, N1498, N799);
nand NAND3 (N1501, N1492, N352, N920);
and AND4 (N1502, N1501, N753, N853, N822);
or OR4 (N1503, N1460, N1042, N133, N215);
and AND3 (N1504, N1494, N1404, N343);
or OR3 (N1505, N1497, N906, N441);
and AND2 (N1506, N1489, N1200);
nand NAND3 (N1507, N1480, N1051, N987);
and AND3 (N1508, N1478, N20, N956);
and AND3 (N1509, N1502, N1383, N293);
nand NAND4 (N1510, N1500, N1488, N48, N1461);
nor NOR3 (N1511, N1507, N1093, N651);
xor XOR2 (N1512, N1496, N1081);
and AND3 (N1513, N1503, N805, N1208);
nand NAND4 (N1514, N1512, N887, N1197, N1466);
xor XOR2 (N1515, N1508, N1389);
nand NAND3 (N1516, N1504, N176, N1103);
nand NAND3 (N1517, N1505, N274, N1436);
xor XOR2 (N1518, N1514, N77);
nor NOR2 (N1519, N1506, N1366);
and AND2 (N1520, N1509, N420);
and AND3 (N1521, N1516, N449, N422);
xor XOR2 (N1522, N1499, N569);
xor XOR2 (N1523, N1519, N294);
nor NOR4 (N1524, N1521, N1189, N648, N467);
and AND4 (N1525, N1513, N1178, N305, N290);
or OR3 (N1526, N1522, N1229, N819);
buf BUF1 (N1527, N1525);
xor XOR2 (N1528, N1511, N726);
nor NOR3 (N1529, N1518, N1122, N1049);
not NOT1 (N1530, N1528);
or OR3 (N1531, N1515, N485, N138);
or OR4 (N1532, N1531, N329, N723, N610);
nor NOR4 (N1533, N1520, N264, N900, N484);
xor XOR2 (N1534, N1530, N707);
nand NAND3 (N1535, N1532, N1428, N1045);
nor NOR2 (N1536, N1533, N971);
buf BUF1 (N1537, N1527);
buf BUF1 (N1538, N1529);
xor XOR2 (N1539, N1535, N1058);
or OR2 (N1540, N1539, N236);
or OR4 (N1541, N1510, N84, N386, N101);
buf BUF1 (N1542, N1534);
not NOT1 (N1543, N1541);
or OR4 (N1544, N1542, N741, N613, N1204);
xor XOR2 (N1545, N1517, N93);
nand NAND4 (N1546, N1538, N262, N282, N738);
nand NAND3 (N1547, N1540, N1434, N1523);
nor NOR3 (N1548, N338, N40, N58);
or OR3 (N1549, N1547, N1205, N961);
xor XOR2 (N1550, N1537, N1108);
buf BUF1 (N1551, N1524);
nor NOR4 (N1552, N1546, N51, N250, N63);
not NOT1 (N1553, N1548);
xor XOR2 (N1554, N1526, N507);
nor NOR3 (N1555, N1552, N774, N154);
buf BUF1 (N1556, N1544);
not NOT1 (N1557, N1553);
xor XOR2 (N1558, N1555, N1288);
and AND2 (N1559, N1554, N401);
buf BUF1 (N1560, N1545);
nor NOR3 (N1561, N1557, N482, N133);
nand NAND4 (N1562, N1549, N16, N1290, N365);
xor XOR2 (N1563, N1559, N1136);
nor NOR2 (N1564, N1543, N775);
xor XOR2 (N1565, N1558, N968);
nor NOR2 (N1566, N1551, N505);
nand NAND2 (N1567, N1536, N1129);
or OR4 (N1568, N1562, N537, N154, N1095);
or OR3 (N1569, N1550, N1503, N434);
or OR2 (N1570, N1563, N1396);
or OR3 (N1571, N1556, N1443, N1181);
nor NOR3 (N1572, N1569, N227, N907);
and AND4 (N1573, N1566, N707, N692, N945);
nand NAND3 (N1574, N1572, N1463, N837);
buf BUF1 (N1575, N1571);
and AND3 (N1576, N1568, N967, N681);
nand NAND3 (N1577, N1565, N1290, N291);
and AND3 (N1578, N1567, N579, N1150);
nor NOR2 (N1579, N1561, N398);
and AND2 (N1580, N1570, N180);
not NOT1 (N1581, N1573);
buf BUF1 (N1582, N1577);
or OR2 (N1583, N1580, N693);
or OR3 (N1584, N1560, N636, N151);
nand NAND2 (N1585, N1582, N1354);
or OR2 (N1586, N1584, N1318);
or OR4 (N1587, N1574, N1195, N1261, N682);
and AND4 (N1588, N1575, N604, N553, N1462);
nor NOR3 (N1589, N1564, N1022, N857);
nor NOR4 (N1590, N1581, N95, N1169, N1418);
nand NAND2 (N1591, N1579, N715);
or OR4 (N1592, N1585, N502, N557, N1478);
and AND2 (N1593, N1588, N753);
not NOT1 (N1594, N1593);
nor NOR4 (N1595, N1586, N923, N1542, N1093);
buf BUF1 (N1596, N1587);
nand NAND3 (N1597, N1594, N372, N1498);
buf BUF1 (N1598, N1589);
not NOT1 (N1599, N1598);
or OR4 (N1600, N1590, N1544, N744, N194);
not NOT1 (N1601, N1597);
buf BUF1 (N1602, N1599);
not NOT1 (N1603, N1600);
and AND4 (N1604, N1591, N182, N539, N176);
buf BUF1 (N1605, N1601);
or OR4 (N1606, N1583, N1265, N1087, N1106);
xor XOR2 (N1607, N1576, N797);
and AND4 (N1608, N1592, N507, N664, N405);
and AND2 (N1609, N1604, N441);
not NOT1 (N1610, N1602);
not NOT1 (N1611, N1608);
xor XOR2 (N1612, N1610, N130);
and AND2 (N1613, N1606, N194);
buf BUF1 (N1614, N1613);
xor XOR2 (N1615, N1603, N175);
nand NAND3 (N1616, N1595, N81, N10);
or OR3 (N1617, N1615, N437, N252);
nor NOR3 (N1618, N1614, N216, N384);
buf BUF1 (N1619, N1611);
nand NAND3 (N1620, N1619, N1405, N581);
xor XOR2 (N1621, N1617, N160);
xor XOR2 (N1622, N1607, N31);
nand NAND2 (N1623, N1609, N584);
xor XOR2 (N1624, N1620, N325);
or OR4 (N1625, N1622, N1076, N686, N767);
buf BUF1 (N1626, N1612);
nand NAND3 (N1627, N1596, N1513, N1199);
and AND2 (N1628, N1616, N603);
or OR3 (N1629, N1627, N1277, N150);
nand NAND2 (N1630, N1618, N131);
nor NOR2 (N1631, N1625, N1136);
nor NOR2 (N1632, N1629, N432);
not NOT1 (N1633, N1631);
xor XOR2 (N1634, N1578, N245);
buf BUF1 (N1635, N1630);
nor NOR3 (N1636, N1634, N1271, N874);
nor NOR2 (N1637, N1621, N53);
or OR2 (N1638, N1633, N870);
nand NAND2 (N1639, N1626, N694);
xor XOR2 (N1640, N1632, N24);
xor XOR2 (N1641, N1628, N1115);
and AND2 (N1642, N1623, N1633);
xor XOR2 (N1643, N1636, N938);
buf BUF1 (N1644, N1638);
not NOT1 (N1645, N1644);
or OR4 (N1646, N1637, N485, N15, N1278);
nand NAND3 (N1647, N1642, N39, N1002);
and AND4 (N1648, N1605, N802, N1335, N91);
buf BUF1 (N1649, N1647);
nand NAND4 (N1650, N1640, N1570, N195, N495);
or OR2 (N1651, N1645, N1591);
not NOT1 (N1652, N1650);
or OR2 (N1653, N1624, N1420);
nor NOR4 (N1654, N1653, N1541, N601, N1304);
buf BUF1 (N1655, N1652);
buf BUF1 (N1656, N1641);
buf BUF1 (N1657, N1651);
xor XOR2 (N1658, N1639, N138);
or OR2 (N1659, N1635, N898);
or OR3 (N1660, N1655, N527, N87);
not NOT1 (N1661, N1660);
nor NOR4 (N1662, N1656, N1197, N15, N1362);
and AND4 (N1663, N1646, N29, N108, N560);
buf BUF1 (N1664, N1661);
not NOT1 (N1665, N1648);
buf BUF1 (N1666, N1665);
nand NAND2 (N1667, N1664, N585);
nor NOR2 (N1668, N1667, N1131);
and AND3 (N1669, N1666, N1665, N42);
and AND3 (N1670, N1654, N421, N76);
nor NOR3 (N1671, N1663, N1411, N218);
nand NAND4 (N1672, N1668, N320, N578, N1276);
buf BUF1 (N1673, N1658);
nand NAND4 (N1674, N1671, N1061, N90, N657);
nand NAND2 (N1675, N1674, N1258);
or OR4 (N1676, N1673, N1592, N1393, N1050);
buf BUF1 (N1677, N1669);
xor XOR2 (N1678, N1643, N464);
and AND2 (N1679, N1675, N503);
nor NOR3 (N1680, N1678, N854, N920);
and AND2 (N1681, N1662, N1638);
nor NOR4 (N1682, N1680, N180, N1067, N710);
nand NAND2 (N1683, N1677, N1307);
nor NOR2 (N1684, N1679, N1609);
buf BUF1 (N1685, N1684);
nand NAND4 (N1686, N1681, N303, N825, N1490);
and AND2 (N1687, N1649, N1450);
nand NAND2 (N1688, N1670, N1407);
buf BUF1 (N1689, N1657);
and AND4 (N1690, N1672, N1134, N342, N1349);
xor XOR2 (N1691, N1686, N1175);
or OR3 (N1692, N1687, N1590, N500);
or OR3 (N1693, N1659, N561, N1303);
nand NAND4 (N1694, N1692, N1330, N1692, N569);
nor NOR4 (N1695, N1683, N686, N178, N864);
nor NOR4 (N1696, N1694, N1175, N1388, N655);
nand NAND4 (N1697, N1693, N1309, N414, N383);
nor NOR2 (N1698, N1688, N1304);
or OR4 (N1699, N1697, N252, N1696, N259);
nor NOR3 (N1700, N1653, N863, N1692);
xor XOR2 (N1701, N1685, N427);
not NOT1 (N1702, N1689);
or OR2 (N1703, N1702, N599);
buf BUF1 (N1704, N1691);
not NOT1 (N1705, N1698);
nand NAND4 (N1706, N1695, N1438, N689, N1238);
not NOT1 (N1707, N1690);
nand NAND3 (N1708, N1703, N564, N1518);
xor XOR2 (N1709, N1701, N472);
nand NAND3 (N1710, N1707, N211, N6);
not NOT1 (N1711, N1708);
nand NAND3 (N1712, N1706, N169, N90);
buf BUF1 (N1713, N1705);
buf BUF1 (N1714, N1712);
nand NAND2 (N1715, N1676, N1427);
xor XOR2 (N1716, N1713, N218);
not NOT1 (N1717, N1682);
nor NOR4 (N1718, N1715, N851, N159, N187);
buf BUF1 (N1719, N1700);
buf BUF1 (N1720, N1714);
nor NOR2 (N1721, N1710, N184);
or OR2 (N1722, N1717, N103);
and AND4 (N1723, N1711, N364, N1711, N160);
buf BUF1 (N1724, N1722);
not NOT1 (N1725, N1716);
buf BUF1 (N1726, N1721);
not NOT1 (N1727, N1720);
nor NOR3 (N1728, N1709, N1082, N191);
and AND4 (N1729, N1699, N448, N1018, N702);
not NOT1 (N1730, N1725);
buf BUF1 (N1731, N1719);
not NOT1 (N1732, N1704);
xor XOR2 (N1733, N1727, N1719);
and AND2 (N1734, N1730, N1348);
xor XOR2 (N1735, N1732, N343);
nand NAND3 (N1736, N1734, N249, N872);
nand NAND3 (N1737, N1736, N1475, N363);
nand NAND4 (N1738, N1718, N262, N1594, N1194);
nor NOR4 (N1739, N1737, N1406, N935, N76);
nand NAND3 (N1740, N1731, N283, N936);
nand NAND2 (N1741, N1723, N1044);
not NOT1 (N1742, N1740);
buf BUF1 (N1743, N1729);
buf BUF1 (N1744, N1742);
buf BUF1 (N1745, N1726);
and AND3 (N1746, N1741, N254, N1425);
not NOT1 (N1747, N1724);
nand NAND4 (N1748, N1745, N1679, N1490, N907);
not NOT1 (N1749, N1744);
xor XOR2 (N1750, N1746, N1707);
not NOT1 (N1751, N1743);
buf BUF1 (N1752, N1748);
buf BUF1 (N1753, N1735);
and AND2 (N1754, N1751, N679);
and AND2 (N1755, N1738, N1262);
buf BUF1 (N1756, N1749);
nor NOR2 (N1757, N1754, N391);
and AND4 (N1758, N1752, N135, N1444, N718);
nand NAND3 (N1759, N1728, N1754, N397);
or OR2 (N1760, N1739, N1432);
xor XOR2 (N1761, N1756, N311);
and AND3 (N1762, N1761, N1282, N1043);
not NOT1 (N1763, N1760);
and AND2 (N1764, N1763, N1606);
or OR2 (N1765, N1758, N304);
and AND2 (N1766, N1755, N934);
and AND3 (N1767, N1766, N359, N988);
buf BUF1 (N1768, N1762);
xor XOR2 (N1769, N1757, N676);
nor NOR3 (N1770, N1769, N1097, N1413);
or OR4 (N1771, N1768, N867, N90, N1582);
or OR3 (N1772, N1764, N339, N418);
nor NOR2 (N1773, N1771, N1073);
not NOT1 (N1774, N1772);
xor XOR2 (N1775, N1765, N981);
nand NAND3 (N1776, N1773, N1620, N626);
buf BUF1 (N1777, N1733);
nand NAND4 (N1778, N1775, N1215, N1213, N1130);
xor XOR2 (N1779, N1747, N241);
buf BUF1 (N1780, N1779);
not NOT1 (N1781, N1753);
and AND4 (N1782, N1759, N512, N1342, N504);
xor XOR2 (N1783, N1770, N1089);
nor NOR4 (N1784, N1781, N1487, N673, N1649);
xor XOR2 (N1785, N1776, N1418);
or OR3 (N1786, N1784, N710, N1228);
nor NOR3 (N1787, N1778, N674, N730);
and AND3 (N1788, N1767, N134, N1340);
or OR2 (N1789, N1750, N1646);
nand NAND3 (N1790, N1783, N396, N1580);
nand NAND2 (N1791, N1786, N1372);
buf BUF1 (N1792, N1785);
not NOT1 (N1793, N1787);
nor NOR2 (N1794, N1774, N1014);
xor XOR2 (N1795, N1793, N754);
buf BUF1 (N1796, N1790);
buf BUF1 (N1797, N1780);
not NOT1 (N1798, N1795);
buf BUF1 (N1799, N1777);
not NOT1 (N1800, N1794);
nand NAND3 (N1801, N1782, N180, N241);
xor XOR2 (N1802, N1799, N473);
xor XOR2 (N1803, N1789, N253);
buf BUF1 (N1804, N1800);
buf BUF1 (N1805, N1791);
buf BUF1 (N1806, N1797);
and AND4 (N1807, N1798, N1429, N1147, N1281);
not NOT1 (N1808, N1806);
nor NOR2 (N1809, N1805, N1673);
xor XOR2 (N1810, N1807, N338);
nand NAND4 (N1811, N1803, N1017, N191, N572);
nor NOR3 (N1812, N1788, N908, N1127);
xor XOR2 (N1813, N1804, N998);
xor XOR2 (N1814, N1811, N11);
and AND4 (N1815, N1796, N555, N41, N395);
or OR4 (N1816, N1813, N168, N1675, N746);
and AND2 (N1817, N1812, N503);
nor NOR2 (N1818, N1810, N1788);
not NOT1 (N1819, N1815);
not NOT1 (N1820, N1816);
nor NOR2 (N1821, N1809, N702);
nand NAND2 (N1822, N1821, N1757);
not NOT1 (N1823, N1819);
nor NOR4 (N1824, N1802, N48, N1100, N1360);
nand NAND3 (N1825, N1818, N1208, N1759);
or OR3 (N1826, N1817, N1276, N573);
nand NAND3 (N1827, N1825, N1179, N1555);
nor NOR3 (N1828, N1808, N1370, N1597);
xor XOR2 (N1829, N1792, N1533);
not NOT1 (N1830, N1824);
xor XOR2 (N1831, N1827, N1571);
nand NAND2 (N1832, N1820, N178);
nand NAND3 (N1833, N1828, N1685, N1030);
buf BUF1 (N1834, N1830);
and AND4 (N1835, N1834, N1444, N1684, N676);
or OR3 (N1836, N1822, N1075, N983);
buf BUF1 (N1837, N1801);
xor XOR2 (N1838, N1832, N1721);
xor XOR2 (N1839, N1838, N709);
and AND3 (N1840, N1836, N1588, N533);
nor NOR2 (N1841, N1826, N1167);
xor XOR2 (N1842, N1814, N196);
nand NAND2 (N1843, N1842, N851);
nor NOR2 (N1844, N1823, N1836);
or OR4 (N1845, N1840, N1459, N1794, N958);
nor NOR3 (N1846, N1845, N500, N415);
or OR2 (N1847, N1844, N1121);
xor XOR2 (N1848, N1843, N1043);
and AND4 (N1849, N1841, N1374, N699, N1694);
nor NOR2 (N1850, N1849, N1115);
buf BUF1 (N1851, N1829);
or OR4 (N1852, N1833, N68, N24, N751);
and AND2 (N1853, N1851, N113);
and AND3 (N1854, N1848, N1711, N1321);
or OR2 (N1855, N1853, N587);
and AND3 (N1856, N1852, N1461, N992);
xor XOR2 (N1857, N1850, N212);
and AND2 (N1858, N1846, N396);
and AND3 (N1859, N1854, N1581, N411);
buf BUF1 (N1860, N1859);
not NOT1 (N1861, N1839);
xor XOR2 (N1862, N1856, N325);
not NOT1 (N1863, N1835);
or OR2 (N1864, N1861, N345);
nand NAND3 (N1865, N1847, N927, N1778);
not NOT1 (N1866, N1857);
buf BUF1 (N1867, N1858);
or OR3 (N1868, N1860, N23, N548);
nor NOR4 (N1869, N1837, N992, N1335, N694);
xor XOR2 (N1870, N1867, N1309);
or OR4 (N1871, N1865, N1788, N1376, N1532);
nand NAND2 (N1872, N1864, N439);
and AND3 (N1873, N1863, N1267, N1192);
not NOT1 (N1874, N1871);
nand NAND2 (N1875, N1868, N1834);
xor XOR2 (N1876, N1862, N1802);
nor NOR3 (N1877, N1872, N1253, N1006);
and AND3 (N1878, N1869, N1365, N1369);
nand NAND2 (N1879, N1866, N780);
nand NAND4 (N1880, N1870, N431, N406, N769);
xor XOR2 (N1881, N1878, N1110);
nand NAND2 (N1882, N1875, N1685);
xor XOR2 (N1883, N1874, N721);
and AND4 (N1884, N1831, N1337, N831, N1608);
nand NAND2 (N1885, N1884, N930);
not NOT1 (N1886, N1876);
nor NOR3 (N1887, N1877, N1486, N567);
nor NOR2 (N1888, N1880, N373);
nand NAND3 (N1889, N1881, N1804, N853);
buf BUF1 (N1890, N1882);
not NOT1 (N1891, N1873);
or OR3 (N1892, N1879, N624, N48);
or OR3 (N1893, N1885, N248, N553);
or OR3 (N1894, N1889, N1023, N1242);
buf BUF1 (N1895, N1890);
or OR3 (N1896, N1887, N115, N1522);
xor XOR2 (N1897, N1891, N1342);
nor NOR4 (N1898, N1892, N1364, N1622, N1403);
xor XOR2 (N1899, N1883, N1636);
or OR4 (N1900, N1894, N327, N1646, N1584);
nor NOR2 (N1901, N1888, N388);
not NOT1 (N1902, N1895);
nor NOR2 (N1903, N1898, N1546);
nor NOR3 (N1904, N1900, N460, N681);
not NOT1 (N1905, N1886);
xor XOR2 (N1906, N1905, N1389);
xor XOR2 (N1907, N1901, N1460);
or OR4 (N1908, N1896, N1521, N1439, N1089);
or OR4 (N1909, N1893, N1741, N1561, N9);
xor XOR2 (N1910, N1909, N916);
nand NAND4 (N1911, N1908, N1493, N43, N609);
nor NOR4 (N1912, N1910, N831, N1150, N504);
or OR3 (N1913, N1907, N699, N1121);
nor NOR3 (N1914, N1906, N38, N548);
and AND4 (N1915, N1912, N331, N210, N1605);
and AND4 (N1916, N1899, N439, N939, N240);
not NOT1 (N1917, N1855);
and AND3 (N1918, N1917, N1008, N792);
buf BUF1 (N1919, N1911);
not NOT1 (N1920, N1919);
xor XOR2 (N1921, N1918, N678);
nor NOR3 (N1922, N1902, N565, N1086);
buf BUF1 (N1923, N1897);
not NOT1 (N1924, N1922);
nand NAND3 (N1925, N1924, N661, N343);
nand NAND4 (N1926, N1913, N933, N199, N1044);
xor XOR2 (N1927, N1914, N388);
not NOT1 (N1928, N1920);
and AND4 (N1929, N1925, N58, N717, N175);
not NOT1 (N1930, N1904);
nand NAND4 (N1931, N1929, N456, N269, N795);
or OR4 (N1932, N1923, N1510, N1084, N728);
nand NAND2 (N1933, N1921, N1504);
not NOT1 (N1934, N1926);
or OR2 (N1935, N1903, N1152);
not NOT1 (N1936, N1933);
or OR4 (N1937, N1935, N1251, N1089, N1090);
xor XOR2 (N1938, N1927, N852);
or OR2 (N1939, N1916, N1081);
or OR4 (N1940, N1938, N1059, N1129, N1446);
nand NAND4 (N1941, N1936, N1132, N671, N1193);
and AND2 (N1942, N1915, N1520);
nand NAND3 (N1943, N1939, N1319, N1441);
and AND3 (N1944, N1930, N1489, N1107);
buf BUF1 (N1945, N1937);
nor NOR2 (N1946, N1944, N561);
nor NOR4 (N1947, N1945, N743, N1146, N1112);
nand NAND4 (N1948, N1928, N1241, N1832, N196);
or OR4 (N1949, N1946, N1845, N1210, N268);
nand NAND2 (N1950, N1932, N1038);
not NOT1 (N1951, N1942);
and AND4 (N1952, N1940, N65, N21, N1364);
buf BUF1 (N1953, N1943);
nand NAND4 (N1954, N1951, N771, N1920, N289);
or OR2 (N1955, N1934, N1586);
nand NAND4 (N1956, N1941, N891, N171, N750);
nand NAND4 (N1957, N1948, N1669, N1642, N1181);
xor XOR2 (N1958, N1952, N1214);
and AND2 (N1959, N1958, N436);
nand NAND2 (N1960, N1959, N1946);
nand NAND3 (N1961, N1955, N1475, N1791);
xor XOR2 (N1962, N1953, N1907);
nand NAND2 (N1963, N1962, N1001);
buf BUF1 (N1964, N1956);
xor XOR2 (N1965, N1960, N271);
xor XOR2 (N1966, N1947, N1180);
nand NAND3 (N1967, N1950, N1857, N1136);
buf BUF1 (N1968, N1967);
or OR2 (N1969, N1957, N567);
nand NAND3 (N1970, N1968, N391, N880);
and AND3 (N1971, N1964, N1841, N1815);
buf BUF1 (N1972, N1966);
xor XOR2 (N1973, N1949, N1398);
not NOT1 (N1974, N1970);
nand NAND4 (N1975, N1973, N1579, N1969, N723);
nand NAND3 (N1976, N1286, N744, N1525);
buf BUF1 (N1977, N1976);
xor XOR2 (N1978, N1961, N1051);
xor XOR2 (N1979, N1954, N73);
nor NOR2 (N1980, N1977, N1665);
not NOT1 (N1981, N1971);
nand NAND3 (N1982, N1978, N1735, N1392);
or OR2 (N1983, N1974, N623);
and AND3 (N1984, N1983, N1505, N446);
not NOT1 (N1985, N1979);
nand NAND2 (N1986, N1980, N224);
and AND3 (N1987, N1985, N566, N399);
nand NAND2 (N1988, N1982, N1981);
nand NAND2 (N1989, N875, N1059);
buf BUF1 (N1990, N1986);
not NOT1 (N1991, N1988);
and AND2 (N1992, N1989, N691);
buf BUF1 (N1993, N1931);
xor XOR2 (N1994, N1984, N1347);
nand NAND4 (N1995, N1987, N402, N252, N1765);
nand NAND2 (N1996, N1992, N1170);
and AND3 (N1997, N1972, N488, N467);
buf BUF1 (N1998, N1990);
and AND4 (N1999, N1994, N1326, N980, N1089);
or OR2 (N2000, N1965, N1848);
not NOT1 (N2001, N1991);
xor XOR2 (N2002, N1975, N1271);
and AND3 (N2003, N1963, N1009, N534);
nand NAND4 (N2004, N1995, N1844, N1857, N433);
buf BUF1 (N2005, N2002);
xor XOR2 (N2006, N2004, N1801);
buf BUF1 (N2007, N1997);
nand NAND2 (N2008, N2007, N1708);
not NOT1 (N2009, N2005);
xor XOR2 (N2010, N2008, N1865);
and AND3 (N2011, N2003, N1604, N770);
buf BUF1 (N2012, N1996);
nor NOR4 (N2013, N2011, N256, N947, N1438);
nand NAND2 (N2014, N2000, N1451);
xor XOR2 (N2015, N2006, N312);
or OR4 (N2016, N2001, N1125, N1595, N644);
or OR2 (N2017, N2015, N1578);
xor XOR2 (N2018, N2010, N430);
buf BUF1 (N2019, N2018);
and AND2 (N2020, N1998, N1323);
and AND2 (N2021, N2013, N202);
nand NAND4 (N2022, N2021, N1877, N775, N767);
and AND4 (N2023, N1993, N760, N260, N267);
nand NAND4 (N2024, N2014, N946, N94, N1442);
xor XOR2 (N2025, N2019, N1316);
xor XOR2 (N2026, N2022, N460);
or OR2 (N2027, N2009, N653);
and AND3 (N2028, N2024, N687, N459);
not NOT1 (N2029, N2012);
nand NAND3 (N2030, N2025, N1502, N1664);
or OR2 (N2031, N2030, N89);
nor NOR2 (N2032, N2028, N740);
nor NOR4 (N2033, N2023, N704, N1312, N936);
nand NAND3 (N2034, N2033, N2005, N1213);
not NOT1 (N2035, N2016);
buf BUF1 (N2036, N2034);
and AND4 (N2037, N2026, N264, N269, N494);
nor NOR4 (N2038, N2036, N1152, N898, N1611);
nor NOR3 (N2039, N2029, N1368, N1575);
nor NOR2 (N2040, N2035, N470);
and AND2 (N2041, N2017, N1385);
nor NOR4 (N2042, N2039, N2006, N1609, N783);
or OR4 (N2043, N2032, N245, N987, N1736);
not NOT1 (N2044, N2027);
nor NOR3 (N2045, N2038, N460, N221);
and AND2 (N2046, N1999, N708);
not NOT1 (N2047, N2042);
and AND2 (N2048, N2045, N140);
xor XOR2 (N2049, N2043, N359);
nand NAND2 (N2050, N2020, N909);
or OR4 (N2051, N2046, N367, N1362, N1874);
nand NAND4 (N2052, N2047, N944, N771, N654);
nor NOR2 (N2053, N2048, N883);
and AND4 (N2054, N2044, N1762, N463, N1159);
nor NOR3 (N2055, N2051, N1313, N373);
or OR4 (N2056, N2055, N1150, N695, N955);
nand NAND4 (N2057, N2040, N1614, N1382, N1850);
buf BUF1 (N2058, N2054);
and AND2 (N2059, N2056, N78);
nand NAND4 (N2060, N2050, N1661, N261, N792);
and AND3 (N2061, N2057, N1694, N666);
buf BUF1 (N2062, N2060);
xor XOR2 (N2063, N2052, N558);
xor XOR2 (N2064, N2053, N91);
or OR2 (N2065, N2062, N1383);
not NOT1 (N2066, N2058);
buf BUF1 (N2067, N2041);
buf BUF1 (N2068, N2031);
nand NAND3 (N2069, N2067, N456, N1158);
buf BUF1 (N2070, N2064);
nand NAND2 (N2071, N2059, N1974);
buf BUF1 (N2072, N2065);
nand NAND4 (N2073, N2071, N1024, N1583, N977);
xor XOR2 (N2074, N2049, N974);
not NOT1 (N2075, N2037);
or OR3 (N2076, N2061, N1255, N761);
buf BUF1 (N2077, N2075);
or OR3 (N2078, N2076, N38, N1687);
or OR4 (N2079, N2078, N542, N1689, N964);
nor NOR2 (N2080, N2066, N1989);
or OR4 (N2081, N2069, N1711, N57, N2009);
nor NOR4 (N2082, N2063, N318, N1215, N1740);
buf BUF1 (N2083, N2072);
nor NOR3 (N2084, N2077, N1136, N543);
and AND3 (N2085, N2082, N1625, N1136);
buf BUF1 (N2086, N2083);
nand NAND3 (N2087, N2081, N2054, N1396);
buf BUF1 (N2088, N2074);
or OR4 (N2089, N2068, N647, N1067, N1261);
and AND2 (N2090, N2089, N976);
and AND2 (N2091, N2090, N493);
or OR3 (N2092, N2087, N482, N920);
nand NAND2 (N2093, N2079, N445);
nor NOR2 (N2094, N2070, N1113);
not NOT1 (N2095, N2091);
xor XOR2 (N2096, N2095, N102);
not NOT1 (N2097, N2084);
nand NAND4 (N2098, N2094, N683, N2094, N1759);
nor NOR3 (N2099, N2086, N677, N1912);
nand NAND4 (N2100, N2099, N471, N287, N127);
not NOT1 (N2101, N2098);
not NOT1 (N2102, N2080);
nor NOR3 (N2103, N2092, N47, N281);
and AND3 (N2104, N2102, N1786, N541);
or OR2 (N2105, N2096, N2097);
and AND2 (N2106, N569, N2011);
or OR4 (N2107, N2105, N1254, N1166, N1564);
buf BUF1 (N2108, N2093);
nor NOR4 (N2109, N2100, N1696, N1868, N1521);
and AND3 (N2110, N2101, N49, N1971);
nor NOR3 (N2111, N2103, N1689, N1433);
xor XOR2 (N2112, N2073, N184);
nand NAND2 (N2113, N2107, N73);
nand NAND3 (N2114, N2108, N1137, N460);
not NOT1 (N2115, N2085);
nand NAND4 (N2116, N2115, N392, N811, N1761);
nor NOR2 (N2117, N2109, N869);
nand NAND3 (N2118, N2112, N1561, N1228);
nor NOR3 (N2119, N2113, N733, N400);
buf BUF1 (N2120, N2110);
nand NAND2 (N2121, N2106, N2107);
or OR4 (N2122, N2116, N1596, N298, N716);
buf BUF1 (N2123, N2119);
xor XOR2 (N2124, N2104, N1078);
nand NAND2 (N2125, N2111, N1535);
xor XOR2 (N2126, N2114, N1310);
buf BUF1 (N2127, N2124);
not NOT1 (N2128, N2088);
buf BUF1 (N2129, N2127);
nor NOR3 (N2130, N2117, N2030, N67);
nor NOR3 (N2131, N2128, N16, N1456);
and AND2 (N2132, N2120, N999);
nand NAND3 (N2133, N2118, N816, N1135);
nand NAND4 (N2134, N2121, N1622, N1909, N38);
buf BUF1 (N2135, N2129);
nor NOR2 (N2136, N2131, N1411);
nor NOR4 (N2137, N2126, N287, N1358, N1584);
or OR4 (N2138, N2136, N2025, N2124, N769);
nand NAND4 (N2139, N2135, N2104, N838, N1081);
or OR2 (N2140, N2138, N1498);
or OR4 (N2141, N2137, N668, N1182, N384);
or OR2 (N2142, N2122, N460);
nand NAND2 (N2143, N2139, N969);
buf BUF1 (N2144, N2133);
and AND3 (N2145, N2134, N1846, N536);
and AND2 (N2146, N2142, N1193);
buf BUF1 (N2147, N2141);
nand NAND3 (N2148, N2147, N970, N1238);
or OR3 (N2149, N2144, N1549, N113);
nor NOR4 (N2150, N2145, N1772, N1175, N14);
nand NAND4 (N2151, N2150, N1547, N1585, N1484);
buf BUF1 (N2152, N2146);
nand NAND4 (N2153, N2149, N1913, N530, N829);
or OR3 (N2154, N2140, N1150, N2012);
nand NAND2 (N2155, N2154, N977);
or OR4 (N2156, N2125, N1013, N1831, N1861);
xor XOR2 (N2157, N2148, N547);
not NOT1 (N2158, N2123);
not NOT1 (N2159, N2156);
not NOT1 (N2160, N2143);
or OR3 (N2161, N2160, N597, N1808);
xor XOR2 (N2162, N2157, N357);
nor NOR4 (N2163, N2151, N993, N1179, N1659);
and AND2 (N2164, N2132, N1994);
xor XOR2 (N2165, N2164, N526);
not NOT1 (N2166, N2155);
not NOT1 (N2167, N2158);
nor NOR3 (N2168, N2167, N1287, N1830);
nor NOR4 (N2169, N2159, N866, N1386, N36);
nor NOR4 (N2170, N2166, N1655, N398, N1485);
and AND4 (N2171, N2152, N1969, N738, N748);
xor XOR2 (N2172, N2170, N981);
xor XOR2 (N2173, N2172, N1197);
xor XOR2 (N2174, N2165, N1583);
nor NOR4 (N2175, N2171, N871, N221, N670);
not NOT1 (N2176, N2175);
and AND3 (N2177, N2153, N1854, N1160);
and AND3 (N2178, N2130, N915, N2144);
buf BUF1 (N2179, N2173);
nand NAND3 (N2180, N2169, N1368, N311);
nand NAND3 (N2181, N2161, N1773, N1350);
not NOT1 (N2182, N2178);
and AND2 (N2183, N2180, N472);
nor NOR3 (N2184, N2177, N1801, N332);
not NOT1 (N2185, N2162);
nand NAND4 (N2186, N2163, N2093, N371, N393);
and AND3 (N2187, N2186, N25, N1247);
xor XOR2 (N2188, N2185, N1683);
buf BUF1 (N2189, N2187);
not NOT1 (N2190, N2168);
nor NOR2 (N2191, N2189, N220);
or OR4 (N2192, N2190, N838, N561, N118);
not NOT1 (N2193, N2192);
and AND2 (N2194, N2193, N287);
or OR4 (N2195, N2181, N1641, N1323, N710);
nand NAND3 (N2196, N2194, N600, N930);
nor NOR3 (N2197, N2179, N1714, N422);
and AND2 (N2198, N2197, N1236);
nor NOR4 (N2199, N2184, N967, N482, N431);
nor NOR4 (N2200, N2176, N1957, N1986, N532);
nand NAND4 (N2201, N2182, N1609, N2057, N1120);
nand NAND3 (N2202, N2188, N674, N492);
and AND4 (N2203, N2200, N578, N1561, N2085);
nor NOR4 (N2204, N2199, N1563, N129, N2151);
not NOT1 (N2205, N2202);
or OR2 (N2206, N2174, N1141);
or OR3 (N2207, N2204, N1695, N1199);
or OR4 (N2208, N2191, N604, N746, N73);
nor NOR4 (N2209, N2195, N1390, N1664, N808);
or OR3 (N2210, N2206, N2134, N1524);
xor XOR2 (N2211, N2196, N1490);
xor XOR2 (N2212, N2203, N214);
nor NOR3 (N2213, N2183, N345, N2163);
xor XOR2 (N2214, N2211, N1316);
nand NAND2 (N2215, N2213, N1307);
nand NAND2 (N2216, N2207, N1653);
nor NOR3 (N2217, N2201, N1792, N333);
and AND3 (N2218, N2209, N2037, N1819);
nor NOR4 (N2219, N2212, N739, N1885, N860);
buf BUF1 (N2220, N2217);
not NOT1 (N2221, N2208);
buf BUF1 (N2222, N2198);
and AND2 (N2223, N2214, N1789);
nor NOR3 (N2224, N2219, N754, N1857);
or OR4 (N2225, N2222, N43, N872, N1837);
nor NOR3 (N2226, N2224, N1713, N1558);
buf BUF1 (N2227, N2225);
not NOT1 (N2228, N2205);
not NOT1 (N2229, N2228);
or OR3 (N2230, N2216, N510, N1941);
not NOT1 (N2231, N2221);
or OR2 (N2232, N2231, N272);
nor NOR2 (N2233, N2220, N700);
xor XOR2 (N2234, N2215, N170);
buf BUF1 (N2235, N2233);
nand NAND2 (N2236, N2230, N945);
and AND2 (N2237, N2218, N1400);
or OR2 (N2238, N2223, N2223);
nor NOR4 (N2239, N2232, N1350, N1724, N1538);
and AND2 (N2240, N2226, N220);
xor XOR2 (N2241, N2237, N871);
nand NAND3 (N2242, N2238, N903, N2223);
and AND2 (N2243, N2235, N954);
nand NAND3 (N2244, N2242, N450, N172);
nor NOR4 (N2245, N2241, N1929, N915, N1448);
buf BUF1 (N2246, N2240);
not NOT1 (N2247, N2210);
not NOT1 (N2248, N2247);
buf BUF1 (N2249, N2245);
buf BUF1 (N2250, N2229);
nand NAND3 (N2251, N2244, N854, N1040);
or OR3 (N2252, N2236, N823, N57);
nand NAND4 (N2253, N2239, N1157, N1785, N411);
or OR2 (N2254, N2251, N763);
nand NAND4 (N2255, N2246, N2063, N1396, N249);
or OR3 (N2256, N2227, N1985, N1985);
buf BUF1 (N2257, N2255);
buf BUF1 (N2258, N2252);
and AND3 (N2259, N2234, N1413, N768);
xor XOR2 (N2260, N2259, N1361);
or OR4 (N2261, N2257, N1178, N2083, N183);
or OR3 (N2262, N2254, N680, N1446);
nor NOR3 (N2263, N2243, N125, N1154);
buf BUF1 (N2264, N2263);
xor XOR2 (N2265, N2248, N1529);
xor XOR2 (N2266, N2250, N1129);
xor XOR2 (N2267, N2249, N301);
or OR3 (N2268, N2256, N2252, N2009);
nand NAND3 (N2269, N2267, N1462, N424);
xor XOR2 (N2270, N2260, N1713);
not NOT1 (N2271, N2269);
nand NAND4 (N2272, N2270, N13, N2072, N640);
nand NAND4 (N2273, N2272, N1478, N2135, N1234);
not NOT1 (N2274, N2253);
buf BUF1 (N2275, N2268);
xor XOR2 (N2276, N2271, N295);
xor XOR2 (N2277, N2276, N2084);
xor XOR2 (N2278, N2274, N1040);
buf BUF1 (N2279, N2278);
nand NAND3 (N2280, N2262, N2259, N2010);
nor NOR3 (N2281, N2277, N469, N2036);
xor XOR2 (N2282, N2258, N186);
buf BUF1 (N2283, N2281);
nor NOR2 (N2284, N2261, N4);
nor NOR4 (N2285, N2266, N969, N2094, N473);
buf BUF1 (N2286, N2265);
or OR4 (N2287, N2280, N1960, N1271, N2162);
nor NOR2 (N2288, N2282, N1793);
nor NOR4 (N2289, N2264, N8, N1361, N1787);
buf BUF1 (N2290, N2287);
buf BUF1 (N2291, N2273);
and AND4 (N2292, N2290, N1265, N1231, N1415);
nor NOR4 (N2293, N2275, N1220, N1664, N1994);
nand NAND2 (N2294, N2284, N1157);
nor NOR4 (N2295, N2293, N74, N1645, N464);
buf BUF1 (N2296, N2289);
and AND3 (N2297, N2285, N1277, N1291);
xor XOR2 (N2298, N2297, N1404);
buf BUF1 (N2299, N2288);
buf BUF1 (N2300, N2298);
nor NOR3 (N2301, N2291, N451, N503);
and AND4 (N2302, N2294, N588, N907, N895);
not NOT1 (N2303, N2300);
nand NAND2 (N2304, N2283, N2219);
and AND3 (N2305, N2303, N1468, N602);
not NOT1 (N2306, N2292);
nor NOR3 (N2307, N2304, N1442, N1330);
xor XOR2 (N2308, N2307, N162);
and AND3 (N2309, N2299, N1104, N1556);
not NOT1 (N2310, N2306);
and AND4 (N2311, N2309, N45, N1877, N673);
nand NAND3 (N2312, N2295, N798, N396);
nor NOR3 (N2313, N2286, N561, N1771);
buf BUF1 (N2314, N2311);
nor NOR2 (N2315, N2313, N841);
buf BUF1 (N2316, N2314);
not NOT1 (N2317, N2296);
or OR2 (N2318, N2301, N657);
nand NAND2 (N2319, N2317, N2136);
buf BUF1 (N2320, N2312);
or OR3 (N2321, N2310, N64, N459);
or OR4 (N2322, N2321, N432, N511, N3);
nor NOR3 (N2323, N2320, N1557, N208);
and AND4 (N2324, N2279, N293, N1995, N1332);
xor XOR2 (N2325, N2305, N2189);
or OR4 (N2326, N2318, N924, N1656, N1253);
and AND3 (N2327, N2315, N1, N2005);
buf BUF1 (N2328, N2326);
xor XOR2 (N2329, N2316, N329);
xor XOR2 (N2330, N2319, N1769);
buf BUF1 (N2331, N2302);
not NOT1 (N2332, N2324);
buf BUF1 (N2333, N2323);
or OR2 (N2334, N2328, N1073);
or OR3 (N2335, N2332, N595, N1403);
buf BUF1 (N2336, N2333);
buf BUF1 (N2337, N2336);
or OR2 (N2338, N2325, N790);
nor NOR2 (N2339, N2338, N1503);
nand NAND4 (N2340, N2308, N1102, N1885, N577);
or OR3 (N2341, N2335, N417, N178);
and AND2 (N2342, N2339, N1679);
and AND4 (N2343, N2337, N2056, N1830, N2133);
not NOT1 (N2344, N2340);
buf BUF1 (N2345, N2344);
nor NOR3 (N2346, N2341, N2115, N1172);
nand NAND4 (N2347, N2345, N2066, N2190, N1436);
and AND2 (N2348, N2342, N2109);
or OR4 (N2349, N2331, N2161, N1327, N811);
buf BUF1 (N2350, N2348);
or OR4 (N2351, N2347, N2232, N685, N1616);
xor XOR2 (N2352, N2346, N381);
nand NAND2 (N2353, N2327, N213);
not NOT1 (N2354, N2343);
nand NAND3 (N2355, N2322, N833, N1071);
nor NOR3 (N2356, N2334, N417, N1760);
nand NAND2 (N2357, N2355, N2222);
xor XOR2 (N2358, N2354, N1295);
or OR2 (N2359, N2329, N139);
or OR2 (N2360, N2330, N432);
buf BUF1 (N2361, N2349);
or OR4 (N2362, N2360, N1353, N2200, N1633);
and AND2 (N2363, N2362, N1855);
nand NAND2 (N2364, N2351, N1180);
or OR4 (N2365, N2363, N2151, N554, N1867);
nor NOR2 (N2366, N2357, N1770);
buf BUF1 (N2367, N2365);
not NOT1 (N2368, N2367);
buf BUF1 (N2369, N2364);
or OR2 (N2370, N2359, N264);
xor XOR2 (N2371, N2356, N617);
xor XOR2 (N2372, N2350, N1392);
nand NAND3 (N2373, N2352, N913, N1393);
nor NOR2 (N2374, N2366, N1790);
not NOT1 (N2375, N2353);
xor XOR2 (N2376, N2369, N396);
or OR3 (N2377, N2375, N1583, N1072);
or OR2 (N2378, N2361, N2026);
xor XOR2 (N2379, N2377, N334);
buf BUF1 (N2380, N2372);
nand NAND3 (N2381, N2379, N956, N2161);
nand NAND2 (N2382, N2378, N2052);
and AND2 (N2383, N2381, N2161);
and AND2 (N2384, N2370, N1570);
nor NOR2 (N2385, N2380, N376);
buf BUF1 (N2386, N2368);
not NOT1 (N2387, N2386);
nand NAND2 (N2388, N2376, N224);
nand NAND3 (N2389, N2383, N2361, N1396);
xor XOR2 (N2390, N2374, N106);
and AND3 (N2391, N2382, N1031, N1741);
nor NOR3 (N2392, N2373, N2201, N99);
nand NAND4 (N2393, N2371, N2112, N1085, N332);
not NOT1 (N2394, N2391);
or OR2 (N2395, N2392, N380);
or OR2 (N2396, N2388, N1538);
not NOT1 (N2397, N2395);
nor NOR3 (N2398, N2389, N555, N1991);
not NOT1 (N2399, N2358);
not NOT1 (N2400, N2385);
xor XOR2 (N2401, N2396, N798);
nor NOR4 (N2402, N2401, N658, N768, N1496);
not NOT1 (N2403, N2400);
and AND4 (N2404, N2393, N1781, N2097, N369);
or OR3 (N2405, N2390, N2352, N330);
xor XOR2 (N2406, N2398, N926);
buf BUF1 (N2407, N2387);
buf BUF1 (N2408, N2399);
and AND2 (N2409, N2405, N2405);
nor NOR3 (N2410, N2404, N1914, N2282);
nand NAND4 (N2411, N2403, N1031, N1812, N1849);
nand NAND2 (N2412, N2394, N370);
xor XOR2 (N2413, N2412, N2318);
nand NAND2 (N2414, N2410, N261);
and AND4 (N2415, N2411, N259, N1876, N1299);
buf BUF1 (N2416, N2402);
xor XOR2 (N2417, N2406, N41);
or OR3 (N2418, N2415, N661, N722);
and AND2 (N2419, N2407, N2108);
nand NAND3 (N2420, N2417, N1806, N1004);
not NOT1 (N2421, N2414);
or OR2 (N2422, N2419, N2086);
not NOT1 (N2423, N2397);
not NOT1 (N2424, N2421);
and AND2 (N2425, N2413, N1915);
nor NOR4 (N2426, N2416, N1456, N1136, N1041);
not NOT1 (N2427, N2425);
nand NAND2 (N2428, N2384, N1270);
buf BUF1 (N2429, N2409);
not NOT1 (N2430, N2424);
nor NOR3 (N2431, N2408, N399, N1130);
nand NAND4 (N2432, N2429, N1969, N1711, N1361);
xor XOR2 (N2433, N2420, N2098);
not NOT1 (N2434, N2428);
or OR4 (N2435, N2433, N2413, N1251, N1031);
nor NOR2 (N2436, N2435, N455);
buf BUF1 (N2437, N2427);
and AND3 (N2438, N2430, N981, N642);
and AND3 (N2439, N2432, N617, N651);
nor NOR3 (N2440, N2418, N2166, N2178);
nor NOR4 (N2441, N2438, N770, N834, N459);
and AND2 (N2442, N2441, N621);
nand NAND3 (N2443, N2434, N2380, N1154);
buf BUF1 (N2444, N2436);
and AND3 (N2445, N2422, N499, N1722);
nand NAND3 (N2446, N2426, N2335, N17);
not NOT1 (N2447, N2442);
and AND4 (N2448, N2444, N203, N323, N1639);
or OR4 (N2449, N2423, N388, N118, N2035);
buf BUF1 (N2450, N2439);
and AND4 (N2451, N2448, N894, N897, N2400);
buf BUF1 (N2452, N2451);
or OR4 (N2453, N2443, N975, N1633, N314);
or OR3 (N2454, N2437, N947, N1241);
xor XOR2 (N2455, N2453, N1367);
and AND3 (N2456, N2431, N698, N2437);
xor XOR2 (N2457, N2454, N224);
and AND2 (N2458, N2449, N1392);
buf BUF1 (N2459, N2445);
not NOT1 (N2460, N2452);
or OR3 (N2461, N2460, N651, N361);
and AND3 (N2462, N2446, N269, N1722);
nand NAND3 (N2463, N2462, N256, N161);
or OR3 (N2464, N2463, N2017, N1392);
nand NAND2 (N2465, N2440, N1565);
nor NOR3 (N2466, N2461, N163, N1408);
nor NOR3 (N2467, N2464, N298, N77);
xor XOR2 (N2468, N2455, N854);
and AND4 (N2469, N2447, N665, N2444, N2151);
xor XOR2 (N2470, N2468, N1399);
buf BUF1 (N2471, N2456);
and AND2 (N2472, N2459, N1725);
nor NOR2 (N2473, N2465, N7);
and AND3 (N2474, N2466, N1248, N1207);
not NOT1 (N2475, N2471);
nor NOR2 (N2476, N2457, N2049);
not NOT1 (N2477, N2450);
nand NAND4 (N2478, N2473, N2247, N390, N884);
nor NOR3 (N2479, N2470, N813, N1471);
buf BUF1 (N2480, N2467);
nand NAND2 (N2481, N2480, N1343);
not NOT1 (N2482, N2458);
buf BUF1 (N2483, N2469);
not NOT1 (N2484, N2475);
buf BUF1 (N2485, N2483);
or OR2 (N2486, N2481, N875);
buf BUF1 (N2487, N2476);
buf BUF1 (N2488, N2474);
not NOT1 (N2489, N2482);
nand NAND4 (N2490, N2478, N480, N1294, N1658);
and AND2 (N2491, N2479, N2106);
and AND3 (N2492, N2489, N1056, N1495);
and AND4 (N2493, N2490, N1918, N2290, N182);
xor XOR2 (N2494, N2493, N497);
buf BUF1 (N2495, N2491);
nand NAND3 (N2496, N2487, N898, N1464);
and AND3 (N2497, N2485, N400, N1662);
nor NOR4 (N2498, N2477, N1430, N2065, N269);
nand NAND2 (N2499, N2496, N110);
or OR3 (N2500, N2488, N2035, N1920);
and AND3 (N2501, N2494, N335, N516);
and AND4 (N2502, N2472, N1731, N451, N820);
nand NAND3 (N2503, N2501, N428, N597);
xor XOR2 (N2504, N2495, N821);
buf BUF1 (N2505, N2502);
nor NOR3 (N2506, N2497, N4, N848);
nor NOR4 (N2507, N2492, N2042, N378, N101);
nor NOR3 (N2508, N2506, N2417, N354);
not NOT1 (N2509, N2484);
buf BUF1 (N2510, N2508);
and AND2 (N2511, N2499, N1169);
or OR4 (N2512, N2498, N1089, N2131, N1437);
or OR4 (N2513, N2486, N889, N1370, N2275);
nor NOR2 (N2514, N2512, N277);
xor XOR2 (N2515, N2511, N1330);
xor XOR2 (N2516, N2513, N2511);
not NOT1 (N2517, N2505);
buf BUF1 (N2518, N2517);
and AND2 (N2519, N2518, N2237);
and AND2 (N2520, N2507, N790);
nand NAND4 (N2521, N2516, N2491, N1983, N837);
xor XOR2 (N2522, N2504, N219);
xor XOR2 (N2523, N2521, N1230);
or OR3 (N2524, N2514, N928, N1164);
xor XOR2 (N2525, N2515, N2064);
not NOT1 (N2526, N2520);
buf BUF1 (N2527, N2526);
nor NOR2 (N2528, N2503, N1162);
buf BUF1 (N2529, N2523);
nor NOR4 (N2530, N2529, N1303, N1788, N2236);
buf BUF1 (N2531, N2525);
not NOT1 (N2532, N2527);
xor XOR2 (N2533, N2522, N1764);
xor XOR2 (N2534, N2531, N928);
nor NOR3 (N2535, N2509, N2270, N1641);
xor XOR2 (N2536, N2533, N1718);
not NOT1 (N2537, N2524);
or OR4 (N2538, N2537, N1556, N2477, N722);
nor NOR4 (N2539, N2519, N602, N195, N1080);
buf BUF1 (N2540, N2535);
not NOT1 (N2541, N2528);
and AND2 (N2542, N2534, N349);
or OR2 (N2543, N2542, N1318);
nand NAND2 (N2544, N2538, N1880);
or OR2 (N2545, N2510, N664);
not NOT1 (N2546, N2539);
buf BUF1 (N2547, N2540);
buf BUF1 (N2548, N2543);
xor XOR2 (N2549, N2532, N65);
and AND3 (N2550, N2548, N207, N992);
and AND2 (N2551, N2545, N2130);
nor NOR4 (N2552, N2541, N971, N2132, N331);
xor XOR2 (N2553, N2550, N2137);
nor NOR2 (N2554, N2552, N2029);
xor XOR2 (N2555, N2547, N923);
xor XOR2 (N2556, N2536, N939);
buf BUF1 (N2557, N2544);
nand NAND2 (N2558, N2546, N609);
buf BUF1 (N2559, N2500);
not NOT1 (N2560, N2530);
nor NOR2 (N2561, N2555, N1044);
and AND2 (N2562, N2560, N578);
nor NOR4 (N2563, N2551, N2173, N125, N1);
nor NOR4 (N2564, N2562, N612, N207, N1929);
xor XOR2 (N2565, N2558, N612);
or OR3 (N2566, N2564, N2537, N189);
nor NOR3 (N2567, N2553, N819, N1612);
or OR4 (N2568, N2566, N175, N1903, N1313);
and AND2 (N2569, N2556, N1215);
xor XOR2 (N2570, N2559, N1537);
or OR4 (N2571, N2570, N953, N1915, N2388);
or OR3 (N2572, N2557, N1810, N2559);
nand NAND2 (N2573, N2554, N702);
xor XOR2 (N2574, N2565, N1573);
and AND2 (N2575, N2573, N2467);
xor XOR2 (N2576, N2549, N2206);
or OR2 (N2577, N2568, N210);
nor NOR3 (N2578, N2563, N1250, N1617);
not NOT1 (N2579, N2575);
and AND3 (N2580, N2572, N240, N1526);
nand NAND3 (N2581, N2576, N2102, N1150);
or OR3 (N2582, N2577, N908, N469);
nand NAND3 (N2583, N2581, N1876, N2087);
xor XOR2 (N2584, N2571, N2551);
not NOT1 (N2585, N2583);
and AND4 (N2586, N2569, N1264, N1023, N1390);
nor NOR4 (N2587, N2574, N794, N1480, N140);
and AND3 (N2588, N2561, N1781, N1727);
nand NAND2 (N2589, N2578, N1228);
or OR4 (N2590, N2586, N2357, N1494, N732);
and AND4 (N2591, N2585, N1951, N735, N942);
nand NAND3 (N2592, N2582, N981, N1959);
nand NAND3 (N2593, N2567, N2228, N2102);
and AND3 (N2594, N2589, N796, N2332);
nor NOR3 (N2595, N2587, N877, N667);
buf BUF1 (N2596, N2595);
nor NOR4 (N2597, N2593, N670, N816, N2232);
xor XOR2 (N2598, N2594, N341);
and AND3 (N2599, N2591, N2288, N832);
xor XOR2 (N2600, N2599, N95);
nor NOR2 (N2601, N2597, N737);
nor NOR3 (N2602, N2600, N784, N75);
buf BUF1 (N2603, N2588);
or OR4 (N2604, N2602, N1630, N2181, N810);
and AND4 (N2605, N2590, N2547, N500, N1720);
nand NAND2 (N2606, N2598, N2076);
not NOT1 (N2607, N2579);
or OR4 (N2608, N2592, N988, N367, N302);
or OR4 (N2609, N2596, N822, N1538, N803);
not NOT1 (N2610, N2604);
nand NAND4 (N2611, N2601, N992, N2601, N2035);
not NOT1 (N2612, N2608);
nand NAND3 (N2613, N2605, N622, N515);
not NOT1 (N2614, N2603);
not NOT1 (N2615, N2607);
nor NOR2 (N2616, N2580, N843);
buf BUF1 (N2617, N2609);
buf BUF1 (N2618, N2611);
not NOT1 (N2619, N2606);
nand NAND2 (N2620, N2610, N241);
and AND2 (N2621, N2615, N360);
buf BUF1 (N2622, N2617);
and AND3 (N2623, N2619, N1055, N960);
nand NAND3 (N2624, N2622, N324, N566);
nand NAND4 (N2625, N2620, N1654, N1101, N910);
or OR4 (N2626, N2625, N1288, N900, N1621);
nand NAND3 (N2627, N2616, N2323, N1952);
xor XOR2 (N2628, N2614, N1963);
and AND4 (N2629, N2628, N725, N518, N2160);
not NOT1 (N2630, N2627);
nand NAND2 (N2631, N2612, N1364);
nor NOR4 (N2632, N2621, N1190, N2033, N1097);
or OR3 (N2633, N2584, N2064, N1338);
nor NOR4 (N2634, N2632, N76, N121, N728);
buf BUF1 (N2635, N2630);
nor NOR2 (N2636, N2635, N621);
nand NAND2 (N2637, N2618, N1471);
or OR2 (N2638, N2634, N1923);
and AND4 (N2639, N2638, N559, N764, N2027);
nand NAND2 (N2640, N2629, N1051);
and AND3 (N2641, N2613, N2255, N1747);
or OR4 (N2642, N2633, N644, N1722, N447);
nor NOR3 (N2643, N2624, N775, N1578);
and AND3 (N2644, N2641, N863, N2075);
or OR4 (N2645, N2631, N1961, N966, N2045);
nand NAND4 (N2646, N2639, N1059, N1607, N1331);
nand NAND3 (N2647, N2637, N1400, N1999);
not NOT1 (N2648, N2626);
nand NAND3 (N2649, N2643, N2000, N930);
xor XOR2 (N2650, N2649, N1803);
or OR4 (N2651, N2642, N2433, N1702, N2296);
nor NOR4 (N2652, N2647, N169, N2081, N2059);
and AND2 (N2653, N2650, N2173);
or OR2 (N2654, N2644, N1333);
nand NAND2 (N2655, N2640, N1043);
xor XOR2 (N2656, N2636, N359);
nand NAND4 (N2657, N2653, N2553, N979, N2009);
or OR4 (N2658, N2645, N2136, N2342, N582);
not NOT1 (N2659, N2648);
nand NAND3 (N2660, N2657, N620, N73);
or OR4 (N2661, N2658, N701, N2230, N1109);
or OR4 (N2662, N2661, N2485, N850, N465);
nor NOR2 (N2663, N2656, N287);
buf BUF1 (N2664, N2663);
nor NOR3 (N2665, N2662, N370, N494);
nor NOR3 (N2666, N2660, N1563, N1018);
xor XOR2 (N2667, N2623, N678);
and AND2 (N2668, N2667, N1405);
nand NAND2 (N2669, N2655, N1673);
and AND3 (N2670, N2659, N1663, N2458);
buf BUF1 (N2671, N2664);
buf BUF1 (N2672, N2668);
xor XOR2 (N2673, N2651, N968);
nor NOR4 (N2674, N2665, N1272, N438, N491);
or OR2 (N2675, N2671, N2136);
buf BUF1 (N2676, N2646);
not NOT1 (N2677, N2669);
not NOT1 (N2678, N2674);
buf BUF1 (N2679, N2676);
nand NAND2 (N2680, N2678, N612);
or OR4 (N2681, N2677, N964, N1706, N984);
xor XOR2 (N2682, N2670, N168);
nand NAND4 (N2683, N2679, N88, N295, N1560);
buf BUF1 (N2684, N2673);
nand NAND2 (N2685, N2652, N433);
buf BUF1 (N2686, N2675);
not NOT1 (N2687, N2685);
and AND4 (N2688, N2683, N731, N332, N1882);
nor NOR3 (N2689, N2681, N1907, N18);
xor XOR2 (N2690, N2682, N1612);
or OR4 (N2691, N2690, N2488, N565, N1416);
xor XOR2 (N2692, N2686, N1643);
nand NAND4 (N2693, N2680, N370, N1342, N421);
nand NAND4 (N2694, N2692, N1727, N321, N1388);
buf BUF1 (N2695, N2666);
not NOT1 (N2696, N2694);
nor NOR2 (N2697, N2689, N2151);
and AND4 (N2698, N2672, N748, N2412, N2363);
not NOT1 (N2699, N2654);
and AND4 (N2700, N2696, N1438, N1051, N261);
not NOT1 (N2701, N2699);
nand NAND4 (N2702, N2701, N433, N2331, N1266);
and AND2 (N2703, N2691, N810);
xor XOR2 (N2704, N2700, N2395);
nor NOR3 (N2705, N2697, N1351, N1806);
nand NAND3 (N2706, N2684, N1018, N2438);
or OR2 (N2707, N2688, N1620);
and AND3 (N2708, N2706, N2081, N2098);
nand NAND3 (N2709, N2698, N2185, N772);
nor NOR2 (N2710, N2709, N1931);
buf BUF1 (N2711, N2704);
and AND2 (N2712, N2708, N561);
nand NAND3 (N2713, N2711, N1594, N135);
nand NAND2 (N2714, N2702, N112);
and AND4 (N2715, N2687, N2225, N800, N2148);
and AND2 (N2716, N2693, N1298);
nand NAND4 (N2717, N2710, N2201, N2273, N512);
nor NOR4 (N2718, N2716, N1106, N9, N452);
or OR2 (N2719, N2713, N2559);
or OR4 (N2720, N2695, N2527, N1734, N2605);
xor XOR2 (N2721, N2720, N2172);
xor XOR2 (N2722, N2703, N616);
xor XOR2 (N2723, N2718, N542);
or OR2 (N2724, N2707, N1556);
not NOT1 (N2725, N2722);
xor XOR2 (N2726, N2725, N1494);
nor NOR2 (N2727, N2712, N2647);
and AND3 (N2728, N2715, N2324, N2685);
xor XOR2 (N2729, N2719, N2091);
or OR2 (N2730, N2717, N2537);
not NOT1 (N2731, N2727);
nor NOR3 (N2732, N2721, N1757, N401);
buf BUF1 (N2733, N2724);
and AND2 (N2734, N2732, N58);
xor XOR2 (N2735, N2731, N1756);
or OR2 (N2736, N2734, N1437);
xor XOR2 (N2737, N2723, N2114);
nor NOR3 (N2738, N2705, N799, N1721);
not NOT1 (N2739, N2736);
and AND2 (N2740, N2735, N871);
xor XOR2 (N2741, N2738, N1312);
nor NOR4 (N2742, N2737, N106, N1805, N1050);
not NOT1 (N2743, N2728);
nand NAND4 (N2744, N2741, N120, N885, N2543);
and AND2 (N2745, N2733, N675);
nand NAND2 (N2746, N2745, N765);
nand NAND3 (N2747, N2729, N335, N2240);
nor NOR2 (N2748, N2739, N393);
and AND3 (N2749, N2714, N937, N1524);
and AND4 (N2750, N2747, N1051, N280, N1874);
nand NAND4 (N2751, N2750, N639, N516, N626);
not NOT1 (N2752, N2740);
and AND3 (N2753, N2752, N2597, N1695);
xor XOR2 (N2754, N2744, N1106);
nor NOR2 (N2755, N2751, N223);
nor NOR3 (N2756, N2754, N1929, N1476);
not NOT1 (N2757, N2743);
or OR2 (N2758, N2749, N564);
xor XOR2 (N2759, N2756, N1139);
and AND2 (N2760, N2759, N2204);
or OR3 (N2761, N2758, N1921, N2556);
xor XOR2 (N2762, N2757, N3);
and AND4 (N2763, N2762, N1229, N2022, N1413);
nor NOR2 (N2764, N2726, N1928);
nor NOR4 (N2765, N2760, N938, N385, N2167);
not NOT1 (N2766, N2761);
nand NAND2 (N2767, N2753, N2316);
or OR4 (N2768, N2766, N852, N571, N1065);
buf BUF1 (N2769, N2768);
and AND3 (N2770, N2765, N2596, N1250);
buf BUF1 (N2771, N2769);
nand NAND2 (N2772, N2771, N1519);
and AND4 (N2773, N2755, N2151, N1973, N1236);
buf BUF1 (N2774, N2742);
nor NOR4 (N2775, N2748, N2033, N1491, N1206);
xor XOR2 (N2776, N2767, N2631);
not NOT1 (N2777, N2774);
xor XOR2 (N2778, N2730, N595);
and AND4 (N2779, N2777, N2501, N1211, N940);
nor NOR2 (N2780, N2779, N2058);
buf BUF1 (N2781, N2764);
buf BUF1 (N2782, N2770);
buf BUF1 (N2783, N2782);
and AND4 (N2784, N2746, N1652, N1981, N2202);
xor XOR2 (N2785, N2773, N1469);
not NOT1 (N2786, N2780);
buf BUF1 (N2787, N2784);
buf BUF1 (N2788, N2781);
xor XOR2 (N2789, N2776, N143);
or OR3 (N2790, N2778, N1593, N143);
buf BUF1 (N2791, N2787);
and AND4 (N2792, N2763, N2154, N799, N2121);
or OR2 (N2793, N2786, N2631);
nand NAND2 (N2794, N2788, N915);
buf BUF1 (N2795, N2783);
nor NOR4 (N2796, N2790, N2253, N1173, N2037);
nor NOR2 (N2797, N2791, N2035);
nor NOR4 (N2798, N2785, N1801, N867, N2747);
and AND3 (N2799, N2789, N728, N698);
and AND2 (N2800, N2797, N2489);
or OR4 (N2801, N2800, N1540, N1172, N755);
xor XOR2 (N2802, N2799, N2141);
xor XOR2 (N2803, N2795, N2487);
not NOT1 (N2804, N2794);
or OR2 (N2805, N2772, N2563);
nand NAND4 (N2806, N2802, N2440, N2742, N687);
buf BUF1 (N2807, N2806);
not NOT1 (N2808, N2805);
and AND3 (N2809, N2801, N621, N1059);
nand NAND4 (N2810, N2798, N2346, N1268, N2710);
nor NOR4 (N2811, N2804, N1931, N810, N774);
buf BUF1 (N2812, N2793);
or OR4 (N2813, N2812, N397, N993, N1112);
or OR4 (N2814, N2792, N1923, N1061, N306);
xor XOR2 (N2815, N2803, N117);
and AND2 (N2816, N2808, N1101);
not NOT1 (N2817, N2815);
buf BUF1 (N2818, N2796);
and AND4 (N2819, N2817, N2614, N324, N2258);
nor NOR2 (N2820, N2810, N732);
nand NAND2 (N2821, N2809, N2714);
and AND3 (N2822, N2814, N1428, N1920);
and AND3 (N2823, N2819, N377, N1755);
or OR3 (N2824, N2811, N320, N477);
buf BUF1 (N2825, N2820);
not NOT1 (N2826, N2818);
xor XOR2 (N2827, N2813, N2104);
and AND4 (N2828, N2821, N2350, N52, N1960);
and AND3 (N2829, N2826, N1499, N1139);
or OR3 (N2830, N2775, N827, N1281);
not NOT1 (N2831, N2807);
buf BUF1 (N2832, N2824);
nor NOR4 (N2833, N2823, N2352, N2312, N1717);
nor NOR3 (N2834, N2833, N1577, N324);
buf BUF1 (N2835, N2832);
and AND2 (N2836, N2835, N569);
xor XOR2 (N2837, N2828, N2450);
or OR4 (N2838, N2822, N1498, N1312, N1417);
buf BUF1 (N2839, N2834);
not NOT1 (N2840, N2830);
nor NOR4 (N2841, N2825, N1783, N2487, N1640);
nand NAND4 (N2842, N2837, N2046, N1358, N2185);
and AND4 (N2843, N2836, N207, N155, N749);
buf BUF1 (N2844, N2841);
xor XOR2 (N2845, N2844, N1439);
not NOT1 (N2846, N2831);
xor XOR2 (N2847, N2845, N901);
nand NAND2 (N2848, N2847, N361);
nand NAND3 (N2849, N2816, N1327, N1168);
or OR4 (N2850, N2838, N868, N1583, N2650);
not NOT1 (N2851, N2849);
and AND3 (N2852, N2851, N1222, N397);
not NOT1 (N2853, N2827);
and AND2 (N2854, N2852, N1047);
xor XOR2 (N2855, N2842, N929);
or OR2 (N2856, N2855, N2430);
buf BUF1 (N2857, N2853);
nand NAND4 (N2858, N2857, N2596, N2272, N879);
and AND3 (N2859, N2839, N2691, N2248);
not NOT1 (N2860, N2843);
nand NAND4 (N2861, N2860, N171, N774, N470);
and AND3 (N2862, N2858, N2491, N2395);
nor NOR4 (N2863, N2859, N2238, N954, N1354);
xor XOR2 (N2864, N2850, N763);
not NOT1 (N2865, N2864);
and AND2 (N2866, N2862, N678);
and AND2 (N2867, N2829, N12);
xor XOR2 (N2868, N2863, N87);
xor XOR2 (N2869, N2840, N680);
xor XOR2 (N2870, N2856, N1368);
not NOT1 (N2871, N2868);
nand NAND2 (N2872, N2867, N2272);
xor XOR2 (N2873, N2848, N2131);
nor NOR3 (N2874, N2866, N802, N2725);
and AND4 (N2875, N2873, N333, N2264, N2316);
nand NAND2 (N2876, N2872, N854);
and AND3 (N2877, N2869, N1327, N268);
and AND4 (N2878, N2870, N1784, N2589, N1875);
nand NAND2 (N2879, N2875, N1452);
and AND4 (N2880, N2879, N1760, N1147, N893);
nand NAND3 (N2881, N2854, N223, N1856);
xor XOR2 (N2882, N2878, N1947);
or OR4 (N2883, N2846, N2331, N1934, N2846);
xor XOR2 (N2884, N2871, N1284);
not NOT1 (N2885, N2861);
xor XOR2 (N2886, N2865, N856);
not NOT1 (N2887, N2876);
or OR4 (N2888, N2884, N699, N2002, N308);
xor XOR2 (N2889, N2874, N340);
xor XOR2 (N2890, N2882, N1822);
or OR4 (N2891, N2885, N960, N231, N2608);
and AND4 (N2892, N2891, N56, N1587, N1408);
or OR2 (N2893, N2890, N2875);
nor NOR3 (N2894, N2892, N939, N576);
buf BUF1 (N2895, N2880);
not NOT1 (N2896, N2895);
or OR3 (N2897, N2877, N820, N2625);
and AND3 (N2898, N2894, N951, N991);
nor NOR2 (N2899, N2883, N817);
nor NOR3 (N2900, N2887, N2446, N2);
not NOT1 (N2901, N2899);
buf BUF1 (N2902, N2900);
nor NOR4 (N2903, N2889, N1818, N1290, N1325);
nor NOR4 (N2904, N2886, N1699, N2900, N1386);
xor XOR2 (N2905, N2898, N2434);
nor NOR3 (N2906, N2896, N2847, N1500);
nor NOR4 (N2907, N2888, N2825, N639, N1877);
xor XOR2 (N2908, N2905, N1938);
buf BUF1 (N2909, N2881);
buf BUF1 (N2910, N2907);
nor NOR2 (N2911, N2910, N1195);
xor XOR2 (N2912, N2903, N993);
buf BUF1 (N2913, N2911);
buf BUF1 (N2914, N2897);
xor XOR2 (N2915, N2912, N1140);
nor NOR3 (N2916, N2908, N2732, N381);
buf BUF1 (N2917, N2914);
xor XOR2 (N2918, N2906, N278);
or OR3 (N2919, N2902, N171, N1221);
not NOT1 (N2920, N2915);
nor NOR3 (N2921, N2919, N1101, N35);
xor XOR2 (N2922, N2913, N470);
xor XOR2 (N2923, N2916, N2095);
xor XOR2 (N2924, N2893, N997);
nor NOR3 (N2925, N2922, N2888, N1083);
buf BUF1 (N2926, N2909);
buf BUF1 (N2927, N2923);
xor XOR2 (N2928, N2927, N603);
xor XOR2 (N2929, N2924, N543);
nor NOR4 (N2930, N2925, N2740, N598, N434);
buf BUF1 (N2931, N2904);
xor XOR2 (N2932, N2931, N2688);
xor XOR2 (N2933, N2921, N2144);
nand NAND3 (N2934, N2920, N311, N232);
and AND2 (N2935, N2933, N1758);
and AND3 (N2936, N2917, N2647, N1796);
buf BUF1 (N2937, N2901);
nand NAND2 (N2938, N2936, N1524);
or OR4 (N2939, N2918, N1398, N1723, N908);
not NOT1 (N2940, N2938);
nand NAND4 (N2941, N2934, N2430, N578, N2052);
not NOT1 (N2942, N2929);
nand NAND3 (N2943, N2928, N2099, N892);
nand NAND3 (N2944, N2935, N728, N1439);
nand NAND2 (N2945, N2930, N2285);
not NOT1 (N2946, N2941);
and AND4 (N2947, N2932, N66, N1375, N1091);
nand NAND3 (N2948, N2947, N958, N2740);
xor XOR2 (N2949, N2942, N762);
xor XOR2 (N2950, N2939, N545);
not NOT1 (N2951, N2937);
or OR4 (N2952, N2943, N342, N420, N307);
not NOT1 (N2953, N2926);
or OR4 (N2954, N2949, N2774, N390, N2343);
nand NAND2 (N2955, N2950, N213);
xor XOR2 (N2956, N2954, N421);
nor NOR3 (N2957, N2944, N713, N2304);
xor XOR2 (N2958, N2957, N868);
buf BUF1 (N2959, N2945);
nand NAND3 (N2960, N2956, N669, N2651);
not NOT1 (N2961, N2959);
nand NAND3 (N2962, N2948, N1279, N2330);
and AND4 (N2963, N2955, N507, N2928, N362);
and AND4 (N2964, N2940, N1617, N827, N457);
buf BUF1 (N2965, N2960);
nand NAND2 (N2966, N2962, N2767);
buf BUF1 (N2967, N2951);
buf BUF1 (N2968, N2946);
or OR3 (N2969, N2953, N416, N1808);
xor XOR2 (N2970, N2963, N1264);
nor NOR4 (N2971, N2966, N1054, N2631, N2839);
buf BUF1 (N2972, N2967);
nor NOR2 (N2973, N2970, N318);
not NOT1 (N2974, N2971);
buf BUF1 (N2975, N2974);
nand NAND4 (N2976, N2961, N1353, N1387, N2710);
nor NOR2 (N2977, N2965, N1466);
not NOT1 (N2978, N2964);
and AND3 (N2979, N2976, N1098, N452);
or OR3 (N2980, N2973, N2616, N559);
buf BUF1 (N2981, N2968);
nor NOR4 (N2982, N2980, N873, N1881, N837);
nand NAND4 (N2983, N2958, N1605, N513, N1208);
buf BUF1 (N2984, N2972);
or OR4 (N2985, N2975, N2735, N690, N1644);
buf BUF1 (N2986, N2977);
and AND3 (N2987, N2978, N421, N1616);
or OR2 (N2988, N2987, N869);
nor NOR3 (N2989, N2969, N459, N579);
buf BUF1 (N2990, N2985);
and AND4 (N2991, N2990, N874, N2419, N847);
nand NAND3 (N2992, N2984, N2898, N2738);
nor NOR2 (N2993, N2952, N2295);
nand NAND2 (N2994, N2986, N2);
and AND3 (N2995, N2994, N2858, N2830);
and AND3 (N2996, N2979, N2570, N1668);
not NOT1 (N2997, N2989);
not NOT1 (N2998, N2992);
xor XOR2 (N2999, N2998, N2691);
buf BUF1 (N3000, N2982);
or OR2 (N3001, N2995, N831);
or OR2 (N3002, N3000, N1902);
not NOT1 (N3003, N2991);
or OR4 (N3004, N3002, N912, N344, N723);
xor XOR2 (N3005, N2999, N1989);
buf BUF1 (N3006, N2981);
or OR3 (N3007, N2997, N2584, N611);
nand NAND4 (N3008, N2988, N583, N1988, N2088);
not NOT1 (N3009, N3006);
nor NOR3 (N3010, N2996, N34, N2998);
buf BUF1 (N3011, N3004);
not NOT1 (N3012, N3008);
not NOT1 (N3013, N3007);
or OR4 (N3014, N3011, N2319, N2869, N1788);
nor NOR3 (N3015, N3014, N2977, N698);
or OR4 (N3016, N3012, N1602, N285, N1284);
xor XOR2 (N3017, N2993, N1596);
xor XOR2 (N3018, N3016, N2699);
xor XOR2 (N3019, N3018, N2818);
buf BUF1 (N3020, N3017);
nor NOR3 (N3021, N3003, N2559, N1440);
xor XOR2 (N3022, N3020, N472);
nor NOR3 (N3023, N3013, N2855, N2947);
or OR3 (N3024, N3010, N951, N2304);
not NOT1 (N3025, N3021);
and AND2 (N3026, N3015, N1733);
nand NAND3 (N3027, N2983, N1714, N1129);
not NOT1 (N3028, N3024);
or OR2 (N3029, N3019, N2559);
nand NAND3 (N3030, N3026, N1796, N2020);
xor XOR2 (N3031, N3029, N532);
and AND3 (N3032, N3022, N831, N2875);
nor NOR3 (N3033, N3030, N639, N2553);
buf BUF1 (N3034, N3027);
and AND4 (N3035, N3009, N1293, N1891, N1382);
or OR3 (N3036, N3031, N2203, N2820);
and AND4 (N3037, N3034, N1910, N2444, N2070);
not NOT1 (N3038, N3023);
not NOT1 (N3039, N3038);
xor XOR2 (N3040, N3025, N181);
nor NOR3 (N3041, N3035, N70, N2339);
nor NOR2 (N3042, N3032, N1642);
nor NOR4 (N3043, N3040, N2512, N2545, N2635);
or OR3 (N3044, N3001, N1000, N2948);
not NOT1 (N3045, N3043);
nor NOR2 (N3046, N3045, N1902);
xor XOR2 (N3047, N3046, N1763);
or OR2 (N3048, N3042, N1657);
xor XOR2 (N3049, N3041, N1247);
xor XOR2 (N3050, N3047, N245);
nor NOR2 (N3051, N3036, N191);
nor NOR4 (N3052, N3051, N1635, N78, N2832);
or OR4 (N3053, N3050, N483, N32, N243);
nand NAND4 (N3054, N3005, N922, N2793, N2739);
or OR4 (N3055, N3044, N1400, N2893, N2556);
xor XOR2 (N3056, N3049, N1579);
nor NOR3 (N3057, N3053, N1570, N987);
nand NAND2 (N3058, N3052, N2673);
buf BUF1 (N3059, N3056);
nor NOR2 (N3060, N3059, N2221);
xor XOR2 (N3061, N3058, N1745);
nand NAND4 (N3062, N3057, N1195, N497, N7);
and AND4 (N3063, N3048, N607, N2633, N1633);
nand NAND2 (N3064, N3055, N597);
nand NAND4 (N3065, N3033, N106, N2943, N2551);
xor XOR2 (N3066, N3028, N956);
and AND4 (N3067, N3054, N10, N1679, N1096);
buf BUF1 (N3068, N3063);
nor NOR2 (N3069, N3039, N503);
or OR4 (N3070, N3064, N267, N1437, N910);
and AND4 (N3071, N3060, N2155, N1555, N550);
not NOT1 (N3072, N3067);
nor NOR4 (N3073, N3072, N2319, N678, N1061);
nand NAND4 (N3074, N3071, N2034, N3058, N1324);
and AND3 (N3075, N3068, N1663, N713);
nor NOR2 (N3076, N3073, N1604);
not NOT1 (N3077, N3074);
not NOT1 (N3078, N3066);
and AND3 (N3079, N3069, N2852, N2777);
nor NOR3 (N3080, N3037, N2887, N2932);
and AND4 (N3081, N3061, N2304, N1488, N2883);
xor XOR2 (N3082, N3076, N1314);
buf BUF1 (N3083, N3065);
nor NOR3 (N3084, N3081, N1023, N1556);
nand NAND4 (N3085, N3079, N2793, N2351, N1668);
and AND2 (N3086, N3070, N1030);
not NOT1 (N3087, N3084);
nor NOR2 (N3088, N3087, N2443);
nor NOR4 (N3089, N3082, N2724, N30, N2609);
buf BUF1 (N3090, N3085);
not NOT1 (N3091, N3080);
nand NAND4 (N3092, N3086, N2744, N1097, N2499);
nor NOR3 (N3093, N3078, N535, N2671);
buf BUF1 (N3094, N3092);
and AND3 (N3095, N3077, N1851, N337);
nor NOR3 (N3096, N3090, N2556, N936);
xor XOR2 (N3097, N3091, N2981);
and AND4 (N3098, N3075, N1613, N1085, N1521);
or OR3 (N3099, N3089, N2281, N3038);
or OR3 (N3100, N3096, N3012, N225);
nor NOR3 (N3101, N3095, N1273, N1855);
buf BUF1 (N3102, N3099);
or OR2 (N3103, N3101, N2475);
not NOT1 (N3104, N3094);
buf BUF1 (N3105, N3103);
or OR4 (N3106, N3062, N2450, N2821, N624);
or OR2 (N3107, N3088, N2104);
and AND3 (N3108, N3107, N2661, N438);
buf BUF1 (N3109, N3093);
buf BUF1 (N3110, N3098);
or OR4 (N3111, N3102, N971, N704, N215);
not NOT1 (N3112, N3083);
buf BUF1 (N3113, N3104);
not NOT1 (N3114, N3111);
buf BUF1 (N3115, N3113);
xor XOR2 (N3116, N3097, N1364);
or OR4 (N3117, N3112, N723, N2096, N1858);
xor XOR2 (N3118, N3109, N1207);
nor NOR2 (N3119, N3100, N746);
nand NAND2 (N3120, N3115, N1071);
xor XOR2 (N3121, N3117, N2741);
xor XOR2 (N3122, N3105, N245);
xor XOR2 (N3123, N3118, N1481);
and AND4 (N3124, N3122, N1538, N1724, N2998);
nor NOR3 (N3125, N3124, N2674, N3026);
nand NAND3 (N3126, N3123, N3029, N2937);
buf BUF1 (N3127, N3121);
nand NAND2 (N3128, N3120, N1233);
and AND2 (N3129, N3127, N495);
nor NOR2 (N3130, N3110, N2012);
xor XOR2 (N3131, N3129, N1209);
buf BUF1 (N3132, N3130);
xor XOR2 (N3133, N3128, N25);
nor NOR2 (N3134, N3114, N1630);
or OR4 (N3135, N3132, N2916, N2006, N1894);
not NOT1 (N3136, N3116);
nor NOR4 (N3137, N3125, N873, N967, N2754);
nand NAND3 (N3138, N3137, N990, N1241);
or OR3 (N3139, N3136, N2370, N3);
buf BUF1 (N3140, N3135);
nor NOR3 (N3141, N3138, N2393, N1762);
not NOT1 (N3142, N3131);
nor NOR3 (N3143, N3140, N2567, N193);
not NOT1 (N3144, N3119);
or OR3 (N3145, N3144, N1176, N2269);
xor XOR2 (N3146, N3106, N979);
or OR3 (N3147, N3143, N241, N2484);
buf BUF1 (N3148, N3108);
nand NAND3 (N3149, N3142, N266, N232);
and AND2 (N3150, N3145, N1034);
or OR3 (N3151, N3150, N2872, N2582);
buf BUF1 (N3152, N3147);
and AND3 (N3153, N3148, N1859, N1773);
buf BUF1 (N3154, N3151);
xor XOR2 (N3155, N3149, N3017);
nor NOR4 (N3156, N3134, N2235, N1512, N820);
xor XOR2 (N3157, N3154, N811);
buf BUF1 (N3158, N3133);
and AND3 (N3159, N3156, N930, N2958);
nand NAND4 (N3160, N3158, N2788, N2579, N1895);
buf BUF1 (N3161, N3153);
not NOT1 (N3162, N3139);
buf BUF1 (N3163, N3159);
buf BUF1 (N3164, N3162);
nand NAND4 (N3165, N3160, N754, N2770, N513);
or OR2 (N3166, N3165, N2329);
and AND2 (N3167, N3146, N2154);
not NOT1 (N3168, N3161);
nor NOR2 (N3169, N3164, N1828);
nor NOR2 (N3170, N3166, N1382);
and AND2 (N3171, N3152, N893);
or OR2 (N3172, N3155, N2564);
and AND2 (N3173, N3126, N1380);
xor XOR2 (N3174, N3167, N2377);
and AND2 (N3175, N3157, N1582);
and AND3 (N3176, N3171, N1684, N1615);
not NOT1 (N3177, N3163);
or OR4 (N3178, N3141, N3155, N1441, N964);
nor NOR2 (N3179, N3177, N1621);
nor NOR4 (N3180, N3169, N771, N621, N1870);
nand NAND2 (N3181, N3174, N2478);
not NOT1 (N3182, N3170);
xor XOR2 (N3183, N3179, N2250);
xor XOR2 (N3184, N3173, N1154);
xor XOR2 (N3185, N3176, N755);
xor XOR2 (N3186, N3183, N2289);
nor NOR4 (N3187, N3180, N192, N1007, N57);
xor XOR2 (N3188, N3182, N2212);
buf BUF1 (N3189, N3181);
buf BUF1 (N3190, N3184);
nor NOR4 (N3191, N3188, N3043, N2805, N1787);
and AND3 (N3192, N3190, N144, N2788);
or OR2 (N3193, N3189, N643);
nor NOR3 (N3194, N3187, N1017, N2198);
not NOT1 (N3195, N3193);
or OR3 (N3196, N3168, N2763, N1823);
and AND3 (N3197, N3196, N2263, N3186);
buf BUF1 (N3198, N122);
xor XOR2 (N3199, N3172, N1453);
not NOT1 (N3200, N3194);
nand NAND4 (N3201, N3192, N2462, N3091, N486);
xor XOR2 (N3202, N3197, N395);
or OR2 (N3203, N3191, N2451);
xor XOR2 (N3204, N3202, N1210);
xor XOR2 (N3205, N3175, N2396);
not NOT1 (N3206, N3195);
and AND2 (N3207, N3199, N383);
nor NOR3 (N3208, N3198, N864, N821);
buf BUF1 (N3209, N3178);
buf BUF1 (N3210, N3204);
xor XOR2 (N3211, N3208, N2250);
nand NAND2 (N3212, N3205, N2652);
buf BUF1 (N3213, N3200);
nor NOR4 (N3214, N3213, N2811, N2079, N3119);
buf BUF1 (N3215, N3185);
or OR4 (N3216, N3209, N1975, N2020, N2418);
nor NOR4 (N3217, N3216, N1491, N2361, N1678);
and AND2 (N3218, N3214, N129);
nor NOR4 (N3219, N3210, N150, N248, N1737);
nor NOR2 (N3220, N3203, N1504);
buf BUF1 (N3221, N3218);
not NOT1 (N3222, N3206);
xor XOR2 (N3223, N3217, N1942);
xor XOR2 (N3224, N3223, N299);
and AND4 (N3225, N3224, N2873, N797, N625);
not NOT1 (N3226, N3225);
nand NAND3 (N3227, N3221, N1628, N2977);
nand NAND4 (N3228, N3219, N2816, N1312, N309);
xor XOR2 (N3229, N3228, N1780);
xor XOR2 (N3230, N3220, N2380);
and AND3 (N3231, N3207, N223, N1022);
xor XOR2 (N3232, N3227, N1462);
or OR4 (N3233, N3226, N1492, N2397, N65);
and AND4 (N3234, N3230, N3061, N1139, N1692);
or OR2 (N3235, N3234, N2703);
buf BUF1 (N3236, N3232);
or OR4 (N3237, N3215, N2980, N46, N2191);
buf BUF1 (N3238, N3229);
nand NAND4 (N3239, N3237, N2846, N2721, N2031);
not NOT1 (N3240, N3233);
nor NOR2 (N3241, N3239, N2503);
xor XOR2 (N3242, N3212, N1393);
xor XOR2 (N3243, N3211, N294);
or OR4 (N3244, N3222, N1656, N2354, N2686);
xor XOR2 (N3245, N3231, N2270);
nor NOR4 (N3246, N3236, N734, N2367, N1393);
xor XOR2 (N3247, N3240, N736);
and AND4 (N3248, N3242, N1298, N2484, N651);
or OR4 (N3249, N3245, N1941, N2300, N487);
or OR2 (N3250, N3241, N2226);
and AND3 (N3251, N3244, N67, N712);
or OR2 (N3252, N3238, N864);
buf BUF1 (N3253, N3252);
xor XOR2 (N3254, N3250, N2082);
or OR2 (N3255, N3249, N1212);
buf BUF1 (N3256, N3248);
or OR3 (N3257, N3255, N211, N2006);
and AND4 (N3258, N3235, N248, N1615, N2963);
nand NAND4 (N3259, N3257, N564, N2176, N71);
or OR2 (N3260, N3259, N141);
buf BUF1 (N3261, N3258);
not NOT1 (N3262, N3253);
and AND3 (N3263, N3254, N3164, N2322);
and AND3 (N3264, N3261, N455, N1031);
nor NOR2 (N3265, N3246, N3066);
buf BUF1 (N3266, N3256);
xor XOR2 (N3267, N3264, N2241);
not NOT1 (N3268, N3251);
nand NAND2 (N3269, N3262, N2041);
xor XOR2 (N3270, N3269, N1280);
nand NAND3 (N3271, N3267, N1876, N1192);
or OR4 (N3272, N3243, N2525, N2297, N1423);
and AND4 (N3273, N3268, N1762, N2317, N861);
or OR2 (N3274, N3201, N1636);
nor NOR3 (N3275, N3273, N1057, N1203);
nor NOR3 (N3276, N3266, N669, N3048);
and AND4 (N3277, N3271, N1313, N2345, N1122);
or OR3 (N3278, N3274, N2879, N1198);
nor NOR2 (N3279, N3276, N2314);
or OR4 (N3280, N3247, N979, N2264, N926);
not NOT1 (N3281, N3275);
buf BUF1 (N3282, N3278);
buf BUF1 (N3283, N3277);
nor NOR2 (N3284, N3281, N1631);
nor NOR2 (N3285, N3283, N86);
or OR3 (N3286, N3285, N1782, N2326);
and AND2 (N3287, N3270, N2007);
buf BUF1 (N3288, N3280);
xor XOR2 (N3289, N3282, N3177);
nor NOR4 (N3290, N3272, N865, N839, N2823);
and AND3 (N3291, N3289, N364, N3228);
nand NAND3 (N3292, N3290, N126, N561);
or OR3 (N3293, N3263, N948, N1140);
buf BUF1 (N3294, N3279);
buf BUF1 (N3295, N3288);
xor XOR2 (N3296, N3260, N2026);
or OR4 (N3297, N3295, N2088, N3223, N359);
buf BUF1 (N3298, N3286);
or OR2 (N3299, N3291, N575);
nor NOR3 (N3300, N3294, N1924, N2048);
not NOT1 (N3301, N3297);
nand NAND4 (N3302, N3298, N3253, N1225, N970);
buf BUF1 (N3303, N3299);
xor XOR2 (N3304, N3300, N3134);
nor NOR4 (N3305, N3304, N1706, N220, N474);
not NOT1 (N3306, N3303);
xor XOR2 (N3307, N3287, N768);
xor XOR2 (N3308, N3296, N916);
and AND2 (N3309, N3284, N754);
buf BUF1 (N3310, N3293);
and AND2 (N3311, N3265, N523);
xor XOR2 (N3312, N3305, N197);
and AND4 (N3313, N3310, N198, N1437, N1748);
xor XOR2 (N3314, N3307, N1991);
not NOT1 (N3315, N3309);
not NOT1 (N3316, N3306);
and AND4 (N3317, N3311, N458, N1084, N1037);
or OR4 (N3318, N3317, N2683, N240, N2511);
not NOT1 (N3319, N3313);
not NOT1 (N3320, N3314);
and AND3 (N3321, N3318, N3000, N183);
nand NAND3 (N3322, N3316, N1583, N3174);
xor XOR2 (N3323, N3319, N1691);
xor XOR2 (N3324, N3308, N1903);
nand NAND2 (N3325, N3323, N614);
and AND4 (N3326, N3292, N68, N595, N1409);
nor NOR4 (N3327, N3324, N2491, N1910, N489);
not NOT1 (N3328, N3325);
nor NOR2 (N3329, N3312, N1888);
nor NOR2 (N3330, N3301, N3174);
or OR2 (N3331, N3320, N3160);
not NOT1 (N3332, N3327);
buf BUF1 (N3333, N3331);
xor XOR2 (N3334, N3328, N453);
nand NAND2 (N3335, N3321, N2447);
or OR4 (N3336, N3326, N1612, N645, N2891);
buf BUF1 (N3337, N3315);
not NOT1 (N3338, N3333);
nand NAND2 (N3339, N3337, N2333);
nor NOR3 (N3340, N3334, N1710, N3272);
and AND4 (N3341, N3340, N2933, N2730, N2993);
nand NAND2 (N3342, N3322, N2277);
nor NOR4 (N3343, N3332, N2845, N3302, N1078);
buf BUF1 (N3344, N1581);
and AND3 (N3345, N3330, N1555, N2977);
nor NOR3 (N3346, N3329, N879, N2758);
and AND2 (N3347, N3345, N841);
nand NAND3 (N3348, N3336, N41, N624);
nand NAND4 (N3349, N3335, N3136, N1580, N2414);
buf BUF1 (N3350, N3349);
and AND4 (N3351, N3338, N3142, N1765, N287);
nor NOR4 (N3352, N3351, N1745, N555, N1723);
nand NAND2 (N3353, N3350, N1564);
nand NAND2 (N3354, N3339, N2352);
xor XOR2 (N3355, N3343, N2503);
nand NAND2 (N3356, N3352, N995);
buf BUF1 (N3357, N3354);
and AND4 (N3358, N3356, N3340, N3311, N1950);
or OR2 (N3359, N3347, N3263);
nor NOR2 (N3360, N3353, N1659);
xor XOR2 (N3361, N3346, N976);
and AND4 (N3362, N3344, N1872, N750, N2892);
or OR3 (N3363, N3362, N474, N1320);
buf BUF1 (N3364, N3342);
buf BUF1 (N3365, N3364);
nand NAND3 (N3366, N3358, N1036, N939);
xor XOR2 (N3367, N3359, N29);
buf BUF1 (N3368, N3341);
nand NAND2 (N3369, N3357, N2041);
not NOT1 (N3370, N3361);
and AND2 (N3371, N3368, N2476);
buf BUF1 (N3372, N3365);
and AND3 (N3373, N3371, N1541, N3115);
and AND2 (N3374, N3369, N2987);
nand NAND3 (N3375, N3355, N3084, N2868);
nand NAND2 (N3376, N3348, N619);
not NOT1 (N3377, N3374);
or OR3 (N3378, N3360, N3035, N3021);
nor NOR2 (N3379, N3378, N2414);
nor NOR2 (N3380, N3375, N1451);
and AND3 (N3381, N3373, N1713, N1370);
and AND2 (N3382, N3372, N941);
not NOT1 (N3383, N3379);
nand NAND4 (N3384, N3366, N1026, N2411, N383);
or OR3 (N3385, N3380, N1647, N919);
nor NOR2 (N3386, N3382, N1225);
nand NAND2 (N3387, N3367, N727);
nand NAND3 (N3388, N3387, N1248, N1707);
or OR3 (N3389, N3386, N3302, N1556);
or OR3 (N3390, N3363, N825, N1388);
and AND3 (N3391, N3377, N2599, N859);
not NOT1 (N3392, N3376);
not NOT1 (N3393, N3392);
xor XOR2 (N3394, N3388, N2220);
buf BUF1 (N3395, N3394);
buf BUF1 (N3396, N3383);
not NOT1 (N3397, N3381);
xor XOR2 (N3398, N3396, N3116);
or OR2 (N3399, N3395, N1233);
or OR2 (N3400, N3384, N2401);
xor XOR2 (N3401, N3391, N2786);
nor NOR3 (N3402, N3397, N3139, N1958);
buf BUF1 (N3403, N3399);
or OR2 (N3404, N3403, N1192);
nor NOR2 (N3405, N3370, N249);
nor NOR3 (N3406, N3398, N685, N2195);
or OR2 (N3407, N3402, N1545);
xor XOR2 (N3408, N3404, N2536);
or OR3 (N3409, N3390, N1646, N1571);
xor XOR2 (N3410, N3408, N2804);
nor NOR2 (N3411, N3406, N549);
not NOT1 (N3412, N3411);
not NOT1 (N3413, N3401);
nor NOR2 (N3414, N3393, N2065);
nand NAND3 (N3415, N3389, N2629, N1629);
and AND2 (N3416, N3407, N271);
xor XOR2 (N3417, N3410, N2792);
nor NOR2 (N3418, N3417, N2297);
nand NAND3 (N3419, N3413, N797, N3344);
and AND3 (N3420, N3412, N2833, N2179);
nor NOR2 (N3421, N3420, N558);
or OR4 (N3422, N3409, N911, N2176, N937);
nand NAND3 (N3423, N3385, N2417, N2058);
not NOT1 (N3424, N3400);
or OR3 (N3425, N3421, N3421, N2020);
or OR4 (N3426, N3405, N1846, N1382, N2538);
buf BUF1 (N3427, N3419);
nor NOR3 (N3428, N3424, N2290, N550);
and AND3 (N3429, N3416, N1859, N1540);
buf BUF1 (N3430, N3422);
not NOT1 (N3431, N3425);
or OR2 (N3432, N3415, N655);
nand NAND3 (N3433, N3414, N735, N591);
not NOT1 (N3434, N3418);
xor XOR2 (N3435, N3427, N848);
buf BUF1 (N3436, N3431);
xor XOR2 (N3437, N3436, N177);
or OR4 (N3438, N3429, N1659, N340, N2791);
nor NOR2 (N3439, N3438, N996);
xor XOR2 (N3440, N3423, N1044);
nor NOR2 (N3441, N3435, N971);
nor NOR4 (N3442, N3432, N3171, N2465, N544);
xor XOR2 (N3443, N3426, N548);
not NOT1 (N3444, N3428);
xor XOR2 (N3445, N3433, N1975);
not NOT1 (N3446, N3443);
nor NOR2 (N3447, N3437, N39);
nand NAND3 (N3448, N3444, N2198, N1907);
nand NAND2 (N3449, N3434, N1218);
xor XOR2 (N3450, N3448, N823);
buf BUF1 (N3451, N3442);
or OR3 (N3452, N3449, N706, N2863);
and AND3 (N3453, N3445, N2818, N133);
and AND4 (N3454, N3430, N912, N3010, N761);
nand NAND4 (N3455, N3452, N1406, N954, N3186);
or OR3 (N3456, N3455, N176, N2018);
not NOT1 (N3457, N3454);
and AND4 (N3458, N3457, N384, N3359, N646);
nand NAND2 (N3459, N3453, N2028);
not NOT1 (N3460, N3450);
not NOT1 (N3461, N3459);
xor XOR2 (N3462, N3460, N2458);
or OR4 (N3463, N3458, N1073, N2482, N1354);
xor XOR2 (N3464, N3446, N1169);
nor NOR2 (N3465, N3462, N2350);
or OR2 (N3466, N3463, N2111);
not NOT1 (N3467, N3441);
or OR2 (N3468, N3465, N1654);
nand NAND4 (N3469, N3466, N1621, N3232, N3049);
nor NOR3 (N3470, N3469, N267, N3051);
not NOT1 (N3471, N3456);
nand NAND3 (N3472, N3440, N1110, N39);
nand NAND2 (N3473, N3464, N2369);
and AND3 (N3474, N3470, N1184, N492);
not NOT1 (N3475, N3473);
buf BUF1 (N3476, N3472);
nand NAND2 (N3477, N3474, N2808);
xor XOR2 (N3478, N3471, N425);
or OR3 (N3479, N3476, N2499, N3027);
nand NAND2 (N3480, N3439, N1994);
nor NOR3 (N3481, N3451, N3394, N2970);
or OR2 (N3482, N3468, N2634);
buf BUF1 (N3483, N3478);
buf BUF1 (N3484, N3477);
not NOT1 (N3485, N3484);
buf BUF1 (N3486, N3447);
or OR4 (N3487, N3483, N1240, N403, N331);
buf BUF1 (N3488, N3487);
not NOT1 (N3489, N3485);
nand NAND3 (N3490, N3475, N1591, N1496);
xor XOR2 (N3491, N3490, N987);
nor NOR3 (N3492, N3467, N597, N2955);
not NOT1 (N3493, N3488);
and AND4 (N3494, N3489, N1400, N243, N1399);
or OR4 (N3495, N3491, N2586, N2485, N149);
or OR3 (N3496, N3493, N1871, N601);
and AND4 (N3497, N3482, N3015, N2201, N2503);
or OR4 (N3498, N3495, N3030, N342, N2502);
xor XOR2 (N3499, N3498, N1934);
not NOT1 (N3500, N3480);
nor NOR2 (N3501, N3486, N1447);
xor XOR2 (N3502, N3461, N691);
buf BUF1 (N3503, N3479);
nor NOR3 (N3504, N3500, N1749, N3266);
xor XOR2 (N3505, N3481, N2479);
or OR4 (N3506, N3494, N2447, N2068, N3031);
buf BUF1 (N3507, N3502);
nor NOR4 (N3508, N3505, N2568, N3244, N2026);
buf BUF1 (N3509, N3503);
nand NAND2 (N3510, N3504, N996);
or OR2 (N3511, N3496, N2889);
or OR2 (N3512, N3510, N553);
or OR4 (N3513, N3509, N78, N783, N2711);
and AND3 (N3514, N3508, N3264, N2866);
buf BUF1 (N3515, N3501);
xor XOR2 (N3516, N3514, N2329);
xor XOR2 (N3517, N3497, N255);
xor XOR2 (N3518, N3492, N813);
or OR3 (N3519, N3499, N94, N644);
buf BUF1 (N3520, N3513);
xor XOR2 (N3521, N3520, N2515);
buf BUF1 (N3522, N3517);
or OR3 (N3523, N3521, N1538, N3027);
or OR4 (N3524, N3512, N547, N365, N1825);
not NOT1 (N3525, N3507);
or OR4 (N3526, N3516, N1847, N1288, N637);
nand NAND3 (N3527, N3518, N238, N2577);
or OR2 (N3528, N3527, N3391);
not NOT1 (N3529, N3506);
nor NOR4 (N3530, N3523, N1808, N119, N2595);
xor XOR2 (N3531, N3524, N2837);
buf BUF1 (N3532, N3515);
not NOT1 (N3533, N3522);
and AND4 (N3534, N3526, N444, N1841, N786);
or OR2 (N3535, N3531, N3175);
or OR2 (N3536, N3511, N3294);
nand NAND4 (N3537, N3519, N2945, N2936, N2828);
xor XOR2 (N3538, N3537, N3373);
and AND3 (N3539, N3530, N2750, N2929);
or OR3 (N3540, N3538, N2128, N1685);
not NOT1 (N3541, N3536);
buf BUF1 (N3542, N3529);
nor NOR4 (N3543, N3542, N1508, N2673, N766);
xor XOR2 (N3544, N3528, N1592);
buf BUF1 (N3545, N3543);
buf BUF1 (N3546, N3541);
xor XOR2 (N3547, N3525, N807);
nor NOR4 (N3548, N3535, N3023, N675, N185);
nor NOR3 (N3549, N3546, N1725, N2177);
or OR2 (N3550, N3545, N599);
xor XOR2 (N3551, N3550, N3458);
not NOT1 (N3552, N3532);
buf BUF1 (N3553, N3540);
nor NOR2 (N3554, N3551, N3153);
nor NOR2 (N3555, N3539, N474);
buf BUF1 (N3556, N3555);
not NOT1 (N3557, N3534);
nor NOR3 (N3558, N3547, N1925, N898);
or OR4 (N3559, N3549, N3204, N195, N3442);
buf BUF1 (N3560, N3554);
xor XOR2 (N3561, N3533, N2033);
not NOT1 (N3562, N3561);
nand NAND4 (N3563, N3556, N507, N707, N1);
xor XOR2 (N3564, N3557, N995);
or OR3 (N3565, N3548, N212, N2019);
xor XOR2 (N3566, N3564, N423);
nand NAND4 (N3567, N3562, N3029, N2318, N3497);
or OR2 (N3568, N3566, N1866);
and AND4 (N3569, N3565, N1030, N1897, N3414);
buf BUF1 (N3570, N3559);
buf BUF1 (N3571, N3552);
or OR2 (N3572, N3553, N1242);
or OR4 (N3573, N3558, N3505, N2575, N1284);
xor XOR2 (N3574, N3569, N2331);
and AND2 (N3575, N3544, N612);
and AND2 (N3576, N3563, N1734);
buf BUF1 (N3577, N3576);
xor XOR2 (N3578, N3568, N1077);
or OR4 (N3579, N3574, N2952, N2472, N2026);
and AND2 (N3580, N3570, N1013);
buf BUF1 (N3581, N3571);
or OR2 (N3582, N3580, N483);
xor XOR2 (N3583, N3579, N1192);
buf BUF1 (N3584, N3573);
xor XOR2 (N3585, N3584, N1553);
or OR3 (N3586, N3560, N313, N2245);
not NOT1 (N3587, N3582);
nor NOR2 (N3588, N3578, N1183);
nor NOR4 (N3589, N3587, N1729, N2326, N1954);
nand NAND4 (N3590, N3586, N1354, N81, N1576);
nand NAND2 (N3591, N3581, N2207);
and AND2 (N3592, N3575, N989);
or OR2 (N3593, N3583, N810);
nor NOR4 (N3594, N3585, N1064, N347, N2296);
buf BUF1 (N3595, N3572);
nand NAND2 (N3596, N3567, N1485);
buf BUF1 (N3597, N3577);
or OR3 (N3598, N3595, N1779, N2509);
nor NOR2 (N3599, N3593, N1616);
and AND4 (N3600, N3594, N51, N1243, N163);
xor XOR2 (N3601, N3592, N626);
or OR4 (N3602, N3597, N2936, N2915, N2727);
xor XOR2 (N3603, N3599, N405);
nor NOR4 (N3604, N3591, N1115, N2453, N1362);
xor XOR2 (N3605, N3596, N214);
not NOT1 (N3606, N3602);
or OR3 (N3607, N3603, N625, N3155);
nor NOR2 (N3608, N3590, N2894);
not NOT1 (N3609, N3588);
nor NOR3 (N3610, N3601, N1748, N1719);
nand NAND3 (N3611, N3598, N3106, N3193);
nor NOR3 (N3612, N3609, N335, N2232);
xor XOR2 (N3613, N3589, N256);
not NOT1 (N3614, N3613);
not NOT1 (N3615, N3604);
xor XOR2 (N3616, N3605, N2130);
nor NOR2 (N3617, N3615, N2741);
not NOT1 (N3618, N3606);
nand NAND4 (N3619, N3612, N2751, N2405, N3300);
or OR3 (N3620, N3610, N51, N625);
buf BUF1 (N3621, N3607);
and AND3 (N3622, N3621, N617, N2734);
nor NOR2 (N3623, N3614, N3105);
buf BUF1 (N3624, N3616);
nand NAND4 (N3625, N3608, N2119, N770, N3482);
and AND3 (N3626, N3623, N802, N961);
nand NAND2 (N3627, N3617, N2900);
nor NOR2 (N3628, N3625, N3110);
not NOT1 (N3629, N3624);
xor XOR2 (N3630, N3626, N940);
nor NOR3 (N3631, N3630, N640, N1745);
buf BUF1 (N3632, N3611);
xor XOR2 (N3633, N3628, N673);
nor NOR3 (N3634, N3633, N860, N3579);
buf BUF1 (N3635, N3634);
buf BUF1 (N3636, N3635);
nor NOR3 (N3637, N3632, N2068, N2276);
xor XOR2 (N3638, N3622, N27);
or OR3 (N3639, N3618, N2719, N1019);
and AND3 (N3640, N3619, N1824, N1243);
nor NOR4 (N3641, N3627, N3572, N470, N355);
and AND3 (N3642, N3631, N273, N2741);
nor NOR3 (N3643, N3629, N451, N1771);
nor NOR2 (N3644, N3638, N271);
nand NAND3 (N3645, N3639, N3063, N1507);
not NOT1 (N3646, N3620);
buf BUF1 (N3647, N3600);
buf BUF1 (N3648, N3641);
xor XOR2 (N3649, N3644, N3648);
buf BUF1 (N3650, N3136);
nor NOR3 (N3651, N3649, N1, N217);
or OR4 (N3652, N3640, N536, N1788, N833);
buf BUF1 (N3653, N3651);
buf BUF1 (N3654, N3645);
and AND2 (N3655, N3653, N239);
buf BUF1 (N3656, N3636);
buf BUF1 (N3657, N3646);
and AND3 (N3658, N3642, N309, N1294);
nand NAND4 (N3659, N3657, N853, N493, N2780);
nand NAND4 (N3660, N3656, N2042, N323, N2610);
buf BUF1 (N3661, N3650);
nand NAND2 (N3662, N3658, N2926);
xor XOR2 (N3663, N3652, N1783);
and AND2 (N3664, N3659, N57);
or OR3 (N3665, N3664, N990, N2183);
nand NAND3 (N3666, N3643, N1181, N1449);
xor XOR2 (N3667, N3662, N2983);
buf BUF1 (N3668, N3661);
nor NOR3 (N3669, N3660, N2343, N1219);
or OR4 (N3670, N3669, N2883, N105, N1240);
xor XOR2 (N3671, N3668, N2197);
nor NOR4 (N3672, N3637, N1829, N154, N3206);
not NOT1 (N3673, N3647);
not NOT1 (N3674, N3670);
nand NAND2 (N3675, N3674, N2918);
and AND3 (N3676, N3663, N2479, N315);
nand NAND2 (N3677, N3654, N68);
nor NOR3 (N3678, N3665, N2721, N1708);
not NOT1 (N3679, N3671);
xor XOR2 (N3680, N3677, N1994);
and AND4 (N3681, N3676, N2162, N2731, N3382);
nand NAND2 (N3682, N3655, N700);
nand NAND4 (N3683, N3681, N886, N919, N144);
nand NAND2 (N3684, N3667, N3378);
nor NOR4 (N3685, N3682, N2107, N453, N1122);
or OR3 (N3686, N3685, N2029, N2650);
not NOT1 (N3687, N3679);
not NOT1 (N3688, N3687);
and AND3 (N3689, N3673, N1533, N2396);
nor NOR2 (N3690, N3675, N2216);
buf BUF1 (N3691, N3672);
xor XOR2 (N3692, N3666, N987);
and AND2 (N3693, N3680, N3684);
nor NOR4 (N3694, N277, N2820, N1653, N3222);
nor NOR4 (N3695, N3678, N2007, N731, N2995);
xor XOR2 (N3696, N3692, N3425);
buf BUF1 (N3697, N3691);
buf BUF1 (N3698, N3695);
nor NOR4 (N3699, N3696, N1829, N2925, N3509);
not NOT1 (N3700, N3688);
or OR4 (N3701, N3690, N1608, N3682, N3259);
and AND2 (N3702, N3698, N1743);
nor NOR4 (N3703, N3700, N1989, N384, N542);
and AND3 (N3704, N3699, N2892, N186);
nand NAND4 (N3705, N3686, N3587, N2178, N2505);
and AND4 (N3706, N3683, N2617, N336, N2726);
xor XOR2 (N3707, N3703, N1409);
and AND3 (N3708, N3706, N957, N2932);
or OR3 (N3709, N3707, N1447, N973);
xor XOR2 (N3710, N3702, N538);
not NOT1 (N3711, N3701);
buf BUF1 (N3712, N3711);
nand NAND2 (N3713, N3697, N404);
or OR3 (N3714, N3713, N535, N327);
nor NOR2 (N3715, N3714, N1430);
or OR4 (N3716, N3709, N280, N1787, N2592);
nand NAND4 (N3717, N3716, N1882, N1739, N3030);
xor XOR2 (N3718, N3708, N2486);
or OR2 (N3719, N3712, N88);
xor XOR2 (N3720, N3717, N2529);
buf BUF1 (N3721, N3693);
not NOT1 (N3722, N3719);
not NOT1 (N3723, N3721);
and AND2 (N3724, N3723, N2273);
nor NOR4 (N3725, N3722, N2191, N98, N1290);
buf BUF1 (N3726, N3704);
not NOT1 (N3727, N3724);
nand NAND3 (N3728, N3720, N1158, N2672);
or OR3 (N3729, N3710, N809, N2061);
buf BUF1 (N3730, N3727);
buf BUF1 (N3731, N3715);
nand NAND2 (N3732, N3689, N2865);
and AND4 (N3733, N3694, N3446, N636, N2130);
nor NOR3 (N3734, N3725, N2479, N222);
buf BUF1 (N3735, N3729);
or OR4 (N3736, N3735, N3079, N21, N564);
or OR3 (N3737, N3718, N1177, N2152);
and AND4 (N3738, N3736, N69, N272, N2361);
and AND2 (N3739, N3734, N1492);
or OR2 (N3740, N3739, N3480);
buf BUF1 (N3741, N3732);
xor XOR2 (N3742, N3738, N2302);
xor XOR2 (N3743, N3728, N3475);
nor NOR3 (N3744, N3733, N2331, N1609);
xor XOR2 (N3745, N3737, N3164);
or OR3 (N3746, N3744, N1437, N2025);
or OR3 (N3747, N3745, N2694, N1314);
or OR3 (N3748, N3730, N1405, N2846);
and AND4 (N3749, N3731, N3508, N2729, N2574);
or OR2 (N3750, N3749, N2208);
nand NAND2 (N3751, N3743, N3312);
nor NOR3 (N3752, N3705, N227, N1379);
nand NAND4 (N3753, N3742, N1732, N2379, N2189);
nor NOR2 (N3754, N3746, N2578);
nor NOR3 (N3755, N3726, N361, N543);
and AND4 (N3756, N3740, N115, N927, N813);
buf BUF1 (N3757, N3741);
buf BUF1 (N3758, N3747);
or OR2 (N3759, N3757, N3482);
nor NOR4 (N3760, N3751, N2050, N3432, N2568);
nor NOR3 (N3761, N3759, N1680, N2750);
xor XOR2 (N3762, N3753, N2678);
xor XOR2 (N3763, N3758, N2915);
not NOT1 (N3764, N3760);
or OR2 (N3765, N3750, N1030);
not NOT1 (N3766, N3754);
or OR2 (N3767, N3764, N2700);
or OR3 (N3768, N3767, N3508, N2720);
xor XOR2 (N3769, N3752, N1694);
and AND4 (N3770, N3763, N2349, N1633, N2019);
not NOT1 (N3771, N3761);
nand NAND2 (N3772, N3769, N3585);
xor XOR2 (N3773, N3768, N1406);
buf BUF1 (N3774, N3765);
or OR2 (N3775, N3772, N3667);
or OR2 (N3776, N3774, N2282);
or OR2 (N3777, N3775, N2957);
nor NOR4 (N3778, N3766, N1199, N1522, N336);
or OR2 (N3779, N3773, N2490);
nand NAND4 (N3780, N3776, N878, N1570, N3092);
and AND2 (N3781, N3778, N2472);
xor XOR2 (N3782, N3781, N2750);
nand NAND4 (N3783, N3777, N597, N1895, N2438);
xor XOR2 (N3784, N3755, N397);
xor XOR2 (N3785, N3771, N824);
or OR4 (N3786, N3785, N2000, N743, N200);
nor NOR2 (N3787, N3784, N1673);
or OR3 (N3788, N3782, N1828, N1661);
not NOT1 (N3789, N3780);
nor NOR3 (N3790, N3770, N2238, N3495);
buf BUF1 (N3791, N3788);
buf BUF1 (N3792, N3783);
buf BUF1 (N3793, N3786);
xor XOR2 (N3794, N3792, N1098);
or OR4 (N3795, N3789, N3195, N1053, N2883);
nor NOR4 (N3796, N3793, N518, N652, N3527);
or OR4 (N3797, N3794, N942, N645, N3698);
xor XOR2 (N3798, N3762, N118);
nand NAND2 (N3799, N3798, N1946);
not NOT1 (N3800, N3748);
or OR3 (N3801, N3800, N3543, N695);
nand NAND3 (N3802, N3799, N2074, N1038);
or OR4 (N3803, N3797, N848, N2210, N1505);
xor XOR2 (N3804, N3791, N3336);
nor NOR2 (N3805, N3756, N1141);
nand NAND4 (N3806, N3803, N921, N2905, N1052);
and AND3 (N3807, N3802, N116, N29);
not NOT1 (N3808, N3790);
buf BUF1 (N3809, N3787);
and AND3 (N3810, N3806, N3194, N717);
buf BUF1 (N3811, N3809);
nor NOR3 (N3812, N3796, N2292, N3703);
xor XOR2 (N3813, N3805, N2945);
or OR4 (N3814, N3801, N569, N716, N1529);
or OR2 (N3815, N3795, N1050);
not NOT1 (N3816, N3810);
buf BUF1 (N3817, N3815);
buf BUF1 (N3818, N3814);
xor XOR2 (N3819, N3818, N1490);
xor XOR2 (N3820, N3808, N3104);
nand NAND3 (N3821, N3804, N1758, N1856);
nand NAND3 (N3822, N3816, N3, N1290);
nor NOR2 (N3823, N3807, N2637);
nor NOR2 (N3824, N3779, N1900);
nor NOR2 (N3825, N3817, N2615);
nor NOR3 (N3826, N3812, N2762, N2039);
buf BUF1 (N3827, N3826);
and AND2 (N3828, N3821, N2224);
nor NOR3 (N3829, N3824, N3486, N701);
not NOT1 (N3830, N3813);
buf BUF1 (N3831, N3823);
not NOT1 (N3832, N3827);
not NOT1 (N3833, N3822);
not NOT1 (N3834, N3811);
nand NAND2 (N3835, N3832, N1607);
or OR4 (N3836, N3834, N623, N3360, N3519);
xor XOR2 (N3837, N3828, N2582);
nand NAND4 (N3838, N3833, N1536, N1940, N3254);
nor NOR3 (N3839, N3825, N2268, N862);
nor NOR4 (N3840, N3839, N2028, N1044, N884);
xor XOR2 (N3841, N3836, N3677);
or OR2 (N3842, N3831, N386);
and AND3 (N3843, N3840, N3667, N3306);
xor XOR2 (N3844, N3837, N2267);
buf BUF1 (N3845, N3843);
nor NOR2 (N3846, N3830, N575);
buf BUF1 (N3847, N3845);
xor XOR2 (N3848, N3838, N3065);
not NOT1 (N3849, N3819);
buf BUF1 (N3850, N3842);
or OR4 (N3851, N3835, N260, N774, N3446);
buf BUF1 (N3852, N3841);
buf BUF1 (N3853, N3848);
or OR2 (N3854, N3844, N174);
xor XOR2 (N3855, N3846, N3025);
xor XOR2 (N3856, N3849, N3655);
or OR2 (N3857, N3847, N3047);
xor XOR2 (N3858, N3852, N2105);
nor NOR2 (N3859, N3858, N3823);
or OR3 (N3860, N3854, N892, N3646);
nor NOR2 (N3861, N3820, N3099);
nor NOR4 (N3862, N3855, N1479, N3657, N1047);
and AND4 (N3863, N3861, N3814, N1802, N875);
nor NOR3 (N3864, N3862, N1569, N2372);
or OR2 (N3865, N3860, N3318);
or OR3 (N3866, N3851, N2660, N2682);
buf BUF1 (N3867, N3850);
xor XOR2 (N3868, N3829, N2886);
not NOT1 (N3869, N3868);
not NOT1 (N3870, N3866);
nand NAND3 (N3871, N3867, N3834, N540);
buf BUF1 (N3872, N3853);
not NOT1 (N3873, N3863);
or OR3 (N3874, N3856, N1960, N3546);
xor XOR2 (N3875, N3871, N446);
not NOT1 (N3876, N3864);
xor XOR2 (N3877, N3872, N2788);
and AND4 (N3878, N3876, N1952, N615, N2626);
not NOT1 (N3879, N3865);
nand NAND3 (N3880, N3878, N2094, N1349);
and AND3 (N3881, N3870, N3056, N2542);
and AND3 (N3882, N3880, N3224, N149);
buf BUF1 (N3883, N3882);
buf BUF1 (N3884, N3869);
or OR3 (N3885, N3857, N504, N3467);
xor XOR2 (N3886, N3881, N359);
nor NOR2 (N3887, N3873, N2450);
not NOT1 (N3888, N3887);
nor NOR4 (N3889, N3875, N1058, N1987, N613);
nor NOR3 (N3890, N3877, N3418, N1793);
xor XOR2 (N3891, N3879, N2578);
xor XOR2 (N3892, N3885, N2608);
and AND3 (N3893, N3889, N1689, N2743);
buf BUF1 (N3894, N3891);
nand NAND2 (N3895, N3893, N3693);
nand NAND2 (N3896, N3890, N2167);
xor XOR2 (N3897, N3896, N1553);
nand NAND2 (N3898, N3892, N2166);
nand NAND3 (N3899, N3883, N3131, N51);
nor NOR4 (N3900, N3886, N1471, N3281, N3341);
nand NAND3 (N3901, N3874, N1821, N1284);
xor XOR2 (N3902, N3884, N3678);
nand NAND4 (N3903, N3898, N3037, N3342, N538);
nand NAND4 (N3904, N3903, N3843, N3824, N2074);
not NOT1 (N3905, N3904);
nand NAND3 (N3906, N3888, N1630, N475);
nand NAND2 (N3907, N3900, N688);
xor XOR2 (N3908, N3897, N1200);
or OR2 (N3909, N3894, N2183);
nor NOR2 (N3910, N3906, N3494);
not NOT1 (N3911, N3905);
nor NOR4 (N3912, N3908, N521, N3739, N3300);
nor NOR3 (N3913, N3911, N1954, N3284);
and AND3 (N3914, N3895, N2001, N657);
nand NAND2 (N3915, N3912, N894);
buf BUF1 (N3916, N3899);
not NOT1 (N3917, N3901);
and AND4 (N3918, N3907, N93, N3171, N3255);
and AND4 (N3919, N3914, N1324, N596, N1153);
buf BUF1 (N3920, N3918);
nand NAND4 (N3921, N3859, N878, N2144, N1448);
nor NOR4 (N3922, N3913, N370, N3411, N2155);
buf BUF1 (N3923, N3916);
nor NOR4 (N3924, N3917, N3093, N2430, N3769);
or OR2 (N3925, N3919, N3373);
xor XOR2 (N3926, N3924, N3138);
and AND2 (N3927, N3902, N2925);
buf BUF1 (N3928, N3925);
not NOT1 (N3929, N3920);
nor NOR4 (N3930, N3909, N1801, N1010, N2262);
and AND3 (N3931, N3929, N3463, N686);
and AND2 (N3932, N3910, N3710);
not NOT1 (N3933, N3923);
xor XOR2 (N3934, N3915, N3752);
buf BUF1 (N3935, N3928);
nand NAND2 (N3936, N3933, N3018);
nand NAND2 (N3937, N3935, N2475);
nand NAND4 (N3938, N3922, N1323, N927, N3110);
buf BUF1 (N3939, N3938);
not NOT1 (N3940, N3936);
buf BUF1 (N3941, N3930);
not NOT1 (N3942, N3932);
nand NAND4 (N3943, N3939, N589, N2807, N3603);
nand NAND3 (N3944, N3926, N2640, N2192);
or OR4 (N3945, N3937, N213, N1053, N846);
or OR4 (N3946, N3931, N3034, N1874, N1480);
xor XOR2 (N3947, N3942, N3686);
and AND3 (N3948, N3945, N1879, N276);
and AND3 (N3949, N3943, N3013, N301);
not NOT1 (N3950, N3948);
buf BUF1 (N3951, N3921);
nand NAND3 (N3952, N3940, N2560, N1550);
not NOT1 (N3953, N3947);
and AND2 (N3954, N3941, N1552);
nor NOR2 (N3955, N3950, N30);
nor NOR4 (N3956, N3955, N1660, N2826, N164);
buf BUF1 (N3957, N3934);
and AND3 (N3958, N3927, N411, N2157);
nand NAND2 (N3959, N3953, N1942);
not NOT1 (N3960, N3952);
and AND3 (N3961, N3954, N402, N3883);
and AND4 (N3962, N3944, N1113, N1430, N791);
nor NOR2 (N3963, N3959, N1302);
not NOT1 (N3964, N3960);
nor NOR3 (N3965, N3951, N2733, N2403);
xor XOR2 (N3966, N3961, N2862);
not NOT1 (N3967, N3946);
xor XOR2 (N3968, N3965, N2203);
xor XOR2 (N3969, N3964, N1374);
nand NAND3 (N3970, N3962, N1295, N2606);
or OR4 (N3971, N3968, N3949, N253, N2431);
nor NOR3 (N3972, N3413, N2950, N2780);
buf BUF1 (N3973, N3957);
buf BUF1 (N3974, N3971);
nor NOR4 (N3975, N3966, N2307, N606, N1188);
xor XOR2 (N3976, N3974, N1875);
and AND3 (N3977, N3956, N2376, N3469);
not NOT1 (N3978, N3976);
nand NAND3 (N3979, N3963, N1196, N3240);
and AND2 (N3980, N3977, N996);
nand NAND3 (N3981, N3978, N1126, N1353);
and AND3 (N3982, N3970, N1826, N474);
nand NAND4 (N3983, N3958, N2531, N2820, N411);
nor NOR3 (N3984, N3982, N674, N1779);
or OR2 (N3985, N3969, N2581);
nand NAND2 (N3986, N3981, N2124);
or OR2 (N3987, N3975, N471);
or OR4 (N3988, N3983, N1363, N3070, N2675);
or OR3 (N3989, N3984, N3931, N1468);
and AND3 (N3990, N3980, N787, N2831);
nand NAND3 (N3991, N3986, N3735, N1894);
and AND4 (N3992, N3987, N2340, N2228, N3304);
or OR2 (N3993, N3990, N1577);
not NOT1 (N3994, N3985);
nand NAND4 (N3995, N3972, N207, N2801, N3402);
nor NOR2 (N3996, N3994, N908);
nor NOR2 (N3997, N3993, N2688);
and AND2 (N3998, N3995, N500);
nor NOR3 (N3999, N3989, N2441, N1540);
or OR3 (N4000, N3992, N1889, N3228);
and AND2 (N4001, N3973, N963);
and AND4 (N4002, N3988, N1022, N1102, N3028);
and AND4 (N4003, N3991, N2588, N3808, N3639);
nand NAND2 (N4004, N4003, N2914);
xor XOR2 (N4005, N3967, N3529);
nand NAND2 (N4006, N4005, N2500);
and AND3 (N4007, N3999, N3542, N3178);
or OR3 (N4008, N3996, N479, N1168);
xor XOR2 (N4009, N3979, N2671);
buf BUF1 (N4010, N3997);
nand NAND4 (N4011, N4007, N1501, N1257, N837);
not NOT1 (N4012, N4011);
or OR2 (N4013, N4012, N1385);
not NOT1 (N4014, N4004);
not NOT1 (N4015, N4009);
nor NOR4 (N4016, N4000, N1175, N1164, N2801);
and AND4 (N4017, N4006, N382, N814, N1823);
xor XOR2 (N4018, N4002, N3839);
buf BUF1 (N4019, N4017);
or OR3 (N4020, N4016, N496, N3953);
and AND3 (N4021, N4014, N2635, N610);
nor NOR3 (N4022, N4019, N2028, N3516);
buf BUF1 (N4023, N4018);
nand NAND2 (N4024, N4013, N3233);
buf BUF1 (N4025, N4001);
buf BUF1 (N4026, N4010);
nor NOR2 (N4027, N4020, N1620);
nor NOR2 (N4028, N4021, N2241);
nor NOR4 (N4029, N4015, N3857, N1727, N568);
xor XOR2 (N4030, N4008, N1996);
nor NOR2 (N4031, N4028, N1593);
or OR2 (N4032, N4025, N420);
or OR3 (N4033, N4031, N3015, N1621);
buf BUF1 (N4034, N4030);
xor XOR2 (N4035, N4023, N1282);
nand NAND2 (N4036, N4024, N40);
not NOT1 (N4037, N4022);
and AND3 (N4038, N4027, N3736, N2569);
and AND3 (N4039, N4029, N1943, N1085);
xor XOR2 (N4040, N4034, N2353);
or OR2 (N4041, N4026, N2349);
buf BUF1 (N4042, N4039);
xor XOR2 (N4043, N4042, N1521);
nand NAND3 (N4044, N4038, N3830, N2948);
xor XOR2 (N4045, N3998, N164);
buf BUF1 (N4046, N4037);
not NOT1 (N4047, N4033);
xor XOR2 (N4048, N4047, N1493);
xor XOR2 (N4049, N4046, N3267);
not NOT1 (N4050, N4043);
xor XOR2 (N4051, N4045, N2193);
and AND3 (N4052, N4048, N2354, N1445);
nor NOR4 (N4053, N4036, N3587, N2364, N2658);
xor XOR2 (N4054, N4049, N2336);
nor NOR4 (N4055, N4032, N2600, N3484, N3266);
and AND2 (N4056, N4050, N3683);
and AND4 (N4057, N4044, N3134, N3007, N2498);
not NOT1 (N4058, N4052);
and AND3 (N4059, N4041, N2131, N2857);
or OR4 (N4060, N4059, N3665, N786, N3193);
nand NAND4 (N4061, N4054, N2598, N3147, N3790);
or OR2 (N4062, N4040, N2966);
nor NOR3 (N4063, N4057, N913, N3042);
not NOT1 (N4064, N4053);
not NOT1 (N4065, N4063);
or OR2 (N4066, N4058, N404);
nand NAND4 (N4067, N4066, N2340, N3382, N2254);
nand NAND3 (N4068, N4067, N4052, N2627);
and AND2 (N4069, N4065, N1734);
not NOT1 (N4070, N4064);
nand NAND3 (N4071, N4056, N1353, N1529);
and AND4 (N4072, N4055, N1962, N2053, N953);
buf BUF1 (N4073, N4069);
or OR4 (N4074, N4062, N3972, N1216, N2994);
or OR3 (N4075, N4061, N545, N2667);
xor XOR2 (N4076, N4051, N1185);
or OR4 (N4077, N4035, N1609, N2365, N1934);
nand NAND3 (N4078, N4070, N3674, N1130);
buf BUF1 (N4079, N4072);
nor NOR4 (N4080, N4073, N2265, N736, N3102);
not NOT1 (N4081, N4068);
not NOT1 (N4082, N4076);
buf BUF1 (N4083, N4074);
not NOT1 (N4084, N4081);
xor XOR2 (N4085, N4077, N208);
buf BUF1 (N4086, N4060);
nor NOR4 (N4087, N4084, N167, N2744, N569);
nand NAND3 (N4088, N4071, N3181, N1440);
not NOT1 (N4089, N4078);
xor XOR2 (N4090, N4088, N1135);
xor XOR2 (N4091, N4089, N95);
xor XOR2 (N4092, N4079, N2193);
not NOT1 (N4093, N4086);
nor NOR4 (N4094, N4080, N1927, N32, N950);
xor XOR2 (N4095, N4087, N3573);
or OR4 (N4096, N4093, N4086, N478, N2619);
and AND3 (N4097, N4083, N705, N2937);
xor XOR2 (N4098, N4094, N2485);
nand NAND3 (N4099, N4091, N1651, N889);
buf BUF1 (N4100, N4085);
not NOT1 (N4101, N4075);
and AND2 (N4102, N4098, N1508);
and AND3 (N4103, N4102, N2026, N3433);
not NOT1 (N4104, N4099);
xor XOR2 (N4105, N4104, N558);
xor XOR2 (N4106, N4100, N1439);
xor XOR2 (N4107, N4101, N610);
not NOT1 (N4108, N4105);
or OR3 (N4109, N4095, N2075, N4051);
buf BUF1 (N4110, N4103);
nor NOR4 (N4111, N4090, N636, N3865, N1082);
buf BUF1 (N4112, N4108);
buf BUF1 (N4113, N4097);
xor XOR2 (N4114, N4112, N2937);
and AND4 (N4115, N4109, N746, N359, N1730);
or OR3 (N4116, N4096, N2857, N275);
not NOT1 (N4117, N4114);
and AND3 (N4118, N4111, N3969, N2441);
nand NAND2 (N4119, N4117, N2537);
and AND2 (N4120, N4110, N1743);
and AND3 (N4121, N4107, N685, N3984);
not NOT1 (N4122, N4082);
and AND4 (N4123, N4121, N295, N3632, N1345);
and AND2 (N4124, N4123, N1173);
and AND2 (N4125, N4124, N3290);
or OR4 (N4126, N4122, N709, N47, N3258);
or OR2 (N4127, N4106, N1457);
or OR4 (N4128, N4125, N636, N3621, N793);
xor XOR2 (N4129, N4092, N991);
nor NOR4 (N4130, N4113, N1825, N2212, N825);
buf BUF1 (N4131, N4127);
buf BUF1 (N4132, N4120);
not NOT1 (N4133, N4118);
nand NAND2 (N4134, N4128, N1222);
nor NOR3 (N4135, N4129, N350, N3509);
xor XOR2 (N4136, N4119, N3559);
nand NAND2 (N4137, N4136, N3730);
xor XOR2 (N4138, N4115, N1246);
not NOT1 (N4139, N4134);
xor XOR2 (N4140, N4138, N1924);
xor XOR2 (N4141, N4140, N2421);
buf BUF1 (N4142, N4133);
xor XOR2 (N4143, N4137, N504);
buf BUF1 (N4144, N4142);
xor XOR2 (N4145, N4143, N1370);
nand NAND3 (N4146, N4141, N1548, N1647);
nand NAND2 (N4147, N4131, N979);
nand NAND2 (N4148, N4116, N1121);
or OR2 (N4149, N4147, N850);
buf BUF1 (N4150, N4132);
nand NAND3 (N4151, N4149, N670, N3295);
buf BUF1 (N4152, N4148);
nand NAND3 (N4153, N4151, N2644, N2310);
xor XOR2 (N4154, N4146, N1870);
and AND3 (N4155, N4145, N635, N1488);
or OR3 (N4156, N4130, N4085, N1163);
buf BUF1 (N4157, N4155);
and AND4 (N4158, N4126, N2254, N199, N3423);
and AND3 (N4159, N4135, N2413, N977);
or OR3 (N4160, N4154, N1654, N3023);
buf BUF1 (N4161, N4144);
or OR3 (N4162, N4139, N4146, N2725);
or OR4 (N4163, N4156, N3168, N2078, N2983);
buf BUF1 (N4164, N4153);
nand NAND2 (N4165, N4163, N3584);
not NOT1 (N4166, N4152);
and AND3 (N4167, N4165, N2676, N1584);
nand NAND2 (N4168, N4164, N2438);
or OR3 (N4169, N4166, N1062, N1860);
buf BUF1 (N4170, N4159);
and AND2 (N4171, N4168, N3330);
nor NOR4 (N4172, N4171, N4168, N3664, N932);
or OR3 (N4173, N4150, N3512, N1643);
not NOT1 (N4174, N4167);
buf BUF1 (N4175, N4161);
xor XOR2 (N4176, N4157, N1015);
xor XOR2 (N4177, N4158, N1834);
or OR4 (N4178, N4175, N3390, N2705, N3875);
xor XOR2 (N4179, N4174, N3257);
nand NAND3 (N4180, N4170, N1038, N943);
xor XOR2 (N4181, N4179, N699);
nand NAND3 (N4182, N4172, N4026, N3222);
or OR4 (N4183, N4162, N2621, N1557, N3596);
nor NOR2 (N4184, N4176, N3020);
or OR3 (N4185, N4169, N3252, N2783);
or OR3 (N4186, N4182, N2556, N3317);
nand NAND3 (N4187, N4186, N3023, N3603);
not NOT1 (N4188, N4173);
nor NOR4 (N4189, N4180, N3012, N2566, N759);
xor XOR2 (N4190, N4160, N4079);
and AND3 (N4191, N4184, N616, N1076);
and AND2 (N4192, N4188, N74);
nor NOR2 (N4193, N4189, N1120);
not NOT1 (N4194, N4185);
nand NAND3 (N4195, N4190, N3879, N3420);
xor XOR2 (N4196, N4187, N3802);
xor XOR2 (N4197, N4181, N893);
nor NOR3 (N4198, N4177, N3477, N1825);
not NOT1 (N4199, N4178);
not NOT1 (N4200, N4183);
nor NOR2 (N4201, N4198, N3709);
buf BUF1 (N4202, N4201);
nand NAND4 (N4203, N4196, N3319, N3702, N3447);
not NOT1 (N4204, N4202);
or OR4 (N4205, N4194, N2163, N1347, N1124);
and AND2 (N4206, N4191, N835);
not NOT1 (N4207, N4197);
nor NOR3 (N4208, N4205, N527, N454);
xor XOR2 (N4209, N4206, N2876);
or OR4 (N4210, N4203, N3170, N1002, N2296);
nand NAND3 (N4211, N4193, N2729, N1619);
buf BUF1 (N4212, N4210);
or OR3 (N4213, N4204, N2419, N2415);
and AND4 (N4214, N4192, N721, N1485, N66);
xor XOR2 (N4215, N4200, N1966);
buf BUF1 (N4216, N4195);
nand NAND4 (N4217, N4199, N3460, N1367, N750);
buf BUF1 (N4218, N4212);
nand NAND2 (N4219, N4208, N2470);
nor NOR3 (N4220, N4216, N4059, N3147);
xor XOR2 (N4221, N4220, N1667);
and AND4 (N4222, N4211, N3129, N1264, N354);
or OR2 (N4223, N4214, N3167);
and AND4 (N4224, N4209, N774, N1939, N3928);
nor NOR4 (N4225, N4224, N480, N1670, N1406);
or OR3 (N4226, N4215, N897, N2808);
nand NAND3 (N4227, N4218, N3390, N1618);
and AND4 (N4228, N4221, N2820, N2624, N262);
nor NOR3 (N4229, N4223, N2726, N784);
xor XOR2 (N4230, N4222, N3792);
xor XOR2 (N4231, N4230, N3883);
nand NAND3 (N4232, N4225, N3020, N1875);
or OR4 (N4233, N4228, N3854, N900, N3340);
not NOT1 (N4234, N4227);
not NOT1 (N4235, N4207);
xor XOR2 (N4236, N4231, N2434);
nor NOR3 (N4237, N4219, N3987, N459);
nand NAND2 (N4238, N4233, N1387);
not NOT1 (N4239, N4229);
buf BUF1 (N4240, N4213);
and AND2 (N4241, N4240, N1244);
and AND3 (N4242, N4234, N1396, N4074);
not NOT1 (N4243, N4242);
xor XOR2 (N4244, N4239, N474);
nand NAND4 (N4245, N4244, N3700, N234, N1262);
and AND4 (N4246, N4237, N1955, N2428, N3482);
xor XOR2 (N4247, N4217, N3397);
nor NOR3 (N4248, N4243, N576, N3508);
buf BUF1 (N4249, N4247);
buf BUF1 (N4250, N4235);
nand NAND4 (N4251, N4226, N674, N2145, N1474);
nand NAND3 (N4252, N4250, N2350, N2780);
not NOT1 (N4253, N4241);
buf BUF1 (N4254, N4238);
buf BUF1 (N4255, N4246);
not NOT1 (N4256, N4251);
not NOT1 (N4257, N4236);
nor NOR3 (N4258, N4256, N1133, N362);
or OR3 (N4259, N4245, N1455, N1853);
and AND3 (N4260, N4249, N471, N3360);
not NOT1 (N4261, N4254);
not NOT1 (N4262, N4253);
and AND3 (N4263, N4255, N3283, N2580);
nor NOR3 (N4264, N4261, N1242, N2572);
xor XOR2 (N4265, N4259, N16);
and AND2 (N4266, N4252, N1466);
not NOT1 (N4267, N4258);
or OR2 (N4268, N4232, N4248);
xor XOR2 (N4269, N4119, N89);
buf BUF1 (N4270, N4262);
nor NOR2 (N4271, N4264, N2232);
xor XOR2 (N4272, N4260, N44);
nand NAND2 (N4273, N4271, N141);
xor XOR2 (N4274, N4263, N291);
not NOT1 (N4275, N4268);
nor NOR2 (N4276, N4275, N2749);
nand NAND4 (N4277, N4274, N1678, N1518, N3454);
xor XOR2 (N4278, N4272, N1424);
nor NOR4 (N4279, N4269, N3595, N2761, N1667);
and AND2 (N4280, N4257, N982);
xor XOR2 (N4281, N4266, N2888);
or OR4 (N4282, N4270, N3106, N2056, N1535);
buf BUF1 (N4283, N4265);
nor NOR3 (N4284, N4267, N3936, N3548);
buf BUF1 (N4285, N4279);
nand NAND4 (N4286, N4277, N4265, N3854, N3910);
buf BUF1 (N4287, N4278);
and AND3 (N4288, N4285, N1248, N2339);
xor XOR2 (N4289, N4288, N703);
buf BUF1 (N4290, N4284);
nand NAND4 (N4291, N4282, N2452, N3757, N877);
not NOT1 (N4292, N4273);
and AND3 (N4293, N4290, N1822, N3392);
not NOT1 (N4294, N4292);
nand NAND4 (N4295, N4289, N3209, N2005, N2264);
or OR4 (N4296, N4287, N2928, N977, N2593);
xor XOR2 (N4297, N4281, N3937);
nor NOR2 (N4298, N4276, N2133);
nor NOR3 (N4299, N4297, N860, N3035);
nor NOR4 (N4300, N4293, N1892, N1831, N513);
or OR3 (N4301, N4294, N562, N197);
and AND3 (N4302, N4283, N1129, N948);
buf BUF1 (N4303, N4302);
buf BUF1 (N4304, N4295);
or OR3 (N4305, N4280, N2211, N3258);
and AND2 (N4306, N4298, N511);
nor NOR4 (N4307, N4299, N3264, N2062, N1617);
xor XOR2 (N4308, N4296, N2583);
not NOT1 (N4309, N4304);
nor NOR2 (N4310, N4303, N2262);
not NOT1 (N4311, N4300);
or OR3 (N4312, N4305, N2358, N3684);
buf BUF1 (N4313, N4286);
not NOT1 (N4314, N4310);
not NOT1 (N4315, N4301);
or OR2 (N4316, N4291, N1372);
or OR4 (N4317, N4316, N3411, N2759, N738);
not NOT1 (N4318, N4317);
and AND2 (N4319, N4311, N2643);
nand NAND2 (N4320, N4312, N1426);
or OR3 (N4321, N4319, N3756, N3146);
nand NAND4 (N4322, N4320, N2307, N3412, N1311);
nand NAND4 (N4323, N4315, N1399, N1712, N3990);
xor XOR2 (N4324, N4322, N41);
and AND2 (N4325, N4324, N4310);
xor XOR2 (N4326, N4325, N1982);
nand NAND3 (N4327, N4313, N321, N4079);
and AND3 (N4328, N4309, N2577, N2769);
nand NAND2 (N4329, N4314, N3594);
nand NAND3 (N4330, N4323, N1831, N4180);
not NOT1 (N4331, N4330);
nand NAND2 (N4332, N4306, N2024);
nand NAND4 (N4333, N4331, N2707, N3108, N2201);
nand NAND2 (N4334, N4307, N4123);
nand NAND3 (N4335, N4329, N1004, N2263);
or OR2 (N4336, N4318, N2517);
xor XOR2 (N4337, N4327, N2440);
xor XOR2 (N4338, N4336, N2803);
buf BUF1 (N4339, N4337);
and AND3 (N4340, N4335, N4172, N3927);
or OR2 (N4341, N4326, N1323);
not NOT1 (N4342, N4339);
not NOT1 (N4343, N4338);
nor NOR2 (N4344, N4332, N3826);
nand NAND2 (N4345, N4340, N3935);
not NOT1 (N4346, N4334);
nand NAND4 (N4347, N4321, N2144, N3323, N673);
and AND3 (N4348, N4342, N1278, N2071);
xor XOR2 (N4349, N4348, N2209);
buf BUF1 (N4350, N4349);
buf BUF1 (N4351, N4350);
not NOT1 (N4352, N4308);
nor NOR3 (N4353, N4345, N3578, N2645);
nand NAND3 (N4354, N4333, N1597, N885);
nand NAND3 (N4355, N4346, N3110, N182);
nor NOR4 (N4356, N4347, N3566, N2100, N2855);
or OR2 (N4357, N4341, N340);
nand NAND4 (N4358, N4357, N3003, N2416, N3987);
nand NAND4 (N4359, N4354, N1084, N1979, N2292);
buf BUF1 (N4360, N4356);
or OR2 (N4361, N4343, N1264);
not NOT1 (N4362, N4360);
and AND4 (N4363, N4361, N602, N2091, N1518);
nand NAND2 (N4364, N4358, N2989);
and AND3 (N4365, N4364, N3926, N13);
buf BUF1 (N4366, N4355);
not NOT1 (N4367, N4344);
xor XOR2 (N4368, N4351, N2641);
xor XOR2 (N4369, N4352, N2703);
and AND3 (N4370, N4359, N3155, N2881);
buf BUF1 (N4371, N4368);
or OR4 (N4372, N4370, N2657, N2586, N4076);
not NOT1 (N4373, N4371);
nand NAND2 (N4374, N4365, N2237);
nand NAND4 (N4375, N4369, N3571, N1158, N3829);
not NOT1 (N4376, N4363);
nor NOR2 (N4377, N4367, N1554);
nand NAND3 (N4378, N4375, N2269, N2106);
xor XOR2 (N4379, N4378, N3228);
and AND2 (N4380, N4353, N4195);
and AND3 (N4381, N4373, N1483, N502);
nor NOR2 (N4382, N4362, N2171);
not NOT1 (N4383, N4379);
buf BUF1 (N4384, N4381);
or OR2 (N4385, N4383, N2327);
nor NOR2 (N4386, N4380, N4229);
nand NAND4 (N4387, N4374, N4100, N3247, N2083);
and AND4 (N4388, N4384, N2076, N2593, N3054);
and AND3 (N4389, N4386, N1519, N2830);
xor XOR2 (N4390, N4372, N3501);
or OR3 (N4391, N4385, N2493, N75);
and AND2 (N4392, N4377, N3336);
xor XOR2 (N4393, N4328, N1342);
nor NOR3 (N4394, N4391, N3885, N209);
nand NAND4 (N4395, N4387, N1083, N2327, N2515);
or OR2 (N4396, N4376, N2668);
nand NAND2 (N4397, N4389, N3101);
xor XOR2 (N4398, N4397, N2573);
xor XOR2 (N4399, N4366, N2082);
xor XOR2 (N4400, N4392, N2611);
buf BUF1 (N4401, N4396);
not NOT1 (N4402, N4398);
or OR2 (N4403, N4400, N2913);
not NOT1 (N4404, N4401);
nand NAND3 (N4405, N4388, N2856, N3169);
not NOT1 (N4406, N4402);
and AND4 (N4407, N4393, N2090, N2848, N3879);
xor XOR2 (N4408, N4382, N1263);
buf BUF1 (N4409, N4394);
and AND3 (N4410, N4407, N2362, N2334);
not NOT1 (N4411, N4390);
not NOT1 (N4412, N4404);
and AND2 (N4413, N4410, N2664);
nand NAND3 (N4414, N4413, N1652, N1543);
not NOT1 (N4415, N4395);
or OR2 (N4416, N4403, N222);
nor NOR3 (N4417, N4415, N1142, N2244);
and AND3 (N4418, N4406, N2278, N3571);
nand NAND3 (N4419, N4416, N3823, N1176);
not NOT1 (N4420, N4408);
xor XOR2 (N4421, N4412, N365);
not NOT1 (N4422, N4414);
nand NAND2 (N4423, N4418, N624);
xor XOR2 (N4424, N4405, N1480);
xor XOR2 (N4425, N4424, N3406);
buf BUF1 (N4426, N4425);
or OR2 (N4427, N4421, N2115);
nand NAND2 (N4428, N4409, N1565);
and AND3 (N4429, N4420, N1081, N3278);
or OR2 (N4430, N4419, N4060);
or OR3 (N4431, N4426, N2124, N3756);
buf BUF1 (N4432, N4427);
buf BUF1 (N4433, N4423);
buf BUF1 (N4434, N4431);
buf BUF1 (N4435, N4399);
and AND3 (N4436, N4434, N3874, N4286);
buf BUF1 (N4437, N4422);
xor XOR2 (N4438, N4428, N1957);
xor XOR2 (N4439, N4438, N3308);
or OR3 (N4440, N4429, N3216, N3771);
nand NAND3 (N4441, N4417, N1965, N650);
not NOT1 (N4442, N4432);
or OR2 (N4443, N4440, N61);
nand NAND3 (N4444, N4411, N534, N1124);
nor NOR3 (N4445, N4430, N1822, N2504);
nand NAND2 (N4446, N4444, N2227);
buf BUF1 (N4447, N4435);
and AND4 (N4448, N4441, N950, N2563, N3793);
and AND2 (N4449, N4448, N2074);
buf BUF1 (N4450, N4449);
or OR3 (N4451, N4447, N3721, N93);
nor NOR3 (N4452, N4445, N2394, N508);
or OR3 (N4453, N4446, N2354, N4258);
xor XOR2 (N4454, N4443, N1177);
or OR3 (N4455, N4452, N913, N265);
nand NAND4 (N4456, N4455, N148, N2356, N4309);
xor XOR2 (N4457, N4439, N2326);
nor NOR2 (N4458, N4442, N3297);
buf BUF1 (N4459, N4436);
or OR4 (N4460, N4457, N4420, N1913, N1680);
nor NOR4 (N4461, N4450, N703, N2968, N1657);
nor NOR4 (N4462, N4456, N2675, N3591, N2608);
nor NOR3 (N4463, N4460, N4198, N492);
and AND2 (N4464, N4433, N33);
not NOT1 (N4465, N4454);
nor NOR2 (N4466, N4465, N2936);
not NOT1 (N4467, N4466);
nand NAND2 (N4468, N4464, N4181);
nor NOR3 (N4469, N4467, N2510, N2201);
nor NOR2 (N4470, N4462, N3824);
nor NOR4 (N4471, N4470, N355, N3503, N53);
xor XOR2 (N4472, N4461, N1800);
not NOT1 (N4473, N4437);
and AND2 (N4474, N4468, N3984);
and AND4 (N4475, N4458, N2027, N4176, N2371);
buf BUF1 (N4476, N4463);
nand NAND2 (N4477, N4471, N1624);
nor NOR4 (N4478, N4473, N96, N2412, N1976);
buf BUF1 (N4479, N4453);
and AND3 (N4480, N4476, N2472, N868);
not NOT1 (N4481, N4459);
nor NOR2 (N4482, N4469, N3982);
and AND2 (N4483, N4479, N4319);
and AND2 (N4484, N4483, N1527);
buf BUF1 (N4485, N4472);
buf BUF1 (N4486, N4478);
nand NAND3 (N4487, N4485, N1242, N3916);
xor XOR2 (N4488, N4487, N2423);
or OR3 (N4489, N4482, N4393, N2075);
buf BUF1 (N4490, N4484);
nand NAND2 (N4491, N4489, N1876);
nand NAND4 (N4492, N4451, N4347, N4161, N4353);
buf BUF1 (N4493, N4477);
and AND4 (N4494, N4491, N9, N1249, N99);
not NOT1 (N4495, N4490);
or OR4 (N4496, N4475, N2414, N1503, N3452);
xor XOR2 (N4497, N4494, N973);
buf BUF1 (N4498, N4496);
and AND4 (N4499, N4498, N2988, N3894, N1510);
nand NAND2 (N4500, N4499, N1068);
nand NAND4 (N4501, N4492, N496, N2165, N1352);
nand NAND2 (N4502, N4501, N2884);
nand NAND2 (N4503, N4493, N3376);
and AND2 (N4504, N4481, N3172);
buf BUF1 (N4505, N4474);
and AND3 (N4506, N4505, N1915, N2823);
or OR4 (N4507, N4500, N2801, N1614, N4494);
or OR4 (N4508, N4506, N3620, N2997, N3280);
nand NAND4 (N4509, N4497, N872, N595, N3655);
or OR4 (N4510, N4503, N3508, N4005, N556);
xor XOR2 (N4511, N4488, N216);
nor NOR3 (N4512, N4504, N1571, N4081);
not NOT1 (N4513, N4502);
nor NOR3 (N4514, N4510, N4324, N1677);
nand NAND4 (N4515, N4511, N2592, N584, N501);
not NOT1 (N4516, N4509);
not NOT1 (N4517, N4486);
nand NAND4 (N4518, N4495, N66, N1459, N2599);
xor XOR2 (N4519, N4508, N537);
xor XOR2 (N4520, N4517, N1749);
and AND3 (N4521, N4520, N1743, N2225);
xor XOR2 (N4522, N4514, N1010);
nand NAND4 (N4523, N4515, N410, N3033, N1985);
nand NAND2 (N4524, N4519, N1751);
and AND3 (N4525, N4507, N3569, N4441);
nand NAND4 (N4526, N4512, N187, N284, N204);
nand NAND2 (N4527, N4521, N3443);
and AND4 (N4528, N4523, N2076, N4441, N2210);
buf BUF1 (N4529, N4528);
xor XOR2 (N4530, N4527, N2488);
xor XOR2 (N4531, N4480, N3324);
nor NOR2 (N4532, N4525, N369);
xor XOR2 (N4533, N4524, N56);
buf BUF1 (N4534, N4526);
not NOT1 (N4535, N4533);
xor XOR2 (N4536, N4531, N451);
buf BUF1 (N4537, N4532);
nor NOR3 (N4538, N4536, N768, N3112);
or OR3 (N4539, N4534, N1148, N2078);
or OR4 (N4540, N4513, N2725, N2145, N713);
or OR3 (N4541, N4540, N1807, N1676);
nand NAND3 (N4542, N4541, N1866, N4225);
nand NAND2 (N4543, N4538, N936);
nor NOR2 (N4544, N4537, N2304);
nor NOR4 (N4545, N4530, N2198, N1356, N2280);
not NOT1 (N4546, N4529);
and AND3 (N4547, N4539, N483, N651);
nand NAND3 (N4548, N4518, N3158, N2141);
not NOT1 (N4549, N4547);
buf BUF1 (N4550, N4548);
not NOT1 (N4551, N4522);
or OR2 (N4552, N4549, N3209);
and AND4 (N4553, N4535, N1210, N3125, N111);
or OR3 (N4554, N4552, N165, N4505);
or OR3 (N4555, N4544, N1141, N1352);
nand NAND4 (N4556, N4551, N4187, N117, N3841);
xor XOR2 (N4557, N4550, N281);
buf BUF1 (N4558, N4557);
or OR4 (N4559, N4553, N316, N3306, N800);
and AND2 (N4560, N4516, N1664);
and AND3 (N4561, N4554, N2680, N1680);
nand NAND3 (N4562, N4556, N4140, N3715);
nand NAND4 (N4563, N4543, N3830, N2918, N869);
nor NOR3 (N4564, N4558, N1371, N885);
xor XOR2 (N4565, N4542, N2220);
buf BUF1 (N4566, N4560);
buf BUF1 (N4567, N4564);
nand NAND2 (N4568, N4546, N3897);
nand NAND2 (N4569, N4563, N4092);
nand NAND4 (N4570, N4561, N1762, N3976, N2693);
not NOT1 (N4571, N4562);
nor NOR3 (N4572, N4568, N2232, N1488);
buf BUF1 (N4573, N4571);
and AND4 (N4574, N4545, N4449, N2876, N2185);
buf BUF1 (N4575, N4574);
and AND2 (N4576, N4555, N3880);
or OR2 (N4577, N4559, N1293);
nor NOR3 (N4578, N4577, N2844, N496);
and AND2 (N4579, N4576, N1626);
not NOT1 (N4580, N4569);
xor XOR2 (N4581, N4566, N1194);
or OR3 (N4582, N4575, N22, N3590);
or OR4 (N4583, N4565, N1506, N3077, N3341);
or OR4 (N4584, N4580, N789, N4149, N1790);
nand NAND4 (N4585, N4583, N3159, N3456, N564);
nor NOR3 (N4586, N4570, N2720, N2649);
or OR4 (N4587, N4586, N3210, N2846, N301);
and AND4 (N4588, N4578, N3934, N1862, N3864);
not NOT1 (N4589, N4588);
or OR4 (N4590, N4581, N4419, N2397, N1355);
and AND3 (N4591, N4582, N2267, N1419);
and AND3 (N4592, N4591, N1805, N2215);
buf BUF1 (N4593, N4590);
not NOT1 (N4594, N4589);
buf BUF1 (N4595, N4587);
and AND3 (N4596, N4593, N4159, N2070);
nand NAND4 (N4597, N4567, N238, N1963, N2294);
or OR3 (N4598, N4584, N2261, N4435);
or OR2 (N4599, N4596, N4067);
nand NAND4 (N4600, N4573, N4365, N4179, N1433);
buf BUF1 (N4601, N4597);
or OR2 (N4602, N4595, N488);
or OR2 (N4603, N4572, N1848);
and AND4 (N4604, N4603, N3223, N3423, N2511);
nand NAND2 (N4605, N4600, N482);
or OR2 (N4606, N4585, N1463);
not NOT1 (N4607, N4598);
nor NOR2 (N4608, N4594, N2030);
buf BUF1 (N4609, N4608);
nor NOR4 (N4610, N4599, N4609, N3346, N475);
nor NOR3 (N4611, N2225, N897, N1729);
or OR2 (N4612, N4610, N1838);
buf BUF1 (N4613, N4592);
not NOT1 (N4614, N4607);
nor NOR4 (N4615, N4579, N4598, N762, N1197);
nand NAND3 (N4616, N4606, N946, N1476);
not NOT1 (N4617, N4604);
nor NOR3 (N4618, N4602, N3592, N4402);
nor NOR2 (N4619, N4618, N1507);
nand NAND2 (N4620, N4611, N3328);
buf BUF1 (N4621, N4614);
xor XOR2 (N4622, N4613, N2357);
not NOT1 (N4623, N4601);
buf BUF1 (N4624, N4623);
nand NAND4 (N4625, N4621, N3739, N1340, N1051);
nor NOR2 (N4626, N4619, N3274);
buf BUF1 (N4627, N4620);
xor XOR2 (N4628, N4615, N2333);
nand NAND2 (N4629, N4622, N4358);
nand NAND3 (N4630, N4605, N4086, N945);
buf BUF1 (N4631, N4629);
and AND4 (N4632, N4624, N3263, N4202, N670);
and AND4 (N4633, N4632, N1257, N4180, N3655);
nand NAND3 (N4634, N4616, N1958, N190);
nand NAND2 (N4635, N4626, N3618);
nor NOR4 (N4636, N4634, N1749, N363, N993);
not NOT1 (N4637, N4627);
xor XOR2 (N4638, N4630, N1084);
not NOT1 (N4639, N4612);
buf BUF1 (N4640, N4631);
and AND2 (N4641, N4633, N4499);
nand NAND4 (N4642, N4636, N3613, N4202, N3464);
not NOT1 (N4643, N4638);
or OR3 (N4644, N4641, N1998, N2806);
nand NAND4 (N4645, N4642, N3670, N1937, N4405);
xor XOR2 (N4646, N4645, N671);
xor XOR2 (N4647, N4625, N2515);
and AND3 (N4648, N4643, N417, N1451);
xor XOR2 (N4649, N4640, N3944);
or OR4 (N4650, N4647, N982, N3346, N2075);
and AND3 (N4651, N4646, N4042, N389);
or OR3 (N4652, N4617, N2028, N2698);
not NOT1 (N4653, N4652);
nor NOR3 (N4654, N4644, N3742, N3966);
or OR4 (N4655, N4635, N1422, N2378, N495);
not NOT1 (N4656, N4653);
nand NAND2 (N4657, N4628, N2665);
xor XOR2 (N4658, N4639, N1857);
or OR4 (N4659, N4648, N2698, N4156, N4392);
xor XOR2 (N4660, N4651, N3037);
nand NAND3 (N4661, N4659, N1897, N212);
nand NAND2 (N4662, N4637, N3133);
buf BUF1 (N4663, N4654);
not NOT1 (N4664, N4657);
buf BUF1 (N4665, N4661);
and AND2 (N4666, N4660, N4021);
xor XOR2 (N4667, N4666, N2992);
xor XOR2 (N4668, N4650, N3376);
xor XOR2 (N4669, N4664, N437);
nand NAND4 (N4670, N4655, N2824, N3238, N71);
xor XOR2 (N4671, N4649, N1027);
or OR3 (N4672, N4671, N1469, N589);
or OR3 (N4673, N4672, N2806, N337);
and AND4 (N4674, N4667, N1538, N828, N1803);
xor XOR2 (N4675, N4668, N199);
or OR2 (N4676, N4662, N3024);
or OR2 (N4677, N4663, N3686);
or OR3 (N4678, N4665, N769, N2388);
xor XOR2 (N4679, N4677, N1136);
not NOT1 (N4680, N4675);
and AND4 (N4681, N4656, N2301, N4631, N2900);
buf BUF1 (N4682, N4680);
nand NAND4 (N4683, N4682, N2571, N460, N4526);
nor NOR4 (N4684, N4658, N2935, N2876, N4461);
nand NAND3 (N4685, N4673, N2581, N4188);
buf BUF1 (N4686, N4670);
not NOT1 (N4687, N4685);
and AND3 (N4688, N4674, N1223, N4545);
xor XOR2 (N4689, N4679, N967);
xor XOR2 (N4690, N4676, N2838);
xor XOR2 (N4691, N4690, N4623);
xor XOR2 (N4692, N4681, N3417);
or OR2 (N4693, N4691, N3014);
nand NAND4 (N4694, N4692, N4282, N501, N1421);
buf BUF1 (N4695, N4684);
nor NOR3 (N4696, N4683, N3258, N4592);
buf BUF1 (N4697, N4694);
xor XOR2 (N4698, N4693, N4532);
or OR2 (N4699, N4695, N2982);
or OR3 (N4700, N4698, N4694, N1971);
or OR3 (N4701, N4687, N3526, N2320);
buf BUF1 (N4702, N4697);
nand NAND2 (N4703, N4669, N3637);
buf BUF1 (N4704, N4700);
not NOT1 (N4705, N4688);
xor XOR2 (N4706, N4699, N3830);
buf BUF1 (N4707, N4704);
or OR4 (N4708, N4689, N949, N1152, N2954);
nand NAND2 (N4709, N4696, N3305);
xor XOR2 (N4710, N4705, N67);
or OR2 (N4711, N4706, N282);
not NOT1 (N4712, N4702);
nor NOR4 (N4713, N4708, N4619, N263, N5);
not NOT1 (N4714, N4711);
not NOT1 (N4715, N4709);
not NOT1 (N4716, N4712);
buf BUF1 (N4717, N4686);
not NOT1 (N4718, N4716);
xor XOR2 (N4719, N4710, N4654);
buf BUF1 (N4720, N4701);
and AND4 (N4721, N4720, N4635, N1902, N2504);
nand NAND2 (N4722, N4721, N1732);
nor NOR2 (N4723, N4718, N4171);
nor NOR2 (N4724, N4707, N3101);
not NOT1 (N4725, N4714);
or OR2 (N4726, N4703, N3208);
nand NAND3 (N4727, N4719, N4539, N827);
or OR4 (N4728, N4723, N1601, N3847, N203);
or OR2 (N4729, N4722, N1825);
buf BUF1 (N4730, N4713);
xor XOR2 (N4731, N4678, N1319);
nor NOR3 (N4732, N4726, N2421, N4477);
xor XOR2 (N4733, N4731, N1111);
buf BUF1 (N4734, N4732);
nand NAND3 (N4735, N4730, N4270, N918);
nand NAND2 (N4736, N4735, N558);
not NOT1 (N4737, N4733);
xor XOR2 (N4738, N4736, N4239);
or OR2 (N4739, N4737, N1451);
nand NAND4 (N4740, N4724, N2324, N4171, N270);
nor NOR4 (N4741, N4738, N103, N3320, N1048);
xor XOR2 (N4742, N4717, N3876);
nand NAND4 (N4743, N4728, N4181, N1552, N2497);
nor NOR3 (N4744, N4739, N2088, N3294);
buf BUF1 (N4745, N4715);
xor XOR2 (N4746, N4743, N1385);
nor NOR4 (N4747, N4740, N1587, N1740, N3966);
and AND3 (N4748, N4729, N2195, N2973);
xor XOR2 (N4749, N4742, N4012);
nand NAND4 (N4750, N4748, N2687, N3913, N2351);
or OR4 (N4751, N4749, N1747, N3536, N1416);
or OR3 (N4752, N4750, N2226, N4240);
or OR4 (N4753, N4725, N3566, N2457, N3398);
or OR4 (N4754, N4727, N1163, N1035, N594);
and AND4 (N4755, N4751, N1381, N1034, N2765);
not NOT1 (N4756, N4754);
or OR4 (N4757, N4744, N1549, N4338, N2503);
nor NOR4 (N4758, N4752, N4357, N3480, N484);
not NOT1 (N4759, N4758);
not NOT1 (N4760, N4757);
not NOT1 (N4761, N4746);
nand NAND2 (N4762, N4747, N3374);
or OR3 (N4763, N4756, N2853, N4134);
or OR4 (N4764, N4761, N341, N41, N1825);
not NOT1 (N4765, N4753);
xor XOR2 (N4766, N4763, N661);
xor XOR2 (N4767, N4760, N902);
or OR4 (N4768, N4741, N597, N3344, N4014);
not NOT1 (N4769, N4734);
buf BUF1 (N4770, N4765);
and AND2 (N4771, N4745, N3986);
nand NAND2 (N4772, N4771, N2805);
nand NAND2 (N4773, N4768, N2377);
xor XOR2 (N4774, N4755, N1306);
xor XOR2 (N4775, N4772, N1852);
xor XOR2 (N4776, N4774, N2122);
not NOT1 (N4777, N4762);
nor NOR2 (N4778, N4767, N2367);
nor NOR3 (N4779, N4778, N4449, N1420);
or OR4 (N4780, N4776, N2137, N244, N3908);
nand NAND2 (N4781, N4770, N2322);
and AND4 (N4782, N4779, N3266, N3453, N2189);
nor NOR3 (N4783, N4759, N1173, N4405);
not NOT1 (N4784, N4780);
not NOT1 (N4785, N4766);
not NOT1 (N4786, N4784);
xor XOR2 (N4787, N4782, N2340);
buf BUF1 (N4788, N4787);
or OR2 (N4789, N4775, N3985);
nand NAND3 (N4790, N4781, N1921, N2961);
and AND3 (N4791, N4786, N1029, N14);
xor XOR2 (N4792, N4791, N4381);
and AND3 (N4793, N4792, N1208, N3283);
nor NOR4 (N4794, N4773, N2728, N1613, N3070);
and AND4 (N4795, N4789, N3510, N1186, N2904);
nor NOR4 (N4796, N4794, N3328, N2945, N4288);
nand NAND4 (N4797, N4788, N1300, N2970, N1457);
xor XOR2 (N4798, N4793, N1808);
not NOT1 (N4799, N4769);
or OR2 (N4800, N4799, N53);
nand NAND3 (N4801, N4800, N2057, N173);
and AND4 (N4802, N4764, N4721, N2222, N1929);
not NOT1 (N4803, N4795);
xor XOR2 (N4804, N4798, N2799);
buf BUF1 (N4805, N4797);
xor XOR2 (N4806, N4804, N1509);
not NOT1 (N4807, N4790);
buf BUF1 (N4808, N4777);
nand NAND2 (N4809, N4807, N3044);
xor XOR2 (N4810, N4801, N1400);
xor XOR2 (N4811, N4802, N268);
buf BUF1 (N4812, N4785);
nor NOR2 (N4813, N4805, N4138);
nor NOR2 (N4814, N4812, N3635);
or OR4 (N4815, N4803, N2357, N2816, N923);
nand NAND4 (N4816, N4815, N1688, N2955, N1563);
not NOT1 (N4817, N4806);
not NOT1 (N4818, N4810);
not NOT1 (N4819, N4817);
not NOT1 (N4820, N4796);
nor NOR2 (N4821, N4816, N4680);
and AND2 (N4822, N4814, N3335);
buf BUF1 (N4823, N4821);
or OR4 (N4824, N4811, N3552, N599, N3586);
and AND3 (N4825, N4820, N3287, N2968);
or OR2 (N4826, N4808, N218);
nand NAND2 (N4827, N4819, N4637);
nor NOR4 (N4828, N4823, N2328, N2502, N3943);
or OR4 (N4829, N4827, N4591, N3142, N3294);
nor NOR2 (N4830, N4829, N4566);
nor NOR3 (N4831, N4822, N2502, N3007);
buf BUF1 (N4832, N4818);
not NOT1 (N4833, N4831);
and AND3 (N4834, N4833, N810, N909);
buf BUF1 (N4835, N4813);
not NOT1 (N4836, N4832);
xor XOR2 (N4837, N4826, N3284);
not NOT1 (N4838, N4836);
and AND3 (N4839, N4828, N3822, N1357);
not NOT1 (N4840, N4838);
not NOT1 (N4841, N4840);
buf BUF1 (N4842, N4825);
xor XOR2 (N4843, N4841, N2476);
xor XOR2 (N4844, N4839, N787);
xor XOR2 (N4845, N4844, N358);
nor NOR2 (N4846, N4783, N4589);
or OR3 (N4847, N4809, N1425, N766);
not NOT1 (N4848, N4843);
or OR4 (N4849, N4846, N1437, N2826, N3315);
buf BUF1 (N4850, N4837);
nand NAND4 (N4851, N4842, N784, N4277, N4078);
nor NOR4 (N4852, N4849, N1932, N3227, N2972);
or OR3 (N4853, N4834, N4148, N1629);
and AND2 (N4854, N4824, N15);
buf BUF1 (N4855, N4848);
and AND2 (N4856, N4851, N1715);
and AND4 (N4857, N4853, N153, N2680, N2007);
not NOT1 (N4858, N4855);
or OR4 (N4859, N4852, N213, N2630, N3465);
nand NAND3 (N4860, N4835, N2566, N152);
nand NAND2 (N4861, N4830, N3835);
nand NAND4 (N4862, N4847, N3182, N3966, N1026);
and AND2 (N4863, N4845, N1351);
and AND4 (N4864, N4859, N1267, N1246, N3901);
buf BUF1 (N4865, N4858);
and AND2 (N4866, N4862, N2498);
nand NAND4 (N4867, N4850, N2470, N2467, N4844);
not NOT1 (N4868, N4861);
not NOT1 (N4869, N4867);
or OR2 (N4870, N4860, N2011);
nand NAND4 (N4871, N4856, N4108, N2987, N3533);
not NOT1 (N4872, N4870);
xor XOR2 (N4873, N4864, N4110);
and AND2 (N4874, N4869, N1102);
and AND2 (N4875, N4872, N625);
xor XOR2 (N4876, N4874, N4356);
not NOT1 (N4877, N4854);
xor XOR2 (N4878, N4868, N4368);
nand NAND2 (N4879, N4866, N2210);
or OR3 (N4880, N4873, N3676, N1862);
and AND4 (N4881, N4863, N1461, N1262, N1827);
not NOT1 (N4882, N4879);
not NOT1 (N4883, N4871);
buf BUF1 (N4884, N4865);
nor NOR4 (N4885, N4881, N2549, N2755, N3419);
nand NAND2 (N4886, N4857, N3144);
and AND4 (N4887, N4886, N2178, N4576, N2567);
nand NAND3 (N4888, N4878, N3377, N4296);
and AND2 (N4889, N4887, N1219);
nor NOR4 (N4890, N4884, N3376, N3256, N469);
or OR3 (N4891, N4885, N3632, N432);
nor NOR2 (N4892, N4882, N1729);
nor NOR4 (N4893, N4889, N4646, N2092, N3910);
or OR4 (N4894, N4877, N181, N4615, N1374);
nand NAND3 (N4895, N4891, N4000, N2115);
not NOT1 (N4896, N4892);
nor NOR2 (N4897, N4893, N1579);
and AND2 (N4898, N4895, N4509);
buf BUF1 (N4899, N4890);
nand NAND4 (N4900, N4897, N2967, N633, N2156);
or OR4 (N4901, N4876, N3374, N1444, N1850);
nor NOR4 (N4902, N4880, N639, N3448, N3285);
nor NOR3 (N4903, N4901, N4879, N1545);
not NOT1 (N4904, N4894);
or OR3 (N4905, N4875, N2462, N3638);
and AND3 (N4906, N4899, N4609, N317);
or OR4 (N4907, N4906, N1805, N1163, N4204);
buf BUF1 (N4908, N4900);
not NOT1 (N4909, N4905);
xor XOR2 (N4910, N4902, N672);
not NOT1 (N4911, N4883);
buf BUF1 (N4912, N4909);
nor NOR2 (N4913, N4908, N2523);
nor NOR2 (N4914, N4898, N4840);
and AND4 (N4915, N4911, N2241, N2260, N4526);
buf BUF1 (N4916, N4914);
nand NAND4 (N4917, N4888, N334, N1552, N1898);
and AND4 (N4918, N4903, N3326, N3810, N1932);
xor XOR2 (N4919, N4910, N300);
xor XOR2 (N4920, N4919, N1358);
or OR3 (N4921, N4907, N1809, N785);
and AND2 (N4922, N4896, N1118);
or OR2 (N4923, N4915, N176);
not NOT1 (N4924, N4904);
or OR3 (N4925, N4923, N1207, N1689);
xor XOR2 (N4926, N4921, N4159);
or OR2 (N4927, N4924, N380);
not NOT1 (N4928, N4917);
xor XOR2 (N4929, N4918, N1011);
xor XOR2 (N4930, N4916, N4833);
buf BUF1 (N4931, N4926);
nor NOR4 (N4932, N4931, N1216, N1211, N1688);
xor XOR2 (N4933, N4932, N1241);
and AND3 (N4934, N4929, N3000, N1395);
or OR4 (N4935, N4927, N2777, N1912, N143);
nor NOR3 (N4936, N4913, N2351, N4074);
nand NAND2 (N4937, N4934, N921);
or OR3 (N4938, N4933, N672, N1077);
xor XOR2 (N4939, N4938, N920);
nand NAND4 (N4940, N4937, N2791, N3107, N1808);
nand NAND2 (N4941, N4940, N1467);
not NOT1 (N4942, N4925);
not NOT1 (N4943, N4941);
buf BUF1 (N4944, N4922);
buf BUF1 (N4945, N4943);
buf BUF1 (N4946, N4936);
nand NAND4 (N4947, N4939, N4911, N1831, N3194);
nand NAND4 (N4948, N4930, N4227, N4786, N1990);
not NOT1 (N4949, N4942);
or OR2 (N4950, N4944, N942);
nand NAND4 (N4951, N4946, N1475, N377, N4464);
not NOT1 (N4952, N4945);
not NOT1 (N4953, N4920);
and AND3 (N4954, N4949, N3712, N1163);
or OR3 (N4955, N4947, N4438, N2917);
xor XOR2 (N4956, N4950, N3686);
or OR2 (N4957, N4935, N3310);
buf BUF1 (N4958, N4928);
nand NAND2 (N4959, N4953, N2258);
or OR3 (N4960, N4959, N4136, N2912);
xor XOR2 (N4961, N4960, N1621);
not NOT1 (N4962, N4954);
and AND3 (N4963, N4948, N1266, N677);
nand NAND2 (N4964, N4951, N1428);
buf BUF1 (N4965, N4961);
buf BUF1 (N4966, N4956);
or OR2 (N4967, N4963, N3997);
nand NAND3 (N4968, N4966, N4664, N28);
xor XOR2 (N4969, N4912, N3490);
or OR3 (N4970, N4958, N2957, N1736);
xor XOR2 (N4971, N4955, N2295);
and AND3 (N4972, N4970, N231, N4000);
xor XOR2 (N4973, N4967, N4386);
nand NAND3 (N4974, N4965, N3716, N187);
xor XOR2 (N4975, N4964, N3388);
buf BUF1 (N4976, N4971);
or OR3 (N4977, N4973, N2456, N4596);
nand NAND2 (N4978, N4968, N2520);
xor XOR2 (N4979, N4969, N1072);
nor NOR3 (N4980, N4975, N1942, N1236);
or OR2 (N4981, N4957, N4891);
buf BUF1 (N4982, N4981);
nand NAND2 (N4983, N4952, N3342);
and AND3 (N4984, N4976, N683, N437);
nor NOR2 (N4985, N4983, N3038);
nor NOR4 (N4986, N4982, N341, N4867, N834);
and AND4 (N4987, N4979, N4829, N2973, N1696);
nor NOR3 (N4988, N4977, N3016, N3030);
or OR2 (N4989, N4962, N1271);
and AND4 (N4990, N4986, N1060, N4814, N685);
or OR2 (N4991, N4987, N4508);
xor XOR2 (N4992, N4974, N2681);
nand NAND3 (N4993, N4972, N760, N2050);
nand NAND3 (N4994, N4992, N2859, N4389);
nand NAND2 (N4995, N4985, N2893);
not NOT1 (N4996, N4991);
nand NAND2 (N4997, N4989, N1205);
not NOT1 (N4998, N4980);
nor NOR3 (N4999, N4993, N3217, N2298);
xor XOR2 (N5000, N4998, N3533);
or OR4 (N5001, N4984, N1292, N1968, N1034);
and AND3 (N5002, N4997, N3642, N992);
not NOT1 (N5003, N4978);
or OR3 (N5004, N5001, N2076, N358);
xor XOR2 (N5005, N5003, N3593);
buf BUF1 (N5006, N4996);
and AND2 (N5007, N4990, N369);
not NOT1 (N5008, N5007);
nand NAND2 (N5009, N5004, N995);
nor NOR2 (N5010, N5000, N3501);
and AND4 (N5011, N5002, N1247, N1149, N1549);
and AND2 (N5012, N5006, N3522);
xor XOR2 (N5013, N5005, N3913);
buf BUF1 (N5014, N5010);
buf BUF1 (N5015, N5014);
xor XOR2 (N5016, N5013, N2911);
not NOT1 (N5017, N4999);
nor NOR2 (N5018, N5009, N2239);
xor XOR2 (N5019, N5017, N2771);
not NOT1 (N5020, N5015);
xor XOR2 (N5021, N5018, N2538);
buf BUF1 (N5022, N5011);
buf BUF1 (N5023, N5008);
nor NOR2 (N5024, N5021, N1182);
not NOT1 (N5025, N5016);
not NOT1 (N5026, N5019);
xor XOR2 (N5027, N5026, N2772);
or OR3 (N5028, N4995, N69, N3940);
nand NAND3 (N5029, N5012, N2113, N1974);
or OR2 (N5030, N5029, N1068);
xor XOR2 (N5031, N5027, N4975);
and AND4 (N5032, N5024, N2209, N2286, N2335);
not NOT1 (N5033, N5025);
buf BUF1 (N5034, N5022);
not NOT1 (N5035, N5031);
not NOT1 (N5036, N5030);
and AND4 (N5037, N5034, N272, N582, N1023);
nor NOR3 (N5038, N5020, N1220, N2582);
and AND2 (N5039, N4988, N709);
not NOT1 (N5040, N5037);
or OR4 (N5041, N5023, N2579, N851, N3483);
not NOT1 (N5042, N5039);
or OR4 (N5043, N5036, N1738, N2615, N1732);
or OR4 (N5044, N5038, N4135, N4887, N4358);
xor XOR2 (N5045, N5028, N958);
xor XOR2 (N5046, N5042, N1401);
buf BUF1 (N5047, N5035);
not NOT1 (N5048, N5044);
nand NAND4 (N5049, N5032, N3237, N419, N463);
or OR2 (N5050, N5041, N1612);
or OR3 (N5051, N5040, N656, N2753);
or OR2 (N5052, N5045, N207);
and AND4 (N5053, N5043, N2243, N3035, N3847);
buf BUF1 (N5054, N5033);
not NOT1 (N5055, N5054);
xor XOR2 (N5056, N5055, N2059);
xor XOR2 (N5057, N5049, N879);
nand NAND2 (N5058, N5048, N946);
buf BUF1 (N5059, N5056);
and AND3 (N5060, N5050, N4779, N2875);
nand NAND4 (N5061, N5058, N747, N1090, N337);
nor NOR4 (N5062, N5060, N1733, N3541, N4257);
or OR4 (N5063, N5061, N3672, N4222, N221);
nand NAND4 (N5064, N5051, N501, N2940, N1912);
xor XOR2 (N5065, N5052, N1489);
or OR3 (N5066, N5063, N1155, N2189);
buf BUF1 (N5067, N5057);
buf BUF1 (N5068, N5059);
or OR4 (N5069, N5064, N2793, N1738, N350);
buf BUF1 (N5070, N5066);
xor XOR2 (N5071, N5069, N598);
buf BUF1 (N5072, N5067);
nand NAND4 (N5073, N5070, N2109, N4784, N4088);
not NOT1 (N5074, N5062);
xor XOR2 (N5075, N5073, N3877);
buf BUF1 (N5076, N5047);
xor XOR2 (N5077, N5075, N4773);
nand NAND2 (N5078, N4994, N1761);
nand NAND3 (N5079, N5053, N1284, N3695);
and AND4 (N5080, N5074, N533, N373, N565);
nor NOR3 (N5081, N5046, N1950, N712);
xor XOR2 (N5082, N5072, N4902);
nand NAND3 (N5083, N5082, N2387, N3472);
nor NOR3 (N5084, N5076, N4406, N3287);
or OR3 (N5085, N5071, N4503, N904);
or OR2 (N5086, N5078, N426);
buf BUF1 (N5087, N5086);
and AND3 (N5088, N5087, N3880, N2129);
buf BUF1 (N5089, N5068);
buf BUF1 (N5090, N5083);
or OR4 (N5091, N5085, N644, N3198, N2779);
or OR3 (N5092, N5065, N4473, N833);
not NOT1 (N5093, N5088);
nand NAND2 (N5094, N5084, N2961);
xor XOR2 (N5095, N5077, N4860);
or OR2 (N5096, N5093, N3116);
buf BUF1 (N5097, N5080);
or OR3 (N5098, N5079, N2968, N3695);
nor NOR4 (N5099, N5096, N2233, N5015, N4895);
and AND2 (N5100, N5097, N236);
not NOT1 (N5101, N5089);
xor XOR2 (N5102, N5092, N4102);
and AND3 (N5103, N5095, N3922, N1273);
nor NOR4 (N5104, N5094, N518, N2759, N3577);
nand NAND3 (N5105, N5090, N3542, N2);
nor NOR3 (N5106, N5102, N1386, N326);
nor NOR3 (N5107, N5100, N826, N3621);
and AND4 (N5108, N5098, N4044, N2447, N1610);
buf BUF1 (N5109, N5091);
nor NOR4 (N5110, N5081, N1030, N4557, N965);
not NOT1 (N5111, N5110);
nand NAND3 (N5112, N5104, N331, N3806);
xor XOR2 (N5113, N5101, N3884);
nor NOR4 (N5114, N5112, N4665, N2246, N1300);
or OR3 (N5115, N5108, N4608, N4372);
buf BUF1 (N5116, N5106);
not NOT1 (N5117, N5113);
and AND2 (N5118, N5116, N979);
not NOT1 (N5119, N5105);
and AND2 (N5120, N5118, N3861);
nand NAND4 (N5121, N5103, N4645, N1156, N503);
not NOT1 (N5122, N5120);
buf BUF1 (N5123, N5099);
not NOT1 (N5124, N5115);
nand NAND2 (N5125, N5117, N3442);
nand NAND3 (N5126, N5121, N3316, N1395);
buf BUF1 (N5127, N5119);
and AND2 (N5128, N5127, N271);
buf BUF1 (N5129, N5122);
nor NOR2 (N5130, N5125, N4736);
buf BUF1 (N5131, N5111);
and AND3 (N5132, N5114, N351, N2736);
nor NOR3 (N5133, N5128, N1369, N2674);
xor XOR2 (N5134, N5130, N1253);
xor XOR2 (N5135, N5126, N419);
buf BUF1 (N5136, N5133);
not NOT1 (N5137, N5123);
xor XOR2 (N5138, N5131, N3566);
or OR4 (N5139, N5124, N3293, N155, N2236);
nor NOR4 (N5140, N5136, N3732, N2137, N1539);
xor XOR2 (N5141, N5139, N4560);
buf BUF1 (N5142, N5141);
and AND4 (N5143, N5109, N2389, N2503, N4078);
not NOT1 (N5144, N5143);
nand NAND2 (N5145, N5134, N3447);
nand NAND2 (N5146, N5140, N2376);
not NOT1 (N5147, N5135);
buf BUF1 (N5148, N5144);
nand NAND3 (N5149, N5137, N5047, N1554);
nand NAND4 (N5150, N5148, N426, N3226, N4315);
xor XOR2 (N5151, N5138, N1213);
nor NOR3 (N5152, N5129, N4566, N2350);
xor XOR2 (N5153, N5145, N1366);
xor XOR2 (N5154, N5150, N2663);
nor NOR2 (N5155, N5107, N4435);
nor NOR3 (N5156, N5149, N469, N4753);
xor XOR2 (N5157, N5155, N684);
buf BUF1 (N5158, N5153);
buf BUF1 (N5159, N5142);
buf BUF1 (N5160, N5152);
or OR2 (N5161, N5160, N3151);
not NOT1 (N5162, N5158);
nor NOR3 (N5163, N5146, N3838, N663);
buf BUF1 (N5164, N5154);
nor NOR4 (N5165, N5151, N888, N1353, N1159);
xor XOR2 (N5166, N5132, N307);
nor NOR4 (N5167, N5166, N3771, N1254, N5066);
xor XOR2 (N5168, N5159, N3850);
and AND4 (N5169, N5163, N475, N4234, N3473);
or OR4 (N5170, N5147, N1241, N2603, N3563);
not NOT1 (N5171, N5168);
xor XOR2 (N5172, N5167, N3301);
not NOT1 (N5173, N5170);
and AND4 (N5174, N5165, N1875, N2192, N1049);
and AND4 (N5175, N5161, N2375, N3052, N707);
nor NOR2 (N5176, N5156, N3190);
buf BUF1 (N5177, N5175);
buf BUF1 (N5178, N5174);
not NOT1 (N5179, N5169);
buf BUF1 (N5180, N5171);
nand NAND2 (N5181, N5164, N236);
nand NAND3 (N5182, N5180, N2246, N632);
nand NAND3 (N5183, N5179, N407, N2141);
buf BUF1 (N5184, N5173);
nor NOR2 (N5185, N5157, N736);
and AND4 (N5186, N5177, N1442, N1164, N234);
and AND2 (N5187, N5183, N510);
buf BUF1 (N5188, N5187);
not NOT1 (N5189, N5184);
nor NOR4 (N5190, N5185, N153, N163, N5081);
buf BUF1 (N5191, N5188);
buf BUF1 (N5192, N5191);
xor XOR2 (N5193, N5176, N1544);
nor NOR3 (N5194, N5178, N2215, N3403);
buf BUF1 (N5195, N5193);
xor XOR2 (N5196, N5181, N994);
nand NAND3 (N5197, N5195, N5123, N216);
or OR4 (N5198, N5194, N18, N1896, N2297);
or OR4 (N5199, N5196, N507, N59, N535);
xor XOR2 (N5200, N5172, N107);
and AND3 (N5201, N5182, N682, N2848);
nand NAND3 (N5202, N5190, N963, N4550);
nand NAND3 (N5203, N5201, N4244, N4418);
xor XOR2 (N5204, N5203, N3847);
xor XOR2 (N5205, N5199, N247);
nor NOR2 (N5206, N5202, N592);
nand NAND2 (N5207, N5204, N5047);
or OR3 (N5208, N5192, N3321, N3449);
nand NAND2 (N5209, N5197, N4744);
not NOT1 (N5210, N5209);
buf BUF1 (N5211, N5206);
and AND4 (N5212, N5189, N2009, N5044, N4789);
nand NAND3 (N5213, N5207, N2649, N3105);
or OR3 (N5214, N5210, N2708, N162);
and AND2 (N5215, N5162, N2301);
or OR2 (N5216, N5208, N3003);
nand NAND4 (N5217, N5215, N793, N328, N5047);
buf BUF1 (N5218, N5205);
nand NAND3 (N5219, N5217, N3, N2655);
not NOT1 (N5220, N5216);
nor NOR4 (N5221, N5220, N2857, N1157, N4319);
nand NAND3 (N5222, N5212, N5104, N3186);
buf BUF1 (N5223, N5200);
or OR3 (N5224, N5223, N3801, N1094);
or OR4 (N5225, N5213, N961, N4612, N2975);
or OR3 (N5226, N5218, N4578, N2571);
buf BUF1 (N5227, N5186);
or OR2 (N5228, N5214, N582);
buf BUF1 (N5229, N5221);
nor NOR3 (N5230, N5227, N2201, N2528);
and AND3 (N5231, N5211, N3330, N5132);
buf BUF1 (N5232, N5224);
xor XOR2 (N5233, N5219, N1925);
buf BUF1 (N5234, N5231);
and AND4 (N5235, N5232, N4764, N3082, N47);
xor XOR2 (N5236, N5228, N4160);
buf BUF1 (N5237, N5225);
nand NAND4 (N5238, N5237, N3526, N543, N1011);
nand NAND2 (N5239, N5222, N3120);
buf BUF1 (N5240, N5238);
nor NOR4 (N5241, N5226, N1832, N3120, N1015);
nand NAND3 (N5242, N5239, N4155, N2102);
and AND2 (N5243, N5233, N1317);
nand NAND2 (N5244, N5234, N2895);
or OR2 (N5245, N5230, N1241);
nand NAND3 (N5246, N5244, N4386, N3036);
not NOT1 (N5247, N5235);
nor NOR3 (N5248, N5246, N905, N1575);
buf BUF1 (N5249, N5245);
and AND4 (N5250, N5240, N3839, N3584, N1588);
nand NAND4 (N5251, N5242, N4388, N5052, N4127);
and AND3 (N5252, N5247, N2864, N4283);
nand NAND4 (N5253, N5249, N816, N4706, N1651);
and AND2 (N5254, N5251, N1841);
or OR2 (N5255, N5248, N4087);
or OR2 (N5256, N5255, N1731);
buf BUF1 (N5257, N5229);
buf BUF1 (N5258, N5253);
buf BUF1 (N5259, N5256);
nor NOR2 (N5260, N5236, N1525);
not NOT1 (N5261, N5250);
or OR3 (N5262, N5198, N5047, N2400);
not NOT1 (N5263, N5258);
nand NAND4 (N5264, N5243, N2398, N4102, N40);
or OR2 (N5265, N5264, N594);
not NOT1 (N5266, N5257);
and AND3 (N5267, N5266, N4019, N1564);
nor NOR4 (N5268, N5252, N4821, N4161, N3009);
and AND4 (N5269, N5263, N3793, N3319, N4172);
and AND4 (N5270, N5260, N4263, N4265, N4357);
not NOT1 (N5271, N5254);
nor NOR3 (N5272, N5270, N2370, N3573);
not NOT1 (N5273, N5259);
xor XOR2 (N5274, N5272, N2571);
buf BUF1 (N5275, N5265);
nor NOR4 (N5276, N5241, N1218, N4912, N5187);
xor XOR2 (N5277, N5261, N2756);
and AND3 (N5278, N5268, N3216, N3894);
and AND3 (N5279, N5278, N2203, N3479);
not NOT1 (N5280, N5267);
buf BUF1 (N5281, N5277);
and AND3 (N5282, N5275, N4960, N2494);
or OR3 (N5283, N5262, N2498, N2842);
not NOT1 (N5284, N5271);
or OR3 (N5285, N5281, N3181, N575);
or OR4 (N5286, N5285, N1153, N639, N913);
nor NOR4 (N5287, N5286, N3858, N3299, N950);
and AND3 (N5288, N5282, N4178, N4796);
nor NOR3 (N5289, N5276, N4910, N1232);
not NOT1 (N5290, N5289);
and AND4 (N5291, N5280, N333, N4646, N687);
nor NOR2 (N5292, N5283, N4440);
not NOT1 (N5293, N5290);
buf BUF1 (N5294, N5291);
and AND4 (N5295, N5273, N2031, N1164, N1536);
xor XOR2 (N5296, N5287, N2857);
buf BUF1 (N5297, N5296);
buf BUF1 (N5298, N5279);
and AND3 (N5299, N5274, N1780, N2158);
buf BUF1 (N5300, N5293);
nor NOR2 (N5301, N5297, N4707);
and AND4 (N5302, N5301, N2966, N702, N4884);
nor NOR4 (N5303, N5294, N3477, N808, N2052);
xor XOR2 (N5304, N5302, N3315);
nor NOR4 (N5305, N5303, N3413, N2858, N1135);
buf BUF1 (N5306, N5300);
buf BUF1 (N5307, N5284);
not NOT1 (N5308, N5299);
not NOT1 (N5309, N5305);
not NOT1 (N5310, N5292);
nor NOR3 (N5311, N5288, N3802, N1370);
nand NAND2 (N5312, N5295, N4467);
and AND4 (N5313, N5298, N5116, N497, N1971);
buf BUF1 (N5314, N5310);
nand NAND4 (N5315, N5312, N920, N2122, N5044);
or OR4 (N5316, N5304, N4461, N4625, N4494);
not NOT1 (N5317, N5311);
nand NAND3 (N5318, N5317, N742, N3722);
buf BUF1 (N5319, N5314);
nor NOR3 (N5320, N5315, N1499, N395);
or OR4 (N5321, N5318, N4886, N5140, N886);
xor XOR2 (N5322, N5320, N1190);
or OR2 (N5323, N5322, N495);
xor XOR2 (N5324, N5307, N193);
nor NOR3 (N5325, N5313, N129, N166);
xor XOR2 (N5326, N5323, N2201);
xor XOR2 (N5327, N5269, N454);
not NOT1 (N5328, N5321);
nor NOR4 (N5329, N5306, N3040, N371, N2337);
not NOT1 (N5330, N5309);
and AND3 (N5331, N5330, N2414, N2114);
buf BUF1 (N5332, N5324);
nand NAND2 (N5333, N5319, N4410);
buf BUF1 (N5334, N5329);
xor XOR2 (N5335, N5328, N4674);
not NOT1 (N5336, N5308);
xor XOR2 (N5337, N5331, N4733);
and AND2 (N5338, N5333, N5278);
xor XOR2 (N5339, N5316, N4407);
or OR4 (N5340, N5335, N807, N3562, N949);
nand NAND4 (N5341, N5336, N2234, N3475, N4055);
xor XOR2 (N5342, N5338, N4037);
nand NAND3 (N5343, N5341, N3762, N352);
or OR2 (N5344, N5342, N1831);
buf BUF1 (N5345, N5337);
not NOT1 (N5346, N5326);
or OR3 (N5347, N5345, N1150, N1216);
xor XOR2 (N5348, N5334, N160);
or OR2 (N5349, N5346, N5012);
or OR3 (N5350, N5349, N1503, N872);
or OR4 (N5351, N5344, N1982, N3939, N996);
buf BUF1 (N5352, N5351);
nor NOR2 (N5353, N5340, N5031);
nand NAND2 (N5354, N5347, N2680);
nand NAND4 (N5355, N5325, N4972, N664, N1405);
buf BUF1 (N5356, N5354);
or OR4 (N5357, N5350, N2971, N732, N1302);
nor NOR3 (N5358, N5339, N2148, N3463);
not NOT1 (N5359, N5353);
nor NOR4 (N5360, N5355, N4724, N4380, N2813);
xor XOR2 (N5361, N5360, N4571);
nor NOR3 (N5362, N5358, N2492, N2090);
and AND3 (N5363, N5332, N5141, N1452);
or OR2 (N5364, N5361, N5015);
xor XOR2 (N5365, N5359, N81);
or OR3 (N5366, N5363, N4382, N1981);
nand NAND3 (N5367, N5352, N4999, N5219);
nor NOR2 (N5368, N5327, N346);
buf BUF1 (N5369, N5362);
or OR2 (N5370, N5369, N2291);
xor XOR2 (N5371, N5348, N2845);
not NOT1 (N5372, N5367);
xor XOR2 (N5373, N5371, N3050);
and AND4 (N5374, N5356, N1906, N4330, N4885);
nand NAND4 (N5375, N5368, N1769, N574, N498);
not NOT1 (N5376, N5364);
nor NOR3 (N5377, N5375, N3474, N4156);
and AND4 (N5378, N5343, N111, N1422, N3770);
xor XOR2 (N5379, N5366, N1383);
or OR4 (N5380, N5370, N5030, N4733, N2874);
xor XOR2 (N5381, N5380, N4239);
nor NOR4 (N5382, N5377, N4654, N3819, N1219);
nand NAND3 (N5383, N5376, N228, N2104);
and AND2 (N5384, N5379, N2608);
xor XOR2 (N5385, N5374, N3411);
buf BUF1 (N5386, N5372);
buf BUF1 (N5387, N5381);
nand NAND3 (N5388, N5385, N5118, N4259);
nand NAND2 (N5389, N5384, N3374);
buf BUF1 (N5390, N5388);
nand NAND2 (N5391, N5387, N1412);
xor XOR2 (N5392, N5386, N4517);
or OR4 (N5393, N5392, N4693, N1677, N4715);
buf BUF1 (N5394, N5389);
or OR2 (N5395, N5391, N2608);
nand NAND2 (N5396, N5395, N2617);
or OR3 (N5397, N5357, N3371, N4499);
xor XOR2 (N5398, N5383, N3311);
nor NOR3 (N5399, N5373, N3599, N2276);
buf BUF1 (N5400, N5399);
nor NOR4 (N5401, N5400, N4706, N5290, N1945);
or OR4 (N5402, N5394, N4706, N742, N310);
and AND4 (N5403, N5393, N4152, N83, N2759);
nand NAND4 (N5404, N5398, N4203, N3828, N1706);
and AND3 (N5405, N5390, N696, N3321);
nand NAND2 (N5406, N5382, N4886);
or OR4 (N5407, N5405, N2080, N2710, N64);
and AND4 (N5408, N5397, N4698, N1754, N2908);
xor XOR2 (N5409, N5402, N3183);
or OR2 (N5410, N5408, N2823);
and AND2 (N5411, N5407, N989);
and AND3 (N5412, N5396, N2020, N4573);
nand NAND2 (N5413, N5365, N1678);
not NOT1 (N5414, N5401);
nand NAND3 (N5415, N5403, N2640, N5393);
nor NOR3 (N5416, N5378, N4140, N2576);
and AND4 (N5417, N5413, N4101, N995, N3712);
and AND2 (N5418, N5404, N5238);
nor NOR2 (N5419, N5411, N1321);
xor XOR2 (N5420, N5406, N4471);
nand NAND2 (N5421, N5420, N5316);
xor XOR2 (N5422, N5419, N210);
not NOT1 (N5423, N5421);
nand NAND2 (N5424, N5422, N4190);
nor NOR4 (N5425, N5418, N514, N3198, N2915);
and AND4 (N5426, N5415, N1152, N1064, N1441);
or OR4 (N5427, N5424, N717, N2623, N2422);
and AND3 (N5428, N5416, N1335, N1048);
nor NOR2 (N5429, N5409, N4834);
xor XOR2 (N5430, N5414, N589);
not NOT1 (N5431, N5425);
nand NAND2 (N5432, N5417, N3925);
xor XOR2 (N5433, N5429, N5421);
nand NAND4 (N5434, N5432, N3952, N3267, N4458);
or OR2 (N5435, N5410, N344);
nand NAND4 (N5436, N5423, N2820, N1784, N3295);
not NOT1 (N5437, N5427);
and AND3 (N5438, N5431, N1055, N517);
nor NOR2 (N5439, N5426, N4684);
nand NAND3 (N5440, N5436, N353, N4134);
xor XOR2 (N5441, N5437, N5243);
xor XOR2 (N5442, N5440, N4814);
or OR2 (N5443, N5433, N1046);
xor XOR2 (N5444, N5441, N1817);
and AND3 (N5445, N5430, N2257, N2068);
nand NAND4 (N5446, N5445, N3770, N2347, N4756);
or OR3 (N5447, N5439, N2727, N4409);
nor NOR3 (N5448, N5435, N634, N4142);
not NOT1 (N5449, N5434);
nor NOR3 (N5450, N5438, N2911, N3586);
xor XOR2 (N5451, N5444, N4926);
nand NAND4 (N5452, N5448, N3425, N2913, N374);
and AND2 (N5453, N5443, N3857);
and AND4 (N5454, N5412, N448, N4600, N1378);
or OR4 (N5455, N5452, N1969, N3908, N2842);
xor XOR2 (N5456, N5442, N2664);
not NOT1 (N5457, N5456);
or OR3 (N5458, N5446, N2485, N4435);
nand NAND4 (N5459, N5454, N2110, N1385, N1642);
or OR4 (N5460, N5447, N1323, N3096, N3435);
nor NOR4 (N5461, N5428, N2838, N4620, N776);
xor XOR2 (N5462, N5460, N2953);
nor NOR3 (N5463, N5455, N3354, N879);
not NOT1 (N5464, N5457);
and AND4 (N5465, N5462, N3054, N3775, N1827);
nor NOR4 (N5466, N5449, N3818, N4490, N2609);
nor NOR4 (N5467, N5453, N5163, N5462, N251);
or OR3 (N5468, N5450, N1333, N1755);
nor NOR4 (N5469, N5461, N2239, N1382, N750);
nor NOR2 (N5470, N5469, N7);
nand NAND4 (N5471, N5463, N3702, N3828, N1069);
xor XOR2 (N5472, N5471, N3241);
buf BUF1 (N5473, N5459);
not NOT1 (N5474, N5466);
buf BUF1 (N5475, N5467);
not NOT1 (N5476, N5470);
and AND4 (N5477, N5468, N4596, N356, N1979);
nor NOR2 (N5478, N5476, N1295);
buf BUF1 (N5479, N5464);
buf BUF1 (N5480, N5479);
and AND3 (N5481, N5478, N2596, N1226);
xor XOR2 (N5482, N5458, N710);
not NOT1 (N5483, N5474);
nor NOR4 (N5484, N5483, N4763, N2557, N557);
not NOT1 (N5485, N5473);
nand NAND3 (N5486, N5482, N393, N1006);
xor XOR2 (N5487, N5486, N482);
xor XOR2 (N5488, N5485, N19);
or OR2 (N5489, N5475, N1725);
nand NAND4 (N5490, N5489, N774, N3295, N2495);
or OR2 (N5491, N5480, N5128);
nand NAND3 (N5492, N5490, N4352, N2890);
or OR2 (N5493, N5465, N1199);
and AND3 (N5494, N5487, N1171, N2927);
or OR2 (N5495, N5484, N2994);
and AND3 (N5496, N5451, N698, N962);
and AND2 (N5497, N5496, N3384);
and AND3 (N5498, N5481, N26, N1804);
and AND3 (N5499, N5493, N3590, N3934);
and AND2 (N5500, N5492, N5100);
or OR2 (N5501, N5472, N4040);
buf BUF1 (N5502, N5494);
nor NOR3 (N5503, N5498, N3053, N4027);
nor NOR4 (N5504, N5500, N4554, N3058, N507);
nor NOR4 (N5505, N5501, N3061, N1277, N430);
and AND2 (N5506, N5495, N3302);
xor XOR2 (N5507, N5504, N1488);
xor XOR2 (N5508, N5503, N4014);
and AND3 (N5509, N5502, N4819, N2645);
nor NOR2 (N5510, N5508, N4743);
xor XOR2 (N5511, N5507, N5088);
and AND3 (N5512, N5491, N4864, N3923);
nor NOR4 (N5513, N5510, N442, N2744, N3700);
nor NOR2 (N5514, N5505, N3925);
and AND4 (N5515, N5511, N730, N2671, N4690);
nor NOR4 (N5516, N5488, N3871, N1576, N1329);
buf BUF1 (N5517, N5509);
and AND2 (N5518, N5517, N1995);
and AND2 (N5519, N5516, N5209);
xor XOR2 (N5520, N5477, N2749);
xor XOR2 (N5521, N5512, N2024);
or OR4 (N5522, N5499, N3434, N884, N5497);
and AND2 (N5523, N1340, N3922);
nor NOR4 (N5524, N5515, N2980, N5220, N4469);
nand NAND3 (N5525, N5514, N2220, N2667);
or OR3 (N5526, N5521, N1924, N1773);
xor XOR2 (N5527, N5520, N15);
buf BUF1 (N5528, N5518);
nand NAND3 (N5529, N5525, N3667, N4715);
and AND3 (N5530, N5528, N1080, N4524);
or OR4 (N5531, N5519, N71, N2198, N1432);
buf BUF1 (N5532, N5524);
or OR4 (N5533, N5531, N5230, N3715, N4100);
nor NOR3 (N5534, N5533, N4193, N2112);
and AND2 (N5535, N5522, N4365);
not NOT1 (N5536, N5535);
or OR2 (N5537, N5506, N4960);
not NOT1 (N5538, N5527);
nor NOR4 (N5539, N5537, N1279, N2157, N3043);
and AND2 (N5540, N5526, N3723);
not NOT1 (N5541, N5540);
or OR3 (N5542, N5529, N4650, N2181);
nand NAND2 (N5543, N5541, N497);
nor NOR3 (N5544, N5536, N1692, N1329);
nand NAND4 (N5545, N5544, N2159, N1433, N2254);
nor NOR3 (N5546, N5542, N4451, N1129);
or OR4 (N5547, N5546, N849, N4015, N5286);
nor NOR4 (N5548, N5532, N1816, N4855, N1732);
xor XOR2 (N5549, N5539, N638);
nand NAND4 (N5550, N5545, N4571, N4356, N3410);
buf BUF1 (N5551, N5550);
or OR2 (N5552, N5547, N2910);
buf BUF1 (N5553, N5513);
buf BUF1 (N5554, N5552);
not NOT1 (N5555, N5554);
nor NOR3 (N5556, N5534, N3329, N629);
or OR2 (N5557, N5538, N4324);
nor NOR4 (N5558, N5549, N2100, N438, N1514);
and AND3 (N5559, N5548, N4037, N962);
buf BUF1 (N5560, N5558);
not NOT1 (N5561, N5555);
buf BUF1 (N5562, N5557);
and AND2 (N5563, N5553, N2791);
and AND3 (N5564, N5551, N3776, N1376);
xor XOR2 (N5565, N5530, N2748);
nand NAND3 (N5566, N5523, N2070, N1922);
or OR3 (N5567, N5564, N3526, N1860);
nor NOR3 (N5568, N5560, N4181, N684);
and AND4 (N5569, N5568, N3873, N3617, N3031);
and AND4 (N5570, N5565, N5113, N1456, N1001);
not NOT1 (N5571, N5562);
or OR3 (N5572, N5569, N2822, N12);
xor XOR2 (N5573, N5559, N530);
xor XOR2 (N5574, N5571, N474);
xor XOR2 (N5575, N5567, N4830);
xor XOR2 (N5576, N5561, N1396);
nor NOR2 (N5577, N5543, N2543);
and AND4 (N5578, N5563, N677, N5231, N968);
nor NOR4 (N5579, N5578, N2737, N3674, N5191);
xor XOR2 (N5580, N5575, N1815);
nand NAND2 (N5581, N5573, N3860);
or OR3 (N5582, N5566, N960, N497);
xor XOR2 (N5583, N5570, N1873);
nor NOR2 (N5584, N5576, N4481);
not NOT1 (N5585, N5574);
not NOT1 (N5586, N5585);
or OR3 (N5587, N5581, N5331, N4243);
nand NAND4 (N5588, N5587, N1837, N2418, N4171);
nand NAND3 (N5589, N5584, N5002, N5054);
buf BUF1 (N5590, N5589);
nand NAND2 (N5591, N5590, N5122);
buf BUF1 (N5592, N5580);
or OR2 (N5593, N5591, N5194);
xor XOR2 (N5594, N5586, N1943);
nor NOR3 (N5595, N5572, N4855, N4133);
xor XOR2 (N5596, N5592, N5542);
and AND4 (N5597, N5588, N4941, N3489, N4965);
buf BUF1 (N5598, N5556);
xor XOR2 (N5599, N5583, N1914);
or OR3 (N5600, N5577, N742, N138);
buf BUF1 (N5601, N5600);
nor NOR4 (N5602, N5579, N3225, N5014, N416);
buf BUF1 (N5603, N5582);
nor NOR4 (N5604, N5595, N1278, N3750, N2495);
or OR4 (N5605, N5598, N1455, N2313, N1691);
buf BUF1 (N5606, N5597);
nand NAND4 (N5607, N5603, N889, N2853, N5575);
nor NOR3 (N5608, N5599, N216, N2696);
xor XOR2 (N5609, N5606, N3152);
not NOT1 (N5610, N5593);
not NOT1 (N5611, N5601);
buf BUF1 (N5612, N5611);
not NOT1 (N5613, N5607);
buf BUF1 (N5614, N5610);
nor NOR2 (N5615, N5602, N4832);
xor XOR2 (N5616, N5596, N1787);
nand NAND2 (N5617, N5616, N3239);
buf BUF1 (N5618, N5612);
nand NAND4 (N5619, N5604, N2850, N2302, N2179);
xor XOR2 (N5620, N5609, N3901);
or OR3 (N5621, N5594, N3154, N2146);
nor NOR4 (N5622, N5618, N5156, N4495, N4565);
nor NOR2 (N5623, N5622, N1144);
not NOT1 (N5624, N5620);
buf BUF1 (N5625, N5614);
nor NOR4 (N5626, N5619, N2837, N3613, N2109);
not NOT1 (N5627, N5617);
nand NAND4 (N5628, N5608, N5619, N1873, N2582);
nor NOR3 (N5629, N5626, N5253, N449);
not NOT1 (N5630, N5605);
nor NOR3 (N5631, N5629, N2402, N784);
nand NAND2 (N5632, N5615, N3054);
and AND4 (N5633, N5627, N1152, N2080, N972);
not NOT1 (N5634, N5632);
xor XOR2 (N5635, N5634, N784);
and AND2 (N5636, N5628, N3690);
or OR2 (N5637, N5633, N2885);
not NOT1 (N5638, N5624);
nand NAND3 (N5639, N5623, N1294, N2850);
or OR4 (N5640, N5631, N304, N5031, N5458);
nor NOR2 (N5641, N5640, N2704);
buf BUF1 (N5642, N5621);
or OR3 (N5643, N5639, N2135, N4776);
not NOT1 (N5644, N5637);
buf BUF1 (N5645, N5638);
and AND4 (N5646, N5613, N5342, N2761, N4734);
xor XOR2 (N5647, N5635, N288);
nand NAND4 (N5648, N5644, N3808, N4502, N447);
or OR2 (N5649, N5645, N5486);
and AND4 (N5650, N5649, N1376, N1033, N2935);
or OR4 (N5651, N5646, N4568, N4716, N983);
buf BUF1 (N5652, N5625);
xor XOR2 (N5653, N5643, N4618);
not NOT1 (N5654, N5648);
nor NOR3 (N5655, N5651, N4615, N1234);
or OR2 (N5656, N5655, N5560);
or OR4 (N5657, N5636, N1072, N1422, N2894);
and AND3 (N5658, N5630, N327, N1745);
not NOT1 (N5659, N5641);
nand NAND4 (N5660, N5652, N4404, N2118, N3551);
or OR2 (N5661, N5660, N1950);
xor XOR2 (N5662, N5642, N793);
and AND4 (N5663, N5658, N4408, N4938, N3462);
xor XOR2 (N5664, N5656, N1853);
and AND3 (N5665, N5653, N3233, N849);
or OR4 (N5666, N5663, N553, N1030, N1603);
nor NOR2 (N5667, N5657, N1257);
nor NOR2 (N5668, N5667, N2612);
nor NOR3 (N5669, N5668, N230, N4302);
buf BUF1 (N5670, N5664);
not NOT1 (N5671, N5650);
or OR4 (N5672, N5662, N222, N567, N2309);
buf BUF1 (N5673, N5647);
nor NOR4 (N5674, N5654, N4475, N5290, N2235);
nand NAND3 (N5675, N5673, N4207, N5531);
and AND3 (N5676, N5675, N219, N340);
nor NOR4 (N5677, N5665, N2731, N90, N4023);
xor XOR2 (N5678, N5666, N555);
buf BUF1 (N5679, N5659);
nand NAND3 (N5680, N5669, N9, N2869);
buf BUF1 (N5681, N5679);
not NOT1 (N5682, N5674);
not NOT1 (N5683, N5680);
nor NOR2 (N5684, N5676, N3789);
xor XOR2 (N5685, N5671, N1661);
or OR3 (N5686, N5670, N4977, N726);
xor XOR2 (N5687, N5683, N3024);
or OR2 (N5688, N5661, N1328);
nand NAND2 (N5689, N5687, N1203);
and AND4 (N5690, N5682, N3998, N5057, N2753);
or OR2 (N5691, N5672, N320);
or OR4 (N5692, N5688, N4561, N525, N1912);
xor XOR2 (N5693, N5692, N1793);
not NOT1 (N5694, N5684);
nand NAND2 (N5695, N5686, N559);
nand NAND3 (N5696, N5677, N1765, N2071);
nand NAND4 (N5697, N5691, N2459, N2817, N1684);
and AND3 (N5698, N5697, N4698, N5628);
buf BUF1 (N5699, N5690);
or OR2 (N5700, N5689, N3467);
not NOT1 (N5701, N5681);
buf BUF1 (N5702, N5701);
nand NAND3 (N5703, N5678, N4275, N5464);
not NOT1 (N5704, N5696);
nor NOR2 (N5705, N5694, N4911);
not NOT1 (N5706, N5700);
nand NAND3 (N5707, N5703, N4443, N666);
nand NAND3 (N5708, N5707, N2986, N5354);
or OR2 (N5709, N5695, N2317);
nor NOR3 (N5710, N5685, N3080, N582);
xor XOR2 (N5711, N5705, N3100);
nor NOR2 (N5712, N5698, N4939);
or OR3 (N5713, N5711, N3862, N173);
buf BUF1 (N5714, N5704);
and AND2 (N5715, N5712, N680);
buf BUF1 (N5716, N5715);
buf BUF1 (N5717, N5693);
nor NOR3 (N5718, N5699, N2134, N2776);
nor NOR2 (N5719, N5713, N2503);
or OR3 (N5720, N5717, N1432, N5494);
not NOT1 (N5721, N5716);
not NOT1 (N5722, N5719);
nor NOR2 (N5723, N5721, N4034);
xor XOR2 (N5724, N5710, N188);
buf BUF1 (N5725, N5722);
nand NAND3 (N5726, N5725, N5185, N1476);
or OR3 (N5727, N5708, N437, N488);
buf BUF1 (N5728, N5720);
xor XOR2 (N5729, N5726, N3520);
xor XOR2 (N5730, N5727, N1637);
nand NAND4 (N5731, N5706, N3096, N994, N2754);
and AND3 (N5732, N5714, N3160, N5637);
and AND4 (N5733, N5709, N2973, N1854, N1694);
nand NAND4 (N5734, N5731, N477, N4727, N5667);
nor NOR3 (N5735, N5718, N794, N4622);
xor XOR2 (N5736, N5730, N4477);
and AND4 (N5737, N5733, N4668, N225, N4255);
nor NOR3 (N5738, N5724, N1209, N3185);
and AND3 (N5739, N5732, N5369, N3068);
nor NOR3 (N5740, N5736, N1314, N113);
nor NOR3 (N5741, N5723, N5264, N2407);
buf BUF1 (N5742, N5739);
or OR4 (N5743, N5728, N3477, N3930, N140);
nand NAND2 (N5744, N5735, N4566);
and AND3 (N5745, N5740, N1603, N2438);
nor NOR3 (N5746, N5745, N5547, N2103);
nand NAND2 (N5747, N5729, N5052);
xor XOR2 (N5748, N5734, N5540);
nand NAND2 (N5749, N5737, N3311);
xor XOR2 (N5750, N5747, N1886);
buf BUF1 (N5751, N5749);
nand NAND4 (N5752, N5744, N4493, N1218, N3861);
or OR2 (N5753, N5750, N4874);
xor XOR2 (N5754, N5753, N2215);
and AND4 (N5755, N5743, N175, N2025, N505);
not NOT1 (N5756, N5746);
buf BUF1 (N5757, N5752);
nor NOR4 (N5758, N5748, N4223, N179, N1831);
nor NOR4 (N5759, N5755, N2716, N2833, N5740);
buf BUF1 (N5760, N5758);
buf BUF1 (N5761, N5757);
nor NOR4 (N5762, N5759, N1421, N5034, N1404);
or OR3 (N5763, N5762, N5249, N5171);
nor NOR4 (N5764, N5751, N4328, N2676, N1791);
buf BUF1 (N5765, N5756);
and AND2 (N5766, N5702, N4889);
buf BUF1 (N5767, N5760);
nand NAND3 (N5768, N5765, N5399, N5148);
not NOT1 (N5769, N5764);
nand NAND3 (N5770, N5742, N1809, N1325);
nand NAND3 (N5771, N5741, N2320, N5532);
nand NAND4 (N5772, N5768, N3288, N4701, N1764);
buf BUF1 (N5773, N5766);
and AND3 (N5774, N5754, N2826, N4272);
xor XOR2 (N5775, N5761, N3774);
nor NOR3 (N5776, N5763, N3890, N4636);
nand NAND4 (N5777, N5770, N1792, N1936, N4659);
nand NAND3 (N5778, N5774, N551, N5191);
not NOT1 (N5779, N5767);
xor XOR2 (N5780, N5769, N960);
not NOT1 (N5781, N5771);
and AND3 (N5782, N5738, N1150, N3556);
and AND3 (N5783, N5780, N5643, N802);
xor XOR2 (N5784, N5777, N2100);
not NOT1 (N5785, N5776);
nor NOR2 (N5786, N5773, N5249);
or OR2 (N5787, N5782, N729);
or OR3 (N5788, N5783, N2887, N1303);
buf BUF1 (N5789, N5785);
or OR4 (N5790, N5788, N1529, N4032, N1346);
nor NOR4 (N5791, N5779, N3118, N1408, N2115);
or OR4 (N5792, N5772, N4362, N2456, N4546);
buf BUF1 (N5793, N5791);
or OR2 (N5794, N5787, N696);
buf BUF1 (N5795, N5790);
nand NAND4 (N5796, N5781, N475, N5063, N2200);
and AND2 (N5797, N5793, N4447);
not NOT1 (N5798, N5796);
nor NOR4 (N5799, N5797, N901, N323, N970);
and AND2 (N5800, N5784, N1642);
buf BUF1 (N5801, N5778);
buf BUF1 (N5802, N5792);
xor XOR2 (N5803, N5786, N1188);
and AND4 (N5804, N5800, N5701, N3242, N3326);
buf BUF1 (N5805, N5799);
nand NAND2 (N5806, N5804, N1402);
and AND2 (N5807, N5806, N2126);
xor XOR2 (N5808, N5803, N2493);
nand NAND2 (N5809, N5794, N3765);
xor XOR2 (N5810, N5809, N1398);
nand NAND2 (N5811, N5801, N5117);
nand NAND3 (N5812, N5789, N1041, N4635);
and AND2 (N5813, N5805, N2848);
buf BUF1 (N5814, N5812);
and AND2 (N5815, N5795, N3238);
not NOT1 (N5816, N5808);
nor NOR4 (N5817, N5802, N942, N3794, N5542);
or OR2 (N5818, N5816, N881);
and AND3 (N5819, N5817, N2307, N934);
buf BUF1 (N5820, N5807);
buf BUF1 (N5821, N5820);
xor XOR2 (N5822, N5821, N5590);
not NOT1 (N5823, N5775);
or OR3 (N5824, N5798, N480, N2499);
xor XOR2 (N5825, N5824, N3365);
and AND4 (N5826, N5813, N2279, N1237, N5548);
not NOT1 (N5827, N5823);
and AND2 (N5828, N5827, N787);
or OR3 (N5829, N5828, N1373, N2409);
xor XOR2 (N5830, N5825, N4663);
buf BUF1 (N5831, N5822);
nor NOR2 (N5832, N5814, N5532);
or OR2 (N5833, N5811, N245);
or OR4 (N5834, N5810, N3620, N1033, N5228);
xor XOR2 (N5835, N5832, N2072);
nor NOR2 (N5836, N5831, N1409);
buf BUF1 (N5837, N5830);
xor XOR2 (N5838, N5835, N5822);
or OR4 (N5839, N5826, N3673, N5461, N5806);
nand NAND3 (N5840, N5829, N1524, N4074);
xor XOR2 (N5841, N5840, N3466);
nand NAND2 (N5842, N5836, N2447);
nor NOR2 (N5843, N5834, N5133);
nor NOR4 (N5844, N5839, N4031, N253, N4578);
xor XOR2 (N5845, N5842, N996);
and AND4 (N5846, N5844, N5073, N524, N2847);
and AND4 (N5847, N5837, N1016, N1789, N3228);
xor XOR2 (N5848, N5845, N2196);
not NOT1 (N5849, N5848);
or OR3 (N5850, N5847, N5364, N3623);
buf BUF1 (N5851, N5833);
nand NAND2 (N5852, N5850, N3414);
xor XOR2 (N5853, N5815, N5059);
and AND2 (N5854, N5838, N1585);
or OR2 (N5855, N5819, N3181);
nor NOR2 (N5856, N5851, N3109);
nor NOR3 (N5857, N5843, N2447, N743);
not NOT1 (N5858, N5855);
or OR4 (N5859, N5852, N4047, N5549, N4366);
not NOT1 (N5860, N5856);
nand NAND4 (N5861, N5860, N4056, N3848, N1204);
not NOT1 (N5862, N5841);
and AND2 (N5863, N5849, N573);
or OR4 (N5864, N5853, N194, N3227, N5229);
buf BUF1 (N5865, N5854);
and AND2 (N5866, N5861, N2247);
xor XOR2 (N5867, N5858, N5364);
xor XOR2 (N5868, N5863, N5449);
not NOT1 (N5869, N5859);
or OR2 (N5870, N5846, N3126);
or OR4 (N5871, N5864, N4393, N79, N3591);
nand NAND4 (N5872, N5868, N4114, N1390, N435);
buf BUF1 (N5873, N5866);
buf BUF1 (N5874, N5873);
nand NAND3 (N5875, N5862, N966, N4321);
buf BUF1 (N5876, N5818);
nor NOR3 (N5877, N5865, N1622, N4208);
and AND3 (N5878, N5867, N5247, N2073);
not NOT1 (N5879, N5876);
buf BUF1 (N5880, N5857);
or OR2 (N5881, N5871, N3803);
nor NOR3 (N5882, N5870, N4951, N1821);
or OR4 (N5883, N5872, N1796, N5060, N3743);
not NOT1 (N5884, N5877);
or OR4 (N5885, N5879, N2864, N383, N2932);
not NOT1 (N5886, N5874);
xor XOR2 (N5887, N5869, N1986);
nor NOR4 (N5888, N5875, N92, N147, N1967);
nand NAND3 (N5889, N5883, N2817, N1145);
or OR2 (N5890, N5878, N120);
not NOT1 (N5891, N5881);
buf BUF1 (N5892, N5885);
xor XOR2 (N5893, N5886, N3363);
not NOT1 (N5894, N5880);
and AND4 (N5895, N5891, N4394, N1946, N4021);
nand NAND2 (N5896, N5890, N5874);
nand NAND2 (N5897, N5893, N1393);
buf BUF1 (N5898, N5889);
buf BUF1 (N5899, N5882);
not NOT1 (N5900, N5894);
and AND2 (N5901, N5888, N2106);
buf BUF1 (N5902, N5896);
or OR3 (N5903, N5899, N3616, N5652);
buf BUF1 (N5904, N5898);
and AND4 (N5905, N5902, N4688, N1861, N5516);
nand NAND2 (N5906, N5900, N3814);
or OR4 (N5907, N5897, N2319, N700, N1736);
nor NOR2 (N5908, N5905, N2008);
or OR2 (N5909, N5908, N4008);
nor NOR3 (N5910, N5887, N259, N1003);
and AND4 (N5911, N5909, N4669, N1115, N1876);
not NOT1 (N5912, N5904);
nor NOR2 (N5913, N5911, N2927);
buf BUF1 (N5914, N5892);
and AND2 (N5915, N5910, N2322);
and AND4 (N5916, N5895, N5407, N3672, N4335);
nor NOR3 (N5917, N5913, N1258, N3823);
buf BUF1 (N5918, N5916);
xor XOR2 (N5919, N5915, N3047);
buf BUF1 (N5920, N5884);
buf BUF1 (N5921, N5912);
or OR2 (N5922, N5914, N5206);
not NOT1 (N5923, N5906);
xor XOR2 (N5924, N5923, N1097);
buf BUF1 (N5925, N5903);
or OR2 (N5926, N5901, N4732);
nor NOR2 (N5927, N5921, N2149);
nand NAND2 (N5928, N5926, N1905);
xor XOR2 (N5929, N5925, N4206);
nor NOR2 (N5930, N5920, N1463);
nor NOR4 (N5931, N5924, N2242, N4915, N1020);
nand NAND4 (N5932, N5919, N4782, N1393, N355);
nand NAND3 (N5933, N5929, N5830, N1951);
nor NOR4 (N5934, N5931, N1558, N3989, N3954);
xor XOR2 (N5935, N5907, N4102);
xor XOR2 (N5936, N5932, N3487);
and AND3 (N5937, N5928, N2507, N696);
nand NAND3 (N5938, N5922, N3055, N4634);
nand NAND3 (N5939, N5934, N1982, N1778);
or OR4 (N5940, N5930, N523, N2671, N2100);
not NOT1 (N5941, N5918);
and AND3 (N5942, N5935, N1819, N4413);
not NOT1 (N5943, N5927);
not NOT1 (N5944, N5942);
buf BUF1 (N5945, N5944);
nand NAND2 (N5946, N5933, N5784);
or OR3 (N5947, N5937, N2023, N4993);
not NOT1 (N5948, N5946);
buf BUF1 (N5949, N5936);
buf BUF1 (N5950, N5917);
or OR3 (N5951, N5947, N1267, N566);
xor XOR2 (N5952, N5939, N4251);
or OR4 (N5953, N5948, N4398, N5338, N4624);
buf BUF1 (N5954, N5951);
buf BUF1 (N5955, N5945);
or OR2 (N5956, N5940, N5364);
buf BUF1 (N5957, N5956);
or OR3 (N5958, N5953, N304, N4803);
and AND3 (N5959, N5952, N5461, N763);
nor NOR4 (N5960, N5938, N1753, N2408, N2051);
not NOT1 (N5961, N5955);
and AND3 (N5962, N5960, N4069, N4706);
or OR2 (N5963, N5957, N4885);
not NOT1 (N5964, N5943);
nand NAND4 (N5965, N5962, N705, N673, N2848);
and AND4 (N5966, N5954, N2923, N1915, N1235);
nand NAND3 (N5967, N5941, N2331, N3565);
and AND2 (N5968, N5967, N3155);
buf BUF1 (N5969, N5949);
nor NOR2 (N5970, N5950, N3873);
buf BUF1 (N5971, N5966);
xor XOR2 (N5972, N5959, N1466);
nand NAND3 (N5973, N5964, N5661, N4256);
and AND4 (N5974, N5972, N4155, N5245, N4857);
and AND4 (N5975, N5970, N1300, N3962, N4536);
or OR4 (N5976, N5968, N2597, N510, N4053);
xor XOR2 (N5977, N5974, N374);
nand NAND3 (N5978, N5976, N5930, N1108);
nand NAND2 (N5979, N5963, N1589);
or OR2 (N5980, N5977, N1891);
buf BUF1 (N5981, N5958);
not NOT1 (N5982, N5971);
xor XOR2 (N5983, N5980, N5242);
and AND2 (N5984, N5969, N1377);
nand NAND3 (N5985, N5965, N3624, N4586);
nor NOR4 (N5986, N5961, N3644, N452, N2681);
nand NAND4 (N5987, N5983, N5967, N4088, N5544);
and AND2 (N5988, N5985, N1197);
or OR2 (N5989, N5982, N4821);
and AND4 (N5990, N5987, N3736, N5256, N1802);
and AND3 (N5991, N5981, N943, N2134);
and AND4 (N5992, N5975, N2453, N4433, N5194);
or OR2 (N5993, N5986, N2762);
not NOT1 (N5994, N5973);
and AND3 (N5995, N5978, N2691, N309);
nor NOR2 (N5996, N5995, N5323);
or OR4 (N5997, N5989, N3073, N3801, N4734);
nor NOR3 (N5998, N5991, N4027, N4985);
nor NOR4 (N5999, N5990, N693, N4977, N5419);
and AND4 (N6000, N5993, N2972, N5380, N4179);
nand NAND2 (N6001, N5994, N5532);
xor XOR2 (N6002, N5984, N2481);
nor NOR2 (N6003, N5999, N698);
nor NOR4 (N6004, N6000, N1739, N1372, N1353);
buf BUF1 (N6005, N6001);
nor NOR4 (N6006, N5979, N4581, N5082, N3461);
nand NAND3 (N6007, N5992, N4438, N5335);
or OR3 (N6008, N6003, N1223, N5668);
buf BUF1 (N6009, N5996);
and AND2 (N6010, N6007, N3296);
nor NOR3 (N6011, N5997, N2577, N1674);
not NOT1 (N6012, N6005);
xor XOR2 (N6013, N6010, N5869);
or OR3 (N6014, N6012, N3262, N4561);
xor XOR2 (N6015, N6011, N5462);
nor NOR3 (N6016, N6004, N1223, N5786);
xor XOR2 (N6017, N6016, N1287);
and AND2 (N6018, N6015, N5371);
nor NOR2 (N6019, N6017, N5873);
nor NOR4 (N6020, N6018, N4845, N4322, N3357);
nand NAND2 (N6021, N5988, N3257);
or OR3 (N6022, N6021, N981, N5091);
or OR3 (N6023, N6008, N4194, N4091);
buf BUF1 (N6024, N6022);
buf BUF1 (N6025, N6020);
nand NAND2 (N6026, N6023, N3484);
buf BUF1 (N6027, N6009);
nand NAND4 (N6028, N6002, N4639, N3026, N488);
and AND2 (N6029, N6028, N4824);
not NOT1 (N6030, N5998);
xor XOR2 (N6031, N6025, N5404);
not NOT1 (N6032, N6014);
not NOT1 (N6033, N6026);
xor XOR2 (N6034, N6019, N4578);
not NOT1 (N6035, N6032);
nand NAND4 (N6036, N6013, N899, N1825, N2246);
xor XOR2 (N6037, N6033, N4153);
buf BUF1 (N6038, N6035);
and AND3 (N6039, N6006, N10, N2498);
nor NOR3 (N6040, N6027, N4133, N3312);
and AND3 (N6041, N6030, N1241, N2196);
nand NAND3 (N6042, N6040, N1119, N1878);
buf BUF1 (N6043, N6041);
nand NAND3 (N6044, N6043, N5192, N5776);
nor NOR3 (N6045, N6024, N2148, N835);
not NOT1 (N6046, N6038);
not NOT1 (N6047, N6037);
nand NAND3 (N6048, N6039, N28, N133);
nand NAND4 (N6049, N6029, N1771, N1416, N2121);
xor XOR2 (N6050, N6034, N2088);
not NOT1 (N6051, N6045);
buf BUF1 (N6052, N6036);
nand NAND2 (N6053, N6046, N2778);
xor XOR2 (N6054, N6031, N1762);
and AND3 (N6055, N6049, N4760, N1138);
buf BUF1 (N6056, N6053);
and AND3 (N6057, N6048, N1180, N3938);
nor NOR2 (N6058, N6055, N3234);
nor NOR4 (N6059, N6058, N4912, N3976, N1718);
not NOT1 (N6060, N6056);
nor NOR3 (N6061, N6042, N4565, N2503);
nor NOR4 (N6062, N6052, N1794, N2181, N4496);
xor XOR2 (N6063, N6061, N2709);
not NOT1 (N6064, N6059);
nor NOR4 (N6065, N6057, N5586, N3200, N4913);
xor XOR2 (N6066, N6065, N4080);
buf BUF1 (N6067, N6062);
and AND2 (N6068, N6054, N467);
nor NOR4 (N6069, N6063, N5850, N3650, N1278);
not NOT1 (N6070, N6050);
nand NAND2 (N6071, N6067, N4628);
or OR2 (N6072, N6069, N1080);
buf BUF1 (N6073, N6064);
not NOT1 (N6074, N6044);
not NOT1 (N6075, N6073);
nand NAND3 (N6076, N6071, N2052, N3476);
buf BUF1 (N6077, N6074);
xor XOR2 (N6078, N6060, N344);
nor NOR3 (N6079, N6075, N5791, N1567);
or OR4 (N6080, N6068, N4154, N3705, N1833);
nand NAND4 (N6081, N6076, N5311, N3722, N5267);
not NOT1 (N6082, N6066);
buf BUF1 (N6083, N6077);
nand NAND3 (N6084, N6070, N351, N610);
nand NAND2 (N6085, N6080, N1178);
nor NOR2 (N6086, N6051, N5968);
buf BUF1 (N6087, N6084);
buf BUF1 (N6088, N6072);
not NOT1 (N6089, N6083);
nor NOR4 (N6090, N6081, N2297, N1350, N3185);
and AND3 (N6091, N6089, N2865, N5120);
buf BUF1 (N6092, N6079);
and AND3 (N6093, N6091, N4367, N4162);
nor NOR3 (N6094, N6085, N2795, N4220);
buf BUF1 (N6095, N6082);
nand NAND3 (N6096, N6047, N3500, N5436);
not NOT1 (N6097, N6095);
not NOT1 (N6098, N6090);
nor NOR3 (N6099, N6087, N4505, N5592);
nor NOR3 (N6100, N6097, N5215, N2080);
and AND3 (N6101, N6099, N2080, N1473);
and AND2 (N6102, N6101, N2584);
nor NOR3 (N6103, N6078, N214, N3761);
or OR4 (N6104, N6086, N4641, N5456, N187);
xor XOR2 (N6105, N6098, N1351);
nand NAND2 (N6106, N6092, N3139);
buf BUF1 (N6107, N6088);
or OR4 (N6108, N6103, N2550, N1473, N3719);
nor NOR4 (N6109, N6105, N5326, N1424, N559);
nand NAND2 (N6110, N6100, N4337);
or OR2 (N6111, N6110, N2214);
xor XOR2 (N6112, N6106, N4478);
or OR2 (N6113, N6107, N1879);
buf BUF1 (N6114, N6096);
nor NOR4 (N6115, N6102, N5008, N5214, N2596);
and AND2 (N6116, N6111, N5034);
xor XOR2 (N6117, N6094, N176);
buf BUF1 (N6118, N6109);
and AND3 (N6119, N6113, N5287, N2814);
xor XOR2 (N6120, N6118, N4342);
buf BUF1 (N6121, N6116);
not NOT1 (N6122, N6117);
nor NOR3 (N6123, N6121, N2640, N2916);
buf BUF1 (N6124, N6120);
nand NAND3 (N6125, N6123, N569, N5521);
or OR4 (N6126, N6125, N4401, N644, N3352);
not NOT1 (N6127, N6114);
and AND3 (N6128, N6104, N1853, N3334);
xor XOR2 (N6129, N6126, N2134);
not NOT1 (N6130, N6129);
xor XOR2 (N6131, N6127, N212);
nand NAND3 (N6132, N6128, N1509, N2269);
or OR2 (N6133, N6112, N6125);
not NOT1 (N6134, N6133);
or OR3 (N6135, N6115, N5189, N695);
not NOT1 (N6136, N6124);
nand NAND2 (N6137, N6119, N5987);
nor NOR2 (N6138, N6134, N1284);
not NOT1 (N6139, N6122);
and AND3 (N6140, N6139, N3106, N615);
not NOT1 (N6141, N6135);
nor NOR4 (N6142, N6131, N3524, N5558, N1613);
nand NAND2 (N6143, N6142, N1578);
or OR4 (N6144, N6130, N914, N4446, N424);
or OR4 (N6145, N6138, N1330, N3378, N1628);
buf BUF1 (N6146, N6144);
xor XOR2 (N6147, N6132, N4282);
not NOT1 (N6148, N6147);
not NOT1 (N6149, N6108);
xor XOR2 (N6150, N6145, N1059);
not NOT1 (N6151, N6143);
or OR2 (N6152, N6150, N4444);
xor XOR2 (N6153, N6093, N1948);
and AND2 (N6154, N6146, N224);
not NOT1 (N6155, N6137);
xor XOR2 (N6156, N6155, N469);
xor XOR2 (N6157, N6141, N150);
buf BUF1 (N6158, N6136);
nor NOR4 (N6159, N6140, N498, N5143, N1209);
nand NAND2 (N6160, N6148, N4218);
or OR2 (N6161, N6152, N1825);
xor XOR2 (N6162, N6159, N4440);
xor XOR2 (N6163, N6160, N6050);
xor XOR2 (N6164, N6161, N3096);
xor XOR2 (N6165, N6164, N1449);
buf BUF1 (N6166, N6163);
nor NOR4 (N6167, N6149, N1338, N1677, N4140);
or OR3 (N6168, N6165, N3994, N5555);
xor XOR2 (N6169, N6153, N1049);
buf BUF1 (N6170, N6156);
or OR2 (N6171, N6162, N1579);
buf BUF1 (N6172, N6151);
xor XOR2 (N6173, N6171, N139);
xor XOR2 (N6174, N6158, N793);
nand NAND2 (N6175, N6170, N4011);
xor XOR2 (N6176, N6172, N2740);
not NOT1 (N6177, N6176);
nor NOR4 (N6178, N6166, N4205, N692, N427);
xor XOR2 (N6179, N6169, N5680);
buf BUF1 (N6180, N6178);
xor XOR2 (N6181, N6177, N6093);
not NOT1 (N6182, N6168);
buf BUF1 (N6183, N6182);
nor NOR3 (N6184, N6180, N2554, N5543);
xor XOR2 (N6185, N6184, N2428);
nor NOR2 (N6186, N6185, N5022);
and AND2 (N6187, N6183, N2555);
buf BUF1 (N6188, N6187);
nor NOR2 (N6189, N6173, N2406);
nor NOR4 (N6190, N6174, N4070, N5531, N5156);
xor XOR2 (N6191, N6175, N2488);
nor NOR4 (N6192, N6190, N906, N2799, N4462);
and AND3 (N6193, N6192, N4688, N5410);
or OR3 (N6194, N6179, N5062, N1203);
or OR4 (N6195, N6193, N5056, N2026, N5508);
nor NOR3 (N6196, N6191, N5581, N2);
nand NAND2 (N6197, N6196, N2447);
and AND3 (N6198, N6181, N5476, N4667);
not NOT1 (N6199, N6189);
nand NAND2 (N6200, N6186, N237);
or OR4 (N6201, N6200, N5692, N2670, N1146);
buf BUF1 (N6202, N6198);
nor NOR3 (N6203, N6157, N1679, N2483);
buf BUF1 (N6204, N6154);
or OR3 (N6205, N6195, N3543, N471);
nor NOR4 (N6206, N6201, N1236, N1525, N819);
xor XOR2 (N6207, N6197, N379);
and AND4 (N6208, N6199, N134, N1492, N4802);
nand NAND2 (N6209, N6202, N1912);
or OR2 (N6210, N6204, N1481);
buf BUF1 (N6211, N6208);
and AND4 (N6212, N6206, N1585, N4491, N3063);
nor NOR4 (N6213, N6210, N3287, N4075, N482);
or OR4 (N6214, N6188, N5751, N331, N5324);
or OR3 (N6215, N6167, N5600, N1493);
not NOT1 (N6216, N6203);
not NOT1 (N6217, N6211);
and AND2 (N6218, N6205, N3323);
buf BUF1 (N6219, N6216);
xor XOR2 (N6220, N6218, N1411);
and AND2 (N6221, N6220, N2310);
nand NAND2 (N6222, N6214, N1075);
or OR3 (N6223, N6221, N1445, N3934);
buf BUF1 (N6224, N6207);
xor XOR2 (N6225, N6194, N3400);
xor XOR2 (N6226, N6225, N1742);
nand NAND4 (N6227, N6223, N2155, N1050, N5338);
not NOT1 (N6228, N6222);
and AND3 (N6229, N6219, N2932, N2222);
not NOT1 (N6230, N6215);
buf BUF1 (N6231, N6213);
and AND4 (N6232, N6228, N2930, N4875, N5939);
xor XOR2 (N6233, N6232, N1423);
not NOT1 (N6234, N6227);
xor XOR2 (N6235, N6234, N6146);
xor XOR2 (N6236, N6212, N1903);
nand NAND3 (N6237, N6236, N5878, N2268);
buf BUF1 (N6238, N6209);
or OR3 (N6239, N6217, N4002, N4149);
buf BUF1 (N6240, N6231);
xor XOR2 (N6241, N6237, N5055);
nand NAND3 (N6242, N6229, N3584, N2242);
nor NOR2 (N6243, N6239, N3918);
nor NOR4 (N6244, N6230, N5628, N240, N4961);
nand NAND4 (N6245, N6235, N1743, N1898, N1342);
buf BUF1 (N6246, N6233);
nor NOR4 (N6247, N6245, N2455, N3136, N2548);
and AND4 (N6248, N6243, N1636, N2685, N5530);
buf BUF1 (N6249, N6224);
buf BUF1 (N6250, N6246);
nand NAND2 (N6251, N6240, N1620);
or OR4 (N6252, N6251, N880, N5697, N1554);
and AND3 (N6253, N6242, N4214, N3148);
not NOT1 (N6254, N6249);
nor NOR4 (N6255, N6254, N2105, N112, N2251);
nor NOR2 (N6256, N6250, N2381);
or OR4 (N6257, N6253, N3989, N2517, N4986);
not NOT1 (N6258, N6256);
xor XOR2 (N6259, N6258, N4710);
not NOT1 (N6260, N6248);
and AND4 (N6261, N6252, N5617, N5313, N529);
xor XOR2 (N6262, N6238, N4038);
nor NOR3 (N6263, N6259, N3230, N5356);
or OR4 (N6264, N6261, N672, N1700, N5716);
xor XOR2 (N6265, N6263, N1753);
not NOT1 (N6266, N6247);
and AND3 (N6267, N6264, N4317, N6122);
xor XOR2 (N6268, N6267, N5875);
buf BUF1 (N6269, N6265);
or OR3 (N6270, N6226, N1224, N2523);
and AND4 (N6271, N6244, N5600, N631, N5645);
nand NAND3 (N6272, N6241, N4607, N1657);
and AND3 (N6273, N6272, N5521, N3499);
nor NOR4 (N6274, N6269, N764, N5277, N2703);
not NOT1 (N6275, N6257);
and AND4 (N6276, N6268, N427, N5980, N4938);
and AND4 (N6277, N6262, N2184, N1578, N5734);
nor NOR4 (N6278, N6276, N1800, N5593, N4558);
nand NAND4 (N6279, N6260, N281, N3651, N3072);
nand NAND4 (N6280, N6279, N4391, N6151, N5703);
buf BUF1 (N6281, N6270);
not NOT1 (N6282, N6271);
and AND3 (N6283, N6277, N2843, N2338);
and AND4 (N6284, N6275, N3948, N2268, N1422);
nor NOR2 (N6285, N6273, N3370);
or OR2 (N6286, N6280, N4715);
not NOT1 (N6287, N6283);
buf BUF1 (N6288, N6287);
buf BUF1 (N6289, N6282);
and AND3 (N6290, N6285, N197, N2972);
nand NAND2 (N6291, N6284, N2742);
xor XOR2 (N6292, N6266, N3804);
and AND2 (N6293, N6286, N5984);
buf BUF1 (N6294, N6274);
xor XOR2 (N6295, N6278, N4972);
buf BUF1 (N6296, N6288);
buf BUF1 (N6297, N6291);
buf BUF1 (N6298, N6292);
not NOT1 (N6299, N6296);
not NOT1 (N6300, N6295);
and AND3 (N6301, N6293, N2202, N3564);
nor NOR2 (N6302, N6300, N795);
nor NOR2 (N6303, N6289, N3934);
or OR3 (N6304, N6281, N1539, N5797);
buf BUF1 (N6305, N6303);
not NOT1 (N6306, N6297);
or OR2 (N6307, N6255, N1601);
nor NOR2 (N6308, N6290, N3148);
nand NAND4 (N6309, N6298, N2635, N3357, N4340);
xor XOR2 (N6310, N6294, N1925);
buf BUF1 (N6311, N6299);
xor XOR2 (N6312, N6307, N5838);
and AND3 (N6313, N6302, N2425, N3192);
nand NAND3 (N6314, N6309, N2851, N5825);
or OR4 (N6315, N6310, N1232, N895, N3931);
or OR4 (N6316, N6314, N548, N2834, N4136);
and AND2 (N6317, N6313, N1070);
buf BUF1 (N6318, N6315);
and AND4 (N6319, N6316, N242, N1279, N2148);
or OR2 (N6320, N6318, N5935);
nor NOR3 (N6321, N6305, N3191, N6060);
or OR3 (N6322, N6319, N4646, N4849);
nand NAND2 (N6323, N6322, N2894);
buf BUF1 (N6324, N6306);
nor NOR4 (N6325, N6323, N3735, N2722, N1706);
buf BUF1 (N6326, N6312);
not NOT1 (N6327, N6326);
nor NOR3 (N6328, N6304, N5584, N6222);
nor NOR4 (N6329, N6328, N1350, N2361, N26);
xor XOR2 (N6330, N6308, N3032);
nand NAND4 (N6331, N6330, N2830, N470, N1558);
not NOT1 (N6332, N6301);
nand NAND3 (N6333, N6324, N4598, N3812);
xor XOR2 (N6334, N6311, N4724);
xor XOR2 (N6335, N6317, N1473);
nand NAND2 (N6336, N6329, N4483);
or OR3 (N6337, N6320, N4233, N3582);
nand NAND3 (N6338, N6321, N1255, N26);
nand NAND2 (N6339, N6325, N1762);
nand NAND2 (N6340, N6327, N3798);
buf BUF1 (N6341, N6334);
xor XOR2 (N6342, N6333, N4333);
nor NOR4 (N6343, N6341, N3770, N3877, N3812);
nor NOR3 (N6344, N6342, N4178, N3015);
and AND4 (N6345, N6336, N2645, N818, N3482);
not NOT1 (N6346, N6345);
nand NAND3 (N6347, N6344, N1677, N4753);
xor XOR2 (N6348, N6332, N1892);
buf BUF1 (N6349, N6347);
not NOT1 (N6350, N6338);
and AND3 (N6351, N6346, N415, N4794);
buf BUF1 (N6352, N6339);
xor XOR2 (N6353, N6337, N4303);
nand NAND4 (N6354, N6349, N3012, N5270, N4426);
nor NOR3 (N6355, N6354, N3414, N5629);
not NOT1 (N6356, N6353);
xor XOR2 (N6357, N6335, N1711);
not NOT1 (N6358, N6343);
or OR2 (N6359, N6331, N2499);
xor XOR2 (N6360, N6348, N4836);
xor XOR2 (N6361, N6350, N2472);
and AND3 (N6362, N6361, N2848, N2867);
or OR3 (N6363, N6352, N5444, N5999);
buf BUF1 (N6364, N6359);
buf BUF1 (N6365, N6360);
xor XOR2 (N6366, N6357, N3926);
not NOT1 (N6367, N6356);
buf BUF1 (N6368, N6366);
nand NAND3 (N6369, N6355, N5280, N5269);
nor NOR3 (N6370, N6367, N5602, N1529);
nand NAND4 (N6371, N6364, N5278, N6253, N4565);
buf BUF1 (N6372, N6351);
not NOT1 (N6373, N6362);
and AND3 (N6374, N6373, N2391, N5417);
buf BUF1 (N6375, N6374);
nor NOR3 (N6376, N6365, N311, N4644);
xor XOR2 (N6377, N6368, N4223);
nand NAND3 (N6378, N6372, N2, N1957);
nand NAND4 (N6379, N6340, N5126, N3514, N4203);
nand NAND4 (N6380, N6378, N1278, N304, N3923);
nand NAND3 (N6381, N6369, N1943, N1449);
buf BUF1 (N6382, N6376);
nor NOR3 (N6383, N6377, N852, N1863);
nand NAND2 (N6384, N6375, N350);
nor NOR3 (N6385, N6363, N5556, N234);
xor XOR2 (N6386, N6370, N5754);
xor XOR2 (N6387, N6385, N2555);
nand NAND3 (N6388, N6381, N4224, N542);
nand NAND4 (N6389, N6388, N102, N1832, N1398);
or OR2 (N6390, N6386, N3973);
nor NOR2 (N6391, N6384, N2396);
nand NAND4 (N6392, N6389, N1236, N6328, N5005);
or OR4 (N6393, N6382, N3586, N1704, N3286);
nand NAND3 (N6394, N6392, N3743, N855);
nor NOR3 (N6395, N6394, N1582, N4298);
xor XOR2 (N6396, N6383, N2622);
and AND4 (N6397, N6380, N6171, N3424, N6064);
xor XOR2 (N6398, N6396, N4234);
nand NAND3 (N6399, N6391, N6390, N2266);
nand NAND4 (N6400, N4759, N851, N4866, N2384);
not NOT1 (N6401, N6399);
not NOT1 (N6402, N6379);
not NOT1 (N6403, N6387);
not NOT1 (N6404, N6403);
nor NOR4 (N6405, N6401, N2787, N4374, N5770);
and AND2 (N6406, N6358, N871);
xor XOR2 (N6407, N6393, N5414);
and AND3 (N6408, N6405, N6131, N2735);
nand NAND4 (N6409, N6400, N3130, N2748, N3913);
xor XOR2 (N6410, N6406, N4384);
not NOT1 (N6411, N6404);
or OR2 (N6412, N6407, N1316);
and AND2 (N6413, N6398, N781);
and AND2 (N6414, N6411, N6170);
xor XOR2 (N6415, N6412, N2566);
and AND2 (N6416, N6402, N5279);
xor XOR2 (N6417, N6371, N3158);
buf BUF1 (N6418, N6414);
buf BUF1 (N6419, N6410);
not NOT1 (N6420, N6418);
buf BUF1 (N6421, N6417);
buf BUF1 (N6422, N6415);
xor XOR2 (N6423, N6422, N4460);
and AND4 (N6424, N6395, N847, N6309, N2733);
nand NAND3 (N6425, N6416, N3432, N1636);
buf BUF1 (N6426, N6419);
and AND3 (N6427, N6397, N1863, N3939);
not NOT1 (N6428, N6423);
and AND4 (N6429, N6428, N4184, N3072, N4455);
xor XOR2 (N6430, N6426, N272);
not NOT1 (N6431, N6421);
xor XOR2 (N6432, N6429, N722);
not NOT1 (N6433, N6431);
not NOT1 (N6434, N6432);
xor XOR2 (N6435, N6424, N1079);
xor XOR2 (N6436, N6425, N4995);
and AND2 (N6437, N6433, N1532);
nor NOR3 (N6438, N6434, N1171, N5835);
not NOT1 (N6439, N6427);
and AND3 (N6440, N6439, N4936, N1622);
nor NOR2 (N6441, N6440, N6115);
and AND4 (N6442, N6436, N357, N3799, N4759);
and AND4 (N6443, N6438, N5742, N3459, N6073);
or OR3 (N6444, N6413, N957, N3421);
nand NAND2 (N6445, N6444, N1167);
xor XOR2 (N6446, N6437, N164);
or OR2 (N6447, N6409, N2733);
buf BUF1 (N6448, N6447);
not NOT1 (N6449, N6420);
nor NOR3 (N6450, N6448, N139, N5058);
or OR2 (N6451, N6450, N2541);
nor NOR4 (N6452, N6430, N4571, N541, N2526);
not NOT1 (N6453, N6452);
or OR3 (N6454, N6443, N1361, N392);
not NOT1 (N6455, N6445);
xor XOR2 (N6456, N6446, N1199);
buf BUF1 (N6457, N6456);
not NOT1 (N6458, N6441);
xor XOR2 (N6459, N6442, N5488);
nand NAND2 (N6460, N6451, N6352);
and AND4 (N6461, N6454, N3852, N3818, N3538);
xor XOR2 (N6462, N6455, N4260);
and AND2 (N6463, N6449, N2546);
nand NAND3 (N6464, N6453, N4849, N4221);
and AND2 (N6465, N6461, N2779);
buf BUF1 (N6466, N6435);
and AND4 (N6467, N6457, N6119, N5989, N3417);
not NOT1 (N6468, N6408);
and AND4 (N6469, N6463, N3143, N184, N343);
nand NAND3 (N6470, N6464, N6102, N667);
nor NOR3 (N6471, N6459, N793, N3223);
and AND2 (N6472, N6467, N3397);
not NOT1 (N6473, N6460);
and AND2 (N6474, N6462, N545);
buf BUF1 (N6475, N6474);
buf BUF1 (N6476, N6466);
nor NOR2 (N6477, N6475, N3415);
or OR3 (N6478, N6472, N979, N4314);
nor NOR3 (N6479, N6478, N5157, N5321);
and AND2 (N6480, N6473, N3822);
nor NOR2 (N6481, N6477, N5212);
and AND3 (N6482, N6465, N1272, N6430);
nand NAND2 (N6483, N6482, N732);
xor XOR2 (N6484, N6458, N4415);
or OR3 (N6485, N6469, N6392, N6162);
not NOT1 (N6486, N6471);
and AND3 (N6487, N6476, N4079, N2033);
nor NOR3 (N6488, N6483, N6443, N5428);
not NOT1 (N6489, N6484);
nand NAND2 (N6490, N6481, N144);
or OR2 (N6491, N6487, N5883);
and AND4 (N6492, N6468, N6470, N4374, N982);
not NOT1 (N6493, N5219);
and AND2 (N6494, N6489, N35);
not NOT1 (N6495, N6492);
xor XOR2 (N6496, N6488, N5869);
nor NOR3 (N6497, N6491, N1091, N965);
nand NAND2 (N6498, N6493, N1843);
and AND4 (N6499, N6490, N2037, N4730, N5432);
buf BUF1 (N6500, N6486);
buf BUF1 (N6501, N6479);
nor NOR2 (N6502, N6485, N2526);
nand NAND2 (N6503, N6502, N5072);
xor XOR2 (N6504, N6496, N682);
not NOT1 (N6505, N6480);
nor NOR2 (N6506, N6500, N4264);
or OR3 (N6507, N6499, N2078, N5288);
or OR3 (N6508, N6505, N6223, N4812);
not NOT1 (N6509, N6494);
not NOT1 (N6510, N6509);
nor NOR4 (N6511, N6498, N5323, N2997, N5603);
not NOT1 (N6512, N6501);
nand NAND3 (N6513, N6508, N1048, N5470);
nand NAND2 (N6514, N6507, N867);
xor XOR2 (N6515, N6514, N5735);
and AND2 (N6516, N6506, N5071);
or OR3 (N6517, N6510, N404, N4984);
xor XOR2 (N6518, N6517, N3955);
nand NAND2 (N6519, N6516, N2418);
nand NAND2 (N6520, N6497, N2407);
buf BUF1 (N6521, N6503);
nor NOR3 (N6522, N6513, N5440, N3297);
xor XOR2 (N6523, N6522, N3908);
and AND4 (N6524, N6520, N4314, N2355, N1827);
xor XOR2 (N6525, N6523, N5004);
or OR2 (N6526, N6504, N2205);
nand NAND2 (N6527, N6521, N2749);
not NOT1 (N6528, N6495);
buf BUF1 (N6529, N6519);
buf BUF1 (N6530, N6515);
nand NAND4 (N6531, N6526, N4569, N3773, N4882);
xor XOR2 (N6532, N6528, N4183);
not NOT1 (N6533, N6527);
nand NAND3 (N6534, N6531, N6298, N2090);
and AND2 (N6535, N6512, N4732);
buf BUF1 (N6536, N6532);
and AND3 (N6537, N6525, N3463, N4291);
or OR3 (N6538, N6536, N2463, N1875);
buf BUF1 (N6539, N6535);
or OR4 (N6540, N6511, N6169, N2681, N946);
not NOT1 (N6541, N6534);
and AND4 (N6542, N6538, N752, N2300, N5027);
buf BUF1 (N6543, N6533);
buf BUF1 (N6544, N6529);
buf BUF1 (N6545, N6544);
xor XOR2 (N6546, N6541, N2747);
nand NAND4 (N6547, N6542, N5019, N2668, N3477);
buf BUF1 (N6548, N6547);
nand NAND3 (N6549, N6548, N2542, N6467);
or OR2 (N6550, N6518, N87);
or OR2 (N6551, N6549, N2385);
buf BUF1 (N6552, N6550);
xor XOR2 (N6553, N6543, N1858);
not NOT1 (N6554, N6545);
and AND2 (N6555, N6546, N1539);
nor NOR3 (N6556, N6552, N5006, N2672);
and AND4 (N6557, N6556, N4119, N1617, N5412);
nor NOR3 (N6558, N6554, N4414, N3114);
buf BUF1 (N6559, N6558);
xor XOR2 (N6560, N6559, N3268);
or OR2 (N6561, N6540, N523);
and AND3 (N6562, N6551, N614, N1678);
nand NAND2 (N6563, N6539, N1100);
nor NOR2 (N6564, N6562, N2802);
nand NAND2 (N6565, N6563, N4188);
or OR3 (N6566, N6553, N6324, N3368);
not NOT1 (N6567, N6566);
or OR3 (N6568, N6560, N5197, N3728);
nor NOR4 (N6569, N6537, N1182, N5353, N2283);
or OR2 (N6570, N6530, N5971);
or OR3 (N6571, N6555, N2811, N979);
buf BUF1 (N6572, N6568);
xor XOR2 (N6573, N6561, N2572);
or OR3 (N6574, N6571, N6215, N1343);
xor XOR2 (N6575, N6574, N3116);
nand NAND4 (N6576, N6572, N6170, N2817, N13);
or OR2 (N6577, N6569, N4703);
or OR3 (N6578, N6576, N4149, N5721);
or OR4 (N6579, N6524, N5031, N727, N853);
or OR4 (N6580, N6575, N3526, N4426, N3202);
not NOT1 (N6581, N6567);
and AND4 (N6582, N6577, N488, N2499, N24);
not NOT1 (N6583, N6565);
or OR4 (N6584, N6573, N3943, N504, N1164);
nor NOR4 (N6585, N6570, N2211, N5435, N3972);
nand NAND4 (N6586, N6564, N3866, N4816, N5037);
xor XOR2 (N6587, N6580, N248);
nand NAND3 (N6588, N6585, N2409, N4170);
not NOT1 (N6589, N6557);
or OR2 (N6590, N6588, N191);
or OR4 (N6591, N6586, N3166, N5688, N2280);
nand NAND2 (N6592, N6587, N4175);
xor XOR2 (N6593, N6584, N5037);
and AND2 (N6594, N6579, N5989);
buf BUF1 (N6595, N6592);
xor XOR2 (N6596, N6590, N1303);
xor XOR2 (N6597, N6583, N924);
and AND2 (N6598, N6589, N5968);
not NOT1 (N6599, N6582);
nand NAND4 (N6600, N6591, N3791, N6226, N1429);
xor XOR2 (N6601, N6600, N2864);
nand NAND3 (N6602, N6578, N5621, N3427);
not NOT1 (N6603, N6594);
nand NAND3 (N6604, N6603, N4974, N6159);
nand NAND2 (N6605, N6604, N4021);
nor NOR2 (N6606, N6601, N5300);
xor XOR2 (N6607, N6593, N468);
nor NOR4 (N6608, N6599, N3369, N4547, N1928);
nor NOR2 (N6609, N6606, N18);
xor XOR2 (N6610, N6598, N2170);
nand NAND2 (N6611, N6607, N2978);
nand NAND4 (N6612, N6609, N3009, N5264, N4960);
nand NAND4 (N6613, N6608, N3992, N4434, N3048);
not NOT1 (N6614, N6581);
or OR4 (N6615, N6611, N128, N6609, N5020);
xor XOR2 (N6616, N6595, N5009);
nor NOR2 (N6617, N6597, N6438);
not NOT1 (N6618, N6613);
not NOT1 (N6619, N6610);
buf BUF1 (N6620, N6605);
or OR3 (N6621, N6596, N291, N3732);
not NOT1 (N6622, N6621);
and AND2 (N6623, N6615, N1759);
xor XOR2 (N6624, N6622, N2340);
nor NOR2 (N6625, N6602, N5649);
nor NOR4 (N6626, N6616, N982, N2893, N5442);
nor NOR2 (N6627, N6619, N4788);
xor XOR2 (N6628, N6627, N3867);
nand NAND2 (N6629, N6618, N618);
and AND4 (N6630, N6626, N3893, N2271, N4635);
buf BUF1 (N6631, N6629);
nand NAND2 (N6632, N6614, N3944);
or OR2 (N6633, N6628, N443);
or OR4 (N6634, N6631, N3318, N3849, N887);
not NOT1 (N6635, N6617);
xor XOR2 (N6636, N6630, N3153);
and AND3 (N6637, N6623, N5627, N4153);
xor XOR2 (N6638, N6625, N6233);
and AND4 (N6639, N6637, N4775, N5950, N1593);
and AND4 (N6640, N6633, N2970, N4817, N1133);
xor XOR2 (N6641, N6632, N3772);
nor NOR2 (N6642, N6624, N4607);
or OR3 (N6643, N6636, N5407, N4669);
buf BUF1 (N6644, N6639);
buf BUF1 (N6645, N6643);
nand NAND4 (N6646, N6634, N5527, N4369, N6304);
xor XOR2 (N6647, N6638, N2230);
nand NAND3 (N6648, N6644, N681, N4185);
not NOT1 (N6649, N6641);
buf BUF1 (N6650, N6612);
and AND2 (N6651, N6620, N4640);
xor XOR2 (N6652, N6648, N1667);
nand NAND4 (N6653, N6650, N132, N2360, N5823);
or OR4 (N6654, N6635, N4620, N4124, N4446);
nor NOR2 (N6655, N6647, N2047);
nand NAND4 (N6656, N6655, N3309, N4044, N240);
nor NOR2 (N6657, N6649, N2126);
xor XOR2 (N6658, N6652, N1297);
or OR4 (N6659, N6658, N4022, N3256, N6170);
nand NAND3 (N6660, N6651, N3174, N2938);
buf BUF1 (N6661, N6654);
nor NOR3 (N6662, N6660, N636, N1414);
and AND4 (N6663, N6640, N5386, N3793, N1649);
xor XOR2 (N6664, N6656, N1067);
or OR3 (N6665, N6659, N4857, N6652);
nand NAND4 (N6666, N6661, N6320, N3447, N6610);
buf BUF1 (N6667, N6646);
or OR2 (N6668, N6667, N4877);
xor XOR2 (N6669, N6645, N381);
nand NAND3 (N6670, N6657, N4889, N3718);
buf BUF1 (N6671, N6669);
xor XOR2 (N6672, N6670, N6541);
or OR4 (N6673, N6671, N2816, N2153, N458);
or OR3 (N6674, N6673, N1083, N4354);
nand NAND4 (N6675, N6666, N4287, N3753, N18);
nor NOR2 (N6676, N6672, N6669);
nand NAND3 (N6677, N6663, N1766, N93);
and AND4 (N6678, N6676, N5174, N3865, N2945);
xor XOR2 (N6679, N6642, N1109);
and AND2 (N6680, N6665, N2439);
nor NOR2 (N6681, N6664, N5675);
or OR2 (N6682, N6680, N620);
not NOT1 (N6683, N6675);
nor NOR2 (N6684, N6678, N3443);
or OR3 (N6685, N6677, N3056, N1286);
xor XOR2 (N6686, N6674, N4383);
or OR3 (N6687, N6686, N553, N5581);
not NOT1 (N6688, N6681);
xor XOR2 (N6689, N6682, N3977);
and AND4 (N6690, N6683, N1627, N2627, N4312);
and AND4 (N6691, N6689, N2935, N2812, N5991);
not NOT1 (N6692, N6668);
not NOT1 (N6693, N6688);
not NOT1 (N6694, N6653);
and AND3 (N6695, N6685, N1976, N2369);
or OR4 (N6696, N6687, N3126, N670, N1543);
not NOT1 (N6697, N6662);
and AND4 (N6698, N6697, N2652, N5476, N2);
nand NAND2 (N6699, N6695, N3769);
nor NOR4 (N6700, N6698, N5336, N6480, N515);
not NOT1 (N6701, N6679);
xor XOR2 (N6702, N6700, N4011);
not NOT1 (N6703, N6701);
not NOT1 (N6704, N6694);
not NOT1 (N6705, N6691);
not NOT1 (N6706, N6692);
not NOT1 (N6707, N6702);
buf BUF1 (N6708, N6699);
xor XOR2 (N6709, N6693, N4011);
nand NAND3 (N6710, N6704, N5450, N5882);
not NOT1 (N6711, N6708);
or OR2 (N6712, N6711, N6230);
nand NAND4 (N6713, N6703, N6709, N356, N1499);
nor NOR4 (N6714, N5575, N3667, N6163, N6003);
and AND3 (N6715, N6690, N3087, N5968);
or OR2 (N6716, N6696, N1585);
not NOT1 (N6717, N6713);
xor XOR2 (N6718, N6706, N4526);
or OR4 (N6719, N6684, N5618, N4032, N6281);
not NOT1 (N6720, N6714);
not NOT1 (N6721, N6705);
buf BUF1 (N6722, N6707);
nand NAND3 (N6723, N6712, N5241, N4388);
not NOT1 (N6724, N6720);
not NOT1 (N6725, N6721);
nand NAND2 (N6726, N6725, N5815);
xor XOR2 (N6727, N6715, N339);
nand NAND4 (N6728, N6726, N4449, N5606, N1046);
nor NOR2 (N6729, N6719, N5759);
or OR2 (N6730, N6722, N2377);
or OR3 (N6731, N6710, N2093, N3406);
buf BUF1 (N6732, N6718);
and AND2 (N6733, N6717, N3240);
nor NOR4 (N6734, N6731, N5811, N118, N2703);
xor XOR2 (N6735, N6723, N6413);
or OR3 (N6736, N6727, N182, N1311);
buf BUF1 (N6737, N6724);
nor NOR2 (N6738, N6716, N517);
nor NOR4 (N6739, N6730, N5693, N866, N5169);
buf BUF1 (N6740, N6729);
nor NOR3 (N6741, N6734, N194, N2270);
xor XOR2 (N6742, N6739, N196);
and AND3 (N6743, N6733, N6430, N273);
buf BUF1 (N6744, N6743);
and AND2 (N6745, N6744, N2222);
and AND3 (N6746, N6735, N6290, N5389);
nand NAND3 (N6747, N6745, N6038, N3604);
buf BUF1 (N6748, N6736);
nor NOR2 (N6749, N6737, N3980);
not NOT1 (N6750, N6741);
nand NAND2 (N6751, N6740, N6072);
nand NAND2 (N6752, N6732, N3967);
and AND2 (N6753, N6749, N5111);
buf BUF1 (N6754, N6751);
and AND3 (N6755, N6754, N3833, N4635);
and AND2 (N6756, N6738, N5364);
not NOT1 (N6757, N6753);
nor NOR4 (N6758, N6752, N2808, N3519, N456);
nand NAND3 (N6759, N6757, N2758, N5176);
not NOT1 (N6760, N6755);
not NOT1 (N6761, N6746);
xor XOR2 (N6762, N6747, N426);
xor XOR2 (N6763, N6748, N6614);
and AND3 (N6764, N6750, N1651, N1959);
or OR2 (N6765, N6760, N4843);
nor NOR4 (N6766, N6762, N5786, N5999, N3839);
not NOT1 (N6767, N6766);
or OR2 (N6768, N6767, N2721);
nand NAND4 (N6769, N6768, N5116, N1382, N6031);
nand NAND3 (N6770, N6742, N1254, N1800);
nor NOR3 (N6771, N6728, N1652, N6232);
and AND2 (N6772, N6761, N5138);
not NOT1 (N6773, N6764);
not NOT1 (N6774, N6773);
not NOT1 (N6775, N6771);
not NOT1 (N6776, N6770);
buf BUF1 (N6777, N6759);
not NOT1 (N6778, N6774);
not NOT1 (N6779, N6769);
nand NAND2 (N6780, N6777, N339);
buf BUF1 (N6781, N6775);
xor XOR2 (N6782, N6763, N3815);
nor NOR4 (N6783, N6758, N2924, N417, N1551);
buf BUF1 (N6784, N6781);
and AND2 (N6785, N6778, N789);
buf BUF1 (N6786, N6765);
nor NOR4 (N6787, N6785, N6225, N5497, N792);
nor NOR4 (N6788, N6784, N3506, N1615, N6240);
nand NAND3 (N6789, N6780, N5885, N4894);
xor XOR2 (N6790, N6756, N5543);
nor NOR4 (N6791, N6788, N3766, N4394, N6139);
not NOT1 (N6792, N6783);
buf BUF1 (N6793, N6786);
or OR3 (N6794, N6790, N4919, N1130);
nand NAND3 (N6795, N6782, N5001, N2547);
nand NAND4 (N6796, N6789, N166, N1605, N142);
not NOT1 (N6797, N6794);
nor NOR2 (N6798, N6797, N132);
xor XOR2 (N6799, N6787, N4411);
not NOT1 (N6800, N6795);
nand NAND2 (N6801, N6793, N1931);
nand NAND4 (N6802, N6800, N1815, N492, N1061);
nor NOR4 (N6803, N6802, N4027, N4289, N3277);
xor XOR2 (N6804, N6792, N1899);
not NOT1 (N6805, N6779);
xor XOR2 (N6806, N6776, N3478);
or OR2 (N6807, N6804, N592);
and AND4 (N6808, N6791, N6374, N3352, N969);
not NOT1 (N6809, N6807);
nor NOR2 (N6810, N6796, N6100);
xor XOR2 (N6811, N6799, N4901);
buf BUF1 (N6812, N6801);
nor NOR3 (N6813, N6803, N4660, N1414);
xor XOR2 (N6814, N6813, N5891);
nor NOR2 (N6815, N6808, N5883);
nor NOR3 (N6816, N6815, N3405, N1557);
nand NAND2 (N6817, N6809, N2456);
not NOT1 (N6818, N6806);
not NOT1 (N6819, N6811);
or OR2 (N6820, N6816, N1311);
buf BUF1 (N6821, N6814);
xor XOR2 (N6822, N6812, N1819);
and AND4 (N6823, N6820, N6399, N1686, N165);
nor NOR4 (N6824, N6818, N2230, N6525, N6813);
not NOT1 (N6825, N6810);
nand NAND3 (N6826, N6805, N5068, N3079);
buf BUF1 (N6827, N6824);
buf BUF1 (N6828, N6819);
nor NOR2 (N6829, N6822, N381);
buf BUF1 (N6830, N6826);
or OR3 (N6831, N6827, N4157, N1957);
buf BUF1 (N6832, N6829);
and AND3 (N6833, N6772, N3150, N859);
or OR2 (N6834, N6828, N2881);
nand NAND2 (N6835, N6833, N1499);
or OR4 (N6836, N6798, N6097, N56, N3257);
xor XOR2 (N6837, N6825, N2551);
or OR4 (N6838, N6831, N2247, N3149, N399);
buf BUF1 (N6839, N6817);
xor XOR2 (N6840, N6830, N5713);
xor XOR2 (N6841, N6837, N319);
or OR2 (N6842, N6821, N5728);
not NOT1 (N6843, N6839);
not NOT1 (N6844, N6838);
buf BUF1 (N6845, N6823);
buf BUF1 (N6846, N6842);
not NOT1 (N6847, N6844);
nor NOR2 (N6848, N6846, N1130);
or OR3 (N6849, N6835, N3398, N3208);
not NOT1 (N6850, N6840);
nand NAND4 (N6851, N6845, N662, N2419, N4183);
xor XOR2 (N6852, N6847, N773);
nor NOR4 (N6853, N6850, N5485, N1611, N924);
nor NOR2 (N6854, N6836, N6562);
or OR2 (N6855, N6849, N905);
nand NAND3 (N6856, N6832, N5628, N1939);
not NOT1 (N6857, N6834);
or OR3 (N6858, N6841, N4907, N6691);
not NOT1 (N6859, N6848);
or OR2 (N6860, N6843, N1359);
buf BUF1 (N6861, N6852);
nand NAND2 (N6862, N6860, N191);
buf BUF1 (N6863, N6858);
buf BUF1 (N6864, N6854);
and AND3 (N6865, N6859, N2960, N3843);
or OR4 (N6866, N6862, N1240, N4979, N3628);
buf BUF1 (N6867, N6863);
xor XOR2 (N6868, N6867, N1415);
xor XOR2 (N6869, N6865, N5542);
nand NAND2 (N6870, N6869, N1480);
nor NOR3 (N6871, N6866, N4189, N5992);
not NOT1 (N6872, N6870);
and AND2 (N6873, N6853, N1052);
and AND4 (N6874, N6857, N3387, N144, N2246);
nand NAND3 (N6875, N6874, N705, N4143);
xor XOR2 (N6876, N6861, N5336);
not NOT1 (N6877, N6872);
nand NAND3 (N6878, N6871, N5730, N4177);
or OR4 (N6879, N6856, N2723, N4992, N4111);
nand NAND4 (N6880, N6873, N5641, N6412, N686);
or OR2 (N6881, N6877, N3959);
buf BUF1 (N6882, N6878);
nand NAND4 (N6883, N6864, N5111, N2577, N1365);
or OR3 (N6884, N6879, N4125, N1958);
or OR3 (N6885, N6868, N3861, N1593);
buf BUF1 (N6886, N6883);
or OR3 (N6887, N6875, N3691, N6783);
xor XOR2 (N6888, N6881, N5025);
nor NOR2 (N6889, N6885, N3214);
not NOT1 (N6890, N6855);
nor NOR2 (N6891, N6888, N5774);
xor XOR2 (N6892, N6886, N1959);
and AND2 (N6893, N6892, N6062);
nor NOR4 (N6894, N6890, N4585, N3429, N5074);
or OR3 (N6895, N6891, N5835, N3520);
or OR2 (N6896, N6884, N520);
not NOT1 (N6897, N6880);
or OR4 (N6898, N6876, N3688, N1506, N6872);
and AND3 (N6899, N6893, N3692, N4449);
nor NOR3 (N6900, N6896, N6683, N4941);
buf BUF1 (N6901, N6895);
nor NOR3 (N6902, N6899, N3284, N533);
nor NOR4 (N6903, N6889, N1982, N4164, N6251);
and AND3 (N6904, N6902, N5867, N6586);
and AND2 (N6905, N6887, N615);
buf BUF1 (N6906, N6904);
and AND3 (N6907, N6898, N2534, N6707);
not NOT1 (N6908, N6907);
nor NOR3 (N6909, N6905, N3879, N1550);
and AND4 (N6910, N6908, N6898, N6654, N5798);
not NOT1 (N6911, N6900);
buf BUF1 (N6912, N6894);
nand NAND2 (N6913, N6901, N407);
buf BUF1 (N6914, N6897);
xor XOR2 (N6915, N6912, N2049);
nand NAND3 (N6916, N6909, N6366, N5392);
and AND2 (N6917, N6851, N5990);
not NOT1 (N6918, N6882);
not NOT1 (N6919, N6914);
and AND4 (N6920, N6916, N1471, N1387, N1607);
nand NAND2 (N6921, N6910, N6054);
xor XOR2 (N6922, N6921, N4693);
not NOT1 (N6923, N6911);
nor NOR4 (N6924, N6913, N5018, N2488, N2919);
and AND2 (N6925, N6917, N4172);
xor XOR2 (N6926, N6906, N5160);
xor XOR2 (N6927, N6915, N4088);
buf BUF1 (N6928, N6924);
nand NAND3 (N6929, N6920, N3344, N1839);
or OR4 (N6930, N6927, N4170, N3620, N2909);
and AND3 (N6931, N6922, N5370, N2856);
xor XOR2 (N6932, N6930, N5994);
not NOT1 (N6933, N6928);
nor NOR4 (N6934, N6918, N2988, N1130, N1948);
buf BUF1 (N6935, N6929);
and AND2 (N6936, N6926, N258);
and AND2 (N6937, N6931, N1620);
xor XOR2 (N6938, N6923, N4476);
or OR4 (N6939, N6925, N3623, N2628, N5042);
not NOT1 (N6940, N6903);
nand NAND2 (N6941, N6938, N4346);
and AND2 (N6942, N6932, N1626);
and AND3 (N6943, N6934, N6500, N3925);
nor NOR3 (N6944, N6935, N5631, N6758);
nor NOR3 (N6945, N6942, N6208, N3062);
nor NOR3 (N6946, N6941, N2021, N3249);
xor XOR2 (N6947, N6937, N3066);
nor NOR3 (N6948, N6933, N605, N6247);
xor XOR2 (N6949, N6947, N5134);
not NOT1 (N6950, N6944);
or OR4 (N6951, N6939, N3323, N6100, N6510);
and AND2 (N6952, N6945, N5107);
nor NOR2 (N6953, N6936, N3013);
buf BUF1 (N6954, N6943);
and AND2 (N6955, N6949, N3531);
and AND2 (N6956, N6946, N4613);
nand NAND4 (N6957, N6954, N1565, N6384, N4073);
and AND4 (N6958, N6957, N879, N4952, N2237);
and AND4 (N6959, N6919, N628, N3548, N1407);
or OR4 (N6960, N6955, N2099, N5282, N5671);
buf BUF1 (N6961, N6953);
xor XOR2 (N6962, N6956, N1716);
nor NOR2 (N6963, N6961, N6373);
nand NAND4 (N6964, N6962, N6184, N4603, N4066);
nand NAND2 (N6965, N6958, N3987);
or OR4 (N6966, N6963, N203, N3338, N3875);
xor XOR2 (N6967, N6959, N1026);
not NOT1 (N6968, N6940);
and AND3 (N6969, N6952, N218, N514);
buf BUF1 (N6970, N6967);
buf BUF1 (N6971, N6969);
nor NOR4 (N6972, N6968, N3183, N5338, N1963);
and AND4 (N6973, N6964, N2996, N6839, N6731);
or OR3 (N6974, N6960, N5001, N6015);
nor NOR3 (N6975, N6966, N2890, N495);
or OR3 (N6976, N6972, N3521, N2990);
not NOT1 (N6977, N6974);
not NOT1 (N6978, N6976);
and AND2 (N6979, N6965, N3763);
or OR3 (N6980, N6950, N1581, N5238);
nor NOR3 (N6981, N6951, N4136, N2375);
xor XOR2 (N6982, N6973, N2772);
nand NAND4 (N6983, N6982, N1395, N1821, N3848);
nand NAND4 (N6984, N6978, N2078, N6610, N4060);
nor NOR3 (N6985, N6948, N1924, N6633);
or OR3 (N6986, N6975, N4685, N4660);
buf BUF1 (N6987, N6985);
buf BUF1 (N6988, N6971);
not NOT1 (N6989, N6984);
and AND3 (N6990, N6977, N293, N632);
not NOT1 (N6991, N6983);
or OR2 (N6992, N6989, N2595);
buf BUF1 (N6993, N6980);
and AND3 (N6994, N6990, N4828, N6690);
and AND4 (N6995, N6970, N3777, N3919, N3500);
buf BUF1 (N6996, N6992);
and AND3 (N6997, N6988, N1739, N1868);
nand NAND2 (N6998, N6981, N4055);
nor NOR2 (N6999, N6991, N993);
and AND2 (N7000, N6998, N6876);
nand NAND4 (N7001, N6986, N1982, N2338, N5029);
buf BUF1 (N7002, N6996);
nand NAND3 (N7003, N7000, N3723, N6415);
or OR4 (N7004, N7003, N1664, N3277, N2734);
buf BUF1 (N7005, N6999);
nor NOR4 (N7006, N7002, N919, N938, N2689);
or OR4 (N7007, N6995, N5287, N3563, N3301);
or OR3 (N7008, N7006, N2446, N6883);
or OR2 (N7009, N7007, N5364);
or OR4 (N7010, N7008, N5357, N6741, N1200);
or OR2 (N7011, N6979, N5381);
buf BUF1 (N7012, N7010);
and AND4 (N7013, N7005, N6920, N5309, N2866);
nor NOR4 (N7014, N7012, N4231, N5098, N1320);
not NOT1 (N7015, N6994);
or OR4 (N7016, N7011, N1209, N3232, N6112);
nor NOR2 (N7017, N7013, N948);
nand NAND3 (N7018, N7017, N2638, N6895);
and AND2 (N7019, N6997, N3822);
or OR3 (N7020, N7015, N443, N1145);
buf BUF1 (N7021, N7004);
nor NOR2 (N7022, N7019, N6163);
nor NOR3 (N7023, N7021, N1816, N523);
and AND3 (N7024, N7018, N2467, N1268);
and AND4 (N7025, N7014, N1345, N5013, N6359);
xor XOR2 (N7026, N7020, N919);
or OR2 (N7027, N6987, N2768);
nor NOR3 (N7028, N7025, N6966, N1806);
or OR2 (N7029, N7024, N3481);
nor NOR2 (N7030, N7016, N3489);
nand NAND4 (N7031, N7027, N3551, N6503, N1673);
or OR4 (N7032, N7001, N715, N4029, N6817);
buf BUF1 (N7033, N7028);
buf BUF1 (N7034, N7022);
not NOT1 (N7035, N7023);
not NOT1 (N7036, N7034);
and AND4 (N7037, N7029, N6682, N6441, N2205);
xor XOR2 (N7038, N7035, N6752);
nor NOR4 (N7039, N7009, N3060, N1391, N2547);
buf BUF1 (N7040, N7030);
nand NAND3 (N7041, N6993, N3782, N1325);
buf BUF1 (N7042, N7037);
xor XOR2 (N7043, N7038, N3849);
nand NAND4 (N7044, N7042, N2440, N1404, N5892);
or OR4 (N7045, N7040, N557, N3606, N1327);
not NOT1 (N7046, N7026);
nor NOR2 (N7047, N7032, N3180);
not NOT1 (N7048, N7036);
nand NAND2 (N7049, N7041, N2533);
and AND3 (N7050, N7043, N7028, N5672);
or OR2 (N7051, N7046, N740);
xor XOR2 (N7052, N7033, N5406);
nor NOR4 (N7053, N7047, N3741, N6182, N6787);
not NOT1 (N7054, N7045);
nand NAND3 (N7055, N7031, N1461, N5840);
buf BUF1 (N7056, N7039);
xor XOR2 (N7057, N7053, N4912);
nor NOR3 (N7058, N7051, N1249, N4179);
xor XOR2 (N7059, N7057, N1358);
and AND4 (N7060, N7055, N553, N2508, N5935);
buf BUF1 (N7061, N7060);
nand NAND3 (N7062, N7049, N101, N6393);
nand NAND4 (N7063, N7050, N4742, N5094, N6771);
or OR2 (N7064, N7052, N1372);
nand NAND4 (N7065, N7059, N3326, N1254, N3548);
not NOT1 (N7066, N7061);
not NOT1 (N7067, N7054);
not NOT1 (N7068, N7056);
nand NAND2 (N7069, N7068, N256);
xor XOR2 (N7070, N7069, N2645);
xor XOR2 (N7071, N7058, N7049);
nand NAND2 (N7072, N7065, N2556);
not NOT1 (N7073, N7072);
xor XOR2 (N7074, N7048, N2314);
buf BUF1 (N7075, N7073);
or OR3 (N7076, N7066, N4533, N3904);
not NOT1 (N7077, N7063);
buf BUF1 (N7078, N7077);
and AND3 (N7079, N7076, N5232, N473);
buf BUF1 (N7080, N7071);
nor NOR4 (N7081, N7080, N722, N1148, N6253);
buf BUF1 (N7082, N7070);
not NOT1 (N7083, N7078);
xor XOR2 (N7084, N7081, N807);
xor XOR2 (N7085, N7084, N4350);
not NOT1 (N7086, N7062);
not NOT1 (N7087, N7044);
nand NAND4 (N7088, N7082, N2181, N5606, N5112);
or OR3 (N7089, N7075, N6310, N3029);
nand NAND2 (N7090, N7079, N2756);
nand NAND4 (N7091, N7090, N6677, N4729, N1418);
nand NAND3 (N7092, N7088, N2260, N6270);
not NOT1 (N7093, N7067);
nand NAND2 (N7094, N7086, N6340);
xor XOR2 (N7095, N7074, N3896);
and AND3 (N7096, N7064, N3892, N4717);
xor XOR2 (N7097, N7085, N4975);
xor XOR2 (N7098, N7087, N73);
buf BUF1 (N7099, N7089);
nor NOR3 (N7100, N7098, N6321, N697);
and AND2 (N7101, N7100, N6980);
buf BUF1 (N7102, N7092);
not NOT1 (N7103, N7093);
xor XOR2 (N7104, N7103, N5053);
not NOT1 (N7105, N7101);
not NOT1 (N7106, N7104);
nand NAND3 (N7107, N7091, N2000, N3841);
or OR3 (N7108, N7097, N4228, N4996);
not NOT1 (N7109, N7105);
buf BUF1 (N7110, N7096);
or OR3 (N7111, N7094, N3274, N3564);
not NOT1 (N7112, N7108);
nand NAND4 (N7113, N7109, N386, N435, N2707);
not NOT1 (N7114, N7112);
not NOT1 (N7115, N7083);
not NOT1 (N7116, N7106);
and AND2 (N7117, N7107, N3508);
not NOT1 (N7118, N7102);
nand NAND2 (N7119, N7099, N1220);
and AND3 (N7120, N7115, N1272, N2706);
not NOT1 (N7121, N7116);
xor XOR2 (N7122, N7117, N3724);
xor XOR2 (N7123, N7113, N2820);
nand NAND2 (N7124, N7118, N2263);
xor XOR2 (N7125, N7110, N6548);
not NOT1 (N7126, N7111);
and AND3 (N7127, N7124, N5679, N4739);
or OR3 (N7128, N7114, N155, N4822);
or OR3 (N7129, N7119, N6394, N5661);
nor NOR4 (N7130, N7121, N4542, N1428, N2603);
buf BUF1 (N7131, N7120);
xor XOR2 (N7132, N7129, N4850);
nor NOR2 (N7133, N7123, N6428);
nor NOR3 (N7134, N7126, N662, N3863);
or OR3 (N7135, N7133, N4831, N1085);
nand NAND4 (N7136, N7122, N4261, N6192, N762);
buf BUF1 (N7137, N7127);
xor XOR2 (N7138, N7137, N6633);
and AND4 (N7139, N7138, N58, N3247, N6283);
not NOT1 (N7140, N7139);
xor XOR2 (N7141, N7095, N1723);
nor NOR2 (N7142, N7125, N1438);
xor XOR2 (N7143, N7140, N2559);
not NOT1 (N7144, N7128);
and AND2 (N7145, N7136, N4599);
or OR4 (N7146, N7132, N6360, N3212, N3297);
or OR3 (N7147, N7134, N5499, N3517);
nand NAND3 (N7148, N7146, N6452, N5778);
or OR3 (N7149, N7142, N3759, N1970);
not NOT1 (N7150, N7147);
buf BUF1 (N7151, N7149);
not NOT1 (N7152, N7131);
nor NOR2 (N7153, N7150, N3130);
not NOT1 (N7154, N7144);
nor NOR2 (N7155, N7145, N2395);
nor NOR4 (N7156, N7154, N622, N6380, N2770);
or OR4 (N7157, N7155, N3957, N2253, N3396);
and AND4 (N7158, N7157, N2858, N977, N6883);
and AND2 (N7159, N7141, N1079);
and AND4 (N7160, N7148, N5331, N2120, N2429);
nand NAND3 (N7161, N7152, N4875, N5256);
not NOT1 (N7162, N7143);
xor XOR2 (N7163, N7135, N3185);
and AND2 (N7164, N7160, N3629);
or OR4 (N7165, N7153, N1896, N3128, N4731);
nand NAND2 (N7166, N7163, N2230);
buf BUF1 (N7167, N7159);
and AND3 (N7168, N7158, N1206, N4037);
not NOT1 (N7169, N7162);
or OR3 (N7170, N7166, N5871, N5005);
buf BUF1 (N7171, N7165);
not NOT1 (N7172, N7151);
or OR4 (N7173, N7172, N4956, N2146, N3755);
or OR3 (N7174, N7168, N4856, N707);
nor NOR3 (N7175, N7156, N6153, N3569);
not NOT1 (N7176, N7173);
nand NAND4 (N7177, N7170, N4571, N5837, N2869);
and AND3 (N7178, N7169, N5957, N6804);
xor XOR2 (N7179, N7178, N3573);
nand NAND2 (N7180, N7164, N3567);
and AND2 (N7181, N7177, N6299);
nand NAND3 (N7182, N7174, N2279, N5989);
nor NOR2 (N7183, N7130, N1465);
nor NOR2 (N7184, N7180, N3875);
nor NOR4 (N7185, N7175, N1545, N3813, N146);
not NOT1 (N7186, N7181);
buf BUF1 (N7187, N7171);
not NOT1 (N7188, N7187);
and AND2 (N7189, N7179, N4748);
buf BUF1 (N7190, N7176);
or OR2 (N7191, N7185, N1769);
buf BUF1 (N7192, N7184);
nand NAND4 (N7193, N7189, N748, N5813, N223);
and AND4 (N7194, N7192, N5973, N6594, N7045);
buf BUF1 (N7195, N7188);
not NOT1 (N7196, N7161);
nand NAND3 (N7197, N7182, N5233, N7106);
or OR3 (N7198, N7191, N4425, N1201);
and AND2 (N7199, N7186, N5456);
buf BUF1 (N7200, N7197);
nand NAND4 (N7201, N7190, N6231, N6417, N1413);
nand NAND4 (N7202, N7193, N152, N5261, N6813);
xor XOR2 (N7203, N7199, N3973);
buf BUF1 (N7204, N7195);
xor XOR2 (N7205, N7203, N3789);
or OR2 (N7206, N7205, N5210);
nand NAND2 (N7207, N7194, N7072);
nand NAND4 (N7208, N7201, N1845, N123, N1953);
buf BUF1 (N7209, N7208);
nor NOR2 (N7210, N7167, N5581);
and AND2 (N7211, N7207, N3898);
or OR3 (N7212, N7196, N2615, N1529);
buf BUF1 (N7213, N7204);
xor XOR2 (N7214, N7200, N1659);
not NOT1 (N7215, N7198);
and AND2 (N7216, N7215, N5968);
buf BUF1 (N7217, N7213);
nor NOR2 (N7218, N7214, N5909);
nand NAND2 (N7219, N7183, N2013);
nand NAND3 (N7220, N7218, N3184, N3726);
not NOT1 (N7221, N7209);
nand NAND3 (N7222, N7212, N6197, N4419);
xor XOR2 (N7223, N7202, N4960);
nor NOR3 (N7224, N7221, N4707, N6292);
nand NAND2 (N7225, N7223, N5425);
nand NAND4 (N7226, N7216, N4878, N4065, N123);
xor XOR2 (N7227, N7226, N2699);
nor NOR2 (N7228, N7220, N6076);
not NOT1 (N7229, N7206);
nand NAND2 (N7230, N7225, N5691);
or OR4 (N7231, N7219, N4180, N4117, N6780);
buf BUF1 (N7232, N7217);
not NOT1 (N7233, N7229);
or OR2 (N7234, N7224, N3962);
nand NAND2 (N7235, N7228, N5032);
nor NOR4 (N7236, N7222, N2119, N5518, N4472);
buf BUF1 (N7237, N7236);
nor NOR2 (N7238, N7230, N960);
nor NOR4 (N7239, N7232, N7070, N4159, N1810);
not NOT1 (N7240, N7238);
not NOT1 (N7241, N7211);
buf BUF1 (N7242, N7233);
and AND3 (N7243, N7241, N4808, N3807);
nand NAND4 (N7244, N7237, N3308, N2870, N2122);
and AND2 (N7245, N7227, N6988);
not NOT1 (N7246, N7242);
nor NOR2 (N7247, N7235, N316);
xor XOR2 (N7248, N7239, N4172);
nand NAND2 (N7249, N7231, N4569);
or OR4 (N7250, N7243, N5421, N528, N4340);
nand NAND2 (N7251, N7245, N4572);
not NOT1 (N7252, N7210);
xor XOR2 (N7253, N7250, N6800);
nor NOR2 (N7254, N7247, N3268);
buf BUF1 (N7255, N7251);
buf BUF1 (N7256, N7249);
or OR4 (N7257, N7240, N4597, N5465, N5413);
not NOT1 (N7258, N7256);
xor XOR2 (N7259, N7258, N4928);
nor NOR2 (N7260, N7246, N3723);
buf BUF1 (N7261, N7259);
and AND2 (N7262, N7234, N5065);
nand NAND4 (N7263, N7260, N4685, N4157, N6212);
xor XOR2 (N7264, N7253, N6743);
not NOT1 (N7265, N7248);
nor NOR4 (N7266, N7265, N2982, N4979, N4037);
xor XOR2 (N7267, N7261, N3037);
nand NAND2 (N7268, N7264, N4049);
xor XOR2 (N7269, N7268, N4061);
or OR2 (N7270, N7267, N6097);
buf BUF1 (N7271, N7252);
xor XOR2 (N7272, N7263, N4547);
xor XOR2 (N7273, N7254, N5566);
and AND4 (N7274, N7269, N4724, N1132, N5942);
and AND3 (N7275, N7262, N6694, N6847);
xor XOR2 (N7276, N7244, N4111);
xor XOR2 (N7277, N7275, N570);
buf BUF1 (N7278, N7257);
or OR3 (N7279, N7276, N6114, N3748);
not NOT1 (N7280, N7274);
xor XOR2 (N7281, N7255, N5637);
not NOT1 (N7282, N7281);
not NOT1 (N7283, N7272);
and AND3 (N7284, N7279, N5027, N7204);
or OR2 (N7285, N7284, N5763);
and AND4 (N7286, N7266, N5765, N2891, N3662);
not NOT1 (N7287, N7278);
and AND3 (N7288, N7277, N4991, N2448);
and AND3 (N7289, N7288, N2981, N3641);
and AND4 (N7290, N7283, N1447, N582, N6398);
and AND3 (N7291, N7282, N5953, N1395);
buf BUF1 (N7292, N7290);
xor XOR2 (N7293, N7273, N3932);
not NOT1 (N7294, N7289);
or OR2 (N7295, N7286, N1545);
or OR2 (N7296, N7295, N6363);
xor XOR2 (N7297, N7271, N588);
nor NOR3 (N7298, N7285, N4805, N1414);
nor NOR3 (N7299, N7292, N495, N7008);
nand NAND3 (N7300, N7296, N6613, N4463);
xor XOR2 (N7301, N7270, N2990);
not NOT1 (N7302, N7291);
and AND4 (N7303, N7293, N4821, N4436, N7211);
and AND3 (N7304, N7280, N6021, N4518);
nand NAND3 (N7305, N7297, N2664, N532);
buf BUF1 (N7306, N7301);
nor NOR4 (N7307, N7298, N3521, N1763, N5415);
xor XOR2 (N7308, N7303, N3826);
and AND2 (N7309, N7306, N2348);
buf BUF1 (N7310, N7299);
not NOT1 (N7311, N7302);
buf BUF1 (N7312, N7305);
and AND3 (N7313, N7307, N3139, N877);
buf BUF1 (N7314, N7294);
xor XOR2 (N7315, N7312, N3097);
xor XOR2 (N7316, N7311, N1694);
or OR3 (N7317, N7287, N1210, N1161);
buf BUF1 (N7318, N7315);
xor XOR2 (N7319, N7316, N1028);
nand NAND4 (N7320, N7310, N158, N4472, N2666);
or OR3 (N7321, N7309, N3657, N2321);
not NOT1 (N7322, N7300);
nor NOR4 (N7323, N7319, N258, N3082, N6903);
or OR3 (N7324, N7308, N3614, N1610);
buf BUF1 (N7325, N7324);
buf BUF1 (N7326, N7323);
nand NAND2 (N7327, N7322, N3790);
or OR3 (N7328, N7326, N2519, N3313);
nor NOR3 (N7329, N7325, N4638, N7036);
buf BUF1 (N7330, N7328);
not NOT1 (N7331, N7317);
nand NAND4 (N7332, N7313, N5235, N6285, N164);
nor NOR2 (N7333, N7318, N7239);
xor XOR2 (N7334, N7314, N1394);
buf BUF1 (N7335, N7321);
nand NAND2 (N7336, N7332, N6941);
not NOT1 (N7337, N7304);
not NOT1 (N7338, N7320);
nor NOR4 (N7339, N7336, N3956, N3482, N2694);
buf BUF1 (N7340, N7330);
xor XOR2 (N7341, N7338, N7180);
xor XOR2 (N7342, N7340, N583);
nand NAND2 (N7343, N7342, N6870);
xor XOR2 (N7344, N7329, N4954);
nor NOR2 (N7345, N7334, N4110);
nor NOR4 (N7346, N7343, N5018, N552, N1251);
nor NOR2 (N7347, N7344, N702);
or OR3 (N7348, N7333, N3195, N2950);
nor NOR4 (N7349, N7348, N7066, N6271, N1431);
not NOT1 (N7350, N7349);
nor NOR2 (N7351, N7339, N2678);
and AND2 (N7352, N7327, N3231);
nand NAND3 (N7353, N7352, N1647, N2351);
xor XOR2 (N7354, N7331, N2066);
and AND4 (N7355, N7346, N4331, N4491, N2000);
or OR4 (N7356, N7355, N4619, N6278, N6377);
buf BUF1 (N7357, N7345);
nand NAND3 (N7358, N7341, N3999, N526);
buf BUF1 (N7359, N7354);
or OR4 (N7360, N7337, N6845, N6428, N4601);
or OR3 (N7361, N7356, N2556, N7353);
nor NOR4 (N7362, N154, N3887, N1358, N6045);
and AND3 (N7363, N7361, N5718, N530);
nand NAND2 (N7364, N7335, N7002);
nand NAND4 (N7365, N7362, N1112, N5983, N5635);
and AND4 (N7366, N7350, N614, N3468, N4769);
nor NOR3 (N7367, N7366, N1069, N1028);
or OR4 (N7368, N7365, N4787, N2010, N3792);
not NOT1 (N7369, N7368);
nor NOR4 (N7370, N7367, N6581, N3977, N2800);
and AND2 (N7371, N7359, N4400);
not NOT1 (N7372, N7358);
not NOT1 (N7373, N7351);
and AND2 (N7374, N7371, N3508);
buf BUF1 (N7375, N7363);
xor XOR2 (N7376, N7364, N628);
nand NAND4 (N7377, N7376, N2457, N1819, N6466);
buf BUF1 (N7378, N7372);
and AND4 (N7379, N7347, N6291, N327, N2997);
nand NAND3 (N7380, N7375, N1162, N4659);
and AND2 (N7381, N7379, N1762);
nor NOR2 (N7382, N7369, N424);
and AND3 (N7383, N7377, N1753, N4271);
xor XOR2 (N7384, N7373, N675);
xor XOR2 (N7385, N7384, N103);
buf BUF1 (N7386, N7370);
not NOT1 (N7387, N7357);
nand NAND4 (N7388, N7378, N5932, N2352, N398);
xor XOR2 (N7389, N7374, N6238);
xor XOR2 (N7390, N7385, N579);
and AND3 (N7391, N7390, N2992, N5318);
or OR3 (N7392, N7389, N5182, N1931);
nand NAND2 (N7393, N7380, N7217);
buf BUF1 (N7394, N7387);
or OR2 (N7395, N7383, N1235);
not NOT1 (N7396, N7391);
nor NOR4 (N7397, N7382, N3256, N648, N4418);
and AND3 (N7398, N7392, N34, N700);
xor XOR2 (N7399, N7396, N4209);
buf BUF1 (N7400, N7398);
or OR2 (N7401, N7399, N7281);
nand NAND2 (N7402, N7395, N7368);
or OR2 (N7403, N7393, N5210);
buf BUF1 (N7404, N7388);
or OR2 (N7405, N7386, N6967);
xor XOR2 (N7406, N7400, N2466);
not NOT1 (N7407, N7381);
xor XOR2 (N7408, N7406, N4561);
or OR3 (N7409, N7407, N972, N5169);
xor XOR2 (N7410, N7402, N6778);
xor XOR2 (N7411, N7401, N2067);
xor XOR2 (N7412, N7408, N2657);
nor NOR3 (N7413, N7404, N1623, N1288);
not NOT1 (N7414, N7411);
not NOT1 (N7415, N7405);
or OR4 (N7416, N7414, N5127, N5662, N5069);
nand NAND4 (N7417, N7416, N7021, N2527, N3663);
not NOT1 (N7418, N7394);
nand NAND2 (N7419, N7403, N224);
and AND3 (N7420, N7410, N2465, N2641);
nor NOR2 (N7421, N7360, N5682);
and AND3 (N7422, N7421, N3511, N7267);
nor NOR4 (N7423, N7419, N7079, N1247, N2278);
or OR4 (N7424, N7412, N221, N4906, N968);
or OR3 (N7425, N7417, N5430, N4798);
and AND4 (N7426, N7422, N6626, N1377, N4282);
and AND2 (N7427, N7418, N1922);
buf BUF1 (N7428, N7426);
xor XOR2 (N7429, N7397, N2398);
not NOT1 (N7430, N7428);
nor NOR3 (N7431, N7423, N3238, N662);
buf BUF1 (N7432, N7420);
xor XOR2 (N7433, N7415, N6134);
or OR4 (N7434, N7433, N3426, N2354, N954);
nand NAND3 (N7435, N7431, N7358, N409);
or OR4 (N7436, N7434, N2007, N3277, N4328);
not NOT1 (N7437, N7432);
buf BUF1 (N7438, N7435);
and AND3 (N7439, N7424, N2328, N6036);
or OR3 (N7440, N7429, N1160, N6795);
xor XOR2 (N7441, N7436, N4054);
nand NAND3 (N7442, N7430, N243, N2515);
buf BUF1 (N7443, N7439);
nor NOR4 (N7444, N7437, N4325, N360, N125);
and AND4 (N7445, N7443, N1205, N6761, N636);
and AND3 (N7446, N7444, N5307, N1324);
or OR2 (N7447, N7409, N1104);
buf BUF1 (N7448, N7425);
and AND4 (N7449, N7441, N4886, N1618, N5834);
nand NAND3 (N7450, N7446, N1967, N6258);
nor NOR4 (N7451, N7413, N7236, N2504, N2853);
not NOT1 (N7452, N7440);
not NOT1 (N7453, N7445);
nand NAND2 (N7454, N7453, N6494);
not NOT1 (N7455, N7452);
not NOT1 (N7456, N7427);
xor XOR2 (N7457, N7447, N7370);
xor XOR2 (N7458, N7448, N2365);
not NOT1 (N7459, N7456);
nor NOR2 (N7460, N7458, N4814);
buf BUF1 (N7461, N7450);
nor NOR2 (N7462, N7459, N1726);
nor NOR2 (N7463, N7461, N1045);
not NOT1 (N7464, N7455);
xor XOR2 (N7465, N7462, N1264);
buf BUF1 (N7466, N7464);
nand NAND3 (N7467, N7460, N91, N233);
xor XOR2 (N7468, N7466, N5727);
nand NAND2 (N7469, N7465, N300);
not NOT1 (N7470, N7469);
not NOT1 (N7471, N7463);
xor XOR2 (N7472, N7457, N1216);
or OR3 (N7473, N7451, N7342, N5208);
not NOT1 (N7474, N7467);
xor XOR2 (N7475, N7473, N445);
xor XOR2 (N7476, N7470, N4871);
not NOT1 (N7477, N7472);
nor NOR2 (N7478, N7474, N2391);
xor XOR2 (N7479, N7468, N14);
or OR2 (N7480, N7476, N1049);
nand NAND2 (N7481, N7442, N2101);
or OR4 (N7482, N7438, N576, N5311, N4586);
buf BUF1 (N7483, N7449);
nand NAND3 (N7484, N7471, N3720, N809);
or OR3 (N7485, N7483, N5656, N3632);
buf BUF1 (N7486, N7479);
xor XOR2 (N7487, N7482, N4868);
and AND2 (N7488, N7477, N7464);
or OR4 (N7489, N7488, N6085, N4221, N6202);
nor NOR3 (N7490, N7484, N6857, N2297);
and AND4 (N7491, N7475, N5823, N1813, N1846);
buf BUF1 (N7492, N7487);
and AND2 (N7493, N7480, N5156);
and AND3 (N7494, N7485, N3373, N5257);
nor NOR3 (N7495, N7493, N6221, N5484);
xor XOR2 (N7496, N7490, N2108);
xor XOR2 (N7497, N7496, N2858);
xor XOR2 (N7498, N7495, N2494);
nand NAND4 (N7499, N7478, N6258, N3219, N1655);
or OR3 (N7500, N7497, N4590, N1688);
and AND4 (N7501, N7494, N2773, N6680, N1776);
nand NAND2 (N7502, N7501, N2775);
not NOT1 (N7503, N7491);
nor NOR2 (N7504, N7503, N1284);
nand NAND4 (N7505, N7504, N5306, N6228, N1193);
nand NAND2 (N7506, N7486, N4586);
or OR4 (N7507, N7481, N6324, N6183, N581);
buf BUF1 (N7508, N7502);
nand NAND2 (N7509, N7498, N345);
not NOT1 (N7510, N7507);
buf BUF1 (N7511, N7506);
buf BUF1 (N7512, N7454);
not NOT1 (N7513, N7509);
and AND2 (N7514, N7499, N1802);
nand NAND3 (N7515, N7510, N1670, N4566);
xor XOR2 (N7516, N7512, N5911);
not NOT1 (N7517, N7508);
nand NAND3 (N7518, N7515, N5333, N3145);
nor NOR4 (N7519, N7511, N4507, N4085, N4541);
nor NOR3 (N7520, N7517, N5131, N69);
and AND3 (N7521, N7500, N3530, N5915);
xor XOR2 (N7522, N7518, N1744);
nor NOR3 (N7523, N7513, N6092, N6751);
or OR4 (N7524, N7521, N6968, N1334, N1039);
not NOT1 (N7525, N7523);
nor NOR2 (N7526, N7524, N3276);
and AND3 (N7527, N7492, N5655, N7153);
nor NOR2 (N7528, N7516, N5201);
buf BUF1 (N7529, N7489);
xor XOR2 (N7530, N7526, N414);
or OR4 (N7531, N7522, N3410, N2561, N3413);
nor NOR3 (N7532, N7525, N2602, N1401);
xor XOR2 (N7533, N7514, N1313);
buf BUF1 (N7534, N7529);
not NOT1 (N7535, N7531);
not NOT1 (N7536, N7505);
or OR4 (N7537, N7533, N2777, N3892, N4446);
not NOT1 (N7538, N7532);
and AND3 (N7539, N7519, N4284, N6439);
buf BUF1 (N7540, N7536);
xor XOR2 (N7541, N7538, N4942);
nand NAND4 (N7542, N7537, N829, N6577, N5801);
nor NOR3 (N7543, N7520, N4990, N4682);
not NOT1 (N7544, N7534);
and AND3 (N7545, N7540, N7028, N826);
buf BUF1 (N7546, N7528);
or OR4 (N7547, N7542, N7468, N2321, N433);
nand NAND3 (N7548, N7544, N6782, N7231);
or OR3 (N7549, N7539, N1280, N7095);
xor XOR2 (N7550, N7546, N2653);
or OR2 (N7551, N7527, N5651);
or OR3 (N7552, N7549, N7452, N5886);
nor NOR2 (N7553, N7535, N272);
xor XOR2 (N7554, N7543, N3795);
nand NAND3 (N7555, N7530, N3282, N3574);
not NOT1 (N7556, N7541);
nor NOR2 (N7557, N7553, N2607);
nor NOR3 (N7558, N7555, N1714, N45);
or OR4 (N7559, N7558, N3275, N1310, N5496);
not NOT1 (N7560, N7548);
and AND3 (N7561, N7550, N1050, N7156);
nand NAND2 (N7562, N7556, N3165);
xor XOR2 (N7563, N7557, N5806);
or OR2 (N7564, N7563, N6006);
nor NOR3 (N7565, N7554, N2091, N114);
and AND4 (N7566, N7559, N7558, N4905, N562);
buf BUF1 (N7567, N7545);
nor NOR4 (N7568, N7566, N112, N4475, N3436);
buf BUF1 (N7569, N7562);
buf BUF1 (N7570, N7551);
or OR2 (N7571, N7547, N3787);
and AND4 (N7572, N7569, N4718, N1188, N3996);
or OR2 (N7573, N7571, N3260);
or OR2 (N7574, N7570, N6299);
nor NOR3 (N7575, N7552, N4127, N5572);
not NOT1 (N7576, N7561);
buf BUF1 (N7577, N7567);
buf BUF1 (N7578, N7565);
buf BUF1 (N7579, N7578);
or OR3 (N7580, N7579, N3337, N5241);
or OR4 (N7581, N7577, N4302, N4182, N6427);
xor XOR2 (N7582, N7573, N7136);
nor NOR4 (N7583, N7564, N7177, N2181, N1842);
nand NAND4 (N7584, N7560, N1801, N3194, N657);
and AND2 (N7585, N7568, N2522);
buf BUF1 (N7586, N7585);
not NOT1 (N7587, N7575);
nand NAND3 (N7588, N7581, N5879, N6924);
not NOT1 (N7589, N7576);
not NOT1 (N7590, N7588);
nor NOR4 (N7591, N7572, N5853, N2424, N2585);
buf BUF1 (N7592, N7589);
not NOT1 (N7593, N7580);
nand NAND3 (N7594, N7584, N2735, N6230);
nand NAND4 (N7595, N7574, N3129, N2468, N4498);
buf BUF1 (N7596, N7592);
nand NAND2 (N7597, N7583, N6315);
buf BUF1 (N7598, N7582);
or OR3 (N7599, N7595, N2742, N6183);
or OR3 (N7600, N7591, N4040, N6049);
and AND2 (N7601, N7586, N5451);
nand NAND2 (N7602, N7594, N1996);
not NOT1 (N7603, N7597);
nand NAND2 (N7604, N7587, N5624);
nor NOR2 (N7605, N7596, N5833);
buf BUF1 (N7606, N7599);
buf BUF1 (N7607, N7602);
or OR3 (N7608, N7605, N86, N6460);
nand NAND2 (N7609, N7604, N5785);
or OR4 (N7610, N7598, N4397, N5108, N3431);
buf BUF1 (N7611, N7609);
not NOT1 (N7612, N7593);
not NOT1 (N7613, N7590);
xor XOR2 (N7614, N7607, N5537);
nand NAND2 (N7615, N7612, N5606);
xor XOR2 (N7616, N7600, N479);
not NOT1 (N7617, N7608);
nand NAND4 (N7618, N7610, N3396, N6592, N7006);
and AND3 (N7619, N7616, N5408, N2404);
or OR3 (N7620, N7613, N2119, N5434);
or OR2 (N7621, N7614, N6895);
xor XOR2 (N7622, N7621, N7288);
and AND3 (N7623, N7617, N5529, N4152);
nor NOR3 (N7624, N7603, N5993, N2774);
xor XOR2 (N7625, N7606, N71);
and AND3 (N7626, N7618, N7551, N5987);
nand NAND4 (N7627, N7601, N4004, N3078, N599);
nand NAND4 (N7628, N7615, N3881, N5682, N7342);
xor XOR2 (N7629, N7619, N4960);
nor NOR2 (N7630, N7626, N5085);
or OR2 (N7631, N7628, N2040);
not NOT1 (N7632, N7611);
buf BUF1 (N7633, N7629);
nor NOR2 (N7634, N7630, N3755);
nand NAND2 (N7635, N7624, N3302);
nand NAND4 (N7636, N7632, N765, N7418, N4093);
buf BUF1 (N7637, N7635);
or OR4 (N7638, N7634, N83, N5198, N1546);
not NOT1 (N7639, N7627);
not NOT1 (N7640, N7636);
xor XOR2 (N7641, N7637, N5671);
xor XOR2 (N7642, N7622, N2824);
nand NAND2 (N7643, N7641, N6534);
buf BUF1 (N7644, N7642);
or OR4 (N7645, N7623, N4222, N5207, N2657);
buf BUF1 (N7646, N7625);
or OR3 (N7647, N7646, N5809, N2655);
nand NAND4 (N7648, N7645, N1420, N5348, N44);
or OR3 (N7649, N7647, N6706, N1763);
nor NOR2 (N7650, N7649, N5942);
buf BUF1 (N7651, N7644);
xor XOR2 (N7652, N7648, N2206);
nand NAND2 (N7653, N7638, N4245);
xor XOR2 (N7654, N7631, N7397);
nor NOR3 (N7655, N7640, N3895, N6498);
xor XOR2 (N7656, N7650, N1732);
xor XOR2 (N7657, N7653, N6234);
xor XOR2 (N7658, N7657, N4826);
nor NOR4 (N7659, N7639, N4253, N5394, N6089);
buf BUF1 (N7660, N7633);
xor XOR2 (N7661, N7659, N291);
or OR2 (N7662, N7658, N5458);
buf BUF1 (N7663, N7620);
nand NAND3 (N7664, N7655, N5009, N6327);
nor NOR2 (N7665, N7660, N314);
or OR3 (N7666, N7662, N3791, N4665);
not NOT1 (N7667, N7651);
and AND3 (N7668, N7663, N4158, N3613);
nand NAND4 (N7669, N7666, N6885, N724, N1396);
nor NOR3 (N7670, N7665, N2782, N5460);
and AND3 (N7671, N7661, N1188, N3718);
and AND2 (N7672, N7656, N2116);
not NOT1 (N7673, N7643);
nand NAND2 (N7674, N7668, N5865);
not NOT1 (N7675, N7669);
and AND2 (N7676, N7654, N3023);
nor NOR4 (N7677, N7670, N6312, N6787, N2740);
or OR4 (N7678, N7671, N2339, N7623, N2602);
nor NOR3 (N7679, N7678, N5819, N6009);
not NOT1 (N7680, N7676);
or OR4 (N7681, N7674, N5341, N4178, N1690);
buf BUF1 (N7682, N7652);
nand NAND3 (N7683, N7664, N6299, N5566);
xor XOR2 (N7684, N7667, N771);
not NOT1 (N7685, N7681);
xor XOR2 (N7686, N7682, N5769);
or OR3 (N7687, N7683, N962, N7625);
nor NOR3 (N7688, N7686, N395, N265);
buf BUF1 (N7689, N7684);
nand NAND4 (N7690, N7679, N4210, N3745, N6784);
and AND2 (N7691, N7687, N1493);
nand NAND4 (N7692, N7677, N1725, N2571, N4193);
and AND3 (N7693, N7685, N1696, N836);
nand NAND2 (N7694, N7689, N4216);
xor XOR2 (N7695, N7672, N3170);
or OR2 (N7696, N7694, N2096);
xor XOR2 (N7697, N7688, N522);
not NOT1 (N7698, N7695);
and AND4 (N7699, N7675, N2721, N4916, N7533);
or OR2 (N7700, N7696, N69);
nand NAND2 (N7701, N7699, N5901);
buf BUF1 (N7702, N7673);
not NOT1 (N7703, N7691);
buf BUF1 (N7704, N7692);
nor NOR3 (N7705, N7697, N634, N3337);
nor NOR3 (N7706, N7704, N6154, N372);
nand NAND2 (N7707, N7690, N5578);
and AND3 (N7708, N7706, N6557, N5294);
nor NOR3 (N7709, N7705, N5960, N4456);
buf BUF1 (N7710, N7693);
buf BUF1 (N7711, N7707);
and AND4 (N7712, N7701, N2112, N6956, N859);
nand NAND3 (N7713, N7710, N5253, N6469);
nand NAND2 (N7714, N7708, N5257);
or OR3 (N7715, N7709, N7029, N451);
buf BUF1 (N7716, N7703);
xor XOR2 (N7717, N7714, N2815);
or OR3 (N7718, N7711, N7602, N1452);
nor NOR3 (N7719, N7716, N67, N3701);
or OR2 (N7720, N7702, N3147);
buf BUF1 (N7721, N7718);
nand NAND3 (N7722, N7713, N1315, N525);
not NOT1 (N7723, N7717);
xor XOR2 (N7724, N7723, N892);
not NOT1 (N7725, N7719);
xor XOR2 (N7726, N7725, N3388);
not NOT1 (N7727, N7700);
buf BUF1 (N7728, N7722);
buf BUF1 (N7729, N7727);
nor NOR3 (N7730, N7712, N6588, N1235);
or OR4 (N7731, N7720, N2264, N4444, N1436);
and AND4 (N7732, N7698, N1570, N1247, N241);
nor NOR2 (N7733, N7729, N1218);
and AND4 (N7734, N7724, N2518, N2438, N2486);
not NOT1 (N7735, N7726);
buf BUF1 (N7736, N7735);
xor XOR2 (N7737, N7734, N2659);
xor XOR2 (N7738, N7731, N7700);
not NOT1 (N7739, N7738);
xor XOR2 (N7740, N7733, N299);
or OR4 (N7741, N7732, N3513, N7218, N6265);
or OR2 (N7742, N7730, N3989);
nor NOR4 (N7743, N7742, N6886, N6118, N3665);
nor NOR4 (N7744, N7680, N7162, N5428, N6715);
not NOT1 (N7745, N7740);
and AND3 (N7746, N7737, N5476, N2589);
or OR4 (N7747, N7739, N709, N1612, N2618);
nor NOR4 (N7748, N7728, N4178, N1605, N4462);
buf BUF1 (N7749, N7715);
nand NAND4 (N7750, N7747, N7360, N4976, N5293);
not NOT1 (N7751, N7743);
nand NAND4 (N7752, N7746, N1995, N4714, N6360);
not NOT1 (N7753, N7749);
nor NOR3 (N7754, N7752, N4110, N907);
and AND4 (N7755, N7753, N556, N636, N6790);
nand NAND2 (N7756, N7741, N686);
nand NAND2 (N7757, N7754, N42);
nor NOR2 (N7758, N7748, N2710);
nand NAND3 (N7759, N7755, N5551, N942);
not NOT1 (N7760, N7757);
or OR4 (N7761, N7760, N2060, N1185, N5776);
not NOT1 (N7762, N7745);
or OR2 (N7763, N7736, N594);
nand NAND2 (N7764, N7762, N3519);
nor NOR3 (N7765, N7744, N7348, N7105);
nand NAND2 (N7766, N7764, N7575);
and AND2 (N7767, N7758, N5968);
or OR4 (N7768, N7751, N6357, N778, N2378);
xor XOR2 (N7769, N7759, N6987);
and AND3 (N7770, N7768, N4745, N374);
xor XOR2 (N7771, N7756, N4836);
not NOT1 (N7772, N7771);
xor XOR2 (N7773, N7767, N4909);
buf BUF1 (N7774, N7770);
not NOT1 (N7775, N7774);
and AND2 (N7776, N7765, N1660);
nand NAND3 (N7777, N7773, N729, N1607);
nor NOR2 (N7778, N7721, N5366);
or OR2 (N7779, N7778, N2256);
nand NAND4 (N7780, N7766, N6877, N3343, N6088);
buf BUF1 (N7781, N7750);
xor XOR2 (N7782, N7763, N2833);
nor NOR3 (N7783, N7780, N6684, N1499);
nand NAND4 (N7784, N7761, N4147, N1758, N2457);
nor NOR3 (N7785, N7783, N2673, N1451);
not NOT1 (N7786, N7776);
not NOT1 (N7787, N7781);
and AND2 (N7788, N7785, N2405);
nor NOR2 (N7789, N7777, N5360);
and AND2 (N7790, N7784, N2041);
and AND3 (N7791, N7782, N4419, N1927);
nor NOR3 (N7792, N7791, N165, N6410);
buf BUF1 (N7793, N7775);
not NOT1 (N7794, N7779);
or OR4 (N7795, N7769, N5578, N5695, N3249);
nand NAND3 (N7796, N7794, N748, N6820);
nor NOR4 (N7797, N7789, N5975, N5736, N1741);
nand NAND2 (N7798, N7788, N6831);
not NOT1 (N7799, N7796);
and AND3 (N7800, N7798, N2493, N5078);
not NOT1 (N7801, N7793);
not NOT1 (N7802, N7772);
or OR2 (N7803, N7797, N4560);
nor NOR2 (N7804, N7799, N5660);
nor NOR2 (N7805, N7790, N2099);
or OR4 (N7806, N7802, N4877, N3530, N4791);
or OR3 (N7807, N7800, N5137, N2833);
nor NOR3 (N7808, N7803, N1703, N5210);
and AND3 (N7809, N7804, N1903, N7401);
xor XOR2 (N7810, N7795, N5725);
nand NAND4 (N7811, N7808, N887, N582, N4074);
xor XOR2 (N7812, N7792, N5025);
not NOT1 (N7813, N7807);
and AND2 (N7814, N7786, N6157);
or OR4 (N7815, N7810, N4392, N7364, N7625);
nand NAND3 (N7816, N7806, N1477, N1603);
xor XOR2 (N7817, N7805, N3485);
xor XOR2 (N7818, N7816, N1975);
or OR4 (N7819, N7814, N2364, N7817, N7279);
buf BUF1 (N7820, N4056);
nor NOR3 (N7821, N7812, N3060, N7265);
or OR2 (N7822, N7811, N4871);
xor XOR2 (N7823, N7787, N5426);
buf BUF1 (N7824, N7820);
xor XOR2 (N7825, N7819, N170);
not NOT1 (N7826, N7824);
xor XOR2 (N7827, N7801, N3878);
and AND3 (N7828, N7821, N3567, N4480);
buf BUF1 (N7829, N7818);
nand NAND2 (N7830, N7823, N920);
buf BUF1 (N7831, N7815);
not NOT1 (N7832, N7826);
nand NAND3 (N7833, N7829, N3974, N3997);
buf BUF1 (N7834, N7825);
xor XOR2 (N7835, N7832, N5697);
not NOT1 (N7836, N7835);
or OR3 (N7837, N7834, N2057, N3375);
and AND2 (N7838, N7833, N5284);
buf BUF1 (N7839, N7837);
nand NAND4 (N7840, N7822, N4079, N2915, N6940);
nor NOR2 (N7841, N7831, N2542);
not NOT1 (N7842, N7840);
and AND3 (N7843, N7841, N4367, N3404);
not NOT1 (N7844, N7813);
nand NAND3 (N7845, N7809, N5995, N6281);
buf BUF1 (N7846, N7838);
xor XOR2 (N7847, N7845, N1134);
nor NOR3 (N7848, N7843, N5411, N7779);
nand NAND3 (N7849, N7847, N7013, N2353);
not NOT1 (N7850, N7844);
buf BUF1 (N7851, N7830);
nand NAND2 (N7852, N7842, N5539);
buf BUF1 (N7853, N7851);
xor XOR2 (N7854, N7846, N7564);
nor NOR3 (N7855, N7849, N796, N4044);
or OR4 (N7856, N7836, N3928, N4096, N3185);
nand NAND3 (N7857, N7827, N3118, N4654);
nor NOR2 (N7858, N7855, N684);
not NOT1 (N7859, N7858);
nor NOR3 (N7860, N7848, N6680, N2808);
not NOT1 (N7861, N7859);
not NOT1 (N7862, N7854);
nand NAND2 (N7863, N7853, N2987);
buf BUF1 (N7864, N7828);
nor NOR4 (N7865, N7852, N7454, N5250, N1727);
nor NOR3 (N7866, N7860, N6686, N7028);
buf BUF1 (N7867, N7857);
nand NAND2 (N7868, N7865, N5154);
nand NAND3 (N7869, N7864, N3835, N1511);
not NOT1 (N7870, N7839);
not NOT1 (N7871, N7863);
xor XOR2 (N7872, N7869, N2186);
nand NAND2 (N7873, N7868, N7169);
or OR2 (N7874, N7873, N1297);
nor NOR4 (N7875, N7850, N6463, N3589, N706);
nor NOR3 (N7876, N7861, N4533, N4947);
or OR2 (N7877, N7856, N6530);
nor NOR3 (N7878, N7870, N6973, N3255);
nor NOR4 (N7879, N7871, N3896, N6453, N3938);
not NOT1 (N7880, N7862);
not NOT1 (N7881, N7878);
nand NAND3 (N7882, N7877, N6543, N6034);
buf BUF1 (N7883, N7882);
not NOT1 (N7884, N7879);
and AND3 (N7885, N7880, N5749, N2153);
and AND3 (N7886, N7875, N6533, N6478);
buf BUF1 (N7887, N7886);
and AND3 (N7888, N7884, N6171, N2938);
xor XOR2 (N7889, N7887, N2194);
and AND3 (N7890, N7883, N366, N2566);
not NOT1 (N7891, N7889);
buf BUF1 (N7892, N7874);
and AND3 (N7893, N7872, N6333, N4163);
not NOT1 (N7894, N7888);
and AND3 (N7895, N7885, N129, N3508);
and AND2 (N7896, N7894, N2688);
nand NAND3 (N7897, N7895, N4518, N2066);
buf BUF1 (N7898, N7876);
nand NAND4 (N7899, N7893, N1986, N6105, N585);
xor XOR2 (N7900, N7899, N5823);
buf BUF1 (N7901, N7896);
not NOT1 (N7902, N7892);
not NOT1 (N7903, N7891);
and AND3 (N7904, N7890, N7296, N1656);
xor XOR2 (N7905, N7867, N7746);
nand NAND3 (N7906, N7881, N3403, N7221);
and AND2 (N7907, N7866, N259);
nand NAND2 (N7908, N7906, N579);
xor XOR2 (N7909, N7898, N3377);
nand NAND3 (N7910, N7909, N4618, N3556);
or OR2 (N7911, N7902, N2129);
xor XOR2 (N7912, N7905, N7884);
buf BUF1 (N7913, N7900);
not NOT1 (N7914, N7911);
nand NAND4 (N7915, N7913, N6054, N116, N7460);
buf BUF1 (N7916, N7907);
not NOT1 (N7917, N7903);
nor NOR2 (N7918, N7914, N2665);
xor XOR2 (N7919, N7904, N1081);
buf BUF1 (N7920, N7918);
not NOT1 (N7921, N7912);
nor NOR3 (N7922, N7910, N6008, N5951);
or OR2 (N7923, N7916, N2020);
and AND2 (N7924, N7908, N2811);
or OR3 (N7925, N7919, N4081, N536);
nor NOR3 (N7926, N7923, N3194, N1462);
not NOT1 (N7927, N7920);
xor XOR2 (N7928, N7924, N5603);
buf BUF1 (N7929, N7915);
and AND4 (N7930, N7927, N2223, N1074, N2324);
and AND2 (N7931, N7925, N202);
and AND3 (N7932, N7929, N7931, N7493);
buf BUF1 (N7933, N7686);
xor XOR2 (N7934, N7917, N5781);
buf BUF1 (N7935, N7932);
nand NAND3 (N7936, N7933, N4494, N2893);
or OR2 (N7937, N7934, N3376);
buf BUF1 (N7938, N7928);
and AND3 (N7939, N7901, N3122, N5307);
or OR4 (N7940, N7922, N4747, N1091, N3344);
buf BUF1 (N7941, N7935);
buf BUF1 (N7942, N7926);
nand NAND4 (N7943, N7937, N6627, N7216, N7688);
nor NOR4 (N7944, N7930, N7901, N1620, N2603);
not NOT1 (N7945, N7939);
xor XOR2 (N7946, N7945, N1639);
nor NOR2 (N7947, N7944, N6832);
or OR2 (N7948, N7921, N3391);
and AND2 (N7949, N7943, N3741);
xor XOR2 (N7950, N7948, N7033);
xor XOR2 (N7951, N7942, N2675);
buf BUF1 (N7952, N7946);
xor XOR2 (N7953, N7949, N3742);
and AND2 (N7954, N7947, N387);
buf BUF1 (N7955, N7941);
or OR3 (N7956, N7940, N7501, N7493);
or OR3 (N7957, N7938, N6813, N2507);
and AND3 (N7958, N7953, N1773, N2372);
xor XOR2 (N7959, N7958, N1820);
and AND2 (N7960, N7955, N1596);
nand NAND2 (N7961, N7897, N3526);
not NOT1 (N7962, N7936);
nand NAND4 (N7963, N7959, N3443, N5578, N1550);
xor XOR2 (N7964, N7951, N3245);
not NOT1 (N7965, N7954);
xor XOR2 (N7966, N7965, N4428);
or OR4 (N7967, N7963, N7330, N1457, N5699);
xor XOR2 (N7968, N7952, N5937);
not NOT1 (N7969, N7961);
nand NAND2 (N7970, N7950, N7092);
and AND3 (N7971, N7964, N5794, N3600);
xor XOR2 (N7972, N7969, N3862);
not NOT1 (N7973, N7966);
nor NOR2 (N7974, N7972, N317);
buf BUF1 (N7975, N7967);
nand NAND2 (N7976, N7957, N2150);
or OR2 (N7977, N7962, N624);
nor NOR2 (N7978, N7975, N819);
xor XOR2 (N7979, N7973, N18);
nand NAND3 (N7980, N7979, N1614, N5612);
and AND4 (N7981, N7970, N4438, N5415, N1995);
nand NAND2 (N7982, N7978, N2735);
nor NOR3 (N7983, N7982, N3606, N2922);
and AND3 (N7984, N7983, N1988, N7177);
or OR3 (N7985, N7984, N4906, N1819);
not NOT1 (N7986, N7977);
nor NOR4 (N7987, N7985, N1878, N2255, N2470);
xor XOR2 (N7988, N7976, N5137);
or OR3 (N7989, N7986, N1958, N500);
not NOT1 (N7990, N7956);
and AND4 (N7991, N7990, N7723, N2087, N1213);
or OR3 (N7992, N7989, N3484, N4539);
not NOT1 (N7993, N7971);
buf BUF1 (N7994, N7987);
xor XOR2 (N7995, N7991, N2422);
nand NAND4 (N7996, N7974, N1761, N3930, N1044);
and AND4 (N7997, N7992, N4329, N7792, N3714);
not NOT1 (N7998, N7995);
buf BUF1 (N7999, N7980);
and AND2 (N8000, N7996, N7892);
nand NAND3 (N8001, N7981, N3041, N896);
nor NOR3 (N8002, N7960, N5144, N7785);
and AND2 (N8003, N7997, N7184);
nand NAND4 (N8004, N8003, N1391, N981, N5428);
and AND2 (N8005, N7998, N5511);
buf BUF1 (N8006, N7993);
and AND3 (N8007, N8000, N662, N3986);
not NOT1 (N8008, N8002);
nor NOR4 (N8009, N8005, N1681, N6857, N1278);
nand NAND4 (N8010, N7994, N6556, N5747, N3060);
nand NAND3 (N8011, N7968, N1526, N116);
buf BUF1 (N8012, N8010);
nand NAND2 (N8013, N8006, N7842);
buf BUF1 (N8014, N8011);
or OR4 (N8015, N8013, N3235, N111, N2716);
buf BUF1 (N8016, N8009);
not NOT1 (N8017, N8014);
buf BUF1 (N8018, N8016);
nor NOR2 (N8019, N8008, N922);
xor XOR2 (N8020, N8015, N6957);
nor NOR3 (N8021, N8001, N1584, N4901);
or OR3 (N8022, N8012, N4971, N3321);
buf BUF1 (N8023, N7999);
xor XOR2 (N8024, N8019, N1472);
nor NOR3 (N8025, N8020, N6138, N5754);
xor XOR2 (N8026, N8024, N7802);
and AND3 (N8027, N8007, N4886, N1790);
and AND2 (N8028, N8004, N868);
or OR4 (N8029, N8021, N6278, N4769, N5121);
or OR3 (N8030, N8029, N3718, N2458);
xor XOR2 (N8031, N8027, N4193);
not NOT1 (N8032, N8031);
buf BUF1 (N8033, N8017);
nor NOR3 (N8034, N8033, N4431, N4354);
xor XOR2 (N8035, N7988, N7795);
buf BUF1 (N8036, N8018);
nand NAND2 (N8037, N8026, N7643);
or OR4 (N8038, N8032, N1728, N301, N584);
nand NAND4 (N8039, N8034, N6485, N3712, N5169);
xor XOR2 (N8040, N8025, N954);
xor XOR2 (N8041, N8035, N3748);
and AND4 (N8042, N8041, N6967, N35, N7927);
nor NOR2 (N8043, N8023, N6965);
buf BUF1 (N8044, N8028);
nor NOR2 (N8045, N8039, N4161);
and AND2 (N8046, N8037, N6857);
xor XOR2 (N8047, N8045, N4608);
buf BUF1 (N8048, N8030);
nand NAND3 (N8049, N8048, N2804, N6888);
nor NOR4 (N8050, N8046, N5074, N6667, N590);
or OR2 (N8051, N8038, N3932);
nand NAND2 (N8052, N8049, N2219);
nor NOR4 (N8053, N8042, N6765, N1215, N3484);
buf BUF1 (N8054, N8040);
xor XOR2 (N8055, N8044, N7690);
or OR3 (N8056, N8022, N4084, N7743);
and AND3 (N8057, N8036, N5271, N104);
buf BUF1 (N8058, N8050);
buf BUF1 (N8059, N8057);
and AND3 (N8060, N8043, N6261, N2401);
not NOT1 (N8061, N8053);
nand NAND4 (N8062, N8051, N1204, N6904, N7331);
not NOT1 (N8063, N8060);
nand NAND2 (N8064, N8052, N6719);
nand NAND3 (N8065, N8058, N6399, N5341);
and AND4 (N8066, N8065, N3826, N6645, N6575);
xor XOR2 (N8067, N8059, N6774);
and AND2 (N8068, N8061, N2152);
xor XOR2 (N8069, N8067, N6064);
nor NOR2 (N8070, N8047, N3268);
xor XOR2 (N8071, N8055, N3616);
or OR2 (N8072, N8068, N5308);
xor XOR2 (N8073, N8070, N6828);
or OR2 (N8074, N8064, N478);
nor NOR4 (N8075, N8073, N4260, N615, N2346);
or OR3 (N8076, N8062, N3661, N5619);
and AND3 (N8077, N8075, N800, N7260);
and AND3 (N8078, N8071, N3103, N2560);
or OR3 (N8079, N8076, N6484, N3360);
xor XOR2 (N8080, N8072, N759);
not NOT1 (N8081, N8063);
not NOT1 (N8082, N8077);
nand NAND2 (N8083, N8078, N5075);
not NOT1 (N8084, N8069);
not NOT1 (N8085, N8074);
and AND2 (N8086, N8054, N6111);
buf BUF1 (N8087, N8085);
and AND2 (N8088, N8082, N6154);
and AND4 (N8089, N8084, N2253, N6845, N145);
nor NOR4 (N8090, N8079, N1970, N3804, N1004);
or OR4 (N8091, N8088, N54, N4629, N7306);
and AND4 (N8092, N8066, N5468, N1989, N5653);
nor NOR2 (N8093, N8086, N3597);
nor NOR2 (N8094, N8083, N5789);
xor XOR2 (N8095, N8089, N888);
xor XOR2 (N8096, N8087, N4891);
xor XOR2 (N8097, N8092, N6952);
buf BUF1 (N8098, N8080);
or OR2 (N8099, N8090, N7674);
or OR4 (N8100, N8056, N1811, N2967, N4152);
xor XOR2 (N8101, N8100, N7401);
nand NAND4 (N8102, N8098, N6209, N6563, N2128);
buf BUF1 (N8103, N8101);
buf BUF1 (N8104, N8097);
or OR4 (N8105, N8081, N8042, N5250, N2244);
and AND3 (N8106, N8091, N3561, N5909);
xor XOR2 (N8107, N8104, N6337);
or OR2 (N8108, N8095, N2735);
and AND4 (N8109, N8093, N5140, N8037, N4740);
or OR3 (N8110, N8096, N1519, N6396);
or OR2 (N8111, N8110, N1110);
nand NAND3 (N8112, N8109, N6628, N174);
or OR3 (N8113, N8106, N461, N6605);
nor NOR2 (N8114, N8099, N972);
buf BUF1 (N8115, N8103);
not NOT1 (N8116, N8105);
buf BUF1 (N8117, N8113);
not NOT1 (N8118, N8094);
and AND4 (N8119, N8118, N6756, N7062, N7839);
buf BUF1 (N8120, N8117);
not NOT1 (N8121, N8102);
buf BUF1 (N8122, N8112);
xor XOR2 (N8123, N8120, N4898);
xor XOR2 (N8124, N8119, N4249);
or OR2 (N8125, N8114, N3362);
or OR2 (N8126, N8115, N5360);
nand NAND4 (N8127, N8126, N5720, N3205, N801);
and AND4 (N8128, N8108, N2096, N2828, N6002);
not NOT1 (N8129, N8124);
or OR3 (N8130, N8127, N5806, N3744);
nand NAND2 (N8131, N8111, N4207);
and AND2 (N8132, N8130, N4384);
nor NOR4 (N8133, N8128, N3660, N6746, N4290);
buf BUF1 (N8134, N8131);
nor NOR2 (N8135, N8132, N7293);
nand NAND4 (N8136, N8125, N2989, N1560, N5100);
not NOT1 (N8137, N8129);
xor XOR2 (N8138, N8116, N4671);
and AND3 (N8139, N8123, N5489, N6757);
nand NAND2 (N8140, N8136, N479);
or OR2 (N8141, N8107, N3023);
buf BUF1 (N8142, N8121);
buf BUF1 (N8143, N8139);
nor NOR2 (N8144, N8133, N6813);
nand NAND2 (N8145, N8134, N3180);
xor XOR2 (N8146, N8140, N321);
xor XOR2 (N8147, N8143, N7556);
or OR3 (N8148, N8135, N6376, N6261);
nand NAND2 (N8149, N8142, N7445);
nor NOR3 (N8150, N8138, N5879, N3347);
not NOT1 (N8151, N8137);
or OR3 (N8152, N8144, N248, N1855);
not NOT1 (N8153, N8151);
nor NOR2 (N8154, N8141, N7389);
or OR2 (N8155, N8147, N3074);
nor NOR3 (N8156, N8150, N7761, N4651);
and AND2 (N8157, N8122, N6075);
xor XOR2 (N8158, N8152, N6236);
nor NOR3 (N8159, N8145, N2192, N443);
nand NAND4 (N8160, N8158, N3887, N5163, N967);
and AND4 (N8161, N8148, N772, N7479, N1526);
not NOT1 (N8162, N8154);
buf BUF1 (N8163, N8159);
xor XOR2 (N8164, N8149, N1240);
xor XOR2 (N8165, N8163, N4540);
xor XOR2 (N8166, N8164, N2818);
or OR2 (N8167, N8162, N6996);
nor NOR4 (N8168, N8160, N4187, N1503, N6816);
nand NAND3 (N8169, N8168, N6204, N4165);
xor XOR2 (N8170, N8155, N408);
and AND4 (N8171, N8156, N4490, N2197, N4838);
and AND2 (N8172, N8171, N6899);
xor XOR2 (N8173, N8167, N8141);
and AND4 (N8174, N8173, N1344, N7274, N3836);
nor NOR2 (N8175, N8172, N6075);
buf BUF1 (N8176, N8174);
nor NOR2 (N8177, N8169, N2086);
and AND4 (N8178, N8146, N7102, N1075, N4887);
and AND3 (N8179, N8175, N4559, N3621);
not NOT1 (N8180, N8170);
xor XOR2 (N8181, N8177, N2649);
nand NAND4 (N8182, N8161, N3848, N4557, N2385);
buf BUF1 (N8183, N8181);
nand NAND2 (N8184, N8176, N186);
xor XOR2 (N8185, N8153, N6431);
not NOT1 (N8186, N8157);
nor NOR4 (N8187, N8178, N3746, N5613, N5428);
xor XOR2 (N8188, N8183, N3808);
xor XOR2 (N8189, N8165, N2533);
and AND3 (N8190, N8182, N4210, N4806);
buf BUF1 (N8191, N8189);
xor XOR2 (N8192, N8179, N5287);
not NOT1 (N8193, N8186);
and AND4 (N8194, N8166, N6480, N6105, N2772);
and AND2 (N8195, N8188, N993);
and AND4 (N8196, N8194, N2874, N6072, N7617);
buf BUF1 (N8197, N8180);
nor NOR2 (N8198, N8190, N8153);
nand NAND4 (N8199, N8185, N6366, N895, N6987);
nand NAND3 (N8200, N8187, N5431, N6290);
xor XOR2 (N8201, N8193, N6370);
xor XOR2 (N8202, N8191, N4007);
nand NAND4 (N8203, N8198, N5563, N7297, N7857);
xor XOR2 (N8204, N8195, N2552);
buf BUF1 (N8205, N8204);
buf BUF1 (N8206, N8196);
nor NOR3 (N8207, N8184, N6411, N6515);
and AND2 (N8208, N8200, N6723);
xor XOR2 (N8209, N8203, N7036);
buf BUF1 (N8210, N8197);
buf BUF1 (N8211, N8199);
xor XOR2 (N8212, N8202, N4524);
nor NOR3 (N8213, N8205, N380, N2277);
xor XOR2 (N8214, N8192, N2114);
and AND4 (N8215, N8210, N6831, N2818, N326);
xor XOR2 (N8216, N8206, N1428);
nand NAND4 (N8217, N8214, N929, N3455, N2398);
or OR4 (N8218, N8201, N5694, N4716, N141);
nand NAND2 (N8219, N8208, N1116);
xor XOR2 (N8220, N8207, N6793);
buf BUF1 (N8221, N8216);
not NOT1 (N8222, N8213);
nor NOR2 (N8223, N8220, N5601);
or OR3 (N8224, N8218, N2025, N6640);
nand NAND3 (N8225, N8223, N288, N6598);
xor XOR2 (N8226, N8222, N1566);
or OR4 (N8227, N8211, N2765, N6017, N2208);
nand NAND2 (N8228, N8227, N1209);
nor NOR3 (N8229, N8209, N3722, N6555);
nand NAND4 (N8230, N8224, N8159, N6428, N1350);
buf BUF1 (N8231, N8215);
xor XOR2 (N8232, N8226, N4884);
xor XOR2 (N8233, N8232, N5914);
xor XOR2 (N8234, N8233, N1561);
buf BUF1 (N8235, N8231);
xor XOR2 (N8236, N8229, N277);
nor NOR3 (N8237, N8236, N2378, N1721);
not NOT1 (N8238, N8230);
xor XOR2 (N8239, N8235, N6393);
buf BUF1 (N8240, N8237);
xor XOR2 (N8241, N8240, N178);
or OR4 (N8242, N8225, N7882, N3214, N8105);
nor NOR4 (N8243, N8221, N2152, N6047, N4789);
nand NAND2 (N8244, N8217, N4739);
not NOT1 (N8245, N8212);
not NOT1 (N8246, N8234);
xor XOR2 (N8247, N8245, N6838);
and AND3 (N8248, N8242, N3417, N7402);
nand NAND2 (N8249, N8228, N1877);
buf BUF1 (N8250, N8247);
not NOT1 (N8251, N8250);
nor NOR2 (N8252, N8244, N5644);
and AND2 (N8253, N8243, N1875);
xor XOR2 (N8254, N8251, N5249);
not NOT1 (N8255, N8249);
xor XOR2 (N8256, N8238, N6215);
or OR2 (N8257, N8239, N6853);
nor NOR2 (N8258, N8253, N2630);
or OR4 (N8259, N8254, N4291, N4774, N5091);
buf BUF1 (N8260, N8248);
not NOT1 (N8261, N8258);
nand NAND2 (N8262, N8261, N6742);
buf BUF1 (N8263, N8262);
xor XOR2 (N8264, N8260, N2176);
not NOT1 (N8265, N8264);
xor XOR2 (N8266, N8265, N1180);
xor XOR2 (N8267, N8263, N6909);
nand NAND2 (N8268, N8267, N1679);
or OR4 (N8269, N8219, N3108, N5777, N2385);
buf BUF1 (N8270, N8269);
buf BUF1 (N8271, N8270);
nor NOR3 (N8272, N8241, N4399, N6650);
not NOT1 (N8273, N8256);
or OR3 (N8274, N8259, N5361, N535);
buf BUF1 (N8275, N8266);
or OR2 (N8276, N8246, N7887);
xor XOR2 (N8277, N8255, N214);
or OR2 (N8278, N8276, N1487);
nand NAND4 (N8279, N8277, N5458, N332, N4878);
and AND3 (N8280, N8271, N5440, N6822);
nand NAND4 (N8281, N8279, N1115, N142, N3545);
or OR3 (N8282, N8273, N3971, N3948);
and AND3 (N8283, N8275, N4776, N7350);
buf BUF1 (N8284, N8281);
buf BUF1 (N8285, N8268);
or OR4 (N8286, N8280, N3438, N4463, N107);
not NOT1 (N8287, N8283);
xor XOR2 (N8288, N8285, N3818);
nor NOR3 (N8289, N8278, N2102, N2072);
xor XOR2 (N8290, N8287, N8240);
or OR3 (N8291, N8288, N6900, N4149);
or OR4 (N8292, N8290, N7486, N6436, N4038);
nor NOR4 (N8293, N8291, N7025, N3826, N3371);
or OR2 (N8294, N8293, N8241);
or OR2 (N8295, N8282, N180);
or OR4 (N8296, N8257, N6092, N1858, N8059);
not NOT1 (N8297, N8295);
xor XOR2 (N8298, N8252, N3332);
xor XOR2 (N8299, N8294, N5807);
nand NAND3 (N8300, N8272, N4322, N682);
nor NOR4 (N8301, N8298, N1474, N3870, N2356);
nand NAND2 (N8302, N8301, N5369);
buf BUF1 (N8303, N8297);
and AND3 (N8304, N8289, N4133, N7754);
and AND3 (N8305, N8292, N1444, N3773);
and AND2 (N8306, N8304, N162);
and AND4 (N8307, N8296, N6767, N6594, N4031);
nor NOR2 (N8308, N8286, N2574);
nand NAND2 (N8309, N8302, N4068);
nand NAND4 (N8310, N8274, N3936, N5845, N4089);
nand NAND4 (N8311, N8303, N5969, N6705, N5567);
xor XOR2 (N8312, N8307, N6437);
not NOT1 (N8313, N8308);
and AND4 (N8314, N8299, N72, N7000, N5078);
nor NOR2 (N8315, N8309, N7259);
not NOT1 (N8316, N8310);
nor NOR4 (N8317, N8316, N7696, N5726, N3663);
not NOT1 (N8318, N8311);
nor NOR3 (N8319, N8318, N7246, N1722);
nor NOR4 (N8320, N8284, N1121, N4533, N8299);
xor XOR2 (N8321, N8314, N2449);
xor XOR2 (N8322, N8305, N3072);
xor XOR2 (N8323, N8320, N5837);
and AND2 (N8324, N8319, N7304);
nor NOR3 (N8325, N8323, N5863, N1977);
and AND3 (N8326, N8312, N4941, N7309);
buf BUF1 (N8327, N8317);
xor XOR2 (N8328, N8327, N6903);
buf BUF1 (N8329, N8322);
xor XOR2 (N8330, N8325, N3878);
and AND3 (N8331, N8330, N690, N953);
and AND2 (N8332, N8321, N966);
buf BUF1 (N8333, N8326);
and AND2 (N8334, N8324, N2576);
xor XOR2 (N8335, N8334, N978);
xor XOR2 (N8336, N8335, N7726);
xor XOR2 (N8337, N8329, N7360);
buf BUF1 (N8338, N8336);
and AND3 (N8339, N8331, N5814, N1661);
nand NAND3 (N8340, N8337, N6780, N2780);
or OR2 (N8341, N8306, N899);
xor XOR2 (N8342, N8328, N3083);
buf BUF1 (N8343, N8342);
buf BUF1 (N8344, N8333);
and AND2 (N8345, N8338, N6567);
or OR3 (N8346, N8332, N1753, N6795);
xor XOR2 (N8347, N8313, N3132);
buf BUF1 (N8348, N8343);
not NOT1 (N8349, N8346);
and AND4 (N8350, N8340, N427, N6264, N5361);
nor NOR2 (N8351, N8348, N1389);
xor XOR2 (N8352, N8341, N3783);
not NOT1 (N8353, N8315);
xor XOR2 (N8354, N8300, N7385);
buf BUF1 (N8355, N8345);
nand NAND3 (N8356, N8351, N1403, N3091);
xor XOR2 (N8357, N8339, N5731);
nand NAND3 (N8358, N8344, N5111, N6703);
nor NOR4 (N8359, N8358, N3407, N6394, N6295);
or OR2 (N8360, N8355, N6173);
or OR3 (N8361, N8353, N742, N8251);
nor NOR4 (N8362, N8350, N2779, N2421, N3649);
and AND3 (N8363, N8349, N4648, N1553);
or OR2 (N8364, N8362, N2914);
not NOT1 (N8365, N8354);
xor XOR2 (N8366, N8360, N3800);
and AND2 (N8367, N8356, N7878);
and AND4 (N8368, N8367, N8272, N3944, N1036);
buf BUF1 (N8369, N8366);
or OR4 (N8370, N8365, N504, N2680, N6140);
and AND4 (N8371, N8361, N1300, N7492, N7383);
or OR2 (N8372, N8369, N2904);
and AND3 (N8373, N8368, N6986, N4677);
xor XOR2 (N8374, N8352, N1192);
or OR4 (N8375, N8373, N1890, N918, N1454);
buf BUF1 (N8376, N8347);
nand NAND3 (N8377, N8363, N7263, N6786);
buf BUF1 (N8378, N8364);
or OR3 (N8379, N8378, N7592, N6781);
nand NAND4 (N8380, N8376, N6378, N6420, N4623);
and AND4 (N8381, N8379, N5255, N4890, N6747);
nor NOR2 (N8382, N8359, N4646);
or OR2 (N8383, N8357, N8297);
xor XOR2 (N8384, N8380, N8305);
nor NOR3 (N8385, N8382, N8199, N2612);
nor NOR2 (N8386, N8372, N5849);
and AND4 (N8387, N8385, N1070, N2866, N4977);
not NOT1 (N8388, N8381);
not NOT1 (N8389, N8371);
nand NAND2 (N8390, N8384, N1201);
not NOT1 (N8391, N8388);
xor XOR2 (N8392, N8383, N5023);
or OR4 (N8393, N8390, N6515, N1964, N1592);
buf BUF1 (N8394, N8389);
nand NAND3 (N8395, N8391, N89, N6328);
nand NAND4 (N8396, N8374, N4709, N2192, N8023);
not NOT1 (N8397, N8394);
or OR2 (N8398, N8386, N5351);
or OR2 (N8399, N8397, N1009);
nand NAND2 (N8400, N8393, N7161);
and AND4 (N8401, N8375, N3881, N3351, N6058);
xor XOR2 (N8402, N8400, N2727);
and AND4 (N8403, N8377, N839, N6019, N1624);
nor NOR4 (N8404, N8387, N588, N2292, N7539);
nand NAND3 (N8405, N8404, N7521, N6624);
nand NAND4 (N8406, N8398, N7962, N2537, N8190);
and AND3 (N8407, N8396, N5981, N5013);
nor NOR3 (N8408, N8407, N1611, N396);
xor XOR2 (N8409, N8395, N3726);
nor NOR3 (N8410, N8409, N6269, N4377);
buf BUF1 (N8411, N8370);
nand NAND4 (N8412, N8402, N3948, N7195, N8229);
nor NOR4 (N8413, N8399, N5733, N7215, N7571);
and AND3 (N8414, N8401, N1676, N5271);
nor NOR4 (N8415, N8411, N2484, N3581, N6172);
xor XOR2 (N8416, N8414, N5799);
and AND3 (N8417, N8405, N2681, N7576);
not NOT1 (N8418, N8413);
not NOT1 (N8419, N8408);
not NOT1 (N8420, N8419);
nor NOR3 (N8421, N8392, N7797, N3808);
buf BUF1 (N8422, N8412);
not NOT1 (N8423, N8415);
xor XOR2 (N8424, N8420, N1524);
nor NOR3 (N8425, N8403, N5888, N1681);
and AND2 (N8426, N8423, N4140);
not NOT1 (N8427, N8425);
nor NOR4 (N8428, N8426, N4132, N5737, N4927);
not NOT1 (N8429, N8421);
nand NAND2 (N8430, N8416, N3497);
and AND2 (N8431, N8428, N298);
and AND3 (N8432, N8418, N1344, N5726);
buf BUF1 (N8433, N8432);
or OR3 (N8434, N8410, N3388, N4254);
nand NAND4 (N8435, N8433, N855, N6468, N684);
buf BUF1 (N8436, N8435);
not NOT1 (N8437, N8430);
buf BUF1 (N8438, N8427);
not NOT1 (N8439, N8436);
buf BUF1 (N8440, N8437);
nand NAND2 (N8441, N8406, N8362);
and AND4 (N8442, N8439, N7091, N1365, N1502);
nor NOR2 (N8443, N8440, N3679);
not NOT1 (N8444, N8434);
nor NOR2 (N8445, N8442, N7339);
and AND3 (N8446, N8443, N851, N2470);
and AND4 (N8447, N8438, N679, N4799, N1623);
buf BUF1 (N8448, N8446);
and AND2 (N8449, N8444, N1703);
not NOT1 (N8450, N8417);
nand NAND2 (N8451, N8424, N632);
and AND2 (N8452, N8429, N645);
xor XOR2 (N8453, N8445, N3261);
nand NAND2 (N8454, N8449, N3379);
nand NAND3 (N8455, N8452, N2000, N6221);
nor NOR4 (N8456, N8450, N7148, N7235, N240);
not NOT1 (N8457, N8453);
buf BUF1 (N8458, N8454);
nor NOR4 (N8459, N8451, N3229, N3859, N5430);
nor NOR3 (N8460, N8422, N6550, N2553);
xor XOR2 (N8461, N8457, N247);
xor XOR2 (N8462, N8431, N8365);
or OR4 (N8463, N8455, N7684, N7649, N3062);
nor NOR4 (N8464, N8441, N8401, N5302, N2366);
and AND2 (N8465, N8461, N3946);
or OR2 (N8466, N8462, N1066);
not NOT1 (N8467, N8465);
xor XOR2 (N8468, N8464, N3745);
xor XOR2 (N8469, N8460, N7143);
and AND3 (N8470, N8467, N6706, N3986);
buf BUF1 (N8471, N8456);
buf BUF1 (N8472, N8468);
and AND4 (N8473, N8469, N1301, N2184, N4342);
not NOT1 (N8474, N8470);
nor NOR3 (N8475, N8448, N5566, N2044);
xor XOR2 (N8476, N8463, N3942);
or OR3 (N8477, N8466, N825, N6121);
nand NAND2 (N8478, N8471, N4892);
and AND4 (N8479, N8473, N2459, N3355, N8386);
not NOT1 (N8480, N8478);
and AND4 (N8481, N8474, N7923, N3399, N2358);
not NOT1 (N8482, N8481);
and AND3 (N8483, N8482, N1683, N3001);
nand NAND3 (N8484, N8472, N4963, N2213);
nor NOR4 (N8485, N8447, N6347, N3663, N5131);
buf BUF1 (N8486, N8479);
nor NOR4 (N8487, N8475, N74, N2482, N4481);
and AND4 (N8488, N8486, N8070, N3314, N7062);
or OR3 (N8489, N8488, N5142, N2085);
not NOT1 (N8490, N8485);
and AND3 (N8491, N8483, N1886, N4474);
and AND4 (N8492, N8487, N3412, N5085, N4664);
not NOT1 (N8493, N8458);
xor XOR2 (N8494, N8492, N948);
buf BUF1 (N8495, N8490);
or OR4 (N8496, N8477, N2906, N6505, N4596);
nor NOR2 (N8497, N8480, N3499);
buf BUF1 (N8498, N8497);
or OR3 (N8499, N8496, N3347, N1879);
nand NAND2 (N8500, N8499, N2954);
and AND4 (N8501, N8491, N725, N5863, N2752);
or OR2 (N8502, N8500, N3136);
xor XOR2 (N8503, N8494, N7368);
buf BUF1 (N8504, N8501);
nor NOR2 (N8505, N8459, N5406);
buf BUF1 (N8506, N8476);
xor XOR2 (N8507, N8505, N568);
or OR3 (N8508, N8503, N7246, N7066);
not NOT1 (N8509, N8508);
and AND3 (N8510, N8484, N7269, N2139);
and AND2 (N8511, N8510, N148);
buf BUF1 (N8512, N8498);
or OR2 (N8513, N8493, N4430);
nand NAND2 (N8514, N8495, N5350);
nand NAND4 (N8515, N8512, N3456, N671, N2767);
or OR3 (N8516, N8511, N2385, N545);
or OR4 (N8517, N8507, N5627, N2034, N4340);
nand NAND3 (N8518, N8506, N8130, N5249);
nand NAND2 (N8519, N8502, N1951);
and AND2 (N8520, N8518, N5613);
buf BUF1 (N8521, N8489);
buf BUF1 (N8522, N8513);
nor NOR3 (N8523, N8509, N8239, N3251);
buf BUF1 (N8524, N8516);
or OR2 (N8525, N8519, N7160);
nand NAND4 (N8526, N8522, N279, N2417, N3652);
xor XOR2 (N8527, N8523, N4403);
xor XOR2 (N8528, N8521, N2661);
xor XOR2 (N8529, N8520, N425);
or OR2 (N8530, N8528, N4938);
nand NAND4 (N8531, N8504, N6173, N4544, N3027);
or OR4 (N8532, N8517, N8133, N5997, N851);
buf BUF1 (N8533, N8532);
nor NOR4 (N8534, N8533, N5127, N2949, N5834);
nor NOR4 (N8535, N8530, N2564, N8369, N8400);
xor XOR2 (N8536, N8526, N5286);
xor XOR2 (N8537, N8525, N3171);
buf BUF1 (N8538, N8515);
and AND3 (N8539, N8534, N98, N1337);
not NOT1 (N8540, N8527);
not NOT1 (N8541, N8540);
xor XOR2 (N8542, N8541, N1880);
nor NOR3 (N8543, N8542, N3016, N3055);
not NOT1 (N8544, N8539);
not NOT1 (N8545, N8535);
buf BUF1 (N8546, N8536);
or OR4 (N8547, N8524, N2569, N5111, N6955);
nand NAND2 (N8548, N8538, N6164);
not NOT1 (N8549, N8544);
nand NAND3 (N8550, N8546, N1596, N6527);
xor XOR2 (N8551, N8549, N6475);
and AND3 (N8552, N8529, N3786, N690);
buf BUF1 (N8553, N8547);
not NOT1 (N8554, N8537);
xor XOR2 (N8555, N8531, N3182);
not NOT1 (N8556, N8551);
nand NAND2 (N8557, N8555, N6625);
nand NAND2 (N8558, N8543, N6568);
nor NOR4 (N8559, N8553, N1645, N421, N7173);
buf BUF1 (N8560, N8556);
xor XOR2 (N8561, N8557, N792);
xor XOR2 (N8562, N8561, N7879);
xor XOR2 (N8563, N8554, N2537);
xor XOR2 (N8564, N8548, N1694);
and AND2 (N8565, N8514, N1589);
and AND2 (N8566, N8560, N449);
or OR2 (N8567, N8550, N6554);
or OR3 (N8568, N8566, N7650, N7819);
or OR3 (N8569, N8552, N4391, N1973);
xor XOR2 (N8570, N8568, N339);
xor XOR2 (N8571, N8563, N5761);
nand NAND3 (N8572, N8559, N2295, N868);
xor XOR2 (N8573, N8545, N4475);
or OR4 (N8574, N8564, N6614, N6321, N1571);
and AND4 (N8575, N8569, N6658, N6519, N1125);
xor XOR2 (N8576, N8571, N4991);
buf BUF1 (N8577, N8562);
not NOT1 (N8578, N8567);
nand NAND3 (N8579, N8558, N7100, N6624);
nor NOR3 (N8580, N8574, N276, N4796);
or OR3 (N8581, N8576, N7544, N7297);
nor NOR4 (N8582, N8581, N4067, N6548, N643);
and AND4 (N8583, N8565, N7769, N4756, N8264);
buf BUF1 (N8584, N8583);
or OR2 (N8585, N8573, N3271);
nor NOR3 (N8586, N8580, N7554, N2551);
nand NAND3 (N8587, N8578, N1702, N6282);
xor XOR2 (N8588, N8584, N2828);
xor XOR2 (N8589, N8586, N873);
or OR2 (N8590, N8579, N5269);
and AND2 (N8591, N8577, N1520);
nand NAND4 (N8592, N8585, N1631, N454, N3208);
not NOT1 (N8593, N8587);
buf BUF1 (N8594, N8570);
and AND4 (N8595, N8575, N5551, N6793, N2881);
and AND3 (N8596, N8589, N4796, N7880);
buf BUF1 (N8597, N8593);
xor XOR2 (N8598, N8596, N5111);
buf BUF1 (N8599, N8588);
or OR4 (N8600, N8599, N5662, N3505, N4894);
or OR3 (N8601, N8572, N8438, N7214);
not NOT1 (N8602, N8598);
and AND3 (N8603, N8602, N5299, N3769);
or OR4 (N8604, N8592, N3357, N2568, N5519);
and AND4 (N8605, N8591, N8047, N1435, N7501);
not NOT1 (N8606, N8603);
nor NOR2 (N8607, N8605, N3107);
not NOT1 (N8608, N8607);
nor NOR2 (N8609, N8600, N1166);
xor XOR2 (N8610, N8608, N5956);
and AND2 (N8611, N8594, N3042);
or OR3 (N8612, N8610, N2982, N3817);
nor NOR2 (N8613, N8611, N4957);
nand NAND4 (N8614, N8612, N3427, N4127, N8292);
nor NOR3 (N8615, N8614, N3167, N5348);
and AND3 (N8616, N8604, N7227, N3683);
xor XOR2 (N8617, N8582, N6771);
xor XOR2 (N8618, N8617, N1564);
nand NAND2 (N8619, N8613, N8069);
nor NOR4 (N8620, N8597, N5303, N2989, N3224);
nand NAND4 (N8621, N8615, N577, N6478, N3235);
buf BUF1 (N8622, N8619);
or OR3 (N8623, N8621, N130, N2631);
nor NOR4 (N8624, N8595, N2042, N2397, N753);
not NOT1 (N8625, N8623);
not NOT1 (N8626, N8624);
nor NOR3 (N8627, N8590, N7752, N6180);
or OR3 (N8628, N8626, N5750, N3779);
not NOT1 (N8629, N8628);
buf BUF1 (N8630, N8616);
xor XOR2 (N8631, N8622, N4023);
and AND2 (N8632, N8631, N3704);
and AND4 (N8633, N8601, N463, N6795, N5882);
nand NAND2 (N8634, N8627, N6806);
xor XOR2 (N8635, N8609, N1554);
or OR4 (N8636, N8635, N8082, N5607, N3727);
or OR3 (N8637, N8629, N4861, N3045);
and AND3 (N8638, N8636, N3024, N3073);
and AND4 (N8639, N8632, N4661, N1720, N4520);
nor NOR2 (N8640, N8639, N6048);
and AND3 (N8641, N8637, N3770, N3654);
nand NAND2 (N8642, N8630, N1853);
xor XOR2 (N8643, N8641, N3886);
and AND4 (N8644, N8634, N5048, N309, N2078);
and AND3 (N8645, N8640, N4454, N926);
nor NOR2 (N8646, N8644, N4433);
not NOT1 (N8647, N8645);
xor XOR2 (N8648, N8606, N415);
and AND4 (N8649, N8620, N3510, N7174, N5054);
xor XOR2 (N8650, N8646, N3567);
buf BUF1 (N8651, N8618);
or OR2 (N8652, N8638, N2333);
nor NOR3 (N8653, N8652, N3640, N7989);
or OR2 (N8654, N8647, N1092);
not NOT1 (N8655, N8651);
nand NAND3 (N8656, N8650, N7652, N5857);
nor NOR3 (N8657, N8633, N6939, N6495);
or OR3 (N8658, N8648, N1182, N1296);
not NOT1 (N8659, N8658);
xor XOR2 (N8660, N8655, N5360);
nand NAND2 (N8661, N8659, N3735);
and AND2 (N8662, N8657, N1168);
xor XOR2 (N8663, N8660, N2489);
xor XOR2 (N8664, N8654, N677);
buf BUF1 (N8665, N8662);
or OR2 (N8666, N8664, N1377);
and AND2 (N8667, N8661, N5401);
buf BUF1 (N8668, N8653);
nand NAND4 (N8669, N8666, N3953, N2202, N239);
not NOT1 (N8670, N8643);
not NOT1 (N8671, N8668);
xor XOR2 (N8672, N8671, N927);
and AND3 (N8673, N8672, N4461, N1304);
buf BUF1 (N8674, N8670);
nor NOR3 (N8675, N8665, N2071, N6458);
xor XOR2 (N8676, N8649, N2851);
nor NOR3 (N8677, N8669, N7313, N6494);
nor NOR4 (N8678, N8642, N1076, N3415, N8394);
and AND3 (N8679, N8673, N6749, N6604);
or OR3 (N8680, N8663, N3219, N1556);
nand NAND4 (N8681, N8679, N323, N5247, N2033);
nand NAND4 (N8682, N8675, N5117, N7943, N3859);
and AND2 (N8683, N8625, N4986);
buf BUF1 (N8684, N8656);
not NOT1 (N8685, N8667);
xor XOR2 (N8686, N8677, N5259);
buf BUF1 (N8687, N8684);
or OR4 (N8688, N8674, N421, N8143, N3740);
nor NOR2 (N8689, N8682, N4286);
nor NOR3 (N8690, N8681, N2920, N8037);
buf BUF1 (N8691, N8688);
xor XOR2 (N8692, N8686, N2169);
not NOT1 (N8693, N8683);
and AND3 (N8694, N8685, N4143, N2541);
or OR4 (N8695, N8678, N3544, N4345, N8496);
nand NAND2 (N8696, N8690, N1852);
and AND2 (N8697, N8691, N8206);
xor XOR2 (N8698, N8692, N7381);
and AND4 (N8699, N8680, N667, N7617, N6785);
nor NOR4 (N8700, N8693, N3937, N3678, N2958);
or OR4 (N8701, N8676, N6673, N3880, N108);
buf BUF1 (N8702, N8695);
and AND3 (N8703, N8697, N5526, N2357);
not NOT1 (N8704, N8696);
and AND2 (N8705, N8700, N4997);
not NOT1 (N8706, N8704);
buf BUF1 (N8707, N8699);
not NOT1 (N8708, N8703);
xor XOR2 (N8709, N8706, N4934);
xor XOR2 (N8710, N8702, N3978);
not NOT1 (N8711, N8707);
not NOT1 (N8712, N8709);
xor XOR2 (N8713, N8701, N83);
and AND2 (N8714, N8708, N7997);
xor XOR2 (N8715, N8711, N3354);
not NOT1 (N8716, N8713);
nor NOR3 (N8717, N8712, N8481, N4889);
not NOT1 (N8718, N8717);
nand NAND4 (N8719, N8694, N4675, N8279, N6386);
or OR2 (N8720, N8714, N7505);
and AND3 (N8721, N8720, N3247, N1719);
nor NOR4 (N8722, N8710, N8480, N4247, N6220);
and AND2 (N8723, N8689, N2966);
and AND4 (N8724, N8721, N2834, N7849, N4871);
not NOT1 (N8725, N8698);
xor XOR2 (N8726, N8725, N4311);
nand NAND3 (N8727, N8715, N4587, N3096);
nand NAND2 (N8728, N8716, N4851);
buf BUF1 (N8729, N8727);
or OR3 (N8730, N8722, N3874, N4233);
and AND4 (N8731, N8728, N8158, N5045, N5391);
nand NAND2 (N8732, N8687, N267);
xor XOR2 (N8733, N8724, N5821);
nand NAND4 (N8734, N8733, N4374, N5446, N1134);
not NOT1 (N8735, N8729);
and AND3 (N8736, N8718, N7642, N7387);
not NOT1 (N8737, N8731);
buf BUF1 (N8738, N8735);
buf BUF1 (N8739, N8734);
buf BUF1 (N8740, N8726);
nand NAND3 (N8741, N8739, N2624, N2089);
or OR3 (N8742, N8736, N4463, N2409);
and AND4 (N8743, N8705, N6669, N1545, N1500);
buf BUF1 (N8744, N8738);
not NOT1 (N8745, N8741);
nand NAND3 (N8746, N8742, N1338, N3146);
and AND4 (N8747, N8719, N134, N3664, N4056);
xor XOR2 (N8748, N8737, N6331);
nand NAND3 (N8749, N8723, N3505, N6242);
or OR2 (N8750, N8748, N2958);
or OR4 (N8751, N8750, N5353, N8093, N1465);
xor XOR2 (N8752, N8745, N2359);
buf BUF1 (N8753, N8732);
xor XOR2 (N8754, N8752, N2701);
xor XOR2 (N8755, N8749, N6639);
or OR4 (N8756, N8754, N2900, N4537, N4535);
nand NAND2 (N8757, N8746, N7225);
nor NOR2 (N8758, N8743, N4523);
nor NOR4 (N8759, N8747, N7164, N6157, N6344);
nand NAND3 (N8760, N8758, N6627, N526);
or OR2 (N8761, N8753, N6298);
xor XOR2 (N8762, N8761, N5917);
xor XOR2 (N8763, N8740, N8443);
nor NOR2 (N8764, N8730, N4756);
or OR3 (N8765, N8764, N8566, N1279);
or OR3 (N8766, N8762, N4357, N428);
buf BUF1 (N8767, N8760);
and AND2 (N8768, N8755, N4573);
and AND4 (N8769, N8765, N1220, N2956, N3697);
or OR4 (N8770, N8767, N4701, N1203, N6114);
nand NAND4 (N8771, N8769, N6101, N5188, N7872);
nor NOR4 (N8772, N8766, N834, N3170, N4834);
buf BUF1 (N8773, N8771);
nor NOR2 (N8774, N8751, N3299);
xor XOR2 (N8775, N8756, N3138);
buf BUF1 (N8776, N8763);
or OR2 (N8777, N8759, N1364);
buf BUF1 (N8778, N8770);
not NOT1 (N8779, N8778);
nor NOR3 (N8780, N8779, N4809, N8708);
and AND2 (N8781, N8773, N8348);
xor XOR2 (N8782, N8774, N1247);
xor XOR2 (N8783, N8780, N2190);
not NOT1 (N8784, N8744);
nor NOR2 (N8785, N8776, N2981);
and AND4 (N8786, N8772, N1957, N4551, N3233);
buf BUF1 (N8787, N8785);
or OR4 (N8788, N8787, N514, N617, N3420);
nor NOR4 (N8789, N8777, N4967, N218, N527);
or OR3 (N8790, N8775, N3124, N1509);
and AND3 (N8791, N8781, N8177, N7441);
and AND4 (N8792, N8788, N5867, N1479, N772);
and AND2 (N8793, N8792, N3813);
and AND3 (N8794, N8782, N5856, N4429);
or OR4 (N8795, N8793, N5602, N8129, N4359);
not NOT1 (N8796, N8784);
xor XOR2 (N8797, N8791, N2889);
xor XOR2 (N8798, N8768, N6689);
not NOT1 (N8799, N8783);
buf BUF1 (N8800, N8799);
nand NAND2 (N8801, N8794, N1367);
nor NOR2 (N8802, N8797, N6019);
not NOT1 (N8803, N8786);
xor XOR2 (N8804, N8796, N573);
nand NAND2 (N8805, N8795, N649);
xor XOR2 (N8806, N8803, N608);
nor NOR3 (N8807, N8806, N2431, N2267);
or OR3 (N8808, N8757, N5408, N5305);
nor NOR2 (N8809, N8800, N1412);
buf BUF1 (N8810, N8789);
xor XOR2 (N8811, N8809, N2346);
and AND4 (N8812, N8790, N1714, N8222, N3446);
not NOT1 (N8813, N8807);
and AND3 (N8814, N8812, N2119, N6531);
nor NOR2 (N8815, N8813, N1910);
xor XOR2 (N8816, N8801, N455);
nand NAND4 (N8817, N8811, N2123, N1354, N237);
and AND2 (N8818, N8804, N6531);
or OR4 (N8819, N8802, N748, N5701, N8619);
not NOT1 (N8820, N8818);
buf BUF1 (N8821, N8810);
nor NOR2 (N8822, N8798, N8494);
or OR2 (N8823, N8814, N7686);
or OR3 (N8824, N8805, N6069, N5356);
buf BUF1 (N8825, N8822);
nand NAND3 (N8826, N8823, N3627, N4555);
and AND4 (N8827, N8821, N5164, N3377, N214);
buf BUF1 (N8828, N8817);
and AND3 (N8829, N8808, N8274, N7443);
nor NOR2 (N8830, N8824, N5030);
and AND2 (N8831, N8820, N825);
buf BUF1 (N8832, N8829);
buf BUF1 (N8833, N8816);
xor XOR2 (N8834, N8826, N5592);
or OR3 (N8835, N8825, N1332, N3309);
buf BUF1 (N8836, N8834);
or OR3 (N8837, N8835, N4454, N3274);
and AND3 (N8838, N8836, N7051, N6331);
xor XOR2 (N8839, N8832, N213);
or OR2 (N8840, N8830, N3962);
nand NAND2 (N8841, N8827, N5321);
buf BUF1 (N8842, N8837);
nand NAND2 (N8843, N8840, N7682);
nand NAND3 (N8844, N8815, N4575, N1848);
not NOT1 (N8845, N8842);
and AND2 (N8846, N8831, N638);
nor NOR3 (N8847, N8828, N3036, N6756);
buf BUF1 (N8848, N8843);
buf BUF1 (N8849, N8844);
nand NAND3 (N8850, N8848, N8745, N2916);
or OR3 (N8851, N8833, N700, N345);
nor NOR2 (N8852, N8851, N7479);
nor NOR3 (N8853, N8847, N5544, N3855);
or OR2 (N8854, N8838, N1574);
or OR4 (N8855, N8853, N8376, N5968, N1731);
buf BUF1 (N8856, N8854);
nor NOR4 (N8857, N8849, N6034, N443, N5209);
or OR2 (N8858, N8846, N3360);
not NOT1 (N8859, N8857);
nor NOR4 (N8860, N8841, N7274, N1359, N7795);
xor XOR2 (N8861, N8852, N3448);
xor XOR2 (N8862, N8839, N6143);
xor XOR2 (N8863, N8850, N8564);
or OR2 (N8864, N8855, N5746);
xor XOR2 (N8865, N8860, N1705);
and AND2 (N8866, N8863, N6207);
xor XOR2 (N8867, N8862, N208);
nor NOR2 (N8868, N8864, N2427);
or OR3 (N8869, N8865, N8429, N7596);
not NOT1 (N8870, N8858);
not NOT1 (N8871, N8859);
xor XOR2 (N8872, N8868, N6862);
xor XOR2 (N8873, N8870, N2282);
and AND3 (N8874, N8866, N3002, N8577);
nand NAND2 (N8875, N8861, N1552);
or OR2 (N8876, N8872, N7000);
xor XOR2 (N8877, N8875, N4807);
not NOT1 (N8878, N8856);
and AND3 (N8879, N8877, N6258, N4198);
not NOT1 (N8880, N8871);
or OR4 (N8881, N8819, N3155, N213, N1939);
or OR2 (N8882, N8874, N5286);
xor XOR2 (N8883, N8880, N1733);
nor NOR3 (N8884, N8881, N3320, N1529);
xor XOR2 (N8885, N8884, N6096);
nor NOR4 (N8886, N8845, N3590, N4000, N3219);
buf BUF1 (N8887, N8883);
not NOT1 (N8888, N8886);
xor XOR2 (N8889, N8867, N4962);
xor XOR2 (N8890, N8887, N5740);
xor XOR2 (N8891, N8879, N148);
xor XOR2 (N8892, N8889, N2906);
or OR3 (N8893, N8888, N514, N7788);
nor NOR4 (N8894, N8893, N4100, N3508, N2169);
nand NAND2 (N8895, N8869, N1346);
or OR3 (N8896, N8882, N8873, N299);
buf BUF1 (N8897, N5730);
xor XOR2 (N8898, N8890, N158);
buf BUF1 (N8899, N8896);
or OR2 (N8900, N8892, N2388);
and AND4 (N8901, N8885, N4107, N2828, N3710);
nor NOR4 (N8902, N8897, N3441, N400, N4377);
nor NOR4 (N8903, N8901, N1739, N3300, N4107);
nor NOR3 (N8904, N8900, N7412, N8479);
not NOT1 (N8905, N8895);
not NOT1 (N8906, N8878);
nand NAND4 (N8907, N8903, N7560, N3737, N3031);
xor XOR2 (N8908, N8902, N7142);
nand NAND2 (N8909, N8898, N8273);
nand NAND2 (N8910, N8899, N523);
nand NAND4 (N8911, N8906, N7884, N812, N5877);
nor NOR2 (N8912, N8905, N1816);
xor XOR2 (N8913, N8891, N6089);
nor NOR2 (N8914, N8908, N6340);
nand NAND2 (N8915, N8911, N719);
buf BUF1 (N8916, N8907);
nor NOR4 (N8917, N8913, N4354, N3557, N4590);
nor NOR3 (N8918, N8912, N2119, N204);
nand NAND4 (N8919, N8909, N4532, N3342, N7398);
xor XOR2 (N8920, N8915, N8184);
buf BUF1 (N8921, N8914);
buf BUF1 (N8922, N8894);
xor XOR2 (N8923, N8920, N7840);
nand NAND3 (N8924, N8917, N4724, N1893);
buf BUF1 (N8925, N8904);
xor XOR2 (N8926, N8923, N7871);
nor NOR4 (N8927, N8926, N529, N684, N895);
not NOT1 (N8928, N8918);
not NOT1 (N8929, N8924);
nor NOR2 (N8930, N8910, N8179);
nor NOR3 (N8931, N8930, N7563, N2473);
nand NAND2 (N8932, N8931, N8694);
not NOT1 (N8933, N8928);
and AND3 (N8934, N8916, N6359, N166);
or OR2 (N8935, N8932, N5475);
and AND2 (N8936, N8876, N7714);
xor XOR2 (N8937, N8934, N7074);
xor XOR2 (N8938, N8935, N7018);
nand NAND2 (N8939, N8922, N5313);
nand NAND2 (N8940, N8919, N7849);
nor NOR4 (N8941, N8936, N2638, N5634, N5399);
nor NOR2 (N8942, N8938, N2581);
or OR3 (N8943, N8927, N1394, N5182);
or OR2 (N8944, N8929, N725);
nand NAND2 (N8945, N8937, N3363);
not NOT1 (N8946, N8939);
not NOT1 (N8947, N8943);
xor XOR2 (N8948, N8921, N5748);
or OR3 (N8949, N8941, N8259, N8866);
or OR4 (N8950, N8948, N6071, N2801, N3715);
and AND4 (N8951, N8933, N4197, N7830, N5619);
not NOT1 (N8952, N8942);
buf BUF1 (N8953, N8951);
not NOT1 (N8954, N8944);
nand NAND3 (N8955, N8952, N7453, N5243);
nand NAND4 (N8956, N8946, N952, N8762, N3154);
not NOT1 (N8957, N8925);
and AND2 (N8958, N8950, N6287);
xor XOR2 (N8959, N8945, N4207);
nand NAND2 (N8960, N8958, N4260);
nand NAND4 (N8961, N8940, N7139, N4621, N3186);
xor XOR2 (N8962, N8947, N2284);
and AND3 (N8963, N8953, N7683, N3143);
xor XOR2 (N8964, N8957, N7690);
and AND2 (N8965, N8949, N1214);
or OR4 (N8966, N8956, N4870, N8509, N235);
nor NOR2 (N8967, N8965, N7028);
nor NOR3 (N8968, N8960, N8400, N6354);
and AND3 (N8969, N8968, N8012, N202);
buf BUF1 (N8970, N8955);
and AND3 (N8971, N8964, N7602, N7875);
xor XOR2 (N8972, N8954, N5055);
or OR3 (N8973, N8972, N1776, N1814);
nand NAND4 (N8974, N8970, N6712, N8681, N6443);
nor NOR2 (N8975, N8974, N2713);
nor NOR3 (N8976, N8969, N210, N1363);
and AND2 (N8977, N8962, N5372);
not NOT1 (N8978, N8961);
buf BUF1 (N8979, N8973);
not NOT1 (N8980, N8976);
not NOT1 (N8981, N8959);
not NOT1 (N8982, N8980);
nand NAND3 (N8983, N8966, N160, N5710);
not NOT1 (N8984, N8963);
and AND4 (N8985, N8975, N1377, N4366, N6100);
nor NOR4 (N8986, N8984, N71, N8103, N6205);
xor XOR2 (N8987, N8983, N8092);
not NOT1 (N8988, N8971);
buf BUF1 (N8989, N8987);
nand NAND4 (N8990, N8967, N4606, N8211, N609);
not NOT1 (N8991, N8982);
nor NOR3 (N8992, N8988, N6521, N7049);
xor XOR2 (N8993, N8985, N4262);
not NOT1 (N8994, N8989);
nand NAND4 (N8995, N8981, N8716, N2922, N1068);
nor NOR2 (N8996, N8977, N3540);
or OR3 (N8997, N8979, N8407, N1954);
or OR2 (N8998, N8990, N7429);
buf BUF1 (N8999, N8993);
or OR4 (N9000, N8997, N8693, N8577, N1416);
nand NAND3 (N9001, N8998, N8395, N1143);
or OR3 (N9002, N8996, N4473, N8122);
xor XOR2 (N9003, N8978, N5847);
nor NOR4 (N9004, N9000, N2549, N7285, N4972);
nand NAND4 (N9005, N8991, N8663, N672, N1143);
xor XOR2 (N9006, N9004, N8114);
nand NAND4 (N9007, N8992, N3856, N444, N7674);
and AND3 (N9008, N9003, N2196, N4772);
buf BUF1 (N9009, N9005);
nand NAND3 (N9010, N9008, N6772, N3876);
nand NAND4 (N9011, N9006, N1698, N3987, N8491);
nor NOR3 (N9012, N8999, N6550, N617);
and AND3 (N9013, N9002, N3878, N5311);
buf BUF1 (N9014, N9011);
not NOT1 (N9015, N8995);
nand NAND4 (N9016, N8994, N6729, N692, N8157);
xor XOR2 (N9017, N9013, N7267);
not NOT1 (N9018, N9016);
xor XOR2 (N9019, N9009, N8873);
not NOT1 (N9020, N9018);
nor NOR4 (N9021, N9017, N4688, N5051, N1933);
nand NAND3 (N9022, N9019, N5408, N7348);
buf BUF1 (N9023, N9014);
not NOT1 (N9024, N8986);
buf BUF1 (N9025, N9010);
nor NOR3 (N9026, N9020, N2549, N4443);
buf BUF1 (N9027, N9024);
nor NOR3 (N9028, N9001, N3685, N5998);
and AND4 (N9029, N9026, N2549, N5015, N1621);
nor NOR3 (N9030, N9028, N2890, N6440);
nand NAND3 (N9031, N9025, N4960, N445);
or OR4 (N9032, N9027, N2738, N8486, N7367);
not NOT1 (N9033, N9022);
buf BUF1 (N9034, N9007);
nand NAND3 (N9035, N9023, N8461, N4207);
nand NAND2 (N9036, N9035, N1233);
xor XOR2 (N9037, N9030, N7556);
buf BUF1 (N9038, N9032);
or OR3 (N9039, N9033, N394, N5954);
or OR3 (N9040, N9012, N5369, N8711);
or OR4 (N9041, N9034, N1681, N6481, N6434);
nand NAND4 (N9042, N9038, N6255, N28, N884);
buf BUF1 (N9043, N9037);
nand NAND2 (N9044, N9040, N2604);
xor XOR2 (N9045, N9015, N5490);
buf BUF1 (N9046, N9041);
buf BUF1 (N9047, N9036);
nand NAND2 (N9048, N9039, N3281);
or OR2 (N9049, N9048, N3049);
buf BUF1 (N9050, N9044);
or OR4 (N9051, N9049, N6026, N3687, N506);
xor XOR2 (N9052, N9051, N1442);
or OR4 (N9053, N9047, N182, N120, N3686);
nand NAND3 (N9054, N9045, N6600, N4044);
nor NOR2 (N9055, N9046, N674);
not NOT1 (N9056, N9050);
nor NOR4 (N9057, N9053, N2706, N7182, N4121);
and AND4 (N9058, N9057, N1815, N4170, N6535);
not NOT1 (N9059, N9052);
xor XOR2 (N9060, N9058, N6066);
xor XOR2 (N9061, N9031, N1626);
xor XOR2 (N9062, N9042, N693);
not NOT1 (N9063, N9055);
nor NOR2 (N9064, N9062, N1677);
xor XOR2 (N9065, N9060, N8639);
xor XOR2 (N9066, N9021, N3318);
or OR3 (N9067, N9065, N8783, N3186);
xor XOR2 (N9068, N9063, N2513);
xor XOR2 (N9069, N9066, N3129);
xor XOR2 (N9070, N9067, N161);
nand NAND3 (N9071, N9069, N4003, N4986);
not NOT1 (N9072, N9043);
not NOT1 (N9073, N9070);
not NOT1 (N9074, N9073);
not NOT1 (N9075, N9071);
buf BUF1 (N9076, N9064);
and AND2 (N9077, N9059, N3584);
buf BUF1 (N9078, N9074);
and AND2 (N9079, N9054, N5724);
and AND3 (N9080, N9068, N8966, N2935);
and AND2 (N9081, N9056, N3812);
not NOT1 (N9082, N9079);
nand NAND4 (N9083, N9078, N1579, N8741, N1987);
nand NAND4 (N9084, N9081, N8689, N3583, N5778);
buf BUF1 (N9085, N9076);
nor NOR3 (N9086, N9075, N5120, N1975);
xor XOR2 (N9087, N9080, N3449);
xor XOR2 (N9088, N9087, N2239);
nor NOR4 (N9089, N9029, N7583, N5599, N1231);
buf BUF1 (N9090, N9083);
nor NOR2 (N9091, N9061, N1818);
not NOT1 (N9092, N9090);
nand NAND3 (N9093, N9088, N8203, N2116);
nor NOR2 (N9094, N9091, N2299);
and AND2 (N9095, N9085, N7166);
buf BUF1 (N9096, N9086);
nor NOR4 (N9097, N9092, N2115, N7479, N4449);
not NOT1 (N9098, N9097);
buf BUF1 (N9099, N9094);
nor NOR4 (N9100, N9084, N294, N1909, N681);
nand NAND3 (N9101, N9096, N4738, N1506);
and AND2 (N9102, N9101, N8897);
and AND3 (N9103, N9093, N9075, N5455);
not NOT1 (N9104, N9077);
or OR2 (N9105, N9095, N4635);
xor XOR2 (N9106, N9098, N3962);
xor XOR2 (N9107, N9082, N6343);
xor XOR2 (N9108, N9105, N3209);
not NOT1 (N9109, N9089);
buf BUF1 (N9110, N9107);
xor XOR2 (N9111, N9110, N8860);
xor XOR2 (N9112, N9100, N1090);
and AND4 (N9113, N9103, N385, N798, N5894);
not NOT1 (N9114, N9113);
or OR3 (N9115, N9111, N4071, N638);
or OR4 (N9116, N9112, N4679, N2154, N3668);
not NOT1 (N9117, N9099);
nand NAND3 (N9118, N9115, N555, N2112);
and AND4 (N9119, N9118, N2791, N5218, N9064);
xor XOR2 (N9120, N9108, N8878);
nand NAND4 (N9121, N9117, N3797, N5849, N5300);
nand NAND3 (N9122, N9072, N6421, N1748);
nor NOR3 (N9123, N9109, N9026, N2154);
nand NAND2 (N9124, N9104, N7041);
nor NOR2 (N9125, N9120, N7821);
or OR2 (N9126, N9123, N846);
not NOT1 (N9127, N9116);
or OR3 (N9128, N9122, N7233, N2000);
xor XOR2 (N9129, N9127, N2875);
or OR3 (N9130, N9114, N6755, N2382);
or OR4 (N9131, N9124, N7206, N3361, N7807);
or OR2 (N9132, N9106, N8225);
buf BUF1 (N9133, N9126);
xor XOR2 (N9134, N9129, N6938);
nor NOR3 (N9135, N9128, N5874, N1060);
nand NAND3 (N9136, N9125, N4356, N5075);
and AND3 (N9137, N9132, N4657, N6314);
nor NOR4 (N9138, N9133, N2867, N2440, N1157);
buf BUF1 (N9139, N9137);
nor NOR4 (N9140, N9134, N6780, N5252, N4420);
buf BUF1 (N9141, N9140);
xor XOR2 (N9142, N9119, N7793);
xor XOR2 (N9143, N9121, N5551);
not NOT1 (N9144, N9139);
nand NAND4 (N9145, N9102, N538, N2390, N1752);
nand NAND3 (N9146, N9131, N3910, N5114);
nand NAND3 (N9147, N9144, N8300, N2212);
or OR2 (N9148, N9146, N9110);
and AND2 (N9149, N9147, N8085);
or OR3 (N9150, N9130, N4131, N4063);
buf BUF1 (N9151, N9142);
xor XOR2 (N9152, N9136, N6850);
xor XOR2 (N9153, N9141, N2436);
or OR4 (N9154, N9148, N3859, N16, N6025);
not NOT1 (N9155, N9151);
or OR2 (N9156, N9154, N8571);
or OR4 (N9157, N9156, N3952, N2208, N838);
nor NOR3 (N9158, N9145, N2429, N2308);
nand NAND4 (N9159, N9149, N2658, N1843, N303);
and AND2 (N9160, N9159, N4577);
nand NAND2 (N9161, N9143, N3086);
not NOT1 (N9162, N9135);
xor XOR2 (N9163, N9138, N1052);
nor NOR3 (N9164, N9157, N7891, N7655);
buf BUF1 (N9165, N9152);
or OR4 (N9166, N9155, N2362, N6195, N6180);
buf BUF1 (N9167, N9162);
buf BUF1 (N9168, N9153);
buf BUF1 (N9169, N9160);
and AND3 (N9170, N9158, N3798, N4602);
xor XOR2 (N9171, N9150, N6830);
nor NOR4 (N9172, N9166, N1112, N6615, N2895);
and AND2 (N9173, N9163, N4350);
nor NOR4 (N9174, N9170, N6664, N2078, N5849);
and AND4 (N9175, N9167, N6967, N4612, N5300);
xor XOR2 (N9176, N9161, N3152);
and AND2 (N9177, N9172, N8806);
or OR2 (N9178, N9176, N2009);
buf BUF1 (N9179, N9169);
not NOT1 (N9180, N9164);
not NOT1 (N9181, N9165);
nor NOR3 (N9182, N9175, N7903, N6313);
not NOT1 (N9183, N9182);
and AND2 (N9184, N9181, N2914);
nand NAND4 (N9185, N9173, N6040, N5809, N8298);
nand NAND2 (N9186, N9180, N8688);
buf BUF1 (N9187, N9171);
or OR2 (N9188, N9185, N7296);
or OR4 (N9189, N9188, N1642, N3029, N3421);
not NOT1 (N9190, N9186);
xor XOR2 (N9191, N9183, N9009);
and AND2 (N9192, N9191, N2057);
or OR3 (N9193, N9178, N1711, N4822);
and AND3 (N9194, N9193, N751, N5143);
xor XOR2 (N9195, N9184, N2972);
and AND3 (N9196, N9189, N3515, N9002);
not NOT1 (N9197, N9194);
and AND2 (N9198, N9179, N2781);
nor NOR3 (N9199, N9195, N1905, N8226);
nor NOR3 (N9200, N9192, N1731, N2503);
and AND3 (N9201, N9174, N6750, N7300);
and AND4 (N9202, N9197, N2226, N8830, N7742);
and AND3 (N9203, N9187, N1124, N2397);
buf BUF1 (N9204, N9196);
nor NOR4 (N9205, N9168, N5795, N6891, N1704);
buf BUF1 (N9206, N9177);
or OR4 (N9207, N9206, N1238, N4643, N7016);
or OR4 (N9208, N9200, N4195, N8263, N1271);
nand NAND2 (N9209, N9203, N5514);
xor XOR2 (N9210, N9205, N982);
or OR4 (N9211, N9190, N1155, N2829, N5891);
and AND4 (N9212, N9201, N7456, N5435, N2269);
and AND3 (N9213, N9199, N7897, N3534);
or OR3 (N9214, N9212, N2534, N6311);
buf BUF1 (N9215, N9209);
not NOT1 (N9216, N9211);
buf BUF1 (N9217, N9207);
not NOT1 (N9218, N9213);
not NOT1 (N9219, N9215);
nor NOR2 (N9220, N9218, N5939);
not NOT1 (N9221, N9219);
and AND3 (N9222, N9220, N3690, N4618);
nor NOR4 (N9223, N9198, N857, N1056, N7597);
not NOT1 (N9224, N9214);
or OR4 (N9225, N9224, N489, N7694, N4550);
xor XOR2 (N9226, N9221, N4393);
or OR4 (N9227, N9204, N295, N6563, N7128);
buf BUF1 (N9228, N9226);
nor NOR4 (N9229, N9217, N1303, N4721, N6382);
nand NAND2 (N9230, N9228, N4422);
nor NOR3 (N9231, N9216, N5631, N6194);
nand NAND4 (N9232, N9210, N3682, N2057, N7509);
nor NOR3 (N9233, N9222, N4784, N1008);
xor XOR2 (N9234, N9208, N3543);
nor NOR3 (N9235, N9227, N1624, N6396);
nand NAND2 (N9236, N9233, N931);
xor XOR2 (N9237, N9225, N2556);
and AND2 (N9238, N9223, N5024);
not NOT1 (N9239, N9229);
nor NOR4 (N9240, N9231, N815, N8988, N6475);
nor NOR4 (N9241, N9237, N8026, N8100, N3939);
and AND4 (N9242, N9238, N1563, N7961, N8623);
nor NOR4 (N9243, N9240, N681, N3563, N2629);
or OR2 (N9244, N9241, N7873);
nor NOR4 (N9245, N9236, N4493, N9116, N8071);
or OR4 (N9246, N9230, N4211, N5087, N4029);
buf BUF1 (N9247, N9234);
or OR3 (N9248, N9247, N3242, N2696);
buf BUF1 (N9249, N9242);
nand NAND3 (N9250, N9232, N5621, N7199);
or OR2 (N9251, N9235, N2269);
not NOT1 (N9252, N9239);
or OR3 (N9253, N9251, N619, N5898);
xor XOR2 (N9254, N9243, N6394);
or OR2 (N9255, N9254, N1788);
or OR2 (N9256, N9253, N7777);
nor NOR4 (N9257, N9245, N711, N2301, N1190);
or OR4 (N9258, N9202, N8710, N5145, N7267);
xor XOR2 (N9259, N9257, N8930);
xor XOR2 (N9260, N9252, N7032);
buf BUF1 (N9261, N9248);
xor XOR2 (N9262, N9259, N7727);
and AND3 (N9263, N9258, N724, N2443);
nand NAND4 (N9264, N9249, N766, N4415, N8140);
or OR4 (N9265, N9250, N3385, N8620, N6115);
or OR3 (N9266, N9256, N5829, N8569);
nand NAND3 (N9267, N9246, N1013, N8136);
nand NAND3 (N9268, N9260, N2944, N8661);
or OR3 (N9269, N9244, N5188, N658);
nor NOR4 (N9270, N9269, N8879, N6548, N434);
xor XOR2 (N9271, N9265, N2172);
and AND3 (N9272, N9270, N7095, N2578);
not NOT1 (N9273, N9271);
xor XOR2 (N9274, N9268, N1309);
buf BUF1 (N9275, N9267);
xor XOR2 (N9276, N9266, N452);
buf BUF1 (N9277, N9273);
xor XOR2 (N9278, N9276, N968);
xor XOR2 (N9279, N9277, N9000);
xor XOR2 (N9280, N9262, N2868);
not NOT1 (N9281, N9263);
xor XOR2 (N9282, N9255, N4685);
nand NAND3 (N9283, N9261, N7718, N1247);
buf BUF1 (N9284, N9274);
buf BUF1 (N9285, N9281);
not NOT1 (N9286, N9278);
and AND2 (N9287, N9283, N2084);
and AND3 (N9288, N9280, N5835, N4283);
xor XOR2 (N9289, N9264, N2260);
not NOT1 (N9290, N9282);
or OR3 (N9291, N9290, N5607, N3104);
or OR3 (N9292, N9287, N8029, N2561);
and AND3 (N9293, N9286, N1886, N4003);
buf BUF1 (N9294, N9275);
not NOT1 (N9295, N9285);
buf BUF1 (N9296, N9293);
xor XOR2 (N9297, N9288, N8000);
and AND2 (N9298, N9291, N8868);
xor XOR2 (N9299, N9292, N6005);
and AND2 (N9300, N9298, N4657);
xor XOR2 (N9301, N9294, N3439);
or OR3 (N9302, N9301, N2953, N3074);
buf BUF1 (N9303, N9272);
nor NOR2 (N9304, N9299, N7135);
or OR3 (N9305, N9295, N5538, N93);
or OR4 (N9306, N9289, N5903, N8283, N7389);
nor NOR2 (N9307, N9300, N8891);
nand NAND3 (N9308, N9304, N4838, N196);
and AND3 (N9309, N9303, N5116, N1630);
or OR4 (N9310, N9309, N5983, N1755, N3856);
or OR2 (N9311, N9296, N4756);
buf BUF1 (N9312, N9306);
xor XOR2 (N9313, N9311, N8237);
not NOT1 (N9314, N9312);
nor NOR3 (N9315, N9305, N870, N8125);
nor NOR2 (N9316, N9310, N6160);
nand NAND3 (N9317, N9279, N1634, N3438);
or OR2 (N9318, N9308, N4106);
or OR2 (N9319, N9307, N7729);
and AND4 (N9320, N9313, N3008, N4373, N2664);
and AND4 (N9321, N9316, N2612, N8757, N3595);
buf BUF1 (N9322, N9320);
and AND3 (N9323, N9302, N4505, N2397);
xor XOR2 (N9324, N9323, N5537);
buf BUF1 (N9325, N9315);
or OR3 (N9326, N9318, N8093, N4758);
and AND4 (N9327, N9324, N1613, N5216, N1015);
and AND3 (N9328, N9297, N4204, N8628);
or OR2 (N9329, N9328, N6975);
buf BUF1 (N9330, N9314);
not NOT1 (N9331, N9326);
or OR3 (N9332, N9331, N893, N5630);
and AND2 (N9333, N9329, N598);
nand NAND3 (N9334, N9327, N6555, N1468);
and AND3 (N9335, N9334, N6773, N6545);
buf BUF1 (N9336, N9332);
xor XOR2 (N9337, N9325, N1623);
or OR3 (N9338, N9337, N6833, N695);
buf BUF1 (N9339, N9319);
nor NOR2 (N9340, N9317, N3557);
and AND2 (N9341, N9336, N3129);
not NOT1 (N9342, N9340);
and AND2 (N9343, N9341, N2357);
xor XOR2 (N9344, N9322, N3106);
nand NAND3 (N9345, N9344, N3385, N2029);
buf BUF1 (N9346, N9335);
nor NOR4 (N9347, N9339, N3048, N4859, N7485);
buf BUF1 (N9348, N9338);
nor NOR2 (N9349, N9346, N2313);
and AND2 (N9350, N9333, N2597);
nand NAND4 (N9351, N9342, N4451, N1963, N7700);
not NOT1 (N9352, N9321);
xor XOR2 (N9353, N9330, N8877);
nor NOR4 (N9354, N9347, N2785, N601, N8048);
xor XOR2 (N9355, N9284, N4974);
buf BUF1 (N9356, N9349);
xor XOR2 (N9357, N9351, N98);
not NOT1 (N9358, N9352);
buf BUF1 (N9359, N9358);
xor XOR2 (N9360, N9357, N984);
or OR3 (N9361, N9348, N4644, N9171);
not NOT1 (N9362, N9343);
or OR3 (N9363, N9362, N2789, N7028);
nor NOR3 (N9364, N9356, N7983, N5200);
and AND3 (N9365, N9364, N6400, N7926);
and AND2 (N9366, N9354, N7948);
not NOT1 (N9367, N9366);
xor XOR2 (N9368, N9359, N2517);
and AND2 (N9369, N9350, N4873);
nand NAND4 (N9370, N9361, N2839, N7016, N1591);
xor XOR2 (N9371, N9370, N294);
not NOT1 (N9372, N9368);
nand NAND2 (N9373, N9371, N6521);
xor XOR2 (N9374, N9360, N5225);
nor NOR4 (N9375, N9372, N8126, N3547, N8801);
buf BUF1 (N9376, N9353);
or OR3 (N9377, N9355, N6176, N8501);
nor NOR2 (N9378, N9373, N8912);
buf BUF1 (N9379, N9377);
nand NAND2 (N9380, N9345, N2265);
and AND2 (N9381, N9374, N1209);
and AND2 (N9382, N9376, N5091);
xor XOR2 (N9383, N9367, N1991);
xor XOR2 (N9384, N9383, N2233);
buf BUF1 (N9385, N9382);
not NOT1 (N9386, N9384);
nand NAND2 (N9387, N9378, N840);
or OR2 (N9388, N9386, N5042);
nand NAND4 (N9389, N9387, N3851, N6080, N2503);
nand NAND2 (N9390, N9363, N6558);
and AND4 (N9391, N9388, N7679, N3707, N8261);
nor NOR3 (N9392, N9385, N916, N974);
nand NAND4 (N9393, N9392, N8139, N8770, N5852);
or OR2 (N9394, N9365, N5961);
buf BUF1 (N9395, N9389);
nor NOR2 (N9396, N9390, N5585);
and AND3 (N9397, N9393, N4411, N1695);
not NOT1 (N9398, N9381);
xor XOR2 (N9399, N9379, N4287);
not NOT1 (N9400, N9369);
or OR4 (N9401, N9396, N3249, N2004, N3958);
nor NOR3 (N9402, N9397, N1616, N2808);
nand NAND4 (N9403, N9400, N9220, N4818, N5298);
buf BUF1 (N9404, N9395);
buf BUF1 (N9405, N9402);
not NOT1 (N9406, N9405);
xor XOR2 (N9407, N9399, N4670);
nand NAND4 (N9408, N9375, N8570, N7497, N1584);
buf BUF1 (N9409, N9380);
not NOT1 (N9410, N9404);
not NOT1 (N9411, N9394);
or OR4 (N9412, N9410, N9350, N2619, N6470);
not NOT1 (N9413, N9406);
buf BUF1 (N9414, N9391);
or OR3 (N9415, N9413, N9236, N1135);
not NOT1 (N9416, N9403);
buf BUF1 (N9417, N9409);
or OR3 (N9418, N9412, N8342, N8236);
buf BUF1 (N9419, N9408);
nor NOR3 (N9420, N9407, N1950, N2138);
nor NOR3 (N9421, N9401, N5276, N1032);
xor XOR2 (N9422, N9420, N4788);
not NOT1 (N9423, N9414);
nor NOR2 (N9424, N9422, N7799);
buf BUF1 (N9425, N9417);
and AND4 (N9426, N9416, N4261, N3629, N509);
nand NAND4 (N9427, N9421, N8932, N1929, N3108);
xor XOR2 (N9428, N9411, N301);
and AND2 (N9429, N9423, N7809);
not NOT1 (N9430, N9429);
not NOT1 (N9431, N9425);
nand NAND2 (N9432, N9427, N5215);
or OR4 (N9433, N9432, N8224, N1426, N5858);
xor XOR2 (N9434, N9428, N1952);
and AND4 (N9435, N9431, N5005, N6927, N7445);
and AND4 (N9436, N9415, N8919, N2173, N9112);
buf BUF1 (N9437, N9419);
buf BUF1 (N9438, N9430);
xor XOR2 (N9439, N9438, N6230);
not NOT1 (N9440, N9437);
and AND4 (N9441, N9424, N9362, N393, N4814);
xor XOR2 (N9442, N9435, N1842);
buf BUF1 (N9443, N9434);
and AND4 (N9444, N9439, N2672, N1663, N4525);
buf BUF1 (N9445, N9398);
or OR3 (N9446, N9441, N5581, N2092);
or OR4 (N9447, N9446, N5363, N5413, N865);
not NOT1 (N9448, N9442);
buf BUF1 (N9449, N9445);
and AND2 (N9450, N9433, N5756);
buf BUF1 (N9451, N9418);
buf BUF1 (N9452, N9436);
not NOT1 (N9453, N9426);
xor XOR2 (N9454, N9448, N4864);
nor NOR4 (N9455, N9454, N3051, N5319, N2222);
xor XOR2 (N9456, N9451, N2110);
and AND2 (N9457, N9453, N6309);
and AND4 (N9458, N9443, N3639, N7413, N7344);
nor NOR4 (N9459, N9455, N5882, N8254, N3502);
or OR3 (N9460, N9458, N6292, N591);
xor XOR2 (N9461, N9460, N6961);
nand NAND3 (N9462, N9452, N5470, N864);
buf BUF1 (N9463, N9462);
and AND3 (N9464, N9463, N1056, N4391);
nand NAND4 (N9465, N9457, N1425, N5002, N9104);
nand NAND4 (N9466, N9464, N5737, N8911, N2705);
buf BUF1 (N9467, N9450);
not NOT1 (N9468, N9459);
nor NOR4 (N9469, N9465, N2406, N7895, N1147);
nand NAND2 (N9470, N9469, N8060);
or OR4 (N9471, N9467, N5373, N3536, N3881);
or OR2 (N9472, N9470, N6514);
xor XOR2 (N9473, N9471, N3656);
not NOT1 (N9474, N9468);
and AND4 (N9475, N9461, N6649, N1415, N1540);
not NOT1 (N9476, N9440);
and AND4 (N9477, N9476, N5789, N2018, N3878);
xor XOR2 (N9478, N9477, N2794);
nor NOR4 (N9479, N9449, N6707, N3072, N8077);
xor XOR2 (N9480, N9478, N7019);
nand NAND4 (N9481, N9474, N3725, N1173, N9314);
or OR4 (N9482, N9480, N1748, N2251, N1520);
or OR4 (N9483, N9475, N1541, N8264, N3645);
or OR4 (N9484, N9482, N3392, N7649, N2733);
nand NAND2 (N9485, N9481, N4176);
buf BUF1 (N9486, N9472);
buf BUF1 (N9487, N9473);
or OR2 (N9488, N9487, N8032);
and AND4 (N9489, N9488, N2016, N2539, N9029);
and AND2 (N9490, N9479, N8565);
nand NAND2 (N9491, N9484, N1694);
nand NAND2 (N9492, N9456, N389);
buf BUF1 (N9493, N9490);
and AND3 (N9494, N9492, N7660, N2438);
buf BUF1 (N9495, N9466);
nor NOR2 (N9496, N9489, N328);
not NOT1 (N9497, N9486);
xor XOR2 (N9498, N9485, N5897);
nand NAND3 (N9499, N9494, N1819, N7228);
xor XOR2 (N9500, N9447, N3525);
buf BUF1 (N9501, N9493);
or OR2 (N9502, N9483, N521);
xor XOR2 (N9503, N9497, N33);
nor NOR2 (N9504, N9491, N7372);
and AND2 (N9505, N9503, N4376);
nand NAND2 (N9506, N9505, N3971);
and AND4 (N9507, N9444, N9249, N4351, N812);
xor XOR2 (N9508, N9502, N6854);
not NOT1 (N9509, N9506);
nand NAND2 (N9510, N9504, N649);
nand NAND2 (N9511, N9508, N7176);
buf BUF1 (N9512, N9511);
or OR4 (N9513, N9496, N2880, N1701, N4927);
not NOT1 (N9514, N9499);
and AND3 (N9515, N9500, N2975, N8790);
not NOT1 (N9516, N9509);
nor NOR4 (N9517, N9507, N2901, N2194, N2089);
nor NOR2 (N9518, N9514, N7145);
nor NOR3 (N9519, N9512, N46, N6600);
nor NOR4 (N9520, N9519, N2765, N9177, N1644);
and AND2 (N9521, N9518, N918);
nor NOR3 (N9522, N9516, N7068, N4689);
buf BUF1 (N9523, N9521);
and AND2 (N9524, N9510, N4882);
xor XOR2 (N9525, N9498, N3672);
or OR2 (N9526, N9524, N8430);
nand NAND4 (N9527, N9523, N6205, N8048, N4581);
nand NAND2 (N9528, N9525, N5719);
or OR3 (N9529, N9520, N873, N6073);
nand NAND4 (N9530, N9515, N965, N4333, N6129);
nand NAND3 (N9531, N9495, N3222, N8905);
buf BUF1 (N9532, N9522);
and AND3 (N9533, N9513, N3409, N7603);
nand NAND2 (N9534, N9526, N1207);
or OR2 (N9535, N9529, N3581);
buf BUF1 (N9536, N9528);
buf BUF1 (N9537, N9535);
xor XOR2 (N9538, N9501, N2222);
nor NOR3 (N9539, N9531, N5509, N3674);
not NOT1 (N9540, N9517);
nand NAND2 (N9541, N9530, N6652);
nor NOR4 (N9542, N9527, N2709, N9014, N1860);
nand NAND4 (N9543, N9533, N163, N8455, N4846);
nand NAND2 (N9544, N9536, N153);
or OR3 (N9545, N9542, N1670, N6811);
nor NOR4 (N9546, N9532, N7396, N9445, N1222);
not NOT1 (N9547, N9544);
xor XOR2 (N9548, N9547, N419);
not NOT1 (N9549, N9545);
and AND2 (N9550, N9546, N5801);
and AND3 (N9551, N9534, N2103, N2305);
nor NOR3 (N9552, N9540, N4259, N6819);
xor XOR2 (N9553, N9543, N5701);
nor NOR3 (N9554, N9548, N459, N4505);
or OR3 (N9555, N9554, N2875, N4827);
xor XOR2 (N9556, N9539, N4261);
nor NOR2 (N9557, N9552, N1311);
nand NAND3 (N9558, N9553, N8717, N4729);
buf BUF1 (N9559, N9556);
or OR3 (N9560, N9551, N2172, N1925);
and AND4 (N9561, N9558, N9367, N8095, N8051);
or OR2 (N9562, N9561, N1503);
and AND2 (N9563, N9555, N3430);
buf BUF1 (N9564, N9541);
xor XOR2 (N9565, N9560, N624);
not NOT1 (N9566, N9537);
nor NOR3 (N9567, N9565, N3415, N751);
not NOT1 (N9568, N9566);
or OR3 (N9569, N9564, N6833, N1837);
and AND3 (N9570, N9567, N127, N3170);
buf BUF1 (N9571, N9569);
nor NOR2 (N9572, N9562, N8143);
not NOT1 (N9573, N9568);
or OR4 (N9574, N9550, N9048, N2115, N7899);
xor XOR2 (N9575, N9559, N1775);
nand NAND2 (N9576, N9572, N4827);
not NOT1 (N9577, N9574);
or OR4 (N9578, N9573, N5583, N4597, N5321);
xor XOR2 (N9579, N9549, N669);
not NOT1 (N9580, N9538);
nand NAND4 (N9581, N9570, N4238, N2170, N558);
not NOT1 (N9582, N9557);
xor XOR2 (N9583, N9577, N3448);
buf BUF1 (N9584, N9583);
or OR4 (N9585, N9578, N470, N2167, N1052);
buf BUF1 (N9586, N9576);
or OR4 (N9587, N9585, N9079, N4287, N4046);
not NOT1 (N9588, N9586);
nor NOR4 (N9589, N9575, N5874, N7216, N9380);
xor XOR2 (N9590, N9563, N7738);
buf BUF1 (N9591, N9584);
buf BUF1 (N9592, N9587);
or OR4 (N9593, N9571, N1465, N2068, N976);
nor NOR3 (N9594, N9580, N2885, N3854);
nand NAND2 (N9595, N9594, N8173);
nor NOR2 (N9596, N9589, N5245);
xor XOR2 (N9597, N9582, N4313);
or OR4 (N9598, N9579, N4732, N3165, N3105);
and AND2 (N9599, N9592, N7020);
and AND3 (N9600, N9588, N6277, N7674);
and AND2 (N9601, N9593, N5687);
xor XOR2 (N9602, N9591, N3828);
nor NOR4 (N9603, N9596, N7142, N2518, N5772);
and AND2 (N9604, N9599, N4244);
buf BUF1 (N9605, N9598);
nand NAND2 (N9606, N9605, N8298);
buf BUF1 (N9607, N9606);
nand NAND4 (N9608, N9590, N1522, N4532, N7627);
nor NOR2 (N9609, N9604, N4580);
nand NAND2 (N9610, N9602, N7687);
nand NAND3 (N9611, N9601, N3528, N681);
and AND4 (N9612, N9608, N45, N7940, N600);
not NOT1 (N9613, N9595);
nand NAND2 (N9614, N9611, N7594);
nand NAND3 (N9615, N9613, N9399, N8477);
nand NAND4 (N9616, N9603, N4700, N5418, N6119);
nor NOR2 (N9617, N9597, N4792);
xor XOR2 (N9618, N9610, N9159);
buf BUF1 (N9619, N9612);
and AND2 (N9620, N9607, N7879);
and AND4 (N9621, N9614, N2870, N8364, N8831);
buf BUF1 (N9622, N9616);
nor NOR2 (N9623, N9615, N2303);
nor NOR3 (N9624, N9623, N7031, N2998);
nand NAND3 (N9625, N9581, N3497, N66);
buf BUF1 (N9626, N9620);
nand NAND3 (N9627, N9617, N8739, N1487);
and AND3 (N9628, N9600, N4426, N8423);
or OR2 (N9629, N9609, N6966);
or OR4 (N9630, N9627, N8937, N5688, N8110);
xor XOR2 (N9631, N9625, N3045);
nor NOR4 (N9632, N9618, N79, N2405, N409);
nor NOR2 (N9633, N9621, N4254);
nand NAND2 (N9634, N9630, N442);
nor NOR4 (N9635, N9631, N4045, N6346, N7972);
xor XOR2 (N9636, N9635, N9494);
not NOT1 (N9637, N9619);
or OR4 (N9638, N9634, N5238, N6600, N2613);
not NOT1 (N9639, N9622);
not NOT1 (N9640, N9636);
nand NAND4 (N9641, N9626, N608, N3707, N491);
and AND3 (N9642, N9638, N8323, N8869);
buf BUF1 (N9643, N9628);
nand NAND3 (N9644, N9632, N221, N7143);
xor XOR2 (N9645, N9644, N539);
buf BUF1 (N9646, N9642);
and AND2 (N9647, N9629, N5496);
or OR2 (N9648, N9624, N8812);
nor NOR2 (N9649, N9648, N3182);
nand NAND2 (N9650, N9637, N7381);
xor XOR2 (N9651, N9647, N1129);
buf BUF1 (N9652, N9651);
not NOT1 (N9653, N9650);
and AND3 (N9654, N9640, N6946, N5014);
or OR2 (N9655, N9641, N331);
or OR2 (N9656, N9639, N5366);
nand NAND2 (N9657, N9633, N3530);
nor NOR4 (N9658, N9657, N9174, N5665, N8628);
nand NAND3 (N9659, N9655, N7535, N3860);
buf BUF1 (N9660, N9649);
nand NAND2 (N9661, N9646, N2120);
buf BUF1 (N9662, N9654);
buf BUF1 (N9663, N9660);
xor XOR2 (N9664, N9663, N7043);
nand NAND4 (N9665, N9659, N7335, N7885, N294);
nor NOR4 (N9666, N9652, N2924, N5634, N4216);
nor NOR2 (N9667, N9658, N6172);
not NOT1 (N9668, N9643);
not NOT1 (N9669, N9645);
xor XOR2 (N9670, N9664, N7215);
and AND3 (N9671, N9661, N7487, N7929);
or OR3 (N9672, N9665, N4464, N1551);
buf BUF1 (N9673, N9662);
xor XOR2 (N9674, N9656, N6222);
not NOT1 (N9675, N9668);
not NOT1 (N9676, N9672);
not NOT1 (N9677, N9670);
xor XOR2 (N9678, N9671, N8804);
or OR4 (N9679, N9666, N9059, N4694, N7612);
and AND3 (N9680, N9673, N5961, N7421);
xor XOR2 (N9681, N9680, N4748);
nor NOR3 (N9682, N9675, N981, N5152);
nand NAND3 (N9683, N9677, N3746, N2047);
or OR3 (N9684, N9681, N4983, N1588);
not NOT1 (N9685, N9653);
or OR3 (N9686, N9676, N7502, N4198);
and AND3 (N9687, N9674, N8211, N9469);
nor NOR4 (N9688, N9686, N2783, N610, N1756);
buf BUF1 (N9689, N9669);
nand NAND4 (N9690, N9678, N345, N9650, N4745);
not NOT1 (N9691, N9667);
not NOT1 (N9692, N9684);
buf BUF1 (N9693, N9689);
nor NOR4 (N9694, N9679, N446, N2369, N5048);
nor NOR3 (N9695, N9687, N3586, N485);
and AND2 (N9696, N9683, N8378);
and AND2 (N9697, N9693, N1135);
xor XOR2 (N9698, N9691, N8320);
buf BUF1 (N9699, N9692);
or OR2 (N9700, N9699, N2146);
nand NAND4 (N9701, N9700, N525, N4149, N2477);
and AND2 (N9702, N9701, N6646);
buf BUF1 (N9703, N9695);
xor XOR2 (N9704, N9703, N281);
not NOT1 (N9705, N9702);
and AND3 (N9706, N9690, N6433, N5650);
not NOT1 (N9707, N9696);
not NOT1 (N9708, N9706);
buf BUF1 (N9709, N9698);
not NOT1 (N9710, N9704);
nor NOR4 (N9711, N9710, N4109, N7179, N9008);
buf BUF1 (N9712, N9694);
xor XOR2 (N9713, N9709, N8041);
and AND3 (N9714, N9685, N3726, N5298);
and AND4 (N9715, N9682, N8506, N6196, N6280);
and AND3 (N9716, N9707, N2742, N3386);
buf BUF1 (N9717, N9708);
nand NAND2 (N9718, N9688, N2262);
and AND3 (N9719, N9716, N1662, N925);
not NOT1 (N9720, N9711);
and AND3 (N9721, N9715, N329, N430);
or OR2 (N9722, N9721, N5558);
not NOT1 (N9723, N9697);
and AND3 (N9724, N9718, N6592, N4594);
nor NOR4 (N9725, N9724, N8939, N39, N3543);
and AND4 (N9726, N9717, N895, N7639, N674);
nand NAND2 (N9727, N9714, N8749);
nor NOR2 (N9728, N9723, N2410);
or OR4 (N9729, N9727, N4103, N1142, N6603);
buf BUF1 (N9730, N9720);
or OR2 (N9731, N9719, N648);
xor XOR2 (N9732, N9725, N6012);
not NOT1 (N9733, N9728);
and AND4 (N9734, N9729, N9730, N792, N1927);
not NOT1 (N9735, N2291);
and AND2 (N9736, N9731, N6154);
or OR2 (N9737, N9733, N3780);
or OR2 (N9738, N9726, N4244);
nand NAND4 (N9739, N9737, N9165, N5803, N4703);
or OR3 (N9740, N9713, N50, N998);
nand NAND2 (N9741, N9712, N7516);
nand NAND2 (N9742, N9722, N5052);
and AND3 (N9743, N9738, N6954, N1963);
not NOT1 (N9744, N9736);
nor NOR4 (N9745, N9740, N8044, N4690, N2069);
nor NOR3 (N9746, N9742, N3164, N9355);
or OR4 (N9747, N9705, N5307, N4486, N8727);
nand NAND3 (N9748, N9735, N2927, N4658);
xor XOR2 (N9749, N9746, N9234);
not NOT1 (N9750, N9749);
buf BUF1 (N9751, N9744);
nor NOR4 (N9752, N9734, N8714, N299, N4913);
or OR3 (N9753, N9745, N2444, N4561);
not NOT1 (N9754, N9753);
nand NAND4 (N9755, N9748, N5414, N4455, N9075);
or OR3 (N9756, N9739, N280, N8167);
nand NAND3 (N9757, N9741, N2330, N8481);
not NOT1 (N9758, N9751);
xor XOR2 (N9759, N9752, N2335);
nand NAND4 (N9760, N9756, N3682, N6988, N9436);
buf BUF1 (N9761, N9760);
buf BUF1 (N9762, N9750);
buf BUF1 (N9763, N9758);
not NOT1 (N9764, N9754);
nor NOR2 (N9765, N9761, N8094);
nand NAND3 (N9766, N9755, N3110, N758);
or OR3 (N9767, N9765, N3291, N8634);
buf BUF1 (N9768, N9763);
nor NOR4 (N9769, N9732, N2739, N2675, N5538);
nand NAND4 (N9770, N9767, N2427, N8744, N9655);
not NOT1 (N9771, N9762);
not NOT1 (N9772, N9747);
xor XOR2 (N9773, N9770, N5074);
or OR3 (N9774, N9759, N5363, N1827);
nand NAND2 (N9775, N9766, N7937);
xor XOR2 (N9776, N9771, N1747);
and AND4 (N9777, N9757, N2594, N8145, N7838);
not NOT1 (N9778, N9776);
buf BUF1 (N9779, N9777);
not NOT1 (N9780, N9764);
buf BUF1 (N9781, N9773);
or OR4 (N9782, N9743, N7545, N3361, N1842);
nor NOR4 (N9783, N9780, N7545, N5553, N7809);
not NOT1 (N9784, N9772);
nor NOR4 (N9785, N9782, N7050, N4538, N4682);
xor XOR2 (N9786, N9778, N2362);
buf BUF1 (N9787, N9769);
nand NAND2 (N9788, N9784, N5544);
nor NOR4 (N9789, N9774, N4255, N7992, N8917);
buf BUF1 (N9790, N9768);
xor XOR2 (N9791, N9783, N7527);
and AND2 (N9792, N9781, N6004);
nor NOR2 (N9793, N9788, N8724);
not NOT1 (N9794, N9793);
nand NAND4 (N9795, N9785, N1573, N3884, N6808);
and AND4 (N9796, N9790, N6005, N6904, N4772);
not NOT1 (N9797, N9786);
and AND3 (N9798, N9795, N3127, N3942);
nand NAND4 (N9799, N9797, N9193, N538, N4898);
or OR3 (N9800, N9791, N6116, N7516);
xor XOR2 (N9801, N9794, N7974);
not NOT1 (N9802, N9779);
buf BUF1 (N9803, N9775);
and AND4 (N9804, N9802, N4517, N4665, N1812);
buf BUF1 (N9805, N9798);
nand NAND3 (N9806, N9801, N7488, N4160);
nand NAND2 (N9807, N9800, N1997);
nor NOR3 (N9808, N9789, N2182, N4020);
buf BUF1 (N9809, N9808);
buf BUF1 (N9810, N9809);
xor XOR2 (N9811, N9804, N1739);
and AND2 (N9812, N9796, N1841);
buf BUF1 (N9813, N9807);
nand NAND3 (N9814, N9805, N5664, N7460);
nor NOR3 (N9815, N9811, N8995, N2543);
and AND4 (N9816, N9810, N995, N2077, N2576);
and AND3 (N9817, N9799, N7282, N1574);
and AND3 (N9818, N9814, N1748, N3623);
xor XOR2 (N9819, N9787, N8202);
xor XOR2 (N9820, N9817, N7797);
nand NAND3 (N9821, N9820, N8801, N2112);
buf BUF1 (N9822, N9806);
nand NAND3 (N9823, N9822, N210, N5164);
not NOT1 (N9824, N9812);
buf BUF1 (N9825, N9823);
buf BUF1 (N9826, N9815);
or OR4 (N9827, N9826, N3971, N7077, N4430);
not NOT1 (N9828, N9818);
nor NOR4 (N9829, N9827, N4939, N2465, N2722);
or OR4 (N9830, N9821, N295, N5666, N9746);
and AND3 (N9831, N9829, N6694, N9348);
buf BUF1 (N9832, N9831);
and AND4 (N9833, N9819, N2294, N1510, N176);
xor XOR2 (N9834, N9792, N1839);
xor XOR2 (N9835, N9813, N3906);
buf BUF1 (N9836, N9803);
or OR4 (N9837, N9835, N4792, N261, N9728);
not NOT1 (N9838, N9828);
xor XOR2 (N9839, N9836, N9518);
or OR2 (N9840, N9838, N6115);
nand NAND3 (N9841, N9840, N6032, N3042);
nor NOR3 (N9842, N9834, N8128, N511);
xor XOR2 (N9843, N9837, N8679);
buf BUF1 (N9844, N9842);
buf BUF1 (N9845, N9843);
or OR3 (N9846, N9844, N8508, N7184);
nand NAND2 (N9847, N9833, N5391);
nor NOR2 (N9848, N9816, N4874);
or OR2 (N9849, N9841, N9751);
not NOT1 (N9850, N9847);
buf BUF1 (N9851, N9849);
or OR4 (N9852, N9824, N991, N6520, N4375);
or OR2 (N9853, N9846, N2688);
and AND4 (N9854, N9853, N9129, N9162, N1142);
nor NOR4 (N9855, N9845, N8857, N9618, N4391);
not NOT1 (N9856, N9852);
nor NOR2 (N9857, N9848, N1756);
nand NAND3 (N9858, N9825, N7195, N5352);
nand NAND2 (N9859, N9858, N6676);
and AND4 (N9860, N9830, N2432, N6007, N184);
and AND2 (N9861, N9851, N2196);
nor NOR3 (N9862, N9850, N3810, N2748);
xor XOR2 (N9863, N9855, N9603);
nand NAND2 (N9864, N9854, N6001);
nor NOR2 (N9865, N9863, N1625);
and AND3 (N9866, N9860, N3021, N3812);
buf BUF1 (N9867, N9866);
or OR3 (N9868, N9859, N6605, N1688);
xor XOR2 (N9869, N9865, N4690);
not NOT1 (N9870, N9861);
nor NOR3 (N9871, N9870, N8106, N7998);
xor XOR2 (N9872, N9871, N5420);
nor NOR3 (N9873, N9839, N8194, N4006);
nand NAND4 (N9874, N9864, N8186, N609, N2930);
and AND2 (N9875, N9868, N6394);
not NOT1 (N9876, N9874);
or OR4 (N9877, N9873, N7703, N4988, N1171);
not NOT1 (N9878, N9856);
and AND3 (N9879, N9876, N8027, N5297);
buf BUF1 (N9880, N9877);
nor NOR2 (N9881, N9875, N170);
not NOT1 (N9882, N9881);
nand NAND3 (N9883, N9857, N3041, N2706);
xor XOR2 (N9884, N9867, N5106);
buf BUF1 (N9885, N9872);
and AND2 (N9886, N9882, N1880);
nand NAND4 (N9887, N9878, N9456, N535, N5961);
buf BUF1 (N9888, N9887);
nor NOR3 (N9889, N9880, N7689, N4983);
nand NAND3 (N9890, N9879, N6171, N6556);
or OR3 (N9891, N9886, N6989, N7418);
buf BUF1 (N9892, N9883);
buf BUF1 (N9893, N9885);
nand NAND4 (N9894, N9890, N3792, N9605, N6274);
nor NOR3 (N9895, N9892, N3225, N8764);
not NOT1 (N9896, N9862);
buf BUF1 (N9897, N9869);
and AND2 (N9898, N9891, N8383);
not NOT1 (N9899, N9832);
or OR2 (N9900, N9899, N7506);
not NOT1 (N9901, N9884);
and AND2 (N9902, N9901, N5271);
and AND2 (N9903, N9893, N9454);
buf BUF1 (N9904, N9900);
not NOT1 (N9905, N9903);
not NOT1 (N9906, N9896);
xor XOR2 (N9907, N9898, N7791);
nand NAND2 (N9908, N9902, N9766);
xor XOR2 (N9909, N9905, N966);
or OR3 (N9910, N9907, N9114, N4634);
nor NOR3 (N9911, N9895, N9714, N4513);
nor NOR4 (N9912, N9908, N8751, N2669, N2604);
xor XOR2 (N9913, N9889, N2148);
and AND4 (N9914, N9910, N1786, N9775, N8526);
nand NAND4 (N9915, N9888, N9016, N4494, N8948);
buf BUF1 (N9916, N9915);
buf BUF1 (N9917, N9913);
or OR2 (N9918, N9911, N4323);
buf BUF1 (N9919, N9912);
nor NOR4 (N9920, N9916, N3093, N3629, N2149);
nor NOR4 (N9921, N9920, N7458, N9473, N207);
not NOT1 (N9922, N9917);
buf BUF1 (N9923, N9922);
nand NAND4 (N9924, N9904, N6020, N2731, N9798);
and AND3 (N9925, N9924, N3937, N6111);
or OR4 (N9926, N9909, N5868, N1026, N9188);
nand NAND4 (N9927, N9918, N8169, N7742, N6635);
and AND3 (N9928, N9894, N3283, N4831);
nor NOR3 (N9929, N9926, N7769, N4446);
and AND3 (N9930, N9906, N8841, N1269);
nand NAND2 (N9931, N9897, N7529);
and AND2 (N9932, N9930, N2043);
and AND3 (N9933, N9921, N479, N4670);
nand NAND3 (N9934, N9927, N3907, N1871);
nor NOR2 (N9935, N9919, N2314);
or OR3 (N9936, N9931, N9837, N5269);
buf BUF1 (N9937, N9936);
buf BUF1 (N9938, N9933);
xor XOR2 (N9939, N9932, N2933);
nand NAND3 (N9940, N9928, N2516, N8208);
nor NOR4 (N9941, N9934, N5039, N2862, N6229);
buf BUF1 (N9942, N9925);
buf BUF1 (N9943, N9929);
buf BUF1 (N9944, N9941);
and AND4 (N9945, N9938, N1347, N5233, N2282);
and AND2 (N9946, N9943, N5382);
buf BUF1 (N9947, N9923);
nor NOR4 (N9948, N9939, N9700, N196, N6919);
not NOT1 (N9949, N9942);
or OR2 (N9950, N9948, N6728);
or OR2 (N9951, N9947, N9692);
or OR2 (N9952, N9945, N7438);
xor XOR2 (N9953, N9914, N4574);
xor XOR2 (N9954, N9944, N7327);
nor NOR3 (N9955, N9952, N3766, N3115);
buf BUF1 (N9956, N9951);
xor XOR2 (N9957, N9946, N6025);
and AND4 (N9958, N9953, N8435, N8458, N1797);
or OR2 (N9959, N9955, N4235);
nand NAND3 (N9960, N9950, N6237, N3330);
nor NOR4 (N9961, N9940, N6658, N7959, N9007);
buf BUF1 (N9962, N9937);
and AND3 (N9963, N9956, N850, N4325);
xor XOR2 (N9964, N9962, N7522);
nand NAND3 (N9965, N9957, N6177, N853);
xor XOR2 (N9966, N9954, N6215);
buf BUF1 (N9967, N9959);
xor XOR2 (N9968, N9964, N7601);
or OR2 (N9969, N9961, N5133);
buf BUF1 (N9970, N9968);
nor NOR4 (N9971, N9935, N7369, N7156, N1508);
xor XOR2 (N9972, N9949, N6009);
nand NAND3 (N9973, N9971, N4370, N3031);
buf BUF1 (N9974, N9973);
buf BUF1 (N9975, N9958);
xor XOR2 (N9976, N9975, N78);
nor NOR3 (N9977, N9960, N8892, N397);
xor XOR2 (N9978, N9969, N8446);
or OR4 (N9979, N9977, N258, N4317, N9593);
buf BUF1 (N9980, N9963);
buf BUF1 (N9981, N9972);
and AND3 (N9982, N9980, N2639, N3006);
nand NAND3 (N9983, N9967, N7867, N3760);
and AND4 (N9984, N9970, N9304, N2739, N2696);
not NOT1 (N9985, N9979);
nor NOR2 (N9986, N9985, N6935);
and AND2 (N9987, N9981, N5738);
nor NOR3 (N9988, N9978, N8977, N5450);
or OR4 (N9989, N9966, N7068, N8793, N125);
nor NOR4 (N9990, N9986, N1952, N7301, N4246);
nand NAND4 (N9991, N9984, N6053, N7222, N3241);
nand NAND2 (N9992, N9990, N3847);
xor XOR2 (N9993, N9992, N4580);
nand NAND4 (N9994, N9982, N5652, N6457, N6550);
nor NOR2 (N9995, N9988, N2055);
nor NOR4 (N9996, N9965, N9939, N1001, N13);
nand NAND4 (N9997, N9974, N3601, N3294, N4679);
xor XOR2 (N9998, N9989, N5167);
or OR3 (N9999, N9976, N616, N5947);
xor XOR2 (N10000, N9998, N9117);
xor XOR2 (N10001, N10000, N8660);
buf BUF1 (N10002, N10001);
not NOT1 (N10003, N9983);
nand NAND4 (N10004, N9997, N7342, N901, N8892);
xor XOR2 (N10005, N9987, N9693);
and AND2 (N10006, N10005, N3442);
xor XOR2 (N10007, N9999, N2383);
xor XOR2 (N10008, N10006, N6608);
buf BUF1 (N10009, N9991);
not NOT1 (N10010, N10008);
xor XOR2 (N10011, N9994, N6191);
and AND4 (N10012, N9996, N7763, N3567, N524);
nand NAND2 (N10013, N10011, N5457);
buf BUF1 (N10014, N10002);
and AND2 (N10015, N10013, N5544);
xor XOR2 (N10016, N10010, N5301);
not NOT1 (N10017, N9995);
or OR4 (N10018, N10004, N1893, N6159, N7872);
nand NAND2 (N10019, N9993, N4891);
not NOT1 (N10020, N10012);
not NOT1 (N10021, N10003);
xor XOR2 (N10022, N10015, N3963);
xor XOR2 (N10023, N10007, N7412);
nand NAND2 (N10024, N10014, N1049);
not NOT1 (N10025, N10020);
nor NOR3 (N10026, N10024, N5063, N4763);
or OR3 (N10027, N10009, N4494, N7687);
nand NAND4 (N10028, N10027, N690, N4828, N92);
nor NOR4 (N10029, N10025, N8292, N6003, N723);
nor NOR4 (N10030, N10026, N3233, N8999, N1266);
or OR4 (N10031, N10017, N8354, N392, N4104);
not NOT1 (N10032, N10016);
or OR4 (N10033, N10022, N6092, N3700, N6004);
not NOT1 (N10034, N10028);
not NOT1 (N10035, N10032);
buf BUF1 (N10036, N10031);
buf BUF1 (N10037, N10023);
buf BUF1 (N10038, N10034);
or OR3 (N10039, N10038, N6617, N1882);
or OR4 (N10040, N10036, N1784, N3246, N1796);
and AND3 (N10041, N10019, N6445, N1438);
buf BUF1 (N10042, N10037);
and AND4 (N10043, N10035, N1221, N7226, N4239);
not NOT1 (N10044, N10039);
nand NAND3 (N10045, N10041, N3705, N1519);
buf BUF1 (N10046, N10040);
buf BUF1 (N10047, N10030);
and AND2 (N10048, N10033, N1089);
nand NAND4 (N10049, N10047, N8119, N3215, N3507);
xor XOR2 (N10050, N10018, N763);
and AND4 (N10051, N10042, N1740, N8173, N7295);
nand NAND2 (N10052, N10043, N860);
and AND4 (N10053, N10046, N8456, N101, N4424);
nand NAND2 (N10054, N10044, N3594);
xor XOR2 (N10055, N10045, N3966);
or OR2 (N10056, N10050, N5747);
buf BUF1 (N10057, N10029);
or OR3 (N10058, N10049, N2753, N6507);
or OR3 (N10059, N10054, N6303, N9600);
xor XOR2 (N10060, N10051, N3940);
nor NOR4 (N10061, N10052, N6406, N3568, N1043);
nand NAND4 (N10062, N10058, N2642, N946, N5394);
xor XOR2 (N10063, N10053, N3676);
and AND3 (N10064, N10021, N3695, N8668);
not NOT1 (N10065, N10056);
nand NAND4 (N10066, N10064, N5226, N1370, N8988);
and AND2 (N10067, N10066, N4142);
xor XOR2 (N10068, N10060, N1009);
nor NOR3 (N10069, N10059, N6862, N6851);
not NOT1 (N10070, N10068);
nor NOR3 (N10071, N10048, N1127, N8987);
or OR2 (N10072, N10069, N7968);
and AND4 (N10073, N10055, N4395, N9999, N3259);
buf BUF1 (N10074, N10067);
buf BUF1 (N10075, N10065);
xor XOR2 (N10076, N10074, N4577);
nor NOR3 (N10077, N10073, N1173, N726);
buf BUF1 (N10078, N10057);
nand NAND4 (N10079, N10077, N3744, N9483, N8900);
nor NOR2 (N10080, N10061, N9869);
and AND2 (N10081, N10076, N8416);
and AND3 (N10082, N10062, N7978, N327);
nand NAND4 (N10083, N10080, N1950, N8471, N1697);
nand NAND3 (N10084, N10063, N3334, N7437);
or OR2 (N10085, N10082, N2423);
and AND3 (N10086, N10071, N3733, N93);
xor XOR2 (N10087, N10072, N1734);
buf BUF1 (N10088, N10081);
xor XOR2 (N10089, N10085, N5696);
and AND3 (N10090, N10087, N6603, N503);
xor XOR2 (N10091, N10084, N443);
or OR2 (N10092, N10083, N5650);
buf BUF1 (N10093, N10079);
buf BUF1 (N10094, N10091);
xor XOR2 (N10095, N10075, N6967);
not NOT1 (N10096, N10095);
nor NOR4 (N10097, N10090, N3033, N6220, N8631);
xor XOR2 (N10098, N10078, N3164);
not NOT1 (N10099, N10088);
xor XOR2 (N10100, N10086, N6141);
buf BUF1 (N10101, N10099);
nor NOR2 (N10102, N10070, N3750);
not NOT1 (N10103, N10096);
and AND2 (N10104, N10093, N1194);
not NOT1 (N10105, N10100);
xor XOR2 (N10106, N10101, N5378);
and AND2 (N10107, N10094, N730);
or OR2 (N10108, N10107, N1754);
buf BUF1 (N10109, N10089);
xor XOR2 (N10110, N10098, N4565);
xor XOR2 (N10111, N10105, N9013);
nand NAND2 (N10112, N10108, N7411);
not NOT1 (N10113, N10110);
nor NOR2 (N10114, N10109, N5610);
xor XOR2 (N10115, N10111, N2038);
buf BUF1 (N10116, N10103);
xor XOR2 (N10117, N10116, N9631);
nor NOR3 (N10118, N10092, N6810, N5223);
nor NOR3 (N10119, N10114, N6048, N1050);
and AND2 (N10120, N10113, N4725);
not NOT1 (N10121, N10112);
xor XOR2 (N10122, N10120, N4183);
nor NOR2 (N10123, N10104, N3360);
nor NOR3 (N10124, N10115, N952, N8253);
nand NAND2 (N10125, N10106, N6034);
and AND2 (N10126, N10125, N319);
nor NOR4 (N10127, N10117, N7577, N8573, N8157);
buf BUF1 (N10128, N10118);
nand NAND4 (N10129, N10124, N9330, N5399, N9402);
buf BUF1 (N10130, N10119);
xor XOR2 (N10131, N10127, N2710);
buf BUF1 (N10132, N10126);
nor NOR2 (N10133, N10102, N903);
nand NAND3 (N10134, N10097, N6498, N5535);
xor XOR2 (N10135, N10130, N6237);
nand NAND3 (N10136, N10123, N1502, N4446);
or OR2 (N10137, N10131, N4404);
nor NOR3 (N10138, N10134, N3401, N462);
buf BUF1 (N10139, N10121);
xor XOR2 (N10140, N10138, N6574);
and AND3 (N10141, N10139, N5801, N3747);
not NOT1 (N10142, N10136);
nand NAND2 (N10143, N10132, N1547);
not NOT1 (N10144, N10137);
and AND2 (N10145, N10135, N4640);
xor XOR2 (N10146, N10128, N6108);
not NOT1 (N10147, N10144);
or OR4 (N10148, N10142, N7986, N2974, N230);
or OR4 (N10149, N10148, N4474, N1880, N5437);
not NOT1 (N10150, N10145);
xor XOR2 (N10151, N10146, N9557);
not NOT1 (N10152, N10122);
xor XOR2 (N10153, N10149, N4930);
buf BUF1 (N10154, N10151);
and AND4 (N10155, N10154, N8616, N9675, N6501);
and AND4 (N10156, N10147, N3055, N6836, N2075);
or OR3 (N10157, N10156, N8527, N10141);
nand NAND3 (N10158, N6653, N8594, N973);
nor NOR2 (N10159, N10158, N2412);
nand NAND3 (N10160, N10159, N9736, N835);
and AND4 (N10161, N10160, N3418, N893, N5992);
buf BUF1 (N10162, N10150);
and AND4 (N10163, N10155, N9008, N5430, N2467);
nand NAND2 (N10164, N10162, N6304);
not NOT1 (N10165, N10152);
nand NAND3 (N10166, N10133, N8204, N3296);
xor XOR2 (N10167, N10163, N8914);
buf BUF1 (N10168, N10153);
and AND2 (N10169, N10157, N5307);
nand NAND4 (N10170, N10143, N3732, N7236, N9542);
buf BUF1 (N10171, N10161);
or OR2 (N10172, N10171, N2546);
or OR2 (N10173, N10129, N6033);
xor XOR2 (N10174, N10168, N7291);
nand NAND4 (N10175, N10164, N6308, N1860, N3342);
nor NOR2 (N10176, N10175, N2347);
buf BUF1 (N10177, N10169);
buf BUF1 (N10178, N10167);
nand NAND4 (N10179, N10173, N9720, N9211, N9776);
and AND2 (N10180, N10177, N1968);
and AND4 (N10181, N10170, N5550, N622, N8644);
or OR3 (N10182, N10181, N8293, N3615);
not NOT1 (N10183, N10174);
nor NOR3 (N10184, N10179, N6985, N6292);
buf BUF1 (N10185, N10183);
nor NOR3 (N10186, N10182, N7681, N434);
buf BUF1 (N10187, N10184);
nor NOR3 (N10188, N10185, N6121, N5703);
nand NAND2 (N10189, N10186, N1151);
xor XOR2 (N10190, N10187, N5016);
or OR3 (N10191, N10190, N452, N5270);
nand NAND2 (N10192, N10189, N3460);
nor NOR2 (N10193, N10140, N9170);
or OR3 (N10194, N10176, N2742, N6151);
and AND4 (N10195, N10166, N2831, N6689, N5998);
or OR2 (N10196, N10165, N9053);
and AND4 (N10197, N10172, N10166, N2141, N6678);
and AND2 (N10198, N10193, N8963);
or OR2 (N10199, N10180, N1481);
xor XOR2 (N10200, N10197, N4809);
buf BUF1 (N10201, N10200);
nor NOR3 (N10202, N10201, N4038, N10019);
or OR3 (N10203, N10188, N2679, N2525);
xor XOR2 (N10204, N10192, N8182);
nor NOR4 (N10205, N10199, N9073, N2340, N4769);
buf BUF1 (N10206, N10195);
nand NAND2 (N10207, N10206, N5150);
not NOT1 (N10208, N10204);
xor XOR2 (N10209, N10208, N8047);
buf BUF1 (N10210, N10194);
buf BUF1 (N10211, N10191);
nor NOR3 (N10212, N10207, N3275, N7538);
and AND4 (N10213, N10178, N10205, N8386, N7219);
or OR4 (N10214, N8084, N6589, N1988, N1508);
or OR4 (N10215, N10210, N6634, N8624, N811);
nor NOR4 (N10216, N10196, N432, N2661, N1333);
or OR4 (N10217, N10198, N3582, N9226, N3469);
not NOT1 (N10218, N10215);
nor NOR2 (N10219, N10214, N4489);
buf BUF1 (N10220, N10217);
or OR2 (N10221, N10213, N7723);
nand NAND2 (N10222, N10203, N1166);
not NOT1 (N10223, N10202);
nor NOR2 (N10224, N10223, N4801);
xor XOR2 (N10225, N10212, N9179);
nor NOR4 (N10226, N10209, N1081, N5851, N10074);
or OR2 (N10227, N10222, N4863);
nand NAND3 (N10228, N10227, N6250, N9021);
xor XOR2 (N10229, N10228, N862);
buf BUF1 (N10230, N10218);
nand NAND4 (N10231, N10211, N6776, N8478, N7672);
xor XOR2 (N10232, N10226, N3401);
xor XOR2 (N10233, N10220, N2500);
not NOT1 (N10234, N10233);
not NOT1 (N10235, N10216);
not NOT1 (N10236, N10221);
nor NOR3 (N10237, N10235, N4015, N2886);
nor NOR2 (N10238, N10232, N485);
xor XOR2 (N10239, N10219, N3639);
not NOT1 (N10240, N10237);
nand NAND4 (N10241, N10224, N1875, N9165, N2341);
not NOT1 (N10242, N10234);
buf BUF1 (N10243, N10242);
and AND4 (N10244, N10236, N3039, N9985, N2804);
nand NAND4 (N10245, N10243, N1462, N8221, N1843);
or OR2 (N10246, N10241, N1056);
xor XOR2 (N10247, N10238, N5813);
xor XOR2 (N10248, N10231, N8867);
nand NAND3 (N10249, N10239, N9653, N9784);
not NOT1 (N10250, N10230);
buf BUF1 (N10251, N10249);
buf BUF1 (N10252, N10251);
nand NAND4 (N10253, N10245, N7124, N2217, N881);
or OR4 (N10254, N10240, N4510, N3276, N2632);
not NOT1 (N10255, N10229);
not NOT1 (N10256, N10254);
and AND2 (N10257, N10247, N1945);
buf BUF1 (N10258, N10250);
xor XOR2 (N10259, N10255, N1656);
nand NAND3 (N10260, N10225, N7136, N948);
or OR2 (N10261, N10252, N6601);
xor XOR2 (N10262, N10256, N5453);
buf BUF1 (N10263, N10246);
xor XOR2 (N10264, N10258, N2612);
and AND4 (N10265, N10263, N6819, N8036, N8597);
nor NOR4 (N10266, N10265, N7671, N3247, N2054);
and AND4 (N10267, N10248, N5763, N57, N7244);
not NOT1 (N10268, N10264);
xor XOR2 (N10269, N10244, N2577);
nand NAND4 (N10270, N10253, N3368, N2282, N492);
nor NOR2 (N10271, N10269, N3346);
nor NOR4 (N10272, N10260, N5810, N5778, N194);
nor NOR3 (N10273, N10270, N6607, N9181);
and AND4 (N10274, N10262, N9315, N4327, N4184);
not NOT1 (N10275, N10273);
buf BUF1 (N10276, N10261);
buf BUF1 (N10277, N10276);
not NOT1 (N10278, N10272);
xor XOR2 (N10279, N10259, N8289);
buf BUF1 (N10280, N10277);
not NOT1 (N10281, N10279);
and AND2 (N10282, N10275, N4684);
and AND2 (N10283, N10282, N5526);
xor XOR2 (N10284, N10283, N140);
nand NAND4 (N10285, N10284, N9878, N7807, N5741);
xor XOR2 (N10286, N10257, N7064);
not NOT1 (N10287, N10278);
or OR3 (N10288, N10274, N1066, N9360);
nand NAND3 (N10289, N10281, N888, N6227);
or OR2 (N10290, N10285, N2438);
not NOT1 (N10291, N10289);
buf BUF1 (N10292, N10290);
nand NAND2 (N10293, N10291, N2855);
nand NAND2 (N10294, N10266, N90);
nor NOR4 (N10295, N10268, N791, N1177, N9193);
or OR4 (N10296, N10295, N9374, N7933, N9863);
xor XOR2 (N10297, N10296, N174);
nand NAND3 (N10298, N10292, N907, N5467);
and AND2 (N10299, N10288, N8426);
or OR4 (N10300, N10297, N9257, N2677, N4498);
buf BUF1 (N10301, N10300);
buf BUF1 (N10302, N10294);
buf BUF1 (N10303, N10287);
buf BUF1 (N10304, N10303);
not NOT1 (N10305, N10271);
or OR2 (N10306, N10304, N7686);
or OR3 (N10307, N10293, N1794, N2458);
and AND4 (N10308, N10306, N6943, N9347, N5829);
and AND3 (N10309, N10280, N9013, N1184);
nor NOR3 (N10310, N10305, N4252, N2971);
nor NOR2 (N10311, N10309, N10086);
nor NOR2 (N10312, N10308, N4404);
not NOT1 (N10313, N10301);
and AND4 (N10314, N10313, N101, N1854, N1048);
and AND3 (N10315, N10298, N7392, N7067);
or OR2 (N10316, N10315, N1584);
buf BUF1 (N10317, N10310);
not NOT1 (N10318, N10311);
not NOT1 (N10319, N10302);
nor NOR3 (N10320, N10307, N7523, N9464);
xor XOR2 (N10321, N10314, N7702);
or OR2 (N10322, N10286, N9683);
and AND2 (N10323, N10321, N9453);
nand NAND3 (N10324, N10312, N9784, N8001);
buf BUF1 (N10325, N10317);
nand NAND2 (N10326, N10267, N7217);
and AND3 (N10327, N10320, N8238, N8159);
nand NAND3 (N10328, N10316, N580, N4664);
nor NOR2 (N10329, N10323, N5821);
and AND4 (N10330, N10299, N1986, N5184, N9915);
nor NOR2 (N10331, N10330, N8268);
and AND4 (N10332, N10328, N3393, N8570, N2560);
xor XOR2 (N10333, N10331, N4403);
buf BUF1 (N10334, N10333);
nand NAND3 (N10335, N10327, N5622, N2836);
buf BUF1 (N10336, N10322);
and AND3 (N10337, N10332, N9114, N5995);
nand NAND2 (N10338, N10334, N895);
not NOT1 (N10339, N10318);
xor XOR2 (N10340, N10326, N10064);
nor NOR2 (N10341, N10340, N1036);
xor XOR2 (N10342, N10324, N6117);
nand NAND2 (N10343, N10337, N5442);
nor NOR3 (N10344, N10338, N2708, N2107);
not NOT1 (N10345, N10341);
and AND2 (N10346, N10343, N6234);
buf BUF1 (N10347, N10336);
nor NOR3 (N10348, N10346, N5064, N8407);
or OR4 (N10349, N10329, N6427, N5783, N695);
or OR4 (N10350, N10335, N8369, N1910, N3912);
nor NOR3 (N10351, N10342, N6935, N2368);
not NOT1 (N10352, N10325);
nor NOR3 (N10353, N10348, N7304, N5731);
not NOT1 (N10354, N10349);
and AND3 (N10355, N10354, N1943, N9845);
buf BUF1 (N10356, N10345);
nand NAND2 (N10357, N10352, N2219);
buf BUF1 (N10358, N10339);
nor NOR3 (N10359, N10344, N6181, N6056);
buf BUF1 (N10360, N10351);
nor NOR2 (N10361, N10353, N5481);
buf BUF1 (N10362, N10319);
or OR4 (N10363, N10356, N8235, N9373, N3116);
nand NAND2 (N10364, N10347, N1793);
or OR2 (N10365, N10362, N10207);
buf BUF1 (N10366, N10365);
or OR2 (N10367, N10358, N1859);
xor XOR2 (N10368, N10357, N9475);
not NOT1 (N10369, N10364);
or OR2 (N10370, N10350, N5584);
or OR2 (N10371, N10360, N6094);
or OR2 (N10372, N10361, N3521);
buf BUF1 (N10373, N10369);
or OR2 (N10374, N10366, N1321);
buf BUF1 (N10375, N10355);
buf BUF1 (N10376, N10371);
and AND2 (N10377, N10359, N8893);
nand NAND4 (N10378, N10375, N2398, N2668, N10359);
nor NOR2 (N10379, N10370, N4753);
nand NAND2 (N10380, N10378, N6454);
or OR2 (N10381, N10368, N2999);
nand NAND2 (N10382, N10380, N2016);
not NOT1 (N10383, N10377);
nand NAND2 (N10384, N10373, N371);
xor XOR2 (N10385, N10374, N10382);
not NOT1 (N10386, N3786);
nand NAND2 (N10387, N10383, N2145);
xor XOR2 (N10388, N10372, N3526);
nor NOR3 (N10389, N10363, N1742, N6922);
buf BUF1 (N10390, N10381);
buf BUF1 (N10391, N10389);
and AND3 (N10392, N10387, N7480, N6690);
nand NAND4 (N10393, N10379, N3564, N6285, N8433);
nand NAND3 (N10394, N10386, N2327, N4014);
buf BUF1 (N10395, N10384);
xor XOR2 (N10396, N10391, N4898);
or OR3 (N10397, N10394, N7943, N3716);
nor NOR4 (N10398, N10392, N3336, N2363, N8461);
or OR3 (N10399, N10367, N2908, N4552);
or OR4 (N10400, N10397, N6802, N3909, N1754);
or OR4 (N10401, N10396, N1286, N1518, N6745);
not NOT1 (N10402, N10395);
or OR3 (N10403, N10398, N4090, N3558);
and AND3 (N10404, N10399, N871, N9709);
buf BUF1 (N10405, N10385);
nor NOR3 (N10406, N10402, N3694, N654);
not NOT1 (N10407, N10388);
or OR3 (N10408, N10401, N10314, N4823);
nand NAND3 (N10409, N10406, N1390, N4553);
not NOT1 (N10410, N10376);
nor NOR3 (N10411, N10410, N8477, N3767);
not NOT1 (N10412, N10408);
xor XOR2 (N10413, N10412, N3540);
xor XOR2 (N10414, N10413, N10281);
and AND2 (N10415, N10404, N6227);
or OR4 (N10416, N10400, N800, N10017, N6363);
nor NOR3 (N10417, N10403, N4797, N9033);
buf BUF1 (N10418, N10415);
buf BUF1 (N10419, N10407);
not NOT1 (N10420, N10419);
xor XOR2 (N10421, N10418, N3971);
nand NAND4 (N10422, N10417, N8741, N8169, N5011);
xor XOR2 (N10423, N10420, N6016);
not NOT1 (N10424, N10390);
nor NOR4 (N10425, N10411, N1787, N5552, N8704);
xor XOR2 (N10426, N10422, N10145);
nand NAND2 (N10427, N10425, N8905);
buf BUF1 (N10428, N10414);
nand NAND4 (N10429, N10416, N4947, N6484, N1384);
xor XOR2 (N10430, N10429, N4329);
not NOT1 (N10431, N10423);
nor NOR4 (N10432, N10431, N5137, N9804, N6695);
or OR4 (N10433, N10424, N5221, N6507, N544);
nand NAND2 (N10434, N10432, N7215);
or OR2 (N10435, N10421, N10078);
nand NAND3 (N10436, N10426, N10183, N6850);
nor NOR4 (N10437, N10436, N9529, N8326, N9433);
nor NOR3 (N10438, N10427, N4831, N7521);
or OR4 (N10439, N10433, N3007, N1606, N6198);
not NOT1 (N10440, N10434);
xor XOR2 (N10441, N10438, N4748);
nand NAND4 (N10442, N10393, N6117, N8645, N7166);
xor XOR2 (N10443, N10435, N1968);
nor NOR3 (N10444, N10409, N5627, N8189);
or OR3 (N10445, N10443, N3797, N91);
xor XOR2 (N10446, N10442, N1663);
and AND3 (N10447, N10439, N720, N3828);
and AND3 (N10448, N10437, N425, N4373);
nand NAND3 (N10449, N10430, N8130, N5549);
nor NOR2 (N10450, N10405, N160);
nand NAND3 (N10451, N10446, N2183, N5550);
and AND3 (N10452, N10440, N4498, N10350);
or OR3 (N10453, N10451, N401, N4221);
and AND3 (N10454, N10452, N9977, N3996);
not NOT1 (N10455, N10428);
nor NOR4 (N10456, N10449, N6397, N8709, N9486);
buf BUF1 (N10457, N10455);
nand NAND2 (N10458, N10441, N4039);
not NOT1 (N10459, N10456);
nand NAND2 (N10460, N10447, N10174);
buf BUF1 (N10461, N10448);
nand NAND4 (N10462, N10457, N4285, N793, N4432);
not NOT1 (N10463, N10459);
nand NAND3 (N10464, N10463, N4439, N2559);
buf BUF1 (N10465, N10461);
nor NOR4 (N10466, N10445, N8082, N5191, N2572);
and AND3 (N10467, N10458, N2299, N382);
buf BUF1 (N10468, N10465);
and AND2 (N10469, N10468, N4805);
xor XOR2 (N10470, N10460, N3603);
nor NOR3 (N10471, N10453, N7863, N1502);
and AND3 (N10472, N10469, N8228, N9544);
nand NAND4 (N10473, N10466, N8326, N1372, N304);
and AND4 (N10474, N10444, N9097, N7399, N823);
or OR3 (N10475, N10464, N4609, N912);
nand NAND3 (N10476, N10474, N2339, N5437);
nor NOR4 (N10477, N10472, N8143, N2379, N10067);
buf BUF1 (N10478, N10454);
nand NAND3 (N10479, N10462, N1881, N4769);
nor NOR3 (N10480, N10476, N7020, N9752);
nor NOR4 (N10481, N10478, N3961, N5409, N8339);
not NOT1 (N10482, N10477);
nand NAND4 (N10483, N10482, N8110, N144, N2653);
nand NAND2 (N10484, N10467, N8249);
not NOT1 (N10485, N10479);
nor NOR4 (N10486, N10473, N5168, N10091, N8557);
not NOT1 (N10487, N10483);
or OR4 (N10488, N10481, N1603, N2366, N9554);
or OR4 (N10489, N10470, N1265, N7238, N5558);
or OR2 (N10490, N10485, N4052);
or OR3 (N10491, N10471, N9950, N7210);
and AND3 (N10492, N10488, N4153, N5562);
xor XOR2 (N10493, N10484, N3733);
and AND4 (N10494, N10492, N5433, N8318, N10075);
nand NAND4 (N10495, N10490, N6621, N9595, N568);
or OR4 (N10496, N10480, N6894, N9673, N2403);
buf BUF1 (N10497, N10495);
not NOT1 (N10498, N10497);
nor NOR3 (N10499, N10487, N8482, N8818);
nand NAND4 (N10500, N10486, N2219, N3116, N2216);
and AND3 (N10501, N10494, N9270, N4921);
nand NAND4 (N10502, N10450, N7053, N9350, N1013);
and AND3 (N10503, N10498, N1828, N3681);
and AND3 (N10504, N10491, N419, N6846);
nand NAND3 (N10505, N10496, N509, N9923);
nor NOR2 (N10506, N10475, N5080);
xor XOR2 (N10507, N10501, N108);
and AND3 (N10508, N10504, N7549, N994);
and AND4 (N10509, N10500, N7124, N7633, N3794);
or OR4 (N10510, N10502, N1997, N2026, N321);
or OR3 (N10511, N10503, N729, N512);
nor NOR4 (N10512, N10506, N584, N4252, N238);
buf BUF1 (N10513, N10512);
and AND2 (N10514, N10493, N2140);
nand NAND4 (N10515, N10505, N4752, N2602, N4194);
nor NOR3 (N10516, N10511, N2295, N5922);
buf BUF1 (N10517, N10510);
and AND2 (N10518, N10516, N5835);
and AND2 (N10519, N10489, N4569);
nor NOR4 (N10520, N10509, N5961, N5541, N2240);
and AND3 (N10521, N10513, N10232, N7099);
nand NAND3 (N10522, N10518, N9084, N6621);
buf BUF1 (N10523, N10499);
buf BUF1 (N10524, N10514);
xor XOR2 (N10525, N10523, N7899);
xor XOR2 (N10526, N10515, N675);
nor NOR4 (N10527, N10525, N10392, N6473, N8447);
and AND3 (N10528, N10517, N9451, N6126);
nor NOR3 (N10529, N10524, N3269, N1707);
xor XOR2 (N10530, N10520, N4040);
nor NOR3 (N10531, N10508, N2540, N9227);
buf BUF1 (N10532, N10528);
xor XOR2 (N10533, N10529, N611);
not NOT1 (N10534, N10531);
nor NOR2 (N10535, N10507, N4778);
nand NAND4 (N10536, N10535, N9395, N2016, N6566);
not NOT1 (N10537, N10536);
not NOT1 (N10538, N10521);
buf BUF1 (N10539, N10519);
buf BUF1 (N10540, N10530);
not NOT1 (N10541, N10538);
and AND4 (N10542, N10532, N600, N3734, N9637);
buf BUF1 (N10543, N10522);
xor XOR2 (N10544, N10533, N8770);
buf BUF1 (N10545, N10527);
nor NOR3 (N10546, N10537, N4652, N7155);
buf BUF1 (N10547, N10545);
xor XOR2 (N10548, N10534, N9859);
nor NOR4 (N10549, N10541, N7839, N9911, N1541);
or OR3 (N10550, N10539, N8405, N8676);
nor NOR3 (N10551, N10540, N10372, N2594);
not NOT1 (N10552, N10550);
and AND3 (N10553, N10548, N7206, N5922);
buf BUF1 (N10554, N10552);
nor NOR4 (N10555, N10542, N10097, N5529, N10346);
not NOT1 (N10556, N10547);
xor XOR2 (N10557, N10551, N1942);
not NOT1 (N10558, N10549);
nor NOR4 (N10559, N10554, N2851, N8445, N7163);
nor NOR4 (N10560, N10559, N2536, N3302, N9495);
and AND4 (N10561, N10553, N996, N1620, N9179);
and AND4 (N10562, N10560, N1486, N6705, N443);
or OR2 (N10563, N10557, N4944);
nor NOR4 (N10564, N10526, N8999, N8526, N6721);
buf BUF1 (N10565, N10564);
buf BUF1 (N10566, N10544);
and AND2 (N10567, N10543, N7865);
nor NOR3 (N10568, N10558, N2541, N5008);
not NOT1 (N10569, N10555);
xor XOR2 (N10570, N10566, N8766);
or OR3 (N10571, N10570, N9046, N4032);
xor XOR2 (N10572, N10561, N2430);
buf BUF1 (N10573, N10568);
xor XOR2 (N10574, N10567, N1849);
buf BUF1 (N10575, N10563);
or OR3 (N10576, N10546, N1848, N9773);
not NOT1 (N10577, N10576);
xor XOR2 (N10578, N10575, N3625);
and AND4 (N10579, N10569, N10244, N5856, N8850);
not NOT1 (N10580, N10562);
nand NAND2 (N10581, N10579, N7806);
nor NOR3 (N10582, N10578, N1229, N7401);
xor XOR2 (N10583, N10571, N7318);
nand NAND4 (N10584, N10580, N88, N7607, N584);
nand NAND4 (N10585, N10577, N4926, N10339, N1108);
or OR4 (N10586, N10572, N9048, N9305, N10112);
or OR4 (N10587, N10565, N9561, N619, N10119);
and AND4 (N10588, N10586, N9942, N1581, N9750);
or OR3 (N10589, N10581, N7798, N6240);
nand NAND4 (N10590, N10582, N7024, N4953, N7949);
and AND4 (N10591, N10574, N1407, N10083, N6440);
not NOT1 (N10592, N10583);
not NOT1 (N10593, N10556);
and AND3 (N10594, N10573, N9380, N1175);
or OR3 (N10595, N10585, N5413, N1300);
not NOT1 (N10596, N10590);
buf BUF1 (N10597, N10584);
xor XOR2 (N10598, N10595, N3339);
buf BUF1 (N10599, N10588);
nor NOR4 (N10600, N10599, N236, N3648, N10060);
xor XOR2 (N10601, N10597, N5841);
not NOT1 (N10602, N10596);
or OR4 (N10603, N10587, N8497, N3113, N3466);
nor NOR2 (N10604, N10602, N5298);
xor XOR2 (N10605, N10593, N3359);
or OR4 (N10606, N10600, N9062, N6156, N3167);
and AND3 (N10607, N10604, N4929, N3045);
xor XOR2 (N10608, N10589, N2703);
nand NAND2 (N10609, N10594, N702);
nand NAND4 (N10610, N10606, N46, N5638, N2691);
nand NAND4 (N10611, N10591, N9370, N6568, N7891);
or OR2 (N10612, N10607, N4094);
not NOT1 (N10613, N10598);
or OR4 (N10614, N10613, N1411, N8100, N9453);
xor XOR2 (N10615, N10608, N4931);
and AND2 (N10616, N10592, N4006);
nand NAND2 (N10617, N10615, N2659);
and AND3 (N10618, N10601, N4629, N26);
xor XOR2 (N10619, N10614, N2421);
buf BUF1 (N10620, N10619);
and AND2 (N10621, N10620, N3679);
nand NAND4 (N10622, N10610, N9097, N566, N4997);
not NOT1 (N10623, N10611);
buf BUF1 (N10624, N10605);
xor XOR2 (N10625, N10609, N2137);
buf BUF1 (N10626, N10623);
not NOT1 (N10627, N10616);
buf BUF1 (N10628, N10627);
not NOT1 (N10629, N10603);
not NOT1 (N10630, N10612);
nor NOR2 (N10631, N10621, N6387);
nand NAND2 (N10632, N10631, N1851);
buf BUF1 (N10633, N10629);
xor XOR2 (N10634, N10632, N858);
or OR2 (N10635, N10617, N10397);
buf BUF1 (N10636, N10618);
buf BUF1 (N10637, N10622);
and AND2 (N10638, N10628, N9177);
buf BUF1 (N10639, N10635);
or OR3 (N10640, N10638, N9190, N3951);
xor XOR2 (N10641, N10624, N293);
and AND2 (N10642, N10639, N14);
and AND2 (N10643, N10640, N8944);
and AND3 (N10644, N10630, N2375, N6289);
xor XOR2 (N10645, N10626, N7937);
nor NOR4 (N10646, N10641, N3424, N3168, N9485);
or OR3 (N10647, N10634, N5405, N6284);
nor NOR4 (N10648, N10633, N4291, N8312, N4189);
and AND3 (N10649, N10637, N7090, N5228);
nand NAND4 (N10650, N10625, N4871, N1770, N9804);
buf BUF1 (N10651, N10647);
nand NAND3 (N10652, N10643, N2085, N4615);
not NOT1 (N10653, N10651);
not NOT1 (N10654, N10650);
buf BUF1 (N10655, N10646);
nor NOR4 (N10656, N10655, N5376, N5325, N8588);
nand NAND3 (N10657, N10654, N10313, N3774);
buf BUF1 (N10658, N10648);
nand NAND2 (N10659, N10636, N10045);
xor XOR2 (N10660, N10657, N1529);
nor NOR3 (N10661, N10659, N3146, N4444);
not NOT1 (N10662, N10642);
nand NAND2 (N10663, N10661, N9043);
nor NOR3 (N10664, N10652, N7189, N4357);
nor NOR4 (N10665, N10663, N6791, N463, N2917);
or OR3 (N10666, N10656, N61, N2676);
xor XOR2 (N10667, N10645, N2348);
nor NOR2 (N10668, N10664, N7638);
not NOT1 (N10669, N10653);
nor NOR2 (N10670, N10662, N8085);
xor XOR2 (N10671, N10665, N5470);
nor NOR3 (N10672, N10660, N9195, N2295);
and AND3 (N10673, N10669, N229, N4036);
not NOT1 (N10674, N10666);
not NOT1 (N10675, N10658);
or OR3 (N10676, N10667, N5786, N8560);
xor XOR2 (N10677, N10673, N4539);
buf BUF1 (N10678, N10670);
or OR2 (N10679, N10644, N7187);
nor NOR3 (N10680, N10675, N1805, N6078);
nor NOR3 (N10681, N10668, N1250, N3198);
buf BUF1 (N10682, N10674);
buf BUF1 (N10683, N10676);
buf BUF1 (N10684, N10680);
not NOT1 (N10685, N10678);
and AND3 (N10686, N10649, N392, N1824);
and AND3 (N10687, N10681, N2405, N4481);
xor XOR2 (N10688, N10684, N3458);
buf BUF1 (N10689, N10685);
nand NAND4 (N10690, N10687, N3793, N10104, N4568);
not NOT1 (N10691, N10677);
nand NAND4 (N10692, N10689, N6207, N10022, N304);
buf BUF1 (N10693, N10679);
buf BUF1 (N10694, N10693);
nand NAND3 (N10695, N10682, N2808, N5241);
buf BUF1 (N10696, N10694);
and AND2 (N10697, N10688, N136);
nor NOR3 (N10698, N10690, N6135, N338);
nor NOR4 (N10699, N10683, N3914, N5144, N4599);
not NOT1 (N10700, N10699);
xor XOR2 (N10701, N10691, N9112);
nand NAND3 (N10702, N10692, N1579, N3294);
buf BUF1 (N10703, N10702);
xor XOR2 (N10704, N10672, N1971);
not NOT1 (N10705, N10700);
nand NAND4 (N10706, N10698, N3764, N1893, N966);
nand NAND2 (N10707, N10704, N3386);
buf BUF1 (N10708, N10686);
buf BUF1 (N10709, N10701);
and AND4 (N10710, N10708, N1097, N6748, N9331);
xor XOR2 (N10711, N10696, N3390);
not NOT1 (N10712, N10707);
nand NAND2 (N10713, N10671, N2059);
xor XOR2 (N10714, N10697, N10462);
not NOT1 (N10715, N10710);
not NOT1 (N10716, N10711);
nand NAND3 (N10717, N10715, N686, N970);
or OR4 (N10718, N10716, N7376, N4864, N739);
and AND2 (N10719, N10703, N5489);
nand NAND2 (N10720, N10705, N9955);
xor XOR2 (N10721, N10695, N6587);
and AND4 (N10722, N10719, N2499, N1602, N9909);
and AND4 (N10723, N10714, N2123, N3089, N9585);
and AND4 (N10724, N10706, N9240, N512, N6678);
buf BUF1 (N10725, N10713);
not NOT1 (N10726, N10721);
nor NOR3 (N10727, N10712, N2842, N5202);
nand NAND3 (N10728, N10724, N5158, N6770);
or OR2 (N10729, N10728, N2141);
nand NAND4 (N10730, N10729, N8219, N2681, N5336);
buf BUF1 (N10731, N10726);
not NOT1 (N10732, N10727);
nor NOR2 (N10733, N10730, N2760);
or OR2 (N10734, N10723, N7737);
nand NAND4 (N10735, N10732, N1437, N893, N8443);
not NOT1 (N10736, N10722);
not NOT1 (N10737, N10725);
or OR4 (N10738, N10720, N6419, N1018, N4182);
xor XOR2 (N10739, N10737, N6683);
nand NAND4 (N10740, N10736, N2627, N4887, N6611);
or OR3 (N10741, N10738, N4801, N3996);
buf BUF1 (N10742, N10733);
nand NAND3 (N10743, N10735, N5775, N9739);
not NOT1 (N10744, N10743);
not NOT1 (N10745, N10742);
and AND3 (N10746, N10718, N8475, N8464);
buf BUF1 (N10747, N10734);
xor XOR2 (N10748, N10740, N3094);
or OR2 (N10749, N10709, N4279);
xor XOR2 (N10750, N10748, N2311);
nand NAND2 (N10751, N10745, N7713);
buf BUF1 (N10752, N10717);
nand NAND3 (N10753, N10731, N4079, N775);
nand NAND2 (N10754, N10752, N5321);
not NOT1 (N10755, N10741);
nand NAND2 (N10756, N10739, N6061);
xor XOR2 (N10757, N10747, N9023);
nor NOR3 (N10758, N10753, N5829, N4765);
and AND3 (N10759, N10755, N2393, N5269);
nor NOR4 (N10760, N10758, N8113, N6426, N8283);
buf BUF1 (N10761, N10749);
nor NOR2 (N10762, N10756, N6895);
buf BUF1 (N10763, N10761);
buf BUF1 (N10764, N10746);
not NOT1 (N10765, N10754);
and AND4 (N10766, N10765, N3605, N3356, N1632);
and AND2 (N10767, N10762, N8957);
buf BUF1 (N10768, N10763);
nor NOR4 (N10769, N10766, N6534, N9142, N2278);
nor NOR4 (N10770, N10751, N1917, N2850, N4061);
xor XOR2 (N10771, N10750, N95);
nor NOR3 (N10772, N10767, N6946, N3121);
xor XOR2 (N10773, N10772, N7924);
xor XOR2 (N10774, N10769, N10718);
or OR4 (N10775, N10760, N7215, N10293, N7971);
buf BUF1 (N10776, N10744);
xor XOR2 (N10777, N10757, N8619);
or OR3 (N10778, N10773, N2892, N10621);
and AND3 (N10779, N10778, N8137, N2818);
xor XOR2 (N10780, N10776, N8959);
nand NAND2 (N10781, N10775, N599);
buf BUF1 (N10782, N10771);
buf BUF1 (N10783, N10768);
nand NAND3 (N10784, N10782, N5578, N2173);
nor NOR3 (N10785, N10780, N1222, N8040);
xor XOR2 (N10786, N10774, N5924);
xor XOR2 (N10787, N10779, N8164);
and AND4 (N10788, N10777, N4482, N245, N2114);
xor XOR2 (N10789, N10784, N6308);
not NOT1 (N10790, N10788);
or OR2 (N10791, N10786, N5147);
nand NAND2 (N10792, N10791, N4891);
not NOT1 (N10793, N10785);
or OR2 (N10794, N10792, N328);
and AND4 (N10795, N10764, N4733, N7630, N5621);
buf BUF1 (N10796, N10790);
or OR3 (N10797, N10783, N1213, N5801);
or OR3 (N10798, N10793, N6305, N8182);
nand NAND4 (N10799, N10759, N120, N5169, N3046);
buf BUF1 (N10800, N10787);
nor NOR2 (N10801, N10770, N2272);
not NOT1 (N10802, N10801);
or OR2 (N10803, N10802, N6534);
buf BUF1 (N10804, N10803);
buf BUF1 (N10805, N10795);
or OR3 (N10806, N10794, N6464, N3820);
xor XOR2 (N10807, N10796, N9852);
nor NOR3 (N10808, N10781, N2995, N5429);
and AND3 (N10809, N10804, N5368, N3003);
nor NOR4 (N10810, N10808, N1825, N8098, N6569);
buf BUF1 (N10811, N10810);
xor XOR2 (N10812, N10807, N660);
nor NOR2 (N10813, N10809, N7699);
buf BUF1 (N10814, N10800);
not NOT1 (N10815, N10813);
or OR4 (N10816, N10806, N928, N5788, N6444);
nand NAND2 (N10817, N10812, N10788);
not NOT1 (N10818, N10799);
not NOT1 (N10819, N10811);
and AND2 (N10820, N10814, N2612);
xor XOR2 (N10821, N10815, N3180);
buf BUF1 (N10822, N10819);
nand NAND2 (N10823, N10822, N6897);
nand NAND4 (N10824, N10817, N9120, N7795, N2383);
xor XOR2 (N10825, N10797, N4804);
or OR2 (N10826, N10818, N5520);
nor NOR2 (N10827, N10821, N1168);
or OR2 (N10828, N10816, N2219);
and AND4 (N10829, N10789, N6415, N6471, N10503);
or OR3 (N10830, N10805, N2297, N5018);
nor NOR3 (N10831, N10798, N1673, N9863);
buf BUF1 (N10832, N10827);
not NOT1 (N10833, N10820);
or OR2 (N10834, N10825, N9234);
nand NAND3 (N10835, N10834, N1417, N1034);
buf BUF1 (N10836, N10835);
xor XOR2 (N10837, N10823, N7838);
not NOT1 (N10838, N10824);
nand NAND2 (N10839, N10831, N9522);
xor XOR2 (N10840, N10839, N3760);
or OR4 (N10841, N10837, N2373, N10382, N1726);
not NOT1 (N10842, N10826);
buf BUF1 (N10843, N10840);
or OR3 (N10844, N10841, N10196, N10671);
buf BUF1 (N10845, N10843);
and AND4 (N10846, N10833, N4751, N7021, N948);
xor XOR2 (N10847, N10832, N2026);
not NOT1 (N10848, N10844);
and AND4 (N10849, N10842, N6053, N8763, N4291);
and AND4 (N10850, N10847, N3074, N6800, N9144);
nand NAND2 (N10851, N10849, N472);
buf BUF1 (N10852, N10836);
xor XOR2 (N10853, N10845, N10024);
nand NAND4 (N10854, N10829, N6714, N5463, N1365);
xor XOR2 (N10855, N10838, N9210);
buf BUF1 (N10856, N10853);
xor XOR2 (N10857, N10851, N5860);
nor NOR2 (N10858, N10854, N8102);
or OR4 (N10859, N10848, N8747, N1523, N10625);
not NOT1 (N10860, N10850);
nand NAND3 (N10861, N10846, N6816, N9627);
xor XOR2 (N10862, N10857, N6114);
not NOT1 (N10863, N10862);
not NOT1 (N10864, N10855);
not NOT1 (N10865, N10864);
nor NOR2 (N10866, N10863, N1404);
xor XOR2 (N10867, N10830, N838);
and AND2 (N10868, N10828, N9019);
xor XOR2 (N10869, N10866, N1203);
nand NAND4 (N10870, N10852, N9388, N7409, N3424);
and AND4 (N10871, N10860, N3849, N8275, N9443);
or OR4 (N10872, N10858, N2391, N8223, N4463);
or OR2 (N10873, N10868, N7191);
not NOT1 (N10874, N10861);
buf BUF1 (N10875, N10867);
not NOT1 (N10876, N10859);
and AND3 (N10877, N10875, N228, N7587);
xor XOR2 (N10878, N10870, N4838);
or OR4 (N10879, N10876, N2246, N10188, N584);
buf BUF1 (N10880, N10856);
xor XOR2 (N10881, N10874, N10512);
nor NOR4 (N10882, N10879, N5390, N6600, N9844);
nand NAND2 (N10883, N10882, N7847);
nor NOR4 (N10884, N10865, N3927, N6091, N9172);
not NOT1 (N10885, N10869);
buf BUF1 (N10886, N10884);
buf BUF1 (N10887, N10886);
nor NOR4 (N10888, N10878, N727, N7052, N8556);
and AND4 (N10889, N10887, N10247, N8568, N7292);
nand NAND3 (N10890, N10881, N7814, N5055);
nor NOR3 (N10891, N10885, N7931, N3036);
and AND3 (N10892, N10890, N8819, N2131);
nor NOR4 (N10893, N10877, N5552, N1004, N6953);
nor NOR3 (N10894, N10893, N1264, N1819);
buf BUF1 (N10895, N10873);
nor NOR3 (N10896, N10883, N8792, N4275);
nand NAND3 (N10897, N10894, N10691, N4264);
and AND4 (N10898, N10888, N5033, N3096, N702);
xor XOR2 (N10899, N10880, N5075);
and AND2 (N10900, N10891, N10591);
nand NAND2 (N10901, N10892, N9336);
nand NAND3 (N10902, N10896, N8139, N4471);
buf BUF1 (N10903, N10902);
not NOT1 (N10904, N10872);
or OR4 (N10905, N10903, N1318, N1136, N1625);
not NOT1 (N10906, N10900);
nand NAND2 (N10907, N10897, N9910);
nor NOR4 (N10908, N10907, N4842, N3362, N2715);
buf BUF1 (N10909, N10895);
buf BUF1 (N10910, N10904);
xor XOR2 (N10911, N10889, N8840);
buf BUF1 (N10912, N10901);
nor NOR2 (N10913, N10909, N9789);
and AND4 (N10914, N10912, N8668, N6123, N1047);
and AND3 (N10915, N10899, N532, N5666);
or OR2 (N10916, N10871, N2501);
buf BUF1 (N10917, N10910);
buf BUF1 (N10918, N10913);
nor NOR3 (N10919, N10906, N189, N4417);
nand NAND4 (N10920, N10898, N3290, N2877, N5691);
buf BUF1 (N10921, N10917);
buf BUF1 (N10922, N10914);
nor NOR3 (N10923, N10911, N1870, N8145);
xor XOR2 (N10924, N10908, N7813);
nand NAND4 (N10925, N10920, N7058, N2111, N1677);
or OR3 (N10926, N10918, N4915, N1910);
nor NOR2 (N10927, N10921, N3433);
buf BUF1 (N10928, N10919);
xor XOR2 (N10929, N10925, N7287);
xor XOR2 (N10930, N10915, N9672);
nor NOR2 (N10931, N10916, N10716);
nand NAND2 (N10932, N10922, N9004);
or OR2 (N10933, N10927, N5022);
xor XOR2 (N10934, N10931, N4406);
nor NOR2 (N10935, N10933, N8129);
not NOT1 (N10936, N10934);
and AND3 (N10937, N10924, N4371, N3110);
or OR2 (N10938, N10926, N5412);
buf BUF1 (N10939, N10932);
or OR2 (N10940, N10936, N5545);
nand NAND2 (N10941, N10937, N5654);
and AND4 (N10942, N10928, N7425, N4242, N4266);
nand NAND3 (N10943, N10905, N8044, N5258);
xor XOR2 (N10944, N10930, N8653);
not NOT1 (N10945, N10942);
nand NAND4 (N10946, N10938, N2938, N397, N4556);
xor XOR2 (N10947, N10935, N1165);
xor XOR2 (N10948, N10940, N10830);
nand NAND3 (N10949, N10943, N7606, N1387);
not NOT1 (N10950, N10944);
buf BUF1 (N10951, N10946);
xor XOR2 (N10952, N10951, N3372);
nor NOR4 (N10953, N10939, N1377, N6508, N2716);
buf BUF1 (N10954, N10941);
not NOT1 (N10955, N10945);
not NOT1 (N10956, N10923);
or OR4 (N10957, N10955, N2690, N2654, N698);
xor XOR2 (N10958, N10947, N5439);
or OR2 (N10959, N10958, N8);
and AND3 (N10960, N10954, N4996, N10432);
or OR3 (N10961, N10956, N345, N6970);
not NOT1 (N10962, N10929);
nand NAND3 (N10963, N10950, N9793, N7171);
or OR3 (N10964, N10957, N6151, N1279);
xor XOR2 (N10965, N10962, N5319);
and AND2 (N10966, N10963, N3374);
nand NAND2 (N10967, N10960, N9458);
xor XOR2 (N10968, N10953, N6192);
nand NAND2 (N10969, N10966, N9352);
buf BUF1 (N10970, N10969);
nand NAND4 (N10971, N10948, N3258, N5638, N7313);
xor XOR2 (N10972, N10965, N5879);
nor NOR3 (N10973, N10961, N3232, N5565);
buf BUF1 (N10974, N10973);
xor XOR2 (N10975, N10968, N1560);
buf BUF1 (N10976, N10949);
xor XOR2 (N10977, N10972, N7302);
nand NAND3 (N10978, N10959, N5256, N9889);
or OR3 (N10979, N10975, N8195, N5033);
nand NAND2 (N10980, N10974, N10833);
or OR4 (N10981, N10970, N5492, N3088, N8761);
or OR3 (N10982, N10978, N6096, N4273);
not NOT1 (N10983, N10982);
or OR3 (N10984, N10952, N399, N9356);
buf BUF1 (N10985, N10971);
buf BUF1 (N10986, N10980);
buf BUF1 (N10987, N10986);
or OR4 (N10988, N10964, N4594, N10960, N4367);
nor NOR4 (N10989, N10977, N8558, N9949, N9198);
not NOT1 (N10990, N10976);
xor XOR2 (N10991, N10983, N2163);
nand NAND2 (N10992, N10979, N2729);
or OR2 (N10993, N10985, N1997);
or OR3 (N10994, N10993, N10107, N4757);
not NOT1 (N10995, N10989);
and AND4 (N10996, N10994, N7351, N8206, N10950);
nor NOR4 (N10997, N10992, N7599, N6589, N5573);
buf BUF1 (N10998, N10984);
nor NOR4 (N10999, N10991, N6318, N10592, N5215);
and AND4 (N11000, N10995, N6796, N3916, N7711);
nand NAND2 (N11001, N10999, N2833);
xor XOR2 (N11002, N11001, N5595);
not NOT1 (N11003, N10997);
not NOT1 (N11004, N11003);
nand NAND2 (N11005, N10998, N8435);
nand NAND2 (N11006, N11000, N6301);
buf BUF1 (N11007, N10981);
xor XOR2 (N11008, N10967, N8292);
or OR4 (N11009, N11008, N7565, N930, N5755);
and AND3 (N11010, N10996, N451, N5952);
or OR3 (N11011, N11005, N9571, N4102);
and AND4 (N11012, N11006, N10852, N2876, N2203);
buf BUF1 (N11013, N11012);
not NOT1 (N11014, N11004);
nor NOR2 (N11015, N10988, N7767);
nand NAND4 (N11016, N11014, N10385, N3122, N6143);
nor NOR4 (N11017, N11016, N3927, N8410, N724);
nand NAND4 (N11018, N10990, N8917, N6723, N3796);
buf BUF1 (N11019, N11010);
nand NAND4 (N11020, N11017, N5397, N5590, N2660);
buf BUF1 (N11021, N11015);
nand NAND3 (N11022, N10987, N7038, N4284);
nor NOR2 (N11023, N11018, N5392);
nand NAND4 (N11024, N11002, N9052, N6303, N3147);
and AND3 (N11025, N11024, N1989, N9450);
nand NAND4 (N11026, N11020, N8880, N3486, N5543);
nand NAND2 (N11027, N11025, N9760);
and AND3 (N11028, N11027, N6724, N9428);
nor NOR4 (N11029, N11028, N4846, N2679, N1982);
nor NOR3 (N11030, N11013, N9623, N7314);
and AND4 (N11031, N11011, N2571, N10352, N1656);
and AND4 (N11032, N11031, N9164, N7521, N854);
and AND3 (N11033, N11021, N5827, N2572);
not NOT1 (N11034, N11033);
nand NAND4 (N11035, N11009, N10621, N2516, N4848);
nand NAND2 (N11036, N11029, N5990);
buf BUF1 (N11037, N11030);
and AND3 (N11038, N11022, N4590, N5535);
xor XOR2 (N11039, N11023, N1974);
and AND4 (N11040, N11026, N5731, N5860, N1102);
or OR4 (N11041, N11007, N5864, N8959, N9941);
or OR4 (N11042, N11034, N2220, N1280, N4256);
or OR2 (N11043, N11038, N1033);
nor NOR2 (N11044, N11039, N9060);
and AND3 (N11045, N11032, N6305, N9872);
nand NAND4 (N11046, N11019, N2698, N871, N762);
not NOT1 (N11047, N11045);
not NOT1 (N11048, N11040);
buf BUF1 (N11049, N11046);
not NOT1 (N11050, N11036);
xor XOR2 (N11051, N11043, N7766);
nor NOR3 (N11052, N11049, N7132, N6080);
and AND2 (N11053, N11052, N6589);
and AND2 (N11054, N11044, N9293);
nor NOR3 (N11055, N11054, N5892, N425);
and AND2 (N11056, N11035, N1269);
xor XOR2 (N11057, N11056, N8136);
or OR2 (N11058, N11051, N10327);
nand NAND3 (N11059, N11041, N9678, N10677);
nand NAND3 (N11060, N11055, N8494, N1586);
or OR4 (N11061, N11060, N4631, N1573, N4828);
not NOT1 (N11062, N11061);
nor NOR3 (N11063, N11037, N8919, N3730);
nor NOR2 (N11064, N11058, N1602);
and AND2 (N11065, N11053, N354);
nand NAND2 (N11066, N11042, N6652);
nand NAND4 (N11067, N11050, N9372, N8379, N3247);
or OR3 (N11068, N11065, N8385, N6327);
nor NOR2 (N11069, N11063, N6456);
not NOT1 (N11070, N11057);
nand NAND3 (N11071, N11048, N8262, N3866);
nand NAND3 (N11072, N11059, N8039, N8052);
xor XOR2 (N11073, N11066, N9189);
buf BUF1 (N11074, N11047);
xor XOR2 (N11075, N11074, N1021);
not NOT1 (N11076, N11070);
not NOT1 (N11077, N11072);
not NOT1 (N11078, N11075);
nand NAND2 (N11079, N11064, N4642);
or OR3 (N11080, N11069, N7279, N5293);
or OR3 (N11081, N11071, N3432, N5648);
nor NOR2 (N11082, N11062, N8761);
nor NOR3 (N11083, N11076, N6618, N4736);
or OR2 (N11084, N11068, N9303);
or OR2 (N11085, N11078, N6939);
nor NOR2 (N11086, N11082, N9838);
nand NAND4 (N11087, N11086, N6897, N8348, N10901);
not NOT1 (N11088, N11087);
buf BUF1 (N11089, N11073);
not NOT1 (N11090, N11079);
buf BUF1 (N11091, N11067);
buf BUF1 (N11092, N11091);
or OR3 (N11093, N11088, N2280, N2559);
and AND2 (N11094, N11083, N2427);
not NOT1 (N11095, N11080);
or OR4 (N11096, N11093, N3008, N7684, N7377);
and AND2 (N11097, N11090, N3947);
not NOT1 (N11098, N11096);
nor NOR2 (N11099, N11081, N11060);
xor XOR2 (N11100, N11097, N4795);
xor XOR2 (N11101, N11089, N5792);
buf BUF1 (N11102, N11098);
buf BUF1 (N11103, N11100);
buf BUF1 (N11104, N11084);
or OR2 (N11105, N11085, N9672);
xor XOR2 (N11106, N11104, N5727);
nand NAND2 (N11107, N11105, N6293);
or OR3 (N11108, N11103, N2163, N5724);
buf BUF1 (N11109, N11107);
buf BUF1 (N11110, N11108);
and AND3 (N11111, N11077, N5116, N2489);
xor XOR2 (N11112, N11110, N3783);
not NOT1 (N11113, N11106);
nor NOR3 (N11114, N11092, N8839, N1094);
nand NAND2 (N11115, N11114, N140);
and AND3 (N11116, N11095, N7139, N8182);
not NOT1 (N11117, N11116);
and AND4 (N11118, N11109, N3461, N9788, N7625);
or OR4 (N11119, N11111, N7215, N7389, N120);
nand NAND2 (N11120, N11118, N8905);
nand NAND2 (N11121, N11094, N7317);
and AND3 (N11122, N11099, N8212, N3976);
and AND2 (N11123, N11102, N3624);
nor NOR4 (N11124, N11119, N8643, N10549, N7641);
nand NAND2 (N11125, N11112, N1724);
and AND2 (N11126, N11124, N2713);
or OR3 (N11127, N11123, N2747, N6204);
and AND2 (N11128, N11125, N8045);
xor XOR2 (N11129, N11120, N5865);
xor XOR2 (N11130, N11127, N2103);
buf BUF1 (N11131, N11130);
nand NAND4 (N11132, N11117, N1869, N9687, N5043);
or OR3 (N11133, N11122, N7300, N6283);
nor NOR4 (N11134, N11113, N10428, N6977, N6868);
or OR3 (N11135, N11128, N6361, N7361);
not NOT1 (N11136, N11133);
not NOT1 (N11137, N11126);
nor NOR2 (N11138, N11129, N451);
and AND4 (N11139, N11131, N5207, N7218, N5250);
not NOT1 (N11140, N11136);
or OR4 (N11141, N11139, N4805, N9300, N8876);
nor NOR2 (N11142, N11121, N8953);
xor XOR2 (N11143, N11134, N976);
or OR3 (N11144, N11137, N5615, N671);
nand NAND4 (N11145, N11141, N900, N6405, N2761);
buf BUF1 (N11146, N11138);
nor NOR4 (N11147, N11132, N2299, N8351, N518);
or OR2 (N11148, N11143, N2906);
buf BUF1 (N11149, N11142);
not NOT1 (N11150, N11135);
not NOT1 (N11151, N11150);
buf BUF1 (N11152, N11101);
xor XOR2 (N11153, N11144, N3777);
or OR3 (N11154, N11147, N1095, N5656);
buf BUF1 (N11155, N11149);
buf BUF1 (N11156, N11145);
not NOT1 (N11157, N11115);
nand NAND4 (N11158, N11140, N5611, N597, N4884);
and AND2 (N11159, N11155, N10880);
not NOT1 (N11160, N11152);
nand NAND3 (N11161, N11157, N8466, N7492);
nor NOR2 (N11162, N11148, N5935);
and AND2 (N11163, N11158, N9935);
xor XOR2 (N11164, N11161, N736);
or OR3 (N11165, N11156, N5436, N8957);
buf BUF1 (N11166, N11163);
xor XOR2 (N11167, N11159, N7965);
and AND4 (N11168, N11146, N6580, N6163, N5025);
nor NOR4 (N11169, N11160, N1092, N8179, N609);
xor XOR2 (N11170, N11154, N3908);
nand NAND2 (N11171, N11170, N135);
buf BUF1 (N11172, N11168);
nand NAND4 (N11173, N11165, N1904, N7511, N2396);
buf BUF1 (N11174, N11166);
nor NOR3 (N11175, N11173, N10446, N10467);
xor XOR2 (N11176, N11162, N8816);
not NOT1 (N11177, N11167);
buf BUF1 (N11178, N11153);
and AND3 (N11179, N11151, N9195, N3781);
and AND2 (N11180, N11178, N3117);
xor XOR2 (N11181, N11175, N10808);
or OR2 (N11182, N11180, N9603);
nor NOR4 (N11183, N11182, N1627, N2968, N6547);
buf BUF1 (N11184, N11171);
or OR3 (N11185, N11164, N8542, N1609);
not NOT1 (N11186, N11183);
xor XOR2 (N11187, N11186, N8306);
buf BUF1 (N11188, N11176);
xor XOR2 (N11189, N11179, N7463);
nor NOR2 (N11190, N11177, N7948);
xor XOR2 (N11191, N11174, N8103);
buf BUF1 (N11192, N11181);
xor XOR2 (N11193, N11185, N4620);
not NOT1 (N11194, N11190);
or OR4 (N11195, N11189, N9073, N9368, N3690);
buf BUF1 (N11196, N11193);
and AND3 (N11197, N11191, N8126, N6725);
not NOT1 (N11198, N11195);
not NOT1 (N11199, N11197);
xor XOR2 (N11200, N11199, N906);
and AND2 (N11201, N11187, N8892);
xor XOR2 (N11202, N11198, N4387);
nor NOR4 (N11203, N11192, N9801, N9184, N3221);
buf BUF1 (N11204, N11196);
not NOT1 (N11205, N11204);
nand NAND2 (N11206, N11201, N6552);
or OR2 (N11207, N11206, N1333);
or OR4 (N11208, N11184, N8493, N5420, N4159);
nor NOR2 (N11209, N11169, N3148);
nor NOR2 (N11210, N11207, N10111);
or OR2 (N11211, N11200, N5979);
nor NOR3 (N11212, N11209, N8376, N1604);
xor XOR2 (N11213, N11212, N6101);
nand NAND4 (N11214, N11211, N8066, N1420, N8511);
buf BUF1 (N11215, N11213);
nand NAND4 (N11216, N11194, N6814, N356, N10842);
or OR2 (N11217, N11202, N3162);
or OR2 (N11218, N11208, N3925);
nand NAND2 (N11219, N11188, N8401);
or OR4 (N11220, N11210, N7821, N6121, N10790);
buf BUF1 (N11221, N11217);
nor NOR4 (N11222, N11221, N613, N10739, N2574);
and AND3 (N11223, N11219, N5427, N4117);
and AND3 (N11224, N11222, N932, N3595);
not NOT1 (N11225, N11224);
and AND4 (N11226, N11220, N3081, N1644, N30);
nand NAND2 (N11227, N11225, N5163);
nor NOR3 (N11228, N11172, N7980, N5061);
and AND4 (N11229, N11223, N2894, N6296, N6356);
nand NAND2 (N11230, N11228, N10092);
nand NAND3 (N11231, N11203, N6282, N1654);
xor XOR2 (N11232, N11226, N1752);
nor NOR3 (N11233, N11227, N474, N4545);
xor XOR2 (N11234, N11218, N6918);
buf BUF1 (N11235, N11234);
and AND4 (N11236, N11232, N8783, N2607, N6616);
buf BUF1 (N11237, N11214);
or OR3 (N11238, N11231, N3052, N5953);
and AND3 (N11239, N11238, N6432, N1935);
nor NOR4 (N11240, N11216, N6304, N5329, N706);
nor NOR2 (N11241, N11205, N7775);
or OR4 (N11242, N11237, N855, N3466, N8365);
nor NOR4 (N11243, N11230, N5009, N9530, N4442);
xor XOR2 (N11244, N11242, N5555);
not NOT1 (N11245, N11215);
not NOT1 (N11246, N11235);
or OR3 (N11247, N11243, N9151, N580);
not NOT1 (N11248, N11247);
xor XOR2 (N11249, N11229, N924);
or OR4 (N11250, N11236, N7001, N5205, N9947);
buf BUF1 (N11251, N11240);
buf BUF1 (N11252, N11233);
nand NAND2 (N11253, N11239, N9403);
and AND2 (N11254, N11248, N4627);
xor XOR2 (N11255, N11245, N1576);
and AND4 (N11256, N11250, N3608, N10558, N10813);
nor NOR2 (N11257, N11254, N1367);
not NOT1 (N11258, N11255);
not NOT1 (N11259, N11244);
and AND4 (N11260, N11258, N4230, N918, N8596);
nor NOR2 (N11261, N11249, N2126);
or OR2 (N11262, N11259, N2737);
nand NAND3 (N11263, N11241, N7761, N1000);
nand NAND3 (N11264, N11253, N7284, N3753);
buf BUF1 (N11265, N11260);
xor XOR2 (N11266, N11246, N1173);
xor XOR2 (N11267, N11265, N307);
and AND2 (N11268, N11263, N3948);
nand NAND2 (N11269, N11262, N9645);
nand NAND2 (N11270, N11252, N8928);
or OR3 (N11271, N11257, N7206, N1944);
or OR3 (N11272, N11268, N4837, N3589);
nand NAND2 (N11273, N11266, N7098);
nand NAND3 (N11274, N11267, N5648, N8276);
not NOT1 (N11275, N11256);
nand NAND4 (N11276, N11272, N10602, N3953, N9747);
nand NAND3 (N11277, N11273, N8226, N4401);
and AND2 (N11278, N11271, N9457);
buf BUF1 (N11279, N11264);
and AND2 (N11280, N11274, N2834);
not NOT1 (N11281, N11270);
not NOT1 (N11282, N11261);
buf BUF1 (N11283, N11275);
and AND3 (N11284, N11276, N3755, N1878);
buf BUF1 (N11285, N11277);
nor NOR2 (N11286, N11281, N7178);
or OR2 (N11287, N11283, N3933);
buf BUF1 (N11288, N11285);
buf BUF1 (N11289, N11279);
not NOT1 (N11290, N11280);
or OR4 (N11291, N11284, N5482, N4039, N6462);
and AND4 (N11292, N11288, N7819, N8759, N10159);
nor NOR2 (N11293, N11291, N7975);
and AND4 (N11294, N11293, N8951, N8770, N6081);
or OR2 (N11295, N11294, N9162);
nor NOR4 (N11296, N11292, N7126, N2575, N10845);
and AND3 (N11297, N11289, N5002, N4209);
nand NAND3 (N11298, N11290, N1401, N5644);
buf BUF1 (N11299, N11287);
and AND3 (N11300, N11251, N9781, N2974);
buf BUF1 (N11301, N11300);
or OR4 (N11302, N11295, N9912, N4532, N637);
and AND2 (N11303, N11299, N5471);
or OR4 (N11304, N11302, N5833, N8145, N8015);
not NOT1 (N11305, N11282);
buf BUF1 (N11306, N11297);
nor NOR3 (N11307, N11298, N374, N837);
nand NAND4 (N11308, N11306, N3755, N7479, N1623);
and AND2 (N11309, N11308, N6165);
or OR3 (N11310, N11296, N10952, N5809);
nand NAND4 (N11311, N11278, N355, N982, N4984);
nor NOR3 (N11312, N11307, N7674, N2687);
buf BUF1 (N11313, N11303);
nand NAND2 (N11314, N11301, N2049);
or OR4 (N11315, N11309, N10831, N5968, N1335);
nor NOR3 (N11316, N11314, N9262, N5203);
and AND3 (N11317, N11269, N1705, N6616);
nand NAND2 (N11318, N11311, N6593);
and AND3 (N11319, N11318, N5172, N4135);
nand NAND3 (N11320, N11286, N1771, N7189);
and AND2 (N11321, N11319, N4189);
or OR4 (N11322, N11317, N9635, N5029, N6589);
or OR2 (N11323, N11304, N11318);
and AND3 (N11324, N11316, N7534, N4158);
and AND2 (N11325, N11320, N1654);
and AND3 (N11326, N11313, N1968, N11179);
and AND3 (N11327, N11321, N9809, N4925);
nand NAND2 (N11328, N11325, N8595);
nor NOR2 (N11329, N11323, N299);
nand NAND4 (N11330, N11326, N925, N6271, N9377);
or OR4 (N11331, N11324, N1655, N7344, N528);
nand NAND4 (N11332, N11329, N10905, N6199, N4388);
nor NOR4 (N11333, N11322, N6385, N9321, N9595);
nor NOR4 (N11334, N11328, N4553, N8677, N211);
nand NAND2 (N11335, N11305, N2846);
not NOT1 (N11336, N11335);
nand NAND2 (N11337, N11336, N8507);
not NOT1 (N11338, N11331);
nor NOR2 (N11339, N11310, N1241);
not NOT1 (N11340, N11330);
nor NOR4 (N11341, N11333, N3444, N69, N3381);
nand NAND3 (N11342, N11327, N3685, N6342);
nand NAND2 (N11343, N11342, N9650);
or OR4 (N11344, N11343, N9112, N9522, N8599);
buf BUF1 (N11345, N11315);
nor NOR2 (N11346, N11344, N7832);
nor NOR4 (N11347, N11338, N7923, N2228, N2428);
or OR4 (N11348, N11346, N2826, N9172, N4920);
xor XOR2 (N11349, N11341, N6576);
nand NAND2 (N11350, N11347, N5854);
nand NAND4 (N11351, N11348, N577, N9865, N10537);
or OR4 (N11352, N11312, N10105, N4302, N3103);
or OR4 (N11353, N11339, N4401, N10520, N7927);
or OR4 (N11354, N11351, N6142, N5503, N6342);
nand NAND4 (N11355, N11354, N11252, N3929, N4021);
nand NAND2 (N11356, N11345, N8008);
buf BUF1 (N11357, N11350);
xor XOR2 (N11358, N11352, N3135);
nor NOR4 (N11359, N11337, N8302, N10733, N3477);
xor XOR2 (N11360, N11355, N9330);
nor NOR3 (N11361, N11349, N9880, N3844);
or OR3 (N11362, N11359, N3708, N8721);
not NOT1 (N11363, N11362);
nor NOR4 (N11364, N11356, N7875, N615, N8650);
nor NOR3 (N11365, N11332, N3450, N4932);
not NOT1 (N11366, N11364);
xor XOR2 (N11367, N11357, N11234);
nor NOR2 (N11368, N11340, N5796);
buf BUF1 (N11369, N11365);
not NOT1 (N11370, N11367);
buf BUF1 (N11371, N11358);
nor NOR4 (N11372, N11368, N4836, N3754, N11136);
nor NOR2 (N11373, N11360, N574);
buf BUF1 (N11374, N11370);
xor XOR2 (N11375, N11373, N1133);
and AND4 (N11376, N11361, N951, N11117, N1593);
and AND3 (N11377, N11353, N3143, N6147);
buf BUF1 (N11378, N11377);
and AND3 (N11379, N11371, N3563, N3196);
nand NAND4 (N11380, N11369, N3779, N7763, N3691);
nor NOR2 (N11381, N11363, N1201);
buf BUF1 (N11382, N11375);
buf BUF1 (N11383, N11381);
nor NOR3 (N11384, N11378, N8786, N580);
nor NOR3 (N11385, N11372, N2802, N7693);
or OR4 (N11386, N11374, N8999, N3071, N2958);
not NOT1 (N11387, N11376);
nor NOR4 (N11388, N11385, N10038, N6270, N7893);
and AND3 (N11389, N11366, N3469, N10608);
and AND3 (N11390, N11379, N7174, N3795);
xor XOR2 (N11391, N11389, N8492);
nand NAND4 (N11392, N11380, N6094, N5431, N10903);
nand NAND4 (N11393, N11388, N2367, N4370, N6230);
buf BUF1 (N11394, N11387);
buf BUF1 (N11395, N11386);
nand NAND4 (N11396, N11383, N939, N11298, N4464);
xor XOR2 (N11397, N11384, N4825);
not NOT1 (N11398, N11393);
nor NOR4 (N11399, N11392, N7089, N1917, N6023);
xor XOR2 (N11400, N11390, N7130);
or OR4 (N11401, N11382, N242, N9147, N4884);
not NOT1 (N11402, N11401);
and AND3 (N11403, N11400, N4093, N3213);
or OR4 (N11404, N11396, N700, N7224, N6664);
nor NOR3 (N11405, N11395, N5332, N6272);
or OR2 (N11406, N11403, N8865);
or OR3 (N11407, N11334, N10295, N8238);
nor NOR4 (N11408, N11402, N1418, N8203, N3773);
xor XOR2 (N11409, N11405, N11071);
or OR4 (N11410, N11399, N9846, N1105, N3440);
and AND2 (N11411, N11398, N1395);
buf BUF1 (N11412, N11394);
nor NOR2 (N11413, N11406, N353);
nor NOR4 (N11414, N11410, N5013, N321, N9933);
nand NAND4 (N11415, N11414, N3522, N1727, N7403);
buf BUF1 (N11416, N11391);
or OR4 (N11417, N11408, N8961, N5429, N312);
nor NOR2 (N11418, N11416, N880);
nor NOR4 (N11419, N11418, N4126, N3818, N9883);
not NOT1 (N11420, N11415);
nor NOR4 (N11421, N11420, N991, N7555, N4539);
xor XOR2 (N11422, N11421, N4505);
nor NOR4 (N11423, N11412, N2021, N7267, N2736);
not NOT1 (N11424, N11417);
nor NOR3 (N11425, N11409, N7317, N4024);
not NOT1 (N11426, N11397);
xor XOR2 (N11427, N11419, N1670);
nor NOR3 (N11428, N11423, N10671, N5694);
nor NOR4 (N11429, N11425, N11076, N7269, N4852);
nor NOR2 (N11430, N11422, N10056);
or OR4 (N11431, N11407, N5493, N2459, N6636);
not NOT1 (N11432, N11429);
buf BUF1 (N11433, N11432);
or OR2 (N11434, N11431, N10283);
nor NOR2 (N11435, N11428, N270);
and AND4 (N11436, N11435, N8294, N1840, N3165);
not NOT1 (N11437, N11430);
or OR3 (N11438, N11424, N9461, N6197);
nor NOR3 (N11439, N11413, N4415, N9846);
nor NOR3 (N11440, N11439, N7059, N4546);
nand NAND4 (N11441, N11438, N4952, N4913, N3739);
xor XOR2 (N11442, N11433, N1714);
nor NOR4 (N11443, N11436, N8357, N4746, N3611);
and AND4 (N11444, N11442, N7642, N3576, N1092);
xor XOR2 (N11445, N11427, N3755);
nand NAND2 (N11446, N11426, N3026);
xor XOR2 (N11447, N11443, N5846);
or OR2 (N11448, N11441, N11255);
or OR2 (N11449, N11447, N6504);
not NOT1 (N11450, N11445);
not NOT1 (N11451, N11404);
nand NAND2 (N11452, N11448, N8764);
not NOT1 (N11453, N11440);
not NOT1 (N11454, N11437);
nor NOR3 (N11455, N11454, N3132, N2331);
nor NOR2 (N11456, N11444, N3163);
xor XOR2 (N11457, N11449, N87);
nor NOR4 (N11458, N11453, N3299, N10166, N4414);
and AND4 (N11459, N11458, N6613, N926, N3762);
or OR4 (N11460, N11446, N5080, N5486, N6905);
buf BUF1 (N11461, N11455);
not NOT1 (N11462, N11460);
nor NOR3 (N11463, N11457, N1696, N10766);
buf BUF1 (N11464, N11451);
and AND4 (N11465, N11464, N10092, N1756, N9600);
or OR2 (N11466, N11411, N6231);
and AND2 (N11467, N11456, N3513);
buf BUF1 (N11468, N11461);
buf BUF1 (N11469, N11450);
xor XOR2 (N11470, N11469, N5127);
nand NAND3 (N11471, N11462, N7402, N10187);
xor XOR2 (N11472, N11467, N5181);
not NOT1 (N11473, N11470);
nand NAND2 (N11474, N11465, N8450);
xor XOR2 (N11475, N11452, N11301);
nand NAND4 (N11476, N11468, N2604, N9654, N4480);
nand NAND3 (N11477, N11474, N10898, N8498);
and AND4 (N11478, N11475, N1534, N8191, N9481);
not NOT1 (N11479, N11477);
and AND3 (N11480, N11459, N313, N581);
nand NAND3 (N11481, N11434, N5329, N9058);
buf BUF1 (N11482, N11479);
buf BUF1 (N11483, N11463);
buf BUF1 (N11484, N11480);
not NOT1 (N11485, N11478);
nand NAND2 (N11486, N11484, N7347);
buf BUF1 (N11487, N11486);
nand NAND3 (N11488, N11482, N10409, N7974);
not NOT1 (N11489, N11473);
xor XOR2 (N11490, N11471, N4710);
or OR2 (N11491, N11488, N8225);
xor XOR2 (N11492, N11489, N662);
nand NAND2 (N11493, N11483, N8374);
nor NOR4 (N11494, N11476, N2503, N1242, N9233);
nand NAND4 (N11495, N11485, N5897, N7660, N5129);
nand NAND4 (N11496, N11494, N11202, N10659, N8441);
buf BUF1 (N11497, N11472);
or OR4 (N11498, N11492, N341, N3597, N9112);
nor NOR4 (N11499, N11466, N522, N4882, N1378);
nor NOR4 (N11500, N11495, N476, N1939, N2509);
buf BUF1 (N11501, N11497);
and AND2 (N11502, N11490, N2477);
not NOT1 (N11503, N11500);
not NOT1 (N11504, N11493);
buf BUF1 (N11505, N11502);
and AND3 (N11506, N11505, N635, N8449);
not NOT1 (N11507, N11503);
nand NAND3 (N11508, N11498, N1825, N307);
nand NAND2 (N11509, N11496, N7503);
xor XOR2 (N11510, N11499, N1760);
and AND3 (N11511, N11507, N697, N9964);
nor NOR4 (N11512, N11491, N10164, N4541, N4431);
not NOT1 (N11513, N11504);
not NOT1 (N11514, N11512);
and AND4 (N11515, N11514, N5616, N3934, N11075);
nand NAND4 (N11516, N11501, N5070, N1523, N9890);
xor XOR2 (N11517, N11510, N9459);
buf BUF1 (N11518, N11517);
buf BUF1 (N11519, N11515);
buf BUF1 (N11520, N11508);
not NOT1 (N11521, N11481);
or OR3 (N11522, N11519, N3243, N2505);
buf BUF1 (N11523, N11518);
or OR3 (N11524, N11513, N8851, N4978);
buf BUF1 (N11525, N11509);
or OR3 (N11526, N11523, N6843, N8591);
not NOT1 (N11527, N11525);
buf BUF1 (N11528, N11524);
not NOT1 (N11529, N11522);
not NOT1 (N11530, N11487);
or OR3 (N11531, N11529, N1441, N7882);
nor NOR4 (N11532, N11506, N2506, N1771, N4927);
xor XOR2 (N11533, N11526, N7773);
or OR4 (N11534, N11516, N6162, N9191, N9858);
nand NAND3 (N11535, N11528, N4038, N8502);
xor XOR2 (N11536, N11530, N10604);
not NOT1 (N11537, N11536);
buf BUF1 (N11538, N11531);
nand NAND4 (N11539, N11537, N2461, N4777, N2127);
buf BUF1 (N11540, N11534);
not NOT1 (N11541, N11527);
nor NOR2 (N11542, N11521, N8969);
buf BUF1 (N11543, N11540);
not NOT1 (N11544, N11543);
nor NOR3 (N11545, N11541, N5524, N6427);
nand NAND3 (N11546, N11535, N1305, N9538);
not NOT1 (N11547, N11511);
not NOT1 (N11548, N11532);
not NOT1 (N11549, N11547);
or OR4 (N11550, N11545, N3473, N10677, N8813);
or OR3 (N11551, N11546, N9465, N5236);
and AND4 (N11552, N11549, N10453, N1000, N1334);
nor NOR4 (N11553, N11548, N5681, N9663, N1306);
not NOT1 (N11554, N11544);
or OR2 (N11555, N11542, N10895);
xor XOR2 (N11556, N11533, N2220);
xor XOR2 (N11557, N11520, N8752);
and AND2 (N11558, N11538, N11062);
nor NOR3 (N11559, N11550, N4691, N8680);
not NOT1 (N11560, N11552);
or OR4 (N11561, N11539, N3872, N268, N416);
and AND3 (N11562, N11551, N9705, N4009);
buf BUF1 (N11563, N11560);
or OR2 (N11564, N11562, N7398);
buf BUF1 (N11565, N11564);
nand NAND4 (N11566, N11557, N3209, N6026, N1790);
and AND2 (N11567, N11563, N2490);
xor XOR2 (N11568, N11566, N2658);
nand NAND2 (N11569, N11558, N4727);
xor XOR2 (N11570, N11556, N9062);
nor NOR4 (N11571, N11570, N11081, N6106, N5673);
not NOT1 (N11572, N11568);
buf BUF1 (N11573, N11553);
nor NOR3 (N11574, N11561, N2569, N6071);
buf BUF1 (N11575, N11573);
or OR3 (N11576, N11575, N129, N5160);
buf BUF1 (N11577, N11571);
nor NOR3 (N11578, N11572, N6369, N8257);
and AND4 (N11579, N11554, N6123, N10007, N2134);
buf BUF1 (N11580, N11567);
or OR2 (N11581, N11580, N7566);
or OR2 (N11582, N11576, N2279);
or OR4 (N11583, N11581, N10669, N2991, N118);
or OR3 (N11584, N11577, N2253, N1522);
nand NAND4 (N11585, N11578, N3219, N6369, N7526);
nand NAND2 (N11586, N11559, N7567);
nor NOR3 (N11587, N11569, N1033, N9548);
nand NAND4 (N11588, N11555, N8602, N4465, N3853);
or OR2 (N11589, N11565, N1024);
nand NAND2 (N11590, N11586, N8246);
xor XOR2 (N11591, N11585, N768);
xor XOR2 (N11592, N11583, N1137);
xor XOR2 (N11593, N11574, N9084);
nor NOR3 (N11594, N11591, N3633, N8384);
or OR3 (N11595, N11592, N8653, N5334);
buf BUF1 (N11596, N11579);
nand NAND3 (N11597, N11596, N234, N10751);
nor NOR3 (N11598, N11595, N5050, N7802);
or OR4 (N11599, N11588, N4004, N9903, N140);
and AND3 (N11600, N11594, N4766, N4058);
nor NOR2 (N11601, N11584, N6337);
nor NOR3 (N11602, N11589, N8151, N7302);
buf BUF1 (N11603, N11601);
buf BUF1 (N11604, N11590);
nand NAND3 (N11605, N11603, N4449, N3457);
or OR2 (N11606, N11593, N2799);
and AND2 (N11607, N11606, N4398);
buf BUF1 (N11608, N11598);
or OR3 (N11609, N11582, N8230, N1108);
buf BUF1 (N11610, N11604);
nand NAND4 (N11611, N11610, N2322, N9978, N2627);
buf BUF1 (N11612, N11608);
buf BUF1 (N11613, N11609);
xor XOR2 (N11614, N11612, N1999);
xor XOR2 (N11615, N11602, N8447);
nand NAND3 (N11616, N11605, N9419, N2268);
and AND2 (N11617, N11587, N10094);
buf BUF1 (N11618, N11599);
not NOT1 (N11619, N11618);
not NOT1 (N11620, N11611);
buf BUF1 (N11621, N11607);
not NOT1 (N11622, N11597);
not NOT1 (N11623, N11622);
and AND3 (N11624, N11614, N7300, N527);
not NOT1 (N11625, N11616);
xor XOR2 (N11626, N11620, N3452);
buf BUF1 (N11627, N11615);
nand NAND3 (N11628, N11626, N9796, N7244);
or OR2 (N11629, N11600, N11273);
nand NAND3 (N11630, N11621, N7537, N3119);
buf BUF1 (N11631, N11627);
and AND2 (N11632, N11625, N882);
and AND3 (N11633, N11629, N207, N4264);
xor XOR2 (N11634, N11624, N10017);
and AND3 (N11635, N11613, N2054, N4963);
and AND3 (N11636, N11633, N10540, N6088);
not NOT1 (N11637, N11631);
nor NOR4 (N11638, N11634, N9830, N8276, N1346);
nand NAND2 (N11639, N11617, N10624);
not NOT1 (N11640, N11632);
and AND2 (N11641, N11637, N8389);
not NOT1 (N11642, N11636);
nor NOR3 (N11643, N11640, N3120, N7986);
buf BUF1 (N11644, N11639);
nor NOR3 (N11645, N11638, N6576, N9524);
or OR2 (N11646, N11628, N10459);
xor XOR2 (N11647, N11643, N5002);
xor XOR2 (N11648, N11646, N7961);
and AND3 (N11649, N11645, N9211, N4173);
or OR4 (N11650, N11630, N8073, N4621, N9138);
nor NOR4 (N11651, N11623, N11113, N11537, N2568);
and AND4 (N11652, N11642, N7822, N10059, N174);
nor NOR2 (N11653, N11651, N10334);
and AND2 (N11654, N11653, N11569);
or OR3 (N11655, N11641, N1155, N11248);
xor XOR2 (N11656, N11650, N4510);
xor XOR2 (N11657, N11649, N1568);
nand NAND4 (N11658, N11648, N6043, N10339, N7471);
nor NOR3 (N11659, N11635, N9171, N9582);
buf BUF1 (N11660, N11655);
xor XOR2 (N11661, N11657, N3383);
nor NOR2 (N11662, N11658, N8734);
nor NOR2 (N11663, N11652, N4356);
buf BUF1 (N11664, N11619);
xor XOR2 (N11665, N11644, N3615);
and AND3 (N11666, N11647, N3172, N2495);
or OR2 (N11667, N11656, N1954);
and AND2 (N11668, N11662, N3272);
xor XOR2 (N11669, N11660, N3676);
and AND4 (N11670, N11668, N912, N3454, N4660);
and AND3 (N11671, N11670, N371, N10281);
and AND4 (N11672, N11659, N1578, N10627, N9183);
xor XOR2 (N11673, N11667, N448);
nand NAND2 (N11674, N11673, N253);
xor XOR2 (N11675, N11672, N718);
buf BUF1 (N11676, N11671);
buf BUF1 (N11677, N11676);
or OR3 (N11678, N11669, N4943, N3231);
buf BUF1 (N11679, N11677);
or OR3 (N11680, N11661, N6266, N4166);
or OR2 (N11681, N11675, N842);
not NOT1 (N11682, N11665);
or OR4 (N11683, N11674, N171, N2364, N2052);
nand NAND3 (N11684, N11678, N7931, N776);
xor XOR2 (N11685, N11684, N1747);
xor XOR2 (N11686, N11679, N5013);
and AND4 (N11687, N11663, N5463, N1627, N4566);
nor NOR2 (N11688, N11654, N8922);
xor XOR2 (N11689, N11664, N7223);
nand NAND2 (N11690, N11688, N11057);
and AND4 (N11691, N11689, N9462, N4678, N10215);
buf BUF1 (N11692, N11666);
nor NOR4 (N11693, N11680, N6418, N9988, N2561);
xor XOR2 (N11694, N11687, N4904);
not NOT1 (N11695, N11693);
buf BUF1 (N11696, N11694);
xor XOR2 (N11697, N11683, N2641);
and AND2 (N11698, N11681, N4884);
nor NOR2 (N11699, N11692, N1218);
nand NAND2 (N11700, N11690, N5716);
buf BUF1 (N11701, N11697);
and AND2 (N11702, N11691, N124);
nor NOR2 (N11703, N11685, N1628);
buf BUF1 (N11704, N11702);
and AND3 (N11705, N11700, N9841, N6161);
buf BUF1 (N11706, N11696);
xor XOR2 (N11707, N11705, N4692);
buf BUF1 (N11708, N11701);
nand NAND3 (N11709, N11703, N432, N2378);
not NOT1 (N11710, N11707);
not NOT1 (N11711, N11709);
nor NOR2 (N11712, N11711, N2146);
and AND2 (N11713, N11708, N2040);
nand NAND3 (N11714, N11698, N8434, N7725);
buf BUF1 (N11715, N11695);
not NOT1 (N11716, N11712);
nand NAND3 (N11717, N11710, N7949, N4966);
nor NOR3 (N11718, N11715, N5436, N2512);
not NOT1 (N11719, N11682);
or OR4 (N11720, N11719, N9551, N1373, N2086);
buf BUF1 (N11721, N11686);
not NOT1 (N11722, N11714);
nor NOR4 (N11723, N11716, N8264, N11670, N5269);
or OR4 (N11724, N11722, N3329, N3063, N5096);
nor NOR3 (N11725, N11706, N8577, N2100);
xor XOR2 (N11726, N11725, N9346);
or OR2 (N11727, N11713, N9505);
buf BUF1 (N11728, N11724);
and AND4 (N11729, N11699, N5498, N3300, N3327);
or OR4 (N11730, N11729, N7476, N4563, N6203);
buf BUF1 (N11731, N11718);
nand NAND4 (N11732, N11721, N1043, N7110, N3978);
buf BUF1 (N11733, N11727);
xor XOR2 (N11734, N11717, N4858);
xor XOR2 (N11735, N11730, N9264);
not NOT1 (N11736, N11720);
xor XOR2 (N11737, N11728, N8549);
buf BUF1 (N11738, N11726);
or OR3 (N11739, N11733, N5407, N3051);
and AND3 (N11740, N11736, N8273, N7015);
xor XOR2 (N11741, N11723, N7493);
nor NOR2 (N11742, N11734, N11610);
and AND2 (N11743, N11731, N3429);
buf BUF1 (N11744, N11738);
not NOT1 (N11745, N11735);
buf BUF1 (N11746, N11740);
and AND3 (N11747, N11744, N11224, N9881);
nor NOR2 (N11748, N11741, N7931);
nor NOR4 (N11749, N11739, N9946, N11632, N9591);
xor XOR2 (N11750, N11743, N1388);
not NOT1 (N11751, N11750);
nor NOR4 (N11752, N11749, N11523, N9609, N1772);
buf BUF1 (N11753, N11745);
nor NOR4 (N11754, N11742, N6157, N9443, N1893);
and AND2 (N11755, N11753, N9026);
xor XOR2 (N11756, N11732, N6289);
buf BUF1 (N11757, N11756);
and AND2 (N11758, N11748, N11627);
and AND2 (N11759, N11737, N2407);
or OR3 (N11760, N11751, N4808, N7541);
and AND3 (N11761, N11704, N2092, N776);
or OR2 (N11762, N11754, N8563);
buf BUF1 (N11763, N11755);
or OR4 (N11764, N11761, N3848, N10927, N9480);
not NOT1 (N11765, N11758);
and AND4 (N11766, N11760, N1863, N692, N9700);
nor NOR4 (N11767, N11765, N2801, N3656, N1981);
nand NAND3 (N11768, N11766, N11066, N9036);
buf BUF1 (N11769, N11746);
nand NAND3 (N11770, N11752, N9893, N10880);
not NOT1 (N11771, N11759);
buf BUF1 (N11772, N11769);
xor XOR2 (N11773, N11747, N465);
nand NAND2 (N11774, N11772, N3197);
buf BUF1 (N11775, N11767);
not NOT1 (N11776, N11774);
not NOT1 (N11777, N11776);
buf BUF1 (N11778, N11770);
or OR3 (N11779, N11763, N9035, N6244);
not NOT1 (N11780, N11779);
not NOT1 (N11781, N11778);
and AND3 (N11782, N11781, N8318, N242);
buf BUF1 (N11783, N11757);
xor XOR2 (N11784, N11782, N8132);
buf BUF1 (N11785, N11773);
nand NAND2 (N11786, N11783, N7517);
nand NAND2 (N11787, N11784, N11356);
buf BUF1 (N11788, N11764);
nor NOR3 (N11789, N11777, N60, N4682);
nor NOR2 (N11790, N11788, N2087);
buf BUF1 (N11791, N11775);
buf BUF1 (N11792, N11791);
or OR2 (N11793, N11785, N544);
not NOT1 (N11794, N11771);
xor XOR2 (N11795, N11789, N4723);
or OR3 (N11796, N11793, N9229, N5597);
and AND4 (N11797, N11786, N4559, N8561, N10504);
and AND4 (N11798, N11780, N4966, N3265, N8774);
buf BUF1 (N11799, N11790);
and AND2 (N11800, N11794, N8142);
nor NOR2 (N11801, N11796, N2430);
and AND3 (N11802, N11768, N9200, N5094);
or OR2 (N11803, N11802, N894);
not NOT1 (N11804, N11799);
not NOT1 (N11805, N11803);
not NOT1 (N11806, N11800);
and AND4 (N11807, N11797, N6475, N5163, N7007);
nand NAND3 (N11808, N11798, N6875, N6299);
nor NOR4 (N11809, N11806, N6056, N2481, N6054);
nand NAND4 (N11810, N11807, N8757, N1079, N917);
not NOT1 (N11811, N11801);
or OR4 (N11812, N11792, N542, N4453, N3317);
and AND4 (N11813, N11795, N6795, N679, N323);
buf BUF1 (N11814, N11809);
nor NOR2 (N11815, N11808, N5120);
or OR2 (N11816, N11810, N9809);
nor NOR4 (N11817, N11816, N5707, N9341, N5649);
buf BUF1 (N11818, N11813);
not NOT1 (N11819, N11818);
not NOT1 (N11820, N11815);
or OR3 (N11821, N11817, N11337, N1341);
or OR3 (N11822, N11819, N724, N8160);
xor XOR2 (N11823, N11820, N7543);
and AND2 (N11824, N11804, N6003);
nand NAND3 (N11825, N11805, N10160, N2572);
nor NOR4 (N11826, N11762, N1618, N1000, N7832);
buf BUF1 (N11827, N11811);
xor XOR2 (N11828, N11787, N8067);
not NOT1 (N11829, N11814);
xor XOR2 (N11830, N11826, N10400);
not NOT1 (N11831, N11825);
nor NOR2 (N11832, N11828, N8348);
nand NAND3 (N11833, N11823, N3794, N342);
nand NAND4 (N11834, N11812, N6420, N3691, N5594);
or OR2 (N11835, N11833, N5835);
or OR4 (N11836, N11831, N1470, N8363, N11310);
or OR2 (N11837, N11832, N8655);
nor NOR4 (N11838, N11830, N6000, N9831, N11489);
nand NAND2 (N11839, N11836, N3663);
xor XOR2 (N11840, N11837, N3771);
nor NOR3 (N11841, N11835, N11220, N11304);
and AND2 (N11842, N11838, N10773);
buf BUF1 (N11843, N11822);
xor XOR2 (N11844, N11841, N2157);
and AND2 (N11845, N11843, N4308);
buf BUF1 (N11846, N11824);
and AND3 (N11847, N11829, N198, N5136);
or OR3 (N11848, N11840, N2247, N8380);
buf BUF1 (N11849, N11834);
not NOT1 (N11850, N11849);
and AND2 (N11851, N11850, N4110);
not NOT1 (N11852, N11847);
or OR3 (N11853, N11845, N11517, N10526);
xor XOR2 (N11854, N11851, N2997);
and AND2 (N11855, N11853, N11465);
or OR2 (N11856, N11855, N6805);
or OR2 (N11857, N11839, N8814);
or OR4 (N11858, N11842, N10920, N9737, N7179);
nand NAND4 (N11859, N11857, N8511, N4818, N8039);
and AND2 (N11860, N11844, N2839);
nand NAND4 (N11861, N11858, N3868, N5555, N4282);
not NOT1 (N11862, N11846);
nand NAND2 (N11863, N11848, N7230);
xor XOR2 (N11864, N11861, N8966);
not NOT1 (N11865, N11862);
buf BUF1 (N11866, N11852);
not NOT1 (N11867, N11856);
nor NOR3 (N11868, N11860, N9012, N7866);
not NOT1 (N11869, N11866);
or OR3 (N11870, N11867, N139, N930);
not NOT1 (N11871, N11869);
nand NAND4 (N11872, N11821, N985, N2626, N11555);
and AND3 (N11873, N11827, N9177, N11250);
nor NOR3 (N11874, N11872, N6511, N10621);
not NOT1 (N11875, N11863);
or OR3 (N11876, N11864, N9984, N7077);
or OR3 (N11877, N11859, N11316, N9490);
and AND3 (N11878, N11874, N9422, N10987);
and AND2 (N11879, N11854, N10082);
or OR3 (N11880, N11875, N10169, N2614);
and AND2 (N11881, N11880, N8233);
and AND2 (N11882, N11870, N1722);
buf BUF1 (N11883, N11881);
not NOT1 (N11884, N11873);
xor XOR2 (N11885, N11877, N3509);
xor XOR2 (N11886, N11879, N597);
not NOT1 (N11887, N11865);
buf BUF1 (N11888, N11886);
xor XOR2 (N11889, N11888, N3556);
and AND3 (N11890, N11883, N3740, N1141);
xor XOR2 (N11891, N11889, N5557);
or OR4 (N11892, N11878, N9916, N65, N10484);
buf BUF1 (N11893, N11887);
buf BUF1 (N11894, N11891);
buf BUF1 (N11895, N11884);
nand NAND2 (N11896, N11892, N939);
buf BUF1 (N11897, N11895);
xor XOR2 (N11898, N11896, N11387);
nand NAND3 (N11899, N11890, N2933, N9080);
nand NAND2 (N11900, N11885, N3643);
nor NOR4 (N11901, N11899, N6751, N4347, N4802);
nor NOR4 (N11902, N11900, N10528, N1045, N579);
or OR4 (N11903, N11901, N7871, N6950, N3740);
nand NAND3 (N11904, N11902, N10379, N7397);
or OR2 (N11905, N11897, N7684);
nand NAND2 (N11906, N11871, N9260);
buf BUF1 (N11907, N11868);
buf BUF1 (N11908, N11893);
and AND2 (N11909, N11908, N9717);
buf BUF1 (N11910, N11882);
not NOT1 (N11911, N11906);
nand NAND3 (N11912, N11911, N8815, N6230);
and AND4 (N11913, N11904, N8398, N5857, N8635);
nor NOR3 (N11914, N11913, N4420, N10312);
not NOT1 (N11915, N11910);
not NOT1 (N11916, N11907);
buf BUF1 (N11917, N11894);
not NOT1 (N11918, N11909);
nor NOR2 (N11919, N11916, N9764);
nor NOR2 (N11920, N11912, N2425);
buf BUF1 (N11921, N11914);
nand NAND2 (N11922, N11921, N10080);
xor XOR2 (N11923, N11917, N11512);
nor NOR2 (N11924, N11918, N9454);
or OR3 (N11925, N11905, N11178, N3766);
not NOT1 (N11926, N11915);
and AND3 (N11927, N11924, N8004, N2746);
not NOT1 (N11928, N11923);
xor XOR2 (N11929, N11903, N9965);
not NOT1 (N11930, N11925);
or OR4 (N11931, N11929, N8219, N4408, N5739);
and AND2 (N11932, N11930, N3202);
nand NAND3 (N11933, N11920, N4469, N7268);
nor NOR2 (N11934, N11927, N8522);
buf BUF1 (N11935, N11928);
or OR4 (N11936, N11926, N4642, N3549, N8256);
not NOT1 (N11937, N11919);
nor NOR3 (N11938, N11936, N1551, N361);
or OR2 (N11939, N11876, N6215);
buf BUF1 (N11940, N11938);
xor XOR2 (N11941, N11933, N281);
and AND4 (N11942, N11922, N5873, N812, N5894);
nand NAND2 (N11943, N11898, N1303);
or OR2 (N11944, N11931, N5441);
xor XOR2 (N11945, N11935, N32);
or OR2 (N11946, N11944, N11299);
and AND4 (N11947, N11941, N8376, N914, N1980);
and AND2 (N11948, N11937, N11778);
buf BUF1 (N11949, N11946);
and AND4 (N11950, N11940, N2260, N1356, N11776);
nor NOR3 (N11951, N11943, N8749, N2339);
nor NOR3 (N11952, N11947, N574, N10437);
nor NOR2 (N11953, N11949, N9551);
nor NOR2 (N11954, N11950, N9782);
or OR4 (N11955, N11939, N6107, N2434, N6335);
xor XOR2 (N11956, N11951, N5740);
nand NAND2 (N11957, N11954, N2501);
nor NOR2 (N11958, N11942, N10010);
or OR3 (N11959, N11958, N4075, N8295);
and AND3 (N11960, N11956, N10996, N7338);
or OR3 (N11961, N11959, N1322, N1646);
or OR3 (N11962, N11952, N10179, N11855);
and AND3 (N11963, N11961, N1528, N1049);
xor XOR2 (N11964, N11960, N6055);
or OR3 (N11965, N11955, N8392, N3668);
xor XOR2 (N11966, N11957, N1434);
nand NAND2 (N11967, N11948, N4374);
nor NOR3 (N11968, N11932, N11821, N8270);
nand NAND3 (N11969, N11962, N8296, N11573);
xor XOR2 (N11970, N11934, N7759);
nand NAND2 (N11971, N11966, N3962);
nor NOR4 (N11972, N11945, N9781, N7910, N1932);
or OR3 (N11973, N11970, N7839, N3271);
buf BUF1 (N11974, N11967);
and AND2 (N11975, N11969, N11706);
not NOT1 (N11976, N11973);
and AND2 (N11977, N11975, N11820);
xor XOR2 (N11978, N11964, N1690);
and AND3 (N11979, N11972, N6972, N2953);
or OR2 (N11980, N11953, N5781);
and AND2 (N11981, N11979, N9916);
not NOT1 (N11982, N11965);
not NOT1 (N11983, N11977);
or OR3 (N11984, N11978, N1768, N4677);
buf BUF1 (N11985, N11982);
xor XOR2 (N11986, N11968, N1562);
not NOT1 (N11987, N11963);
or OR2 (N11988, N11976, N9201);
and AND2 (N11989, N11981, N11680);
buf BUF1 (N11990, N11980);
and AND2 (N11991, N11974, N10262);
nand NAND4 (N11992, N11985, N6501, N2111, N11188);
xor XOR2 (N11993, N11984, N1352);
buf BUF1 (N11994, N11993);
not NOT1 (N11995, N11992);
and AND4 (N11996, N11986, N7692, N11141, N9123);
not NOT1 (N11997, N11994);
and AND3 (N11998, N11971, N6447, N11476);
or OR3 (N11999, N11988, N2944, N3865);
nand NAND4 (N12000, N11998, N4422, N3754, N966);
not NOT1 (N12001, N11991);
buf BUF1 (N12002, N12001);
nor NOR4 (N12003, N11983, N9015, N808, N1312);
nor NOR3 (N12004, N11997, N3684, N11468);
buf BUF1 (N12005, N11995);
nand NAND2 (N12006, N11999, N8419);
or OR2 (N12007, N12002, N11186);
not NOT1 (N12008, N12004);
nand NAND4 (N12009, N11987, N4141, N8772, N10737);
xor XOR2 (N12010, N12006, N4043);
nand NAND2 (N12011, N12005, N9101);
buf BUF1 (N12012, N12007);
or OR4 (N12013, N12011, N8434, N9328, N3136);
nor NOR4 (N12014, N11990, N1926, N9861, N1885);
and AND4 (N12015, N12014, N10150, N2069, N2634);
xor XOR2 (N12016, N12010, N10590);
nand NAND3 (N12017, N12016, N8552, N5680);
nand NAND3 (N12018, N11989, N10657, N4223);
nand NAND2 (N12019, N12013, N11330);
xor XOR2 (N12020, N12015, N7705);
nand NAND3 (N12021, N12008, N6960, N4946);
not NOT1 (N12022, N12017);
buf BUF1 (N12023, N12018);
xor XOR2 (N12024, N11996, N3798);
xor XOR2 (N12025, N12022, N3180);
not NOT1 (N12026, N12012);
nor NOR2 (N12027, N12009, N2946);
not NOT1 (N12028, N12023);
nand NAND3 (N12029, N12020, N1678, N10194);
not NOT1 (N12030, N12019);
nand NAND3 (N12031, N12025, N7333, N5993);
not NOT1 (N12032, N12003);
xor XOR2 (N12033, N12028, N332);
not NOT1 (N12034, N12032);
and AND3 (N12035, N12000, N10920, N7359);
or OR3 (N12036, N12033, N1158, N5812);
and AND2 (N12037, N12021, N7425);
not NOT1 (N12038, N12035);
or OR4 (N12039, N12029, N2973, N8755, N9955);
and AND4 (N12040, N12037, N3626, N10539, N9784);
or OR2 (N12041, N12026, N10264);
not NOT1 (N12042, N12038);
and AND3 (N12043, N12041, N6732, N6073);
buf BUF1 (N12044, N12027);
not NOT1 (N12045, N12031);
and AND2 (N12046, N12024, N9466);
xor XOR2 (N12047, N12045, N1237);
or OR4 (N12048, N12034, N5411, N7955, N2798);
nor NOR2 (N12049, N12043, N180);
or OR4 (N12050, N12040, N6969, N6466, N2094);
and AND3 (N12051, N12046, N4360, N7872);
or OR4 (N12052, N12049, N2085, N7502, N10659);
and AND2 (N12053, N12039, N1027);
not NOT1 (N12054, N12030);
not NOT1 (N12055, N12052);
buf BUF1 (N12056, N12051);
nand NAND3 (N12057, N12036, N9114, N942);
nand NAND3 (N12058, N12055, N5003, N10445);
buf BUF1 (N12059, N12054);
not NOT1 (N12060, N12058);
or OR2 (N12061, N12060, N9244);
not NOT1 (N12062, N12056);
not NOT1 (N12063, N12062);
or OR3 (N12064, N12042, N253, N846);
buf BUF1 (N12065, N12061);
xor XOR2 (N12066, N12057, N7786);
buf BUF1 (N12067, N12064);
nand NAND3 (N12068, N12065, N4310, N1929);
xor XOR2 (N12069, N12053, N3736);
nor NOR3 (N12070, N12047, N2961, N11468);
nor NOR4 (N12071, N12070, N534, N9101, N1775);
not NOT1 (N12072, N12044);
nor NOR2 (N12073, N12067, N2785);
nor NOR3 (N12074, N12059, N5803, N6861);
not NOT1 (N12075, N12072);
nand NAND4 (N12076, N12073, N4797, N9658, N2835);
not NOT1 (N12077, N12048);
and AND4 (N12078, N12076, N2815, N1382, N9258);
nor NOR4 (N12079, N12071, N2577, N7711, N630);
buf BUF1 (N12080, N12069);
nor NOR2 (N12081, N12079, N8000);
buf BUF1 (N12082, N12081);
nor NOR2 (N12083, N12050, N5934);
nor NOR4 (N12084, N12066, N1501, N11000, N6422);
nand NAND4 (N12085, N12074, N612, N6661, N7719);
buf BUF1 (N12086, N12077);
buf BUF1 (N12087, N12082);
not NOT1 (N12088, N12086);
buf BUF1 (N12089, N12063);
or OR4 (N12090, N12085, N5943, N10282, N8071);
nor NOR3 (N12091, N12090, N8578, N8766);
nor NOR3 (N12092, N12078, N11137, N2081);
and AND2 (N12093, N12091, N7116);
nand NAND3 (N12094, N12087, N5375, N6392);
and AND4 (N12095, N12089, N1404, N6400, N7191);
xor XOR2 (N12096, N12084, N9140);
nand NAND3 (N12097, N12080, N4151, N1728);
and AND3 (N12098, N12095, N9571, N7240);
and AND2 (N12099, N12088, N1955);
xor XOR2 (N12100, N12075, N8122);
buf BUF1 (N12101, N12092);
buf BUF1 (N12102, N12097);
not NOT1 (N12103, N12068);
or OR3 (N12104, N12093, N9343, N777);
or OR4 (N12105, N12083, N11369, N3881, N2693);
not NOT1 (N12106, N12103);
or OR3 (N12107, N12094, N10495, N1066);
nor NOR4 (N12108, N12098, N11194, N5562, N4642);
and AND3 (N12109, N12096, N9021, N4053);
and AND2 (N12110, N12102, N11123);
nand NAND2 (N12111, N12109, N10642);
nand NAND2 (N12112, N12101, N5982);
xor XOR2 (N12113, N12105, N4932);
not NOT1 (N12114, N12104);
not NOT1 (N12115, N12108);
or OR2 (N12116, N12114, N2022);
buf BUF1 (N12117, N12111);
or OR3 (N12118, N12106, N2655, N6356);
not NOT1 (N12119, N12117);
nand NAND4 (N12120, N12116, N5870, N10245, N10957);
nand NAND4 (N12121, N12119, N8456, N125, N7191);
and AND2 (N12122, N12121, N228);
not NOT1 (N12123, N12113);
nand NAND2 (N12124, N12100, N9776);
not NOT1 (N12125, N12099);
nor NOR3 (N12126, N12110, N808, N11180);
and AND4 (N12127, N12115, N10444, N9341, N454);
or OR3 (N12128, N12127, N2435, N3659);
xor XOR2 (N12129, N12126, N3476);
xor XOR2 (N12130, N12125, N797);
nor NOR3 (N12131, N12128, N1470, N6015);
or OR2 (N12132, N12112, N9989);
not NOT1 (N12133, N12129);
buf BUF1 (N12134, N12118);
not NOT1 (N12135, N12134);
xor XOR2 (N12136, N12124, N3511);
buf BUF1 (N12137, N12123);
buf BUF1 (N12138, N12107);
not NOT1 (N12139, N12133);
and AND2 (N12140, N12122, N6559);
nor NOR2 (N12141, N12139, N6293);
buf BUF1 (N12142, N12120);
not NOT1 (N12143, N12130);
not NOT1 (N12144, N12142);
and AND3 (N12145, N12140, N5142, N10397);
nand NAND4 (N12146, N12136, N11148, N3506, N7522);
not NOT1 (N12147, N12143);
or OR2 (N12148, N12135, N4914);
nor NOR2 (N12149, N12146, N2831);
not NOT1 (N12150, N12144);
not NOT1 (N12151, N12145);
and AND2 (N12152, N12147, N771);
or OR4 (N12153, N12141, N8932, N10250, N5612);
and AND2 (N12154, N12131, N10834);
not NOT1 (N12155, N12153);
and AND3 (N12156, N12150, N7732, N5303);
not NOT1 (N12157, N12148);
nor NOR3 (N12158, N12151, N6073, N8508);
or OR4 (N12159, N12152, N10829, N2414, N10720);
or OR3 (N12160, N12159, N3981, N2250);
not NOT1 (N12161, N12138);
buf BUF1 (N12162, N12155);
not NOT1 (N12163, N12161);
nor NOR2 (N12164, N12149, N3508);
nor NOR4 (N12165, N12156, N12119, N11642, N8429);
buf BUF1 (N12166, N12137);
and AND2 (N12167, N12157, N5071);
or OR3 (N12168, N12160, N12055, N6446);
xor XOR2 (N12169, N12163, N8127);
or OR2 (N12170, N12132, N8659);
xor XOR2 (N12171, N12165, N10946);
or OR2 (N12172, N12164, N2177);
buf BUF1 (N12173, N12169);
or OR4 (N12174, N12166, N5061, N8905, N11063);
nand NAND4 (N12175, N12171, N2112, N715, N9007);
nand NAND2 (N12176, N12173, N8230);
or OR3 (N12177, N12172, N6044, N4408);
nand NAND4 (N12178, N12176, N5171, N4048, N6965);
not NOT1 (N12179, N12168);
nand NAND2 (N12180, N12162, N6234);
not NOT1 (N12181, N12158);
nor NOR4 (N12182, N12154, N4158, N7690, N6029);
and AND3 (N12183, N12175, N9306, N11545);
nor NOR3 (N12184, N12177, N647, N315);
buf BUF1 (N12185, N12170);
xor XOR2 (N12186, N12182, N1188);
and AND4 (N12187, N12174, N10117, N2086, N9285);
or OR2 (N12188, N12185, N11416);
xor XOR2 (N12189, N12187, N9299);
buf BUF1 (N12190, N12181);
or OR4 (N12191, N12167, N10935, N4901, N10871);
not NOT1 (N12192, N12186);
and AND2 (N12193, N12189, N9790);
or OR2 (N12194, N12192, N10794);
nand NAND4 (N12195, N12178, N5678, N9480, N2863);
buf BUF1 (N12196, N12184);
nand NAND4 (N12197, N12195, N8735, N10971, N11367);
xor XOR2 (N12198, N12191, N2393);
buf BUF1 (N12199, N12198);
buf BUF1 (N12200, N12196);
buf BUF1 (N12201, N12200);
xor XOR2 (N12202, N12188, N2600);
nand NAND4 (N12203, N12179, N11486, N11122, N6054);
and AND4 (N12204, N12194, N11580, N10255, N10034);
and AND3 (N12205, N12197, N7891, N8819);
and AND3 (N12206, N12204, N5807, N6194);
or OR4 (N12207, N12190, N6092, N3709, N5321);
nor NOR4 (N12208, N12183, N5493, N7887, N4926);
nor NOR4 (N12209, N12205, N2471, N10983, N2352);
not NOT1 (N12210, N12193);
buf BUF1 (N12211, N12199);
buf BUF1 (N12212, N12209);
not NOT1 (N12213, N12207);
buf BUF1 (N12214, N12203);
nor NOR3 (N12215, N12180, N9584, N10279);
and AND4 (N12216, N12215, N6293, N1319, N7699);
or OR3 (N12217, N12211, N9417, N770);
or OR4 (N12218, N12214, N7874, N1341, N4656);
nand NAND3 (N12219, N12212, N11694, N2183);
not NOT1 (N12220, N12201);
nor NOR4 (N12221, N12213, N8763, N921, N12007);
xor XOR2 (N12222, N12220, N2112);
or OR2 (N12223, N12210, N11808);
not NOT1 (N12224, N12222);
nor NOR3 (N12225, N12216, N6931, N8297);
buf BUF1 (N12226, N12217);
buf BUF1 (N12227, N12225);
and AND3 (N12228, N12219, N1552, N7373);
or OR4 (N12229, N12224, N11669, N11559, N5400);
nand NAND3 (N12230, N12223, N6936, N11334);
or OR2 (N12231, N12221, N9031);
buf BUF1 (N12232, N12227);
and AND3 (N12233, N12226, N264, N5443);
xor XOR2 (N12234, N12202, N10664);
or OR2 (N12235, N12230, N6969);
or OR2 (N12236, N12229, N8353);
nand NAND4 (N12237, N12232, N4304, N5814, N9545);
xor XOR2 (N12238, N12228, N934);
nand NAND3 (N12239, N12235, N36, N7331);
not NOT1 (N12240, N12233);
xor XOR2 (N12241, N12239, N447);
or OR3 (N12242, N12234, N9665, N8151);
buf BUF1 (N12243, N12238);
not NOT1 (N12244, N12206);
or OR2 (N12245, N12208, N6138);
xor XOR2 (N12246, N12242, N1847);
nor NOR4 (N12247, N12245, N6425, N931, N8551);
or OR2 (N12248, N12244, N5599);
buf BUF1 (N12249, N12231);
xor XOR2 (N12250, N12240, N481);
buf BUF1 (N12251, N12248);
nor NOR2 (N12252, N12243, N262);
nor NOR3 (N12253, N12252, N808, N7840);
and AND2 (N12254, N12251, N6019);
buf BUF1 (N12255, N12253);
nor NOR4 (N12256, N12249, N7805, N2970, N6528);
buf BUF1 (N12257, N12237);
nor NOR2 (N12258, N12254, N11288);
not NOT1 (N12259, N12256);
nor NOR2 (N12260, N12246, N2789);
nand NAND3 (N12261, N12250, N8729, N739);
nor NOR2 (N12262, N12236, N7512);
nand NAND3 (N12263, N12258, N7860, N4013);
not NOT1 (N12264, N12263);
and AND3 (N12265, N12218, N7900, N4156);
and AND2 (N12266, N12247, N9182);
and AND3 (N12267, N12259, N9838, N3838);
nand NAND2 (N12268, N12262, N4868);
nor NOR4 (N12269, N12260, N3845, N1117, N1827);
or OR2 (N12270, N12261, N11700);
not NOT1 (N12271, N12270);
nor NOR2 (N12272, N12271, N459);
and AND2 (N12273, N12269, N5127);
not NOT1 (N12274, N12272);
nor NOR4 (N12275, N12273, N6819, N1458, N7483);
buf BUF1 (N12276, N12274);
nor NOR3 (N12277, N12257, N6979, N8687);
nor NOR3 (N12278, N12267, N9428, N324);
nor NOR3 (N12279, N12278, N6165, N1619);
and AND3 (N12280, N12279, N4869, N8404);
buf BUF1 (N12281, N12241);
xor XOR2 (N12282, N12277, N6251);
xor XOR2 (N12283, N12268, N4754);
or OR2 (N12284, N12255, N6214);
or OR2 (N12285, N12281, N4001);
nor NOR4 (N12286, N12264, N2587, N7691, N4987);
or OR3 (N12287, N12265, N994, N5861);
and AND3 (N12288, N12276, N4986, N10910);
and AND3 (N12289, N12266, N1519, N8611);
and AND3 (N12290, N12288, N10872, N4783);
or OR3 (N12291, N12290, N1124, N346);
or OR4 (N12292, N12275, N10590, N10478, N11205);
nand NAND2 (N12293, N12284, N7307);
or OR4 (N12294, N12293, N11785, N2013, N9552);
buf BUF1 (N12295, N12292);
nor NOR4 (N12296, N12282, N3123, N5146, N6248);
not NOT1 (N12297, N12289);
not NOT1 (N12298, N12285);
nor NOR2 (N12299, N12283, N11590);
buf BUF1 (N12300, N12280);
nor NOR2 (N12301, N12295, N11065);
xor XOR2 (N12302, N12298, N1716);
buf BUF1 (N12303, N12286);
nor NOR2 (N12304, N12297, N2914);
xor XOR2 (N12305, N12304, N5752);
not NOT1 (N12306, N12291);
nand NAND2 (N12307, N12305, N332);
nand NAND3 (N12308, N12296, N9043, N2571);
buf BUF1 (N12309, N12301);
buf BUF1 (N12310, N12306);
and AND4 (N12311, N12309, N5774, N3100, N6270);
xor XOR2 (N12312, N12300, N4872);
nor NOR3 (N12313, N12308, N326, N3741);
xor XOR2 (N12314, N12307, N7192);
not NOT1 (N12315, N12312);
or OR3 (N12316, N12311, N1794, N10112);
nor NOR4 (N12317, N12315, N1201, N11269, N1298);
and AND4 (N12318, N12317, N11666, N4012, N6177);
nor NOR2 (N12319, N12302, N9325);
xor XOR2 (N12320, N12313, N8486);
xor XOR2 (N12321, N12319, N4835);
or OR3 (N12322, N12321, N1119, N6391);
nor NOR3 (N12323, N12310, N10096, N8435);
or OR2 (N12324, N12320, N251);
not NOT1 (N12325, N12287);
and AND4 (N12326, N12323, N5780, N3237, N419);
nand NAND3 (N12327, N12322, N9987, N7541);
or OR2 (N12328, N12303, N11941);
not NOT1 (N12329, N12318);
xor XOR2 (N12330, N12316, N7063);
nand NAND4 (N12331, N12324, N3268, N3032, N6993);
and AND3 (N12332, N12328, N9151, N1863);
nand NAND2 (N12333, N12326, N2272);
or OR4 (N12334, N12332, N8228, N153, N445);
nand NAND4 (N12335, N12329, N3250, N2272, N8863);
or OR2 (N12336, N12333, N2712);
nand NAND2 (N12337, N12334, N11871);
nor NOR4 (N12338, N12294, N4254, N6387, N5188);
nand NAND4 (N12339, N12314, N7224, N310, N6101);
nor NOR4 (N12340, N12339, N11627, N3950, N8790);
buf BUF1 (N12341, N12336);
buf BUF1 (N12342, N12340);
buf BUF1 (N12343, N12299);
xor XOR2 (N12344, N12342, N4206);
nand NAND3 (N12345, N12327, N2303, N3940);
buf BUF1 (N12346, N12330);
nand NAND2 (N12347, N12338, N3681);
xor XOR2 (N12348, N12325, N11148);
nor NOR4 (N12349, N12344, N10857, N7043, N1381);
buf BUF1 (N12350, N12346);
nand NAND2 (N12351, N12335, N6179);
nor NOR2 (N12352, N12351, N10479);
buf BUF1 (N12353, N12349);
xor XOR2 (N12354, N12345, N10208);
or OR3 (N12355, N12350, N3143, N7654);
and AND2 (N12356, N12348, N11666);
xor XOR2 (N12357, N12354, N7447);
not NOT1 (N12358, N12352);
and AND4 (N12359, N12357, N12335, N9509, N2368);
nand NAND3 (N12360, N12353, N311, N5413);
buf BUF1 (N12361, N12341);
nor NOR4 (N12362, N12337, N4608, N6236, N5258);
or OR4 (N12363, N12355, N8882, N6033, N6062);
and AND3 (N12364, N12360, N5291, N7425);
not NOT1 (N12365, N12364);
not NOT1 (N12366, N12365);
nor NOR4 (N12367, N12343, N3618, N8974, N7633);
or OR2 (N12368, N12363, N790);
buf BUF1 (N12369, N12356);
nor NOR3 (N12370, N12367, N2070, N7935);
and AND4 (N12371, N12362, N10613, N5665, N1801);
nor NOR3 (N12372, N12358, N11831, N7877);
nand NAND4 (N12373, N12361, N4393, N8496, N249);
nor NOR2 (N12374, N12373, N143);
not NOT1 (N12375, N12368);
and AND4 (N12376, N12372, N11895, N10843, N3352);
or OR2 (N12377, N12369, N3940);
nand NAND2 (N12378, N12376, N4961);
nor NOR4 (N12379, N12370, N2170, N2917, N2231);
not NOT1 (N12380, N12371);
xor XOR2 (N12381, N12374, N1744);
buf BUF1 (N12382, N12366);
nor NOR3 (N12383, N12347, N749, N5857);
nor NOR4 (N12384, N12377, N2985, N1139, N10110);
nor NOR2 (N12385, N12379, N7829);
nand NAND4 (N12386, N12385, N9101, N6295, N2328);
nand NAND2 (N12387, N12386, N3829);
buf BUF1 (N12388, N12384);
nor NOR4 (N12389, N12381, N1347, N7771, N12293);
nor NOR4 (N12390, N12382, N4020, N5041, N9850);
not NOT1 (N12391, N12380);
nand NAND3 (N12392, N12378, N7079, N7373);
nand NAND3 (N12393, N12387, N1838, N9538);
nor NOR2 (N12394, N12391, N1675);
not NOT1 (N12395, N12383);
nor NOR2 (N12396, N12392, N9167);
nand NAND4 (N12397, N12396, N8472, N24, N7832);
buf BUF1 (N12398, N12395);
not NOT1 (N12399, N12359);
and AND2 (N12400, N12398, N9565);
nand NAND2 (N12401, N12397, N6174);
buf BUF1 (N12402, N12389);
xor XOR2 (N12403, N12402, N4789);
and AND2 (N12404, N12388, N1552);
nor NOR4 (N12405, N12375, N8180, N12181, N3881);
xor XOR2 (N12406, N12401, N3814);
or OR4 (N12407, N12403, N10197, N11485, N6550);
nand NAND4 (N12408, N12399, N11352, N3969, N2368);
not NOT1 (N12409, N12408);
and AND4 (N12410, N12404, N6554, N7753, N6072);
xor XOR2 (N12411, N12405, N7298);
nor NOR4 (N12412, N12400, N12126, N11498, N7054);
and AND4 (N12413, N12409, N76, N12033, N1740);
nand NAND3 (N12414, N12394, N11014, N2924);
and AND3 (N12415, N12406, N8834, N10075);
or OR3 (N12416, N12412, N11208, N6394);
and AND2 (N12417, N12390, N3770);
nand NAND3 (N12418, N12416, N9221, N7215);
nor NOR2 (N12419, N12418, N203);
buf BUF1 (N12420, N12411);
not NOT1 (N12421, N12417);
and AND4 (N12422, N12421, N7678, N3901, N7950);
not NOT1 (N12423, N12407);
or OR2 (N12424, N12419, N992);
not NOT1 (N12425, N12393);
nor NOR4 (N12426, N12425, N2448, N10250, N4672);
and AND2 (N12427, N12426, N5199);
buf BUF1 (N12428, N12420);
nand NAND3 (N12429, N12410, N9929, N11221);
and AND2 (N12430, N12423, N12327);
nor NOR4 (N12431, N12428, N12299, N7642, N12138);
not NOT1 (N12432, N12424);
not NOT1 (N12433, N12422);
or OR3 (N12434, N12413, N4415, N6751);
and AND3 (N12435, N12427, N2343, N5585);
buf BUF1 (N12436, N12435);
or OR3 (N12437, N12415, N11209, N11854);
buf BUF1 (N12438, N12331);
not NOT1 (N12439, N12429);
nand NAND2 (N12440, N12436, N2066);
nand NAND4 (N12441, N12438, N4548, N5339, N2851);
not NOT1 (N12442, N12441);
buf BUF1 (N12443, N12442);
nor NOR4 (N12444, N12433, N8460, N8007, N11476);
nor NOR4 (N12445, N12443, N9604, N8709, N7173);
xor XOR2 (N12446, N12431, N6148);
or OR2 (N12447, N12430, N11912);
nand NAND2 (N12448, N12434, N10153);
nor NOR4 (N12449, N12445, N3656, N9777, N340);
nand NAND4 (N12450, N12446, N8616, N1083, N3081);
buf BUF1 (N12451, N12444);
and AND2 (N12452, N12448, N1818);
nand NAND4 (N12453, N12450, N12138, N7314, N9461);
nand NAND3 (N12454, N12432, N10065, N11267);
xor XOR2 (N12455, N12439, N2558);
or OR2 (N12456, N12451, N5683);
xor XOR2 (N12457, N12454, N6272);
buf BUF1 (N12458, N12449);
nor NOR2 (N12459, N12453, N10787);
xor XOR2 (N12460, N12437, N4491);
not NOT1 (N12461, N12459);
and AND4 (N12462, N12457, N10268, N10443, N12208);
nand NAND4 (N12463, N12414, N4054, N6320, N8192);
and AND4 (N12464, N12447, N11313, N12157, N10634);
buf BUF1 (N12465, N12456);
xor XOR2 (N12466, N12461, N4280);
not NOT1 (N12467, N12466);
nand NAND4 (N12468, N12440, N150, N8349, N6543);
not NOT1 (N12469, N12460);
or OR3 (N12470, N12462, N7036, N9099);
buf BUF1 (N12471, N12467);
nor NOR3 (N12472, N12470, N6989, N8337);
and AND2 (N12473, N12468, N10339);
xor XOR2 (N12474, N12464, N4510);
xor XOR2 (N12475, N12463, N8484);
xor XOR2 (N12476, N12452, N4176);
xor XOR2 (N12477, N12473, N10994);
nand NAND3 (N12478, N12458, N8852, N3815);
xor XOR2 (N12479, N12478, N3547);
nand NAND3 (N12480, N12475, N10109, N10229);
xor XOR2 (N12481, N12471, N6271);
and AND2 (N12482, N12481, N10951);
and AND3 (N12483, N12477, N1967, N347);
not NOT1 (N12484, N12469);
not NOT1 (N12485, N12474);
nand NAND4 (N12486, N12465, N10513, N861, N3294);
nand NAND4 (N12487, N12479, N2995, N11993, N5133);
nand NAND2 (N12488, N12484, N5998);
xor XOR2 (N12489, N12483, N445);
nand NAND3 (N12490, N12480, N11799, N4848);
xor XOR2 (N12491, N12455, N7117);
or OR2 (N12492, N12486, N8128);
xor XOR2 (N12493, N12487, N6498);
and AND2 (N12494, N12489, N11485);
not NOT1 (N12495, N12476);
nand NAND3 (N12496, N12490, N4418, N11174);
or OR2 (N12497, N12494, N468);
or OR2 (N12498, N12493, N6109);
not NOT1 (N12499, N12495);
and AND2 (N12500, N12497, N950);
not NOT1 (N12501, N12488);
or OR3 (N12502, N12501, N10189, N6412);
nand NAND4 (N12503, N12500, N4004, N8557, N988);
not NOT1 (N12504, N12491);
xor XOR2 (N12505, N12496, N2578);
nand NAND3 (N12506, N12503, N4139, N2209);
and AND2 (N12507, N12492, N11456);
nand NAND3 (N12508, N12472, N12341, N7188);
xor XOR2 (N12509, N12506, N4369);
buf BUF1 (N12510, N12504);
buf BUF1 (N12511, N12498);
or OR3 (N12512, N12508, N6823, N11147);
nand NAND4 (N12513, N12485, N11256, N3436, N6517);
and AND2 (N12514, N12499, N164);
and AND4 (N12515, N12512, N10014, N6018, N11177);
not NOT1 (N12516, N12505);
not NOT1 (N12517, N12509);
xor XOR2 (N12518, N12516, N11092);
nand NAND3 (N12519, N12510, N8623, N8746);
xor XOR2 (N12520, N12507, N5372);
nand NAND4 (N12521, N12502, N3799, N11734, N10637);
buf BUF1 (N12522, N12519);
xor XOR2 (N12523, N12482, N9702);
nand NAND3 (N12524, N12523, N11579, N11351);
nor NOR2 (N12525, N12518, N6129);
or OR4 (N12526, N12524, N2775, N10782, N4145);
nand NAND3 (N12527, N12522, N8680, N10181);
buf BUF1 (N12528, N12526);
xor XOR2 (N12529, N12521, N673);
buf BUF1 (N12530, N12525);
not NOT1 (N12531, N12514);
or OR2 (N12532, N12515, N1027);
or OR3 (N12533, N12517, N3395, N3551);
and AND2 (N12534, N12530, N7910);
buf BUF1 (N12535, N12532);
xor XOR2 (N12536, N12529, N2485);
nor NOR4 (N12537, N12534, N11772, N518, N7325);
xor XOR2 (N12538, N12528, N11112);
or OR2 (N12539, N12533, N10228);
and AND4 (N12540, N12513, N9382, N3066, N1725);
nand NAND3 (N12541, N12535, N8129, N1709);
nor NOR3 (N12542, N12538, N1849, N1256);
xor XOR2 (N12543, N12539, N12201);
buf BUF1 (N12544, N12536);
and AND2 (N12545, N12543, N6999);
or OR3 (N12546, N12520, N155, N7671);
and AND3 (N12547, N12537, N8325, N6237);
and AND3 (N12548, N12527, N3012, N614);
xor XOR2 (N12549, N12542, N11893);
nand NAND3 (N12550, N12549, N8504, N4294);
nor NOR3 (N12551, N12547, N2669, N10798);
and AND4 (N12552, N12545, N11882, N3399, N10260);
buf BUF1 (N12553, N12548);
xor XOR2 (N12554, N12541, N4963);
and AND2 (N12555, N12511, N5615);
not NOT1 (N12556, N12554);
buf BUF1 (N12557, N12556);
nor NOR2 (N12558, N12551, N5218);
nor NOR3 (N12559, N12553, N6624, N9848);
not NOT1 (N12560, N12555);
and AND2 (N12561, N12552, N7377);
and AND4 (N12562, N12550, N4105, N9612, N1663);
nor NOR3 (N12563, N12540, N10936, N12037);
nand NAND3 (N12564, N12557, N5042, N362);
nand NAND3 (N12565, N12561, N1948, N1802);
xor XOR2 (N12566, N12546, N829);
not NOT1 (N12567, N12562);
buf BUF1 (N12568, N12544);
or OR2 (N12569, N12560, N5153);
and AND3 (N12570, N12566, N2335, N10474);
xor XOR2 (N12571, N12568, N596);
and AND4 (N12572, N12563, N394, N8158, N2632);
and AND3 (N12573, N12564, N9422, N2769);
buf BUF1 (N12574, N12571);
buf BUF1 (N12575, N12565);
nand NAND4 (N12576, N12575, N4792, N9925, N1313);
nor NOR2 (N12577, N12558, N2301);
buf BUF1 (N12578, N12570);
nand NAND2 (N12579, N12577, N9552);
xor XOR2 (N12580, N12569, N7284);
not NOT1 (N12581, N12572);
and AND2 (N12582, N12574, N10024);
or OR2 (N12583, N12559, N1953);
buf BUF1 (N12584, N12583);
or OR4 (N12585, N12582, N3934, N7307, N10827);
or OR3 (N12586, N12578, N9896, N6973);
xor XOR2 (N12587, N12531, N11010);
and AND3 (N12588, N12580, N1321, N10589);
buf BUF1 (N12589, N12581);
nand NAND3 (N12590, N12584, N11760, N3664);
and AND3 (N12591, N12590, N11862, N9369);
xor XOR2 (N12592, N12591, N769);
or OR4 (N12593, N12567, N2324, N1899, N10885);
nor NOR3 (N12594, N12586, N11153, N3330);
not NOT1 (N12595, N12579);
buf BUF1 (N12596, N12589);
buf BUF1 (N12597, N12576);
and AND3 (N12598, N12585, N2370, N1617);
or OR3 (N12599, N12598, N3206, N11007);
nand NAND2 (N12600, N12594, N2832);
nand NAND3 (N12601, N12596, N5598, N9410);
xor XOR2 (N12602, N12592, N3844);
nor NOR2 (N12603, N12573, N6910);
or OR3 (N12604, N12602, N11626, N7419);
not NOT1 (N12605, N12599);
buf BUF1 (N12606, N12605);
and AND2 (N12607, N12600, N12554);
xor XOR2 (N12608, N12604, N5359);
nand NAND3 (N12609, N12593, N5474, N10403);
and AND2 (N12610, N12587, N7406);
or OR2 (N12611, N12588, N4765);
or OR2 (N12612, N12606, N4874);
nand NAND4 (N12613, N12595, N3656, N9859, N6074);
or OR4 (N12614, N12611, N4289, N2437, N10242);
not NOT1 (N12615, N12613);
nand NAND2 (N12616, N12615, N4420);
and AND3 (N12617, N12603, N5147, N752);
nor NOR3 (N12618, N12607, N8915, N12296);
and AND3 (N12619, N12597, N231, N10006);
nand NAND2 (N12620, N12614, N12057);
and AND4 (N12621, N12610, N1016, N2335, N10384);
buf BUF1 (N12622, N12601);
buf BUF1 (N12623, N12616);
or OR3 (N12624, N12608, N1408, N7588);
buf BUF1 (N12625, N12609);
buf BUF1 (N12626, N12618);
xor XOR2 (N12627, N12617, N2265);
buf BUF1 (N12628, N12622);
or OR4 (N12629, N12628, N11334, N1515, N3930);
and AND3 (N12630, N12627, N12091, N5618);
or OR4 (N12631, N12619, N10195, N10147, N129);
and AND2 (N12632, N12623, N1908);
xor XOR2 (N12633, N12631, N11555);
xor XOR2 (N12634, N12629, N8932);
xor XOR2 (N12635, N12630, N7731);
nand NAND3 (N12636, N12632, N8060, N6256);
xor XOR2 (N12637, N12626, N8250);
nor NOR2 (N12638, N12637, N3385);
and AND3 (N12639, N12634, N3910, N3196);
nand NAND3 (N12640, N12633, N3617, N541);
not NOT1 (N12641, N12639);
nand NAND4 (N12642, N12635, N3284, N1598, N3166);
buf BUF1 (N12643, N12624);
xor XOR2 (N12644, N12621, N565);
nor NOR2 (N12645, N12636, N11549);
not NOT1 (N12646, N12612);
xor XOR2 (N12647, N12641, N2910);
buf BUF1 (N12648, N12642);
buf BUF1 (N12649, N12645);
xor XOR2 (N12650, N12647, N3164);
or OR2 (N12651, N12638, N10115);
or OR3 (N12652, N12643, N1095, N6919);
xor XOR2 (N12653, N12625, N2565);
xor XOR2 (N12654, N12652, N5463);
not NOT1 (N12655, N12653);
and AND3 (N12656, N12655, N4855, N8531);
buf BUF1 (N12657, N12646);
or OR3 (N12658, N12648, N11821, N12261);
nand NAND2 (N12659, N12644, N11205);
nor NOR3 (N12660, N12656, N10996, N9995);
xor XOR2 (N12661, N12657, N9529);
or OR3 (N12662, N12654, N7486, N12408);
and AND2 (N12663, N12660, N6094);
nor NOR3 (N12664, N12661, N7628, N12421);
and AND2 (N12665, N12658, N9907);
nor NOR2 (N12666, N12649, N550);
xor XOR2 (N12667, N12663, N1921);
nand NAND4 (N12668, N12620, N418, N305, N1243);
nand NAND3 (N12669, N12664, N2084, N9419);
nand NAND3 (N12670, N12650, N10985, N11489);
nor NOR4 (N12671, N12659, N7461, N3382, N5334);
nor NOR3 (N12672, N12671, N1851, N8409);
xor XOR2 (N12673, N12640, N1939);
nor NOR4 (N12674, N12673, N12200, N11197, N7689);
and AND4 (N12675, N12670, N794, N1105, N7017);
not NOT1 (N12676, N12668);
nor NOR4 (N12677, N12662, N3158, N1690, N2303);
nand NAND3 (N12678, N12672, N6471, N4341);
or OR4 (N12679, N12651, N11675, N1968, N11438);
buf BUF1 (N12680, N12677);
nor NOR4 (N12681, N12665, N10200, N11674, N8356);
nand NAND3 (N12682, N12679, N9578, N1862);
nand NAND3 (N12683, N12674, N11669, N12193);
buf BUF1 (N12684, N12678);
nor NOR4 (N12685, N12682, N6048, N2017, N10837);
buf BUF1 (N12686, N12684);
and AND4 (N12687, N12676, N6161, N7228, N11820);
not NOT1 (N12688, N12686);
nand NAND4 (N12689, N12667, N9130, N7006, N1441);
nand NAND4 (N12690, N12689, N5922, N10545, N5691);
and AND2 (N12691, N12685, N6921);
xor XOR2 (N12692, N12675, N6418);
xor XOR2 (N12693, N12688, N2015);
or OR4 (N12694, N12666, N3816, N11038, N4830);
and AND2 (N12695, N12693, N11880);
xor XOR2 (N12696, N12687, N10549);
buf BUF1 (N12697, N12681);
not NOT1 (N12698, N12691);
and AND4 (N12699, N12697, N4910, N7789, N7485);
buf BUF1 (N12700, N12669);
and AND4 (N12701, N12695, N10789, N8236, N5622);
buf BUF1 (N12702, N12701);
nand NAND4 (N12703, N12702, N11879, N6271, N5718);
buf BUF1 (N12704, N12703);
not NOT1 (N12705, N12694);
nand NAND4 (N12706, N12698, N1627, N6020, N11979);
buf BUF1 (N12707, N12700);
nand NAND4 (N12708, N12705, N10947, N9101, N4617);
and AND4 (N12709, N12706, N905, N5618, N152);
buf BUF1 (N12710, N12696);
buf BUF1 (N12711, N12680);
and AND3 (N12712, N12708, N4485, N8970);
nand NAND3 (N12713, N12699, N376, N11899);
nand NAND2 (N12714, N12690, N4782);
and AND3 (N12715, N12692, N8873, N5804);
not NOT1 (N12716, N12715);
buf BUF1 (N12717, N12704);
buf BUF1 (N12718, N12713);
not NOT1 (N12719, N12716);
and AND3 (N12720, N12719, N2423, N11713);
buf BUF1 (N12721, N12718);
or OR4 (N12722, N12711, N8054, N10170, N12117);
buf BUF1 (N12723, N12720);
or OR3 (N12724, N12722, N8057, N5577);
not NOT1 (N12725, N12710);
not NOT1 (N12726, N12725);
nand NAND2 (N12727, N12712, N5372);
or OR3 (N12728, N12724, N9528, N762);
or OR3 (N12729, N12709, N12684, N4320);
or OR3 (N12730, N12723, N11151, N2745);
nor NOR2 (N12731, N12727, N10804);
nor NOR2 (N12732, N12714, N6026);
xor XOR2 (N12733, N12732, N4180);
xor XOR2 (N12734, N12683, N174);
nand NAND4 (N12735, N12731, N3074, N7976, N3745);
not NOT1 (N12736, N12730);
buf BUF1 (N12737, N12726);
and AND2 (N12738, N12717, N4174);
nor NOR4 (N12739, N12737, N3937, N9387, N10211);
and AND2 (N12740, N12734, N11255);
xor XOR2 (N12741, N12733, N9274);
nor NOR3 (N12742, N12739, N8108, N10224);
or OR2 (N12743, N12742, N3918);
and AND4 (N12744, N12743, N1470, N11414, N11388);
buf BUF1 (N12745, N12728);
xor XOR2 (N12746, N12741, N4695);
buf BUF1 (N12747, N12707);
not NOT1 (N12748, N12744);
or OR3 (N12749, N12748, N8279, N5051);
not NOT1 (N12750, N12747);
not NOT1 (N12751, N12735);
and AND2 (N12752, N12729, N11754);
nand NAND2 (N12753, N12738, N3181);
nand NAND3 (N12754, N12753, N6478, N7134);
and AND4 (N12755, N12752, N1007, N5666, N3297);
and AND4 (N12756, N12750, N6191, N10395, N3316);
or OR4 (N12757, N12721, N3915, N11663, N3243);
or OR4 (N12758, N12745, N3477, N10276, N3245);
not NOT1 (N12759, N12749);
nand NAND2 (N12760, N12759, N9678);
buf BUF1 (N12761, N12760);
nand NAND3 (N12762, N12761, N11046, N1023);
not NOT1 (N12763, N12754);
nor NOR3 (N12764, N12757, N10229, N9865);
or OR4 (N12765, N12751, N3060, N3217, N5706);
xor XOR2 (N12766, N12765, N5091);
not NOT1 (N12767, N12740);
buf BUF1 (N12768, N12756);
nand NAND4 (N12769, N12755, N567, N3927, N12037);
xor XOR2 (N12770, N12762, N4394);
or OR2 (N12771, N12736, N11269);
nor NOR3 (N12772, N12769, N875, N6294);
nor NOR3 (N12773, N12746, N10129, N7853);
not NOT1 (N12774, N12764);
and AND4 (N12775, N12766, N5205, N6085, N1270);
not NOT1 (N12776, N12770);
nand NAND3 (N12777, N12763, N9634, N622);
xor XOR2 (N12778, N12772, N4965);
not NOT1 (N12779, N12777);
buf BUF1 (N12780, N12758);
xor XOR2 (N12781, N12776, N553);
or OR3 (N12782, N12773, N12122, N5384);
nand NAND4 (N12783, N12768, N11102, N1532, N8355);
and AND2 (N12784, N12775, N578);
or OR4 (N12785, N12767, N10840, N5925, N8681);
nor NOR4 (N12786, N12783, N451, N3631, N3537);
or OR4 (N12787, N12781, N9420, N5651, N6824);
nand NAND4 (N12788, N12774, N3312, N8299, N4640);
and AND4 (N12789, N12780, N10132, N10451, N7268);
not NOT1 (N12790, N12778);
nand NAND3 (N12791, N12790, N3598, N2703);
xor XOR2 (N12792, N12791, N9445);
or OR3 (N12793, N12779, N6329, N8864);
or OR2 (N12794, N12793, N5289);
buf BUF1 (N12795, N12794);
and AND3 (N12796, N12788, N3364, N2886);
not NOT1 (N12797, N12771);
xor XOR2 (N12798, N12797, N11660);
not NOT1 (N12799, N12785);
xor XOR2 (N12800, N12795, N3007);
and AND4 (N12801, N12798, N9619, N1598, N9178);
xor XOR2 (N12802, N12792, N4488);
nor NOR4 (N12803, N12799, N896, N2734, N3100);
nor NOR2 (N12804, N12786, N7491);
or OR2 (N12805, N12787, N11072);
nand NAND4 (N12806, N12803, N11053, N2644, N281);
xor XOR2 (N12807, N12806, N7186);
nand NAND4 (N12808, N12784, N2673, N4896, N10656);
nand NAND2 (N12809, N12796, N3573);
xor XOR2 (N12810, N12805, N12516);
nor NOR3 (N12811, N12809, N7916, N8116);
nor NOR2 (N12812, N12802, N4814);
not NOT1 (N12813, N12789);
or OR3 (N12814, N12801, N10912, N7748);
xor XOR2 (N12815, N12804, N10911);
or OR3 (N12816, N12812, N7635, N8177);
xor XOR2 (N12817, N12813, N7969);
and AND4 (N12818, N12807, N10691, N9701, N5251);
nor NOR4 (N12819, N12818, N4339, N9237, N11860);
nand NAND3 (N12820, N12800, N11789, N977);
and AND2 (N12821, N12819, N5322);
buf BUF1 (N12822, N12821);
buf BUF1 (N12823, N12817);
nand NAND4 (N12824, N12810, N6282, N11220, N1919);
or OR3 (N12825, N12824, N272, N11173);
or OR3 (N12826, N12814, N2321, N9987);
not NOT1 (N12827, N12823);
and AND2 (N12828, N12811, N5332);
nand NAND4 (N12829, N12816, N10069, N1082, N6494);
nor NOR3 (N12830, N12826, N7489, N12196);
nand NAND2 (N12831, N12820, N5788);
or OR4 (N12832, N12829, N33, N3641, N5755);
nor NOR2 (N12833, N12815, N5085);
not NOT1 (N12834, N12833);
and AND2 (N12835, N12822, N4702);
xor XOR2 (N12836, N12825, N2664);
nand NAND2 (N12837, N12782, N11437);
nand NAND4 (N12838, N12834, N6430, N3299, N10442);
not NOT1 (N12839, N12830);
xor XOR2 (N12840, N12836, N12009);
not NOT1 (N12841, N12828);
nor NOR4 (N12842, N12827, N9853, N11741, N418);
nand NAND2 (N12843, N12842, N12710);
not NOT1 (N12844, N12843);
or OR2 (N12845, N12838, N12112);
or OR3 (N12846, N12831, N7598, N211);
xor XOR2 (N12847, N12832, N9632);
and AND3 (N12848, N12839, N12280, N7034);
xor XOR2 (N12849, N12846, N11755);
and AND4 (N12850, N12808, N3922, N7914, N5066);
not NOT1 (N12851, N12841);
xor XOR2 (N12852, N12844, N282);
or OR2 (N12853, N12835, N10617);
xor XOR2 (N12854, N12851, N106);
nand NAND2 (N12855, N12853, N10815);
and AND2 (N12856, N12848, N9607);
buf BUF1 (N12857, N12849);
or OR2 (N12858, N12840, N7248);
and AND3 (N12859, N12855, N12287, N7247);
buf BUF1 (N12860, N12854);
or OR4 (N12861, N12858, N1698, N12157, N8416);
nand NAND3 (N12862, N12850, N11787, N3760);
buf BUF1 (N12863, N12847);
or OR2 (N12864, N12860, N3532);
and AND2 (N12865, N12863, N5563);
buf BUF1 (N12866, N12861);
nor NOR3 (N12867, N12866, N3511, N5964);
xor XOR2 (N12868, N12857, N3487);
or OR4 (N12869, N12868, N8438, N10005, N11859);
not NOT1 (N12870, N12867);
or OR2 (N12871, N12865, N10540);
or OR3 (N12872, N12864, N3570, N2857);
and AND3 (N12873, N12869, N8611, N4128);
not NOT1 (N12874, N12870);
nand NAND4 (N12875, N12856, N7577, N3191, N8920);
and AND4 (N12876, N12871, N11224, N4121, N12775);
nor NOR2 (N12877, N12872, N10287);
or OR4 (N12878, N12876, N6970, N805, N5537);
and AND4 (N12879, N12874, N4974, N4572, N4499);
buf BUF1 (N12880, N12875);
buf BUF1 (N12881, N12852);
and AND3 (N12882, N12878, N1615, N9435);
xor XOR2 (N12883, N12877, N12568);
not NOT1 (N12884, N12862);
xor XOR2 (N12885, N12884, N11756);
nor NOR2 (N12886, N12837, N4604);
nand NAND4 (N12887, N12885, N2874, N3741, N7450);
buf BUF1 (N12888, N12859);
xor XOR2 (N12889, N12887, N4880);
not NOT1 (N12890, N12888);
xor XOR2 (N12891, N12880, N12137);
and AND3 (N12892, N12890, N6281, N3641);
nand NAND4 (N12893, N12891, N27, N5049, N8539);
buf BUF1 (N12894, N12889);
not NOT1 (N12895, N12873);
not NOT1 (N12896, N12895);
or OR3 (N12897, N12893, N145, N7510);
and AND3 (N12898, N12892, N1919, N12436);
and AND2 (N12899, N12898, N12613);
and AND2 (N12900, N12899, N10924);
not NOT1 (N12901, N12886);
xor XOR2 (N12902, N12879, N6097);
xor XOR2 (N12903, N12900, N12608);
nand NAND3 (N12904, N12902, N12287, N4598);
xor XOR2 (N12905, N12883, N10026);
nor NOR3 (N12906, N12896, N3195, N2745);
and AND4 (N12907, N12901, N8269, N5760, N10669);
nor NOR4 (N12908, N12904, N7888, N10586, N4755);
not NOT1 (N12909, N12907);
xor XOR2 (N12910, N12909, N5563);
xor XOR2 (N12911, N12905, N1968);
or OR4 (N12912, N12908, N9257, N10180, N5105);
and AND4 (N12913, N12906, N10222, N4146, N10887);
or OR3 (N12914, N12910, N9837, N3641);
and AND2 (N12915, N12912, N9317);
buf BUF1 (N12916, N12897);
and AND4 (N12917, N12915, N3725, N2073, N37);
or OR4 (N12918, N12845, N1683, N8506, N12355);
nand NAND3 (N12919, N12911, N5540, N9697);
or OR3 (N12920, N12881, N12916, N1689);
xor XOR2 (N12921, N4492, N12744);
buf BUF1 (N12922, N12913);
or OR4 (N12923, N12882, N2842, N8562, N2244);
not NOT1 (N12924, N12922);
xor XOR2 (N12925, N12923, N9253);
not NOT1 (N12926, N12919);
and AND3 (N12927, N12894, N3754, N9973);
nor NOR4 (N12928, N12920, N8010, N507, N5371);
buf BUF1 (N12929, N12903);
and AND4 (N12930, N12918, N10556, N1663, N12426);
and AND2 (N12931, N12914, N3658);
xor XOR2 (N12932, N12930, N6662);
nand NAND2 (N12933, N12926, N10095);
not NOT1 (N12934, N12931);
xor XOR2 (N12935, N12934, N8832);
not NOT1 (N12936, N12935);
or OR2 (N12937, N12928, N10181);
buf BUF1 (N12938, N12925);
nand NAND4 (N12939, N12936, N5192, N4232, N9727);
buf BUF1 (N12940, N12929);
or OR4 (N12941, N12917, N7631, N40, N9341);
xor XOR2 (N12942, N12932, N7691);
nand NAND2 (N12943, N12938, N6480);
not NOT1 (N12944, N12940);
nand NAND4 (N12945, N12924, N8010, N8813, N7421);
and AND2 (N12946, N12945, N1723);
buf BUF1 (N12947, N12921);
nand NAND3 (N12948, N12927, N8691, N1895);
nor NOR4 (N12949, N12943, N5074, N12149, N5800);
buf BUF1 (N12950, N12946);
nor NOR4 (N12951, N12947, N6736, N9743, N7676);
xor XOR2 (N12952, N12948, N11652);
buf BUF1 (N12953, N12933);
nand NAND3 (N12954, N12950, N8786, N8086);
not NOT1 (N12955, N12951);
buf BUF1 (N12956, N12949);
buf BUF1 (N12957, N12942);
nor NOR4 (N12958, N12957, N8256, N7162, N3120);
nand NAND4 (N12959, N12953, N914, N288, N1792);
buf BUF1 (N12960, N12937);
nand NAND4 (N12961, N12960, N3110, N6323, N3142);
buf BUF1 (N12962, N12956);
buf BUF1 (N12963, N12962);
not NOT1 (N12964, N12959);
and AND4 (N12965, N12961, N11570, N7716, N10591);
not NOT1 (N12966, N12954);
buf BUF1 (N12967, N12952);
nand NAND2 (N12968, N12939, N4813);
buf BUF1 (N12969, N12964);
xor XOR2 (N12970, N12963, N12394);
xor XOR2 (N12971, N12941, N1131);
and AND3 (N12972, N12968, N6487, N6967);
buf BUF1 (N12973, N12969);
nor NOR3 (N12974, N12958, N8271, N7889);
buf BUF1 (N12975, N12966);
nand NAND2 (N12976, N12974, N3436);
buf BUF1 (N12977, N12965);
xor XOR2 (N12978, N12977, N1669);
or OR3 (N12979, N12967, N7150, N2385);
nand NAND3 (N12980, N12976, N5467, N6146);
not NOT1 (N12981, N12970);
or OR4 (N12982, N12981, N12712, N6062, N11216);
or OR3 (N12983, N12979, N5083, N5770);
and AND2 (N12984, N12980, N4023);
xor XOR2 (N12985, N12971, N8859);
and AND2 (N12986, N12955, N6061);
xor XOR2 (N12987, N12985, N9456);
and AND4 (N12988, N12982, N12344, N4743, N11262);
buf BUF1 (N12989, N12984);
and AND4 (N12990, N12987, N4696, N4833, N12315);
xor XOR2 (N12991, N12986, N12224);
xor XOR2 (N12992, N12990, N2372);
nand NAND3 (N12993, N12992, N6633, N211);
buf BUF1 (N12994, N12983);
or OR3 (N12995, N12973, N10252, N8644);
or OR2 (N12996, N12988, N11212);
and AND2 (N12997, N12994, N2070);
and AND4 (N12998, N12972, N10436, N8617, N3034);
not NOT1 (N12999, N12991);
not NOT1 (N13000, N12998);
xor XOR2 (N13001, N12978, N4105);
and AND2 (N13002, N12996, N9933);
xor XOR2 (N13003, N12993, N7876);
nand NAND2 (N13004, N13002, N6245);
or OR3 (N13005, N13000, N7440, N11350);
nand NAND2 (N13006, N13005, N5398);
nand NAND4 (N13007, N13004, N10986, N7371, N4773);
xor XOR2 (N13008, N12975, N12626);
xor XOR2 (N13009, N13001, N2407);
buf BUF1 (N13010, N13008);
buf BUF1 (N13011, N12989);
not NOT1 (N13012, N13011);
nand NAND3 (N13013, N13003, N11208, N12049);
buf BUF1 (N13014, N12999);
or OR2 (N13015, N13009, N3413);
nand NAND2 (N13016, N13013, N4576);
not NOT1 (N13017, N12944);
nor NOR3 (N13018, N13007, N477, N11835);
nand NAND2 (N13019, N13015, N6739);
and AND3 (N13020, N13017, N10432, N8549);
xor XOR2 (N13021, N13016, N6962);
buf BUF1 (N13022, N13019);
nor NOR3 (N13023, N13021, N11558, N2061);
and AND4 (N13024, N13010, N3146, N9671, N2815);
or OR3 (N13025, N13012, N11636, N9677);
nand NAND4 (N13026, N12995, N4172, N1698, N10405);
or OR2 (N13027, N13024, N1715);
buf BUF1 (N13028, N13025);
or OR2 (N13029, N13026, N5838);
xor XOR2 (N13030, N12997, N4213);
xor XOR2 (N13031, N13028, N10075);
or OR3 (N13032, N13006, N8295, N138);
buf BUF1 (N13033, N13029);
nand NAND2 (N13034, N13020, N8505);
xor XOR2 (N13035, N13027, N12691);
nand NAND3 (N13036, N13023, N1863, N5477);
and AND4 (N13037, N13035, N7084, N4108, N10318);
nand NAND4 (N13038, N13037, N4737, N7621, N7567);
nand NAND3 (N13039, N13018, N7376, N2098);
and AND3 (N13040, N13034, N6655, N6573);
not NOT1 (N13041, N13022);
not NOT1 (N13042, N13030);
buf BUF1 (N13043, N13031);
or OR4 (N13044, N13014, N11647, N7744, N11944);
buf BUF1 (N13045, N13044);
xor XOR2 (N13046, N13040, N10137);
or OR2 (N13047, N13045, N2749);
and AND2 (N13048, N13046, N4257);
or OR4 (N13049, N13038, N2196, N6906, N1313);
buf BUF1 (N13050, N13039);
buf BUF1 (N13051, N13050);
nand NAND2 (N13052, N13051, N6110);
xor XOR2 (N13053, N13049, N1337);
nor NOR3 (N13054, N13047, N10821, N6058);
nor NOR3 (N13055, N13054, N10183, N3409);
nand NAND2 (N13056, N13041, N2829);
or OR3 (N13057, N13043, N7381, N8954);
xor XOR2 (N13058, N13052, N148);
or OR4 (N13059, N13048, N10672, N1721, N4784);
and AND3 (N13060, N13058, N4594, N2869);
nand NAND4 (N13061, N13036, N8646, N931, N429);
and AND2 (N13062, N13042, N11200);
buf BUF1 (N13063, N13059);
nor NOR4 (N13064, N13055, N12452, N8124, N10671);
nor NOR3 (N13065, N13056, N9196, N3126);
nor NOR4 (N13066, N13033, N3528, N5024, N5029);
and AND3 (N13067, N13032, N7331, N9080);
nor NOR4 (N13068, N13067, N5923, N1990, N3996);
or OR2 (N13069, N13068, N7559);
xor XOR2 (N13070, N13060, N8970);
xor XOR2 (N13071, N13063, N11712);
buf BUF1 (N13072, N13069);
or OR4 (N13073, N13065, N5992, N7648, N2015);
not NOT1 (N13074, N13057);
nor NOR4 (N13075, N13070, N12099, N852, N6284);
buf BUF1 (N13076, N13062);
or OR2 (N13077, N13071, N12807);
not NOT1 (N13078, N13075);
not NOT1 (N13079, N13078);
xor XOR2 (N13080, N13076, N4527);
xor XOR2 (N13081, N13077, N10561);
and AND2 (N13082, N13080, N6927);
nand NAND2 (N13083, N13066, N9055);
or OR2 (N13084, N13082, N2802);
xor XOR2 (N13085, N13083, N12933);
nor NOR4 (N13086, N13064, N12403, N3503, N7920);
nor NOR4 (N13087, N13074, N10951, N5823, N6339);
nand NAND2 (N13088, N13086, N10594);
not NOT1 (N13089, N13087);
xor XOR2 (N13090, N13079, N3261);
and AND2 (N13091, N13089, N5365);
and AND4 (N13092, N13091, N6644, N4510, N2336);
nor NOR4 (N13093, N13084, N11614, N5219, N10886);
and AND3 (N13094, N13093, N12946, N11708);
buf BUF1 (N13095, N13061);
not NOT1 (N13096, N13095);
buf BUF1 (N13097, N13092);
not NOT1 (N13098, N13090);
or OR3 (N13099, N13073, N12334, N11111);
nor NOR4 (N13100, N13096, N4316, N6652, N7375);
buf BUF1 (N13101, N13097);
and AND4 (N13102, N13101, N959, N6618, N12639);
not NOT1 (N13103, N13094);
and AND3 (N13104, N13103, N2045, N7584);
and AND4 (N13105, N13072, N1495, N10337, N11098);
xor XOR2 (N13106, N13104, N1892);
not NOT1 (N13107, N13098);
nand NAND4 (N13108, N13099, N1359, N5409, N7800);
xor XOR2 (N13109, N13106, N4287);
buf BUF1 (N13110, N13105);
xor XOR2 (N13111, N13109, N4635);
and AND3 (N13112, N13107, N7618, N4207);
or OR2 (N13113, N13100, N4839);
not NOT1 (N13114, N13111);
and AND4 (N13115, N13085, N7954, N8910, N12601);
nand NAND4 (N13116, N13088, N13095, N5612, N7836);
not NOT1 (N13117, N13114);
xor XOR2 (N13118, N13108, N8804);
xor XOR2 (N13119, N13115, N5275);
and AND2 (N13120, N13081, N12540);
or OR2 (N13121, N13053, N4560);
or OR2 (N13122, N13110, N2688);
or OR4 (N13123, N13118, N8193, N5284, N9540);
nor NOR4 (N13124, N13117, N10475, N5043, N10879);
xor XOR2 (N13125, N13120, N6772);
xor XOR2 (N13126, N13102, N2987);
and AND4 (N13127, N13119, N6748, N3083, N5150);
not NOT1 (N13128, N13121);
xor XOR2 (N13129, N13126, N3407);
buf BUF1 (N13130, N13116);
xor XOR2 (N13131, N13112, N4238);
and AND3 (N13132, N13125, N12816, N11993);
xor XOR2 (N13133, N13127, N6906);
or OR3 (N13134, N13131, N2265, N10526);
xor XOR2 (N13135, N13132, N5696);
or OR2 (N13136, N13122, N2364);
and AND2 (N13137, N13123, N9447);
not NOT1 (N13138, N13129);
not NOT1 (N13139, N13136);
buf BUF1 (N13140, N13138);
not NOT1 (N13141, N13124);
nor NOR2 (N13142, N13133, N9163);
nor NOR4 (N13143, N13135, N12292, N4975, N4716);
nand NAND3 (N13144, N13137, N2311, N5197);
buf BUF1 (N13145, N13128);
nor NOR4 (N13146, N13140, N10131, N7213, N7979);
nor NOR4 (N13147, N13144, N2713, N9643, N4882);
and AND3 (N13148, N13113, N9620, N12782);
and AND2 (N13149, N13146, N8271);
or OR3 (N13150, N13139, N11580, N7291);
and AND4 (N13151, N13141, N11560, N13098, N1999);
and AND3 (N13152, N13145, N8984, N11396);
buf BUF1 (N13153, N13149);
and AND4 (N13154, N13147, N6616, N3298, N1191);
and AND3 (N13155, N13152, N5276, N401);
or OR2 (N13156, N13143, N1689);
and AND2 (N13157, N13156, N8895);
buf BUF1 (N13158, N13157);
or OR2 (N13159, N13153, N12732);
and AND4 (N13160, N13159, N1657, N8940, N6285);
and AND2 (N13161, N13148, N5266);
nor NOR4 (N13162, N13151, N12836, N6061, N3231);
not NOT1 (N13163, N13160);
buf BUF1 (N13164, N13150);
buf BUF1 (N13165, N13134);
buf BUF1 (N13166, N13162);
or OR2 (N13167, N13166, N1543);
or OR4 (N13168, N13154, N2465, N10528, N9774);
xor XOR2 (N13169, N13161, N11373);
nand NAND3 (N13170, N13164, N470, N781);
not NOT1 (N13171, N13167);
nor NOR4 (N13172, N13165, N1860, N13121, N7915);
or OR4 (N13173, N13168, N10484, N2383, N12997);
nand NAND2 (N13174, N13169, N10848);
xor XOR2 (N13175, N13172, N619);
and AND2 (N13176, N13173, N4281);
or OR2 (N13177, N13142, N11323);
nor NOR3 (N13178, N13174, N12359, N8170);
xor XOR2 (N13179, N13130, N12861);
xor XOR2 (N13180, N13155, N8256);
nor NOR4 (N13181, N13163, N2286, N6110, N7190);
nor NOR2 (N13182, N13177, N516);
not NOT1 (N13183, N13179);
or OR3 (N13184, N13170, N10598, N5448);
nand NAND4 (N13185, N13182, N6006, N12176, N7299);
and AND3 (N13186, N13176, N11769, N2292);
and AND2 (N13187, N13186, N6393);
xor XOR2 (N13188, N13158, N8537);
not NOT1 (N13189, N13181);
xor XOR2 (N13190, N13171, N7324);
buf BUF1 (N13191, N13180);
buf BUF1 (N13192, N13191);
or OR3 (N13193, N13178, N3414, N4556);
nor NOR3 (N13194, N13185, N5395, N2232);
not NOT1 (N13195, N13192);
and AND3 (N13196, N13175, N5151, N1030);
nor NOR4 (N13197, N13183, N7405, N586, N4228);
not NOT1 (N13198, N13188);
and AND2 (N13199, N13190, N6608);
nor NOR3 (N13200, N13193, N12256, N11755);
nand NAND2 (N13201, N13184, N3033);
or OR4 (N13202, N13198, N13118, N12924, N7009);
not NOT1 (N13203, N13189);
xor XOR2 (N13204, N13199, N12767);
or OR2 (N13205, N13203, N8394);
nand NAND3 (N13206, N13204, N6241, N9478);
buf BUF1 (N13207, N13202);
nand NAND3 (N13208, N13187, N7310, N7336);
nor NOR4 (N13209, N13207, N6282, N10728, N11457);
and AND4 (N13210, N13196, N4732, N967, N3256);
nor NOR3 (N13211, N13200, N11560, N6910);
nor NOR3 (N13212, N13195, N6378, N298);
nor NOR4 (N13213, N13194, N8959, N1379, N67);
or OR2 (N13214, N13211, N3487);
not NOT1 (N13215, N13205);
buf BUF1 (N13216, N13197);
or OR2 (N13217, N13214, N9040);
and AND3 (N13218, N13201, N9055, N12119);
not NOT1 (N13219, N13213);
nor NOR3 (N13220, N13208, N5185, N10154);
xor XOR2 (N13221, N13210, N6995);
and AND3 (N13222, N13215, N7167, N10464);
nor NOR3 (N13223, N13209, N11353, N4431);
and AND2 (N13224, N13223, N3764);
nand NAND3 (N13225, N13218, N9138, N9046);
nor NOR2 (N13226, N13217, N11347);
nand NAND3 (N13227, N13226, N9851, N2121);
or OR2 (N13228, N13224, N4035);
buf BUF1 (N13229, N13221);
nand NAND2 (N13230, N13219, N10435);
nand NAND2 (N13231, N13216, N4079);
not NOT1 (N13232, N13225);
nor NOR3 (N13233, N13232, N7116, N1373);
and AND4 (N13234, N13222, N2545, N6307, N6376);
not NOT1 (N13235, N13230);
xor XOR2 (N13236, N13233, N8069);
xor XOR2 (N13237, N13234, N9254);
or OR4 (N13238, N13212, N5962, N9818, N6346);
buf BUF1 (N13239, N13228);
xor XOR2 (N13240, N13235, N2964);
buf BUF1 (N13241, N13238);
or OR2 (N13242, N13220, N19);
nor NOR2 (N13243, N13227, N13133);
not NOT1 (N13244, N13241);
buf BUF1 (N13245, N13242);
buf BUF1 (N13246, N13229);
xor XOR2 (N13247, N13231, N7252);
not NOT1 (N13248, N13239);
not NOT1 (N13249, N13245);
buf BUF1 (N13250, N13243);
nor NOR2 (N13251, N13249, N9703);
nor NOR3 (N13252, N13244, N8292, N12567);
buf BUF1 (N13253, N13251);
nand NAND2 (N13254, N13253, N7112);
buf BUF1 (N13255, N13248);
nor NOR3 (N13256, N13240, N11034, N278);
not NOT1 (N13257, N13237);
xor XOR2 (N13258, N13246, N8721);
buf BUF1 (N13259, N13247);
buf BUF1 (N13260, N13258);
or OR2 (N13261, N13206, N7303);
not NOT1 (N13262, N13250);
not NOT1 (N13263, N13236);
xor XOR2 (N13264, N13254, N6955);
or OR2 (N13265, N13262, N12337);
and AND2 (N13266, N13255, N12816);
or OR4 (N13267, N13261, N12845, N610, N8938);
or OR4 (N13268, N13257, N3198, N5146, N11665);
and AND3 (N13269, N13265, N12819, N7504);
nor NOR3 (N13270, N13267, N10965, N6544);
nand NAND3 (N13271, N13266, N6096, N10722);
buf BUF1 (N13272, N13260);
and AND4 (N13273, N13263, N3855, N7195, N7820);
xor XOR2 (N13274, N13259, N7848);
nor NOR3 (N13275, N13271, N3504, N8451);
nor NOR2 (N13276, N13272, N4199);
xor XOR2 (N13277, N13275, N10897);
xor XOR2 (N13278, N13269, N10010);
buf BUF1 (N13279, N13277);
and AND3 (N13280, N13274, N3836, N6854);
or OR4 (N13281, N13273, N6490, N2654, N1232);
nand NAND3 (N13282, N13270, N8716, N3411);
nor NOR2 (N13283, N13252, N7880);
nand NAND2 (N13284, N13278, N7406);
nand NAND4 (N13285, N13283, N10606, N9570, N9765);
and AND2 (N13286, N13285, N12296);
not NOT1 (N13287, N13281);
not NOT1 (N13288, N13284);
xor XOR2 (N13289, N13268, N8944);
nor NOR2 (N13290, N13264, N3587);
not NOT1 (N13291, N13287);
nor NOR3 (N13292, N13280, N280, N1398);
nand NAND2 (N13293, N13286, N7112);
nor NOR4 (N13294, N13292, N4822, N11478, N1574);
xor XOR2 (N13295, N13276, N714);
not NOT1 (N13296, N13291);
and AND2 (N13297, N13290, N10502);
xor XOR2 (N13298, N13279, N4034);
or OR4 (N13299, N13295, N11352, N1694, N994);
xor XOR2 (N13300, N13299, N10319);
nand NAND3 (N13301, N13293, N10249, N9231);
nor NOR4 (N13302, N13301, N2539, N1144, N5903);
buf BUF1 (N13303, N13294);
xor XOR2 (N13304, N13300, N6987);
xor XOR2 (N13305, N13256, N8668);
nand NAND3 (N13306, N13289, N6022, N11658);
and AND3 (N13307, N13298, N6467, N12065);
and AND3 (N13308, N13304, N12953, N6387);
nand NAND2 (N13309, N13296, N5536);
not NOT1 (N13310, N13302);
or OR4 (N13311, N13288, N7806, N6883, N5810);
not NOT1 (N13312, N13303);
nor NOR4 (N13313, N13305, N11784, N3154, N1551);
not NOT1 (N13314, N13308);
xor XOR2 (N13315, N13314, N13202);
not NOT1 (N13316, N13309);
not NOT1 (N13317, N13311);
nand NAND3 (N13318, N13282, N4005, N9759);
and AND4 (N13319, N13297, N11299, N3879, N525);
xor XOR2 (N13320, N13313, N11558);
nand NAND3 (N13321, N13307, N681, N4944);
buf BUF1 (N13322, N13319);
nand NAND4 (N13323, N13312, N10575, N670, N580);
and AND3 (N13324, N13315, N3610, N1223);
nand NAND3 (N13325, N13321, N8810, N9855);
nor NOR2 (N13326, N13322, N3651);
nand NAND3 (N13327, N13316, N12309, N12047);
nor NOR3 (N13328, N13317, N10316, N8867);
buf BUF1 (N13329, N13327);
not NOT1 (N13330, N13323);
xor XOR2 (N13331, N13320, N11932);
buf BUF1 (N13332, N13318);
nand NAND4 (N13333, N13332, N3984, N6496, N7566);
not NOT1 (N13334, N13330);
buf BUF1 (N13335, N13324);
buf BUF1 (N13336, N13326);
and AND2 (N13337, N13333, N9748);
nor NOR4 (N13338, N13328, N5370, N728, N11199);
not NOT1 (N13339, N13336);
nor NOR2 (N13340, N13310, N9682);
or OR4 (N13341, N13329, N2848, N3578, N1842);
nor NOR2 (N13342, N13339, N3084);
or OR2 (N13343, N13337, N7381);
and AND2 (N13344, N13342, N6041);
nand NAND4 (N13345, N13343, N7589, N11959, N8665);
not NOT1 (N13346, N13306);
xor XOR2 (N13347, N13331, N3061);
or OR3 (N13348, N13341, N11918, N5852);
nor NOR2 (N13349, N13338, N2272);
or OR4 (N13350, N13346, N3859, N1374, N6464);
buf BUF1 (N13351, N13345);
buf BUF1 (N13352, N13325);
buf BUF1 (N13353, N13335);
or OR4 (N13354, N13349, N5607, N5771, N4323);
buf BUF1 (N13355, N13351);
or OR2 (N13356, N13344, N5638);
buf BUF1 (N13357, N13334);
and AND3 (N13358, N13350, N1804, N11569);
nor NOR3 (N13359, N13352, N8176, N716);
nor NOR4 (N13360, N13356, N11501, N12403, N772);
and AND3 (N13361, N13348, N9525, N12036);
and AND4 (N13362, N13358, N1926, N8348, N9938);
or OR4 (N13363, N13360, N3949, N4246, N3001);
nand NAND3 (N13364, N13354, N6557, N3620);
buf BUF1 (N13365, N13361);
not NOT1 (N13366, N13362);
and AND3 (N13367, N13366, N9417, N5680);
and AND2 (N13368, N13363, N8242);
and AND3 (N13369, N13365, N12701, N5738);
nor NOR3 (N13370, N13367, N9917, N12772);
or OR3 (N13371, N13359, N8817, N7350);
and AND2 (N13372, N13357, N4331);
nor NOR2 (N13373, N13369, N982);
or OR3 (N13374, N13353, N7901, N9022);
not NOT1 (N13375, N13374);
not NOT1 (N13376, N13364);
not NOT1 (N13377, N13340);
not NOT1 (N13378, N13371);
buf BUF1 (N13379, N13378);
buf BUF1 (N13380, N13370);
nand NAND2 (N13381, N13377, N12865);
nor NOR2 (N13382, N13376, N3343);
or OR4 (N13383, N13380, N320, N5589, N961);
nand NAND3 (N13384, N13381, N7940, N11984);
nor NOR3 (N13385, N13383, N12858, N12885);
nand NAND3 (N13386, N13347, N1473, N7673);
not NOT1 (N13387, N13385);
buf BUF1 (N13388, N13372);
and AND4 (N13389, N13387, N10739, N1730, N132);
xor XOR2 (N13390, N13386, N1219);
and AND4 (N13391, N13389, N8868, N6031, N3706);
and AND3 (N13392, N13375, N12408, N8207);
xor XOR2 (N13393, N13355, N2568);
buf BUF1 (N13394, N13382);
nor NOR3 (N13395, N13373, N4148, N10668);
and AND4 (N13396, N13394, N7437, N11755, N8699);
buf BUF1 (N13397, N13388);
xor XOR2 (N13398, N13396, N9579);
not NOT1 (N13399, N13379);
not NOT1 (N13400, N13368);
or OR3 (N13401, N13384, N8103, N12470);
not NOT1 (N13402, N13393);
or OR4 (N13403, N13401, N10216, N3495, N6746);
nand NAND3 (N13404, N13390, N8118, N9919);
buf BUF1 (N13405, N13392);
and AND4 (N13406, N13400, N6826, N5355, N11298);
and AND4 (N13407, N13403, N9139, N12198, N11526);
or OR3 (N13408, N13406, N682, N9527);
nor NOR3 (N13409, N13398, N4885, N4501);
xor XOR2 (N13410, N13409, N11607);
not NOT1 (N13411, N13395);
or OR3 (N13412, N13408, N4392, N7676);
or OR4 (N13413, N13407, N11992, N4255, N12709);
buf BUF1 (N13414, N13402);
and AND4 (N13415, N13410, N2550, N10564, N3594);
nor NOR3 (N13416, N13397, N6730, N4040);
not NOT1 (N13417, N13405);
not NOT1 (N13418, N13404);
buf BUF1 (N13419, N13411);
and AND4 (N13420, N13414, N1760, N582, N6632);
nand NAND2 (N13421, N13420, N12312);
xor XOR2 (N13422, N13399, N9853);
and AND4 (N13423, N13419, N3633, N9262, N8366);
not NOT1 (N13424, N13422);
not NOT1 (N13425, N13424);
and AND4 (N13426, N13425, N5292, N11368, N11434);
and AND2 (N13427, N13421, N11425);
and AND3 (N13428, N13416, N1739, N12903);
nand NAND2 (N13429, N13418, N1339);
or OR3 (N13430, N13428, N8828, N684);
not NOT1 (N13431, N13423);
nor NOR4 (N13432, N13430, N5703, N7776, N9916);
not NOT1 (N13433, N13426);
not NOT1 (N13434, N13417);
nor NOR3 (N13435, N13427, N3473, N6363);
buf BUF1 (N13436, N13434);
nand NAND4 (N13437, N13413, N10219, N6790, N2011);
nand NAND4 (N13438, N13437, N4797, N8069, N3423);
nor NOR3 (N13439, N13436, N7081, N5336);
nor NOR3 (N13440, N13391, N11196, N1319);
or OR4 (N13441, N13412, N6675, N4147, N4145);
nand NAND4 (N13442, N13441, N11656, N6395, N1124);
buf BUF1 (N13443, N13442);
buf BUF1 (N13444, N13440);
nor NOR4 (N13445, N13439, N1138, N2980, N5240);
nand NAND4 (N13446, N13415, N1551, N3230, N8374);
xor XOR2 (N13447, N13429, N6311);
nand NAND2 (N13448, N13445, N3646);
nand NAND2 (N13449, N13431, N3599);
and AND3 (N13450, N13443, N11165, N13412);
not NOT1 (N13451, N13446);
xor XOR2 (N13452, N13432, N2852);
and AND4 (N13453, N13451, N10890, N3375, N12854);
nor NOR2 (N13454, N13447, N8306);
or OR3 (N13455, N13449, N4756, N7338);
xor XOR2 (N13456, N13433, N4411);
xor XOR2 (N13457, N13450, N2189);
nand NAND4 (N13458, N13438, N11607, N10591, N262);
not NOT1 (N13459, N13453);
xor XOR2 (N13460, N13454, N7345);
not NOT1 (N13461, N13456);
or OR2 (N13462, N13457, N5262);
not NOT1 (N13463, N13435);
or OR3 (N13464, N13461, N3523, N3730);
not NOT1 (N13465, N13460);
nand NAND2 (N13466, N13458, N4612);
buf BUF1 (N13467, N13462);
xor XOR2 (N13468, N13467, N5376);
nor NOR2 (N13469, N13463, N6340);
nor NOR2 (N13470, N13466, N11353);
and AND2 (N13471, N13464, N6312);
not NOT1 (N13472, N13455);
and AND4 (N13473, N13472, N8041, N6082, N10926);
nand NAND2 (N13474, N13470, N10840);
and AND2 (N13475, N13473, N10588);
and AND3 (N13476, N13469, N12152, N1178);
xor XOR2 (N13477, N13452, N12326);
xor XOR2 (N13478, N13459, N9085);
nor NOR4 (N13479, N13477, N1441, N9290, N5869);
nor NOR3 (N13480, N13444, N560, N13283);
xor XOR2 (N13481, N13471, N3763);
buf BUF1 (N13482, N13465);
nor NOR3 (N13483, N13478, N3095, N10867);
nor NOR3 (N13484, N13482, N4996, N2126);
buf BUF1 (N13485, N13480);
not NOT1 (N13486, N13479);
xor XOR2 (N13487, N13486, N11519);
xor XOR2 (N13488, N13475, N8439);
buf BUF1 (N13489, N13485);
nor NOR4 (N13490, N13474, N8341, N10743, N9796);
not NOT1 (N13491, N13489);
not NOT1 (N13492, N13484);
nor NOR4 (N13493, N13490, N10213, N8330, N4590);
buf BUF1 (N13494, N13488);
nor NOR4 (N13495, N13491, N1290, N10676, N9537);
buf BUF1 (N13496, N13492);
nor NOR4 (N13497, N13493, N12596, N8801, N8201);
buf BUF1 (N13498, N13481);
or OR4 (N13499, N13448, N8004, N11624, N4603);
xor XOR2 (N13500, N13476, N7423);
nand NAND4 (N13501, N13468, N5173, N12582, N5185);
nor NOR2 (N13502, N13499, N4985);
and AND4 (N13503, N13498, N1505, N997, N8658);
xor XOR2 (N13504, N13497, N584);
and AND3 (N13505, N13501, N3951, N10355);
not NOT1 (N13506, N13495);
nor NOR2 (N13507, N13496, N11787);
nand NAND3 (N13508, N13500, N1856, N7676);
xor XOR2 (N13509, N13508, N3573);
not NOT1 (N13510, N13487);
buf BUF1 (N13511, N13494);
and AND2 (N13512, N13509, N6096);
nand NAND3 (N13513, N13505, N3129, N5005);
nand NAND2 (N13514, N13513, N3402);
not NOT1 (N13515, N13483);
nor NOR4 (N13516, N13510, N12575, N3049, N12243);
or OR3 (N13517, N13502, N2228, N9465);
or OR2 (N13518, N13511, N13041);
or OR2 (N13519, N13512, N8426);
not NOT1 (N13520, N13518);
not NOT1 (N13521, N13514);
nor NOR2 (N13522, N13504, N9822);
nor NOR2 (N13523, N13507, N11829);
and AND4 (N13524, N13520, N11074, N11961, N10185);
nand NAND2 (N13525, N13506, N12181);
xor XOR2 (N13526, N13517, N7535);
not NOT1 (N13527, N13521);
xor XOR2 (N13528, N13527, N5232);
nor NOR3 (N13529, N13522, N5323, N10477);
xor XOR2 (N13530, N13528, N2322);
not NOT1 (N13531, N13529);
not NOT1 (N13532, N13519);
xor XOR2 (N13533, N13516, N9116);
nor NOR2 (N13534, N13523, N9815);
or OR3 (N13535, N13530, N11303, N6466);
not NOT1 (N13536, N13525);
xor XOR2 (N13537, N13526, N6418);
and AND2 (N13538, N13503, N2094);
nand NAND4 (N13539, N13531, N12405, N4631, N13037);
or OR2 (N13540, N13538, N11923);
nand NAND3 (N13541, N13534, N1001, N4158);
buf BUF1 (N13542, N13540);
and AND2 (N13543, N13542, N4419);
and AND2 (N13544, N13543, N940);
or OR4 (N13545, N13532, N847, N10792, N3873);
xor XOR2 (N13546, N13515, N10315);
not NOT1 (N13547, N13533);
buf BUF1 (N13548, N13545);
nand NAND4 (N13549, N13536, N2405, N5876, N8327);
buf BUF1 (N13550, N13539);
nand NAND2 (N13551, N13541, N4007);
not NOT1 (N13552, N13537);
buf BUF1 (N13553, N13547);
or OR2 (N13554, N13551, N10737);
or OR3 (N13555, N13544, N11781, N2225);
and AND4 (N13556, N13524, N3909, N9393, N6002);
not NOT1 (N13557, N13552);
and AND3 (N13558, N13546, N4950, N1503);
and AND3 (N13559, N13548, N1203, N4593);
or OR3 (N13560, N13554, N9490, N3482);
nand NAND2 (N13561, N13535, N583);
xor XOR2 (N13562, N13559, N6404);
or OR2 (N13563, N13557, N7367);
or OR4 (N13564, N13550, N1570, N1852, N4376);
buf BUF1 (N13565, N13560);
buf BUF1 (N13566, N13561);
xor XOR2 (N13567, N13558, N12202);
and AND2 (N13568, N13564, N12436);
or OR4 (N13569, N13562, N10442, N6510, N347);
and AND2 (N13570, N13565, N10175);
and AND4 (N13571, N13569, N11835, N10128, N1422);
not NOT1 (N13572, N13556);
nand NAND2 (N13573, N13571, N8007);
or OR2 (N13574, N13573, N4623);
nand NAND4 (N13575, N13566, N1445, N2368, N10747);
xor XOR2 (N13576, N13553, N5713);
xor XOR2 (N13577, N13567, N6560);
buf BUF1 (N13578, N13549);
nand NAND4 (N13579, N13578, N3846, N5551, N10971);
xor XOR2 (N13580, N13577, N4273);
nor NOR2 (N13581, N13575, N3961);
xor XOR2 (N13582, N13581, N4705);
and AND2 (N13583, N13572, N5029);
or OR4 (N13584, N13563, N3077, N4655, N12728);
and AND3 (N13585, N13580, N10255, N5438);
and AND3 (N13586, N13579, N11871, N12034);
and AND3 (N13587, N13585, N8083, N4287);
and AND3 (N13588, N13586, N11534, N10146);
xor XOR2 (N13589, N13568, N7843);
and AND3 (N13590, N13576, N1369, N1465);
xor XOR2 (N13591, N13587, N4127);
buf BUF1 (N13592, N13574);
buf BUF1 (N13593, N13588);
nand NAND2 (N13594, N13590, N8391);
buf BUF1 (N13595, N13555);
nand NAND4 (N13596, N13583, N13558, N8911, N7607);
not NOT1 (N13597, N13582);
nor NOR3 (N13598, N13597, N7874, N12711);
buf BUF1 (N13599, N13596);
nor NOR2 (N13600, N13584, N9749);
and AND2 (N13601, N13589, N4730);
or OR4 (N13602, N13601, N4505, N11682, N4899);
and AND3 (N13603, N13598, N5635, N9395);
nand NAND2 (N13604, N13592, N5164);
or OR4 (N13605, N13595, N3392, N295, N3287);
nand NAND4 (N13606, N13593, N7719, N10760, N12088);
nor NOR4 (N13607, N13602, N2233, N3015, N11129);
not NOT1 (N13608, N13600);
xor XOR2 (N13609, N13604, N4607);
or OR4 (N13610, N13606, N9342, N6824, N9778);
nand NAND2 (N13611, N13605, N13496);
nor NOR4 (N13612, N13594, N9670, N4496, N12617);
xor XOR2 (N13613, N13599, N4187);
or OR4 (N13614, N13611, N7089, N3514, N2392);
not NOT1 (N13615, N13613);
nor NOR2 (N13616, N13615, N6228);
not NOT1 (N13617, N13614);
buf BUF1 (N13618, N13616);
or OR2 (N13619, N13610, N9297);
and AND2 (N13620, N13591, N2547);
xor XOR2 (N13621, N13617, N13259);
xor XOR2 (N13622, N13607, N13179);
or OR2 (N13623, N13612, N9398);
buf BUF1 (N13624, N13621);
nor NOR3 (N13625, N13603, N4688, N8778);
xor XOR2 (N13626, N13623, N5772);
and AND2 (N13627, N13609, N8625);
buf BUF1 (N13628, N13627);
not NOT1 (N13629, N13570);
xor XOR2 (N13630, N13608, N7414);
or OR4 (N13631, N13620, N3704, N8473, N2878);
not NOT1 (N13632, N13629);
buf BUF1 (N13633, N13625);
and AND3 (N13634, N13628, N8734, N10956);
or OR3 (N13635, N13619, N1647, N325);
nand NAND3 (N13636, N13626, N949, N5708);
not NOT1 (N13637, N13618);
not NOT1 (N13638, N13634);
nand NAND2 (N13639, N13630, N3816);
nor NOR2 (N13640, N13632, N5778);
xor XOR2 (N13641, N13640, N13590);
or OR4 (N13642, N13624, N5155, N12991, N12614);
nor NOR4 (N13643, N13641, N2246, N1639, N6529);
and AND2 (N13644, N13631, N4105);
nor NOR2 (N13645, N13636, N11722);
not NOT1 (N13646, N13635);
buf BUF1 (N13647, N13637);
or OR3 (N13648, N13638, N3687, N2207);
buf BUF1 (N13649, N13622);
nand NAND3 (N13650, N13643, N3704, N5627);
and AND3 (N13651, N13650, N4520, N9784);
buf BUF1 (N13652, N13647);
not NOT1 (N13653, N13649);
and AND2 (N13654, N13648, N9003);
not NOT1 (N13655, N13653);
and AND4 (N13656, N13639, N2405, N1434, N11411);
nor NOR3 (N13657, N13645, N5877, N8421);
buf BUF1 (N13658, N13655);
not NOT1 (N13659, N13657);
nand NAND4 (N13660, N13658, N8110, N12060, N1954);
xor XOR2 (N13661, N13654, N7427);
nand NAND2 (N13662, N13646, N8807);
not NOT1 (N13663, N13662);
not NOT1 (N13664, N13656);
xor XOR2 (N13665, N13652, N13607);
xor XOR2 (N13666, N13659, N12991);
and AND4 (N13667, N13661, N10477, N11352, N1121);
nor NOR4 (N13668, N13664, N5452, N81, N13140);
or OR3 (N13669, N13642, N7039, N5181);
and AND2 (N13670, N13667, N11008);
or OR2 (N13671, N13644, N3830);
buf BUF1 (N13672, N13663);
or OR4 (N13673, N13660, N9192, N8688, N82);
not NOT1 (N13674, N13670);
or OR2 (N13675, N13666, N9337);
or OR2 (N13676, N13673, N8742);
and AND2 (N13677, N13671, N11598);
buf BUF1 (N13678, N13633);
nand NAND2 (N13679, N13651, N12919);
and AND3 (N13680, N13669, N10239, N286);
xor XOR2 (N13681, N13672, N299);
nor NOR2 (N13682, N13675, N1890);
nor NOR2 (N13683, N13682, N5135);
or OR2 (N13684, N13674, N1334);
nor NOR3 (N13685, N13676, N12992, N9929);
and AND3 (N13686, N13683, N3276, N8152);
or OR4 (N13687, N13680, N3474, N2603, N917);
buf BUF1 (N13688, N13685);
nor NOR2 (N13689, N13679, N13400);
and AND2 (N13690, N13668, N12714);
or OR4 (N13691, N13689, N9027, N4662, N7522);
buf BUF1 (N13692, N13690);
xor XOR2 (N13693, N13665, N1167);
nand NAND3 (N13694, N13692, N6558, N13116);
or OR3 (N13695, N13678, N12521, N3202);
not NOT1 (N13696, N13695);
or OR4 (N13697, N13677, N10371, N12484, N3521);
nand NAND4 (N13698, N13681, N2378, N3954, N2102);
nor NOR3 (N13699, N13694, N1888, N5594);
nor NOR4 (N13700, N13693, N8407, N264, N11786);
and AND2 (N13701, N13696, N5994);
or OR4 (N13702, N13684, N3618, N1494, N13250);
not NOT1 (N13703, N13697);
buf BUF1 (N13704, N13687);
nor NOR4 (N13705, N13699, N1450, N3090, N11280);
nand NAND4 (N13706, N13691, N466, N2151, N7851);
buf BUF1 (N13707, N13700);
or OR4 (N13708, N13701, N1446, N10845, N3477);
and AND4 (N13709, N13705, N5999, N3046, N1692);
and AND3 (N13710, N13702, N5842, N11172);
or OR3 (N13711, N13688, N13134, N1682);
or OR3 (N13712, N13709, N9, N2939);
nand NAND3 (N13713, N13706, N59, N8043);
and AND3 (N13714, N13698, N7343, N2849);
buf BUF1 (N13715, N13712);
nand NAND2 (N13716, N13708, N11654);
or OR4 (N13717, N13713, N5662, N3811, N8854);
or OR4 (N13718, N13716, N11922, N13116, N3365);
nand NAND3 (N13719, N13710, N12142, N12295);
nand NAND2 (N13720, N13719, N889);
not NOT1 (N13721, N13704);
not NOT1 (N13722, N13703);
nand NAND4 (N13723, N13720, N8409, N10996, N10953);
buf BUF1 (N13724, N13721);
or OR3 (N13725, N13717, N7908, N9918);
xor XOR2 (N13726, N13711, N5422);
buf BUF1 (N13727, N13722);
and AND3 (N13728, N13714, N8292, N11419);
xor XOR2 (N13729, N13725, N2109);
or OR3 (N13730, N13729, N1618, N4809);
or OR2 (N13731, N13707, N5158);
or OR3 (N13732, N13724, N4128, N12552);
not NOT1 (N13733, N13726);
nand NAND2 (N13734, N13727, N5130);
buf BUF1 (N13735, N13723);
not NOT1 (N13736, N13730);
and AND2 (N13737, N13732, N9578);
not NOT1 (N13738, N13737);
and AND3 (N13739, N13735, N11109, N13227);
nand NAND4 (N13740, N13733, N4527, N6456, N1090);
and AND2 (N13741, N13736, N7191);
xor XOR2 (N13742, N13739, N5384);
not NOT1 (N13743, N13715);
or OR4 (N13744, N13743, N5029, N10531, N9456);
not NOT1 (N13745, N13744);
nand NAND2 (N13746, N13686, N3059);
buf BUF1 (N13747, N13734);
buf BUF1 (N13748, N13742);
xor XOR2 (N13749, N13718, N11660);
buf BUF1 (N13750, N13728);
buf BUF1 (N13751, N13745);
and AND4 (N13752, N13749, N9267, N6744, N9657);
and AND2 (N13753, N13731, N10262);
nor NOR3 (N13754, N13750, N7169, N4006);
xor XOR2 (N13755, N13748, N12538);
nand NAND3 (N13756, N13752, N3507, N3295);
not NOT1 (N13757, N13747);
buf BUF1 (N13758, N13741);
not NOT1 (N13759, N13756);
nor NOR4 (N13760, N13738, N2152, N7597, N12040);
or OR4 (N13761, N13753, N5858, N131, N8592);
nor NOR2 (N13762, N13760, N1945);
xor XOR2 (N13763, N13757, N10416);
buf BUF1 (N13764, N13759);
buf BUF1 (N13765, N13740);
nand NAND3 (N13766, N13765, N3002, N3205);
not NOT1 (N13767, N13755);
nor NOR2 (N13768, N13758, N10274);
xor XOR2 (N13769, N13746, N8998);
nor NOR3 (N13770, N13763, N11914, N6229);
not NOT1 (N13771, N13766);
buf BUF1 (N13772, N13767);
not NOT1 (N13773, N13761);
and AND3 (N13774, N13769, N12772, N6126);
xor XOR2 (N13775, N13770, N9374);
buf BUF1 (N13776, N13751);
and AND4 (N13777, N13764, N2814, N5145, N726);
nand NAND2 (N13778, N13776, N6820);
and AND3 (N13779, N13773, N5314, N6999);
xor XOR2 (N13780, N13772, N8646);
buf BUF1 (N13781, N13768);
and AND4 (N13782, N13779, N8176, N11960, N5295);
or OR2 (N13783, N13771, N8273);
buf BUF1 (N13784, N13781);
or OR3 (N13785, N13762, N10335, N7040);
nand NAND4 (N13786, N13780, N13333, N3953, N11888);
nor NOR4 (N13787, N13778, N1432, N11068, N895);
xor XOR2 (N13788, N13783, N3504);
nor NOR4 (N13789, N13774, N11652, N950, N9441);
buf BUF1 (N13790, N13777);
nand NAND2 (N13791, N13788, N13301);
nand NAND4 (N13792, N13789, N12957, N1964, N7318);
xor XOR2 (N13793, N13784, N422);
nor NOR2 (N13794, N13787, N5333);
buf BUF1 (N13795, N13792);
or OR4 (N13796, N13794, N5801, N665, N12673);
not NOT1 (N13797, N13791);
and AND4 (N13798, N13785, N5800, N10853, N6858);
xor XOR2 (N13799, N13786, N6809);
nand NAND4 (N13800, N13796, N4121, N8738, N5350);
buf BUF1 (N13801, N13793);
nand NAND3 (N13802, N13754, N12300, N6583);
not NOT1 (N13803, N13790);
and AND3 (N13804, N13795, N12413, N3461);
xor XOR2 (N13805, N13803, N2386);
not NOT1 (N13806, N13797);
xor XOR2 (N13807, N13800, N8010);
nand NAND3 (N13808, N13798, N8028, N12459);
nand NAND2 (N13809, N13801, N4193);
xor XOR2 (N13810, N13809, N10886);
xor XOR2 (N13811, N13802, N3402);
buf BUF1 (N13812, N13810);
nor NOR3 (N13813, N13806, N8841, N13299);
buf BUF1 (N13814, N13811);
nand NAND3 (N13815, N13807, N5699, N11023);
buf BUF1 (N13816, N13775);
xor XOR2 (N13817, N13812, N5758);
and AND2 (N13818, N13805, N1806);
nand NAND4 (N13819, N13813, N2079, N9202, N13343);
not NOT1 (N13820, N13819);
or OR4 (N13821, N13804, N3426, N1460, N1334);
or OR2 (N13822, N13808, N10910);
or OR3 (N13823, N13814, N10862, N9838);
nor NOR3 (N13824, N13823, N11591, N11984);
nor NOR2 (N13825, N13821, N8523);
nand NAND4 (N13826, N13820, N7693, N8186, N10571);
not NOT1 (N13827, N13818);
not NOT1 (N13828, N13822);
or OR4 (N13829, N13828, N965, N13218, N13389);
or OR4 (N13830, N13826, N2295, N3426, N5144);
buf BUF1 (N13831, N13829);
and AND4 (N13832, N13825, N10124, N674, N9307);
buf BUF1 (N13833, N13815);
and AND4 (N13834, N13816, N5893, N3398, N5520);
nor NOR4 (N13835, N13817, N5535, N3354, N6210);
and AND3 (N13836, N13799, N12091, N3741);
nand NAND4 (N13837, N13833, N2791, N8957, N8058);
not NOT1 (N13838, N13824);
buf BUF1 (N13839, N13837);
buf BUF1 (N13840, N13827);
xor XOR2 (N13841, N13840, N5343);
nand NAND3 (N13842, N13835, N3631, N5071);
and AND2 (N13843, N13841, N2011);
and AND4 (N13844, N13782, N10578, N9657, N7775);
or OR2 (N13845, N13839, N7536);
not NOT1 (N13846, N13838);
xor XOR2 (N13847, N13836, N13414);
nor NOR4 (N13848, N13832, N12988, N7489, N187);
or OR2 (N13849, N13831, N4387);
buf BUF1 (N13850, N13849);
or OR4 (N13851, N13843, N7096, N12291, N7687);
nor NOR3 (N13852, N13850, N11086, N99);
not NOT1 (N13853, N13846);
nor NOR2 (N13854, N13848, N3990);
xor XOR2 (N13855, N13854, N2435);
and AND4 (N13856, N13853, N7889, N3430, N9055);
buf BUF1 (N13857, N13855);
not NOT1 (N13858, N13842);
and AND2 (N13859, N13851, N10971);
buf BUF1 (N13860, N13857);
or OR2 (N13861, N13847, N1467);
and AND3 (N13862, N13852, N10445, N8969);
buf BUF1 (N13863, N13860);
nand NAND3 (N13864, N13862, N999, N9687);
buf BUF1 (N13865, N13858);
and AND3 (N13866, N13856, N7438, N8001);
nor NOR3 (N13867, N13865, N12133, N1778);
buf BUF1 (N13868, N13866);
buf BUF1 (N13869, N13861);
or OR4 (N13870, N13864, N4539, N13200, N6634);
not NOT1 (N13871, N13870);
and AND3 (N13872, N13830, N2496, N13821);
nor NOR4 (N13873, N13872, N2764, N4784, N7546);
xor XOR2 (N13874, N13845, N11752);
nand NAND4 (N13875, N13859, N10433, N6587, N9123);
buf BUF1 (N13876, N13868);
buf BUF1 (N13877, N13873);
nor NOR3 (N13878, N13874, N8959, N8781);
not NOT1 (N13879, N13877);
not NOT1 (N13880, N13876);
or OR2 (N13881, N13867, N7533);
xor XOR2 (N13882, N13875, N225);
or OR3 (N13883, N13834, N11264, N728);
nand NAND3 (N13884, N13863, N1527, N6363);
or OR4 (N13885, N13844, N1904, N6648, N7151);
not NOT1 (N13886, N13878);
and AND3 (N13887, N13879, N1192, N4673);
and AND3 (N13888, N13880, N7385, N6733);
nor NOR2 (N13889, N13881, N7290);
or OR4 (N13890, N13883, N10854, N8273, N5577);
and AND4 (N13891, N13869, N13120, N5685, N417);
buf BUF1 (N13892, N13888);
not NOT1 (N13893, N13890);
buf BUF1 (N13894, N13884);
nor NOR4 (N13895, N13894, N10744, N6098, N5232);
and AND2 (N13896, N13887, N11545);
and AND4 (N13897, N13882, N13399, N1454, N9274);
buf BUF1 (N13898, N13896);
nand NAND2 (N13899, N13889, N9743);
or OR2 (N13900, N13885, N3571);
xor XOR2 (N13901, N13899, N8871);
nand NAND4 (N13902, N13900, N12012, N9822, N12934);
buf BUF1 (N13903, N13902);
xor XOR2 (N13904, N13898, N10998);
and AND2 (N13905, N13891, N12703);
nor NOR3 (N13906, N13903, N234, N5507);
xor XOR2 (N13907, N13893, N2882);
not NOT1 (N13908, N13904);
buf BUF1 (N13909, N13886);
buf BUF1 (N13910, N13907);
and AND2 (N13911, N13908, N2780);
nor NOR3 (N13912, N13910, N10557, N8188);
nor NOR3 (N13913, N13897, N12982, N2978);
not NOT1 (N13914, N13906);
and AND4 (N13915, N13901, N13359, N9012, N12707);
and AND3 (N13916, N13915, N2410, N11064);
or OR3 (N13917, N13916, N1696, N1684);
buf BUF1 (N13918, N13914);
buf BUF1 (N13919, N13917);
and AND4 (N13920, N13918, N1122, N11061, N13768);
and AND2 (N13921, N13920, N10660);
not NOT1 (N13922, N13905);
nand NAND2 (N13923, N13921, N6566);
nor NOR2 (N13924, N13871, N11504);
or OR3 (N13925, N13895, N9946, N5720);
nand NAND3 (N13926, N13919, N9231, N1365);
or OR3 (N13927, N13913, N1026, N8209);
nor NOR2 (N13928, N13909, N1852);
buf BUF1 (N13929, N13925);
or OR3 (N13930, N13912, N2629, N6896);
nand NAND2 (N13931, N13922, N8045);
nor NOR4 (N13932, N13929, N2883, N9857, N12094);
not NOT1 (N13933, N13924);
or OR4 (N13934, N13911, N6436, N5659, N8061);
xor XOR2 (N13935, N13923, N3380);
xor XOR2 (N13936, N13935, N5790);
nor NOR4 (N13937, N13892, N11804, N3858, N7043);
and AND4 (N13938, N13937, N217, N2201, N5771);
xor XOR2 (N13939, N13936, N13362);
xor XOR2 (N13940, N13933, N3493);
or OR2 (N13941, N13932, N2783);
nor NOR4 (N13942, N13928, N5252, N9392, N153);
not NOT1 (N13943, N13940);
buf BUF1 (N13944, N13943);
xor XOR2 (N13945, N13942, N6465);
xor XOR2 (N13946, N13927, N8631);
not NOT1 (N13947, N13941);
nand NAND4 (N13948, N13944, N12534, N12999, N12816);
not NOT1 (N13949, N13947);
and AND4 (N13950, N13938, N2592, N6174, N5782);
not NOT1 (N13951, N13945);
buf BUF1 (N13952, N13939);
xor XOR2 (N13953, N13926, N7657);
or OR4 (N13954, N13949, N5576, N6446, N6593);
or OR2 (N13955, N13931, N48);
xor XOR2 (N13956, N13952, N10438);
xor XOR2 (N13957, N13934, N6013);
or OR3 (N13958, N13954, N10095, N6188);
xor XOR2 (N13959, N13946, N419);
buf BUF1 (N13960, N13955);
buf BUF1 (N13961, N13948);
buf BUF1 (N13962, N13951);
buf BUF1 (N13963, N13961);
nand NAND2 (N13964, N13953, N2584);
or OR2 (N13965, N13958, N11863);
buf BUF1 (N13966, N13959);
buf BUF1 (N13967, N13965);
xor XOR2 (N13968, N13930, N13241);
nand NAND4 (N13969, N13956, N12791, N6448, N13390);
nor NOR3 (N13970, N13960, N8182, N10392);
and AND4 (N13971, N13962, N13709, N1699, N12075);
and AND4 (N13972, N13967, N11138, N7860, N12609);
nor NOR4 (N13973, N13950, N10417, N4671, N560);
or OR4 (N13974, N13970, N6455, N13300, N13321);
buf BUF1 (N13975, N13969);
buf BUF1 (N13976, N13966);
not NOT1 (N13977, N13957);
xor XOR2 (N13978, N13971, N12610);
not NOT1 (N13979, N13975);
xor XOR2 (N13980, N13973, N6701);
xor XOR2 (N13981, N13977, N8943);
xor XOR2 (N13982, N13981, N7756);
or OR3 (N13983, N13979, N13870, N1826);
or OR2 (N13984, N13976, N5303);
xor XOR2 (N13985, N13982, N12555);
xor XOR2 (N13986, N13974, N5163);
not NOT1 (N13987, N13983);
and AND2 (N13988, N13968, N541);
xor XOR2 (N13989, N13964, N151);
nor NOR4 (N13990, N13984, N3462, N12693, N5561);
nand NAND2 (N13991, N13972, N3696);
not NOT1 (N13992, N13986);
or OR2 (N13993, N13992, N9618);
xor XOR2 (N13994, N13985, N8802);
nand NAND4 (N13995, N13989, N10321, N4859, N6052);
nand NAND4 (N13996, N13987, N6486, N11581, N10713);
nor NOR4 (N13997, N13990, N1452, N6509, N3419);
xor XOR2 (N13998, N13995, N4468);
xor XOR2 (N13999, N13994, N1797);
nand NAND4 (N14000, N13963, N10511, N566, N7126);
and AND2 (N14001, N13988, N13319);
xor XOR2 (N14002, N13978, N13456);
nand NAND2 (N14003, N13996, N1426);
and AND3 (N14004, N13993, N11626, N9416);
buf BUF1 (N14005, N13997);
xor XOR2 (N14006, N13998, N6230);
buf BUF1 (N14007, N13980);
nand NAND4 (N14008, N14003, N9387, N3472, N12097);
and AND4 (N14009, N14008, N11404, N5448, N4943);
buf BUF1 (N14010, N14005);
nor NOR4 (N14011, N14009, N9767, N11809, N7282);
nor NOR3 (N14012, N14000, N13805, N6466);
not NOT1 (N14013, N14010);
and AND2 (N14014, N14002, N2597);
nor NOR2 (N14015, N14012, N3282);
nor NOR4 (N14016, N14011, N395, N5572, N4076);
nand NAND2 (N14017, N14007, N4006);
and AND2 (N14018, N14006, N3605);
nand NAND4 (N14019, N14014, N175, N6034, N4838);
nor NOR4 (N14020, N14004, N13546, N6691, N1332);
not NOT1 (N14021, N14017);
not NOT1 (N14022, N14015);
or OR3 (N14023, N14021, N11591, N6601);
and AND3 (N14024, N13999, N10285, N4526);
buf BUF1 (N14025, N14024);
not NOT1 (N14026, N14019);
and AND2 (N14027, N14013, N7490);
and AND2 (N14028, N14022, N1962);
buf BUF1 (N14029, N14025);
or OR2 (N14030, N14027, N4463);
buf BUF1 (N14031, N14030);
and AND2 (N14032, N14023, N6428);
not NOT1 (N14033, N14032);
xor XOR2 (N14034, N14018, N9361);
and AND3 (N14035, N14028, N12454, N1165);
buf BUF1 (N14036, N14034);
xor XOR2 (N14037, N14020, N1253);
and AND4 (N14038, N14001, N11802, N1864, N7580);
buf BUF1 (N14039, N14038);
nand NAND4 (N14040, N14031, N9127, N5725, N4751);
or OR2 (N14041, N13991, N11660);
xor XOR2 (N14042, N14033, N10836);
nor NOR2 (N14043, N14035, N14013);
xor XOR2 (N14044, N14016, N8258);
or OR2 (N14045, N14041, N10869);
nor NOR2 (N14046, N14036, N289);
buf BUF1 (N14047, N14043);
not NOT1 (N14048, N14029);
buf BUF1 (N14049, N14042);
nand NAND4 (N14050, N14037, N2400, N13484, N9006);
and AND2 (N14051, N14048, N11989);
or OR2 (N14052, N14050, N2965);
xor XOR2 (N14053, N14051, N11027);
or OR3 (N14054, N14045, N3294, N3198);
not NOT1 (N14055, N14052);
and AND4 (N14056, N14049, N2516, N3413, N8316);
buf BUF1 (N14057, N14039);
nand NAND3 (N14058, N14057, N11926, N5526);
and AND3 (N14059, N14055, N12985, N9230);
not NOT1 (N14060, N14058);
not NOT1 (N14061, N14026);
buf BUF1 (N14062, N14056);
buf BUF1 (N14063, N14054);
buf BUF1 (N14064, N14059);
nor NOR3 (N14065, N14044, N10163, N6480);
and AND3 (N14066, N14047, N5437, N4707);
nor NOR2 (N14067, N14046, N2832);
nand NAND3 (N14068, N14062, N3484, N8428);
and AND4 (N14069, N14060, N8899, N4528, N13907);
nor NOR3 (N14070, N14064, N13195, N8250);
and AND2 (N14071, N14063, N9091);
or OR3 (N14072, N14068, N6930, N12920);
or OR3 (N14073, N14072, N4802, N7764);
or OR2 (N14074, N14053, N5148);
or OR4 (N14075, N14061, N10193, N8580, N5870);
xor XOR2 (N14076, N14071, N4510);
buf BUF1 (N14077, N14073);
or OR3 (N14078, N14040, N11505, N10965);
buf BUF1 (N14079, N14065);
and AND2 (N14080, N14079, N10070);
buf BUF1 (N14081, N14074);
buf BUF1 (N14082, N14077);
not NOT1 (N14083, N14080);
or OR3 (N14084, N14083, N2241, N2074);
xor XOR2 (N14085, N14081, N12411);
nand NAND3 (N14086, N14078, N5906, N9593);
xor XOR2 (N14087, N14067, N3216);
xor XOR2 (N14088, N14082, N12038);
xor XOR2 (N14089, N14086, N11573);
xor XOR2 (N14090, N14088, N3575);
buf BUF1 (N14091, N14070);
nand NAND4 (N14092, N14075, N5273, N9150, N7335);
not NOT1 (N14093, N14085);
and AND3 (N14094, N14091, N12270, N4);
xor XOR2 (N14095, N14092, N9867);
buf BUF1 (N14096, N14084);
nand NAND3 (N14097, N14095, N10963, N8913);
or OR2 (N14098, N14090, N4252);
buf BUF1 (N14099, N14097);
not NOT1 (N14100, N14094);
not NOT1 (N14101, N14100);
and AND4 (N14102, N14093, N459, N12107, N4824);
and AND3 (N14103, N14066, N11374, N2617);
nand NAND4 (N14104, N14098, N9540, N12808, N5314);
not NOT1 (N14105, N14104);
nor NOR2 (N14106, N14096, N11171);
nand NAND4 (N14107, N14087, N12373, N7208, N2505);
or OR3 (N14108, N14099, N731, N3993);
and AND2 (N14109, N14103, N5803);
xor XOR2 (N14110, N14109, N1295);
nand NAND3 (N14111, N14101, N5368, N12035);
buf BUF1 (N14112, N14069);
nand NAND2 (N14113, N14112, N8767);
not NOT1 (N14114, N14113);
buf BUF1 (N14115, N14107);
not NOT1 (N14116, N14114);
not NOT1 (N14117, N14111);
or OR2 (N14118, N14089, N13493);
buf BUF1 (N14119, N14105);
and AND4 (N14120, N14116, N13461, N344, N2896);
xor XOR2 (N14121, N14120, N609);
buf BUF1 (N14122, N14117);
or OR3 (N14123, N14121, N6144, N2346);
or OR3 (N14124, N14115, N10014, N2914);
not NOT1 (N14125, N14118);
buf BUF1 (N14126, N14123);
and AND4 (N14127, N14124, N6156, N5876, N10679);
xor XOR2 (N14128, N14127, N13137);
or OR4 (N14129, N14128, N8193, N11837, N5892);
and AND4 (N14130, N14129, N8986, N13395, N6523);
buf BUF1 (N14131, N14125);
xor XOR2 (N14132, N14126, N3953);
not NOT1 (N14133, N14132);
or OR3 (N14134, N14106, N11404, N8273);
buf BUF1 (N14135, N14130);
xor XOR2 (N14136, N14135, N7542);
or OR3 (N14137, N14108, N2553, N9891);
xor XOR2 (N14138, N14133, N448);
buf BUF1 (N14139, N14102);
not NOT1 (N14140, N14137);
and AND2 (N14141, N14122, N11270);
or OR2 (N14142, N14110, N12858);
or OR3 (N14143, N14142, N13448, N11894);
buf BUF1 (N14144, N14139);
buf BUF1 (N14145, N14140);
nor NOR2 (N14146, N14141, N5737);
and AND2 (N14147, N14131, N5442);
and AND3 (N14148, N14147, N5644, N9503);
buf BUF1 (N14149, N14148);
not NOT1 (N14150, N14076);
not NOT1 (N14151, N14136);
nand NAND2 (N14152, N14149, N8122);
not NOT1 (N14153, N14151);
xor XOR2 (N14154, N14145, N6806);
nor NOR4 (N14155, N14153, N1294, N9557, N8683);
buf BUF1 (N14156, N14146);
not NOT1 (N14157, N14152);
buf BUF1 (N14158, N14138);
not NOT1 (N14159, N14119);
or OR3 (N14160, N14159, N13596, N11372);
buf BUF1 (N14161, N14157);
buf BUF1 (N14162, N14150);
nor NOR4 (N14163, N14156, N7829, N10451, N13311);
xor XOR2 (N14164, N14155, N2956);
not NOT1 (N14165, N14154);
not NOT1 (N14166, N14134);
not NOT1 (N14167, N14161);
nor NOR2 (N14168, N14158, N8155);
not NOT1 (N14169, N14166);
and AND3 (N14170, N14143, N13300, N4181);
not NOT1 (N14171, N14165);
xor XOR2 (N14172, N14168, N10642);
not NOT1 (N14173, N14163);
nor NOR3 (N14174, N14172, N4400, N8604);
xor XOR2 (N14175, N14170, N5104);
and AND4 (N14176, N14174, N9503, N9380, N7188);
and AND4 (N14177, N14169, N3955, N9333, N7297);
nand NAND3 (N14178, N14160, N2282, N8842);
or OR2 (N14179, N14167, N7924);
not NOT1 (N14180, N14178);
or OR4 (N14181, N14175, N793, N7979, N3084);
and AND3 (N14182, N14176, N13797, N770);
nor NOR2 (N14183, N14180, N511);
nor NOR3 (N14184, N14179, N9771, N5903);
nand NAND2 (N14185, N14182, N2488);
not NOT1 (N14186, N14171);
and AND2 (N14187, N14186, N13836);
or OR2 (N14188, N14162, N11207);
nand NAND4 (N14189, N14188, N8326, N11675, N11935);
xor XOR2 (N14190, N14185, N6958);
and AND3 (N14191, N14190, N9849, N915);
xor XOR2 (N14192, N14181, N6958);
and AND2 (N14193, N14191, N11402);
nand NAND4 (N14194, N14189, N1003, N3586, N12624);
nand NAND2 (N14195, N14184, N729);
buf BUF1 (N14196, N14144);
and AND3 (N14197, N14196, N11893, N1651);
nor NOR2 (N14198, N14164, N12301);
or OR4 (N14199, N14198, N4742, N11157, N6943);
or OR4 (N14200, N14187, N12184, N12118, N8009);
buf BUF1 (N14201, N14195);
or OR3 (N14202, N14201, N9819, N11349);
xor XOR2 (N14203, N14200, N12067);
buf BUF1 (N14204, N14197);
nand NAND3 (N14205, N14177, N1592, N12067);
not NOT1 (N14206, N14192);
and AND3 (N14207, N14194, N12273, N4229);
buf BUF1 (N14208, N14199);
nand NAND3 (N14209, N14173, N10891, N10399);
not NOT1 (N14210, N14205);
xor XOR2 (N14211, N14183, N12628);
xor XOR2 (N14212, N14209, N14194);
and AND2 (N14213, N14208, N3313);
buf BUF1 (N14214, N14206);
nand NAND3 (N14215, N14212, N4958, N9263);
nand NAND3 (N14216, N14215, N13891, N8643);
not NOT1 (N14217, N14213);
and AND3 (N14218, N14202, N5354, N9833);
not NOT1 (N14219, N14211);
xor XOR2 (N14220, N14193, N4200);
buf BUF1 (N14221, N14214);
xor XOR2 (N14222, N14220, N1003);
nand NAND2 (N14223, N14222, N8971);
nor NOR4 (N14224, N14217, N8247, N3406, N13435);
or OR2 (N14225, N14219, N4600);
nor NOR3 (N14226, N14207, N2993, N5766);
and AND2 (N14227, N14216, N11016);
and AND2 (N14228, N14210, N6742);
buf BUF1 (N14229, N14203);
buf BUF1 (N14230, N14204);
buf BUF1 (N14231, N14221);
not NOT1 (N14232, N14227);
xor XOR2 (N14233, N14228, N2974);
and AND3 (N14234, N14225, N6716, N13902);
buf BUF1 (N14235, N14224);
not NOT1 (N14236, N14234);
and AND2 (N14237, N14231, N9213);
buf BUF1 (N14238, N14223);
xor XOR2 (N14239, N14237, N13588);
nor NOR3 (N14240, N14239, N11212, N3434);
xor XOR2 (N14241, N14240, N12517);
buf BUF1 (N14242, N14241);
and AND4 (N14243, N14238, N13605, N6225, N7170);
or OR2 (N14244, N14226, N7396);
buf BUF1 (N14245, N14230);
or OR3 (N14246, N14233, N2934, N13500);
xor XOR2 (N14247, N14229, N13562);
nand NAND4 (N14248, N14236, N7745, N3056, N8026);
buf BUF1 (N14249, N14232);
or OR3 (N14250, N14244, N11015, N3340);
buf BUF1 (N14251, N14245);
xor XOR2 (N14252, N14250, N4237);
nand NAND3 (N14253, N14246, N11361, N9928);
nand NAND3 (N14254, N14253, N9384, N11273);
xor XOR2 (N14255, N14247, N8782);
buf BUF1 (N14256, N14242);
nand NAND4 (N14257, N14256, N2151, N6063, N12871);
nor NOR3 (N14258, N14252, N876, N992);
nor NOR3 (N14259, N14255, N8073, N950);
nand NAND2 (N14260, N14254, N5841);
nand NAND3 (N14261, N14257, N13045, N8924);
xor XOR2 (N14262, N14218, N10962);
nand NAND3 (N14263, N14243, N2076, N5341);
xor XOR2 (N14264, N14261, N13617);
xor XOR2 (N14265, N14235, N2339);
nor NOR3 (N14266, N14260, N1075, N8847);
xor XOR2 (N14267, N14262, N13364);
xor XOR2 (N14268, N14258, N5243);
buf BUF1 (N14269, N14265);
and AND4 (N14270, N14249, N6951, N6862, N13235);
xor XOR2 (N14271, N14269, N2478);
nor NOR2 (N14272, N14259, N8857);
not NOT1 (N14273, N14272);
not NOT1 (N14274, N14271);
xor XOR2 (N14275, N14270, N10105);
and AND2 (N14276, N14267, N10334);
or OR3 (N14277, N14264, N743, N9834);
xor XOR2 (N14278, N14263, N8301);
or OR3 (N14279, N14277, N7834, N12645);
buf BUF1 (N14280, N14251);
xor XOR2 (N14281, N14268, N13828);
nor NOR3 (N14282, N14275, N588, N7875);
or OR2 (N14283, N14266, N7007);
buf BUF1 (N14284, N14273);
or OR4 (N14285, N14248, N203, N12177, N13412);
xor XOR2 (N14286, N14285, N7274);
xor XOR2 (N14287, N14282, N5002);
nor NOR3 (N14288, N14274, N10651, N1787);
nor NOR2 (N14289, N14278, N10966);
nand NAND3 (N14290, N14280, N6040, N2788);
or OR3 (N14291, N14289, N8366, N11276);
buf BUF1 (N14292, N14287);
nor NOR4 (N14293, N14291, N5377, N10964, N2162);
not NOT1 (N14294, N14288);
not NOT1 (N14295, N14292);
buf BUF1 (N14296, N14295);
or OR4 (N14297, N14284, N2208, N10166, N8973);
not NOT1 (N14298, N14286);
nor NOR4 (N14299, N14290, N576, N702, N13171);
nor NOR2 (N14300, N14299, N1911);
not NOT1 (N14301, N14276);
nand NAND2 (N14302, N14279, N11975);
buf BUF1 (N14303, N14298);
nand NAND3 (N14304, N14283, N1135, N2411);
and AND2 (N14305, N14304, N388);
buf BUF1 (N14306, N14293);
nand NAND2 (N14307, N14303, N11608);
buf BUF1 (N14308, N14307);
not NOT1 (N14309, N14297);
nor NOR2 (N14310, N14309, N4840);
nor NOR4 (N14311, N14302, N12703, N8847, N11118);
not NOT1 (N14312, N14311);
xor XOR2 (N14313, N14312, N13390);
nand NAND3 (N14314, N14301, N11252, N7604);
and AND2 (N14315, N14300, N3329);
nand NAND4 (N14316, N14296, N9492, N9860, N10607);
and AND2 (N14317, N14294, N2352);
nand NAND3 (N14318, N14308, N4039, N2757);
not NOT1 (N14319, N14281);
and AND4 (N14320, N14317, N6322, N8469, N10514);
nor NOR4 (N14321, N14314, N4417, N13863, N8080);
not NOT1 (N14322, N14305);
or OR2 (N14323, N14318, N1409);
xor XOR2 (N14324, N14320, N5453);
nor NOR2 (N14325, N14319, N11335);
not NOT1 (N14326, N14323);
xor XOR2 (N14327, N14322, N11737);
nor NOR2 (N14328, N14316, N5377);
xor XOR2 (N14329, N14315, N3043);
or OR3 (N14330, N14306, N12068, N2265);
not NOT1 (N14331, N14328);
nor NOR4 (N14332, N14330, N9963, N7281, N7699);
or OR2 (N14333, N14327, N10151);
nor NOR4 (N14334, N14332, N10605, N13049, N4503);
or OR4 (N14335, N14321, N2719, N9742, N1001);
nand NAND4 (N14336, N14324, N12842, N7699, N6157);
xor XOR2 (N14337, N14336, N12475);
not NOT1 (N14338, N14337);
xor XOR2 (N14339, N14334, N5239);
not NOT1 (N14340, N14329);
or OR4 (N14341, N14326, N10624, N6943, N5893);
xor XOR2 (N14342, N14340, N1600);
nand NAND3 (N14343, N14339, N11289, N13653);
nor NOR2 (N14344, N14341, N1052);
xor XOR2 (N14345, N14338, N6393);
or OR2 (N14346, N14325, N8333);
and AND4 (N14347, N14335, N1875, N1812, N4738);
nor NOR4 (N14348, N14347, N1037, N9451, N1400);
and AND3 (N14349, N14343, N7813, N8484);
not NOT1 (N14350, N14349);
nand NAND3 (N14351, N14350, N6994, N5003);
not NOT1 (N14352, N14344);
and AND4 (N14353, N14331, N8018, N8602, N4697);
nand NAND2 (N14354, N14348, N7246);
nor NOR4 (N14355, N14351, N11522, N159, N8518);
and AND2 (N14356, N14333, N3835);
nor NOR2 (N14357, N14342, N9997);
and AND3 (N14358, N14310, N14097, N3290);
and AND4 (N14359, N14313, N14078, N5683, N10109);
or OR4 (N14360, N14357, N8914, N210, N11316);
or OR2 (N14361, N14346, N7443);
and AND2 (N14362, N14345, N1562);
nor NOR4 (N14363, N14360, N8707, N1822, N7803);
not NOT1 (N14364, N14354);
nor NOR3 (N14365, N14353, N1495, N1816);
not NOT1 (N14366, N14355);
not NOT1 (N14367, N14363);
buf BUF1 (N14368, N14365);
xor XOR2 (N14369, N14361, N4624);
nand NAND3 (N14370, N14362, N6841, N658);
nor NOR2 (N14371, N14352, N8130);
buf BUF1 (N14372, N14367);
not NOT1 (N14373, N14359);
not NOT1 (N14374, N14370);
xor XOR2 (N14375, N14369, N7794);
and AND2 (N14376, N14375, N12246);
nor NOR2 (N14377, N14358, N1147);
and AND3 (N14378, N14364, N14184, N8731);
xor XOR2 (N14379, N14378, N12642);
not NOT1 (N14380, N14366);
buf BUF1 (N14381, N14368);
and AND3 (N14382, N14377, N10197, N3385);
not NOT1 (N14383, N14376);
nor NOR2 (N14384, N14379, N1119);
not NOT1 (N14385, N14382);
buf BUF1 (N14386, N14384);
nand NAND4 (N14387, N14372, N1948, N13436, N4377);
xor XOR2 (N14388, N14386, N13081);
nand NAND2 (N14389, N14371, N3781);
and AND3 (N14390, N14356, N3186, N8079);
xor XOR2 (N14391, N14388, N1390);
xor XOR2 (N14392, N14383, N10022);
or OR2 (N14393, N14390, N6765);
buf BUF1 (N14394, N14393);
nand NAND2 (N14395, N14380, N6370);
nor NOR4 (N14396, N14387, N436, N6321, N8401);
not NOT1 (N14397, N14389);
not NOT1 (N14398, N14397);
and AND2 (N14399, N14374, N4449);
and AND3 (N14400, N14392, N8735, N4681);
buf BUF1 (N14401, N14391);
buf BUF1 (N14402, N14385);
buf BUF1 (N14403, N14381);
not NOT1 (N14404, N14402);
not NOT1 (N14405, N14403);
xor XOR2 (N14406, N14373, N14275);
buf BUF1 (N14407, N14405);
or OR4 (N14408, N14399, N6208, N4136, N4972);
buf BUF1 (N14409, N14404);
and AND3 (N14410, N14401, N8573, N9726);
and AND2 (N14411, N14406, N807);
nor NOR2 (N14412, N14411, N1870);
nor NOR2 (N14413, N14407, N1359);
and AND2 (N14414, N14396, N4488);
buf BUF1 (N14415, N14394);
buf BUF1 (N14416, N14398);
not NOT1 (N14417, N14412);
buf BUF1 (N14418, N14416);
xor XOR2 (N14419, N14413, N1999);
xor XOR2 (N14420, N14410, N8879);
and AND4 (N14421, N14414, N13101, N1437, N14198);
buf BUF1 (N14422, N14395);
xor XOR2 (N14423, N14419, N2580);
and AND4 (N14424, N14420, N4937, N11512, N5828);
buf BUF1 (N14425, N14424);
buf BUF1 (N14426, N14422);
nand NAND3 (N14427, N14415, N7045, N11135);
xor XOR2 (N14428, N14426, N13254);
nor NOR3 (N14429, N14418, N12269, N4910);
or OR4 (N14430, N14409, N6825, N2307, N7394);
nand NAND2 (N14431, N14400, N6237);
nor NOR4 (N14432, N14431, N8253, N1721, N9822);
nor NOR2 (N14433, N14421, N407);
buf BUF1 (N14434, N14433);
nor NOR4 (N14435, N14417, N204, N3980, N4899);
nand NAND4 (N14436, N14423, N2914, N10799, N717);
xor XOR2 (N14437, N14435, N8515);
not NOT1 (N14438, N14434);
and AND2 (N14439, N14437, N7279);
nand NAND2 (N14440, N14436, N13423);
or OR2 (N14441, N14438, N10272);
not NOT1 (N14442, N14425);
not NOT1 (N14443, N14408);
not NOT1 (N14444, N14443);
xor XOR2 (N14445, N14440, N12817);
and AND2 (N14446, N14445, N1793);
nand NAND3 (N14447, N14444, N812, N1482);
and AND2 (N14448, N14446, N511);
not NOT1 (N14449, N14432);
and AND2 (N14450, N14442, N2802);
not NOT1 (N14451, N14447);
xor XOR2 (N14452, N14427, N7444);
not NOT1 (N14453, N14430);
buf BUF1 (N14454, N14451);
not NOT1 (N14455, N14450);
or OR4 (N14456, N14455, N2431, N4031, N3513);
nand NAND2 (N14457, N14439, N12498);
not NOT1 (N14458, N14452);
not NOT1 (N14459, N14429);
buf BUF1 (N14460, N14449);
nand NAND3 (N14461, N14441, N6808, N3046);
and AND4 (N14462, N14460, N261, N4579, N10791);
not NOT1 (N14463, N14458);
buf BUF1 (N14464, N14462);
buf BUF1 (N14465, N14456);
buf BUF1 (N14466, N14457);
nand NAND4 (N14467, N14461, N10213, N7966, N568);
or OR3 (N14468, N14466, N2755, N6310);
nor NOR2 (N14469, N14453, N8008);
nand NAND2 (N14470, N14448, N2812);
xor XOR2 (N14471, N14459, N3835);
and AND3 (N14472, N14465, N3332, N9567);
nand NAND3 (N14473, N14428, N4710, N130);
nor NOR4 (N14474, N14454, N11590, N13589, N3069);
and AND2 (N14475, N14467, N3121);
nor NOR2 (N14476, N14471, N11834);
xor XOR2 (N14477, N14464, N12355);
nor NOR2 (N14478, N14474, N8041);
nor NOR4 (N14479, N14470, N1749, N5300, N350);
not NOT1 (N14480, N14476);
nor NOR4 (N14481, N14463, N304, N12437, N4096);
nand NAND3 (N14482, N14469, N7110, N6704);
or OR4 (N14483, N14475, N11522, N8141, N5817);
not NOT1 (N14484, N14481);
buf BUF1 (N14485, N14479);
and AND2 (N14486, N14480, N9174);
or OR3 (N14487, N14484, N8962, N141);
and AND4 (N14488, N14478, N13511, N3690, N5125);
buf BUF1 (N14489, N14483);
buf BUF1 (N14490, N14485);
nor NOR3 (N14491, N14482, N12644, N12223);
not NOT1 (N14492, N14473);
not NOT1 (N14493, N14486);
or OR2 (N14494, N14491, N13233);
nor NOR4 (N14495, N14488, N14373, N8510, N3816);
nor NOR2 (N14496, N14472, N7897);
nor NOR2 (N14497, N14489, N9754);
not NOT1 (N14498, N14487);
buf BUF1 (N14499, N14468);
buf BUF1 (N14500, N14494);
xor XOR2 (N14501, N14493, N3987);
nor NOR4 (N14502, N14496, N3548, N6353, N5664);
nor NOR3 (N14503, N14498, N14069, N5402);
nor NOR3 (N14504, N14501, N1740, N65);
and AND3 (N14505, N14490, N2009, N4300);
not NOT1 (N14506, N14504);
and AND4 (N14507, N14497, N9495, N1265, N10811);
not NOT1 (N14508, N14500);
not NOT1 (N14509, N14495);
and AND4 (N14510, N14505, N547, N1625, N9510);
nor NOR4 (N14511, N14508, N2897, N8892, N8389);
nand NAND4 (N14512, N14477, N3016, N2795, N12310);
buf BUF1 (N14513, N14503);
not NOT1 (N14514, N14499);
not NOT1 (N14515, N14509);
xor XOR2 (N14516, N14512, N9206);
not NOT1 (N14517, N14515);
or OR2 (N14518, N14517, N4699);
nor NOR3 (N14519, N14506, N6888, N7384);
not NOT1 (N14520, N14507);
nand NAND2 (N14521, N14514, N10418);
and AND3 (N14522, N14502, N13175, N13533);
and AND3 (N14523, N14522, N8445, N2824);
and AND2 (N14524, N14516, N8313);
buf BUF1 (N14525, N14510);
or OR2 (N14526, N14524, N1838);
nand NAND2 (N14527, N14526, N6106);
buf BUF1 (N14528, N14513);
not NOT1 (N14529, N14520);
and AND2 (N14530, N14528, N12162);
buf BUF1 (N14531, N14530);
nand NAND4 (N14532, N14519, N5656, N14093, N201);
buf BUF1 (N14533, N14529);
not NOT1 (N14534, N14492);
or OR4 (N14535, N14525, N9190, N136, N5315);
or OR4 (N14536, N14535, N6867, N1997, N2172);
xor XOR2 (N14537, N14536, N9473);
buf BUF1 (N14538, N14534);
nor NOR4 (N14539, N14537, N10150, N4194, N10922);
and AND4 (N14540, N14523, N10372, N5990, N11337);
xor XOR2 (N14541, N14527, N5258);
xor XOR2 (N14542, N14539, N6514);
and AND2 (N14543, N14532, N3553);
and AND2 (N14544, N14543, N5513);
or OR2 (N14545, N14540, N115);
xor XOR2 (N14546, N14511, N8603);
xor XOR2 (N14547, N14533, N13081);
or OR2 (N14548, N14546, N4083);
nand NAND3 (N14549, N14541, N8153, N12298);
or OR4 (N14550, N14548, N4436, N4928, N10061);
or OR3 (N14551, N14531, N3625, N10928);
not NOT1 (N14552, N14538);
xor XOR2 (N14553, N14542, N10402);
buf BUF1 (N14554, N14544);
nor NOR4 (N14555, N14549, N5054, N14489, N13524);
buf BUF1 (N14556, N14555);
buf BUF1 (N14557, N14551);
nand NAND2 (N14558, N14557, N11712);
buf BUF1 (N14559, N14550);
and AND3 (N14560, N14518, N8586, N9955);
not NOT1 (N14561, N14560);
not NOT1 (N14562, N14547);
xor XOR2 (N14563, N14554, N6930);
nand NAND3 (N14564, N14521, N9363, N5036);
xor XOR2 (N14565, N14559, N3260);
xor XOR2 (N14566, N14553, N8207);
nand NAND3 (N14567, N14563, N282, N1733);
xor XOR2 (N14568, N14561, N10097);
not NOT1 (N14569, N14564);
and AND2 (N14570, N14558, N6042);
nand NAND4 (N14571, N14552, N6162, N7064, N6642);
or OR3 (N14572, N14567, N8322, N62);
buf BUF1 (N14573, N14571);
nor NOR2 (N14574, N14545, N7605);
and AND4 (N14575, N14568, N9911, N8279, N8964);
and AND3 (N14576, N14566, N6255, N13727);
or OR4 (N14577, N14573, N4716, N4566, N11671);
and AND2 (N14578, N14577, N6443);
or OR3 (N14579, N14575, N6254, N7362);
nor NOR2 (N14580, N14570, N8238);
not NOT1 (N14581, N14572);
buf BUF1 (N14582, N14562);
not NOT1 (N14583, N14556);
or OR4 (N14584, N14569, N2954, N13980, N9308);
nor NOR4 (N14585, N14574, N2057, N4502, N6020);
and AND4 (N14586, N14576, N10844, N691, N14387);
xor XOR2 (N14587, N14582, N4036);
and AND2 (N14588, N14581, N1578);
not NOT1 (N14589, N14584);
nor NOR4 (N14590, N14578, N10837, N1172, N6748);
buf BUF1 (N14591, N14590);
and AND3 (N14592, N14565, N13497, N13944);
and AND3 (N14593, N14580, N7066, N6449);
not NOT1 (N14594, N14588);
buf BUF1 (N14595, N14594);
or OR2 (N14596, N14591, N3666);
buf BUF1 (N14597, N14583);
xor XOR2 (N14598, N14596, N3426);
not NOT1 (N14599, N14598);
not NOT1 (N14600, N14597);
buf BUF1 (N14601, N14585);
buf BUF1 (N14602, N14601);
nor NOR3 (N14603, N14595, N9223, N3075);
and AND4 (N14604, N14600, N11875, N2192, N12871);
or OR4 (N14605, N14587, N7073, N9106, N7097);
or OR2 (N14606, N14579, N745);
buf BUF1 (N14607, N14603);
nor NOR2 (N14608, N14604, N8507);
xor XOR2 (N14609, N14589, N9417);
nand NAND2 (N14610, N14606, N10805);
nor NOR2 (N14611, N14607, N4876);
nand NAND3 (N14612, N14609, N9772, N11524);
buf BUF1 (N14613, N14592);
nor NOR4 (N14614, N14613, N242, N9776, N7713);
nor NOR3 (N14615, N14610, N3606, N8867);
or OR3 (N14616, N14615, N8093, N9295);
xor XOR2 (N14617, N14599, N3771);
and AND2 (N14618, N14616, N5598);
not NOT1 (N14619, N14586);
and AND3 (N14620, N14619, N12843, N4212);
xor XOR2 (N14621, N14618, N2341);
not NOT1 (N14622, N14611);
nor NOR2 (N14623, N14608, N14353);
buf BUF1 (N14624, N14605);
nand NAND3 (N14625, N14617, N4422, N3365);
nor NOR4 (N14626, N14624, N2852, N10949, N648);
buf BUF1 (N14627, N14625);
or OR3 (N14628, N14614, N368, N13752);
buf BUF1 (N14629, N14628);
nor NOR2 (N14630, N14602, N13057);
buf BUF1 (N14631, N14627);
xor XOR2 (N14632, N14621, N1191);
nor NOR4 (N14633, N14626, N13037, N7843, N12365);
and AND4 (N14634, N14622, N8729, N3182, N14295);
nand NAND2 (N14635, N14631, N6036);
or OR3 (N14636, N14623, N9781, N14275);
xor XOR2 (N14637, N14630, N6847);
nand NAND3 (N14638, N14636, N1554, N7919);
or OR4 (N14639, N14612, N6979, N11791, N8385);
nand NAND2 (N14640, N14632, N1152);
nand NAND2 (N14641, N14593, N5733);
and AND4 (N14642, N14640, N4780, N11816, N13291);
not NOT1 (N14643, N14634);
or OR4 (N14644, N14620, N10080, N10810, N11304);
nor NOR3 (N14645, N14638, N10873, N2784);
nor NOR3 (N14646, N14645, N1186, N2244);
not NOT1 (N14647, N14635);
xor XOR2 (N14648, N14646, N160);
or OR4 (N14649, N14648, N4537, N7099, N12314);
nor NOR2 (N14650, N14641, N7583);
nor NOR2 (N14651, N14642, N10529);
nor NOR2 (N14652, N14643, N14056);
not NOT1 (N14653, N14644);
nor NOR2 (N14654, N14649, N1939);
and AND4 (N14655, N14629, N9834, N4416, N13439);
nand NAND2 (N14656, N14652, N9042);
or OR3 (N14657, N14651, N9349, N7434);
not NOT1 (N14658, N14637);
and AND4 (N14659, N14639, N10105, N9515, N9965);
and AND2 (N14660, N14650, N6195);
xor XOR2 (N14661, N14655, N13795);
xor XOR2 (N14662, N14659, N5917);
or OR3 (N14663, N14661, N6089, N240);
xor XOR2 (N14664, N14633, N9133);
or OR3 (N14665, N14658, N12133, N7285);
not NOT1 (N14666, N14660);
not NOT1 (N14667, N14663);
nand NAND2 (N14668, N14666, N5733);
xor XOR2 (N14669, N14664, N4954);
xor XOR2 (N14670, N14653, N11700);
xor XOR2 (N14671, N14654, N12090);
not NOT1 (N14672, N14662);
nand NAND2 (N14673, N14665, N2426);
and AND3 (N14674, N14656, N7173, N13655);
xor XOR2 (N14675, N14673, N6673);
nor NOR2 (N14676, N14670, N4085);
buf BUF1 (N14677, N14674);
not NOT1 (N14678, N14647);
or OR4 (N14679, N14672, N24, N11035, N3895);
buf BUF1 (N14680, N14667);
nand NAND4 (N14681, N14679, N7518, N107, N10454);
or OR4 (N14682, N14681, N557, N4826, N3805);
not NOT1 (N14683, N14669);
not NOT1 (N14684, N14683);
xor XOR2 (N14685, N14676, N11471);
nand NAND4 (N14686, N14682, N11555, N12909, N11509);
nor NOR4 (N14687, N14686, N8492, N1784, N3336);
nor NOR3 (N14688, N14677, N13422, N3197);
buf BUF1 (N14689, N14688);
xor XOR2 (N14690, N14684, N13540);
or OR3 (N14691, N14668, N6306, N12814);
nand NAND3 (N14692, N14689, N10909, N3223);
not NOT1 (N14693, N14678);
not NOT1 (N14694, N14692);
buf BUF1 (N14695, N14671);
buf BUF1 (N14696, N14693);
xor XOR2 (N14697, N14685, N7190);
xor XOR2 (N14698, N14690, N9207);
xor XOR2 (N14699, N14687, N1269);
buf BUF1 (N14700, N14698);
buf BUF1 (N14701, N14691);
nand NAND2 (N14702, N14680, N3581);
nand NAND3 (N14703, N14694, N6984, N4997);
nand NAND4 (N14704, N14675, N1028, N6428, N10262);
xor XOR2 (N14705, N14696, N9755);
or OR4 (N14706, N14702, N14603, N13098, N8302);
nor NOR3 (N14707, N14697, N8980, N7985);
xor XOR2 (N14708, N14703, N1529);
nand NAND3 (N14709, N14699, N1421, N5541);
or OR4 (N14710, N14701, N2378, N11913, N7131);
xor XOR2 (N14711, N14710, N5992);
not NOT1 (N14712, N14657);
or OR3 (N14713, N14705, N7383, N10010);
not NOT1 (N14714, N14704);
buf BUF1 (N14715, N14711);
and AND4 (N14716, N14700, N13989, N11496, N13576);
and AND2 (N14717, N14709, N10795);
and AND4 (N14718, N14712, N7060, N2070, N13260);
nor NOR2 (N14719, N14717, N1478);
xor XOR2 (N14720, N14716, N7842);
nand NAND2 (N14721, N14715, N12276);
not NOT1 (N14722, N14721);
or OR4 (N14723, N14713, N829, N8262, N979);
xor XOR2 (N14724, N14695, N6226);
nand NAND4 (N14725, N14720, N6904, N359, N13902);
xor XOR2 (N14726, N14714, N12972);
or OR3 (N14727, N14725, N12655, N13531);
or OR3 (N14728, N14708, N8516, N2724);
buf BUF1 (N14729, N14724);
or OR4 (N14730, N14728, N8462, N13701, N5003);
nand NAND3 (N14731, N14729, N9667, N4953);
nor NOR2 (N14732, N14722, N7674);
xor XOR2 (N14733, N14719, N3230);
nor NOR4 (N14734, N14726, N6052, N5036, N340);
not NOT1 (N14735, N14730);
and AND2 (N14736, N14733, N7211);
not NOT1 (N14737, N14735);
or OR3 (N14738, N14723, N6886, N10759);
nor NOR3 (N14739, N14732, N3896, N14661);
not NOT1 (N14740, N14706);
not NOT1 (N14741, N14737);
not NOT1 (N14742, N14707);
nand NAND4 (N14743, N14718, N5411, N1793, N8294);
buf BUF1 (N14744, N14740);
xor XOR2 (N14745, N14744, N11912);
nand NAND2 (N14746, N14742, N11425);
nand NAND2 (N14747, N14739, N13735);
or OR4 (N14748, N14747, N9081, N1399, N916);
or OR4 (N14749, N14745, N1310, N11551, N13677);
and AND2 (N14750, N14743, N12497);
or OR4 (N14751, N14734, N12400, N1561, N6537);
or OR2 (N14752, N14741, N7682);
and AND4 (N14753, N14752, N5426, N9604, N248);
or OR3 (N14754, N14749, N2443, N2766);
and AND3 (N14755, N14736, N11419, N2574);
nand NAND2 (N14756, N14748, N6977);
not NOT1 (N14757, N14754);
nor NOR4 (N14758, N14755, N7372, N2568, N2677);
buf BUF1 (N14759, N14727);
nand NAND2 (N14760, N14759, N11079);
buf BUF1 (N14761, N14751);
or OR4 (N14762, N14750, N4576, N1974, N5662);
not NOT1 (N14763, N14758);
xor XOR2 (N14764, N14761, N13607);
xor XOR2 (N14765, N14756, N2411);
xor XOR2 (N14766, N14765, N2846);
nor NOR2 (N14767, N14746, N13478);
and AND2 (N14768, N14762, N511);
not NOT1 (N14769, N14768);
and AND2 (N14770, N14766, N1733);
not NOT1 (N14771, N14764);
xor XOR2 (N14772, N14767, N3865);
nand NAND4 (N14773, N14753, N8268, N13127, N4776);
nor NOR3 (N14774, N14738, N3327, N6462);
not NOT1 (N14775, N14770);
nor NOR3 (N14776, N14773, N11163, N13198);
or OR4 (N14777, N14763, N2834, N3122, N3282);
not NOT1 (N14778, N14772);
not NOT1 (N14779, N14731);
not NOT1 (N14780, N14757);
not NOT1 (N14781, N14779);
nor NOR2 (N14782, N14777, N1014);
buf BUF1 (N14783, N14781);
or OR3 (N14784, N14774, N449, N12480);
buf BUF1 (N14785, N14760);
not NOT1 (N14786, N14780);
not NOT1 (N14787, N14776);
xor XOR2 (N14788, N14783, N3099);
xor XOR2 (N14789, N14782, N6262);
buf BUF1 (N14790, N14787);
nor NOR3 (N14791, N14789, N2619, N4002);
and AND3 (N14792, N14790, N7091, N8706);
nor NOR4 (N14793, N14784, N11166, N1209, N12263);
or OR3 (N14794, N14788, N3109, N3275);
nand NAND4 (N14795, N14791, N11774, N13221, N3316);
nand NAND3 (N14796, N14794, N10962, N10609);
not NOT1 (N14797, N14775);
nor NOR2 (N14798, N14769, N4742);
or OR2 (N14799, N14796, N3182);
xor XOR2 (N14800, N14798, N11263);
xor XOR2 (N14801, N14786, N11981);
nor NOR3 (N14802, N14771, N12275, N14610);
buf BUF1 (N14803, N14802);
xor XOR2 (N14804, N14801, N1250);
and AND3 (N14805, N14795, N13638, N4359);
and AND4 (N14806, N14800, N5236, N2213, N9229);
xor XOR2 (N14807, N14806, N9870);
xor XOR2 (N14808, N14792, N7866);
xor XOR2 (N14809, N14808, N11641);
nor NOR2 (N14810, N14809, N14440);
or OR2 (N14811, N14803, N4545);
buf BUF1 (N14812, N14807);
nand NAND4 (N14813, N14797, N8710, N6971, N5113);
nor NOR4 (N14814, N14785, N10899, N9761, N11107);
or OR2 (N14815, N14810, N4329);
xor XOR2 (N14816, N14812, N11884);
or OR3 (N14817, N14799, N1795, N13531);
not NOT1 (N14818, N14813);
or OR4 (N14819, N14814, N299, N2810, N4487);
not NOT1 (N14820, N14793);
nand NAND4 (N14821, N14805, N8730, N4814, N11917);
or OR3 (N14822, N14815, N4059, N4401);
nand NAND4 (N14823, N14811, N8329, N8712, N10092);
nor NOR4 (N14824, N14821, N14660, N5438, N10444);
buf BUF1 (N14825, N14816);
and AND2 (N14826, N14817, N5039);
or OR2 (N14827, N14824, N1921);
or OR4 (N14828, N14820, N7211, N9913, N4700);
not NOT1 (N14829, N14825);
or OR2 (N14830, N14826, N7063);
not NOT1 (N14831, N14804);
nor NOR3 (N14832, N14827, N10829, N7203);
not NOT1 (N14833, N14828);
nand NAND2 (N14834, N14778, N2769);
buf BUF1 (N14835, N14822);
xor XOR2 (N14836, N14830, N9589);
buf BUF1 (N14837, N14834);
and AND2 (N14838, N14819, N10637);
xor XOR2 (N14839, N14836, N8);
xor XOR2 (N14840, N14831, N3303);
or OR2 (N14841, N14832, N5663);
nand NAND4 (N14842, N14818, N1909, N1717, N14431);
or OR3 (N14843, N14840, N3731, N971);
and AND2 (N14844, N14833, N8737);
or OR3 (N14845, N14835, N11902, N1858);
buf BUF1 (N14846, N14843);
not NOT1 (N14847, N14838);
or OR3 (N14848, N14839, N1744, N5113);
nor NOR2 (N14849, N14829, N11683);
not NOT1 (N14850, N14847);
nor NOR3 (N14851, N14848, N14408, N7589);
nor NOR4 (N14852, N14850, N5822, N8305, N522);
buf BUF1 (N14853, N14837);
and AND4 (N14854, N14823, N13393, N2411, N10719);
or OR3 (N14855, N14841, N5555, N10164);
buf BUF1 (N14856, N14845);
buf BUF1 (N14857, N14851);
xor XOR2 (N14858, N14852, N1495);
not NOT1 (N14859, N14854);
nor NOR2 (N14860, N14849, N837);
nand NAND3 (N14861, N14853, N4606, N10614);
xor XOR2 (N14862, N14861, N14741);
nand NAND3 (N14863, N14855, N2027, N7265);
nand NAND4 (N14864, N14842, N7679, N2421, N8193);
nor NOR4 (N14865, N14864, N5832, N10109, N10257);
buf BUF1 (N14866, N14859);
nor NOR2 (N14867, N14846, N4847);
and AND4 (N14868, N14867, N8996, N4778, N2382);
and AND2 (N14869, N14856, N9986);
or OR4 (N14870, N14860, N14125, N4155, N774);
buf BUF1 (N14871, N14857);
nand NAND4 (N14872, N14868, N12670, N12809, N5220);
xor XOR2 (N14873, N14870, N8016);
xor XOR2 (N14874, N14858, N8670);
nor NOR3 (N14875, N14874, N3436, N9394);
and AND3 (N14876, N14862, N5117, N1725);
nor NOR2 (N14877, N14872, N3197);
buf BUF1 (N14878, N14869);
not NOT1 (N14879, N14875);
buf BUF1 (N14880, N14865);
not NOT1 (N14881, N14871);
nand NAND3 (N14882, N14866, N9874, N8009);
nor NOR4 (N14883, N14876, N14574, N4798, N9205);
not NOT1 (N14884, N14880);
not NOT1 (N14885, N14877);
or OR3 (N14886, N14879, N12399, N1805);
xor XOR2 (N14887, N14844, N2410);
nor NOR2 (N14888, N14887, N8757);
and AND4 (N14889, N14878, N6029, N2121, N6911);
nor NOR4 (N14890, N14863, N1163, N11835, N1414);
and AND4 (N14891, N14882, N11248, N580, N6239);
and AND4 (N14892, N14891, N1578, N2358, N6979);
nand NAND4 (N14893, N14890, N8231, N911, N7444);
xor XOR2 (N14894, N14886, N10624);
and AND3 (N14895, N14881, N1485, N4771);
or OR3 (N14896, N14884, N2326, N2125);
xor XOR2 (N14897, N14883, N9434);
not NOT1 (N14898, N14889);
and AND2 (N14899, N14885, N8447);
nand NAND2 (N14900, N14896, N556);
nor NOR2 (N14901, N14894, N13685);
not NOT1 (N14902, N14873);
and AND4 (N14903, N14898, N321, N11715, N4836);
not NOT1 (N14904, N14893);
and AND4 (N14905, N14904, N6931, N12006, N1503);
not NOT1 (N14906, N14905);
and AND4 (N14907, N14902, N1117, N1514, N5337);
xor XOR2 (N14908, N14903, N5157);
or OR3 (N14909, N14895, N7511, N7077);
or OR2 (N14910, N14901, N14708);
nand NAND4 (N14911, N14888, N10570, N1936, N2309);
and AND2 (N14912, N14907, N8742);
xor XOR2 (N14913, N14892, N8312);
buf BUF1 (N14914, N14909);
xor XOR2 (N14915, N14911, N1391);
or OR4 (N14916, N14900, N10136, N8222, N6383);
buf BUF1 (N14917, N14899);
buf BUF1 (N14918, N14908);
or OR3 (N14919, N14915, N1748, N2999);
xor XOR2 (N14920, N14918, N4509);
buf BUF1 (N14921, N14897);
buf BUF1 (N14922, N14919);
buf BUF1 (N14923, N14912);
xor XOR2 (N14924, N14922, N7312);
nand NAND3 (N14925, N14921, N10518, N12518);
or OR2 (N14926, N14906, N562);
and AND3 (N14927, N14916, N13082, N9736);
not NOT1 (N14928, N14925);
not NOT1 (N14929, N14926);
nor NOR3 (N14930, N14924, N9300, N1733);
or OR3 (N14931, N14928, N13772, N5332);
xor XOR2 (N14932, N14910, N9451);
xor XOR2 (N14933, N14932, N12924);
nor NOR4 (N14934, N14933, N5418, N1525, N11115);
nand NAND2 (N14935, N14929, N6020);
or OR4 (N14936, N14935, N4598, N14140, N13277);
nor NOR3 (N14937, N14930, N10740, N603);
buf BUF1 (N14938, N14931);
xor XOR2 (N14939, N14938, N10744);
and AND2 (N14940, N14920, N6381);
nor NOR3 (N14941, N14939, N6078, N68);
nand NAND2 (N14942, N14917, N8547);
nand NAND3 (N14943, N14927, N3364, N6771);
buf BUF1 (N14944, N14914);
xor XOR2 (N14945, N14923, N6816);
or OR2 (N14946, N14940, N14739);
buf BUF1 (N14947, N14936);
xor XOR2 (N14948, N14913, N14740);
or OR2 (N14949, N14943, N3061);
and AND4 (N14950, N14946, N14646, N1295, N9900);
or OR3 (N14951, N14942, N14296, N4840);
nand NAND2 (N14952, N14934, N4820);
and AND2 (N14953, N14945, N5233);
and AND4 (N14954, N14937, N8330, N7103, N6459);
or OR2 (N14955, N14948, N3431);
xor XOR2 (N14956, N14950, N4962);
not NOT1 (N14957, N14953);
or OR3 (N14958, N14957, N10184, N3542);
buf BUF1 (N14959, N14944);
nor NOR4 (N14960, N14959, N9952, N2407, N479);
not NOT1 (N14961, N14949);
xor XOR2 (N14962, N14954, N5026);
or OR3 (N14963, N14952, N3771, N7150);
buf BUF1 (N14964, N14947);
nand NAND3 (N14965, N14955, N14127, N10385);
xor XOR2 (N14966, N14958, N4739);
or OR4 (N14967, N14956, N10340, N503, N9754);
not NOT1 (N14968, N14960);
nand NAND2 (N14969, N14968, N6101);
not NOT1 (N14970, N14951);
buf BUF1 (N14971, N14970);
xor XOR2 (N14972, N14963, N14678);
not NOT1 (N14973, N14962);
buf BUF1 (N14974, N14969);
buf BUF1 (N14975, N14972);
xor XOR2 (N14976, N14964, N2966);
xor XOR2 (N14977, N14965, N12895);
nand NAND3 (N14978, N14977, N5450, N13273);
or OR3 (N14979, N14978, N12331, N5994);
and AND2 (N14980, N14973, N4848);
or OR2 (N14981, N14961, N9219);
not NOT1 (N14982, N14975);
nand NAND2 (N14983, N14974, N5713);
xor XOR2 (N14984, N14971, N7713);
nor NOR2 (N14985, N14966, N1804);
and AND3 (N14986, N14981, N2784, N4317);
and AND4 (N14987, N14983, N9913, N6556, N1986);
nor NOR3 (N14988, N14979, N3482, N17);
buf BUF1 (N14989, N14982);
and AND3 (N14990, N14986, N10095, N1592);
or OR2 (N14991, N14967, N12953);
and AND3 (N14992, N14941, N10714, N11023);
and AND3 (N14993, N14990, N5567, N3949);
xor XOR2 (N14994, N14985, N8145);
xor XOR2 (N14995, N14993, N2018);
nand NAND2 (N14996, N14976, N412);
buf BUF1 (N14997, N14987);
buf BUF1 (N14998, N14984);
buf BUF1 (N14999, N14991);
xor XOR2 (N15000, N14992, N3996);
or OR2 (N15001, N14988, N10441);
nor NOR3 (N15002, N14997, N10841, N392);
or OR2 (N15003, N15001, N3630);
nand NAND4 (N15004, N15002, N2839, N4198, N3938);
buf BUF1 (N15005, N14999);
buf BUF1 (N15006, N15004);
not NOT1 (N15007, N15006);
or OR3 (N15008, N15007, N9530, N7733);
buf BUF1 (N15009, N14994);
xor XOR2 (N15010, N15000, N14907);
nor NOR2 (N15011, N15009, N416);
nor NOR3 (N15012, N14996, N7077, N12218);
not NOT1 (N15013, N15011);
buf BUF1 (N15014, N15003);
nand NAND3 (N15015, N14989, N11838, N1994);
nor NOR3 (N15016, N15005, N3546, N5538);
nor NOR2 (N15017, N15008, N5741);
or OR4 (N15018, N15010, N13292, N4429, N12144);
xor XOR2 (N15019, N15016, N7952);
nand NAND2 (N15020, N14998, N12088);
not NOT1 (N15021, N15015);
nand NAND3 (N15022, N15014, N12248, N5079);
and AND3 (N15023, N14980, N14989, N11158);
or OR2 (N15024, N15022, N4323);
and AND3 (N15025, N14995, N6645, N14106);
or OR2 (N15026, N15013, N12302);
or OR2 (N15027, N15019, N5370);
nand NAND3 (N15028, N15021, N14025, N8953);
xor XOR2 (N15029, N15017, N9705);
nand NAND2 (N15030, N15023, N5537);
and AND4 (N15031, N15024, N3474, N12018, N6474);
and AND2 (N15032, N15027, N9640);
nor NOR3 (N15033, N15030, N12865, N740);
nor NOR3 (N15034, N15018, N7, N5204);
xor XOR2 (N15035, N15025, N3247);
or OR3 (N15036, N15028, N10368, N12751);
buf BUF1 (N15037, N15033);
nor NOR2 (N15038, N15035, N7648);
nor NOR3 (N15039, N15029, N1426, N9566);
or OR4 (N15040, N15012, N6151, N6101, N5227);
nor NOR3 (N15041, N15036, N2953, N14383);
xor XOR2 (N15042, N15040, N11817);
buf BUF1 (N15043, N15041);
xor XOR2 (N15044, N15043, N5032);
nor NOR4 (N15045, N15044, N9234, N5258, N10821);
buf BUF1 (N15046, N15037);
not NOT1 (N15047, N15031);
nor NOR3 (N15048, N15020, N1739, N14323);
nand NAND2 (N15049, N15047, N3989);
not NOT1 (N15050, N15045);
buf BUF1 (N15051, N15050);
and AND4 (N15052, N15038, N9294, N5958, N7207);
xor XOR2 (N15053, N15042, N3832);
or OR4 (N15054, N15051, N4683, N4825, N1540);
buf BUF1 (N15055, N15053);
buf BUF1 (N15056, N15054);
xor XOR2 (N15057, N15034, N5199);
and AND3 (N15058, N15049, N9406, N6559);
xor XOR2 (N15059, N15039, N2003);
xor XOR2 (N15060, N15056, N14393);
nand NAND2 (N15061, N15059, N1991);
or OR4 (N15062, N15055, N14144, N5873, N2557);
nor NOR4 (N15063, N15048, N3650, N5493, N13695);
nor NOR2 (N15064, N15061, N14965);
nand NAND4 (N15065, N15062, N8433, N6639, N2646);
not NOT1 (N15066, N15052);
or OR4 (N15067, N15058, N6009, N11884, N12722);
buf BUF1 (N15068, N15065);
buf BUF1 (N15069, N15063);
nor NOR2 (N15070, N15060, N8510);
and AND4 (N15071, N15032, N6745, N2494, N6742);
nor NOR2 (N15072, N15067, N1832);
nand NAND3 (N15073, N15046, N9489, N13432);
not NOT1 (N15074, N15073);
xor XOR2 (N15075, N15057, N4239);
nor NOR4 (N15076, N15070, N11604, N1069, N5057);
nor NOR4 (N15077, N15026, N5482, N8213, N4102);
nand NAND4 (N15078, N15068, N3989, N8742, N4191);
and AND2 (N15079, N15076, N14861);
or OR4 (N15080, N15069, N228, N2580, N7683);
nor NOR3 (N15081, N15066, N9393, N9908);
not NOT1 (N15082, N15071);
xor XOR2 (N15083, N15082, N14531);
or OR4 (N15084, N15077, N8804, N5837, N4156);
nor NOR3 (N15085, N15064, N12200, N5247);
not NOT1 (N15086, N15080);
nand NAND4 (N15087, N15075, N12959, N9142, N13645);
or OR4 (N15088, N15078, N1088, N13365, N14204);
nor NOR4 (N15089, N15088, N12683, N6414, N4772);
nor NOR3 (N15090, N15081, N8623, N10604);
xor XOR2 (N15091, N15086, N7275);
buf BUF1 (N15092, N15087);
nor NOR4 (N15093, N15084, N6220, N7538, N4890);
xor XOR2 (N15094, N15092, N10218);
nor NOR3 (N15095, N15094, N4090, N11298);
nor NOR4 (N15096, N15072, N617, N766, N9901);
buf BUF1 (N15097, N15091);
nor NOR4 (N15098, N15089, N12554, N1685, N3531);
and AND4 (N15099, N15098, N14813, N5030, N588);
and AND4 (N15100, N15099, N3188, N12812, N2441);
xor XOR2 (N15101, N15090, N7738);
nor NOR3 (N15102, N15083, N7548, N11397);
nor NOR2 (N15103, N15100, N813);
buf BUF1 (N15104, N15103);
buf BUF1 (N15105, N15079);
nand NAND3 (N15106, N15102, N8823, N14252);
or OR4 (N15107, N15101, N4508, N4230, N14935);
nor NOR3 (N15108, N15104, N11140, N7314);
xor XOR2 (N15109, N15093, N1109);
not NOT1 (N15110, N15108);
xor XOR2 (N15111, N15106, N9141);
buf BUF1 (N15112, N15111);
not NOT1 (N15113, N15085);
nor NOR3 (N15114, N15113, N9936, N10369);
and AND2 (N15115, N15097, N10158);
or OR3 (N15116, N15115, N7124, N6309);
xor XOR2 (N15117, N15095, N537);
xor XOR2 (N15118, N15105, N11129);
nor NOR2 (N15119, N15114, N15010);
not NOT1 (N15120, N15074);
buf BUF1 (N15121, N15120);
nor NOR4 (N15122, N15118, N8653, N1217, N12032);
and AND4 (N15123, N15116, N10801, N11611, N8162);
nand NAND3 (N15124, N15122, N14609, N10733);
xor XOR2 (N15125, N15123, N9906);
nand NAND4 (N15126, N15096, N4861, N8911, N10419);
not NOT1 (N15127, N15107);
not NOT1 (N15128, N15121);
or OR3 (N15129, N15125, N9890, N8362);
xor XOR2 (N15130, N15124, N13535);
buf BUF1 (N15131, N15112);
or OR4 (N15132, N15130, N4621, N6004, N9573);
not NOT1 (N15133, N15127);
buf BUF1 (N15134, N15128);
or OR2 (N15135, N15109, N10185);
or OR2 (N15136, N15126, N10308);
nand NAND2 (N15137, N15129, N3970);
buf BUF1 (N15138, N15137);
or OR4 (N15139, N15132, N478, N3319, N1359);
xor XOR2 (N15140, N15131, N91);
not NOT1 (N15141, N15110);
nand NAND2 (N15142, N15117, N712);
not NOT1 (N15143, N15142);
nand NAND3 (N15144, N15141, N8603, N13393);
nor NOR3 (N15145, N15134, N3592, N6261);
nand NAND2 (N15146, N15140, N6135);
xor XOR2 (N15147, N15143, N5916);
or OR3 (N15148, N15135, N11065, N10783);
nand NAND2 (N15149, N15138, N2869);
nor NOR4 (N15150, N15146, N12316, N11889, N2714);
nand NAND2 (N15151, N15148, N479);
xor XOR2 (N15152, N15149, N3790);
buf BUF1 (N15153, N15119);
nor NOR4 (N15154, N15151, N10151, N10647, N1193);
xor XOR2 (N15155, N15133, N7956);
nor NOR2 (N15156, N15136, N2772);
not NOT1 (N15157, N15144);
or OR3 (N15158, N15153, N1507, N9351);
not NOT1 (N15159, N15156);
nor NOR4 (N15160, N15152, N6826, N11154, N1297);
not NOT1 (N15161, N15155);
and AND3 (N15162, N15150, N11170, N388);
or OR2 (N15163, N15154, N13433);
nand NAND4 (N15164, N15145, N6414, N3952, N4945);
nor NOR3 (N15165, N15159, N6684, N7071);
and AND2 (N15166, N15158, N7131);
and AND2 (N15167, N15161, N8530);
nand NAND4 (N15168, N15165, N10425, N14966, N2588);
or OR3 (N15169, N15164, N11233, N7054);
or OR4 (N15170, N15157, N15072, N4371, N13783);
buf BUF1 (N15171, N15162);
nand NAND2 (N15172, N15171, N8149);
not NOT1 (N15173, N15160);
xor XOR2 (N15174, N15167, N11783);
nor NOR2 (N15175, N15139, N5550);
or OR2 (N15176, N15170, N10958);
xor XOR2 (N15177, N15175, N342);
and AND3 (N15178, N15147, N6313, N7154);
or OR3 (N15179, N15168, N7274, N2002);
buf BUF1 (N15180, N15178);
not NOT1 (N15181, N15180);
or OR3 (N15182, N15172, N2118, N8238);
xor XOR2 (N15183, N15181, N3694);
or OR4 (N15184, N15174, N3241, N12839, N6693);
buf BUF1 (N15185, N15184);
not NOT1 (N15186, N15179);
xor XOR2 (N15187, N15176, N15161);
or OR3 (N15188, N15187, N8024, N12095);
not NOT1 (N15189, N15185);
not NOT1 (N15190, N15186);
nor NOR3 (N15191, N15177, N5004, N982);
buf BUF1 (N15192, N15191);
nand NAND3 (N15193, N15192, N7863, N820);
not NOT1 (N15194, N15193);
xor XOR2 (N15195, N15163, N10917);
not NOT1 (N15196, N15173);
nor NOR4 (N15197, N15195, N4745, N10398, N11675);
not NOT1 (N15198, N15166);
buf BUF1 (N15199, N15169);
buf BUF1 (N15200, N15198);
buf BUF1 (N15201, N15199);
or OR2 (N15202, N15188, N14844);
nor NOR4 (N15203, N15194, N4134, N4690, N3453);
buf BUF1 (N15204, N15183);
not NOT1 (N15205, N15189);
nor NOR4 (N15206, N15204, N1083, N9775, N10951);
and AND4 (N15207, N15190, N9208, N8872, N3452);
or OR3 (N15208, N15206, N4903, N2614);
and AND4 (N15209, N15208, N1841, N3718, N13520);
nor NOR4 (N15210, N15207, N5033, N12162, N12991);
not NOT1 (N15211, N15209);
not NOT1 (N15212, N15201);
or OR4 (N15213, N15211, N3874, N4058, N11763);
buf BUF1 (N15214, N15210);
buf BUF1 (N15215, N15205);
and AND2 (N15216, N15196, N274);
and AND2 (N15217, N15214, N4525);
nor NOR2 (N15218, N15213, N1133);
and AND2 (N15219, N15212, N14358);
or OR4 (N15220, N15182, N10518, N5623, N46);
and AND4 (N15221, N15215, N309, N9584, N14886);
or OR4 (N15222, N15221, N4141, N10312, N4647);
nand NAND4 (N15223, N15202, N3206, N982, N1211);
or OR3 (N15224, N15222, N1469, N48);
or OR3 (N15225, N15224, N14642, N5918);
or OR2 (N15226, N15203, N6718);
nor NOR4 (N15227, N15216, N4339, N9191, N8888);
or OR4 (N15228, N15220, N2244, N1123, N4300);
xor XOR2 (N15229, N15197, N1423);
not NOT1 (N15230, N15229);
not NOT1 (N15231, N15228);
and AND2 (N15232, N15230, N604);
and AND4 (N15233, N15217, N677, N7351, N12812);
nor NOR3 (N15234, N15226, N12224, N1714);
nand NAND4 (N15235, N15231, N11139, N8260, N9809);
nand NAND4 (N15236, N15219, N203, N9216, N3790);
nor NOR3 (N15237, N15227, N212, N493);
nor NOR4 (N15238, N15223, N1063, N3782, N14907);
xor XOR2 (N15239, N15232, N2855);
nand NAND4 (N15240, N15236, N6770, N12573, N12577);
xor XOR2 (N15241, N15240, N2888);
nor NOR4 (N15242, N15218, N1851, N7124, N3647);
not NOT1 (N15243, N15237);
buf BUF1 (N15244, N15238);
not NOT1 (N15245, N15200);
and AND3 (N15246, N15239, N12324, N11492);
xor XOR2 (N15247, N15244, N5029);
nand NAND3 (N15248, N15246, N2979, N4147);
xor XOR2 (N15249, N15225, N5582);
xor XOR2 (N15250, N15241, N1934);
nor NOR2 (N15251, N15247, N11455);
xor XOR2 (N15252, N15251, N15131);
buf BUF1 (N15253, N15235);
buf BUF1 (N15254, N15233);
not NOT1 (N15255, N15248);
xor XOR2 (N15256, N15250, N6379);
not NOT1 (N15257, N15245);
nand NAND3 (N15258, N15254, N3060, N14922);
nor NOR2 (N15259, N15242, N6746);
or OR3 (N15260, N15243, N69, N3318);
nand NAND4 (N15261, N15234, N11061, N2821, N2635);
nor NOR2 (N15262, N15257, N14853);
or OR2 (N15263, N15249, N11638);
buf BUF1 (N15264, N15255);
nor NOR4 (N15265, N15261, N10930, N154, N7231);
and AND4 (N15266, N15264, N8005, N1451, N3656);
buf BUF1 (N15267, N15252);
and AND4 (N15268, N15263, N1439, N9542, N14207);
or OR4 (N15269, N15259, N12453, N2067, N6451);
not NOT1 (N15270, N15260);
nand NAND4 (N15271, N15269, N11165, N14617, N7752);
nand NAND2 (N15272, N15258, N10235);
nand NAND4 (N15273, N15253, N5108, N4191, N4804);
or OR3 (N15274, N15271, N2339, N7032);
xor XOR2 (N15275, N15266, N12431);
xor XOR2 (N15276, N15274, N2171);
not NOT1 (N15277, N15273);
nor NOR2 (N15278, N15268, N10399);
nand NAND3 (N15279, N15275, N5398, N9043);
not NOT1 (N15280, N15277);
nand NAND3 (N15281, N15262, N1268, N11039);
or OR2 (N15282, N15276, N11904);
and AND2 (N15283, N15256, N4955);
buf BUF1 (N15284, N15281);
not NOT1 (N15285, N15280);
and AND2 (N15286, N15265, N10056);
or OR2 (N15287, N15284, N12038);
nor NOR4 (N15288, N15287, N4516, N10238, N12556);
buf BUF1 (N15289, N15272);
xor XOR2 (N15290, N15283, N8230);
buf BUF1 (N15291, N15286);
xor XOR2 (N15292, N15290, N8245);
buf BUF1 (N15293, N15288);
not NOT1 (N15294, N15293);
and AND4 (N15295, N15289, N1234, N6763, N2245);
xor XOR2 (N15296, N15278, N9465);
nand NAND4 (N15297, N15270, N3529, N10228, N9304);
or OR2 (N15298, N15279, N12012);
nor NOR2 (N15299, N15267, N14291);
not NOT1 (N15300, N15296);
or OR4 (N15301, N15291, N9902, N9392, N12086);
or OR2 (N15302, N15301, N7332);
nand NAND4 (N15303, N15302, N2451, N4736, N12247);
xor XOR2 (N15304, N15292, N9435);
buf BUF1 (N15305, N15282);
or OR3 (N15306, N15297, N10039, N2705);
and AND2 (N15307, N15295, N14016);
and AND4 (N15308, N15298, N3520, N8070, N14837);
nand NAND3 (N15309, N15294, N6981, N1654);
and AND3 (N15310, N15304, N15214, N1870);
nor NOR3 (N15311, N15305, N12848, N10222);
nand NAND4 (N15312, N15303, N10167, N6524, N7230);
nand NAND2 (N15313, N15309, N6839);
nor NOR4 (N15314, N15310, N4865, N418, N11856);
buf BUF1 (N15315, N15314);
xor XOR2 (N15316, N15312, N12026);
and AND3 (N15317, N15308, N10321, N13203);
nor NOR2 (N15318, N15306, N6695);
not NOT1 (N15319, N15285);
xor XOR2 (N15320, N15318, N5624);
and AND3 (N15321, N15316, N5705, N13797);
and AND4 (N15322, N15315, N7035, N12309, N2761);
nand NAND4 (N15323, N15317, N8292, N14259, N5064);
or OR4 (N15324, N15323, N3397, N10638, N690);
xor XOR2 (N15325, N15300, N681);
buf BUF1 (N15326, N15307);
nor NOR4 (N15327, N15326, N14506, N14770, N10278);
and AND4 (N15328, N15320, N8701, N5412, N5304);
or OR4 (N15329, N15322, N10233, N7711, N4977);
buf BUF1 (N15330, N15327);
or OR2 (N15331, N15311, N5617);
nand NAND2 (N15332, N15321, N2094);
nand NAND4 (N15333, N15299, N256, N11504, N10059);
and AND2 (N15334, N15333, N10572);
or OR2 (N15335, N15328, N9711);
nand NAND4 (N15336, N15329, N5035, N13400, N9420);
buf BUF1 (N15337, N15324);
and AND4 (N15338, N15313, N5952, N2259, N2231);
and AND3 (N15339, N15336, N14425, N11760);
or OR3 (N15340, N15334, N13788, N6149);
nand NAND4 (N15341, N15325, N6073, N1257, N5127);
nor NOR3 (N15342, N15337, N2815, N9989);
not NOT1 (N15343, N15339);
not NOT1 (N15344, N15342);
and AND3 (N15345, N15319, N12783, N14889);
or OR3 (N15346, N15332, N1278, N9894);
or OR4 (N15347, N15343, N14229, N8191, N12120);
nand NAND3 (N15348, N15338, N10051, N679);
not NOT1 (N15349, N15348);
nor NOR4 (N15350, N15346, N13668, N9033, N14029);
not NOT1 (N15351, N15341);
nor NOR4 (N15352, N15335, N12884, N3241, N4933);
or OR2 (N15353, N15352, N7501);
nand NAND4 (N15354, N15347, N6904, N6440, N14101);
buf BUF1 (N15355, N15349);
buf BUF1 (N15356, N15355);
not NOT1 (N15357, N15331);
xor XOR2 (N15358, N15330, N10415);
nor NOR3 (N15359, N15356, N11514, N1572);
not NOT1 (N15360, N15351);
and AND3 (N15361, N15359, N5330, N14961);
xor XOR2 (N15362, N15358, N1456);
and AND4 (N15363, N15344, N2930, N11079, N14311);
nor NOR2 (N15364, N15353, N1851);
or OR3 (N15365, N15357, N7032, N12287);
nand NAND3 (N15366, N15345, N10428, N14597);
or OR4 (N15367, N15361, N12814, N10380, N1404);
xor XOR2 (N15368, N15360, N3107);
not NOT1 (N15369, N15340);
and AND3 (N15370, N15362, N14959, N1317);
or OR4 (N15371, N15350, N8073, N8775, N8194);
not NOT1 (N15372, N15363);
nand NAND4 (N15373, N15368, N14666, N9680, N11251);
not NOT1 (N15374, N15369);
or OR2 (N15375, N15373, N10799);
nor NOR3 (N15376, N15366, N5007, N9637);
buf BUF1 (N15377, N15371);
buf BUF1 (N15378, N15376);
buf BUF1 (N15379, N15374);
nor NOR3 (N15380, N15370, N12674, N10397);
not NOT1 (N15381, N15354);
or OR2 (N15382, N15372, N14773);
xor XOR2 (N15383, N15367, N13712);
nor NOR3 (N15384, N15381, N6856, N11106);
nand NAND3 (N15385, N15364, N7751, N9542);
or OR3 (N15386, N15375, N6037, N3354);
or OR4 (N15387, N15380, N8422, N3140, N9049);
or OR3 (N15388, N15384, N3014, N13776);
or OR2 (N15389, N15387, N4104);
xor XOR2 (N15390, N15383, N1150);
buf BUF1 (N15391, N15390);
nand NAND3 (N15392, N15385, N15382, N5553);
buf BUF1 (N15393, N8397);
and AND4 (N15394, N15365, N15106, N9631, N4686);
not NOT1 (N15395, N15393);
xor XOR2 (N15396, N15389, N13129);
and AND4 (N15397, N15377, N5918, N12177, N7791);
or OR3 (N15398, N15386, N1257, N11837);
not NOT1 (N15399, N15391);
buf BUF1 (N15400, N15378);
or OR3 (N15401, N15388, N5397, N14717);
nor NOR4 (N15402, N15399, N6566, N14614, N1841);
nor NOR3 (N15403, N15401, N6157, N6920);
buf BUF1 (N15404, N15379);
buf BUF1 (N15405, N15398);
not NOT1 (N15406, N15392);
nor NOR3 (N15407, N15402, N5480, N202);
and AND2 (N15408, N15397, N12558);
xor XOR2 (N15409, N15406, N5226);
or OR2 (N15410, N15409, N10365);
or OR2 (N15411, N15407, N774);
xor XOR2 (N15412, N15411, N8198);
xor XOR2 (N15413, N15400, N7342);
or OR4 (N15414, N15405, N8919, N12373, N11884);
buf BUF1 (N15415, N15396);
nor NOR4 (N15416, N15394, N3959, N11447, N11783);
or OR2 (N15417, N15412, N14280);
not NOT1 (N15418, N15413);
buf BUF1 (N15419, N15410);
not NOT1 (N15420, N15416);
buf BUF1 (N15421, N15395);
xor XOR2 (N15422, N15414, N13632);
nor NOR3 (N15423, N15404, N10834, N187);
and AND3 (N15424, N15418, N4534, N9697);
nand NAND3 (N15425, N15419, N7025, N2524);
nand NAND3 (N15426, N15420, N6914, N10533);
xor XOR2 (N15427, N15417, N3585);
nor NOR3 (N15428, N15415, N12759, N13519);
not NOT1 (N15429, N15421);
or OR3 (N15430, N15425, N6920, N15252);
or OR3 (N15431, N15428, N2814, N5434);
buf BUF1 (N15432, N15431);
nor NOR2 (N15433, N15427, N9558);
and AND2 (N15434, N15424, N4605);
xor XOR2 (N15435, N15430, N5605);
or OR4 (N15436, N15435, N13689, N4957, N3543);
and AND4 (N15437, N15423, N10176, N6945, N1423);
and AND4 (N15438, N15434, N6974, N4690, N86);
nor NOR2 (N15439, N15433, N3364);
xor XOR2 (N15440, N15439, N3810);
not NOT1 (N15441, N15440);
nor NOR2 (N15442, N15422, N3336);
nor NOR2 (N15443, N15437, N1557);
nor NOR4 (N15444, N15408, N10914, N11743, N14590);
or OR4 (N15445, N15442, N6528, N5956, N7077);
xor XOR2 (N15446, N15436, N4596);
or OR4 (N15447, N15426, N12892, N5541, N7410);
and AND4 (N15448, N15446, N9564, N3879, N2724);
buf BUF1 (N15449, N15441);
not NOT1 (N15450, N15443);
xor XOR2 (N15451, N15448, N720);
or OR4 (N15452, N15403, N7600, N5378, N7135);
not NOT1 (N15453, N15451);
or OR2 (N15454, N15444, N8772);
xor XOR2 (N15455, N15429, N13494);
not NOT1 (N15456, N15453);
or OR3 (N15457, N15450, N2841, N1402);
and AND2 (N15458, N15449, N12174);
or OR2 (N15459, N15457, N9044);
buf BUF1 (N15460, N15456);
and AND3 (N15461, N15438, N11436, N9422);
xor XOR2 (N15462, N15458, N867);
or OR4 (N15463, N15462, N583, N9662, N1834);
nor NOR4 (N15464, N15459, N9729, N1619, N2454);
buf BUF1 (N15465, N15464);
and AND4 (N15466, N15461, N15245, N5431, N2587);
and AND4 (N15467, N15452, N2389, N7841, N9310);
nand NAND2 (N15468, N15455, N1314);
or OR4 (N15469, N15447, N12365, N1941, N1205);
not NOT1 (N15470, N15432);
nand NAND4 (N15471, N15460, N857, N506, N10407);
nor NOR4 (N15472, N15470, N3578, N3905, N10927);
xor XOR2 (N15473, N15454, N3632);
or OR4 (N15474, N15466, N2084, N8646, N4296);
not NOT1 (N15475, N15469);
nand NAND3 (N15476, N15474, N13374, N7551);
buf BUF1 (N15477, N15475);
not NOT1 (N15478, N15477);
xor XOR2 (N15479, N15473, N2331);
not NOT1 (N15480, N15463);
or OR2 (N15481, N15467, N11617);
or OR4 (N15482, N15476, N542, N13526, N7828);
nand NAND3 (N15483, N15468, N1243, N691);
nor NOR3 (N15484, N15478, N2572, N5237);
xor XOR2 (N15485, N15445, N12003);
and AND4 (N15486, N15465, N11764, N9887, N179);
xor XOR2 (N15487, N15472, N13442);
nor NOR3 (N15488, N15485, N4105, N4126);
and AND2 (N15489, N15480, N2524);
nor NOR2 (N15490, N15483, N12682);
not NOT1 (N15491, N15488);
buf BUF1 (N15492, N15486);
or OR4 (N15493, N15487, N2384, N3562, N9596);
xor XOR2 (N15494, N15489, N9659);
or OR3 (N15495, N15484, N7833, N3181);
buf BUF1 (N15496, N15493);
or OR4 (N15497, N15479, N15330, N6456, N14075);
xor XOR2 (N15498, N15471, N12839);
not NOT1 (N15499, N15494);
buf BUF1 (N15500, N15490);
or OR4 (N15501, N15500, N5075, N7777, N9190);
xor XOR2 (N15502, N15495, N10996);
and AND3 (N15503, N15502, N11307, N6585);
buf BUF1 (N15504, N15482);
or OR2 (N15505, N15481, N8623);
nor NOR2 (N15506, N15497, N8572);
xor XOR2 (N15507, N15505, N9183);
xor XOR2 (N15508, N15492, N6916);
not NOT1 (N15509, N15508);
or OR4 (N15510, N15501, N723, N10272, N10957);
buf BUF1 (N15511, N15491);
xor XOR2 (N15512, N15507, N12127);
xor XOR2 (N15513, N15510, N13063);
nand NAND2 (N15514, N15509, N6408);
or OR3 (N15515, N15504, N8217, N3751);
xor XOR2 (N15516, N15515, N4801);
not NOT1 (N15517, N15511);
or OR3 (N15518, N15503, N13003, N15072);
buf BUF1 (N15519, N15513);
and AND2 (N15520, N15498, N3470);
xor XOR2 (N15521, N15520, N15036);
nor NOR4 (N15522, N15512, N7391, N14927, N12931);
nor NOR3 (N15523, N15506, N11540, N1000);
nor NOR4 (N15524, N15523, N14615, N7169, N310);
nor NOR4 (N15525, N15514, N4343, N13238, N12779);
nand NAND4 (N15526, N15519, N9059, N8765, N9041);
and AND2 (N15527, N15524, N151);
buf BUF1 (N15528, N15526);
or OR3 (N15529, N15499, N6180, N2037);
nor NOR3 (N15530, N15496, N4781, N3015);
nand NAND3 (N15531, N15522, N1327, N14932);
and AND2 (N15532, N15518, N1646);
or OR3 (N15533, N15521, N10450, N14512);
or OR2 (N15534, N15528, N1564);
not NOT1 (N15535, N15532);
and AND3 (N15536, N15529, N9533, N10287);
buf BUF1 (N15537, N15531);
xor XOR2 (N15538, N15535, N3766);
or OR2 (N15539, N15533, N8361);
nand NAND2 (N15540, N15527, N12226);
not NOT1 (N15541, N15537);
xor XOR2 (N15542, N15538, N9292);
nand NAND2 (N15543, N15540, N7635);
not NOT1 (N15544, N15541);
nand NAND4 (N15545, N15534, N8990, N7238, N119);
or OR3 (N15546, N15517, N4453, N14896);
or OR2 (N15547, N15516, N4225);
not NOT1 (N15548, N15539);
nor NOR4 (N15549, N15543, N10550, N7246, N10926);
buf BUF1 (N15550, N15548);
xor XOR2 (N15551, N15549, N11363);
not NOT1 (N15552, N15546);
buf BUF1 (N15553, N15552);
nor NOR2 (N15554, N15544, N11918);
buf BUF1 (N15555, N15536);
nor NOR3 (N15556, N15545, N724, N961);
xor XOR2 (N15557, N15556, N7332);
nand NAND2 (N15558, N15551, N11776);
not NOT1 (N15559, N15525);
and AND4 (N15560, N15550, N3690, N10362, N7769);
buf BUF1 (N15561, N15560);
buf BUF1 (N15562, N15542);
not NOT1 (N15563, N15554);
and AND4 (N15564, N15555, N7586, N9999, N10320);
xor XOR2 (N15565, N15530, N9148);
nand NAND4 (N15566, N15547, N6888, N14704, N7017);
xor XOR2 (N15567, N15559, N14504);
nand NAND2 (N15568, N15558, N1622);
or OR4 (N15569, N15566, N11698, N12164, N4171);
buf BUF1 (N15570, N15569);
not NOT1 (N15571, N15561);
buf BUF1 (N15572, N15571);
nand NAND4 (N15573, N15567, N4907, N9680, N2911);
nand NAND3 (N15574, N15562, N70, N10140);
nor NOR3 (N15575, N15557, N9628, N12360);
buf BUF1 (N15576, N15574);
not NOT1 (N15577, N15572);
not NOT1 (N15578, N15564);
and AND4 (N15579, N15563, N15185, N7443, N359);
and AND4 (N15580, N15575, N337, N13030, N616);
xor XOR2 (N15581, N15577, N5559);
not NOT1 (N15582, N15573);
buf BUF1 (N15583, N15582);
xor XOR2 (N15584, N15570, N11752);
buf BUF1 (N15585, N15584);
buf BUF1 (N15586, N15580);
nand NAND4 (N15587, N15585, N13669, N14747, N555);
or OR2 (N15588, N15568, N8427);
or OR3 (N15589, N15553, N786, N5534);
buf BUF1 (N15590, N15581);
or OR3 (N15591, N15565, N4897, N3659);
buf BUF1 (N15592, N15576);
or OR2 (N15593, N15586, N1988);
not NOT1 (N15594, N15583);
xor XOR2 (N15595, N15587, N2570);
nand NAND4 (N15596, N15589, N8679, N1673, N12881);
xor XOR2 (N15597, N15596, N14094);
or OR3 (N15598, N15588, N1967, N2260);
xor XOR2 (N15599, N15592, N8278);
not NOT1 (N15600, N15597);
nand NAND3 (N15601, N15600, N2786, N3067);
nor NOR2 (N15602, N15593, N13472);
nand NAND4 (N15603, N15591, N5361, N11662, N3532);
or OR2 (N15604, N15599, N14108);
buf BUF1 (N15605, N15594);
or OR4 (N15606, N15598, N6882, N4266, N9867);
nand NAND4 (N15607, N15606, N5859, N11637, N8923);
not NOT1 (N15608, N15603);
nand NAND4 (N15609, N15608, N10344, N6941, N13392);
not NOT1 (N15610, N15578);
and AND4 (N15611, N15579, N12551, N2947, N15052);
xor XOR2 (N15612, N15607, N14523);
not NOT1 (N15613, N15590);
and AND3 (N15614, N15595, N7384, N2650);
xor XOR2 (N15615, N15605, N5008);
and AND3 (N15616, N15612, N1441, N8011);
xor XOR2 (N15617, N15610, N6302);
nor NOR4 (N15618, N15601, N3379, N5414, N5338);
and AND3 (N15619, N15609, N12230, N1048);
nor NOR3 (N15620, N15602, N10393, N12497);
nand NAND2 (N15621, N15614, N5150);
nor NOR2 (N15622, N15613, N1742);
not NOT1 (N15623, N15620);
not NOT1 (N15624, N15611);
and AND4 (N15625, N15617, N15104, N9648, N15162);
xor XOR2 (N15626, N15621, N486);
or OR3 (N15627, N15616, N5961, N11186);
nor NOR3 (N15628, N15604, N2387, N8799);
or OR3 (N15629, N15625, N806, N7019);
nand NAND2 (N15630, N15624, N14585);
buf BUF1 (N15631, N15618);
buf BUF1 (N15632, N15627);
buf BUF1 (N15633, N15619);
xor XOR2 (N15634, N15633, N13231);
or OR4 (N15635, N15634, N4581, N7487, N8128);
and AND4 (N15636, N15635, N12832, N14611, N11508);
nand NAND2 (N15637, N15628, N13688);
nor NOR4 (N15638, N15615, N2270, N15563, N12924);
nor NOR2 (N15639, N15631, N14576);
and AND3 (N15640, N15638, N6362, N4814);
xor XOR2 (N15641, N15637, N7807);
not NOT1 (N15642, N15641);
nand NAND2 (N15643, N15639, N927);
not NOT1 (N15644, N15626);
not NOT1 (N15645, N15630);
buf BUF1 (N15646, N15644);
nand NAND2 (N15647, N15646, N2424);
buf BUF1 (N15648, N15645);
nor NOR4 (N15649, N15647, N5838, N5052, N780);
nor NOR4 (N15650, N15642, N2550, N8967, N10453);
xor XOR2 (N15651, N15632, N861);
buf BUF1 (N15652, N15629);
buf BUF1 (N15653, N15643);
not NOT1 (N15654, N15636);
xor XOR2 (N15655, N15650, N5169);
or OR4 (N15656, N15651, N1471, N6650, N8236);
not NOT1 (N15657, N15623);
buf BUF1 (N15658, N15652);
buf BUF1 (N15659, N15648);
not NOT1 (N15660, N15649);
or OR4 (N15661, N15657, N8224, N14959, N9161);
buf BUF1 (N15662, N15660);
buf BUF1 (N15663, N15656);
and AND2 (N15664, N15659, N13731);
and AND4 (N15665, N15653, N454, N255, N7205);
xor XOR2 (N15666, N15655, N12510);
buf BUF1 (N15667, N15662);
or OR3 (N15668, N15640, N9655, N3055);
nand NAND2 (N15669, N15666, N2081);
nand NAND2 (N15670, N15661, N953);
xor XOR2 (N15671, N15668, N120);
nand NAND2 (N15672, N15658, N9889);
xor XOR2 (N15673, N15622, N8924);
or OR2 (N15674, N15667, N7736);
or OR3 (N15675, N15669, N5208, N1272);
or OR4 (N15676, N15674, N13915, N4563, N7755);
or OR3 (N15677, N15672, N1475, N15207);
or OR3 (N15678, N15654, N3511, N9563);
nor NOR2 (N15679, N15678, N5534);
and AND3 (N15680, N15665, N1019, N2395);
xor XOR2 (N15681, N15664, N7398);
not NOT1 (N15682, N15681);
not NOT1 (N15683, N15671);
xor XOR2 (N15684, N15675, N3396);
nand NAND4 (N15685, N15663, N4202, N14734, N3045);
nor NOR2 (N15686, N15683, N1869);
buf BUF1 (N15687, N15670);
nor NOR2 (N15688, N15679, N5589);
buf BUF1 (N15689, N15688);
not NOT1 (N15690, N15689);
not NOT1 (N15691, N15687);
xor XOR2 (N15692, N15691, N991);
and AND4 (N15693, N15682, N7714, N12080, N13505);
not NOT1 (N15694, N15673);
xor XOR2 (N15695, N15676, N4484);
nand NAND3 (N15696, N15677, N10719, N4941);
or OR4 (N15697, N15685, N2172, N7681, N5641);
xor XOR2 (N15698, N15697, N3247);
buf BUF1 (N15699, N15680);
buf BUF1 (N15700, N15686);
and AND3 (N15701, N15692, N7578, N11591);
or OR3 (N15702, N15684, N8820, N8334);
and AND4 (N15703, N15702, N1624, N14035, N7509);
buf BUF1 (N15704, N15696);
and AND4 (N15705, N15694, N6870, N10585, N4943);
nor NOR2 (N15706, N15703, N4134);
and AND2 (N15707, N15698, N14300);
nor NOR3 (N15708, N15695, N1189, N199);
nand NAND4 (N15709, N15693, N12988, N7228, N13507);
xor XOR2 (N15710, N15690, N2572);
or OR4 (N15711, N15706, N4029, N320, N8081);
buf BUF1 (N15712, N15709);
nor NOR2 (N15713, N15708, N15318);
nor NOR2 (N15714, N15704, N11887);
or OR3 (N15715, N15705, N7905, N9868);
and AND2 (N15716, N15715, N6556);
buf BUF1 (N15717, N15707);
buf BUF1 (N15718, N15713);
buf BUF1 (N15719, N15716);
not NOT1 (N15720, N15712);
xor XOR2 (N15721, N15717, N10294);
not NOT1 (N15722, N15714);
and AND2 (N15723, N15720, N8678);
or OR2 (N15724, N15700, N9566);
and AND2 (N15725, N15723, N8694);
nor NOR3 (N15726, N15699, N12093, N8651);
xor XOR2 (N15727, N15726, N14038);
and AND3 (N15728, N15711, N7110, N13945);
nor NOR3 (N15729, N15719, N13417, N151);
xor XOR2 (N15730, N15722, N8777);
and AND4 (N15731, N15729, N149, N5433, N12677);
nand NAND3 (N15732, N15710, N917, N3227);
and AND2 (N15733, N15727, N10538);
xor XOR2 (N15734, N15733, N15512);
nand NAND2 (N15735, N15731, N11526);
or OR4 (N15736, N15701, N6900, N4130, N7937);
and AND2 (N15737, N15732, N10701);
or OR3 (N15738, N15725, N10605, N1989);
not NOT1 (N15739, N15730);
xor XOR2 (N15740, N15728, N13304);
and AND3 (N15741, N15724, N9933, N10918);
buf BUF1 (N15742, N15739);
and AND2 (N15743, N15737, N7338);
or OR3 (N15744, N15738, N5631, N4428);
and AND4 (N15745, N15734, N14001, N2149, N6401);
xor XOR2 (N15746, N15744, N5322);
buf BUF1 (N15747, N15736);
buf BUF1 (N15748, N15745);
not NOT1 (N15749, N15747);
nand NAND2 (N15750, N15743, N15586);
nand NAND2 (N15751, N15740, N13478);
not NOT1 (N15752, N15721);
buf BUF1 (N15753, N15751);
and AND2 (N15754, N15746, N11990);
nor NOR2 (N15755, N15735, N792);
and AND4 (N15756, N15752, N2927, N3252, N12058);
xor XOR2 (N15757, N15748, N14636);
nand NAND3 (N15758, N15741, N12134, N1870);
xor XOR2 (N15759, N15749, N2214);
nand NAND2 (N15760, N15718, N12849);
and AND2 (N15761, N15742, N12998);
and AND2 (N15762, N15754, N269);
nand NAND3 (N15763, N15762, N10028, N1536);
or OR3 (N15764, N15763, N5321, N4143);
xor XOR2 (N15765, N15760, N2091);
not NOT1 (N15766, N15765);
nor NOR4 (N15767, N15755, N12915, N440, N13806);
and AND3 (N15768, N15758, N830, N12594);
buf BUF1 (N15769, N15753);
xor XOR2 (N15770, N15764, N1524);
nand NAND4 (N15771, N15768, N610, N2872, N15692);
nand NAND3 (N15772, N15769, N11912, N7887);
not NOT1 (N15773, N15767);
or OR4 (N15774, N15766, N11871, N3545, N2924);
and AND3 (N15775, N15750, N9766, N2508);
or OR4 (N15776, N15774, N4467, N1567, N1030);
or OR2 (N15777, N15759, N6756);
and AND4 (N15778, N15770, N1709, N3638, N13405);
buf BUF1 (N15779, N15757);
xor XOR2 (N15780, N15775, N289);
or OR3 (N15781, N15780, N6544, N1933);
or OR4 (N15782, N15772, N8822, N8663, N6711);
xor XOR2 (N15783, N15782, N12360);
not NOT1 (N15784, N15778);
not NOT1 (N15785, N15784);
nand NAND2 (N15786, N15779, N14585);
buf BUF1 (N15787, N15786);
nand NAND4 (N15788, N15776, N6734, N5068, N3142);
nor NOR4 (N15789, N15777, N10505, N9037, N5742);
buf BUF1 (N15790, N15781);
or OR3 (N15791, N15756, N10724, N5890);
nand NAND2 (N15792, N15789, N8804);
xor XOR2 (N15793, N15790, N10662);
nor NOR4 (N15794, N15783, N13626, N8276, N5766);
nor NOR4 (N15795, N15785, N5457, N10394, N12409);
xor XOR2 (N15796, N15771, N15667);
or OR2 (N15797, N15791, N5245);
nor NOR4 (N15798, N15793, N2994, N6466, N8838);
nor NOR3 (N15799, N15797, N15156, N2829);
xor XOR2 (N15800, N15792, N14803);
not NOT1 (N15801, N15800);
xor XOR2 (N15802, N15773, N15706);
not NOT1 (N15803, N15761);
nand NAND3 (N15804, N15802, N9463, N2346);
nor NOR3 (N15805, N15787, N5982, N13079);
nand NAND3 (N15806, N15794, N15433, N9787);
xor XOR2 (N15807, N15801, N6665);
and AND4 (N15808, N15807, N6348, N451, N13247);
xor XOR2 (N15809, N15799, N12489);
or OR3 (N15810, N15806, N11531, N11093);
or OR3 (N15811, N15804, N14137, N3137);
or OR3 (N15812, N15810, N1812, N15199);
nand NAND4 (N15813, N15805, N644, N6611, N11218);
xor XOR2 (N15814, N15788, N2843);
nor NOR4 (N15815, N15803, N8494, N11614, N2469);
and AND3 (N15816, N15808, N9437, N2357);
buf BUF1 (N15817, N15813);
buf BUF1 (N15818, N15817);
buf BUF1 (N15819, N15812);
nor NOR3 (N15820, N15818, N15705, N1630);
buf BUF1 (N15821, N15819);
or OR4 (N15822, N15796, N7487, N12433, N4981);
nor NOR2 (N15823, N15795, N307);
and AND3 (N15824, N15811, N12443, N8629);
nand NAND4 (N15825, N15823, N4264, N13935, N9419);
nor NOR3 (N15826, N15816, N3584, N11976);
not NOT1 (N15827, N15825);
or OR4 (N15828, N15814, N4104, N2068, N8973);
and AND2 (N15829, N15815, N11510);
nor NOR4 (N15830, N15826, N11936, N4943, N5483);
and AND4 (N15831, N15830, N9041, N4473, N14906);
and AND2 (N15832, N15822, N2426);
and AND3 (N15833, N15821, N15201, N5353);
nand NAND2 (N15834, N15798, N9955);
nand NAND2 (N15835, N15809, N12320);
not NOT1 (N15836, N15835);
nand NAND2 (N15837, N15824, N12197);
nand NAND3 (N15838, N15836, N13913, N3950);
or OR2 (N15839, N15838, N4924);
or OR2 (N15840, N15837, N7341);
or OR2 (N15841, N15831, N3381);
nor NOR4 (N15842, N15839, N8691, N13494, N15499);
or OR4 (N15843, N15828, N7694, N13402, N5703);
nand NAND2 (N15844, N15820, N5471);
and AND3 (N15845, N15843, N3733, N13576);
nor NOR4 (N15846, N15841, N11458, N14228, N1687);
or OR4 (N15847, N15834, N8607, N11273, N15456);
and AND3 (N15848, N15840, N8320, N653);
nor NOR3 (N15849, N15833, N15295, N4914);
buf BUF1 (N15850, N15827);
nand NAND4 (N15851, N15844, N2601, N592, N11343);
or OR3 (N15852, N15850, N8804, N9343);
nor NOR2 (N15853, N15832, N6811);
xor XOR2 (N15854, N15847, N11955);
or OR2 (N15855, N15829, N9315);
xor XOR2 (N15856, N15848, N10789);
nor NOR2 (N15857, N15852, N4777);
not NOT1 (N15858, N15856);
and AND4 (N15859, N15849, N9627, N7398, N12410);
nor NOR4 (N15860, N15858, N3181, N3756, N11552);
not NOT1 (N15861, N15853);
buf BUF1 (N15862, N15851);
or OR3 (N15863, N15862, N950, N1803);
xor XOR2 (N15864, N15855, N9863);
not NOT1 (N15865, N15859);
nand NAND2 (N15866, N15863, N2278);
nor NOR3 (N15867, N15846, N8412, N11970);
nor NOR3 (N15868, N15842, N3239, N15063);
and AND3 (N15869, N15845, N13176, N8204);
nor NOR2 (N15870, N15861, N301);
and AND2 (N15871, N15868, N2632);
and AND3 (N15872, N15860, N963, N5486);
or OR4 (N15873, N15871, N12432, N4398, N9444);
or OR2 (N15874, N15866, N4222);
not NOT1 (N15875, N15870);
and AND2 (N15876, N15874, N7963);
or OR3 (N15877, N15875, N2628, N1898);
and AND2 (N15878, N15854, N1351);
nor NOR2 (N15879, N15872, N212);
and AND4 (N15880, N15864, N445, N11236, N3225);
or OR4 (N15881, N15878, N8204, N5623, N3172);
xor XOR2 (N15882, N15881, N7034);
not NOT1 (N15883, N15877);
xor XOR2 (N15884, N15883, N12999);
xor XOR2 (N15885, N15869, N3762);
nor NOR2 (N15886, N15873, N2712);
xor XOR2 (N15887, N15867, N1652);
nor NOR4 (N15888, N15884, N10612, N6203, N4756);
nor NOR3 (N15889, N15879, N1436, N12298);
nand NAND4 (N15890, N15857, N9680, N3035, N7568);
nor NOR4 (N15891, N15887, N699, N1533, N10411);
or OR3 (N15892, N15888, N13192, N8372);
or OR4 (N15893, N15892, N6279, N2860, N14878);
or OR2 (N15894, N15882, N4817);
buf BUF1 (N15895, N15889);
nand NAND3 (N15896, N15865, N4044, N9049);
nand NAND2 (N15897, N15886, N2512);
nand NAND4 (N15898, N15894, N3122, N12514, N15530);
buf BUF1 (N15899, N15876);
nand NAND4 (N15900, N15890, N7121, N13237, N5004);
and AND3 (N15901, N15898, N3539, N15321);
not NOT1 (N15902, N15896);
nand NAND4 (N15903, N15902, N15551, N8687, N7610);
or OR2 (N15904, N15897, N1697);
and AND3 (N15905, N15891, N14138, N15846);
nor NOR3 (N15906, N15903, N14516, N10558);
nor NOR2 (N15907, N15880, N1411);
buf BUF1 (N15908, N15885);
nand NAND4 (N15909, N15906, N5095, N13272, N1041);
and AND3 (N15910, N15908, N13124, N14301);
xor XOR2 (N15911, N15901, N12694);
not NOT1 (N15912, N15895);
nor NOR2 (N15913, N15905, N11514);
and AND4 (N15914, N15899, N10520, N14139, N8085);
xor XOR2 (N15915, N15912, N5757);
nand NAND4 (N15916, N15910, N11870, N8172, N14254);
nand NAND3 (N15917, N15911, N8175, N15416);
nand NAND3 (N15918, N15909, N15505, N13610);
and AND4 (N15919, N15916, N5696, N9109, N4952);
nor NOR3 (N15920, N15917, N2014, N7213);
buf BUF1 (N15921, N15907);
xor XOR2 (N15922, N15900, N10096);
nand NAND3 (N15923, N15919, N2387, N7292);
buf BUF1 (N15924, N15913);
nor NOR4 (N15925, N15918, N13284, N24, N6683);
nand NAND4 (N15926, N15924, N4739, N10728, N14395);
buf BUF1 (N15927, N15920);
buf BUF1 (N15928, N15921);
buf BUF1 (N15929, N15928);
buf BUF1 (N15930, N15923);
xor XOR2 (N15931, N15893, N8658);
not NOT1 (N15932, N15929);
and AND3 (N15933, N15931, N1492, N4950);
nand NAND4 (N15934, N15930, N14096, N15252, N10203);
nand NAND4 (N15935, N15904, N5823, N955, N3439);
and AND2 (N15936, N15934, N3695);
buf BUF1 (N15937, N15933);
and AND4 (N15938, N15927, N8932, N15388, N12155);
xor XOR2 (N15939, N15937, N8598);
nand NAND3 (N15940, N15925, N1913, N2552);
buf BUF1 (N15941, N15915);
nor NOR4 (N15942, N15941, N2744, N9993, N5083);
not NOT1 (N15943, N15935);
and AND2 (N15944, N15932, N15419);
buf BUF1 (N15945, N15926);
xor XOR2 (N15946, N15922, N3457);
nor NOR2 (N15947, N15914, N5432);
and AND3 (N15948, N15936, N1152, N3166);
and AND4 (N15949, N15940, N9547, N14456, N15544);
buf BUF1 (N15950, N15949);
not NOT1 (N15951, N15939);
buf BUF1 (N15952, N15938);
xor XOR2 (N15953, N15948, N13622);
not NOT1 (N15954, N15944);
nor NOR3 (N15955, N15954, N12760, N9672);
or OR3 (N15956, N15947, N2910, N9595);
nor NOR4 (N15957, N15946, N9823, N12945, N13020);
xor XOR2 (N15958, N15950, N10531);
and AND2 (N15959, N15945, N2513);
or OR2 (N15960, N15943, N700);
buf BUF1 (N15961, N15952);
nand NAND2 (N15962, N15958, N8258);
nand NAND2 (N15963, N15959, N9298);
not NOT1 (N15964, N15953);
xor XOR2 (N15965, N15955, N2083);
xor XOR2 (N15966, N15963, N7832);
not NOT1 (N15967, N15956);
nand NAND3 (N15968, N15960, N1844, N5977);
xor XOR2 (N15969, N15961, N6195);
xor XOR2 (N15970, N15951, N3355);
and AND4 (N15971, N15957, N2798, N1231, N8385);
not NOT1 (N15972, N15962);
nand NAND4 (N15973, N15964, N812, N15888, N4220);
and AND2 (N15974, N15967, N5377);
buf BUF1 (N15975, N15972);
not NOT1 (N15976, N15974);
not NOT1 (N15977, N15968);
or OR2 (N15978, N15965, N15217);
not NOT1 (N15979, N15977);
and AND3 (N15980, N15979, N10401, N8496);
or OR4 (N15981, N15969, N6623, N14994, N2261);
nand NAND3 (N15982, N15975, N13116, N14353);
buf BUF1 (N15983, N15966);
and AND2 (N15984, N15976, N13715);
not NOT1 (N15985, N15984);
not NOT1 (N15986, N15942);
or OR3 (N15987, N15985, N12753, N1625);
or OR3 (N15988, N15983, N13733, N14013);
or OR4 (N15989, N15986, N10120, N5538, N13201);
not NOT1 (N15990, N15988);
xor XOR2 (N15991, N15989, N13634);
not NOT1 (N15992, N15978);
nor NOR4 (N15993, N15990, N11927, N13715, N14868);
not NOT1 (N15994, N15993);
buf BUF1 (N15995, N15973);
and AND2 (N15996, N15980, N12332);
xor XOR2 (N15997, N15996, N15951);
not NOT1 (N15998, N15982);
not NOT1 (N15999, N15994);
not NOT1 (N16000, N15981);
buf BUF1 (N16001, N16000);
nor NOR4 (N16002, N15998, N8181, N15182, N7485);
nand NAND3 (N16003, N16002, N273, N396);
buf BUF1 (N16004, N15992);
nor NOR4 (N16005, N15970, N10752, N7957, N2247);
not NOT1 (N16006, N15991);
and AND3 (N16007, N15995, N6867, N9980);
or OR4 (N16008, N16001, N11401, N1968, N6675);
not NOT1 (N16009, N16005);
or OR4 (N16010, N16006, N5819, N1851, N11224);
endmodule