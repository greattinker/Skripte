// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N2497,N2513,N2510,N2509,N2516,N2512,N2506,N2515,N2507,N2517;

xor XOR2 (N18, N4, N9);
xor XOR2 (N19, N2, N16);
not NOT1 (N20, N12);
not NOT1 (N21, N5);
or OR2 (N22, N12, N19);
and AND2 (N23, N1, N19);
and AND3 (N24, N14, N16, N10);
xor XOR2 (N25, N10, N18);
or OR4 (N26, N15, N24, N21, N5);
xor XOR2 (N27, N22, N9);
nor NOR3 (N28, N27, N13, N8);
not NOT1 (N29, N14);
xor XOR2 (N30, N18, N13);
not NOT1 (N31, N15);
buf BUF1 (N32, N3);
not NOT1 (N33, N9);
buf BUF1 (N34, N28);
and AND2 (N35, N29, N15);
and AND2 (N36, N31, N28);
nand NAND4 (N37, N26, N11, N21, N3);
not NOT1 (N38, N35);
or OR3 (N39, N25, N12, N37);
not NOT1 (N40, N13);
nand NAND3 (N41, N32, N7, N6);
nor NOR4 (N42, N41, N23, N20, N26);
nand NAND3 (N43, N9, N9, N42);
or OR4 (N44, N9, N7, N26, N39);
nor NOR2 (N45, N18, N41);
not NOT1 (N46, N5);
not NOT1 (N47, N33);
not NOT1 (N48, N40);
not NOT1 (N49, N30);
xor XOR2 (N50, N36, N22);
nor NOR4 (N51, N50, N3, N24, N6);
and AND4 (N52, N38, N37, N18, N46);
buf BUF1 (N53, N18);
nand NAND3 (N54, N45, N1, N31);
nand NAND2 (N55, N47, N16);
xor XOR2 (N56, N44, N38);
and AND2 (N57, N56, N13);
not NOT1 (N58, N53);
nand NAND4 (N59, N52, N54, N58, N47);
xor XOR2 (N60, N39, N23);
nand NAND3 (N61, N26, N55, N13);
or OR2 (N62, N48, N46);
and AND4 (N63, N15, N35, N45, N43);
not NOT1 (N64, N37);
not NOT1 (N65, N34);
xor XOR2 (N66, N49, N5);
not NOT1 (N67, N63);
xor XOR2 (N68, N61, N46);
nand NAND4 (N69, N60, N44, N9, N9);
not NOT1 (N70, N67);
or OR3 (N71, N70, N70, N32);
nand NAND2 (N72, N68, N36);
buf BUF1 (N73, N57);
buf BUF1 (N74, N65);
not NOT1 (N75, N72);
or OR2 (N76, N51, N32);
not NOT1 (N77, N75);
or OR3 (N78, N71, N49, N5);
buf BUF1 (N79, N62);
or OR2 (N80, N73, N3);
xor XOR2 (N81, N74, N78);
nand NAND2 (N82, N36, N17);
nand NAND4 (N83, N80, N8, N29, N62);
buf BUF1 (N84, N64);
nor NOR4 (N85, N83, N54, N18, N32);
not NOT1 (N86, N76);
or OR4 (N87, N79, N30, N45, N44);
or OR2 (N88, N82, N85);
nand NAND4 (N89, N40, N2, N18, N7);
or OR2 (N90, N89, N83);
nand NAND2 (N91, N90, N1);
buf BUF1 (N92, N87);
buf BUF1 (N93, N86);
nor NOR3 (N94, N84, N8, N61);
not NOT1 (N95, N93);
nand NAND2 (N96, N91, N86);
buf BUF1 (N97, N59);
buf BUF1 (N98, N66);
xor XOR2 (N99, N95, N74);
xor XOR2 (N100, N88, N93);
or OR4 (N101, N97, N36, N27, N68);
nor NOR2 (N102, N94, N57);
xor XOR2 (N103, N102, N75);
or OR4 (N104, N77, N66, N30, N73);
nand NAND3 (N105, N98, N79, N34);
or OR4 (N106, N100, N75, N45, N70);
xor XOR2 (N107, N103, N36);
or OR4 (N108, N104, N42, N52, N58);
xor XOR2 (N109, N108, N64);
and AND2 (N110, N69, N22);
not NOT1 (N111, N105);
and AND3 (N112, N111, N62, N46);
nand NAND2 (N113, N99, N52);
buf BUF1 (N114, N81);
and AND2 (N115, N106, N27);
nand NAND3 (N116, N115, N80, N29);
nand NAND3 (N117, N109, N62, N43);
not NOT1 (N118, N101);
and AND4 (N119, N117, N1, N50, N84);
nand NAND3 (N120, N92, N24, N39);
and AND2 (N121, N114, N117);
or OR4 (N122, N107, N103, N28, N1);
nand NAND4 (N123, N110, N55, N73, N117);
nor NOR4 (N124, N112, N73, N107, N96);
nor NOR3 (N125, N71, N96, N109);
not NOT1 (N126, N113);
nand NAND4 (N127, N118, N14, N115, N3);
nor NOR3 (N128, N126, N11, N56);
and AND3 (N129, N122, N58, N31);
nor NOR3 (N130, N129, N87, N18);
or OR3 (N131, N116, N67, N82);
xor XOR2 (N132, N119, N118);
xor XOR2 (N133, N120, N28);
or OR4 (N134, N124, N64, N93, N63);
or OR2 (N135, N132, N108);
buf BUF1 (N136, N133);
buf BUF1 (N137, N136);
not NOT1 (N138, N128);
xor XOR2 (N139, N123, N15);
nor NOR2 (N140, N130, N116);
buf BUF1 (N141, N137);
not NOT1 (N142, N131);
not NOT1 (N143, N121);
nor NOR3 (N144, N127, N106, N23);
or OR3 (N145, N143, N108, N89);
nor NOR4 (N146, N140, N120, N88, N117);
or OR2 (N147, N134, N130);
not NOT1 (N148, N144);
not NOT1 (N149, N145);
xor XOR2 (N150, N139, N127);
buf BUF1 (N151, N146);
nand NAND4 (N152, N138, N15, N135, N81);
and AND4 (N153, N130, N150, N103, N151);
or OR4 (N154, N47, N15, N130, N78);
xor XOR2 (N155, N140, N140);
xor XOR2 (N156, N142, N92);
or OR4 (N157, N141, N102, N117, N143);
not NOT1 (N158, N153);
nand NAND2 (N159, N125, N156);
not NOT1 (N160, N28);
xor XOR2 (N161, N158, N92);
not NOT1 (N162, N148);
xor XOR2 (N163, N147, N69);
nor NOR3 (N164, N154, N24, N157);
and AND3 (N165, N74, N70, N67);
nand NAND4 (N166, N165, N64, N135, N150);
nor NOR4 (N167, N149, N12, N79, N121);
not NOT1 (N168, N160);
buf BUF1 (N169, N168);
not NOT1 (N170, N152);
not NOT1 (N171, N164);
nor NOR2 (N172, N169, N162);
and AND3 (N173, N151, N39, N68);
xor XOR2 (N174, N155, N50);
nand NAND4 (N175, N173, N156, N128, N168);
nor NOR2 (N176, N171, N83);
nand NAND3 (N177, N175, N37, N56);
nand NAND2 (N178, N172, N53);
xor XOR2 (N179, N163, N132);
nor NOR3 (N180, N166, N66, N1);
xor XOR2 (N181, N167, N162);
nor NOR4 (N182, N179, N144, N52, N8);
xor XOR2 (N183, N170, N148);
xor XOR2 (N184, N183, N90);
xor XOR2 (N185, N181, N65);
and AND3 (N186, N185, N148, N78);
not NOT1 (N187, N182);
buf BUF1 (N188, N180);
buf BUF1 (N189, N187);
not NOT1 (N190, N188);
and AND4 (N191, N176, N126, N177, N97);
nor NOR3 (N192, N98, N26, N119);
nand NAND4 (N193, N174, N124, N40, N5);
nor NOR4 (N194, N159, N176, N97, N77);
nor NOR3 (N195, N192, N128, N158);
xor XOR2 (N196, N178, N100);
or OR2 (N197, N184, N19);
nor NOR4 (N198, N190, N130, N57, N68);
or OR4 (N199, N189, N192, N183, N42);
or OR4 (N200, N191, N192, N189, N69);
buf BUF1 (N201, N161);
xor XOR2 (N202, N200, N134);
or OR2 (N203, N197, N87);
and AND2 (N204, N198, N186);
or OR3 (N205, N95, N78, N91);
or OR2 (N206, N204, N21);
buf BUF1 (N207, N203);
not NOT1 (N208, N196);
or OR2 (N209, N193, N143);
or OR2 (N210, N205, N99);
and AND4 (N211, N194, N53, N194, N117);
not NOT1 (N212, N208);
nor NOR2 (N213, N211, N12);
not NOT1 (N214, N206);
nor NOR4 (N215, N214, N207, N16, N15);
not NOT1 (N216, N24);
and AND4 (N217, N201, N206, N90, N11);
not NOT1 (N218, N212);
not NOT1 (N219, N210);
or OR4 (N220, N202, N125, N155, N163);
not NOT1 (N221, N219);
or OR2 (N222, N218, N102);
buf BUF1 (N223, N209);
and AND3 (N224, N221, N164, N190);
nand NAND2 (N225, N223, N168);
nor NOR2 (N226, N225, N213);
nor NOR2 (N227, N1, N17);
nor NOR4 (N228, N220, N146, N93, N9);
xor XOR2 (N229, N217, N197);
xor XOR2 (N230, N224, N66);
xor XOR2 (N231, N229, N204);
nand NAND2 (N232, N222, N114);
nor NOR4 (N233, N216, N209, N191, N190);
nor NOR2 (N234, N233, N197);
or OR2 (N235, N226, N12);
nor NOR2 (N236, N232, N189);
or OR2 (N237, N199, N144);
or OR4 (N238, N234, N174, N148, N13);
and AND4 (N239, N231, N58, N24, N102);
nand NAND4 (N240, N235, N221, N136, N163);
or OR3 (N241, N237, N202, N134);
xor XOR2 (N242, N228, N7);
nor NOR2 (N243, N240, N108);
nand NAND3 (N244, N241, N32, N149);
and AND2 (N245, N215, N15);
not NOT1 (N246, N245);
buf BUF1 (N247, N227);
nand NAND3 (N248, N230, N152, N200);
buf BUF1 (N249, N239);
or OR3 (N250, N236, N45, N65);
nor NOR3 (N251, N247, N31, N203);
buf BUF1 (N252, N242);
xor XOR2 (N253, N250, N70);
nand NAND2 (N254, N243, N58);
nand NAND4 (N255, N246, N156, N211, N94);
nor NOR2 (N256, N255, N65);
nand NAND3 (N257, N254, N115, N253);
or OR3 (N258, N243, N187, N179);
nand NAND4 (N259, N256, N96, N36, N104);
nor NOR4 (N260, N257, N15, N34, N244);
and AND3 (N261, N26, N211, N226);
buf BUF1 (N262, N260);
buf BUF1 (N263, N249);
buf BUF1 (N264, N251);
and AND3 (N265, N248, N103, N245);
xor XOR2 (N266, N265, N35);
xor XOR2 (N267, N238, N251);
not NOT1 (N268, N252);
or OR4 (N269, N268, N121, N243, N173);
and AND2 (N270, N266, N203);
and AND4 (N271, N263, N62, N220, N143);
not NOT1 (N272, N259);
nor NOR3 (N273, N262, N115, N88);
buf BUF1 (N274, N264);
xor XOR2 (N275, N274, N101);
or OR4 (N276, N261, N163, N226, N70);
and AND4 (N277, N273, N93, N180, N72);
xor XOR2 (N278, N269, N88);
xor XOR2 (N279, N276, N41);
xor XOR2 (N280, N277, N122);
or OR2 (N281, N279, N161);
not NOT1 (N282, N270);
or OR2 (N283, N258, N149);
not NOT1 (N284, N280);
nand NAND4 (N285, N281, N60, N283, N249);
buf BUF1 (N286, N177);
not NOT1 (N287, N285);
or OR3 (N288, N267, N97, N195);
buf BUF1 (N289, N267);
not NOT1 (N290, N271);
buf BUF1 (N291, N278);
or OR3 (N292, N291, N247, N108);
nand NAND4 (N293, N272, N105, N99, N251);
nor NOR2 (N294, N286, N30);
buf BUF1 (N295, N282);
not NOT1 (N296, N295);
xor XOR2 (N297, N293, N254);
nand NAND2 (N298, N297, N88);
nand NAND3 (N299, N287, N225, N241);
nand NAND4 (N300, N296, N295, N169, N108);
nor NOR3 (N301, N292, N146, N232);
nor NOR2 (N302, N275, N127);
not NOT1 (N303, N288);
or OR4 (N304, N303, N262, N1, N11);
nor NOR4 (N305, N302, N205, N239, N106);
nand NAND2 (N306, N305, N8);
buf BUF1 (N307, N298);
xor XOR2 (N308, N307, N82);
nor NOR2 (N309, N294, N136);
and AND2 (N310, N306, N146);
or OR4 (N311, N299, N265, N129, N239);
not NOT1 (N312, N310);
nand NAND2 (N313, N289, N246);
and AND4 (N314, N301, N41, N235, N136);
or OR2 (N315, N308, N258);
xor XOR2 (N316, N304, N245);
not NOT1 (N317, N314);
xor XOR2 (N318, N313, N302);
and AND4 (N319, N317, N197, N274, N82);
nand NAND4 (N320, N309, N263, N271, N284);
nand NAND4 (N321, N15, N52, N76, N312);
or OR4 (N322, N22, N132, N128, N147);
or OR4 (N323, N290, N234, N194, N164);
buf BUF1 (N324, N300);
and AND3 (N325, N324, N93, N306);
xor XOR2 (N326, N319, N230);
xor XOR2 (N327, N311, N181);
buf BUF1 (N328, N320);
nor NOR3 (N329, N328, N215, N167);
buf BUF1 (N330, N315);
or OR2 (N331, N322, N106);
and AND2 (N332, N329, N216);
not NOT1 (N333, N316);
xor XOR2 (N334, N331, N315);
or OR3 (N335, N321, N308, N23);
or OR2 (N336, N335, N292);
nand NAND2 (N337, N326, N89);
or OR4 (N338, N325, N78, N274, N316);
buf BUF1 (N339, N323);
xor XOR2 (N340, N338, N96);
xor XOR2 (N341, N333, N93);
xor XOR2 (N342, N334, N3);
xor XOR2 (N343, N342, N140);
and AND3 (N344, N337, N142, N248);
xor XOR2 (N345, N340, N37);
xor XOR2 (N346, N341, N187);
nor NOR3 (N347, N327, N345, N198);
and AND3 (N348, N282, N344, N218);
or OR3 (N349, N195, N62, N229);
xor XOR2 (N350, N339, N160);
not NOT1 (N351, N350);
or OR3 (N352, N347, N268, N236);
nand NAND3 (N353, N348, N78, N271);
and AND3 (N354, N349, N353, N19);
or OR4 (N355, N78, N312, N39, N220);
buf BUF1 (N356, N330);
or OR2 (N357, N352, N115);
xor XOR2 (N358, N346, N281);
xor XOR2 (N359, N332, N89);
xor XOR2 (N360, N358, N282);
nand NAND4 (N361, N343, N108, N3, N280);
not NOT1 (N362, N318);
and AND4 (N363, N336, N60, N243, N79);
not NOT1 (N364, N351);
buf BUF1 (N365, N357);
buf BUF1 (N366, N356);
nor NOR4 (N367, N366, N283, N191, N129);
buf BUF1 (N368, N361);
nor NOR2 (N369, N359, N230);
not NOT1 (N370, N363);
and AND4 (N371, N369, N297, N200, N318);
nand NAND4 (N372, N367, N269, N289, N228);
nor NOR2 (N373, N370, N320);
nor NOR4 (N374, N365, N297, N305, N248);
nand NAND2 (N375, N373, N233);
xor XOR2 (N376, N375, N290);
nor NOR4 (N377, N360, N273, N344, N112);
buf BUF1 (N378, N362);
nor NOR4 (N379, N372, N316, N133, N7);
and AND3 (N380, N376, N180, N346);
nor NOR4 (N381, N354, N154, N228, N133);
not NOT1 (N382, N381);
nand NAND4 (N383, N382, N340, N99, N259);
xor XOR2 (N384, N378, N8);
buf BUF1 (N385, N374);
not NOT1 (N386, N355);
nor NOR4 (N387, N383, N272, N343, N311);
xor XOR2 (N388, N371, N278);
xor XOR2 (N389, N368, N372);
and AND3 (N390, N385, N175, N49);
and AND2 (N391, N388, N362);
buf BUF1 (N392, N391);
nor NOR2 (N393, N387, N101);
nand NAND4 (N394, N393, N346, N146, N195);
nand NAND3 (N395, N386, N24, N215);
buf BUF1 (N396, N395);
nand NAND4 (N397, N389, N49, N184, N106);
nor NOR3 (N398, N397, N147, N273);
xor XOR2 (N399, N377, N299);
and AND2 (N400, N390, N374);
and AND3 (N401, N384, N13, N233);
xor XOR2 (N402, N380, N277);
not NOT1 (N403, N394);
or OR2 (N404, N400, N243);
not NOT1 (N405, N379);
nor NOR4 (N406, N398, N181, N320, N17);
or OR2 (N407, N402, N117);
or OR4 (N408, N403, N355, N167, N353);
and AND4 (N409, N408, N126, N140, N294);
nand NAND3 (N410, N364, N406, N249);
or OR2 (N411, N186, N109);
nand NAND4 (N412, N405, N78, N118, N5);
nand NAND4 (N413, N396, N320, N351, N336);
nand NAND2 (N414, N409, N403);
buf BUF1 (N415, N407);
and AND2 (N416, N414, N235);
or OR3 (N417, N416, N279, N323);
nor NOR2 (N418, N401, N201);
xor XOR2 (N419, N410, N41);
and AND3 (N420, N418, N416, N44);
nor NOR3 (N421, N413, N351, N309);
nand NAND4 (N422, N412, N296, N259, N390);
and AND2 (N423, N419, N99);
or OR2 (N424, N415, N352);
not NOT1 (N425, N411);
buf BUF1 (N426, N417);
and AND3 (N427, N426, N86, N380);
and AND3 (N428, N399, N32, N179);
nand NAND4 (N429, N427, N319, N358, N110);
nor NOR3 (N430, N423, N28, N322);
xor XOR2 (N431, N392, N313);
and AND3 (N432, N431, N266, N114);
buf BUF1 (N433, N429);
xor XOR2 (N434, N422, N288);
nor NOR2 (N435, N421, N417);
not NOT1 (N436, N425);
and AND4 (N437, N436, N239, N405, N217);
nand NAND4 (N438, N432, N347, N260, N301);
nor NOR4 (N439, N434, N66, N351, N181);
nand NAND3 (N440, N430, N157, N234);
and AND3 (N441, N404, N81, N382);
nor NOR4 (N442, N420, N71, N218, N282);
nand NAND3 (N443, N439, N246, N307);
nand NAND3 (N444, N433, N205, N199);
or OR4 (N445, N440, N345, N116, N204);
nand NAND4 (N446, N442, N138, N417, N14);
and AND4 (N447, N424, N341, N72, N333);
and AND3 (N448, N444, N292, N118);
xor XOR2 (N449, N445, N178);
nand NAND2 (N450, N435, N137);
buf BUF1 (N451, N448);
xor XOR2 (N452, N437, N200);
and AND3 (N453, N450, N11, N135);
nor NOR2 (N454, N441, N315);
not NOT1 (N455, N447);
and AND2 (N456, N453, N55);
or OR2 (N457, N454, N308);
or OR4 (N458, N446, N433, N52, N50);
not NOT1 (N459, N455);
and AND2 (N460, N456, N226);
nor NOR4 (N461, N428, N236, N66, N144);
nand NAND3 (N462, N443, N126, N203);
or OR4 (N463, N449, N188, N180, N175);
buf BUF1 (N464, N462);
buf BUF1 (N465, N458);
nor NOR3 (N466, N452, N247, N344);
nor NOR3 (N467, N457, N307, N466);
not NOT1 (N468, N49);
or OR4 (N469, N467, N310, N253, N466);
xor XOR2 (N470, N469, N428);
xor XOR2 (N471, N459, N379);
xor XOR2 (N472, N463, N61);
not NOT1 (N473, N464);
not NOT1 (N474, N473);
not NOT1 (N475, N468);
and AND4 (N476, N471, N74, N425, N29);
and AND3 (N477, N451, N317, N259);
buf BUF1 (N478, N472);
and AND4 (N479, N460, N265, N369, N167);
buf BUF1 (N480, N478);
nand NAND3 (N481, N477, N197, N106);
or OR2 (N482, N476, N331);
buf BUF1 (N483, N482);
xor XOR2 (N484, N461, N43);
buf BUF1 (N485, N481);
not NOT1 (N486, N480);
buf BUF1 (N487, N485);
or OR4 (N488, N483, N337, N131, N306);
and AND4 (N489, N479, N174, N158, N289);
nand NAND3 (N490, N486, N240, N312);
xor XOR2 (N491, N490, N252);
buf BUF1 (N492, N491);
buf BUF1 (N493, N474);
or OR2 (N494, N489, N31);
and AND4 (N495, N488, N115, N306, N131);
buf BUF1 (N496, N494);
or OR4 (N497, N484, N468, N276, N261);
nor NOR3 (N498, N475, N37, N112);
buf BUF1 (N499, N492);
nand NAND4 (N500, N496, N356, N284, N266);
nand NAND3 (N501, N500, N120, N197);
nand NAND3 (N502, N438, N377, N468);
and AND4 (N503, N487, N163, N306, N107);
not NOT1 (N504, N499);
and AND4 (N505, N504, N412, N73, N339);
and AND4 (N506, N503, N201, N139, N435);
and AND4 (N507, N502, N354, N188, N145);
or OR4 (N508, N498, N229, N190, N248);
xor XOR2 (N509, N505, N119);
or OR2 (N510, N501, N18);
xor XOR2 (N511, N509, N77);
nand NAND4 (N512, N493, N84, N306, N109);
nand NAND2 (N513, N465, N99);
nand NAND4 (N514, N512, N437, N342, N46);
or OR2 (N515, N510, N360);
nand NAND3 (N516, N508, N166, N233);
xor XOR2 (N517, N470, N54);
nand NAND4 (N518, N515, N517, N407, N417);
and AND3 (N519, N278, N93, N129);
nor NOR3 (N520, N513, N250, N146);
nand NAND3 (N521, N507, N242, N147);
and AND2 (N522, N518, N444);
or OR4 (N523, N521, N349, N491, N407);
nor NOR4 (N524, N520, N335, N161, N190);
nand NAND3 (N525, N522, N5, N325);
not NOT1 (N526, N523);
nor NOR3 (N527, N511, N18, N261);
nand NAND4 (N528, N516, N314, N507, N67);
nand NAND4 (N529, N495, N243, N268, N300);
or OR2 (N530, N506, N166);
buf BUF1 (N531, N524);
nor NOR2 (N532, N531, N472);
nor NOR2 (N533, N530, N506);
not NOT1 (N534, N528);
or OR2 (N535, N534, N158);
and AND2 (N536, N533, N188);
nand NAND4 (N537, N535, N198, N206, N493);
nor NOR2 (N538, N519, N301);
not NOT1 (N539, N529);
xor XOR2 (N540, N532, N209);
xor XOR2 (N541, N526, N56);
and AND4 (N542, N540, N159, N532, N14);
and AND4 (N543, N514, N402, N139, N223);
or OR4 (N544, N497, N529, N103, N138);
nor NOR3 (N545, N527, N355, N455);
xor XOR2 (N546, N539, N280);
nor NOR2 (N547, N544, N398);
buf BUF1 (N548, N542);
or OR3 (N549, N541, N273, N301);
not NOT1 (N550, N549);
or OR2 (N551, N538, N491);
nor NOR4 (N552, N545, N293, N334, N159);
xor XOR2 (N553, N548, N364);
xor XOR2 (N554, N537, N124);
nand NAND3 (N555, N547, N497, N237);
and AND3 (N556, N551, N179, N130);
not NOT1 (N557, N555);
or OR2 (N558, N536, N424);
buf BUF1 (N559, N543);
xor XOR2 (N560, N559, N404);
and AND3 (N561, N552, N307, N273);
and AND3 (N562, N560, N57, N147);
not NOT1 (N563, N561);
xor XOR2 (N564, N562, N171);
nand NAND4 (N565, N563, N397, N171, N558);
xor XOR2 (N566, N87, N510);
or OR4 (N567, N553, N545, N543, N342);
not NOT1 (N568, N554);
buf BUF1 (N569, N550);
and AND3 (N570, N546, N39, N155);
nor NOR4 (N571, N556, N149, N36, N532);
nand NAND4 (N572, N571, N164, N469, N172);
nor NOR3 (N573, N572, N202, N561);
not NOT1 (N574, N567);
xor XOR2 (N575, N570, N51);
nor NOR3 (N576, N569, N154, N142);
nor NOR2 (N577, N576, N165);
nor NOR4 (N578, N525, N533, N555, N371);
buf BUF1 (N579, N573);
and AND3 (N580, N557, N578, N343);
nor NOR2 (N581, N569, N67);
and AND3 (N582, N574, N448, N318);
nand NAND4 (N583, N582, N476, N175, N418);
nand NAND2 (N584, N580, N532);
nand NAND2 (N585, N568, N472);
buf BUF1 (N586, N564);
nand NAND2 (N587, N586, N371);
not NOT1 (N588, N583);
or OR2 (N589, N577, N128);
nor NOR3 (N590, N575, N310, N443);
not NOT1 (N591, N566);
buf BUF1 (N592, N588);
or OR2 (N593, N579, N447);
nand NAND4 (N594, N581, N67, N314, N390);
not NOT1 (N595, N565);
xor XOR2 (N596, N584, N241);
xor XOR2 (N597, N596, N430);
or OR4 (N598, N592, N188, N412, N222);
xor XOR2 (N599, N587, N202);
not NOT1 (N600, N589);
nor NOR3 (N601, N585, N242, N181);
and AND2 (N602, N593, N420);
xor XOR2 (N603, N597, N304);
not NOT1 (N604, N598);
or OR4 (N605, N595, N331, N349, N70);
buf BUF1 (N606, N601);
and AND2 (N607, N600, N550);
not NOT1 (N608, N604);
or OR4 (N609, N602, N207, N64, N411);
buf BUF1 (N610, N609);
nand NAND4 (N611, N603, N3, N262, N195);
xor XOR2 (N612, N599, N332);
xor XOR2 (N613, N606, N282);
buf BUF1 (N614, N613);
nand NAND4 (N615, N591, N555, N494, N471);
not NOT1 (N616, N611);
or OR2 (N617, N614, N380);
xor XOR2 (N618, N594, N134);
nor NOR4 (N619, N608, N86, N275, N35);
and AND2 (N620, N610, N336);
xor XOR2 (N621, N612, N136);
nand NAND2 (N622, N616, N132);
and AND3 (N623, N615, N149, N20);
and AND4 (N624, N605, N476, N212, N295);
nand NAND2 (N625, N617, N135);
not NOT1 (N626, N624);
nor NOR3 (N627, N619, N411, N69);
xor XOR2 (N628, N620, N490);
not NOT1 (N629, N622);
buf BUF1 (N630, N623);
nand NAND4 (N631, N630, N145, N448, N178);
not NOT1 (N632, N590);
nand NAND2 (N633, N629, N2);
nand NAND2 (N634, N618, N431);
buf BUF1 (N635, N625);
not NOT1 (N636, N632);
buf BUF1 (N637, N626);
xor XOR2 (N638, N633, N429);
nor NOR3 (N639, N637, N480, N65);
and AND3 (N640, N638, N289, N245);
xor XOR2 (N641, N634, N141);
buf BUF1 (N642, N631);
not NOT1 (N643, N641);
and AND4 (N644, N639, N471, N423, N63);
xor XOR2 (N645, N607, N224);
nor NOR2 (N646, N636, N490);
and AND2 (N647, N640, N340);
xor XOR2 (N648, N647, N152);
xor XOR2 (N649, N635, N362);
or OR4 (N650, N643, N127, N550, N274);
nor NOR3 (N651, N649, N627, N248);
or OR3 (N652, N284, N422, N424);
buf BUF1 (N653, N621);
or OR2 (N654, N653, N281);
buf BUF1 (N655, N648);
nor NOR2 (N656, N628, N196);
or OR2 (N657, N652, N298);
or OR2 (N658, N645, N558);
or OR4 (N659, N656, N253, N37, N618);
or OR2 (N660, N657, N76);
xor XOR2 (N661, N655, N285);
xor XOR2 (N662, N659, N408);
not NOT1 (N663, N651);
xor XOR2 (N664, N650, N552);
buf BUF1 (N665, N654);
nand NAND2 (N666, N665, N116);
and AND2 (N667, N662, N353);
xor XOR2 (N668, N642, N664);
and AND4 (N669, N148, N589, N568, N645);
or OR3 (N670, N658, N347, N33);
nand NAND3 (N671, N669, N372, N416);
buf BUF1 (N672, N663);
not NOT1 (N673, N660);
or OR3 (N674, N646, N200, N28);
xor XOR2 (N675, N661, N406);
xor XOR2 (N676, N670, N352);
buf BUF1 (N677, N666);
buf BUF1 (N678, N673);
nor NOR2 (N679, N676, N490);
nand NAND3 (N680, N667, N336, N270);
nand NAND2 (N681, N677, N91);
or OR2 (N682, N679, N188);
nand NAND4 (N683, N644, N471, N511, N63);
nand NAND3 (N684, N683, N335, N377);
not NOT1 (N685, N682);
not NOT1 (N686, N684);
buf BUF1 (N687, N686);
and AND2 (N688, N687, N657);
nor NOR3 (N689, N672, N381, N279);
not NOT1 (N690, N674);
not NOT1 (N691, N689);
buf BUF1 (N692, N671);
nor NOR2 (N693, N688, N428);
nor NOR2 (N694, N691, N51);
not NOT1 (N695, N693);
and AND4 (N696, N678, N215, N227, N351);
nand NAND4 (N697, N694, N146, N523, N472);
or OR2 (N698, N680, N541);
and AND2 (N699, N698, N118);
and AND3 (N700, N681, N202, N17);
not NOT1 (N701, N685);
and AND4 (N702, N700, N603, N7, N666);
xor XOR2 (N703, N692, N678);
xor XOR2 (N704, N702, N409);
and AND4 (N705, N703, N456, N316, N356);
and AND4 (N706, N705, N637, N389, N397);
xor XOR2 (N707, N696, N530);
buf BUF1 (N708, N668);
and AND3 (N709, N697, N108, N386);
buf BUF1 (N710, N706);
xor XOR2 (N711, N695, N677);
buf BUF1 (N712, N710);
buf BUF1 (N713, N709);
nand NAND2 (N714, N690, N299);
and AND4 (N715, N714, N302, N47, N14);
nor NOR4 (N716, N715, N626, N369, N425);
buf BUF1 (N717, N711);
nand NAND4 (N718, N704, N126, N186, N448);
nand NAND4 (N719, N712, N504, N497, N114);
nor NOR4 (N720, N713, N47, N698, N19);
and AND2 (N721, N719, N704);
xor XOR2 (N722, N707, N546);
nor NOR4 (N723, N718, N304, N421, N117);
not NOT1 (N724, N723);
xor XOR2 (N725, N722, N194);
nand NAND3 (N726, N724, N518, N656);
buf BUF1 (N727, N708);
or OR4 (N728, N675, N190, N396, N462);
or OR4 (N729, N721, N693, N121, N136);
xor XOR2 (N730, N716, N436);
not NOT1 (N731, N699);
nor NOR2 (N732, N720, N238);
or OR3 (N733, N725, N415, N216);
buf BUF1 (N734, N701);
and AND4 (N735, N717, N140, N734, N344);
nand NAND2 (N736, N176, N464);
and AND3 (N737, N727, N495, N727);
not NOT1 (N738, N737);
buf BUF1 (N739, N730);
nand NAND4 (N740, N733, N110, N154, N408);
nor NOR3 (N741, N729, N84, N576);
and AND4 (N742, N736, N425, N445, N434);
xor XOR2 (N743, N741, N149);
nor NOR2 (N744, N732, N457);
buf BUF1 (N745, N739);
and AND3 (N746, N742, N122, N370);
nand NAND3 (N747, N735, N310, N310);
and AND4 (N748, N728, N575, N322, N620);
and AND4 (N749, N745, N204, N222, N515);
nand NAND3 (N750, N749, N499, N134);
not NOT1 (N751, N747);
nor NOR4 (N752, N740, N361, N745, N491);
and AND4 (N753, N751, N31, N19, N750);
xor XOR2 (N754, N72, N209);
buf BUF1 (N755, N753);
and AND4 (N756, N744, N72, N190, N284);
not NOT1 (N757, N748);
and AND4 (N758, N743, N387, N305, N53);
or OR4 (N759, N746, N183, N650, N339);
nand NAND3 (N760, N726, N590, N731);
buf BUF1 (N761, N31);
buf BUF1 (N762, N758);
nor NOR4 (N763, N754, N265, N260, N122);
not NOT1 (N764, N752);
not NOT1 (N765, N763);
nand NAND2 (N766, N762, N293);
or OR4 (N767, N755, N128, N406, N662);
xor XOR2 (N768, N759, N633);
nand NAND3 (N769, N756, N384, N250);
and AND3 (N770, N766, N699, N358);
nor NOR4 (N771, N757, N499, N310, N238);
or OR3 (N772, N770, N358, N279);
not NOT1 (N773, N772);
nand NAND4 (N774, N767, N722, N708, N625);
or OR3 (N775, N769, N107, N38);
xor XOR2 (N776, N774, N562);
nand NAND3 (N777, N773, N667, N656);
and AND3 (N778, N777, N86, N110);
xor XOR2 (N779, N771, N715);
and AND2 (N780, N778, N278);
nand NAND3 (N781, N775, N340, N578);
xor XOR2 (N782, N779, N716);
and AND4 (N783, N776, N769, N479, N433);
or OR2 (N784, N768, N374);
nand NAND2 (N785, N780, N640);
nor NOR3 (N786, N781, N313, N99);
not NOT1 (N787, N765);
xor XOR2 (N788, N761, N412);
nand NAND3 (N789, N783, N172, N409);
or OR4 (N790, N785, N203, N173, N484);
or OR2 (N791, N764, N614);
xor XOR2 (N792, N738, N470);
buf BUF1 (N793, N791);
or OR2 (N794, N792, N697);
nor NOR4 (N795, N789, N500, N600, N327);
and AND3 (N796, N790, N292, N225);
nand NAND2 (N797, N782, N690);
nor NOR2 (N798, N786, N635);
xor XOR2 (N799, N798, N436);
nor NOR2 (N800, N799, N382);
buf BUF1 (N801, N760);
not NOT1 (N802, N795);
nand NAND4 (N803, N794, N622, N323, N253);
buf BUF1 (N804, N796);
xor XOR2 (N805, N801, N323);
xor XOR2 (N806, N797, N575);
or OR2 (N807, N784, N215);
xor XOR2 (N808, N806, N294);
nor NOR2 (N809, N807, N163);
xor XOR2 (N810, N809, N572);
nand NAND2 (N811, N810, N99);
and AND2 (N812, N793, N77);
nor NOR4 (N813, N802, N668, N803, N92);
xor XOR2 (N814, N349, N676);
buf BUF1 (N815, N812);
nor NOR2 (N816, N800, N189);
not NOT1 (N817, N811);
and AND4 (N818, N813, N103, N306, N273);
nor NOR4 (N819, N804, N150, N205, N621);
buf BUF1 (N820, N819);
not NOT1 (N821, N805);
or OR2 (N822, N817, N97);
nand NAND3 (N823, N821, N749, N459);
and AND2 (N824, N788, N145);
not NOT1 (N825, N824);
nand NAND4 (N826, N825, N433, N711, N105);
or OR3 (N827, N815, N81, N28);
and AND4 (N828, N816, N260, N64, N527);
nor NOR4 (N829, N808, N752, N58, N814);
not NOT1 (N830, N572);
or OR3 (N831, N822, N230, N90);
not NOT1 (N832, N829);
nand NAND2 (N833, N820, N646);
and AND3 (N834, N787, N474, N44);
xor XOR2 (N835, N831, N135);
xor XOR2 (N836, N832, N29);
and AND4 (N837, N823, N185, N708, N79);
not NOT1 (N838, N827);
nor NOR3 (N839, N835, N155, N645);
xor XOR2 (N840, N828, N426);
xor XOR2 (N841, N839, N526);
nor NOR2 (N842, N836, N6);
xor XOR2 (N843, N830, N584);
not NOT1 (N844, N841);
nor NOR3 (N845, N842, N527, N399);
not NOT1 (N846, N838);
or OR3 (N847, N840, N419, N481);
nand NAND2 (N848, N818, N843);
nor NOR2 (N849, N792, N614);
xor XOR2 (N850, N834, N257);
nand NAND4 (N851, N847, N763, N365, N451);
buf BUF1 (N852, N846);
nand NAND4 (N853, N849, N372, N327, N715);
not NOT1 (N854, N851);
not NOT1 (N855, N844);
and AND2 (N856, N852, N670);
and AND3 (N857, N853, N56, N86);
buf BUF1 (N858, N854);
and AND4 (N859, N857, N703, N810, N840);
and AND4 (N860, N833, N579, N676, N508);
and AND4 (N861, N860, N653, N618, N496);
and AND3 (N862, N826, N709, N818);
nand NAND2 (N863, N858, N6);
and AND3 (N864, N859, N159, N458);
or OR2 (N865, N856, N535);
nand NAND4 (N866, N855, N773, N253, N723);
or OR3 (N867, N845, N116, N583);
buf BUF1 (N868, N861);
or OR2 (N869, N862, N171);
not NOT1 (N870, N865);
nand NAND4 (N871, N866, N353, N232, N779);
or OR2 (N872, N837, N34);
nor NOR3 (N873, N848, N533, N721);
or OR4 (N874, N871, N153, N290, N202);
nor NOR4 (N875, N869, N390, N788, N288);
and AND4 (N876, N864, N440, N329, N486);
and AND4 (N877, N874, N791, N681, N101);
buf BUF1 (N878, N877);
and AND4 (N879, N867, N675, N730, N259);
and AND4 (N880, N879, N365, N848, N219);
nand NAND3 (N881, N878, N485, N176);
xor XOR2 (N882, N873, N619);
not NOT1 (N883, N880);
and AND3 (N884, N868, N30, N813);
and AND2 (N885, N872, N162);
and AND4 (N886, N885, N86, N762, N872);
or OR3 (N887, N881, N314, N824);
xor XOR2 (N888, N887, N212);
nand NAND4 (N889, N883, N519, N731, N208);
buf BUF1 (N890, N884);
xor XOR2 (N891, N882, N686);
nand NAND2 (N892, N891, N532);
and AND3 (N893, N876, N529, N408);
nor NOR2 (N894, N863, N39);
and AND3 (N895, N890, N82, N551);
and AND3 (N896, N870, N40, N253);
nor NOR4 (N897, N893, N875, N787, N529);
buf BUF1 (N898, N823);
and AND3 (N899, N850, N802, N662);
nand NAND3 (N900, N892, N679, N755);
not NOT1 (N901, N896);
xor XOR2 (N902, N901, N328);
buf BUF1 (N903, N899);
nor NOR2 (N904, N903, N881);
nand NAND2 (N905, N888, N893);
nand NAND2 (N906, N894, N159);
nor NOR2 (N907, N897, N209);
or OR3 (N908, N902, N904, N464);
nand NAND2 (N909, N18, N758);
nand NAND3 (N910, N907, N95, N314);
buf BUF1 (N911, N900);
or OR3 (N912, N909, N253, N593);
or OR2 (N913, N895, N616);
not NOT1 (N914, N906);
nor NOR4 (N915, N913, N326, N511, N349);
xor XOR2 (N916, N915, N778);
and AND2 (N917, N886, N404);
and AND4 (N918, N908, N448, N559, N204);
and AND3 (N919, N914, N491, N46);
and AND4 (N920, N918, N711, N919, N417);
nor NOR2 (N921, N861, N790);
not NOT1 (N922, N916);
not NOT1 (N923, N912);
xor XOR2 (N924, N898, N519);
xor XOR2 (N925, N923, N264);
buf BUF1 (N926, N925);
nor NOR3 (N927, N924, N369, N358);
and AND4 (N928, N922, N758, N15, N227);
nand NAND3 (N929, N917, N273, N326);
or OR4 (N930, N929, N581, N599, N120);
nand NAND2 (N931, N921, N115);
not NOT1 (N932, N911);
not NOT1 (N933, N928);
xor XOR2 (N934, N927, N553);
buf BUF1 (N935, N889);
nand NAND3 (N936, N910, N295, N290);
not NOT1 (N937, N926);
nand NAND4 (N938, N920, N857, N768, N217);
not NOT1 (N939, N930);
nand NAND3 (N940, N936, N366, N445);
and AND3 (N941, N935, N822, N734);
not NOT1 (N942, N940);
or OR3 (N943, N942, N713, N173);
xor XOR2 (N944, N932, N396);
and AND2 (N945, N939, N134);
and AND2 (N946, N938, N913);
nand NAND2 (N947, N933, N646);
or OR3 (N948, N947, N186, N732);
buf BUF1 (N949, N945);
not NOT1 (N950, N931);
buf BUF1 (N951, N937);
and AND4 (N952, N905, N601, N430, N799);
or OR3 (N953, N941, N481, N2);
buf BUF1 (N954, N953);
xor XOR2 (N955, N934, N799);
nand NAND3 (N956, N944, N381, N911);
xor XOR2 (N957, N951, N887);
nor NOR2 (N958, N956, N407);
nor NOR4 (N959, N955, N833, N937, N656);
or OR3 (N960, N950, N843, N941);
nor NOR2 (N961, N952, N123);
and AND4 (N962, N957, N5, N99, N889);
buf BUF1 (N963, N943);
not NOT1 (N964, N962);
or OR2 (N965, N949, N34);
nand NAND4 (N966, N961, N15, N912, N617);
or OR3 (N967, N959, N34, N871);
nand NAND2 (N968, N966, N187);
nand NAND2 (N969, N964, N854);
not NOT1 (N970, N954);
nor NOR2 (N971, N969, N194);
buf BUF1 (N972, N970);
or OR4 (N973, N946, N934, N412, N274);
nand NAND4 (N974, N971, N603, N828, N388);
nand NAND2 (N975, N960, N708);
or OR2 (N976, N965, N93);
not NOT1 (N977, N973);
nor NOR3 (N978, N967, N260, N341);
nand NAND3 (N979, N974, N665, N552);
nor NOR2 (N980, N975, N364);
and AND2 (N981, N977, N783);
buf BUF1 (N982, N981);
nand NAND2 (N983, N976, N918);
buf BUF1 (N984, N948);
buf BUF1 (N985, N983);
and AND4 (N986, N968, N460, N429, N385);
or OR2 (N987, N978, N867);
not NOT1 (N988, N963);
nor NOR3 (N989, N980, N135, N436);
not NOT1 (N990, N989);
and AND3 (N991, N958, N65, N620);
or OR3 (N992, N984, N223, N728);
or OR2 (N993, N987, N721);
nor NOR4 (N994, N992, N637, N190, N97);
nand NAND4 (N995, N972, N620, N109, N249);
nand NAND2 (N996, N991, N170);
nand NAND3 (N997, N985, N947, N300);
nand NAND2 (N998, N982, N863);
nand NAND3 (N999, N986, N98, N617);
nor NOR4 (N1000, N993, N928, N971, N24);
or OR3 (N1001, N979, N783, N654);
nand NAND2 (N1002, N1001, N280);
not NOT1 (N1003, N988);
buf BUF1 (N1004, N999);
nor NOR4 (N1005, N998, N717, N593, N126);
xor XOR2 (N1006, N1003, N593);
xor XOR2 (N1007, N1002, N524);
not NOT1 (N1008, N1004);
nand NAND2 (N1009, N996, N865);
nor NOR3 (N1010, N995, N928, N700);
and AND2 (N1011, N1000, N265);
nand NAND3 (N1012, N1011, N174, N7);
xor XOR2 (N1013, N994, N459);
nor NOR2 (N1014, N1006, N64);
or OR4 (N1015, N1009, N834, N426, N354);
xor XOR2 (N1016, N1008, N345);
or OR4 (N1017, N1016, N874, N923, N562);
nand NAND3 (N1018, N1013, N878, N860);
nor NOR4 (N1019, N1014, N697, N466, N159);
and AND4 (N1020, N1012, N800, N810, N824);
buf BUF1 (N1021, N1010);
not NOT1 (N1022, N1021);
not NOT1 (N1023, N1018);
buf BUF1 (N1024, N1022);
or OR3 (N1025, N1024, N898, N952);
nand NAND3 (N1026, N1023, N109, N1013);
nor NOR4 (N1027, N990, N865, N14, N882);
nor NOR2 (N1028, N1027, N548);
nor NOR3 (N1029, N1019, N734, N47);
nor NOR4 (N1030, N1029, N878, N851, N132);
xor XOR2 (N1031, N997, N24);
xor XOR2 (N1032, N1031, N330);
xor XOR2 (N1033, N1020, N648);
not NOT1 (N1034, N1032);
nand NAND4 (N1035, N1026, N114, N840, N671);
buf BUF1 (N1036, N1034);
and AND3 (N1037, N1017, N206, N976);
xor XOR2 (N1038, N1007, N430);
xor XOR2 (N1039, N1005, N88);
and AND4 (N1040, N1035, N595, N355, N867);
not NOT1 (N1041, N1039);
nand NAND4 (N1042, N1041, N899, N785, N161);
buf BUF1 (N1043, N1038);
buf BUF1 (N1044, N1042);
nand NAND4 (N1045, N1030, N240, N413, N523);
nor NOR4 (N1046, N1028, N412, N820, N773);
nor NOR2 (N1047, N1015, N471);
buf BUF1 (N1048, N1045);
nand NAND4 (N1049, N1043, N1037, N260, N502);
nand NAND3 (N1050, N159, N246, N515);
not NOT1 (N1051, N1047);
buf BUF1 (N1052, N1044);
nor NOR3 (N1053, N1049, N194, N413);
nor NOR4 (N1054, N1025, N26, N1004, N123);
xor XOR2 (N1055, N1052, N260);
or OR3 (N1056, N1033, N473, N975);
xor XOR2 (N1057, N1056, N210);
xor XOR2 (N1058, N1055, N662);
and AND4 (N1059, N1053, N259, N689, N57);
not NOT1 (N1060, N1057);
and AND4 (N1061, N1046, N368, N795, N817);
or OR2 (N1062, N1054, N476);
nor NOR3 (N1063, N1048, N324, N648);
buf BUF1 (N1064, N1051);
not NOT1 (N1065, N1050);
xor XOR2 (N1066, N1062, N161);
or OR3 (N1067, N1065, N290, N455);
or OR3 (N1068, N1036, N610, N921);
nor NOR4 (N1069, N1067, N374, N135, N736);
not NOT1 (N1070, N1069);
nand NAND2 (N1071, N1061, N284);
not NOT1 (N1072, N1058);
or OR3 (N1073, N1066, N197, N304);
xor XOR2 (N1074, N1040, N328);
nor NOR2 (N1075, N1063, N187);
and AND2 (N1076, N1064, N611);
xor XOR2 (N1077, N1073, N982);
nand NAND3 (N1078, N1059, N847, N846);
and AND3 (N1079, N1070, N772, N812);
or OR3 (N1080, N1077, N663, N610);
nand NAND3 (N1081, N1071, N646, N188);
nand NAND3 (N1082, N1060, N288, N180);
buf BUF1 (N1083, N1074);
nor NOR4 (N1084, N1068, N11, N369, N291);
or OR4 (N1085, N1072, N1046, N663, N358);
xor XOR2 (N1086, N1085, N737);
xor XOR2 (N1087, N1079, N154);
buf BUF1 (N1088, N1086);
and AND3 (N1089, N1078, N702, N969);
buf BUF1 (N1090, N1082);
buf BUF1 (N1091, N1075);
not NOT1 (N1092, N1087);
and AND4 (N1093, N1076, N754, N407, N819);
xor XOR2 (N1094, N1080, N345);
nor NOR3 (N1095, N1090, N432, N372);
xor XOR2 (N1096, N1093, N523);
nand NAND3 (N1097, N1084, N87, N1016);
or OR4 (N1098, N1089, N53, N74, N795);
or OR2 (N1099, N1081, N540);
nor NOR2 (N1100, N1094, N128);
nor NOR4 (N1101, N1092, N858, N1024, N756);
nor NOR2 (N1102, N1083, N41);
or OR2 (N1103, N1102, N412);
and AND3 (N1104, N1096, N527, N155);
not NOT1 (N1105, N1098);
buf BUF1 (N1106, N1103);
and AND4 (N1107, N1091, N491, N658, N154);
nor NOR3 (N1108, N1097, N449, N265);
xor XOR2 (N1109, N1108, N366);
nand NAND4 (N1110, N1095, N140, N593, N432);
nand NAND4 (N1111, N1109, N169, N998, N8);
xor XOR2 (N1112, N1088, N754);
or OR4 (N1113, N1101, N129, N468, N612);
nand NAND3 (N1114, N1100, N448, N499);
nand NAND4 (N1115, N1111, N1062, N134, N920);
nand NAND3 (N1116, N1114, N374, N1016);
or OR2 (N1117, N1106, N1104);
and AND2 (N1118, N594, N1035);
nand NAND4 (N1119, N1116, N410, N11, N910);
nand NAND4 (N1120, N1113, N923, N1055, N886);
buf BUF1 (N1121, N1118);
and AND4 (N1122, N1110, N746, N15, N938);
and AND4 (N1123, N1105, N980, N596, N801);
xor XOR2 (N1124, N1115, N573);
or OR4 (N1125, N1122, N1049, N791, N285);
nor NOR2 (N1126, N1121, N49);
nor NOR3 (N1127, N1125, N718, N1089);
nand NAND2 (N1128, N1119, N715);
xor XOR2 (N1129, N1112, N119);
nand NAND2 (N1130, N1120, N325);
nor NOR3 (N1131, N1099, N707, N400);
and AND2 (N1132, N1127, N457);
nand NAND4 (N1133, N1129, N635, N483, N946);
and AND3 (N1134, N1107, N882, N983);
nand NAND3 (N1135, N1130, N1003, N552);
nand NAND3 (N1136, N1123, N914, N972);
xor XOR2 (N1137, N1131, N925);
and AND3 (N1138, N1117, N423, N530);
not NOT1 (N1139, N1133);
not NOT1 (N1140, N1136);
and AND4 (N1141, N1126, N1000, N720, N669);
or OR4 (N1142, N1128, N1132, N537, N144);
buf BUF1 (N1143, N553);
nor NOR4 (N1144, N1140, N356, N870, N161);
and AND2 (N1145, N1135, N832);
or OR2 (N1146, N1134, N397);
nor NOR3 (N1147, N1142, N471, N219);
buf BUF1 (N1148, N1145);
and AND2 (N1149, N1141, N30);
buf BUF1 (N1150, N1137);
not NOT1 (N1151, N1147);
nor NOR2 (N1152, N1144, N261);
or OR2 (N1153, N1139, N673);
buf BUF1 (N1154, N1153);
not NOT1 (N1155, N1150);
buf BUF1 (N1156, N1138);
not NOT1 (N1157, N1151);
nor NOR3 (N1158, N1152, N332, N505);
not NOT1 (N1159, N1148);
not NOT1 (N1160, N1154);
not NOT1 (N1161, N1149);
xor XOR2 (N1162, N1155, N1095);
buf BUF1 (N1163, N1160);
buf BUF1 (N1164, N1146);
buf BUF1 (N1165, N1156);
buf BUF1 (N1166, N1165);
nor NOR4 (N1167, N1163, N147, N1101, N1058);
nor NOR2 (N1168, N1124, N237);
or OR2 (N1169, N1164, N587);
and AND3 (N1170, N1143, N868, N144);
nand NAND4 (N1171, N1158, N777, N330, N390);
xor XOR2 (N1172, N1157, N148);
nand NAND3 (N1173, N1166, N719, N195);
buf BUF1 (N1174, N1172);
nand NAND4 (N1175, N1159, N939, N1016, N925);
not NOT1 (N1176, N1162);
nor NOR3 (N1177, N1169, N109, N1059);
and AND4 (N1178, N1177, N635, N1000, N1153);
not NOT1 (N1179, N1175);
xor XOR2 (N1180, N1173, N1133);
not NOT1 (N1181, N1167);
nor NOR3 (N1182, N1170, N754, N489);
buf BUF1 (N1183, N1168);
nor NOR4 (N1184, N1181, N573, N746, N1176);
nor NOR3 (N1185, N965, N923, N924);
not NOT1 (N1186, N1182);
not NOT1 (N1187, N1184);
nor NOR4 (N1188, N1171, N538, N225, N288);
xor XOR2 (N1189, N1180, N686);
xor XOR2 (N1190, N1179, N714);
nand NAND2 (N1191, N1186, N826);
and AND3 (N1192, N1174, N344, N358);
nand NAND2 (N1193, N1187, N1013);
nor NOR4 (N1194, N1190, N372, N725, N623);
nand NAND4 (N1195, N1191, N294, N1021, N512);
nor NOR2 (N1196, N1189, N699);
xor XOR2 (N1197, N1185, N1188);
or OR2 (N1198, N706, N986);
xor XOR2 (N1199, N1194, N56);
nand NAND3 (N1200, N1192, N576, N393);
and AND3 (N1201, N1198, N408, N440);
and AND2 (N1202, N1201, N117);
nand NAND3 (N1203, N1196, N52, N164);
xor XOR2 (N1204, N1199, N388);
xor XOR2 (N1205, N1200, N1160);
and AND2 (N1206, N1178, N431);
buf BUF1 (N1207, N1203);
buf BUF1 (N1208, N1202);
buf BUF1 (N1209, N1195);
nor NOR3 (N1210, N1161, N39, N748);
xor XOR2 (N1211, N1209, N14);
and AND3 (N1212, N1193, N787, N977);
and AND3 (N1213, N1204, N72, N1182);
and AND3 (N1214, N1197, N1053, N128);
buf BUF1 (N1215, N1210);
buf BUF1 (N1216, N1206);
xor XOR2 (N1217, N1211, N1071);
and AND3 (N1218, N1214, N737, N348);
or OR4 (N1219, N1217, N302, N558, N938);
buf BUF1 (N1220, N1213);
buf BUF1 (N1221, N1205);
xor XOR2 (N1222, N1219, N124);
not NOT1 (N1223, N1183);
not NOT1 (N1224, N1207);
nand NAND3 (N1225, N1220, N511, N94);
xor XOR2 (N1226, N1218, N905);
xor XOR2 (N1227, N1212, N1222);
and AND4 (N1228, N1003, N1135, N1036, N1107);
nor NOR3 (N1229, N1215, N349, N599);
nor NOR4 (N1230, N1228, N126, N1167, N105);
xor XOR2 (N1231, N1216, N493);
buf BUF1 (N1232, N1208);
nor NOR2 (N1233, N1231, N84);
nor NOR2 (N1234, N1232, N137);
nand NAND4 (N1235, N1233, N107, N438, N721);
or OR3 (N1236, N1234, N89, N1181);
xor XOR2 (N1237, N1227, N275);
or OR4 (N1238, N1224, N794, N324, N379);
nand NAND2 (N1239, N1235, N741);
nor NOR3 (N1240, N1225, N1124, N207);
nand NAND4 (N1241, N1230, N404, N414, N219);
xor XOR2 (N1242, N1229, N846);
nor NOR2 (N1243, N1223, N514);
or OR4 (N1244, N1237, N13, N572, N549);
xor XOR2 (N1245, N1241, N230);
not NOT1 (N1246, N1244);
and AND3 (N1247, N1238, N1131, N1102);
or OR2 (N1248, N1239, N607);
buf BUF1 (N1249, N1247);
or OR2 (N1250, N1246, N560);
buf BUF1 (N1251, N1245);
xor XOR2 (N1252, N1243, N622);
nor NOR4 (N1253, N1221, N161, N347, N389);
xor XOR2 (N1254, N1240, N374);
nand NAND2 (N1255, N1236, N649);
nand NAND2 (N1256, N1242, N512);
or OR3 (N1257, N1249, N334, N459);
nand NAND4 (N1258, N1257, N153, N685, N484);
xor XOR2 (N1259, N1250, N423);
not NOT1 (N1260, N1253);
xor XOR2 (N1261, N1259, N211);
or OR3 (N1262, N1261, N522, N882);
nor NOR2 (N1263, N1258, N174);
not NOT1 (N1264, N1251);
xor XOR2 (N1265, N1252, N1234);
buf BUF1 (N1266, N1256);
and AND2 (N1267, N1248, N1082);
nand NAND3 (N1268, N1264, N25, N801);
and AND4 (N1269, N1263, N558, N1041, N437);
nor NOR4 (N1270, N1262, N56, N1013, N768);
nand NAND4 (N1271, N1255, N253, N147, N238);
nor NOR3 (N1272, N1268, N609, N128);
not NOT1 (N1273, N1226);
and AND4 (N1274, N1273, N28, N728, N414);
nor NOR3 (N1275, N1254, N1188, N766);
nor NOR3 (N1276, N1275, N1116, N1087);
xor XOR2 (N1277, N1260, N650);
nand NAND4 (N1278, N1277, N1124, N648, N1181);
xor XOR2 (N1279, N1271, N32);
buf BUF1 (N1280, N1267);
and AND3 (N1281, N1274, N1266, N950);
or OR3 (N1282, N356, N315, N401);
or OR2 (N1283, N1272, N290);
not NOT1 (N1284, N1270);
buf BUF1 (N1285, N1265);
or OR2 (N1286, N1285, N705);
or OR4 (N1287, N1279, N43, N557, N832);
nor NOR4 (N1288, N1284, N952, N32, N994);
and AND4 (N1289, N1276, N423, N605, N1215);
nor NOR4 (N1290, N1287, N275, N624, N366);
nand NAND4 (N1291, N1269, N24, N79, N507);
nor NOR4 (N1292, N1281, N90, N1095, N839);
nor NOR3 (N1293, N1291, N943, N1060);
or OR3 (N1294, N1286, N1211, N376);
not NOT1 (N1295, N1294);
and AND4 (N1296, N1295, N159, N468, N857);
buf BUF1 (N1297, N1282);
nor NOR4 (N1298, N1290, N1164, N678, N316);
and AND4 (N1299, N1289, N979, N692, N795);
not NOT1 (N1300, N1299);
and AND3 (N1301, N1296, N172, N804);
not NOT1 (N1302, N1292);
nor NOR4 (N1303, N1300, N1012, N931, N305);
buf BUF1 (N1304, N1283);
nand NAND3 (N1305, N1301, N1139, N654);
and AND3 (N1306, N1298, N717, N599);
nor NOR2 (N1307, N1302, N1233);
buf BUF1 (N1308, N1306);
buf BUF1 (N1309, N1305);
buf BUF1 (N1310, N1307);
xor XOR2 (N1311, N1293, N293);
or OR3 (N1312, N1309, N1222, N248);
and AND4 (N1313, N1304, N621, N563, N215);
nor NOR2 (N1314, N1280, N1209);
not NOT1 (N1315, N1278);
not NOT1 (N1316, N1288);
and AND2 (N1317, N1303, N809);
or OR2 (N1318, N1311, N453);
or OR3 (N1319, N1310, N865, N540);
buf BUF1 (N1320, N1317);
buf BUF1 (N1321, N1316);
or OR2 (N1322, N1314, N1155);
and AND3 (N1323, N1319, N682, N565);
and AND3 (N1324, N1315, N462, N866);
xor XOR2 (N1325, N1321, N474);
nand NAND2 (N1326, N1297, N88);
and AND2 (N1327, N1313, N791);
and AND2 (N1328, N1322, N775);
or OR4 (N1329, N1308, N156, N1107, N1121);
nor NOR3 (N1330, N1324, N646, N838);
or OR4 (N1331, N1312, N136, N1137, N1052);
not NOT1 (N1332, N1328);
xor XOR2 (N1333, N1323, N821);
buf BUF1 (N1334, N1327);
buf BUF1 (N1335, N1330);
or OR4 (N1336, N1334, N1117, N1035, N303);
not NOT1 (N1337, N1318);
not NOT1 (N1338, N1337);
xor XOR2 (N1339, N1331, N345);
not NOT1 (N1340, N1338);
and AND3 (N1341, N1332, N307, N190);
buf BUF1 (N1342, N1340);
xor XOR2 (N1343, N1339, N1055);
or OR2 (N1344, N1326, N1183);
or OR3 (N1345, N1333, N808, N1086);
or OR2 (N1346, N1342, N634);
and AND4 (N1347, N1320, N443, N1301, N755);
nor NOR3 (N1348, N1343, N1121, N93);
nand NAND3 (N1349, N1335, N115, N93);
nor NOR2 (N1350, N1349, N1146);
nor NOR2 (N1351, N1347, N1138);
or OR2 (N1352, N1341, N294);
not NOT1 (N1353, N1329);
not NOT1 (N1354, N1336);
xor XOR2 (N1355, N1325, N1261);
and AND2 (N1356, N1352, N484);
nor NOR2 (N1357, N1346, N10);
or OR3 (N1358, N1344, N1025, N483);
not NOT1 (N1359, N1356);
xor XOR2 (N1360, N1348, N406);
xor XOR2 (N1361, N1358, N579);
buf BUF1 (N1362, N1359);
not NOT1 (N1363, N1350);
buf BUF1 (N1364, N1362);
or OR4 (N1365, N1363, N589, N1260, N1188);
or OR4 (N1366, N1353, N1256, N361, N116);
buf BUF1 (N1367, N1354);
not NOT1 (N1368, N1360);
not NOT1 (N1369, N1367);
xor XOR2 (N1370, N1368, N1007);
not NOT1 (N1371, N1370);
xor XOR2 (N1372, N1361, N173);
buf BUF1 (N1373, N1355);
buf BUF1 (N1374, N1345);
or OR2 (N1375, N1372, N932);
and AND4 (N1376, N1366, N1132, N222, N402);
xor XOR2 (N1377, N1357, N68);
or OR4 (N1378, N1373, N600, N281, N1244);
nor NOR2 (N1379, N1369, N275);
and AND4 (N1380, N1379, N568, N466, N738);
nand NAND2 (N1381, N1375, N80);
xor XOR2 (N1382, N1378, N1333);
not NOT1 (N1383, N1374);
or OR3 (N1384, N1381, N682, N920);
xor XOR2 (N1385, N1364, N664);
and AND3 (N1386, N1377, N236, N543);
nor NOR3 (N1387, N1385, N784, N188);
xor XOR2 (N1388, N1384, N1364);
not NOT1 (N1389, N1365);
nor NOR3 (N1390, N1351, N589, N718);
xor XOR2 (N1391, N1389, N477);
nor NOR2 (N1392, N1388, N1329);
not NOT1 (N1393, N1382);
or OR2 (N1394, N1391, N997);
not NOT1 (N1395, N1392);
buf BUF1 (N1396, N1393);
buf BUF1 (N1397, N1383);
nand NAND2 (N1398, N1394, N1006);
nand NAND2 (N1399, N1376, N930);
or OR4 (N1400, N1390, N1019, N1356, N236);
or OR3 (N1401, N1396, N773, N97);
or OR2 (N1402, N1386, N400);
not NOT1 (N1403, N1380);
not NOT1 (N1404, N1399);
xor XOR2 (N1405, N1397, N802);
or OR3 (N1406, N1401, N852, N960);
buf BUF1 (N1407, N1371);
and AND2 (N1408, N1395, N273);
xor XOR2 (N1409, N1403, N410);
not NOT1 (N1410, N1409);
and AND4 (N1411, N1405, N1340, N1021, N629);
not NOT1 (N1412, N1410);
nand NAND3 (N1413, N1387, N550, N397);
xor XOR2 (N1414, N1412, N428);
nor NOR4 (N1415, N1414, N550, N830, N181);
and AND4 (N1416, N1411, N334, N993, N636);
nand NAND2 (N1417, N1406, N462);
and AND2 (N1418, N1413, N924);
not NOT1 (N1419, N1402);
buf BUF1 (N1420, N1417);
buf BUF1 (N1421, N1420);
and AND3 (N1422, N1400, N580, N865);
nand NAND2 (N1423, N1407, N655);
and AND4 (N1424, N1398, N955, N237, N359);
not NOT1 (N1425, N1418);
xor XOR2 (N1426, N1421, N225);
or OR4 (N1427, N1415, N1060, N776, N1202);
nand NAND2 (N1428, N1425, N143);
buf BUF1 (N1429, N1416);
not NOT1 (N1430, N1427);
and AND4 (N1431, N1408, N1205, N1318, N351);
nand NAND3 (N1432, N1422, N429, N549);
xor XOR2 (N1433, N1424, N919);
xor XOR2 (N1434, N1404, N835);
or OR2 (N1435, N1433, N497);
and AND2 (N1436, N1423, N592);
not NOT1 (N1437, N1429);
nor NOR3 (N1438, N1430, N731, N298);
and AND2 (N1439, N1437, N811);
buf BUF1 (N1440, N1432);
or OR2 (N1441, N1431, N1359);
xor XOR2 (N1442, N1441, N547);
buf BUF1 (N1443, N1442);
nand NAND2 (N1444, N1419, N440);
nor NOR4 (N1445, N1435, N153, N655, N852);
and AND3 (N1446, N1444, N1243, N863);
buf BUF1 (N1447, N1434);
nand NAND3 (N1448, N1438, N188, N162);
not NOT1 (N1449, N1448);
not NOT1 (N1450, N1436);
and AND3 (N1451, N1446, N1188, N204);
not NOT1 (N1452, N1440);
buf BUF1 (N1453, N1443);
xor XOR2 (N1454, N1453, N174);
or OR2 (N1455, N1450, N725);
nor NOR3 (N1456, N1449, N444, N28);
buf BUF1 (N1457, N1451);
xor XOR2 (N1458, N1452, N8);
buf BUF1 (N1459, N1454);
nor NOR3 (N1460, N1426, N1007, N839);
xor XOR2 (N1461, N1447, N345);
nor NOR4 (N1462, N1457, N757, N196, N453);
and AND2 (N1463, N1439, N991);
nor NOR4 (N1464, N1460, N474, N339, N43);
nor NOR3 (N1465, N1463, N682, N551);
not NOT1 (N1466, N1465);
xor XOR2 (N1467, N1464, N332);
and AND4 (N1468, N1462, N1452, N536, N1272);
buf BUF1 (N1469, N1467);
and AND4 (N1470, N1428, N798, N385, N1254);
and AND3 (N1471, N1455, N1229, N39);
or OR4 (N1472, N1458, N1034, N1023, N595);
nor NOR2 (N1473, N1472, N915);
nor NOR3 (N1474, N1456, N499, N1262);
xor XOR2 (N1475, N1466, N1171);
nand NAND2 (N1476, N1470, N149);
buf BUF1 (N1477, N1474);
nand NAND3 (N1478, N1461, N734, N784);
buf BUF1 (N1479, N1468);
and AND3 (N1480, N1475, N392, N1054);
or OR2 (N1481, N1478, N1308);
or OR2 (N1482, N1481, N630);
nor NOR4 (N1483, N1479, N1317, N1151, N1429);
not NOT1 (N1484, N1482);
not NOT1 (N1485, N1476);
buf BUF1 (N1486, N1484);
buf BUF1 (N1487, N1473);
nor NOR3 (N1488, N1485, N547, N533);
buf BUF1 (N1489, N1486);
nor NOR4 (N1490, N1480, N1230, N1246, N270);
buf BUF1 (N1491, N1483);
not NOT1 (N1492, N1488);
buf BUF1 (N1493, N1471);
nor NOR4 (N1494, N1445, N60, N301, N970);
not NOT1 (N1495, N1459);
nand NAND4 (N1496, N1493, N225, N646, N365);
xor XOR2 (N1497, N1490, N1405);
xor XOR2 (N1498, N1497, N1096);
buf BUF1 (N1499, N1491);
and AND4 (N1500, N1477, N1270, N212, N1039);
or OR4 (N1501, N1494, N921, N976, N350);
buf BUF1 (N1502, N1499);
or OR3 (N1503, N1469, N167, N683);
xor XOR2 (N1504, N1496, N688);
nand NAND2 (N1505, N1498, N605);
or OR3 (N1506, N1503, N1025, N1066);
nand NAND4 (N1507, N1501, N223, N1170, N429);
and AND4 (N1508, N1495, N1264, N760, N1449);
xor XOR2 (N1509, N1489, N1404);
nor NOR3 (N1510, N1504, N31, N518);
xor XOR2 (N1511, N1502, N209);
nor NOR4 (N1512, N1509, N510, N701, N1312);
and AND4 (N1513, N1487, N741, N325, N39);
or OR2 (N1514, N1513, N733);
or OR2 (N1515, N1492, N931);
and AND2 (N1516, N1507, N786);
not NOT1 (N1517, N1508);
xor XOR2 (N1518, N1510, N1452);
xor XOR2 (N1519, N1515, N310);
nand NAND3 (N1520, N1511, N926, N903);
or OR3 (N1521, N1505, N973, N533);
xor XOR2 (N1522, N1521, N915);
and AND3 (N1523, N1516, N600, N594);
xor XOR2 (N1524, N1523, N826);
and AND4 (N1525, N1514, N26, N860, N1485);
nor NOR3 (N1526, N1520, N996, N847);
nand NAND3 (N1527, N1525, N241, N644);
nand NAND3 (N1528, N1506, N1423, N331);
xor XOR2 (N1529, N1500, N766);
nand NAND3 (N1530, N1524, N1225, N1052);
nand NAND4 (N1531, N1526, N384, N919, N437);
nand NAND4 (N1532, N1528, N76, N1127, N582);
buf BUF1 (N1533, N1532);
or OR3 (N1534, N1533, N46, N1518);
nand NAND4 (N1535, N135, N287, N1530, N1182);
not NOT1 (N1536, N39);
buf BUF1 (N1537, N1527);
nand NAND2 (N1538, N1512, N220);
not NOT1 (N1539, N1529);
or OR4 (N1540, N1539, N813, N777, N502);
xor XOR2 (N1541, N1517, N1306);
xor XOR2 (N1542, N1534, N76);
and AND3 (N1543, N1522, N1171, N1129);
nor NOR4 (N1544, N1541, N992, N845, N1111);
not NOT1 (N1545, N1542);
buf BUF1 (N1546, N1543);
nor NOR3 (N1547, N1537, N235, N1395);
and AND3 (N1548, N1536, N610, N898);
buf BUF1 (N1549, N1538);
not NOT1 (N1550, N1549);
nor NOR4 (N1551, N1550, N1126, N66, N923);
buf BUF1 (N1552, N1535);
not NOT1 (N1553, N1548);
xor XOR2 (N1554, N1551, N519);
buf BUF1 (N1555, N1553);
xor XOR2 (N1556, N1554, N1449);
xor XOR2 (N1557, N1556, N41);
nand NAND4 (N1558, N1552, N585, N1138, N783);
buf BUF1 (N1559, N1531);
nor NOR4 (N1560, N1546, N924, N245, N1483);
nor NOR4 (N1561, N1555, N646, N1250, N229);
buf BUF1 (N1562, N1545);
buf BUF1 (N1563, N1559);
nor NOR2 (N1564, N1544, N541);
nor NOR4 (N1565, N1519, N232, N886, N1478);
and AND2 (N1566, N1561, N152);
and AND2 (N1567, N1562, N1380);
nor NOR3 (N1568, N1566, N632, N1320);
xor XOR2 (N1569, N1547, N943);
not NOT1 (N1570, N1563);
buf BUF1 (N1571, N1557);
nor NOR4 (N1572, N1568, N318, N1373, N597);
nand NAND4 (N1573, N1558, N182, N898, N895);
xor XOR2 (N1574, N1572, N579);
or OR3 (N1575, N1574, N591, N112);
buf BUF1 (N1576, N1540);
buf BUF1 (N1577, N1564);
and AND3 (N1578, N1575, N500, N631);
or OR2 (N1579, N1573, N1139);
nand NAND3 (N1580, N1567, N1515, N990);
not NOT1 (N1581, N1565);
xor XOR2 (N1582, N1579, N21);
nand NAND4 (N1583, N1578, N1035, N429, N522);
or OR2 (N1584, N1560, N483);
or OR2 (N1585, N1583, N1);
buf BUF1 (N1586, N1576);
or OR3 (N1587, N1581, N118, N1025);
and AND4 (N1588, N1570, N1429, N1243, N255);
not NOT1 (N1589, N1584);
nand NAND2 (N1590, N1577, N819);
not NOT1 (N1591, N1589);
not NOT1 (N1592, N1588);
or OR4 (N1593, N1587, N1245, N984, N760);
or OR4 (N1594, N1580, N424, N214, N650);
xor XOR2 (N1595, N1582, N512);
xor XOR2 (N1596, N1591, N1174);
xor XOR2 (N1597, N1571, N1183);
nor NOR3 (N1598, N1596, N791, N1469);
nand NAND4 (N1599, N1594, N868, N26, N205);
not NOT1 (N1600, N1598);
or OR2 (N1601, N1585, N999);
or OR2 (N1602, N1597, N197);
not NOT1 (N1603, N1590);
buf BUF1 (N1604, N1603);
and AND4 (N1605, N1593, N520, N1526, N318);
nor NOR3 (N1606, N1586, N384, N1097);
not NOT1 (N1607, N1602);
not NOT1 (N1608, N1599);
buf BUF1 (N1609, N1569);
xor XOR2 (N1610, N1592, N760);
nor NOR2 (N1611, N1605, N547);
and AND3 (N1612, N1608, N1063, N968);
nand NAND2 (N1613, N1611, N526);
buf BUF1 (N1614, N1601);
nand NAND4 (N1615, N1604, N362, N1166, N707);
or OR4 (N1616, N1615, N1570, N1525, N1135);
buf BUF1 (N1617, N1609);
buf BUF1 (N1618, N1595);
buf BUF1 (N1619, N1617);
buf BUF1 (N1620, N1606);
not NOT1 (N1621, N1618);
buf BUF1 (N1622, N1612);
not NOT1 (N1623, N1613);
nand NAND2 (N1624, N1622, N1130);
nor NOR2 (N1625, N1620, N1171);
buf BUF1 (N1626, N1610);
or OR3 (N1627, N1614, N356, N828);
nand NAND2 (N1628, N1627, N537);
xor XOR2 (N1629, N1619, N1499);
nor NOR2 (N1630, N1623, N1309);
and AND4 (N1631, N1629, N406, N1510, N914);
or OR4 (N1632, N1624, N459, N1409, N585);
not NOT1 (N1633, N1626);
buf BUF1 (N1634, N1631);
buf BUF1 (N1635, N1625);
not NOT1 (N1636, N1621);
not NOT1 (N1637, N1628);
nor NOR4 (N1638, N1634, N1408, N787, N295);
not NOT1 (N1639, N1638);
nand NAND2 (N1640, N1639, N1078);
xor XOR2 (N1641, N1607, N662);
or OR2 (N1642, N1630, N891);
not NOT1 (N1643, N1632);
nor NOR2 (N1644, N1616, N1015);
xor XOR2 (N1645, N1633, N169);
buf BUF1 (N1646, N1641);
nand NAND3 (N1647, N1646, N594, N215);
buf BUF1 (N1648, N1635);
and AND4 (N1649, N1644, N618, N1115, N398);
not NOT1 (N1650, N1600);
or OR4 (N1651, N1642, N738, N1448, N1093);
or OR3 (N1652, N1643, N1393, N931);
and AND4 (N1653, N1648, N492, N930, N174);
buf BUF1 (N1654, N1640);
nor NOR4 (N1655, N1636, N866, N1616, N517);
xor XOR2 (N1656, N1637, N248);
nor NOR3 (N1657, N1645, N329, N898);
and AND3 (N1658, N1655, N1171, N889);
and AND4 (N1659, N1649, N590, N744, N1176);
xor XOR2 (N1660, N1659, N1602);
nand NAND4 (N1661, N1660, N720, N857, N336);
or OR4 (N1662, N1656, N143, N1479, N801);
xor XOR2 (N1663, N1650, N342);
not NOT1 (N1664, N1653);
or OR3 (N1665, N1647, N438, N557);
nand NAND2 (N1666, N1654, N10);
nand NAND3 (N1667, N1652, N219, N829);
xor XOR2 (N1668, N1661, N1411);
or OR2 (N1669, N1667, N148);
or OR4 (N1670, N1651, N1042, N210, N1418);
or OR4 (N1671, N1658, N148, N1433, N1347);
or OR2 (N1672, N1666, N1542);
xor XOR2 (N1673, N1662, N390);
xor XOR2 (N1674, N1665, N375);
nor NOR4 (N1675, N1669, N983, N498, N1194);
or OR3 (N1676, N1664, N1357, N1306);
xor XOR2 (N1677, N1675, N759);
nor NOR3 (N1678, N1657, N446, N719);
or OR3 (N1679, N1672, N1296, N732);
nor NOR3 (N1680, N1663, N1095, N717);
xor XOR2 (N1681, N1676, N132);
xor XOR2 (N1682, N1677, N3);
nor NOR4 (N1683, N1671, N390, N838, N1204);
or OR2 (N1684, N1670, N1672);
or OR3 (N1685, N1681, N128, N1624);
buf BUF1 (N1686, N1674);
xor XOR2 (N1687, N1678, N347);
xor XOR2 (N1688, N1679, N1605);
and AND4 (N1689, N1668, N560, N1347, N476);
nor NOR4 (N1690, N1684, N1173, N842, N417);
or OR2 (N1691, N1685, N57);
and AND3 (N1692, N1682, N773, N540);
nor NOR4 (N1693, N1688, N932, N523, N1397);
and AND4 (N1694, N1693, N1020, N1461, N35);
or OR2 (N1695, N1687, N628);
buf BUF1 (N1696, N1673);
not NOT1 (N1697, N1683);
nand NAND2 (N1698, N1680, N585);
not NOT1 (N1699, N1691);
and AND4 (N1700, N1686, N630, N684, N267);
or OR3 (N1701, N1698, N353, N203);
or OR2 (N1702, N1692, N1503);
and AND2 (N1703, N1689, N1409);
and AND3 (N1704, N1697, N1423, N706);
buf BUF1 (N1705, N1700);
not NOT1 (N1706, N1703);
and AND2 (N1707, N1699, N502);
or OR3 (N1708, N1696, N1296, N1526);
buf BUF1 (N1709, N1707);
nor NOR3 (N1710, N1708, N1572, N36);
or OR4 (N1711, N1706, N674, N1312, N53);
xor XOR2 (N1712, N1701, N545);
nor NOR2 (N1713, N1712, N472);
buf BUF1 (N1714, N1705);
xor XOR2 (N1715, N1695, N734);
and AND3 (N1716, N1713, N622, N247);
buf BUF1 (N1717, N1690);
and AND4 (N1718, N1710, N119, N182, N528);
nor NOR4 (N1719, N1711, N414, N38, N1474);
nand NAND2 (N1720, N1716, N96);
or OR3 (N1721, N1718, N417, N1699);
xor XOR2 (N1722, N1709, N1253);
not NOT1 (N1723, N1715);
and AND4 (N1724, N1723, N786, N714, N931);
nand NAND3 (N1725, N1721, N649, N1580);
buf BUF1 (N1726, N1719);
nor NOR4 (N1727, N1722, N418, N1145, N301);
xor XOR2 (N1728, N1702, N1232);
and AND2 (N1729, N1728, N526);
buf BUF1 (N1730, N1727);
xor XOR2 (N1731, N1694, N806);
not NOT1 (N1732, N1726);
and AND4 (N1733, N1725, N674, N589, N250);
xor XOR2 (N1734, N1731, N594);
nor NOR2 (N1735, N1733, N1671);
and AND3 (N1736, N1734, N1687, N946);
and AND4 (N1737, N1736, N1293, N299, N167);
xor XOR2 (N1738, N1720, N943);
nand NAND4 (N1739, N1714, N849, N99, N726);
or OR4 (N1740, N1732, N1315, N304, N892);
nand NAND2 (N1741, N1737, N640);
or OR2 (N1742, N1740, N693);
not NOT1 (N1743, N1729);
and AND3 (N1744, N1704, N1414, N13);
nand NAND3 (N1745, N1724, N304, N803);
nand NAND4 (N1746, N1741, N86, N983, N91);
and AND2 (N1747, N1743, N895);
xor XOR2 (N1748, N1747, N506);
xor XOR2 (N1749, N1748, N630);
nor NOR3 (N1750, N1735, N965, N292);
xor XOR2 (N1751, N1749, N900);
and AND4 (N1752, N1750, N815, N507, N1472);
xor XOR2 (N1753, N1751, N341);
buf BUF1 (N1754, N1738);
and AND4 (N1755, N1752, N353, N1160, N58);
or OR4 (N1756, N1753, N892, N532, N1203);
or OR4 (N1757, N1717, N477, N994, N765);
and AND4 (N1758, N1754, N463, N407, N1197);
nand NAND4 (N1759, N1755, N121, N927, N829);
nand NAND3 (N1760, N1758, N488, N1554);
nand NAND3 (N1761, N1730, N241, N1709);
not NOT1 (N1762, N1761);
nand NAND2 (N1763, N1744, N876);
nand NAND3 (N1764, N1760, N1460, N209);
and AND2 (N1765, N1757, N779);
buf BUF1 (N1766, N1756);
or OR3 (N1767, N1766, N1184, N1511);
or OR3 (N1768, N1762, N55, N386);
nand NAND4 (N1769, N1764, N1004, N1617, N1450);
not NOT1 (N1770, N1763);
nand NAND4 (N1771, N1769, N981, N691, N1068);
nand NAND3 (N1772, N1759, N404, N379);
nand NAND4 (N1773, N1746, N383, N1130, N885);
not NOT1 (N1774, N1765);
and AND2 (N1775, N1767, N1597);
nand NAND3 (N1776, N1775, N1204, N1408);
not NOT1 (N1777, N1739);
xor XOR2 (N1778, N1768, N886);
or OR4 (N1779, N1776, N524, N1018, N1404);
not NOT1 (N1780, N1774);
nand NAND4 (N1781, N1780, N648, N1231, N60);
buf BUF1 (N1782, N1745);
nand NAND2 (N1783, N1777, N1497);
or OR2 (N1784, N1770, N540);
buf BUF1 (N1785, N1784);
buf BUF1 (N1786, N1742);
xor XOR2 (N1787, N1778, N899);
or OR3 (N1788, N1783, N356, N1522);
buf BUF1 (N1789, N1781);
buf BUF1 (N1790, N1789);
xor XOR2 (N1791, N1771, N417);
nand NAND3 (N1792, N1788, N155, N334);
not NOT1 (N1793, N1773);
buf BUF1 (N1794, N1779);
nand NAND2 (N1795, N1772, N1629);
nand NAND3 (N1796, N1792, N1596, N1281);
nand NAND4 (N1797, N1790, N1335, N1106, N1172);
not NOT1 (N1798, N1782);
and AND4 (N1799, N1797, N588, N60, N1540);
xor XOR2 (N1800, N1798, N1450);
buf BUF1 (N1801, N1800);
xor XOR2 (N1802, N1786, N1656);
or OR4 (N1803, N1787, N249, N1090, N688);
nand NAND4 (N1804, N1796, N417, N974, N766);
and AND2 (N1805, N1785, N869);
buf BUF1 (N1806, N1793);
buf BUF1 (N1807, N1803);
or OR4 (N1808, N1794, N253, N1692, N1434);
buf BUF1 (N1809, N1802);
nor NOR2 (N1810, N1804, N552);
and AND2 (N1811, N1808, N1483);
xor XOR2 (N1812, N1809, N1762);
buf BUF1 (N1813, N1807);
xor XOR2 (N1814, N1795, N221);
buf BUF1 (N1815, N1801);
not NOT1 (N1816, N1812);
or OR4 (N1817, N1811, N673, N1394, N1065);
not NOT1 (N1818, N1791);
xor XOR2 (N1819, N1816, N1512);
buf BUF1 (N1820, N1815);
buf BUF1 (N1821, N1799);
buf BUF1 (N1822, N1806);
nand NAND4 (N1823, N1819, N486, N1017, N231);
or OR4 (N1824, N1821, N575, N1687, N1669);
buf BUF1 (N1825, N1813);
and AND3 (N1826, N1822, N449, N245);
buf BUF1 (N1827, N1818);
buf BUF1 (N1828, N1805);
or OR2 (N1829, N1823, N722);
not NOT1 (N1830, N1820);
not NOT1 (N1831, N1810);
xor XOR2 (N1832, N1828, N857);
nor NOR3 (N1833, N1827, N1012, N258);
nand NAND2 (N1834, N1831, N39);
or OR2 (N1835, N1833, N851);
and AND4 (N1836, N1834, N1, N367, N551);
not NOT1 (N1837, N1825);
nor NOR4 (N1838, N1837, N558, N506, N1067);
nor NOR4 (N1839, N1838, N378, N276, N1787);
nand NAND4 (N1840, N1826, N1738, N1335, N743);
and AND4 (N1841, N1830, N309, N1536, N1081);
nand NAND3 (N1842, N1841, N1505, N1017);
xor XOR2 (N1843, N1814, N332);
xor XOR2 (N1844, N1829, N1179);
buf BUF1 (N1845, N1824);
buf BUF1 (N1846, N1836);
nor NOR3 (N1847, N1844, N1671, N1616);
nor NOR3 (N1848, N1845, N459, N1739);
xor XOR2 (N1849, N1839, N1637);
buf BUF1 (N1850, N1843);
or OR2 (N1851, N1850, N489);
not NOT1 (N1852, N1835);
and AND2 (N1853, N1817, N1363);
xor XOR2 (N1854, N1842, N1354);
not NOT1 (N1855, N1851);
buf BUF1 (N1856, N1847);
buf BUF1 (N1857, N1849);
nor NOR2 (N1858, N1856, N1726);
and AND2 (N1859, N1852, N491);
nand NAND2 (N1860, N1853, N1381);
buf BUF1 (N1861, N1832);
and AND2 (N1862, N1854, N272);
or OR4 (N1863, N1860, N1025, N462, N648);
xor XOR2 (N1864, N1840, N1361);
not NOT1 (N1865, N1859);
nand NAND3 (N1866, N1857, N156, N1649);
not NOT1 (N1867, N1861);
buf BUF1 (N1868, N1848);
nor NOR4 (N1869, N1858, N1861, N1277, N357);
and AND4 (N1870, N1862, N708, N290, N412);
not NOT1 (N1871, N1869);
or OR2 (N1872, N1866, N569);
or OR3 (N1873, N1872, N1814, N1228);
xor XOR2 (N1874, N1855, N158);
or OR2 (N1875, N1871, N239);
buf BUF1 (N1876, N1864);
or OR2 (N1877, N1846, N1448);
nand NAND3 (N1878, N1863, N1220, N1599);
and AND3 (N1879, N1870, N1458, N751);
and AND3 (N1880, N1876, N1121, N1793);
buf BUF1 (N1881, N1879);
xor XOR2 (N1882, N1875, N1457);
nor NOR2 (N1883, N1868, N863);
nor NOR2 (N1884, N1865, N1191);
xor XOR2 (N1885, N1883, N334);
nand NAND4 (N1886, N1877, N985, N1788, N1463);
or OR3 (N1887, N1880, N1471, N1700);
and AND3 (N1888, N1873, N1645, N761);
and AND2 (N1889, N1886, N652);
not NOT1 (N1890, N1888);
or OR3 (N1891, N1867, N994, N1506);
xor XOR2 (N1892, N1884, N1232);
not NOT1 (N1893, N1882);
not NOT1 (N1894, N1892);
nor NOR2 (N1895, N1893, N1032);
buf BUF1 (N1896, N1891);
xor XOR2 (N1897, N1889, N154);
or OR4 (N1898, N1874, N501, N1436, N1186);
nor NOR3 (N1899, N1885, N521, N1789);
or OR2 (N1900, N1897, N1297);
xor XOR2 (N1901, N1900, N1247);
and AND3 (N1902, N1898, N1201, N450);
or OR3 (N1903, N1895, N1749, N1517);
buf BUF1 (N1904, N1878);
nand NAND3 (N1905, N1903, N490, N1268);
or OR2 (N1906, N1890, N1733);
xor XOR2 (N1907, N1894, N1322);
buf BUF1 (N1908, N1904);
xor XOR2 (N1909, N1907, N1675);
nor NOR3 (N1910, N1908, N674, N1678);
not NOT1 (N1911, N1896);
nor NOR3 (N1912, N1911, N857, N1109);
not NOT1 (N1913, N1901);
and AND3 (N1914, N1902, N1616, N1463);
not NOT1 (N1915, N1881);
buf BUF1 (N1916, N1914);
buf BUF1 (N1917, N1913);
buf BUF1 (N1918, N1905);
not NOT1 (N1919, N1909);
or OR3 (N1920, N1916, N1415, N1056);
xor XOR2 (N1921, N1899, N1161);
not NOT1 (N1922, N1918);
nand NAND4 (N1923, N1906, N1519, N70, N295);
xor XOR2 (N1924, N1920, N654);
nand NAND3 (N1925, N1910, N1603, N1881);
nor NOR4 (N1926, N1921, N245, N1147, N1053);
xor XOR2 (N1927, N1922, N1614);
not NOT1 (N1928, N1926);
not NOT1 (N1929, N1927);
buf BUF1 (N1930, N1928);
or OR2 (N1931, N1924, N1580);
nand NAND2 (N1932, N1931, N994);
not NOT1 (N1933, N1930);
and AND3 (N1934, N1919, N1043, N393);
xor XOR2 (N1935, N1887, N79);
or OR3 (N1936, N1917, N1124, N1499);
nor NOR2 (N1937, N1934, N1844);
nor NOR3 (N1938, N1937, N1909, N319);
and AND2 (N1939, N1912, N108);
nand NAND3 (N1940, N1933, N370, N627);
nand NAND4 (N1941, N1939, N1573, N1244, N806);
nor NOR2 (N1942, N1941, N1751);
and AND2 (N1943, N1940, N339);
not NOT1 (N1944, N1935);
or OR2 (N1945, N1929, N1151);
or OR4 (N1946, N1944, N302, N1877, N747);
buf BUF1 (N1947, N1938);
and AND3 (N1948, N1946, N1508, N1831);
not NOT1 (N1949, N1936);
nand NAND4 (N1950, N1915, N407, N617, N1408);
buf BUF1 (N1951, N1943);
buf BUF1 (N1952, N1932);
or OR3 (N1953, N1948, N782, N1260);
nor NOR2 (N1954, N1947, N329);
nand NAND3 (N1955, N1923, N511, N1750);
xor XOR2 (N1956, N1925, N1903);
nor NOR2 (N1957, N1953, N485);
buf BUF1 (N1958, N1951);
nand NAND2 (N1959, N1942, N335);
buf BUF1 (N1960, N1957);
and AND4 (N1961, N1959, N1612, N78, N1056);
not NOT1 (N1962, N1961);
and AND2 (N1963, N1958, N1852);
xor XOR2 (N1964, N1962, N951);
not NOT1 (N1965, N1955);
not NOT1 (N1966, N1950);
nand NAND3 (N1967, N1945, N220, N1441);
buf BUF1 (N1968, N1949);
and AND4 (N1969, N1956, N253, N1615, N1036);
not NOT1 (N1970, N1954);
and AND4 (N1971, N1960, N1772, N48, N1204);
nor NOR2 (N1972, N1965, N542);
nor NOR2 (N1973, N1968, N995);
xor XOR2 (N1974, N1967, N873);
buf BUF1 (N1975, N1970);
or OR4 (N1976, N1973, N1144, N326, N1489);
nand NAND4 (N1977, N1966, N1130, N736, N811);
xor XOR2 (N1978, N1969, N1884);
xor XOR2 (N1979, N1974, N1643);
xor XOR2 (N1980, N1964, N236);
nor NOR3 (N1981, N1971, N1626, N410);
and AND3 (N1982, N1976, N991, N1785);
or OR3 (N1983, N1952, N1540, N1288);
nand NAND4 (N1984, N1972, N66, N1659, N1213);
nand NAND3 (N1985, N1975, N364, N1710);
nand NAND2 (N1986, N1985, N442);
nand NAND2 (N1987, N1984, N1669);
or OR2 (N1988, N1978, N1664);
nand NAND4 (N1989, N1982, N1286, N1434, N1321);
not NOT1 (N1990, N1980);
nor NOR2 (N1991, N1983, N96);
or OR4 (N1992, N1990, N726, N451, N1478);
or OR2 (N1993, N1991, N228);
buf BUF1 (N1994, N1987);
nand NAND3 (N1995, N1979, N1254, N72);
and AND4 (N1996, N1986, N478, N129, N508);
nand NAND4 (N1997, N1992, N1083, N1721, N770);
nand NAND2 (N1998, N1993, N1611);
and AND2 (N1999, N1988, N1563);
not NOT1 (N2000, N1998);
nor NOR4 (N2001, N1996, N1544, N1328, N717);
not NOT1 (N2002, N1977);
nor NOR3 (N2003, N1999, N1438, N685);
or OR4 (N2004, N1997, N96, N1584, N1085);
buf BUF1 (N2005, N2000);
buf BUF1 (N2006, N1994);
buf BUF1 (N2007, N2004);
nand NAND3 (N2008, N1963, N1262, N1722);
or OR3 (N2009, N2007, N1981, N1306);
or OR2 (N2010, N530, N1243);
xor XOR2 (N2011, N1989, N1041);
and AND2 (N2012, N2001, N1406);
not NOT1 (N2013, N2009);
not NOT1 (N2014, N2013);
and AND2 (N2015, N2008, N876);
nand NAND2 (N2016, N2010, N1006);
nand NAND4 (N2017, N1995, N588, N368, N1337);
or OR2 (N2018, N2012, N1767);
nor NOR2 (N2019, N2018, N650);
nand NAND2 (N2020, N2006, N958);
xor XOR2 (N2021, N2005, N456);
not NOT1 (N2022, N2017);
xor XOR2 (N2023, N2020, N1334);
or OR3 (N2024, N2014, N1701, N1355);
nand NAND3 (N2025, N2015, N746, N371);
or OR2 (N2026, N2025, N1869);
not NOT1 (N2027, N2023);
not NOT1 (N2028, N2019);
not NOT1 (N2029, N2026);
buf BUF1 (N2030, N2028);
and AND4 (N2031, N2024, N538, N875, N632);
or OR3 (N2032, N2003, N2025, N476);
nand NAND4 (N2033, N2021, N1179, N1536, N1684);
not NOT1 (N2034, N2030);
and AND3 (N2035, N2029, N71, N1142);
not NOT1 (N2036, N2033);
buf BUF1 (N2037, N2002);
nor NOR4 (N2038, N2035, N239, N719, N118);
or OR3 (N2039, N2011, N526, N3);
or OR4 (N2040, N2027, N1450, N1075, N1377);
nand NAND4 (N2041, N2022, N648, N322, N1447);
and AND3 (N2042, N2036, N1206, N1329);
not NOT1 (N2043, N2038);
not NOT1 (N2044, N2016);
and AND3 (N2045, N2042, N600, N655);
nand NAND2 (N2046, N2040, N1779);
xor XOR2 (N2047, N2046, N315);
xor XOR2 (N2048, N2041, N300);
xor XOR2 (N2049, N2045, N421);
nand NAND3 (N2050, N2037, N95, N1444);
or OR2 (N2051, N2049, N449);
xor XOR2 (N2052, N2032, N300);
xor XOR2 (N2053, N2052, N259);
or OR3 (N2054, N2039, N1875, N1729);
nand NAND4 (N2055, N2050, N213, N1108, N81);
not NOT1 (N2056, N2051);
nand NAND4 (N2057, N2047, N319, N1130, N1853);
or OR4 (N2058, N2053, N206, N1625, N1169);
nand NAND4 (N2059, N2044, N1432, N1471, N821);
or OR3 (N2060, N2048, N1048, N809);
or OR2 (N2061, N2034, N1632);
or OR3 (N2062, N2054, N69, N328);
buf BUF1 (N2063, N2057);
buf BUF1 (N2064, N2062);
nor NOR4 (N2065, N2031, N1279, N1105, N247);
xor XOR2 (N2066, N2061, N256);
or OR2 (N2067, N2065, N1334);
and AND2 (N2068, N2064, N1559);
nor NOR4 (N2069, N2058, N1509, N1676, N1270);
or OR2 (N2070, N2069, N1113);
buf BUF1 (N2071, N2060);
nor NOR3 (N2072, N2059, N1323, N267);
nand NAND2 (N2073, N2043, N1145);
nor NOR3 (N2074, N2071, N696, N1386);
not NOT1 (N2075, N2073);
or OR2 (N2076, N2056, N58);
and AND4 (N2077, N2063, N247, N1296, N426);
or OR3 (N2078, N2076, N1239, N1355);
and AND4 (N2079, N2070, N1934, N1366, N793);
not NOT1 (N2080, N2077);
nor NOR2 (N2081, N2055, N1239);
and AND2 (N2082, N2080, N110);
nand NAND2 (N2083, N2079, N1908);
or OR2 (N2084, N2068, N1418);
and AND3 (N2085, N2084, N1673, N521);
xor XOR2 (N2086, N2074, N2073);
nand NAND3 (N2087, N2066, N34, N1311);
nand NAND4 (N2088, N2078, N676, N1169, N1997);
not NOT1 (N2089, N2075);
xor XOR2 (N2090, N2082, N886);
nand NAND2 (N2091, N2072, N604);
and AND3 (N2092, N2088, N1629, N1148);
nand NAND2 (N2093, N2067, N747);
buf BUF1 (N2094, N2083);
and AND4 (N2095, N2081, N1630, N35, N1132);
not NOT1 (N2096, N2095);
and AND2 (N2097, N2091, N1999);
and AND4 (N2098, N2087, N1177, N405, N728);
or OR3 (N2099, N2094, N580, N326);
or OR4 (N2100, N2089, N647, N719, N2017);
nor NOR3 (N2101, N2096, N745, N1342);
buf BUF1 (N2102, N2097);
and AND4 (N2103, N2102, N401, N1618, N250);
xor XOR2 (N2104, N2098, N479);
buf BUF1 (N2105, N2099);
xor XOR2 (N2106, N2090, N619);
buf BUF1 (N2107, N2086);
nand NAND4 (N2108, N2105, N673, N601, N1119);
not NOT1 (N2109, N2092);
nor NOR2 (N2110, N2104, N1700);
and AND3 (N2111, N2085, N1937, N452);
not NOT1 (N2112, N2107);
or OR2 (N2113, N2111, N143);
and AND3 (N2114, N2110, N368, N7);
xor XOR2 (N2115, N2108, N1231);
buf BUF1 (N2116, N2103);
nor NOR2 (N2117, N2114, N42);
or OR4 (N2118, N2117, N762, N800, N1743);
buf BUF1 (N2119, N2116);
nand NAND3 (N2120, N2106, N742, N1113);
or OR4 (N2121, N2100, N1719, N410, N1152);
or OR4 (N2122, N2121, N445, N1695, N1462);
buf BUF1 (N2123, N2119);
buf BUF1 (N2124, N2115);
and AND3 (N2125, N2112, N523, N1185);
nor NOR2 (N2126, N2093, N1028);
buf BUF1 (N2127, N2124);
and AND4 (N2128, N2101, N70, N912, N1619);
buf BUF1 (N2129, N2126);
not NOT1 (N2130, N2125);
or OR4 (N2131, N2120, N1361, N1540, N673);
and AND4 (N2132, N2128, N1804, N1550, N588);
buf BUF1 (N2133, N2129);
nand NAND2 (N2134, N2127, N801);
and AND4 (N2135, N2131, N1006, N1986, N759);
xor XOR2 (N2136, N2118, N1468);
nand NAND2 (N2137, N2136, N1223);
buf BUF1 (N2138, N2113);
xor XOR2 (N2139, N2137, N421);
not NOT1 (N2140, N2133);
nor NOR2 (N2141, N2139, N1024);
and AND2 (N2142, N2122, N809);
or OR4 (N2143, N2142, N1618, N1064, N377);
not NOT1 (N2144, N2130);
nand NAND2 (N2145, N2123, N1876);
xor XOR2 (N2146, N2132, N1645);
and AND4 (N2147, N2140, N2060, N896, N1701);
or OR2 (N2148, N2145, N1120);
xor XOR2 (N2149, N2109, N912);
nand NAND2 (N2150, N2134, N1677);
and AND3 (N2151, N2141, N879, N1877);
nor NOR2 (N2152, N2138, N1453);
buf BUF1 (N2153, N2135);
and AND2 (N2154, N2151, N151);
nor NOR2 (N2155, N2147, N1169);
and AND2 (N2156, N2152, N166);
xor XOR2 (N2157, N2143, N796);
xor XOR2 (N2158, N2146, N1119);
and AND2 (N2159, N2154, N1407);
nor NOR4 (N2160, N2144, N360, N179, N1056);
and AND2 (N2161, N2160, N1974);
not NOT1 (N2162, N2155);
not NOT1 (N2163, N2157);
nor NOR3 (N2164, N2153, N1752, N1696);
xor XOR2 (N2165, N2156, N130);
nand NAND3 (N2166, N2158, N1279, N310);
nand NAND3 (N2167, N2150, N506, N773);
buf BUF1 (N2168, N2161);
and AND4 (N2169, N2165, N111, N898, N1762);
nor NOR3 (N2170, N2162, N38, N82);
and AND2 (N2171, N2148, N1955);
nand NAND2 (N2172, N2171, N536);
xor XOR2 (N2173, N2170, N414);
nor NOR2 (N2174, N2163, N1400);
nor NOR2 (N2175, N2159, N114);
or OR4 (N2176, N2149, N979, N2167, N1682);
and AND2 (N2177, N1425, N518);
buf BUF1 (N2178, N2173);
nand NAND2 (N2179, N2168, N1600);
not NOT1 (N2180, N2169);
nor NOR4 (N2181, N2174, N1167, N1551, N799);
xor XOR2 (N2182, N2176, N754);
nor NOR4 (N2183, N2175, N2148, N288, N447);
or OR2 (N2184, N2178, N1901);
xor XOR2 (N2185, N2182, N808);
and AND3 (N2186, N2184, N543, N1302);
xor XOR2 (N2187, N2183, N1701);
nand NAND2 (N2188, N2179, N2121);
xor XOR2 (N2189, N2166, N1043);
or OR4 (N2190, N2185, N849, N1865, N1909);
nor NOR4 (N2191, N2187, N858, N713, N835);
or OR4 (N2192, N2191, N1818, N1569, N1576);
nand NAND2 (N2193, N2181, N140);
nand NAND3 (N2194, N2189, N1260, N1254);
not NOT1 (N2195, N2188);
or OR2 (N2196, N2195, N1026);
nor NOR2 (N2197, N2192, N739);
not NOT1 (N2198, N2196);
or OR4 (N2199, N2190, N56, N1180, N1433);
and AND4 (N2200, N2186, N620, N1561, N1506);
xor XOR2 (N2201, N2200, N1465);
not NOT1 (N2202, N2197);
and AND2 (N2203, N2198, N1618);
or OR4 (N2204, N2177, N63, N664, N86);
or OR4 (N2205, N2199, N1022, N1719, N1890);
not NOT1 (N2206, N2205);
xor XOR2 (N2207, N2180, N1242);
buf BUF1 (N2208, N2203);
buf BUF1 (N2209, N2201);
and AND2 (N2210, N2164, N424);
xor XOR2 (N2211, N2204, N1366);
nor NOR3 (N2212, N2206, N1105, N771);
nand NAND4 (N2213, N2202, N71, N744, N1743);
not NOT1 (N2214, N2213);
or OR3 (N2215, N2210, N150, N72);
not NOT1 (N2216, N2212);
nand NAND2 (N2217, N2216, N314);
not NOT1 (N2218, N2215);
nor NOR3 (N2219, N2193, N168, N1796);
nand NAND4 (N2220, N2209, N54, N1704, N758);
not NOT1 (N2221, N2218);
not NOT1 (N2222, N2208);
buf BUF1 (N2223, N2194);
nor NOR2 (N2224, N2223, N1974);
nor NOR4 (N2225, N2214, N695, N1832, N1622);
nor NOR3 (N2226, N2211, N1579, N2060);
buf BUF1 (N2227, N2222);
and AND2 (N2228, N2220, N1189);
xor XOR2 (N2229, N2227, N417);
nor NOR2 (N2230, N2217, N1963);
and AND2 (N2231, N2219, N1023);
not NOT1 (N2232, N2231);
and AND3 (N2233, N2224, N410, N1552);
nor NOR3 (N2234, N2221, N854, N931);
nand NAND3 (N2235, N2172, N311, N1718);
or OR4 (N2236, N2225, N389, N1887, N990);
nand NAND4 (N2237, N2207, N421, N2045, N87);
and AND2 (N2238, N2236, N1824);
not NOT1 (N2239, N2238);
not NOT1 (N2240, N2232);
nand NAND2 (N2241, N2226, N654);
xor XOR2 (N2242, N2230, N1845);
xor XOR2 (N2243, N2239, N707);
nand NAND4 (N2244, N2235, N2217, N1448, N267);
xor XOR2 (N2245, N2229, N540);
nand NAND4 (N2246, N2237, N1695, N1299, N116);
xor XOR2 (N2247, N2244, N1059);
not NOT1 (N2248, N2241);
nor NOR2 (N2249, N2247, N1355);
xor XOR2 (N2250, N2243, N952);
and AND2 (N2251, N2250, N1042);
not NOT1 (N2252, N2228);
nand NAND3 (N2253, N2251, N1023, N1032);
nand NAND2 (N2254, N2246, N2136);
xor XOR2 (N2255, N2252, N779);
buf BUF1 (N2256, N2248);
nor NOR2 (N2257, N2234, N1090);
or OR4 (N2258, N2245, N311, N663, N1035);
and AND3 (N2259, N2258, N844, N1059);
nand NAND4 (N2260, N2242, N869, N1398, N610);
and AND3 (N2261, N2254, N327, N1121);
xor XOR2 (N2262, N2255, N1694);
or OR2 (N2263, N2240, N1742);
and AND2 (N2264, N2233, N1004);
or OR4 (N2265, N2249, N1404, N653, N2055);
and AND3 (N2266, N2265, N299, N1011);
or OR4 (N2267, N2257, N840, N1422, N74);
xor XOR2 (N2268, N2256, N120);
and AND4 (N2269, N2253, N2080, N417, N641);
nor NOR2 (N2270, N2268, N1864);
and AND4 (N2271, N2260, N999, N1378, N498);
nand NAND2 (N2272, N2259, N253);
buf BUF1 (N2273, N2262);
nand NAND4 (N2274, N2271, N247, N617, N1745);
nand NAND3 (N2275, N2266, N967, N2193);
not NOT1 (N2276, N2269);
xor XOR2 (N2277, N2264, N1497);
nor NOR4 (N2278, N2275, N844, N852, N1677);
or OR4 (N2279, N2263, N1258, N1490, N2151);
nand NAND4 (N2280, N2272, N225, N2102, N1461);
buf BUF1 (N2281, N2277);
xor XOR2 (N2282, N2278, N1351);
xor XOR2 (N2283, N2281, N1857);
nor NOR4 (N2284, N2274, N257, N346, N1978);
nand NAND4 (N2285, N2282, N66, N1164, N1627);
or OR3 (N2286, N2261, N2223, N1138);
nor NOR4 (N2287, N2280, N45, N801, N1272);
buf BUF1 (N2288, N2267);
buf BUF1 (N2289, N2279);
nand NAND2 (N2290, N2273, N1084);
or OR3 (N2291, N2283, N274, N800);
buf BUF1 (N2292, N2291);
and AND2 (N2293, N2286, N1142);
xor XOR2 (N2294, N2289, N2018);
buf BUF1 (N2295, N2284);
xor XOR2 (N2296, N2287, N752);
buf BUF1 (N2297, N2276);
buf BUF1 (N2298, N2296);
xor XOR2 (N2299, N2285, N1039);
or OR4 (N2300, N2294, N498, N346, N1505);
not NOT1 (N2301, N2288);
buf BUF1 (N2302, N2290);
or OR4 (N2303, N2299, N1486, N1691, N1595);
xor XOR2 (N2304, N2293, N1526);
nand NAND4 (N2305, N2300, N1097, N953, N113);
or OR2 (N2306, N2298, N100);
buf BUF1 (N2307, N2295);
nand NAND4 (N2308, N2307, N850, N1148, N1738);
nand NAND4 (N2309, N2308, N377, N284, N597);
nand NAND2 (N2310, N2302, N1507);
xor XOR2 (N2311, N2297, N1823);
nand NAND4 (N2312, N2310, N1847, N424, N171);
nand NAND2 (N2313, N2303, N109);
and AND3 (N2314, N2270, N90, N651);
and AND4 (N2315, N2305, N1049, N112, N267);
and AND2 (N2316, N2301, N1425);
buf BUF1 (N2317, N2312);
and AND2 (N2318, N2313, N495);
nor NOR3 (N2319, N2311, N1118, N1407);
buf BUF1 (N2320, N2319);
buf BUF1 (N2321, N2318);
xor XOR2 (N2322, N2309, N359);
xor XOR2 (N2323, N2314, N391);
not NOT1 (N2324, N2306);
nand NAND4 (N2325, N2315, N361, N161, N79);
and AND4 (N2326, N2292, N982, N572, N222);
buf BUF1 (N2327, N2325);
or OR3 (N2328, N2324, N629, N427);
nor NOR3 (N2329, N2321, N214, N574);
nor NOR4 (N2330, N2316, N363, N843, N1384);
xor XOR2 (N2331, N2320, N2147);
and AND2 (N2332, N2326, N2044);
nor NOR3 (N2333, N2327, N349, N1831);
xor XOR2 (N2334, N2323, N2241);
not NOT1 (N2335, N2330);
and AND2 (N2336, N2331, N592);
not NOT1 (N2337, N2333);
and AND3 (N2338, N2322, N1743, N1930);
not NOT1 (N2339, N2332);
xor XOR2 (N2340, N2334, N563);
xor XOR2 (N2341, N2338, N1264);
not NOT1 (N2342, N2341);
nand NAND3 (N2343, N2342, N581, N1985);
nor NOR4 (N2344, N2317, N201, N164, N1260);
not NOT1 (N2345, N2344);
or OR2 (N2346, N2345, N204);
xor XOR2 (N2347, N2329, N2114);
nand NAND3 (N2348, N2346, N1482, N1224);
or OR4 (N2349, N2347, N1452, N2261, N439);
not NOT1 (N2350, N2337);
nor NOR3 (N2351, N2350, N2217, N143);
nor NOR2 (N2352, N2336, N1581);
or OR4 (N2353, N2352, N795, N1046, N1238);
nor NOR2 (N2354, N2351, N954);
and AND2 (N2355, N2328, N2211);
or OR2 (N2356, N2355, N1707);
buf BUF1 (N2357, N2304);
nor NOR4 (N2358, N2335, N585, N83, N1827);
xor XOR2 (N2359, N2340, N61);
nand NAND3 (N2360, N2354, N1539, N690);
buf BUF1 (N2361, N2353);
or OR2 (N2362, N2343, N1023);
and AND4 (N2363, N2358, N974, N785, N1213);
nor NOR3 (N2364, N2361, N1169, N2065);
or OR4 (N2365, N2357, N157, N1300, N654);
buf BUF1 (N2366, N2359);
or OR2 (N2367, N2363, N409);
buf BUF1 (N2368, N2349);
and AND2 (N2369, N2365, N1649);
xor XOR2 (N2370, N2368, N915);
not NOT1 (N2371, N2367);
nand NAND4 (N2372, N2339, N1169, N443, N1963);
buf BUF1 (N2373, N2372);
or OR4 (N2374, N2366, N1473, N822, N1528);
or OR4 (N2375, N2370, N376, N778, N2174);
buf BUF1 (N2376, N2374);
nand NAND4 (N2377, N2371, N1241, N19, N879);
buf BUF1 (N2378, N2356);
buf BUF1 (N2379, N2348);
xor XOR2 (N2380, N2377, N917);
buf BUF1 (N2381, N2379);
nor NOR2 (N2382, N2378, N1822);
xor XOR2 (N2383, N2362, N107);
nand NAND3 (N2384, N2375, N1207, N2159);
not NOT1 (N2385, N2380);
or OR3 (N2386, N2383, N553, N344);
and AND2 (N2387, N2381, N1515);
not NOT1 (N2388, N2376);
buf BUF1 (N2389, N2364);
xor XOR2 (N2390, N2373, N1287);
buf BUF1 (N2391, N2386);
or OR3 (N2392, N2390, N1529, N149);
nor NOR2 (N2393, N2385, N408);
and AND2 (N2394, N2392, N962);
xor XOR2 (N2395, N2391, N1645);
xor XOR2 (N2396, N2382, N738);
not NOT1 (N2397, N2396);
nor NOR3 (N2398, N2384, N1032, N277);
and AND4 (N2399, N2393, N1401, N1356, N1341);
buf BUF1 (N2400, N2399);
and AND4 (N2401, N2395, N752, N1178, N997);
not NOT1 (N2402, N2401);
buf BUF1 (N2403, N2397);
not NOT1 (N2404, N2387);
xor XOR2 (N2405, N2360, N745);
xor XOR2 (N2406, N2403, N2357);
xor XOR2 (N2407, N2394, N1263);
not NOT1 (N2408, N2404);
and AND3 (N2409, N2406, N2130, N360);
xor XOR2 (N2410, N2402, N176);
and AND4 (N2411, N2400, N880, N1831, N252);
and AND3 (N2412, N2398, N402, N130);
nand NAND2 (N2413, N2412, N515);
xor XOR2 (N2414, N2369, N1686);
not NOT1 (N2415, N2388);
nand NAND3 (N2416, N2407, N1128, N689);
nor NOR2 (N2417, N2409, N193);
and AND2 (N2418, N2416, N1717);
xor XOR2 (N2419, N2414, N1051);
or OR4 (N2420, N2419, N1578, N1408, N1545);
nand NAND3 (N2421, N2417, N325, N2148);
xor XOR2 (N2422, N2420, N427);
not NOT1 (N2423, N2410);
nand NAND3 (N2424, N2389, N2212, N1380);
buf BUF1 (N2425, N2413);
not NOT1 (N2426, N2411);
xor XOR2 (N2427, N2425, N2077);
buf BUF1 (N2428, N2423);
nand NAND2 (N2429, N2422, N2343);
and AND2 (N2430, N2428, N1230);
nor NOR2 (N2431, N2421, N1559);
buf BUF1 (N2432, N2408);
xor XOR2 (N2433, N2415, N1339);
and AND4 (N2434, N2427, N2157, N950, N491);
nand NAND2 (N2435, N2433, N286);
not NOT1 (N2436, N2431);
xor XOR2 (N2437, N2429, N1787);
xor XOR2 (N2438, N2434, N2369);
nor NOR3 (N2439, N2436, N905, N2027);
and AND3 (N2440, N2439, N309, N1930);
and AND2 (N2441, N2424, N606);
and AND2 (N2442, N2441, N793);
nand NAND2 (N2443, N2426, N498);
not NOT1 (N2444, N2418);
nor NOR2 (N2445, N2435, N1943);
xor XOR2 (N2446, N2444, N217);
nand NAND3 (N2447, N2437, N791, N48);
or OR4 (N2448, N2405, N1190, N141, N1351);
xor XOR2 (N2449, N2448, N1251);
xor XOR2 (N2450, N2440, N828);
and AND4 (N2451, N2447, N945, N850, N1697);
nand NAND2 (N2452, N2443, N2415);
nor NOR2 (N2453, N2450, N1340);
buf BUF1 (N2454, N2430);
buf BUF1 (N2455, N2451);
and AND4 (N2456, N2452, N818, N187, N61);
nor NOR3 (N2457, N2456, N2060, N2242);
nand NAND4 (N2458, N2454, N2406, N2194, N2216);
and AND3 (N2459, N2457, N923, N1562);
not NOT1 (N2460, N2446);
buf BUF1 (N2461, N2459);
buf BUF1 (N2462, N2438);
nor NOR3 (N2463, N2455, N469, N1679);
buf BUF1 (N2464, N2461);
xor XOR2 (N2465, N2445, N119);
buf BUF1 (N2466, N2464);
and AND4 (N2467, N2458, N516, N1301, N302);
nand NAND4 (N2468, N2460, N2202, N32, N2183);
and AND3 (N2469, N2432, N702, N444);
nand NAND4 (N2470, N2465, N1020, N1212, N461);
and AND3 (N2471, N2469, N2455, N1047);
or OR2 (N2472, N2462, N513);
and AND3 (N2473, N2463, N1274, N2416);
xor XOR2 (N2474, N2466, N851);
nand NAND3 (N2475, N2449, N65, N1547);
not NOT1 (N2476, N2471);
buf BUF1 (N2477, N2473);
and AND3 (N2478, N2474, N717, N1978);
nor NOR4 (N2479, N2470, N2047, N1435, N1813);
or OR4 (N2480, N2475, N2174, N1927, N1523);
and AND3 (N2481, N2467, N358, N757);
and AND2 (N2482, N2481, N1940);
nand NAND2 (N2483, N2472, N766);
nand NAND2 (N2484, N2478, N545);
nand NAND4 (N2485, N2480, N574, N2455, N2458);
not NOT1 (N2486, N2453);
or OR4 (N2487, N2477, N637, N1241, N554);
and AND4 (N2488, N2442, N530, N768, N265);
nand NAND2 (N2489, N2476, N1433);
and AND2 (N2490, N2487, N1730);
not NOT1 (N2491, N2483);
buf BUF1 (N2492, N2489);
nor NOR4 (N2493, N2484, N1828, N2154, N801);
or OR2 (N2494, N2491, N2076);
and AND4 (N2495, N2492, N349, N2239, N1036);
or OR3 (N2496, N2493, N58, N1087);
or OR2 (N2497, N2490, N1080);
and AND2 (N2498, N2495, N178);
buf BUF1 (N2499, N2488);
buf BUF1 (N2500, N2499);
buf BUF1 (N2501, N2468);
buf BUF1 (N2502, N2496);
buf BUF1 (N2503, N2500);
nand NAND2 (N2504, N2486, N340);
xor XOR2 (N2505, N2498, N373);
nor NOR2 (N2506, N2494, N1190);
xor XOR2 (N2507, N2502, N889);
buf BUF1 (N2508, N2504);
nand NAND4 (N2509, N2485, N2322, N260, N94);
and AND3 (N2510, N2503, N1838, N657);
buf BUF1 (N2511, N2508);
nand NAND4 (N2512, N2479, N1555, N1831, N1081);
buf BUF1 (N2513, N2482);
not NOT1 (N2514, N2505);
or OR3 (N2515, N2514, N330, N778);
nor NOR2 (N2516, N2501, N787);
and AND4 (N2517, N2511, N2097, N1533, N2429);
endmodule