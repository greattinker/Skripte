// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;

output N312,N300,N309,N295,N301,N305,N311,N310,N288,N313;

or OR3 (N14, N1, N7, N3);
or OR2 (N15, N14, N11);
nand NAND3 (N16, N13, N3, N2);
nand NAND2 (N17, N12, N16);
buf BUF1 (N18, N6);
nand NAND2 (N19, N1, N1);
not NOT1 (N20, N4);
and AND3 (N21, N7, N3, N8);
not NOT1 (N22, N16);
or OR2 (N23, N6, N5);
xor XOR2 (N24, N11, N14);
nand NAND3 (N25, N6, N1, N11);
nand NAND2 (N26, N21, N4);
buf BUF1 (N27, N24);
or OR3 (N28, N27, N18, N3);
buf BUF1 (N29, N28);
nor NOR3 (N30, N9, N21, N8);
xor XOR2 (N31, N30, N1);
not NOT1 (N32, N19);
nand NAND3 (N33, N23, N14, N3);
nor NOR3 (N34, N22, N18, N28);
buf BUF1 (N35, N20);
not NOT1 (N36, N34);
nor NOR4 (N37, N32, N2, N6, N12);
nor NOR3 (N38, N26, N10, N16);
not NOT1 (N39, N17);
nand NAND4 (N40, N38, N2, N35, N9);
nand NAND4 (N41, N31, N13, N3, N26);
buf BUF1 (N42, N26);
not NOT1 (N43, N41);
buf BUF1 (N44, N29);
and AND4 (N45, N25, N26, N29, N44);
and AND2 (N46, N9, N14);
or OR3 (N47, N40, N11, N27);
not NOT1 (N48, N39);
nor NOR4 (N49, N46, N27, N41, N19);
not NOT1 (N50, N48);
or OR4 (N51, N43, N42, N29, N10);
or OR3 (N52, N16, N24, N5);
not NOT1 (N53, N49);
buf BUF1 (N54, N52);
xor XOR2 (N55, N54, N28);
xor XOR2 (N56, N47, N1);
xor XOR2 (N57, N37, N7);
nor NOR4 (N58, N15, N23, N49, N35);
and AND4 (N59, N51, N52, N19, N3);
xor XOR2 (N60, N53, N22);
or OR3 (N61, N33, N4, N11);
nand NAND3 (N62, N56, N54, N61);
xor XOR2 (N63, N26, N34);
and AND2 (N64, N63, N23);
or OR4 (N65, N55, N54, N23, N9);
xor XOR2 (N66, N50, N24);
xor XOR2 (N67, N58, N51);
nand NAND2 (N68, N57, N20);
nand NAND4 (N69, N68, N25, N37, N46);
nor NOR3 (N70, N69, N31, N39);
buf BUF1 (N71, N67);
nor NOR3 (N72, N64, N16, N59);
xor XOR2 (N73, N38, N18);
or OR3 (N74, N66, N5, N1);
nand NAND4 (N75, N71, N30, N33, N54);
buf BUF1 (N76, N70);
nor NOR2 (N77, N75, N9);
nor NOR4 (N78, N77, N13, N55, N29);
or OR3 (N79, N45, N76, N55);
nor NOR3 (N80, N9, N48, N34);
nor NOR2 (N81, N36, N10);
or OR3 (N82, N65, N47, N47);
not NOT1 (N83, N72);
nor NOR2 (N84, N74, N7);
nor NOR3 (N85, N80, N57, N47);
or OR4 (N86, N78, N47, N11, N1);
nor NOR3 (N87, N60, N37, N3);
not NOT1 (N88, N79);
nand NAND2 (N89, N85, N33);
and AND3 (N90, N73, N56, N53);
nand NAND3 (N91, N90, N50, N31);
nand NAND4 (N92, N84, N86, N69, N23);
buf BUF1 (N93, N56);
buf BUF1 (N94, N93);
xor XOR2 (N95, N88, N7);
xor XOR2 (N96, N83, N50);
buf BUF1 (N97, N91);
nand NAND4 (N98, N92, N58, N64, N66);
or OR4 (N99, N98, N96, N18, N15);
nor NOR2 (N100, N69, N81);
and AND3 (N101, N34, N47, N20);
buf BUF1 (N102, N100);
nand NAND3 (N103, N62, N53, N33);
buf BUF1 (N104, N82);
or OR3 (N105, N95, N46, N56);
and AND3 (N106, N102, N103, N16);
buf BUF1 (N107, N21);
xor XOR2 (N108, N105, N99);
xor XOR2 (N109, N1, N51);
not NOT1 (N110, N108);
not NOT1 (N111, N94);
nand NAND2 (N112, N111, N99);
nor NOR3 (N113, N110, N69, N41);
nor NOR2 (N114, N97, N49);
buf BUF1 (N115, N109);
not NOT1 (N116, N101);
nand NAND2 (N117, N104, N31);
nor NOR4 (N118, N89, N103, N98, N27);
buf BUF1 (N119, N107);
nor NOR2 (N120, N114, N69);
or OR2 (N121, N117, N3);
and AND2 (N122, N87, N44);
or OR4 (N123, N121, N112, N49, N28);
not NOT1 (N124, N5);
not NOT1 (N125, N120);
nand NAND4 (N126, N124, N97, N64, N32);
buf BUF1 (N127, N123);
nor NOR4 (N128, N116, N59, N60, N98);
xor XOR2 (N129, N126, N53);
not NOT1 (N130, N125);
and AND4 (N131, N122, N61, N12, N72);
and AND4 (N132, N113, N60, N30, N109);
buf BUF1 (N133, N127);
buf BUF1 (N134, N133);
or OR2 (N135, N128, N35);
xor XOR2 (N136, N130, N89);
xor XOR2 (N137, N135, N89);
nand NAND4 (N138, N136, N73, N10, N115);
xor XOR2 (N139, N135, N14);
or OR4 (N140, N138, N69, N9, N7);
and AND2 (N141, N118, N85);
not NOT1 (N142, N132);
buf BUF1 (N143, N139);
or OR3 (N144, N142, N3, N33);
not NOT1 (N145, N144);
and AND4 (N146, N140, N112, N76, N90);
or OR2 (N147, N137, N142);
nor NOR2 (N148, N143, N35);
and AND4 (N149, N119, N42, N99, N62);
or OR2 (N150, N146, N96);
or OR2 (N151, N147, N24);
nand NAND4 (N152, N149, N113, N21, N132);
not NOT1 (N153, N129);
or OR3 (N154, N152, N126, N74);
not NOT1 (N155, N134);
xor XOR2 (N156, N151, N35);
not NOT1 (N157, N153);
xor XOR2 (N158, N141, N109);
not NOT1 (N159, N155);
nor NOR3 (N160, N148, N52, N112);
xor XOR2 (N161, N150, N138);
or OR3 (N162, N131, N59, N161);
not NOT1 (N163, N152);
nand NAND2 (N164, N163, N114);
or OR2 (N165, N154, N47);
not NOT1 (N166, N159);
not NOT1 (N167, N157);
nor NOR4 (N168, N156, N137, N36, N154);
nor NOR4 (N169, N166, N131, N10, N166);
not NOT1 (N170, N145);
xor XOR2 (N171, N106, N22);
and AND3 (N172, N162, N108, N52);
not NOT1 (N173, N164);
nor NOR2 (N174, N158, N7);
or OR4 (N175, N170, N46, N63, N166);
or OR2 (N176, N169, N42);
and AND3 (N177, N174, N55, N38);
buf BUF1 (N178, N176);
or OR2 (N179, N171, N175);
and AND3 (N180, N112, N42, N75);
or OR4 (N181, N165, N28, N14, N50);
xor XOR2 (N182, N178, N146);
nand NAND2 (N183, N167, N91);
and AND4 (N184, N177, N163, N23, N143);
not NOT1 (N185, N182);
nand NAND3 (N186, N184, N55, N107);
and AND2 (N187, N181, N146);
and AND4 (N188, N160, N47, N70, N113);
nand NAND2 (N189, N172, N63);
not NOT1 (N190, N185);
nand NAND4 (N191, N189, N77, N35, N34);
nor NOR2 (N192, N180, N136);
nor NOR2 (N193, N183, N21);
not NOT1 (N194, N193);
buf BUF1 (N195, N186);
not NOT1 (N196, N194);
not NOT1 (N197, N191);
xor XOR2 (N198, N188, N104);
not NOT1 (N199, N179);
nand NAND2 (N200, N195, N43);
or OR4 (N201, N197, N193, N15, N166);
nand NAND3 (N202, N199, N171, N108);
or OR3 (N203, N196, N5, N174);
xor XOR2 (N204, N173, N1);
buf BUF1 (N205, N168);
and AND2 (N206, N203, N86);
or OR2 (N207, N204, N126);
or OR4 (N208, N201, N167, N137, N127);
nor NOR2 (N209, N187, N33);
buf BUF1 (N210, N208);
nand NAND4 (N211, N192, N37, N111, N53);
xor XOR2 (N212, N207, N189);
not NOT1 (N213, N202);
nor NOR2 (N214, N190, N177);
buf BUF1 (N215, N210);
not NOT1 (N216, N206);
xor XOR2 (N217, N212, N36);
nand NAND2 (N218, N216, N102);
buf BUF1 (N219, N205);
not NOT1 (N220, N198);
nand NAND2 (N221, N211, N63);
buf BUF1 (N222, N200);
and AND2 (N223, N214, N196);
nor NOR2 (N224, N218, N3);
not NOT1 (N225, N213);
and AND3 (N226, N223, N212, N223);
xor XOR2 (N227, N215, N157);
nor NOR2 (N228, N225, N20);
and AND2 (N229, N224, N183);
nand NAND2 (N230, N226, N149);
and AND2 (N231, N230, N59);
or OR2 (N232, N220, N178);
buf BUF1 (N233, N209);
and AND3 (N234, N228, N140, N86);
xor XOR2 (N235, N227, N105);
not NOT1 (N236, N222);
not NOT1 (N237, N232);
not NOT1 (N238, N231);
nor NOR3 (N239, N233, N200, N53);
xor XOR2 (N240, N229, N85);
or OR2 (N241, N238, N94);
or OR2 (N242, N240, N138);
or OR4 (N243, N242, N185, N201, N8);
and AND4 (N244, N236, N201, N194, N110);
nor NOR3 (N245, N221, N239, N220);
xor XOR2 (N246, N64, N154);
nor NOR4 (N247, N234, N51, N195, N119);
or OR4 (N248, N219, N153, N119, N159);
or OR2 (N249, N245, N195);
not NOT1 (N250, N246);
and AND4 (N251, N235, N194, N97, N29);
and AND2 (N252, N249, N211);
nand NAND2 (N253, N250, N211);
or OR4 (N254, N237, N156, N96, N222);
or OR4 (N255, N253, N22, N45, N227);
or OR2 (N256, N252, N132);
nor NOR3 (N257, N247, N51, N164);
nor NOR2 (N258, N241, N189);
or OR2 (N259, N243, N144);
nand NAND3 (N260, N256, N64, N88);
xor XOR2 (N261, N217, N247);
xor XOR2 (N262, N248, N103);
nor NOR3 (N263, N260, N154, N109);
and AND3 (N264, N259, N102, N17);
nand NAND3 (N265, N262, N251, N208);
nor NOR3 (N266, N257, N169, N186);
buf BUF1 (N267, N204);
nand NAND3 (N268, N258, N107, N242);
and AND4 (N269, N261, N251, N88, N76);
nand NAND2 (N270, N269, N208);
xor XOR2 (N271, N255, N145);
nor NOR3 (N272, N254, N117, N180);
nand NAND4 (N273, N272, N4, N69, N94);
and AND4 (N274, N264, N67, N110, N256);
buf BUF1 (N275, N273);
buf BUF1 (N276, N263);
or OR3 (N277, N275, N216, N158);
nor NOR4 (N278, N267, N72, N26, N79);
nand NAND2 (N279, N278, N43);
nor NOR2 (N280, N274, N190);
not NOT1 (N281, N271);
xor XOR2 (N282, N281, N53);
xor XOR2 (N283, N268, N45);
not NOT1 (N284, N283);
buf BUF1 (N285, N282);
buf BUF1 (N286, N279);
or OR2 (N287, N265, N50);
nand NAND3 (N288, N284, N237, N256);
xor XOR2 (N289, N287, N76);
xor XOR2 (N290, N266, N220);
not NOT1 (N291, N244);
not NOT1 (N292, N289);
or OR2 (N293, N276, N138);
and AND3 (N294, N277, N273, N222);
nand NAND4 (N295, N294, N159, N89, N91);
not NOT1 (N296, N292);
nor NOR4 (N297, N280, N1, N24, N296);
and AND2 (N298, N7, N272);
buf BUF1 (N299, N286);
xor XOR2 (N300, N297, N263);
xor XOR2 (N301, N285, N238);
xor XOR2 (N302, N298, N278);
or OR4 (N303, N293, N11, N181, N33);
not NOT1 (N304, N303);
nor NOR2 (N305, N299, N111);
buf BUF1 (N306, N270);
or OR4 (N307, N304, N283, N185, N154);
nand NAND3 (N308, N306, N67, N21);
or OR2 (N309, N291, N281);
or OR2 (N310, N302, N53);
or OR3 (N311, N307, N308, N7);
nand NAND2 (N312, N33, N86);
not NOT1 (N313, N290);
endmodule