// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N514,N504,N509,N515,N510,N513,N505,N512,N516,N517;

nor NOR4 (N18, N9, N12, N4, N17);
or OR3 (N19, N8, N5, N8);
or OR2 (N20, N8, N17);
nand NAND3 (N21, N10, N7, N1);
or OR3 (N22, N9, N21, N9);
not NOT1 (N23, N12);
and AND4 (N24, N4, N14, N18, N19);
xor XOR2 (N25, N6, N11);
and AND3 (N26, N9, N22, N13);
nand NAND2 (N27, N23, N26);
and AND4 (N28, N18, N9, N14, N6);
xor XOR2 (N29, N4, N20);
buf BUF1 (N30, N28);
and AND2 (N31, N15, N10);
nand NAND2 (N32, N26, N28);
and AND4 (N33, N2, N2, N21, N20);
not NOT1 (N34, N5);
nand NAND4 (N35, N27, N32, N20, N20);
and AND3 (N36, N13, N20, N6);
nor NOR3 (N37, N29, N21, N8);
xor XOR2 (N38, N28, N31);
xor XOR2 (N39, N9, N13);
and AND2 (N40, N25, N39);
not NOT1 (N41, N25);
nor NOR2 (N42, N24, N28);
buf BUF1 (N43, N37);
nand NAND2 (N44, N42, N11);
or OR3 (N45, N41, N24, N8);
nand NAND3 (N46, N44, N28, N24);
or OR4 (N47, N38, N5, N7, N27);
xor XOR2 (N48, N35, N14);
buf BUF1 (N49, N30);
nand NAND2 (N50, N46, N46);
xor XOR2 (N51, N33, N28);
or OR3 (N52, N36, N26, N12);
not NOT1 (N53, N50);
nor NOR4 (N54, N53, N17, N23, N14);
or OR3 (N55, N52, N33, N4);
or OR2 (N56, N55, N43);
and AND2 (N57, N43, N34);
buf BUF1 (N58, N57);
nor NOR4 (N59, N6, N12, N8, N10);
and AND4 (N60, N54, N28, N28, N23);
nand NAND3 (N61, N45, N29, N38);
not NOT1 (N62, N40);
or OR3 (N63, N48, N24, N4);
xor XOR2 (N64, N56, N52);
and AND2 (N65, N59, N47);
nor NOR2 (N66, N48, N59);
nand NAND4 (N67, N66, N13, N50, N20);
nor NOR3 (N68, N60, N26, N21);
xor XOR2 (N69, N58, N30);
nand NAND3 (N70, N62, N33, N41);
and AND4 (N71, N67, N49, N6, N26);
buf BUF1 (N72, N8);
buf BUF1 (N73, N65);
xor XOR2 (N74, N70, N25);
and AND4 (N75, N61, N23, N25, N32);
buf BUF1 (N76, N63);
nand NAND3 (N77, N69, N13, N33);
or OR4 (N78, N64, N73, N65, N57);
nand NAND4 (N79, N10, N15, N68, N54);
not NOT1 (N80, N37);
xor XOR2 (N81, N75, N22);
nor NOR4 (N82, N79, N11, N1, N17);
or OR3 (N83, N76, N3, N82);
xor XOR2 (N84, N66, N27);
xor XOR2 (N85, N74, N7);
nand NAND2 (N86, N83, N54);
nor NOR4 (N87, N85, N63, N24, N84);
nand NAND4 (N88, N12, N4, N6, N70);
not NOT1 (N89, N88);
not NOT1 (N90, N78);
nor NOR4 (N91, N81, N38, N29, N84);
not NOT1 (N92, N71);
and AND4 (N93, N89, N26, N86, N49);
buf BUF1 (N94, N4);
or OR4 (N95, N72, N85, N44, N47);
xor XOR2 (N96, N91, N59);
or OR3 (N97, N87, N19, N25);
buf BUF1 (N98, N80);
and AND4 (N99, N90, N42, N62, N49);
not NOT1 (N100, N93);
not NOT1 (N101, N51);
and AND4 (N102, N100, N37, N52, N29);
nor NOR2 (N103, N96, N83);
nor NOR3 (N104, N99, N72, N79);
and AND2 (N105, N98, N1);
nor NOR4 (N106, N92, N50, N80, N28);
nand NAND3 (N107, N101, N85, N56);
nand NAND4 (N108, N105, N15, N61, N44);
nor NOR2 (N109, N107, N51);
xor XOR2 (N110, N109, N83);
nand NAND4 (N111, N97, N100, N32, N101);
xor XOR2 (N112, N111, N76);
nor NOR2 (N113, N77, N63);
and AND2 (N114, N112, N99);
nor NOR4 (N115, N104, N83, N66, N10);
not NOT1 (N116, N108);
buf BUF1 (N117, N115);
or OR3 (N118, N94, N16, N24);
not NOT1 (N119, N106);
buf BUF1 (N120, N103);
not NOT1 (N121, N116);
xor XOR2 (N122, N117, N117);
nand NAND2 (N123, N110, N22);
or OR2 (N124, N95, N12);
and AND3 (N125, N102, N83, N22);
and AND4 (N126, N119, N17, N43, N20);
nand NAND4 (N127, N125, N9, N2, N74);
or OR2 (N128, N124, N88);
or OR2 (N129, N118, N60);
and AND4 (N130, N126, N48, N126, N98);
xor XOR2 (N131, N122, N44);
buf BUF1 (N132, N128);
nand NAND2 (N133, N132, N91);
xor XOR2 (N134, N113, N56);
xor XOR2 (N135, N123, N94);
nand NAND4 (N136, N133, N97, N89, N6);
nor NOR3 (N137, N136, N2, N133);
not NOT1 (N138, N134);
and AND3 (N139, N131, N107, N69);
xor XOR2 (N140, N127, N34);
nand NAND2 (N141, N121, N44);
buf BUF1 (N142, N135);
xor XOR2 (N143, N139, N46);
or OR4 (N144, N129, N135, N93, N54);
and AND2 (N145, N138, N139);
or OR2 (N146, N130, N27);
nor NOR3 (N147, N146, N2, N123);
or OR2 (N148, N143, N61);
xor XOR2 (N149, N144, N80);
buf BUF1 (N150, N149);
buf BUF1 (N151, N147);
nor NOR3 (N152, N148, N91, N50);
xor XOR2 (N153, N140, N139);
and AND2 (N154, N145, N83);
not NOT1 (N155, N151);
not NOT1 (N156, N137);
not NOT1 (N157, N155);
nand NAND2 (N158, N153, N36);
nand NAND2 (N159, N152, N63);
and AND2 (N160, N159, N23);
not NOT1 (N161, N158);
and AND4 (N162, N142, N45, N127, N68);
nor NOR2 (N163, N162, N83);
xor XOR2 (N164, N156, N37);
or OR3 (N165, N161, N125, N14);
nand NAND2 (N166, N163, N71);
and AND2 (N167, N154, N11);
xor XOR2 (N168, N164, N151);
not NOT1 (N169, N120);
nor NOR3 (N170, N165, N102, N114);
buf BUF1 (N171, N13);
xor XOR2 (N172, N157, N84);
buf BUF1 (N173, N160);
buf BUF1 (N174, N150);
or OR3 (N175, N166, N31, N5);
nand NAND3 (N176, N167, N129, N36);
xor XOR2 (N177, N173, N77);
xor XOR2 (N178, N174, N149);
and AND2 (N179, N177, N25);
and AND4 (N180, N178, N156, N56, N169);
buf BUF1 (N181, N169);
buf BUF1 (N182, N180);
nand NAND2 (N183, N179, N4);
buf BUF1 (N184, N141);
and AND3 (N185, N183, N144, N77);
not NOT1 (N186, N176);
buf BUF1 (N187, N181);
and AND4 (N188, N170, N118, N69, N61);
or OR2 (N189, N175, N175);
buf BUF1 (N190, N185);
or OR4 (N191, N172, N183, N74, N137);
nand NAND3 (N192, N182, N185, N55);
buf BUF1 (N193, N184);
not NOT1 (N194, N186);
nand NAND4 (N195, N187, N122, N104, N145);
and AND4 (N196, N194, N26, N158, N175);
and AND4 (N197, N192, N160, N161, N178);
and AND3 (N198, N190, N103, N96);
nor NOR2 (N199, N189, N130);
and AND4 (N200, N168, N126, N94, N13);
not NOT1 (N201, N171);
xor XOR2 (N202, N200, N102);
and AND3 (N203, N202, N164, N92);
not NOT1 (N204, N198);
xor XOR2 (N205, N193, N3);
nor NOR4 (N206, N201, N93, N88, N89);
nand NAND4 (N207, N188, N159, N44, N75);
buf BUF1 (N208, N206);
or OR3 (N209, N207, N27, N99);
buf BUF1 (N210, N208);
and AND3 (N211, N196, N120, N16);
or OR2 (N212, N205, N12);
not NOT1 (N213, N210);
nor NOR4 (N214, N213, N138, N167, N9);
and AND2 (N215, N214, N150);
nand NAND4 (N216, N204, N164, N79, N91);
and AND2 (N217, N195, N44);
nand NAND4 (N218, N211, N13, N99, N29);
or OR3 (N219, N218, N63, N157);
or OR4 (N220, N203, N116, N5, N6);
not NOT1 (N221, N215);
or OR2 (N222, N216, N194);
or OR2 (N223, N220, N158);
and AND4 (N224, N212, N102, N166, N44);
or OR4 (N225, N224, N209, N43, N118);
buf BUF1 (N226, N181);
not NOT1 (N227, N197);
nor NOR2 (N228, N199, N7);
xor XOR2 (N229, N221, N182);
xor XOR2 (N230, N229, N146);
buf BUF1 (N231, N227);
nand NAND2 (N232, N231, N31);
nand NAND2 (N233, N230, N172);
nand NAND3 (N234, N191, N31, N166);
nand NAND2 (N235, N232, N128);
nand NAND2 (N236, N228, N47);
buf BUF1 (N237, N223);
nor NOR4 (N238, N225, N3, N107, N154);
buf BUF1 (N239, N222);
nand NAND4 (N240, N238, N43, N124, N22);
nand NAND2 (N241, N237, N103);
xor XOR2 (N242, N240, N99);
and AND2 (N243, N219, N65);
nand NAND4 (N244, N236, N227, N237, N20);
or OR4 (N245, N226, N38, N48, N148);
not NOT1 (N246, N241);
nor NOR3 (N247, N244, N204, N190);
and AND2 (N248, N235, N31);
nand NAND2 (N249, N246, N42);
buf BUF1 (N250, N245);
nand NAND2 (N251, N217, N125);
or OR3 (N252, N249, N216, N94);
and AND4 (N253, N243, N113, N127, N133);
not NOT1 (N254, N252);
buf BUF1 (N255, N251);
nand NAND3 (N256, N253, N43, N77);
nor NOR4 (N257, N233, N82, N18, N65);
and AND3 (N258, N247, N82, N159);
not NOT1 (N259, N250);
nand NAND3 (N260, N259, N160, N52);
nor NOR4 (N261, N258, N195, N84, N74);
and AND2 (N262, N242, N228);
buf BUF1 (N263, N257);
nor NOR3 (N264, N260, N39, N217);
buf BUF1 (N265, N264);
and AND4 (N266, N254, N249, N205, N87);
not NOT1 (N267, N261);
nor NOR2 (N268, N265, N7);
buf BUF1 (N269, N266);
not NOT1 (N270, N268);
buf BUF1 (N271, N255);
and AND3 (N272, N270, N1, N232);
nand NAND2 (N273, N263, N103);
buf BUF1 (N274, N272);
buf BUF1 (N275, N269);
or OR4 (N276, N256, N33, N169, N23);
or OR2 (N277, N273, N121);
and AND4 (N278, N271, N260, N141, N252);
nor NOR3 (N279, N234, N158, N61);
not NOT1 (N280, N267);
and AND4 (N281, N274, N223, N143, N11);
xor XOR2 (N282, N262, N168);
and AND4 (N283, N239, N276, N191, N107);
nor NOR2 (N284, N211, N77);
nand NAND2 (N285, N282, N150);
xor XOR2 (N286, N281, N267);
not NOT1 (N287, N283);
not NOT1 (N288, N280);
not NOT1 (N289, N278);
not NOT1 (N290, N288);
nor NOR2 (N291, N284, N5);
nor NOR3 (N292, N279, N127, N252);
not NOT1 (N293, N248);
buf BUF1 (N294, N293);
xor XOR2 (N295, N294, N238);
buf BUF1 (N296, N275);
and AND2 (N297, N290, N178);
buf BUF1 (N298, N296);
buf BUF1 (N299, N285);
and AND4 (N300, N287, N91, N203, N232);
or OR4 (N301, N300, N267, N179, N283);
xor XOR2 (N302, N297, N206);
and AND3 (N303, N291, N162, N52);
or OR2 (N304, N277, N165);
nor NOR2 (N305, N303, N121);
nor NOR2 (N306, N292, N213);
buf BUF1 (N307, N286);
not NOT1 (N308, N304);
xor XOR2 (N309, N302, N59);
not NOT1 (N310, N308);
xor XOR2 (N311, N306, N100);
xor XOR2 (N312, N289, N253);
or OR3 (N313, N311, N171, N154);
xor XOR2 (N314, N298, N254);
and AND3 (N315, N312, N177, N252);
and AND4 (N316, N309, N54, N94, N182);
buf BUF1 (N317, N316);
not NOT1 (N318, N317);
buf BUF1 (N319, N295);
buf BUF1 (N320, N319);
nor NOR3 (N321, N310, N54, N229);
and AND3 (N322, N321, N291, N250);
not NOT1 (N323, N301);
nand NAND3 (N324, N299, N92, N37);
xor XOR2 (N325, N318, N234);
or OR2 (N326, N322, N148);
and AND4 (N327, N314, N130, N168, N87);
nand NAND3 (N328, N323, N229, N285);
buf BUF1 (N329, N326);
buf BUF1 (N330, N313);
and AND3 (N331, N315, N70, N234);
xor XOR2 (N332, N328, N94);
nor NOR2 (N333, N305, N250);
nor NOR4 (N334, N320, N250, N194, N312);
buf BUF1 (N335, N333);
buf BUF1 (N336, N331);
or OR2 (N337, N336, N232);
and AND2 (N338, N325, N159);
not NOT1 (N339, N307);
nand NAND4 (N340, N330, N219, N260, N140);
or OR3 (N341, N332, N290, N86);
or OR3 (N342, N340, N288, N118);
nand NAND3 (N343, N341, N313, N234);
and AND2 (N344, N327, N339);
nor NOR2 (N345, N57, N289);
and AND2 (N346, N343, N246);
nor NOR4 (N347, N335, N335, N159, N24);
nor NOR4 (N348, N342, N109, N129, N162);
buf BUF1 (N349, N345);
or OR2 (N350, N338, N304);
nand NAND2 (N351, N349, N343);
xor XOR2 (N352, N324, N79);
and AND2 (N353, N344, N227);
nand NAND3 (N354, N337, N64, N95);
nand NAND2 (N355, N352, N259);
and AND2 (N356, N354, N252);
not NOT1 (N357, N350);
buf BUF1 (N358, N334);
xor XOR2 (N359, N347, N289);
xor XOR2 (N360, N329, N294);
nor NOR3 (N361, N348, N190, N168);
not NOT1 (N362, N351);
and AND3 (N363, N361, N15, N48);
not NOT1 (N364, N358);
nand NAND3 (N365, N364, N88, N141);
or OR4 (N366, N357, N202, N3, N209);
not NOT1 (N367, N365);
nand NAND3 (N368, N360, N83, N326);
not NOT1 (N369, N359);
buf BUF1 (N370, N363);
nor NOR4 (N371, N366, N11, N209, N48);
not NOT1 (N372, N346);
nor NOR3 (N373, N368, N167, N37);
nand NAND4 (N374, N371, N243, N125, N356);
or OR4 (N375, N2, N137, N251, N148);
not NOT1 (N376, N367);
xor XOR2 (N377, N375, N79);
and AND2 (N378, N362, N136);
nand NAND4 (N379, N355, N256, N54, N204);
xor XOR2 (N380, N370, N305);
xor XOR2 (N381, N376, N76);
and AND2 (N382, N377, N335);
nor NOR2 (N383, N369, N144);
xor XOR2 (N384, N372, N165);
buf BUF1 (N385, N373);
and AND2 (N386, N378, N30);
or OR4 (N387, N385, N350, N123, N247);
and AND4 (N388, N384, N212, N39, N294);
nand NAND3 (N389, N382, N118, N206);
or OR2 (N390, N381, N322);
and AND3 (N391, N390, N215, N304);
nand NAND2 (N392, N391, N266);
or OR2 (N393, N388, N212);
and AND3 (N394, N387, N235, N172);
xor XOR2 (N395, N392, N328);
nand NAND2 (N396, N374, N235);
or OR4 (N397, N396, N119, N353, N300);
nor NOR2 (N398, N139, N14);
not NOT1 (N399, N395);
xor XOR2 (N400, N386, N132);
nor NOR3 (N401, N393, N33, N39);
nor NOR4 (N402, N379, N53, N117, N36);
nor NOR2 (N403, N389, N153);
or OR4 (N404, N401, N15, N340, N176);
not NOT1 (N405, N398);
or OR3 (N406, N399, N166, N145);
buf BUF1 (N407, N405);
or OR4 (N408, N404, N407, N346, N47);
buf BUF1 (N409, N229);
not NOT1 (N410, N406);
nor NOR3 (N411, N400, N298, N136);
or OR2 (N412, N383, N191);
buf BUF1 (N413, N411);
not NOT1 (N414, N408);
or OR3 (N415, N413, N99, N25);
nor NOR4 (N416, N380, N377, N390, N132);
nand NAND3 (N417, N397, N73, N99);
nor NOR3 (N418, N410, N97, N162);
and AND3 (N419, N402, N244, N6);
xor XOR2 (N420, N415, N290);
or OR4 (N421, N420, N324, N285, N265);
and AND4 (N422, N419, N101, N167, N182);
not NOT1 (N423, N421);
and AND3 (N424, N409, N204, N247);
buf BUF1 (N425, N423);
and AND4 (N426, N418, N374, N145, N31);
nand NAND4 (N427, N394, N368, N264, N156);
or OR4 (N428, N422, N9, N386, N195);
buf BUF1 (N429, N426);
buf BUF1 (N430, N416);
xor XOR2 (N431, N414, N72);
not NOT1 (N432, N424);
and AND4 (N433, N427, N278, N152, N353);
and AND3 (N434, N417, N402, N292);
nand NAND2 (N435, N434, N57);
or OR4 (N436, N435, N183, N266, N341);
buf BUF1 (N437, N425);
and AND4 (N438, N431, N206, N395, N198);
not NOT1 (N439, N437);
buf BUF1 (N440, N438);
not NOT1 (N441, N412);
or OR4 (N442, N440, N199, N201, N57);
or OR3 (N443, N428, N43, N24);
xor XOR2 (N444, N430, N157);
xor XOR2 (N445, N433, N296);
buf BUF1 (N446, N403);
nor NOR2 (N447, N443, N110);
or OR3 (N448, N432, N185, N22);
and AND2 (N449, N445, N9);
nor NOR3 (N450, N449, N394, N66);
or OR2 (N451, N429, N382);
nand NAND2 (N452, N451, N29);
or OR2 (N453, N446, N130);
and AND4 (N454, N448, N192, N250, N427);
nor NOR4 (N455, N439, N21, N156, N315);
nor NOR2 (N456, N444, N405);
nand NAND3 (N457, N447, N218, N405);
xor XOR2 (N458, N442, N251);
or OR2 (N459, N441, N256);
nor NOR2 (N460, N458, N114);
or OR2 (N461, N457, N381);
xor XOR2 (N462, N450, N61);
not NOT1 (N463, N436);
nand NAND2 (N464, N461, N447);
and AND4 (N465, N452, N348, N343, N386);
buf BUF1 (N466, N456);
xor XOR2 (N467, N463, N256);
nor NOR2 (N468, N465, N389);
not NOT1 (N469, N467);
not NOT1 (N470, N464);
buf BUF1 (N471, N454);
nand NAND3 (N472, N470, N166, N50);
nor NOR2 (N473, N466, N260);
buf BUF1 (N474, N459);
nand NAND4 (N475, N462, N167, N172, N212);
nor NOR3 (N476, N472, N441, N429);
not NOT1 (N477, N453);
and AND4 (N478, N455, N304, N390, N400);
nor NOR4 (N479, N478, N245, N179, N306);
not NOT1 (N480, N460);
buf BUF1 (N481, N474);
nor NOR2 (N482, N468, N15);
buf BUF1 (N483, N480);
and AND2 (N484, N482, N5);
or OR2 (N485, N469, N263);
and AND2 (N486, N473, N6);
buf BUF1 (N487, N477);
and AND4 (N488, N485, N220, N266, N367);
xor XOR2 (N489, N481, N163);
or OR3 (N490, N488, N213, N65);
and AND3 (N491, N476, N306, N187);
and AND3 (N492, N491, N138, N51);
xor XOR2 (N493, N490, N467);
and AND3 (N494, N487, N256, N122);
not NOT1 (N495, N475);
and AND4 (N496, N483, N421, N491, N111);
xor XOR2 (N497, N493, N306);
not NOT1 (N498, N486);
nand NAND4 (N499, N494, N233, N383, N316);
and AND2 (N500, N492, N97);
nand NAND2 (N501, N479, N401);
buf BUF1 (N502, N484);
nand NAND2 (N503, N502, N416);
nand NAND2 (N504, N503, N287);
and AND3 (N505, N501, N271, N297);
nor NOR3 (N506, N500, N484, N56);
not NOT1 (N507, N506);
or OR4 (N508, N471, N340, N282, N182);
not NOT1 (N509, N508);
not NOT1 (N510, N498);
buf BUF1 (N511, N489);
or OR4 (N512, N497, N275, N307, N179);
buf BUF1 (N513, N495);
nor NOR3 (N514, N496, N342, N270);
nor NOR4 (N515, N511, N371, N347, N21);
not NOT1 (N516, N499);
xor XOR2 (N517, N507, N63);
endmodule