// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N990,N1012,N1004,N1000,N1006,N1011,N1010,N1013,N980,N1015;

and AND4 (N16, N6, N3, N6, N5);
xor XOR2 (N17, N7, N4);
nand NAND3 (N18, N15, N6, N1);
xor XOR2 (N19, N14, N4);
or OR4 (N20, N16, N7, N8, N17);
buf BUF1 (N21, N16);
nor NOR3 (N22, N8, N19, N3);
nor NOR2 (N23, N13, N9);
or OR2 (N24, N11, N15);
buf BUF1 (N25, N16);
not NOT1 (N26, N19);
nand NAND2 (N27, N25, N17);
or OR4 (N28, N15, N16, N20, N10);
or OR3 (N29, N8, N26, N7);
nor NOR4 (N30, N7, N18, N16, N7);
or OR4 (N31, N27, N12, N9, N7);
buf BUF1 (N32, N4);
xor XOR2 (N33, N5, N32);
or OR3 (N34, N22, N28, N5);
xor XOR2 (N35, N28, N18);
xor XOR2 (N36, N25, N23);
or OR2 (N37, N12, N30);
not NOT1 (N38, N26);
buf BUF1 (N39, N24);
buf BUF1 (N40, N31);
nor NOR4 (N41, N21, N35, N29, N38);
and AND2 (N42, N31, N4);
or OR3 (N43, N16, N39, N41);
nor NOR4 (N44, N19, N15, N3, N30);
or OR4 (N45, N10, N4, N10, N9);
not NOT1 (N46, N16);
nand NAND4 (N47, N37, N24, N29, N37);
buf BUF1 (N48, N46);
and AND2 (N49, N36, N33);
buf BUF1 (N50, N1);
or OR4 (N51, N43, N33, N11, N9);
buf BUF1 (N52, N40);
xor XOR2 (N53, N45, N13);
and AND2 (N54, N53, N35);
or OR4 (N55, N47, N16, N37, N12);
buf BUF1 (N56, N51);
not NOT1 (N57, N52);
nor NOR4 (N58, N54, N30, N25, N23);
xor XOR2 (N59, N55, N45);
and AND4 (N60, N56, N6, N51, N11);
not NOT1 (N61, N60);
not NOT1 (N62, N48);
not NOT1 (N63, N49);
buf BUF1 (N64, N58);
and AND3 (N65, N62, N15, N63);
or OR4 (N66, N60, N51, N30, N22);
nor NOR4 (N67, N66, N34, N59, N59);
and AND4 (N68, N35, N44, N9, N22);
buf BUF1 (N69, N32);
not NOT1 (N70, N25);
not NOT1 (N71, N65);
and AND4 (N72, N68, N3, N30, N32);
nand NAND4 (N73, N70, N13, N19, N38);
xor XOR2 (N74, N42, N14);
or OR2 (N75, N57, N29);
and AND2 (N76, N75, N61);
or OR4 (N77, N57, N42, N39, N54);
nor NOR2 (N78, N73, N12);
nand NAND2 (N79, N77, N78);
or OR3 (N80, N31, N45, N8);
or OR3 (N81, N76, N60, N62);
not NOT1 (N82, N69);
buf BUF1 (N83, N71);
and AND2 (N84, N74, N31);
nor NOR3 (N85, N84, N72, N18);
xor XOR2 (N86, N78, N81);
buf BUF1 (N87, N19);
or OR3 (N88, N50, N17, N13);
and AND3 (N89, N88, N51, N24);
nor NOR3 (N90, N79, N88, N86);
nand NAND4 (N91, N13, N50, N8, N19);
nor NOR4 (N92, N82, N69, N3, N50);
buf BUF1 (N93, N87);
or OR3 (N94, N93, N29, N89);
and AND3 (N95, N16, N67, N55);
nand NAND4 (N96, N17, N28, N12, N26);
or OR4 (N97, N92, N90, N94, N59);
nand NAND4 (N98, N45, N57, N93, N96);
and AND2 (N99, N27, N62);
nor NOR4 (N100, N3, N75, N66, N44);
and AND4 (N101, N85, N44, N74, N5);
or OR2 (N102, N91, N6);
buf BUF1 (N103, N99);
or OR4 (N104, N101, N14, N80, N50);
and AND4 (N105, N25, N94, N22, N45);
buf BUF1 (N106, N100);
and AND4 (N107, N106, N31, N22, N76);
buf BUF1 (N108, N102);
not NOT1 (N109, N83);
nand NAND4 (N110, N98, N79, N91, N85);
not NOT1 (N111, N104);
buf BUF1 (N112, N110);
not NOT1 (N113, N107);
or OR2 (N114, N95, N23);
nand NAND2 (N115, N109, N80);
nand NAND3 (N116, N105, N92, N5);
nand NAND4 (N117, N116, N116, N23, N116);
not NOT1 (N118, N112);
and AND4 (N119, N113, N65, N114, N55);
or OR2 (N120, N118, N76);
buf BUF1 (N121, N109);
or OR3 (N122, N111, N93, N28);
buf BUF1 (N123, N64);
or OR3 (N124, N120, N13, N3);
and AND2 (N125, N119, N102);
nor NOR2 (N126, N122, N81);
nor NOR3 (N127, N123, N123, N53);
and AND4 (N128, N121, N105, N49, N102);
buf BUF1 (N129, N115);
buf BUF1 (N130, N125);
not NOT1 (N131, N128);
or OR3 (N132, N117, N9, N1);
buf BUF1 (N133, N132);
nor NOR3 (N134, N126, N47, N77);
buf BUF1 (N135, N108);
nor NOR2 (N136, N135, N79);
or OR2 (N137, N129, N15);
nor NOR4 (N138, N133, N99, N126, N105);
nand NAND3 (N139, N136, N85, N6);
and AND4 (N140, N137, N12, N71, N82);
xor XOR2 (N141, N134, N8);
not NOT1 (N142, N103);
or OR3 (N143, N97, N5, N2);
nor NOR4 (N144, N140, N126, N52, N61);
nand NAND3 (N145, N139, N83, N141);
not NOT1 (N146, N37);
nand NAND2 (N147, N145, N30);
nor NOR3 (N148, N138, N65, N113);
and AND2 (N149, N147, N111);
nor NOR2 (N150, N143, N44);
not NOT1 (N151, N142);
nand NAND2 (N152, N144, N26);
xor XOR2 (N153, N124, N111);
nor NOR3 (N154, N153, N9, N95);
nand NAND3 (N155, N131, N10, N56);
nor NOR4 (N156, N154, N83, N109, N67);
nor NOR2 (N157, N146, N20);
nor NOR2 (N158, N148, N134);
xor XOR2 (N159, N149, N60);
not NOT1 (N160, N155);
or OR4 (N161, N151, N84, N68, N5);
and AND4 (N162, N152, N102, N81, N99);
or OR3 (N163, N159, N57, N108);
not NOT1 (N164, N127);
not NOT1 (N165, N164);
nand NAND2 (N166, N157, N20);
nor NOR4 (N167, N165, N70, N93, N46);
nand NAND4 (N168, N167, N78, N77, N65);
nand NAND2 (N169, N160, N49);
nor NOR4 (N170, N169, N129, N60, N13);
buf BUF1 (N171, N156);
and AND3 (N172, N166, N73, N80);
not NOT1 (N173, N150);
or OR2 (N174, N172, N117);
buf BUF1 (N175, N161);
xor XOR2 (N176, N173, N71);
nor NOR2 (N177, N174, N11);
nand NAND2 (N178, N130, N115);
nor NOR2 (N179, N170, N126);
nand NAND4 (N180, N177, N76, N35, N94);
xor XOR2 (N181, N175, N47);
or OR2 (N182, N162, N114);
nand NAND4 (N183, N181, N135, N138, N6);
xor XOR2 (N184, N168, N116);
or OR4 (N185, N176, N42, N100, N45);
buf BUF1 (N186, N179);
or OR4 (N187, N183, N107, N61, N171);
or OR3 (N188, N84, N110, N171);
buf BUF1 (N189, N178);
not NOT1 (N190, N180);
and AND4 (N191, N182, N46, N143, N37);
nor NOR2 (N192, N186, N59);
and AND2 (N193, N191, N27);
nor NOR3 (N194, N184, N114, N108);
or OR4 (N195, N189, N40, N126, N127);
xor XOR2 (N196, N187, N50);
or OR3 (N197, N158, N22, N68);
xor XOR2 (N198, N185, N92);
buf BUF1 (N199, N163);
xor XOR2 (N200, N193, N71);
and AND3 (N201, N190, N4, N15);
nor NOR4 (N202, N194, N101, N36, N64);
xor XOR2 (N203, N199, N194);
xor XOR2 (N204, N197, N95);
xor XOR2 (N205, N203, N143);
not NOT1 (N206, N204);
not NOT1 (N207, N195);
not NOT1 (N208, N188);
buf BUF1 (N209, N208);
and AND2 (N210, N201, N57);
or OR3 (N211, N202, N37, N150);
and AND4 (N212, N198, N16, N166, N191);
xor XOR2 (N213, N196, N154);
nor NOR4 (N214, N211, N95, N80, N21);
buf BUF1 (N215, N209);
nand NAND3 (N216, N205, N35, N147);
nor NOR3 (N217, N192, N105, N19);
and AND4 (N218, N207, N125, N82, N118);
xor XOR2 (N219, N217, N95);
and AND4 (N220, N213, N30, N70, N146);
not NOT1 (N221, N219);
or OR4 (N222, N206, N21, N198, N67);
xor XOR2 (N223, N215, N189);
buf BUF1 (N224, N218);
xor XOR2 (N225, N214, N162);
xor XOR2 (N226, N220, N184);
not NOT1 (N227, N225);
not NOT1 (N228, N227);
buf BUF1 (N229, N224);
buf BUF1 (N230, N210);
or OR4 (N231, N200, N18, N56, N48);
not NOT1 (N232, N221);
not NOT1 (N233, N229);
xor XOR2 (N234, N212, N167);
and AND4 (N235, N226, N234, N107, N158);
or OR4 (N236, N178, N132, N16, N149);
nor NOR4 (N237, N216, N204, N162, N173);
or OR3 (N238, N232, N226, N131);
xor XOR2 (N239, N222, N11);
xor XOR2 (N240, N231, N59);
or OR4 (N241, N236, N83, N50, N112);
not NOT1 (N242, N228);
or OR2 (N243, N237, N183);
nand NAND3 (N244, N238, N56, N45);
nor NOR2 (N245, N240, N146);
and AND3 (N246, N245, N22, N95);
and AND4 (N247, N246, N46, N52, N5);
nand NAND2 (N248, N241, N54);
xor XOR2 (N249, N239, N114);
or OR4 (N250, N249, N88, N83, N10);
nand NAND3 (N251, N250, N128, N220);
xor XOR2 (N252, N244, N137);
or OR4 (N253, N242, N100, N231, N91);
or OR4 (N254, N223, N59, N244, N118);
nand NAND4 (N255, N253, N182, N168, N38);
buf BUF1 (N256, N251);
xor XOR2 (N257, N256, N251);
nor NOR2 (N258, N243, N167);
nand NAND4 (N259, N258, N22, N100, N81);
xor XOR2 (N260, N252, N59);
nand NAND2 (N261, N257, N111);
nand NAND4 (N262, N233, N79, N201, N177);
nand NAND4 (N263, N255, N30, N137, N7);
buf BUF1 (N264, N261);
nand NAND2 (N265, N248, N25);
nand NAND2 (N266, N254, N179);
buf BUF1 (N267, N230);
or OR2 (N268, N267, N249);
nand NAND3 (N269, N265, N9, N130);
not NOT1 (N270, N264);
xor XOR2 (N271, N247, N14);
nor NOR4 (N272, N259, N262, N264, N125);
not NOT1 (N273, N75);
or OR4 (N274, N260, N171, N228, N258);
not NOT1 (N275, N263);
nor NOR4 (N276, N235, N261, N198, N186);
or OR2 (N277, N269, N15);
or OR3 (N278, N271, N132, N52);
not NOT1 (N279, N277);
not NOT1 (N280, N275);
nor NOR3 (N281, N280, N138, N32);
buf BUF1 (N282, N273);
or OR3 (N283, N272, N128, N74);
not NOT1 (N284, N266);
not NOT1 (N285, N284);
nand NAND2 (N286, N285, N151);
not NOT1 (N287, N279);
xor XOR2 (N288, N270, N156);
xor XOR2 (N289, N278, N143);
or OR3 (N290, N281, N256, N207);
or OR4 (N291, N268, N50, N43, N155);
nor NOR2 (N292, N290, N153);
or OR2 (N293, N274, N145);
buf BUF1 (N294, N288);
buf BUF1 (N295, N293);
or OR4 (N296, N282, N186, N221, N39);
buf BUF1 (N297, N283);
not NOT1 (N298, N287);
xor XOR2 (N299, N292, N40);
nor NOR3 (N300, N291, N175, N248);
xor XOR2 (N301, N286, N176);
not NOT1 (N302, N300);
nand NAND2 (N303, N297, N301);
nand NAND4 (N304, N49, N247, N2, N71);
and AND2 (N305, N302, N60);
nor NOR4 (N306, N296, N164, N45, N276);
nor NOR2 (N307, N113, N223);
xor XOR2 (N308, N295, N45);
nor NOR2 (N309, N289, N238);
or OR3 (N310, N308, N37, N59);
or OR3 (N311, N303, N173, N40);
buf BUF1 (N312, N298);
or OR3 (N313, N307, N150, N18);
buf BUF1 (N314, N310);
and AND2 (N315, N306, N301);
nand NAND3 (N316, N315, N237, N89);
buf BUF1 (N317, N311);
buf BUF1 (N318, N314);
buf BUF1 (N319, N318);
nor NOR2 (N320, N319, N250);
buf BUF1 (N321, N320);
buf BUF1 (N322, N317);
or OR2 (N323, N313, N228);
nor NOR3 (N324, N305, N106, N165);
xor XOR2 (N325, N323, N266);
xor XOR2 (N326, N304, N241);
xor XOR2 (N327, N326, N271);
or OR2 (N328, N299, N265);
xor XOR2 (N329, N322, N277);
nor NOR3 (N330, N316, N64, N272);
and AND4 (N331, N329, N275, N126, N119);
not NOT1 (N332, N327);
nor NOR2 (N333, N332, N111);
or OR4 (N334, N325, N223, N237, N86);
nor NOR2 (N335, N324, N110);
nand NAND4 (N336, N331, N331, N207, N180);
and AND4 (N337, N321, N44, N325, N31);
nor NOR2 (N338, N328, N200);
nand NAND4 (N339, N312, N68, N65, N3);
nand NAND3 (N340, N330, N2, N70);
nand NAND3 (N341, N336, N51, N150);
xor XOR2 (N342, N309, N204);
or OR3 (N343, N333, N35, N277);
nand NAND4 (N344, N343, N21, N151, N32);
buf BUF1 (N345, N340);
not NOT1 (N346, N335);
nor NOR2 (N347, N339, N34);
not NOT1 (N348, N338);
xor XOR2 (N349, N294, N304);
nand NAND2 (N350, N345, N89);
not NOT1 (N351, N348);
not NOT1 (N352, N337);
and AND3 (N353, N351, N304, N163);
xor XOR2 (N354, N353, N249);
buf BUF1 (N355, N347);
xor XOR2 (N356, N355, N102);
and AND4 (N357, N346, N319, N198, N157);
not NOT1 (N358, N344);
buf BUF1 (N359, N350);
not NOT1 (N360, N342);
nor NOR2 (N361, N354, N253);
nand NAND4 (N362, N341, N243, N204, N143);
xor XOR2 (N363, N349, N355);
buf BUF1 (N364, N360);
nand NAND4 (N365, N362, N319, N321, N257);
not NOT1 (N366, N361);
not NOT1 (N367, N364);
nand NAND2 (N368, N365, N181);
or OR3 (N369, N356, N116, N335);
not NOT1 (N370, N368);
nand NAND3 (N371, N352, N303, N217);
and AND4 (N372, N369, N266, N339, N292);
xor XOR2 (N373, N358, N338);
buf BUF1 (N374, N372);
or OR3 (N375, N334, N357, N56);
xor XOR2 (N376, N86, N186);
or OR3 (N377, N371, N22, N144);
not NOT1 (N378, N374);
not NOT1 (N379, N367);
not NOT1 (N380, N375);
buf BUF1 (N381, N378);
and AND3 (N382, N379, N16, N169);
and AND4 (N383, N370, N157, N184, N208);
nor NOR2 (N384, N363, N78);
or OR3 (N385, N359, N237, N218);
and AND4 (N386, N382, N197, N80, N1);
nand NAND4 (N387, N377, N357, N80, N27);
nor NOR4 (N388, N385, N329, N74, N54);
not NOT1 (N389, N376);
and AND4 (N390, N384, N83, N138, N245);
and AND4 (N391, N386, N68, N388, N223);
nand NAND3 (N392, N1, N168, N163);
buf BUF1 (N393, N387);
or OR3 (N394, N383, N34, N371);
buf BUF1 (N395, N380);
xor XOR2 (N396, N393, N380);
and AND2 (N397, N394, N32);
nor NOR4 (N398, N381, N126, N49, N30);
not NOT1 (N399, N366);
nand NAND3 (N400, N396, N286, N29);
or OR3 (N401, N391, N136, N132);
buf BUF1 (N402, N390);
not NOT1 (N403, N389);
and AND3 (N404, N395, N112, N150);
or OR3 (N405, N398, N266, N214);
nor NOR4 (N406, N405, N253, N324, N352);
not NOT1 (N407, N404);
and AND3 (N408, N406, N328, N54);
buf BUF1 (N409, N397);
xor XOR2 (N410, N408, N285);
buf BUF1 (N411, N403);
not NOT1 (N412, N373);
buf BUF1 (N413, N407);
or OR2 (N414, N410, N408);
or OR3 (N415, N411, N61, N218);
not NOT1 (N416, N409);
not NOT1 (N417, N401);
buf BUF1 (N418, N392);
not NOT1 (N419, N418);
and AND2 (N420, N402, N297);
buf BUF1 (N421, N419);
nor NOR2 (N422, N413, N136);
buf BUF1 (N423, N412);
xor XOR2 (N424, N422, N124);
buf BUF1 (N425, N420);
or OR2 (N426, N399, N386);
nor NOR4 (N427, N416, N349, N319, N319);
not NOT1 (N428, N400);
xor XOR2 (N429, N427, N350);
or OR3 (N430, N414, N299, N188);
and AND3 (N431, N421, N68, N354);
or OR2 (N432, N415, N348);
nand NAND2 (N433, N423, N8);
and AND2 (N434, N430, N324);
or OR2 (N435, N431, N280);
xor XOR2 (N436, N432, N115);
and AND2 (N437, N434, N177);
nor NOR2 (N438, N428, N417);
nor NOR4 (N439, N87, N379, N309, N152);
not NOT1 (N440, N435);
xor XOR2 (N441, N437, N111);
nand NAND3 (N442, N425, N16, N74);
not NOT1 (N443, N429);
nor NOR3 (N444, N426, N60, N311);
nor NOR2 (N445, N439, N26);
and AND3 (N446, N433, N117, N290);
nor NOR2 (N447, N441, N77);
nand NAND3 (N448, N444, N115, N162);
xor XOR2 (N449, N443, N160);
not NOT1 (N450, N436);
or OR2 (N451, N448, N157);
nor NOR2 (N452, N438, N14);
or OR4 (N453, N424, N123, N26, N217);
nor NOR4 (N454, N453, N70, N204, N118);
buf BUF1 (N455, N440);
or OR3 (N456, N445, N338, N436);
or OR3 (N457, N449, N446, N415);
xor XOR2 (N458, N55, N37);
not NOT1 (N459, N458);
and AND2 (N460, N459, N211);
nor NOR3 (N461, N451, N384, N124);
nand NAND3 (N462, N457, N360, N24);
not NOT1 (N463, N452);
xor XOR2 (N464, N460, N22);
not NOT1 (N465, N447);
xor XOR2 (N466, N455, N336);
and AND2 (N467, N463, N106);
not NOT1 (N468, N442);
buf BUF1 (N469, N468);
xor XOR2 (N470, N461, N316);
xor XOR2 (N471, N462, N435);
nand NAND3 (N472, N465, N454, N289);
nand NAND3 (N473, N322, N424, N163);
and AND2 (N474, N471, N47);
buf BUF1 (N475, N467);
nand NAND4 (N476, N475, N34, N170, N319);
buf BUF1 (N477, N456);
or OR3 (N478, N466, N198, N40);
nand NAND4 (N479, N464, N372, N266, N294);
nand NAND2 (N480, N476, N173);
not NOT1 (N481, N473);
nand NAND3 (N482, N481, N477, N148);
not NOT1 (N483, N295);
or OR3 (N484, N472, N216, N232);
and AND2 (N485, N469, N156);
buf BUF1 (N486, N483);
or OR4 (N487, N474, N190, N199, N189);
buf BUF1 (N488, N485);
or OR2 (N489, N479, N61);
not NOT1 (N490, N486);
or OR2 (N491, N450, N376);
xor XOR2 (N492, N489, N304);
buf BUF1 (N493, N491);
xor XOR2 (N494, N470, N81);
xor XOR2 (N495, N478, N22);
or OR2 (N496, N487, N92);
and AND2 (N497, N482, N320);
not NOT1 (N498, N497);
nand NAND3 (N499, N480, N365, N401);
or OR3 (N500, N488, N266, N112);
xor XOR2 (N501, N498, N18);
not NOT1 (N502, N499);
xor XOR2 (N503, N494, N41);
or OR3 (N504, N496, N434, N149);
nor NOR3 (N505, N492, N165, N474);
not NOT1 (N506, N495);
or OR4 (N507, N505, N166, N497, N149);
buf BUF1 (N508, N500);
nand NAND2 (N509, N507, N44);
buf BUF1 (N510, N504);
not NOT1 (N511, N490);
nand NAND4 (N512, N501, N397, N493, N460);
buf BUF1 (N513, N17);
nand NAND2 (N514, N513, N506);
or OR4 (N515, N83, N432, N511, N170);
nor NOR4 (N516, N273, N348, N195, N346);
xor XOR2 (N517, N515, N306);
xor XOR2 (N518, N512, N272);
not NOT1 (N519, N517);
or OR3 (N520, N508, N103, N129);
nand NAND2 (N521, N502, N80);
xor XOR2 (N522, N510, N284);
buf BUF1 (N523, N521);
buf BUF1 (N524, N514);
xor XOR2 (N525, N509, N114);
buf BUF1 (N526, N503);
and AND4 (N527, N522, N22, N322, N3);
or OR2 (N528, N523, N246);
or OR4 (N529, N516, N22, N60, N88);
not NOT1 (N530, N519);
xor XOR2 (N531, N527, N343);
or OR2 (N532, N525, N378);
buf BUF1 (N533, N529);
or OR2 (N534, N530, N35);
and AND2 (N535, N520, N440);
buf BUF1 (N536, N526);
or OR2 (N537, N531, N239);
xor XOR2 (N538, N528, N481);
nor NOR3 (N539, N537, N519, N174);
and AND4 (N540, N484, N51, N115, N444);
nand NAND3 (N541, N534, N530, N411);
buf BUF1 (N542, N539);
xor XOR2 (N543, N535, N352);
nand NAND2 (N544, N538, N88);
not NOT1 (N545, N542);
buf BUF1 (N546, N544);
buf BUF1 (N547, N540);
and AND3 (N548, N543, N48, N50);
buf BUF1 (N549, N533);
nand NAND3 (N550, N532, N421, N331);
not NOT1 (N551, N541);
not NOT1 (N552, N546);
nor NOR3 (N553, N549, N346, N209);
nand NAND4 (N554, N550, N163, N160, N198);
buf BUF1 (N555, N553);
not NOT1 (N556, N545);
and AND4 (N557, N547, N546, N446, N275);
buf BUF1 (N558, N536);
buf BUF1 (N559, N554);
buf BUF1 (N560, N557);
nand NAND4 (N561, N558, N222, N276, N482);
not NOT1 (N562, N548);
not NOT1 (N563, N518);
and AND4 (N564, N562, N153, N110, N371);
or OR4 (N565, N555, N452, N158, N164);
not NOT1 (N566, N560);
not NOT1 (N567, N552);
nand NAND3 (N568, N565, N423, N132);
buf BUF1 (N569, N567);
or OR2 (N570, N551, N62);
and AND3 (N571, N566, N84, N225);
or OR2 (N572, N559, N166);
or OR2 (N573, N568, N64);
nor NOR2 (N574, N572, N77);
not NOT1 (N575, N524);
or OR4 (N576, N563, N124, N97, N454);
nor NOR3 (N577, N570, N169, N67);
nand NAND2 (N578, N576, N425);
xor XOR2 (N579, N571, N541);
and AND3 (N580, N556, N450, N103);
buf BUF1 (N581, N575);
or OR4 (N582, N578, N133, N326, N114);
nor NOR2 (N583, N579, N451);
not NOT1 (N584, N581);
or OR4 (N585, N584, N261, N252, N205);
xor XOR2 (N586, N582, N95);
and AND3 (N587, N586, N472, N45);
buf BUF1 (N588, N574);
xor XOR2 (N589, N573, N18);
nand NAND3 (N590, N588, N494, N522);
nand NAND4 (N591, N580, N242, N324, N274);
xor XOR2 (N592, N583, N91);
not NOT1 (N593, N587);
buf BUF1 (N594, N564);
and AND4 (N595, N594, N372, N135, N455);
or OR4 (N596, N561, N354, N504, N450);
and AND2 (N597, N595, N77);
xor XOR2 (N598, N589, N324);
xor XOR2 (N599, N592, N355);
and AND2 (N600, N599, N267);
nor NOR4 (N601, N590, N272, N103, N83);
xor XOR2 (N602, N577, N466);
nor NOR3 (N603, N601, N309, N121);
not NOT1 (N604, N600);
nor NOR2 (N605, N585, N358);
and AND3 (N606, N598, N163, N404);
nor NOR2 (N607, N569, N221);
and AND3 (N608, N596, N281, N309);
nor NOR3 (N609, N605, N501, N552);
nand NAND2 (N610, N593, N438);
or OR3 (N611, N609, N543, N22);
nor NOR3 (N612, N604, N49, N245);
and AND3 (N613, N610, N587, N167);
nand NAND3 (N614, N611, N285, N164);
xor XOR2 (N615, N612, N592);
not NOT1 (N616, N613);
nor NOR2 (N617, N606, N424);
nand NAND3 (N618, N597, N262, N278);
buf BUF1 (N619, N617);
or OR2 (N620, N616, N158);
nand NAND2 (N621, N615, N148);
nand NAND2 (N622, N607, N254);
buf BUF1 (N623, N602);
not NOT1 (N624, N620);
and AND2 (N625, N614, N271);
and AND4 (N626, N621, N471, N428, N406);
nor NOR2 (N627, N622, N560);
or OR3 (N628, N623, N517, N195);
not NOT1 (N629, N624);
or OR3 (N630, N618, N502, N619);
nor NOR4 (N631, N597, N269, N239, N473);
nand NAND2 (N632, N625, N532);
not NOT1 (N633, N627);
and AND3 (N634, N591, N545, N457);
buf BUF1 (N635, N632);
or OR4 (N636, N628, N196, N269, N425);
xor XOR2 (N637, N630, N168);
nor NOR2 (N638, N634, N341);
and AND4 (N639, N603, N236, N275, N75);
nand NAND2 (N640, N635, N77);
buf BUF1 (N641, N638);
not NOT1 (N642, N637);
buf BUF1 (N643, N642);
nor NOR2 (N644, N631, N163);
not NOT1 (N645, N608);
nor NOR2 (N646, N626, N288);
nand NAND4 (N647, N639, N214, N413, N276);
or OR4 (N648, N647, N241, N272, N64);
and AND3 (N649, N641, N176, N487);
or OR3 (N650, N645, N526, N356);
or OR4 (N651, N649, N240, N209, N339);
or OR3 (N652, N629, N562, N410);
or OR3 (N653, N640, N116, N588);
or OR2 (N654, N633, N645);
xor XOR2 (N655, N644, N1);
and AND2 (N656, N655, N76);
nor NOR4 (N657, N648, N598, N553, N236);
xor XOR2 (N658, N652, N380);
and AND2 (N659, N643, N561);
buf BUF1 (N660, N657);
xor XOR2 (N661, N659, N145);
and AND4 (N662, N651, N11, N289, N648);
buf BUF1 (N663, N662);
nand NAND2 (N664, N646, N233);
and AND2 (N665, N661, N633);
or OR4 (N666, N664, N502, N293, N297);
or OR2 (N667, N654, N426);
and AND4 (N668, N666, N221, N105, N558);
nor NOR3 (N669, N667, N634, N514);
or OR4 (N670, N636, N114, N268, N665);
nor NOR2 (N671, N38, N154);
not NOT1 (N672, N668);
or OR4 (N673, N653, N4, N370, N18);
and AND4 (N674, N650, N548, N605, N102);
xor XOR2 (N675, N656, N208);
nor NOR3 (N676, N669, N614, N563);
or OR2 (N677, N658, N177);
not NOT1 (N678, N660);
and AND2 (N679, N670, N307);
nand NAND4 (N680, N663, N259, N592, N359);
nor NOR3 (N681, N672, N60, N296);
and AND4 (N682, N673, N263, N642, N227);
buf BUF1 (N683, N678);
not NOT1 (N684, N680);
nand NAND4 (N685, N684, N427, N528, N635);
nand NAND3 (N686, N671, N541, N597);
nand NAND4 (N687, N682, N344, N45, N60);
not NOT1 (N688, N675);
xor XOR2 (N689, N681, N529);
and AND2 (N690, N687, N18);
not NOT1 (N691, N686);
or OR3 (N692, N690, N54, N134);
nor NOR2 (N693, N688, N327);
nand NAND4 (N694, N683, N378, N604, N14);
nor NOR4 (N695, N685, N690, N347, N521);
nor NOR3 (N696, N693, N631, N602);
nand NAND4 (N697, N694, N298, N338, N628);
nand NAND4 (N698, N679, N440, N655, N16);
not NOT1 (N699, N691);
nand NAND3 (N700, N676, N592, N600);
nor NOR2 (N701, N692, N605);
and AND3 (N702, N700, N101, N105);
nor NOR2 (N703, N697, N225);
and AND2 (N704, N696, N172);
not NOT1 (N705, N701);
not NOT1 (N706, N699);
nand NAND2 (N707, N674, N427);
and AND4 (N708, N705, N309, N613, N632);
or OR2 (N709, N677, N468);
buf BUF1 (N710, N708);
buf BUF1 (N711, N704);
not NOT1 (N712, N706);
and AND2 (N713, N702, N81);
xor XOR2 (N714, N695, N102);
nor NOR4 (N715, N698, N77, N456, N514);
buf BUF1 (N716, N709);
or OR4 (N717, N712, N175, N129, N419);
not NOT1 (N718, N716);
and AND3 (N719, N718, N140, N473);
and AND2 (N720, N714, N207);
and AND4 (N721, N719, N277, N54, N451);
not NOT1 (N722, N710);
or OR2 (N723, N722, N326);
nand NAND4 (N724, N717, N412, N324, N478);
nor NOR2 (N725, N723, N96);
nand NAND2 (N726, N707, N664);
and AND4 (N727, N715, N693, N261, N275);
and AND4 (N728, N727, N478, N630, N602);
xor XOR2 (N729, N720, N375);
buf BUF1 (N730, N729);
nand NAND3 (N731, N689, N197, N390);
nor NOR3 (N732, N725, N277, N189);
xor XOR2 (N733, N721, N564);
not NOT1 (N734, N713);
not NOT1 (N735, N728);
nand NAND2 (N736, N734, N364);
not NOT1 (N737, N730);
nand NAND4 (N738, N736, N676, N677, N351);
buf BUF1 (N739, N703);
or OR2 (N740, N732, N503);
or OR2 (N741, N731, N27);
nand NAND4 (N742, N735, N195, N128, N620);
nor NOR3 (N743, N742, N203, N447);
buf BUF1 (N744, N740);
nand NAND3 (N745, N724, N536, N129);
and AND4 (N746, N744, N614, N21, N542);
or OR3 (N747, N738, N291, N432);
xor XOR2 (N748, N739, N663);
xor XOR2 (N749, N741, N469);
nor NOR3 (N750, N726, N724, N603);
and AND3 (N751, N737, N132, N121);
and AND2 (N752, N743, N677);
not NOT1 (N753, N747);
not NOT1 (N754, N750);
or OR4 (N755, N753, N133, N15, N249);
or OR2 (N756, N754, N133);
and AND3 (N757, N752, N617, N628);
nand NAND4 (N758, N711, N501, N441, N747);
and AND2 (N759, N733, N62);
not NOT1 (N760, N756);
nor NOR4 (N761, N746, N22, N465, N449);
xor XOR2 (N762, N748, N477);
nor NOR4 (N763, N745, N342, N277, N317);
buf BUF1 (N764, N762);
xor XOR2 (N765, N755, N539);
not NOT1 (N766, N760);
not NOT1 (N767, N761);
or OR3 (N768, N758, N574, N115);
or OR4 (N769, N757, N624, N313, N192);
nand NAND2 (N770, N759, N706);
nand NAND3 (N771, N751, N337, N345);
or OR3 (N772, N766, N188, N750);
and AND4 (N773, N770, N277, N363, N226);
or OR2 (N774, N767, N471);
or OR3 (N775, N772, N332, N682);
nor NOR2 (N776, N769, N191);
xor XOR2 (N777, N749, N10);
or OR4 (N778, N768, N673, N518, N208);
buf BUF1 (N779, N765);
and AND3 (N780, N774, N683, N163);
nand NAND3 (N781, N775, N527, N543);
or OR4 (N782, N763, N210, N625, N64);
nor NOR2 (N783, N781, N391);
buf BUF1 (N784, N779);
not NOT1 (N785, N776);
buf BUF1 (N786, N784);
nand NAND4 (N787, N780, N4, N126, N422);
and AND4 (N788, N783, N419, N455, N679);
xor XOR2 (N789, N787, N395);
or OR2 (N790, N789, N590);
not NOT1 (N791, N778);
nand NAND2 (N792, N791, N584);
buf BUF1 (N793, N786);
buf BUF1 (N794, N785);
and AND3 (N795, N788, N151, N69);
or OR4 (N796, N790, N133, N350, N475);
nor NOR4 (N797, N795, N427, N250, N194);
buf BUF1 (N798, N797);
buf BUF1 (N799, N793);
buf BUF1 (N800, N782);
or OR2 (N801, N799, N120);
nand NAND3 (N802, N798, N474, N43);
xor XOR2 (N803, N801, N573);
buf BUF1 (N804, N796);
nand NAND3 (N805, N777, N261, N12);
not NOT1 (N806, N794);
not NOT1 (N807, N773);
or OR4 (N808, N804, N570, N509, N504);
buf BUF1 (N809, N803);
not NOT1 (N810, N792);
or OR2 (N811, N764, N574);
buf BUF1 (N812, N811);
or OR3 (N813, N800, N73, N386);
and AND3 (N814, N808, N614, N565);
nand NAND2 (N815, N809, N17);
or OR2 (N816, N771, N125);
buf BUF1 (N817, N806);
nand NAND3 (N818, N812, N264, N165);
nor NOR3 (N819, N816, N473, N258);
or OR2 (N820, N802, N478);
and AND3 (N821, N805, N440, N84);
nand NAND2 (N822, N813, N618);
xor XOR2 (N823, N819, N569);
xor XOR2 (N824, N823, N755);
and AND3 (N825, N820, N397, N718);
nor NOR4 (N826, N824, N505, N735, N199);
nand NAND4 (N827, N817, N70, N757, N700);
nor NOR2 (N828, N818, N91);
and AND4 (N829, N810, N96, N610, N188);
nand NAND4 (N830, N828, N295, N18, N64);
not NOT1 (N831, N815);
not NOT1 (N832, N830);
nor NOR3 (N833, N807, N698, N72);
or OR4 (N834, N831, N301, N196, N375);
nand NAND4 (N835, N821, N405, N489, N799);
buf BUF1 (N836, N835);
and AND3 (N837, N822, N401, N466);
xor XOR2 (N838, N833, N420);
nand NAND4 (N839, N827, N425, N822, N538);
nand NAND2 (N840, N825, N519);
buf BUF1 (N841, N837);
buf BUF1 (N842, N840);
and AND2 (N843, N829, N351);
and AND4 (N844, N841, N781, N773, N616);
nand NAND2 (N845, N826, N677);
or OR4 (N846, N832, N294, N838, N75);
buf BUF1 (N847, N648);
nor NOR4 (N848, N839, N693, N258, N255);
buf BUF1 (N849, N843);
and AND2 (N850, N834, N605);
nand NAND2 (N851, N848, N48);
nand NAND2 (N852, N842, N139);
xor XOR2 (N853, N836, N281);
or OR2 (N854, N851, N155);
xor XOR2 (N855, N852, N733);
xor XOR2 (N856, N845, N560);
buf BUF1 (N857, N847);
nand NAND3 (N858, N857, N663, N101);
not NOT1 (N859, N850);
and AND4 (N860, N814, N327, N33, N606);
nor NOR4 (N861, N855, N856, N151, N586);
nand NAND4 (N862, N124, N690, N619, N850);
or OR3 (N863, N844, N531, N649);
and AND2 (N864, N862, N405);
and AND3 (N865, N854, N781, N84);
buf BUF1 (N866, N849);
not NOT1 (N867, N853);
or OR2 (N868, N866, N171);
and AND2 (N869, N859, N676);
not NOT1 (N870, N860);
nor NOR3 (N871, N846, N190, N540);
and AND4 (N872, N861, N755, N824, N50);
not NOT1 (N873, N871);
and AND2 (N874, N858, N535);
and AND3 (N875, N863, N743, N671);
nand NAND3 (N876, N869, N704, N75);
xor XOR2 (N877, N865, N94);
buf BUF1 (N878, N872);
or OR4 (N879, N877, N170, N141, N790);
or OR2 (N880, N875, N111);
or OR4 (N881, N868, N349, N414, N34);
not NOT1 (N882, N867);
nand NAND3 (N883, N864, N525, N601);
nand NAND3 (N884, N878, N102, N244);
xor XOR2 (N885, N870, N198);
not NOT1 (N886, N884);
xor XOR2 (N887, N886, N279);
nand NAND4 (N888, N885, N209, N136, N867);
and AND2 (N889, N881, N17);
xor XOR2 (N890, N874, N326);
xor XOR2 (N891, N889, N295);
or OR4 (N892, N882, N71, N25, N638);
or OR2 (N893, N876, N129);
nor NOR3 (N894, N879, N578, N205);
nor NOR4 (N895, N883, N853, N334, N474);
nor NOR3 (N896, N887, N617, N145);
nand NAND3 (N897, N890, N817, N735);
or OR3 (N898, N891, N719, N752);
or OR2 (N899, N873, N793);
buf BUF1 (N900, N898);
not NOT1 (N901, N888);
nor NOR3 (N902, N892, N534, N760);
not NOT1 (N903, N897);
not NOT1 (N904, N894);
or OR3 (N905, N901, N558, N878);
xor XOR2 (N906, N896, N609);
or OR2 (N907, N906, N399);
not NOT1 (N908, N900);
nor NOR4 (N909, N895, N885, N62, N369);
nand NAND4 (N910, N899, N264, N591, N731);
or OR2 (N911, N880, N377);
xor XOR2 (N912, N907, N844);
buf BUF1 (N913, N912);
xor XOR2 (N914, N911, N795);
or OR4 (N915, N913, N381, N43, N284);
or OR2 (N916, N893, N402);
buf BUF1 (N917, N902);
and AND3 (N918, N909, N418, N698);
buf BUF1 (N919, N916);
nand NAND4 (N920, N914, N447, N846, N124);
nand NAND3 (N921, N908, N501, N656);
buf BUF1 (N922, N921);
nand NAND2 (N923, N922, N78);
not NOT1 (N924, N923);
buf BUF1 (N925, N910);
not NOT1 (N926, N925);
or OR2 (N927, N924, N864);
nor NOR2 (N928, N926, N824);
or OR3 (N929, N917, N175, N562);
xor XOR2 (N930, N919, N160);
or OR4 (N931, N930, N115, N279, N889);
nand NAND4 (N932, N915, N383, N682, N67);
nor NOR3 (N933, N928, N293, N473);
not NOT1 (N934, N904);
buf BUF1 (N935, N927);
nand NAND2 (N936, N903, N371);
xor XOR2 (N937, N933, N402);
or OR4 (N938, N932, N678, N793, N364);
or OR4 (N939, N920, N883, N93, N567);
and AND4 (N940, N905, N45, N399, N938);
xor XOR2 (N941, N29, N198);
nor NOR3 (N942, N918, N582, N175);
and AND4 (N943, N941, N365, N822, N736);
not NOT1 (N944, N937);
not NOT1 (N945, N936);
and AND4 (N946, N931, N304, N650, N330);
and AND3 (N947, N935, N855, N838);
xor XOR2 (N948, N940, N695);
nand NAND3 (N949, N929, N443, N688);
not NOT1 (N950, N942);
and AND2 (N951, N934, N230);
or OR4 (N952, N951, N385, N445, N598);
xor XOR2 (N953, N952, N180);
nor NOR3 (N954, N939, N812, N467);
nand NAND4 (N955, N947, N21, N557, N581);
and AND2 (N956, N955, N144);
nand NAND3 (N957, N950, N247, N295);
nor NOR4 (N958, N943, N617, N282, N743);
nand NAND4 (N959, N946, N426, N321, N395);
and AND4 (N960, N944, N233, N629, N276);
nor NOR2 (N961, N958, N4);
xor XOR2 (N962, N956, N172);
xor XOR2 (N963, N962, N163);
and AND3 (N964, N948, N671, N314);
nor NOR4 (N965, N960, N777, N666, N327);
nor NOR3 (N966, N945, N60, N190);
nand NAND2 (N967, N949, N455);
not NOT1 (N968, N965);
nand NAND3 (N969, N963, N324, N897);
or OR4 (N970, N969, N239, N399, N489);
xor XOR2 (N971, N966, N596);
and AND2 (N972, N967, N760);
nand NAND2 (N973, N954, N694);
xor XOR2 (N974, N953, N383);
nor NOR3 (N975, N973, N752, N478);
and AND2 (N976, N975, N71);
not NOT1 (N977, N961);
buf BUF1 (N978, N964);
nand NAND2 (N979, N968, N84);
not NOT1 (N980, N978);
xor XOR2 (N981, N971, N571);
not NOT1 (N982, N979);
xor XOR2 (N983, N981, N399);
buf BUF1 (N984, N974);
nand NAND2 (N985, N959, N855);
or OR2 (N986, N985, N540);
nor NOR4 (N987, N977, N916, N171, N819);
not NOT1 (N988, N976);
buf BUF1 (N989, N988);
and AND2 (N990, N983, N118);
nor NOR4 (N991, N972, N860, N899, N872);
nor NOR3 (N992, N982, N50, N116);
and AND3 (N993, N989, N991, N440);
nor NOR2 (N994, N505, N423);
and AND4 (N995, N957, N113, N75, N204);
not NOT1 (N996, N984);
and AND3 (N997, N992, N578, N412);
buf BUF1 (N998, N994);
nand NAND4 (N999, N998, N321, N752, N29);
nand NAND4 (N1000, N995, N353, N51, N506);
buf BUF1 (N1001, N999);
xor XOR2 (N1002, N993, N416);
xor XOR2 (N1003, N996, N991);
not NOT1 (N1004, N986);
nand NAND4 (N1005, N1003, N538, N119, N645);
and AND4 (N1006, N1002, N109, N746, N236);
not NOT1 (N1007, N987);
or OR4 (N1008, N1005, N994, N970, N507);
xor XOR2 (N1009, N1007, N426);
xor XOR2 (N1010, N748, N617);
and AND2 (N1011, N1001, N702);
not NOT1 (N1012, N1008);
nor NOR2 (N1013, N1009, N531);
not NOT1 (N1014, N997);
xor XOR2 (N1015, N1014, N872);
endmodule