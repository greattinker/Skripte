// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N310,N305,N313,N290,N293,N312,N304,N311,N309,N314;

nand NAND2 (N15, N6, N8);
xor XOR2 (N16, N5, N9);
nor NOR4 (N17, N2, N2, N6, N2);
not NOT1 (N18, N6);
nor NOR2 (N19, N15, N4);
nand NAND2 (N20, N13, N6);
xor XOR2 (N21, N6, N12);
and AND4 (N22, N10, N15, N16, N8);
or OR2 (N23, N7, N13);
and AND3 (N24, N8, N2, N13);
or OR4 (N25, N9, N1, N21, N8);
and AND2 (N26, N18, N4);
nor NOR3 (N27, N24, N21, N13);
nor NOR2 (N28, N17, N27);
buf BUF1 (N29, N1);
or OR3 (N30, N11, N17, N7);
or OR3 (N31, N28, N6, N2);
xor XOR2 (N32, N12, N1);
and AND3 (N33, N31, N22, N21);
not NOT1 (N34, N32);
and AND3 (N35, N20, N8, N2);
or OR4 (N36, N28, N18, N5, N9);
xor XOR2 (N37, N34, N12);
xor XOR2 (N38, N37, N6);
or OR4 (N39, N35, N1, N26, N13);
not NOT1 (N40, N39);
buf BUF1 (N41, N29);
not NOT1 (N42, N16);
buf BUF1 (N43, N38);
nor NOR4 (N44, N19, N9, N19, N14);
nand NAND2 (N45, N33, N19);
nand NAND3 (N46, N42, N8, N39);
xor XOR2 (N47, N23, N4);
nand NAND3 (N48, N41, N12, N33);
not NOT1 (N49, N47);
buf BUF1 (N50, N36);
not NOT1 (N51, N40);
nand NAND2 (N52, N49, N29);
or OR4 (N53, N50, N15, N42, N39);
not NOT1 (N54, N43);
nand NAND3 (N55, N44, N14, N46);
buf BUF1 (N56, N12);
and AND4 (N57, N45, N4, N46, N25);
and AND2 (N58, N52, N39);
and AND3 (N59, N46, N1, N31);
nand NAND3 (N60, N58, N59, N28);
nor NOR2 (N61, N50, N46);
not NOT1 (N62, N57);
xor XOR2 (N63, N61, N60);
xor XOR2 (N64, N61, N43);
xor XOR2 (N65, N55, N14);
or OR4 (N66, N48, N13, N31, N22);
buf BUF1 (N67, N63);
and AND4 (N68, N54, N12, N63, N38);
or OR4 (N69, N68, N14, N60, N23);
xor XOR2 (N70, N51, N35);
buf BUF1 (N71, N70);
nor NOR2 (N72, N56, N39);
and AND4 (N73, N72, N1, N28, N64);
buf BUF1 (N74, N56);
nor NOR2 (N75, N65, N20);
not NOT1 (N76, N74);
xor XOR2 (N77, N69, N68);
nor NOR2 (N78, N30, N71);
nor NOR4 (N79, N51, N2, N63, N32);
and AND3 (N80, N77, N46, N60);
nand NAND4 (N81, N76, N27, N36, N17);
nor NOR3 (N82, N79, N49, N41);
nor NOR3 (N83, N73, N45, N20);
nor NOR4 (N84, N82, N68, N77, N47);
not NOT1 (N85, N53);
and AND4 (N86, N84, N12, N5, N67);
nand NAND2 (N87, N21, N24);
or OR4 (N88, N85, N17, N23, N75);
buf BUF1 (N89, N34);
nor NOR2 (N90, N83, N17);
not NOT1 (N91, N62);
not NOT1 (N92, N78);
xor XOR2 (N93, N92, N2);
buf BUF1 (N94, N89);
or OR3 (N95, N90, N62, N77);
not NOT1 (N96, N87);
not NOT1 (N97, N86);
or OR2 (N98, N96, N72);
nand NAND4 (N99, N93, N46, N46, N31);
nor NOR4 (N100, N98, N90, N66, N47);
xor XOR2 (N101, N63, N9);
nand NAND4 (N102, N94, N101, N61, N35);
not NOT1 (N103, N27);
xor XOR2 (N104, N91, N102);
and AND2 (N105, N26, N27);
not NOT1 (N106, N95);
nor NOR4 (N107, N88, N21, N85, N76);
nand NAND4 (N108, N100, N79, N43, N17);
xor XOR2 (N109, N103, N81);
not NOT1 (N110, N36);
and AND3 (N111, N107, N57, N17);
nand NAND4 (N112, N99, N51, N53, N9);
nor NOR3 (N113, N112, N88, N71);
not NOT1 (N114, N108);
or OR2 (N115, N113, N29);
nor NOR2 (N116, N106, N35);
nand NAND3 (N117, N111, N95, N48);
nor NOR2 (N118, N110, N22);
and AND3 (N119, N117, N34, N54);
nor NOR2 (N120, N115, N34);
nand NAND4 (N121, N104, N80, N101, N94);
and AND3 (N122, N17, N107, N36);
xor XOR2 (N123, N114, N16);
or OR2 (N124, N121, N59);
buf BUF1 (N125, N97);
nand NAND3 (N126, N120, N11, N108);
or OR3 (N127, N116, N40, N22);
buf BUF1 (N128, N122);
xor XOR2 (N129, N125, N50);
and AND4 (N130, N127, N27, N122, N21);
nor NOR3 (N131, N129, N112, N94);
buf BUF1 (N132, N123);
nor NOR2 (N133, N124, N58);
nand NAND4 (N134, N132, N76, N94, N114);
xor XOR2 (N135, N126, N8);
nand NAND3 (N136, N118, N121, N124);
and AND4 (N137, N133, N42, N10, N25);
xor XOR2 (N138, N109, N12);
buf BUF1 (N139, N136);
and AND2 (N140, N139, N79);
buf BUF1 (N141, N135);
and AND2 (N142, N137, N63);
buf BUF1 (N143, N119);
nor NOR2 (N144, N131, N76);
buf BUF1 (N145, N142);
buf BUF1 (N146, N128);
buf BUF1 (N147, N130);
nor NOR4 (N148, N144, N54, N13, N136);
nand NAND3 (N149, N143, N20, N80);
not NOT1 (N150, N148);
not NOT1 (N151, N134);
not NOT1 (N152, N146);
or OR2 (N153, N147, N35);
buf BUF1 (N154, N152);
or OR4 (N155, N138, N100, N33, N147);
or OR4 (N156, N151, N104, N147, N9);
buf BUF1 (N157, N156);
nor NOR4 (N158, N157, N141, N92, N88);
or OR3 (N159, N147, N96, N9);
buf BUF1 (N160, N149);
xor XOR2 (N161, N155, N67);
not NOT1 (N162, N145);
or OR2 (N163, N153, N85);
nor NOR2 (N164, N158, N80);
nand NAND3 (N165, N164, N21, N156);
nand NAND3 (N166, N161, N91, N129);
not NOT1 (N167, N166);
nor NOR3 (N168, N163, N125, N129);
nor NOR2 (N169, N105, N48);
nand NAND4 (N170, N169, N3, N145, N87);
and AND3 (N171, N170, N86, N157);
buf BUF1 (N172, N140);
nand NAND3 (N173, N162, N158, N113);
not NOT1 (N174, N165);
nor NOR4 (N175, N154, N128, N150, N170);
xor XOR2 (N176, N99, N165);
xor XOR2 (N177, N160, N96);
and AND2 (N178, N167, N69);
nand NAND2 (N179, N172, N124);
nor NOR2 (N180, N174, N163);
nor NOR3 (N181, N168, N11, N122);
and AND3 (N182, N178, N28, N75);
and AND2 (N183, N177, N172);
buf BUF1 (N184, N176);
not NOT1 (N185, N175);
or OR2 (N186, N184, N182);
nand NAND4 (N187, N17, N86, N70, N14);
nand NAND2 (N188, N180, N30);
buf BUF1 (N189, N183);
nor NOR3 (N190, N181, N44, N159);
xor XOR2 (N191, N180, N28);
nand NAND2 (N192, N190, N191);
and AND3 (N193, N33, N104, N108);
or OR2 (N194, N193, N82);
not NOT1 (N195, N189);
and AND2 (N196, N173, N77);
xor XOR2 (N197, N185, N111);
xor XOR2 (N198, N179, N168);
buf BUF1 (N199, N194);
nor NOR4 (N200, N197, N149, N119, N99);
xor XOR2 (N201, N187, N16);
and AND4 (N202, N188, N118, N42, N197);
buf BUF1 (N203, N200);
buf BUF1 (N204, N201);
not NOT1 (N205, N203);
or OR4 (N206, N195, N162, N128, N31);
buf BUF1 (N207, N205);
or OR4 (N208, N192, N68, N55, N112);
and AND3 (N209, N202, N163, N117);
xor XOR2 (N210, N186, N79);
nor NOR2 (N211, N207, N88);
xor XOR2 (N212, N210, N175);
or OR3 (N213, N211, N40, N136);
not NOT1 (N214, N208);
nor NOR2 (N215, N213, N209);
xor XOR2 (N216, N26, N179);
xor XOR2 (N217, N216, N68);
buf BUF1 (N218, N171);
or OR4 (N219, N199, N196, N146, N158);
nor NOR4 (N220, N147, N84, N90, N25);
nor NOR4 (N221, N204, N101, N50, N71);
nand NAND4 (N222, N221, N16, N36, N14);
not NOT1 (N223, N220);
or OR4 (N224, N223, N129, N178, N216);
or OR4 (N225, N206, N149, N54, N50);
and AND3 (N226, N214, N77, N157);
buf BUF1 (N227, N217);
and AND2 (N228, N227, N32);
not NOT1 (N229, N218);
nand NAND2 (N230, N225, N130);
or OR3 (N231, N229, N12, N5);
xor XOR2 (N232, N226, N74);
nand NAND2 (N233, N198, N185);
buf BUF1 (N234, N224);
xor XOR2 (N235, N212, N210);
or OR4 (N236, N231, N186, N22, N93);
and AND2 (N237, N219, N186);
or OR4 (N238, N234, N232, N49, N197);
nor NOR2 (N239, N205, N207);
buf BUF1 (N240, N228);
and AND3 (N241, N236, N206, N124);
nor NOR4 (N242, N230, N225, N166, N198);
xor XOR2 (N243, N239, N41);
nor NOR4 (N244, N222, N74, N91, N112);
nand NAND4 (N245, N235, N129, N119, N118);
buf BUF1 (N246, N241);
xor XOR2 (N247, N237, N208);
xor XOR2 (N248, N240, N236);
buf BUF1 (N249, N215);
and AND3 (N250, N242, N143, N98);
or OR3 (N251, N243, N155, N192);
and AND4 (N252, N245, N199, N143, N144);
xor XOR2 (N253, N252, N181);
buf BUF1 (N254, N244);
nand NAND3 (N255, N251, N246, N191);
buf BUF1 (N256, N140);
nand NAND3 (N257, N255, N102, N178);
buf BUF1 (N258, N247);
or OR4 (N259, N257, N148, N120, N158);
or OR3 (N260, N238, N149, N223);
nand NAND2 (N261, N258, N199);
nor NOR3 (N262, N256, N244, N1);
and AND4 (N263, N250, N257, N206, N213);
not NOT1 (N264, N249);
and AND4 (N265, N248, N129, N12, N33);
and AND2 (N266, N233, N136);
and AND2 (N267, N253, N237);
or OR4 (N268, N265, N126, N262, N107);
not NOT1 (N269, N49);
and AND4 (N270, N259, N178, N156, N113);
or OR3 (N271, N266, N249, N260);
nor NOR3 (N272, N242, N168, N189);
and AND2 (N273, N271, N54);
and AND3 (N274, N261, N145, N41);
and AND3 (N275, N272, N38, N100);
xor XOR2 (N276, N273, N89);
or OR3 (N277, N275, N275, N239);
xor XOR2 (N278, N269, N40);
xor XOR2 (N279, N264, N118);
or OR4 (N280, N276, N186, N56, N151);
nand NAND2 (N281, N270, N146);
xor XOR2 (N282, N274, N149);
nor NOR3 (N283, N281, N115, N227);
nor NOR3 (N284, N268, N85, N216);
nand NAND4 (N285, N279, N81, N232, N268);
not NOT1 (N286, N285);
nand NAND4 (N287, N280, N15, N118, N221);
and AND2 (N288, N284, N164);
or OR2 (N289, N278, N192);
nor NOR3 (N290, N289, N105, N234);
xor XOR2 (N291, N254, N236);
or OR3 (N292, N267, N266, N213);
and AND2 (N293, N291, N158);
and AND3 (N294, N282, N162, N245);
buf BUF1 (N295, N277);
buf BUF1 (N296, N286);
xor XOR2 (N297, N294, N123);
and AND2 (N298, N292, N214);
and AND2 (N299, N288, N152);
nor NOR4 (N300, N299, N275, N206, N189);
nand NAND3 (N301, N287, N233, N228);
nand NAND3 (N302, N296, N301, N212);
xor XOR2 (N303, N186, N247);
buf BUF1 (N304, N297);
buf BUF1 (N305, N303);
nor NOR2 (N306, N263, N299);
buf BUF1 (N307, N302);
or OR4 (N308, N295, N25, N301, N107);
nor NOR2 (N309, N298, N36);
buf BUF1 (N310, N283);
nor NOR4 (N311, N307, N294, N11, N121);
nand NAND2 (N312, N306, N289);
xor XOR2 (N313, N300, N64);
xor XOR2 (N314, N308, N173);
endmodule