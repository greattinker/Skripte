// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N2508,N2487,N2492,N2497,N2504,N2507,N2499,N2505,N2509,N2510;

xor XOR2 (N11, N2, N10);
not NOT1 (N12, N3);
xor XOR2 (N13, N12, N6);
nand NAND2 (N14, N6, N2);
nor NOR3 (N15, N14, N6, N14);
and AND4 (N16, N4, N14, N9, N4);
xor XOR2 (N17, N14, N15);
buf BUF1 (N18, N9);
nor NOR4 (N19, N4, N2, N12, N11);
nor NOR4 (N20, N18, N19, N17, N5);
not NOT1 (N21, N14);
xor XOR2 (N22, N13, N6);
nand NAND2 (N23, N6, N1);
nor NOR2 (N24, N14, N7);
xor XOR2 (N25, N15, N13);
and AND4 (N26, N2, N25, N13, N18);
or OR2 (N27, N7, N3);
or OR4 (N28, N15, N11, N27, N23);
and AND2 (N29, N8, N20);
not NOT1 (N30, N10);
nand NAND3 (N31, N19, N2, N6);
or OR3 (N32, N12, N27, N17);
nand NAND4 (N33, N30, N21, N12, N4);
not NOT1 (N34, N10);
nand NAND2 (N35, N16, N15);
buf BUF1 (N36, N22);
or OR2 (N37, N33, N13);
or OR4 (N38, N35, N8, N25, N14);
not NOT1 (N39, N34);
nor NOR3 (N40, N24, N38, N20);
nand NAND4 (N41, N18, N20, N21, N39);
or OR4 (N42, N4, N12, N10, N37);
or OR4 (N43, N12, N18, N29, N14);
nor NOR2 (N44, N4, N8);
xor XOR2 (N45, N41, N43);
not NOT1 (N46, N21);
or OR4 (N47, N40, N26, N42, N40);
buf BUF1 (N48, N45);
buf BUF1 (N49, N46);
and AND3 (N50, N43, N24, N22);
and AND4 (N51, N23, N21, N21, N12);
not NOT1 (N52, N50);
xor XOR2 (N53, N48, N30);
nand NAND2 (N54, N32, N15);
nor NOR3 (N55, N31, N45, N40);
buf BUF1 (N56, N47);
xor XOR2 (N57, N51, N55);
buf BUF1 (N58, N44);
buf BUF1 (N59, N32);
and AND2 (N60, N52, N34);
not NOT1 (N61, N53);
nor NOR4 (N62, N28, N19, N32, N5);
xor XOR2 (N63, N60, N40);
xor XOR2 (N64, N62, N16);
nand NAND3 (N65, N59, N5, N24);
buf BUF1 (N66, N49);
nand NAND2 (N67, N58, N41);
buf BUF1 (N68, N63);
nand NAND4 (N69, N36, N30, N51, N32);
nor NOR2 (N70, N66, N22);
not NOT1 (N71, N65);
nand NAND3 (N72, N70, N60, N68);
xor XOR2 (N73, N38, N72);
nor NOR4 (N74, N41, N35, N35, N29);
or OR3 (N75, N69, N11, N34);
buf BUF1 (N76, N67);
nor NOR4 (N77, N74, N76, N32, N53);
nand NAND2 (N78, N11, N44);
xor XOR2 (N79, N57, N70);
nor NOR2 (N80, N77, N9);
nor NOR3 (N81, N75, N57, N54);
or OR2 (N82, N73, N39);
not NOT1 (N83, N42);
or OR3 (N84, N71, N39, N73);
nand NAND4 (N85, N84, N51, N32, N16);
buf BUF1 (N86, N61);
nor NOR4 (N87, N78, N73, N33, N42);
and AND3 (N88, N81, N17, N45);
nor NOR4 (N89, N88, N5, N31, N86);
nand NAND2 (N90, N68, N12);
xor XOR2 (N91, N64, N60);
not NOT1 (N92, N82);
buf BUF1 (N93, N56);
and AND3 (N94, N90, N2, N39);
nand NAND3 (N95, N92, N40, N5);
not NOT1 (N96, N87);
xor XOR2 (N97, N95, N85);
xor XOR2 (N98, N87, N11);
not NOT1 (N99, N93);
and AND2 (N100, N94, N51);
nor NOR2 (N101, N79, N48);
nor NOR2 (N102, N91, N15);
not NOT1 (N103, N101);
nor NOR4 (N104, N100, N43, N17, N89);
not NOT1 (N105, N38);
buf BUF1 (N106, N80);
nand NAND2 (N107, N97, N44);
xor XOR2 (N108, N105, N18);
or OR3 (N109, N83, N14, N61);
or OR2 (N110, N103, N3);
buf BUF1 (N111, N108);
not NOT1 (N112, N109);
nor NOR3 (N113, N104, N94, N34);
or OR2 (N114, N113, N3);
buf BUF1 (N115, N107);
and AND2 (N116, N96, N29);
nand NAND3 (N117, N112, N27, N60);
nor NOR3 (N118, N98, N64, N18);
and AND2 (N119, N110, N48);
nor NOR4 (N120, N117, N68, N2, N90);
buf BUF1 (N121, N120);
or OR4 (N122, N111, N3, N73, N110);
and AND4 (N123, N102, N59, N28, N69);
nor NOR4 (N124, N122, N107, N73, N45);
buf BUF1 (N125, N118);
nand NAND2 (N126, N119, N64);
nor NOR3 (N127, N106, N111, N11);
nor NOR2 (N128, N126, N111);
or OR4 (N129, N127, N97, N52, N84);
buf BUF1 (N130, N123);
nand NAND4 (N131, N125, N38, N104, N30);
buf BUF1 (N132, N130);
and AND3 (N133, N99, N107, N10);
or OR2 (N134, N114, N71);
and AND3 (N135, N121, N11, N106);
not NOT1 (N136, N132);
or OR2 (N137, N135, N95);
nor NOR3 (N138, N133, N131, N55);
nand NAND2 (N139, N88, N15);
and AND2 (N140, N134, N14);
and AND2 (N141, N140, N21);
and AND4 (N142, N128, N110, N123, N130);
nand NAND4 (N143, N137, N10, N83, N6);
or OR4 (N144, N141, N53, N90, N85);
nand NAND2 (N145, N115, N58);
nor NOR3 (N146, N143, N97, N95);
or OR4 (N147, N136, N132, N135, N111);
or OR3 (N148, N142, N67, N129);
or OR3 (N149, N47, N133, N7);
nand NAND2 (N150, N149, N27);
not NOT1 (N151, N144);
nand NAND4 (N152, N147, N150, N93, N122);
xor XOR2 (N153, N92, N147);
or OR4 (N154, N153, N97, N101, N80);
or OR3 (N155, N116, N20, N19);
and AND4 (N156, N124, N48, N135, N10);
buf BUF1 (N157, N146);
nor NOR4 (N158, N154, N84, N57, N21);
buf BUF1 (N159, N152);
or OR4 (N160, N159, N140, N12, N124);
buf BUF1 (N161, N151);
xor XOR2 (N162, N158, N131);
nand NAND4 (N163, N161, N123, N118, N91);
nand NAND4 (N164, N145, N63, N40, N128);
buf BUF1 (N165, N148);
nand NAND4 (N166, N163, N42, N38, N100);
buf BUF1 (N167, N156);
nand NAND4 (N168, N167, N99, N39, N130);
or OR2 (N169, N139, N48);
not NOT1 (N170, N169);
or OR4 (N171, N155, N24, N138, N15);
nor NOR3 (N172, N23, N45, N37);
and AND3 (N173, N164, N69, N56);
and AND4 (N174, N166, N164, N146, N59);
nand NAND4 (N175, N173, N92, N107, N61);
not NOT1 (N176, N174);
or OR4 (N177, N165, N94, N112, N5);
nand NAND3 (N178, N177, N137, N32);
xor XOR2 (N179, N171, N159);
nor NOR2 (N180, N172, N158);
xor XOR2 (N181, N176, N96);
nor NOR2 (N182, N175, N105);
nand NAND2 (N183, N157, N37);
xor XOR2 (N184, N179, N160);
xor XOR2 (N185, N135, N171);
not NOT1 (N186, N178);
xor XOR2 (N187, N168, N169);
nand NAND2 (N188, N162, N77);
nor NOR2 (N189, N181, N101);
xor XOR2 (N190, N184, N122);
xor XOR2 (N191, N185, N120);
and AND4 (N192, N189, N47, N4, N65);
xor XOR2 (N193, N170, N126);
and AND3 (N194, N180, N18, N83);
nor NOR4 (N195, N191, N59, N111, N110);
or OR4 (N196, N190, N65, N172, N62);
xor XOR2 (N197, N195, N189);
or OR2 (N198, N192, N82);
xor XOR2 (N199, N194, N92);
xor XOR2 (N200, N188, N10);
nand NAND3 (N201, N200, N132, N117);
xor XOR2 (N202, N187, N1);
nor NOR2 (N203, N182, N169);
or OR2 (N204, N199, N17);
and AND2 (N205, N196, N56);
xor XOR2 (N206, N198, N168);
xor XOR2 (N207, N205, N119);
nand NAND4 (N208, N197, N33, N24, N64);
and AND4 (N209, N203, N196, N171, N69);
not NOT1 (N210, N202);
or OR4 (N211, N186, N55, N147, N152);
nand NAND2 (N212, N206, N151);
xor XOR2 (N213, N212, N98);
buf BUF1 (N214, N208);
xor XOR2 (N215, N211, N127);
nand NAND2 (N216, N210, N105);
not NOT1 (N217, N207);
not NOT1 (N218, N214);
not NOT1 (N219, N193);
nor NOR2 (N220, N209, N16);
nand NAND2 (N221, N215, N125);
nor NOR2 (N222, N219, N158);
and AND2 (N223, N222, N55);
not NOT1 (N224, N217);
and AND2 (N225, N220, N6);
not NOT1 (N226, N225);
or OR4 (N227, N204, N178, N192, N83);
nor NOR4 (N228, N227, N187, N222, N30);
or OR3 (N229, N216, N81, N53);
or OR4 (N230, N183, N140, N194, N168);
nor NOR4 (N231, N223, N140, N9, N148);
or OR4 (N232, N228, N187, N194, N102);
nand NAND4 (N233, N213, N2, N41, N52);
xor XOR2 (N234, N221, N78);
not NOT1 (N235, N201);
buf BUF1 (N236, N226);
or OR3 (N237, N231, N197, N173);
xor XOR2 (N238, N233, N5);
and AND3 (N239, N224, N172, N158);
nor NOR2 (N240, N239, N52);
xor XOR2 (N241, N218, N11);
nand NAND2 (N242, N241, N88);
nand NAND3 (N243, N238, N212, N197);
or OR2 (N244, N242, N165);
not NOT1 (N245, N237);
xor XOR2 (N246, N236, N192);
not NOT1 (N247, N234);
buf BUF1 (N248, N245);
and AND2 (N249, N232, N45);
not NOT1 (N250, N240);
nor NOR3 (N251, N247, N75, N209);
nand NAND4 (N252, N251, N92, N127, N191);
not NOT1 (N253, N248);
or OR2 (N254, N246, N223);
nand NAND4 (N255, N254, N215, N46, N169);
nand NAND3 (N256, N253, N3, N49);
and AND3 (N257, N250, N127, N126);
nand NAND2 (N258, N229, N217);
xor XOR2 (N259, N258, N72);
or OR4 (N260, N244, N133, N209, N95);
not NOT1 (N261, N249);
buf BUF1 (N262, N256);
and AND3 (N263, N261, N61, N226);
nor NOR3 (N264, N252, N26, N221);
xor XOR2 (N265, N260, N49);
nor NOR4 (N266, N235, N81, N124, N23);
and AND2 (N267, N265, N23);
buf BUF1 (N268, N262);
nor NOR3 (N269, N243, N144, N19);
not NOT1 (N270, N267);
nand NAND3 (N271, N268, N175, N233);
xor XOR2 (N272, N266, N76);
xor XOR2 (N273, N257, N191);
or OR4 (N274, N271, N38, N241, N194);
nor NOR4 (N275, N263, N215, N168, N97);
nor NOR2 (N276, N269, N178);
and AND4 (N277, N259, N61, N185, N275);
not NOT1 (N278, N275);
xor XOR2 (N279, N277, N132);
nand NAND4 (N280, N273, N105, N106, N60);
nand NAND2 (N281, N279, N104);
nor NOR3 (N282, N272, N242, N61);
and AND4 (N283, N278, N111, N63, N5);
buf BUF1 (N284, N281);
xor XOR2 (N285, N283, N246);
or OR3 (N286, N282, N48, N74);
and AND4 (N287, N255, N133, N42, N90);
or OR2 (N288, N280, N223);
xor XOR2 (N289, N274, N208);
not NOT1 (N290, N230);
buf BUF1 (N291, N287);
or OR2 (N292, N264, N2);
buf BUF1 (N293, N291);
nand NAND3 (N294, N284, N196, N57);
buf BUF1 (N295, N289);
buf BUF1 (N296, N270);
not NOT1 (N297, N286);
or OR4 (N298, N292, N91, N254, N85);
not NOT1 (N299, N298);
or OR4 (N300, N294, N28, N45, N266);
xor XOR2 (N301, N295, N210);
nor NOR2 (N302, N285, N218);
buf BUF1 (N303, N301);
and AND2 (N304, N296, N83);
xor XOR2 (N305, N302, N87);
and AND2 (N306, N300, N76);
or OR3 (N307, N306, N306, N153);
or OR4 (N308, N304, N3, N78, N258);
or OR3 (N309, N288, N227, N161);
nand NAND2 (N310, N299, N152);
xor XOR2 (N311, N310, N175);
and AND3 (N312, N290, N5, N207);
nand NAND3 (N313, N307, N251, N118);
nand NAND2 (N314, N276, N38);
and AND2 (N315, N314, N160);
nand NAND3 (N316, N309, N156, N194);
or OR2 (N317, N297, N169);
or OR3 (N318, N317, N33, N98);
or OR2 (N319, N318, N88);
not NOT1 (N320, N312);
or OR3 (N321, N313, N25, N299);
nor NOR2 (N322, N315, N194);
nand NAND3 (N323, N293, N35, N315);
or OR2 (N324, N320, N212);
xor XOR2 (N325, N321, N7);
and AND4 (N326, N308, N192, N200, N276);
buf BUF1 (N327, N322);
xor XOR2 (N328, N311, N301);
not NOT1 (N329, N325);
not NOT1 (N330, N305);
and AND4 (N331, N323, N295, N55, N173);
or OR4 (N332, N326, N137, N70, N149);
or OR4 (N333, N332, N133, N310, N300);
not NOT1 (N334, N333);
buf BUF1 (N335, N328);
nand NAND2 (N336, N327, N138);
not NOT1 (N337, N330);
nor NOR2 (N338, N329, N297);
nor NOR3 (N339, N336, N301, N134);
and AND4 (N340, N324, N232, N34, N123);
or OR3 (N341, N331, N248, N171);
buf BUF1 (N342, N340);
and AND3 (N343, N319, N332, N280);
not NOT1 (N344, N335);
not NOT1 (N345, N337);
nor NOR3 (N346, N339, N291, N3);
nand NAND3 (N347, N342, N259, N195);
and AND2 (N348, N344, N130);
nand NAND3 (N349, N347, N3, N323);
nor NOR2 (N350, N303, N15);
not NOT1 (N351, N334);
xor XOR2 (N352, N351, N291);
nand NAND3 (N353, N349, N104, N76);
not NOT1 (N354, N350);
buf BUF1 (N355, N338);
and AND4 (N356, N352, N22, N216, N326);
buf BUF1 (N357, N348);
nor NOR2 (N358, N316, N138);
xor XOR2 (N359, N356, N165);
nand NAND2 (N360, N343, N54);
xor XOR2 (N361, N353, N161);
xor XOR2 (N362, N354, N185);
nand NAND3 (N363, N341, N180, N233);
not NOT1 (N364, N346);
not NOT1 (N365, N357);
nand NAND4 (N366, N361, N38, N279, N129);
or OR2 (N367, N362, N173);
not NOT1 (N368, N364);
or OR4 (N369, N363, N52, N88, N24);
and AND3 (N370, N360, N215, N105);
nand NAND4 (N371, N365, N56, N115, N23);
or OR4 (N372, N355, N149, N120, N253);
nor NOR2 (N373, N366, N362);
nor NOR2 (N374, N359, N48);
and AND2 (N375, N367, N82);
buf BUF1 (N376, N369);
buf BUF1 (N377, N358);
or OR3 (N378, N373, N365, N122);
not NOT1 (N379, N370);
nand NAND4 (N380, N371, N61, N168, N170);
or OR2 (N381, N380, N105);
xor XOR2 (N382, N345, N214);
xor XOR2 (N383, N381, N251);
and AND2 (N384, N376, N126);
buf BUF1 (N385, N374);
or OR2 (N386, N377, N310);
nand NAND2 (N387, N372, N77);
and AND2 (N388, N383, N220);
not NOT1 (N389, N387);
and AND4 (N390, N388, N64, N174, N3);
and AND4 (N391, N390, N295, N368, N342);
or OR4 (N392, N339, N31, N171, N262);
not NOT1 (N393, N392);
nand NAND4 (N394, N386, N184, N326, N234);
xor XOR2 (N395, N375, N36);
nand NAND3 (N396, N379, N280, N176);
buf BUF1 (N397, N395);
nand NAND3 (N398, N394, N353, N122);
or OR4 (N399, N396, N192, N25, N370);
or OR2 (N400, N384, N22);
or OR2 (N401, N399, N242);
not NOT1 (N402, N391);
and AND3 (N403, N385, N90, N141);
and AND4 (N404, N397, N230, N287, N252);
xor XOR2 (N405, N402, N351);
nand NAND4 (N406, N405, N60, N227, N66);
nand NAND4 (N407, N382, N385, N285, N162);
buf BUF1 (N408, N401);
not NOT1 (N409, N398);
or OR4 (N410, N393, N202, N281, N122);
nor NOR2 (N411, N389, N38);
nand NAND2 (N412, N400, N296);
not NOT1 (N413, N411);
or OR3 (N414, N409, N225, N153);
nand NAND2 (N415, N406, N364);
or OR4 (N416, N413, N185, N315, N85);
buf BUF1 (N417, N412);
nand NAND2 (N418, N407, N38);
xor XOR2 (N419, N408, N180);
xor XOR2 (N420, N415, N34);
or OR2 (N421, N418, N95);
and AND2 (N422, N410, N366);
not NOT1 (N423, N417);
buf BUF1 (N424, N403);
nor NOR4 (N425, N404, N249, N238, N268);
nand NAND3 (N426, N416, N404, N29);
or OR2 (N427, N422, N336);
buf BUF1 (N428, N414);
or OR2 (N429, N419, N427);
nand NAND4 (N430, N81, N21, N136, N156);
nand NAND2 (N431, N420, N359);
buf BUF1 (N432, N424);
or OR3 (N433, N428, N292, N406);
not NOT1 (N434, N430);
and AND4 (N435, N426, N272, N295, N380);
xor XOR2 (N436, N435, N37);
nand NAND2 (N437, N434, N292);
buf BUF1 (N438, N378);
nand NAND2 (N439, N423, N62);
or OR4 (N440, N421, N206, N390, N141);
buf BUF1 (N441, N425);
not NOT1 (N442, N438);
buf BUF1 (N443, N437);
nor NOR2 (N444, N433, N53);
and AND4 (N445, N440, N79, N306, N214);
or OR2 (N446, N445, N383);
xor XOR2 (N447, N446, N377);
not NOT1 (N448, N431);
nand NAND4 (N449, N439, N376, N124, N153);
or OR2 (N450, N442, N65);
and AND3 (N451, N441, N405, N439);
nand NAND2 (N452, N432, N175);
buf BUF1 (N453, N444);
and AND2 (N454, N448, N67);
nor NOR2 (N455, N447, N410);
buf BUF1 (N456, N451);
not NOT1 (N457, N453);
buf BUF1 (N458, N457);
xor XOR2 (N459, N436, N204);
nand NAND4 (N460, N459, N365, N158, N220);
nor NOR2 (N461, N449, N176);
and AND3 (N462, N443, N110, N245);
nor NOR4 (N463, N456, N35, N430, N285);
or OR2 (N464, N455, N381);
not NOT1 (N465, N461);
buf BUF1 (N466, N465);
xor XOR2 (N467, N466, N50);
nor NOR3 (N468, N454, N65, N303);
and AND4 (N469, N458, N427, N376, N416);
nor NOR2 (N470, N429, N438);
not NOT1 (N471, N460);
or OR4 (N472, N463, N400, N45, N354);
and AND4 (N473, N468, N281, N83, N61);
nor NOR3 (N474, N467, N189, N17);
nand NAND2 (N475, N474, N55);
buf BUF1 (N476, N475);
buf BUF1 (N477, N462);
nor NOR2 (N478, N450, N108);
buf BUF1 (N479, N472);
or OR4 (N480, N471, N436, N395, N205);
buf BUF1 (N481, N464);
xor XOR2 (N482, N477, N368);
not NOT1 (N483, N479);
buf BUF1 (N484, N473);
buf BUF1 (N485, N483);
and AND4 (N486, N452, N336, N5, N290);
buf BUF1 (N487, N469);
not NOT1 (N488, N482);
and AND2 (N489, N476, N305);
or OR3 (N490, N486, N430, N100);
nor NOR4 (N491, N470, N354, N92, N319);
xor XOR2 (N492, N490, N453);
buf BUF1 (N493, N485);
xor XOR2 (N494, N484, N267);
xor XOR2 (N495, N481, N492);
or OR2 (N496, N45, N19);
nand NAND2 (N497, N491, N78);
nand NAND4 (N498, N494, N399, N317, N421);
nand NAND2 (N499, N498, N55);
nor NOR3 (N500, N496, N145, N42);
or OR2 (N501, N487, N50);
xor XOR2 (N502, N478, N476);
or OR2 (N503, N495, N72);
nand NAND2 (N504, N503, N462);
xor XOR2 (N505, N493, N122);
and AND3 (N506, N480, N22, N118);
nand NAND3 (N507, N504, N367, N356);
and AND3 (N508, N489, N304, N396);
nor NOR3 (N509, N505, N12, N187);
buf BUF1 (N510, N500);
and AND2 (N511, N502, N422);
nor NOR4 (N512, N510, N487, N393, N439);
nand NAND4 (N513, N506, N76, N404, N391);
and AND2 (N514, N501, N393);
not NOT1 (N515, N488);
or OR2 (N516, N511, N68);
and AND3 (N517, N515, N200, N420);
nand NAND3 (N518, N514, N218, N98);
nor NOR2 (N519, N517, N42);
buf BUF1 (N520, N512);
and AND2 (N521, N508, N71);
nor NOR4 (N522, N518, N268, N384, N421);
not NOT1 (N523, N521);
and AND4 (N524, N509, N152, N276, N347);
or OR3 (N525, N519, N268, N156);
not NOT1 (N526, N507);
and AND3 (N527, N497, N311, N377);
nand NAND2 (N528, N524, N184);
or OR4 (N529, N522, N38, N32, N523);
buf BUF1 (N530, N104);
nor NOR4 (N531, N513, N230, N525, N166);
and AND3 (N532, N346, N117, N204);
buf BUF1 (N533, N532);
and AND2 (N534, N531, N264);
buf BUF1 (N535, N530);
nor NOR2 (N536, N526, N263);
buf BUF1 (N537, N533);
nand NAND3 (N538, N529, N142, N84);
and AND3 (N539, N516, N265, N415);
or OR3 (N540, N499, N190, N380);
buf BUF1 (N541, N535);
nor NOR3 (N542, N520, N285, N464);
nor NOR2 (N543, N541, N334);
or OR2 (N544, N534, N234);
nand NAND3 (N545, N540, N352, N179);
xor XOR2 (N546, N539, N242);
or OR4 (N547, N537, N342, N490, N47);
and AND3 (N548, N547, N40, N296);
nand NAND4 (N549, N542, N400, N269, N40);
or OR3 (N550, N544, N74, N292);
buf BUF1 (N551, N548);
or OR3 (N552, N527, N141, N495);
nor NOR4 (N553, N528, N266, N494, N5);
not NOT1 (N554, N552);
buf BUF1 (N555, N546);
xor XOR2 (N556, N555, N426);
and AND3 (N557, N543, N441, N192);
or OR3 (N558, N557, N292, N220);
nand NAND2 (N559, N536, N283);
nor NOR4 (N560, N549, N484, N337, N246);
not NOT1 (N561, N559);
buf BUF1 (N562, N545);
or OR2 (N563, N551, N166);
or OR4 (N564, N550, N219, N179, N279);
and AND3 (N565, N553, N160, N452);
not NOT1 (N566, N565);
nor NOR2 (N567, N556, N410);
xor XOR2 (N568, N560, N85);
nor NOR4 (N569, N568, N53, N352, N290);
not NOT1 (N570, N566);
buf BUF1 (N571, N569);
nor NOR4 (N572, N538, N49, N259, N180);
xor XOR2 (N573, N567, N392);
or OR3 (N574, N563, N143, N359);
not NOT1 (N575, N573);
and AND4 (N576, N554, N392, N556, N340);
not NOT1 (N577, N570);
nand NAND3 (N578, N577, N147, N455);
or OR2 (N579, N564, N440);
buf BUF1 (N580, N571);
nor NOR3 (N581, N576, N246, N186);
not NOT1 (N582, N572);
nand NAND4 (N583, N558, N50, N287, N246);
and AND2 (N584, N580, N211);
and AND4 (N585, N561, N185, N156, N556);
buf BUF1 (N586, N579);
buf BUF1 (N587, N581);
nor NOR3 (N588, N575, N169, N100);
not NOT1 (N589, N583);
nor NOR2 (N590, N578, N193);
buf BUF1 (N591, N584);
or OR2 (N592, N582, N15);
not NOT1 (N593, N585);
not NOT1 (N594, N574);
or OR4 (N595, N589, N457, N458, N392);
or OR2 (N596, N587, N220);
xor XOR2 (N597, N562, N286);
or OR3 (N598, N594, N575, N166);
nand NAND3 (N599, N591, N575, N482);
buf BUF1 (N600, N586);
xor XOR2 (N601, N588, N278);
or OR3 (N602, N596, N483, N243);
and AND2 (N603, N590, N437);
or OR2 (N604, N598, N554);
nor NOR3 (N605, N604, N303, N89);
xor XOR2 (N606, N599, N491);
nand NAND2 (N607, N602, N541);
and AND4 (N608, N603, N102, N387, N343);
buf BUF1 (N609, N607);
or OR2 (N610, N601, N587);
and AND3 (N611, N592, N122, N403);
buf BUF1 (N612, N610);
and AND4 (N613, N593, N83, N566, N409);
and AND4 (N614, N595, N348, N537, N450);
and AND4 (N615, N605, N498, N53, N558);
and AND3 (N616, N611, N32, N268);
nand NAND3 (N617, N612, N329, N610);
nor NOR2 (N618, N617, N350);
nor NOR4 (N619, N597, N250, N76, N71);
nand NAND4 (N620, N613, N586, N60, N547);
buf BUF1 (N621, N619);
or OR2 (N622, N608, N5);
xor XOR2 (N623, N615, N497);
or OR2 (N624, N620, N311);
or OR3 (N625, N624, N583, N362);
nor NOR3 (N626, N616, N234, N316);
and AND4 (N627, N622, N525, N495, N186);
or OR4 (N628, N618, N26, N439, N242);
nor NOR4 (N629, N628, N511, N413, N189);
or OR2 (N630, N627, N356);
nand NAND3 (N631, N626, N516, N485);
not NOT1 (N632, N609);
buf BUF1 (N633, N621);
or OR3 (N634, N625, N573, N63);
or OR3 (N635, N632, N20, N271);
nor NOR2 (N636, N633, N351);
or OR2 (N637, N636, N362);
xor XOR2 (N638, N623, N631);
xor XOR2 (N639, N279, N53);
nand NAND4 (N640, N630, N223, N86, N509);
nand NAND3 (N641, N629, N26, N544);
buf BUF1 (N642, N635);
not NOT1 (N643, N638);
buf BUF1 (N644, N643);
not NOT1 (N645, N614);
nand NAND2 (N646, N637, N612);
buf BUF1 (N647, N639);
nor NOR2 (N648, N600, N445);
xor XOR2 (N649, N634, N201);
and AND2 (N650, N606, N333);
nor NOR2 (N651, N650, N646);
and AND4 (N652, N16, N77, N38, N119);
nand NAND2 (N653, N649, N552);
xor XOR2 (N654, N644, N523);
and AND2 (N655, N642, N412);
and AND2 (N656, N654, N163);
not NOT1 (N657, N656);
xor XOR2 (N658, N655, N33);
xor XOR2 (N659, N645, N584);
nor NOR3 (N660, N657, N619, N314);
buf BUF1 (N661, N640);
buf BUF1 (N662, N647);
buf BUF1 (N663, N658);
nor NOR2 (N664, N653, N578);
nor NOR3 (N665, N661, N372, N211);
or OR2 (N666, N641, N118);
buf BUF1 (N667, N651);
nand NAND2 (N668, N665, N555);
not NOT1 (N669, N660);
xor XOR2 (N670, N659, N228);
xor XOR2 (N671, N667, N415);
or OR3 (N672, N662, N270, N152);
or OR3 (N673, N666, N535, N41);
buf BUF1 (N674, N664);
nand NAND4 (N675, N663, N268, N17, N533);
or OR3 (N676, N674, N239, N201);
xor XOR2 (N677, N673, N542);
not NOT1 (N678, N669);
nand NAND2 (N679, N678, N504);
nand NAND3 (N680, N652, N205, N367);
xor XOR2 (N681, N679, N148);
nand NAND4 (N682, N676, N347, N427, N624);
or OR4 (N683, N680, N582, N289, N138);
and AND4 (N684, N671, N573, N308, N328);
or OR2 (N685, N677, N409);
and AND2 (N686, N682, N611);
nor NOR2 (N687, N672, N217);
buf BUF1 (N688, N685);
not NOT1 (N689, N668);
buf BUF1 (N690, N681);
or OR2 (N691, N688, N53);
not NOT1 (N692, N691);
or OR4 (N693, N689, N353, N426, N69);
nor NOR2 (N694, N648, N611);
not NOT1 (N695, N692);
not NOT1 (N696, N675);
not NOT1 (N697, N687);
or OR2 (N698, N694, N73);
and AND3 (N699, N690, N632, N428);
nand NAND4 (N700, N693, N139, N6, N302);
buf BUF1 (N701, N697);
nor NOR3 (N702, N698, N139, N611);
buf BUF1 (N703, N699);
or OR3 (N704, N686, N62, N439);
buf BUF1 (N705, N702);
not NOT1 (N706, N695);
buf BUF1 (N707, N683);
xor XOR2 (N708, N700, N65);
buf BUF1 (N709, N696);
buf BUF1 (N710, N701);
not NOT1 (N711, N704);
buf BUF1 (N712, N684);
or OR4 (N713, N712, N391, N458, N649);
buf BUF1 (N714, N703);
and AND2 (N715, N707, N652);
nor NOR4 (N716, N706, N291, N197, N72);
or OR4 (N717, N708, N177, N283, N241);
or OR4 (N718, N715, N456, N611, N595);
or OR2 (N719, N709, N172);
buf BUF1 (N720, N713);
nor NOR4 (N721, N718, N522, N660, N628);
and AND3 (N722, N705, N250, N6);
nand NAND2 (N723, N710, N561);
nand NAND4 (N724, N716, N542, N235, N328);
nand NAND4 (N725, N717, N724, N614, N277);
nor NOR3 (N726, N50, N146, N261);
not NOT1 (N727, N670);
buf BUF1 (N728, N721);
nor NOR3 (N729, N727, N297, N317);
and AND4 (N730, N725, N207, N192, N587);
nor NOR4 (N731, N729, N551, N167, N86);
nor NOR4 (N732, N711, N340, N331, N532);
xor XOR2 (N733, N731, N537);
not NOT1 (N734, N723);
nand NAND4 (N735, N714, N577, N530, N26);
nand NAND4 (N736, N735, N67, N145, N168);
nor NOR4 (N737, N734, N702, N145, N713);
nor NOR3 (N738, N726, N676, N618);
xor XOR2 (N739, N728, N495);
and AND2 (N740, N736, N701);
xor XOR2 (N741, N732, N648);
buf BUF1 (N742, N722);
buf BUF1 (N743, N730);
or OR4 (N744, N733, N264, N555, N467);
and AND4 (N745, N744, N601, N435, N521);
and AND4 (N746, N720, N634, N53, N227);
xor XOR2 (N747, N740, N180);
buf BUF1 (N748, N719);
buf BUF1 (N749, N737);
or OR4 (N750, N743, N614, N479, N351);
xor XOR2 (N751, N738, N657);
xor XOR2 (N752, N747, N396);
buf BUF1 (N753, N741);
buf BUF1 (N754, N752);
and AND4 (N755, N750, N610, N492, N132);
and AND2 (N756, N745, N263);
nand NAND4 (N757, N754, N694, N681, N214);
xor XOR2 (N758, N746, N394);
or OR4 (N759, N742, N621, N580, N136);
or OR3 (N760, N739, N501, N202);
xor XOR2 (N761, N760, N743);
and AND3 (N762, N756, N133, N570);
buf BUF1 (N763, N749);
nor NOR4 (N764, N758, N153, N465, N224);
buf BUF1 (N765, N755);
or OR2 (N766, N765, N378);
buf BUF1 (N767, N748);
nand NAND4 (N768, N763, N82, N761, N503);
buf BUF1 (N769, N73);
and AND4 (N770, N753, N189, N474, N559);
and AND3 (N771, N759, N137, N459);
and AND3 (N772, N771, N337, N521);
nor NOR4 (N773, N764, N414, N267, N148);
xor XOR2 (N774, N768, N21);
nand NAND4 (N775, N766, N119, N148, N2);
nand NAND4 (N776, N751, N6, N425, N29);
not NOT1 (N777, N770);
nor NOR4 (N778, N773, N249, N412, N563);
nor NOR3 (N779, N767, N40, N209);
nor NOR3 (N780, N774, N634, N28);
nor NOR3 (N781, N776, N428, N445);
nor NOR3 (N782, N762, N706, N487);
xor XOR2 (N783, N777, N412);
xor XOR2 (N784, N781, N608);
and AND2 (N785, N780, N267);
buf BUF1 (N786, N784);
not NOT1 (N787, N785);
not NOT1 (N788, N786);
or OR2 (N789, N775, N137);
buf BUF1 (N790, N772);
nand NAND3 (N791, N779, N588, N34);
xor XOR2 (N792, N791, N348);
nand NAND2 (N793, N787, N686);
or OR2 (N794, N793, N225);
nor NOR3 (N795, N757, N174, N487);
nand NAND4 (N796, N789, N342, N437, N156);
nand NAND2 (N797, N792, N256);
nand NAND4 (N798, N794, N2, N497, N354);
nor NOR3 (N799, N798, N235, N60);
or OR3 (N800, N795, N362, N612);
and AND2 (N801, N783, N544);
xor XOR2 (N802, N799, N166);
nor NOR3 (N803, N797, N621, N177);
or OR2 (N804, N796, N138);
or OR2 (N805, N782, N384);
or OR2 (N806, N788, N709);
and AND2 (N807, N806, N221);
and AND3 (N808, N803, N160, N9);
or OR3 (N809, N807, N402, N519);
buf BUF1 (N810, N778);
xor XOR2 (N811, N790, N655);
xor XOR2 (N812, N808, N196);
buf BUF1 (N813, N812);
xor XOR2 (N814, N811, N795);
xor XOR2 (N815, N804, N512);
or OR3 (N816, N814, N39, N583);
nor NOR4 (N817, N800, N300, N57, N147);
or OR2 (N818, N769, N713);
xor XOR2 (N819, N810, N347);
not NOT1 (N820, N818);
nand NAND3 (N821, N809, N587, N638);
buf BUF1 (N822, N821);
and AND2 (N823, N802, N361);
or OR4 (N824, N823, N106, N663, N682);
buf BUF1 (N825, N805);
or OR4 (N826, N816, N23, N528, N114);
or OR4 (N827, N813, N380, N97, N9);
buf BUF1 (N828, N817);
nor NOR3 (N829, N827, N670, N14);
not NOT1 (N830, N828);
buf BUF1 (N831, N815);
and AND4 (N832, N820, N797, N81, N539);
buf BUF1 (N833, N826);
xor XOR2 (N834, N801, N723);
and AND4 (N835, N830, N205, N771, N349);
xor XOR2 (N836, N822, N592);
xor XOR2 (N837, N829, N310);
and AND2 (N838, N825, N101);
xor XOR2 (N839, N824, N775);
and AND3 (N840, N838, N187, N476);
nor NOR3 (N841, N836, N668, N546);
buf BUF1 (N842, N831);
and AND2 (N843, N837, N796);
or OR2 (N844, N839, N127);
nand NAND2 (N845, N842, N541);
buf BUF1 (N846, N832);
not NOT1 (N847, N845);
and AND2 (N848, N833, N628);
nand NAND3 (N849, N848, N610, N800);
nand NAND2 (N850, N841, N274);
not NOT1 (N851, N840);
not NOT1 (N852, N844);
nor NOR2 (N853, N846, N813);
nor NOR3 (N854, N851, N452, N236);
and AND4 (N855, N843, N9, N600, N333);
not NOT1 (N856, N834);
xor XOR2 (N857, N854, N831);
nor NOR2 (N858, N849, N460);
not NOT1 (N859, N835);
buf BUF1 (N860, N856);
and AND3 (N861, N847, N169, N546);
nor NOR2 (N862, N857, N636);
and AND4 (N863, N860, N455, N629, N415);
buf BUF1 (N864, N819);
or OR4 (N865, N858, N210, N495, N714);
or OR2 (N866, N863, N42);
not NOT1 (N867, N850);
nand NAND3 (N868, N862, N729, N686);
buf BUF1 (N869, N855);
or OR2 (N870, N859, N268);
and AND2 (N871, N852, N818);
nor NOR4 (N872, N868, N772, N348, N473);
or OR4 (N873, N871, N865, N716, N830);
not NOT1 (N874, N406);
and AND2 (N875, N866, N747);
or OR4 (N876, N870, N601, N227, N358);
xor XOR2 (N877, N869, N629);
or OR2 (N878, N864, N595);
not NOT1 (N879, N872);
xor XOR2 (N880, N878, N768);
xor XOR2 (N881, N877, N736);
not NOT1 (N882, N861);
not NOT1 (N883, N867);
or OR4 (N884, N880, N157, N367, N778);
or OR3 (N885, N884, N504, N754);
not NOT1 (N886, N874);
buf BUF1 (N887, N881);
nand NAND4 (N888, N853, N161, N434, N297);
nor NOR4 (N889, N875, N66, N824, N285);
nand NAND4 (N890, N885, N868, N762, N844);
not NOT1 (N891, N882);
nor NOR2 (N892, N873, N255);
nor NOR4 (N893, N876, N876, N77, N235);
nor NOR2 (N894, N892, N627);
nor NOR3 (N895, N879, N733, N229);
xor XOR2 (N896, N893, N381);
or OR3 (N897, N894, N394, N342);
xor XOR2 (N898, N886, N694);
buf BUF1 (N899, N887);
or OR3 (N900, N888, N591, N496);
nor NOR3 (N901, N896, N254, N134);
or OR3 (N902, N891, N430, N605);
not NOT1 (N903, N898);
and AND4 (N904, N900, N228, N435, N202);
or OR2 (N905, N902, N403);
nand NAND4 (N906, N899, N901, N306, N774);
or OR3 (N907, N328, N248, N55);
nor NOR3 (N908, N907, N137, N600);
not NOT1 (N909, N906);
not NOT1 (N910, N889);
nor NOR4 (N911, N905, N76, N93, N37);
and AND2 (N912, N895, N371);
or OR4 (N913, N890, N830, N694, N466);
nand NAND2 (N914, N903, N207);
not NOT1 (N915, N912);
and AND3 (N916, N910, N645, N224);
or OR4 (N917, N913, N549, N338, N364);
or OR3 (N918, N883, N900, N803);
or OR3 (N919, N897, N521, N294);
and AND4 (N920, N918, N769, N575, N816);
nor NOR4 (N921, N904, N434, N516, N425);
and AND4 (N922, N914, N308, N395, N515);
and AND2 (N923, N920, N104);
buf BUF1 (N924, N923);
nand NAND3 (N925, N917, N639, N497);
not NOT1 (N926, N911);
nor NOR4 (N927, N924, N880, N528, N164);
not NOT1 (N928, N927);
xor XOR2 (N929, N925, N39);
and AND2 (N930, N921, N473);
buf BUF1 (N931, N922);
not NOT1 (N932, N916);
xor XOR2 (N933, N932, N758);
nor NOR3 (N934, N909, N488, N389);
not NOT1 (N935, N931);
nor NOR2 (N936, N929, N620);
not NOT1 (N937, N915);
xor XOR2 (N938, N934, N84);
or OR2 (N939, N919, N877);
not NOT1 (N940, N937);
buf BUF1 (N941, N928);
and AND2 (N942, N938, N553);
xor XOR2 (N943, N926, N861);
nand NAND3 (N944, N943, N783, N915);
nor NOR3 (N945, N941, N703, N852);
or OR2 (N946, N940, N141);
nand NAND3 (N947, N939, N99, N395);
or OR4 (N948, N930, N357, N113, N876);
and AND3 (N949, N947, N407, N636);
and AND4 (N950, N933, N310, N66, N753);
nand NAND3 (N951, N908, N706, N672);
and AND3 (N952, N936, N212, N258);
and AND3 (N953, N949, N726, N546);
buf BUF1 (N954, N944);
or OR3 (N955, N954, N818, N431);
or OR2 (N956, N950, N49);
nor NOR3 (N957, N955, N359, N535);
nor NOR4 (N958, N956, N497, N339, N211);
buf BUF1 (N959, N952);
or OR4 (N960, N946, N55, N353, N48);
or OR2 (N961, N953, N414);
nor NOR4 (N962, N959, N332, N432, N762);
xor XOR2 (N963, N935, N496);
nand NAND4 (N964, N945, N725, N314, N252);
not NOT1 (N965, N951);
not NOT1 (N966, N961);
nor NOR3 (N967, N964, N627, N306);
and AND2 (N968, N966, N155);
or OR3 (N969, N948, N192, N246);
and AND4 (N970, N965, N183, N969, N875);
nand NAND4 (N971, N852, N24, N94, N200);
xor XOR2 (N972, N967, N794);
or OR2 (N973, N972, N96);
and AND4 (N974, N957, N212, N160, N478);
and AND3 (N975, N973, N441, N335);
or OR4 (N976, N970, N248, N253, N448);
and AND2 (N977, N976, N502);
or OR2 (N978, N942, N543);
not NOT1 (N979, N975);
nor NOR2 (N980, N978, N515);
buf BUF1 (N981, N971);
nand NAND3 (N982, N963, N686, N818);
not NOT1 (N983, N981);
nor NOR4 (N984, N974, N713, N437, N199);
and AND2 (N985, N962, N68);
or OR3 (N986, N968, N589, N364);
nor NOR4 (N987, N982, N438, N766, N378);
xor XOR2 (N988, N984, N705);
buf BUF1 (N989, N985);
or OR3 (N990, N960, N130, N385);
and AND2 (N991, N980, N790);
xor XOR2 (N992, N977, N298);
or OR4 (N993, N990, N477, N987, N662);
nor NOR2 (N994, N96, N145);
and AND2 (N995, N993, N909);
and AND3 (N996, N994, N484, N545);
xor XOR2 (N997, N983, N626);
and AND4 (N998, N979, N790, N311, N935);
nand NAND3 (N999, N996, N187, N704);
buf BUF1 (N1000, N958);
nand NAND4 (N1001, N999, N101, N122, N467);
nor NOR2 (N1002, N988, N151);
nand NAND2 (N1003, N1002, N540);
and AND2 (N1004, N1000, N395);
nor NOR2 (N1005, N992, N973);
not NOT1 (N1006, N1005);
or OR4 (N1007, N1001, N311, N770, N73);
buf BUF1 (N1008, N991);
buf BUF1 (N1009, N1003);
and AND4 (N1010, N997, N729, N346, N446);
buf BUF1 (N1011, N1004);
or OR3 (N1012, N1009, N397, N467);
buf BUF1 (N1013, N1011);
not NOT1 (N1014, N1008);
or OR4 (N1015, N1014, N441, N698, N201);
nand NAND4 (N1016, N1007, N288, N286, N814);
and AND2 (N1017, N1013, N510);
or OR2 (N1018, N1012, N226);
xor XOR2 (N1019, N1016, N113);
buf BUF1 (N1020, N1017);
nand NAND4 (N1021, N1020, N46, N68, N283);
or OR4 (N1022, N995, N990, N62, N886);
and AND2 (N1023, N1010, N592);
buf BUF1 (N1024, N1023);
nor NOR2 (N1025, N989, N919);
and AND2 (N1026, N1018, N739);
buf BUF1 (N1027, N1022);
not NOT1 (N1028, N1024);
buf BUF1 (N1029, N998);
and AND3 (N1030, N1029, N371, N379);
not NOT1 (N1031, N1028);
and AND2 (N1032, N1025, N224);
or OR3 (N1033, N1030, N1004, N881);
or OR3 (N1034, N1019, N511, N142);
xor XOR2 (N1035, N1006, N36);
buf BUF1 (N1036, N1015);
xor XOR2 (N1037, N1035, N821);
or OR4 (N1038, N1031, N399, N38, N755);
and AND4 (N1039, N1021, N700, N885, N805);
buf BUF1 (N1040, N986);
or OR3 (N1041, N1037, N956, N186);
and AND2 (N1042, N1027, N468);
nor NOR4 (N1043, N1038, N656, N325, N285);
or OR3 (N1044, N1042, N175, N693);
xor XOR2 (N1045, N1032, N235);
nand NAND2 (N1046, N1039, N1040);
nand NAND4 (N1047, N173, N739, N628, N831);
not NOT1 (N1048, N1047);
not NOT1 (N1049, N1043);
buf BUF1 (N1050, N1045);
or OR2 (N1051, N1041, N883);
nor NOR2 (N1052, N1033, N902);
xor XOR2 (N1053, N1044, N837);
and AND3 (N1054, N1051, N47, N285);
xor XOR2 (N1055, N1049, N81);
nand NAND3 (N1056, N1055, N193, N1025);
xor XOR2 (N1057, N1056, N340);
and AND2 (N1058, N1026, N283);
xor XOR2 (N1059, N1057, N277);
buf BUF1 (N1060, N1050);
xor XOR2 (N1061, N1054, N141);
xor XOR2 (N1062, N1034, N10);
nor NOR3 (N1063, N1061, N696, N918);
nor NOR3 (N1064, N1048, N441, N440);
buf BUF1 (N1065, N1063);
or OR4 (N1066, N1060, N1011, N158, N689);
and AND3 (N1067, N1062, N614, N825);
not NOT1 (N1068, N1065);
or OR2 (N1069, N1068, N653);
nor NOR3 (N1070, N1069, N365, N224);
and AND2 (N1071, N1059, N849);
nand NAND4 (N1072, N1053, N828, N609, N114);
not NOT1 (N1073, N1064);
or OR3 (N1074, N1072, N120, N107);
and AND3 (N1075, N1058, N195, N580);
buf BUF1 (N1076, N1067);
or OR4 (N1077, N1071, N24, N250, N370);
buf BUF1 (N1078, N1073);
nand NAND4 (N1079, N1075, N781, N931, N1064);
not NOT1 (N1080, N1074);
xor XOR2 (N1081, N1079, N1080);
xor XOR2 (N1082, N993, N803);
not NOT1 (N1083, N1046);
nor NOR3 (N1084, N1077, N679, N54);
or OR3 (N1085, N1083, N389, N639);
or OR4 (N1086, N1078, N1035, N218, N1037);
and AND4 (N1087, N1086, N681, N934, N843);
nand NAND3 (N1088, N1076, N958, N773);
buf BUF1 (N1089, N1082);
nor NOR2 (N1090, N1085, N992);
nand NAND3 (N1091, N1084, N421, N862);
buf BUF1 (N1092, N1091);
not NOT1 (N1093, N1088);
or OR4 (N1094, N1052, N885, N372, N526);
or OR3 (N1095, N1036, N797, N551);
not NOT1 (N1096, N1092);
not NOT1 (N1097, N1070);
and AND2 (N1098, N1097, N1032);
not NOT1 (N1099, N1087);
buf BUF1 (N1100, N1098);
nor NOR4 (N1101, N1089, N945, N143, N1000);
xor XOR2 (N1102, N1081, N530);
and AND2 (N1103, N1096, N399);
xor XOR2 (N1104, N1099, N281);
and AND3 (N1105, N1100, N756, N243);
and AND4 (N1106, N1090, N657, N50, N351);
nand NAND2 (N1107, N1103, N968);
nor NOR4 (N1108, N1101, N172, N348, N977);
buf BUF1 (N1109, N1102);
xor XOR2 (N1110, N1093, N631);
or OR4 (N1111, N1066, N1090, N548, N581);
and AND3 (N1112, N1110, N579, N572);
and AND3 (N1113, N1095, N160, N248);
and AND3 (N1114, N1107, N465, N583);
nand NAND3 (N1115, N1094, N450, N351);
nand NAND3 (N1116, N1113, N150, N633);
nand NAND4 (N1117, N1106, N268, N792, N894);
or OR4 (N1118, N1112, N28, N496, N277);
buf BUF1 (N1119, N1114);
not NOT1 (N1120, N1119);
nand NAND4 (N1121, N1108, N306, N413, N614);
nor NOR2 (N1122, N1116, N67);
nand NAND4 (N1123, N1122, N755, N346, N949);
nor NOR2 (N1124, N1109, N1067);
buf BUF1 (N1125, N1105);
nand NAND3 (N1126, N1125, N363, N103);
not NOT1 (N1127, N1120);
and AND3 (N1128, N1118, N528, N220);
and AND3 (N1129, N1121, N96, N918);
nand NAND4 (N1130, N1127, N278, N290, N60);
nor NOR4 (N1131, N1111, N337, N542, N56);
buf BUF1 (N1132, N1124);
buf BUF1 (N1133, N1130);
xor XOR2 (N1134, N1115, N170);
not NOT1 (N1135, N1134);
buf BUF1 (N1136, N1104);
nor NOR3 (N1137, N1129, N257, N74);
nor NOR3 (N1138, N1131, N635, N53);
buf BUF1 (N1139, N1132);
or OR3 (N1140, N1136, N13, N506);
or OR2 (N1141, N1140, N88);
xor XOR2 (N1142, N1141, N480);
nand NAND2 (N1143, N1139, N638);
buf BUF1 (N1144, N1138);
and AND3 (N1145, N1137, N417, N221);
xor XOR2 (N1146, N1135, N294);
nor NOR2 (N1147, N1126, N44);
and AND4 (N1148, N1143, N1075, N646, N710);
xor XOR2 (N1149, N1142, N415);
and AND2 (N1150, N1133, N370);
not NOT1 (N1151, N1148);
xor XOR2 (N1152, N1150, N128);
xor XOR2 (N1153, N1145, N278);
nor NOR4 (N1154, N1151, N806, N1066, N890);
nor NOR3 (N1155, N1152, N1142, N637);
not NOT1 (N1156, N1149);
buf BUF1 (N1157, N1154);
nor NOR2 (N1158, N1156, N886);
or OR3 (N1159, N1128, N429, N393);
nand NAND2 (N1160, N1158, N962);
buf BUF1 (N1161, N1159);
buf BUF1 (N1162, N1123);
nor NOR4 (N1163, N1153, N1028, N1076, N152);
nand NAND2 (N1164, N1144, N279);
not NOT1 (N1165, N1146);
and AND3 (N1166, N1160, N1055, N654);
not NOT1 (N1167, N1165);
buf BUF1 (N1168, N1166);
not NOT1 (N1169, N1162);
or OR4 (N1170, N1169, N160, N998, N708);
xor XOR2 (N1171, N1163, N370);
nand NAND2 (N1172, N1155, N1105);
not NOT1 (N1173, N1164);
nor NOR2 (N1174, N1117, N21);
xor XOR2 (N1175, N1168, N10);
buf BUF1 (N1176, N1175);
xor XOR2 (N1177, N1170, N573);
not NOT1 (N1178, N1172);
and AND2 (N1179, N1177, N877);
buf BUF1 (N1180, N1157);
buf BUF1 (N1181, N1180);
nor NOR4 (N1182, N1179, N425, N403, N81);
nand NAND3 (N1183, N1178, N701, N853);
xor XOR2 (N1184, N1171, N469);
not NOT1 (N1185, N1173);
buf BUF1 (N1186, N1181);
nand NAND2 (N1187, N1182, N541);
not NOT1 (N1188, N1147);
nand NAND4 (N1189, N1176, N351, N50, N158);
not NOT1 (N1190, N1183);
xor XOR2 (N1191, N1188, N1106);
nor NOR3 (N1192, N1189, N1044, N400);
and AND2 (N1193, N1161, N828);
buf BUF1 (N1194, N1192);
or OR2 (N1195, N1190, N14);
nor NOR4 (N1196, N1174, N1040, N697, N223);
xor XOR2 (N1197, N1191, N120);
nor NOR3 (N1198, N1187, N269, N1019);
nor NOR2 (N1199, N1184, N766);
not NOT1 (N1200, N1199);
and AND3 (N1201, N1198, N307, N974);
nand NAND3 (N1202, N1201, N200, N408);
xor XOR2 (N1203, N1196, N263);
buf BUF1 (N1204, N1202);
nand NAND4 (N1205, N1203, N742, N646, N1191);
nand NAND2 (N1206, N1204, N221);
and AND4 (N1207, N1185, N1016, N620, N1095);
xor XOR2 (N1208, N1207, N197);
or OR2 (N1209, N1208, N548);
xor XOR2 (N1210, N1200, N141);
xor XOR2 (N1211, N1195, N1100);
xor XOR2 (N1212, N1186, N354);
nor NOR4 (N1213, N1212, N671, N924, N568);
nor NOR4 (N1214, N1211, N662, N840, N781);
not NOT1 (N1215, N1214);
xor XOR2 (N1216, N1215, N812);
and AND4 (N1217, N1213, N140, N532, N149);
and AND2 (N1218, N1206, N174);
not NOT1 (N1219, N1218);
nor NOR3 (N1220, N1210, N736, N192);
and AND3 (N1221, N1205, N908, N674);
and AND2 (N1222, N1216, N548);
and AND3 (N1223, N1167, N606, N633);
and AND3 (N1224, N1219, N1060, N332);
buf BUF1 (N1225, N1194);
and AND2 (N1226, N1224, N605);
xor XOR2 (N1227, N1221, N1094);
xor XOR2 (N1228, N1220, N974);
buf BUF1 (N1229, N1227);
nor NOR3 (N1230, N1193, N454, N487);
xor XOR2 (N1231, N1229, N25);
nand NAND2 (N1232, N1223, N62);
xor XOR2 (N1233, N1222, N1073);
not NOT1 (N1234, N1226);
nand NAND4 (N1235, N1234, N671, N1197, N962);
nor NOR2 (N1236, N295, N845);
and AND3 (N1237, N1235, N645, N1229);
and AND4 (N1238, N1233, N1211, N289, N409);
not NOT1 (N1239, N1225);
buf BUF1 (N1240, N1236);
and AND4 (N1241, N1237, N1066, N266, N896);
or OR4 (N1242, N1238, N378, N1200, N1104);
or OR3 (N1243, N1209, N852, N267);
not NOT1 (N1244, N1217);
nor NOR3 (N1245, N1231, N395, N647);
xor XOR2 (N1246, N1228, N513);
not NOT1 (N1247, N1232);
and AND4 (N1248, N1247, N1205, N963, N729);
xor XOR2 (N1249, N1241, N1074);
and AND4 (N1250, N1245, N930, N154, N194);
not NOT1 (N1251, N1250);
xor XOR2 (N1252, N1248, N365);
nor NOR3 (N1253, N1252, N5, N410);
and AND3 (N1254, N1251, N557, N1147);
nand NAND4 (N1255, N1239, N1071, N164, N818);
or OR4 (N1256, N1230, N1158, N856, N1139);
nor NOR4 (N1257, N1242, N115, N389, N311);
xor XOR2 (N1258, N1246, N139);
and AND4 (N1259, N1240, N1038, N918, N159);
xor XOR2 (N1260, N1244, N47);
buf BUF1 (N1261, N1258);
xor XOR2 (N1262, N1243, N1049);
and AND3 (N1263, N1257, N113, N481);
xor XOR2 (N1264, N1263, N682);
not NOT1 (N1265, N1256);
not NOT1 (N1266, N1265);
xor XOR2 (N1267, N1259, N1224);
xor XOR2 (N1268, N1260, N209);
nor NOR3 (N1269, N1253, N128, N223);
xor XOR2 (N1270, N1267, N589);
nor NOR3 (N1271, N1264, N758, N120);
not NOT1 (N1272, N1271);
nand NAND4 (N1273, N1270, N97, N611, N1148);
xor XOR2 (N1274, N1262, N543);
or OR2 (N1275, N1274, N565);
xor XOR2 (N1276, N1266, N142);
xor XOR2 (N1277, N1275, N7);
nand NAND4 (N1278, N1255, N19, N765, N623);
or OR2 (N1279, N1272, N777);
and AND4 (N1280, N1273, N259, N967, N627);
xor XOR2 (N1281, N1277, N1035);
buf BUF1 (N1282, N1278);
and AND4 (N1283, N1280, N53, N207, N1105);
xor XOR2 (N1284, N1269, N422);
nand NAND3 (N1285, N1284, N920, N268);
xor XOR2 (N1286, N1249, N1217);
or OR4 (N1287, N1283, N190, N1270, N42);
and AND3 (N1288, N1286, N694, N612);
buf BUF1 (N1289, N1261);
or OR3 (N1290, N1282, N673, N51);
and AND3 (N1291, N1268, N329, N733);
nand NAND4 (N1292, N1281, N779, N956, N1216);
or OR3 (N1293, N1285, N933, N498);
or OR4 (N1294, N1287, N1052, N65, N989);
xor XOR2 (N1295, N1289, N74);
nor NOR4 (N1296, N1292, N753, N99, N32);
and AND3 (N1297, N1288, N20, N1290);
nand NAND4 (N1298, N114, N263, N865, N667);
nor NOR4 (N1299, N1298, N196, N32, N1017);
xor XOR2 (N1300, N1294, N621);
and AND3 (N1301, N1291, N590, N1133);
not NOT1 (N1302, N1254);
buf BUF1 (N1303, N1301);
not NOT1 (N1304, N1297);
nand NAND2 (N1305, N1276, N1217);
buf BUF1 (N1306, N1296);
not NOT1 (N1307, N1295);
not NOT1 (N1308, N1305);
xor XOR2 (N1309, N1302, N1010);
buf BUF1 (N1310, N1293);
nor NOR3 (N1311, N1299, N265, N182);
nand NAND2 (N1312, N1304, N255);
or OR4 (N1313, N1309, N1153, N327, N137);
and AND4 (N1314, N1307, N224, N233, N228);
nand NAND2 (N1315, N1310, N708);
and AND3 (N1316, N1311, N451, N22);
buf BUF1 (N1317, N1312);
nor NOR3 (N1318, N1316, N1013, N678);
nand NAND4 (N1319, N1318, N726, N683, N124);
nand NAND2 (N1320, N1300, N1205);
nor NOR4 (N1321, N1320, N175, N536, N207);
nand NAND2 (N1322, N1321, N1072);
not NOT1 (N1323, N1319);
and AND4 (N1324, N1306, N12, N491, N908);
nor NOR3 (N1325, N1317, N491, N193);
xor XOR2 (N1326, N1323, N232);
xor XOR2 (N1327, N1326, N699);
xor XOR2 (N1328, N1308, N776);
nor NOR2 (N1329, N1303, N640);
and AND3 (N1330, N1279, N878, N1033);
nor NOR2 (N1331, N1329, N1068);
nor NOR3 (N1332, N1314, N427, N666);
and AND4 (N1333, N1327, N539, N1026, N876);
buf BUF1 (N1334, N1330);
nor NOR3 (N1335, N1325, N402, N1089);
and AND2 (N1336, N1328, N431);
buf BUF1 (N1337, N1334);
xor XOR2 (N1338, N1333, N614);
nor NOR2 (N1339, N1332, N1013);
buf BUF1 (N1340, N1336);
and AND3 (N1341, N1322, N1039, N417);
buf BUF1 (N1342, N1331);
xor XOR2 (N1343, N1342, N430);
nor NOR4 (N1344, N1341, N1094, N571, N204);
buf BUF1 (N1345, N1343);
buf BUF1 (N1346, N1339);
xor XOR2 (N1347, N1313, N1322);
xor XOR2 (N1348, N1347, N1260);
xor XOR2 (N1349, N1340, N778);
and AND3 (N1350, N1337, N744, N1023);
buf BUF1 (N1351, N1315);
nor NOR2 (N1352, N1338, N845);
nor NOR3 (N1353, N1324, N824, N268);
xor XOR2 (N1354, N1352, N508);
xor XOR2 (N1355, N1354, N311);
or OR2 (N1356, N1350, N156);
or OR2 (N1357, N1355, N1316);
nor NOR2 (N1358, N1348, N329);
not NOT1 (N1359, N1351);
nor NOR2 (N1360, N1356, N72);
or OR4 (N1361, N1344, N75, N19, N673);
nor NOR2 (N1362, N1346, N47);
not NOT1 (N1363, N1361);
nand NAND4 (N1364, N1349, N914, N835, N468);
or OR2 (N1365, N1357, N1237);
not NOT1 (N1366, N1363);
nand NAND2 (N1367, N1360, N1013);
not NOT1 (N1368, N1367);
not NOT1 (N1369, N1364);
xor XOR2 (N1370, N1365, N14);
xor XOR2 (N1371, N1359, N289);
xor XOR2 (N1372, N1366, N1125);
nor NOR2 (N1373, N1369, N609);
or OR2 (N1374, N1373, N483);
and AND2 (N1375, N1372, N171);
or OR3 (N1376, N1371, N342, N630);
not NOT1 (N1377, N1353);
nor NOR4 (N1378, N1335, N152, N1125, N43);
nor NOR2 (N1379, N1378, N860);
nand NAND3 (N1380, N1362, N1070, N1166);
buf BUF1 (N1381, N1377);
xor XOR2 (N1382, N1368, N1047);
or OR3 (N1383, N1379, N567, N1086);
nand NAND4 (N1384, N1345, N1256, N659, N171);
and AND3 (N1385, N1384, N873, N343);
nor NOR3 (N1386, N1381, N836, N885);
or OR4 (N1387, N1382, N1160, N538, N763);
nand NAND4 (N1388, N1380, N85, N369, N57);
xor XOR2 (N1389, N1386, N466);
buf BUF1 (N1390, N1376);
not NOT1 (N1391, N1383);
nor NOR3 (N1392, N1385, N840, N1158);
buf BUF1 (N1393, N1375);
or OR4 (N1394, N1358, N663, N630, N617);
not NOT1 (N1395, N1389);
not NOT1 (N1396, N1394);
or OR4 (N1397, N1374, N443, N986, N427);
buf BUF1 (N1398, N1388);
buf BUF1 (N1399, N1370);
or OR4 (N1400, N1387, N53, N950, N1247);
or OR2 (N1401, N1392, N727);
nor NOR2 (N1402, N1400, N1180);
buf BUF1 (N1403, N1401);
or OR3 (N1404, N1402, N894, N318);
nand NAND3 (N1405, N1390, N588, N1088);
and AND4 (N1406, N1397, N449, N1353, N1076);
xor XOR2 (N1407, N1398, N877);
or OR4 (N1408, N1404, N681, N946, N147);
not NOT1 (N1409, N1405);
buf BUF1 (N1410, N1393);
nor NOR3 (N1411, N1410, N67, N826);
buf BUF1 (N1412, N1409);
nand NAND3 (N1413, N1403, N719, N793);
or OR4 (N1414, N1413, N1206, N18, N372);
not NOT1 (N1415, N1407);
and AND3 (N1416, N1395, N585, N1381);
nand NAND4 (N1417, N1411, N245, N749, N296);
xor XOR2 (N1418, N1415, N1141);
and AND4 (N1419, N1408, N897, N451, N133);
buf BUF1 (N1420, N1419);
nor NOR2 (N1421, N1396, N430);
and AND2 (N1422, N1420, N779);
and AND3 (N1423, N1414, N899, N1066);
buf BUF1 (N1424, N1422);
nor NOR2 (N1425, N1421, N65);
and AND4 (N1426, N1418, N510, N1152, N1085);
and AND3 (N1427, N1412, N803, N1036);
and AND3 (N1428, N1416, N827, N315);
and AND2 (N1429, N1399, N9);
not NOT1 (N1430, N1429);
nand NAND2 (N1431, N1423, N1100);
and AND4 (N1432, N1417, N376, N943, N19);
and AND3 (N1433, N1391, N938, N1361);
nor NOR2 (N1434, N1433, N154);
xor XOR2 (N1435, N1430, N55);
nand NAND2 (N1436, N1431, N1009);
nand NAND3 (N1437, N1434, N211, N23);
nor NOR4 (N1438, N1436, N33, N618, N655);
nor NOR2 (N1439, N1406, N189);
nand NAND3 (N1440, N1435, N475, N1260);
and AND4 (N1441, N1432, N1124, N1006, N786);
xor XOR2 (N1442, N1439, N1117);
buf BUF1 (N1443, N1437);
xor XOR2 (N1444, N1438, N541);
nand NAND2 (N1445, N1440, N371);
and AND2 (N1446, N1424, N1117);
not NOT1 (N1447, N1426);
or OR4 (N1448, N1447, N6, N497, N805);
buf BUF1 (N1449, N1446);
nor NOR2 (N1450, N1442, N1261);
nor NOR4 (N1451, N1428, N507, N275, N1285);
and AND4 (N1452, N1448, N279, N349, N18);
xor XOR2 (N1453, N1445, N351);
not NOT1 (N1454, N1443);
or OR4 (N1455, N1454, N192, N881, N706);
not NOT1 (N1456, N1455);
not NOT1 (N1457, N1456);
xor XOR2 (N1458, N1453, N493);
nor NOR2 (N1459, N1427, N349);
nand NAND4 (N1460, N1451, N1100, N326, N955);
or OR2 (N1461, N1460, N462);
nand NAND4 (N1462, N1425, N482, N1299, N234);
or OR2 (N1463, N1449, N1327);
or OR4 (N1464, N1452, N1081, N883, N482);
xor XOR2 (N1465, N1459, N1081);
nor NOR2 (N1466, N1461, N535);
xor XOR2 (N1467, N1462, N1397);
nand NAND2 (N1468, N1457, N496);
buf BUF1 (N1469, N1466);
nor NOR2 (N1470, N1465, N1003);
not NOT1 (N1471, N1463);
or OR4 (N1472, N1468, N549, N95, N996);
not NOT1 (N1473, N1444);
buf BUF1 (N1474, N1473);
nor NOR4 (N1475, N1472, N1318, N703, N490);
buf BUF1 (N1476, N1471);
nor NOR4 (N1477, N1464, N705, N1056, N204);
buf BUF1 (N1478, N1450);
nor NOR2 (N1479, N1458, N317);
nand NAND3 (N1480, N1467, N1290, N490);
and AND3 (N1481, N1478, N250, N269);
or OR4 (N1482, N1469, N697, N583, N558);
nand NAND4 (N1483, N1474, N402, N1105, N603);
nand NAND2 (N1484, N1480, N965);
and AND2 (N1485, N1470, N612);
and AND4 (N1486, N1479, N1318, N297, N1095);
buf BUF1 (N1487, N1482);
not NOT1 (N1488, N1485);
xor XOR2 (N1489, N1486, N1342);
and AND3 (N1490, N1475, N1222, N556);
buf BUF1 (N1491, N1476);
or OR2 (N1492, N1477, N1190);
and AND3 (N1493, N1488, N38, N87);
nor NOR4 (N1494, N1487, N343, N1072, N81);
not NOT1 (N1495, N1491);
and AND3 (N1496, N1495, N200, N310);
xor XOR2 (N1497, N1496, N952);
or OR2 (N1498, N1493, N1461);
nand NAND2 (N1499, N1497, N34);
nand NAND3 (N1500, N1483, N1058, N193);
nand NAND3 (N1501, N1499, N538, N301);
or OR2 (N1502, N1489, N274);
nor NOR3 (N1503, N1500, N253, N596);
nor NOR4 (N1504, N1498, N581, N1129, N688);
buf BUF1 (N1505, N1502);
xor XOR2 (N1506, N1505, N980);
xor XOR2 (N1507, N1492, N637);
not NOT1 (N1508, N1481);
xor XOR2 (N1509, N1494, N1061);
xor XOR2 (N1510, N1504, N967);
nor NOR4 (N1511, N1506, N127, N498, N352);
or OR3 (N1512, N1503, N1074, N305);
and AND4 (N1513, N1509, N79, N1186, N1304);
not NOT1 (N1514, N1510);
and AND4 (N1515, N1501, N414, N1253, N1092);
not NOT1 (N1516, N1514);
not NOT1 (N1517, N1508);
not NOT1 (N1518, N1512);
and AND2 (N1519, N1518, N698);
or OR4 (N1520, N1513, N218, N645, N1426);
xor XOR2 (N1521, N1519, N1375);
nand NAND2 (N1522, N1520, N435);
nand NAND2 (N1523, N1507, N449);
nand NAND3 (N1524, N1517, N947, N926);
not NOT1 (N1525, N1515);
or OR2 (N1526, N1522, N392);
not NOT1 (N1527, N1511);
not NOT1 (N1528, N1526);
buf BUF1 (N1529, N1525);
or OR3 (N1530, N1484, N26, N1464);
or OR4 (N1531, N1530, N417, N660, N1057);
xor XOR2 (N1532, N1521, N330);
xor XOR2 (N1533, N1516, N503);
buf BUF1 (N1534, N1527);
not NOT1 (N1535, N1534);
or OR2 (N1536, N1490, N274);
not NOT1 (N1537, N1532);
or OR4 (N1538, N1523, N759, N822, N1128);
buf BUF1 (N1539, N1528);
not NOT1 (N1540, N1536);
or OR4 (N1541, N1535, N921, N838, N1390);
buf BUF1 (N1542, N1529);
xor XOR2 (N1543, N1540, N904);
xor XOR2 (N1544, N1524, N723);
or OR4 (N1545, N1531, N358, N873, N699);
and AND2 (N1546, N1537, N732);
nor NOR3 (N1547, N1533, N791, N248);
xor XOR2 (N1548, N1547, N1443);
xor XOR2 (N1549, N1548, N1539);
nor NOR4 (N1550, N805, N1250, N788, N1252);
nand NAND4 (N1551, N1546, N7, N1326, N758);
xor XOR2 (N1552, N1543, N434);
nor NOR2 (N1553, N1551, N1180);
or OR3 (N1554, N1541, N476, N1315);
xor XOR2 (N1555, N1538, N1125);
and AND2 (N1556, N1545, N1552);
or OR2 (N1557, N778, N1136);
and AND4 (N1558, N1556, N1322, N820, N417);
buf BUF1 (N1559, N1549);
not NOT1 (N1560, N1555);
buf BUF1 (N1561, N1544);
buf BUF1 (N1562, N1542);
xor XOR2 (N1563, N1557, N1160);
nand NAND4 (N1564, N1550, N1440, N286, N1213);
buf BUF1 (N1565, N1564);
not NOT1 (N1566, N1559);
nand NAND2 (N1567, N1553, N496);
and AND2 (N1568, N1566, N886);
nor NOR3 (N1569, N1563, N347, N736);
buf BUF1 (N1570, N1569);
buf BUF1 (N1571, N1560);
nor NOR4 (N1572, N1568, N453, N708, N658);
nor NOR4 (N1573, N1441, N1300, N828, N467);
nor NOR4 (N1574, N1572, N340, N144, N769);
not NOT1 (N1575, N1574);
nand NAND3 (N1576, N1562, N1306, N1556);
or OR3 (N1577, N1565, N1246, N442);
nand NAND2 (N1578, N1570, N320);
nand NAND3 (N1579, N1573, N813, N1400);
nand NAND2 (N1580, N1554, N282);
not NOT1 (N1581, N1579);
and AND3 (N1582, N1577, N718, N989);
and AND2 (N1583, N1558, N466);
nand NAND3 (N1584, N1567, N65, N1256);
and AND3 (N1585, N1571, N765, N1227);
or OR3 (N1586, N1561, N134, N83);
or OR3 (N1587, N1581, N36, N891);
nor NOR4 (N1588, N1587, N1174, N843, N1572);
xor XOR2 (N1589, N1576, N622);
not NOT1 (N1590, N1589);
nand NAND2 (N1591, N1584, N378);
nor NOR4 (N1592, N1583, N1545, N509, N756);
buf BUF1 (N1593, N1591);
nand NAND4 (N1594, N1586, N1202, N296, N884);
buf BUF1 (N1595, N1585);
and AND2 (N1596, N1578, N346);
or OR3 (N1597, N1592, N1096, N1215);
nand NAND2 (N1598, N1596, N1073);
not NOT1 (N1599, N1597);
nand NAND3 (N1600, N1582, N1064, N1365);
nand NAND4 (N1601, N1588, N230, N25, N12);
nor NOR4 (N1602, N1599, N1467, N147, N70);
buf BUF1 (N1603, N1598);
buf BUF1 (N1604, N1600);
nand NAND4 (N1605, N1602, N731, N478, N905);
nor NOR4 (N1606, N1604, N595, N1441, N767);
and AND4 (N1607, N1605, N651, N1253, N986);
nand NAND3 (N1608, N1575, N646, N1516);
nand NAND2 (N1609, N1593, N1103);
not NOT1 (N1610, N1607);
buf BUF1 (N1611, N1595);
buf BUF1 (N1612, N1601);
xor XOR2 (N1613, N1590, N1463);
not NOT1 (N1614, N1594);
xor XOR2 (N1615, N1611, N1508);
nor NOR3 (N1616, N1612, N1501, N1110);
not NOT1 (N1617, N1608);
xor XOR2 (N1618, N1617, N453);
nor NOR3 (N1619, N1613, N274, N867);
not NOT1 (N1620, N1606);
nor NOR2 (N1621, N1616, N1130);
nor NOR4 (N1622, N1609, N936, N922, N572);
and AND4 (N1623, N1603, N1566, N1105, N148);
xor XOR2 (N1624, N1618, N403);
nor NOR4 (N1625, N1620, N173, N1057, N1448);
buf BUF1 (N1626, N1624);
xor XOR2 (N1627, N1614, N264);
buf BUF1 (N1628, N1619);
or OR4 (N1629, N1628, N1557, N1035, N1081);
buf BUF1 (N1630, N1610);
nor NOR3 (N1631, N1625, N1222, N1283);
and AND3 (N1632, N1630, N1425, N1566);
and AND3 (N1633, N1629, N1534, N1354);
not NOT1 (N1634, N1580);
and AND3 (N1635, N1632, N606, N445);
buf BUF1 (N1636, N1635);
xor XOR2 (N1637, N1631, N1444);
or OR4 (N1638, N1622, N1032, N1134, N224);
and AND3 (N1639, N1638, N358, N1565);
nor NOR2 (N1640, N1637, N1301);
or OR3 (N1641, N1626, N336, N798);
nor NOR4 (N1642, N1634, N794, N344, N1409);
buf BUF1 (N1643, N1627);
and AND2 (N1644, N1636, N304);
or OR4 (N1645, N1644, N268, N1093, N134);
nor NOR2 (N1646, N1640, N356);
buf BUF1 (N1647, N1642);
or OR4 (N1648, N1641, N308, N177, N222);
and AND4 (N1649, N1648, N1279, N757, N766);
buf BUF1 (N1650, N1615);
not NOT1 (N1651, N1645);
or OR2 (N1652, N1651, N133);
buf BUF1 (N1653, N1647);
not NOT1 (N1654, N1653);
and AND4 (N1655, N1646, N1117, N411, N731);
nand NAND2 (N1656, N1650, N360);
nor NOR2 (N1657, N1652, N30);
and AND4 (N1658, N1639, N500, N547, N820);
buf BUF1 (N1659, N1643);
nor NOR4 (N1660, N1623, N1137, N725, N720);
and AND3 (N1661, N1621, N795, N759);
xor XOR2 (N1662, N1633, N487);
not NOT1 (N1663, N1660);
not NOT1 (N1664, N1659);
buf BUF1 (N1665, N1663);
buf BUF1 (N1666, N1654);
and AND2 (N1667, N1665, N1479);
or OR3 (N1668, N1658, N939, N499);
nor NOR4 (N1669, N1656, N1227, N1450, N237);
xor XOR2 (N1670, N1657, N116);
buf BUF1 (N1671, N1664);
or OR4 (N1672, N1669, N1518, N335, N1581);
not NOT1 (N1673, N1671);
and AND2 (N1674, N1667, N203);
or OR4 (N1675, N1666, N1116, N1305, N1336);
xor XOR2 (N1676, N1655, N1575);
or OR4 (N1677, N1675, N119, N1395, N994);
xor XOR2 (N1678, N1674, N1018);
xor XOR2 (N1679, N1676, N1019);
and AND3 (N1680, N1678, N1204, N1637);
and AND3 (N1681, N1672, N984, N744);
not NOT1 (N1682, N1681);
buf BUF1 (N1683, N1680);
buf BUF1 (N1684, N1670);
buf BUF1 (N1685, N1649);
and AND2 (N1686, N1661, N1293);
xor XOR2 (N1687, N1679, N690);
buf BUF1 (N1688, N1683);
or OR4 (N1689, N1662, N450, N1468, N670);
nand NAND3 (N1690, N1673, N1163, N246);
or OR2 (N1691, N1690, N757);
nand NAND3 (N1692, N1686, N733, N128);
and AND4 (N1693, N1682, N1598, N182, N605);
nor NOR2 (N1694, N1688, N592);
buf BUF1 (N1695, N1692);
nand NAND3 (N1696, N1687, N729, N979);
and AND4 (N1697, N1695, N322, N956, N530);
buf BUF1 (N1698, N1693);
not NOT1 (N1699, N1691);
or OR3 (N1700, N1668, N1085, N1459);
nand NAND4 (N1701, N1697, N876, N335, N351);
xor XOR2 (N1702, N1701, N1486);
xor XOR2 (N1703, N1700, N1676);
buf BUF1 (N1704, N1677);
not NOT1 (N1705, N1703);
nand NAND2 (N1706, N1699, N468);
or OR4 (N1707, N1705, N587, N1676, N695);
or OR3 (N1708, N1698, N269, N358);
xor XOR2 (N1709, N1689, N735);
and AND3 (N1710, N1704, N410, N1108);
not NOT1 (N1711, N1685);
xor XOR2 (N1712, N1709, N1325);
and AND4 (N1713, N1696, N1180, N860, N521);
or OR4 (N1714, N1694, N856, N834, N704);
nand NAND2 (N1715, N1711, N833);
nor NOR3 (N1716, N1706, N447, N974);
or OR3 (N1717, N1713, N427, N375);
xor XOR2 (N1718, N1716, N733);
nor NOR2 (N1719, N1718, N928);
nor NOR2 (N1720, N1714, N840);
nor NOR4 (N1721, N1707, N1295, N1638, N467);
nor NOR4 (N1722, N1712, N93, N1494, N589);
nor NOR2 (N1723, N1710, N1211);
nand NAND3 (N1724, N1715, N758, N350);
not NOT1 (N1725, N1721);
nand NAND3 (N1726, N1717, N180, N1556);
or OR2 (N1727, N1725, N404);
buf BUF1 (N1728, N1720);
buf BUF1 (N1729, N1728);
not NOT1 (N1730, N1708);
nand NAND3 (N1731, N1702, N1392, N679);
and AND4 (N1732, N1684, N677, N1048, N522);
or OR3 (N1733, N1727, N164, N1597);
and AND3 (N1734, N1724, N246, N1589);
nor NOR4 (N1735, N1733, N1149, N1681, N1135);
or OR3 (N1736, N1719, N362, N1216);
nor NOR2 (N1737, N1730, N1555);
and AND2 (N1738, N1729, N773);
or OR4 (N1739, N1723, N1602, N1465, N1703);
or OR3 (N1740, N1739, N1543, N9);
nand NAND4 (N1741, N1740, N787, N793, N264);
and AND4 (N1742, N1736, N1326, N1427, N1025);
or OR2 (N1743, N1738, N1381);
not NOT1 (N1744, N1741);
nand NAND4 (N1745, N1732, N224, N1535, N1259);
nand NAND2 (N1746, N1734, N1029);
nand NAND2 (N1747, N1722, N1126);
nand NAND4 (N1748, N1743, N1277, N1551, N1410);
nand NAND4 (N1749, N1726, N1495, N496, N1093);
buf BUF1 (N1750, N1745);
nor NOR4 (N1751, N1737, N1652, N1563, N975);
not NOT1 (N1752, N1731);
xor XOR2 (N1753, N1750, N364);
xor XOR2 (N1754, N1753, N684);
xor XOR2 (N1755, N1748, N420);
or OR4 (N1756, N1755, N540, N286, N711);
nand NAND3 (N1757, N1746, N248, N1182);
or OR4 (N1758, N1752, N737, N772, N991);
and AND2 (N1759, N1758, N1107);
buf BUF1 (N1760, N1757);
and AND3 (N1761, N1754, N883, N890);
and AND3 (N1762, N1751, N277, N297);
not NOT1 (N1763, N1735);
nor NOR4 (N1764, N1742, N750, N268, N1412);
not NOT1 (N1765, N1760);
and AND2 (N1766, N1744, N1423);
not NOT1 (N1767, N1761);
not NOT1 (N1768, N1765);
buf BUF1 (N1769, N1764);
or OR3 (N1770, N1769, N296, N1386);
buf BUF1 (N1771, N1768);
or OR3 (N1772, N1756, N1253, N191);
nor NOR2 (N1773, N1759, N624);
or OR2 (N1774, N1771, N1117);
and AND3 (N1775, N1762, N544, N185);
nand NAND3 (N1776, N1774, N1596, N489);
xor XOR2 (N1777, N1749, N280);
and AND2 (N1778, N1747, N418);
and AND3 (N1779, N1767, N1194, N1399);
nand NAND2 (N1780, N1775, N150);
xor XOR2 (N1781, N1766, N1425);
not NOT1 (N1782, N1763);
xor XOR2 (N1783, N1770, N170);
or OR3 (N1784, N1782, N29, N1703);
not NOT1 (N1785, N1772);
nand NAND3 (N1786, N1779, N284, N1558);
buf BUF1 (N1787, N1783);
not NOT1 (N1788, N1776);
or OR3 (N1789, N1785, N476, N991);
or OR3 (N1790, N1773, N494, N441);
nor NOR4 (N1791, N1786, N24, N1725, N863);
and AND4 (N1792, N1778, N912, N679, N458);
xor XOR2 (N1793, N1790, N394);
nand NAND3 (N1794, N1791, N721, N386);
buf BUF1 (N1795, N1789);
and AND2 (N1796, N1792, N1722);
nand NAND4 (N1797, N1780, N166, N1391, N1072);
nor NOR3 (N1798, N1795, N431, N5);
xor XOR2 (N1799, N1777, N1177);
buf BUF1 (N1800, N1784);
xor XOR2 (N1801, N1788, N209);
buf BUF1 (N1802, N1794);
not NOT1 (N1803, N1797);
and AND4 (N1804, N1801, N1602, N154, N449);
and AND3 (N1805, N1781, N351, N30);
and AND4 (N1806, N1803, N334, N383, N622);
nor NOR2 (N1807, N1798, N1022);
buf BUF1 (N1808, N1807);
and AND3 (N1809, N1805, N1605, N1756);
xor XOR2 (N1810, N1796, N757);
buf BUF1 (N1811, N1799);
nor NOR2 (N1812, N1810, N1104);
not NOT1 (N1813, N1787);
xor XOR2 (N1814, N1808, N943);
not NOT1 (N1815, N1804);
buf BUF1 (N1816, N1811);
buf BUF1 (N1817, N1814);
nand NAND2 (N1818, N1802, N1248);
buf BUF1 (N1819, N1809);
xor XOR2 (N1820, N1800, N1456);
or OR4 (N1821, N1818, N62, N1570, N1000);
nand NAND4 (N1822, N1819, N523, N1733, N955);
not NOT1 (N1823, N1793);
buf BUF1 (N1824, N1822);
xor XOR2 (N1825, N1820, N1280);
nor NOR2 (N1826, N1812, N1121);
xor XOR2 (N1827, N1817, N323);
nor NOR4 (N1828, N1827, N1294, N1552, N490);
xor XOR2 (N1829, N1828, N1455);
xor XOR2 (N1830, N1821, N970);
xor XOR2 (N1831, N1823, N977);
xor XOR2 (N1832, N1829, N17);
buf BUF1 (N1833, N1816);
not NOT1 (N1834, N1832);
nand NAND3 (N1835, N1826, N1196, N238);
nor NOR3 (N1836, N1825, N1631, N250);
nand NAND3 (N1837, N1815, N252, N1105);
not NOT1 (N1838, N1824);
and AND3 (N1839, N1834, N1719, N863);
or OR4 (N1840, N1837, N811, N1363, N388);
not NOT1 (N1841, N1838);
buf BUF1 (N1842, N1840);
nand NAND2 (N1843, N1839, N1769);
not NOT1 (N1844, N1841);
nor NOR3 (N1845, N1813, N1428, N1575);
nor NOR3 (N1846, N1842, N1041, N1444);
and AND4 (N1847, N1844, N868, N376, N1189);
not NOT1 (N1848, N1843);
nand NAND4 (N1849, N1847, N1042, N711, N1197);
not NOT1 (N1850, N1831);
buf BUF1 (N1851, N1835);
xor XOR2 (N1852, N1806, N562);
nand NAND2 (N1853, N1845, N302);
xor XOR2 (N1854, N1836, N1232);
or OR4 (N1855, N1851, N653, N435, N1575);
buf BUF1 (N1856, N1854);
or OR3 (N1857, N1855, N1658, N1526);
nand NAND2 (N1858, N1853, N1025);
nand NAND4 (N1859, N1833, N1739, N519, N1112);
xor XOR2 (N1860, N1849, N490);
nand NAND3 (N1861, N1859, N1809, N1064);
not NOT1 (N1862, N1852);
buf BUF1 (N1863, N1862);
nand NAND3 (N1864, N1850, N1646, N69);
xor XOR2 (N1865, N1846, N482);
xor XOR2 (N1866, N1860, N865);
buf BUF1 (N1867, N1866);
nor NOR3 (N1868, N1830, N455, N654);
not NOT1 (N1869, N1858);
or OR4 (N1870, N1863, N1111, N399, N263);
nor NOR2 (N1871, N1870, N910);
xor XOR2 (N1872, N1856, N1162);
or OR2 (N1873, N1857, N303);
nor NOR3 (N1874, N1869, N1546, N1073);
or OR4 (N1875, N1865, N1215, N315, N1282);
not NOT1 (N1876, N1864);
buf BUF1 (N1877, N1873);
or OR4 (N1878, N1876, N1283, N1735, N1528);
xor XOR2 (N1879, N1861, N363);
or OR4 (N1880, N1879, N287, N1291, N1566);
buf BUF1 (N1881, N1872);
or OR2 (N1882, N1880, N1153);
nand NAND3 (N1883, N1848, N216, N720);
not NOT1 (N1884, N1874);
nor NOR2 (N1885, N1883, N1762);
nor NOR4 (N1886, N1877, N1556, N1266, N844);
not NOT1 (N1887, N1871);
not NOT1 (N1888, N1887);
nor NOR4 (N1889, N1884, N718, N1825, N887);
nand NAND3 (N1890, N1867, N1874, N136);
or OR4 (N1891, N1882, N478, N768, N751);
and AND2 (N1892, N1891, N511);
not NOT1 (N1893, N1890);
not NOT1 (N1894, N1868);
buf BUF1 (N1895, N1885);
buf BUF1 (N1896, N1875);
xor XOR2 (N1897, N1888, N728);
buf BUF1 (N1898, N1895);
buf BUF1 (N1899, N1881);
and AND4 (N1900, N1899, N83, N1207, N1120);
nand NAND2 (N1901, N1900, N531);
nand NAND2 (N1902, N1896, N906);
and AND3 (N1903, N1897, N1721, N1148);
and AND2 (N1904, N1886, N468);
or OR3 (N1905, N1893, N906, N384);
and AND3 (N1906, N1904, N26, N1573);
not NOT1 (N1907, N1894);
not NOT1 (N1908, N1889);
nor NOR4 (N1909, N1901, N203, N668, N1585);
buf BUF1 (N1910, N1892);
or OR3 (N1911, N1905, N352, N1229);
or OR4 (N1912, N1878, N1062, N856, N1264);
xor XOR2 (N1913, N1908, N1379);
xor XOR2 (N1914, N1909, N668);
xor XOR2 (N1915, N1914, N582);
nor NOR3 (N1916, N1903, N1733, N749);
xor XOR2 (N1917, N1912, N543);
buf BUF1 (N1918, N1915);
buf BUF1 (N1919, N1913);
buf BUF1 (N1920, N1911);
and AND4 (N1921, N1910, N1703, N1747, N593);
buf BUF1 (N1922, N1921);
buf BUF1 (N1923, N1919);
xor XOR2 (N1924, N1923, N1621);
not NOT1 (N1925, N1902);
or OR4 (N1926, N1922, N714, N1524, N1634);
nand NAND4 (N1927, N1898, N565, N1531, N1664);
nor NOR4 (N1928, N1925, N1924, N404, N1873);
nor NOR2 (N1929, N369, N1491);
nor NOR4 (N1930, N1916, N323, N505, N877);
buf BUF1 (N1931, N1907);
nand NAND2 (N1932, N1928, N1374);
and AND2 (N1933, N1918, N412);
and AND3 (N1934, N1906, N1201, N718);
and AND3 (N1935, N1932, N1541, N76);
nand NAND2 (N1936, N1930, N1456);
or OR4 (N1937, N1920, N897, N485, N20);
nand NAND2 (N1938, N1931, N1559);
nand NAND2 (N1939, N1935, N1345);
nand NAND4 (N1940, N1917, N9, N691, N1592);
and AND2 (N1941, N1934, N1026);
nand NAND3 (N1942, N1939, N1405, N375);
and AND4 (N1943, N1937, N1340, N1497, N98);
xor XOR2 (N1944, N1942, N1545);
not NOT1 (N1945, N1936);
or OR3 (N1946, N1938, N1237, N105);
or OR3 (N1947, N1926, N82, N238);
or OR2 (N1948, N1929, N1076);
nor NOR3 (N1949, N1927, N13, N920);
nor NOR3 (N1950, N1933, N1694, N1019);
xor XOR2 (N1951, N1943, N466);
or OR4 (N1952, N1944, N550, N39, N1558);
nor NOR2 (N1953, N1950, N273);
buf BUF1 (N1954, N1949);
buf BUF1 (N1955, N1952);
not NOT1 (N1956, N1945);
buf BUF1 (N1957, N1953);
nor NOR4 (N1958, N1947, N1023, N413, N1805);
not NOT1 (N1959, N1941);
xor XOR2 (N1960, N1958, N986);
not NOT1 (N1961, N1954);
not NOT1 (N1962, N1955);
or OR2 (N1963, N1959, N216);
xor XOR2 (N1964, N1956, N633);
or OR2 (N1965, N1948, N791);
nand NAND3 (N1966, N1962, N1879, N580);
nor NOR2 (N1967, N1963, N1138);
nor NOR4 (N1968, N1964, N740, N1926, N904);
nor NOR3 (N1969, N1965, N1726, N1685);
nor NOR3 (N1970, N1951, N1778, N1117);
xor XOR2 (N1971, N1960, N526);
and AND2 (N1972, N1946, N1323);
xor XOR2 (N1973, N1966, N391);
and AND2 (N1974, N1970, N361);
nor NOR4 (N1975, N1967, N699, N1089, N1210);
buf BUF1 (N1976, N1971);
or OR3 (N1977, N1957, N1580, N651);
buf BUF1 (N1978, N1972);
or OR2 (N1979, N1940, N1291);
buf BUF1 (N1980, N1968);
nor NOR2 (N1981, N1975, N688);
nand NAND2 (N1982, N1974, N404);
buf BUF1 (N1983, N1979);
buf BUF1 (N1984, N1976);
nand NAND4 (N1985, N1961, N677, N331, N1600);
nand NAND3 (N1986, N1980, N77, N89);
xor XOR2 (N1987, N1977, N631);
nand NAND4 (N1988, N1983, N1170, N412, N129);
nor NOR2 (N1989, N1987, N1772);
nor NOR2 (N1990, N1988, N1407);
nor NOR2 (N1991, N1985, N1442);
not NOT1 (N1992, N1981);
buf BUF1 (N1993, N1984);
buf BUF1 (N1994, N1969);
buf BUF1 (N1995, N1973);
nand NAND3 (N1996, N1993, N930, N552);
or OR3 (N1997, N1996, N1695, N1026);
or OR4 (N1998, N1982, N761, N1901, N1289);
nand NAND3 (N1999, N1986, N1019, N990);
not NOT1 (N2000, N1990);
or OR4 (N2001, N1992, N87, N1165, N1294);
nand NAND4 (N2002, N2000, N1540, N1534, N119);
or OR2 (N2003, N1989, N1411);
not NOT1 (N2004, N1978);
buf BUF1 (N2005, N1997);
xor XOR2 (N2006, N1995, N1611);
buf BUF1 (N2007, N2003);
buf BUF1 (N2008, N1998);
not NOT1 (N2009, N1999);
nand NAND4 (N2010, N2004, N234, N1946, N1469);
nand NAND4 (N2011, N2006, N199, N897, N1932);
nand NAND2 (N2012, N1994, N49);
nand NAND3 (N2013, N2001, N1418, N1422);
nand NAND3 (N2014, N2012, N477, N520);
xor XOR2 (N2015, N2013, N306);
or OR4 (N2016, N2009, N1403, N773, N1943);
xor XOR2 (N2017, N1991, N1240);
or OR3 (N2018, N2015, N299, N1459);
and AND2 (N2019, N2014, N805);
nand NAND4 (N2020, N2002, N552, N27, N1199);
or OR3 (N2021, N2016, N1085, N247);
not NOT1 (N2022, N2011);
buf BUF1 (N2023, N2005);
xor XOR2 (N2024, N2010, N1771);
nand NAND2 (N2025, N2019, N800);
and AND4 (N2026, N2024, N1328, N1565, N513);
not NOT1 (N2027, N2023);
and AND4 (N2028, N2008, N157, N446, N242);
and AND2 (N2029, N2022, N1288);
not NOT1 (N2030, N2007);
and AND2 (N2031, N2030, N56);
buf BUF1 (N2032, N2018);
and AND3 (N2033, N2026, N1482, N77);
or OR3 (N2034, N2033, N1116, N160);
nor NOR4 (N2035, N2034, N157, N1522, N407);
not NOT1 (N2036, N2021);
or OR4 (N2037, N2031, N729, N1184, N578);
not NOT1 (N2038, N2029);
nand NAND3 (N2039, N2027, N608, N15);
nor NOR2 (N2040, N2037, N1354);
and AND2 (N2041, N2038, N189);
not NOT1 (N2042, N2028);
nand NAND4 (N2043, N2039, N1464, N1835, N1447);
nand NAND3 (N2044, N2042, N1249, N6);
or OR3 (N2045, N2041, N554, N1043);
buf BUF1 (N2046, N2045);
nand NAND4 (N2047, N2043, N556, N1574, N232);
nor NOR3 (N2048, N2046, N656, N677);
buf BUF1 (N2049, N2036);
nor NOR3 (N2050, N2044, N586, N384);
nand NAND2 (N2051, N2020, N253);
nor NOR4 (N2052, N2035, N471, N1485, N794);
or OR3 (N2053, N2051, N1705, N1396);
and AND4 (N2054, N2050, N1253, N735, N543);
or OR4 (N2055, N2025, N87, N655, N1547);
xor XOR2 (N2056, N2054, N1371);
not NOT1 (N2057, N2032);
nand NAND4 (N2058, N2056, N184, N1610, N562);
nor NOR4 (N2059, N2057, N1633, N878, N1910);
nand NAND4 (N2060, N2047, N715, N1650, N935);
or OR3 (N2061, N2040, N9, N1623);
not NOT1 (N2062, N2053);
buf BUF1 (N2063, N2049);
xor XOR2 (N2064, N2058, N332);
buf BUF1 (N2065, N2063);
and AND4 (N2066, N2048, N2064, N532, N867);
nand NAND3 (N2067, N1473, N567, N1343);
not NOT1 (N2068, N2059);
buf BUF1 (N2069, N2061);
nand NAND2 (N2070, N2017, N1563);
nand NAND4 (N2071, N2070, N920, N238, N693);
not NOT1 (N2072, N2068);
nand NAND3 (N2073, N2055, N236, N557);
nor NOR3 (N2074, N2071, N1161, N1760);
nand NAND4 (N2075, N2073, N293, N704, N371);
nand NAND4 (N2076, N2069, N1316, N121, N965);
or OR2 (N2077, N2075, N301);
not NOT1 (N2078, N2077);
buf BUF1 (N2079, N2074);
nand NAND3 (N2080, N2062, N1820, N369);
buf BUF1 (N2081, N2078);
xor XOR2 (N2082, N2072, N708);
not NOT1 (N2083, N2079);
or OR4 (N2084, N2081, N1401, N2026, N588);
xor XOR2 (N2085, N2067, N1698);
nor NOR3 (N2086, N2076, N1748, N951);
nor NOR4 (N2087, N2080, N85, N1274, N1);
not NOT1 (N2088, N2087);
nor NOR4 (N2089, N2052, N607, N507, N1746);
nor NOR2 (N2090, N2065, N1808);
nand NAND2 (N2091, N2060, N1119);
and AND2 (N2092, N2086, N1795);
and AND2 (N2093, N2082, N1018);
not NOT1 (N2094, N2084);
not NOT1 (N2095, N2088);
and AND3 (N2096, N2083, N377, N684);
nand NAND2 (N2097, N2092, N1456);
nand NAND3 (N2098, N2095, N459, N1671);
and AND2 (N2099, N2089, N1264);
not NOT1 (N2100, N2090);
nand NAND2 (N2101, N2097, N1724);
buf BUF1 (N2102, N2094);
not NOT1 (N2103, N2093);
buf BUF1 (N2104, N2102);
not NOT1 (N2105, N2096);
and AND4 (N2106, N2099, N2012, N1503, N263);
or OR2 (N2107, N2105, N603);
nand NAND2 (N2108, N2100, N722);
xor XOR2 (N2109, N2091, N1655);
not NOT1 (N2110, N2085);
buf BUF1 (N2111, N2108);
or OR4 (N2112, N2098, N2007, N1961, N800);
nor NOR2 (N2113, N2111, N182);
buf BUF1 (N2114, N2112);
nand NAND3 (N2115, N2101, N1770, N270);
nand NAND3 (N2116, N2115, N936, N1485);
nand NAND3 (N2117, N2110, N1479, N2044);
xor XOR2 (N2118, N2116, N942);
xor XOR2 (N2119, N2106, N28);
nor NOR3 (N2120, N2107, N1582, N207);
not NOT1 (N2121, N2104);
nor NOR2 (N2122, N2121, N2024);
nor NOR4 (N2123, N2109, N1822, N1269, N735);
not NOT1 (N2124, N2114);
or OR4 (N2125, N2117, N466, N1348, N1968);
or OR2 (N2126, N2122, N183);
or OR2 (N2127, N2123, N1925);
not NOT1 (N2128, N2113);
xor XOR2 (N2129, N2127, N309);
xor XOR2 (N2130, N2125, N1579);
buf BUF1 (N2131, N2128);
nand NAND4 (N2132, N2124, N761, N32, N295);
buf BUF1 (N2133, N2066);
and AND2 (N2134, N2118, N1357);
not NOT1 (N2135, N2103);
buf BUF1 (N2136, N2119);
and AND3 (N2137, N2136, N980, N789);
buf BUF1 (N2138, N2131);
xor XOR2 (N2139, N2137, N1823);
not NOT1 (N2140, N2138);
or OR3 (N2141, N2134, N865, N1350);
buf BUF1 (N2142, N2135);
or OR2 (N2143, N2132, N1971);
xor XOR2 (N2144, N2140, N1226);
nand NAND2 (N2145, N2133, N107);
nand NAND4 (N2146, N2139, N784, N1368, N338);
nand NAND2 (N2147, N2141, N1273);
nor NOR3 (N2148, N2143, N1300, N1166);
and AND4 (N2149, N2145, N1592, N1999, N255);
and AND4 (N2150, N2126, N1139, N751, N1975);
xor XOR2 (N2151, N2144, N1490);
buf BUF1 (N2152, N2148);
nor NOR4 (N2153, N2120, N1704, N1184, N1086);
or OR3 (N2154, N2153, N2033, N1401);
nor NOR4 (N2155, N2147, N418, N912, N15);
nor NOR3 (N2156, N2155, N996, N418);
or OR4 (N2157, N2149, N763, N470, N1263);
and AND3 (N2158, N2142, N516, N1143);
nand NAND3 (N2159, N2151, N2061, N493);
xor XOR2 (N2160, N2150, N1908);
and AND3 (N2161, N2129, N1298, N1077);
and AND2 (N2162, N2130, N1003);
or OR2 (N2163, N2162, N1013);
or OR4 (N2164, N2146, N936, N289, N265);
buf BUF1 (N2165, N2158);
or OR4 (N2166, N2159, N1088, N1253, N1085);
and AND2 (N2167, N2165, N1860);
nor NOR2 (N2168, N2161, N839);
buf BUF1 (N2169, N2160);
or OR4 (N2170, N2169, N1423, N415, N1542);
nand NAND3 (N2171, N2156, N1340, N304);
or OR4 (N2172, N2168, N986, N1642, N1723);
buf BUF1 (N2173, N2163);
xor XOR2 (N2174, N2172, N1623);
or OR4 (N2175, N2170, N1399, N573, N939);
or OR3 (N2176, N2173, N374, N1570);
buf BUF1 (N2177, N2171);
and AND2 (N2178, N2177, N1767);
xor XOR2 (N2179, N2178, N426);
buf BUF1 (N2180, N2179);
nor NOR2 (N2181, N2166, N467);
not NOT1 (N2182, N2175);
and AND2 (N2183, N2180, N469);
or OR3 (N2184, N2176, N1585, N1942);
buf BUF1 (N2185, N2184);
or OR4 (N2186, N2152, N1153, N549, N1726);
buf BUF1 (N2187, N2167);
xor XOR2 (N2188, N2187, N905);
nand NAND3 (N2189, N2157, N297, N548);
or OR3 (N2190, N2189, N1169, N1340);
nor NOR2 (N2191, N2154, N1968);
and AND2 (N2192, N2174, N1911);
or OR3 (N2193, N2190, N2159, N557);
and AND3 (N2194, N2188, N447, N195);
not NOT1 (N2195, N2185);
or OR4 (N2196, N2192, N1756, N328, N347);
or OR4 (N2197, N2182, N655, N176, N2075);
xor XOR2 (N2198, N2164, N1515);
xor XOR2 (N2199, N2181, N527);
not NOT1 (N2200, N2191);
xor XOR2 (N2201, N2200, N2160);
nor NOR4 (N2202, N2196, N1979, N1841, N267);
buf BUF1 (N2203, N2197);
not NOT1 (N2204, N2193);
or OR3 (N2205, N2202, N1911, N615);
not NOT1 (N2206, N2204);
or OR4 (N2207, N2199, N852, N901, N1748);
xor XOR2 (N2208, N2206, N1615);
nor NOR4 (N2209, N2198, N365, N609, N972);
nor NOR3 (N2210, N2186, N656, N1436);
nor NOR3 (N2211, N2207, N1639, N1532);
not NOT1 (N2212, N2205);
xor XOR2 (N2213, N2210, N943);
nor NOR3 (N2214, N2201, N1785, N1268);
not NOT1 (N2215, N2208);
xor XOR2 (N2216, N2209, N186);
nand NAND3 (N2217, N2194, N732, N1090);
xor XOR2 (N2218, N2215, N1792);
and AND3 (N2219, N2211, N1256, N1963);
buf BUF1 (N2220, N2213);
or OR3 (N2221, N2220, N1795, N2077);
or OR2 (N2222, N2195, N1949);
nand NAND2 (N2223, N2219, N1226);
nand NAND2 (N2224, N2212, N1831);
nand NAND2 (N2225, N2221, N1045);
xor XOR2 (N2226, N2183, N2056);
nor NOR2 (N2227, N2218, N840);
nor NOR3 (N2228, N2214, N2036, N1032);
nand NAND3 (N2229, N2225, N1479, N1401);
nor NOR2 (N2230, N2227, N1164);
nand NAND2 (N2231, N2222, N895);
or OR3 (N2232, N2229, N1300, N511);
nand NAND2 (N2233, N2224, N1900);
not NOT1 (N2234, N2230);
nor NOR4 (N2235, N2203, N476, N857, N456);
buf BUF1 (N2236, N2232);
and AND2 (N2237, N2217, N687);
nand NAND2 (N2238, N2236, N1089);
nand NAND3 (N2239, N2228, N1605, N1727);
or OR3 (N2240, N2226, N579, N1154);
nor NOR4 (N2241, N2223, N1371, N410, N1192);
nor NOR4 (N2242, N2237, N1779, N543, N1740);
and AND2 (N2243, N2241, N2190);
buf BUF1 (N2244, N2238);
nand NAND2 (N2245, N2233, N635);
xor XOR2 (N2246, N2231, N897);
not NOT1 (N2247, N2243);
buf BUF1 (N2248, N2239);
not NOT1 (N2249, N2245);
nand NAND3 (N2250, N2234, N744, N323);
nand NAND3 (N2251, N2247, N117, N1861);
xor XOR2 (N2252, N2240, N644);
and AND4 (N2253, N2248, N1531, N264, N1264);
buf BUF1 (N2254, N2252);
not NOT1 (N2255, N2253);
nor NOR3 (N2256, N2244, N1961, N1182);
nand NAND4 (N2257, N2246, N566, N369, N997);
or OR4 (N2258, N2257, N1134, N1989, N2135);
xor XOR2 (N2259, N2258, N507);
not NOT1 (N2260, N2249);
not NOT1 (N2261, N2256);
not NOT1 (N2262, N2260);
not NOT1 (N2263, N2216);
nand NAND3 (N2264, N2254, N156, N329);
nand NAND2 (N2265, N2259, N2167);
or OR3 (N2266, N2265, N689, N1848);
buf BUF1 (N2267, N2261);
buf BUF1 (N2268, N2242);
or OR2 (N2269, N2263, N334);
buf BUF1 (N2270, N2262);
xor XOR2 (N2271, N2267, N1245);
buf BUF1 (N2272, N2271);
or OR2 (N2273, N2255, N137);
or OR2 (N2274, N2269, N1734);
nor NOR4 (N2275, N2266, N940, N1362, N242);
or OR3 (N2276, N2268, N2240, N1804);
not NOT1 (N2277, N2270);
buf BUF1 (N2278, N2277);
or OR2 (N2279, N2250, N1031);
or OR2 (N2280, N2278, N1196);
or OR3 (N2281, N2273, N656, N653);
and AND2 (N2282, N2264, N385);
xor XOR2 (N2283, N2282, N1464);
xor XOR2 (N2284, N2272, N1433);
nor NOR2 (N2285, N2251, N102);
nor NOR3 (N2286, N2284, N16, N828);
or OR3 (N2287, N2276, N2202, N948);
nand NAND2 (N2288, N2275, N1054);
or OR3 (N2289, N2281, N1554, N955);
and AND2 (N2290, N2287, N789);
or OR4 (N2291, N2289, N328, N321, N494);
and AND4 (N2292, N2285, N62, N567, N410);
nand NAND4 (N2293, N2286, N1615, N1110, N1202);
and AND2 (N2294, N2288, N1668);
or OR3 (N2295, N2293, N1569, N1392);
xor XOR2 (N2296, N2295, N1062);
xor XOR2 (N2297, N2274, N564);
or OR3 (N2298, N2291, N2174, N226);
and AND4 (N2299, N2235, N121, N58, N1241);
xor XOR2 (N2300, N2296, N596);
buf BUF1 (N2301, N2280);
nand NAND4 (N2302, N2300, N2130, N679, N862);
or OR4 (N2303, N2298, N1051, N354, N1913);
and AND4 (N2304, N2299, N2290, N344, N1112);
buf BUF1 (N2305, N2135);
nor NOR2 (N2306, N2292, N92);
xor XOR2 (N2307, N2305, N1082);
xor XOR2 (N2308, N2302, N1574);
nand NAND4 (N2309, N2308, N577, N1870, N1602);
nand NAND4 (N2310, N2307, N85, N2219, N1134);
and AND2 (N2311, N2306, N1712);
and AND3 (N2312, N2303, N422, N821);
or OR3 (N2313, N2279, N1771, N934);
nand NAND2 (N2314, N2301, N1776);
not NOT1 (N2315, N2314);
xor XOR2 (N2316, N2297, N7);
not NOT1 (N2317, N2312);
or OR4 (N2318, N2311, N2254, N111, N64);
and AND2 (N2319, N2283, N1814);
not NOT1 (N2320, N2319);
nand NAND3 (N2321, N2304, N969, N1719);
and AND3 (N2322, N2317, N1220, N2157);
or OR4 (N2323, N2318, N823, N2219, N979);
xor XOR2 (N2324, N2316, N795);
not NOT1 (N2325, N2315);
not NOT1 (N2326, N2310);
nor NOR4 (N2327, N2294, N1749, N1372, N1852);
and AND4 (N2328, N2323, N2080, N1772, N2195);
nor NOR3 (N2329, N2325, N2005, N51);
nand NAND4 (N2330, N2309, N642, N2050, N32);
xor XOR2 (N2331, N2321, N1174);
nor NOR2 (N2332, N2330, N441);
or OR3 (N2333, N2324, N1536, N1140);
or OR4 (N2334, N2327, N176, N522, N1391);
nand NAND2 (N2335, N2329, N369);
xor XOR2 (N2336, N2322, N273);
not NOT1 (N2337, N2328);
buf BUF1 (N2338, N2332);
buf BUF1 (N2339, N2313);
and AND2 (N2340, N2320, N2148);
and AND2 (N2341, N2340, N1279);
xor XOR2 (N2342, N2333, N1244);
xor XOR2 (N2343, N2337, N488);
and AND3 (N2344, N2343, N120, N1782);
nor NOR3 (N2345, N2344, N1570, N638);
xor XOR2 (N2346, N2342, N63);
nor NOR4 (N2347, N2331, N1419, N491, N102);
and AND2 (N2348, N2347, N946);
buf BUF1 (N2349, N2346);
nor NOR2 (N2350, N2349, N722);
or OR2 (N2351, N2339, N524);
nor NOR3 (N2352, N2350, N2301, N1766);
xor XOR2 (N2353, N2351, N633);
nand NAND4 (N2354, N2338, N1695, N82, N2109);
nand NAND2 (N2355, N2345, N1958);
not NOT1 (N2356, N2326);
nand NAND3 (N2357, N2352, N1360, N197);
or OR2 (N2358, N2336, N755);
or OR2 (N2359, N2341, N1411);
or OR2 (N2360, N2353, N928);
nor NOR2 (N2361, N2354, N2142);
and AND2 (N2362, N2335, N1135);
nor NOR2 (N2363, N2358, N750);
buf BUF1 (N2364, N2359);
nand NAND4 (N2365, N2364, N862, N634, N1558);
xor XOR2 (N2366, N2355, N258);
or OR4 (N2367, N2362, N1547, N2152, N2216);
xor XOR2 (N2368, N2366, N893);
not NOT1 (N2369, N2363);
nor NOR3 (N2370, N2368, N1976, N545);
buf BUF1 (N2371, N2370);
not NOT1 (N2372, N2334);
nand NAND4 (N2373, N2369, N292, N1805, N2026);
buf BUF1 (N2374, N2373);
not NOT1 (N2375, N2348);
or OR3 (N2376, N2374, N1662, N2339);
and AND4 (N2377, N2376, N1362, N1450, N2029);
not NOT1 (N2378, N2360);
nand NAND2 (N2379, N2367, N1335);
xor XOR2 (N2380, N2375, N2377);
nand NAND3 (N2381, N2353, N1025, N809);
xor XOR2 (N2382, N2380, N66);
nor NOR3 (N2383, N2372, N1694, N1654);
xor XOR2 (N2384, N2383, N1551);
xor XOR2 (N2385, N2378, N823);
not NOT1 (N2386, N2385);
buf BUF1 (N2387, N2384);
xor XOR2 (N2388, N2379, N2076);
or OR2 (N2389, N2381, N1077);
xor XOR2 (N2390, N2388, N1180);
xor XOR2 (N2391, N2361, N2375);
and AND2 (N2392, N2391, N1198);
or OR2 (N2393, N2356, N1799);
nand NAND2 (N2394, N2389, N73);
and AND2 (N2395, N2392, N2283);
and AND2 (N2396, N2390, N1243);
nor NOR2 (N2397, N2396, N2272);
xor XOR2 (N2398, N2371, N2076);
xor XOR2 (N2399, N2386, N1333);
not NOT1 (N2400, N2393);
or OR3 (N2401, N2382, N1115, N1851);
xor XOR2 (N2402, N2395, N13);
and AND2 (N2403, N2394, N178);
or OR2 (N2404, N2398, N472);
not NOT1 (N2405, N2402);
nand NAND3 (N2406, N2397, N803, N1862);
nor NOR3 (N2407, N2387, N1035, N814);
buf BUF1 (N2408, N2400);
and AND2 (N2409, N2407, N1693);
and AND2 (N2410, N2365, N324);
or OR3 (N2411, N2401, N2367, N1267);
nor NOR4 (N2412, N2403, N976, N1094, N799);
or OR2 (N2413, N2410, N14);
buf BUF1 (N2414, N2357);
nand NAND4 (N2415, N2411, N101, N1293, N1111);
or OR4 (N2416, N2409, N236, N311, N1120);
not NOT1 (N2417, N2408);
nand NAND3 (N2418, N2399, N105, N407);
nand NAND4 (N2419, N2413, N1342, N71, N789);
nor NOR2 (N2420, N2412, N275);
not NOT1 (N2421, N2406);
or OR4 (N2422, N2421, N876, N845, N773);
nor NOR3 (N2423, N2404, N1503, N1521);
buf BUF1 (N2424, N2423);
not NOT1 (N2425, N2417);
and AND2 (N2426, N2419, N2325);
not NOT1 (N2427, N2405);
nor NOR2 (N2428, N2414, N1892);
nand NAND4 (N2429, N2427, N1744, N233, N876);
nand NAND2 (N2430, N2424, N1452);
nand NAND4 (N2431, N2430, N1282, N1833, N1943);
nand NAND3 (N2432, N2420, N1283, N2261);
xor XOR2 (N2433, N2428, N1477);
nor NOR2 (N2434, N2433, N1303);
xor XOR2 (N2435, N2416, N1186);
xor XOR2 (N2436, N2431, N2358);
xor XOR2 (N2437, N2434, N78);
not NOT1 (N2438, N2436);
and AND4 (N2439, N2425, N647, N2268, N367);
buf BUF1 (N2440, N2437);
buf BUF1 (N2441, N2415);
nor NOR3 (N2442, N2429, N2188, N782);
and AND2 (N2443, N2432, N1427);
or OR2 (N2444, N2442, N1030);
or OR2 (N2445, N2443, N191);
or OR2 (N2446, N2444, N1744);
nor NOR3 (N2447, N2438, N253, N259);
and AND4 (N2448, N2445, N1068, N677, N43);
and AND2 (N2449, N2448, N1896);
xor XOR2 (N2450, N2418, N563);
xor XOR2 (N2451, N2440, N1936);
not NOT1 (N2452, N2435);
xor XOR2 (N2453, N2447, N386);
buf BUF1 (N2454, N2449);
nand NAND2 (N2455, N2451, N956);
or OR2 (N2456, N2446, N1830);
and AND2 (N2457, N2456, N166);
nor NOR2 (N2458, N2455, N797);
not NOT1 (N2459, N2422);
buf BUF1 (N2460, N2452);
buf BUF1 (N2461, N2457);
not NOT1 (N2462, N2458);
not NOT1 (N2463, N2459);
nand NAND4 (N2464, N2462, N2343, N1940, N1894);
buf BUF1 (N2465, N2464);
not NOT1 (N2466, N2426);
or OR4 (N2467, N2441, N1744, N1703, N1967);
xor XOR2 (N2468, N2453, N2428);
and AND3 (N2469, N2466, N1845, N186);
not NOT1 (N2470, N2469);
xor XOR2 (N2471, N2450, N1320);
and AND2 (N2472, N2470, N2425);
xor XOR2 (N2473, N2465, N491);
xor XOR2 (N2474, N2472, N1299);
nor NOR3 (N2475, N2474, N943, N694);
buf BUF1 (N2476, N2460);
and AND4 (N2477, N2473, N1385, N242, N2221);
or OR2 (N2478, N2467, N534);
or OR4 (N2479, N2471, N1152, N1584, N1695);
or OR4 (N2480, N2461, N2358, N77, N482);
or OR2 (N2481, N2476, N44);
buf BUF1 (N2482, N2454);
buf BUF1 (N2483, N2468);
nand NAND2 (N2484, N2475, N216);
not NOT1 (N2485, N2481);
not NOT1 (N2486, N2477);
nor NOR4 (N2487, N2479, N643, N141, N749);
nand NAND2 (N2488, N2482, N635);
and AND3 (N2489, N2439, N1745, N1966);
or OR4 (N2490, N2463, N360, N975, N1847);
or OR2 (N2491, N2490, N2108);
and AND2 (N2492, N2485, N2491);
or OR2 (N2493, N2464, N1430);
not NOT1 (N2494, N2489);
not NOT1 (N2495, N2484);
nor NOR3 (N2496, N2493, N47, N145);
nor NOR4 (N2497, N2478, N2452, N1695, N233);
and AND3 (N2498, N2486, N964, N1278);
buf BUF1 (N2499, N2480);
nand NAND2 (N2500, N2498, N1081);
xor XOR2 (N2501, N2496, N2006);
and AND4 (N2502, N2500, N696, N1361, N1667);
nand NAND4 (N2503, N2495, N2284, N1010, N2464);
buf BUF1 (N2504, N2503);
or OR2 (N2505, N2483, N746);
buf BUF1 (N2506, N2502);
not NOT1 (N2507, N2488);
xor XOR2 (N2508, N2501, N2320);
or OR3 (N2509, N2506, N1379, N1417);
or OR2 (N2510, N2494, N1365);
endmodule