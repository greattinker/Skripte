// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N6405,N6397,N6422,N6412,N6417,N6418,N6414,N6420,N6421,N6423;

buf BUF1 (N24, N19);
xor XOR2 (N25, N17, N2);
xor XOR2 (N26, N24, N24);
nand NAND4 (N27, N23, N9, N7, N12);
buf BUF1 (N28, N6);
or OR4 (N29, N23, N18, N22, N11);
or OR4 (N30, N12, N18, N11, N12);
nor NOR4 (N31, N19, N21, N3, N7);
or OR2 (N32, N12, N1);
not NOT1 (N33, N26);
xor XOR2 (N34, N3, N3);
buf BUF1 (N35, N5);
or OR4 (N36, N32, N6, N1, N18);
not NOT1 (N37, N33);
not NOT1 (N38, N28);
or OR4 (N39, N31, N17, N8, N2);
and AND4 (N40, N29, N12, N36, N39);
and AND3 (N41, N9, N18, N7);
buf BUF1 (N42, N1);
nor NOR3 (N43, N37, N24, N26);
nand NAND2 (N44, N27, N43);
nand NAND2 (N45, N16, N3);
buf BUF1 (N46, N42);
buf BUF1 (N47, N35);
and AND2 (N48, N30, N25);
nand NAND2 (N49, N32, N27);
and AND2 (N50, N40, N11);
nor NOR4 (N51, N46, N6, N49, N22);
and AND3 (N52, N45, N22, N11);
or OR2 (N53, N35, N30);
not NOT1 (N54, N34);
nor NOR4 (N55, N54, N12, N33, N44);
nor NOR4 (N56, N5, N13, N46, N46);
or OR3 (N57, N41, N54, N33);
nand NAND3 (N58, N50, N2, N56);
nor NOR4 (N59, N31, N27, N24, N33);
or OR3 (N60, N57, N52, N29);
not NOT1 (N61, N12);
or OR2 (N62, N61, N42);
xor XOR2 (N63, N51, N13);
and AND2 (N64, N53, N59);
not NOT1 (N65, N29);
nor NOR2 (N66, N60, N2);
not NOT1 (N67, N66);
not NOT1 (N68, N38);
nor NOR4 (N69, N55, N62, N17, N62);
nand NAND4 (N70, N9, N48, N2, N54);
xor XOR2 (N71, N14, N43);
buf BUF1 (N72, N65);
nand NAND4 (N73, N72, N3, N50, N10);
nand NAND3 (N74, N64, N34, N68);
nor NOR3 (N75, N52, N32, N42);
nand NAND3 (N76, N67, N50, N52);
nor NOR2 (N77, N76, N9);
nand NAND4 (N78, N63, N70, N75, N28);
nor NOR3 (N79, N27, N49, N21);
buf BUF1 (N80, N12);
xor XOR2 (N81, N78, N65);
xor XOR2 (N82, N69, N53);
buf BUF1 (N83, N77);
nor NOR3 (N84, N71, N30, N9);
and AND4 (N85, N74, N68, N58, N58);
xor XOR2 (N86, N41, N21);
or OR4 (N87, N86, N39, N28, N50);
buf BUF1 (N88, N87);
or OR2 (N89, N84, N65);
or OR3 (N90, N82, N74, N24);
not NOT1 (N91, N79);
buf BUF1 (N92, N91);
nor NOR2 (N93, N83, N35);
or OR4 (N94, N93, N91, N24, N20);
nor NOR3 (N95, N92, N85, N90);
buf BUF1 (N96, N12);
nand NAND2 (N97, N29, N85);
not NOT1 (N98, N81);
nor NOR2 (N99, N80, N7);
not NOT1 (N100, N89);
nand NAND4 (N101, N99, N55, N2, N91);
or OR4 (N102, N73, N10, N92, N54);
nor NOR4 (N103, N97, N18, N76, N96);
nor NOR4 (N104, N13, N33, N90, N51);
nand NAND3 (N105, N95, N16, N88);
and AND4 (N106, N102, N60, N66, N69);
buf BUF1 (N107, N95);
not NOT1 (N108, N106);
nand NAND3 (N109, N94, N36, N87);
and AND2 (N110, N101, N18);
not NOT1 (N111, N98);
nor NOR4 (N112, N100, N61, N18, N58);
not NOT1 (N113, N109);
and AND2 (N114, N107, N97);
not NOT1 (N115, N110);
not NOT1 (N116, N112);
nand NAND2 (N117, N116, N87);
xor XOR2 (N118, N115, N42);
nor NOR3 (N119, N105, N35, N98);
buf BUF1 (N120, N114);
and AND4 (N121, N120, N89, N100, N27);
nand NAND4 (N122, N108, N121, N108, N11);
nor NOR4 (N123, N55, N23, N68, N56);
nand NAND4 (N124, N118, N4, N4, N70);
and AND4 (N125, N117, N107, N90, N101);
nand NAND2 (N126, N119, N99);
or OR3 (N127, N47, N6, N25);
and AND4 (N128, N126, N107, N58, N87);
nor NOR2 (N129, N122, N126);
buf BUF1 (N130, N124);
and AND4 (N131, N127, N58, N74, N49);
nand NAND4 (N132, N129, N83, N101, N47);
xor XOR2 (N133, N128, N27);
and AND4 (N134, N111, N56, N49, N54);
buf BUF1 (N135, N131);
nand NAND2 (N136, N103, N80);
xor XOR2 (N137, N135, N34);
nor NOR4 (N138, N137, N126, N79, N44);
and AND3 (N139, N125, N23, N90);
and AND2 (N140, N130, N94);
nand NAND2 (N141, N133, N53);
not NOT1 (N142, N123);
nand NAND4 (N143, N138, N79, N43, N94);
xor XOR2 (N144, N139, N13);
buf BUF1 (N145, N132);
nand NAND4 (N146, N145, N47, N82, N107);
or OR3 (N147, N142, N105, N1);
xor XOR2 (N148, N134, N123);
not NOT1 (N149, N147);
nor NOR4 (N150, N149, N64, N76, N128);
xor XOR2 (N151, N140, N10);
nor NOR2 (N152, N143, N73);
buf BUF1 (N153, N144);
nand NAND2 (N154, N150, N65);
xor XOR2 (N155, N148, N142);
buf BUF1 (N156, N153);
nand NAND2 (N157, N151, N91);
not NOT1 (N158, N152);
not NOT1 (N159, N136);
or OR4 (N160, N156, N127, N47, N81);
nand NAND2 (N161, N154, N67);
xor XOR2 (N162, N159, N28);
nor NOR3 (N163, N158, N1, N70);
and AND4 (N164, N157, N1, N75, N58);
or OR4 (N165, N162, N66, N149, N133);
xor XOR2 (N166, N160, N17);
not NOT1 (N167, N113);
or OR2 (N168, N166, N6);
not NOT1 (N169, N168);
xor XOR2 (N170, N167, N93);
and AND3 (N171, N165, N131, N69);
not NOT1 (N172, N161);
nor NOR4 (N173, N172, N37, N117, N93);
and AND4 (N174, N104, N29, N20, N94);
not NOT1 (N175, N170);
or OR2 (N176, N141, N105);
not NOT1 (N177, N163);
buf BUF1 (N178, N173);
and AND4 (N179, N169, N131, N41, N109);
buf BUF1 (N180, N174);
nand NAND2 (N181, N180, N169);
or OR2 (N182, N155, N115);
not NOT1 (N183, N176);
xor XOR2 (N184, N178, N162);
not NOT1 (N185, N179);
xor XOR2 (N186, N175, N91);
or OR3 (N187, N183, N32, N79);
or OR2 (N188, N181, N32);
buf BUF1 (N189, N177);
buf BUF1 (N190, N146);
not NOT1 (N191, N164);
xor XOR2 (N192, N186, N7);
and AND3 (N193, N189, N180, N62);
nor NOR3 (N194, N171, N157, N144);
and AND2 (N195, N194, N180);
or OR3 (N196, N185, N101, N39);
or OR4 (N197, N195, N63, N114, N105);
xor XOR2 (N198, N193, N47);
and AND2 (N199, N188, N129);
nor NOR4 (N200, N192, N112, N11, N168);
nand NAND3 (N201, N198, N82, N189);
buf BUF1 (N202, N200);
nor NOR4 (N203, N196, N36, N135, N190);
not NOT1 (N204, N203);
nand NAND3 (N205, N15, N5, N144);
or OR2 (N206, N197, N125);
nor NOR3 (N207, N202, N115, N190);
buf BUF1 (N208, N182);
buf BUF1 (N209, N187);
buf BUF1 (N210, N207);
nor NOR3 (N211, N184, N41, N102);
buf BUF1 (N212, N201);
nor NOR3 (N213, N205, N87, N9);
nand NAND2 (N214, N213, N110);
not NOT1 (N215, N214);
and AND2 (N216, N209, N123);
buf BUF1 (N217, N208);
nor NOR2 (N218, N212, N197);
nor NOR3 (N219, N210, N52, N139);
nand NAND4 (N220, N204, N91, N91, N10);
xor XOR2 (N221, N206, N164);
or OR2 (N222, N199, N35);
nor NOR2 (N223, N217, N18);
not NOT1 (N224, N222);
buf BUF1 (N225, N218);
nand NAND4 (N226, N219, N187, N103, N125);
not NOT1 (N227, N211);
not NOT1 (N228, N227);
or OR4 (N229, N221, N104, N122, N201);
or OR3 (N230, N223, N137, N189);
buf BUF1 (N231, N215);
and AND2 (N232, N224, N57);
xor XOR2 (N233, N216, N93);
not NOT1 (N234, N229);
xor XOR2 (N235, N230, N74);
not NOT1 (N236, N226);
or OR3 (N237, N191, N191, N36);
or OR2 (N238, N233, N133);
or OR3 (N239, N232, N171, N100);
nand NAND3 (N240, N228, N154, N184);
buf BUF1 (N241, N235);
buf BUF1 (N242, N238);
nor NOR4 (N243, N225, N79, N27, N38);
buf BUF1 (N244, N234);
buf BUF1 (N245, N239);
or OR2 (N246, N244, N68);
not NOT1 (N247, N240);
and AND2 (N248, N243, N172);
or OR2 (N249, N246, N139);
not NOT1 (N250, N220);
buf BUF1 (N251, N250);
not NOT1 (N252, N249);
xor XOR2 (N253, N241, N245);
buf BUF1 (N254, N17);
or OR2 (N255, N248, N29);
buf BUF1 (N256, N251);
or OR4 (N257, N254, N164, N3, N145);
buf BUF1 (N258, N252);
not NOT1 (N259, N242);
not NOT1 (N260, N253);
or OR4 (N261, N256, N8, N119, N80);
and AND4 (N262, N260, N100, N112, N251);
xor XOR2 (N263, N255, N220);
xor XOR2 (N264, N259, N260);
nor NOR3 (N265, N262, N167, N213);
and AND2 (N266, N257, N125);
or OR4 (N267, N258, N209, N107, N251);
or OR4 (N268, N265, N230, N262, N21);
not NOT1 (N269, N263);
not NOT1 (N270, N247);
buf BUF1 (N271, N268);
buf BUF1 (N272, N261);
nor NOR2 (N273, N237, N250);
buf BUF1 (N274, N236);
not NOT1 (N275, N270);
buf BUF1 (N276, N272);
and AND4 (N277, N269, N80, N156, N58);
buf BUF1 (N278, N273);
and AND2 (N279, N231, N146);
nor NOR3 (N280, N275, N253, N83);
buf BUF1 (N281, N278);
or OR2 (N282, N271, N137);
buf BUF1 (N283, N280);
not NOT1 (N284, N281);
xor XOR2 (N285, N276, N27);
xor XOR2 (N286, N266, N97);
nand NAND3 (N287, N267, N114, N83);
nor NOR3 (N288, N286, N20, N161);
or OR4 (N289, N287, N183, N21, N67);
nand NAND4 (N290, N285, N40, N189, N222);
and AND3 (N291, N288, N80, N98);
not NOT1 (N292, N282);
and AND3 (N293, N289, N43, N132);
xor XOR2 (N294, N284, N123);
and AND3 (N295, N293, N111, N116);
not NOT1 (N296, N283);
xor XOR2 (N297, N292, N91);
buf BUF1 (N298, N296);
xor XOR2 (N299, N264, N82);
and AND4 (N300, N291, N188, N23, N119);
buf BUF1 (N301, N299);
not NOT1 (N302, N295);
and AND3 (N303, N277, N25, N241);
xor XOR2 (N304, N297, N214);
or OR4 (N305, N279, N9, N157, N118);
nand NAND4 (N306, N274, N186, N227, N171);
nor NOR2 (N307, N294, N5);
not NOT1 (N308, N306);
not NOT1 (N309, N298);
nand NAND4 (N310, N309, N264, N239, N112);
buf BUF1 (N311, N303);
nand NAND3 (N312, N290, N212, N88);
xor XOR2 (N313, N304, N4);
nand NAND4 (N314, N300, N49, N73, N58);
not NOT1 (N315, N314);
or OR3 (N316, N302, N30, N177);
xor XOR2 (N317, N315, N24);
nor NOR2 (N318, N305, N130);
buf BUF1 (N319, N313);
buf BUF1 (N320, N316);
and AND4 (N321, N307, N153, N197, N185);
or OR3 (N322, N301, N46, N52);
buf BUF1 (N323, N311);
nand NAND3 (N324, N321, N174, N306);
xor XOR2 (N325, N324, N172);
buf BUF1 (N326, N323);
buf BUF1 (N327, N320);
xor XOR2 (N328, N312, N154);
and AND3 (N329, N310, N27, N62);
nor NOR2 (N330, N326, N125);
nor NOR3 (N331, N318, N159, N323);
or OR4 (N332, N331, N277, N278, N160);
nor NOR2 (N333, N330, N327);
xor XOR2 (N334, N121, N147);
and AND3 (N335, N329, N68, N188);
and AND4 (N336, N322, N146, N113, N292);
nor NOR2 (N337, N332, N144);
nor NOR3 (N338, N336, N334, N330);
buf BUF1 (N339, N273);
nand NAND4 (N340, N319, N132, N74, N312);
nor NOR2 (N341, N317, N230);
and AND4 (N342, N333, N28, N62, N143);
buf BUF1 (N343, N328);
nor NOR4 (N344, N335, N88, N315, N9);
nor NOR4 (N345, N340, N259, N251, N196);
or OR4 (N346, N325, N124, N330, N140);
or OR3 (N347, N345, N251, N21);
buf BUF1 (N348, N344);
and AND2 (N349, N342, N264);
xor XOR2 (N350, N308, N280);
buf BUF1 (N351, N341);
xor XOR2 (N352, N350, N50);
and AND3 (N353, N351, N150, N33);
xor XOR2 (N354, N337, N127);
and AND3 (N355, N338, N211, N137);
nor NOR3 (N356, N353, N146, N156);
nand NAND2 (N357, N346, N300);
xor XOR2 (N358, N356, N253);
nand NAND3 (N359, N354, N292, N215);
xor XOR2 (N360, N349, N150);
and AND3 (N361, N355, N354, N333);
nor NOR2 (N362, N343, N15);
or OR2 (N363, N347, N217);
nor NOR4 (N364, N339, N301, N167, N205);
nand NAND3 (N365, N362, N198, N331);
nand NAND2 (N366, N365, N290);
or OR2 (N367, N348, N137);
buf BUF1 (N368, N363);
and AND3 (N369, N366, N295, N228);
nand NAND3 (N370, N369, N348, N284);
and AND4 (N371, N360, N32, N134, N296);
or OR3 (N372, N371, N320, N307);
not NOT1 (N373, N357);
nand NAND2 (N374, N373, N129);
not NOT1 (N375, N372);
buf BUF1 (N376, N375);
not NOT1 (N377, N359);
nand NAND3 (N378, N358, N326, N93);
xor XOR2 (N379, N374, N99);
nor NOR3 (N380, N368, N43, N236);
buf BUF1 (N381, N364);
xor XOR2 (N382, N377, N372);
and AND2 (N383, N370, N154);
not NOT1 (N384, N367);
buf BUF1 (N385, N361);
buf BUF1 (N386, N378);
xor XOR2 (N387, N386, N190);
not NOT1 (N388, N381);
nand NAND2 (N389, N382, N368);
nand NAND3 (N390, N379, N212, N212);
buf BUF1 (N391, N380);
or OR3 (N392, N391, N295, N376);
buf BUF1 (N393, N355);
not NOT1 (N394, N388);
or OR2 (N395, N385, N343);
not NOT1 (N396, N384);
nor NOR2 (N397, N395, N151);
nand NAND3 (N398, N393, N300, N337);
or OR2 (N399, N398, N278);
xor XOR2 (N400, N387, N209);
or OR3 (N401, N352, N179, N377);
nor NOR3 (N402, N400, N268, N82);
or OR3 (N403, N402, N393, N159);
and AND4 (N404, N396, N276, N3, N46);
xor XOR2 (N405, N404, N188);
buf BUF1 (N406, N389);
and AND3 (N407, N392, N82, N171);
nor NOR2 (N408, N406, N95);
or OR3 (N409, N390, N366, N396);
nand NAND4 (N410, N394, N174, N252, N342);
not NOT1 (N411, N383);
nor NOR3 (N412, N405, N258, N268);
and AND3 (N413, N408, N275, N359);
nand NAND4 (N414, N399, N384, N253, N246);
buf BUF1 (N415, N412);
not NOT1 (N416, N410);
buf BUF1 (N417, N407);
or OR3 (N418, N403, N286, N292);
and AND4 (N419, N397, N54, N124, N403);
nor NOR3 (N420, N414, N50, N77);
nor NOR4 (N421, N401, N83, N406, N377);
nor NOR2 (N422, N419, N347);
or OR4 (N423, N422, N185, N103, N296);
nor NOR4 (N424, N417, N232, N231, N38);
or OR2 (N425, N415, N340);
xor XOR2 (N426, N411, N262);
xor XOR2 (N427, N409, N396);
nand NAND3 (N428, N427, N362, N25);
not NOT1 (N429, N421);
or OR2 (N430, N416, N425);
nand NAND2 (N431, N374, N116);
xor XOR2 (N432, N424, N262);
buf BUF1 (N433, N418);
nand NAND2 (N434, N426, N329);
and AND3 (N435, N432, N69, N159);
or OR2 (N436, N423, N287);
nand NAND4 (N437, N433, N18, N171, N159);
xor XOR2 (N438, N431, N108);
nand NAND3 (N439, N413, N424, N308);
nor NOR4 (N440, N439, N116, N148, N128);
xor XOR2 (N441, N429, N148);
nor NOR4 (N442, N438, N346, N330, N436);
xor XOR2 (N443, N90, N1);
nand NAND4 (N444, N434, N273, N7, N138);
and AND3 (N445, N442, N193, N154);
nor NOR4 (N446, N440, N359, N15, N202);
nand NAND4 (N447, N420, N301, N85, N222);
or OR4 (N448, N428, N148, N242, N262);
not NOT1 (N449, N447);
not NOT1 (N450, N437);
not NOT1 (N451, N441);
and AND4 (N452, N430, N387, N381, N408);
and AND4 (N453, N450, N355, N97, N447);
buf BUF1 (N454, N451);
nand NAND2 (N455, N454, N376);
xor XOR2 (N456, N435, N246);
nand NAND4 (N457, N452, N102, N139, N396);
and AND4 (N458, N448, N394, N159, N153);
not NOT1 (N459, N443);
or OR4 (N460, N444, N317, N155, N443);
xor XOR2 (N461, N460, N334);
buf BUF1 (N462, N456);
buf BUF1 (N463, N449);
nand NAND3 (N464, N455, N219, N60);
not NOT1 (N465, N458);
xor XOR2 (N466, N453, N435);
xor XOR2 (N467, N463, N333);
nor NOR4 (N468, N466, N241, N75, N244);
nand NAND4 (N469, N464, N54, N332, N394);
nand NAND4 (N470, N465, N66, N136, N273);
or OR4 (N471, N457, N248, N169, N288);
or OR4 (N472, N461, N411, N398, N170);
buf BUF1 (N473, N470);
and AND2 (N474, N446, N457);
buf BUF1 (N475, N459);
not NOT1 (N476, N475);
xor XOR2 (N477, N462, N12);
not NOT1 (N478, N476);
and AND3 (N479, N472, N405, N13);
nand NAND4 (N480, N477, N75, N411, N300);
or OR4 (N481, N445, N22, N74, N265);
buf BUF1 (N482, N473);
buf BUF1 (N483, N481);
nor NOR2 (N484, N468, N24);
or OR2 (N485, N469, N39);
buf BUF1 (N486, N485);
buf BUF1 (N487, N483);
nand NAND3 (N488, N478, N484, N244);
xor XOR2 (N489, N379, N348);
not NOT1 (N490, N482);
buf BUF1 (N491, N467);
and AND3 (N492, N486, N150, N89);
xor XOR2 (N493, N487, N112);
nor NOR3 (N494, N489, N392, N203);
not NOT1 (N495, N492);
and AND4 (N496, N480, N320, N203, N417);
xor XOR2 (N497, N496, N188);
xor XOR2 (N498, N488, N286);
nor NOR3 (N499, N494, N428, N401);
nand NAND4 (N500, N471, N458, N278, N309);
or OR4 (N501, N479, N94, N110, N485);
or OR3 (N502, N495, N224, N411);
and AND2 (N503, N491, N278);
xor XOR2 (N504, N498, N365);
xor XOR2 (N505, N500, N409);
or OR4 (N506, N497, N129, N284, N453);
nor NOR2 (N507, N503, N402);
buf BUF1 (N508, N504);
nand NAND4 (N509, N508, N373, N12, N122);
nor NOR2 (N510, N505, N466);
buf BUF1 (N511, N502);
xor XOR2 (N512, N511, N306);
or OR4 (N513, N510, N165, N412, N313);
nand NAND4 (N514, N499, N34, N122, N121);
nor NOR2 (N515, N506, N364);
nor NOR2 (N516, N493, N149);
xor XOR2 (N517, N507, N235);
nor NOR4 (N518, N501, N116, N414, N222);
or OR2 (N519, N517, N124);
buf BUF1 (N520, N515);
not NOT1 (N521, N518);
buf BUF1 (N522, N519);
not NOT1 (N523, N520);
or OR3 (N524, N509, N97, N103);
nor NOR2 (N525, N512, N57);
not NOT1 (N526, N516);
not NOT1 (N527, N523);
nor NOR4 (N528, N527, N442, N29, N135);
xor XOR2 (N529, N528, N192);
and AND3 (N530, N490, N250, N257);
nand NAND2 (N531, N522, N457);
xor XOR2 (N532, N531, N312);
nand NAND3 (N533, N525, N158, N365);
buf BUF1 (N534, N532);
buf BUF1 (N535, N529);
not NOT1 (N536, N526);
and AND2 (N537, N534, N408);
xor XOR2 (N538, N521, N94);
xor XOR2 (N539, N536, N9);
or OR2 (N540, N537, N82);
buf BUF1 (N541, N514);
not NOT1 (N542, N513);
nor NOR2 (N543, N535, N58);
not NOT1 (N544, N533);
or OR2 (N545, N543, N250);
and AND2 (N546, N539, N528);
and AND3 (N547, N541, N539, N200);
or OR3 (N548, N542, N503, N337);
buf BUF1 (N549, N538);
nor NOR4 (N550, N547, N328, N275, N145);
nand NAND3 (N551, N550, N184, N435);
and AND3 (N552, N548, N479, N129);
nand NAND3 (N553, N530, N277, N491);
not NOT1 (N554, N544);
and AND2 (N555, N546, N295);
xor XOR2 (N556, N545, N196);
or OR2 (N557, N555, N381);
buf BUF1 (N558, N524);
not NOT1 (N559, N558);
nand NAND3 (N560, N552, N399, N201);
or OR3 (N561, N474, N419, N546);
buf BUF1 (N562, N557);
nor NOR4 (N563, N556, N120, N502, N444);
not NOT1 (N564, N540);
nand NAND2 (N565, N551, N412);
buf BUF1 (N566, N560);
buf BUF1 (N567, N564);
or OR3 (N568, N549, N387, N244);
nand NAND2 (N569, N559, N318);
or OR3 (N570, N553, N311, N58);
nand NAND3 (N571, N569, N564, N171);
and AND4 (N572, N565, N364, N349, N403);
or OR3 (N573, N568, N451, N315);
or OR2 (N574, N563, N468);
nand NAND4 (N575, N572, N358, N150, N247);
nor NOR3 (N576, N566, N516, N17);
and AND4 (N577, N570, N284, N457, N130);
xor XOR2 (N578, N574, N412);
nand NAND3 (N579, N573, N263, N304);
not NOT1 (N580, N579);
nor NOR2 (N581, N571, N419);
not NOT1 (N582, N567);
not NOT1 (N583, N554);
or OR4 (N584, N561, N482, N514, N326);
nand NAND4 (N585, N575, N361, N433, N459);
nor NOR2 (N586, N562, N388);
buf BUF1 (N587, N578);
and AND3 (N588, N587, N330, N569);
xor XOR2 (N589, N576, N58);
nor NOR3 (N590, N581, N524, N5);
and AND2 (N591, N584, N477);
nand NAND3 (N592, N588, N530, N309);
nor NOR3 (N593, N586, N396, N554);
and AND2 (N594, N577, N73);
xor XOR2 (N595, N585, N291);
nor NOR4 (N596, N593, N15, N65, N574);
buf BUF1 (N597, N592);
or OR2 (N598, N591, N330);
or OR2 (N599, N582, N400);
nor NOR2 (N600, N589, N326);
and AND3 (N601, N594, N509, N130);
and AND2 (N602, N601, N544);
or OR2 (N603, N583, N79);
not NOT1 (N604, N602);
buf BUF1 (N605, N604);
nor NOR3 (N606, N590, N256, N442);
nor NOR2 (N607, N598, N309);
nor NOR4 (N608, N597, N534, N288, N137);
nor NOR4 (N609, N607, N246, N37, N409);
xor XOR2 (N610, N606, N282);
nand NAND2 (N611, N603, N157);
nor NOR3 (N612, N611, N307, N366);
and AND4 (N613, N612, N401, N532, N61);
buf BUF1 (N614, N595);
or OR3 (N615, N613, N215, N465);
nand NAND4 (N616, N580, N79, N347, N475);
xor XOR2 (N617, N608, N399);
not NOT1 (N618, N610);
or OR4 (N619, N617, N142, N37, N551);
or OR4 (N620, N599, N483, N75, N356);
and AND3 (N621, N614, N539, N481);
not NOT1 (N622, N605);
and AND2 (N623, N600, N330);
nor NOR4 (N624, N621, N527, N260, N286);
and AND4 (N625, N618, N301, N450, N493);
or OR2 (N626, N624, N460);
not NOT1 (N627, N626);
xor XOR2 (N628, N609, N205);
and AND2 (N629, N628, N63);
or OR4 (N630, N616, N165, N250, N353);
buf BUF1 (N631, N625);
nor NOR2 (N632, N620, N257);
or OR3 (N633, N623, N171, N425);
and AND3 (N634, N632, N103, N40);
nand NAND2 (N635, N633, N123);
and AND4 (N636, N615, N458, N175, N288);
and AND3 (N637, N631, N194, N546);
or OR4 (N638, N629, N240, N374, N284);
or OR2 (N639, N635, N399);
nor NOR4 (N640, N637, N145, N61, N532);
nor NOR3 (N641, N622, N202, N576);
and AND3 (N642, N634, N235, N69);
not NOT1 (N643, N596);
nand NAND3 (N644, N639, N209, N159);
nor NOR4 (N645, N627, N557, N145, N88);
nand NAND4 (N646, N636, N441, N567, N90);
not NOT1 (N647, N630);
nand NAND2 (N648, N638, N563);
and AND2 (N649, N642, N393);
not NOT1 (N650, N648);
and AND3 (N651, N641, N631, N232);
nor NOR4 (N652, N644, N265, N409, N454);
xor XOR2 (N653, N651, N302);
and AND4 (N654, N652, N306, N379, N362);
not NOT1 (N655, N653);
buf BUF1 (N656, N645);
buf BUF1 (N657, N643);
buf BUF1 (N658, N646);
or OR4 (N659, N658, N632, N644, N480);
buf BUF1 (N660, N640);
nor NOR4 (N661, N647, N459, N328, N479);
nand NAND2 (N662, N660, N293);
or OR3 (N663, N661, N575, N545);
and AND2 (N664, N657, N455);
nand NAND4 (N665, N663, N598, N7, N352);
nand NAND3 (N666, N662, N362, N593);
and AND3 (N667, N664, N436, N291);
nor NOR4 (N668, N665, N376, N254, N606);
not NOT1 (N669, N649);
nand NAND4 (N670, N656, N377, N235, N195);
buf BUF1 (N671, N670);
nor NOR4 (N672, N655, N463, N217, N201);
and AND2 (N673, N654, N343);
or OR2 (N674, N667, N278);
buf BUF1 (N675, N668);
not NOT1 (N676, N650);
and AND2 (N677, N674, N173);
and AND3 (N678, N659, N648, N614);
and AND3 (N679, N676, N575, N527);
and AND3 (N680, N677, N419, N500);
and AND4 (N681, N666, N110, N188, N535);
not NOT1 (N682, N680);
nor NOR2 (N683, N673, N58);
xor XOR2 (N684, N681, N75);
nor NOR4 (N685, N679, N241, N238, N452);
buf BUF1 (N686, N675);
and AND4 (N687, N686, N77, N333, N139);
xor XOR2 (N688, N678, N295);
buf BUF1 (N689, N619);
buf BUF1 (N690, N687);
not NOT1 (N691, N683);
not NOT1 (N692, N691);
or OR2 (N693, N671, N609);
nand NAND2 (N694, N685, N225);
or OR4 (N695, N690, N661, N262, N441);
xor XOR2 (N696, N695, N580);
not NOT1 (N697, N669);
not NOT1 (N698, N697);
not NOT1 (N699, N694);
buf BUF1 (N700, N698);
not NOT1 (N701, N684);
and AND3 (N702, N696, N655, N540);
buf BUF1 (N703, N682);
nand NAND2 (N704, N699, N113);
buf BUF1 (N705, N702);
not NOT1 (N706, N689);
not NOT1 (N707, N688);
nand NAND2 (N708, N705, N29);
nand NAND3 (N709, N672, N464, N45);
not NOT1 (N710, N704);
nor NOR4 (N711, N700, N363, N532, N672);
xor XOR2 (N712, N711, N20);
and AND3 (N713, N709, N193, N491);
buf BUF1 (N714, N710);
nand NAND4 (N715, N706, N35, N240, N16);
not NOT1 (N716, N701);
nand NAND2 (N717, N703, N565);
not NOT1 (N718, N713);
and AND4 (N719, N692, N163, N222, N30);
xor XOR2 (N720, N716, N656);
buf BUF1 (N721, N718);
not NOT1 (N722, N721);
xor XOR2 (N723, N717, N562);
or OR4 (N724, N707, N343, N720, N448);
not NOT1 (N725, N195);
not NOT1 (N726, N693);
nand NAND4 (N727, N722, N171, N678, N265);
and AND2 (N728, N714, N390);
or OR2 (N729, N708, N498);
buf BUF1 (N730, N719);
nand NAND4 (N731, N723, N507, N597, N162);
or OR4 (N732, N724, N409, N299, N15);
buf BUF1 (N733, N729);
or OR4 (N734, N726, N233, N187, N711);
buf BUF1 (N735, N727);
not NOT1 (N736, N731);
not NOT1 (N737, N730);
or OR2 (N738, N734, N194);
and AND3 (N739, N725, N634, N339);
and AND3 (N740, N737, N567, N338);
nand NAND2 (N741, N733, N417);
buf BUF1 (N742, N736);
xor XOR2 (N743, N739, N267);
nor NOR3 (N744, N741, N609, N505);
and AND4 (N745, N740, N47, N187, N85);
xor XOR2 (N746, N744, N505);
nor NOR4 (N747, N728, N370, N122, N375);
or OR2 (N748, N747, N247);
nand NAND4 (N749, N742, N39, N237, N416);
nand NAND4 (N750, N743, N734, N473, N329);
buf BUF1 (N751, N738);
xor XOR2 (N752, N746, N191);
xor XOR2 (N753, N751, N179);
not NOT1 (N754, N712);
nand NAND4 (N755, N732, N685, N272, N45);
nor NOR4 (N756, N735, N360, N91, N119);
xor XOR2 (N757, N748, N503);
nor NOR2 (N758, N752, N69);
not NOT1 (N759, N749);
and AND2 (N760, N755, N551);
buf BUF1 (N761, N756);
xor XOR2 (N762, N754, N452);
nand NAND2 (N763, N760, N606);
or OR3 (N764, N757, N82, N314);
not NOT1 (N765, N763);
nand NAND2 (N766, N753, N226);
not NOT1 (N767, N715);
nand NAND3 (N768, N762, N651, N661);
buf BUF1 (N769, N759);
and AND2 (N770, N768, N131);
or OR4 (N771, N767, N174, N625, N255);
not NOT1 (N772, N745);
nand NAND4 (N773, N765, N19, N224, N549);
nor NOR4 (N774, N772, N314, N580, N52);
not NOT1 (N775, N774);
xor XOR2 (N776, N775, N489);
and AND3 (N777, N750, N431, N495);
and AND4 (N778, N764, N284, N727, N625);
not NOT1 (N779, N773);
and AND4 (N780, N771, N116, N617, N513);
nand NAND2 (N781, N779, N33);
xor XOR2 (N782, N780, N327);
buf BUF1 (N783, N776);
xor XOR2 (N784, N769, N670);
and AND2 (N785, N782, N32);
nand NAND3 (N786, N777, N586, N741);
nand NAND3 (N787, N770, N480, N55);
not NOT1 (N788, N784);
and AND3 (N789, N781, N673, N82);
not NOT1 (N790, N786);
xor XOR2 (N791, N778, N233);
xor XOR2 (N792, N758, N768);
and AND3 (N793, N766, N611, N415);
not NOT1 (N794, N788);
and AND4 (N795, N794, N305, N531, N581);
xor XOR2 (N796, N785, N270);
and AND2 (N797, N793, N165);
nand NAND2 (N798, N789, N115);
or OR2 (N799, N790, N163);
nor NOR2 (N800, N797, N779);
xor XOR2 (N801, N791, N230);
buf BUF1 (N802, N796);
xor XOR2 (N803, N795, N735);
or OR3 (N804, N798, N664, N533);
buf BUF1 (N805, N792);
xor XOR2 (N806, N802, N714);
nand NAND3 (N807, N804, N555, N645);
nand NAND4 (N808, N800, N162, N77, N397);
or OR2 (N809, N806, N727);
xor XOR2 (N810, N799, N309);
xor XOR2 (N811, N803, N436);
nand NAND4 (N812, N801, N724, N601, N63);
nor NOR2 (N813, N805, N386);
buf BUF1 (N814, N807);
xor XOR2 (N815, N761, N389);
xor XOR2 (N816, N813, N755);
not NOT1 (N817, N787);
buf BUF1 (N818, N812);
buf BUF1 (N819, N808);
xor XOR2 (N820, N816, N127);
not NOT1 (N821, N809);
not NOT1 (N822, N810);
or OR3 (N823, N811, N418, N118);
buf BUF1 (N824, N818);
or OR2 (N825, N824, N13);
buf BUF1 (N826, N783);
xor XOR2 (N827, N817, N657);
nand NAND4 (N828, N822, N753, N109, N470);
or OR3 (N829, N826, N357, N716);
xor XOR2 (N830, N828, N677);
nor NOR3 (N831, N820, N339, N194);
not NOT1 (N832, N829);
nand NAND2 (N833, N819, N311);
not NOT1 (N834, N833);
xor XOR2 (N835, N823, N630);
buf BUF1 (N836, N832);
and AND2 (N837, N836, N603);
buf BUF1 (N838, N825);
nand NAND3 (N839, N837, N404, N45);
nor NOR3 (N840, N830, N504, N354);
or OR4 (N841, N840, N152, N99, N624);
nor NOR4 (N842, N835, N377, N332, N722);
xor XOR2 (N843, N827, N798);
xor XOR2 (N844, N839, N802);
or OR3 (N845, N834, N384, N76);
buf BUF1 (N846, N845);
or OR4 (N847, N815, N468, N275, N767);
xor XOR2 (N848, N814, N797);
xor XOR2 (N849, N848, N648);
and AND4 (N850, N842, N345, N100, N196);
and AND3 (N851, N849, N34, N398);
nand NAND3 (N852, N851, N549, N592);
nor NOR4 (N853, N838, N216, N311, N770);
or OR4 (N854, N852, N626, N66, N813);
not NOT1 (N855, N854);
xor XOR2 (N856, N821, N505);
buf BUF1 (N857, N850);
not NOT1 (N858, N841);
nor NOR4 (N859, N844, N490, N257, N471);
nand NAND3 (N860, N831, N856, N800);
not NOT1 (N861, N169);
nor NOR3 (N862, N859, N488, N182);
buf BUF1 (N863, N861);
and AND3 (N864, N855, N776, N646);
and AND2 (N865, N858, N382);
not NOT1 (N866, N864);
nand NAND4 (N867, N853, N734, N591, N386);
and AND3 (N868, N865, N471, N864);
buf BUF1 (N869, N843);
xor XOR2 (N870, N868, N804);
and AND2 (N871, N870, N608);
nor NOR3 (N872, N866, N231, N827);
or OR2 (N873, N863, N449);
buf BUF1 (N874, N869);
buf BUF1 (N875, N871);
and AND3 (N876, N875, N364, N49);
nand NAND4 (N877, N860, N543, N451, N741);
or OR4 (N878, N872, N518, N535, N42);
xor XOR2 (N879, N846, N577);
or OR3 (N880, N874, N396, N742);
not NOT1 (N881, N880);
and AND4 (N882, N881, N454, N765, N368);
xor XOR2 (N883, N882, N20);
or OR4 (N884, N862, N46, N747, N294);
not NOT1 (N885, N879);
buf BUF1 (N886, N883);
and AND3 (N887, N885, N520, N248);
nor NOR3 (N888, N847, N194, N852);
or OR3 (N889, N857, N764, N578);
not NOT1 (N890, N873);
buf BUF1 (N891, N876);
not NOT1 (N892, N887);
or OR3 (N893, N892, N476, N282);
or OR2 (N894, N884, N519);
or OR2 (N895, N890, N801);
not NOT1 (N896, N886);
and AND3 (N897, N867, N777, N779);
buf BUF1 (N898, N894);
xor XOR2 (N899, N895, N691);
and AND2 (N900, N896, N326);
and AND3 (N901, N897, N55, N26);
nor NOR4 (N902, N901, N457, N851, N637);
and AND4 (N903, N878, N470, N502, N265);
and AND4 (N904, N889, N69, N301, N72);
buf BUF1 (N905, N900);
xor XOR2 (N906, N899, N803);
and AND3 (N907, N891, N696, N32);
and AND3 (N908, N902, N747, N302);
or OR4 (N909, N905, N853, N189, N94);
xor XOR2 (N910, N907, N335);
xor XOR2 (N911, N877, N54);
xor XOR2 (N912, N909, N679);
not NOT1 (N913, N910);
nand NAND2 (N914, N903, N910);
nor NOR2 (N915, N912, N446);
buf BUF1 (N916, N898);
nand NAND4 (N917, N893, N525, N68, N133);
or OR4 (N918, N914, N374, N822, N717);
nor NOR2 (N919, N906, N154);
not NOT1 (N920, N908);
nand NAND4 (N921, N904, N181, N33, N552);
not NOT1 (N922, N888);
nand NAND2 (N923, N919, N383);
xor XOR2 (N924, N918, N232);
xor XOR2 (N925, N922, N39);
xor XOR2 (N926, N925, N371);
not NOT1 (N927, N921);
nand NAND2 (N928, N911, N136);
or OR3 (N929, N927, N240, N117);
buf BUF1 (N930, N917);
or OR2 (N931, N928, N642);
not NOT1 (N932, N924);
buf BUF1 (N933, N923);
not NOT1 (N934, N913);
nand NAND2 (N935, N933, N615);
nand NAND2 (N936, N915, N353);
or OR3 (N937, N930, N662, N161);
xor XOR2 (N938, N935, N621);
or OR4 (N939, N936, N223, N937, N885);
buf BUF1 (N940, N508);
and AND3 (N941, N929, N229, N474);
buf BUF1 (N942, N939);
nand NAND2 (N943, N932, N500);
not NOT1 (N944, N920);
not NOT1 (N945, N943);
buf BUF1 (N946, N944);
xor XOR2 (N947, N942, N841);
not NOT1 (N948, N945);
and AND2 (N949, N948, N66);
buf BUF1 (N950, N934);
and AND2 (N951, N949, N769);
xor XOR2 (N952, N950, N210);
buf BUF1 (N953, N926);
buf BUF1 (N954, N938);
xor XOR2 (N955, N947, N299);
nand NAND3 (N956, N954, N798, N441);
nor NOR4 (N957, N956, N4, N360, N214);
not NOT1 (N958, N946);
or OR4 (N959, N955, N66, N687, N257);
xor XOR2 (N960, N916, N808);
nor NOR2 (N961, N960, N714);
and AND2 (N962, N951, N293);
buf BUF1 (N963, N952);
buf BUF1 (N964, N958);
buf BUF1 (N965, N940);
not NOT1 (N966, N961);
and AND4 (N967, N959, N324, N379, N557);
not NOT1 (N968, N963);
nand NAND2 (N969, N964, N650);
not NOT1 (N970, N968);
not NOT1 (N971, N941);
buf BUF1 (N972, N969);
buf BUF1 (N973, N970);
buf BUF1 (N974, N962);
nand NAND3 (N975, N971, N643, N234);
buf BUF1 (N976, N931);
or OR4 (N977, N973, N396, N147, N60);
xor XOR2 (N978, N966, N599);
not NOT1 (N979, N965);
buf BUF1 (N980, N977);
buf BUF1 (N981, N953);
and AND4 (N982, N975, N256, N341, N249);
nor NOR4 (N983, N978, N354, N923, N307);
nor NOR2 (N984, N981, N256);
not NOT1 (N985, N980);
buf BUF1 (N986, N979);
or OR4 (N987, N967, N342, N821, N249);
buf BUF1 (N988, N982);
buf BUF1 (N989, N984);
buf BUF1 (N990, N983);
and AND2 (N991, N986, N121);
nand NAND4 (N992, N972, N497, N748, N860);
nor NOR4 (N993, N988, N385, N583, N850);
nor NOR2 (N994, N957, N544);
buf BUF1 (N995, N976);
not NOT1 (N996, N993);
and AND3 (N997, N995, N441, N613);
and AND4 (N998, N974, N827, N377, N131);
nor NOR4 (N999, N996, N536, N349, N628);
buf BUF1 (N1000, N992);
buf BUF1 (N1001, N985);
and AND2 (N1002, N987, N183);
nand NAND2 (N1003, N1002, N745);
or OR2 (N1004, N989, N633);
and AND3 (N1005, N997, N695, N9);
xor XOR2 (N1006, N990, N771);
xor XOR2 (N1007, N1000, N454);
and AND3 (N1008, N999, N771, N834);
xor XOR2 (N1009, N1004, N974);
or OR3 (N1010, N1007, N384, N1009);
and AND3 (N1011, N424, N971, N391);
and AND2 (N1012, N1010, N941);
or OR4 (N1013, N1003, N32, N423, N928);
not NOT1 (N1014, N998);
or OR4 (N1015, N1012, N862, N641, N151);
buf BUF1 (N1016, N1005);
or OR2 (N1017, N994, N256);
not NOT1 (N1018, N1011);
or OR3 (N1019, N1013, N801, N98);
buf BUF1 (N1020, N1019);
nor NOR4 (N1021, N1016, N698, N787, N814);
or OR2 (N1022, N1018, N1002);
buf BUF1 (N1023, N991);
nand NAND3 (N1024, N1021, N880, N304);
nand NAND2 (N1025, N1022, N1004);
nor NOR2 (N1026, N1006, N898);
and AND4 (N1027, N1017, N208, N55, N432);
and AND4 (N1028, N1020, N33, N535, N37);
or OR2 (N1029, N1001, N924);
and AND2 (N1030, N1029, N744);
xor XOR2 (N1031, N1014, N840);
and AND4 (N1032, N1030, N856, N157, N54);
nand NAND2 (N1033, N1015, N338);
or OR4 (N1034, N1023, N776, N259, N382);
xor XOR2 (N1035, N1032, N668);
nand NAND4 (N1036, N1008, N752, N958, N333);
or OR3 (N1037, N1028, N414, N969);
not NOT1 (N1038, N1035);
and AND2 (N1039, N1037, N127);
or OR3 (N1040, N1031, N640, N485);
not NOT1 (N1041, N1025);
xor XOR2 (N1042, N1034, N704);
buf BUF1 (N1043, N1026);
nand NAND2 (N1044, N1039, N91);
nand NAND3 (N1045, N1027, N399, N540);
buf BUF1 (N1046, N1044);
xor XOR2 (N1047, N1036, N36);
or OR4 (N1048, N1046, N529, N407, N179);
nor NOR4 (N1049, N1041, N104, N910, N494);
buf BUF1 (N1050, N1033);
nor NOR4 (N1051, N1040, N734, N655, N420);
xor XOR2 (N1052, N1038, N706);
not NOT1 (N1053, N1052);
buf BUF1 (N1054, N1051);
buf BUF1 (N1055, N1047);
nand NAND3 (N1056, N1053, N239, N809);
and AND2 (N1057, N1048, N873);
buf BUF1 (N1058, N1055);
nor NOR2 (N1059, N1057, N505);
nor NOR4 (N1060, N1059, N492, N207, N618);
and AND4 (N1061, N1054, N109, N48, N9);
not NOT1 (N1062, N1061);
or OR2 (N1063, N1060, N1000);
nor NOR4 (N1064, N1045, N827, N1001, N658);
xor XOR2 (N1065, N1058, N104);
buf BUF1 (N1066, N1049);
or OR2 (N1067, N1065, N448);
nor NOR3 (N1068, N1043, N542, N21);
buf BUF1 (N1069, N1056);
not NOT1 (N1070, N1069);
buf BUF1 (N1071, N1024);
nand NAND4 (N1072, N1071, N845, N841, N80);
and AND2 (N1073, N1067, N152);
nor NOR3 (N1074, N1068, N270, N621);
xor XOR2 (N1075, N1064, N722);
buf BUF1 (N1076, N1075);
nand NAND3 (N1077, N1076, N739, N1004);
nand NAND4 (N1078, N1077, N492, N398, N581);
not NOT1 (N1079, N1066);
nand NAND3 (N1080, N1050, N623, N446);
and AND4 (N1081, N1079, N327, N129, N832);
nor NOR4 (N1082, N1062, N687, N219, N511);
not NOT1 (N1083, N1080);
nand NAND3 (N1084, N1073, N1077, N567);
nor NOR4 (N1085, N1078, N1067, N749, N702);
nor NOR2 (N1086, N1072, N981);
nor NOR2 (N1087, N1081, N606);
nor NOR2 (N1088, N1063, N740);
nand NAND3 (N1089, N1088, N169, N655);
buf BUF1 (N1090, N1070);
nand NAND3 (N1091, N1074, N426, N530);
buf BUF1 (N1092, N1085);
not NOT1 (N1093, N1090);
not NOT1 (N1094, N1042);
and AND3 (N1095, N1094, N1089, N790);
xor XOR2 (N1096, N772, N822);
xor XOR2 (N1097, N1095, N151);
buf BUF1 (N1098, N1084);
xor XOR2 (N1099, N1092, N664);
xor XOR2 (N1100, N1098, N110);
xor XOR2 (N1101, N1100, N246);
buf BUF1 (N1102, N1091);
nor NOR4 (N1103, N1101, N316, N544, N832);
xor XOR2 (N1104, N1097, N257);
and AND3 (N1105, N1093, N750, N746);
buf BUF1 (N1106, N1099);
nand NAND2 (N1107, N1096, N995);
buf BUF1 (N1108, N1083);
or OR3 (N1109, N1106, N58, N810);
not NOT1 (N1110, N1107);
nor NOR3 (N1111, N1103, N398, N21);
not NOT1 (N1112, N1082);
nand NAND2 (N1113, N1110, N943);
buf BUF1 (N1114, N1111);
nor NOR3 (N1115, N1113, N131, N721);
nand NAND4 (N1116, N1109, N859, N224, N1091);
not NOT1 (N1117, N1115);
or OR3 (N1118, N1104, N1103, N36);
or OR3 (N1119, N1102, N1114, N632);
buf BUF1 (N1120, N1107);
buf BUF1 (N1121, N1086);
and AND4 (N1122, N1112, N627, N314, N847);
not NOT1 (N1123, N1118);
or OR4 (N1124, N1122, N321, N835, N134);
and AND4 (N1125, N1121, N187, N67, N721);
or OR4 (N1126, N1119, N567, N889, N517);
xor XOR2 (N1127, N1123, N1020);
nand NAND4 (N1128, N1116, N1027, N440, N1094);
not NOT1 (N1129, N1105);
not NOT1 (N1130, N1127);
nor NOR2 (N1131, N1108, N49);
xor XOR2 (N1132, N1130, N132);
or OR2 (N1133, N1125, N604);
not NOT1 (N1134, N1117);
nor NOR4 (N1135, N1120, N371, N1023, N746);
and AND2 (N1136, N1128, N1067);
and AND3 (N1137, N1134, N565, N10);
nand NAND3 (N1138, N1129, N666, N82);
and AND4 (N1139, N1131, N119, N66, N846);
nand NAND4 (N1140, N1136, N840, N376, N116);
and AND3 (N1141, N1135, N825, N834);
not NOT1 (N1142, N1124);
or OR3 (N1143, N1132, N194, N451);
xor XOR2 (N1144, N1133, N75);
nand NAND4 (N1145, N1137, N1101, N334, N1041);
not NOT1 (N1146, N1144);
nor NOR4 (N1147, N1142, N727, N109, N475);
nor NOR2 (N1148, N1140, N635);
buf BUF1 (N1149, N1126);
not NOT1 (N1150, N1146);
buf BUF1 (N1151, N1149);
or OR2 (N1152, N1139, N878);
or OR4 (N1153, N1138, N1111, N1087, N91);
nor NOR4 (N1154, N569, N742, N868, N193);
nand NAND2 (N1155, N1141, N962);
and AND3 (N1156, N1151, N582, N410);
xor XOR2 (N1157, N1148, N758);
nand NAND4 (N1158, N1153, N821, N195, N1155);
or OR3 (N1159, N162, N873, N924);
and AND3 (N1160, N1145, N22, N844);
nor NOR3 (N1161, N1143, N951, N960);
or OR2 (N1162, N1147, N136);
nand NAND2 (N1163, N1162, N171);
buf BUF1 (N1164, N1160);
not NOT1 (N1165, N1150);
and AND4 (N1166, N1165, N92, N560, N552);
or OR2 (N1167, N1156, N105);
buf BUF1 (N1168, N1167);
not NOT1 (N1169, N1161);
nor NOR4 (N1170, N1154, N916, N787, N119);
nand NAND3 (N1171, N1168, N1049, N1093);
xor XOR2 (N1172, N1152, N826);
nor NOR2 (N1173, N1172, N672);
buf BUF1 (N1174, N1170);
xor XOR2 (N1175, N1163, N337);
buf BUF1 (N1176, N1171);
or OR3 (N1177, N1176, N290, N409);
nand NAND4 (N1178, N1173, N414, N383, N354);
or OR2 (N1179, N1174, N1031);
nor NOR3 (N1180, N1158, N893, N882);
buf BUF1 (N1181, N1177);
buf BUF1 (N1182, N1159);
buf BUF1 (N1183, N1179);
and AND4 (N1184, N1182, N315, N106, N844);
nand NAND2 (N1185, N1175, N626);
nand NAND3 (N1186, N1184, N456, N417);
and AND3 (N1187, N1157, N982, N765);
and AND2 (N1188, N1186, N569);
not NOT1 (N1189, N1183);
not NOT1 (N1190, N1166);
not NOT1 (N1191, N1185);
xor XOR2 (N1192, N1188, N431);
nand NAND4 (N1193, N1187, N394, N100, N863);
xor XOR2 (N1194, N1193, N818);
not NOT1 (N1195, N1194);
not NOT1 (N1196, N1178);
or OR2 (N1197, N1196, N926);
buf BUF1 (N1198, N1190);
and AND3 (N1199, N1198, N1080, N636);
or OR2 (N1200, N1169, N434);
not NOT1 (N1201, N1197);
nand NAND2 (N1202, N1181, N179);
buf BUF1 (N1203, N1202);
nand NAND4 (N1204, N1201, N603, N941, N443);
or OR2 (N1205, N1189, N758);
buf BUF1 (N1206, N1180);
not NOT1 (N1207, N1206);
nand NAND3 (N1208, N1207, N258, N640);
and AND2 (N1209, N1208, N954);
or OR2 (N1210, N1203, N413);
not NOT1 (N1211, N1164);
xor XOR2 (N1212, N1210, N217);
xor XOR2 (N1213, N1200, N355);
not NOT1 (N1214, N1192);
and AND3 (N1215, N1213, N94, N1138);
xor XOR2 (N1216, N1191, N451);
and AND3 (N1217, N1211, N668, N629);
nor NOR2 (N1218, N1212, N1132);
nor NOR2 (N1219, N1214, N429);
xor XOR2 (N1220, N1195, N992);
or OR4 (N1221, N1220, N729, N1048, N1025);
and AND4 (N1222, N1205, N877, N205, N307);
buf BUF1 (N1223, N1222);
nand NAND3 (N1224, N1216, N772, N487);
or OR3 (N1225, N1217, N401, N251);
or OR2 (N1226, N1219, N332);
nor NOR3 (N1227, N1221, N745, N1226);
not NOT1 (N1228, N678);
nand NAND4 (N1229, N1215, N104, N279, N1159);
buf BUF1 (N1230, N1209);
not NOT1 (N1231, N1230);
xor XOR2 (N1232, N1224, N25);
and AND3 (N1233, N1229, N485, N372);
nor NOR2 (N1234, N1223, N1022);
nand NAND3 (N1235, N1234, N1070, N26);
buf BUF1 (N1236, N1204);
xor XOR2 (N1237, N1199, N73);
nand NAND2 (N1238, N1227, N1010);
buf BUF1 (N1239, N1237);
not NOT1 (N1240, N1238);
not NOT1 (N1241, N1228);
xor XOR2 (N1242, N1240, N1095);
nor NOR2 (N1243, N1231, N487);
nand NAND2 (N1244, N1232, N53);
xor XOR2 (N1245, N1233, N604);
buf BUF1 (N1246, N1242);
nand NAND4 (N1247, N1236, N970, N577, N1211);
xor XOR2 (N1248, N1245, N535);
not NOT1 (N1249, N1247);
buf BUF1 (N1250, N1248);
buf BUF1 (N1251, N1241);
nand NAND2 (N1252, N1225, N81);
or OR3 (N1253, N1239, N742, N1140);
or OR3 (N1254, N1252, N692, N56);
xor XOR2 (N1255, N1235, N1187);
xor XOR2 (N1256, N1255, N264);
not NOT1 (N1257, N1246);
nor NOR4 (N1258, N1256, N369, N1171, N897);
or OR4 (N1259, N1218, N436, N365, N860);
buf BUF1 (N1260, N1254);
nor NOR3 (N1261, N1259, N604, N819);
buf BUF1 (N1262, N1251);
buf BUF1 (N1263, N1253);
or OR2 (N1264, N1258, N283);
buf BUF1 (N1265, N1261);
and AND3 (N1266, N1257, N216, N1171);
nand NAND4 (N1267, N1243, N1204, N411, N726);
and AND3 (N1268, N1260, N829, N698);
xor XOR2 (N1269, N1268, N1095);
and AND4 (N1270, N1244, N85, N299, N445);
not NOT1 (N1271, N1270);
buf BUF1 (N1272, N1250);
not NOT1 (N1273, N1262);
or OR3 (N1274, N1249, N883, N161);
nor NOR4 (N1275, N1272, N574, N1188, N266);
nor NOR4 (N1276, N1264, N1182, N261, N249);
buf BUF1 (N1277, N1269);
buf BUF1 (N1278, N1267);
nor NOR4 (N1279, N1277, N10, N1219, N202);
nand NAND3 (N1280, N1275, N151, N19);
or OR2 (N1281, N1273, N146);
not NOT1 (N1282, N1263);
xor XOR2 (N1283, N1265, N386);
or OR4 (N1284, N1266, N277, N840, N605);
nand NAND2 (N1285, N1283, N107);
nand NAND2 (N1286, N1278, N784);
nand NAND2 (N1287, N1279, N980);
and AND2 (N1288, N1282, N833);
nor NOR4 (N1289, N1271, N824, N1004, N629);
nor NOR4 (N1290, N1281, N1092, N257, N69);
buf BUF1 (N1291, N1286);
and AND2 (N1292, N1288, N934);
or OR2 (N1293, N1289, N163);
xor XOR2 (N1294, N1293, N163);
nand NAND3 (N1295, N1285, N997, N263);
xor XOR2 (N1296, N1287, N1073);
nand NAND4 (N1297, N1295, N1225, N329, N1212);
buf BUF1 (N1298, N1297);
buf BUF1 (N1299, N1280);
nand NAND4 (N1300, N1296, N636, N113, N24);
nor NOR4 (N1301, N1284, N295, N621, N18);
xor XOR2 (N1302, N1276, N408);
nand NAND3 (N1303, N1300, N872, N272);
nand NAND2 (N1304, N1299, N179);
or OR3 (N1305, N1274, N635, N1080);
nor NOR4 (N1306, N1290, N1282, N461, N1214);
nand NAND2 (N1307, N1294, N300);
or OR3 (N1308, N1298, N192, N1140);
nor NOR3 (N1309, N1304, N519, N18);
nand NAND2 (N1310, N1308, N1227);
nand NAND3 (N1311, N1307, N1248, N219);
nand NAND4 (N1312, N1303, N563, N612, N1196);
xor XOR2 (N1313, N1310, N543);
and AND3 (N1314, N1305, N252, N462);
nand NAND3 (N1315, N1309, N44, N612);
nand NAND4 (N1316, N1311, N66, N654, N929);
not NOT1 (N1317, N1291);
xor XOR2 (N1318, N1314, N291);
nor NOR3 (N1319, N1302, N535, N303);
nor NOR2 (N1320, N1318, N312);
nor NOR4 (N1321, N1301, N913, N430, N226);
nand NAND2 (N1322, N1312, N481);
and AND2 (N1323, N1306, N348);
buf BUF1 (N1324, N1320);
nand NAND4 (N1325, N1292, N634, N586, N572);
not NOT1 (N1326, N1315);
nand NAND3 (N1327, N1325, N318, N344);
xor XOR2 (N1328, N1322, N715);
nand NAND3 (N1329, N1328, N684, N214);
or OR2 (N1330, N1327, N506);
nand NAND4 (N1331, N1313, N12, N380, N9);
and AND4 (N1332, N1324, N586, N622, N25);
and AND4 (N1333, N1329, N248, N954, N800);
buf BUF1 (N1334, N1317);
nor NOR4 (N1335, N1333, N659, N174, N29);
and AND3 (N1336, N1331, N823, N372);
and AND2 (N1337, N1330, N551);
not NOT1 (N1338, N1336);
xor XOR2 (N1339, N1323, N1079);
buf BUF1 (N1340, N1316);
buf BUF1 (N1341, N1334);
or OR4 (N1342, N1321, N1183, N780, N232);
not NOT1 (N1343, N1342);
not NOT1 (N1344, N1319);
nor NOR2 (N1345, N1344, N48);
or OR3 (N1346, N1345, N1001, N1039);
buf BUF1 (N1347, N1340);
buf BUF1 (N1348, N1346);
and AND2 (N1349, N1332, N1337);
not NOT1 (N1350, N1055);
or OR4 (N1351, N1326, N1232, N519, N867);
or OR2 (N1352, N1351, N977);
buf BUF1 (N1353, N1343);
and AND3 (N1354, N1348, N450, N758);
nor NOR4 (N1355, N1335, N965, N146, N1288);
nand NAND4 (N1356, N1339, N472, N1187, N1153);
and AND2 (N1357, N1353, N434);
xor XOR2 (N1358, N1354, N742);
or OR2 (N1359, N1347, N352);
not NOT1 (N1360, N1359);
nor NOR4 (N1361, N1358, N119, N662, N1313);
xor XOR2 (N1362, N1352, N512);
and AND4 (N1363, N1362, N427, N117, N487);
and AND2 (N1364, N1341, N65);
nand NAND3 (N1365, N1349, N1168, N849);
nand NAND2 (N1366, N1357, N65);
or OR4 (N1367, N1365, N16, N1265, N288);
nor NOR4 (N1368, N1360, N1062, N627, N1152);
not NOT1 (N1369, N1363);
buf BUF1 (N1370, N1350);
not NOT1 (N1371, N1338);
and AND3 (N1372, N1355, N900, N367);
or OR4 (N1373, N1364, N1053, N552, N570);
and AND4 (N1374, N1372, N1117, N803, N487);
buf BUF1 (N1375, N1369);
nor NOR2 (N1376, N1374, N591);
xor XOR2 (N1377, N1356, N744);
xor XOR2 (N1378, N1370, N386);
buf BUF1 (N1379, N1368);
not NOT1 (N1380, N1377);
and AND2 (N1381, N1361, N236);
nand NAND4 (N1382, N1367, N677, N573, N72);
not NOT1 (N1383, N1373);
and AND2 (N1384, N1375, N1008);
nand NAND3 (N1385, N1383, N1070, N1271);
nand NAND3 (N1386, N1385, N400, N774);
and AND4 (N1387, N1378, N1151, N1198, N905);
and AND3 (N1388, N1384, N1381, N30);
and AND2 (N1389, N41, N995);
and AND4 (N1390, N1380, N311, N35, N361);
and AND3 (N1391, N1387, N907, N879);
or OR4 (N1392, N1371, N1288, N443, N77);
nor NOR2 (N1393, N1389, N99);
and AND3 (N1394, N1390, N506, N1105);
not NOT1 (N1395, N1392);
nand NAND4 (N1396, N1379, N886, N1317, N118);
or OR3 (N1397, N1366, N962, N866);
or OR3 (N1398, N1376, N655, N179);
or OR2 (N1399, N1398, N1233);
nor NOR4 (N1400, N1391, N277, N174, N433);
xor XOR2 (N1401, N1382, N259);
xor XOR2 (N1402, N1397, N472);
xor XOR2 (N1403, N1400, N877);
nand NAND4 (N1404, N1399, N408, N1182, N1181);
not NOT1 (N1405, N1402);
not NOT1 (N1406, N1401);
xor XOR2 (N1407, N1393, N174);
and AND4 (N1408, N1403, N1018, N287, N394);
or OR3 (N1409, N1396, N1279, N196);
and AND4 (N1410, N1404, N1047, N369, N791);
not NOT1 (N1411, N1407);
nor NOR4 (N1412, N1394, N294, N132, N1228);
xor XOR2 (N1413, N1409, N300);
not NOT1 (N1414, N1411);
nor NOR4 (N1415, N1406, N1255, N896, N387);
xor XOR2 (N1416, N1405, N684);
nor NOR3 (N1417, N1413, N457, N1320);
not NOT1 (N1418, N1414);
nor NOR3 (N1419, N1417, N1084, N770);
nand NAND2 (N1420, N1388, N888);
and AND2 (N1421, N1410, N1048);
nor NOR4 (N1422, N1421, N870, N539, N1021);
not NOT1 (N1423, N1395);
and AND4 (N1424, N1412, N1169, N1204, N1350);
not NOT1 (N1425, N1423);
buf BUF1 (N1426, N1424);
xor XOR2 (N1427, N1420, N1087);
buf BUF1 (N1428, N1419);
xor XOR2 (N1429, N1426, N681);
or OR2 (N1430, N1408, N1245);
buf BUF1 (N1431, N1422);
and AND3 (N1432, N1431, N748, N1238);
nor NOR3 (N1433, N1432, N271, N416);
nand NAND2 (N1434, N1433, N242);
xor XOR2 (N1435, N1427, N1125);
not NOT1 (N1436, N1386);
or OR2 (N1437, N1416, N772);
or OR2 (N1438, N1418, N177);
buf BUF1 (N1439, N1429);
or OR4 (N1440, N1430, N360, N405, N29);
nor NOR3 (N1441, N1438, N65, N351);
not NOT1 (N1442, N1428);
nand NAND2 (N1443, N1434, N211);
not NOT1 (N1444, N1437);
or OR2 (N1445, N1442, N413);
not NOT1 (N1446, N1441);
xor XOR2 (N1447, N1439, N1368);
nand NAND3 (N1448, N1445, N763, N919);
not NOT1 (N1449, N1435);
or OR2 (N1450, N1444, N1301);
and AND4 (N1451, N1443, N962, N342, N1136);
and AND3 (N1452, N1425, N1110, N747);
xor XOR2 (N1453, N1415, N1449);
not NOT1 (N1454, N84);
and AND4 (N1455, N1450, N1103, N351, N565);
buf BUF1 (N1456, N1455);
not NOT1 (N1457, N1452);
and AND3 (N1458, N1440, N277, N1167);
or OR3 (N1459, N1446, N808, N1165);
buf BUF1 (N1460, N1458);
and AND2 (N1461, N1459, N727);
and AND4 (N1462, N1436, N317, N1159, N1185);
and AND2 (N1463, N1447, N251);
xor XOR2 (N1464, N1456, N126);
xor XOR2 (N1465, N1460, N139);
buf BUF1 (N1466, N1463);
nor NOR3 (N1467, N1462, N439, N882);
not NOT1 (N1468, N1457);
nor NOR2 (N1469, N1448, N302);
nand NAND3 (N1470, N1467, N1263, N427);
nand NAND3 (N1471, N1470, N934, N1347);
buf BUF1 (N1472, N1453);
xor XOR2 (N1473, N1471, N47);
not NOT1 (N1474, N1466);
xor XOR2 (N1475, N1474, N27);
nor NOR2 (N1476, N1475, N1393);
and AND3 (N1477, N1476, N135, N1053);
nor NOR2 (N1478, N1461, N1069);
or OR2 (N1479, N1477, N1131);
xor XOR2 (N1480, N1478, N1411);
or OR4 (N1481, N1472, N1113, N288, N493);
not NOT1 (N1482, N1454);
nor NOR4 (N1483, N1451, N992, N654, N1466);
nand NAND2 (N1484, N1464, N602);
buf BUF1 (N1485, N1480);
and AND2 (N1486, N1481, N1311);
or OR3 (N1487, N1473, N975, N260);
xor XOR2 (N1488, N1479, N1391);
xor XOR2 (N1489, N1486, N1398);
buf BUF1 (N1490, N1468);
buf BUF1 (N1491, N1488);
xor XOR2 (N1492, N1483, N1430);
or OR3 (N1493, N1487, N1322, N629);
or OR2 (N1494, N1465, N969);
nand NAND3 (N1495, N1489, N681, N421);
buf BUF1 (N1496, N1482);
nand NAND3 (N1497, N1493, N941, N1407);
buf BUF1 (N1498, N1494);
and AND3 (N1499, N1497, N1120, N825);
nand NAND3 (N1500, N1469, N335, N347);
and AND4 (N1501, N1498, N142, N1306, N687);
and AND4 (N1502, N1491, N201, N929, N876);
or OR2 (N1503, N1484, N449);
not NOT1 (N1504, N1502);
xor XOR2 (N1505, N1500, N1483);
not NOT1 (N1506, N1499);
or OR2 (N1507, N1496, N567);
and AND3 (N1508, N1505, N634, N536);
xor XOR2 (N1509, N1507, N1124);
xor XOR2 (N1510, N1509, N906);
or OR2 (N1511, N1504, N241);
nand NAND2 (N1512, N1503, N745);
xor XOR2 (N1513, N1510, N846);
not NOT1 (N1514, N1485);
nor NOR2 (N1515, N1508, N1168);
nand NAND4 (N1516, N1512, N1343, N1288, N1289);
not NOT1 (N1517, N1506);
nand NAND4 (N1518, N1514, N1299, N753, N873);
and AND4 (N1519, N1518, N124, N1232, N1454);
xor XOR2 (N1520, N1515, N1323);
nor NOR2 (N1521, N1520, N1032);
nor NOR3 (N1522, N1513, N740, N119);
not NOT1 (N1523, N1490);
not NOT1 (N1524, N1519);
not NOT1 (N1525, N1495);
or OR3 (N1526, N1511, N1094, N700);
not NOT1 (N1527, N1516);
nor NOR2 (N1528, N1525, N47);
and AND4 (N1529, N1517, N640, N594, N301);
nand NAND4 (N1530, N1492, N1360, N75, N565);
xor XOR2 (N1531, N1524, N956);
nor NOR2 (N1532, N1523, N1418);
or OR3 (N1533, N1529, N209, N1149);
and AND3 (N1534, N1530, N49, N112);
and AND3 (N1535, N1531, N75, N1406);
nor NOR2 (N1536, N1521, N839);
buf BUF1 (N1537, N1501);
not NOT1 (N1538, N1535);
nor NOR4 (N1539, N1528, N332, N916, N853);
or OR3 (N1540, N1537, N266, N1039);
not NOT1 (N1541, N1526);
nor NOR3 (N1542, N1534, N1119, N135);
xor XOR2 (N1543, N1542, N571);
not NOT1 (N1544, N1540);
nor NOR2 (N1545, N1541, N388);
xor XOR2 (N1546, N1539, N1206);
nand NAND3 (N1547, N1538, N1270, N1272);
not NOT1 (N1548, N1543);
and AND4 (N1549, N1546, N1321, N688, N21);
or OR2 (N1550, N1545, N606);
nand NAND3 (N1551, N1549, N553, N1379);
or OR4 (N1552, N1551, N400, N12, N913);
or OR3 (N1553, N1548, N565, N145);
and AND3 (N1554, N1522, N255, N23);
xor XOR2 (N1555, N1536, N1384);
or OR3 (N1556, N1547, N309, N551);
and AND3 (N1557, N1556, N687, N117);
nor NOR3 (N1558, N1527, N1014, N702);
not NOT1 (N1559, N1532);
and AND3 (N1560, N1550, N491, N747);
nand NAND4 (N1561, N1560, N1004, N943, N986);
nor NOR2 (N1562, N1555, N1201);
and AND2 (N1563, N1554, N707);
nand NAND2 (N1564, N1544, N1547);
xor XOR2 (N1565, N1557, N207);
and AND4 (N1566, N1564, N1148, N816, N534);
and AND4 (N1567, N1559, N241, N412, N1075);
nor NOR4 (N1568, N1565, N590, N106, N302);
nand NAND2 (N1569, N1561, N682);
nand NAND2 (N1570, N1558, N1482);
not NOT1 (N1571, N1553);
nor NOR2 (N1572, N1571, N1204);
xor XOR2 (N1573, N1570, N518);
not NOT1 (N1574, N1562);
buf BUF1 (N1575, N1574);
nor NOR4 (N1576, N1566, N599, N946, N839);
nor NOR2 (N1577, N1569, N594);
or OR4 (N1578, N1572, N296, N473, N513);
xor XOR2 (N1579, N1533, N132);
nor NOR3 (N1580, N1579, N206, N919);
xor XOR2 (N1581, N1563, N1249);
or OR2 (N1582, N1575, N208);
and AND2 (N1583, N1552, N145);
xor XOR2 (N1584, N1581, N405);
xor XOR2 (N1585, N1576, N1502);
nor NOR2 (N1586, N1573, N1290);
nand NAND4 (N1587, N1568, N1126, N1545, N594);
buf BUF1 (N1588, N1583);
buf BUF1 (N1589, N1588);
nor NOR2 (N1590, N1586, N1193);
buf BUF1 (N1591, N1589);
buf BUF1 (N1592, N1587);
xor XOR2 (N1593, N1590, N575);
nor NOR2 (N1594, N1578, N643);
or OR4 (N1595, N1580, N1163, N1532, N180);
xor XOR2 (N1596, N1592, N153);
and AND2 (N1597, N1585, N1092);
not NOT1 (N1598, N1593);
nand NAND4 (N1599, N1567, N1424, N871, N1525);
nor NOR4 (N1600, N1582, N1440, N1124, N1263);
and AND3 (N1601, N1599, N1386, N1421);
xor XOR2 (N1602, N1598, N1437);
or OR3 (N1603, N1577, N314, N1214);
nor NOR2 (N1604, N1600, N1140);
xor XOR2 (N1605, N1601, N1064);
nor NOR3 (N1606, N1591, N554, N195);
nor NOR3 (N1607, N1596, N303, N976);
buf BUF1 (N1608, N1604);
and AND2 (N1609, N1607, N652);
or OR3 (N1610, N1602, N1414, N811);
and AND3 (N1611, N1603, N257, N811);
nand NAND3 (N1612, N1610, N1232, N345);
xor XOR2 (N1613, N1584, N95);
nor NOR3 (N1614, N1611, N1423, N351);
nor NOR2 (N1615, N1613, N1242);
nor NOR3 (N1616, N1606, N720, N390);
not NOT1 (N1617, N1594);
buf BUF1 (N1618, N1617);
and AND3 (N1619, N1609, N12, N428);
nor NOR4 (N1620, N1619, N706, N1538, N252);
and AND3 (N1621, N1620, N327, N200);
xor XOR2 (N1622, N1612, N1529);
or OR4 (N1623, N1622, N93, N813, N61);
or OR2 (N1624, N1621, N1086);
nand NAND4 (N1625, N1595, N1285, N900, N1108);
nand NAND2 (N1626, N1618, N650);
nand NAND2 (N1627, N1626, N1624);
or OR4 (N1628, N1589, N1321, N1578, N1532);
not NOT1 (N1629, N1614);
nand NAND4 (N1630, N1605, N1319, N746, N1260);
nand NAND3 (N1631, N1630, N838, N1297);
buf BUF1 (N1632, N1623);
buf BUF1 (N1633, N1631);
nor NOR2 (N1634, N1625, N281);
and AND3 (N1635, N1629, N570, N747);
xor XOR2 (N1636, N1616, N622);
or OR2 (N1637, N1615, N1407);
and AND4 (N1638, N1597, N948, N746, N895);
nor NOR2 (N1639, N1633, N602);
not NOT1 (N1640, N1634);
nand NAND3 (N1641, N1635, N200, N345);
nor NOR3 (N1642, N1636, N943, N372);
and AND4 (N1643, N1632, N1010, N606, N935);
and AND4 (N1644, N1638, N510, N768, N1608);
xor XOR2 (N1645, N1129, N963);
buf BUF1 (N1646, N1641);
buf BUF1 (N1647, N1628);
and AND2 (N1648, N1647, N1629);
and AND2 (N1649, N1640, N1354);
buf BUF1 (N1650, N1645);
xor XOR2 (N1651, N1646, N1055);
xor XOR2 (N1652, N1642, N1226);
not NOT1 (N1653, N1643);
not NOT1 (N1654, N1644);
xor XOR2 (N1655, N1639, N1485);
or OR2 (N1656, N1637, N596);
not NOT1 (N1657, N1656);
and AND2 (N1658, N1648, N1469);
or OR2 (N1659, N1650, N1133);
nor NOR3 (N1660, N1651, N1023, N619);
or OR3 (N1661, N1627, N846, N1637);
nand NAND4 (N1662, N1654, N1547, N79, N1402);
buf BUF1 (N1663, N1653);
buf BUF1 (N1664, N1659);
or OR4 (N1665, N1649, N724, N1148, N1574);
nor NOR3 (N1666, N1660, N200, N1555);
not NOT1 (N1667, N1661);
or OR3 (N1668, N1655, N1430, N307);
and AND3 (N1669, N1666, N548, N1446);
buf BUF1 (N1670, N1663);
xor XOR2 (N1671, N1668, N1059);
nor NOR3 (N1672, N1665, N676, N464);
nand NAND2 (N1673, N1672, N407);
and AND3 (N1674, N1662, N754, N830);
nand NAND3 (N1675, N1664, N475, N821);
xor XOR2 (N1676, N1669, N815);
or OR2 (N1677, N1670, N1184);
buf BUF1 (N1678, N1671);
buf BUF1 (N1679, N1658);
xor XOR2 (N1680, N1657, N392);
not NOT1 (N1681, N1677);
buf BUF1 (N1682, N1652);
buf BUF1 (N1683, N1682);
nand NAND3 (N1684, N1667, N1578, N774);
xor XOR2 (N1685, N1673, N1120);
xor XOR2 (N1686, N1674, N125);
and AND4 (N1687, N1685, N997, N1462, N344);
xor XOR2 (N1688, N1681, N299);
nor NOR2 (N1689, N1684, N300);
nand NAND4 (N1690, N1678, N291, N1373, N1096);
nand NAND4 (N1691, N1687, N664, N50, N662);
buf BUF1 (N1692, N1683);
or OR3 (N1693, N1675, N1628, N26);
xor XOR2 (N1694, N1690, N828);
xor XOR2 (N1695, N1680, N1678);
xor XOR2 (N1696, N1693, N1136);
nand NAND3 (N1697, N1694, N879, N1082);
or OR3 (N1698, N1676, N782, N1362);
buf BUF1 (N1699, N1679);
nor NOR3 (N1700, N1697, N1280, N793);
nand NAND2 (N1701, N1689, N1448);
nor NOR2 (N1702, N1695, N1277);
and AND2 (N1703, N1692, N241);
not NOT1 (N1704, N1686);
or OR3 (N1705, N1691, N625, N1257);
buf BUF1 (N1706, N1699);
or OR3 (N1707, N1704, N1189, N396);
and AND4 (N1708, N1696, N1444, N64, N37);
buf BUF1 (N1709, N1698);
or OR4 (N1710, N1700, N210, N801, N1390);
or OR4 (N1711, N1709, N387, N862, N680);
buf BUF1 (N1712, N1703);
nand NAND2 (N1713, N1711, N695);
and AND3 (N1714, N1713, N93, N575);
not NOT1 (N1715, N1714);
nand NAND4 (N1716, N1702, N31, N950, N249);
not NOT1 (N1717, N1705);
nand NAND3 (N1718, N1708, N482, N620);
nor NOR4 (N1719, N1712, N1518, N1635, N674);
nand NAND4 (N1720, N1715, N1349, N76, N1501);
and AND4 (N1721, N1717, N137, N1476, N1696);
and AND4 (N1722, N1716, N56, N64, N613);
nor NOR2 (N1723, N1688, N10);
or OR3 (N1724, N1701, N341, N1342);
buf BUF1 (N1725, N1724);
nand NAND2 (N1726, N1706, N1127);
nor NOR2 (N1727, N1723, N349);
nand NAND2 (N1728, N1725, N223);
nor NOR3 (N1729, N1718, N460, N1670);
and AND2 (N1730, N1719, N340);
not NOT1 (N1731, N1710);
and AND3 (N1732, N1730, N467, N1398);
xor XOR2 (N1733, N1728, N655);
or OR3 (N1734, N1733, N322, N910);
nor NOR4 (N1735, N1731, N8, N1423, N83);
not NOT1 (N1736, N1721);
nand NAND2 (N1737, N1720, N1662);
and AND3 (N1738, N1735, N883, N1407);
not NOT1 (N1739, N1707);
buf BUF1 (N1740, N1739);
nor NOR3 (N1741, N1726, N740, N272);
or OR2 (N1742, N1722, N118);
xor XOR2 (N1743, N1732, N470);
buf BUF1 (N1744, N1736);
and AND4 (N1745, N1744, N688, N688, N1207);
nor NOR3 (N1746, N1740, N398, N475);
nor NOR4 (N1747, N1746, N613, N659, N432);
not NOT1 (N1748, N1743);
xor XOR2 (N1749, N1727, N143);
xor XOR2 (N1750, N1738, N706);
or OR2 (N1751, N1734, N549);
xor XOR2 (N1752, N1729, N1466);
nand NAND3 (N1753, N1747, N1445, N188);
nand NAND2 (N1754, N1742, N1121);
not NOT1 (N1755, N1745);
and AND2 (N1756, N1741, N912);
or OR4 (N1757, N1755, N685, N385, N1630);
xor XOR2 (N1758, N1757, N515);
nand NAND3 (N1759, N1756, N731, N941);
xor XOR2 (N1760, N1754, N853);
xor XOR2 (N1761, N1759, N713);
buf BUF1 (N1762, N1751);
not NOT1 (N1763, N1750);
xor XOR2 (N1764, N1758, N811);
or OR4 (N1765, N1752, N1470, N991, N374);
nand NAND4 (N1766, N1749, N1096, N454, N1512);
and AND2 (N1767, N1748, N376);
buf BUF1 (N1768, N1737);
not NOT1 (N1769, N1768);
and AND2 (N1770, N1766, N872);
xor XOR2 (N1771, N1760, N1699);
buf BUF1 (N1772, N1764);
or OR4 (N1773, N1770, N1088, N559, N1486);
xor XOR2 (N1774, N1763, N764);
and AND2 (N1775, N1769, N1463);
buf BUF1 (N1776, N1753);
xor XOR2 (N1777, N1761, N448);
and AND3 (N1778, N1776, N338, N787);
nor NOR3 (N1779, N1767, N1680, N1440);
xor XOR2 (N1780, N1772, N622);
xor XOR2 (N1781, N1778, N961);
buf BUF1 (N1782, N1781);
nand NAND3 (N1783, N1774, N1049, N1216);
not NOT1 (N1784, N1780);
nor NOR2 (N1785, N1773, N1194);
and AND4 (N1786, N1775, N42, N1417, N1160);
not NOT1 (N1787, N1785);
nand NAND3 (N1788, N1783, N316, N709);
xor XOR2 (N1789, N1777, N913);
buf BUF1 (N1790, N1784);
or OR3 (N1791, N1789, N17, N409);
nor NOR2 (N1792, N1790, N19);
nor NOR4 (N1793, N1787, N659, N722, N1443);
buf BUF1 (N1794, N1771);
nand NAND3 (N1795, N1788, N1466, N44);
nor NOR4 (N1796, N1782, N593, N606, N1506);
xor XOR2 (N1797, N1791, N651);
nand NAND3 (N1798, N1792, N361, N120);
buf BUF1 (N1799, N1795);
nand NAND2 (N1800, N1765, N1671);
buf BUF1 (N1801, N1800);
nor NOR2 (N1802, N1796, N700);
and AND2 (N1803, N1779, N225);
nor NOR3 (N1804, N1797, N1565, N1263);
nor NOR3 (N1805, N1802, N815, N553);
nor NOR3 (N1806, N1762, N292, N971);
nand NAND3 (N1807, N1805, N1693, N454);
not NOT1 (N1808, N1803);
xor XOR2 (N1809, N1806, N609);
and AND4 (N1810, N1794, N616, N349, N1537);
and AND2 (N1811, N1807, N213);
xor XOR2 (N1812, N1811, N1293);
xor XOR2 (N1813, N1786, N250);
not NOT1 (N1814, N1813);
nor NOR2 (N1815, N1810, N953);
and AND2 (N1816, N1814, N1689);
and AND2 (N1817, N1812, N1056);
not NOT1 (N1818, N1809);
buf BUF1 (N1819, N1799);
and AND3 (N1820, N1801, N122, N1172);
xor XOR2 (N1821, N1820, N741);
xor XOR2 (N1822, N1798, N287);
buf BUF1 (N1823, N1816);
or OR3 (N1824, N1821, N1371, N33);
nand NAND4 (N1825, N1808, N783, N37, N702);
nor NOR2 (N1826, N1819, N1528);
and AND4 (N1827, N1825, N1318, N1793, N384);
or OR4 (N1828, N872, N552, N385, N356);
and AND2 (N1829, N1824, N487);
or OR4 (N1830, N1822, N283, N357, N1105);
and AND3 (N1831, N1818, N1422, N297);
xor XOR2 (N1832, N1829, N656);
or OR4 (N1833, N1817, N1345, N1560, N1568);
or OR4 (N1834, N1826, N1705, N1829, N752);
and AND2 (N1835, N1830, N1231);
nor NOR3 (N1836, N1828, N647, N250);
and AND4 (N1837, N1815, N1701, N1246, N651);
xor XOR2 (N1838, N1804, N664);
not NOT1 (N1839, N1831);
buf BUF1 (N1840, N1838);
buf BUF1 (N1841, N1827);
xor XOR2 (N1842, N1840, N489);
nand NAND3 (N1843, N1833, N1050, N1667);
not NOT1 (N1844, N1841);
nand NAND3 (N1845, N1844, N1402, N226);
nor NOR2 (N1846, N1839, N1788);
not NOT1 (N1847, N1835);
nand NAND2 (N1848, N1836, N67);
nand NAND4 (N1849, N1846, N9, N1224, N1178);
nand NAND4 (N1850, N1823, N439, N1531, N1029);
xor XOR2 (N1851, N1832, N1664);
not NOT1 (N1852, N1848);
or OR3 (N1853, N1850, N288, N1184);
and AND3 (N1854, N1853, N637, N561);
nor NOR2 (N1855, N1843, N271);
not NOT1 (N1856, N1845);
nand NAND4 (N1857, N1851, N126, N1266, N488);
xor XOR2 (N1858, N1842, N641);
nor NOR2 (N1859, N1837, N1126);
nor NOR2 (N1860, N1847, N1149);
xor XOR2 (N1861, N1834, N1082);
nand NAND2 (N1862, N1861, N467);
nand NAND3 (N1863, N1858, N1707, N1251);
and AND2 (N1864, N1857, N1468);
nor NOR4 (N1865, N1856, N853, N1836, N823);
or OR2 (N1866, N1854, N1840);
xor XOR2 (N1867, N1863, N417);
nor NOR4 (N1868, N1866, N1055, N635, N877);
nand NAND4 (N1869, N1852, N785, N1285, N364);
nand NAND2 (N1870, N1865, N1139);
buf BUF1 (N1871, N1868);
nor NOR3 (N1872, N1849, N86, N1442);
xor XOR2 (N1873, N1870, N1260);
nand NAND2 (N1874, N1867, N1080);
not NOT1 (N1875, N1860);
not NOT1 (N1876, N1872);
buf BUF1 (N1877, N1876);
and AND2 (N1878, N1864, N332);
xor XOR2 (N1879, N1874, N1418);
nand NAND2 (N1880, N1875, N448);
nor NOR4 (N1881, N1855, N734, N554, N1539);
xor XOR2 (N1882, N1859, N181);
nor NOR3 (N1883, N1878, N325, N1310);
or OR2 (N1884, N1873, N338);
nor NOR3 (N1885, N1884, N21, N419);
and AND3 (N1886, N1883, N1388, N1539);
nand NAND4 (N1887, N1869, N1528, N1828, N1237);
nand NAND4 (N1888, N1882, N1390, N777, N117);
and AND4 (N1889, N1881, N765, N905, N1654);
or OR2 (N1890, N1889, N91);
nand NAND4 (N1891, N1890, N821, N228, N1535);
or OR3 (N1892, N1891, N721, N1766);
nand NAND4 (N1893, N1877, N426, N416, N944);
buf BUF1 (N1894, N1871);
and AND2 (N1895, N1880, N364);
buf BUF1 (N1896, N1895);
buf BUF1 (N1897, N1892);
xor XOR2 (N1898, N1896, N329);
nor NOR3 (N1899, N1897, N1176, N1204);
or OR4 (N1900, N1893, N794, N11, N973);
xor XOR2 (N1901, N1879, N229);
nor NOR2 (N1902, N1887, N564);
or OR4 (N1903, N1886, N204, N1238, N874);
and AND4 (N1904, N1888, N640, N1534, N742);
buf BUF1 (N1905, N1901);
nand NAND3 (N1906, N1905, N935, N616);
xor XOR2 (N1907, N1894, N453);
or OR2 (N1908, N1902, N1359);
nand NAND3 (N1909, N1885, N1685, N347);
buf BUF1 (N1910, N1862);
and AND4 (N1911, N1910, N439, N1184, N1046);
nand NAND2 (N1912, N1903, N1406);
buf BUF1 (N1913, N1911);
or OR2 (N1914, N1906, N122);
and AND3 (N1915, N1913, N541, N575);
or OR2 (N1916, N1909, N642);
or OR3 (N1917, N1915, N959, N1781);
nand NAND3 (N1918, N1917, N477, N1642);
buf BUF1 (N1919, N1907);
buf BUF1 (N1920, N1908);
not NOT1 (N1921, N1899);
not NOT1 (N1922, N1900);
or OR3 (N1923, N1921, N647, N322);
xor XOR2 (N1924, N1904, N23);
nor NOR4 (N1925, N1914, N114, N544, N916);
or OR3 (N1926, N1923, N841, N985);
nor NOR3 (N1927, N1918, N1074, N1413);
and AND3 (N1928, N1924, N1447, N721);
and AND4 (N1929, N1925, N12, N1081, N1836);
xor XOR2 (N1930, N1927, N633);
and AND2 (N1931, N1916, N638);
nand NAND3 (N1932, N1919, N635, N1670);
xor XOR2 (N1933, N1929, N837);
nor NOR2 (N1934, N1912, N1294);
or OR3 (N1935, N1934, N1405, N1084);
nor NOR4 (N1936, N1928, N289, N168, N983);
and AND2 (N1937, N1935, N715);
not NOT1 (N1938, N1898);
nor NOR4 (N1939, N1932, N699, N104, N1126);
nand NAND3 (N1940, N1936, N1804, N433);
not NOT1 (N1941, N1937);
xor XOR2 (N1942, N1926, N265);
nand NAND2 (N1943, N1941, N513);
or OR2 (N1944, N1940, N1330);
nand NAND4 (N1945, N1922, N1444, N1943, N715);
or OR2 (N1946, N1018, N1757);
buf BUF1 (N1947, N1942);
nor NOR2 (N1948, N1945, N1037);
xor XOR2 (N1949, N1933, N748);
nor NOR4 (N1950, N1931, N991, N764, N649);
xor XOR2 (N1951, N1920, N1342);
or OR4 (N1952, N1948, N1067, N438, N682);
nand NAND4 (N1953, N1947, N266, N794, N1926);
not NOT1 (N1954, N1951);
or OR3 (N1955, N1950, N578, N1699);
not NOT1 (N1956, N1952);
xor XOR2 (N1957, N1946, N1435);
xor XOR2 (N1958, N1939, N1150);
buf BUF1 (N1959, N1938);
not NOT1 (N1960, N1944);
nor NOR3 (N1961, N1949, N1642, N1704);
and AND3 (N1962, N1960, N852, N1176);
nor NOR3 (N1963, N1953, N969, N104);
nor NOR4 (N1964, N1956, N1084, N1077, N414);
buf BUF1 (N1965, N1963);
buf BUF1 (N1966, N1954);
or OR4 (N1967, N1965, N1489, N1158, N270);
xor XOR2 (N1968, N1967, N1832);
buf BUF1 (N1969, N1958);
and AND3 (N1970, N1930, N143, N831);
nor NOR4 (N1971, N1966, N64, N1209, N1794);
or OR4 (N1972, N1955, N1171, N931, N166);
nor NOR3 (N1973, N1972, N107, N39);
xor XOR2 (N1974, N1962, N560);
nor NOR2 (N1975, N1957, N67);
nor NOR3 (N1976, N1975, N1074, N1080);
or OR4 (N1977, N1974, N1468, N1579, N1020);
buf BUF1 (N1978, N1968);
nor NOR3 (N1979, N1977, N625, N1778);
and AND4 (N1980, N1959, N359, N1746, N1818);
buf BUF1 (N1981, N1969);
nor NOR4 (N1982, N1961, N1280, N1692, N939);
or OR4 (N1983, N1982, N1280, N1922, N115);
and AND4 (N1984, N1978, N55, N1211, N1080);
or OR4 (N1985, N1983, N649, N1230, N70);
buf BUF1 (N1986, N1970);
nor NOR4 (N1987, N1976, N1016, N89, N817);
xor XOR2 (N1988, N1979, N1793);
nor NOR4 (N1989, N1988, N1876, N668, N1734);
buf BUF1 (N1990, N1981);
not NOT1 (N1991, N1987);
nand NAND2 (N1992, N1980, N679);
and AND3 (N1993, N1992, N1867, N308);
xor XOR2 (N1994, N1964, N552);
xor XOR2 (N1995, N1973, N250);
not NOT1 (N1996, N1985);
and AND2 (N1997, N1990, N1517);
nor NOR4 (N1998, N1995, N1366, N1806, N777);
xor XOR2 (N1999, N1984, N1652);
xor XOR2 (N2000, N1994, N1813);
not NOT1 (N2001, N1999);
xor XOR2 (N2002, N1998, N1305);
nor NOR2 (N2003, N1993, N363);
or OR2 (N2004, N1971, N433);
nor NOR3 (N2005, N2002, N969, N139);
and AND3 (N2006, N1996, N484, N1916);
buf BUF1 (N2007, N2004);
and AND3 (N2008, N2000, N105, N709);
nand NAND2 (N2009, N2001, N222);
xor XOR2 (N2010, N1989, N1375);
buf BUF1 (N2011, N1986);
nor NOR3 (N2012, N1997, N371, N1399);
xor XOR2 (N2013, N2007, N912);
xor XOR2 (N2014, N2003, N1252);
and AND4 (N2015, N2010, N1546, N1266, N457);
xor XOR2 (N2016, N2011, N1182);
xor XOR2 (N2017, N2009, N211);
nand NAND4 (N2018, N2017, N1151, N1756, N654);
and AND4 (N2019, N2006, N876, N565, N1877);
not NOT1 (N2020, N2019);
xor XOR2 (N2021, N2005, N1738);
or OR2 (N2022, N2018, N314);
or OR3 (N2023, N2008, N991, N298);
or OR4 (N2024, N1991, N1982, N114, N982);
not NOT1 (N2025, N2021);
or OR2 (N2026, N2014, N32);
and AND3 (N2027, N2016, N351, N15);
or OR2 (N2028, N2012, N1553);
buf BUF1 (N2029, N2020);
not NOT1 (N2030, N2023);
nand NAND4 (N2031, N2025, N360, N1867, N1124);
nor NOR4 (N2032, N2029, N618, N1757, N1875);
or OR3 (N2033, N2031, N902, N731);
nor NOR4 (N2034, N2030, N1505, N1296, N913);
or OR3 (N2035, N2015, N1878, N1410);
xor XOR2 (N2036, N2034, N333);
and AND3 (N2037, N2033, N230, N2026);
not NOT1 (N2038, N1905);
or OR4 (N2039, N2038, N112, N1709, N998);
not NOT1 (N2040, N2022);
and AND3 (N2041, N2027, N744, N1426);
not NOT1 (N2042, N2037);
or OR3 (N2043, N2039, N1984, N1251);
or OR3 (N2044, N2042, N698, N435);
not NOT1 (N2045, N2035);
not NOT1 (N2046, N2041);
not NOT1 (N2047, N2024);
nor NOR3 (N2048, N2043, N142, N1934);
or OR4 (N2049, N2028, N1627, N1296, N33);
nand NAND4 (N2050, N2046, N36, N728, N923);
nand NAND3 (N2051, N2040, N1159, N1868);
nand NAND3 (N2052, N2032, N439, N542);
nor NOR4 (N2053, N2036, N1866, N427, N1174);
not NOT1 (N2054, N2050);
not NOT1 (N2055, N2054);
not NOT1 (N2056, N2044);
buf BUF1 (N2057, N2051);
nand NAND4 (N2058, N2057, N2006, N1544, N1619);
buf BUF1 (N2059, N2055);
nor NOR3 (N2060, N2059, N1025, N1917);
or OR4 (N2061, N2047, N6, N1567, N1769);
buf BUF1 (N2062, N2061);
and AND2 (N2063, N2049, N1323);
nor NOR4 (N2064, N2063, N314, N1878, N866);
nor NOR2 (N2065, N2062, N606);
or OR2 (N2066, N2052, N850);
or OR2 (N2067, N2058, N470);
nor NOR3 (N2068, N2066, N1962, N58);
xor XOR2 (N2069, N2048, N1402);
not NOT1 (N2070, N2053);
or OR4 (N2071, N2067, N1371, N1341, N582);
not NOT1 (N2072, N2068);
and AND3 (N2073, N2069, N1279, N1791);
or OR3 (N2074, N2064, N1854, N867);
xor XOR2 (N2075, N2065, N2029);
nand NAND3 (N2076, N2071, N671, N574);
buf BUF1 (N2077, N2072);
nand NAND3 (N2078, N2073, N1660, N1526);
buf BUF1 (N2079, N2060);
nand NAND3 (N2080, N2079, N2048, N1454);
not NOT1 (N2081, N2070);
or OR4 (N2082, N2075, N519, N1189, N282);
nand NAND3 (N2083, N2082, N365, N123);
and AND4 (N2084, N2074, N1051, N1266, N147);
nand NAND3 (N2085, N2076, N734, N1612);
and AND4 (N2086, N2013, N1692, N1060, N569);
nor NOR4 (N2087, N2085, N1595, N1134, N1334);
and AND3 (N2088, N2056, N1457, N1221);
nand NAND2 (N2089, N2088, N846);
or OR3 (N2090, N2081, N1028, N1105);
nor NOR3 (N2091, N2083, N1762, N1455);
nor NOR3 (N2092, N2080, N1563, N1463);
not NOT1 (N2093, N2090);
or OR4 (N2094, N2078, N61, N543, N465);
and AND2 (N2095, N2092, N600);
xor XOR2 (N2096, N2087, N1876);
and AND2 (N2097, N2077, N2079);
xor XOR2 (N2098, N2097, N1938);
or OR3 (N2099, N2045, N1385, N1188);
not NOT1 (N2100, N2086);
buf BUF1 (N2101, N2091);
or OR3 (N2102, N2101, N47, N1685);
not NOT1 (N2103, N2102);
and AND3 (N2104, N2103, N905, N969);
nor NOR3 (N2105, N2089, N215, N2002);
nor NOR4 (N2106, N2105, N88, N106, N1748);
buf BUF1 (N2107, N2096);
nand NAND3 (N2108, N2098, N1633, N207);
buf BUF1 (N2109, N2094);
not NOT1 (N2110, N2104);
nand NAND2 (N2111, N2100, N1172);
buf BUF1 (N2112, N2107);
and AND4 (N2113, N2109, N870, N1720, N702);
not NOT1 (N2114, N2108);
xor XOR2 (N2115, N2114, N440);
and AND3 (N2116, N2095, N1072, N1846);
buf BUF1 (N2117, N2116);
xor XOR2 (N2118, N2117, N1577);
nor NOR3 (N2119, N2112, N880, N833);
buf BUF1 (N2120, N2115);
buf BUF1 (N2121, N2120);
not NOT1 (N2122, N2084);
xor XOR2 (N2123, N2111, N1318);
nand NAND3 (N2124, N2110, N1361, N1647);
buf BUF1 (N2125, N2093);
not NOT1 (N2126, N2118);
or OR3 (N2127, N2121, N1931, N2106);
not NOT1 (N2128, N357);
nor NOR2 (N2129, N2099, N1368);
nand NAND3 (N2130, N2122, N262, N545);
nor NOR3 (N2131, N2128, N1140, N1211);
xor XOR2 (N2132, N2125, N1214);
nor NOR4 (N2133, N2119, N217, N1837, N201);
nor NOR3 (N2134, N2127, N634, N1477);
nand NAND4 (N2135, N2126, N1965, N832, N1068);
nor NOR4 (N2136, N2133, N1783, N627, N141);
xor XOR2 (N2137, N2132, N509);
nand NAND2 (N2138, N2136, N779);
nor NOR4 (N2139, N2138, N107, N656, N2039);
and AND3 (N2140, N2134, N1166, N1852);
nor NOR2 (N2141, N2131, N1426);
buf BUF1 (N2142, N2139);
nor NOR4 (N2143, N2141, N631, N85, N1026);
nand NAND4 (N2144, N2135, N1126, N1638, N196);
or OR3 (N2145, N2140, N765, N1716);
xor XOR2 (N2146, N2124, N1573);
nand NAND2 (N2147, N2113, N2108);
or OR3 (N2148, N2147, N1330, N684);
nor NOR2 (N2149, N2143, N868);
not NOT1 (N2150, N2145);
not NOT1 (N2151, N2146);
xor XOR2 (N2152, N2123, N1889);
and AND4 (N2153, N2144, N1204, N776, N356);
xor XOR2 (N2154, N2151, N2085);
nor NOR4 (N2155, N2137, N407, N1865, N1519);
buf BUF1 (N2156, N2142);
nand NAND4 (N2157, N2154, N673, N509, N107);
nor NOR2 (N2158, N2152, N1779);
xor XOR2 (N2159, N2150, N323);
nor NOR4 (N2160, N2157, N326, N194, N1874);
not NOT1 (N2161, N2160);
not NOT1 (N2162, N2148);
xor XOR2 (N2163, N2129, N1580);
xor XOR2 (N2164, N2162, N1393);
buf BUF1 (N2165, N2163);
or OR2 (N2166, N2164, N308);
not NOT1 (N2167, N2130);
xor XOR2 (N2168, N2167, N660);
xor XOR2 (N2169, N2168, N976);
xor XOR2 (N2170, N2153, N251);
xor XOR2 (N2171, N2161, N994);
and AND4 (N2172, N2169, N193, N1293, N2042);
buf BUF1 (N2173, N2172);
nand NAND3 (N2174, N2165, N2061, N1505);
buf BUF1 (N2175, N2156);
xor XOR2 (N2176, N2174, N1461);
not NOT1 (N2177, N2159);
and AND3 (N2178, N2158, N365, N604);
or OR2 (N2179, N2176, N376);
nor NOR4 (N2180, N2149, N2178, N1863, N2057);
xor XOR2 (N2181, N473, N1885);
not NOT1 (N2182, N2179);
buf BUF1 (N2183, N2173);
or OR4 (N2184, N2170, N669, N1159, N1256);
and AND2 (N2185, N2183, N917);
nand NAND2 (N2186, N2185, N1069);
xor XOR2 (N2187, N2155, N1468);
buf BUF1 (N2188, N2184);
not NOT1 (N2189, N2177);
nor NOR2 (N2190, N2186, N721);
buf BUF1 (N2191, N2190);
nand NAND4 (N2192, N2166, N1525, N705, N460);
and AND4 (N2193, N2191, N855, N355, N606);
not NOT1 (N2194, N2187);
or OR4 (N2195, N2175, N1131, N1468, N1235);
or OR2 (N2196, N2195, N962);
nor NOR2 (N2197, N2196, N241);
nor NOR4 (N2198, N2188, N1629, N1031, N441);
or OR4 (N2199, N2198, N629, N1132, N1711);
nor NOR3 (N2200, N2189, N1748, N1810);
nand NAND3 (N2201, N2171, N677, N1106);
nand NAND3 (N2202, N2197, N577, N1334);
or OR3 (N2203, N2202, N124, N547);
and AND4 (N2204, N2200, N2134, N433, N1887);
and AND4 (N2205, N2181, N1719, N506, N1380);
or OR3 (N2206, N2182, N1847, N1578);
or OR4 (N2207, N2205, N144, N895, N685);
or OR3 (N2208, N2203, N1101, N999);
buf BUF1 (N2209, N2206);
nor NOR3 (N2210, N2180, N1857, N56);
xor XOR2 (N2211, N2209, N2121);
or OR3 (N2212, N2199, N449, N332);
not NOT1 (N2213, N2212);
buf BUF1 (N2214, N2201);
nor NOR4 (N2215, N2204, N2077, N448, N1172);
buf BUF1 (N2216, N2207);
nor NOR2 (N2217, N2194, N1247);
or OR4 (N2218, N2211, N2176, N1235, N1552);
nand NAND3 (N2219, N2214, N1695, N1962);
nand NAND4 (N2220, N2210, N1219, N766, N1850);
not NOT1 (N2221, N2219);
and AND4 (N2222, N2221, N589, N1693, N243);
xor XOR2 (N2223, N2216, N1115);
xor XOR2 (N2224, N2218, N907);
nand NAND2 (N2225, N2192, N2138);
not NOT1 (N2226, N2225);
not NOT1 (N2227, N2213);
xor XOR2 (N2228, N2215, N1139);
and AND4 (N2229, N2208, N571, N1330, N1398);
xor XOR2 (N2230, N2222, N586);
buf BUF1 (N2231, N2224);
nor NOR4 (N2232, N2228, N593, N2131, N1054);
buf BUF1 (N2233, N2227);
nand NAND4 (N2234, N2229, N1181, N140, N284);
not NOT1 (N2235, N2223);
nor NOR3 (N2236, N2220, N996, N1217);
and AND4 (N2237, N2234, N974, N1724, N27);
not NOT1 (N2238, N2237);
nand NAND2 (N2239, N2233, N1268);
nand NAND2 (N2240, N2238, N6);
nand NAND2 (N2241, N2226, N1333);
not NOT1 (N2242, N2241);
buf BUF1 (N2243, N2230);
nand NAND3 (N2244, N2232, N403, N1431);
buf BUF1 (N2245, N2242);
nor NOR2 (N2246, N2235, N132);
nor NOR4 (N2247, N2236, N1409, N635, N2117);
nand NAND3 (N2248, N2244, N1070, N1377);
buf BUF1 (N2249, N2239);
and AND3 (N2250, N2246, N178, N905);
xor XOR2 (N2251, N2217, N2171);
nor NOR3 (N2252, N2231, N1978, N327);
or OR2 (N2253, N2240, N1519);
and AND4 (N2254, N2247, N772, N1448, N294);
nor NOR2 (N2255, N2249, N1254);
or OR4 (N2256, N2253, N1635, N91, N1828);
not NOT1 (N2257, N2193);
xor XOR2 (N2258, N2256, N1876);
buf BUF1 (N2259, N2250);
not NOT1 (N2260, N2255);
buf BUF1 (N2261, N2258);
nor NOR2 (N2262, N2261, N1805);
and AND3 (N2263, N2257, N1276, N579);
not NOT1 (N2264, N2254);
nand NAND3 (N2265, N2251, N1938, N696);
nand NAND3 (N2266, N2262, N471, N429);
nand NAND2 (N2267, N2264, N1374);
and AND2 (N2268, N2260, N2029);
buf BUF1 (N2269, N2267);
nand NAND4 (N2270, N2259, N234, N2150, N2027);
nor NOR3 (N2271, N2243, N1700, N484);
or OR2 (N2272, N2265, N1550);
or OR4 (N2273, N2266, N2237, N429, N1901);
buf BUF1 (N2274, N2273);
xor XOR2 (N2275, N2271, N1757);
not NOT1 (N2276, N2245);
buf BUF1 (N2277, N2276);
and AND3 (N2278, N2248, N1161, N1688);
and AND4 (N2279, N2270, N70, N2055, N1688);
buf BUF1 (N2280, N2277);
not NOT1 (N2281, N2279);
xor XOR2 (N2282, N2263, N273);
not NOT1 (N2283, N2272);
xor XOR2 (N2284, N2280, N2188);
nor NOR3 (N2285, N2275, N1103, N485);
nor NOR4 (N2286, N2285, N2246, N1256, N1517);
or OR2 (N2287, N2252, N1563);
buf BUF1 (N2288, N2281);
nor NOR3 (N2289, N2269, N23, N2266);
xor XOR2 (N2290, N2268, N1768);
and AND3 (N2291, N2284, N520, N2082);
xor XOR2 (N2292, N2289, N858);
buf BUF1 (N2293, N2291);
nor NOR2 (N2294, N2293, N364);
buf BUF1 (N2295, N2290);
nor NOR4 (N2296, N2286, N1870, N1948, N1572);
and AND2 (N2297, N2282, N1824);
and AND2 (N2298, N2287, N453);
or OR3 (N2299, N2283, N1773, N2094);
not NOT1 (N2300, N2278);
or OR4 (N2301, N2298, N670, N1771, N504);
nor NOR2 (N2302, N2301, N775);
not NOT1 (N2303, N2274);
buf BUF1 (N2304, N2299);
xor XOR2 (N2305, N2288, N1100);
buf BUF1 (N2306, N2300);
or OR2 (N2307, N2292, N618);
not NOT1 (N2308, N2294);
not NOT1 (N2309, N2305);
buf BUF1 (N2310, N2307);
nand NAND2 (N2311, N2306, N230);
nor NOR2 (N2312, N2297, N1849);
nand NAND4 (N2313, N2303, N107, N555, N585);
nand NAND4 (N2314, N2311, N2191, N246, N1823);
and AND4 (N2315, N2309, N1646, N757, N1546);
and AND4 (N2316, N2315, N204, N787, N2257);
nor NOR4 (N2317, N2304, N697, N1186, N60);
or OR3 (N2318, N2302, N478, N619);
or OR4 (N2319, N2310, N1942, N657, N104);
or OR4 (N2320, N2318, N623, N1905, N1198);
not NOT1 (N2321, N2312);
or OR4 (N2322, N2296, N110, N1943, N259);
buf BUF1 (N2323, N2308);
nand NAND2 (N2324, N2323, N147);
nand NAND2 (N2325, N2322, N2289);
or OR4 (N2326, N2325, N1994, N1493, N289);
or OR4 (N2327, N2314, N1580, N387, N1299);
nor NOR3 (N2328, N2321, N487, N1928);
nor NOR3 (N2329, N2317, N721, N2258);
nor NOR3 (N2330, N2326, N2296, N754);
xor XOR2 (N2331, N2328, N1977);
nand NAND4 (N2332, N2329, N1524, N776, N1693);
nor NOR4 (N2333, N2319, N2187, N577, N1750);
or OR2 (N2334, N2295, N1567);
xor XOR2 (N2335, N2330, N2105);
nor NOR3 (N2336, N2332, N62, N2077);
xor XOR2 (N2337, N2316, N1019);
or OR4 (N2338, N2324, N696, N502, N1556);
nor NOR2 (N2339, N2327, N1557);
or OR4 (N2340, N2339, N1185, N2198, N2253);
nand NAND3 (N2341, N2337, N910, N1935);
buf BUF1 (N2342, N2335);
and AND3 (N2343, N2320, N250, N2190);
xor XOR2 (N2344, N2333, N1488);
nand NAND4 (N2345, N2313, N1491, N817, N906);
and AND3 (N2346, N2331, N1322, N878);
xor XOR2 (N2347, N2336, N602);
xor XOR2 (N2348, N2343, N576);
nand NAND2 (N2349, N2348, N434);
buf BUF1 (N2350, N2338);
nor NOR4 (N2351, N2346, N2336, N514, N1779);
or OR2 (N2352, N2344, N1256);
nand NAND2 (N2353, N2345, N1189);
nand NAND2 (N2354, N2353, N1744);
buf BUF1 (N2355, N2350);
or OR2 (N2356, N2340, N1035);
or OR3 (N2357, N2342, N495, N1781);
or OR3 (N2358, N2356, N6, N684);
xor XOR2 (N2359, N2357, N891);
nand NAND4 (N2360, N2358, N923, N1562, N991);
or OR4 (N2361, N2354, N121, N1934, N927);
nand NAND4 (N2362, N2360, N2361, N1372, N21);
and AND3 (N2363, N2272, N1746, N1036);
nor NOR2 (N2364, N2362, N996);
nor NOR2 (N2365, N2341, N1557);
nand NAND4 (N2366, N2364, N1634, N1679, N158);
or OR3 (N2367, N2351, N751, N2279);
nand NAND4 (N2368, N2365, N737, N2327, N1023);
xor XOR2 (N2369, N2366, N788);
buf BUF1 (N2370, N2352);
buf BUF1 (N2371, N2369);
nor NOR4 (N2372, N2349, N1297, N1886, N58);
xor XOR2 (N2373, N2363, N1680);
and AND3 (N2374, N2334, N283, N527);
nand NAND4 (N2375, N2374, N1608, N1700, N705);
buf BUF1 (N2376, N2375);
xor XOR2 (N2377, N2367, N1610);
or OR4 (N2378, N2377, N1129, N777, N81);
nor NOR2 (N2379, N2347, N535);
nand NAND4 (N2380, N2355, N238, N1984, N192);
nand NAND3 (N2381, N2368, N1187, N146);
nor NOR2 (N2382, N2373, N2184);
nor NOR3 (N2383, N2370, N1172, N1062);
nand NAND4 (N2384, N2372, N1389, N202, N137);
not NOT1 (N2385, N2381);
and AND3 (N2386, N2384, N1293, N1836);
nand NAND2 (N2387, N2376, N1909);
nor NOR4 (N2388, N2380, N2139, N1974, N1194);
nor NOR2 (N2389, N2371, N1932);
or OR2 (N2390, N2389, N223);
xor XOR2 (N2391, N2359, N1299);
and AND2 (N2392, N2385, N720);
and AND2 (N2393, N2392, N365);
not NOT1 (N2394, N2388);
not NOT1 (N2395, N2391);
nand NAND4 (N2396, N2393, N1510, N979, N1059);
nor NOR3 (N2397, N2379, N2291, N2145);
and AND4 (N2398, N2390, N965, N1990, N2164);
or OR4 (N2399, N2398, N1422, N49, N807);
xor XOR2 (N2400, N2399, N924);
nor NOR3 (N2401, N2383, N737, N951);
and AND3 (N2402, N2387, N1662, N1201);
and AND4 (N2403, N2400, N512, N672, N1433);
buf BUF1 (N2404, N2402);
buf BUF1 (N2405, N2378);
xor XOR2 (N2406, N2401, N1094);
not NOT1 (N2407, N2394);
xor XOR2 (N2408, N2382, N1813);
xor XOR2 (N2409, N2397, N424);
nand NAND4 (N2410, N2395, N332, N1401, N93);
buf BUF1 (N2411, N2386);
nor NOR2 (N2412, N2406, N2180);
nand NAND2 (N2413, N2410, N840);
nor NOR4 (N2414, N2396, N2164, N1306, N766);
and AND3 (N2415, N2403, N2286, N1989);
nand NAND3 (N2416, N2411, N1805, N1459);
nand NAND2 (N2417, N2405, N1438);
nand NAND2 (N2418, N2412, N654);
not NOT1 (N2419, N2408);
xor XOR2 (N2420, N2414, N1048);
and AND4 (N2421, N2409, N2335, N251, N1186);
buf BUF1 (N2422, N2413);
nand NAND2 (N2423, N2419, N1909);
nor NOR4 (N2424, N2418, N392, N182, N488);
not NOT1 (N2425, N2424);
nand NAND2 (N2426, N2425, N433);
or OR3 (N2427, N2415, N889, N800);
xor XOR2 (N2428, N2422, N964);
and AND3 (N2429, N2427, N774, N1562);
and AND2 (N2430, N2429, N182);
nand NAND2 (N2431, N2423, N816);
nor NOR4 (N2432, N2420, N792, N2042, N1817);
nor NOR3 (N2433, N2417, N157, N395);
xor XOR2 (N2434, N2431, N2213);
buf BUF1 (N2435, N2404);
not NOT1 (N2436, N2432);
or OR3 (N2437, N2436, N638, N2092);
and AND4 (N2438, N2430, N2212, N2420, N1902);
not NOT1 (N2439, N2421);
nor NOR4 (N2440, N2407, N815, N2360, N1256);
or OR2 (N2441, N2433, N1640);
not NOT1 (N2442, N2438);
and AND4 (N2443, N2442, N1333, N1028, N2421);
xor XOR2 (N2444, N2435, N1860);
buf BUF1 (N2445, N2443);
nor NOR4 (N2446, N2441, N1253, N569, N1675);
xor XOR2 (N2447, N2437, N1761);
and AND4 (N2448, N2444, N907, N833, N648);
xor XOR2 (N2449, N2428, N2045);
not NOT1 (N2450, N2434);
nand NAND2 (N2451, N2450, N1026);
or OR2 (N2452, N2448, N754);
not NOT1 (N2453, N2449);
and AND3 (N2454, N2426, N813, N2126);
nor NOR2 (N2455, N2447, N508);
xor XOR2 (N2456, N2440, N405);
and AND3 (N2457, N2455, N1642, N776);
not NOT1 (N2458, N2457);
not NOT1 (N2459, N2445);
buf BUF1 (N2460, N2456);
nor NOR2 (N2461, N2439, N307);
nand NAND4 (N2462, N2453, N399, N1299, N2445);
xor XOR2 (N2463, N2452, N2333);
not NOT1 (N2464, N2463);
buf BUF1 (N2465, N2458);
buf BUF1 (N2466, N2451);
buf BUF1 (N2467, N2446);
not NOT1 (N2468, N2459);
and AND4 (N2469, N2462, N2443, N336, N882);
or OR2 (N2470, N2416, N2221);
nand NAND2 (N2471, N2466, N7);
buf BUF1 (N2472, N2469);
xor XOR2 (N2473, N2454, N119);
or OR3 (N2474, N2467, N248, N592);
nor NOR2 (N2475, N2461, N593);
and AND2 (N2476, N2468, N2318);
buf BUF1 (N2477, N2473);
xor XOR2 (N2478, N2464, N924);
and AND4 (N2479, N2470, N1800, N1602, N2193);
xor XOR2 (N2480, N2478, N1782);
or OR2 (N2481, N2472, N528);
buf BUF1 (N2482, N2477);
nand NAND4 (N2483, N2481, N1775, N1408, N1390);
nand NAND3 (N2484, N2476, N2151, N2075);
not NOT1 (N2485, N2471);
or OR2 (N2486, N2475, N2378);
or OR3 (N2487, N2486, N385, N467);
not NOT1 (N2488, N2482);
buf BUF1 (N2489, N2474);
or OR4 (N2490, N2479, N2197, N966, N2210);
or OR4 (N2491, N2480, N2155, N1560, N1537);
nor NOR2 (N2492, N2460, N790);
or OR2 (N2493, N2483, N1765);
xor XOR2 (N2494, N2492, N1925);
and AND2 (N2495, N2490, N289);
not NOT1 (N2496, N2491);
xor XOR2 (N2497, N2488, N813);
not NOT1 (N2498, N2497);
buf BUF1 (N2499, N2493);
or OR4 (N2500, N2498, N1811, N2480, N1523);
nor NOR3 (N2501, N2495, N487, N481);
xor XOR2 (N2502, N2500, N1199);
nor NOR2 (N2503, N2494, N1762);
nand NAND2 (N2504, N2503, N853);
xor XOR2 (N2505, N2484, N1999);
xor XOR2 (N2506, N2499, N1952);
nand NAND2 (N2507, N2465, N2426);
buf BUF1 (N2508, N2496);
or OR2 (N2509, N2507, N2201);
nand NAND4 (N2510, N2508, N2112, N628, N1125);
or OR3 (N2511, N2510, N876, N1462);
nor NOR2 (N2512, N2489, N1082);
nand NAND2 (N2513, N2506, N2252);
nand NAND2 (N2514, N2487, N2189);
xor XOR2 (N2515, N2501, N674);
buf BUF1 (N2516, N2509);
buf BUF1 (N2517, N2511);
and AND3 (N2518, N2513, N101, N395);
and AND4 (N2519, N2485, N1504, N781, N104);
not NOT1 (N2520, N2516);
and AND3 (N2521, N2519, N941, N600);
xor XOR2 (N2522, N2518, N1343);
xor XOR2 (N2523, N2505, N2496);
and AND4 (N2524, N2502, N340, N979, N509);
xor XOR2 (N2525, N2521, N1470);
or OR4 (N2526, N2514, N528, N578, N856);
and AND2 (N2527, N2520, N553);
not NOT1 (N2528, N2524);
or OR4 (N2529, N2525, N1391, N2255, N2297);
nor NOR3 (N2530, N2512, N1546, N125);
or OR4 (N2531, N2523, N821, N1992, N1470);
or OR2 (N2532, N2531, N1141);
xor XOR2 (N2533, N2515, N1070);
buf BUF1 (N2534, N2529);
nor NOR2 (N2535, N2517, N1439);
xor XOR2 (N2536, N2528, N1106);
and AND2 (N2537, N2530, N2042);
xor XOR2 (N2538, N2537, N695);
nor NOR3 (N2539, N2522, N1258, N737);
or OR3 (N2540, N2536, N1919, N140);
not NOT1 (N2541, N2535);
xor XOR2 (N2542, N2534, N296);
nand NAND2 (N2543, N2542, N1167);
nand NAND4 (N2544, N2539, N2474, N1820, N1804);
and AND4 (N2545, N2541, N2241, N789, N622);
nor NOR4 (N2546, N2532, N1946, N1299, N2300);
not NOT1 (N2547, N2538);
xor XOR2 (N2548, N2546, N1359);
nand NAND3 (N2549, N2545, N703, N640);
xor XOR2 (N2550, N2533, N785);
and AND2 (N2551, N2549, N83);
not NOT1 (N2552, N2547);
or OR2 (N2553, N2527, N1090);
not NOT1 (N2554, N2526);
buf BUF1 (N2555, N2540);
nand NAND4 (N2556, N2548, N1201, N63, N1082);
not NOT1 (N2557, N2504);
nand NAND2 (N2558, N2555, N698);
and AND4 (N2559, N2557, N1251, N1772, N341);
nor NOR2 (N2560, N2559, N1183);
or OR3 (N2561, N2544, N1702, N1780);
nor NOR3 (N2562, N2551, N651, N1607);
xor XOR2 (N2563, N2558, N1716);
nor NOR4 (N2564, N2553, N44, N1632, N492);
and AND4 (N2565, N2564, N1763, N388, N2144);
xor XOR2 (N2566, N2552, N1018);
buf BUF1 (N2567, N2561);
xor XOR2 (N2568, N2560, N2452);
buf BUF1 (N2569, N2568);
and AND4 (N2570, N2543, N1003, N202, N886);
xor XOR2 (N2571, N2554, N1901);
not NOT1 (N2572, N2556);
not NOT1 (N2573, N2567);
nor NOR3 (N2574, N2569, N324, N596);
nand NAND3 (N2575, N2566, N458, N396);
and AND3 (N2576, N2563, N1215, N2147);
buf BUF1 (N2577, N2565);
nand NAND3 (N2578, N2570, N2565, N2062);
or OR4 (N2579, N2575, N1199, N809, N1431);
and AND3 (N2580, N2562, N283, N74);
xor XOR2 (N2581, N2573, N888);
nor NOR4 (N2582, N2580, N949, N947, N1518);
or OR2 (N2583, N2581, N1969);
buf BUF1 (N2584, N2572);
or OR4 (N2585, N2584, N1051, N2467, N1757);
nand NAND4 (N2586, N2579, N1505, N1644, N2131);
not NOT1 (N2587, N2571);
or OR3 (N2588, N2582, N386, N1435);
and AND2 (N2589, N2550, N1570);
not NOT1 (N2590, N2588);
xor XOR2 (N2591, N2590, N1121);
nand NAND3 (N2592, N2587, N2169, N747);
not NOT1 (N2593, N2583);
xor XOR2 (N2594, N2586, N1486);
buf BUF1 (N2595, N2578);
and AND4 (N2596, N2585, N2216, N1625, N1337);
nor NOR4 (N2597, N2596, N2197, N2209, N744);
buf BUF1 (N2598, N2595);
not NOT1 (N2599, N2593);
or OR4 (N2600, N2598, N1962, N1686, N703);
nor NOR3 (N2601, N2599, N2143, N695);
or OR4 (N2602, N2600, N1785, N2164, N1562);
not NOT1 (N2603, N2576);
nor NOR2 (N2604, N2597, N1709);
or OR3 (N2605, N2603, N178, N791);
or OR4 (N2606, N2594, N1612, N2024, N1278);
not NOT1 (N2607, N2601);
or OR2 (N2608, N2574, N1576);
or OR4 (N2609, N2606, N2182, N2431, N1956);
not NOT1 (N2610, N2602);
xor XOR2 (N2611, N2605, N2303);
or OR2 (N2612, N2607, N2141);
nand NAND3 (N2613, N2610, N2086, N209);
nand NAND4 (N2614, N2577, N770, N1123, N1801);
and AND3 (N2615, N2591, N622, N378);
or OR2 (N2616, N2612, N195);
nand NAND3 (N2617, N2608, N430, N2531);
and AND3 (N2618, N2613, N968, N820);
buf BUF1 (N2619, N2609);
and AND2 (N2620, N2615, N2334);
buf BUF1 (N2621, N2617);
and AND4 (N2622, N2589, N2106, N126, N1958);
not NOT1 (N2623, N2618);
nor NOR2 (N2624, N2622, N2097);
xor XOR2 (N2625, N2614, N878);
nor NOR3 (N2626, N2624, N261, N668);
not NOT1 (N2627, N2616);
or OR2 (N2628, N2626, N1052);
xor XOR2 (N2629, N2623, N1952);
or OR2 (N2630, N2611, N1628);
nand NAND3 (N2631, N2621, N490, N233);
xor XOR2 (N2632, N2627, N2317);
not NOT1 (N2633, N2604);
nand NAND3 (N2634, N2630, N872, N471);
and AND4 (N2635, N2632, N2124, N1773, N938);
xor XOR2 (N2636, N2592, N1246);
nand NAND4 (N2637, N2629, N876, N182, N2506);
nand NAND2 (N2638, N2635, N6);
and AND2 (N2639, N2634, N861);
nand NAND3 (N2640, N2619, N98, N1938);
xor XOR2 (N2641, N2633, N795);
and AND2 (N2642, N2641, N1433);
nand NAND3 (N2643, N2636, N549, N1721);
xor XOR2 (N2644, N2628, N403);
and AND2 (N2645, N2631, N1291);
xor XOR2 (N2646, N2644, N2546);
and AND4 (N2647, N2642, N396, N2439, N1291);
not NOT1 (N2648, N2647);
or OR2 (N2649, N2645, N436);
xor XOR2 (N2650, N2638, N1884);
or OR3 (N2651, N2625, N2533, N387);
buf BUF1 (N2652, N2620);
not NOT1 (N2653, N2643);
nor NOR3 (N2654, N2652, N1122, N2447);
or OR4 (N2655, N2651, N856, N1483, N1334);
xor XOR2 (N2656, N2655, N1349);
not NOT1 (N2657, N2654);
nor NOR2 (N2658, N2639, N1222);
nor NOR3 (N2659, N2653, N1298, N1300);
nor NOR3 (N2660, N2659, N186, N1490);
buf BUF1 (N2661, N2660);
nand NAND2 (N2662, N2648, N1378);
and AND4 (N2663, N2661, N578, N1498, N1047);
xor XOR2 (N2664, N2637, N1635);
or OR3 (N2665, N2663, N301, N2627);
or OR3 (N2666, N2646, N2514, N1355);
buf BUF1 (N2667, N2664);
not NOT1 (N2668, N2666);
xor XOR2 (N2669, N2657, N1070);
nor NOR2 (N2670, N2668, N478);
xor XOR2 (N2671, N2662, N479);
buf BUF1 (N2672, N2658);
and AND2 (N2673, N2671, N1403);
and AND3 (N2674, N2650, N938, N2043);
or OR3 (N2675, N2674, N1604, N325);
or OR2 (N2676, N2670, N1842);
and AND2 (N2677, N2665, N66);
xor XOR2 (N2678, N2672, N1688);
buf BUF1 (N2679, N2669);
or OR4 (N2680, N2679, N6, N878, N2520);
and AND3 (N2681, N2673, N340, N306);
nand NAND3 (N2682, N2649, N2058, N749);
not NOT1 (N2683, N2675);
not NOT1 (N2684, N2656);
buf BUF1 (N2685, N2677);
nor NOR4 (N2686, N2678, N2023, N1556, N2589);
nand NAND3 (N2687, N2676, N190, N2177);
or OR4 (N2688, N2640, N1610, N979, N2473);
xor XOR2 (N2689, N2683, N2283);
or OR2 (N2690, N2688, N2472);
not NOT1 (N2691, N2687);
not NOT1 (N2692, N2680);
and AND4 (N2693, N2692, N875, N2483, N2373);
and AND4 (N2694, N2681, N2327, N509, N2071);
not NOT1 (N2695, N2684);
buf BUF1 (N2696, N2691);
nand NAND3 (N2697, N2696, N901, N2631);
xor XOR2 (N2698, N2690, N2170);
not NOT1 (N2699, N2693);
not NOT1 (N2700, N2685);
nor NOR3 (N2701, N2695, N2084, N2046);
xor XOR2 (N2702, N2686, N620);
nor NOR2 (N2703, N2689, N135);
or OR4 (N2704, N2697, N642, N2635, N1012);
nor NOR4 (N2705, N2694, N1325, N632, N749);
nand NAND2 (N2706, N2667, N43);
nor NOR2 (N2707, N2702, N1245);
xor XOR2 (N2708, N2703, N2316);
and AND3 (N2709, N2700, N1353, N1188);
nand NAND2 (N2710, N2699, N2111);
or OR2 (N2711, N2706, N2421);
or OR4 (N2712, N2709, N2457, N2367, N2603);
xor XOR2 (N2713, N2682, N1648);
nor NOR2 (N2714, N2698, N1349);
nor NOR2 (N2715, N2704, N2317);
buf BUF1 (N2716, N2705);
buf BUF1 (N2717, N2708);
xor XOR2 (N2718, N2713, N2393);
xor XOR2 (N2719, N2718, N500);
or OR4 (N2720, N2701, N1070, N358, N2185);
and AND2 (N2721, N2707, N2245);
and AND4 (N2722, N2714, N1805, N284, N2287);
and AND3 (N2723, N2717, N863, N376);
nor NOR3 (N2724, N2723, N1738, N681);
buf BUF1 (N2725, N2716);
nor NOR3 (N2726, N2720, N1740, N698);
not NOT1 (N2727, N2722);
buf BUF1 (N2728, N2719);
buf BUF1 (N2729, N2715);
not NOT1 (N2730, N2712);
and AND4 (N2731, N2725, N301, N916, N1271);
and AND4 (N2732, N2729, N843, N760, N2574);
xor XOR2 (N2733, N2732, N1614);
or OR3 (N2734, N2721, N1685, N1922);
nor NOR4 (N2735, N2731, N1592, N233, N1293);
buf BUF1 (N2736, N2734);
nand NAND4 (N2737, N2730, N972, N1802, N420);
nand NAND4 (N2738, N2727, N1574, N356, N997);
buf BUF1 (N2739, N2736);
or OR4 (N2740, N2738, N539, N2509, N1271);
or OR4 (N2741, N2724, N1408, N1366, N669);
or OR4 (N2742, N2710, N406, N1284, N1166);
and AND4 (N2743, N2728, N1975, N996, N2559);
not NOT1 (N2744, N2740);
xor XOR2 (N2745, N2733, N2740);
not NOT1 (N2746, N2726);
nand NAND3 (N2747, N2745, N1265, N1310);
or OR4 (N2748, N2739, N1688, N2616, N1041);
xor XOR2 (N2749, N2743, N2295);
buf BUF1 (N2750, N2711);
xor XOR2 (N2751, N2735, N2685);
xor XOR2 (N2752, N2737, N408);
xor XOR2 (N2753, N2749, N873);
xor XOR2 (N2754, N2746, N1538);
not NOT1 (N2755, N2747);
nor NOR2 (N2756, N2751, N829);
not NOT1 (N2757, N2756);
not NOT1 (N2758, N2754);
buf BUF1 (N2759, N2753);
buf BUF1 (N2760, N2744);
xor XOR2 (N2761, N2750, N1504);
nor NOR2 (N2762, N2748, N905);
or OR2 (N2763, N2760, N1437);
xor XOR2 (N2764, N2742, N920);
and AND4 (N2765, N2752, N2111, N1667, N1182);
not NOT1 (N2766, N2758);
and AND3 (N2767, N2765, N2464, N2563);
nand NAND2 (N2768, N2761, N689);
not NOT1 (N2769, N2762);
not NOT1 (N2770, N2768);
xor XOR2 (N2771, N2741, N239);
and AND2 (N2772, N2766, N1112);
or OR4 (N2773, N2769, N248, N2009, N989);
or OR4 (N2774, N2772, N762, N1368, N2370);
or OR2 (N2775, N2763, N1783);
or OR4 (N2776, N2755, N2554, N2501, N1252);
xor XOR2 (N2777, N2759, N1137);
nand NAND2 (N2778, N2776, N935);
or OR3 (N2779, N2770, N1614, N1066);
xor XOR2 (N2780, N2775, N737);
nand NAND3 (N2781, N2767, N405, N2017);
nor NOR2 (N2782, N2777, N373);
not NOT1 (N2783, N2757);
nand NAND4 (N2784, N2782, N1531, N2330, N2041);
xor XOR2 (N2785, N2764, N251);
nand NAND3 (N2786, N2774, N1231, N1220);
and AND4 (N2787, N2781, N921, N1046, N2675);
or OR3 (N2788, N2784, N1300, N2689);
not NOT1 (N2789, N2771);
xor XOR2 (N2790, N2780, N918);
not NOT1 (N2791, N2788);
not NOT1 (N2792, N2778);
nand NAND4 (N2793, N2786, N2285, N1258, N2339);
nand NAND2 (N2794, N2783, N2617);
nor NOR4 (N2795, N2773, N1929, N69, N2441);
not NOT1 (N2796, N2794);
not NOT1 (N2797, N2779);
buf BUF1 (N2798, N2785);
buf BUF1 (N2799, N2791);
and AND2 (N2800, N2796, N2781);
or OR4 (N2801, N2799, N2072, N897, N294);
or OR2 (N2802, N2798, N2541);
or OR4 (N2803, N2793, N1168, N1183, N882);
buf BUF1 (N2804, N2802);
nor NOR4 (N2805, N2800, N2366, N1285, N72);
or OR3 (N2806, N2789, N1421, N1436);
nand NAND4 (N2807, N2801, N2790, N212, N628);
buf BUF1 (N2808, N2734);
and AND3 (N2809, N2806, N288, N590);
nand NAND2 (N2810, N2797, N141);
not NOT1 (N2811, N2795);
nand NAND2 (N2812, N2803, N2628);
nand NAND4 (N2813, N2792, N461, N2644, N959);
not NOT1 (N2814, N2808);
xor XOR2 (N2815, N2787, N2462);
or OR2 (N2816, N2804, N1213);
nor NOR2 (N2817, N2815, N560);
not NOT1 (N2818, N2813);
or OR4 (N2819, N2805, N414, N2429, N2541);
not NOT1 (N2820, N2807);
nor NOR3 (N2821, N2819, N986, N2170);
nand NAND4 (N2822, N2812, N1678, N740, N2295);
and AND2 (N2823, N2818, N1083);
xor XOR2 (N2824, N2809, N1095);
xor XOR2 (N2825, N2811, N1295);
not NOT1 (N2826, N2816);
not NOT1 (N2827, N2814);
xor XOR2 (N2828, N2822, N1582);
nand NAND3 (N2829, N2823, N2003, N473);
buf BUF1 (N2830, N2810);
not NOT1 (N2831, N2826);
nand NAND3 (N2832, N2830, N2366, N182);
or OR3 (N2833, N2820, N2689, N824);
not NOT1 (N2834, N2829);
and AND2 (N2835, N2833, N2019);
nand NAND4 (N2836, N2828, N21, N2591, N1317);
or OR3 (N2837, N2821, N658, N1185);
and AND4 (N2838, N2834, N1278, N2792, N2747);
xor XOR2 (N2839, N2831, N1835);
nor NOR3 (N2840, N2817, N2318, N2818);
nand NAND3 (N2841, N2839, N899, N2090);
buf BUF1 (N2842, N2836);
xor XOR2 (N2843, N2832, N2283);
buf BUF1 (N2844, N2837);
nor NOR3 (N2845, N2840, N1404, N672);
xor XOR2 (N2846, N2843, N1397);
buf BUF1 (N2847, N2845);
or OR3 (N2848, N2842, N2795, N2370);
and AND4 (N2849, N2847, N648, N423, N1987);
and AND4 (N2850, N2838, N680, N456, N644);
buf BUF1 (N2851, N2850);
xor XOR2 (N2852, N2824, N2628);
not NOT1 (N2853, N2835);
not NOT1 (N2854, N2848);
or OR2 (N2855, N2844, N2700);
or OR4 (N2856, N2851, N626, N230, N798);
nor NOR2 (N2857, N2846, N1358);
nand NAND2 (N2858, N2825, N2158);
or OR4 (N2859, N2849, N944, N2237, N760);
xor XOR2 (N2860, N2859, N153);
nor NOR2 (N2861, N2856, N429);
xor XOR2 (N2862, N2852, N1971);
or OR3 (N2863, N2853, N203, N1464);
not NOT1 (N2864, N2861);
nor NOR4 (N2865, N2827, N2227, N725, N1317);
not NOT1 (N2866, N2863);
nand NAND3 (N2867, N2864, N1061, N1490);
buf BUF1 (N2868, N2855);
buf BUF1 (N2869, N2866);
not NOT1 (N2870, N2854);
nand NAND2 (N2871, N2862, N431);
not NOT1 (N2872, N2871);
nor NOR4 (N2873, N2858, N1915, N1044, N372);
not NOT1 (N2874, N2870);
or OR3 (N2875, N2841, N1568, N872);
and AND4 (N2876, N2873, N624, N2293, N2560);
xor XOR2 (N2877, N2875, N2743);
buf BUF1 (N2878, N2872);
or OR3 (N2879, N2869, N2719, N1714);
buf BUF1 (N2880, N2868);
or OR4 (N2881, N2874, N182, N2708, N2451);
nand NAND4 (N2882, N2879, N387, N2054, N1669);
not NOT1 (N2883, N2867);
xor XOR2 (N2884, N2857, N2596);
nand NAND4 (N2885, N2882, N1154, N2493, N2199);
not NOT1 (N2886, N2880);
buf BUF1 (N2887, N2860);
xor XOR2 (N2888, N2883, N1429);
xor XOR2 (N2889, N2884, N1826);
and AND2 (N2890, N2865, N1698);
not NOT1 (N2891, N2877);
xor XOR2 (N2892, N2881, N2554);
or OR3 (N2893, N2891, N1674, N1858);
nand NAND4 (N2894, N2890, N2691, N843, N1969);
nor NOR2 (N2895, N2885, N1612);
and AND2 (N2896, N2888, N160);
or OR2 (N2897, N2878, N1329);
not NOT1 (N2898, N2892);
nor NOR4 (N2899, N2876, N2090, N2497, N468);
nor NOR4 (N2900, N2899, N1160, N1530, N2772);
not NOT1 (N2901, N2898);
xor XOR2 (N2902, N2889, N878);
xor XOR2 (N2903, N2897, N321);
and AND3 (N2904, N2896, N1429, N2083);
nand NAND4 (N2905, N2886, N2809, N1959, N1341);
or OR3 (N2906, N2900, N2194, N1085);
or OR2 (N2907, N2895, N401);
xor XOR2 (N2908, N2904, N2157);
or OR2 (N2909, N2894, N2689);
buf BUF1 (N2910, N2909);
not NOT1 (N2911, N2901);
or OR3 (N2912, N2905, N2133, N2058);
or OR3 (N2913, N2911, N2029, N294);
xor XOR2 (N2914, N2913, N2142);
xor XOR2 (N2915, N2914, N974);
or OR2 (N2916, N2903, N24);
not NOT1 (N2917, N2910);
buf BUF1 (N2918, N2915);
nand NAND3 (N2919, N2912, N1011, N968);
or OR3 (N2920, N2917, N152, N2810);
or OR2 (N2921, N2919, N2607);
not NOT1 (N2922, N2902);
nand NAND2 (N2923, N2907, N2548);
xor XOR2 (N2924, N2906, N686);
nand NAND3 (N2925, N2908, N432, N1851);
and AND3 (N2926, N2921, N370, N2315);
or OR3 (N2927, N2887, N2424, N514);
nand NAND3 (N2928, N2923, N2813, N1331);
xor XOR2 (N2929, N2920, N97);
nand NAND3 (N2930, N2922, N1206, N359);
not NOT1 (N2931, N2930);
and AND3 (N2932, N2929, N1241, N2241);
xor XOR2 (N2933, N2927, N616);
nand NAND4 (N2934, N2925, N2879, N2175, N1983);
or OR4 (N2935, N2928, N2648, N1645, N2093);
nor NOR2 (N2936, N2918, N2890);
nor NOR4 (N2937, N2916, N614, N1801, N2442);
and AND2 (N2938, N2932, N2861);
not NOT1 (N2939, N2938);
nor NOR2 (N2940, N2931, N104);
xor XOR2 (N2941, N2937, N2464);
xor XOR2 (N2942, N2941, N1776);
and AND2 (N2943, N2939, N1105);
buf BUF1 (N2944, N2893);
buf BUF1 (N2945, N2933);
nand NAND2 (N2946, N2934, N484);
xor XOR2 (N2947, N2924, N1698);
and AND3 (N2948, N2940, N1573, N1829);
nor NOR4 (N2949, N2936, N655, N2018, N1031);
and AND4 (N2950, N2944, N639, N1305, N2690);
nand NAND3 (N2951, N2949, N1188, N257);
and AND2 (N2952, N2951, N838);
or OR3 (N2953, N2942, N2539, N1492);
nor NOR3 (N2954, N2935, N1335, N2419);
nor NOR4 (N2955, N2954, N853, N2101, N2180);
and AND2 (N2956, N2950, N2451);
not NOT1 (N2957, N2952);
nand NAND4 (N2958, N2955, N1160, N1773, N1479);
and AND4 (N2959, N2948, N2132, N953, N859);
nor NOR2 (N2960, N2943, N1571);
and AND2 (N2961, N2946, N2005);
or OR3 (N2962, N2961, N1276, N840);
buf BUF1 (N2963, N2947);
nand NAND2 (N2964, N2959, N2910);
buf BUF1 (N2965, N2958);
nor NOR3 (N2966, N2965, N167, N915);
buf BUF1 (N2967, N2966);
or OR4 (N2968, N2960, N915, N2205, N2176);
xor XOR2 (N2969, N2953, N56);
and AND3 (N2970, N2957, N1847, N407);
not NOT1 (N2971, N2963);
not NOT1 (N2972, N2971);
not NOT1 (N2973, N2968);
and AND2 (N2974, N2926, N122);
nor NOR2 (N2975, N2964, N2944);
or OR4 (N2976, N2974, N1164, N1345, N1831);
not NOT1 (N2977, N2945);
and AND3 (N2978, N2970, N2079, N2087);
not NOT1 (N2979, N2975);
nor NOR2 (N2980, N2967, N1862);
buf BUF1 (N2981, N2976);
buf BUF1 (N2982, N2980);
and AND4 (N2983, N2977, N1704, N1064, N2361);
nand NAND2 (N2984, N2978, N2710);
nor NOR3 (N2985, N2981, N2783, N2001);
buf BUF1 (N2986, N2956);
buf BUF1 (N2987, N2982);
and AND2 (N2988, N2962, N2119);
and AND4 (N2989, N2973, N16, N2562, N528);
xor XOR2 (N2990, N2979, N2167);
or OR3 (N2991, N2987, N1044, N1883);
nand NAND3 (N2992, N2990, N2737, N79);
nand NAND2 (N2993, N2969, N2433);
and AND2 (N2994, N2985, N2379);
buf BUF1 (N2995, N2992);
buf BUF1 (N2996, N2986);
xor XOR2 (N2997, N2984, N2792);
nor NOR2 (N2998, N2996, N1422);
xor XOR2 (N2999, N2991, N2498);
nand NAND3 (N3000, N2999, N1654, N591);
nand NAND4 (N3001, N3000, N1746, N346, N1364);
xor XOR2 (N3002, N2998, N75);
nor NOR4 (N3003, N2989, N2232, N2153, N52);
not NOT1 (N3004, N3002);
and AND2 (N3005, N2993, N758);
nand NAND4 (N3006, N3004, N334, N2928, N618);
nor NOR3 (N3007, N2988, N2754, N1922);
or OR4 (N3008, N2983, N2505, N2637, N1639);
buf BUF1 (N3009, N2995);
buf BUF1 (N3010, N3009);
xor XOR2 (N3011, N2972, N1616);
nor NOR3 (N3012, N2994, N2065, N1635);
or OR2 (N3013, N3008, N2484);
nand NAND2 (N3014, N3003, N2723);
or OR4 (N3015, N3010, N2394, N2372, N2797);
nand NAND4 (N3016, N3001, N846, N1547, N2959);
buf BUF1 (N3017, N3007);
xor XOR2 (N3018, N3006, N854);
nand NAND2 (N3019, N3013, N2320);
xor XOR2 (N3020, N3016, N1871);
nand NAND3 (N3021, N3019, N1301, N2644);
nand NAND2 (N3022, N3015, N2987);
buf BUF1 (N3023, N3018);
nand NAND3 (N3024, N3017, N1441, N945);
nor NOR4 (N3025, N3021, N2345, N2099, N629);
and AND4 (N3026, N3014, N2752, N932, N128);
nor NOR3 (N3027, N3005, N2143, N2361);
and AND2 (N3028, N3024, N1753);
nand NAND4 (N3029, N3020, N1944, N2676, N2906);
and AND2 (N3030, N3011, N1278);
buf BUF1 (N3031, N2997);
or OR3 (N3032, N3028, N1076, N514);
or OR3 (N3033, N3030, N2299, N2965);
and AND3 (N3034, N3026, N844, N696);
xor XOR2 (N3035, N3025, N343);
or OR2 (N3036, N3033, N142);
or OR3 (N3037, N3012, N2664, N2190);
or OR3 (N3038, N3023, N2161, N59);
or OR4 (N3039, N3037, N126, N1162, N405);
nand NAND4 (N3040, N3027, N278, N826, N2658);
nor NOR2 (N3041, N3031, N2261);
not NOT1 (N3042, N3035);
buf BUF1 (N3043, N3032);
or OR2 (N3044, N3022, N1267);
nor NOR2 (N3045, N3040, N2288);
xor XOR2 (N3046, N3029, N2167);
not NOT1 (N3047, N3045);
xor XOR2 (N3048, N3042, N1757);
xor XOR2 (N3049, N3041, N1760);
nand NAND4 (N3050, N3039, N1661, N272, N1527);
and AND2 (N3051, N3036, N1879);
nand NAND3 (N3052, N3043, N2628, N2357);
nor NOR4 (N3053, N3049, N1755, N50, N55);
nand NAND4 (N3054, N3048, N2455, N2254, N2709);
nor NOR4 (N3055, N3053, N1007, N101, N1722);
nor NOR4 (N3056, N3047, N420, N2670, N11);
not NOT1 (N3057, N3038);
or OR3 (N3058, N3051, N1579, N2152);
buf BUF1 (N3059, N3057);
nor NOR2 (N3060, N3050, N1595);
not NOT1 (N3061, N3055);
nor NOR4 (N3062, N3054, N228, N2921, N2202);
or OR3 (N3063, N3062, N2373, N2056);
nor NOR3 (N3064, N3046, N1796, N744);
not NOT1 (N3065, N3034);
xor XOR2 (N3066, N3058, N1232);
not NOT1 (N3067, N3056);
nand NAND3 (N3068, N3066, N631, N1364);
buf BUF1 (N3069, N3068);
nor NOR2 (N3070, N3059, N2048);
xor XOR2 (N3071, N3060, N2929);
xor XOR2 (N3072, N3061, N438);
nand NAND4 (N3073, N3063, N551, N1097, N2948);
nand NAND3 (N3074, N3070, N2717, N2128);
or OR4 (N3075, N3073, N2321, N1499, N2783);
not NOT1 (N3076, N3075);
nor NOR4 (N3077, N3067, N2671, N2313, N2219);
not NOT1 (N3078, N3071);
nor NOR2 (N3079, N3044, N1568);
or OR3 (N3080, N3072, N1349, N984);
nand NAND3 (N3081, N3077, N301, N1468);
or OR3 (N3082, N3078, N1095, N2648);
not NOT1 (N3083, N3081);
buf BUF1 (N3084, N3079);
or OR2 (N3085, N3064, N1695);
not NOT1 (N3086, N3069);
buf BUF1 (N3087, N3084);
not NOT1 (N3088, N3083);
not NOT1 (N3089, N3085);
nand NAND3 (N3090, N3076, N2078, N2240);
nand NAND2 (N3091, N3052, N1594);
not NOT1 (N3092, N3080);
nor NOR4 (N3093, N3089, N1523, N1774, N1590);
not NOT1 (N3094, N3082);
and AND3 (N3095, N3090, N601, N1843);
nor NOR3 (N3096, N3094, N1149, N173);
nor NOR2 (N3097, N3092, N166);
nand NAND3 (N3098, N3065, N2416, N1439);
or OR3 (N3099, N3074, N1871, N11);
buf BUF1 (N3100, N3096);
not NOT1 (N3101, N3086);
not NOT1 (N3102, N3091);
nor NOR4 (N3103, N3101, N2409, N2119, N214);
and AND4 (N3104, N3099, N788, N1129, N581);
nand NAND3 (N3105, N3097, N351, N370);
buf BUF1 (N3106, N3103);
or OR3 (N3107, N3093, N1312, N1916);
xor XOR2 (N3108, N3087, N322);
not NOT1 (N3109, N3105);
and AND4 (N3110, N3109, N2629, N902, N2671);
nand NAND4 (N3111, N3107, N903, N2203, N2027);
or OR2 (N3112, N3095, N2661);
nand NAND2 (N3113, N3106, N1883);
xor XOR2 (N3114, N3112, N3018);
buf BUF1 (N3115, N3100);
not NOT1 (N3116, N3113);
nor NOR2 (N3117, N3098, N427);
nor NOR2 (N3118, N3088, N1419);
buf BUF1 (N3119, N3102);
nand NAND4 (N3120, N3108, N2801, N1317, N2766);
or OR2 (N3121, N3116, N331);
not NOT1 (N3122, N3114);
nor NOR4 (N3123, N3122, N806, N971, N1960);
not NOT1 (N3124, N3115);
nor NOR3 (N3125, N3118, N1718, N280);
nand NAND3 (N3126, N3104, N476, N2694);
and AND3 (N3127, N3121, N1763, N1049);
and AND3 (N3128, N3119, N565, N596);
nand NAND4 (N3129, N3111, N1698, N272, N2302);
nand NAND3 (N3130, N3124, N284, N700);
nor NOR3 (N3131, N3129, N728, N3036);
nor NOR2 (N3132, N3117, N1098);
or OR4 (N3133, N3127, N517, N2339, N1764);
buf BUF1 (N3134, N3120);
xor XOR2 (N3135, N3131, N3045);
buf BUF1 (N3136, N3135);
nand NAND2 (N3137, N3133, N2785);
not NOT1 (N3138, N3126);
nor NOR2 (N3139, N3125, N3093);
xor XOR2 (N3140, N3137, N1714);
nor NOR3 (N3141, N3132, N1041, N310);
and AND4 (N3142, N3123, N821, N1501, N413);
buf BUF1 (N3143, N3130);
xor XOR2 (N3144, N3140, N2347);
nand NAND2 (N3145, N3134, N1628);
buf BUF1 (N3146, N3142);
or OR4 (N3147, N3141, N3012, N2430, N348);
xor XOR2 (N3148, N3144, N2530);
nand NAND4 (N3149, N3143, N750, N889, N1353);
nor NOR3 (N3150, N3128, N290, N1458);
xor XOR2 (N3151, N3110, N402);
and AND4 (N3152, N3146, N373, N2809, N623);
xor XOR2 (N3153, N3151, N141);
or OR4 (N3154, N3149, N2361, N826, N52);
buf BUF1 (N3155, N3139);
nor NOR4 (N3156, N3154, N2079, N588, N292);
not NOT1 (N3157, N3155);
and AND2 (N3158, N3157, N1465);
nor NOR2 (N3159, N3158, N392);
not NOT1 (N3160, N3159);
xor XOR2 (N3161, N3138, N577);
xor XOR2 (N3162, N3152, N625);
not NOT1 (N3163, N3145);
xor XOR2 (N3164, N3162, N6);
or OR2 (N3165, N3156, N2319);
not NOT1 (N3166, N3136);
and AND2 (N3167, N3163, N2607);
not NOT1 (N3168, N3148);
buf BUF1 (N3169, N3164);
or OR2 (N3170, N3150, N388);
not NOT1 (N3171, N3166);
and AND3 (N3172, N3167, N598, N1004);
nand NAND2 (N3173, N3161, N2504);
and AND2 (N3174, N3171, N2927);
and AND2 (N3175, N3165, N1716);
nor NOR4 (N3176, N3160, N1537, N1063, N2768);
nor NOR3 (N3177, N3147, N321, N3002);
nor NOR2 (N3178, N3176, N3001);
or OR2 (N3179, N3173, N2164);
not NOT1 (N3180, N3179);
nand NAND2 (N3181, N3168, N2522);
not NOT1 (N3182, N3172);
nor NOR3 (N3183, N3178, N2519, N2055);
not NOT1 (N3184, N3174);
xor XOR2 (N3185, N3181, N2761);
and AND2 (N3186, N3177, N1187);
or OR2 (N3187, N3182, N2481);
or OR2 (N3188, N3170, N2785);
or OR2 (N3189, N3187, N754);
xor XOR2 (N3190, N3189, N1711);
buf BUF1 (N3191, N3185);
nor NOR2 (N3192, N3190, N1423);
or OR3 (N3193, N3191, N2846, N722);
nand NAND2 (N3194, N3193, N2420);
nand NAND2 (N3195, N3184, N1894);
nand NAND3 (N3196, N3188, N3042, N1042);
xor XOR2 (N3197, N3186, N2247);
or OR2 (N3198, N3180, N3140);
buf BUF1 (N3199, N3195);
and AND4 (N3200, N3183, N2132, N2184, N2716);
buf BUF1 (N3201, N3196);
not NOT1 (N3202, N3198);
buf BUF1 (N3203, N3200);
and AND3 (N3204, N3201, N473, N1199);
buf BUF1 (N3205, N3204);
not NOT1 (N3206, N3153);
and AND3 (N3207, N3206, N780, N96);
nor NOR2 (N3208, N3175, N2592);
or OR4 (N3209, N3197, N2476, N1597, N903);
xor XOR2 (N3210, N3169, N2863);
not NOT1 (N3211, N3199);
nor NOR4 (N3212, N3208, N2701, N2596, N939);
xor XOR2 (N3213, N3205, N97);
or OR4 (N3214, N3213, N1128, N1463, N2260);
buf BUF1 (N3215, N3203);
buf BUF1 (N3216, N3194);
nor NOR2 (N3217, N3216, N344);
or OR3 (N3218, N3210, N2610, N1281);
xor XOR2 (N3219, N3218, N2663);
not NOT1 (N3220, N3192);
buf BUF1 (N3221, N3209);
and AND4 (N3222, N3217, N681, N2378, N421);
xor XOR2 (N3223, N3215, N678);
and AND2 (N3224, N3222, N628);
nor NOR4 (N3225, N3224, N1666, N1558, N3087);
xor XOR2 (N3226, N3219, N967);
xor XOR2 (N3227, N3226, N2476);
xor XOR2 (N3228, N3227, N1873);
buf BUF1 (N3229, N3202);
and AND2 (N3230, N3211, N2003);
xor XOR2 (N3231, N3214, N1633);
nand NAND3 (N3232, N3220, N533, N770);
xor XOR2 (N3233, N3231, N1937);
and AND2 (N3234, N3229, N2401);
nand NAND4 (N3235, N3228, N2830, N1891, N2204);
and AND4 (N3236, N3221, N1519, N856, N1376);
and AND4 (N3237, N3223, N1042, N2601, N3170);
buf BUF1 (N3238, N3236);
nand NAND3 (N3239, N3232, N349, N2612);
and AND4 (N3240, N3239, N1524, N1112, N129);
nand NAND2 (N3241, N3212, N1123);
and AND3 (N3242, N3235, N112, N1922);
not NOT1 (N3243, N3238);
or OR4 (N3244, N3225, N2247, N322, N1430);
buf BUF1 (N3245, N3243);
xor XOR2 (N3246, N3245, N2272);
nand NAND2 (N3247, N3233, N700);
nor NOR2 (N3248, N3207, N1623);
buf BUF1 (N3249, N3240);
nor NOR4 (N3250, N3246, N1739, N1582, N2658);
buf BUF1 (N3251, N3249);
nand NAND3 (N3252, N3234, N2497, N1549);
not NOT1 (N3253, N3237);
xor XOR2 (N3254, N3247, N2832);
nor NOR3 (N3255, N3241, N1482, N1588);
not NOT1 (N3256, N3251);
xor XOR2 (N3257, N3250, N371);
or OR2 (N3258, N3242, N1127);
or OR4 (N3259, N3248, N2276, N2258, N1581);
nand NAND2 (N3260, N3230, N2584);
buf BUF1 (N3261, N3254);
not NOT1 (N3262, N3253);
nor NOR2 (N3263, N3261, N1855);
buf BUF1 (N3264, N3252);
and AND2 (N3265, N3244, N296);
not NOT1 (N3266, N3256);
nor NOR4 (N3267, N3262, N2533, N758, N2327);
nand NAND4 (N3268, N3258, N2193, N2705, N1884);
or OR2 (N3269, N3267, N2193);
or OR3 (N3270, N3265, N3145, N98);
buf BUF1 (N3271, N3257);
nand NAND4 (N3272, N3255, N2636, N2819, N2015);
buf BUF1 (N3273, N3270);
nor NOR2 (N3274, N3260, N2935);
not NOT1 (N3275, N3269);
xor XOR2 (N3276, N3263, N51);
or OR2 (N3277, N3264, N1835);
or OR2 (N3278, N3271, N1328);
nor NOR3 (N3279, N3278, N1025, N3004);
nand NAND3 (N3280, N3273, N319, N632);
buf BUF1 (N3281, N3280);
nand NAND4 (N3282, N3268, N2179, N1084, N217);
xor XOR2 (N3283, N3276, N2833);
xor XOR2 (N3284, N3274, N1038);
buf BUF1 (N3285, N3281);
nor NOR2 (N3286, N3259, N1872);
nand NAND3 (N3287, N3279, N1930, N2932);
buf BUF1 (N3288, N3287);
xor XOR2 (N3289, N3283, N1660);
and AND2 (N3290, N3289, N2268);
xor XOR2 (N3291, N3288, N1711);
nor NOR2 (N3292, N3282, N3103);
xor XOR2 (N3293, N3286, N3165);
not NOT1 (N3294, N3266);
nand NAND3 (N3295, N3284, N412, N2694);
nor NOR3 (N3296, N3290, N1208, N504);
and AND4 (N3297, N3285, N214, N1038, N1472);
nand NAND3 (N3298, N3275, N2684, N1043);
nor NOR2 (N3299, N3291, N1676);
or OR2 (N3300, N3277, N612);
and AND2 (N3301, N3296, N2595);
not NOT1 (N3302, N3295);
nand NAND4 (N3303, N3300, N2139, N2611, N1243);
xor XOR2 (N3304, N3297, N1706);
buf BUF1 (N3305, N3303);
and AND3 (N3306, N3292, N759, N2229);
xor XOR2 (N3307, N3304, N2132);
nand NAND2 (N3308, N3305, N1322);
xor XOR2 (N3309, N3306, N607);
and AND2 (N3310, N3301, N183);
not NOT1 (N3311, N3310);
or OR4 (N3312, N3298, N2965, N1675, N1693);
nor NOR3 (N3313, N3293, N1658, N1083);
not NOT1 (N3314, N3311);
nor NOR3 (N3315, N3309, N2592, N912);
xor XOR2 (N3316, N3294, N1794);
nor NOR4 (N3317, N3299, N3150, N542, N306);
and AND2 (N3318, N3314, N2154);
or OR4 (N3319, N3272, N43, N3030, N3015);
nand NAND4 (N3320, N3312, N1461, N1225, N3022);
xor XOR2 (N3321, N3320, N1781);
buf BUF1 (N3322, N3313);
buf BUF1 (N3323, N3315);
or OR2 (N3324, N3302, N604);
nor NOR4 (N3325, N3307, N246, N476, N3245);
or OR2 (N3326, N3319, N2322);
or OR3 (N3327, N3324, N3197, N2263);
xor XOR2 (N3328, N3318, N1059);
nor NOR3 (N3329, N3317, N1866, N664);
or OR4 (N3330, N3316, N360, N1036, N2290);
xor XOR2 (N3331, N3321, N2035);
and AND2 (N3332, N3330, N1308);
buf BUF1 (N3333, N3308);
or OR2 (N3334, N3327, N2017);
buf BUF1 (N3335, N3322);
xor XOR2 (N3336, N3331, N2602);
not NOT1 (N3337, N3335);
buf BUF1 (N3338, N3328);
nand NAND3 (N3339, N3325, N1609, N3287);
or OR4 (N3340, N3332, N1586, N1616, N1148);
xor XOR2 (N3341, N3323, N2229);
nor NOR2 (N3342, N3337, N27);
and AND4 (N3343, N3334, N2162, N818, N2921);
nand NAND4 (N3344, N3336, N2319, N1897, N728);
or OR2 (N3345, N3339, N1314);
xor XOR2 (N3346, N3341, N1839);
nor NOR3 (N3347, N3345, N1036, N199);
or OR2 (N3348, N3343, N2508);
xor XOR2 (N3349, N3344, N1828);
nor NOR3 (N3350, N3348, N3017, N1860);
xor XOR2 (N3351, N3333, N2782);
nand NAND3 (N3352, N3338, N3075, N2732);
xor XOR2 (N3353, N3342, N3258);
and AND4 (N3354, N3326, N1741, N3272, N2550);
not NOT1 (N3355, N3354);
xor XOR2 (N3356, N3329, N692);
buf BUF1 (N3357, N3351);
or OR4 (N3358, N3356, N1307, N236, N658);
and AND3 (N3359, N3352, N2691, N1182);
or OR3 (N3360, N3355, N1044, N1487);
nor NOR3 (N3361, N3360, N3084, N2199);
xor XOR2 (N3362, N3349, N886);
nor NOR2 (N3363, N3347, N1901);
not NOT1 (N3364, N3340);
or OR2 (N3365, N3364, N2678);
and AND2 (N3366, N3357, N572);
and AND2 (N3367, N3359, N2671);
xor XOR2 (N3368, N3346, N1566);
and AND4 (N3369, N3358, N543, N555, N64);
or OR3 (N3370, N3366, N1256, N1439);
not NOT1 (N3371, N3368);
not NOT1 (N3372, N3363);
nand NAND3 (N3373, N3370, N2744, N3048);
and AND4 (N3374, N3372, N1305, N1338, N654);
nand NAND3 (N3375, N3367, N1995, N1036);
buf BUF1 (N3376, N3374);
and AND4 (N3377, N3365, N2483, N2198, N2040);
nor NOR2 (N3378, N3350, N2082);
xor XOR2 (N3379, N3353, N1177);
and AND2 (N3380, N3377, N3033);
xor XOR2 (N3381, N3376, N3082);
or OR3 (N3382, N3381, N2223, N2280);
buf BUF1 (N3383, N3379);
or OR4 (N3384, N3380, N2958, N2070, N3258);
and AND2 (N3385, N3373, N465);
buf BUF1 (N3386, N3384);
nor NOR4 (N3387, N3383, N2760, N2311, N316);
xor XOR2 (N3388, N3371, N1976);
nor NOR3 (N3389, N3387, N2963, N1324);
not NOT1 (N3390, N3389);
not NOT1 (N3391, N3361);
buf BUF1 (N3392, N3390);
and AND3 (N3393, N3391, N1888, N330);
nand NAND2 (N3394, N3388, N1289);
nor NOR2 (N3395, N3382, N3135);
and AND3 (N3396, N3393, N535, N2638);
nand NAND3 (N3397, N3395, N111, N2600);
xor XOR2 (N3398, N3386, N601);
nand NAND3 (N3399, N3378, N2823, N2390);
and AND3 (N3400, N3385, N2392, N2097);
and AND3 (N3401, N3362, N286, N2560);
not NOT1 (N3402, N3392);
not NOT1 (N3403, N3398);
and AND3 (N3404, N3399, N1709, N2512);
nand NAND2 (N3405, N3401, N2243);
or OR2 (N3406, N3396, N2246);
or OR4 (N3407, N3400, N2659, N375, N380);
or OR4 (N3408, N3403, N815, N2546, N1991);
xor XOR2 (N3409, N3406, N1035);
not NOT1 (N3410, N3404);
buf BUF1 (N3411, N3407);
not NOT1 (N3412, N3405);
or OR4 (N3413, N3369, N742, N794, N2381);
buf BUF1 (N3414, N3413);
nor NOR4 (N3415, N3411, N684, N2556, N1666);
nand NAND2 (N3416, N3397, N1824);
not NOT1 (N3417, N3412);
nand NAND2 (N3418, N3408, N3316);
or OR3 (N3419, N3394, N2338, N13);
not NOT1 (N3420, N3410);
buf BUF1 (N3421, N3409);
and AND3 (N3422, N3415, N3051, N276);
or OR3 (N3423, N3414, N998, N1527);
or OR2 (N3424, N3418, N1299);
buf BUF1 (N3425, N3422);
nor NOR4 (N3426, N3419, N2805, N3404, N1396);
not NOT1 (N3427, N3375);
xor XOR2 (N3428, N3402, N3217);
xor XOR2 (N3429, N3427, N1579);
not NOT1 (N3430, N3421);
buf BUF1 (N3431, N3423);
buf BUF1 (N3432, N3424);
not NOT1 (N3433, N3428);
xor XOR2 (N3434, N3431, N2352);
buf BUF1 (N3435, N3434);
xor XOR2 (N3436, N3430, N2845);
not NOT1 (N3437, N3417);
nor NOR3 (N3438, N3425, N471, N804);
not NOT1 (N3439, N3436);
and AND4 (N3440, N3429, N2097, N1916, N1233);
xor XOR2 (N3441, N3433, N1445);
or OR3 (N3442, N3420, N2206, N174);
not NOT1 (N3443, N3442);
nor NOR2 (N3444, N3426, N1853);
not NOT1 (N3445, N3432);
buf BUF1 (N3446, N3440);
nor NOR3 (N3447, N3435, N523, N1788);
nand NAND2 (N3448, N3445, N1649);
or OR4 (N3449, N3443, N3281, N2601, N1861);
xor XOR2 (N3450, N3444, N2821);
or OR4 (N3451, N3437, N2055, N687, N2142);
nand NAND4 (N3452, N3441, N1355, N1215, N435);
xor XOR2 (N3453, N3447, N2504);
buf BUF1 (N3454, N3438);
nor NOR3 (N3455, N3448, N574, N1167);
buf BUF1 (N3456, N3452);
and AND3 (N3457, N3450, N2862, N1304);
not NOT1 (N3458, N3446);
or OR2 (N3459, N3458, N784);
nand NAND3 (N3460, N3454, N1914, N2050);
nor NOR4 (N3461, N3460, N3217, N1013, N2415);
nor NOR2 (N3462, N3457, N26);
nor NOR3 (N3463, N3461, N2889, N2067);
and AND3 (N3464, N3462, N2380, N3141);
buf BUF1 (N3465, N3459);
nand NAND4 (N3466, N3455, N3040, N1551, N2340);
and AND4 (N3467, N3463, N1941, N3064, N3036);
or OR2 (N3468, N3453, N1204);
not NOT1 (N3469, N3465);
buf BUF1 (N3470, N3467);
nand NAND4 (N3471, N3449, N2170, N1872, N2430);
not NOT1 (N3472, N3451);
nand NAND2 (N3473, N3468, N88);
buf BUF1 (N3474, N3469);
and AND2 (N3475, N3474, N244);
buf BUF1 (N3476, N3466);
buf BUF1 (N3477, N3439);
and AND2 (N3478, N3472, N613);
not NOT1 (N3479, N3475);
xor XOR2 (N3480, N3416, N529);
and AND4 (N3481, N3470, N545, N2722, N694);
xor XOR2 (N3482, N3478, N2834);
not NOT1 (N3483, N3479);
and AND2 (N3484, N3483, N2353);
nand NAND4 (N3485, N3464, N3296, N2552, N798);
or OR3 (N3486, N3471, N741, N419);
nor NOR4 (N3487, N3481, N1742, N2303, N2308);
nand NAND4 (N3488, N3480, N1433, N2517, N3027);
buf BUF1 (N3489, N3485);
buf BUF1 (N3490, N3476);
nor NOR2 (N3491, N3473, N3119);
xor XOR2 (N3492, N3482, N1625);
xor XOR2 (N3493, N3486, N3397);
and AND4 (N3494, N3489, N3128, N991, N2406);
nor NOR3 (N3495, N3488, N69, N942);
xor XOR2 (N3496, N3490, N3009);
or OR3 (N3497, N3487, N209, N1209);
and AND2 (N3498, N3493, N3283);
buf BUF1 (N3499, N3456);
not NOT1 (N3500, N3499);
not NOT1 (N3501, N3500);
not NOT1 (N3502, N3496);
nor NOR3 (N3503, N3477, N2957, N1419);
nand NAND4 (N3504, N3494, N3450, N3332, N1586);
or OR4 (N3505, N3492, N3209, N2827, N2676);
xor XOR2 (N3506, N3505, N542);
and AND3 (N3507, N3502, N1839, N2205);
nor NOR2 (N3508, N3498, N1622);
not NOT1 (N3509, N3507);
and AND3 (N3510, N3491, N2270, N3326);
xor XOR2 (N3511, N3509, N969);
buf BUF1 (N3512, N3484);
buf BUF1 (N3513, N3503);
nor NOR4 (N3514, N3497, N3466, N2232, N1645);
and AND2 (N3515, N3508, N224);
xor XOR2 (N3516, N3511, N575);
and AND2 (N3517, N3504, N430);
or OR4 (N3518, N3516, N667, N2908, N3090);
or OR2 (N3519, N3518, N2045);
not NOT1 (N3520, N3512);
buf BUF1 (N3521, N3519);
and AND2 (N3522, N3521, N460);
xor XOR2 (N3523, N3501, N730);
nand NAND3 (N3524, N3495, N1166, N2859);
xor XOR2 (N3525, N3524, N1996);
buf BUF1 (N3526, N3515);
nand NAND4 (N3527, N3526, N1621, N647, N2488);
not NOT1 (N3528, N3506);
not NOT1 (N3529, N3523);
nor NOR3 (N3530, N3525, N2930, N3256);
nand NAND2 (N3531, N3530, N946);
or OR4 (N3532, N3513, N3345, N1962, N2365);
nand NAND2 (N3533, N3532, N2278);
nor NOR3 (N3534, N3527, N963, N116);
nand NAND3 (N3535, N3522, N2225, N1154);
nor NOR3 (N3536, N3533, N3406, N171);
and AND4 (N3537, N3514, N1996, N2486, N2211);
xor XOR2 (N3538, N3531, N1261);
and AND2 (N3539, N3517, N462);
xor XOR2 (N3540, N3535, N2357);
or OR4 (N3541, N3529, N1057, N1073, N2075);
and AND4 (N3542, N3538, N3218, N3031, N105);
buf BUF1 (N3543, N3541);
buf BUF1 (N3544, N3510);
nand NAND2 (N3545, N3539, N3365);
and AND3 (N3546, N3540, N2220, N228);
or OR4 (N3547, N3542, N3158, N362, N2053);
and AND2 (N3548, N3537, N2900);
or OR4 (N3549, N3520, N3246, N3378, N2463);
buf BUF1 (N3550, N3545);
xor XOR2 (N3551, N3547, N1284);
not NOT1 (N3552, N3550);
nor NOR4 (N3553, N3548, N865, N2446, N1137);
xor XOR2 (N3554, N3536, N3001);
or OR4 (N3555, N3551, N1981, N3436, N2566);
not NOT1 (N3556, N3552);
buf BUF1 (N3557, N3528);
nand NAND2 (N3558, N3554, N2811);
nand NAND2 (N3559, N3557, N268);
not NOT1 (N3560, N3549);
not NOT1 (N3561, N3534);
not NOT1 (N3562, N3559);
nor NOR2 (N3563, N3561, N1690);
not NOT1 (N3564, N3544);
xor XOR2 (N3565, N3546, N2454);
or OR4 (N3566, N3543, N625, N993, N3109);
nor NOR2 (N3567, N3565, N2469);
and AND4 (N3568, N3562, N1334, N2314, N912);
buf BUF1 (N3569, N3567);
not NOT1 (N3570, N3563);
and AND3 (N3571, N3555, N1872, N2673);
nor NOR2 (N3572, N3553, N834);
and AND4 (N3573, N3572, N3263, N1195, N3307);
nor NOR2 (N3574, N3570, N2459);
or OR3 (N3575, N3564, N1946, N2246);
or OR4 (N3576, N3568, N668, N540, N33);
and AND2 (N3577, N3569, N2204);
not NOT1 (N3578, N3577);
or OR3 (N3579, N3574, N2034, N381);
buf BUF1 (N3580, N3566);
xor XOR2 (N3581, N3560, N336);
buf BUF1 (N3582, N3573);
and AND4 (N3583, N3576, N2682, N1717, N2225);
nand NAND3 (N3584, N3578, N1160, N2875);
or OR2 (N3585, N3580, N3147);
xor XOR2 (N3586, N3558, N1969);
nor NOR4 (N3587, N3575, N12, N1831, N188);
not NOT1 (N3588, N3556);
and AND3 (N3589, N3587, N3243, N1680);
nor NOR4 (N3590, N3581, N1774, N1296, N1514);
nor NOR4 (N3591, N3579, N411, N2529, N3406);
xor XOR2 (N3592, N3586, N578);
nand NAND3 (N3593, N3588, N329, N1751);
not NOT1 (N3594, N3571);
xor XOR2 (N3595, N3584, N3276);
buf BUF1 (N3596, N3585);
not NOT1 (N3597, N3582);
buf BUF1 (N3598, N3597);
and AND4 (N3599, N3593, N2548, N703, N1071);
or OR2 (N3600, N3598, N1941);
xor XOR2 (N3601, N3592, N522);
or OR3 (N3602, N3596, N2687, N490);
xor XOR2 (N3603, N3600, N373);
xor XOR2 (N3604, N3602, N2265);
nand NAND4 (N3605, N3603, N1699, N1443, N2942);
nand NAND3 (N3606, N3604, N1002, N2570);
xor XOR2 (N3607, N3601, N3460);
or OR4 (N3608, N3590, N2556, N3497, N3059);
and AND2 (N3609, N3595, N132);
nand NAND4 (N3610, N3594, N677, N2198, N2050);
and AND3 (N3611, N3599, N3499, N1938);
xor XOR2 (N3612, N3583, N529);
xor XOR2 (N3613, N3609, N951);
nand NAND4 (N3614, N3605, N2904, N715, N867);
not NOT1 (N3615, N3614);
xor XOR2 (N3616, N3612, N1940);
and AND3 (N3617, N3589, N196, N2102);
not NOT1 (N3618, N3608);
nor NOR3 (N3619, N3616, N464, N1332);
and AND3 (N3620, N3613, N3078, N2555);
nor NOR3 (N3621, N3618, N1471, N2562);
buf BUF1 (N3622, N3619);
nand NAND3 (N3623, N3622, N692, N1975);
nor NOR3 (N3624, N3623, N731, N3312);
and AND4 (N3625, N3610, N1355, N3040, N2574);
xor XOR2 (N3626, N3617, N1327);
nor NOR4 (N3627, N3606, N3394, N522, N349);
not NOT1 (N3628, N3611);
nor NOR2 (N3629, N3615, N3295);
nor NOR4 (N3630, N3624, N3323, N639, N1558);
buf BUF1 (N3631, N3626);
nor NOR2 (N3632, N3631, N1375);
or OR4 (N3633, N3627, N2957, N532, N883);
xor XOR2 (N3634, N3591, N3304);
and AND4 (N3635, N3633, N1787, N74, N393);
and AND3 (N3636, N3607, N1064, N2713);
nand NAND3 (N3637, N3625, N2084, N2502);
nand NAND3 (N3638, N3632, N1173, N1517);
or OR3 (N3639, N3634, N1604, N1429);
nor NOR4 (N3640, N3635, N2834, N555, N1331);
xor XOR2 (N3641, N3620, N314);
and AND4 (N3642, N3630, N1278, N946, N3526);
nand NAND4 (N3643, N3636, N185, N2748, N1847);
xor XOR2 (N3644, N3629, N249);
or OR4 (N3645, N3641, N2552, N2061, N2277);
xor XOR2 (N3646, N3637, N2787);
and AND3 (N3647, N3640, N2684, N2119);
or OR2 (N3648, N3639, N1730);
and AND4 (N3649, N3628, N234, N440, N3155);
nand NAND3 (N3650, N3646, N1115, N1416);
nor NOR3 (N3651, N3650, N2226, N2361);
and AND3 (N3652, N3651, N2646, N2021);
nand NAND4 (N3653, N3649, N478, N3298, N3439);
or OR4 (N3654, N3645, N984, N2902, N1367);
or OR4 (N3655, N3642, N1695, N2425, N1184);
nor NOR4 (N3656, N3654, N260, N3433, N1835);
xor XOR2 (N3657, N3652, N1668);
and AND4 (N3658, N3648, N3451, N812, N1666);
and AND3 (N3659, N3653, N771, N1477);
buf BUF1 (N3660, N3638);
buf BUF1 (N3661, N3621);
nand NAND4 (N3662, N3657, N3239, N58, N660);
or OR4 (N3663, N3655, N1768, N2323, N183);
or OR4 (N3664, N3661, N3647, N1692, N3470);
xor XOR2 (N3665, N2928, N2463);
nand NAND2 (N3666, N3660, N2417);
nor NOR4 (N3667, N3659, N3243, N293, N3001);
buf BUF1 (N3668, N3662);
buf BUF1 (N3669, N3668);
buf BUF1 (N3670, N3644);
nor NOR4 (N3671, N3663, N3376, N2214, N314);
not NOT1 (N3672, N3669);
and AND3 (N3673, N3666, N996, N1119);
or OR3 (N3674, N3665, N2046, N32);
and AND2 (N3675, N3674, N329);
and AND4 (N3676, N3656, N25, N2151, N218);
or OR3 (N3677, N3676, N2422, N2241);
nor NOR4 (N3678, N3675, N3499, N777, N783);
buf BUF1 (N3679, N3670);
and AND2 (N3680, N3664, N966);
not NOT1 (N3681, N3658);
buf BUF1 (N3682, N3672);
and AND3 (N3683, N3671, N2875, N3606);
buf BUF1 (N3684, N3681);
buf BUF1 (N3685, N3673);
buf BUF1 (N3686, N3682);
and AND3 (N3687, N3684, N1118, N2167);
xor XOR2 (N3688, N3683, N3216);
xor XOR2 (N3689, N3678, N2928);
nor NOR4 (N3690, N3689, N3145, N2918, N2160);
xor XOR2 (N3691, N3687, N2242);
not NOT1 (N3692, N3643);
nor NOR2 (N3693, N3685, N2033);
not NOT1 (N3694, N3677);
or OR3 (N3695, N3686, N2712, N783);
nor NOR3 (N3696, N3695, N1023, N435);
xor XOR2 (N3697, N3679, N2935);
nand NAND4 (N3698, N3694, N1769, N3220, N1536);
xor XOR2 (N3699, N3696, N3316);
not NOT1 (N3700, N3688);
nor NOR2 (N3701, N3693, N3004);
not NOT1 (N3702, N3690);
nor NOR3 (N3703, N3699, N1276, N554);
buf BUF1 (N3704, N3700);
buf BUF1 (N3705, N3697);
or OR2 (N3706, N3698, N644);
xor XOR2 (N3707, N3705, N2802);
xor XOR2 (N3708, N3702, N578);
buf BUF1 (N3709, N3680);
xor XOR2 (N3710, N3709, N433);
not NOT1 (N3711, N3708);
or OR4 (N3712, N3710, N408, N2916, N2134);
not NOT1 (N3713, N3667);
xor XOR2 (N3714, N3703, N634);
xor XOR2 (N3715, N3692, N1464);
nand NAND3 (N3716, N3713, N1041, N1781);
xor XOR2 (N3717, N3715, N1577);
nor NOR3 (N3718, N3704, N1427, N2972);
or OR3 (N3719, N3691, N2293, N3201);
and AND2 (N3720, N3716, N532);
not NOT1 (N3721, N3719);
buf BUF1 (N3722, N3718);
nand NAND2 (N3723, N3722, N2045);
or OR3 (N3724, N3707, N2603, N673);
buf BUF1 (N3725, N3712);
and AND4 (N3726, N3711, N2555, N439, N1775);
nor NOR4 (N3727, N3720, N2892, N2358, N2448);
nor NOR4 (N3728, N3706, N3582, N1063, N7);
and AND4 (N3729, N3723, N1740, N1302, N3164);
xor XOR2 (N3730, N3726, N680);
not NOT1 (N3731, N3727);
xor XOR2 (N3732, N3721, N1447);
and AND2 (N3733, N3714, N2124);
and AND4 (N3734, N3724, N2232, N427, N2087);
not NOT1 (N3735, N3732);
and AND3 (N3736, N3725, N3060, N2267);
or OR2 (N3737, N3728, N83);
and AND3 (N3738, N3731, N3409, N2634);
not NOT1 (N3739, N3730);
nor NOR4 (N3740, N3739, N1002, N2142, N2056);
or OR3 (N3741, N3729, N2968, N2138);
nor NOR3 (N3742, N3735, N1366, N442);
buf BUF1 (N3743, N3740);
not NOT1 (N3744, N3741);
buf BUF1 (N3745, N3743);
xor XOR2 (N3746, N3738, N145);
xor XOR2 (N3747, N3733, N842);
nand NAND2 (N3748, N3745, N133);
xor XOR2 (N3749, N3747, N1152);
and AND4 (N3750, N3701, N1917, N3238, N1251);
not NOT1 (N3751, N3742);
buf BUF1 (N3752, N3717);
and AND3 (N3753, N3749, N2038, N2816);
and AND3 (N3754, N3737, N598, N1920);
nor NOR2 (N3755, N3754, N3209);
nor NOR2 (N3756, N3744, N404);
xor XOR2 (N3757, N3750, N634);
xor XOR2 (N3758, N3757, N1886);
or OR2 (N3759, N3746, N1388);
xor XOR2 (N3760, N3751, N2385);
nand NAND2 (N3761, N3755, N394);
nor NOR4 (N3762, N3759, N2161, N3680, N1664);
or OR2 (N3763, N3762, N1540);
buf BUF1 (N3764, N3734);
and AND3 (N3765, N3753, N2448, N2873);
buf BUF1 (N3766, N3756);
not NOT1 (N3767, N3766);
and AND4 (N3768, N3760, N3035, N72, N2110);
not NOT1 (N3769, N3764);
xor XOR2 (N3770, N3768, N3647);
buf BUF1 (N3771, N3765);
buf BUF1 (N3772, N3736);
and AND2 (N3773, N3758, N394);
or OR2 (N3774, N3748, N873);
nor NOR3 (N3775, N3770, N2079, N1466);
and AND2 (N3776, N3773, N3010);
buf BUF1 (N3777, N3774);
or OR4 (N3778, N3771, N2157, N2718, N2269);
not NOT1 (N3779, N3775);
or OR4 (N3780, N3763, N2252, N2014, N882);
not NOT1 (N3781, N3752);
nor NOR4 (N3782, N3767, N997, N3731, N39);
buf BUF1 (N3783, N3780);
nand NAND2 (N3784, N3779, N3712);
xor XOR2 (N3785, N3761, N2304);
nor NOR3 (N3786, N3785, N1481, N3554);
nand NAND4 (N3787, N3776, N3523, N3547, N943);
xor XOR2 (N3788, N3781, N1560);
nor NOR2 (N3789, N3772, N666);
not NOT1 (N3790, N3783);
and AND4 (N3791, N3789, N3447, N1563, N1119);
xor XOR2 (N3792, N3782, N2506);
buf BUF1 (N3793, N3787);
and AND2 (N3794, N3778, N2734);
xor XOR2 (N3795, N3769, N820);
buf BUF1 (N3796, N3791);
or OR3 (N3797, N3795, N2942, N1387);
buf BUF1 (N3798, N3797);
or OR3 (N3799, N3793, N104, N2035);
or OR3 (N3800, N3794, N2160, N1474);
buf BUF1 (N3801, N3800);
or OR4 (N3802, N3801, N3681, N1299, N916);
or OR2 (N3803, N3784, N862);
buf BUF1 (N3804, N3790);
and AND2 (N3805, N3792, N2027);
nand NAND3 (N3806, N3803, N3433, N2242);
not NOT1 (N3807, N3796);
or OR4 (N3808, N3807, N3397, N2455, N3386);
or OR3 (N3809, N3804, N1136, N3603);
buf BUF1 (N3810, N3809);
nand NAND3 (N3811, N3798, N666, N3623);
buf BUF1 (N3812, N3786);
nand NAND2 (N3813, N3806, N2870);
xor XOR2 (N3814, N3788, N1416);
xor XOR2 (N3815, N3799, N2373);
and AND3 (N3816, N3815, N730, N213);
xor XOR2 (N3817, N3808, N2236);
xor XOR2 (N3818, N3814, N2346);
buf BUF1 (N3819, N3812);
nand NAND4 (N3820, N3816, N19, N915, N3399);
buf BUF1 (N3821, N3777);
nand NAND4 (N3822, N3820, N3220, N3609, N3613);
and AND4 (N3823, N3819, N2641, N3778, N2712);
and AND4 (N3824, N3802, N3231, N1654, N3798);
and AND4 (N3825, N3822, N3339, N663, N1125);
buf BUF1 (N3826, N3813);
nor NOR3 (N3827, N3810, N1333, N1066);
or OR3 (N3828, N3826, N3482, N870);
or OR2 (N3829, N3825, N940);
and AND3 (N3830, N3818, N1025, N299);
not NOT1 (N3831, N3823);
or OR4 (N3832, N3811, N2387, N183, N1344);
or OR3 (N3833, N3829, N546, N255);
buf BUF1 (N3834, N3830);
nand NAND4 (N3835, N3805, N1150, N3217, N2361);
xor XOR2 (N3836, N3821, N403);
xor XOR2 (N3837, N3834, N1822);
not NOT1 (N3838, N3827);
xor XOR2 (N3839, N3817, N2896);
not NOT1 (N3840, N3839);
nor NOR4 (N3841, N3840, N3335, N498, N1857);
not NOT1 (N3842, N3837);
nor NOR2 (N3843, N3833, N3634);
buf BUF1 (N3844, N3841);
nand NAND4 (N3845, N3835, N1233, N1617, N853);
nor NOR4 (N3846, N3836, N891, N1331, N1697);
not NOT1 (N3847, N3832);
or OR4 (N3848, N3845, N1095, N1636, N505);
nor NOR3 (N3849, N3848, N1925, N717);
nor NOR3 (N3850, N3842, N1476, N3331);
xor XOR2 (N3851, N3828, N323);
nor NOR2 (N3852, N3844, N45);
buf BUF1 (N3853, N3831);
buf BUF1 (N3854, N3850);
not NOT1 (N3855, N3846);
not NOT1 (N3856, N3838);
and AND2 (N3857, N3824, N3189);
not NOT1 (N3858, N3854);
not NOT1 (N3859, N3855);
xor XOR2 (N3860, N3851, N412);
nand NAND2 (N3861, N3852, N1952);
not NOT1 (N3862, N3853);
nor NOR4 (N3863, N3859, N3610, N2393, N2211);
and AND2 (N3864, N3847, N3162);
not NOT1 (N3865, N3864);
xor XOR2 (N3866, N3849, N214);
and AND4 (N3867, N3857, N1144, N2068, N762);
nor NOR3 (N3868, N3867, N3240, N2326);
xor XOR2 (N3869, N3868, N2649);
buf BUF1 (N3870, N3858);
and AND2 (N3871, N3865, N1937);
and AND3 (N3872, N3862, N2563, N2687);
buf BUF1 (N3873, N3870);
xor XOR2 (N3874, N3872, N2852);
and AND3 (N3875, N3873, N1090, N2267);
not NOT1 (N3876, N3861);
not NOT1 (N3877, N3869);
or OR4 (N3878, N3860, N1857, N946, N852);
buf BUF1 (N3879, N3875);
not NOT1 (N3880, N3843);
nand NAND4 (N3881, N3856, N2921, N3709, N2212);
nor NOR4 (N3882, N3863, N3087, N3708, N2958);
nand NAND2 (N3883, N3866, N2692);
xor XOR2 (N3884, N3882, N2461);
buf BUF1 (N3885, N3876);
or OR3 (N3886, N3879, N2811, N1897);
nand NAND2 (N3887, N3886, N1789);
nand NAND3 (N3888, N3874, N1656, N3474);
and AND2 (N3889, N3885, N1552);
xor XOR2 (N3890, N3883, N1376);
buf BUF1 (N3891, N3884);
xor XOR2 (N3892, N3888, N2986);
not NOT1 (N3893, N3889);
nor NOR2 (N3894, N3893, N422);
buf BUF1 (N3895, N3887);
nand NAND3 (N3896, N3880, N2859, N300);
xor XOR2 (N3897, N3871, N612);
buf BUF1 (N3898, N3895);
nand NAND2 (N3899, N3891, N2450);
buf BUF1 (N3900, N3898);
buf BUF1 (N3901, N3897);
buf BUF1 (N3902, N3894);
xor XOR2 (N3903, N3890, N1724);
and AND3 (N3904, N3896, N1617, N2514);
nor NOR4 (N3905, N3892, N446, N2834, N2272);
not NOT1 (N3906, N3899);
xor XOR2 (N3907, N3878, N2537);
or OR3 (N3908, N3901, N1167, N750);
not NOT1 (N3909, N3905);
not NOT1 (N3910, N3881);
nor NOR3 (N3911, N3910, N2034, N182);
not NOT1 (N3912, N3902);
nor NOR2 (N3913, N3900, N757);
nand NAND3 (N3914, N3903, N2870, N1183);
nand NAND2 (N3915, N3904, N3515);
xor XOR2 (N3916, N3911, N1146);
buf BUF1 (N3917, N3913);
nor NOR2 (N3918, N3907, N1929);
buf BUF1 (N3919, N3918);
nor NOR3 (N3920, N3912, N283, N1918);
nor NOR4 (N3921, N3919, N2455, N2101, N3061);
and AND4 (N3922, N3921, N2892, N906, N804);
or OR4 (N3923, N3906, N1346, N353, N2549);
and AND4 (N3924, N3922, N1767, N1974, N76);
not NOT1 (N3925, N3914);
and AND3 (N3926, N3908, N2525, N2811);
and AND4 (N3927, N3925, N3211, N2349, N2011);
nor NOR2 (N3928, N3877, N714);
nand NAND2 (N3929, N3909, N3892);
and AND2 (N3930, N3928, N357);
nor NOR3 (N3931, N3917, N1940, N3329);
nand NAND2 (N3932, N3930, N2938);
nand NAND2 (N3933, N3920, N2163);
xor XOR2 (N3934, N3923, N1940);
and AND3 (N3935, N3931, N2446, N2607);
and AND2 (N3936, N3926, N212);
not NOT1 (N3937, N3932);
nor NOR3 (N3938, N3927, N3336, N1489);
not NOT1 (N3939, N3929);
or OR2 (N3940, N3934, N2385);
and AND3 (N3941, N3935, N3564, N3031);
buf BUF1 (N3942, N3940);
buf BUF1 (N3943, N3937);
and AND3 (N3944, N3939, N2683, N819);
nand NAND3 (N3945, N3943, N87, N1207);
xor XOR2 (N3946, N3924, N338);
nand NAND3 (N3947, N3941, N1005, N1514);
and AND2 (N3948, N3942, N2742);
or OR4 (N3949, N3916, N1443, N2311, N2608);
not NOT1 (N3950, N3946);
nand NAND4 (N3951, N3915, N1261, N3037, N3570);
xor XOR2 (N3952, N3948, N540);
nand NAND3 (N3953, N3947, N3368, N2661);
buf BUF1 (N3954, N3951);
nand NAND3 (N3955, N3950, N3360, N2712);
and AND2 (N3956, N3938, N11);
or OR3 (N3957, N3953, N1963, N3948);
nand NAND2 (N3958, N3956, N2275);
or OR3 (N3959, N3958, N490, N2271);
or OR3 (N3960, N3955, N3049, N373);
nand NAND4 (N3961, N3952, N2634, N2217, N3454);
not NOT1 (N3962, N3960);
or OR4 (N3963, N3944, N1194, N1387, N3463);
xor XOR2 (N3964, N3962, N2200);
or OR3 (N3965, N3957, N2465, N1598);
buf BUF1 (N3966, N3936);
buf BUF1 (N3967, N3945);
or OR2 (N3968, N3965, N348);
nor NOR2 (N3969, N3961, N2530);
not NOT1 (N3970, N3964);
xor XOR2 (N3971, N3970, N281);
nand NAND2 (N3972, N3954, N2975);
and AND2 (N3973, N3963, N703);
xor XOR2 (N3974, N3969, N3451);
or OR3 (N3975, N3971, N2119, N1025);
or OR3 (N3976, N3972, N528, N2878);
not NOT1 (N3977, N3967);
nor NOR2 (N3978, N3968, N3420);
xor XOR2 (N3979, N3975, N3899);
not NOT1 (N3980, N3966);
xor XOR2 (N3981, N3959, N3826);
or OR2 (N3982, N3979, N2588);
nor NOR3 (N3983, N3977, N734, N2643);
nor NOR3 (N3984, N3933, N1089, N2133);
xor XOR2 (N3985, N3980, N1492);
nand NAND2 (N3986, N3976, N1252);
not NOT1 (N3987, N3983);
not NOT1 (N3988, N3949);
buf BUF1 (N3989, N3987);
and AND3 (N3990, N3986, N1499, N3023);
and AND3 (N3991, N3981, N184, N2561);
nand NAND2 (N3992, N3982, N1850);
not NOT1 (N3993, N3991);
xor XOR2 (N3994, N3992, N846);
buf BUF1 (N3995, N3984);
nand NAND4 (N3996, N3973, N1405, N215, N2345);
and AND4 (N3997, N3996, N2029, N1648, N2265);
xor XOR2 (N3998, N3985, N910);
buf BUF1 (N3999, N3974);
and AND3 (N4000, N3978, N2951, N549);
nand NAND4 (N4001, N3998, N1319, N2721, N2608);
xor XOR2 (N4002, N3999, N1074);
buf BUF1 (N4003, N3990);
xor XOR2 (N4004, N4003, N1322);
nor NOR3 (N4005, N3989, N1362, N3039);
nor NOR2 (N4006, N4002, N3952);
buf BUF1 (N4007, N3988);
nand NAND4 (N4008, N4006, N2112, N1755, N2360);
or OR3 (N4009, N4001, N1712, N1859);
nor NOR4 (N4010, N4000, N1364, N638, N2873);
not NOT1 (N4011, N4005);
buf BUF1 (N4012, N4008);
buf BUF1 (N4013, N4011);
not NOT1 (N4014, N3994);
nand NAND4 (N4015, N4009, N2030, N2901, N570);
and AND4 (N4016, N4012, N3238, N1275, N2655);
buf BUF1 (N4017, N4010);
or OR3 (N4018, N3993, N3247, N2679);
not NOT1 (N4019, N3997);
and AND4 (N4020, N3995, N2410, N189, N475);
buf BUF1 (N4021, N4013);
or OR4 (N4022, N4016, N2341, N1933, N396);
nor NOR3 (N4023, N4018, N837, N2672);
nand NAND4 (N4024, N4015, N2350, N1575, N3491);
and AND3 (N4025, N4019, N1543, N3018);
or OR4 (N4026, N4014, N1596, N765, N1046);
nor NOR2 (N4027, N4004, N1023);
nor NOR2 (N4028, N4023, N482);
nor NOR4 (N4029, N4020, N520, N1201, N1044);
nor NOR4 (N4030, N4024, N1681, N179, N2419);
nor NOR4 (N4031, N4030, N1101, N591, N537);
and AND3 (N4032, N4031, N3053, N2904);
nand NAND2 (N4033, N4029, N2920);
not NOT1 (N4034, N4033);
not NOT1 (N4035, N4026);
and AND3 (N4036, N4007, N313, N2286);
nor NOR3 (N4037, N4022, N2837, N160);
not NOT1 (N4038, N4037);
xor XOR2 (N4039, N4032, N1194);
xor XOR2 (N4040, N4038, N3129);
or OR2 (N4041, N4034, N3180);
not NOT1 (N4042, N4035);
and AND3 (N4043, N4027, N1491, N396);
nand NAND4 (N4044, N4028, N1548, N1795, N1299);
or OR2 (N4045, N4042, N1439);
nor NOR3 (N4046, N4025, N2102, N3799);
nand NAND2 (N4047, N4039, N2262);
nor NOR2 (N4048, N4047, N656);
or OR2 (N4049, N4048, N471);
xor XOR2 (N4050, N4045, N1836);
nand NAND3 (N4051, N4040, N1631, N3050);
xor XOR2 (N4052, N4050, N1608);
or OR2 (N4053, N4049, N1449);
nor NOR2 (N4054, N4051, N1991);
nand NAND4 (N4055, N4036, N1008, N623, N1815);
not NOT1 (N4056, N4054);
xor XOR2 (N4057, N4046, N8);
and AND2 (N4058, N4053, N1839);
not NOT1 (N4059, N4055);
nand NAND3 (N4060, N4056, N1625, N2347);
or OR3 (N4061, N4021, N267, N2171);
buf BUF1 (N4062, N4060);
nand NAND4 (N4063, N4043, N2756, N414, N1763);
and AND3 (N4064, N4058, N1139, N605);
and AND3 (N4065, N4062, N3491, N2148);
buf BUF1 (N4066, N4063);
nor NOR4 (N4067, N4017, N648, N2075, N3639);
xor XOR2 (N4068, N4065, N4059);
nand NAND3 (N4069, N1516, N2328, N1707);
xor XOR2 (N4070, N4066, N1013);
not NOT1 (N4071, N4069);
not NOT1 (N4072, N4057);
xor XOR2 (N4073, N4072, N2029);
buf BUF1 (N4074, N4070);
nor NOR3 (N4075, N4074, N3772, N1717);
and AND3 (N4076, N4071, N2226, N3780);
nand NAND2 (N4077, N4073, N496);
and AND3 (N4078, N4075, N3367, N3604);
and AND2 (N4079, N4068, N1509);
xor XOR2 (N4080, N4052, N394);
nand NAND2 (N4081, N4067, N1165);
nor NOR2 (N4082, N4044, N3482);
nor NOR4 (N4083, N4077, N1320, N515, N2996);
not NOT1 (N4084, N4041);
or OR3 (N4085, N4064, N524, N2184);
nand NAND3 (N4086, N4079, N946, N2518);
nor NOR2 (N4087, N4082, N494);
buf BUF1 (N4088, N4085);
and AND4 (N4089, N4086, N1009, N608, N316);
buf BUF1 (N4090, N4087);
nor NOR3 (N4091, N4080, N3555, N1398);
nor NOR3 (N4092, N4076, N513, N2648);
nor NOR3 (N4093, N4092, N1181, N346);
nand NAND2 (N4094, N4088, N1436);
and AND2 (N4095, N4078, N1288);
nor NOR2 (N4096, N4089, N2730);
or OR2 (N4097, N4091, N498);
nor NOR2 (N4098, N4094, N974);
xor XOR2 (N4099, N4097, N746);
or OR3 (N4100, N4096, N858, N1380);
or OR2 (N4101, N4093, N3792);
nand NAND2 (N4102, N4083, N3530);
nor NOR2 (N4103, N4095, N3943);
nor NOR4 (N4104, N4100, N515, N489, N3253);
or OR2 (N4105, N4103, N2542);
nor NOR2 (N4106, N4081, N3353);
xor XOR2 (N4107, N4106, N1008);
xor XOR2 (N4108, N4102, N3410);
nand NAND3 (N4109, N4061, N1334, N2960);
not NOT1 (N4110, N4101);
not NOT1 (N4111, N4099);
or OR2 (N4112, N4107, N3040);
not NOT1 (N4113, N4110);
nand NAND3 (N4114, N4108, N1986, N1045);
nor NOR2 (N4115, N4105, N2435);
xor XOR2 (N4116, N4114, N2605);
nand NAND3 (N4117, N4111, N678, N642);
nor NOR4 (N4118, N4116, N3126, N975, N2960);
or OR3 (N4119, N4098, N2767, N3769);
not NOT1 (N4120, N4104);
buf BUF1 (N4121, N4115);
not NOT1 (N4122, N4117);
nor NOR2 (N4123, N4121, N96);
or OR4 (N4124, N4084, N2764, N3761, N374);
or OR2 (N4125, N4120, N1708);
or OR3 (N4126, N4119, N3100, N3578);
nor NOR3 (N4127, N4126, N3190, N2784);
nand NAND2 (N4128, N4124, N305);
nand NAND4 (N4129, N4118, N220, N1264, N552);
buf BUF1 (N4130, N4109);
nor NOR4 (N4131, N4090, N2473, N2676, N3870);
nor NOR2 (N4132, N4127, N634);
xor XOR2 (N4133, N4123, N3643);
xor XOR2 (N4134, N4131, N112);
not NOT1 (N4135, N4130);
not NOT1 (N4136, N4134);
buf BUF1 (N4137, N4132);
nor NOR3 (N4138, N4129, N1595, N2227);
or OR2 (N4139, N4125, N587);
nand NAND2 (N4140, N4138, N3349);
buf BUF1 (N4141, N4137);
buf BUF1 (N4142, N4135);
nand NAND3 (N4143, N4139, N1492, N4118);
buf BUF1 (N4144, N4113);
nand NAND3 (N4145, N4122, N3678, N1825);
xor XOR2 (N4146, N4142, N1613);
not NOT1 (N4147, N4140);
buf BUF1 (N4148, N4128);
nand NAND4 (N4149, N4147, N3881, N2790, N1062);
nand NAND3 (N4150, N4112, N674, N3513);
buf BUF1 (N4151, N4149);
nand NAND2 (N4152, N4151, N3287);
or OR2 (N4153, N4146, N747);
not NOT1 (N4154, N4136);
nand NAND2 (N4155, N4143, N2051);
buf BUF1 (N4156, N4152);
or OR2 (N4157, N4155, N3460);
and AND2 (N4158, N4156, N3996);
nor NOR2 (N4159, N4154, N793);
nand NAND4 (N4160, N4133, N3424, N1053, N1029);
buf BUF1 (N4161, N4145);
not NOT1 (N4162, N4148);
and AND2 (N4163, N4159, N2433);
xor XOR2 (N4164, N4150, N2880);
buf BUF1 (N4165, N4144);
or OR3 (N4166, N4153, N1558, N99);
or OR3 (N4167, N4163, N879, N1935);
buf BUF1 (N4168, N4164);
buf BUF1 (N4169, N4167);
not NOT1 (N4170, N4161);
nand NAND2 (N4171, N4157, N590);
and AND3 (N4172, N4158, N4126, N3012);
nand NAND4 (N4173, N4141, N119, N2498, N1559);
xor XOR2 (N4174, N4173, N3737);
xor XOR2 (N4175, N4166, N1890);
not NOT1 (N4176, N4174);
nand NAND4 (N4177, N4175, N522, N109, N4114);
or OR3 (N4178, N4171, N3513, N1683);
or OR4 (N4179, N4169, N749, N2130, N1707);
nand NAND2 (N4180, N4170, N2523);
and AND4 (N4181, N4179, N780, N1643, N2852);
xor XOR2 (N4182, N4176, N1461);
nand NAND4 (N4183, N4162, N173, N2465, N2759);
not NOT1 (N4184, N4181);
nand NAND4 (N4185, N4184, N3815, N1878, N897);
xor XOR2 (N4186, N4172, N2987);
or OR4 (N4187, N4183, N3174, N1816, N2826);
not NOT1 (N4188, N4177);
not NOT1 (N4189, N4188);
not NOT1 (N4190, N4165);
buf BUF1 (N4191, N4190);
or OR3 (N4192, N4185, N3967, N3993);
nor NOR4 (N4193, N4160, N3509, N3499, N1519);
and AND2 (N4194, N4192, N3396);
buf BUF1 (N4195, N4186);
not NOT1 (N4196, N4187);
xor XOR2 (N4197, N4193, N4001);
not NOT1 (N4198, N4182);
or OR4 (N4199, N4189, N3425, N1821, N1752);
nand NAND2 (N4200, N4178, N1777);
or OR2 (N4201, N4168, N1631);
and AND3 (N4202, N4200, N2732, N2930);
or OR2 (N4203, N4194, N1039);
buf BUF1 (N4204, N4203);
not NOT1 (N4205, N4197);
and AND4 (N4206, N4205, N1443, N3542, N1528);
nand NAND4 (N4207, N4199, N1970, N1370, N2087);
and AND2 (N4208, N4180, N334);
or OR2 (N4209, N4208, N3356);
nor NOR3 (N4210, N4202, N632, N1349);
nand NAND3 (N4211, N4206, N1304, N1443);
nor NOR3 (N4212, N4211, N3685, N3);
or OR3 (N4213, N4212, N768, N1237);
and AND3 (N4214, N4191, N140, N4212);
xor XOR2 (N4215, N4195, N2563);
nand NAND2 (N4216, N4198, N3057);
nor NOR2 (N4217, N4210, N2630);
nand NAND2 (N4218, N4217, N570);
nand NAND2 (N4219, N4201, N406);
buf BUF1 (N4220, N4213);
and AND2 (N4221, N4214, N808);
not NOT1 (N4222, N4220);
or OR3 (N4223, N4222, N2707, N2759);
nand NAND3 (N4224, N4223, N333, N1421);
xor XOR2 (N4225, N4221, N146);
nand NAND4 (N4226, N4207, N3767, N2787, N2764);
buf BUF1 (N4227, N4225);
not NOT1 (N4228, N4226);
not NOT1 (N4229, N4215);
nand NAND4 (N4230, N4229, N1047, N4132, N587);
or OR2 (N4231, N4204, N3023);
buf BUF1 (N4232, N4228);
buf BUF1 (N4233, N4224);
nor NOR3 (N4234, N4216, N3957, N1772);
xor XOR2 (N4235, N4218, N3119);
buf BUF1 (N4236, N4230);
and AND2 (N4237, N4219, N843);
xor XOR2 (N4238, N4233, N2645);
nor NOR3 (N4239, N4209, N1106, N3255);
xor XOR2 (N4240, N4196, N1550);
nor NOR4 (N4241, N4236, N1094, N1582, N2935);
and AND4 (N4242, N4231, N3211, N365, N743);
nor NOR4 (N4243, N4238, N884, N2683, N3238);
or OR3 (N4244, N4234, N1228, N3101);
nand NAND3 (N4245, N4235, N2692, N3095);
nor NOR4 (N4246, N4237, N1402, N571, N1750);
nand NAND3 (N4247, N4244, N1133, N3381);
not NOT1 (N4248, N4242);
and AND3 (N4249, N4246, N2322, N2810);
and AND3 (N4250, N4239, N549, N3858);
and AND4 (N4251, N4241, N1938, N4212, N3720);
not NOT1 (N4252, N4243);
nor NOR3 (N4253, N4249, N3344, N3258);
nand NAND3 (N4254, N4240, N2195, N315);
and AND2 (N4255, N4245, N2288);
buf BUF1 (N4256, N4251);
xor XOR2 (N4257, N4232, N1186);
and AND3 (N4258, N4257, N3785, N1678);
nand NAND2 (N4259, N4227, N3441);
nand NAND4 (N4260, N4258, N2185, N2339, N3945);
and AND3 (N4261, N4250, N1085, N1160);
xor XOR2 (N4262, N4252, N3426);
or OR3 (N4263, N4261, N2667, N3474);
buf BUF1 (N4264, N4256);
and AND3 (N4265, N4264, N3047, N4261);
not NOT1 (N4266, N4247);
nand NAND3 (N4267, N4262, N831, N123);
nor NOR4 (N4268, N4260, N770, N268, N3632);
nor NOR4 (N4269, N4259, N2571, N110, N4152);
xor XOR2 (N4270, N4254, N3954);
xor XOR2 (N4271, N4265, N3801);
nand NAND4 (N4272, N4270, N1699, N2446, N2318);
and AND4 (N4273, N4263, N589, N2581, N2534);
nand NAND2 (N4274, N4273, N1598);
buf BUF1 (N4275, N4266);
nor NOR3 (N4276, N4255, N1253, N802);
xor XOR2 (N4277, N4276, N425);
or OR2 (N4278, N4274, N4052);
or OR2 (N4279, N4269, N2451);
and AND3 (N4280, N4272, N2605, N122);
nor NOR4 (N4281, N4267, N2516, N3602, N835);
not NOT1 (N4282, N4277);
nand NAND2 (N4283, N4280, N1912);
xor XOR2 (N4284, N4279, N2632);
nand NAND2 (N4285, N4268, N523);
or OR4 (N4286, N4281, N1085, N1865, N273);
xor XOR2 (N4287, N4285, N2024);
nor NOR3 (N4288, N4271, N1229, N1584);
nor NOR4 (N4289, N4253, N2431, N3457, N3226);
nand NAND4 (N4290, N4275, N273, N1927, N2644);
not NOT1 (N4291, N4289);
nor NOR2 (N4292, N4291, N1581);
nor NOR3 (N4293, N4278, N3980, N1229);
nand NAND4 (N4294, N4290, N1061, N281, N70);
and AND2 (N4295, N4282, N879);
and AND2 (N4296, N4284, N1687);
and AND3 (N4297, N4287, N2187, N627);
nand NAND3 (N4298, N4295, N3500, N3624);
not NOT1 (N4299, N4248);
xor XOR2 (N4300, N4293, N1888);
not NOT1 (N4301, N4296);
nand NAND3 (N4302, N4300, N476, N567);
and AND4 (N4303, N4301, N1311, N3169, N1232);
nand NAND2 (N4304, N4297, N612);
and AND4 (N4305, N4303, N2016, N759, N2064);
not NOT1 (N4306, N4286);
xor XOR2 (N4307, N4298, N2809);
nor NOR4 (N4308, N4292, N1051, N2580, N3619);
nor NOR3 (N4309, N4307, N4149, N1820);
or OR4 (N4310, N4305, N3061, N2923, N1666);
xor XOR2 (N4311, N4288, N3530);
nand NAND2 (N4312, N4310, N133);
xor XOR2 (N4313, N4283, N1708);
nand NAND3 (N4314, N4309, N2403, N1767);
nor NOR2 (N4315, N4313, N2136);
or OR4 (N4316, N4308, N302, N1088, N904);
xor XOR2 (N4317, N4314, N4205);
nor NOR3 (N4318, N4312, N1003, N2446);
xor XOR2 (N4319, N4302, N2384);
and AND3 (N4320, N4294, N3761, N2206);
nor NOR2 (N4321, N4304, N3258);
xor XOR2 (N4322, N4320, N3179);
or OR2 (N4323, N4306, N862);
nor NOR2 (N4324, N4321, N948);
not NOT1 (N4325, N4315);
buf BUF1 (N4326, N4299);
nor NOR3 (N4327, N4325, N3658, N2308);
or OR4 (N4328, N4326, N2639, N4182, N2427);
or OR3 (N4329, N4316, N2097, N1528);
nand NAND3 (N4330, N4322, N1263, N2421);
and AND4 (N4331, N4330, N2457, N236, N1326);
xor XOR2 (N4332, N4328, N4318);
nor NOR4 (N4333, N2484, N1063, N2254, N56);
or OR2 (N4334, N4324, N277);
and AND2 (N4335, N4332, N2828);
not NOT1 (N4336, N4319);
or OR2 (N4337, N4335, N3534);
xor XOR2 (N4338, N4334, N4204);
xor XOR2 (N4339, N4311, N2987);
nand NAND2 (N4340, N4338, N2685);
or OR3 (N4341, N4331, N3522, N1159);
xor XOR2 (N4342, N4317, N2744);
nor NOR4 (N4343, N4341, N4336, N3349, N1415);
nand NAND2 (N4344, N824, N723);
nand NAND4 (N4345, N4339, N1940, N167, N2006);
or OR3 (N4346, N4337, N1163, N4016);
and AND4 (N4347, N4333, N589, N3046, N2793);
nor NOR3 (N4348, N4340, N829, N756);
nand NAND3 (N4349, N4345, N1087, N2927);
and AND3 (N4350, N4327, N4178, N2578);
xor XOR2 (N4351, N4349, N997);
buf BUF1 (N4352, N4343);
nand NAND4 (N4353, N4342, N2270, N865, N1063);
not NOT1 (N4354, N4348);
or OR2 (N4355, N4351, N4213);
nand NAND4 (N4356, N4354, N1866, N3284, N1984);
and AND3 (N4357, N4353, N1117, N2463);
nor NOR4 (N4358, N4356, N1551, N1963, N206);
or OR3 (N4359, N4350, N988, N4312);
nor NOR2 (N4360, N4329, N2973);
or OR2 (N4361, N4346, N1318);
nand NAND3 (N4362, N4361, N3081, N2251);
xor XOR2 (N4363, N4358, N2381);
or OR3 (N4364, N4357, N2415, N3001);
nor NOR4 (N4365, N4362, N2267, N4226, N3621);
nand NAND4 (N4366, N4360, N3561, N401, N1668);
or OR3 (N4367, N4323, N821, N2191);
xor XOR2 (N4368, N4366, N1209);
nor NOR4 (N4369, N4355, N1337, N3683, N830);
xor XOR2 (N4370, N4364, N3930);
and AND3 (N4371, N4352, N4354, N3726);
xor XOR2 (N4372, N4365, N2645);
buf BUF1 (N4373, N4367);
nor NOR4 (N4374, N4370, N1293, N1844, N2141);
nand NAND3 (N4375, N4369, N4369, N1386);
buf BUF1 (N4376, N4375);
nand NAND4 (N4377, N4372, N225, N1816, N2030);
not NOT1 (N4378, N4374);
not NOT1 (N4379, N4378);
or OR4 (N4380, N4347, N2028, N1907, N361);
not NOT1 (N4381, N4373);
xor XOR2 (N4382, N4377, N4169);
not NOT1 (N4383, N4363);
xor XOR2 (N4384, N4383, N2694);
not NOT1 (N4385, N4359);
xor XOR2 (N4386, N4344, N656);
buf BUF1 (N4387, N4376);
nor NOR3 (N4388, N4380, N1912, N715);
or OR2 (N4389, N4371, N3766);
nor NOR2 (N4390, N4382, N1380);
not NOT1 (N4391, N4368);
not NOT1 (N4392, N4390);
and AND2 (N4393, N4388, N1739);
nor NOR3 (N4394, N4384, N4060, N1500);
and AND4 (N4395, N4394, N3930, N1484, N3880);
not NOT1 (N4396, N4386);
or OR4 (N4397, N4396, N281, N3127, N1284);
xor XOR2 (N4398, N4391, N870);
and AND2 (N4399, N4387, N4081);
and AND3 (N4400, N4379, N1333, N3355);
or OR3 (N4401, N4395, N881, N4208);
not NOT1 (N4402, N4401);
nand NAND3 (N4403, N4400, N3688, N695);
nor NOR3 (N4404, N4402, N4215, N2221);
not NOT1 (N4405, N4381);
xor XOR2 (N4406, N4385, N308);
xor XOR2 (N4407, N4406, N3651);
nor NOR4 (N4408, N4397, N3240, N2506, N328);
nand NAND2 (N4409, N4392, N1568);
and AND4 (N4410, N4398, N2307, N148, N1056);
xor XOR2 (N4411, N4389, N249);
nor NOR2 (N4412, N4410, N1484);
nor NOR3 (N4413, N4399, N3037, N1347);
and AND3 (N4414, N4393, N513, N2129);
and AND3 (N4415, N4409, N189, N3171);
nor NOR3 (N4416, N4408, N2607, N3594);
buf BUF1 (N4417, N4412);
nand NAND3 (N4418, N4405, N1048, N667);
and AND2 (N4419, N4404, N4249);
nand NAND2 (N4420, N4419, N4173);
and AND3 (N4421, N4411, N3608, N3664);
or OR3 (N4422, N4407, N1972, N1719);
nor NOR4 (N4423, N4421, N1148, N1939, N3282);
or OR3 (N4424, N4418, N4008, N2165);
not NOT1 (N4425, N4414);
and AND3 (N4426, N4420, N890, N3624);
or OR4 (N4427, N4413, N1026, N3128, N3081);
or OR2 (N4428, N4422, N2413);
and AND3 (N4429, N4417, N1793, N491);
nor NOR4 (N4430, N4416, N2385, N1927, N2764);
buf BUF1 (N4431, N4403);
not NOT1 (N4432, N4429);
not NOT1 (N4433, N4427);
or OR4 (N4434, N4423, N3916, N2965, N1913);
and AND3 (N4435, N4433, N605, N1488);
and AND2 (N4436, N4426, N3041);
xor XOR2 (N4437, N4424, N1886);
or OR4 (N4438, N4425, N2862, N3450, N4047);
buf BUF1 (N4439, N4434);
not NOT1 (N4440, N4437);
buf BUF1 (N4441, N4432);
nor NOR3 (N4442, N4431, N1751, N1469);
and AND2 (N4443, N4415, N2120);
nand NAND3 (N4444, N4435, N844, N3189);
nor NOR2 (N4445, N4440, N2217);
nand NAND4 (N4446, N4428, N1487, N201, N3018);
and AND4 (N4447, N4444, N3016, N1062, N3098);
not NOT1 (N4448, N4439);
not NOT1 (N4449, N4447);
nor NOR4 (N4450, N4448, N1467, N2820, N4287);
and AND2 (N4451, N4441, N1084);
xor XOR2 (N4452, N4430, N836);
xor XOR2 (N4453, N4442, N470);
nor NOR4 (N4454, N4450, N1231, N4092, N2918);
or OR2 (N4455, N4454, N3499);
xor XOR2 (N4456, N4453, N2187);
nor NOR3 (N4457, N4452, N3240, N341);
not NOT1 (N4458, N4457);
nor NOR4 (N4459, N4451, N2356, N1853, N303);
not NOT1 (N4460, N4443);
not NOT1 (N4461, N4460);
nand NAND4 (N4462, N4446, N3849, N1986, N2624);
or OR4 (N4463, N4462, N2034, N2179, N3104);
buf BUF1 (N4464, N4449);
or OR4 (N4465, N4463, N3506, N2187, N1676);
not NOT1 (N4466, N4461);
xor XOR2 (N4467, N4438, N4072);
nor NOR4 (N4468, N4456, N4369, N1081, N1560);
and AND3 (N4469, N4445, N2801, N1393);
buf BUF1 (N4470, N4455);
nor NOR4 (N4471, N4468, N399, N2069, N4041);
xor XOR2 (N4472, N4465, N503);
buf BUF1 (N4473, N4459);
buf BUF1 (N4474, N4471);
or OR4 (N4475, N4467, N472, N2404, N2127);
buf BUF1 (N4476, N4458);
and AND4 (N4477, N4473, N711, N1183, N3607);
nand NAND3 (N4478, N4475, N1336, N149);
or OR3 (N4479, N4474, N1831, N587);
and AND4 (N4480, N4464, N3386, N2180, N3941);
and AND3 (N4481, N4477, N4373, N2332);
xor XOR2 (N4482, N4481, N2865);
and AND4 (N4483, N4479, N3775, N955, N2826);
or OR2 (N4484, N4480, N3764);
not NOT1 (N4485, N4472);
nor NOR4 (N4486, N4484, N1640, N3916, N2671);
not NOT1 (N4487, N4478);
and AND3 (N4488, N4483, N2716, N1394);
not NOT1 (N4489, N4487);
and AND4 (N4490, N4469, N2195, N594, N3032);
not NOT1 (N4491, N4436);
not NOT1 (N4492, N4490);
not NOT1 (N4493, N4486);
not NOT1 (N4494, N4466);
or OR3 (N4495, N4492, N2088, N1352);
or OR2 (N4496, N4482, N433);
nand NAND3 (N4497, N4488, N2260, N238);
and AND4 (N4498, N4495, N1672, N4327, N925);
xor XOR2 (N4499, N4489, N1938);
or OR3 (N4500, N4476, N2418, N4174);
nor NOR3 (N4501, N4493, N2386, N177);
nor NOR3 (N4502, N4494, N631, N1691);
not NOT1 (N4503, N4491);
nand NAND3 (N4504, N4485, N1464, N453);
not NOT1 (N4505, N4502);
not NOT1 (N4506, N4504);
xor XOR2 (N4507, N4506, N1399);
not NOT1 (N4508, N4497);
nand NAND4 (N4509, N4498, N1930, N2936, N3685);
or OR4 (N4510, N4509, N646, N1008, N1412);
not NOT1 (N4511, N4499);
nand NAND2 (N4512, N4470, N3251);
not NOT1 (N4513, N4512);
xor XOR2 (N4514, N4513, N288);
or OR4 (N4515, N4500, N1333, N2160, N3275);
nor NOR3 (N4516, N4501, N2358, N3892);
and AND3 (N4517, N4511, N1708, N2811);
not NOT1 (N4518, N4516);
xor XOR2 (N4519, N4515, N1155);
xor XOR2 (N4520, N4507, N1879);
nand NAND3 (N4521, N4510, N4017, N925);
buf BUF1 (N4522, N4503);
nand NAND4 (N4523, N4508, N3127, N3282, N1583);
or OR2 (N4524, N4518, N504);
buf BUF1 (N4525, N4524);
and AND3 (N4526, N4525, N2434, N2837);
nor NOR3 (N4527, N4505, N3305, N2517);
not NOT1 (N4528, N4496);
not NOT1 (N4529, N4528);
nor NOR3 (N4530, N4526, N2569, N2638);
not NOT1 (N4531, N4527);
not NOT1 (N4532, N4531);
nor NOR3 (N4533, N4514, N3216, N2182);
or OR4 (N4534, N4532, N2915, N1990, N57);
buf BUF1 (N4535, N4522);
nand NAND3 (N4536, N4523, N2211, N511);
nand NAND3 (N4537, N4536, N274, N3877);
buf BUF1 (N4538, N4521);
buf BUF1 (N4539, N4520);
buf BUF1 (N4540, N4535);
nand NAND4 (N4541, N4539, N1375, N3813, N3805);
and AND3 (N4542, N4541, N1700, N3708);
xor XOR2 (N4543, N4542, N3844);
or OR4 (N4544, N4517, N1159, N797, N1632);
or OR3 (N4545, N4538, N151, N2545);
xor XOR2 (N4546, N4533, N3241);
and AND2 (N4547, N4545, N3787);
buf BUF1 (N4548, N4537);
and AND3 (N4549, N4544, N4213, N3056);
buf BUF1 (N4550, N4534);
nor NOR4 (N4551, N4547, N3749, N2418, N4229);
buf BUF1 (N4552, N4530);
and AND4 (N4553, N4549, N3053, N690, N1184);
and AND4 (N4554, N4519, N1117, N1451, N351);
nand NAND4 (N4555, N4529, N1472, N1198, N4137);
and AND4 (N4556, N4555, N77, N882, N4519);
and AND3 (N4557, N4548, N1563, N1981);
xor XOR2 (N4558, N4553, N1289);
buf BUF1 (N4559, N4540);
not NOT1 (N4560, N4557);
and AND4 (N4561, N4546, N2613, N3738, N3611);
buf BUF1 (N4562, N4543);
xor XOR2 (N4563, N4560, N760);
nor NOR2 (N4564, N4561, N3081);
nor NOR4 (N4565, N4564, N295, N656, N3196);
nor NOR2 (N4566, N4552, N2012);
nor NOR4 (N4567, N4563, N4224, N1100, N4461);
xor XOR2 (N4568, N4551, N1780);
xor XOR2 (N4569, N4568, N673);
nand NAND3 (N4570, N4550, N4218, N230);
nor NOR2 (N4571, N4566, N3129);
and AND2 (N4572, N4554, N485);
or OR2 (N4573, N4567, N3041);
nor NOR2 (N4574, N4570, N840);
buf BUF1 (N4575, N4572);
nor NOR2 (N4576, N4574, N3194);
or OR4 (N4577, N4573, N921, N3899, N4426);
not NOT1 (N4578, N4569);
or OR2 (N4579, N4559, N3042);
buf BUF1 (N4580, N4577);
buf BUF1 (N4581, N4576);
and AND3 (N4582, N4565, N594, N882);
buf BUF1 (N4583, N4571);
buf BUF1 (N4584, N4581);
not NOT1 (N4585, N4575);
and AND4 (N4586, N4556, N2034, N1904, N4563);
not NOT1 (N4587, N4579);
or OR4 (N4588, N4562, N2459, N904, N446);
and AND4 (N4589, N4582, N353, N349, N729);
nand NAND3 (N4590, N4583, N4419, N2163);
and AND4 (N4591, N4578, N3604, N988, N2084);
nor NOR3 (N4592, N4586, N2449, N3677);
or OR2 (N4593, N4558, N2561);
xor XOR2 (N4594, N4590, N2236);
xor XOR2 (N4595, N4594, N2147);
or OR4 (N4596, N4595, N2675, N2619, N3054);
or OR2 (N4597, N4593, N827);
or OR3 (N4598, N4584, N4141, N4055);
nor NOR4 (N4599, N4580, N804, N2714, N718);
nand NAND4 (N4600, N4589, N496, N1811, N247);
nand NAND4 (N4601, N4588, N886, N4093, N2395);
not NOT1 (N4602, N4585);
and AND3 (N4603, N4601, N691, N3487);
buf BUF1 (N4604, N4603);
buf BUF1 (N4605, N4599);
and AND4 (N4606, N4600, N3023, N1252, N233);
nand NAND4 (N4607, N4592, N4337, N2125, N2819);
nor NOR4 (N4608, N4604, N3505, N4258, N3808);
buf BUF1 (N4609, N4591);
xor XOR2 (N4610, N4597, N3198);
xor XOR2 (N4611, N4606, N268);
or OR4 (N4612, N4605, N1068, N4486, N1423);
or OR3 (N4613, N4609, N4095, N187);
nand NAND2 (N4614, N4602, N4523);
xor XOR2 (N4615, N4607, N1904);
and AND2 (N4616, N4613, N1016);
nand NAND2 (N4617, N4610, N960);
nand NAND2 (N4618, N4616, N812);
nand NAND2 (N4619, N4614, N2994);
xor XOR2 (N4620, N4619, N2660);
nand NAND2 (N4621, N4617, N2096);
buf BUF1 (N4622, N4596);
buf BUF1 (N4623, N4621);
not NOT1 (N4624, N4587);
or OR2 (N4625, N4623, N4497);
not NOT1 (N4626, N4622);
buf BUF1 (N4627, N4598);
and AND4 (N4628, N4618, N1233, N399, N3197);
nor NOR2 (N4629, N4626, N4413);
nand NAND3 (N4630, N4629, N1646, N548);
nor NOR3 (N4631, N4611, N1543, N4515);
and AND3 (N4632, N4615, N1896, N671);
nand NAND3 (N4633, N4612, N3665, N3385);
xor XOR2 (N4634, N4608, N4014);
xor XOR2 (N4635, N4625, N1783);
and AND3 (N4636, N4633, N1484, N507);
xor XOR2 (N4637, N4634, N462);
nand NAND2 (N4638, N4632, N4237);
xor XOR2 (N4639, N4635, N4247);
buf BUF1 (N4640, N4620);
or OR3 (N4641, N4628, N187, N3208);
buf BUF1 (N4642, N4624);
or OR3 (N4643, N4630, N4115, N3336);
buf BUF1 (N4644, N4640);
nand NAND4 (N4645, N4643, N4187, N3325, N3899);
and AND4 (N4646, N4636, N1057, N860, N2645);
nor NOR3 (N4647, N4642, N3247, N2026);
xor XOR2 (N4648, N4646, N2935);
and AND3 (N4649, N4641, N2700, N148);
buf BUF1 (N4650, N4649);
xor XOR2 (N4651, N4631, N1141);
nand NAND4 (N4652, N4645, N3699, N2360, N4610);
or OR2 (N4653, N4648, N3972);
buf BUF1 (N4654, N4650);
buf BUF1 (N4655, N4653);
not NOT1 (N4656, N4647);
and AND3 (N4657, N4654, N3452, N4628);
xor XOR2 (N4658, N4638, N325);
and AND3 (N4659, N4637, N3619, N646);
nor NOR2 (N4660, N4644, N2868);
and AND4 (N4661, N4658, N272, N3253, N4388);
nand NAND4 (N4662, N4655, N3622, N4314, N330);
nor NOR2 (N4663, N4662, N4008);
and AND4 (N4664, N4660, N534, N633, N2453);
or OR2 (N4665, N4659, N766);
xor XOR2 (N4666, N4652, N745);
xor XOR2 (N4667, N4663, N2742);
xor XOR2 (N4668, N4665, N4040);
nor NOR4 (N4669, N4667, N2941, N2766, N4549);
nor NOR3 (N4670, N4656, N282, N1701);
nand NAND2 (N4671, N4661, N4633);
xor XOR2 (N4672, N4670, N1303);
or OR2 (N4673, N4657, N354);
nor NOR4 (N4674, N4651, N1848, N4140, N1949);
nand NAND2 (N4675, N4671, N166);
nand NAND2 (N4676, N4673, N3585);
nor NOR4 (N4677, N4674, N3443, N1304, N1979);
not NOT1 (N4678, N4639);
nand NAND2 (N4679, N4666, N1127);
nor NOR2 (N4680, N4668, N1268);
buf BUF1 (N4681, N4672);
nor NOR2 (N4682, N4678, N4185);
not NOT1 (N4683, N4664);
and AND3 (N4684, N4680, N3676, N736);
not NOT1 (N4685, N4681);
nand NAND4 (N4686, N4685, N948, N4530, N583);
xor XOR2 (N4687, N4682, N4164);
and AND4 (N4688, N4676, N1869, N961, N3418);
buf BUF1 (N4689, N4675);
nand NAND4 (N4690, N4687, N2296, N1978, N359);
xor XOR2 (N4691, N4688, N2584);
and AND3 (N4692, N4689, N1939, N1996);
not NOT1 (N4693, N4669);
xor XOR2 (N4694, N4693, N2214);
nor NOR3 (N4695, N4683, N2509, N1275);
not NOT1 (N4696, N4692);
xor XOR2 (N4697, N4679, N2056);
not NOT1 (N4698, N4695);
buf BUF1 (N4699, N4627);
or OR2 (N4700, N4698, N3696);
nor NOR4 (N4701, N4690, N3319, N3379, N330);
or OR4 (N4702, N4686, N3134, N2457, N3795);
nand NAND3 (N4703, N4701, N2862, N2709);
and AND2 (N4704, N4696, N4618);
xor XOR2 (N4705, N4699, N4051);
or OR4 (N4706, N4694, N3817, N3776, N175);
not NOT1 (N4707, N4705);
nand NAND3 (N4708, N4704, N2593, N2426);
or OR4 (N4709, N4703, N2381, N2522, N3532);
or OR3 (N4710, N4700, N3277, N912);
nor NOR4 (N4711, N4691, N3015, N2279, N2698);
nand NAND4 (N4712, N4710, N1484, N4199, N1124);
buf BUF1 (N4713, N4712);
buf BUF1 (N4714, N4684);
or OR4 (N4715, N4713, N3715, N4455, N390);
and AND2 (N4716, N4706, N2447);
and AND2 (N4717, N4711, N1290);
nor NOR4 (N4718, N4708, N3147, N4281, N191);
or OR4 (N4719, N4718, N1240, N2187, N4478);
xor XOR2 (N4720, N4697, N1053);
buf BUF1 (N4721, N4714);
nor NOR3 (N4722, N4702, N3139, N3420);
and AND2 (N4723, N4715, N2939);
buf BUF1 (N4724, N4719);
or OR2 (N4725, N4717, N4225);
and AND4 (N4726, N4722, N2065, N898, N4484);
buf BUF1 (N4727, N4726);
nand NAND2 (N4728, N4707, N1565);
nor NOR2 (N4729, N4716, N1133);
xor XOR2 (N4730, N4724, N829);
buf BUF1 (N4731, N4725);
xor XOR2 (N4732, N4730, N1432);
or OR3 (N4733, N4732, N2706, N446);
and AND4 (N4734, N4677, N2372, N3609, N3087);
xor XOR2 (N4735, N4728, N4338);
nand NAND3 (N4736, N4729, N3018, N3097);
not NOT1 (N4737, N4720);
nor NOR4 (N4738, N4709, N4635, N2366, N1791);
buf BUF1 (N4739, N4727);
or OR4 (N4740, N4738, N583, N1330, N3681);
not NOT1 (N4741, N4740);
xor XOR2 (N4742, N4734, N2364);
nor NOR3 (N4743, N4721, N502, N3387);
nor NOR4 (N4744, N4742, N3154, N3150, N1678);
buf BUF1 (N4745, N4743);
and AND2 (N4746, N4723, N1092);
or OR3 (N4747, N4746, N4288, N1445);
nor NOR2 (N4748, N4735, N969);
not NOT1 (N4749, N4736);
nand NAND2 (N4750, N4745, N3153);
xor XOR2 (N4751, N4748, N2101);
and AND3 (N4752, N4749, N151, N3184);
or OR2 (N4753, N4737, N3605);
xor XOR2 (N4754, N4753, N1461);
and AND4 (N4755, N4733, N1254, N3157, N1520);
nor NOR3 (N4756, N4731, N1897, N3962);
or OR3 (N4757, N4744, N2649, N1591);
nor NOR3 (N4758, N4757, N942, N3195);
buf BUF1 (N4759, N4752);
not NOT1 (N4760, N4756);
buf BUF1 (N4761, N4758);
or OR2 (N4762, N4739, N556);
nand NAND2 (N4763, N4754, N1569);
and AND2 (N4764, N4747, N4749);
buf BUF1 (N4765, N4762);
xor XOR2 (N4766, N4764, N597);
nand NAND4 (N4767, N4765, N3946, N2653, N4142);
not NOT1 (N4768, N4766);
xor XOR2 (N4769, N4767, N917);
xor XOR2 (N4770, N4763, N678);
nor NOR4 (N4771, N4741, N1967, N381, N1708);
nor NOR4 (N4772, N4751, N1135, N815, N455);
buf BUF1 (N4773, N4769);
not NOT1 (N4774, N4771);
and AND2 (N4775, N4772, N3112);
and AND2 (N4776, N4770, N821);
buf BUF1 (N4777, N4759);
nand NAND4 (N4778, N4773, N4586, N524, N2465);
nand NAND3 (N4779, N4755, N711, N2815);
not NOT1 (N4780, N4778);
nand NAND3 (N4781, N4761, N3960, N3619);
buf BUF1 (N4782, N4777);
nor NOR4 (N4783, N4750, N1875, N4209, N3871);
and AND3 (N4784, N4775, N1479, N1160);
not NOT1 (N4785, N4784);
and AND4 (N4786, N4780, N4310, N4311, N4110);
xor XOR2 (N4787, N4783, N3564);
buf BUF1 (N4788, N4782);
buf BUF1 (N4789, N4787);
and AND2 (N4790, N4788, N3879);
xor XOR2 (N4791, N4790, N4535);
buf BUF1 (N4792, N4789);
or OR3 (N4793, N4791, N1957, N2903);
or OR3 (N4794, N4786, N1466, N2491);
not NOT1 (N4795, N4781);
buf BUF1 (N4796, N4774);
not NOT1 (N4797, N4792);
nor NOR4 (N4798, N4793, N4537, N2638, N4755);
or OR4 (N4799, N4795, N3577, N4371, N2759);
not NOT1 (N4800, N4794);
xor XOR2 (N4801, N4796, N2509);
or OR2 (N4802, N4768, N2258);
or OR3 (N4803, N4799, N4336, N2141);
xor XOR2 (N4804, N4803, N1919);
and AND3 (N4805, N4779, N2563, N1467);
nor NOR3 (N4806, N4797, N2326, N884);
nand NAND2 (N4807, N4804, N3363);
buf BUF1 (N4808, N4798);
or OR4 (N4809, N4808, N1839, N2274, N598);
nor NOR2 (N4810, N4802, N245);
not NOT1 (N4811, N4760);
xor XOR2 (N4812, N4785, N3600);
and AND2 (N4813, N4811, N2570);
or OR3 (N4814, N4813, N520, N1298);
buf BUF1 (N4815, N4809);
buf BUF1 (N4816, N4806);
and AND3 (N4817, N4815, N3532, N1738);
nor NOR2 (N4818, N4816, N1411);
or OR2 (N4819, N4805, N3466);
nor NOR4 (N4820, N4818, N3734, N4799, N3117);
xor XOR2 (N4821, N4810, N2202);
nor NOR3 (N4822, N4819, N948, N2686);
nor NOR3 (N4823, N4807, N1090, N4181);
nand NAND2 (N4824, N4814, N825);
or OR2 (N4825, N4817, N2168);
and AND4 (N4826, N4823, N672, N3357, N4685);
not NOT1 (N4827, N4776);
nand NAND3 (N4828, N4800, N3947, N4099);
nand NAND3 (N4829, N4824, N755, N1103);
or OR4 (N4830, N4828, N1419, N2126, N3301);
xor XOR2 (N4831, N4801, N3393);
not NOT1 (N4832, N4831);
buf BUF1 (N4833, N4832);
and AND3 (N4834, N4833, N3051, N1673);
and AND4 (N4835, N4821, N1952, N1353, N4733);
xor XOR2 (N4836, N4826, N530);
buf BUF1 (N4837, N4822);
nor NOR3 (N4838, N4827, N1360, N3476);
buf BUF1 (N4839, N4825);
nand NAND2 (N4840, N4837, N4829);
buf BUF1 (N4841, N1049);
nand NAND3 (N4842, N4839, N3520, N3170);
not NOT1 (N4843, N4840);
nand NAND4 (N4844, N4834, N1115, N4069, N3309);
or OR3 (N4845, N4830, N1064, N2513);
buf BUF1 (N4846, N4843);
and AND4 (N4847, N4841, N1759, N2823, N2388);
buf BUF1 (N4848, N4842);
nand NAND3 (N4849, N4846, N2778, N2269);
nor NOR4 (N4850, N4820, N4799, N2554, N1579);
buf BUF1 (N4851, N4849);
xor XOR2 (N4852, N4812, N3764);
and AND4 (N4853, N4847, N1110, N2103, N3530);
buf BUF1 (N4854, N4848);
not NOT1 (N4855, N4851);
xor XOR2 (N4856, N4838, N2840);
not NOT1 (N4857, N4845);
and AND2 (N4858, N4853, N2882);
or OR4 (N4859, N4858, N3771, N3121, N4034);
xor XOR2 (N4860, N4850, N2939);
not NOT1 (N4861, N4844);
nand NAND3 (N4862, N4835, N3693, N1337);
and AND2 (N4863, N4852, N422);
and AND4 (N4864, N4861, N2521, N1832, N953);
buf BUF1 (N4865, N4862);
xor XOR2 (N4866, N4856, N1754);
xor XOR2 (N4867, N4866, N3908);
nand NAND3 (N4868, N4863, N286, N3877);
buf BUF1 (N4869, N4868);
not NOT1 (N4870, N4855);
nor NOR3 (N4871, N4859, N2672, N4360);
nor NOR4 (N4872, N4854, N1709, N4326, N466);
buf BUF1 (N4873, N4857);
xor XOR2 (N4874, N4871, N379);
nand NAND2 (N4875, N4870, N2532);
nor NOR2 (N4876, N4874, N1454);
nand NAND3 (N4877, N4876, N1822, N4071);
nor NOR2 (N4878, N4873, N2656);
xor XOR2 (N4879, N4836, N81);
nand NAND2 (N4880, N4877, N58);
or OR4 (N4881, N4875, N1145, N2136, N48);
or OR3 (N4882, N4879, N4271, N731);
nand NAND2 (N4883, N4881, N4749);
nand NAND2 (N4884, N4867, N2680);
and AND2 (N4885, N4872, N2627);
not NOT1 (N4886, N4880);
nor NOR4 (N4887, N4864, N4235, N1702, N4604);
buf BUF1 (N4888, N4886);
nand NAND2 (N4889, N4885, N2874);
buf BUF1 (N4890, N4887);
not NOT1 (N4891, N4888);
nor NOR4 (N4892, N4891, N3276, N4067, N600);
or OR3 (N4893, N4884, N933, N4293);
xor XOR2 (N4894, N4865, N2934);
or OR2 (N4895, N4860, N3443);
buf BUF1 (N4896, N4893);
nor NOR3 (N4897, N4896, N3279, N4259);
or OR3 (N4898, N4889, N4583, N3998);
and AND4 (N4899, N4869, N3787, N39, N2036);
xor XOR2 (N4900, N4897, N3854);
or OR4 (N4901, N4878, N920, N1072, N1712);
or OR2 (N4902, N4895, N2796);
nand NAND2 (N4903, N4898, N4065);
not NOT1 (N4904, N4902);
xor XOR2 (N4905, N4892, N3383);
buf BUF1 (N4906, N4883);
or OR2 (N4907, N4904, N4539);
buf BUF1 (N4908, N4903);
or OR4 (N4909, N4900, N3045, N3125, N3708);
nand NAND2 (N4910, N4890, N1114);
xor XOR2 (N4911, N4906, N4519);
or OR4 (N4912, N4909, N665, N4474, N4411);
or OR4 (N4913, N4908, N2564, N2957, N3447);
and AND4 (N4914, N4899, N2725, N1990, N3533);
not NOT1 (N4915, N4882);
buf BUF1 (N4916, N4915);
nand NAND4 (N4917, N4916, N3325, N4810, N4645);
buf BUF1 (N4918, N4905);
or OR2 (N4919, N4913, N4394);
buf BUF1 (N4920, N4914);
nor NOR4 (N4921, N4920, N1235, N4606, N4418);
nand NAND2 (N4922, N4912, N1657);
or OR2 (N4923, N4922, N2641);
xor XOR2 (N4924, N4894, N453);
xor XOR2 (N4925, N4919, N4168);
nor NOR4 (N4926, N4925, N3994, N3764, N1717);
or OR4 (N4927, N4923, N4755, N4182, N3735);
buf BUF1 (N4928, N4910);
xor XOR2 (N4929, N4907, N1179);
nand NAND3 (N4930, N4924, N208, N2490);
and AND4 (N4931, N4928, N2679, N4546, N3114);
or OR4 (N4932, N4926, N4061, N1088, N1401);
buf BUF1 (N4933, N4917);
not NOT1 (N4934, N4931);
nor NOR2 (N4935, N4930, N2177);
or OR2 (N4936, N4932, N3183);
not NOT1 (N4937, N4929);
and AND3 (N4938, N4936, N1289, N2321);
buf BUF1 (N4939, N4933);
or OR4 (N4940, N4918, N117, N2052, N785);
nor NOR2 (N4941, N4935, N4002);
not NOT1 (N4942, N4927);
and AND2 (N4943, N4934, N2012);
nand NAND3 (N4944, N4943, N3297, N4351);
nor NOR2 (N4945, N4911, N1182);
or OR2 (N4946, N4938, N1999);
nor NOR2 (N4947, N4901, N854);
buf BUF1 (N4948, N4940);
nor NOR3 (N4949, N4944, N1503, N4334);
buf BUF1 (N4950, N4946);
not NOT1 (N4951, N4941);
not NOT1 (N4952, N4948);
and AND4 (N4953, N4952, N287, N3179, N4922);
nor NOR2 (N4954, N4942, N3707);
or OR4 (N4955, N4950, N4911, N4718, N3954);
not NOT1 (N4956, N4945);
not NOT1 (N4957, N4954);
nor NOR3 (N4958, N4951, N1634, N3737);
xor XOR2 (N4959, N4957, N1302);
buf BUF1 (N4960, N4921);
and AND2 (N4961, N4949, N4300);
nand NAND3 (N4962, N4937, N3324, N4475);
xor XOR2 (N4963, N4962, N3466);
and AND2 (N4964, N4956, N4577);
or OR2 (N4965, N4959, N4231);
not NOT1 (N4966, N4960);
buf BUF1 (N4967, N4961);
not NOT1 (N4968, N4947);
buf BUF1 (N4969, N4967);
nand NAND2 (N4970, N4953, N3579);
xor XOR2 (N4971, N4963, N65);
xor XOR2 (N4972, N4971, N2048);
nand NAND3 (N4973, N4965, N3818, N573);
buf BUF1 (N4974, N4972);
nor NOR2 (N4975, N4969, N1874);
or OR3 (N4976, N4958, N3247, N4088);
nand NAND3 (N4977, N4964, N2292, N3434);
not NOT1 (N4978, N4973);
nor NOR2 (N4979, N4955, N1593);
nand NAND2 (N4980, N4977, N3909);
or OR2 (N4981, N4976, N2338);
or OR4 (N4982, N4975, N647, N1547, N600);
and AND2 (N4983, N4974, N3181);
buf BUF1 (N4984, N4939);
not NOT1 (N4985, N4968);
nor NOR3 (N4986, N4981, N3215, N4909);
not NOT1 (N4987, N4985);
not NOT1 (N4988, N4984);
xor XOR2 (N4989, N4966, N3002);
buf BUF1 (N4990, N4970);
buf BUF1 (N4991, N4979);
nand NAND2 (N4992, N4988, N902);
nor NOR3 (N4993, N4989, N4105, N2830);
nand NAND3 (N4994, N4980, N3515, N4147);
nand NAND4 (N4995, N4987, N4076, N3156, N1777);
not NOT1 (N4996, N4978);
nand NAND2 (N4997, N4996, N1821);
xor XOR2 (N4998, N4990, N4007);
xor XOR2 (N4999, N4983, N1177);
or OR3 (N5000, N4998, N3229, N229);
xor XOR2 (N5001, N4997, N812);
and AND4 (N5002, N4994, N4798, N2362, N2234);
and AND4 (N5003, N4991, N1330, N3694, N1739);
buf BUF1 (N5004, N5001);
xor XOR2 (N5005, N5004, N2892);
and AND2 (N5006, N4993, N2003);
nor NOR2 (N5007, N4995, N3799);
nor NOR3 (N5008, N5006, N2514, N273);
or OR4 (N5009, N5008, N1891, N87, N4254);
buf BUF1 (N5010, N5003);
or OR3 (N5011, N5010, N431, N1356);
nor NOR4 (N5012, N5002, N3928, N4041, N4472);
and AND3 (N5013, N5000, N275, N1907);
nor NOR4 (N5014, N5005, N4593, N2404, N2309);
and AND4 (N5015, N5012, N421, N1242, N1890);
not NOT1 (N5016, N4986);
xor XOR2 (N5017, N5009, N2581);
buf BUF1 (N5018, N5015);
not NOT1 (N5019, N5016);
not NOT1 (N5020, N5013);
or OR4 (N5021, N5019, N82, N4228, N496);
nor NOR3 (N5022, N5014, N2844, N3596);
nand NAND4 (N5023, N4999, N4029, N981, N3161);
not NOT1 (N5024, N5018);
nand NAND4 (N5025, N5024, N47, N4409, N4673);
nor NOR4 (N5026, N5022, N2792, N2906, N3946);
or OR3 (N5027, N5020, N3986, N1368);
nand NAND3 (N5028, N5027, N2818, N4715);
or OR4 (N5029, N5011, N1759, N953, N814);
nor NOR2 (N5030, N5026, N19);
not NOT1 (N5031, N4982);
xor XOR2 (N5032, N5025, N4200);
not NOT1 (N5033, N5029);
not NOT1 (N5034, N5007);
nand NAND2 (N5035, N5030, N368);
or OR4 (N5036, N5023, N2776, N3180, N1111);
nor NOR2 (N5037, N5033, N2693);
not NOT1 (N5038, N5017);
buf BUF1 (N5039, N5038);
or OR2 (N5040, N4992, N52);
buf BUF1 (N5041, N5036);
nand NAND3 (N5042, N5040, N1299, N459);
not NOT1 (N5043, N5037);
nor NOR2 (N5044, N5043, N449);
not NOT1 (N5045, N5034);
buf BUF1 (N5046, N5035);
not NOT1 (N5047, N5045);
buf BUF1 (N5048, N5039);
nor NOR2 (N5049, N5047, N3384);
or OR2 (N5050, N5044, N3278);
nor NOR4 (N5051, N5041, N4991, N1336, N2758);
nand NAND4 (N5052, N5042, N2081, N4775, N848);
not NOT1 (N5053, N5048);
nor NOR4 (N5054, N5031, N1024, N2847, N785);
nor NOR2 (N5055, N5049, N4915);
not NOT1 (N5056, N5028);
and AND4 (N5057, N5032, N2327, N1515, N3685);
nor NOR4 (N5058, N5054, N4882, N3939, N4292);
buf BUF1 (N5059, N5058);
xor XOR2 (N5060, N5053, N246);
buf BUF1 (N5061, N5050);
nor NOR3 (N5062, N5059, N3430, N3769);
or OR3 (N5063, N5057, N4065, N2884);
buf BUF1 (N5064, N5060);
xor XOR2 (N5065, N5063, N1087);
and AND2 (N5066, N5062, N4283);
or OR3 (N5067, N5021, N2021, N1584);
xor XOR2 (N5068, N5051, N3864);
buf BUF1 (N5069, N5065);
buf BUF1 (N5070, N5046);
or OR3 (N5071, N5061, N1506, N1422);
nand NAND2 (N5072, N5067, N2777);
and AND2 (N5073, N5069, N4745);
or OR2 (N5074, N5066, N1166);
and AND2 (N5075, N5064, N2564);
and AND4 (N5076, N5074, N3393, N4747, N4153);
buf BUF1 (N5077, N5076);
and AND4 (N5078, N5070, N3347, N2490, N3698);
nor NOR3 (N5079, N5068, N2603, N1849);
nor NOR4 (N5080, N5055, N3498, N313, N2916);
xor XOR2 (N5081, N5079, N5050);
nor NOR2 (N5082, N5071, N1791);
and AND2 (N5083, N5077, N4819);
nor NOR4 (N5084, N5083, N1267, N1133, N4651);
xor XOR2 (N5085, N5056, N1418);
not NOT1 (N5086, N5080);
not NOT1 (N5087, N5075);
or OR3 (N5088, N5085, N3, N3320);
nand NAND2 (N5089, N5073, N1916);
not NOT1 (N5090, N5082);
not NOT1 (N5091, N5084);
or OR2 (N5092, N5078, N4403);
not NOT1 (N5093, N5090);
xor XOR2 (N5094, N5086, N4546);
and AND4 (N5095, N5091, N61, N2637, N4673);
or OR3 (N5096, N5081, N415, N4243);
buf BUF1 (N5097, N5087);
not NOT1 (N5098, N5093);
nand NAND2 (N5099, N5092, N2818);
nand NAND2 (N5100, N5096, N3288);
nand NAND4 (N5101, N5052, N1328, N613, N1225);
or OR4 (N5102, N5094, N1813, N520, N1806);
buf BUF1 (N5103, N5072);
buf BUF1 (N5104, N5100);
nor NOR2 (N5105, N5098, N4639);
and AND2 (N5106, N5104, N2051);
nand NAND3 (N5107, N5099, N3496, N4036);
buf BUF1 (N5108, N5095);
and AND3 (N5109, N5102, N3181, N2077);
and AND3 (N5110, N5105, N494, N1029);
nor NOR4 (N5111, N5107, N2360, N3979, N2004);
and AND2 (N5112, N5101, N796);
xor XOR2 (N5113, N5110, N4440);
not NOT1 (N5114, N5112);
xor XOR2 (N5115, N5108, N1753);
or OR4 (N5116, N5097, N1765, N105, N2057);
or OR3 (N5117, N5115, N3204, N2101);
nand NAND4 (N5118, N5117, N2579, N2238, N4001);
nor NOR2 (N5119, N5113, N1713);
nand NAND4 (N5120, N5119, N4078, N4396, N2371);
buf BUF1 (N5121, N5114);
nand NAND2 (N5122, N5118, N1725);
nand NAND3 (N5123, N5120, N2392, N3379);
nor NOR2 (N5124, N5109, N4678);
or OR2 (N5125, N5122, N1413);
buf BUF1 (N5126, N5121);
nand NAND3 (N5127, N5123, N4181, N3859);
nand NAND2 (N5128, N5116, N4433);
buf BUF1 (N5129, N5111);
buf BUF1 (N5130, N5129);
buf BUF1 (N5131, N5103);
not NOT1 (N5132, N5128);
or OR3 (N5133, N5130, N3121, N91);
and AND2 (N5134, N5127, N3877);
and AND3 (N5135, N5125, N708, N3276);
and AND3 (N5136, N5135, N4201, N2688);
or OR3 (N5137, N5106, N3596, N3657);
not NOT1 (N5138, N5126);
nor NOR4 (N5139, N5131, N4708, N2690, N2732);
xor XOR2 (N5140, N5133, N4769);
nand NAND4 (N5141, N5139, N4418, N2965, N3645);
not NOT1 (N5142, N5132);
xor XOR2 (N5143, N5136, N5087);
nor NOR4 (N5144, N5143, N3339, N2354, N3099);
buf BUF1 (N5145, N5088);
or OR2 (N5146, N5089, N1936);
nand NAND3 (N5147, N5142, N4517, N3125);
nor NOR4 (N5148, N5145, N2113, N3476, N1788);
xor XOR2 (N5149, N5147, N2620);
nand NAND4 (N5150, N5146, N35, N4510, N3838);
nor NOR2 (N5151, N5137, N4605);
or OR2 (N5152, N5144, N2416);
not NOT1 (N5153, N5148);
and AND3 (N5154, N5149, N1985, N4171);
not NOT1 (N5155, N5140);
buf BUF1 (N5156, N5153);
buf BUF1 (N5157, N5154);
not NOT1 (N5158, N5152);
or OR3 (N5159, N5158, N4813, N44);
xor XOR2 (N5160, N5155, N1736);
xor XOR2 (N5161, N5141, N1406);
xor XOR2 (N5162, N5124, N1842);
xor XOR2 (N5163, N5134, N959);
not NOT1 (N5164, N5157);
nor NOR2 (N5165, N5161, N2736);
not NOT1 (N5166, N5162);
or OR2 (N5167, N5163, N5075);
nand NAND3 (N5168, N5164, N3688, N2857);
xor XOR2 (N5169, N5165, N1419);
not NOT1 (N5170, N5168);
and AND3 (N5171, N5170, N3839, N447);
nor NOR4 (N5172, N5138, N1227, N1277, N888);
nor NOR4 (N5173, N5156, N232, N2246, N3117);
xor XOR2 (N5174, N5166, N5024);
not NOT1 (N5175, N5167);
nand NAND3 (N5176, N5159, N1929, N1832);
or OR2 (N5177, N5151, N3537);
nor NOR3 (N5178, N5174, N2178, N4970);
nor NOR3 (N5179, N5160, N3927, N2697);
nand NAND4 (N5180, N5177, N215, N2923, N4593);
not NOT1 (N5181, N5178);
nand NAND3 (N5182, N5180, N3805, N5169);
not NOT1 (N5183, N2611);
buf BUF1 (N5184, N5172);
xor XOR2 (N5185, N5184, N1321);
not NOT1 (N5186, N5182);
not NOT1 (N5187, N5171);
not NOT1 (N5188, N5179);
buf BUF1 (N5189, N5187);
or OR2 (N5190, N5186, N4977);
xor XOR2 (N5191, N5173, N2892);
not NOT1 (N5192, N5189);
nor NOR2 (N5193, N5175, N794);
xor XOR2 (N5194, N5176, N3055);
and AND4 (N5195, N5190, N1195, N2984, N3272);
nor NOR4 (N5196, N5183, N1211, N3643, N40);
xor XOR2 (N5197, N5191, N3509);
buf BUF1 (N5198, N5195);
nor NOR2 (N5199, N5188, N2736);
nand NAND3 (N5200, N5196, N560, N1179);
not NOT1 (N5201, N5181);
nor NOR2 (N5202, N5197, N1398);
nand NAND4 (N5203, N5150, N1939, N4649, N4428);
or OR4 (N5204, N5200, N4991, N3868, N4830);
or OR4 (N5205, N5201, N2183, N688, N4818);
nand NAND4 (N5206, N5202, N3348, N211, N4637);
nand NAND4 (N5207, N5206, N53, N666, N2667);
xor XOR2 (N5208, N5207, N4009);
nand NAND3 (N5209, N5208, N4018, N4396);
and AND4 (N5210, N5194, N5179, N2263, N3577);
not NOT1 (N5211, N5203);
not NOT1 (N5212, N5192);
nor NOR4 (N5213, N5204, N2854, N4243, N701);
nand NAND4 (N5214, N5211, N4113, N216, N625);
nand NAND4 (N5215, N5212, N2530, N652, N4544);
buf BUF1 (N5216, N5185);
buf BUF1 (N5217, N5214);
not NOT1 (N5218, N5210);
nand NAND2 (N5219, N5216, N1258);
nand NAND3 (N5220, N5198, N4539, N1535);
and AND4 (N5221, N5213, N4674, N4953, N2091);
and AND3 (N5222, N5209, N1658, N160);
buf BUF1 (N5223, N5205);
xor XOR2 (N5224, N5217, N3112);
nand NAND3 (N5225, N5223, N2603, N2418);
not NOT1 (N5226, N5225);
buf BUF1 (N5227, N5220);
buf BUF1 (N5228, N5193);
not NOT1 (N5229, N5224);
not NOT1 (N5230, N5227);
xor XOR2 (N5231, N5218, N1789);
xor XOR2 (N5232, N5231, N931);
or OR4 (N5233, N5230, N2637, N3538, N4790);
nand NAND3 (N5234, N5215, N3435, N4372);
and AND2 (N5235, N5226, N1090);
and AND2 (N5236, N5219, N4300);
not NOT1 (N5237, N5199);
nor NOR4 (N5238, N5222, N4964, N1845, N2214);
nand NAND3 (N5239, N5237, N3439, N4092);
and AND3 (N5240, N5235, N1952, N3629);
buf BUF1 (N5241, N5228);
or OR4 (N5242, N5239, N1782, N4868, N1514);
xor XOR2 (N5243, N5229, N4950);
buf BUF1 (N5244, N5232);
not NOT1 (N5245, N5238);
buf BUF1 (N5246, N5242);
and AND2 (N5247, N5236, N252);
not NOT1 (N5248, N5245);
or OR2 (N5249, N5248, N773);
nand NAND2 (N5250, N5246, N1764);
not NOT1 (N5251, N5241);
nand NAND3 (N5252, N5221, N2890, N1247);
buf BUF1 (N5253, N5247);
or OR4 (N5254, N5251, N4832, N4770, N3830);
nor NOR2 (N5255, N5240, N40);
xor XOR2 (N5256, N5250, N3848);
buf BUF1 (N5257, N5249);
nor NOR3 (N5258, N5254, N4970, N2110);
and AND4 (N5259, N5234, N2097, N1249, N4163);
nand NAND3 (N5260, N5244, N5089, N3476);
or OR3 (N5261, N5233, N3608, N5254);
buf BUF1 (N5262, N5243);
not NOT1 (N5263, N5253);
xor XOR2 (N5264, N5259, N1348);
nand NAND3 (N5265, N5258, N2226, N2130);
buf BUF1 (N5266, N5257);
nor NOR4 (N5267, N5264, N1919, N5069, N3750);
and AND4 (N5268, N5263, N292, N3633, N1963);
buf BUF1 (N5269, N5267);
nand NAND3 (N5270, N5255, N145, N4643);
not NOT1 (N5271, N5265);
nand NAND3 (N5272, N5261, N751, N2698);
and AND2 (N5273, N5269, N5135);
buf BUF1 (N5274, N5266);
or OR4 (N5275, N5252, N4759, N4130, N5188);
and AND3 (N5276, N5274, N2700, N1528);
xor XOR2 (N5277, N5262, N3177);
not NOT1 (N5278, N5256);
nor NOR2 (N5279, N5268, N399);
xor XOR2 (N5280, N5279, N3182);
nand NAND2 (N5281, N5280, N2884);
buf BUF1 (N5282, N5271);
xor XOR2 (N5283, N5278, N1370);
nor NOR3 (N5284, N5260, N2784, N364);
buf BUF1 (N5285, N5273);
or OR2 (N5286, N5285, N2479);
not NOT1 (N5287, N5286);
xor XOR2 (N5288, N5276, N2178);
buf BUF1 (N5289, N5272);
nand NAND4 (N5290, N5275, N4086, N5157, N238);
nand NAND3 (N5291, N5290, N3448, N3477);
nor NOR4 (N5292, N5277, N4140, N3827, N1199);
xor XOR2 (N5293, N5291, N3595);
nor NOR4 (N5294, N5293, N3338, N679, N3460);
not NOT1 (N5295, N5294);
xor XOR2 (N5296, N5282, N5112);
nor NOR2 (N5297, N5289, N2743);
buf BUF1 (N5298, N5287);
or OR3 (N5299, N5283, N380, N2648);
xor XOR2 (N5300, N5299, N5176);
not NOT1 (N5301, N5297);
nor NOR3 (N5302, N5298, N3439, N431);
or OR2 (N5303, N5270, N4227);
buf BUF1 (N5304, N5281);
or OR3 (N5305, N5295, N3529, N3319);
or OR2 (N5306, N5284, N4635);
and AND3 (N5307, N5301, N4914, N957);
not NOT1 (N5308, N5288);
nor NOR2 (N5309, N5302, N939);
and AND2 (N5310, N5308, N4895);
or OR4 (N5311, N5307, N3497, N3227, N4082);
nand NAND3 (N5312, N5304, N1573, N3986);
not NOT1 (N5313, N5305);
not NOT1 (N5314, N5300);
not NOT1 (N5315, N5296);
and AND2 (N5316, N5292, N449);
not NOT1 (N5317, N5306);
and AND2 (N5318, N5316, N206);
nand NAND3 (N5319, N5312, N5178, N3952);
nand NAND2 (N5320, N5309, N1522);
buf BUF1 (N5321, N5311);
not NOT1 (N5322, N5310);
nor NOR3 (N5323, N5315, N3490, N1494);
or OR2 (N5324, N5320, N1846);
and AND3 (N5325, N5322, N1413, N2873);
or OR3 (N5326, N5325, N1699, N2626);
not NOT1 (N5327, N5317);
xor XOR2 (N5328, N5318, N1338);
nand NAND2 (N5329, N5324, N1110);
and AND4 (N5330, N5327, N3089, N721, N4551);
nand NAND4 (N5331, N5321, N4603, N1634, N2129);
buf BUF1 (N5332, N5330);
not NOT1 (N5333, N5323);
buf BUF1 (N5334, N5313);
or OR4 (N5335, N5329, N592, N4338, N4410);
not NOT1 (N5336, N5303);
and AND4 (N5337, N5332, N3069, N3843, N3379);
buf BUF1 (N5338, N5335);
xor XOR2 (N5339, N5326, N3262);
nand NAND2 (N5340, N5338, N2160);
nand NAND4 (N5341, N5314, N551, N614, N3652);
xor XOR2 (N5342, N5333, N2754);
nor NOR3 (N5343, N5331, N784, N4227);
xor XOR2 (N5344, N5341, N82);
not NOT1 (N5345, N5337);
buf BUF1 (N5346, N5345);
nand NAND4 (N5347, N5344, N266, N4825, N584);
and AND4 (N5348, N5319, N627, N92, N249);
and AND4 (N5349, N5339, N3264, N3672, N2165);
buf BUF1 (N5350, N5340);
or OR2 (N5351, N5334, N1891);
nand NAND4 (N5352, N5336, N913, N3317, N5328);
not NOT1 (N5353, N319);
buf BUF1 (N5354, N5350);
not NOT1 (N5355, N5343);
and AND2 (N5356, N5346, N1935);
nand NAND4 (N5357, N5354, N2508, N5206, N3274);
nor NOR2 (N5358, N5357, N4627);
and AND2 (N5359, N5353, N833);
and AND2 (N5360, N5348, N4853);
nor NOR4 (N5361, N5356, N4374, N3803, N1935);
xor XOR2 (N5362, N5352, N2134);
not NOT1 (N5363, N5351);
nor NOR3 (N5364, N5342, N3941, N165);
nor NOR4 (N5365, N5349, N1438, N1911, N2674);
and AND3 (N5366, N5358, N105, N2530);
nand NAND3 (N5367, N5361, N3519, N1802);
or OR2 (N5368, N5364, N4769);
nor NOR2 (N5369, N5362, N23);
nand NAND4 (N5370, N5365, N4841, N525, N1821);
and AND3 (N5371, N5363, N1614, N3265);
nor NOR2 (N5372, N5367, N1300);
not NOT1 (N5373, N5371);
not NOT1 (N5374, N5355);
not NOT1 (N5375, N5372);
buf BUF1 (N5376, N5373);
nor NOR2 (N5377, N5369, N5041);
and AND2 (N5378, N5374, N800);
xor XOR2 (N5379, N5378, N2945);
buf BUF1 (N5380, N5366);
not NOT1 (N5381, N5380);
xor XOR2 (N5382, N5370, N4043);
xor XOR2 (N5383, N5376, N1302);
buf BUF1 (N5384, N5383);
nand NAND4 (N5385, N5375, N246, N4126, N2130);
nand NAND2 (N5386, N5377, N5384);
and AND3 (N5387, N798, N1341, N3116);
xor XOR2 (N5388, N5382, N4672);
nand NAND3 (N5389, N5388, N1079, N3141);
nor NOR3 (N5390, N5368, N2312, N4411);
nand NAND3 (N5391, N5389, N1120, N427);
nand NAND2 (N5392, N5379, N1472);
nand NAND4 (N5393, N5387, N1673, N2132, N1196);
xor XOR2 (N5394, N5347, N2529);
buf BUF1 (N5395, N5390);
not NOT1 (N5396, N5393);
nand NAND4 (N5397, N5386, N1753, N4069, N2490);
xor XOR2 (N5398, N5359, N4404);
buf BUF1 (N5399, N5398);
not NOT1 (N5400, N5391);
buf BUF1 (N5401, N5397);
nor NOR4 (N5402, N5395, N5236, N1262, N1803);
and AND4 (N5403, N5385, N1700, N4018, N4137);
not NOT1 (N5404, N5400);
nor NOR2 (N5405, N5381, N2196);
buf BUF1 (N5406, N5399);
nand NAND2 (N5407, N5401, N407);
nand NAND3 (N5408, N5403, N729, N2752);
or OR2 (N5409, N5394, N1781);
or OR3 (N5410, N5404, N4135, N1603);
buf BUF1 (N5411, N5392);
buf BUF1 (N5412, N5402);
xor XOR2 (N5413, N5406, N3397);
nand NAND2 (N5414, N5409, N1607);
nand NAND2 (N5415, N5408, N2642);
xor XOR2 (N5416, N5396, N920);
not NOT1 (N5417, N5407);
buf BUF1 (N5418, N5416);
and AND2 (N5419, N5415, N4387);
nand NAND4 (N5420, N5414, N2164, N990, N3699);
xor XOR2 (N5421, N5419, N3855);
nand NAND3 (N5422, N5418, N5382, N1134);
not NOT1 (N5423, N5417);
or OR2 (N5424, N5360, N3117);
xor XOR2 (N5425, N5411, N362);
xor XOR2 (N5426, N5422, N3740);
xor XOR2 (N5427, N5413, N901);
nor NOR4 (N5428, N5423, N1878, N414, N2699);
nand NAND2 (N5429, N5421, N5263);
nor NOR4 (N5430, N5420, N4471, N573, N980);
xor XOR2 (N5431, N5429, N151);
xor XOR2 (N5432, N5430, N3006);
or OR3 (N5433, N5426, N5026, N1749);
not NOT1 (N5434, N5433);
nand NAND2 (N5435, N5425, N209);
buf BUF1 (N5436, N5427);
or OR2 (N5437, N5405, N54);
and AND2 (N5438, N5436, N244);
nand NAND3 (N5439, N5434, N3218, N1130);
and AND3 (N5440, N5435, N1200, N4900);
or OR3 (N5441, N5431, N3277, N108);
nor NOR2 (N5442, N5424, N1705);
xor XOR2 (N5443, N5438, N505);
nor NOR3 (N5444, N5412, N2477, N1318);
buf BUF1 (N5445, N5428);
not NOT1 (N5446, N5439);
nor NOR4 (N5447, N5432, N2270, N1579, N1284);
xor XOR2 (N5448, N5443, N495);
nor NOR2 (N5449, N5445, N2068);
buf BUF1 (N5450, N5447);
xor XOR2 (N5451, N5442, N2248);
or OR2 (N5452, N5450, N1153);
buf BUF1 (N5453, N5449);
or OR2 (N5454, N5444, N3297);
and AND3 (N5455, N5448, N2059, N187);
xor XOR2 (N5456, N5441, N2310);
nand NAND2 (N5457, N5455, N1310);
or OR2 (N5458, N5437, N48);
xor XOR2 (N5459, N5440, N3944);
nand NAND3 (N5460, N5456, N1493, N686);
xor XOR2 (N5461, N5460, N1860);
or OR2 (N5462, N5461, N3668);
nor NOR3 (N5463, N5451, N2383, N2160);
nor NOR3 (N5464, N5453, N2699, N1345);
not NOT1 (N5465, N5463);
nand NAND2 (N5466, N5464, N3364);
not NOT1 (N5467, N5462);
nand NAND2 (N5468, N5458, N3933);
nand NAND3 (N5469, N5468, N1298, N50);
and AND2 (N5470, N5446, N4200);
nand NAND3 (N5471, N5459, N4690, N1999);
buf BUF1 (N5472, N5470);
nor NOR2 (N5473, N5452, N825);
nand NAND3 (N5474, N5471, N867, N1165);
xor XOR2 (N5475, N5465, N4174);
xor XOR2 (N5476, N5454, N3599);
xor XOR2 (N5477, N5476, N2784);
xor XOR2 (N5478, N5474, N3416);
xor XOR2 (N5479, N5472, N4152);
not NOT1 (N5480, N5479);
not NOT1 (N5481, N5480);
buf BUF1 (N5482, N5477);
buf BUF1 (N5483, N5466);
xor XOR2 (N5484, N5483, N1554);
or OR2 (N5485, N5469, N2266);
not NOT1 (N5486, N5485);
or OR3 (N5487, N5457, N1171, N1963);
not NOT1 (N5488, N5478);
and AND4 (N5489, N5473, N2135, N4622, N3804);
not NOT1 (N5490, N5484);
and AND3 (N5491, N5481, N1752, N2901);
and AND3 (N5492, N5487, N4794, N1742);
or OR3 (N5493, N5482, N1068, N1415);
nand NAND4 (N5494, N5467, N388, N252, N1650);
not NOT1 (N5495, N5491);
not NOT1 (N5496, N5493);
nor NOR2 (N5497, N5496, N924);
xor XOR2 (N5498, N5497, N352);
not NOT1 (N5499, N5492);
buf BUF1 (N5500, N5498);
xor XOR2 (N5501, N5500, N4250);
or OR2 (N5502, N5494, N1919);
and AND2 (N5503, N5475, N3286);
xor XOR2 (N5504, N5486, N2209);
xor XOR2 (N5505, N5490, N2618);
not NOT1 (N5506, N5410);
or OR2 (N5507, N5501, N3124);
or OR3 (N5508, N5488, N103, N1253);
buf BUF1 (N5509, N5508);
buf BUF1 (N5510, N5499);
xor XOR2 (N5511, N5502, N1913);
xor XOR2 (N5512, N5507, N1064);
not NOT1 (N5513, N5509);
or OR4 (N5514, N5505, N1123, N2623, N5111);
buf BUF1 (N5515, N5506);
and AND2 (N5516, N5513, N868);
buf BUF1 (N5517, N5489);
nor NOR4 (N5518, N5511, N240, N3065, N797);
buf BUF1 (N5519, N5504);
and AND4 (N5520, N5518, N274, N4820, N4459);
xor XOR2 (N5521, N5516, N4006);
nor NOR3 (N5522, N5512, N1343, N5066);
nand NAND3 (N5523, N5521, N5432, N3622);
not NOT1 (N5524, N5522);
not NOT1 (N5525, N5495);
nor NOR2 (N5526, N5523, N4866);
and AND2 (N5527, N5514, N88);
buf BUF1 (N5528, N5519);
buf BUF1 (N5529, N5524);
xor XOR2 (N5530, N5526, N4992);
buf BUF1 (N5531, N5529);
xor XOR2 (N5532, N5530, N5001);
nand NAND4 (N5533, N5517, N5281, N36, N1745);
not NOT1 (N5534, N5503);
nand NAND3 (N5535, N5510, N1448, N1067);
buf BUF1 (N5536, N5535);
nand NAND3 (N5537, N5533, N3264, N2389);
nor NOR3 (N5538, N5528, N1042, N4292);
and AND3 (N5539, N5515, N3662, N5187);
nor NOR2 (N5540, N5537, N680);
not NOT1 (N5541, N5525);
buf BUF1 (N5542, N5539);
nand NAND3 (N5543, N5532, N1750, N5011);
not NOT1 (N5544, N5531);
or OR3 (N5545, N5544, N3769, N3286);
and AND4 (N5546, N5540, N2048, N1659, N1213);
not NOT1 (N5547, N5534);
buf BUF1 (N5548, N5543);
or OR4 (N5549, N5536, N5475, N979, N175);
or OR2 (N5550, N5527, N211);
buf BUF1 (N5551, N5542);
nand NAND4 (N5552, N5546, N4302, N1562, N4113);
not NOT1 (N5553, N5520);
buf BUF1 (N5554, N5549);
not NOT1 (N5555, N5541);
not NOT1 (N5556, N5552);
buf BUF1 (N5557, N5548);
nor NOR4 (N5558, N5551, N4484, N3064, N5060);
or OR4 (N5559, N5545, N2202, N4432, N1080);
or OR2 (N5560, N5558, N61);
nand NAND4 (N5561, N5560, N3541, N780, N4070);
and AND2 (N5562, N5547, N3963);
not NOT1 (N5563, N5538);
buf BUF1 (N5564, N5554);
buf BUF1 (N5565, N5564);
xor XOR2 (N5566, N5550, N1510);
buf BUF1 (N5567, N5555);
buf BUF1 (N5568, N5562);
not NOT1 (N5569, N5568);
not NOT1 (N5570, N5566);
nor NOR2 (N5571, N5561, N4403);
and AND3 (N5572, N5565, N5133, N4199);
xor XOR2 (N5573, N5563, N3537);
nor NOR4 (N5574, N5567, N2324, N1401, N4730);
buf BUF1 (N5575, N5556);
nor NOR3 (N5576, N5575, N2986, N3847);
xor XOR2 (N5577, N5557, N1748);
xor XOR2 (N5578, N5570, N1606);
xor XOR2 (N5579, N5577, N4722);
nor NOR2 (N5580, N5578, N1121);
or OR2 (N5581, N5580, N3175);
not NOT1 (N5582, N5572);
and AND3 (N5583, N5574, N911, N3933);
and AND4 (N5584, N5573, N1519, N4068, N5252);
nand NAND2 (N5585, N5582, N3483);
nor NOR4 (N5586, N5569, N80, N2947, N4555);
xor XOR2 (N5587, N5559, N3255);
not NOT1 (N5588, N5584);
not NOT1 (N5589, N5579);
buf BUF1 (N5590, N5585);
and AND3 (N5591, N5553, N1756, N3256);
nand NAND3 (N5592, N5590, N3763, N3813);
nor NOR2 (N5593, N5576, N2225);
not NOT1 (N5594, N5586);
nand NAND2 (N5595, N5589, N5001);
buf BUF1 (N5596, N5571);
not NOT1 (N5597, N5583);
nand NAND4 (N5598, N5597, N1937, N1351, N1409);
xor XOR2 (N5599, N5581, N4029);
nor NOR2 (N5600, N5595, N1306);
not NOT1 (N5601, N5593);
xor XOR2 (N5602, N5588, N3824);
not NOT1 (N5603, N5602);
or OR2 (N5604, N5591, N4376);
xor XOR2 (N5605, N5592, N984);
not NOT1 (N5606, N5603);
nor NOR3 (N5607, N5596, N2031, N4570);
nor NOR4 (N5608, N5605, N1799, N187, N1541);
nor NOR4 (N5609, N5587, N4397, N433, N4998);
or OR2 (N5610, N5606, N1804);
nand NAND2 (N5611, N5607, N1587);
and AND4 (N5612, N5610, N3474, N4497, N3169);
not NOT1 (N5613, N5601);
or OR2 (N5614, N5599, N4668);
nor NOR4 (N5615, N5608, N4203, N3142, N1811);
nor NOR4 (N5616, N5615, N4971, N1736, N3595);
nand NAND4 (N5617, N5612, N2568, N5552, N2748);
and AND4 (N5618, N5616, N3766, N2382, N244);
not NOT1 (N5619, N5613);
xor XOR2 (N5620, N5598, N2979);
xor XOR2 (N5621, N5619, N2156);
buf BUF1 (N5622, N5618);
nor NOR3 (N5623, N5604, N3416, N160);
xor XOR2 (N5624, N5609, N3095);
not NOT1 (N5625, N5614);
xor XOR2 (N5626, N5594, N892);
not NOT1 (N5627, N5625);
not NOT1 (N5628, N5611);
xor XOR2 (N5629, N5622, N2135);
xor XOR2 (N5630, N5623, N308);
not NOT1 (N5631, N5621);
buf BUF1 (N5632, N5627);
or OR2 (N5633, N5626, N4738);
xor XOR2 (N5634, N5633, N914);
nand NAND3 (N5635, N5632, N3172, N1994);
nand NAND3 (N5636, N5630, N376, N2751);
or OR4 (N5637, N5636, N711, N1990, N5097);
or OR4 (N5638, N5629, N2646, N4525, N3401);
nor NOR4 (N5639, N5637, N1663, N4860, N533);
and AND4 (N5640, N5634, N3966, N3176, N742);
xor XOR2 (N5641, N5639, N3148);
xor XOR2 (N5642, N5617, N1233);
not NOT1 (N5643, N5640);
and AND3 (N5644, N5642, N4367, N2964);
or OR4 (N5645, N5644, N4879, N5085, N558);
and AND3 (N5646, N5638, N3192, N3589);
or OR2 (N5647, N5628, N1767);
nand NAND3 (N5648, N5631, N1054, N1166);
or OR4 (N5649, N5645, N982, N4851, N61);
nand NAND4 (N5650, N5643, N3499, N3934, N1321);
buf BUF1 (N5651, N5635);
nor NOR4 (N5652, N5641, N1851, N3387, N2630);
buf BUF1 (N5653, N5649);
nand NAND2 (N5654, N5651, N3605);
xor XOR2 (N5655, N5648, N2052);
or OR4 (N5656, N5647, N1626, N5341, N1515);
or OR4 (N5657, N5646, N4952, N631, N2416);
or OR2 (N5658, N5654, N2546);
nand NAND4 (N5659, N5657, N4438, N665, N3342);
nor NOR2 (N5660, N5658, N2507);
xor XOR2 (N5661, N5659, N5450);
xor XOR2 (N5662, N5653, N1204);
nand NAND3 (N5663, N5655, N93, N515);
xor XOR2 (N5664, N5661, N1773);
xor XOR2 (N5665, N5624, N3962);
nor NOR4 (N5666, N5660, N2124, N5129, N2236);
and AND3 (N5667, N5656, N2889, N3668);
not NOT1 (N5668, N5652);
and AND3 (N5669, N5650, N5254, N964);
xor XOR2 (N5670, N5666, N5523);
nor NOR2 (N5671, N5620, N957);
or OR3 (N5672, N5663, N866, N2025);
and AND4 (N5673, N5669, N402, N2888, N4139);
or OR2 (N5674, N5673, N109);
xor XOR2 (N5675, N5667, N4885);
xor XOR2 (N5676, N5600, N129);
nor NOR3 (N5677, N5672, N1905, N1206);
not NOT1 (N5678, N5674);
and AND3 (N5679, N5678, N1312, N4485);
xor XOR2 (N5680, N5675, N1202);
nand NAND4 (N5681, N5680, N4667, N2438, N5429);
and AND3 (N5682, N5668, N1865, N3867);
not NOT1 (N5683, N5679);
xor XOR2 (N5684, N5665, N250);
nand NAND4 (N5685, N5671, N877, N4165, N3009);
not NOT1 (N5686, N5682);
xor XOR2 (N5687, N5670, N5254);
nand NAND2 (N5688, N5684, N4680);
not NOT1 (N5689, N5676);
xor XOR2 (N5690, N5662, N4828);
nand NAND2 (N5691, N5686, N3885);
not NOT1 (N5692, N5690);
xor XOR2 (N5693, N5688, N5367);
not NOT1 (N5694, N5677);
xor XOR2 (N5695, N5687, N1954);
xor XOR2 (N5696, N5694, N2567);
buf BUF1 (N5697, N5692);
nand NAND2 (N5698, N5696, N4302);
not NOT1 (N5699, N5693);
and AND3 (N5700, N5681, N384, N736);
and AND3 (N5701, N5691, N1314, N8);
or OR3 (N5702, N5698, N2699, N5163);
and AND3 (N5703, N5697, N339, N2562);
xor XOR2 (N5704, N5685, N580);
and AND3 (N5705, N5695, N2781, N4523);
nor NOR3 (N5706, N5703, N351, N806);
nand NAND4 (N5707, N5683, N2579, N1184, N4210);
nand NAND2 (N5708, N5664, N2724);
xor XOR2 (N5709, N5702, N4968);
and AND4 (N5710, N5707, N3544, N5101, N2448);
buf BUF1 (N5711, N5710);
or OR2 (N5712, N5709, N2769);
nor NOR3 (N5713, N5701, N3710, N3900);
or OR4 (N5714, N5700, N2321, N4135, N2930);
not NOT1 (N5715, N5704);
nand NAND4 (N5716, N5706, N4020, N56, N921);
nand NAND2 (N5717, N5689, N487);
or OR2 (N5718, N5717, N2188);
nor NOR3 (N5719, N5712, N1306, N4922);
and AND2 (N5720, N5714, N875);
buf BUF1 (N5721, N5718);
xor XOR2 (N5722, N5711, N5449);
or OR4 (N5723, N5719, N424, N4241, N3367);
nand NAND4 (N5724, N5715, N2531, N1907, N2745);
or OR2 (N5725, N5705, N3663);
and AND4 (N5726, N5724, N886, N2595, N512);
buf BUF1 (N5727, N5722);
xor XOR2 (N5728, N5723, N4919);
nand NAND3 (N5729, N5699, N3198, N3306);
nand NAND4 (N5730, N5726, N1133, N469, N391);
buf BUF1 (N5731, N5716);
and AND4 (N5732, N5729, N297, N3593, N992);
xor XOR2 (N5733, N5708, N3626);
buf BUF1 (N5734, N5727);
nor NOR2 (N5735, N5721, N18);
xor XOR2 (N5736, N5713, N2783);
xor XOR2 (N5737, N5734, N1476);
and AND3 (N5738, N5735, N1068, N695);
buf BUF1 (N5739, N5736);
or OR4 (N5740, N5737, N2902, N4898, N2012);
xor XOR2 (N5741, N5739, N583);
and AND4 (N5742, N5740, N3409, N572, N487);
nand NAND3 (N5743, N5742, N2105, N3848);
and AND3 (N5744, N5720, N20, N4465);
xor XOR2 (N5745, N5741, N4353);
xor XOR2 (N5746, N5738, N545);
buf BUF1 (N5747, N5728);
not NOT1 (N5748, N5733);
not NOT1 (N5749, N5731);
or OR2 (N5750, N5748, N3561);
buf BUF1 (N5751, N5732);
nor NOR4 (N5752, N5730, N4631, N1075, N5267);
nor NOR4 (N5753, N5746, N3218, N1722, N4998);
or OR4 (N5754, N5751, N4055, N1257, N3365);
nor NOR2 (N5755, N5754, N1441);
xor XOR2 (N5756, N5744, N4209);
nor NOR2 (N5757, N5743, N2520);
and AND3 (N5758, N5747, N4813, N3592);
and AND4 (N5759, N5757, N2828, N1511, N3277);
and AND4 (N5760, N5756, N2695, N4918, N1588);
buf BUF1 (N5761, N5758);
not NOT1 (N5762, N5749);
xor XOR2 (N5763, N5762, N3449);
and AND4 (N5764, N5725, N2751, N5412, N5029);
not NOT1 (N5765, N5750);
nand NAND3 (N5766, N5755, N3192, N2703);
and AND4 (N5767, N5752, N3545, N5585, N26);
buf BUF1 (N5768, N5767);
buf BUF1 (N5769, N5766);
and AND2 (N5770, N5761, N5306);
xor XOR2 (N5771, N5768, N115);
or OR4 (N5772, N5753, N813, N5096, N1336);
nor NOR4 (N5773, N5765, N3714, N4237, N3369);
buf BUF1 (N5774, N5769);
xor XOR2 (N5775, N5745, N809);
buf BUF1 (N5776, N5771);
xor XOR2 (N5777, N5772, N5239);
or OR4 (N5778, N5764, N625, N4175, N3310);
nor NOR2 (N5779, N5770, N5177);
not NOT1 (N5780, N5777);
xor XOR2 (N5781, N5774, N3636);
buf BUF1 (N5782, N5775);
nand NAND3 (N5783, N5781, N2589, N2150);
and AND2 (N5784, N5778, N3443);
or OR2 (N5785, N5759, N1850);
not NOT1 (N5786, N5782);
and AND2 (N5787, N5760, N756);
nand NAND3 (N5788, N5780, N2930, N1649);
nand NAND3 (N5789, N5783, N370, N3695);
not NOT1 (N5790, N5789);
xor XOR2 (N5791, N5786, N1037);
nand NAND2 (N5792, N5787, N5198);
buf BUF1 (N5793, N5779);
nand NAND4 (N5794, N5773, N3275, N3709, N1622);
nand NAND4 (N5795, N5784, N5781, N5355, N4724);
and AND2 (N5796, N5790, N2572);
xor XOR2 (N5797, N5796, N5553);
xor XOR2 (N5798, N5797, N2382);
or OR2 (N5799, N5794, N3787);
not NOT1 (N5800, N5788);
xor XOR2 (N5801, N5793, N4636);
buf BUF1 (N5802, N5801);
xor XOR2 (N5803, N5791, N2457);
buf BUF1 (N5804, N5776);
xor XOR2 (N5805, N5795, N3145);
nand NAND2 (N5806, N5763, N1992);
nand NAND3 (N5807, N5799, N2638, N1657);
xor XOR2 (N5808, N5800, N333);
or OR4 (N5809, N5798, N2001, N3631, N3190);
not NOT1 (N5810, N5804);
not NOT1 (N5811, N5785);
not NOT1 (N5812, N5809);
or OR3 (N5813, N5803, N4293, N3013);
buf BUF1 (N5814, N5810);
buf BUF1 (N5815, N5807);
not NOT1 (N5816, N5808);
buf BUF1 (N5817, N5816);
buf BUF1 (N5818, N5811);
not NOT1 (N5819, N5817);
nor NOR2 (N5820, N5814, N36);
xor XOR2 (N5821, N5802, N3908);
buf BUF1 (N5822, N5805);
and AND3 (N5823, N5812, N3462, N126);
nor NOR3 (N5824, N5818, N4079, N5778);
xor XOR2 (N5825, N5820, N5608);
xor XOR2 (N5826, N5806, N1859);
or OR2 (N5827, N5823, N2906);
not NOT1 (N5828, N5819);
nor NOR3 (N5829, N5813, N881, N3654);
or OR3 (N5830, N5828, N2387, N4430);
and AND4 (N5831, N5824, N159, N5725, N1407);
not NOT1 (N5832, N5821);
or OR4 (N5833, N5815, N5450, N3537, N4745);
nand NAND3 (N5834, N5831, N1737, N1064);
and AND3 (N5835, N5832, N327, N1253);
or OR3 (N5836, N5792, N2077, N4053);
and AND2 (N5837, N5825, N4721);
and AND4 (N5838, N5834, N2471, N1999, N4032);
and AND3 (N5839, N5822, N4754, N4974);
buf BUF1 (N5840, N5833);
and AND3 (N5841, N5826, N2846, N168);
or OR2 (N5842, N5841, N5634);
and AND2 (N5843, N5830, N3491);
nor NOR3 (N5844, N5842, N2755, N1217);
xor XOR2 (N5845, N5843, N5659);
buf BUF1 (N5846, N5844);
not NOT1 (N5847, N5839);
or OR4 (N5848, N5827, N1650, N146, N1298);
or OR4 (N5849, N5848, N1960, N4088, N4004);
and AND2 (N5850, N5836, N3291);
xor XOR2 (N5851, N5837, N5825);
nand NAND4 (N5852, N5845, N3494, N2136, N71);
or OR2 (N5853, N5835, N2272);
nor NOR2 (N5854, N5852, N5803);
or OR4 (N5855, N5850, N3666, N1960, N5398);
buf BUF1 (N5856, N5847);
nor NOR4 (N5857, N5856, N4067, N3108, N3674);
buf BUF1 (N5858, N5857);
nand NAND4 (N5859, N5854, N5092, N3788, N5619);
nand NAND4 (N5860, N5858, N4285, N2978, N673);
nor NOR2 (N5861, N5849, N3448);
nand NAND3 (N5862, N5860, N1159, N3509);
buf BUF1 (N5863, N5829);
xor XOR2 (N5864, N5863, N1962);
nor NOR2 (N5865, N5838, N32);
or OR2 (N5866, N5861, N665);
buf BUF1 (N5867, N5853);
and AND2 (N5868, N5851, N5058);
not NOT1 (N5869, N5867);
buf BUF1 (N5870, N5840);
nor NOR4 (N5871, N5866, N809, N148, N2180);
or OR2 (N5872, N5855, N588);
or OR4 (N5873, N5846, N1725, N1420, N4051);
nor NOR4 (N5874, N5859, N1295, N2942, N2489);
nand NAND4 (N5875, N5874, N224, N1377, N65);
xor XOR2 (N5876, N5868, N4946);
nor NOR3 (N5877, N5870, N2774, N2383);
nand NAND3 (N5878, N5869, N2269, N194);
not NOT1 (N5879, N5864);
nor NOR3 (N5880, N5862, N1828, N4393);
nand NAND3 (N5881, N5873, N2725, N5161);
buf BUF1 (N5882, N5879);
not NOT1 (N5883, N5865);
not NOT1 (N5884, N5883);
not NOT1 (N5885, N5871);
not NOT1 (N5886, N5876);
nor NOR4 (N5887, N5875, N62, N3087, N441);
nor NOR3 (N5888, N5884, N1245, N3526);
buf BUF1 (N5889, N5881);
xor XOR2 (N5890, N5889, N1747);
nor NOR4 (N5891, N5878, N3488, N4762, N3236);
nand NAND4 (N5892, N5882, N3960, N3268, N5065);
nand NAND3 (N5893, N5892, N3383, N305);
nand NAND3 (N5894, N5886, N517, N5801);
buf BUF1 (N5895, N5880);
not NOT1 (N5896, N5893);
not NOT1 (N5897, N5872);
not NOT1 (N5898, N5877);
not NOT1 (N5899, N5885);
nand NAND2 (N5900, N5896, N1900);
not NOT1 (N5901, N5900);
nor NOR3 (N5902, N5891, N2317, N5120);
nor NOR2 (N5903, N5897, N4844);
buf BUF1 (N5904, N5894);
xor XOR2 (N5905, N5888, N4909);
and AND4 (N5906, N5904, N2182, N5815, N5050);
nor NOR4 (N5907, N5905, N5556, N2324, N234);
nand NAND3 (N5908, N5898, N2061, N5384);
or OR3 (N5909, N5902, N1752, N5141);
not NOT1 (N5910, N5906);
and AND3 (N5911, N5903, N4739, N4089);
not NOT1 (N5912, N5907);
nor NOR2 (N5913, N5908, N4594);
xor XOR2 (N5914, N5909, N1262);
nor NOR2 (N5915, N5895, N5184);
and AND2 (N5916, N5890, N1339);
nand NAND3 (N5917, N5910, N5438, N209);
buf BUF1 (N5918, N5917);
nor NOR2 (N5919, N5901, N797);
buf BUF1 (N5920, N5887);
xor XOR2 (N5921, N5919, N2877);
not NOT1 (N5922, N5899);
nor NOR3 (N5923, N5912, N3941, N1953);
and AND2 (N5924, N5922, N2695);
nand NAND4 (N5925, N5915, N2955, N3623, N892);
not NOT1 (N5926, N5921);
not NOT1 (N5927, N5923);
nand NAND2 (N5928, N5920, N5780);
not NOT1 (N5929, N5916);
nor NOR4 (N5930, N5913, N148, N2135, N707);
buf BUF1 (N5931, N5928);
xor XOR2 (N5932, N5930, N1503);
nor NOR4 (N5933, N5914, N5762, N304, N1758);
nand NAND3 (N5934, N5933, N783, N3808);
nand NAND2 (N5935, N5934, N4062);
buf BUF1 (N5936, N5931);
nor NOR4 (N5937, N5936, N5486, N5267, N1100);
nand NAND2 (N5938, N5935, N2576);
buf BUF1 (N5939, N5911);
or OR2 (N5940, N5925, N1481);
not NOT1 (N5941, N5918);
nand NAND2 (N5942, N5941, N5244);
nor NOR2 (N5943, N5940, N3377);
or OR2 (N5944, N5939, N3103);
not NOT1 (N5945, N5929);
nand NAND4 (N5946, N5945, N5662, N5419, N5017);
nand NAND2 (N5947, N5937, N2403);
nand NAND2 (N5948, N5946, N5227);
buf BUF1 (N5949, N5938);
or OR3 (N5950, N5947, N2872, N3530);
nand NAND3 (N5951, N5948, N4788, N4945);
xor XOR2 (N5952, N5950, N1118);
and AND3 (N5953, N5926, N3305, N5587);
nand NAND2 (N5954, N5943, N457);
or OR2 (N5955, N5942, N1040);
or OR2 (N5956, N5944, N3045);
and AND2 (N5957, N5932, N518);
and AND3 (N5958, N5951, N1290, N3074);
xor XOR2 (N5959, N5924, N141);
nor NOR2 (N5960, N5949, N668);
or OR2 (N5961, N5957, N3525);
and AND4 (N5962, N5953, N4447, N786, N2947);
xor XOR2 (N5963, N5952, N3033);
and AND2 (N5964, N5961, N2057);
not NOT1 (N5965, N5959);
buf BUF1 (N5966, N5958);
nor NOR3 (N5967, N5966, N4160, N977);
nand NAND2 (N5968, N5954, N4452);
xor XOR2 (N5969, N5965, N5322);
nand NAND2 (N5970, N5964, N2603);
not NOT1 (N5971, N5963);
not NOT1 (N5972, N5970);
and AND4 (N5973, N5972, N2748, N4446, N3694);
not NOT1 (N5974, N5968);
buf BUF1 (N5975, N5962);
buf BUF1 (N5976, N5971);
and AND2 (N5977, N5956, N5974);
nand NAND3 (N5978, N2405, N3779, N5973);
or OR3 (N5979, N3247, N5276, N4623);
nor NOR3 (N5980, N5969, N2722, N4729);
xor XOR2 (N5981, N5979, N5548);
nand NAND2 (N5982, N5975, N3215);
xor XOR2 (N5983, N5978, N1311);
nor NOR3 (N5984, N5960, N3568, N4553);
xor XOR2 (N5985, N5981, N2961);
buf BUF1 (N5986, N5967);
and AND2 (N5987, N5984, N32);
xor XOR2 (N5988, N5927, N5671);
xor XOR2 (N5989, N5980, N222);
nand NAND4 (N5990, N5989, N1267, N3085, N3338);
xor XOR2 (N5991, N5988, N3914);
buf BUF1 (N5992, N5991);
nor NOR2 (N5993, N5992, N569);
nor NOR2 (N5994, N5993, N382);
or OR2 (N5995, N5977, N2611);
and AND3 (N5996, N5986, N619, N5678);
and AND2 (N5997, N5983, N2777);
xor XOR2 (N5998, N5976, N382);
nor NOR4 (N5999, N5990, N840, N3114, N3804);
nor NOR3 (N6000, N5982, N281, N2509);
nor NOR3 (N6001, N6000, N3351, N5548);
nand NAND4 (N6002, N5994, N4721, N1979, N3845);
xor XOR2 (N6003, N5999, N1385);
nand NAND2 (N6004, N5997, N5332);
and AND4 (N6005, N5996, N5720, N2619, N1380);
nor NOR3 (N6006, N5985, N1646, N1639);
buf BUF1 (N6007, N5987);
not NOT1 (N6008, N6001);
or OR4 (N6009, N6008, N233, N3771, N5054);
nor NOR4 (N6010, N6003, N5842, N1086, N3380);
buf BUF1 (N6011, N6002);
xor XOR2 (N6012, N5998, N3689);
not NOT1 (N6013, N6009);
nor NOR2 (N6014, N6007, N4276);
buf BUF1 (N6015, N6004);
not NOT1 (N6016, N6015);
nand NAND2 (N6017, N5955, N5138);
and AND3 (N6018, N6012, N5389, N4346);
or OR4 (N6019, N6016, N681, N4320, N3236);
or OR2 (N6020, N6019, N5573);
nor NOR4 (N6021, N6011, N4609, N401, N1833);
nand NAND4 (N6022, N6020, N2056, N4890, N2460);
xor XOR2 (N6023, N6021, N4543);
and AND3 (N6024, N6022, N4503, N5682);
buf BUF1 (N6025, N6023);
and AND4 (N6026, N6014, N3217, N2563, N5495);
nor NOR4 (N6027, N6024, N5907, N2128, N2243);
nand NAND2 (N6028, N6013, N3507);
and AND4 (N6029, N6025, N639, N4137, N5155);
nand NAND3 (N6030, N6006, N3805, N4022);
xor XOR2 (N6031, N6028, N5107);
nand NAND2 (N6032, N6026, N4671);
not NOT1 (N6033, N6005);
buf BUF1 (N6034, N6010);
and AND3 (N6035, N6034, N12, N5029);
nand NAND2 (N6036, N6031, N650);
and AND2 (N6037, N6027, N1039);
xor XOR2 (N6038, N6018, N6023);
and AND4 (N6039, N6035, N2961, N109, N523);
buf BUF1 (N6040, N6030);
nor NOR3 (N6041, N6032, N2594, N2835);
nand NAND4 (N6042, N6039, N2427, N356, N1859);
buf BUF1 (N6043, N6041);
or OR4 (N6044, N5995, N3719, N5089, N526);
not NOT1 (N6045, N6036);
not NOT1 (N6046, N6029);
nor NOR2 (N6047, N6044, N4068);
nand NAND4 (N6048, N6037, N6008, N2742, N5877);
nand NAND4 (N6049, N6017, N5403, N1602, N5092);
xor XOR2 (N6050, N6043, N149);
not NOT1 (N6051, N6047);
buf BUF1 (N6052, N6046);
or OR4 (N6053, N6038, N447, N2706, N5640);
buf BUF1 (N6054, N6052);
or OR4 (N6055, N6033, N4156, N2930, N1801);
nor NOR2 (N6056, N6050, N1732);
nor NOR3 (N6057, N6048, N320, N5792);
buf BUF1 (N6058, N6049);
not NOT1 (N6059, N6054);
or OR2 (N6060, N6045, N2656);
or OR4 (N6061, N6059, N3688, N1881, N3032);
nand NAND3 (N6062, N6056, N2459, N3816);
nand NAND3 (N6063, N6060, N665, N2271);
not NOT1 (N6064, N6053);
or OR4 (N6065, N6042, N1739, N4889, N5734);
nand NAND3 (N6066, N6061, N3189, N2386);
not NOT1 (N6067, N6055);
buf BUF1 (N6068, N6066);
or OR3 (N6069, N6063, N864, N4790);
xor XOR2 (N6070, N6069, N4489);
xor XOR2 (N6071, N6067, N3675);
not NOT1 (N6072, N6071);
xor XOR2 (N6073, N6051, N2892);
xor XOR2 (N6074, N6058, N894);
nand NAND4 (N6075, N6065, N1994, N1821, N52);
nand NAND2 (N6076, N6068, N3377);
and AND4 (N6077, N6057, N4351, N3767, N2614);
or OR3 (N6078, N6076, N2883, N345);
and AND2 (N6079, N6062, N2994);
not NOT1 (N6080, N6073);
nand NAND4 (N6081, N6075, N2731, N6038, N5311);
buf BUF1 (N6082, N6078);
nand NAND3 (N6083, N6072, N3157, N5303);
and AND4 (N6084, N6074, N6047, N2304, N4276);
xor XOR2 (N6085, N6070, N4951);
buf BUF1 (N6086, N6064);
xor XOR2 (N6087, N6040, N1713);
xor XOR2 (N6088, N6077, N1684);
or OR3 (N6089, N6081, N6072, N3271);
not NOT1 (N6090, N6080);
xor XOR2 (N6091, N6085, N5100);
or OR4 (N6092, N6086, N1116, N6072, N5082);
and AND2 (N6093, N6082, N3997);
xor XOR2 (N6094, N6088, N2003);
nor NOR4 (N6095, N6084, N4173, N4554, N4317);
buf BUF1 (N6096, N6090);
not NOT1 (N6097, N6094);
buf BUF1 (N6098, N6096);
xor XOR2 (N6099, N6083, N2989);
xor XOR2 (N6100, N6087, N2871);
nor NOR3 (N6101, N6097, N1143, N3897);
xor XOR2 (N6102, N6095, N5548);
not NOT1 (N6103, N6102);
nor NOR4 (N6104, N6093, N2164, N5357, N1193);
nor NOR2 (N6105, N6103, N1767);
nand NAND2 (N6106, N6079, N4824);
or OR2 (N6107, N6105, N1835);
nor NOR2 (N6108, N6091, N2853);
not NOT1 (N6109, N6107);
or OR2 (N6110, N6101, N4115);
or OR3 (N6111, N6092, N4166, N2310);
xor XOR2 (N6112, N6110, N2228);
buf BUF1 (N6113, N6089);
nor NOR3 (N6114, N6113, N4027, N2103);
or OR4 (N6115, N6112, N415, N4541, N3321);
not NOT1 (N6116, N6115);
or OR4 (N6117, N6104, N5655, N2850, N633);
not NOT1 (N6118, N6117);
buf BUF1 (N6119, N6116);
buf BUF1 (N6120, N6108);
or OR2 (N6121, N6118, N1125);
not NOT1 (N6122, N6120);
nor NOR4 (N6123, N6119, N2453, N5396, N4995);
nand NAND2 (N6124, N6123, N5158);
nand NAND2 (N6125, N6106, N206);
xor XOR2 (N6126, N6109, N5886);
buf BUF1 (N6127, N6121);
buf BUF1 (N6128, N6126);
not NOT1 (N6129, N6099);
nor NOR4 (N6130, N6098, N948, N4256, N3944);
buf BUF1 (N6131, N6128);
or OR3 (N6132, N6130, N419, N2663);
and AND3 (N6133, N6129, N1906, N3316);
xor XOR2 (N6134, N6132, N3815);
or OR4 (N6135, N6100, N5317, N2595, N5893);
not NOT1 (N6136, N6134);
xor XOR2 (N6137, N6131, N249);
nand NAND3 (N6138, N6114, N3747, N2541);
or OR3 (N6139, N6127, N2160, N77);
not NOT1 (N6140, N6137);
nand NAND4 (N6141, N6122, N2342, N5604, N6076);
or OR3 (N6142, N6111, N5523, N5460);
nor NOR4 (N6143, N6133, N5444, N3232, N5004);
buf BUF1 (N6144, N6140);
and AND3 (N6145, N6141, N4505, N868);
nand NAND2 (N6146, N6125, N1474);
buf BUF1 (N6147, N6124);
not NOT1 (N6148, N6145);
and AND3 (N6149, N6135, N3673, N34);
or OR3 (N6150, N6139, N6023, N3233);
nor NOR4 (N6151, N6136, N4730, N3808, N3564);
nand NAND4 (N6152, N6150, N2763, N3964, N4360);
or OR2 (N6153, N6151, N4795);
xor XOR2 (N6154, N6138, N5761);
xor XOR2 (N6155, N6143, N1197);
not NOT1 (N6156, N6148);
or OR2 (N6157, N6154, N1672);
buf BUF1 (N6158, N6146);
or OR2 (N6159, N6147, N235);
xor XOR2 (N6160, N6153, N5716);
nor NOR4 (N6161, N6159, N5585, N5330, N2476);
buf BUF1 (N6162, N6156);
and AND2 (N6163, N6160, N548);
nor NOR3 (N6164, N6142, N2956, N3679);
nor NOR4 (N6165, N6162, N4308, N3985, N2137);
and AND4 (N6166, N6158, N4723, N1961, N3168);
nand NAND2 (N6167, N6161, N3087);
not NOT1 (N6168, N6164);
not NOT1 (N6169, N6149);
xor XOR2 (N6170, N6169, N335);
or OR2 (N6171, N6163, N3834);
xor XOR2 (N6172, N6171, N6089);
xor XOR2 (N6173, N6152, N37);
nor NOR3 (N6174, N6168, N228, N3300);
buf BUF1 (N6175, N6174);
nor NOR3 (N6176, N6166, N1174, N3413);
or OR2 (N6177, N6176, N2768);
xor XOR2 (N6178, N6144, N4259);
nand NAND4 (N6179, N6173, N5674, N3794, N398);
nor NOR3 (N6180, N6170, N6118, N5762);
and AND4 (N6181, N6155, N3178, N3706, N5943);
or OR2 (N6182, N6181, N4816);
buf BUF1 (N6183, N6178);
buf BUF1 (N6184, N6182);
or OR4 (N6185, N6172, N5793, N3072, N5078);
nand NAND3 (N6186, N6180, N2872, N5527);
not NOT1 (N6187, N6157);
and AND2 (N6188, N6185, N4747);
not NOT1 (N6189, N6184);
xor XOR2 (N6190, N6188, N3595);
nand NAND2 (N6191, N6167, N5265);
nor NOR2 (N6192, N6186, N4718);
nand NAND4 (N6193, N6175, N1146, N4769, N864);
and AND3 (N6194, N6179, N1584, N1839);
not NOT1 (N6195, N6193);
buf BUF1 (N6196, N6194);
xor XOR2 (N6197, N6191, N2690);
and AND3 (N6198, N6165, N2601, N936);
buf BUF1 (N6199, N6192);
nor NOR2 (N6200, N6183, N6056);
or OR4 (N6201, N6198, N5901, N2976, N1512);
nand NAND4 (N6202, N6195, N4054, N4427, N4754);
not NOT1 (N6203, N6189);
nor NOR2 (N6204, N6190, N3056);
nand NAND2 (N6205, N6203, N1405);
nand NAND4 (N6206, N6200, N509, N950, N507);
or OR4 (N6207, N6197, N2227, N676, N3180);
or OR4 (N6208, N6199, N3773, N770, N1650);
buf BUF1 (N6209, N6206);
buf BUF1 (N6210, N6201);
or OR2 (N6211, N6205, N4191);
buf BUF1 (N6212, N6208);
nand NAND2 (N6213, N6202, N3947);
not NOT1 (N6214, N6177);
and AND2 (N6215, N6187, N4638);
buf BUF1 (N6216, N6215);
or OR4 (N6217, N6204, N5151, N5686, N2527);
xor XOR2 (N6218, N6211, N4591);
nand NAND2 (N6219, N6210, N5748);
xor XOR2 (N6220, N6219, N5306);
and AND3 (N6221, N6220, N6069, N1623);
and AND4 (N6222, N6207, N3589, N3625, N3534);
nand NAND2 (N6223, N6218, N4199);
xor XOR2 (N6224, N6213, N2180);
not NOT1 (N6225, N6222);
buf BUF1 (N6226, N6221);
nand NAND4 (N6227, N6212, N1306, N5483, N3277);
nor NOR3 (N6228, N6216, N4927, N486);
nand NAND3 (N6229, N6224, N2661, N4627);
and AND3 (N6230, N6217, N2165, N3824);
not NOT1 (N6231, N6209);
and AND2 (N6232, N6228, N5662);
xor XOR2 (N6233, N6230, N5862);
nor NOR3 (N6234, N6227, N4509, N1278);
nand NAND4 (N6235, N6214, N998, N5526, N4739);
and AND3 (N6236, N6234, N1131, N5171);
buf BUF1 (N6237, N6229);
or OR2 (N6238, N6232, N3167);
not NOT1 (N6239, N6226);
xor XOR2 (N6240, N6235, N1478);
not NOT1 (N6241, N6240);
nor NOR4 (N6242, N6237, N325, N2804, N4780);
or OR4 (N6243, N6241, N3539, N86, N1856);
nand NAND3 (N6244, N6223, N1179, N5854);
nor NOR2 (N6245, N6238, N648);
nand NAND2 (N6246, N6243, N840);
or OR3 (N6247, N6244, N4916, N3823);
buf BUF1 (N6248, N6196);
nand NAND3 (N6249, N6246, N2312, N3397);
and AND2 (N6250, N6225, N6025);
nand NAND2 (N6251, N6239, N4329);
buf BUF1 (N6252, N6242);
xor XOR2 (N6253, N6245, N1228);
nand NAND3 (N6254, N6252, N1620, N3707);
xor XOR2 (N6255, N6247, N5140);
or OR4 (N6256, N6233, N5021, N1413, N4429);
nand NAND3 (N6257, N6254, N2733, N1929);
nor NOR2 (N6258, N6253, N6121);
nor NOR3 (N6259, N6255, N4589, N323);
nand NAND4 (N6260, N6257, N4792, N2327, N1498);
nand NAND3 (N6261, N6248, N798, N5463);
xor XOR2 (N6262, N6261, N5893);
nand NAND2 (N6263, N6262, N3022);
nand NAND3 (N6264, N6236, N1917, N802);
buf BUF1 (N6265, N6259);
and AND4 (N6266, N6263, N4028, N1007, N5163);
or OR2 (N6267, N6260, N3506);
xor XOR2 (N6268, N6231, N2510);
buf BUF1 (N6269, N6266);
nand NAND3 (N6270, N6251, N2701, N4351);
nand NAND3 (N6271, N6270, N4881, N5851);
nand NAND2 (N6272, N6256, N3924);
xor XOR2 (N6273, N6264, N1828);
buf BUF1 (N6274, N6272);
and AND3 (N6275, N6268, N3639, N964);
nor NOR2 (N6276, N6250, N2620);
nand NAND4 (N6277, N6269, N3870, N1349, N4078);
not NOT1 (N6278, N6267);
not NOT1 (N6279, N6276);
nand NAND3 (N6280, N6271, N5688, N1994);
not NOT1 (N6281, N6249);
and AND2 (N6282, N6273, N5722);
not NOT1 (N6283, N6274);
or OR3 (N6284, N6277, N402, N3568);
xor XOR2 (N6285, N6284, N2358);
xor XOR2 (N6286, N6279, N3856);
and AND3 (N6287, N6275, N3100, N3556);
or OR4 (N6288, N6285, N4742, N5907, N5360);
nand NAND4 (N6289, N6286, N2773, N4200, N2449);
nor NOR3 (N6290, N6280, N4721, N2985);
not NOT1 (N6291, N6287);
nor NOR4 (N6292, N6289, N2576, N5654, N278);
not NOT1 (N6293, N6265);
nand NAND4 (N6294, N6291, N1427, N6281, N5960);
and AND4 (N6295, N4537, N2968, N1981, N5039);
not NOT1 (N6296, N6282);
xor XOR2 (N6297, N6292, N3945);
and AND2 (N6298, N6295, N611);
not NOT1 (N6299, N6296);
not NOT1 (N6300, N6278);
nor NOR4 (N6301, N6288, N5992, N3653, N2011);
and AND4 (N6302, N6301, N5121, N178, N642);
nand NAND4 (N6303, N6258, N4306, N5250, N3240);
nor NOR3 (N6304, N6294, N3699, N331);
nor NOR3 (N6305, N6293, N4263, N6177);
or OR2 (N6306, N6302, N2111);
xor XOR2 (N6307, N6299, N150);
not NOT1 (N6308, N6306);
nand NAND3 (N6309, N6290, N2483, N3040);
buf BUF1 (N6310, N6308);
xor XOR2 (N6311, N6304, N1398);
not NOT1 (N6312, N6297);
nand NAND2 (N6313, N6303, N5419);
not NOT1 (N6314, N6311);
xor XOR2 (N6315, N6313, N5902);
not NOT1 (N6316, N6315);
nor NOR2 (N6317, N6309, N1911);
buf BUF1 (N6318, N6300);
nor NOR3 (N6319, N6298, N2685, N4825);
nor NOR4 (N6320, N6314, N2643, N3062, N2632);
nand NAND3 (N6321, N6318, N3957, N3689);
nand NAND2 (N6322, N6321, N336);
nand NAND3 (N6323, N6322, N6012, N1647);
nand NAND2 (N6324, N6310, N5234);
xor XOR2 (N6325, N6323, N3172);
nor NOR3 (N6326, N6283, N1572, N1730);
xor XOR2 (N6327, N6312, N5164);
nand NAND3 (N6328, N6316, N4437, N5845);
nand NAND2 (N6329, N6307, N1478);
not NOT1 (N6330, N6327);
or OR3 (N6331, N6319, N5434, N5571);
nand NAND3 (N6332, N6328, N866, N2661);
xor XOR2 (N6333, N6329, N221);
buf BUF1 (N6334, N6324);
not NOT1 (N6335, N6330);
nand NAND2 (N6336, N6325, N4417);
xor XOR2 (N6337, N6305, N5402);
buf BUF1 (N6338, N6334);
nor NOR4 (N6339, N6317, N3337, N1741, N3331);
and AND2 (N6340, N6338, N1696);
xor XOR2 (N6341, N6336, N3364);
nor NOR4 (N6342, N6341, N5134, N1742, N5196);
or OR2 (N6343, N6332, N2191);
xor XOR2 (N6344, N6335, N3428);
nand NAND4 (N6345, N6326, N2456, N1198, N3020);
nor NOR4 (N6346, N6337, N5259, N5752, N2105);
xor XOR2 (N6347, N6346, N2315);
or OR3 (N6348, N6333, N4296, N5896);
and AND3 (N6349, N6343, N2856, N2150);
buf BUF1 (N6350, N6340);
or OR2 (N6351, N6349, N1703);
buf BUF1 (N6352, N6320);
and AND2 (N6353, N6345, N5809);
buf BUF1 (N6354, N6353);
buf BUF1 (N6355, N6331);
and AND4 (N6356, N6342, N1538, N6339, N4556);
buf BUF1 (N6357, N6061);
nor NOR2 (N6358, N6354, N5272);
xor XOR2 (N6359, N6352, N1359);
and AND2 (N6360, N6344, N5191);
and AND4 (N6361, N6348, N5106, N5384, N3515);
or OR3 (N6362, N6360, N1520, N4869);
xor XOR2 (N6363, N6355, N515);
nand NAND4 (N6364, N6351, N4233, N1310, N2229);
nor NOR3 (N6365, N6362, N6203, N4817);
not NOT1 (N6366, N6347);
nor NOR4 (N6367, N6357, N5804, N700, N5495);
xor XOR2 (N6368, N6366, N4981);
or OR4 (N6369, N6359, N4843, N4957, N2316);
not NOT1 (N6370, N6367);
or OR3 (N6371, N6368, N4159, N711);
nand NAND2 (N6372, N6370, N1516);
nand NAND2 (N6373, N6356, N4157);
nor NOR2 (N6374, N6373, N2065);
nor NOR3 (N6375, N6358, N3647, N5883);
not NOT1 (N6376, N6375);
or OR3 (N6377, N6365, N3397, N158);
xor XOR2 (N6378, N6363, N1050);
nand NAND2 (N6379, N6374, N706);
and AND2 (N6380, N6379, N6307);
xor XOR2 (N6381, N6378, N368);
and AND2 (N6382, N6380, N2976);
or OR4 (N6383, N6369, N5065, N949, N4534);
xor XOR2 (N6384, N6376, N5163);
not NOT1 (N6385, N6371);
buf BUF1 (N6386, N6382);
not NOT1 (N6387, N6372);
nand NAND2 (N6388, N6384, N1086);
buf BUF1 (N6389, N6381);
and AND4 (N6390, N6361, N2234, N2912, N1919);
or OR4 (N6391, N6377, N3329, N3028, N6211);
nand NAND4 (N6392, N6389, N4062, N2864, N6268);
not NOT1 (N6393, N6391);
nand NAND4 (N6394, N6393, N5487, N314, N2808);
buf BUF1 (N6395, N6386);
and AND2 (N6396, N6394, N445);
xor XOR2 (N6397, N6364, N2191);
buf BUF1 (N6398, N6350);
buf BUF1 (N6399, N6395);
nand NAND2 (N6400, N6385, N2834);
or OR3 (N6401, N6396, N4763, N1245);
buf BUF1 (N6402, N6400);
xor XOR2 (N6403, N6398, N6264);
nor NOR4 (N6404, N6388, N4334, N5524, N698);
nand NAND2 (N6405, N6402, N6045);
or OR4 (N6406, N6390, N1952, N3984, N4363);
buf BUF1 (N6407, N6383);
buf BUF1 (N6408, N6387);
xor XOR2 (N6409, N6401, N5802);
and AND4 (N6410, N6392, N254, N4539, N1115);
nor NOR3 (N6411, N6408, N4622, N4718);
and AND2 (N6412, N6403, N575);
and AND2 (N6413, N6404, N1366);
nor NOR2 (N6414, N6399, N4390);
or OR4 (N6415, N6410, N1248, N5883, N6314);
nor NOR3 (N6416, N6409, N35, N6323);
xor XOR2 (N6417, N6415, N6333);
nor NOR2 (N6418, N6411, N5176);
xor XOR2 (N6419, N6407, N874);
buf BUF1 (N6420, N6406);
not NOT1 (N6421, N6416);
nor NOR4 (N6422, N6413, N5042, N4570, N4182);
xor XOR2 (N6423, N6419, N5423);
endmodule