// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N3515,N3517,N3510,N3489,N3514,N3513,N3503,N3494,N3516,N3518;

buf BUF1 (N19, N12);
nand NAND4 (N20, N18, N14, N13, N4);
nor NOR4 (N21, N14, N6, N18, N15);
nor NOR4 (N22, N15, N3, N1, N4);
nand NAND3 (N23, N15, N8, N16);
and AND2 (N24, N6, N16);
not NOT1 (N25, N1);
and AND4 (N26, N1, N5, N6, N24);
and AND4 (N27, N14, N16, N14, N7);
xor XOR2 (N28, N17, N12);
and AND2 (N29, N10, N9);
not NOT1 (N30, N21);
not NOT1 (N31, N20);
not NOT1 (N32, N29);
buf BUF1 (N33, N31);
buf BUF1 (N34, N33);
nor NOR3 (N35, N26, N15, N32);
buf BUF1 (N36, N16);
nor NOR3 (N37, N30, N34, N14);
not NOT1 (N38, N15);
buf BUF1 (N39, N25);
nand NAND3 (N40, N23, N32, N30);
or OR2 (N41, N35, N9);
buf BUF1 (N42, N28);
not NOT1 (N43, N36);
or OR2 (N44, N22, N30);
nand NAND4 (N45, N44, N44, N16, N18);
and AND4 (N46, N43, N29, N29, N7);
and AND3 (N47, N39, N15, N44);
nor NOR2 (N48, N19, N35);
and AND4 (N49, N42, N39, N38, N27);
buf BUF1 (N50, N22);
xor XOR2 (N51, N15, N29);
not NOT1 (N52, N46);
or OR2 (N53, N51, N9);
xor XOR2 (N54, N52, N11);
or OR2 (N55, N48, N13);
buf BUF1 (N56, N49);
nand NAND3 (N57, N55, N1, N24);
nor NOR4 (N58, N53, N16, N55, N47);
or OR3 (N59, N37, N40, N20);
and AND3 (N60, N48, N2, N22);
nor NOR4 (N61, N52, N59, N10, N5);
or OR3 (N62, N26, N55, N33);
not NOT1 (N63, N58);
buf BUF1 (N64, N54);
buf BUF1 (N65, N45);
nor NOR3 (N66, N65, N3, N48);
or OR2 (N67, N66, N48);
and AND2 (N68, N67, N16);
and AND3 (N69, N62, N32, N68);
xor XOR2 (N70, N54, N13);
xor XOR2 (N71, N41, N53);
buf BUF1 (N72, N56);
and AND2 (N73, N64, N9);
buf BUF1 (N74, N63);
nand NAND2 (N75, N70, N35);
xor XOR2 (N76, N72, N2);
nand NAND4 (N77, N50, N28, N34, N59);
not NOT1 (N78, N60);
nor NOR4 (N79, N75, N49, N46, N19);
or OR3 (N80, N73, N19, N31);
and AND3 (N81, N61, N53, N60);
nand NAND4 (N82, N71, N46, N34, N57);
nor NOR2 (N83, N74, N33);
buf BUF1 (N84, N15);
and AND2 (N85, N79, N71);
not NOT1 (N86, N84);
nor NOR2 (N87, N76, N85);
nor NOR4 (N88, N6, N48, N13, N18);
buf BUF1 (N89, N78);
nand NAND2 (N90, N88, N17);
nand NAND3 (N91, N90, N2, N8);
or OR2 (N92, N91, N69);
and AND4 (N93, N48, N46, N68, N52);
not NOT1 (N94, N77);
not NOT1 (N95, N92);
xor XOR2 (N96, N81, N95);
xor XOR2 (N97, N70, N76);
not NOT1 (N98, N83);
not NOT1 (N99, N80);
or OR2 (N100, N96, N5);
or OR4 (N101, N86, N42, N30, N91);
nand NAND3 (N102, N87, N28, N42);
or OR3 (N103, N98, N51, N61);
nor NOR4 (N104, N99, N100, N37, N21);
xor XOR2 (N105, N102, N82);
nand NAND3 (N106, N64, N20, N26);
nor NOR4 (N107, N79, N15, N27, N56);
xor XOR2 (N108, N103, N71);
nor NOR3 (N109, N104, N43, N88);
nor NOR3 (N110, N106, N79, N95);
not NOT1 (N111, N105);
nand NAND3 (N112, N101, N49, N56);
nand NAND4 (N113, N107, N57, N93, N85);
or OR3 (N114, N74, N113, N27);
nand NAND3 (N115, N103, N82, N81);
and AND4 (N116, N114, N33, N15, N18);
nand NAND2 (N117, N115, N41);
buf BUF1 (N118, N97);
nand NAND3 (N119, N108, N42, N58);
and AND3 (N120, N110, N65, N67);
nor NOR2 (N121, N118, N97);
buf BUF1 (N122, N120);
or OR2 (N123, N122, N10);
xor XOR2 (N124, N112, N37);
nor NOR3 (N125, N117, N35, N19);
not NOT1 (N126, N94);
nor NOR2 (N127, N125, N11);
and AND2 (N128, N116, N10);
nor NOR2 (N129, N127, N8);
nor NOR2 (N130, N109, N27);
buf BUF1 (N131, N130);
not NOT1 (N132, N89);
not NOT1 (N133, N132);
and AND4 (N134, N131, N85, N34, N33);
nor NOR4 (N135, N133, N6, N131, N32);
and AND4 (N136, N111, N14, N66, N24);
nor NOR2 (N137, N134, N25);
or OR4 (N138, N121, N129, N110, N24);
xor XOR2 (N139, N102, N23);
nand NAND4 (N140, N137, N40, N56, N78);
nand NAND2 (N141, N138, N11);
and AND3 (N142, N136, N27, N133);
xor XOR2 (N143, N139, N131);
nand NAND3 (N144, N126, N84, N63);
or OR2 (N145, N128, N3);
nand NAND3 (N146, N135, N74, N101);
and AND4 (N147, N145, N24, N85, N127);
or OR2 (N148, N143, N133);
not NOT1 (N149, N148);
nor NOR3 (N150, N140, N112, N58);
or OR4 (N151, N123, N50, N132, N108);
nand NAND2 (N152, N141, N69);
not NOT1 (N153, N152);
not NOT1 (N154, N144);
buf BUF1 (N155, N150);
and AND4 (N156, N155, N119, N55, N108);
nand NAND3 (N157, N36, N80, N54);
not NOT1 (N158, N156);
nor NOR4 (N159, N147, N69, N60, N84);
and AND2 (N160, N151, N113);
buf BUF1 (N161, N146);
or OR3 (N162, N149, N113, N95);
or OR4 (N163, N154, N135, N76, N151);
not NOT1 (N164, N124);
nand NAND4 (N165, N142, N14, N74, N9);
xor XOR2 (N166, N165, N18);
xor XOR2 (N167, N159, N147);
not NOT1 (N168, N163);
buf BUF1 (N169, N166);
or OR4 (N170, N160, N91, N81, N9);
nor NOR2 (N171, N158, N83);
or OR2 (N172, N164, N99);
buf BUF1 (N173, N157);
not NOT1 (N174, N162);
buf BUF1 (N175, N168);
not NOT1 (N176, N167);
xor XOR2 (N177, N171, N41);
nand NAND3 (N178, N175, N25, N109);
xor XOR2 (N179, N153, N144);
not NOT1 (N180, N179);
xor XOR2 (N181, N178, N106);
nand NAND2 (N182, N177, N167);
not NOT1 (N183, N174);
and AND2 (N184, N176, N66);
nand NAND2 (N185, N182, N76);
not NOT1 (N186, N183);
and AND4 (N187, N184, N176, N72, N28);
buf BUF1 (N188, N169);
or OR2 (N189, N173, N181);
nor NOR3 (N190, N72, N113, N94);
or OR4 (N191, N188, N182, N112, N67);
nor NOR4 (N192, N190, N191, N70, N5);
and AND3 (N193, N183, N137, N47);
nor NOR2 (N194, N192, N165);
nor NOR4 (N195, N185, N123, N170, N11);
buf BUF1 (N196, N135);
nor NOR2 (N197, N189, N184);
buf BUF1 (N198, N180);
or OR3 (N199, N195, N78, N170);
and AND4 (N200, N194, N2, N140, N99);
or OR3 (N201, N186, N109, N87);
or OR2 (N202, N193, N54);
or OR3 (N203, N198, N93, N135);
not NOT1 (N204, N196);
xor XOR2 (N205, N200, N156);
nor NOR4 (N206, N201, N94, N165, N74);
and AND4 (N207, N187, N154, N64, N59);
and AND2 (N208, N204, N167);
or OR4 (N209, N207, N195, N127, N9);
buf BUF1 (N210, N172);
buf BUF1 (N211, N210);
and AND3 (N212, N199, N133, N27);
nor NOR4 (N213, N205, N88, N151, N188);
nor NOR3 (N214, N197, N37, N4);
nor NOR4 (N215, N203, N161, N38, N25);
not NOT1 (N216, N163);
xor XOR2 (N217, N208, N171);
nor NOR3 (N218, N215, N128, N74);
nor NOR3 (N219, N213, N52, N31);
and AND3 (N220, N209, N140, N195);
not NOT1 (N221, N202);
not NOT1 (N222, N218);
or OR2 (N223, N211, N147);
and AND2 (N224, N206, N123);
xor XOR2 (N225, N223, N44);
and AND3 (N226, N219, N191, N186);
nor NOR2 (N227, N214, N84);
xor XOR2 (N228, N224, N112);
nor NOR4 (N229, N225, N151, N199, N73);
nor NOR2 (N230, N229, N218);
xor XOR2 (N231, N227, N72);
and AND2 (N232, N216, N49);
nand NAND3 (N233, N221, N181, N37);
not NOT1 (N234, N230);
buf BUF1 (N235, N217);
buf BUF1 (N236, N212);
and AND4 (N237, N234, N218, N10, N15);
and AND3 (N238, N226, N171, N170);
and AND4 (N239, N238, N17, N82, N201);
nor NOR4 (N240, N232, N96, N92, N82);
xor XOR2 (N241, N235, N177);
buf BUF1 (N242, N233);
nor NOR2 (N243, N222, N221);
or OR4 (N244, N242, N190, N6, N188);
and AND2 (N245, N241, N112);
and AND3 (N246, N220, N33, N131);
nor NOR2 (N247, N243, N222);
nand NAND2 (N248, N239, N27);
and AND2 (N249, N246, N108);
buf BUF1 (N250, N248);
or OR3 (N251, N245, N187, N120);
and AND2 (N252, N250, N212);
nand NAND3 (N253, N244, N70, N97);
not NOT1 (N254, N247);
not NOT1 (N255, N253);
or OR3 (N256, N252, N57, N253);
nor NOR4 (N257, N249, N57, N190, N24);
not NOT1 (N258, N231);
and AND2 (N259, N257, N66);
buf BUF1 (N260, N237);
nand NAND4 (N261, N251, N77, N102, N249);
and AND3 (N262, N261, N62, N251);
nor NOR3 (N263, N260, N164, N218);
or OR3 (N264, N240, N187, N41);
and AND2 (N265, N254, N213);
buf BUF1 (N266, N256);
and AND2 (N267, N228, N241);
nand NAND3 (N268, N265, N85, N67);
not NOT1 (N269, N236);
xor XOR2 (N270, N263, N268);
xor XOR2 (N271, N188, N68);
and AND4 (N272, N266, N207, N249, N189);
not NOT1 (N273, N267);
and AND2 (N274, N271, N83);
nand NAND3 (N275, N255, N166, N23);
nor NOR3 (N276, N275, N194, N76);
nand NAND2 (N277, N270, N94);
buf BUF1 (N278, N262);
and AND2 (N279, N258, N91);
and AND4 (N280, N279, N91, N31, N141);
nand NAND4 (N281, N259, N181, N194, N232);
and AND2 (N282, N277, N157);
buf BUF1 (N283, N282);
xor XOR2 (N284, N264, N226);
buf BUF1 (N285, N280);
or OR4 (N286, N274, N25, N109, N33);
buf BUF1 (N287, N281);
or OR4 (N288, N283, N48, N2, N151);
nand NAND4 (N289, N286, N129, N55, N66);
or OR3 (N290, N272, N24, N4);
xor XOR2 (N291, N273, N124);
and AND3 (N292, N269, N23, N266);
or OR3 (N293, N289, N263, N154);
and AND4 (N294, N284, N242, N143, N185);
nor NOR3 (N295, N278, N12, N230);
and AND3 (N296, N290, N102, N269);
and AND3 (N297, N296, N103, N146);
nor NOR3 (N298, N287, N13, N252);
buf BUF1 (N299, N276);
xor XOR2 (N300, N285, N95);
buf BUF1 (N301, N300);
nor NOR4 (N302, N288, N59, N136, N120);
or OR2 (N303, N301, N38);
buf BUF1 (N304, N293);
or OR4 (N305, N304, N294, N234, N298);
not NOT1 (N306, N138);
nand NAND4 (N307, N141, N292, N255, N206);
not NOT1 (N308, N228);
buf BUF1 (N309, N297);
or OR3 (N310, N309, N97, N101);
nand NAND4 (N311, N305, N294, N121, N80);
not NOT1 (N312, N308);
xor XOR2 (N313, N311, N247);
buf BUF1 (N314, N299);
xor XOR2 (N315, N313, N292);
xor XOR2 (N316, N303, N255);
or OR2 (N317, N307, N313);
nand NAND3 (N318, N306, N204, N241);
not NOT1 (N319, N291);
buf BUF1 (N320, N295);
nand NAND4 (N321, N315, N89, N274, N195);
nand NAND2 (N322, N310, N258);
nand NAND3 (N323, N316, N136, N186);
and AND4 (N324, N317, N263, N165, N8);
xor XOR2 (N325, N324, N29);
buf BUF1 (N326, N318);
and AND4 (N327, N319, N205, N269, N214);
nor NOR2 (N328, N320, N29);
not NOT1 (N329, N312);
buf BUF1 (N330, N323);
xor XOR2 (N331, N322, N317);
xor XOR2 (N332, N330, N214);
nor NOR4 (N333, N326, N55, N55, N54);
nor NOR4 (N334, N328, N25, N91, N234);
nor NOR2 (N335, N334, N30);
nor NOR2 (N336, N314, N271);
and AND3 (N337, N329, N268, N195);
nor NOR2 (N338, N332, N302);
not NOT1 (N339, N108);
or OR2 (N340, N339, N150);
not NOT1 (N341, N331);
buf BUF1 (N342, N327);
xor XOR2 (N343, N340, N340);
or OR2 (N344, N342, N329);
xor XOR2 (N345, N343, N62);
nor NOR4 (N346, N337, N92, N100, N280);
not NOT1 (N347, N341);
or OR3 (N348, N325, N241, N5);
and AND2 (N349, N348, N294);
nand NAND2 (N350, N346, N157);
nor NOR3 (N351, N336, N128, N223);
or OR2 (N352, N350, N165);
xor XOR2 (N353, N344, N87);
nand NAND3 (N354, N335, N106, N151);
or OR2 (N355, N349, N77);
nor NOR4 (N356, N333, N276, N74, N8);
not NOT1 (N357, N353);
nand NAND2 (N358, N357, N34);
and AND4 (N359, N355, N19, N201, N139);
and AND3 (N360, N354, N245, N267);
xor XOR2 (N361, N345, N102);
or OR4 (N362, N356, N29, N121, N83);
nor NOR2 (N363, N352, N260);
nor NOR2 (N364, N360, N20);
buf BUF1 (N365, N321);
buf BUF1 (N366, N365);
not NOT1 (N367, N366);
and AND2 (N368, N361, N342);
and AND3 (N369, N358, N203, N56);
and AND2 (N370, N362, N74);
or OR4 (N371, N364, N13, N118, N80);
nand NAND4 (N372, N370, N365, N135, N305);
xor XOR2 (N373, N347, N372);
not NOT1 (N374, N63);
xor XOR2 (N375, N367, N284);
nand NAND4 (N376, N369, N254, N354, N71);
nand NAND3 (N377, N368, N22, N295);
not NOT1 (N378, N338);
or OR3 (N379, N374, N217, N112);
xor XOR2 (N380, N377, N50);
or OR3 (N381, N379, N158, N285);
not NOT1 (N382, N380);
buf BUF1 (N383, N373);
not NOT1 (N384, N363);
nor NOR2 (N385, N359, N210);
nand NAND2 (N386, N381, N206);
or OR4 (N387, N351, N229, N60, N3);
xor XOR2 (N388, N375, N268);
buf BUF1 (N389, N385);
or OR2 (N390, N387, N111);
nand NAND4 (N391, N376, N350, N3, N229);
not NOT1 (N392, N382);
or OR4 (N393, N383, N201, N363, N206);
xor XOR2 (N394, N384, N111);
xor XOR2 (N395, N393, N312);
and AND4 (N396, N386, N196, N165, N105);
and AND4 (N397, N378, N22, N264, N226);
nor NOR4 (N398, N390, N194, N251, N309);
nor NOR4 (N399, N397, N101, N70, N62);
and AND3 (N400, N388, N277, N192);
nand NAND3 (N401, N371, N173, N34);
buf BUF1 (N402, N392);
nor NOR2 (N403, N394, N261);
not NOT1 (N404, N402);
buf BUF1 (N405, N389);
and AND3 (N406, N395, N159, N224);
nand NAND3 (N407, N404, N321, N174);
or OR2 (N408, N400, N170);
xor XOR2 (N409, N407, N315);
nor NOR2 (N410, N409, N307);
not NOT1 (N411, N399);
nand NAND2 (N412, N391, N220);
xor XOR2 (N413, N411, N342);
and AND4 (N414, N410, N362, N48, N3);
xor XOR2 (N415, N398, N88);
and AND3 (N416, N414, N385, N305);
not NOT1 (N417, N406);
nor NOR2 (N418, N412, N5);
nand NAND4 (N419, N418, N265, N260, N226);
not NOT1 (N420, N417);
nor NOR2 (N421, N420, N411);
or OR3 (N422, N415, N276, N415);
nor NOR2 (N423, N416, N358);
not NOT1 (N424, N421);
or OR4 (N425, N405, N246, N134, N350);
xor XOR2 (N426, N422, N125);
nor NOR2 (N427, N413, N287);
xor XOR2 (N428, N425, N211);
not NOT1 (N429, N428);
nor NOR4 (N430, N426, N159, N212, N360);
and AND3 (N431, N401, N383, N371);
or OR4 (N432, N419, N325, N101, N28);
nor NOR2 (N433, N427, N299);
xor XOR2 (N434, N423, N172);
or OR2 (N435, N430, N351);
not NOT1 (N436, N403);
buf BUF1 (N437, N396);
xor XOR2 (N438, N434, N211);
xor XOR2 (N439, N429, N251);
xor XOR2 (N440, N438, N99);
xor XOR2 (N441, N433, N124);
nor NOR4 (N442, N435, N409, N158, N284);
or OR4 (N443, N432, N214, N164, N375);
and AND2 (N444, N436, N401);
nand NAND2 (N445, N443, N159);
xor XOR2 (N446, N439, N55);
nand NAND2 (N447, N440, N63);
not NOT1 (N448, N446);
or OR3 (N449, N445, N114, N444);
and AND3 (N450, N169, N13, N25);
xor XOR2 (N451, N442, N44);
not NOT1 (N452, N408);
xor XOR2 (N453, N431, N382);
xor XOR2 (N454, N453, N41);
not NOT1 (N455, N451);
and AND2 (N456, N448, N378);
not NOT1 (N457, N437);
not NOT1 (N458, N450);
nor NOR3 (N459, N458, N59, N98);
buf BUF1 (N460, N441);
nor NOR2 (N461, N456, N22);
and AND3 (N462, N455, N427, N196);
nor NOR2 (N463, N462, N379);
and AND3 (N464, N457, N210, N119);
nor NOR4 (N465, N464, N253, N257, N305);
xor XOR2 (N466, N459, N148);
buf BUF1 (N467, N424);
not NOT1 (N468, N460);
xor XOR2 (N469, N449, N283);
buf BUF1 (N470, N465);
xor XOR2 (N471, N469, N392);
nand NAND3 (N472, N447, N219, N351);
nand NAND2 (N473, N467, N230);
or OR4 (N474, N468, N186, N239, N367);
and AND3 (N475, N463, N248, N83);
xor XOR2 (N476, N472, N213);
xor XOR2 (N477, N474, N69);
buf BUF1 (N478, N470);
not NOT1 (N479, N478);
not NOT1 (N480, N476);
nand NAND2 (N481, N461, N374);
and AND2 (N482, N452, N122);
buf BUF1 (N483, N475);
xor XOR2 (N484, N483, N30);
or OR3 (N485, N481, N77, N219);
buf BUF1 (N486, N454);
xor XOR2 (N487, N479, N457);
and AND2 (N488, N471, N160);
nand NAND2 (N489, N485, N397);
or OR4 (N490, N480, N165, N123, N290);
or OR2 (N491, N490, N476);
nor NOR4 (N492, N484, N191, N108, N314);
or OR2 (N493, N477, N35);
nor NOR3 (N494, N492, N413, N25);
not NOT1 (N495, N488);
or OR2 (N496, N466, N234);
nand NAND4 (N497, N473, N73, N197, N193);
buf BUF1 (N498, N487);
or OR2 (N499, N496, N287);
nor NOR2 (N500, N499, N82);
nand NAND4 (N501, N482, N56, N121, N411);
or OR2 (N502, N495, N54);
not NOT1 (N503, N493);
and AND4 (N504, N503, N155, N218, N421);
buf BUF1 (N505, N486);
not NOT1 (N506, N489);
or OR4 (N507, N498, N278, N128, N238);
buf BUF1 (N508, N500);
or OR2 (N509, N501, N268);
nand NAND3 (N510, N494, N428, N103);
or OR4 (N511, N497, N57, N242, N31);
or OR3 (N512, N510, N204, N271);
and AND2 (N513, N506, N369);
xor XOR2 (N514, N512, N195);
and AND3 (N515, N509, N135, N136);
or OR2 (N516, N491, N73);
nand NAND4 (N517, N514, N473, N424, N93);
and AND3 (N518, N505, N365, N129);
xor XOR2 (N519, N507, N468);
nand NAND3 (N520, N516, N505, N420);
xor XOR2 (N521, N518, N32);
xor XOR2 (N522, N511, N48);
not NOT1 (N523, N522);
and AND4 (N524, N523, N381, N276, N148);
and AND4 (N525, N521, N387, N510, N412);
nand NAND4 (N526, N508, N293, N17, N127);
nor NOR2 (N527, N519, N259);
nor NOR2 (N528, N513, N67);
nor NOR2 (N529, N504, N14);
xor XOR2 (N530, N502, N94);
nand NAND3 (N531, N528, N513, N185);
nand NAND2 (N532, N526, N316);
nand NAND3 (N533, N527, N488, N274);
or OR3 (N534, N530, N330, N419);
nor NOR2 (N535, N531, N4);
nand NAND4 (N536, N525, N381, N450, N146);
xor XOR2 (N537, N524, N271);
not NOT1 (N538, N515);
or OR2 (N539, N535, N264);
not NOT1 (N540, N536);
not NOT1 (N541, N534);
xor XOR2 (N542, N541, N120);
and AND4 (N543, N517, N426, N97, N97);
nand NAND3 (N544, N539, N408, N270);
buf BUF1 (N545, N520);
and AND2 (N546, N538, N339);
nand NAND2 (N547, N544, N422);
nor NOR4 (N548, N546, N252, N401, N62);
not NOT1 (N549, N543);
nand NAND3 (N550, N549, N36, N92);
or OR3 (N551, N545, N315, N533);
nor NOR3 (N552, N428, N301, N160);
and AND2 (N553, N552, N233);
and AND2 (N554, N532, N524);
buf BUF1 (N555, N551);
buf BUF1 (N556, N550);
xor XOR2 (N557, N537, N235);
xor XOR2 (N558, N555, N158);
xor XOR2 (N559, N557, N84);
xor XOR2 (N560, N548, N218);
or OR4 (N561, N553, N107, N489, N136);
xor XOR2 (N562, N547, N450);
and AND4 (N563, N559, N155, N426, N251);
not NOT1 (N564, N562);
and AND4 (N565, N542, N22, N474, N187);
not NOT1 (N566, N556);
xor XOR2 (N567, N563, N397);
not NOT1 (N568, N540);
xor XOR2 (N569, N566, N560);
buf BUF1 (N570, N189);
or OR4 (N571, N569, N39, N488, N475);
nor NOR3 (N572, N564, N100, N24);
buf BUF1 (N573, N554);
buf BUF1 (N574, N573);
nor NOR4 (N575, N558, N146, N428, N238);
nand NAND4 (N576, N529, N352, N557, N463);
nor NOR4 (N577, N572, N336, N292, N277);
and AND2 (N578, N575, N438);
nand NAND2 (N579, N568, N415);
and AND3 (N580, N574, N179, N442);
xor XOR2 (N581, N561, N449);
buf BUF1 (N582, N580);
xor XOR2 (N583, N581, N548);
xor XOR2 (N584, N582, N437);
xor XOR2 (N585, N584, N327);
not NOT1 (N586, N578);
nand NAND4 (N587, N567, N348, N525, N426);
or OR2 (N588, N587, N7);
nand NAND2 (N589, N586, N394);
or OR3 (N590, N583, N388, N295);
nand NAND2 (N591, N585, N72);
buf BUF1 (N592, N576);
nand NAND3 (N593, N571, N65, N119);
not NOT1 (N594, N590);
nor NOR2 (N595, N592, N354);
buf BUF1 (N596, N593);
buf BUF1 (N597, N591);
buf BUF1 (N598, N594);
xor XOR2 (N599, N597, N555);
not NOT1 (N600, N589);
nand NAND4 (N601, N588, N119, N416, N518);
nand NAND3 (N602, N600, N218, N213);
nor NOR3 (N603, N579, N178, N168);
or OR2 (N604, N595, N584);
buf BUF1 (N605, N596);
buf BUF1 (N606, N601);
buf BUF1 (N607, N606);
or OR2 (N608, N565, N444);
or OR2 (N609, N599, N370);
buf BUF1 (N610, N605);
nand NAND4 (N611, N607, N173, N486, N51);
buf BUF1 (N612, N609);
xor XOR2 (N613, N570, N228);
and AND2 (N614, N603, N78);
xor XOR2 (N615, N598, N53);
nand NAND3 (N616, N614, N294, N574);
buf BUF1 (N617, N613);
nand NAND4 (N618, N602, N78, N74, N219);
xor XOR2 (N619, N616, N501);
xor XOR2 (N620, N618, N121);
or OR3 (N621, N608, N379, N299);
not NOT1 (N622, N577);
xor XOR2 (N623, N620, N122);
nor NOR4 (N624, N622, N376, N444, N288);
xor XOR2 (N625, N624, N361);
not NOT1 (N626, N612);
not NOT1 (N627, N626);
nor NOR4 (N628, N611, N306, N536, N469);
buf BUF1 (N629, N619);
buf BUF1 (N630, N627);
nand NAND3 (N631, N610, N101, N595);
and AND2 (N632, N628, N199);
and AND4 (N633, N615, N116, N263, N357);
xor XOR2 (N634, N632, N273);
buf BUF1 (N635, N630);
xor XOR2 (N636, N617, N148);
buf BUF1 (N637, N636);
nand NAND4 (N638, N625, N299, N52, N398);
and AND4 (N639, N638, N428, N593, N463);
or OR3 (N640, N631, N567, N612);
or OR2 (N641, N639, N299);
xor XOR2 (N642, N634, N608);
not NOT1 (N643, N633);
buf BUF1 (N644, N604);
and AND3 (N645, N640, N458, N563);
xor XOR2 (N646, N623, N325);
nand NAND4 (N647, N641, N577, N461, N233);
xor XOR2 (N648, N646, N592);
xor XOR2 (N649, N645, N532);
and AND2 (N650, N642, N253);
xor XOR2 (N651, N649, N223);
xor XOR2 (N652, N643, N181);
buf BUF1 (N653, N644);
nand NAND2 (N654, N651, N480);
nand NAND4 (N655, N652, N170, N443, N181);
nand NAND3 (N656, N650, N568, N61);
or OR4 (N657, N635, N79, N128, N354);
nor NOR2 (N658, N637, N422);
or OR2 (N659, N656, N523);
not NOT1 (N660, N659);
and AND2 (N661, N657, N55);
nand NAND4 (N662, N655, N433, N312, N659);
not NOT1 (N663, N662);
and AND2 (N664, N658, N10);
xor XOR2 (N665, N653, N597);
and AND3 (N666, N648, N371, N574);
xor XOR2 (N667, N647, N93);
buf BUF1 (N668, N661);
buf BUF1 (N669, N665);
and AND4 (N670, N629, N244, N407, N134);
or OR3 (N671, N664, N453, N2);
and AND3 (N672, N666, N308, N542);
nand NAND4 (N673, N670, N491, N215, N351);
not NOT1 (N674, N673);
nand NAND4 (N675, N668, N628, N35, N315);
or OR4 (N676, N674, N436, N627, N230);
nor NOR4 (N677, N654, N394, N237, N36);
nor NOR2 (N678, N675, N43);
nor NOR4 (N679, N672, N530, N84, N105);
and AND4 (N680, N676, N170, N245, N550);
or OR3 (N681, N621, N310, N458);
buf BUF1 (N682, N677);
or OR2 (N683, N679, N155);
not NOT1 (N684, N660);
nor NOR2 (N685, N682, N558);
xor XOR2 (N686, N685, N300);
nor NOR2 (N687, N671, N548);
and AND2 (N688, N687, N617);
buf BUF1 (N689, N686);
not NOT1 (N690, N667);
nor NOR4 (N691, N690, N181, N560, N641);
and AND2 (N692, N684, N672);
nor NOR3 (N693, N678, N276, N8);
or OR2 (N694, N691, N84);
xor XOR2 (N695, N663, N681);
or OR4 (N696, N609, N179, N219, N299);
or OR4 (N697, N696, N511, N676, N252);
not NOT1 (N698, N697);
or OR3 (N699, N683, N245, N210);
nand NAND4 (N700, N680, N200, N600, N255);
not NOT1 (N701, N669);
nor NOR4 (N702, N694, N700, N377, N187);
nor NOR4 (N703, N669, N552, N476, N404);
buf BUF1 (N704, N695);
nor NOR3 (N705, N699, N646, N359);
and AND3 (N706, N705, N351, N459);
nor NOR2 (N707, N703, N240);
nand NAND2 (N708, N702, N426);
xor XOR2 (N709, N707, N234);
xor XOR2 (N710, N709, N65);
not NOT1 (N711, N701);
not NOT1 (N712, N708);
not NOT1 (N713, N712);
or OR3 (N714, N713, N481, N22);
xor XOR2 (N715, N693, N227);
xor XOR2 (N716, N706, N193);
and AND2 (N717, N689, N98);
not NOT1 (N718, N711);
nand NAND2 (N719, N717, N563);
and AND2 (N720, N692, N254);
and AND2 (N721, N704, N115);
nor NOR2 (N722, N719, N149);
not NOT1 (N723, N698);
and AND3 (N724, N722, N84, N335);
nand NAND4 (N725, N714, N203, N188, N418);
nand NAND4 (N726, N710, N342, N492, N8);
nand NAND4 (N727, N718, N622, N235, N645);
not NOT1 (N728, N720);
and AND3 (N729, N715, N135, N647);
buf BUF1 (N730, N729);
xor XOR2 (N731, N688, N703);
nand NAND3 (N732, N727, N224, N491);
and AND3 (N733, N732, N272, N695);
xor XOR2 (N734, N725, N14);
xor XOR2 (N735, N724, N25);
not NOT1 (N736, N733);
xor XOR2 (N737, N721, N283);
not NOT1 (N738, N728);
and AND4 (N739, N734, N21, N652, N260);
xor XOR2 (N740, N730, N590);
and AND4 (N741, N740, N500, N192, N341);
or OR2 (N742, N723, N478);
nor NOR4 (N743, N716, N209, N657, N42);
xor XOR2 (N744, N735, N688);
xor XOR2 (N745, N736, N167);
nand NAND2 (N746, N742, N155);
xor XOR2 (N747, N741, N604);
nand NAND3 (N748, N745, N554, N426);
and AND3 (N749, N748, N604, N643);
and AND4 (N750, N739, N735, N205, N188);
buf BUF1 (N751, N749);
nand NAND3 (N752, N738, N741, N337);
buf BUF1 (N753, N751);
and AND3 (N754, N744, N655, N151);
buf BUF1 (N755, N737);
and AND4 (N756, N753, N208, N636, N710);
buf BUF1 (N757, N731);
nand NAND3 (N758, N746, N752, N122);
nor NOR4 (N759, N738, N708, N563, N369);
xor XOR2 (N760, N754, N161);
not NOT1 (N761, N756);
not NOT1 (N762, N759);
and AND4 (N763, N761, N676, N293, N70);
nand NAND2 (N764, N726, N291);
or OR2 (N765, N762, N451);
and AND4 (N766, N747, N738, N639, N385);
buf BUF1 (N767, N764);
or OR4 (N768, N765, N658, N505, N598);
and AND2 (N769, N766, N66);
not NOT1 (N770, N750);
or OR2 (N771, N767, N515);
or OR4 (N772, N758, N380, N727, N197);
or OR3 (N773, N768, N267, N604);
buf BUF1 (N774, N743);
or OR4 (N775, N763, N695, N419, N379);
nand NAND4 (N776, N769, N203, N370, N427);
or OR4 (N777, N776, N104, N678, N750);
not NOT1 (N778, N771);
xor XOR2 (N779, N770, N461);
nand NAND3 (N780, N773, N471, N684);
or OR3 (N781, N778, N492, N141);
and AND4 (N782, N777, N467, N286, N716);
and AND2 (N783, N772, N521);
nor NOR3 (N784, N781, N2, N307);
or OR2 (N785, N775, N244);
not NOT1 (N786, N780);
buf BUF1 (N787, N774);
xor XOR2 (N788, N779, N321);
not NOT1 (N789, N783);
or OR4 (N790, N757, N543, N164, N526);
xor XOR2 (N791, N787, N709);
and AND2 (N792, N760, N250);
xor XOR2 (N793, N782, N688);
or OR4 (N794, N792, N578, N103, N760);
nand NAND4 (N795, N784, N562, N673, N653);
nand NAND3 (N796, N790, N369, N387);
xor XOR2 (N797, N796, N374);
buf BUF1 (N798, N794);
not NOT1 (N799, N795);
or OR3 (N800, N788, N447, N251);
nor NOR2 (N801, N789, N420);
nand NAND2 (N802, N791, N446);
buf BUF1 (N803, N793);
xor XOR2 (N804, N755, N70);
xor XOR2 (N805, N804, N550);
nor NOR3 (N806, N801, N528, N148);
buf BUF1 (N807, N802);
xor XOR2 (N808, N786, N688);
nor NOR4 (N809, N803, N251, N763, N673);
nor NOR3 (N810, N797, N494, N543);
and AND3 (N811, N799, N746, N698);
nand NAND3 (N812, N785, N405, N232);
nand NAND3 (N813, N805, N312, N476);
and AND4 (N814, N809, N9, N301, N539);
not NOT1 (N815, N810);
buf BUF1 (N816, N815);
buf BUF1 (N817, N814);
or OR4 (N818, N811, N816, N666, N654);
nand NAND2 (N819, N590, N256);
nand NAND4 (N820, N798, N117, N204, N289);
and AND4 (N821, N807, N280, N486, N111);
buf BUF1 (N822, N813);
and AND4 (N823, N820, N464, N155, N635);
buf BUF1 (N824, N812);
not NOT1 (N825, N819);
or OR2 (N826, N817, N781);
buf BUF1 (N827, N821);
and AND3 (N828, N808, N400, N657);
nor NOR4 (N829, N806, N470, N147, N740);
nor NOR2 (N830, N829, N719);
xor XOR2 (N831, N825, N204);
not NOT1 (N832, N822);
or OR2 (N833, N831, N659);
buf BUF1 (N834, N827);
or OR2 (N835, N828, N382);
buf BUF1 (N836, N830);
nor NOR4 (N837, N836, N322, N511, N468);
nand NAND4 (N838, N826, N17, N33, N837);
not NOT1 (N839, N456);
nand NAND3 (N840, N824, N532, N221);
and AND3 (N841, N800, N514, N308);
xor XOR2 (N842, N823, N4);
nor NOR4 (N843, N842, N339, N659, N23);
nand NAND2 (N844, N841, N652);
and AND3 (N845, N832, N664, N111);
or OR3 (N846, N840, N420, N74);
buf BUF1 (N847, N818);
nor NOR2 (N848, N834, N718);
buf BUF1 (N849, N843);
buf BUF1 (N850, N847);
nor NOR2 (N851, N845, N59);
and AND4 (N852, N838, N742, N755, N755);
xor XOR2 (N853, N835, N220);
xor XOR2 (N854, N853, N246);
nand NAND3 (N855, N852, N280, N249);
buf BUF1 (N856, N846);
xor XOR2 (N857, N844, N521);
buf BUF1 (N858, N851);
or OR2 (N859, N856, N197);
nor NOR4 (N860, N855, N273, N424, N447);
nor NOR4 (N861, N839, N562, N701, N260);
buf BUF1 (N862, N849);
not NOT1 (N863, N858);
or OR4 (N864, N863, N524, N164, N294);
buf BUF1 (N865, N848);
nand NAND4 (N866, N864, N380, N588, N858);
and AND3 (N867, N861, N328, N519);
or OR4 (N868, N854, N519, N566, N131);
or OR4 (N869, N865, N750, N643, N14);
or OR3 (N870, N850, N860, N37);
not NOT1 (N871, N258);
nor NOR4 (N872, N869, N343, N838, N474);
nor NOR3 (N873, N872, N600, N658);
buf BUF1 (N874, N833);
nor NOR3 (N875, N874, N675, N519);
or OR3 (N876, N870, N203, N534);
nor NOR4 (N877, N876, N21, N209, N144);
nand NAND4 (N878, N868, N311, N503, N703);
xor XOR2 (N879, N871, N768);
nand NAND4 (N880, N862, N261, N698, N145);
and AND4 (N881, N877, N364, N12, N66);
nor NOR4 (N882, N880, N807, N32, N415);
xor XOR2 (N883, N867, N93);
xor XOR2 (N884, N857, N668);
not NOT1 (N885, N881);
nand NAND3 (N886, N873, N578, N672);
nand NAND2 (N887, N882, N14);
not NOT1 (N888, N885);
nand NAND4 (N889, N866, N177, N86, N727);
nand NAND3 (N890, N884, N418, N65);
nand NAND2 (N891, N879, N583);
xor XOR2 (N892, N891, N260);
nand NAND4 (N893, N878, N106, N294, N212);
nor NOR3 (N894, N875, N563, N690);
or OR3 (N895, N886, N482, N243);
buf BUF1 (N896, N883);
not NOT1 (N897, N887);
xor XOR2 (N898, N888, N344);
or OR2 (N899, N892, N748);
not NOT1 (N900, N896);
or OR2 (N901, N859, N42);
xor XOR2 (N902, N899, N671);
not NOT1 (N903, N895);
nand NAND4 (N904, N901, N172, N741, N146);
not NOT1 (N905, N902);
xor XOR2 (N906, N904, N546);
and AND3 (N907, N889, N813, N573);
not NOT1 (N908, N894);
or OR2 (N909, N900, N455);
and AND3 (N910, N909, N43, N719);
not NOT1 (N911, N908);
xor XOR2 (N912, N906, N294);
buf BUF1 (N913, N912);
and AND4 (N914, N897, N346, N629, N405);
nor NOR4 (N915, N903, N901, N380, N481);
xor XOR2 (N916, N890, N574);
and AND2 (N917, N905, N518);
xor XOR2 (N918, N907, N173);
nor NOR3 (N919, N913, N245, N97);
nand NAND4 (N920, N893, N544, N99, N324);
and AND3 (N921, N915, N444, N794);
xor XOR2 (N922, N918, N204);
xor XOR2 (N923, N917, N766);
buf BUF1 (N924, N923);
not NOT1 (N925, N920);
nor NOR3 (N926, N910, N12, N207);
buf BUF1 (N927, N916);
nor NOR3 (N928, N919, N16, N79);
buf BUF1 (N929, N924);
and AND2 (N930, N911, N780);
or OR2 (N931, N922, N817);
xor XOR2 (N932, N930, N881);
and AND2 (N933, N914, N814);
buf BUF1 (N934, N927);
nand NAND4 (N935, N928, N843, N524, N916);
not NOT1 (N936, N925);
xor XOR2 (N937, N926, N122);
and AND2 (N938, N937, N751);
and AND2 (N939, N929, N885);
xor XOR2 (N940, N898, N897);
nand NAND3 (N941, N936, N782, N914);
nor NOR4 (N942, N938, N522, N323, N52);
and AND2 (N943, N931, N334);
or OR4 (N944, N939, N312, N33, N805);
buf BUF1 (N945, N943);
or OR3 (N946, N945, N289, N170);
nor NOR3 (N947, N932, N712, N838);
xor XOR2 (N948, N942, N35);
buf BUF1 (N949, N933);
nand NAND2 (N950, N940, N332);
buf BUF1 (N951, N950);
xor XOR2 (N952, N941, N65);
xor XOR2 (N953, N949, N350);
nor NOR3 (N954, N947, N821, N194);
xor XOR2 (N955, N952, N143);
nor NOR2 (N956, N955, N307);
and AND2 (N957, N954, N886);
not NOT1 (N958, N944);
nand NAND2 (N959, N957, N929);
xor XOR2 (N960, N953, N252);
nor NOR4 (N961, N935, N748, N530, N168);
nand NAND4 (N962, N946, N722, N351, N450);
buf BUF1 (N963, N961);
not NOT1 (N964, N956);
nand NAND2 (N965, N963, N57);
and AND4 (N966, N948, N856, N272, N339);
nor NOR4 (N967, N964, N239, N622, N123);
buf BUF1 (N968, N959);
xor XOR2 (N969, N958, N321);
and AND3 (N970, N968, N181, N267);
xor XOR2 (N971, N969, N52);
or OR3 (N972, N965, N293, N48);
nand NAND3 (N973, N967, N325, N331);
nor NOR2 (N974, N934, N734);
and AND4 (N975, N970, N118, N578, N477);
or OR2 (N976, N974, N555);
nor NOR4 (N977, N971, N950, N934, N843);
and AND4 (N978, N921, N382, N235, N807);
nand NAND4 (N979, N951, N546, N804, N68);
xor XOR2 (N980, N975, N935);
not NOT1 (N981, N977);
or OR4 (N982, N966, N347, N930, N679);
or OR4 (N983, N981, N660, N646, N977);
not NOT1 (N984, N982);
nand NAND3 (N985, N976, N381, N135);
buf BUF1 (N986, N985);
xor XOR2 (N987, N960, N731);
or OR4 (N988, N984, N13, N177, N695);
buf BUF1 (N989, N962);
nor NOR4 (N990, N986, N706, N521, N496);
nand NAND3 (N991, N987, N23, N842);
nand NAND3 (N992, N988, N207, N334);
nor NOR3 (N993, N979, N98, N426);
buf BUF1 (N994, N991);
or OR3 (N995, N973, N835, N133);
xor XOR2 (N996, N994, N649);
nor NOR2 (N997, N992, N577);
not NOT1 (N998, N978);
nor NOR3 (N999, N997, N639, N818);
nand NAND4 (N1000, N996, N28, N330, N280);
nor NOR2 (N1001, N989, N241);
xor XOR2 (N1002, N993, N787);
buf BUF1 (N1003, N990);
xor XOR2 (N1004, N983, N260);
xor XOR2 (N1005, N980, N546);
not NOT1 (N1006, N999);
buf BUF1 (N1007, N995);
or OR2 (N1008, N1005, N897);
nor NOR3 (N1009, N998, N868, N888);
nand NAND4 (N1010, N972, N970, N923, N116);
not NOT1 (N1011, N1009);
not NOT1 (N1012, N1001);
and AND2 (N1013, N1002, N20);
nand NAND4 (N1014, N1006, N835, N214, N99);
or OR2 (N1015, N1012, N933);
xor XOR2 (N1016, N1010, N903);
and AND3 (N1017, N1016, N779, N536);
buf BUF1 (N1018, N1013);
xor XOR2 (N1019, N1007, N812);
nor NOR4 (N1020, N1018, N491, N474, N643);
nor NOR4 (N1021, N1020, N805, N748, N872);
buf BUF1 (N1022, N1019);
or OR2 (N1023, N1008, N244);
or OR3 (N1024, N1000, N298, N514);
xor XOR2 (N1025, N1023, N603);
nand NAND4 (N1026, N1015, N276, N432, N894);
nand NAND3 (N1027, N1024, N309, N790);
xor XOR2 (N1028, N1026, N880);
nand NAND3 (N1029, N1011, N294, N415);
not NOT1 (N1030, N1014);
nand NAND3 (N1031, N1030, N545, N402);
nor NOR3 (N1032, N1027, N769, N497);
and AND3 (N1033, N1029, N887, N1002);
buf BUF1 (N1034, N1025);
nor NOR4 (N1035, N1017, N1025, N152, N480);
not NOT1 (N1036, N1003);
nand NAND3 (N1037, N1028, N921, N299);
xor XOR2 (N1038, N1034, N869);
or OR2 (N1039, N1038, N1036);
or OR3 (N1040, N958, N1033, N974);
nor NOR3 (N1041, N209, N240, N176);
xor XOR2 (N1042, N1041, N749);
not NOT1 (N1043, N1039);
not NOT1 (N1044, N1031);
buf BUF1 (N1045, N1044);
nand NAND3 (N1046, N1004, N1028, N1);
nor NOR3 (N1047, N1040, N4, N348);
nand NAND3 (N1048, N1035, N810, N390);
nand NAND3 (N1049, N1045, N1024, N1034);
buf BUF1 (N1050, N1047);
and AND2 (N1051, N1037, N299);
buf BUF1 (N1052, N1048);
and AND3 (N1053, N1050, N469, N104);
buf BUF1 (N1054, N1049);
nor NOR4 (N1055, N1053, N412, N324, N863);
buf BUF1 (N1056, N1021);
not NOT1 (N1057, N1054);
nor NOR3 (N1058, N1057, N876, N144);
buf BUF1 (N1059, N1032);
or OR3 (N1060, N1055, N437, N643);
and AND4 (N1061, N1022, N905, N1030, N176);
or OR2 (N1062, N1043, N776);
xor XOR2 (N1063, N1056, N641);
not NOT1 (N1064, N1062);
xor XOR2 (N1065, N1042, N452);
xor XOR2 (N1066, N1061, N171);
and AND2 (N1067, N1064, N1019);
xor XOR2 (N1068, N1051, N545);
nand NAND3 (N1069, N1066, N485, N136);
nor NOR4 (N1070, N1046, N989, N156, N1027);
not NOT1 (N1071, N1059);
or OR3 (N1072, N1068, N39, N300);
and AND4 (N1073, N1058, N177, N358, N322);
buf BUF1 (N1074, N1065);
buf BUF1 (N1075, N1074);
and AND4 (N1076, N1063, N48, N856, N644);
not NOT1 (N1077, N1067);
or OR4 (N1078, N1052, N117, N894, N491);
xor XOR2 (N1079, N1069, N411);
buf BUF1 (N1080, N1075);
and AND2 (N1081, N1071, N269);
or OR2 (N1082, N1080, N587);
or OR2 (N1083, N1081, N505);
buf BUF1 (N1084, N1070);
and AND4 (N1085, N1083, N590, N431, N345);
or OR2 (N1086, N1072, N278);
nor NOR3 (N1087, N1084, N240, N69);
or OR2 (N1088, N1076, N342);
xor XOR2 (N1089, N1088, N518);
not NOT1 (N1090, N1079);
and AND4 (N1091, N1085, N967, N425, N568);
and AND2 (N1092, N1077, N474);
not NOT1 (N1093, N1089);
nand NAND3 (N1094, N1082, N1064, N974);
buf BUF1 (N1095, N1073);
or OR4 (N1096, N1060, N181, N422, N37);
nand NAND4 (N1097, N1092, N742, N42, N751);
not NOT1 (N1098, N1087);
nor NOR3 (N1099, N1093, N911, N869);
and AND2 (N1100, N1096, N485);
nand NAND4 (N1101, N1091, N909, N896, N58);
buf BUF1 (N1102, N1100);
and AND4 (N1103, N1099, N784, N13, N661);
and AND2 (N1104, N1098, N820);
xor XOR2 (N1105, N1101, N126);
xor XOR2 (N1106, N1095, N976);
nor NOR2 (N1107, N1104, N257);
xor XOR2 (N1108, N1097, N156);
or OR3 (N1109, N1108, N126, N1);
and AND2 (N1110, N1086, N578);
nand NAND3 (N1111, N1078, N742, N632);
nor NOR2 (N1112, N1103, N604);
nand NAND3 (N1113, N1105, N612, N428);
or OR4 (N1114, N1106, N989, N10, N297);
xor XOR2 (N1115, N1107, N1067);
or OR3 (N1116, N1094, N580, N848);
buf BUF1 (N1117, N1112);
nand NAND4 (N1118, N1116, N762, N992, N827);
nand NAND2 (N1119, N1114, N1051);
buf BUF1 (N1120, N1111);
and AND2 (N1121, N1102, N629);
nor NOR4 (N1122, N1120, N883, N118, N325);
or OR2 (N1123, N1113, N1033);
not NOT1 (N1124, N1119);
nand NAND4 (N1125, N1121, N758, N723, N775);
nor NOR4 (N1126, N1122, N644, N1023, N586);
xor XOR2 (N1127, N1123, N511);
buf BUF1 (N1128, N1117);
not NOT1 (N1129, N1115);
and AND2 (N1130, N1090, N426);
and AND2 (N1131, N1128, N1037);
xor XOR2 (N1132, N1125, N921);
xor XOR2 (N1133, N1130, N617);
or OR2 (N1134, N1132, N48);
buf BUF1 (N1135, N1133);
xor XOR2 (N1136, N1109, N341);
or OR2 (N1137, N1131, N484);
nand NAND3 (N1138, N1135, N830, N403);
xor XOR2 (N1139, N1124, N15);
and AND4 (N1140, N1110, N1134, N1075, N1100);
buf BUF1 (N1141, N22);
and AND2 (N1142, N1140, N596);
and AND4 (N1143, N1139, N25, N906, N428);
buf BUF1 (N1144, N1137);
nor NOR3 (N1145, N1144, N1073, N397);
buf BUF1 (N1146, N1129);
nor NOR2 (N1147, N1146, N799);
and AND2 (N1148, N1127, N1032);
buf BUF1 (N1149, N1141);
nand NAND3 (N1150, N1138, N139, N949);
nor NOR3 (N1151, N1148, N977, N196);
and AND4 (N1152, N1118, N886, N517, N408);
xor XOR2 (N1153, N1142, N162);
not NOT1 (N1154, N1143);
nand NAND2 (N1155, N1145, N836);
or OR3 (N1156, N1152, N443, N342);
not NOT1 (N1157, N1154);
xor XOR2 (N1158, N1150, N1016);
nand NAND2 (N1159, N1153, N984);
nand NAND2 (N1160, N1126, N630);
buf BUF1 (N1161, N1159);
nor NOR4 (N1162, N1149, N85, N716, N986);
and AND3 (N1163, N1151, N521, N171);
buf BUF1 (N1164, N1163);
not NOT1 (N1165, N1156);
nand NAND2 (N1166, N1160, N949);
and AND3 (N1167, N1158, N584, N942);
nand NAND4 (N1168, N1164, N821, N795, N1136);
xor XOR2 (N1169, N639, N807);
not NOT1 (N1170, N1147);
not NOT1 (N1171, N1168);
nor NOR4 (N1172, N1165, N974, N990, N510);
not NOT1 (N1173, N1170);
nand NAND4 (N1174, N1157, N612, N947, N1146);
and AND2 (N1175, N1161, N187);
or OR3 (N1176, N1166, N562, N1057);
xor XOR2 (N1177, N1169, N296);
and AND2 (N1178, N1162, N372);
or OR2 (N1179, N1178, N469);
nor NOR3 (N1180, N1175, N547, N122);
nor NOR2 (N1181, N1180, N367);
buf BUF1 (N1182, N1155);
nor NOR4 (N1183, N1167, N287, N625, N699);
not NOT1 (N1184, N1183);
or OR2 (N1185, N1177, N777);
not NOT1 (N1186, N1184);
or OR2 (N1187, N1186, N277);
or OR3 (N1188, N1172, N1065, N8);
nor NOR4 (N1189, N1171, N1003, N148, N191);
and AND4 (N1190, N1182, N473, N1180, N287);
not NOT1 (N1191, N1179);
nand NAND4 (N1192, N1185, N1171, N763, N885);
or OR2 (N1193, N1191, N220);
nand NAND3 (N1194, N1176, N1052, N490);
xor XOR2 (N1195, N1187, N845);
and AND3 (N1196, N1188, N46, N12);
and AND2 (N1197, N1192, N636);
or OR2 (N1198, N1181, N1008);
or OR4 (N1199, N1193, N293, N480, N928);
xor XOR2 (N1200, N1196, N669);
nand NAND4 (N1201, N1200, N994, N233, N882);
and AND2 (N1202, N1189, N797);
and AND4 (N1203, N1198, N252, N387, N747);
nor NOR4 (N1204, N1174, N858, N870, N702);
and AND4 (N1205, N1199, N841, N1199, N260);
nand NAND3 (N1206, N1205, N574, N287);
nand NAND4 (N1207, N1206, N683, N1001, N622);
nand NAND4 (N1208, N1204, N205, N1080, N654);
buf BUF1 (N1209, N1202);
not NOT1 (N1210, N1197);
xor XOR2 (N1211, N1194, N1081);
or OR3 (N1212, N1190, N856, N340);
not NOT1 (N1213, N1211);
or OR3 (N1214, N1213, N361, N137);
not NOT1 (N1215, N1207);
nand NAND3 (N1216, N1209, N886, N908);
nor NOR3 (N1217, N1212, N836, N286);
nor NOR3 (N1218, N1210, N556, N691);
nor NOR2 (N1219, N1201, N1156);
xor XOR2 (N1220, N1203, N342);
and AND4 (N1221, N1208, N13, N533, N524);
buf BUF1 (N1222, N1215);
buf BUF1 (N1223, N1219);
not NOT1 (N1224, N1217);
xor XOR2 (N1225, N1214, N287);
nand NAND4 (N1226, N1222, N1185, N751, N217);
nand NAND2 (N1227, N1224, N23);
xor XOR2 (N1228, N1220, N42);
or OR2 (N1229, N1218, N890);
and AND2 (N1230, N1195, N686);
buf BUF1 (N1231, N1227);
xor XOR2 (N1232, N1228, N714);
xor XOR2 (N1233, N1229, N805);
not NOT1 (N1234, N1173);
buf BUF1 (N1235, N1234);
nor NOR4 (N1236, N1235, N142, N483, N1014);
nor NOR3 (N1237, N1221, N1141, N163);
xor XOR2 (N1238, N1225, N329);
nand NAND4 (N1239, N1230, N1211, N779, N593);
buf BUF1 (N1240, N1239);
not NOT1 (N1241, N1237);
buf BUF1 (N1242, N1226);
not NOT1 (N1243, N1223);
xor XOR2 (N1244, N1236, N1014);
and AND2 (N1245, N1238, N1019);
buf BUF1 (N1246, N1233);
not NOT1 (N1247, N1240);
xor XOR2 (N1248, N1216, N842);
or OR4 (N1249, N1242, N801, N870, N461);
and AND3 (N1250, N1231, N1115, N577);
or OR3 (N1251, N1243, N1130, N403);
and AND4 (N1252, N1245, N401, N780, N38);
xor XOR2 (N1253, N1251, N1231);
nor NOR2 (N1254, N1244, N1104);
and AND2 (N1255, N1246, N1069);
or OR2 (N1256, N1253, N842);
not NOT1 (N1257, N1241);
not NOT1 (N1258, N1232);
nor NOR3 (N1259, N1254, N1179, N538);
nor NOR2 (N1260, N1255, N824);
nor NOR4 (N1261, N1259, N617, N263, N51);
not NOT1 (N1262, N1256);
not NOT1 (N1263, N1262);
xor XOR2 (N1264, N1260, N1203);
buf BUF1 (N1265, N1263);
not NOT1 (N1266, N1249);
not NOT1 (N1267, N1247);
or OR2 (N1268, N1250, N390);
and AND3 (N1269, N1252, N457, N953);
nor NOR2 (N1270, N1266, N238);
xor XOR2 (N1271, N1269, N1098);
buf BUF1 (N1272, N1257);
nand NAND3 (N1273, N1268, N595, N141);
xor XOR2 (N1274, N1273, N993);
and AND4 (N1275, N1272, N1207, N313, N1020);
xor XOR2 (N1276, N1261, N1185);
xor XOR2 (N1277, N1274, N1196);
or OR3 (N1278, N1271, N569, N255);
xor XOR2 (N1279, N1270, N548);
or OR2 (N1280, N1267, N278);
xor XOR2 (N1281, N1258, N768);
or OR4 (N1282, N1275, N120, N110, N505);
or OR4 (N1283, N1276, N647, N186, N849);
not NOT1 (N1284, N1279);
nand NAND3 (N1285, N1283, N1041, N581);
nand NAND4 (N1286, N1284, N935, N1077, N604);
xor XOR2 (N1287, N1264, N821);
nand NAND2 (N1288, N1278, N272);
nand NAND2 (N1289, N1277, N892);
nor NOR2 (N1290, N1281, N1220);
not NOT1 (N1291, N1265);
nor NOR4 (N1292, N1288, N683, N750, N289);
xor XOR2 (N1293, N1286, N144);
and AND4 (N1294, N1289, N105, N89, N111);
buf BUF1 (N1295, N1280);
xor XOR2 (N1296, N1282, N306);
xor XOR2 (N1297, N1287, N558);
or OR3 (N1298, N1296, N366, N1289);
and AND3 (N1299, N1285, N229, N532);
nand NAND2 (N1300, N1295, N526);
not NOT1 (N1301, N1293);
nand NAND4 (N1302, N1292, N585, N338, N647);
not NOT1 (N1303, N1290);
not NOT1 (N1304, N1298);
nor NOR4 (N1305, N1304, N222, N978, N1255);
and AND3 (N1306, N1291, N274, N274);
xor XOR2 (N1307, N1305, N768);
or OR2 (N1308, N1301, N688);
and AND2 (N1309, N1294, N386);
and AND3 (N1310, N1303, N672, N860);
nand NAND3 (N1311, N1306, N391, N740);
nor NOR3 (N1312, N1299, N740, N1166);
nor NOR3 (N1313, N1307, N388, N751);
not NOT1 (N1314, N1302);
nand NAND2 (N1315, N1248, N1074);
buf BUF1 (N1316, N1297);
nand NAND3 (N1317, N1315, N823, N724);
nand NAND4 (N1318, N1308, N200, N179, N734);
nand NAND2 (N1319, N1317, N94);
nor NOR4 (N1320, N1319, N698, N871, N444);
and AND3 (N1321, N1313, N809, N302);
xor XOR2 (N1322, N1314, N369);
buf BUF1 (N1323, N1309);
xor XOR2 (N1324, N1310, N568);
nand NAND2 (N1325, N1311, N1080);
buf BUF1 (N1326, N1300);
or OR3 (N1327, N1323, N1324, N38);
and AND3 (N1328, N100, N184, N289);
xor XOR2 (N1329, N1327, N610);
nor NOR2 (N1330, N1329, N994);
nor NOR3 (N1331, N1312, N769, N1107);
nand NAND2 (N1332, N1331, N382);
buf BUF1 (N1333, N1320);
buf BUF1 (N1334, N1333);
nor NOR3 (N1335, N1321, N138, N1105);
and AND4 (N1336, N1325, N228, N565, N1169);
buf BUF1 (N1337, N1318);
nand NAND3 (N1338, N1328, N1164, N731);
nand NAND2 (N1339, N1326, N732);
or OR4 (N1340, N1339, N474, N129, N724);
xor XOR2 (N1341, N1330, N525);
nand NAND3 (N1342, N1316, N690, N1324);
not NOT1 (N1343, N1338);
and AND3 (N1344, N1337, N1040, N1172);
or OR4 (N1345, N1332, N423, N1330, N1212);
nand NAND2 (N1346, N1342, N1012);
not NOT1 (N1347, N1336);
or OR2 (N1348, N1347, N651);
buf BUF1 (N1349, N1343);
nand NAND4 (N1350, N1335, N3, N1112, N699);
not NOT1 (N1351, N1344);
nand NAND4 (N1352, N1322, N619, N377, N697);
nor NOR3 (N1353, N1348, N1300, N903);
nand NAND3 (N1354, N1353, N1023, N439);
nand NAND4 (N1355, N1354, N205, N152, N1028);
and AND3 (N1356, N1355, N305, N438);
or OR4 (N1357, N1349, N926, N1099, N899);
nor NOR3 (N1358, N1334, N629, N201);
buf BUF1 (N1359, N1357);
nor NOR4 (N1360, N1346, N1274, N169, N1332);
or OR3 (N1361, N1356, N647, N613);
xor XOR2 (N1362, N1360, N699);
nand NAND3 (N1363, N1361, N1122, N990);
buf BUF1 (N1364, N1352);
not NOT1 (N1365, N1350);
nand NAND2 (N1366, N1362, N1024);
or OR2 (N1367, N1366, N112);
and AND2 (N1368, N1359, N978);
buf BUF1 (N1369, N1363);
buf BUF1 (N1370, N1340);
buf BUF1 (N1371, N1341);
nor NOR3 (N1372, N1371, N154, N246);
nor NOR3 (N1373, N1368, N160, N984);
nand NAND4 (N1374, N1351, N859, N962, N299);
not NOT1 (N1375, N1345);
nor NOR3 (N1376, N1369, N1188, N621);
nand NAND2 (N1377, N1376, N244);
nor NOR3 (N1378, N1358, N245, N203);
xor XOR2 (N1379, N1370, N768);
xor XOR2 (N1380, N1364, N304);
nor NOR4 (N1381, N1379, N471, N771, N496);
nor NOR4 (N1382, N1375, N1123, N809, N905);
not NOT1 (N1383, N1381);
not NOT1 (N1384, N1373);
nand NAND3 (N1385, N1384, N1034, N1134);
or OR4 (N1386, N1367, N454, N776, N829);
buf BUF1 (N1387, N1372);
nor NOR3 (N1388, N1386, N857, N1203);
nor NOR3 (N1389, N1387, N668, N248);
and AND4 (N1390, N1385, N1023, N1367, N1205);
buf BUF1 (N1391, N1382);
xor XOR2 (N1392, N1378, N255);
and AND3 (N1393, N1390, N998, N1374);
nand NAND3 (N1394, N1379, N784, N730);
not NOT1 (N1395, N1394);
not NOT1 (N1396, N1377);
not NOT1 (N1397, N1395);
nand NAND3 (N1398, N1396, N829, N1305);
nand NAND4 (N1399, N1383, N1286, N963, N659);
or OR4 (N1400, N1380, N852, N322, N686);
and AND2 (N1401, N1389, N433);
not NOT1 (N1402, N1365);
or OR4 (N1403, N1397, N927, N177, N37);
nand NAND2 (N1404, N1392, N371);
nand NAND4 (N1405, N1398, N658, N1018, N11);
and AND3 (N1406, N1404, N1120, N949);
not NOT1 (N1407, N1402);
not NOT1 (N1408, N1405);
buf BUF1 (N1409, N1399);
and AND4 (N1410, N1388, N1084, N283, N1298);
and AND3 (N1411, N1407, N783, N30);
buf BUF1 (N1412, N1401);
xor XOR2 (N1413, N1393, N347);
xor XOR2 (N1414, N1391, N189);
buf BUF1 (N1415, N1412);
or OR3 (N1416, N1415, N1187, N1134);
buf BUF1 (N1417, N1410);
nor NOR4 (N1418, N1417, N514, N1140, N1069);
nand NAND4 (N1419, N1409, N169, N1286, N103);
xor XOR2 (N1420, N1403, N1344);
xor XOR2 (N1421, N1413, N587);
xor XOR2 (N1422, N1418, N874);
not NOT1 (N1423, N1408);
or OR3 (N1424, N1419, N1144, N873);
not NOT1 (N1425, N1416);
and AND4 (N1426, N1406, N301, N384, N97);
not NOT1 (N1427, N1400);
buf BUF1 (N1428, N1421);
buf BUF1 (N1429, N1411);
nand NAND3 (N1430, N1427, N1074, N310);
buf BUF1 (N1431, N1420);
and AND2 (N1432, N1426, N497);
buf BUF1 (N1433, N1432);
nand NAND3 (N1434, N1425, N1118, N497);
nor NOR3 (N1435, N1428, N1128, N249);
or OR3 (N1436, N1433, N327, N294);
or OR2 (N1437, N1435, N516);
not NOT1 (N1438, N1424);
not NOT1 (N1439, N1438);
not NOT1 (N1440, N1429);
buf BUF1 (N1441, N1422);
nor NOR4 (N1442, N1441, N158, N862, N180);
buf BUF1 (N1443, N1442);
not NOT1 (N1444, N1440);
buf BUF1 (N1445, N1434);
and AND2 (N1446, N1443, N396);
nand NAND3 (N1447, N1444, N947, N96);
nor NOR2 (N1448, N1439, N655);
or OR2 (N1449, N1448, N17);
xor XOR2 (N1450, N1445, N545);
xor XOR2 (N1451, N1414, N363);
nand NAND3 (N1452, N1423, N337, N1309);
buf BUF1 (N1453, N1446);
or OR4 (N1454, N1430, N1357, N808, N1324);
xor XOR2 (N1455, N1454, N1286);
xor XOR2 (N1456, N1431, N211);
nand NAND2 (N1457, N1450, N965);
nand NAND3 (N1458, N1436, N648, N1271);
and AND2 (N1459, N1457, N1167);
not NOT1 (N1460, N1458);
not NOT1 (N1461, N1459);
or OR2 (N1462, N1456, N1078);
xor XOR2 (N1463, N1452, N682);
and AND3 (N1464, N1455, N146, N1072);
nor NOR2 (N1465, N1460, N1152);
nand NAND4 (N1466, N1462, N120, N227, N1238);
buf BUF1 (N1467, N1464);
nor NOR2 (N1468, N1467, N560);
buf BUF1 (N1469, N1461);
nand NAND4 (N1470, N1447, N944, N543, N380);
and AND2 (N1471, N1449, N1311);
not NOT1 (N1472, N1468);
and AND2 (N1473, N1465, N1010);
not NOT1 (N1474, N1471);
not NOT1 (N1475, N1473);
and AND3 (N1476, N1470, N534, N137);
buf BUF1 (N1477, N1466);
and AND2 (N1478, N1474, N1198);
and AND4 (N1479, N1476, N1369, N939, N691);
buf BUF1 (N1480, N1477);
nor NOR3 (N1481, N1479, N215, N543);
and AND2 (N1482, N1475, N749);
and AND3 (N1483, N1478, N1041, N1219);
not NOT1 (N1484, N1483);
or OR4 (N1485, N1469, N1221, N190, N1418);
and AND3 (N1486, N1484, N225, N133);
not NOT1 (N1487, N1453);
nor NOR4 (N1488, N1487, N173, N662, N446);
xor XOR2 (N1489, N1485, N928);
and AND4 (N1490, N1482, N211, N212, N555);
not NOT1 (N1491, N1472);
nor NOR4 (N1492, N1437, N843, N747, N106);
or OR4 (N1493, N1481, N1133, N1231, N1101);
and AND3 (N1494, N1480, N1021, N210);
buf BUF1 (N1495, N1494);
and AND4 (N1496, N1491, N459, N1085, N1160);
or OR2 (N1497, N1451, N811);
nand NAND4 (N1498, N1489, N863, N1009, N477);
xor XOR2 (N1499, N1495, N511);
nor NOR4 (N1500, N1490, N1184, N1101, N159);
and AND2 (N1501, N1492, N502);
or OR4 (N1502, N1500, N1250, N861, N1300);
nand NAND3 (N1503, N1493, N897, N624);
buf BUF1 (N1504, N1497);
not NOT1 (N1505, N1503);
and AND4 (N1506, N1486, N77, N191, N804);
buf BUF1 (N1507, N1463);
and AND3 (N1508, N1505, N842, N1413);
not NOT1 (N1509, N1501);
and AND4 (N1510, N1508, N963, N1411, N26);
nor NOR2 (N1511, N1507, N914);
buf BUF1 (N1512, N1509);
buf BUF1 (N1513, N1502);
buf BUF1 (N1514, N1498);
and AND3 (N1515, N1510, N409, N1251);
buf BUF1 (N1516, N1496);
xor XOR2 (N1517, N1511, N441);
nor NOR2 (N1518, N1515, N785);
nor NOR3 (N1519, N1513, N850, N111);
not NOT1 (N1520, N1512);
and AND4 (N1521, N1488, N959, N1007, N44);
xor XOR2 (N1522, N1506, N760);
xor XOR2 (N1523, N1516, N457);
and AND4 (N1524, N1520, N311, N1424, N1081);
nand NAND2 (N1525, N1514, N333);
or OR3 (N1526, N1523, N1204, N701);
xor XOR2 (N1527, N1525, N476);
not NOT1 (N1528, N1521);
nor NOR2 (N1529, N1517, N1196);
nor NOR4 (N1530, N1504, N1354, N1034, N817);
buf BUF1 (N1531, N1526);
or OR4 (N1532, N1524, N78, N1439, N300);
buf BUF1 (N1533, N1531);
not NOT1 (N1534, N1519);
nor NOR3 (N1535, N1528, N1483, N142);
nand NAND4 (N1536, N1532, N248, N725, N1398);
or OR3 (N1537, N1534, N714, N923);
nand NAND2 (N1538, N1530, N1523);
nor NOR4 (N1539, N1529, N394, N173, N1141);
nor NOR4 (N1540, N1538, N905, N816, N1034);
not NOT1 (N1541, N1522);
nor NOR2 (N1542, N1540, N1465);
nand NAND3 (N1543, N1542, N276, N1255);
buf BUF1 (N1544, N1527);
and AND2 (N1545, N1541, N1129);
nand NAND4 (N1546, N1545, N1164, N1457, N820);
or OR2 (N1547, N1543, N1018);
not NOT1 (N1548, N1537);
or OR2 (N1549, N1499, N1375);
and AND3 (N1550, N1539, N1418, N575);
not NOT1 (N1551, N1549);
buf BUF1 (N1552, N1535);
not NOT1 (N1553, N1552);
nand NAND4 (N1554, N1548, N944, N881, N1040);
nand NAND2 (N1555, N1553, N769);
or OR3 (N1556, N1550, N1176, N1394);
and AND3 (N1557, N1551, N773, N1489);
nand NAND3 (N1558, N1533, N322, N438);
xor XOR2 (N1559, N1556, N297);
or OR2 (N1560, N1555, N848);
not NOT1 (N1561, N1536);
xor XOR2 (N1562, N1561, N1197);
and AND4 (N1563, N1546, N912, N1157, N907);
not NOT1 (N1564, N1560);
or OR3 (N1565, N1554, N1217, N628);
nand NAND4 (N1566, N1518, N231, N1383, N402);
nor NOR3 (N1567, N1563, N352, N813);
nor NOR4 (N1568, N1558, N109, N332, N1081);
or OR4 (N1569, N1547, N503, N1562, N1096);
not NOT1 (N1570, N455);
xor XOR2 (N1571, N1570, N1251);
or OR4 (N1572, N1568, N395, N219, N654);
or OR3 (N1573, N1564, N1021, N1362);
or OR4 (N1574, N1572, N186, N1030, N1327);
or OR2 (N1575, N1569, N127);
not NOT1 (N1576, N1571);
buf BUF1 (N1577, N1575);
not NOT1 (N1578, N1577);
xor XOR2 (N1579, N1557, N541);
nor NOR3 (N1580, N1574, N1005, N765);
nand NAND3 (N1581, N1559, N1148, N1171);
xor XOR2 (N1582, N1581, N736);
and AND3 (N1583, N1544, N996, N998);
buf BUF1 (N1584, N1565);
nor NOR2 (N1585, N1566, N1002);
or OR4 (N1586, N1585, N173, N1330, N541);
xor XOR2 (N1587, N1567, N65);
nand NAND2 (N1588, N1579, N1356);
xor XOR2 (N1589, N1578, N258);
or OR3 (N1590, N1583, N877, N22);
nor NOR4 (N1591, N1589, N662, N1043, N1504);
xor XOR2 (N1592, N1582, N200);
xor XOR2 (N1593, N1591, N1420);
and AND4 (N1594, N1593, N1577, N615, N198);
nor NOR4 (N1595, N1588, N1, N1097, N568);
and AND3 (N1596, N1587, N335, N512);
and AND2 (N1597, N1573, N643);
not NOT1 (N1598, N1580);
nor NOR3 (N1599, N1594, N416, N554);
not NOT1 (N1600, N1592);
nor NOR3 (N1601, N1586, N999, N468);
not NOT1 (N1602, N1576);
and AND2 (N1603, N1598, N1131);
and AND4 (N1604, N1602, N989, N76, N1512);
buf BUF1 (N1605, N1595);
buf BUF1 (N1606, N1597);
and AND3 (N1607, N1600, N371, N1503);
or OR2 (N1608, N1607, N324);
not NOT1 (N1609, N1605);
nor NOR2 (N1610, N1599, N546);
not NOT1 (N1611, N1604);
xor XOR2 (N1612, N1584, N1534);
or OR3 (N1613, N1608, N60, N1290);
nand NAND2 (N1614, N1596, N1152);
nand NAND2 (N1615, N1611, N534);
xor XOR2 (N1616, N1615, N1484);
nand NAND3 (N1617, N1601, N299, N852);
or OR4 (N1618, N1610, N811, N879, N1258);
nor NOR2 (N1619, N1617, N207);
nor NOR3 (N1620, N1606, N1239, N1266);
buf BUF1 (N1621, N1603);
or OR2 (N1622, N1612, N323);
buf BUF1 (N1623, N1616);
xor XOR2 (N1624, N1614, N439);
xor XOR2 (N1625, N1590, N617);
not NOT1 (N1626, N1622);
not NOT1 (N1627, N1613);
or OR2 (N1628, N1620, N1340);
buf BUF1 (N1629, N1618);
or OR2 (N1630, N1626, N1288);
xor XOR2 (N1631, N1630, N762);
buf BUF1 (N1632, N1628);
buf BUF1 (N1633, N1629);
nor NOR3 (N1634, N1621, N591, N706);
and AND2 (N1635, N1627, N1606);
or OR2 (N1636, N1631, N582);
and AND4 (N1637, N1636, N1304, N1275, N217);
nand NAND4 (N1638, N1634, N181, N1045, N505);
not NOT1 (N1639, N1619);
buf BUF1 (N1640, N1632);
nor NOR3 (N1641, N1639, N378, N263);
nand NAND3 (N1642, N1609, N962, N470);
and AND4 (N1643, N1624, N162, N1587, N974);
not NOT1 (N1644, N1641);
and AND3 (N1645, N1633, N1434, N943);
and AND2 (N1646, N1637, N608);
or OR2 (N1647, N1643, N616);
and AND4 (N1648, N1646, N643, N1491, N870);
xor XOR2 (N1649, N1642, N548);
or OR2 (N1650, N1649, N1571);
not NOT1 (N1651, N1650);
not NOT1 (N1652, N1644);
nand NAND3 (N1653, N1640, N885, N945);
or OR3 (N1654, N1638, N1393, N1485);
not NOT1 (N1655, N1625);
buf BUF1 (N1656, N1654);
nand NAND3 (N1657, N1647, N1286, N281);
nor NOR4 (N1658, N1648, N1570, N393, N72);
xor XOR2 (N1659, N1656, N1120);
or OR3 (N1660, N1655, N689, N186);
buf BUF1 (N1661, N1651);
or OR4 (N1662, N1660, N1289, N343, N1329);
or OR4 (N1663, N1658, N828, N1524, N95);
nor NOR2 (N1664, N1645, N1237);
nand NAND3 (N1665, N1663, N1266, N1146);
nor NOR4 (N1666, N1623, N225, N81, N595);
nor NOR4 (N1667, N1665, N568, N1193, N248);
and AND3 (N1668, N1657, N963, N644);
buf BUF1 (N1669, N1667);
and AND4 (N1670, N1653, N504, N1392, N372);
buf BUF1 (N1671, N1662);
and AND4 (N1672, N1664, N1011, N1128, N906);
or OR4 (N1673, N1672, N87, N331, N230);
xor XOR2 (N1674, N1666, N961);
buf BUF1 (N1675, N1671);
and AND4 (N1676, N1670, N931, N801, N10);
xor XOR2 (N1677, N1661, N1519);
nor NOR4 (N1678, N1668, N1284, N1643, N819);
xor XOR2 (N1679, N1676, N929);
buf BUF1 (N1680, N1673);
nand NAND2 (N1681, N1675, N343);
xor XOR2 (N1682, N1635, N311);
nor NOR2 (N1683, N1680, N23);
not NOT1 (N1684, N1678);
nor NOR4 (N1685, N1684, N418, N253, N1605);
and AND4 (N1686, N1682, N199, N1492, N931);
nor NOR2 (N1687, N1683, N25);
xor XOR2 (N1688, N1679, N901);
and AND2 (N1689, N1685, N127);
nand NAND3 (N1690, N1652, N1439, N1521);
buf BUF1 (N1691, N1690);
nand NAND2 (N1692, N1659, N421);
nor NOR2 (N1693, N1681, N1285);
or OR3 (N1694, N1693, N1691, N1596);
nand NAND4 (N1695, N1276, N1541, N1308, N976);
buf BUF1 (N1696, N1692);
xor XOR2 (N1697, N1686, N323);
not NOT1 (N1698, N1696);
nand NAND2 (N1699, N1695, N771);
xor XOR2 (N1700, N1694, N1250);
and AND3 (N1701, N1699, N1364, N1558);
and AND2 (N1702, N1674, N668);
buf BUF1 (N1703, N1687);
and AND2 (N1704, N1688, N392);
or OR2 (N1705, N1703, N1008);
not NOT1 (N1706, N1700);
buf BUF1 (N1707, N1669);
and AND2 (N1708, N1701, N613);
xor XOR2 (N1709, N1704, N1683);
and AND2 (N1710, N1689, N780);
and AND4 (N1711, N1707, N1115, N1201, N107);
or OR3 (N1712, N1705, N123, N1341);
not NOT1 (N1713, N1697);
nand NAND3 (N1714, N1698, N153, N61);
xor XOR2 (N1715, N1708, N1233);
and AND2 (N1716, N1709, N322);
nor NOR3 (N1717, N1706, N1433, N971);
not NOT1 (N1718, N1712);
xor XOR2 (N1719, N1714, N974);
not NOT1 (N1720, N1710);
buf BUF1 (N1721, N1720);
and AND4 (N1722, N1702, N596, N1627, N11);
and AND4 (N1723, N1721, N876, N170, N1071);
nor NOR4 (N1724, N1713, N939, N87, N875);
or OR3 (N1725, N1719, N1287, N1258);
or OR4 (N1726, N1724, N874, N265, N1040);
buf BUF1 (N1727, N1716);
or OR2 (N1728, N1718, N332);
or OR4 (N1729, N1726, N1515, N912, N1045);
or OR4 (N1730, N1677, N1245, N1439, N222);
or OR2 (N1731, N1729, N212);
or OR2 (N1732, N1728, N670);
xor XOR2 (N1733, N1727, N1334);
and AND2 (N1734, N1725, N1675);
and AND2 (N1735, N1722, N862);
not NOT1 (N1736, N1715);
buf BUF1 (N1737, N1711);
or OR3 (N1738, N1717, N225, N1461);
nor NOR3 (N1739, N1736, N462, N28);
buf BUF1 (N1740, N1733);
and AND4 (N1741, N1735, N925, N1152, N787);
xor XOR2 (N1742, N1741, N106);
buf BUF1 (N1743, N1731);
not NOT1 (N1744, N1737);
not NOT1 (N1745, N1732);
not NOT1 (N1746, N1723);
and AND2 (N1747, N1740, N1508);
xor XOR2 (N1748, N1738, N995);
and AND4 (N1749, N1748, N1433, N1523, N618);
xor XOR2 (N1750, N1739, N1077);
nor NOR4 (N1751, N1747, N1631, N7, N891);
not NOT1 (N1752, N1746);
or OR2 (N1753, N1743, N1687);
or OR2 (N1754, N1752, N621);
nand NAND3 (N1755, N1751, N272, N742);
not NOT1 (N1756, N1745);
xor XOR2 (N1757, N1744, N810);
nor NOR2 (N1758, N1730, N351);
nand NAND3 (N1759, N1755, N1423, N788);
nor NOR2 (N1760, N1759, N730);
or OR3 (N1761, N1749, N58, N1057);
not NOT1 (N1762, N1756);
nand NAND4 (N1763, N1753, N830, N798, N530);
nor NOR3 (N1764, N1760, N265, N1172);
nor NOR4 (N1765, N1762, N1705, N1565, N1529);
or OR2 (N1766, N1754, N1319);
or OR4 (N1767, N1757, N1279, N928, N410);
not NOT1 (N1768, N1758);
nor NOR4 (N1769, N1750, N482, N89, N445);
and AND3 (N1770, N1763, N1413, N720);
or OR3 (N1771, N1761, N541, N1299);
buf BUF1 (N1772, N1767);
buf BUF1 (N1773, N1768);
not NOT1 (N1774, N1764);
or OR4 (N1775, N1769, N544, N238, N1673);
and AND3 (N1776, N1742, N674, N584);
and AND4 (N1777, N1774, N760, N1572, N237);
buf BUF1 (N1778, N1776);
not NOT1 (N1779, N1772);
and AND2 (N1780, N1770, N1727);
nor NOR2 (N1781, N1773, N320);
nand NAND3 (N1782, N1777, N773, N920);
not NOT1 (N1783, N1778);
and AND4 (N1784, N1783, N122, N1089, N1156);
nand NAND3 (N1785, N1782, N1631, N420);
or OR4 (N1786, N1734, N1347, N769, N554);
xor XOR2 (N1787, N1786, N1377);
not NOT1 (N1788, N1784);
xor XOR2 (N1789, N1766, N1454);
not NOT1 (N1790, N1771);
and AND4 (N1791, N1787, N1089, N495, N512);
buf BUF1 (N1792, N1781);
not NOT1 (N1793, N1765);
nor NOR2 (N1794, N1788, N752);
not NOT1 (N1795, N1779);
or OR2 (N1796, N1792, N1336);
nand NAND3 (N1797, N1791, N937, N599);
xor XOR2 (N1798, N1793, N892);
or OR2 (N1799, N1795, N599);
buf BUF1 (N1800, N1790);
nor NOR2 (N1801, N1797, N594);
nand NAND4 (N1802, N1799, N991, N1772, N620);
nand NAND4 (N1803, N1798, N1088, N1156, N167);
not NOT1 (N1804, N1789);
or OR2 (N1805, N1780, N153);
nor NOR3 (N1806, N1805, N574, N1209);
buf BUF1 (N1807, N1806);
not NOT1 (N1808, N1794);
or OR4 (N1809, N1796, N695, N1620, N356);
and AND2 (N1810, N1808, N1355);
or OR2 (N1811, N1802, N1452);
nand NAND3 (N1812, N1807, N1327, N1349);
not NOT1 (N1813, N1810);
buf BUF1 (N1814, N1804);
nand NAND4 (N1815, N1803, N1149, N745, N11);
not NOT1 (N1816, N1813);
nor NOR3 (N1817, N1775, N1203, N1035);
nor NOR3 (N1818, N1814, N457, N237);
and AND3 (N1819, N1815, N1433, N1002);
xor XOR2 (N1820, N1811, N1282);
xor XOR2 (N1821, N1818, N1432);
buf BUF1 (N1822, N1819);
nor NOR2 (N1823, N1821, N886);
buf BUF1 (N1824, N1820);
xor XOR2 (N1825, N1822, N872);
nand NAND4 (N1826, N1812, N1449, N1497, N964);
or OR4 (N1827, N1785, N723, N575, N1762);
and AND2 (N1828, N1801, N1381);
or OR3 (N1829, N1827, N1253, N1584);
nor NOR4 (N1830, N1826, N39, N910, N830);
buf BUF1 (N1831, N1823);
not NOT1 (N1832, N1831);
buf BUF1 (N1833, N1832);
and AND2 (N1834, N1825, N231);
and AND4 (N1835, N1828, N1461, N367, N1491);
not NOT1 (N1836, N1833);
xor XOR2 (N1837, N1816, N771);
xor XOR2 (N1838, N1817, N751);
and AND3 (N1839, N1837, N316, N500);
buf BUF1 (N1840, N1834);
not NOT1 (N1841, N1840);
buf BUF1 (N1842, N1800);
xor XOR2 (N1843, N1824, N1583);
xor XOR2 (N1844, N1835, N1281);
and AND3 (N1845, N1829, N1445, N664);
or OR2 (N1846, N1842, N1145);
nand NAND2 (N1847, N1841, N1074);
buf BUF1 (N1848, N1830);
not NOT1 (N1849, N1845);
not NOT1 (N1850, N1847);
buf BUF1 (N1851, N1850);
not NOT1 (N1852, N1843);
xor XOR2 (N1853, N1848, N1818);
xor XOR2 (N1854, N1844, N1834);
not NOT1 (N1855, N1838);
or OR2 (N1856, N1836, N1710);
xor XOR2 (N1857, N1809, N954);
buf BUF1 (N1858, N1851);
nand NAND4 (N1859, N1855, N488, N863, N1617);
xor XOR2 (N1860, N1856, N592);
nor NOR2 (N1861, N1839, N1010);
or OR3 (N1862, N1859, N715, N1569);
and AND2 (N1863, N1849, N1520);
not NOT1 (N1864, N1863);
not NOT1 (N1865, N1846);
not NOT1 (N1866, N1860);
nand NAND2 (N1867, N1854, N1265);
xor XOR2 (N1868, N1865, N885);
nor NOR4 (N1869, N1867, N592, N1722, N1488);
nand NAND2 (N1870, N1864, N1522);
and AND2 (N1871, N1868, N1218);
or OR4 (N1872, N1857, N539, N1638, N842);
buf BUF1 (N1873, N1858);
or OR4 (N1874, N1862, N66, N987, N101);
or OR2 (N1875, N1870, N1685);
or OR3 (N1876, N1873, N961, N472);
or OR2 (N1877, N1869, N1749);
nand NAND3 (N1878, N1874, N1610, N1273);
not NOT1 (N1879, N1878);
nand NAND3 (N1880, N1872, N470, N562);
xor XOR2 (N1881, N1861, N47);
not NOT1 (N1882, N1876);
nor NOR2 (N1883, N1879, N1086);
not NOT1 (N1884, N1875);
xor XOR2 (N1885, N1882, N429);
buf BUF1 (N1886, N1852);
buf BUF1 (N1887, N1853);
nor NOR3 (N1888, N1883, N1379, N1611);
xor XOR2 (N1889, N1887, N413);
or OR2 (N1890, N1884, N314);
xor XOR2 (N1891, N1890, N1782);
nor NOR3 (N1892, N1881, N1257, N973);
not NOT1 (N1893, N1886);
nor NOR3 (N1894, N1893, N1636, N1519);
or OR2 (N1895, N1894, N751);
not NOT1 (N1896, N1891);
xor XOR2 (N1897, N1885, N1491);
or OR3 (N1898, N1895, N1000, N1738);
or OR3 (N1899, N1880, N1507, N1538);
nor NOR4 (N1900, N1871, N1838, N647, N272);
or OR2 (N1901, N1899, N1165);
and AND3 (N1902, N1900, N656, N582);
or OR2 (N1903, N1888, N951);
or OR4 (N1904, N1889, N683, N724, N1426);
nor NOR2 (N1905, N1877, N394);
or OR4 (N1906, N1896, N870, N1868, N1738);
or OR4 (N1907, N1892, N353, N119, N1752);
buf BUF1 (N1908, N1898);
and AND4 (N1909, N1905, N386, N173, N1286);
or OR4 (N1910, N1897, N570, N81, N439);
buf BUF1 (N1911, N1866);
and AND3 (N1912, N1902, N1070, N865);
nor NOR2 (N1913, N1904, N255);
xor XOR2 (N1914, N1913, N488);
or OR4 (N1915, N1908, N993, N1573, N1830);
xor XOR2 (N1916, N1911, N1237);
nor NOR2 (N1917, N1914, N123);
nand NAND2 (N1918, N1917, N889);
nor NOR3 (N1919, N1909, N362, N700);
xor XOR2 (N1920, N1915, N1240);
buf BUF1 (N1921, N1919);
and AND2 (N1922, N1916, N274);
nand NAND3 (N1923, N1906, N916, N755);
nand NAND4 (N1924, N1912, N1031, N813, N376);
and AND4 (N1925, N1920, N1779, N1417, N1519);
nand NAND2 (N1926, N1924, N1376);
or OR3 (N1927, N1910, N952, N436);
not NOT1 (N1928, N1922);
buf BUF1 (N1929, N1925);
and AND4 (N1930, N1929, N608, N778, N1591);
nand NAND4 (N1931, N1928, N1532, N1119, N1159);
or OR3 (N1932, N1927, N6, N1172);
xor XOR2 (N1933, N1930, N630);
nand NAND4 (N1934, N1932, N1086, N726, N713);
buf BUF1 (N1935, N1903);
and AND3 (N1936, N1901, N504, N1375);
xor XOR2 (N1937, N1926, N339);
and AND4 (N1938, N1921, N1834, N1068, N1514);
buf BUF1 (N1939, N1933);
buf BUF1 (N1940, N1937);
not NOT1 (N1941, N1918);
buf BUF1 (N1942, N1936);
nand NAND2 (N1943, N1931, N742);
not NOT1 (N1944, N1935);
nand NAND3 (N1945, N1944, N1500, N762);
or OR4 (N1946, N1945, N1549, N557, N460);
nor NOR3 (N1947, N1946, N944, N1500);
not NOT1 (N1948, N1939);
not NOT1 (N1949, N1947);
nor NOR4 (N1950, N1938, N1282, N1191, N550);
not NOT1 (N1951, N1949);
buf BUF1 (N1952, N1942);
xor XOR2 (N1953, N1934, N223);
or OR3 (N1954, N1952, N789, N1588);
not NOT1 (N1955, N1950);
nor NOR3 (N1956, N1954, N582, N528);
not NOT1 (N1957, N1940);
buf BUF1 (N1958, N1907);
buf BUF1 (N1959, N1923);
or OR4 (N1960, N1943, N1708, N1144, N1029);
nor NOR2 (N1961, N1951, N1052);
or OR3 (N1962, N1959, N885, N1419);
not NOT1 (N1963, N1955);
buf BUF1 (N1964, N1957);
nor NOR3 (N1965, N1960, N69, N1140);
buf BUF1 (N1966, N1962);
and AND4 (N1967, N1956, N1158, N1329, N611);
nand NAND4 (N1968, N1965, N1441, N54, N613);
and AND3 (N1969, N1964, N476, N1169);
xor XOR2 (N1970, N1968, N337);
xor XOR2 (N1971, N1966, N1154);
buf BUF1 (N1972, N1970);
buf BUF1 (N1973, N1953);
nand NAND3 (N1974, N1941, N1891, N1630);
or OR2 (N1975, N1972, N1007);
or OR4 (N1976, N1971, N1626, N190, N1416);
nor NOR2 (N1977, N1958, N13);
and AND2 (N1978, N1973, N888);
not NOT1 (N1979, N1969);
nor NOR3 (N1980, N1961, N1111, N1756);
not NOT1 (N1981, N1978);
or OR4 (N1982, N1974, N32, N1478, N1675);
or OR4 (N1983, N1975, N950, N1973, N1717);
not NOT1 (N1984, N1982);
or OR2 (N1985, N1976, N863);
not NOT1 (N1986, N1967);
nand NAND3 (N1987, N1977, N911, N369);
or OR3 (N1988, N1981, N1589, N1048);
nand NAND2 (N1989, N1963, N559);
and AND4 (N1990, N1984, N447, N259, N1925);
xor XOR2 (N1991, N1989, N1276);
nor NOR3 (N1992, N1980, N1508, N721);
buf BUF1 (N1993, N1991);
nand NAND2 (N1994, N1985, N972);
xor XOR2 (N1995, N1993, N43);
not NOT1 (N1996, N1995);
and AND2 (N1997, N1979, N1842);
buf BUF1 (N1998, N1988);
or OR3 (N1999, N1983, N650, N1362);
or OR4 (N2000, N1999, N1246, N1956, N1498);
not NOT1 (N2001, N1998);
or OR2 (N2002, N1994, N1649);
xor XOR2 (N2003, N1990, N1324);
and AND4 (N2004, N1996, N719, N624, N1176);
xor XOR2 (N2005, N2001, N123);
not NOT1 (N2006, N1987);
or OR3 (N2007, N2004, N1343, N1427);
nor NOR2 (N2008, N2000, N1120);
nand NAND3 (N2009, N1997, N1739, N421);
xor XOR2 (N2010, N1948, N179);
nand NAND4 (N2011, N2009, N1078, N1685, N36);
xor XOR2 (N2012, N2008, N1915);
xor XOR2 (N2013, N1992, N1028);
nor NOR3 (N2014, N2003, N637, N270);
buf BUF1 (N2015, N2010);
not NOT1 (N2016, N2014);
buf BUF1 (N2017, N2015);
not NOT1 (N2018, N2006);
or OR3 (N2019, N2012, N660, N1516);
buf BUF1 (N2020, N2007);
and AND2 (N2021, N1986, N188);
nand NAND4 (N2022, N2011, N1621, N1781, N1451);
nor NOR3 (N2023, N2018, N703, N4);
nor NOR2 (N2024, N2016, N1542);
and AND4 (N2025, N2024, N1841, N1036, N1205);
or OR2 (N2026, N2020, N47);
xor XOR2 (N2027, N2021, N466);
not NOT1 (N2028, N2005);
buf BUF1 (N2029, N2026);
nor NOR3 (N2030, N2002, N539, N771);
and AND2 (N2031, N2028, N1662);
nand NAND2 (N2032, N2029, N1791);
or OR4 (N2033, N2019, N872, N46, N573);
or OR3 (N2034, N2017, N1874, N1882);
or OR2 (N2035, N2025, N1303);
and AND3 (N2036, N2030, N665, N1467);
and AND4 (N2037, N2013, N511, N1641, N1367);
and AND2 (N2038, N2033, N962);
xor XOR2 (N2039, N2023, N125);
nand NAND3 (N2040, N2027, N983, N766);
xor XOR2 (N2041, N2034, N294);
nor NOR2 (N2042, N2041, N954);
xor XOR2 (N2043, N2037, N1565);
nor NOR2 (N2044, N2039, N1932);
nand NAND4 (N2045, N2035, N329, N926, N1167);
not NOT1 (N2046, N2045);
not NOT1 (N2047, N2046);
or OR4 (N2048, N2044, N1889, N1145, N384);
or OR2 (N2049, N2043, N429);
or OR3 (N2050, N2031, N590, N439);
not NOT1 (N2051, N2022);
not NOT1 (N2052, N2047);
not NOT1 (N2053, N2052);
or OR4 (N2054, N2036, N1840, N832, N1982);
xor XOR2 (N2055, N2049, N496);
or OR2 (N2056, N2048, N775);
and AND4 (N2057, N2053, N1370, N953, N1);
nor NOR3 (N2058, N2038, N1230, N1722);
nand NAND2 (N2059, N2040, N664);
nor NOR4 (N2060, N2051, N229, N942, N670);
and AND4 (N2061, N2059, N1093, N1989, N1815);
xor XOR2 (N2062, N2061, N2017);
nand NAND2 (N2063, N2062, N1201);
buf BUF1 (N2064, N2032);
nor NOR2 (N2065, N2050, N580);
and AND2 (N2066, N2054, N947);
xor XOR2 (N2067, N2063, N716);
or OR3 (N2068, N2067, N1914, N823);
nand NAND4 (N2069, N2058, N755, N1164, N702);
buf BUF1 (N2070, N2057);
and AND2 (N2071, N2069, N438);
nand NAND2 (N2072, N2071, N1780);
buf BUF1 (N2073, N2065);
nand NAND3 (N2074, N2055, N1866, N316);
xor XOR2 (N2075, N2068, N1163);
and AND2 (N2076, N2066, N1399);
nand NAND3 (N2077, N2074, N1568, N272);
xor XOR2 (N2078, N2042, N1236);
not NOT1 (N2079, N2064);
nor NOR2 (N2080, N2056, N521);
or OR3 (N2081, N2077, N1740, N1247);
buf BUF1 (N2082, N2073);
nor NOR4 (N2083, N2070, N319, N1966, N1614);
or OR2 (N2084, N2081, N550);
buf BUF1 (N2085, N2075);
or OR3 (N2086, N2060, N384, N1964);
not NOT1 (N2087, N2085);
xor XOR2 (N2088, N2082, N1802);
nor NOR2 (N2089, N2078, N13);
buf BUF1 (N2090, N2088);
or OR2 (N2091, N2086, N2058);
nor NOR4 (N2092, N2072, N1470, N511, N821);
and AND3 (N2093, N2090, N1646, N199);
xor XOR2 (N2094, N2084, N1281);
buf BUF1 (N2095, N2091);
or OR3 (N2096, N2076, N1718, N1936);
nand NAND3 (N2097, N2079, N757, N85);
not NOT1 (N2098, N2092);
nand NAND2 (N2099, N2089, N946);
xor XOR2 (N2100, N2097, N30);
nand NAND4 (N2101, N2099, N369, N350, N1879);
xor XOR2 (N2102, N2087, N1966);
or OR2 (N2103, N2095, N161);
buf BUF1 (N2104, N2101);
xor XOR2 (N2105, N2103, N924);
nand NAND3 (N2106, N2083, N181, N1724);
xor XOR2 (N2107, N2100, N1737);
and AND4 (N2108, N2107, N1025, N18, N861);
buf BUF1 (N2109, N2105);
and AND3 (N2110, N2104, N257, N251);
xor XOR2 (N2111, N2093, N671);
nand NAND4 (N2112, N2098, N202, N453, N1079);
nand NAND4 (N2113, N2110, N1816, N1306, N2068);
nand NAND4 (N2114, N2111, N1284, N1898, N1848);
nand NAND4 (N2115, N2080, N1321, N269, N1592);
nor NOR3 (N2116, N2114, N1712, N431);
buf BUF1 (N2117, N2106);
nand NAND2 (N2118, N2116, N1952);
nor NOR3 (N2119, N2115, N8, N987);
not NOT1 (N2120, N2119);
and AND4 (N2121, N2102, N1105, N1645, N843);
xor XOR2 (N2122, N2096, N55);
or OR3 (N2123, N2121, N1475, N1779);
and AND2 (N2124, N2117, N393);
and AND4 (N2125, N2094, N1504, N146, N2064);
not NOT1 (N2126, N2113);
xor XOR2 (N2127, N2123, N356);
buf BUF1 (N2128, N2124);
xor XOR2 (N2129, N2112, N2046);
nor NOR3 (N2130, N2128, N686, N934);
or OR3 (N2131, N2118, N1161, N1640);
xor XOR2 (N2132, N2120, N928);
and AND2 (N2133, N2132, N1443);
not NOT1 (N2134, N2130);
and AND4 (N2135, N2126, N1987, N2099, N1430);
xor XOR2 (N2136, N2133, N845);
nand NAND3 (N2137, N2109, N648, N874);
xor XOR2 (N2138, N2125, N205);
xor XOR2 (N2139, N2129, N203);
nor NOR2 (N2140, N2139, N1482);
xor XOR2 (N2141, N2138, N644);
buf BUF1 (N2142, N2137);
nand NAND4 (N2143, N2127, N311, N1011, N15);
buf BUF1 (N2144, N2122);
not NOT1 (N2145, N2134);
buf BUF1 (N2146, N2140);
buf BUF1 (N2147, N2135);
and AND3 (N2148, N2147, N589, N122);
and AND3 (N2149, N2144, N1698, N1103);
not NOT1 (N2150, N2136);
and AND2 (N2151, N2143, N1347);
nor NOR2 (N2152, N2142, N122);
xor XOR2 (N2153, N2131, N381);
or OR2 (N2154, N2153, N1340);
buf BUF1 (N2155, N2148);
nor NOR4 (N2156, N2146, N88, N1286, N1668);
nand NAND4 (N2157, N2108, N745, N169, N2072);
and AND3 (N2158, N2154, N2120, N1017);
nand NAND3 (N2159, N2151, N1061, N985);
xor XOR2 (N2160, N2145, N1960);
and AND3 (N2161, N2155, N990, N1378);
xor XOR2 (N2162, N2149, N1596);
xor XOR2 (N2163, N2159, N65);
nor NOR2 (N2164, N2162, N2093);
nand NAND2 (N2165, N2141, N833);
and AND3 (N2166, N2164, N1408, N1861);
nor NOR4 (N2167, N2157, N756, N1465, N666);
xor XOR2 (N2168, N2165, N2124);
xor XOR2 (N2169, N2168, N2105);
or OR2 (N2170, N2161, N490);
nand NAND4 (N2171, N2150, N899, N2167, N28);
xor XOR2 (N2172, N1680, N494);
or OR3 (N2173, N2169, N1194, N950);
buf BUF1 (N2174, N2172);
buf BUF1 (N2175, N2156);
nand NAND3 (N2176, N2171, N778, N282);
nand NAND2 (N2177, N2160, N373);
nor NOR3 (N2178, N2173, N1793, N2174);
and AND4 (N2179, N1069, N688, N1668, N83);
not NOT1 (N2180, N2178);
xor XOR2 (N2181, N2177, N2118);
xor XOR2 (N2182, N2158, N1342);
or OR3 (N2183, N2166, N2068, N1683);
xor XOR2 (N2184, N2175, N975);
and AND4 (N2185, N2152, N370, N1625, N503);
nand NAND2 (N2186, N2184, N1912);
nor NOR3 (N2187, N2170, N8, N31);
not NOT1 (N2188, N2176);
or OR3 (N2189, N2187, N1893, N103);
nor NOR3 (N2190, N2180, N50, N2145);
nor NOR3 (N2191, N2163, N1008, N122);
and AND2 (N2192, N2181, N1815);
buf BUF1 (N2193, N2190);
xor XOR2 (N2194, N2189, N722);
nand NAND3 (N2195, N2183, N898, N324);
nor NOR2 (N2196, N2191, N1418);
not NOT1 (N2197, N2194);
nor NOR4 (N2198, N2196, N717, N26, N148);
or OR3 (N2199, N2197, N1164, N712);
xor XOR2 (N2200, N2199, N340);
nand NAND2 (N2201, N2179, N2016);
and AND4 (N2202, N2188, N1761, N1051, N27);
not NOT1 (N2203, N2192);
or OR3 (N2204, N2202, N1333, N679);
nand NAND3 (N2205, N2201, N409, N1930);
or OR2 (N2206, N2205, N1142);
nor NOR3 (N2207, N2185, N346, N2109);
or OR3 (N2208, N2206, N544, N960);
xor XOR2 (N2209, N2200, N1746);
and AND4 (N2210, N2209, N782, N599, N1733);
nor NOR4 (N2211, N2204, N437, N2092, N1032);
or OR4 (N2212, N2208, N125, N1763, N1190);
nor NOR2 (N2213, N2203, N2060);
not NOT1 (N2214, N2195);
xor XOR2 (N2215, N2212, N8);
xor XOR2 (N2216, N2210, N1982);
or OR3 (N2217, N2214, N797, N743);
buf BUF1 (N2218, N2207);
not NOT1 (N2219, N2198);
xor XOR2 (N2220, N2218, N1714);
nand NAND3 (N2221, N2219, N2153, N1570);
xor XOR2 (N2222, N2220, N2196);
and AND4 (N2223, N2186, N1621, N208, N441);
xor XOR2 (N2224, N2213, N2219);
buf BUF1 (N2225, N2211);
or OR2 (N2226, N2223, N1483);
and AND3 (N2227, N2193, N802, N721);
and AND2 (N2228, N2222, N611);
or OR3 (N2229, N2225, N99, N707);
not NOT1 (N2230, N2229);
xor XOR2 (N2231, N2216, N820);
or OR4 (N2232, N2231, N668, N1459, N101);
or OR4 (N2233, N2224, N1132, N144, N776);
or OR4 (N2234, N2215, N326, N442, N1580);
not NOT1 (N2235, N2232);
xor XOR2 (N2236, N2228, N1303);
and AND2 (N2237, N2217, N1348);
not NOT1 (N2238, N2235);
buf BUF1 (N2239, N2238);
nor NOR2 (N2240, N2182, N567);
and AND2 (N2241, N2236, N1437);
xor XOR2 (N2242, N2226, N463);
buf BUF1 (N2243, N2227);
not NOT1 (N2244, N2242);
buf BUF1 (N2245, N2240);
buf BUF1 (N2246, N2233);
nor NOR4 (N2247, N2246, N954, N850, N1649);
not NOT1 (N2248, N2234);
buf BUF1 (N2249, N2221);
and AND2 (N2250, N2244, N311);
xor XOR2 (N2251, N2245, N661);
nor NOR2 (N2252, N2243, N667);
xor XOR2 (N2253, N2251, N520);
nor NOR4 (N2254, N2239, N2225, N854, N701);
nand NAND3 (N2255, N2249, N2208, N1275);
buf BUF1 (N2256, N2254);
xor XOR2 (N2257, N2252, N857);
nand NAND3 (N2258, N2248, N167, N925);
xor XOR2 (N2259, N2257, N113);
buf BUF1 (N2260, N2247);
buf BUF1 (N2261, N2230);
xor XOR2 (N2262, N2260, N1981);
nand NAND2 (N2263, N2262, N394);
nor NOR3 (N2264, N2258, N1341, N229);
not NOT1 (N2265, N2237);
xor XOR2 (N2266, N2259, N1174);
not NOT1 (N2267, N2253);
nor NOR3 (N2268, N2267, N1831, N49);
and AND3 (N2269, N2241, N1158, N2025);
nor NOR3 (N2270, N2266, N751, N1207);
nand NAND3 (N2271, N2261, N1702, N1250);
xor XOR2 (N2272, N2255, N1807);
nand NAND3 (N2273, N2272, N2133, N595);
nand NAND4 (N2274, N2268, N1621, N480, N380);
buf BUF1 (N2275, N2269);
and AND4 (N2276, N2271, N632, N1074, N1181);
xor XOR2 (N2277, N2264, N1167);
nor NOR3 (N2278, N2273, N1509, N767);
not NOT1 (N2279, N2265);
not NOT1 (N2280, N2256);
nand NAND2 (N2281, N2263, N104);
buf BUF1 (N2282, N2279);
nand NAND2 (N2283, N2281, N2097);
not NOT1 (N2284, N2274);
nand NAND2 (N2285, N2284, N692);
or OR4 (N2286, N2250, N151, N1419, N1875);
and AND2 (N2287, N2270, N308);
xor XOR2 (N2288, N2282, N372);
nor NOR2 (N2289, N2287, N1544);
or OR4 (N2290, N2278, N1201, N323, N1084);
nor NOR4 (N2291, N2277, N231, N1565, N188);
nand NAND4 (N2292, N2290, N138, N164, N150);
not NOT1 (N2293, N2276);
not NOT1 (N2294, N2283);
nand NAND3 (N2295, N2285, N2007, N432);
buf BUF1 (N2296, N2291);
xor XOR2 (N2297, N2296, N2049);
or OR3 (N2298, N2292, N1585, N2118);
xor XOR2 (N2299, N2289, N2090);
and AND4 (N2300, N2295, N1368, N2042, N1992);
nand NAND3 (N2301, N2288, N1536, N2197);
xor XOR2 (N2302, N2299, N1873);
or OR3 (N2303, N2280, N1812, N586);
xor XOR2 (N2304, N2302, N1410);
nand NAND4 (N2305, N2297, N545, N1764, N2071);
and AND4 (N2306, N2286, N2227, N1639, N272);
not NOT1 (N2307, N2298);
and AND4 (N2308, N2300, N474, N1671, N2194);
or OR3 (N2309, N2308, N1621, N108);
nor NOR4 (N2310, N2294, N2308, N317, N1878);
xor XOR2 (N2311, N2309, N1920);
nor NOR2 (N2312, N2303, N767);
xor XOR2 (N2313, N2307, N773);
not NOT1 (N2314, N2306);
nor NOR2 (N2315, N2312, N773);
nor NOR2 (N2316, N2275, N811);
buf BUF1 (N2317, N2315);
nor NOR4 (N2318, N2317, N2046, N922, N779);
nor NOR2 (N2319, N2318, N790);
or OR2 (N2320, N2310, N1590);
buf BUF1 (N2321, N2319);
buf BUF1 (N2322, N2314);
or OR3 (N2323, N2304, N1887, N2047);
and AND2 (N2324, N2323, N1465);
xor XOR2 (N2325, N2301, N1851);
buf BUF1 (N2326, N2322);
nand NAND4 (N2327, N2293, N304, N517, N1314);
or OR3 (N2328, N2326, N636, N2265);
nor NOR2 (N2329, N2321, N856);
nand NAND4 (N2330, N2329, N2207, N1151, N409);
not NOT1 (N2331, N2325);
buf BUF1 (N2332, N2324);
and AND4 (N2333, N2332, N454, N408, N603);
nor NOR2 (N2334, N2328, N1370);
or OR3 (N2335, N2333, N1609, N896);
and AND4 (N2336, N2311, N530, N1370, N121);
nor NOR3 (N2337, N2316, N1262, N1933);
and AND4 (N2338, N2334, N2028, N1868, N1511);
or OR3 (N2339, N2330, N191, N709);
and AND2 (N2340, N2327, N712);
and AND4 (N2341, N2340, N1491, N553, N921);
or OR3 (N2342, N2335, N2162, N1157);
xor XOR2 (N2343, N2305, N198);
nor NOR4 (N2344, N2331, N1454, N292, N2090);
or OR3 (N2345, N2339, N1207, N626);
xor XOR2 (N2346, N2337, N1240);
and AND4 (N2347, N2344, N692, N191, N1959);
buf BUF1 (N2348, N2336);
not NOT1 (N2349, N2341);
xor XOR2 (N2350, N2343, N735);
not NOT1 (N2351, N2348);
buf BUF1 (N2352, N2347);
not NOT1 (N2353, N2350);
xor XOR2 (N2354, N2313, N1324);
not NOT1 (N2355, N2351);
and AND2 (N2356, N2352, N187);
nor NOR3 (N2357, N2345, N1364, N653);
buf BUF1 (N2358, N2342);
buf BUF1 (N2359, N2349);
nor NOR2 (N2360, N2355, N2293);
and AND4 (N2361, N2357, N284, N1206, N1123);
or OR4 (N2362, N2360, N1667, N1256, N327);
and AND4 (N2363, N2359, N24, N311, N1657);
or OR3 (N2364, N2338, N71, N1729);
xor XOR2 (N2365, N2361, N122);
buf BUF1 (N2366, N2365);
nor NOR3 (N2367, N2358, N1221, N438);
not NOT1 (N2368, N2364);
not NOT1 (N2369, N2367);
nand NAND2 (N2370, N2353, N2257);
not NOT1 (N2371, N2346);
xor XOR2 (N2372, N2368, N1695);
buf BUF1 (N2373, N2354);
not NOT1 (N2374, N2363);
nor NOR2 (N2375, N2366, N1936);
and AND4 (N2376, N2362, N642, N2348, N2335);
buf BUF1 (N2377, N2356);
buf BUF1 (N2378, N2376);
not NOT1 (N2379, N2378);
and AND4 (N2380, N2372, N164, N310, N1503);
buf BUF1 (N2381, N2380);
xor XOR2 (N2382, N2374, N2138);
not NOT1 (N2383, N2369);
or OR3 (N2384, N2375, N33, N974);
buf BUF1 (N2385, N2379);
xor XOR2 (N2386, N2381, N2062);
nand NAND3 (N2387, N2377, N1291, N2144);
nor NOR4 (N2388, N2384, N781, N1414, N574);
not NOT1 (N2389, N2383);
not NOT1 (N2390, N2386);
not NOT1 (N2391, N2382);
buf BUF1 (N2392, N2388);
or OR4 (N2393, N2371, N743, N2029, N425);
nand NAND2 (N2394, N2390, N1728);
or OR4 (N2395, N2373, N547, N278, N459);
and AND4 (N2396, N2394, N757, N219, N1461);
or OR3 (N2397, N2389, N375, N635);
buf BUF1 (N2398, N2387);
or OR2 (N2399, N2393, N1439);
or OR2 (N2400, N2320, N2358);
nand NAND4 (N2401, N2392, N1809, N2159, N1589);
not NOT1 (N2402, N2398);
nor NOR4 (N2403, N2385, N1186, N452, N1211);
nand NAND4 (N2404, N2370, N1443, N2239, N2096);
nand NAND2 (N2405, N2400, N1294);
buf BUF1 (N2406, N2397);
and AND4 (N2407, N2401, N1889, N2040, N2353);
or OR3 (N2408, N2391, N2097, N680);
nand NAND4 (N2409, N2395, N1917, N1272, N2253);
nor NOR2 (N2410, N2405, N1329);
buf BUF1 (N2411, N2403);
buf BUF1 (N2412, N2407);
nand NAND2 (N2413, N2399, N1744);
nor NOR3 (N2414, N2408, N807, N1395);
xor XOR2 (N2415, N2404, N185);
not NOT1 (N2416, N2410);
nor NOR4 (N2417, N2413, N2409, N1909, N1167);
nand NAND2 (N2418, N707, N568);
xor XOR2 (N2419, N2411, N10);
xor XOR2 (N2420, N2402, N84);
nor NOR4 (N2421, N2412, N374, N2164, N2047);
nor NOR4 (N2422, N2418, N209, N1658, N719);
buf BUF1 (N2423, N2416);
nand NAND4 (N2424, N2414, N561, N453, N1049);
xor XOR2 (N2425, N2423, N1783);
nand NAND3 (N2426, N2396, N76, N1618);
nand NAND4 (N2427, N2425, N357, N2154, N1496);
or OR2 (N2428, N2424, N1694);
not NOT1 (N2429, N2421);
or OR2 (N2430, N2415, N500);
not NOT1 (N2431, N2429);
xor XOR2 (N2432, N2422, N1573);
and AND4 (N2433, N2430, N159, N106, N1914);
buf BUF1 (N2434, N2426);
nor NOR4 (N2435, N2428, N951, N1054, N2392);
buf BUF1 (N2436, N2417);
and AND2 (N2437, N2432, N1882);
and AND3 (N2438, N2419, N2359, N437);
not NOT1 (N2439, N2420);
nor NOR2 (N2440, N2431, N2369);
not NOT1 (N2441, N2438);
xor XOR2 (N2442, N2435, N62);
nand NAND2 (N2443, N2440, N1855);
xor XOR2 (N2444, N2427, N27);
buf BUF1 (N2445, N2434);
nand NAND3 (N2446, N2433, N1617, N179);
not NOT1 (N2447, N2443);
not NOT1 (N2448, N2436);
not NOT1 (N2449, N2442);
nand NAND3 (N2450, N2444, N2198, N1232);
and AND2 (N2451, N2406, N1408);
buf BUF1 (N2452, N2445);
and AND4 (N2453, N2450, N1617, N356, N2443);
not NOT1 (N2454, N2449);
and AND4 (N2455, N2447, N353, N1735, N2358);
buf BUF1 (N2456, N2446);
nand NAND4 (N2457, N2453, N352, N1828, N1240);
nand NAND4 (N2458, N2457, N1152, N493, N205);
nand NAND4 (N2459, N2455, N1515, N1685, N1167);
or OR4 (N2460, N2459, N1702, N2380, N217);
buf BUF1 (N2461, N2441);
nand NAND3 (N2462, N2451, N1410, N673);
nand NAND3 (N2463, N2439, N1436, N1915);
nor NOR4 (N2464, N2454, N1137, N1150, N330);
buf BUF1 (N2465, N2460);
buf BUF1 (N2466, N2452);
not NOT1 (N2467, N2465);
xor XOR2 (N2468, N2448, N1829);
or OR2 (N2469, N2437, N590);
nor NOR3 (N2470, N2463, N568, N1128);
not NOT1 (N2471, N2470);
buf BUF1 (N2472, N2466);
or OR2 (N2473, N2461, N675);
buf BUF1 (N2474, N2469);
nor NOR2 (N2475, N2464, N134);
buf BUF1 (N2476, N2468);
nand NAND3 (N2477, N2458, N11, N389);
nand NAND2 (N2478, N2471, N451);
nand NAND3 (N2479, N2472, N319, N2250);
nor NOR2 (N2480, N2477, N2015);
not NOT1 (N2481, N2478);
nor NOR3 (N2482, N2475, N212, N1933);
nand NAND2 (N2483, N2482, N923);
xor XOR2 (N2484, N2473, N892);
xor XOR2 (N2485, N2456, N783);
or OR2 (N2486, N2481, N1861);
xor XOR2 (N2487, N2467, N2486);
nor NOR2 (N2488, N2354, N375);
not NOT1 (N2489, N2484);
or OR3 (N2490, N2485, N1653, N1339);
not NOT1 (N2491, N2476);
nand NAND4 (N2492, N2479, N2196, N697, N2227);
and AND2 (N2493, N2474, N1227);
xor XOR2 (N2494, N2483, N904);
buf BUF1 (N2495, N2480);
buf BUF1 (N2496, N2487);
or OR3 (N2497, N2492, N2281, N832);
buf BUF1 (N2498, N2490);
or OR4 (N2499, N2497, N1030, N1174, N1528);
buf BUF1 (N2500, N2462);
or OR2 (N2501, N2488, N1233);
buf BUF1 (N2502, N2491);
nand NAND4 (N2503, N2502, N1946, N1870, N2253);
nor NOR4 (N2504, N2503, N16, N1796, N94);
not NOT1 (N2505, N2495);
nand NAND2 (N2506, N2500, N2081);
not NOT1 (N2507, N2493);
xor XOR2 (N2508, N2489, N210);
xor XOR2 (N2509, N2494, N213);
buf BUF1 (N2510, N2499);
nor NOR4 (N2511, N2506, N207, N570, N2341);
nand NAND3 (N2512, N2507, N439, N2310);
nor NOR2 (N2513, N2496, N683);
xor XOR2 (N2514, N2505, N718);
xor XOR2 (N2515, N2513, N2458);
nor NOR4 (N2516, N2501, N1971, N2049, N1157);
nand NAND4 (N2517, N2509, N1109, N764, N549);
not NOT1 (N2518, N2517);
and AND4 (N2519, N2508, N1066, N2504, N1346);
nand NAND4 (N2520, N782, N1659, N1210, N528);
and AND4 (N2521, N2510, N2287, N1916, N611);
nand NAND4 (N2522, N2514, N368, N1087, N2340);
nand NAND4 (N2523, N2522, N862, N2260, N2514);
buf BUF1 (N2524, N2516);
nor NOR3 (N2525, N2521, N761, N441);
nand NAND2 (N2526, N2515, N1980);
and AND4 (N2527, N2518, N1035, N1061, N1392);
nand NAND4 (N2528, N2523, N2333, N1015, N568);
xor XOR2 (N2529, N2511, N1299);
xor XOR2 (N2530, N2526, N131);
xor XOR2 (N2531, N2520, N878);
nor NOR4 (N2532, N2530, N990, N1564, N2270);
nand NAND3 (N2533, N2524, N1720, N2134);
and AND4 (N2534, N2531, N1017, N2457, N278);
or OR3 (N2535, N2533, N861, N2046);
nor NOR2 (N2536, N2528, N1987);
buf BUF1 (N2537, N2525);
nor NOR4 (N2538, N2519, N1171, N1460, N2223);
or OR3 (N2539, N2512, N1869, N2164);
not NOT1 (N2540, N2539);
and AND3 (N2541, N2532, N1094, N1842);
nor NOR4 (N2542, N2536, N1521, N1807, N2210);
not NOT1 (N2543, N2527);
nor NOR4 (N2544, N2541, N1714, N420, N4);
nand NAND4 (N2545, N2537, N750, N1380, N1918);
nor NOR3 (N2546, N2540, N1432, N1862);
not NOT1 (N2547, N2545);
nor NOR2 (N2548, N2544, N1193);
nand NAND3 (N2549, N2548, N2449, N1428);
buf BUF1 (N2550, N2534);
or OR4 (N2551, N2543, N1812, N1210, N1929);
xor XOR2 (N2552, N2542, N401);
or OR4 (N2553, N2538, N2125, N2375, N1533);
not NOT1 (N2554, N2547);
xor XOR2 (N2555, N2498, N2467);
buf BUF1 (N2556, N2551);
xor XOR2 (N2557, N2550, N752);
not NOT1 (N2558, N2556);
buf BUF1 (N2559, N2546);
not NOT1 (N2560, N2553);
nor NOR2 (N2561, N2552, N940);
buf BUF1 (N2562, N2558);
buf BUF1 (N2563, N2557);
nor NOR4 (N2564, N2562, N1925, N749, N2395);
and AND2 (N2565, N2560, N1930);
not NOT1 (N2566, N2549);
or OR4 (N2567, N2554, N23, N932, N2396);
not NOT1 (N2568, N2567);
nor NOR3 (N2569, N2564, N1272, N266);
buf BUF1 (N2570, N2568);
and AND2 (N2571, N2529, N1023);
nor NOR2 (N2572, N2569, N1971);
and AND3 (N2573, N2535, N402, N2459);
or OR4 (N2574, N2572, N1105, N1318, N2002);
buf BUF1 (N2575, N2570);
or OR4 (N2576, N2555, N2331, N1634, N1623);
xor XOR2 (N2577, N2561, N484);
and AND3 (N2578, N2573, N1611, N194);
nor NOR2 (N2579, N2575, N106);
not NOT1 (N2580, N2576);
buf BUF1 (N2581, N2577);
and AND2 (N2582, N2566, N656);
and AND2 (N2583, N2559, N1205);
not NOT1 (N2584, N2582);
or OR4 (N2585, N2584, N2513, N18, N652);
and AND4 (N2586, N2579, N108, N707, N210);
and AND3 (N2587, N2586, N1145, N2503);
not NOT1 (N2588, N2581);
nor NOR4 (N2589, N2580, N1467, N124, N1781);
or OR2 (N2590, N2578, N575);
not NOT1 (N2591, N2563);
not NOT1 (N2592, N2565);
buf BUF1 (N2593, N2574);
nand NAND3 (N2594, N2592, N20, N2255);
buf BUF1 (N2595, N2594);
buf BUF1 (N2596, N2589);
or OR2 (N2597, N2571, N1037);
not NOT1 (N2598, N2588);
nor NOR2 (N2599, N2593, N2531);
or OR4 (N2600, N2590, N1447, N1421, N866);
nand NAND3 (N2601, N2600, N285, N719);
or OR3 (N2602, N2583, N29, N919);
and AND4 (N2603, N2585, N2104, N267, N595);
nor NOR4 (N2604, N2597, N1902, N333, N2401);
not NOT1 (N2605, N2603);
nor NOR2 (N2606, N2604, N2485);
nor NOR2 (N2607, N2606, N2353);
not NOT1 (N2608, N2591);
buf BUF1 (N2609, N2587);
xor XOR2 (N2610, N2599, N2488);
xor XOR2 (N2611, N2609, N1066);
xor XOR2 (N2612, N2601, N164);
buf BUF1 (N2613, N2605);
buf BUF1 (N2614, N2613);
nor NOR3 (N2615, N2614, N1273, N1608);
xor XOR2 (N2616, N2611, N155);
or OR3 (N2617, N2615, N1619, N517);
and AND4 (N2618, N2607, N1501, N136, N1211);
not NOT1 (N2619, N2596);
not NOT1 (N2620, N2617);
and AND4 (N2621, N2618, N2464, N1432, N1460);
nor NOR3 (N2622, N2620, N2054, N2070);
xor XOR2 (N2623, N2608, N2325);
and AND3 (N2624, N2612, N184, N1903);
nand NAND2 (N2625, N2621, N2488);
nand NAND4 (N2626, N2616, N986, N2509, N1064);
nor NOR2 (N2627, N2625, N305);
or OR3 (N2628, N2626, N1278, N1281);
not NOT1 (N2629, N2628);
and AND2 (N2630, N2602, N95);
and AND3 (N2631, N2624, N1807, N272);
and AND4 (N2632, N2619, N617, N2290, N143);
nand NAND3 (N2633, N2598, N2086, N294);
nand NAND2 (N2634, N2595, N996);
or OR3 (N2635, N2610, N1254, N930);
xor XOR2 (N2636, N2622, N1037);
not NOT1 (N2637, N2631);
buf BUF1 (N2638, N2623);
nor NOR3 (N2639, N2630, N1999, N976);
xor XOR2 (N2640, N2638, N632);
buf BUF1 (N2641, N2627);
not NOT1 (N2642, N2634);
and AND3 (N2643, N2632, N915, N2161);
buf BUF1 (N2644, N2641);
xor XOR2 (N2645, N2642, N1949);
nand NAND3 (N2646, N2635, N2161, N1602);
and AND4 (N2647, N2629, N512, N1972, N199);
nand NAND2 (N2648, N2646, N1223);
and AND4 (N2649, N2647, N2455, N1558, N188);
and AND3 (N2650, N2643, N2434, N138);
and AND4 (N2651, N2633, N1452, N2233, N1159);
nand NAND2 (N2652, N2651, N20);
or OR4 (N2653, N2652, N876, N1006, N409);
nor NOR4 (N2654, N2648, N237, N1073, N1083);
and AND3 (N2655, N2654, N1728, N380);
nand NAND3 (N2656, N2649, N1500, N361);
buf BUF1 (N2657, N2645);
nand NAND4 (N2658, N2655, N1057, N2081, N2087);
or OR4 (N2659, N2636, N2070, N1304, N629);
not NOT1 (N2660, N2637);
and AND3 (N2661, N2650, N807, N1811);
and AND3 (N2662, N2658, N1099, N155);
buf BUF1 (N2663, N2639);
and AND4 (N2664, N2644, N716, N770, N2589);
not NOT1 (N2665, N2657);
not NOT1 (N2666, N2653);
and AND2 (N2667, N2656, N791);
nand NAND4 (N2668, N2664, N1522, N575, N1129);
buf BUF1 (N2669, N2666);
and AND3 (N2670, N2667, N2576, N1092);
xor XOR2 (N2671, N2661, N54);
and AND4 (N2672, N2670, N931, N1584, N48);
buf BUF1 (N2673, N2663);
nand NAND3 (N2674, N2660, N1470, N535);
nand NAND3 (N2675, N2668, N2569, N1795);
not NOT1 (N2676, N2659);
not NOT1 (N2677, N2674);
nand NAND2 (N2678, N2669, N1026);
buf BUF1 (N2679, N2676);
and AND4 (N2680, N2675, N1353, N1116, N2098);
nand NAND4 (N2681, N2680, N1791, N768, N307);
xor XOR2 (N2682, N2679, N1348);
nand NAND2 (N2683, N2682, N1358);
nor NOR2 (N2684, N2678, N639);
nand NAND2 (N2685, N2640, N1248);
xor XOR2 (N2686, N2672, N1278);
buf BUF1 (N2687, N2683);
nor NOR4 (N2688, N2677, N2649, N2287, N1652);
xor XOR2 (N2689, N2665, N1511);
buf BUF1 (N2690, N2662);
nand NAND4 (N2691, N2671, N464, N1976, N479);
and AND3 (N2692, N2687, N2050, N886);
nor NOR2 (N2693, N2692, N1030);
nor NOR3 (N2694, N2686, N2482, N1358);
or OR2 (N2695, N2689, N1782);
nand NAND3 (N2696, N2688, N759, N2322);
nand NAND4 (N2697, N2695, N1584, N1114, N2631);
nand NAND3 (N2698, N2685, N1996, N2158);
and AND4 (N2699, N2690, N1399, N2454, N395);
nor NOR3 (N2700, N2696, N1589, N1147);
not NOT1 (N2701, N2698);
nor NOR3 (N2702, N2701, N344, N2466);
not NOT1 (N2703, N2681);
and AND3 (N2704, N2684, N107, N1527);
or OR3 (N2705, N2703, N2501, N2381);
or OR4 (N2706, N2691, N669, N871, N1773);
and AND4 (N2707, N2694, N568, N1373, N1620);
nand NAND2 (N2708, N2673, N977);
nor NOR2 (N2709, N2704, N768);
or OR2 (N2710, N2708, N509);
nand NAND3 (N2711, N2707, N398, N2690);
buf BUF1 (N2712, N2709);
nand NAND3 (N2713, N2706, N1172, N264);
nand NAND3 (N2714, N2711, N1563, N183);
and AND3 (N2715, N2700, N2057, N2167);
xor XOR2 (N2716, N2715, N1021);
or OR2 (N2717, N2702, N2340);
or OR3 (N2718, N2714, N1636, N725);
xor XOR2 (N2719, N2710, N814);
or OR2 (N2720, N2718, N1678);
buf BUF1 (N2721, N2716);
xor XOR2 (N2722, N2719, N1159);
or OR4 (N2723, N2705, N87, N1345, N208);
not NOT1 (N2724, N2693);
not NOT1 (N2725, N2721);
nand NAND3 (N2726, N2712, N1717, N713);
not NOT1 (N2727, N2723);
nand NAND3 (N2728, N2699, N2431, N797);
or OR4 (N2729, N2726, N2075, N2615, N1261);
and AND2 (N2730, N2728, N1123);
or OR4 (N2731, N2697, N1850, N285, N2043);
or OR2 (N2732, N2731, N2323);
xor XOR2 (N2733, N2717, N988);
buf BUF1 (N2734, N2724);
nand NAND4 (N2735, N2729, N1964, N1833, N2385);
or OR2 (N2736, N2722, N1704);
and AND4 (N2737, N2713, N2468, N1141, N858);
buf BUF1 (N2738, N2732);
xor XOR2 (N2739, N2725, N2492);
or OR3 (N2740, N2738, N1050, N2047);
not NOT1 (N2741, N2739);
buf BUF1 (N2742, N2733);
or OR3 (N2743, N2737, N2566, N1636);
buf BUF1 (N2744, N2742);
or OR3 (N2745, N2730, N1159, N861);
and AND2 (N2746, N2744, N2387);
and AND2 (N2747, N2734, N2264);
not NOT1 (N2748, N2746);
xor XOR2 (N2749, N2741, N1178);
or OR3 (N2750, N2735, N2359, N1417);
not NOT1 (N2751, N2720);
buf BUF1 (N2752, N2727);
and AND3 (N2753, N2747, N1194, N510);
not NOT1 (N2754, N2748);
or OR2 (N2755, N2740, N103);
buf BUF1 (N2756, N2750);
or OR3 (N2757, N2752, N2550, N115);
nand NAND4 (N2758, N2743, N1203, N1288, N1721);
nor NOR3 (N2759, N2757, N2663, N972);
buf BUF1 (N2760, N2759);
nand NAND4 (N2761, N2749, N1591, N1760, N1140);
xor XOR2 (N2762, N2755, N2677);
and AND3 (N2763, N2754, N2270, N896);
nand NAND2 (N2764, N2736, N2594);
xor XOR2 (N2765, N2764, N301);
or OR2 (N2766, N2745, N528);
or OR3 (N2767, N2761, N568, N1030);
nor NOR4 (N2768, N2765, N2431, N2028, N695);
xor XOR2 (N2769, N2753, N1734);
not NOT1 (N2770, N2760);
buf BUF1 (N2771, N2766);
or OR4 (N2772, N2756, N210, N1136, N2092);
and AND4 (N2773, N2769, N1898, N519, N1565);
and AND2 (N2774, N2768, N1488);
or OR4 (N2775, N2772, N1232, N197, N1579);
nand NAND4 (N2776, N2762, N465, N1246, N1444);
nand NAND4 (N2777, N2776, N812, N2666, N1580);
nor NOR4 (N2778, N2773, N1167, N420, N211);
or OR4 (N2779, N2775, N2336, N916, N699);
xor XOR2 (N2780, N2778, N144);
or OR4 (N2781, N2767, N2459, N1220, N996);
or OR4 (N2782, N2774, N1438, N102, N532);
buf BUF1 (N2783, N2770);
buf BUF1 (N2784, N2780);
and AND2 (N2785, N2758, N911);
nand NAND2 (N2786, N2771, N1580);
buf BUF1 (N2787, N2777);
not NOT1 (N2788, N2763);
nand NAND4 (N2789, N2783, N2434, N2422, N2086);
buf BUF1 (N2790, N2786);
xor XOR2 (N2791, N2790, N2255);
nand NAND3 (N2792, N2785, N1516, N733);
buf BUF1 (N2793, N2788);
or OR4 (N2794, N2792, N1727, N1252, N2181);
not NOT1 (N2795, N2782);
not NOT1 (N2796, N2787);
not NOT1 (N2797, N2793);
xor XOR2 (N2798, N2797, N344);
buf BUF1 (N2799, N2779);
nand NAND2 (N2800, N2789, N1652);
nor NOR2 (N2801, N2798, N579);
nor NOR2 (N2802, N2751, N301);
not NOT1 (N2803, N2801);
not NOT1 (N2804, N2799);
not NOT1 (N2805, N2804);
not NOT1 (N2806, N2805);
not NOT1 (N2807, N2795);
buf BUF1 (N2808, N2781);
and AND2 (N2809, N2791, N1042);
and AND2 (N2810, N2796, N162);
nand NAND2 (N2811, N2806, N1799);
nor NOR4 (N2812, N2811, N2112, N2695, N2791);
and AND3 (N2813, N2784, N206, N1194);
nor NOR4 (N2814, N2794, N919, N1429, N1681);
not NOT1 (N2815, N2808);
not NOT1 (N2816, N2810);
nand NAND2 (N2817, N2803, N1742);
nand NAND2 (N2818, N2809, N2042);
or OR4 (N2819, N2812, N1807, N514, N12);
nor NOR3 (N2820, N2814, N2604, N879);
or OR4 (N2821, N2813, N2284, N1595, N915);
buf BUF1 (N2822, N2802);
nor NOR4 (N2823, N2821, N1024, N77, N742);
not NOT1 (N2824, N2817);
xor XOR2 (N2825, N2823, N1934);
buf BUF1 (N2826, N2815);
nor NOR3 (N2827, N2819, N1510, N1655);
buf BUF1 (N2828, N2822);
xor XOR2 (N2829, N2828, N1983);
nor NOR2 (N2830, N2824, N390);
nand NAND3 (N2831, N2827, N2007, N1405);
xor XOR2 (N2832, N2820, N1109);
nor NOR2 (N2833, N2826, N1127);
xor XOR2 (N2834, N2831, N2588);
nand NAND2 (N2835, N2825, N1311);
and AND3 (N2836, N2816, N2809, N1661);
not NOT1 (N2837, N2835);
nand NAND3 (N2838, N2837, N1815, N549);
or OR2 (N2839, N2829, N468);
and AND2 (N2840, N2830, N2189);
xor XOR2 (N2841, N2832, N2605);
and AND4 (N2842, N2838, N1517, N1608, N2461);
not NOT1 (N2843, N2841);
xor XOR2 (N2844, N2800, N859);
not NOT1 (N2845, N2844);
nand NAND3 (N2846, N2836, N2223, N1434);
and AND2 (N2847, N2818, N1711);
buf BUF1 (N2848, N2833);
and AND3 (N2849, N2845, N1358, N1922);
buf BUF1 (N2850, N2849);
buf BUF1 (N2851, N2834);
nand NAND4 (N2852, N2842, N768, N1847, N2666);
not NOT1 (N2853, N2847);
not NOT1 (N2854, N2848);
nor NOR2 (N2855, N2850, N2749);
or OR2 (N2856, N2843, N1945);
and AND4 (N2857, N2851, N1014, N1172, N510);
nor NOR2 (N2858, N2839, N2218);
buf BUF1 (N2859, N2858);
xor XOR2 (N2860, N2840, N2371);
xor XOR2 (N2861, N2855, N614);
nor NOR2 (N2862, N2856, N231);
buf BUF1 (N2863, N2846);
not NOT1 (N2864, N2853);
not NOT1 (N2865, N2854);
xor XOR2 (N2866, N2862, N2029);
not NOT1 (N2867, N2863);
xor XOR2 (N2868, N2807, N1850);
xor XOR2 (N2869, N2865, N719);
or OR2 (N2870, N2857, N2420);
xor XOR2 (N2871, N2860, N1677);
buf BUF1 (N2872, N2871);
and AND2 (N2873, N2859, N2529);
buf BUF1 (N2874, N2864);
nor NOR3 (N2875, N2868, N1725, N2358);
xor XOR2 (N2876, N2875, N2404);
nand NAND2 (N2877, N2861, N2258);
xor XOR2 (N2878, N2869, N1358);
nand NAND4 (N2879, N2874, N499, N2312, N410);
buf BUF1 (N2880, N2876);
nor NOR4 (N2881, N2878, N2024, N2179, N527);
xor XOR2 (N2882, N2866, N1076);
nand NAND4 (N2883, N2873, N1326, N1623, N2441);
and AND3 (N2884, N2879, N700, N1174);
or OR2 (N2885, N2881, N413);
buf BUF1 (N2886, N2867);
or OR4 (N2887, N2872, N2851, N930, N2779);
xor XOR2 (N2888, N2870, N2075);
not NOT1 (N2889, N2880);
and AND4 (N2890, N2889, N1249, N1925, N1128);
not NOT1 (N2891, N2886);
nor NOR2 (N2892, N2890, N2805);
nor NOR2 (N2893, N2883, N1848);
xor XOR2 (N2894, N2882, N1413);
nor NOR2 (N2895, N2877, N2468);
xor XOR2 (N2896, N2891, N1432);
nand NAND4 (N2897, N2895, N2651, N1394, N230);
not NOT1 (N2898, N2888);
not NOT1 (N2899, N2896);
and AND4 (N2900, N2884, N1749, N2314, N2247);
nand NAND3 (N2901, N2887, N212, N2813);
and AND2 (N2902, N2892, N1702);
xor XOR2 (N2903, N2898, N1660);
or OR4 (N2904, N2903, N587, N1141, N2151);
nor NOR2 (N2905, N2893, N1486);
or OR2 (N2906, N2897, N1787);
and AND4 (N2907, N2899, N1470, N1791, N2166);
nor NOR4 (N2908, N2905, N1594, N967, N151);
nor NOR3 (N2909, N2902, N1824, N828);
and AND4 (N2910, N2906, N831, N884, N299);
buf BUF1 (N2911, N2885);
xor XOR2 (N2912, N2901, N2274);
nor NOR4 (N2913, N2852, N2497, N1741, N1893);
and AND4 (N2914, N2913, N2546, N995, N2154);
and AND4 (N2915, N2909, N1087, N157, N1856);
buf BUF1 (N2916, N2894);
xor XOR2 (N2917, N2900, N473);
xor XOR2 (N2918, N2910, N1104);
or OR2 (N2919, N2915, N1643);
buf BUF1 (N2920, N2916);
not NOT1 (N2921, N2918);
and AND4 (N2922, N2904, N732, N961, N2761);
and AND3 (N2923, N2917, N1410, N1865);
nor NOR2 (N2924, N2921, N2025);
and AND4 (N2925, N2920, N797, N2879, N836);
or OR4 (N2926, N2924, N486, N2851, N1711);
buf BUF1 (N2927, N2926);
and AND2 (N2928, N2923, N376);
xor XOR2 (N2929, N2911, N1552);
nand NAND2 (N2930, N2929, N2742);
or OR4 (N2931, N2928, N202, N814, N1232);
and AND2 (N2932, N2922, N726);
not NOT1 (N2933, N2912);
nor NOR4 (N2934, N2930, N1768, N1708, N1158);
not NOT1 (N2935, N2927);
nand NAND2 (N2936, N2932, N2927);
buf BUF1 (N2937, N2935);
nor NOR4 (N2938, N2907, N2768, N2896, N2864);
not NOT1 (N2939, N2925);
and AND2 (N2940, N2939, N108);
nand NAND3 (N2941, N2919, N129, N516);
nor NOR3 (N2942, N2936, N2125, N2902);
nor NOR3 (N2943, N2914, N2922, N608);
or OR3 (N2944, N2937, N1913, N27);
buf BUF1 (N2945, N2942);
or OR3 (N2946, N2941, N1356, N1186);
nor NOR2 (N2947, N2908, N2921);
nand NAND2 (N2948, N2946, N1234);
or OR2 (N2949, N2944, N1233);
buf BUF1 (N2950, N2934);
xor XOR2 (N2951, N2933, N1543);
not NOT1 (N2952, N2943);
xor XOR2 (N2953, N2940, N26);
and AND4 (N2954, N2938, N248, N966, N1710);
and AND3 (N2955, N2953, N1914, N2118);
buf BUF1 (N2956, N2951);
buf BUF1 (N2957, N2952);
buf BUF1 (N2958, N2956);
buf BUF1 (N2959, N2958);
xor XOR2 (N2960, N2949, N957);
and AND3 (N2961, N2945, N1436, N439);
nand NAND2 (N2962, N2948, N1771);
xor XOR2 (N2963, N2955, N1197);
xor XOR2 (N2964, N2959, N2016);
nand NAND4 (N2965, N2961, N998, N2067, N2459);
nand NAND3 (N2966, N2965, N1676, N2812);
and AND2 (N2967, N2963, N2239);
nor NOR4 (N2968, N2966, N1331, N391, N1529);
or OR2 (N2969, N2960, N1331);
nand NAND3 (N2970, N2947, N99, N2814);
xor XOR2 (N2971, N2954, N2934);
nand NAND2 (N2972, N2957, N882);
or OR3 (N2973, N2950, N2098, N1430);
nor NOR2 (N2974, N2962, N2287);
and AND3 (N2975, N2972, N419, N2886);
and AND4 (N2976, N2931, N1693, N624, N2835);
xor XOR2 (N2977, N2969, N1004);
nand NAND2 (N2978, N2971, N798);
not NOT1 (N2979, N2976);
buf BUF1 (N2980, N2974);
nor NOR2 (N2981, N2977, N1172);
buf BUF1 (N2982, N2968);
xor XOR2 (N2983, N2979, N2399);
nor NOR2 (N2984, N2975, N452);
nand NAND3 (N2985, N2980, N211, N1354);
nand NAND4 (N2986, N2985, N63, N2169, N2648);
nor NOR2 (N2987, N2964, N2931);
xor XOR2 (N2988, N2970, N396);
and AND4 (N2989, N2983, N2615, N2466, N1672);
and AND2 (N2990, N2987, N1651);
nor NOR3 (N2991, N2967, N2973, N1893);
xor XOR2 (N2992, N2758, N642);
and AND3 (N2993, N2991, N747, N839);
and AND3 (N2994, N2982, N1765, N150);
not NOT1 (N2995, N2994);
buf BUF1 (N2996, N2995);
buf BUF1 (N2997, N2984);
xor XOR2 (N2998, N2997, N1619);
buf BUF1 (N2999, N2996);
nand NAND3 (N3000, N2990, N1002, N1870);
nor NOR3 (N3001, N2981, N2511, N818);
not NOT1 (N3002, N2992);
nor NOR3 (N3003, N3000, N840, N720);
nor NOR3 (N3004, N2989, N941, N400);
not NOT1 (N3005, N3004);
buf BUF1 (N3006, N2986);
not NOT1 (N3007, N3003);
nand NAND3 (N3008, N3001, N1506, N2452);
not NOT1 (N3009, N3007);
nand NAND2 (N3010, N3009, N2606);
buf BUF1 (N3011, N3010);
nor NOR3 (N3012, N3006, N1721, N635);
xor XOR2 (N3013, N2993, N2849);
and AND3 (N3014, N2988, N840, N2925);
nor NOR4 (N3015, N3002, N1914, N2781, N2351);
xor XOR2 (N3016, N3008, N2355);
not NOT1 (N3017, N2999);
and AND3 (N3018, N3016, N2158, N2441);
and AND3 (N3019, N3005, N2852, N932);
nor NOR2 (N3020, N3015, N1872);
not NOT1 (N3021, N3011);
nor NOR4 (N3022, N3021, N2507, N2990, N1803);
nand NAND2 (N3023, N3019, N299);
and AND2 (N3024, N3018, N2823);
not NOT1 (N3025, N2998);
xor XOR2 (N3026, N2978, N1197);
or OR2 (N3027, N3022, N1040);
nand NAND4 (N3028, N3026, N2257, N2090, N1590);
and AND3 (N3029, N3024, N1715, N1894);
not NOT1 (N3030, N3027);
or OR3 (N3031, N3028, N2424, N582);
nand NAND2 (N3032, N3020, N1200);
nor NOR2 (N3033, N3017, N815);
nand NAND4 (N3034, N3031, N216, N2747, N2896);
buf BUF1 (N3035, N3013);
or OR2 (N3036, N3034, N1989);
and AND4 (N3037, N3032, N1019, N43, N899);
buf BUF1 (N3038, N3030);
buf BUF1 (N3039, N3014);
and AND2 (N3040, N3039, N737);
nand NAND4 (N3041, N3036, N2970, N2393, N58);
nand NAND4 (N3042, N3035, N162, N747, N2884);
xor XOR2 (N3043, N3025, N2656);
nand NAND2 (N3044, N3042, N1348);
nand NAND2 (N3045, N3012, N1158);
buf BUF1 (N3046, N3037);
buf BUF1 (N3047, N3033);
nor NOR2 (N3048, N3038, N1865);
or OR2 (N3049, N3023, N325);
nor NOR2 (N3050, N3043, N145);
nor NOR3 (N3051, N3049, N651, N2380);
and AND3 (N3052, N3048, N2706, N1908);
xor XOR2 (N3053, N3051, N1426);
and AND2 (N3054, N3047, N3017);
or OR3 (N3055, N3052, N24, N1120);
xor XOR2 (N3056, N3046, N1948);
xor XOR2 (N3057, N3045, N2532);
nor NOR2 (N3058, N3044, N2545);
not NOT1 (N3059, N3054);
or OR4 (N3060, N3053, N2177, N1330, N27);
nor NOR2 (N3061, N3050, N2011);
or OR4 (N3062, N3041, N1857, N1987, N2738);
nand NAND4 (N3063, N3060, N20, N1062, N482);
or OR2 (N3064, N3040, N826);
nor NOR2 (N3065, N3029, N1876);
not NOT1 (N3066, N3062);
and AND4 (N3067, N3061, N2626, N1183, N2955);
nand NAND4 (N3068, N3066, N771, N2475, N1421);
nand NAND4 (N3069, N3056, N862, N1208, N2317);
xor XOR2 (N3070, N3068, N1113);
buf BUF1 (N3071, N3064);
or OR2 (N3072, N3067, N911);
and AND2 (N3073, N3069, N394);
buf BUF1 (N3074, N3072);
not NOT1 (N3075, N3071);
or OR4 (N3076, N3055, N2273, N610, N704);
not NOT1 (N3077, N3074);
nor NOR2 (N3078, N3059, N545);
or OR2 (N3079, N3065, N2279);
not NOT1 (N3080, N3058);
nor NOR2 (N3081, N3076, N29);
buf BUF1 (N3082, N3079);
not NOT1 (N3083, N3070);
and AND4 (N3084, N3082, N176, N1312, N2103);
xor XOR2 (N3085, N3083, N953);
xor XOR2 (N3086, N3057, N1724);
xor XOR2 (N3087, N3084, N1359);
buf BUF1 (N3088, N3081);
buf BUF1 (N3089, N3085);
nand NAND3 (N3090, N3073, N2619, N1854);
xor XOR2 (N3091, N3089, N1261);
nand NAND2 (N3092, N3090, N1236);
not NOT1 (N3093, N3088);
or OR4 (N3094, N3086, N2198, N2925, N1609);
not NOT1 (N3095, N3077);
not NOT1 (N3096, N3075);
nor NOR4 (N3097, N3094, N696, N2776, N2551);
buf BUF1 (N3098, N3093);
buf BUF1 (N3099, N3087);
nand NAND2 (N3100, N3063, N1269);
xor XOR2 (N3101, N3098, N1318);
buf BUF1 (N3102, N3101);
nor NOR4 (N3103, N3095, N686, N2545, N1993);
xor XOR2 (N3104, N3103, N872);
not NOT1 (N3105, N3104);
or OR2 (N3106, N3102, N2252);
nor NOR2 (N3107, N3097, N521);
nand NAND4 (N3108, N3107, N1644, N2791, N1384);
buf BUF1 (N3109, N3092);
nand NAND3 (N3110, N3078, N400, N694);
or OR3 (N3111, N3106, N2516, N2612);
nor NOR3 (N3112, N3091, N1423, N3061);
not NOT1 (N3113, N3096);
buf BUF1 (N3114, N3099);
xor XOR2 (N3115, N3080, N2875);
xor XOR2 (N3116, N3105, N357);
not NOT1 (N3117, N3114);
nor NOR2 (N3118, N3111, N1028);
nor NOR2 (N3119, N3118, N2169);
buf BUF1 (N3120, N3100);
and AND3 (N3121, N3116, N2841, N1418);
or OR4 (N3122, N3109, N283, N2276, N808);
nand NAND3 (N3123, N3112, N3022, N2848);
and AND4 (N3124, N3123, N708, N204, N2328);
and AND4 (N3125, N3110, N3089, N1355, N1674);
or OR3 (N3126, N3121, N997, N100);
not NOT1 (N3127, N3126);
nand NAND2 (N3128, N3115, N2756);
buf BUF1 (N3129, N3125);
or OR4 (N3130, N3117, N1761, N602, N1462);
nand NAND4 (N3131, N3108, N502, N337, N957);
nor NOR2 (N3132, N3131, N721);
nand NAND3 (N3133, N3129, N574, N226);
and AND4 (N3134, N3119, N278, N2665, N1343);
buf BUF1 (N3135, N3120);
buf BUF1 (N3136, N3127);
buf BUF1 (N3137, N3133);
and AND2 (N3138, N3137, N2472);
xor XOR2 (N3139, N3138, N100);
or OR3 (N3140, N3124, N1561, N1483);
xor XOR2 (N3141, N3132, N445);
nand NAND2 (N3142, N3135, N720);
not NOT1 (N3143, N3142);
nor NOR3 (N3144, N3113, N1621, N2678);
not NOT1 (N3145, N3141);
or OR2 (N3146, N3140, N1251);
or OR3 (N3147, N3146, N867, N1614);
not NOT1 (N3148, N3144);
or OR4 (N3149, N3139, N253, N481, N1153);
or OR3 (N3150, N3148, N675, N223);
nand NAND3 (N3151, N3122, N2243, N2319);
nor NOR4 (N3152, N3145, N1391, N2585, N1397);
nand NAND2 (N3153, N3150, N1913);
nand NAND4 (N3154, N3149, N242, N187, N2595);
or OR4 (N3155, N3134, N92, N2734, N2699);
or OR4 (N3156, N3130, N497, N2101, N2144);
not NOT1 (N3157, N3151);
and AND3 (N3158, N3157, N2198, N2804);
nand NAND4 (N3159, N3153, N732, N2179, N1113);
and AND3 (N3160, N3147, N2513, N836);
or OR2 (N3161, N3128, N2985);
nand NAND3 (N3162, N3160, N6, N3141);
not NOT1 (N3163, N3143);
xor XOR2 (N3164, N3158, N2525);
and AND3 (N3165, N3161, N1778, N1691);
not NOT1 (N3166, N3156);
not NOT1 (N3167, N3136);
buf BUF1 (N3168, N3162);
not NOT1 (N3169, N3168);
not NOT1 (N3170, N3154);
buf BUF1 (N3171, N3159);
nor NOR4 (N3172, N3170, N2384, N411, N803);
nor NOR2 (N3173, N3164, N1036);
not NOT1 (N3174, N3169);
or OR2 (N3175, N3165, N939);
or OR2 (N3176, N3166, N1188);
buf BUF1 (N3177, N3155);
and AND3 (N3178, N3172, N438, N1549);
not NOT1 (N3179, N3173);
not NOT1 (N3180, N3177);
buf BUF1 (N3181, N3175);
or OR3 (N3182, N3180, N179, N1195);
and AND3 (N3183, N3167, N1971, N1025);
or OR3 (N3184, N3182, N2999, N2021);
xor XOR2 (N3185, N3163, N61);
or OR2 (N3186, N3184, N694);
nand NAND4 (N3187, N3174, N293, N1636, N2698);
and AND2 (N3188, N3179, N536);
and AND4 (N3189, N3187, N2205, N2497, N215);
xor XOR2 (N3190, N3189, N1064);
or OR3 (N3191, N3176, N1985, N644);
not NOT1 (N3192, N3183);
xor XOR2 (N3193, N3188, N1186);
and AND2 (N3194, N3186, N280);
xor XOR2 (N3195, N3171, N2184);
buf BUF1 (N3196, N3178);
and AND2 (N3197, N3181, N2141);
nand NAND2 (N3198, N3191, N1966);
nor NOR4 (N3199, N3185, N1900, N2980, N815);
buf BUF1 (N3200, N3198);
xor XOR2 (N3201, N3200, N2964);
buf BUF1 (N3202, N3197);
buf BUF1 (N3203, N3202);
or OR4 (N3204, N3192, N2343, N1458, N761);
and AND4 (N3205, N3199, N1143, N125, N1771);
nand NAND4 (N3206, N3196, N3024, N1063, N2284);
or OR4 (N3207, N3203, N2348, N177, N1806);
xor XOR2 (N3208, N3204, N885);
nand NAND4 (N3209, N3190, N1090, N102, N1223);
not NOT1 (N3210, N3206);
not NOT1 (N3211, N3193);
and AND3 (N3212, N3210, N725, N1904);
not NOT1 (N3213, N3209);
xor XOR2 (N3214, N3201, N1503);
xor XOR2 (N3215, N3208, N602);
or OR3 (N3216, N3213, N761, N543);
not NOT1 (N3217, N3211);
buf BUF1 (N3218, N3152);
or OR3 (N3219, N3195, N2787, N935);
nand NAND3 (N3220, N3212, N1129, N2682);
nand NAND2 (N3221, N3220, N1153);
not NOT1 (N3222, N3216);
not NOT1 (N3223, N3219);
buf BUF1 (N3224, N3215);
not NOT1 (N3225, N3194);
not NOT1 (N3226, N3224);
nor NOR4 (N3227, N3226, N1791, N1406, N2337);
and AND4 (N3228, N3222, N3017, N1379, N3195);
not NOT1 (N3229, N3227);
and AND2 (N3230, N3218, N1360);
buf BUF1 (N3231, N3221);
or OR3 (N3232, N3217, N1232, N491);
xor XOR2 (N3233, N3228, N2460);
nor NOR3 (N3234, N3223, N2578, N506);
nand NAND3 (N3235, N3225, N1118, N1258);
and AND3 (N3236, N3214, N1308, N2858);
not NOT1 (N3237, N3233);
xor XOR2 (N3238, N3207, N2390);
or OR2 (N3239, N3237, N2202);
and AND3 (N3240, N3239, N1227, N200);
nor NOR3 (N3241, N3240, N1297, N1752);
buf BUF1 (N3242, N3232);
not NOT1 (N3243, N3234);
nand NAND3 (N3244, N3241, N2095, N2155);
buf BUF1 (N3245, N3235);
nand NAND4 (N3246, N3242, N1099, N1776, N2878);
not NOT1 (N3247, N3246);
and AND3 (N3248, N3205, N3194, N937);
not NOT1 (N3249, N3243);
not NOT1 (N3250, N3238);
not NOT1 (N3251, N3230);
buf BUF1 (N3252, N3249);
not NOT1 (N3253, N3231);
and AND3 (N3254, N3244, N886, N2242);
and AND4 (N3255, N3252, N1624, N1166, N788);
or OR3 (N3256, N3254, N1527, N2277);
buf BUF1 (N3257, N3229);
xor XOR2 (N3258, N3257, N54);
nor NOR2 (N3259, N3256, N15);
nor NOR3 (N3260, N3236, N541, N2486);
not NOT1 (N3261, N3259);
or OR3 (N3262, N3245, N16, N2085);
nor NOR4 (N3263, N3250, N2332, N986, N410);
or OR4 (N3264, N3261, N653, N466, N3118);
not NOT1 (N3265, N3260);
buf BUF1 (N3266, N3255);
nand NAND2 (N3267, N3251, N457);
nor NOR2 (N3268, N3265, N2913);
not NOT1 (N3269, N3264);
not NOT1 (N3270, N3258);
nand NAND3 (N3271, N3253, N3074, N3053);
nor NOR3 (N3272, N3263, N2096, N420);
nor NOR3 (N3273, N3248, N2927, N3097);
not NOT1 (N3274, N3268);
xor XOR2 (N3275, N3270, N320);
not NOT1 (N3276, N3247);
and AND4 (N3277, N3276, N590, N450, N1534);
nor NOR4 (N3278, N3267, N2447, N2092, N2378);
nor NOR2 (N3279, N3273, N110);
buf BUF1 (N3280, N3266);
or OR3 (N3281, N3272, N2342, N2870);
nor NOR4 (N3282, N3279, N514, N3082, N3179);
not NOT1 (N3283, N3282);
buf BUF1 (N3284, N3278);
or OR3 (N3285, N3262, N457, N580);
not NOT1 (N3286, N3277);
and AND3 (N3287, N3274, N605, N318);
xor XOR2 (N3288, N3275, N1597);
or OR4 (N3289, N3284, N272, N380, N478);
and AND3 (N3290, N3289, N1283, N3118);
nor NOR3 (N3291, N3281, N318, N2140);
nand NAND2 (N3292, N3269, N1664);
nor NOR4 (N3293, N3291, N2710, N494, N2591);
xor XOR2 (N3294, N3271, N1996);
nand NAND3 (N3295, N3288, N653, N151);
and AND3 (N3296, N3287, N3069, N906);
nor NOR3 (N3297, N3280, N1964, N1953);
and AND3 (N3298, N3297, N2144, N833);
buf BUF1 (N3299, N3294);
not NOT1 (N3300, N3292);
nand NAND4 (N3301, N3283, N2510, N1842, N2908);
nor NOR4 (N3302, N3295, N2587, N714, N1043);
xor XOR2 (N3303, N3290, N1751);
buf BUF1 (N3304, N3300);
buf BUF1 (N3305, N3296);
nor NOR2 (N3306, N3302, N2794);
or OR2 (N3307, N3293, N2450);
buf BUF1 (N3308, N3307);
nand NAND3 (N3309, N3299, N1432, N1542);
or OR3 (N3310, N3308, N1751, N2526);
nand NAND3 (N3311, N3304, N1239, N1436);
xor XOR2 (N3312, N3285, N3251);
nor NOR4 (N3313, N3311, N2986, N667, N2143);
nand NAND4 (N3314, N3312, N3009, N70, N825);
nor NOR4 (N3315, N3303, N2795, N1068, N2517);
nor NOR3 (N3316, N3313, N1136, N783);
nand NAND3 (N3317, N3314, N2200, N1055);
or OR3 (N3318, N3286, N1516, N2916);
nor NOR3 (N3319, N3316, N1608, N401);
and AND3 (N3320, N3319, N1660, N1153);
nor NOR4 (N3321, N3320, N2775, N426, N2481);
xor XOR2 (N3322, N3310, N922);
buf BUF1 (N3323, N3301);
buf BUF1 (N3324, N3306);
nor NOR2 (N3325, N3305, N965);
or OR3 (N3326, N3317, N1116, N681);
not NOT1 (N3327, N3315);
nand NAND2 (N3328, N3324, N913);
nor NOR4 (N3329, N3327, N2678, N750, N3057);
nand NAND2 (N3330, N3323, N60);
or OR4 (N3331, N3326, N2211, N1123, N1695);
buf BUF1 (N3332, N3328);
nor NOR4 (N3333, N3331, N1861, N1846, N3021);
or OR3 (N3334, N3332, N514, N1074);
nor NOR4 (N3335, N3325, N988, N2230, N160);
and AND2 (N3336, N3321, N3007);
not NOT1 (N3337, N3298);
xor XOR2 (N3338, N3334, N2352);
nand NAND2 (N3339, N3338, N1531);
or OR3 (N3340, N3336, N2006, N2070);
nor NOR3 (N3341, N3339, N2444, N295);
not NOT1 (N3342, N3337);
nor NOR2 (N3343, N3329, N2731);
xor XOR2 (N3344, N3343, N1977);
and AND4 (N3345, N3322, N1279, N1531, N3236);
and AND2 (N3346, N3345, N1026);
not NOT1 (N3347, N3335);
nand NAND2 (N3348, N3340, N3277);
and AND3 (N3349, N3333, N3090, N241);
buf BUF1 (N3350, N3344);
nand NAND3 (N3351, N3330, N407, N726);
buf BUF1 (N3352, N3346);
buf BUF1 (N3353, N3351);
or OR3 (N3354, N3348, N1782, N1474);
nor NOR2 (N3355, N3349, N2025);
nor NOR4 (N3356, N3354, N3084, N2348, N2062);
and AND2 (N3357, N3342, N3124);
nor NOR2 (N3358, N3353, N462);
nand NAND3 (N3359, N3350, N138, N2564);
nand NAND3 (N3360, N3347, N1714, N1014);
nand NAND4 (N3361, N3358, N3131, N2, N3052);
and AND4 (N3362, N3357, N730, N1393, N2905);
xor XOR2 (N3363, N3309, N2561);
buf BUF1 (N3364, N3362);
buf BUF1 (N3365, N3360);
and AND2 (N3366, N3361, N1257);
nand NAND3 (N3367, N3365, N1904, N1277);
or OR4 (N3368, N3355, N1843, N517, N3045);
not NOT1 (N3369, N3352);
buf BUF1 (N3370, N3369);
nand NAND4 (N3371, N3368, N1526, N2858, N3016);
nor NOR3 (N3372, N3370, N899, N417);
or OR2 (N3373, N3371, N2831);
and AND2 (N3374, N3363, N595);
buf BUF1 (N3375, N3367);
or OR3 (N3376, N3341, N440, N1547);
and AND2 (N3377, N3364, N2530);
and AND3 (N3378, N3359, N1821, N2833);
buf BUF1 (N3379, N3372);
nand NAND2 (N3380, N3366, N3127);
buf BUF1 (N3381, N3374);
buf BUF1 (N3382, N3379);
nand NAND3 (N3383, N3375, N2725, N2374);
and AND3 (N3384, N3378, N2386, N643);
not NOT1 (N3385, N3381);
buf BUF1 (N3386, N3377);
buf BUF1 (N3387, N3384);
not NOT1 (N3388, N3386);
buf BUF1 (N3389, N3385);
not NOT1 (N3390, N3389);
xor XOR2 (N3391, N3376, N3234);
nand NAND2 (N3392, N3382, N10);
or OR3 (N3393, N3391, N2712, N2392);
not NOT1 (N3394, N3388);
and AND2 (N3395, N3380, N569);
buf BUF1 (N3396, N3392);
nor NOR4 (N3397, N3318, N1837, N92, N61);
not NOT1 (N3398, N3394);
nor NOR2 (N3399, N3387, N2622);
and AND2 (N3400, N3396, N2998);
or OR2 (N3401, N3393, N28);
not NOT1 (N3402, N3398);
not NOT1 (N3403, N3383);
nand NAND2 (N3404, N3397, N2999);
and AND4 (N3405, N3399, N2465, N274, N519);
and AND3 (N3406, N3401, N2830, N1450);
nor NOR3 (N3407, N3373, N3295, N1244);
nor NOR4 (N3408, N3402, N1283, N2661, N1642);
and AND4 (N3409, N3403, N2959, N2236, N917);
nor NOR3 (N3410, N3404, N2769, N1785);
and AND2 (N3411, N3405, N666);
nand NAND3 (N3412, N3408, N2051, N888);
nand NAND2 (N3413, N3412, N3314);
xor XOR2 (N3414, N3356, N494);
not NOT1 (N3415, N3411);
nand NAND3 (N3416, N3395, N2235, N2088);
buf BUF1 (N3417, N3414);
nor NOR2 (N3418, N3413, N2933);
and AND4 (N3419, N3417, N3376, N2260, N602);
nand NAND3 (N3420, N3409, N2335, N2423);
nor NOR4 (N3421, N3390, N1958, N884, N3298);
nor NOR4 (N3422, N3419, N730, N74, N107);
nor NOR4 (N3423, N3420, N586, N2656, N17);
buf BUF1 (N3424, N3416);
and AND3 (N3425, N3410, N3172, N2604);
buf BUF1 (N3426, N3400);
not NOT1 (N3427, N3418);
buf BUF1 (N3428, N3423);
not NOT1 (N3429, N3427);
not NOT1 (N3430, N3426);
buf BUF1 (N3431, N3406);
xor XOR2 (N3432, N3421, N3365);
or OR4 (N3433, N3424, N1955, N3134, N1033);
nor NOR2 (N3434, N3415, N643);
buf BUF1 (N3435, N3434);
and AND2 (N3436, N3429, N2731);
nand NAND3 (N3437, N3407, N2757, N1140);
nand NAND3 (N3438, N3425, N24, N897);
buf BUF1 (N3439, N3437);
not NOT1 (N3440, N3430);
xor XOR2 (N3441, N3433, N2408);
buf BUF1 (N3442, N3436);
and AND3 (N3443, N3442, N970, N2181);
and AND4 (N3444, N3435, N2132, N2807, N2563);
buf BUF1 (N3445, N3444);
or OR2 (N3446, N3441, N2275);
nand NAND3 (N3447, N3440, N2450, N1986);
and AND3 (N3448, N3428, N346, N247);
nor NOR3 (N3449, N3432, N1440, N2491);
or OR3 (N3450, N3445, N2149, N935);
not NOT1 (N3451, N3443);
xor XOR2 (N3452, N3450, N33);
and AND3 (N3453, N3448, N3395, N2340);
buf BUF1 (N3454, N3447);
or OR4 (N3455, N3451, N1148, N1005, N436);
xor XOR2 (N3456, N3431, N871);
or OR4 (N3457, N3422, N2013, N1684, N517);
and AND4 (N3458, N3455, N1445, N190, N7);
xor XOR2 (N3459, N3449, N2472);
nor NOR2 (N3460, N3457, N514);
or OR4 (N3461, N3453, N2143, N587, N1451);
nand NAND3 (N3462, N3456, N1761, N1246);
nand NAND2 (N3463, N3438, N1589);
or OR2 (N3464, N3460, N2021);
xor XOR2 (N3465, N3459, N1029);
xor XOR2 (N3466, N3454, N1513);
nand NAND3 (N3467, N3465, N1428, N773);
not NOT1 (N3468, N3458);
or OR2 (N3469, N3464, N2616);
and AND2 (N3470, N3446, N1244);
not NOT1 (N3471, N3468);
not NOT1 (N3472, N3470);
nand NAND3 (N3473, N3439, N1627, N278);
not NOT1 (N3474, N3467);
nor NOR4 (N3475, N3473, N3198, N718, N572);
not NOT1 (N3476, N3466);
nor NOR3 (N3477, N3461, N1780, N388);
and AND3 (N3478, N3469, N821, N1718);
not NOT1 (N3479, N3476);
or OR3 (N3480, N3462, N2739, N3424);
nand NAND2 (N3481, N3474, N2412);
xor XOR2 (N3482, N3475, N2764);
nor NOR2 (N3483, N3452, N368);
or OR4 (N3484, N3482, N2121, N132, N1594);
buf BUF1 (N3485, N3483);
xor XOR2 (N3486, N3480, N1887);
or OR4 (N3487, N3481, N652, N2005, N2657);
and AND3 (N3488, N3479, N2221, N265);
buf BUF1 (N3489, N3488);
nand NAND4 (N3490, N3485, N3157, N3249, N1277);
nand NAND3 (N3491, N3487, N2310, N2863);
not NOT1 (N3492, N3477);
or OR3 (N3493, N3490, N3369, N1908);
or OR2 (N3494, N3492, N1799);
nand NAND2 (N3495, N3478, N898);
and AND3 (N3496, N3463, N3417, N1425);
nor NOR2 (N3497, N3484, N2590);
nor NOR3 (N3498, N3493, N1489, N1877);
and AND3 (N3499, N3472, N256, N2238);
and AND3 (N3500, N3495, N2048, N2881);
and AND4 (N3501, N3491, N827, N1271, N2360);
and AND3 (N3502, N3499, N1829, N3339);
nand NAND2 (N3503, N3500, N1695);
buf BUF1 (N3504, N3502);
buf BUF1 (N3505, N3497);
and AND3 (N3506, N3501, N597, N493);
nor NOR4 (N3507, N3498, N1397, N2814, N1285);
or OR2 (N3508, N3506, N3458);
or OR2 (N3509, N3486, N946);
nand NAND4 (N3510, N3507, N1778, N1137, N1974);
xor XOR2 (N3511, N3504, N2473);
nor NOR2 (N3512, N3511, N1974);
nand NAND3 (N3513, N3496, N786, N1164);
or OR2 (N3514, N3471, N2637);
not NOT1 (N3515, N3509);
nor NOR3 (N3516, N3508, N2282, N940);
buf BUF1 (N3517, N3512);
nand NAND3 (N3518, N3505, N1782, N421);
endmodule