// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N3510,N3508,N3491,N3509,N3503,N3507,N3483,N3504,N3496,N3512;

nand NAND3 (N13, N3, N8, N11);
buf BUF1 (N14, N6);
buf BUF1 (N15, N5);
or OR4 (N16, N4, N3, N11, N12);
nor NOR4 (N17, N2, N13, N16, N8);
buf BUF1 (N18, N14);
nand NAND2 (N19, N2, N5);
xor XOR2 (N20, N1, N9);
nand NAND3 (N21, N3, N6, N14);
xor XOR2 (N22, N1, N21);
nor NOR3 (N23, N20, N1, N16);
xor XOR2 (N24, N19, N1);
xor XOR2 (N25, N5, N1);
nor NOR2 (N26, N1, N23);
nor NOR3 (N27, N12, N21, N11);
nand NAND3 (N28, N20, N18, N5);
nor NOR4 (N29, N2, N12, N22, N16);
xor XOR2 (N30, N24, N8);
or OR4 (N31, N16, N21, N3, N1);
nand NAND4 (N32, N22, N31, N31, N21);
nand NAND4 (N33, N31, N25, N19, N16);
not NOT1 (N34, N26);
xor XOR2 (N35, N20, N19);
nand NAND3 (N36, N35, N32, N11);
not NOT1 (N37, N22);
nand NAND4 (N38, N33, N3, N23, N32);
buf BUF1 (N39, N15);
nand NAND3 (N40, N27, N39, N34);
buf BUF1 (N41, N17);
xor XOR2 (N42, N35, N39);
xor XOR2 (N43, N38, N17);
buf BUF1 (N44, N25);
xor XOR2 (N45, N28, N42);
buf BUF1 (N46, N25);
nor NOR4 (N47, N41, N2, N24, N35);
nand NAND3 (N48, N44, N29, N17);
buf BUF1 (N49, N25);
buf BUF1 (N50, N36);
xor XOR2 (N51, N37, N16);
not NOT1 (N52, N50);
or OR2 (N53, N51, N6);
buf BUF1 (N54, N52);
not NOT1 (N55, N48);
buf BUF1 (N56, N40);
xor XOR2 (N57, N47, N32);
nor NOR2 (N58, N45, N4);
and AND4 (N59, N30, N52, N55, N46);
xor XOR2 (N60, N24, N5);
nand NAND3 (N61, N14, N15, N15);
and AND2 (N62, N58, N10);
buf BUF1 (N63, N57);
buf BUF1 (N64, N54);
buf BUF1 (N65, N61);
nor NOR2 (N66, N43, N59);
nand NAND3 (N67, N26, N6, N49);
and AND4 (N68, N45, N20, N35, N10);
nor NOR2 (N69, N66, N21);
or OR2 (N70, N63, N9);
buf BUF1 (N71, N65);
or OR4 (N72, N67, N34, N55, N29);
and AND3 (N73, N70, N22, N59);
nor NOR3 (N74, N53, N50, N10);
buf BUF1 (N75, N60);
nor NOR4 (N76, N71, N71, N11, N28);
nand NAND3 (N77, N75, N70, N64);
buf BUF1 (N78, N67);
xor XOR2 (N79, N69, N7);
xor XOR2 (N80, N77, N4);
and AND2 (N81, N73, N54);
buf BUF1 (N82, N56);
not NOT1 (N83, N68);
and AND2 (N84, N82, N5);
nand NAND3 (N85, N78, N70, N64);
xor XOR2 (N86, N76, N29);
buf BUF1 (N87, N74);
or OR4 (N88, N85, N1, N73, N7);
not NOT1 (N89, N83);
not NOT1 (N90, N72);
nor NOR2 (N91, N80, N89);
and AND4 (N92, N4, N88, N20, N61);
or OR3 (N93, N85, N91, N88);
buf BUF1 (N94, N62);
buf BUF1 (N95, N50);
nor NOR2 (N96, N92, N3);
and AND2 (N97, N96, N64);
or OR3 (N98, N87, N71, N37);
not NOT1 (N99, N79);
not NOT1 (N100, N94);
buf BUF1 (N101, N93);
nand NAND4 (N102, N84, N99, N60, N91);
or OR4 (N103, N2, N81, N49, N33);
nor NOR2 (N104, N17, N43);
xor XOR2 (N105, N97, N68);
xor XOR2 (N106, N105, N93);
buf BUF1 (N107, N90);
buf BUF1 (N108, N107);
xor XOR2 (N109, N106, N62);
or OR3 (N110, N101, N104, N74);
or OR2 (N111, N84, N73);
or OR4 (N112, N110, N74, N14, N75);
not NOT1 (N113, N103);
nor NOR3 (N114, N98, N38, N1);
nand NAND4 (N115, N108, N87, N34, N49);
or OR3 (N116, N109, N8, N35);
nor NOR3 (N117, N112, N70, N27);
not NOT1 (N118, N113);
buf BUF1 (N119, N115);
xor XOR2 (N120, N111, N17);
xor XOR2 (N121, N86, N66);
nand NAND3 (N122, N114, N39, N102);
buf BUF1 (N123, N99);
nor NOR2 (N124, N117, N57);
nand NAND2 (N125, N118, N66);
and AND4 (N126, N116, N47, N34, N83);
nand NAND4 (N127, N122, N69, N119, N123);
or OR2 (N128, N75, N71);
or OR3 (N129, N21, N32, N35);
and AND2 (N130, N129, N82);
not NOT1 (N131, N125);
nor NOR4 (N132, N127, N128, N52, N32);
xor XOR2 (N133, N66, N97);
nand NAND3 (N134, N121, N61, N68);
xor XOR2 (N135, N134, N19);
and AND3 (N136, N135, N111, N120);
nand NAND4 (N137, N8, N65, N85, N101);
not NOT1 (N138, N133);
nor NOR4 (N139, N131, N3, N11, N113);
nor NOR4 (N140, N95, N97, N5, N9);
nor NOR2 (N141, N137, N66);
nand NAND4 (N142, N139, N128, N94, N116);
xor XOR2 (N143, N142, N115);
not NOT1 (N144, N132);
nand NAND2 (N145, N100, N91);
or OR4 (N146, N141, N131, N129, N47);
nor NOR3 (N147, N138, N116, N65);
xor XOR2 (N148, N126, N140);
nor NOR2 (N149, N110, N31);
buf BUF1 (N150, N143);
or OR3 (N151, N148, N7, N85);
and AND4 (N152, N124, N136, N138, N44);
buf BUF1 (N153, N14);
nand NAND3 (N154, N145, N116, N66);
and AND2 (N155, N154, N149);
nand NAND3 (N156, N93, N128, N1);
nor NOR3 (N157, N153, N58, N152);
nor NOR3 (N158, N13, N25, N98);
nor NOR3 (N159, N150, N138, N84);
buf BUF1 (N160, N155);
xor XOR2 (N161, N158, N69);
nand NAND4 (N162, N146, N21, N87, N31);
or OR4 (N163, N156, N83, N137, N87);
xor XOR2 (N164, N130, N9);
xor XOR2 (N165, N144, N28);
nand NAND2 (N166, N161, N114);
not NOT1 (N167, N157);
buf BUF1 (N168, N162);
nand NAND3 (N169, N168, N109, N70);
not NOT1 (N170, N160);
buf BUF1 (N171, N164);
and AND3 (N172, N147, N7, N41);
and AND2 (N173, N170, N120);
buf BUF1 (N174, N165);
nand NAND2 (N175, N163, N32);
nand NAND2 (N176, N169, N56);
nand NAND3 (N177, N167, N33, N13);
xor XOR2 (N178, N171, N25);
not NOT1 (N179, N173);
xor XOR2 (N180, N174, N99);
and AND4 (N181, N159, N151, N171, N99);
not NOT1 (N182, N120);
not NOT1 (N183, N175);
xor XOR2 (N184, N178, N176);
buf BUF1 (N185, N163);
nor NOR4 (N186, N166, N146, N41, N114);
or OR2 (N187, N185, N77);
buf BUF1 (N188, N186);
xor XOR2 (N189, N180, N46);
and AND3 (N190, N187, N48, N15);
buf BUF1 (N191, N183);
nor NOR4 (N192, N172, N54, N183, N140);
not NOT1 (N193, N177);
xor XOR2 (N194, N193, N158);
and AND2 (N195, N190, N11);
buf BUF1 (N196, N181);
or OR2 (N197, N188, N188);
not NOT1 (N198, N184);
xor XOR2 (N199, N198, N152);
xor XOR2 (N200, N192, N93);
xor XOR2 (N201, N191, N99);
xor XOR2 (N202, N197, N9);
or OR2 (N203, N200, N166);
nand NAND4 (N204, N179, N183, N194, N80);
not NOT1 (N205, N152);
buf BUF1 (N206, N195);
nor NOR3 (N207, N204, N1, N131);
nor NOR4 (N208, N205, N79, N197, N95);
buf BUF1 (N209, N202);
not NOT1 (N210, N196);
nor NOR2 (N211, N182, N58);
nand NAND3 (N212, N189, N148, N190);
not NOT1 (N213, N207);
not NOT1 (N214, N208);
nor NOR4 (N215, N211, N96, N81, N166);
or OR3 (N216, N210, N112, N167);
buf BUF1 (N217, N215);
not NOT1 (N218, N199);
nand NAND3 (N219, N214, N69, N156);
nand NAND3 (N220, N217, N121, N182);
and AND3 (N221, N218, N86, N22);
or OR3 (N222, N209, N192, N107);
not NOT1 (N223, N219);
and AND4 (N224, N212, N166, N70, N117);
and AND2 (N225, N203, N107);
or OR4 (N226, N206, N87, N173, N180);
buf BUF1 (N227, N221);
xor XOR2 (N228, N201, N169);
nand NAND4 (N229, N226, N119, N72, N45);
nand NAND3 (N230, N228, N74, N183);
nor NOR3 (N231, N229, N170, N57);
nand NAND2 (N232, N220, N39);
or OR4 (N233, N223, N101, N195, N10);
and AND4 (N234, N224, N203, N72, N15);
nand NAND3 (N235, N213, N4, N211);
and AND3 (N236, N232, N12, N174);
not NOT1 (N237, N225);
nor NOR2 (N238, N233, N183);
nor NOR4 (N239, N230, N84, N131, N135);
nand NAND4 (N240, N231, N87, N52, N164);
nor NOR4 (N241, N240, N41, N196, N108);
nor NOR3 (N242, N234, N89, N169);
xor XOR2 (N243, N241, N132);
and AND4 (N244, N239, N95, N193, N180);
nor NOR4 (N245, N216, N7, N21, N113);
xor XOR2 (N246, N244, N37);
nor NOR2 (N247, N245, N134);
and AND4 (N248, N246, N43, N229, N57);
not NOT1 (N249, N243);
nand NAND4 (N250, N236, N94, N86, N39);
buf BUF1 (N251, N235);
nor NOR3 (N252, N242, N28, N190);
buf BUF1 (N253, N252);
xor XOR2 (N254, N227, N23);
or OR2 (N255, N250, N59);
nand NAND3 (N256, N254, N68, N59);
not NOT1 (N257, N251);
nand NAND4 (N258, N257, N19, N178, N123);
and AND4 (N259, N248, N58, N219, N7);
xor XOR2 (N260, N238, N89);
or OR2 (N261, N237, N106);
or OR2 (N262, N253, N215);
or OR4 (N263, N262, N54, N145, N231);
and AND4 (N264, N258, N254, N23, N143);
nor NOR2 (N265, N256, N152);
not NOT1 (N266, N255);
buf BUF1 (N267, N265);
not NOT1 (N268, N264);
or OR2 (N269, N260, N2);
and AND2 (N270, N266, N196);
nor NOR2 (N271, N268, N55);
nand NAND2 (N272, N247, N104);
nand NAND2 (N273, N267, N43);
not NOT1 (N274, N259);
nand NAND3 (N275, N271, N151, N260);
and AND2 (N276, N269, N187);
xor XOR2 (N277, N275, N167);
xor XOR2 (N278, N249, N69);
and AND3 (N279, N274, N11, N148);
or OR3 (N280, N270, N61, N146);
xor XOR2 (N281, N276, N72);
or OR3 (N282, N278, N73, N255);
not NOT1 (N283, N282);
or OR2 (N284, N281, N119);
nor NOR4 (N285, N261, N261, N45, N265);
or OR2 (N286, N222, N155);
not NOT1 (N287, N280);
buf BUF1 (N288, N286);
or OR4 (N289, N284, N153, N111, N147);
nor NOR3 (N290, N279, N31, N80);
not NOT1 (N291, N287);
or OR3 (N292, N291, N94, N190);
buf BUF1 (N293, N273);
buf BUF1 (N294, N263);
and AND4 (N295, N293, N248, N222, N247);
nand NAND2 (N296, N283, N207);
buf BUF1 (N297, N289);
nor NOR2 (N298, N288, N96);
nand NAND4 (N299, N296, N116, N34, N207);
nor NOR3 (N300, N294, N166, N189);
or OR2 (N301, N297, N295);
not NOT1 (N302, N44);
not NOT1 (N303, N292);
and AND4 (N304, N272, N141, N254, N57);
xor XOR2 (N305, N277, N12);
not NOT1 (N306, N300);
or OR2 (N307, N302, N204);
or OR4 (N308, N305, N185, N45, N19);
and AND4 (N309, N303, N176, N284, N23);
and AND3 (N310, N298, N63, N171);
or OR4 (N311, N306, N21, N273, N203);
nand NAND4 (N312, N309, N34, N88, N302);
buf BUF1 (N313, N285);
nand NAND3 (N314, N301, N113, N152);
not NOT1 (N315, N290);
not NOT1 (N316, N314);
or OR4 (N317, N304, N72, N122, N303);
buf BUF1 (N318, N308);
nand NAND2 (N319, N312, N86);
or OR3 (N320, N318, N193, N112);
or OR4 (N321, N317, N201, N173, N16);
xor XOR2 (N322, N311, N304);
nand NAND4 (N323, N321, N279, N192, N8);
not NOT1 (N324, N322);
xor XOR2 (N325, N323, N173);
nor NOR3 (N326, N299, N129, N70);
not NOT1 (N327, N307);
nand NAND2 (N328, N324, N180);
and AND3 (N329, N326, N116, N165);
not NOT1 (N330, N320);
nand NAND4 (N331, N327, N163, N273, N257);
not NOT1 (N332, N310);
nor NOR4 (N333, N332, N248, N242, N240);
or OR3 (N334, N329, N182, N306);
or OR2 (N335, N333, N160);
not NOT1 (N336, N334);
or OR3 (N337, N313, N73, N156);
xor XOR2 (N338, N315, N215);
and AND4 (N339, N328, N110, N56, N107);
buf BUF1 (N340, N335);
nand NAND2 (N341, N339, N234);
nand NAND4 (N342, N319, N205, N340, N21);
nor NOR4 (N343, N289, N145, N235, N156);
nor NOR4 (N344, N331, N246, N241, N204);
xor XOR2 (N345, N336, N88);
xor XOR2 (N346, N338, N187);
nor NOR3 (N347, N345, N306, N174);
nand NAND2 (N348, N316, N141);
and AND3 (N349, N346, N257, N190);
buf BUF1 (N350, N347);
and AND3 (N351, N342, N288, N57);
xor XOR2 (N352, N343, N321);
not NOT1 (N353, N351);
nand NAND2 (N354, N348, N255);
buf BUF1 (N355, N330);
and AND4 (N356, N350, N171, N84, N191);
nor NOR3 (N357, N337, N96, N328);
xor XOR2 (N358, N354, N230);
nand NAND3 (N359, N356, N158, N43);
nor NOR4 (N360, N352, N251, N244, N35);
xor XOR2 (N361, N341, N32);
buf BUF1 (N362, N349);
not NOT1 (N363, N360);
and AND3 (N364, N355, N107, N105);
nor NOR2 (N365, N325, N160);
and AND3 (N366, N365, N149, N259);
nor NOR2 (N367, N353, N87);
not NOT1 (N368, N362);
nor NOR3 (N369, N359, N280, N255);
buf BUF1 (N370, N358);
nor NOR2 (N371, N366, N111);
and AND4 (N372, N368, N28, N214, N199);
not NOT1 (N373, N370);
not NOT1 (N374, N357);
and AND3 (N375, N361, N189, N264);
or OR2 (N376, N372, N355);
and AND2 (N377, N367, N177);
and AND3 (N378, N376, N226, N15);
or OR3 (N379, N363, N233, N75);
xor XOR2 (N380, N379, N216);
nand NAND4 (N381, N364, N217, N354, N218);
nor NOR4 (N382, N344, N73, N162, N22);
buf BUF1 (N383, N381);
xor XOR2 (N384, N369, N188);
and AND3 (N385, N373, N128, N160);
nor NOR4 (N386, N374, N211, N362, N92);
nand NAND2 (N387, N382, N14);
nand NAND4 (N388, N384, N40, N200, N322);
buf BUF1 (N389, N371);
and AND3 (N390, N378, N65, N281);
xor XOR2 (N391, N386, N153);
and AND3 (N392, N387, N213, N325);
xor XOR2 (N393, N377, N353);
nor NOR2 (N394, N385, N11);
and AND4 (N395, N393, N362, N324, N224);
not NOT1 (N396, N383);
xor XOR2 (N397, N396, N168);
xor XOR2 (N398, N395, N303);
buf BUF1 (N399, N380);
and AND4 (N400, N399, N99, N264, N265);
and AND3 (N401, N391, N163, N59);
xor XOR2 (N402, N392, N303);
xor XOR2 (N403, N388, N277);
or OR4 (N404, N402, N383, N394, N2);
nand NAND4 (N405, N40, N199, N280, N316);
and AND3 (N406, N398, N83, N282);
buf BUF1 (N407, N403);
and AND2 (N408, N390, N387);
xor XOR2 (N409, N407, N183);
nand NAND4 (N410, N397, N70, N311, N368);
xor XOR2 (N411, N409, N151);
xor XOR2 (N412, N404, N187);
or OR3 (N413, N375, N178, N42);
and AND3 (N414, N412, N221, N129);
or OR3 (N415, N410, N5, N326);
not NOT1 (N416, N415);
and AND3 (N417, N416, N199, N181);
xor XOR2 (N418, N406, N210);
or OR3 (N419, N405, N35, N15);
not NOT1 (N420, N417);
nand NAND4 (N421, N411, N369, N31, N299);
buf BUF1 (N422, N421);
nor NOR4 (N423, N419, N88, N260, N97);
xor XOR2 (N424, N413, N377);
and AND4 (N425, N420, N132, N320, N332);
xor XOR2 (N426, N425, N284);
nor NOR2 (N427, N426, N375);
xor XOR2 (N428, N400, N80);
buf BUF1 (N429, N427);
and AND4 (N430, N401, N371, N259, N142);
buf BUF1 (N431, N422);
nand NAND4 (N432, N431, N152, N216, N382);
and AND2 (N433, N424, N293);
nor NOR4 (N434, N432, N87, N289, N106);
buf BUF1 (N435, N408);
and AND3 (N436, N434, N358, N386);
not NOT1 (N437, N433);
nor NOR2 (N438, N436, N197);
nand NAND4 (N439, N428, N111, N276, N423);
xor XOR2 (N440, N233, N176);
not NOT1 (N441, N389);
xor XOR2 (N442, N437, N152);
or OR4 (N443, N440, N367, N355, N39);
nor NOR3 (N444, N430, N190, N289);
nand NAND4 (N445, N438, N146, N200, N439);
or OR2 (N446, N124, N312);
and AND3 (N447, N445, N149, N74);
or OR2 (N448, N429, N361);
buf BUF1 (N449, N435);
or OR4 (N450, N418, N323, N413, N86);
nand NAND2 (N451, N449, N56);
not NOT1 (N452, N447);
not NOT1 (N453, N452);
nand NAND4 (N454, N442, N43, N142, N376);
or OR3 (N455, N448, N148, N254);
nand NAND2 (N456, N443, N36);
buf BUF1 (N457, N455);
and AND2 (N458, N453, N168);
nor NOR2 (N459, N450, N3);
nor NOR3 (N460, N459, N329, N231);
not NOT1 (N461, N456);
xor XOR2 (N462, N457, N343);
nand NAND4 (N463, N414, N186, N17, N230);
nor NOR3 (N464, N462, N400, N145);
nor NOR3 (N465, N446, N311, N319);
and AND4 (N466, N441, N325, N2, N212);
nor NOR2 (N467, N465, N177);
xor XOR2 (N468, N458, N156);
buf BUF1 (N469, N468);
or OR3 (N470, N467, N373, N100);
nor NOR3 (N471, N454, N66, N258);
not NOT1 (N472, N461);
buf BUF1 (N473, N471);
nor NOR4 (N474, N444, N99, N374, N419);
buf BUF1 (N475, N466);
and AND2 (N476, N472, N351);
and AND2 (N477, N476, N394);
buf BUF1 (N478, N451);
xor XOR2 (N479, N464, N95);
not NOT1 (N480, N473);
buf BUF1 (N481, N479);
xor XOR2 (N482, N477, N264);
not NOT1 (N483, N474);
nor NOR4 (N484, N469, N300, N301, N293);
nor NOR2 (N485, N475, N7);
nor NOR4 (N486, N460, N80, N121, N438);
buf BUF1 (N487, N484);
and AND4 (N488, N483, N465, N125, N29);
not NOT1 (N489, N485);
xor XOR2 (N490, N480, N8);
or OR2 (N491, N463, N167);
nor NOR4 (N492, N481, N76, N319, N154);
nor NOR4 (N493, N478, N380, N179, N149);
nand NAND4 (N494, N482, N473, N54, N37);
not NOT1 (N495, N491);
xor XOR2 (N496, N487, N122);
xor XOR2 (N497, N486, N130);
xor XOR2 (N498, N489, N312);
xor XOR2 (N499, N493, N391);
not NOT1 (N500, N495);
and AND3 (N501, N492, N256, N141);
not NOT1 (N502, N490);
not NOT1 (N503, N488);
nor NOR4 (N504, N499, N83, N458, N328);
xor XOR2 (N505, N502, N257);
and AND3 (N506, N503, N422, N477);
xor XOR2 (N507, N505, N249);
nor NOR4 (N508, N498, N349, N130, N497);
buf BUF1 (N509, N3);
nor NOR2 (N510, N507, N136);
nor NOR4 (N511, N509, N161, N187, N251);
or OR4 (N512, N470, N22, N59, N14);
or OR2 (N513, N508, N244);
and AND3 (N514, N506, N65, N81);
xor XOR2 (N515, N500, N11);
nor NOR2 (N516, N513, N14);
xor XOR2 (N517, N494, N54);
nor NOR2 (N518, N496, N57);
not NOT1 (N519, N504);
not NOT1 (N520, N511);
nor NOR2 (N521, N516, N432);
buf BUF1 (N522, N520);
nor NOR4 (N523, N510, N496, N236, N367);
not NOT1 (N524, N519);
nand NAND4 (N525, N521, N427, N107, N483);
not NOT1 (N526, N515);
or OR3 (N527, N518, N480, N361);
nand NAND3 (N528, N526, N41, N433);
not NOT1 (N529, N514);
not NOT1 (N530, N522);
buf BUF1 (N531, N530);
buf BUF1 (N532, N528);
nand NAND4 (N533, N501, N450, N509, N230);
or OR3 (N534, N531, N374, N384);
nor NOR3 (N535, N517, N493, N423);
buf BUF1 (N536, N523);
buf BUF1 (N537, N525);
and AND4 (N538, N532, N87, N140, N336);
or OR2 (N539, N512, N488);
nand NAND2 (N540, N534, N164);
xor XOR2 (N541, N540, N119);
xor XOR2 (N542, N535, N23);
and AND4 (N543, N537, N501, N327, N366);
nor NOR4 (N544, N538, N463, N352, N104);
nor NOR3 (N545, N529, N166, N440);
nor NOR2 (N546, N536, N337);
and AND2 (N547, N541, N490);
or OR4 (N548, N544, N32, N260, N4);
buf BUF1 (N549, N548);
nor NOR2 (N550, N533, N183);
or OR2 (N551, N545, N280);
nand NAND2 (N552, N551, N167);
or OR3 (N553, N549, N393, N148);
buf BUF1 (N554, N553);
nor NOR2 (N555, N524, N325);
not NOT1 (N556, N554);
nand NAND3 (N557, N550, N509, N427);
or OR3 (N558, N546, N212, N116);
not NOT1 (N559, N555);
and AND4 (N560, N547, N545, N73, N57);
or OR4 (N561, N559, N47, N360, N314);
nor NOR3 (N562, N561, N224, N159);
nand NAND2 (N563, N560, N332);
nor NOR4 (N564, N558, N363, N110, N126);
not NOT1 (N565, N563);
xor XOR2 (N566, N562, N374);
or OR3 (N567, N552, N94, N307);
or OR4 (N568, N557, N422, N235, N44);
not NOT1 (N569, N568);
xor XOR2 (N570, N567, N332);
not NOT1 (N571, N542);
and AND3 (N572, N565, N273, N434);
not NOT1 (N573, N527);
or OR4 (N574, N556, N23, N347, N24);
and AND4 (N575, N572, N328, N35, N471);
not NOT1 (N576, N569);
not NOT1 (N577, N539);
and AND2 (N578, N564, N236);
buf BUF1 (N579, N577);
buf BUF1 (N580, N578);
nor NOR4 (N581, N566, N514, N509, N338);
buf BUF1 (N582, N543);
nor NOR2 (N583, N581, N461);
not NOT1 (N584, N570);
buf BUF1 (N585, N573);
or OR3 (N586, N571, N579, N34);
or OR3 (N587, N539, N26, N537);
nand NAND4 (N588, N576, N578, N121, N67);
xor XOR2 (N589, N584, N59);
xor XOR2 (N590, N589, N284);
not NOT1 (N591, N590);
buf BUF1 (N592, N585);
and AND4 (N593, N592, N577, N188, N92);
xor XOR2 (N594, N583, N533);
xor XOR2 (N595, N574, N154);
and AND3 (N596, N580, N79, N201);
nand NAND2 (N597, N593, N8);
not NOT1 (N598, N587);
or OR3 (N599, N575, N411, N42);
or OR2 (N600, N598, N402);
buf BUF1 (N601, N599);
not NOT1 (N602, N595);
xor XOR2 (N603, N591, N392);
or OR4 (N604, N594, N11, N34, N486);
not NOT1 (N605, N601);
nand NAND3 (N606, N588, N128, N40);
or OR4 (N607, N602, N282, N494, N148);
not NOT1 (N608, N604);
nand NAND2 (N609, N608, N306);
nand NAND4 (N610, N586, N207, N128, N207);
xor XOR2 (N611, N603, N121);
buf BUF1 (N612, N596);
not NOT1 (N613, N597);
nor NOR4 (N614, N600, N213, N588, N175);
buf BUF1 (N615, N605);
and AND3 (N616, N615, N435, N198);
xor XOR2 (N617, N607, N12);
not NOT1 (N618, N614);
or OR3 (N619, N610, N388, N511);
or OR2 (N620, N616, N379);
xor XOR2 (N621, N617, N471);
not NOT1 (N622, N619);
xor XOR2 (N623, N609, N297);
not NOT1 (N624, N623);
xor XOR2 (N625, N620, N518);
xor XOR2 (N626, N612, N449);
not NOT1 (N627, N618);
not NOT1 (N628, N627);
buf BUF1 (N629, N606);
or OR4 (N630, N626, N403, N588, N18);
nor NOR2 (N631, N622, N242);
buf BUF1 (N632, N611);
nand NAND2 (N633, N625, N566);
xor XOR2 (N634, N624, N565);
buf BUF1 (N635, N628);
nand NAND4 (N636, N631, N35, N158, N342);
nor NOR4 (N637, N633, N17, N505, N50);
and AND3 (N638, N630, N159, N634);
and AND2 (N639, N225, N634);
and AND4 (N640, N629, N41, N126, N204);
or OR4 (N641, N637, N566, N111, N301);
not NOT1 (N642, N641);
and AND3 (N643, N635, N621, N207);
or OR3 (N644, N214, N183, N389);
nor NOR2 (N645, N613, N363);
or OR3 (N646, N638, N92, N513);
or OR2 (N647, N632, N564);
nor NOR3 (N648, N640, N182, N28);
nand NAND2 (N649, N643, N259);
buf BUF1 (N650, N648);
xor XOR2 (N651, N639, N533);
and AND3 (N652, N650, N170, N589);
nor NOR4 (N653, N646, N541, N118, N250);
nand NAND3 (N654, N651, N337, N482);
nor NOR3 (N655, N652, N140, N319);
nand NAND4 (N656, N655, N319, N190, N331);
xor XOR2 (N657, N644, N409);
nand NAND3 (N658, N653, N257, N392);
buf BUF1 (N659, N649);
not NOT1 (N660, N656);
not NOT1 (N661, N657);
xor XOR2 (N662, N658, N7);
not NOT1 (N663, N662);
not NOT1 (N664, N642);
not NOT1 (N665, N582);
buf BUF1 (N666, N664);
not NOT1 (N667, N661);
xor XOR2 (N668, N645, N552);
not NOT1 (N669, N659);
not NOT1 (N670, N666);
xor XOR2 (N671, N636, N598);
not NOT1 (N672, N671);
nand NAND3 (N673, N647, N366, N141);
xor XOR2 (N674, N660, N460);
buf BUF1 (N675, N667);
or OR4 (N676, N674, N37, N331, N403);
nand NAND3 (N677, N669, N518, N109);
nand NAND4 (N678, N663, N303, N442, N463);
buf BUF1 (N679, N675);
and AND4 (N680, N678, N322, N588, N634);
nor NOR4 (N681, N670, N463, N10, N416);
nor NOR3 (N682, N672, N216, N429);
not NOT1 (N683, N679);
nor NOR3 (N684, N680, N138, N134);
xor XOR2 (N685, N673, N175);
xor XOR2 (N686, N683, N181);
or OR3 (N687, N686, N237, N282);
nor NOR2 (N688, N681, N545);
not NOT1 (N689, N665);
or OR2 (N690, N682, N202);
buf BUF1 (N691, N688);
nor NOR4 (N692, N691, N552, N63, N601);
and AND4 (N693, N687, N278, N362, N278);
nand NAND3 (N694, N676, N467, N590);
nand NAND4 (N695, N690, N691, N273, N382);
and AND4 (N696, N693, N574, N677, N11);
or OR3 (N697, N562, N104, N60);
or OR3 (N698, N685, N326, N416);
buf BUF1 (N699, N668);
and AND2 (N700, N699, N524);
nand NAND4 (N701, N695, N167, N203, N197);
nand NAND2 (N702, N697, N40);
buf BUF1 (N703, N689);
xor XOR2 (N704, N698, N267);
or OR3 (N705, N684, N633, N632);
buf BUF1 (N706, N704);
and AND4 (N707, N692, N498, N643, N577);
xor XOR2 (N708, N705, N393);
buf BUF1 (N709, N702);
nand NAND2 (N710, N706, N650);
and AND3 (N711, N654, N507, N557);
and AND3 (N712, N696, N517, N92);
or OR4 (N713, N707, N94, N408, N331);
and AND3 (N714, N708, N356, N125);
nor NOR4 (N715, N701, N88, N610, N304);
buf BUF1 (N716, N709);
or OR2 (N717, N715, N692);
nor NOR2 (N718, N694, N311);
nand NAND3 (N719, N700, N50, N586);
nand NAND4 (N720, N713, N655, N658, N387);
not NOT1 (N721, N711);
nor NOR4 (N722, N720, N150, N673, N464);
or OR3 (N723, N716, N300, N51);
xor XOR2 (N724, N714, N715);
nor NOR2 (N725, N719, N163);
or OR2 (N726, N712, N371);
and AND3 (N727, N722, N498, N4);
and AND2 (N728, N718, N290);
and AND2 (N729, N710, N167);
or OR3 (N730, N729, N114, N430);
not NOT1 (N731, N727);
nor NOR3 (N732, N721, N100, N358);
and AND4 (N733, N717, N328, N732, N458);
not NOT1 (N734, N525);
nor NOR4 (N735, N731, N255, N299, N256);
or OR3 (N736, N725, N220, N733);
and AND4 (N737, N437, N385, N656, N461);
nand NAND4 (N738, N735, N711, N147, N596);
buf BUF1 (N739, N724);
xor XOR2 (N740, N737, N543);
buf BUF1 (N741, N703);
and AND3 (N742, N726, N90, N120);
and AND4 (N743, N723, N239, N453, N480);
buf BUF1 (N744, N736);
xor XOR2 (N745, N741, N463);
or OR3 (N746, N728, N212, N670);
buf BUF1 (N747, N739);
nor NOR3 (N748, N734, N66, N72);
not NOT1 (N749, N744);
nand NAND2 (N750, N746, N25);
or OR2 (N751, N748, N304);
nor NOR4 (N752, N738, N440, N465, N378);
and AND3 (N753, N749, N304, N98);
and AND3 (N754, N752, N454, N374);
and AND2 (N755, N747, N279);
buf BUF1 (N756, N750);
or OR4 (N757, N745, N512, N229, N675);
buf BUF1 (N758, N730);
buf BUF1 (N759, N751);
nand NAND2 (N760, N759, N203);
or OR4 (N761, N753, N643, N732, N701);
nor NOR3 (N762, N756, N434, N445);
nor NOR3 (N763, N742, N271, N554);
and AND2 (N764, N754, N640);
and AND3 (N765, N755, N56, N457);
and AND3 (N766, N765, N307, N83);
nor NOR3 (N767, N760, N204, N182);
or OR4 (N768, N757, N513, N342, N387);
xor XOR2 (N769, N761, N217);
nor NOR2 (N770, N740, N505);
and AND3 (N771, N743, N352, N523);
buf BUF1 (N772, N770);
buf BUF1 (N773, N766);
nor NOR4 (N774, N762, N411, N314, N348);
nor NOR3 (N775, N767, N205, N170);
xor XOR2 (N776, N758, N428);
nand NAND4 (N777, N768, N614, N267, N509);
xor XOR2 (N778, N777, N163);
xor XOR2 (N779, N774, N665);
nor NOR2 (N780, N779, N243);
not NOT1 (N781, N778);
buf BUF1 (N782, N775);
xor XOR2 (N783, N763, N716);
not NOT1 (N784, N782);
nor NOR4 (N785, N773, N555, N458, N330);
nand NAND2 (N786, N781, N62);
xor XOR2 (N787, N780, N661);
nor NOR4 (N788, N769, N301, N117, N23);
xor XOR2 (N789, N764, N647);
not NOT1 (N790, N785);
or OR4 (N791, N789, N653, N748, N339);
or OR2 (N792, N783, N632);
nand NAND4 (N793, N792, N499, N643, N131);
or OR4 (N794, N784, N620, N596, N133);
and AND2 (N795, N788, N711);
or OR2 (N796, N787, N333);
xor XOR2 (N797, N791, N652);
or OR3 (N798, N786, N83, N79);
nor NOR3 (N799, N797, N602, N175);
nand NAND3 (N800, N798, N433, N317);
not NOT1 (N801, N776);
not NOT1 (N802, N795);
or OR3 (N803, N794, N253, N593);
or OR3 (N804, N772, N294, N356);
xor XOR2 (N805, N799, N779);
not NOT1 (N806, N804);
and AND2 (N807, N796, N448);
not NOT1 (N808, N790);
xor XOR2 (N809, N793, N183);
nor NOR4 (N810, N771, N284, N497, N695);
xor XOR2 (N811, N801, N468);
nand NAND3 (N812, N802, N790, N493);
xor XOR2 (N813, N810, N438);
not NOT1 (N814, N807);
not NOT1 (N815, N814);
or OR2 (N816, N812, N347);
or OR4 (N817, N813, N93, N145, N401);
buf BUF1 (N818, N815);
and AND4 (N819, N818, N742, N146, N347);
xor XOR2 (N820, N808, N240);
buf BUF1 (N821, N806);
xor XOR2 (N822, N820, N300);
or OR3 (N823, N819, N466, N231);
xor XOR2 (N824, N822, N88);
xor XOR2 (N825, N821, N21);
and AND3 (N826, N816, N480, N796);
buf BUF1 (N827, N805);
nand NAND2 (N828, N811, N385);
nand NAND4 (N829, N824, N178, N382, N40);
xor XOR2 (N830, N817, N269);
buf BUF1 (N831, N826);
or OR2 (N832, N828, N692);
and AND4 (N833, N829, N765, N585, N250);
buf BUF1 (N834, N809);
xor XOR2 (N835, N830, N197);
and AND2 (N836, N800, N642);
nor NOR2 (N837, N831, N604);
nand NAND3 (N838, N833, N362, N666);
nor NOR2 (N839, N827, N803);
nor NOR4 (N840, N621, N276, N463, N753);
nor NOR3 (N841, N837, N407, N664);
or OR2 (N842, N841, N723);
or OR3 (N843, N825, N87, N836);
nor NOR3 (N844, N840, N587, N290);
buf BUF1 (N845, N725);
xor XOR2 (N846, N844, N164);
buf BUF1 (N847, N834);
buf BUF1 (N848, N823);
and AND3 (N849, N845, N203, N552);
buf BUF1 (N850, N832);
not NOT1 (N851, N850);
buf BUF1 (N852, N848);
not NOT1 (N853, N839);
xor XOR2 (N854, N842, N125);
not NOT1 (N855, N835);
and AND2 (N856, N849, N613);
and AND2 (N857, N854, N46);
buf BUF1 (N858, N838);
not NOT1 (N859, N858);
and AND2 (N860, N843, N285);
xor XOR2 (N861, N856, N717);
buf BUF1 (N862, N859);
buf BUF1 (N863, N860);
xor XOR2 (N864, N846, N265);
nand NAND3 (N865, N861, N757, N474);
nor NOR3 (N866, N855, N592, N283);
buf BUF1 (N867, N853);
nand NAND4 (N868, N851, N186, N518, N268);
nand NAND3 (N869, N866, N418, N406);
not NOT1 (N870, N862);
not NOT1 (N871, N852);
or OR3 (N872, N867, N614, N384);
nor NOR2 (N873, N864, N50);
xor XOR2 (N874, N872, N799);
nand NAND2 (N875, N869, N629);
xor XOR2 (N876, N847, N846);
buf BUF1 (N877, N875);
and AND2 (N878, N877, N37);
nor NOR3 (N879, N878, N700, N409);
nand NAND4 (N880, N876, N418, N328, N34);
xor XOR2 (N881, N880, N271);
nand NAND2 (N882, N873, N88);
nor NOR2 (N883, N882, N426);
and AND2 (N884, N863, N327);
xor XOR2 (N885, N865, N758);
and AND4 (N886, N883, N620, N122, N388);
nor NOR3 (N887, N871, N846, N822);
or OR2 (N888, N879, N506);
xor XOR2 (N889, N888, N467);
or OR3 (N890, N881, N95, N377);
and AND2 (N891, N885, N600);
xor XOR2 (N892, N857, N1);
buf BUF1 (N893, N884);
nand NAND4 (N894, N887, N444, N246, N442);
xor XOR2 (N895, N890, N855);
xor XOR2 (N896, N889, N45);
and AND3 (N897, N894, N873, N157);
xor XOR2 (N898, N893, N775);
and AND4 (N899, N874, N422, N845, N197);
xor XOR2 (N900, N891, N95);
buf BUF1 (N901, N870);
nand NAND4 (N902, N895, N223, N670, N340);
buf BUF1 (N903, N892);
buf BUF1 (N904, N886);
buf BUF1 (N905, N903);
or OR2 (N906, N901, N492);
buf BUF1 (N907, N904);
or OR3 (N908, N897, N843, N382);
nor NOR4 (N909, N900, N411, N210, N755);
buf BUF1 (N910, N905);
and AND2 (N911, N910, N1);
and AND4 (N912, N898, N446, N582, N178);
nand NAND2 (N913, N907, N122);
nand NAND4 (N914, N911, N568, N734, N434);
xor XOR2 (N915, N902, N227);
xor XOR2 (N916, N912, N428);
not NOT1 (N917, N915);
and AND4 (N918, N908, N830, N43, N124);
nand NAND3 (N919, N896, N813, N520);
and AND2 (N920, N906, N222);
not NOT1 (N921, N918);
nor NOR4 (N922, N917, N102, N8, N31);
not NOT1 (N923, N916);
and AND2 (N924, N920, N420);
nand NAND4 (N925, N919, N153, N90, N182);
nand NAND2 (N926, N925, N870);
buf BUF1 (N927, N922);
nor NOR4 (N928, N927, N861, N449, N617);
buf BUF1 (N929, N923);
nand NAND3 (N930, N913, N178, N516);
and AND4 (N931, N921, N243, N353, N89);
nor NOR2 (N932, N931, N176);
xor XOR2 (N933, N899, N210);
xor XOR2 (N934, N914, N223);
nor NOR3 (N935, N926, N216, N408);
nor NOR4 (N936, N935, N35, N434, N258);
buf BUF1 (N937, N928);
not NOT1 (N938, N936);
or OR3 (N939, N924, N444, N186);
xor XOR2 (N940, N929, N692);
or OR4 (N941, N909, N320, N172, N201);
nor NOR3 (N942, N939, N436, N535);
nand NAND2 (N943, N940, N33);
buf BUF1 (N944, N868);
not NOT1 (N945, N937);
not NOT1 (N946, N932);
buf BUF1 (N947, N945);
buf BUF1 (N948, N930);
and AND3 (N949, N946, N503, N538);
and AND4 (N950, N944, N102, N746, N321);
or OR3 (N951, N938, N774, N277);
and AND2 (N952, N949, N44);
not NOT1 (N953, N941);
xor XOR2 (N954, N933, N458);
nand NAND4 (N955, N950, N101, N906, N321);
nand NAND3 (N956, N954, N668, N907);
and AND2 (N957, N953, N445);
nor NOR2 (N958, N951, N596);
nand NAND4 (N959, N956, N886, N282, N244);
xor XOR2 (N960, N959, N766);
or OR4 (N961, N942, N435, N402, N683);
xor XOR2 (N962, N948, N225);
and AND2 (N963, N962, N368);
xor XOR2 (N964, N943, N669);
not NOT1 (N965, N964);
or OR4 (N966, N934, N230, N349, N542);
buf BUF1 (N967, N961);
xor XOR2 (N968, N952, N357);
nand NAND4 (N969, N958, N604, N947, N755);
nor NOR2 (N970, N893, N854);
not NOT1 (N971, N957);
and AND4 (N972, N970, N459, N553, N630);
or OR4 (N973, N966, N770, N517, N708);
or OR2 (N974, N963, N430);
buf BUF1 (N975, N965);
buf BUF1 (N976, N973);
not NOT1 (N977, N955);
or OR3 (N978, N977, N719, N450);
and AND2 (N979, N974, N490);
not NOT1 (N980, N967);
xor XOR2 (N981, N975, N688);
and AND2 (N982, N978, N871);
and AND2 (N983, N976, N899);
and AND4 (N984, N983, N338, N808, N36);
nor NOR3 (N985, N982, N167, N392);
not NOT1 (N986, N971);
buf BUF1 (N987, N986);
or OR4 (N988, N969, N280, N328, N186);
nor NOR3 (N989, N984, N410, N44);
xor XOR2 (N990, N988, N459);
and AND2 (N991, N972, N23);
or OR3 (N992, N989, N962, N579);
not NOT1 (N993, N992);
nor NOR2 (N994, N990, N17);
and AND3 (N995, N993, N918, N458);
xor XOR2 (N996, N995, N828);
not NOT1 (N997, N994);
not NOT1 (N998, N968);
and AND4 (N999, N991, N396, N888, N358);
and AND4 (N1000, N998, N115, N955, N869);
nand NAND4 (N1001, N979, N721, N531, N534);
nor NOR2 (N1002, N1000, N42);
nor NOR2 (N1003, N1002, N154);
not NOT1 (N1004, N1003);
not NOT1 (N1005, N999);
or OR4 (N1006, N1005, N958, N767, N455);
xor XOR2 (N1007, N985, N979);
not NOT1 (N1008, N981);
nor NOR4 (N1009, N996, N322, N244, N198);
and AND2 (N1010, N1007, N693);
buf BUF1 (N1011, N1006);
xor XOR2 (N1012, N1001, N173);
and AND2 (N1013, N960, N504);
buf BUF1 (N1014, N1009);
buf BUF1 (N1015, N1008);
nand NAND3 (N1016, N997, N103, N242);
xor XOR2 (N1017, N980, N99);
and AND2 (N1018, N1014, N757);
nor NOR2 (N1019, N1010, N935);
or OR4 (N1020, N1004, N200, N667, N776);
xor XOR2 (N1021, N987, N936);
and AND3 (N1022, N1013, N506, N532);
nand NAND2 (N1023, N1022, N825);
not NOT1 (N1024, N1020);
nor NOR3 (N1025, N1023, N469, N622);
or OR3 (N1026, N1016, N917, N433);
nand NAND4 (N1027, N1019, N835, N243, N887);
buf BUF1 (N1028, N1021);
nor NOR2 (N1029, N1011, N780);
or OR4 (N1030, N1017, N309, N261, N1002);
nor NOR3 (N1031, N1012, N656, N967);
not NOT1 (N1032, N1025);
or OR4 (N1033, N1031, N942, N287, N988);
and AND2 (N1034, N1028, N514);
xor XOR2 (N1035, N1032, N341);
buf BUF1 (N1036, N1015);
not NOT1 (N1037, N1018);
nand NAND3 (N1038, N1036, N33, N817);
or OR3 (N1039, N1029, N777, N881);
not NOT1 (N1040, N1027);
nand NAND2 (N1041, N1039, N732);
not NOT1 (N1042, N1034);
buf BUF1 (N1043, N1038);
not NOT1 (N1044, N1037);
xor XOR2 (N1045, N1040, N159);
and AND2 (N1046, N1043, N646);
not NOT1 (N1047, N1042);
and AND4 (N1048, N1044, N812, N338, N986);
nand NAND2 (N1049, N1048, N1012);
xor XOR2 (N1050, N1033, N623);
nor NOR3 (N1051, N1049, N44, N945);
or OR2 (N1052, N1050, N425);
or OR4 (N1053, N1051, N513, N704, N639);
not NOT1 (N1054, N1035);
nor NOR3 (N1055, N1053, N283, N999);
not NOT1 (N1056, N1055);
buf BUF1 (N1057, N1045);
xor XOR2 (N1058, N1052, N946);
buf BUF1 (N1059, N1026);
xor XOR2 (N1060, N1030, N876);
not NOT1 (N1061, N1047);
and AND2 (N1062, N1061, N474);
and AND3 (N1063, N1041, N557, N461);
or OR4 (N1064, N1060, N318, N698, N292);
or OR2 (N1065, N1058, N259);
xor XOR2 (N1066, N1059, N815);
not NOT1 (N1067, N1057);
and AND4 (N1068, N1063, N264, N793, N825);
and AND3 (N1069, N1046, N963, N58);
not NOT1 (N1070, N1062);
not NOT1 (N1071, N1064);
nand NAND3 (N1072, N1065, N982, N376);
nor NOR4 (N1073, N1024, N619, N946, N221);
buf BUF1 (N1074, N1054);
not NOT1 (N1075, N1071);
and AND3 (N1076, N1074, N434, N224);
not NOT1 (N1077, N1069);
not NOT1 (N1078, N1067);
not NOT1 (N1079, N1070);
nor NOR2 (N1080, N1066, N28);
nand NAND4 (N1081, N1080, N223, N873, N988);
or OR3 (N1082, N1068, N534, N860);
buf BUF1 (N1083, N1073);
or OR3 (N1084, N1079, N522, N156);
and AND3 (N1085, N1084, N446, N1043);
and AND3 (N1086, N1076, N215, N910);
buf BUF1 (N1087, N1085);
xor XOR2 (N1088, N1077, N870);
nand NAND3 (N1089, N1087, N319, N392);
xor XOR2 (N1090, N1078, N143);
buf BUF1 (N1091, N1082);
nand NAND4 (N1092, N1089, N548, N451, N353);
or OR3 (N1093, N1083, N593, N1032);
buf BUF1 (N1094, N1075);
nand NAND3 (N1095, N1056, N264, N758);
xor XOR2 (N1096, N1081, N469);
not NOT1 (N1097, N1096);
or OR2 (N1098, N1093, N977);
and AND2 (N1099, N1072, N528);
nand NAND4 (N1100, N1090, N1078, N922, N391);
xor XOR2 (N1101, N1092, N671);
and AND2 (N1102, N1088, N780);
buf BUF1 (N1103, N1102);
buf BUF1 (N1104, N1094);
nor NOR3 (N1105, N1091, N370, N517);
or OR3 (N1106, N1104, N315, N341);
or OR3 (N1107, N1099, N506, N1054);
buf BUF1 (N1108, N1097);
xor XOR2 (N1109, N1108, N162);
nor NOR4 (N1110, N1103, N351, N157, N686);
not NOT1 (N1111, N1100);
not NOT1 (N1112, N1106);
nor NOR2 (N1113, N1112, N349);
nand NAND3 (N1114, N1105, N206, N301);
xor XOR2 (N1115, N1107, N804);
not NOT1 (N1116, N1113);
and AND4 (N1117, N1095, N832, N607, N568);
not NOT1 (N1118, N1116);
nand NAND3 (N1119, N1111, N681, N642);
buf BUF1 (N1120, N1114);
nand NAND4 (N1121, N1117, N791, N977, N766);
xor XOR2 (N1122, N1121, N951);
nand NAND2 (N1123, N1101, N320);
and AND2 (N1124, N1086, N588);
not NOT1 (N1125, N1110);
buf BUF1 (N1126, N1109);
nand NAND4 (N1127, N1115, N702, N590, N1024);
not NOT1 (N1128, N1098);
not NOT1 (N1129, N1127);
or OR3 (N1130, N1118, N606, N417);
buf BUF1 (N1131, N1120);
xor XOR2 (N1132, N1125, N644);
not NOT1 (N1133, N1129);
and AND3 (N1134, N1128, N995, N513);
xor XOR2 (N1135, N1123, N138);
buf BUF1 (N1136, N1130);
not NOT1 (N1137, N1124);
nand NAND2 (N1138, N1137, N454);
buf BUF1 (N1139, N1134);
or OR3 (N1140, N1122, N236, N659);
nor NOR2 (N1141, N1132, N876);
buf BUF1 (N1142, N1133);
not NOT1 (N1143, N1142);
xor XOR2 (N1144, N1126, N101);
not NOT1 (N1145, N1131);
nor NOR4 (N1146, N1138, N122, N470, N638);
nand NAND2 (N1147, N1139, N1048);
not NOT1 (N1148, N1119);
nor NOR3 (N1149, N1146, N1033, N413);
not NOT1 (N1150, N1149);
xor XOR2 (N1151, N1143, N966);
and AND4 (N1152, N1144, N102, N251, N369);
xor XOR2 (N1153, N1135, N815);
xor XOR2 (N1154, N1145, N134);
nand NAND4 (N1155, N1141, N73, N35, N884);
nand NAND3 (N1156, N1140, N1016, N410);
nor NOR4 (N1157, N1153, N873, N660, N189);
buf BUF1 (N1158, N1136);
buf BUF1 (N1159, N1152);
buf BUF1 (N1160, N1155);
or OR3 (N1161, N1147, N522, N935);
and AND4 (N1162, N1148, N1034, N342, N556);
xor XOR2 (N1163, N1154, N486);
and AND3 (N1164, N1157, N273, N561);
not NOT1 (N1165, N1158);
or OR3 (N1166, N1159, N245, N705);
nand NAND3 (N1167, N1150, N200, N816);
nor NOR3 (N1168, N1156, N278, N600);
and AND3 (N1169, N1151, N311, N708);
not NOT1 (N1170, N1162);
or OR3 (N1171, N1161, N759, N766);
not NOT1 (N1172, N1171);
nor NOR4 (N1173, N1169, N660, N462, N782);
buf BUF1 (N1174, N1166);
and AND4 (N1175, N1160, N592, N637, N147);
xor XOR2 (N1176, N1168, N561);
and AND4 (N1177, N1172, N188, N179, N1134);
or OR4 (N1178, N1177, N31, N183, N783);
nand NAND3 (N1179, N1165, N887, N404);
xor XOR2 (N1180, N1173, N928);
buf BUF1 (N1181, N1163);
buf BUF1 (N1182, N1174);
and AND3 (N1183, N1182, N338, N19);
or OR2 (N1184, N1176, N290);
nor NOR2 (N1185, N1183, N902);
xor XOR2 (N1186, N1167, N77);
xor XOR2 (N1187, N1175, N327);
nor NOR4 (N1188, N1185, N317, N42, N422);
and AND4 (N1189, N1180, N995, N1036, N712);
nor NOR4 (N1190, N1178, N870, N723, N838);
or OR3 (N1191, N1190, N970, N573);
and AND2 (N1192, N1188, N571);
nor NOR2 (N1193, N1186, N901);
or OR3 (N1194, N1192, N699, N1059);
buf BUF1 (N1195, N1179);
buf BUF1 (N1196, N1170);
buf BUF1 (N1197, N1191);
not NOT1 (N1198, N1189);
buf BUF1 (N1199, N1194);
not NOT1 (N1200, N1193);
nand NAND4 (N1201, N1199, N246, N935, N556);
nand NAND2 (N1202, N1198, N413);
xor XOR2 (N1203, N1201, N69);
and AND4 (N1204, N1164, N752, N654, N1035);
not NOT1 (N1205, N1202);
and AND3 (N1206, N1187, N584, N635);
nand NAND2 (N1207, N1204, N500);
xor XOR2 (N1208, N1206, N617);
buf BUF1 (N1209, N1181);
buf BUF1 (N1210, N1196);
and AND3 (N1211, N1210, N1031, N883);
nand NAND3 (N1212, N1205, N891, N856);
not NOT1 (N1213, N1195);
or OR3 (N1214, N1184, N862, N534);
and AND2 (N1215, N1212, N977);
buf BUF1 (N1216, N1209);
nor NOR3 (N1217, N1216, N461, N82);
nor NOR3 (N1218, N1213, N191, N486);
nand NAND3 (N1219, N1211, N370, N663);
buf BUF1 (N1220, N1208);
nor NOR2 (N1221, N1215, N726);
and AND3 (N1222, N1219, N74, N1027);
nand NAND4 (N1223, N1218, N555, N423, N603);
nand NAND2 (N1224, N1221, N471);
or OR3 (N1225, N1214, N471, N1007);
not NOT1 (N1226, N1224);
buf BUF1 (N1227, N1223);
or OR3 (N1228, N1207, N1058, N231);
or OR3 (N1229, N1217, N216, N873);
xor XOR2 (N1230, N1226, N631);
nor NOR4 (N1231, N1225, N251, N389, N1198);
or OR2 (N1232, N1228, N625);
buf BUF1 (N1233, N1232);
xor XOR2 (N1234, N1229, N366);
or OR4 (N1235, N1203, N927, N800, N1169);
or OR2 (N1236, N1233, N698);
nor NOR2 (N1237, N1235, N1118);
and AND3 (N1238, N1236, N1107, N28);
buf BUF1 (N1239, N1200);
and AND2 (N1240, N1230, N1064);
not NOT1 (N1241, N1239);
and AND2 (N1242, N1220, N150);
not NOT1 (N1243, N1227);
buf BUF1 (N1244, N1231);
or OR2 (N1245, N1237, N74);
and AND4 (N1246, N1242, N947, N28, N799);
nor NOR4 (N1247, N1246, N753, N857, N1241);
nand NAND2 (N1248, N565, N557);
and AND2 (N1249, N1222, N583);
xor XOR2 (N1250, N1244, N350);
and AND3 (N1251, N1248, N726, N9);
nor NOR2 (N1252, N1238, N845);
nor NOR3 (N1253, N1252, N607, N140);
buf BUF1 (N1254, N1247);
and AND2 (N1255, N1254, N388);
and AND4 (N1256, N1250, N298, N702, N970);
and AND2 (N1257, N1197, N767);
not NOT1 (N1258, N1249);
xor XOR2 (N1259, N1234, N643);
not NOT1 (N1260, N1245);
and AND3 (N1261, N1255, N269, N248);
or OR3 (N1262, N1240, N1115, N1218);
not NOT1 (N1263, N1258);
buf BUF1 (N1264, N1262);
not NOT1 (N1265, N1257);
nor NOR3 (N1266, N1256, N458, N497);
or OR3 (N1267, N1243, N472, N992);
nand NAND3 (N1268, N1266, N180, N1158);
xor XOR2 (N1269, N1259, N941);
nand NAND3 (N1270, N1253, N533, N107);
and AND2 (N1271, N1267, N690);
or OR4 (N1272, N1264, N171, N50, N774);
not NOT1 (N1273, N1265);
not NOT1 (N1274, N1261);
and AND4 (N1275, N1270, N1080, N251, N1090);
nand NAND4 (N1276, N1271, N470, N102, N347);
not NOT1 (N1277, N1274);
and AND4 (N1278, N1251, N731, N71, N225);
not NOT1 (N1279, N1272);
not NOT1 (N1280, N1273);
xor XOR2 (N1281, N1278, N244);
and AND4 (N1282, N1268, N132, N110, N364);
nor NOR3 (N1283, N1277, N973, N550);
buf BUF1 (N1284, N1280);
buf BUF1 (N1285, N1269);
xor XOR2 (N1286, N1285, N1208);
xor XOR2 (N1287, N1276, N263);
not NOT1 (N1288, N1284);
and AND3 (N1289, N1263, N1118, N728);
nor NOR2 (N1290, N1288, N957);
buf BUF1 (N1291, N1283);
nor NOR2 (N1292, N1291, N737);
buf BUF1 (N1293, N1292);
xor XOR2 (N1294, N1275, N150);
xor XOR2 (N1295, N1281, N739);
or OR4 (N1296, N1295, N230, N872, N208);
nor NOR2 (N1297, N1287, N833);
or OR2 (N1298, N1286, N1147);
not NOT1 (N1299, N1279);
xor XOR2 (N1300, N1296, N357);
nand NAND3 (N1301, N1294, N944, N322);
or OR2 (N1302, N1298, N681);
buf BUF1 (N1303, N1260);
not NOT1 (N1304, N1290);
nor NOR3 (N1305, N1293, N721, N856);
buf BUF1 (N1306, N1303);
and AND2 (N1307, N1301, N103);
buf BUF1 (N1308, N1297);
buf BUF1 (N1309, N1289);
or OR2 (N1310, N1282, N178);
or OR4 (N1311, N1307, N1218, N246, N602);
xor XOR2 (N1312, N1306, N1182);
or OR4 (N1313, N1299, N1027, N576, N270);
nand NAND3 (N1314, N1304, N911, N674);
nand NAND2 (N1315, N1305, N615);
xor XOR2 (N1316, N1302, N138);
nor NOR2 (N1317, N1316, N298);
or OR3 (N1318, N1300, N1064, N235);
xor XOR2 (N1319, N1317, N955);
or OR3 (N1320, N1314, N1166, N542);
buf BUF1 (N1321, N1310);
nor NOR4 (N1322, N1308, N979, N858, N934);
xor XOR2 (N1323, N1315, N349);
not NOT1 (N1324, N1319);
xor XOR2 (N1325, N1312, N767);
xor XOR2 (N1326, N1318, N116);
nand NAND4 (N1327, N1323, N651, N134, N526);
not NOT1 (N1328, N1326);
not NOT1 (N1329, N1309);
nand NAND4 (N1330, N1311, N1214, N1014, N58);
not NOT1 (N1331, N1322);
or OR4 (N1332, N1313, N1184, N403, N539);
not NOT1 (N1333, N1328);
buf BUF1 (N1334, N1321);
nand NAND4 (N1335, N1334, N337, N135, N472);
buf BUF1 (N1336, N1332);
or OR3 (N1337, N1325, N316, N1291);
buf BUF1 (N1338, N1327);
or OR2 (N1339, N1329, N1078);
buf BUF1 (N1340, N1337);
or OR2 (N1341, N1339, N1013);
nor NOR4 (N1342, N1333, N1138, N1083, N61);
not NOT1 (N1343, N1338);
and AND2 (N1344, N1343, N483);
xor XOR2 (N1345, N1336, N594);
or OR2 (N1346, N1342, N323);
buf BUF1 (N1347, N1345);
not NOT1 (N1348, N1344);
or OR4 (N1349, N1324, N1234, N922, N21);
nand NAND4 (N1350, N1330, N697, N1182, N394);
buf BUF1 (N1351, N1341);
buf BUF1 (N1352, N1351);
not NOT1 (N1353, N1335);
xor XOR2 (N1354, N1347, N1140);
nor NOR2 (N1355, N1348, N1315);
and AND3 (N1356, N1353, N154, N226);
or OR4 (N1357, N1320, N1086, N528, N55);
or OR4 (N1358, N1354, N1154, N219, N1025);
or OR2 (N1359, N1355, N1058);
nor NOR3 (N1360, N1356, N304, N1256);
buf BUF1 (N1361, N1360);
nor NOR2 (N1362, N1349, N864);
nor NOR4 (N1363, N1362, N385, N420, N716);
xor XOR2 (N1364, N1352, N1184);
nand NAND2 (N1365, N1359, N1038);
or OR3 (N1366, N1331, N1267, N166);
or OR4 (N1367, N1346, N569, N990, N742);
and AND3 (N1368, N1363, N539, N862);
buf BUF1 (N1369, N1364);
not NOT1 (N1370, N1361);
nor NOR4 (N1371, N1366, N311, N1297, N265);
nor NOR3 (N1372, N1367, N779, N671);
not NOT1 (N1373, N1371);
buf BUF1 (N1374, N1358);
or OR3 (N1375, N1372, N558, N1131);
nor NOR3 (N1376, N1369, N342, N69);
nand NAND4 (N1377, N1376, N2, N897, N513);
and AND2 (N1378, N1350, N596);
or OR3 (N1379, N1370, N693, N1012);
and AND2 (N1380, N1357, N76);
nand NAND2 (N1381, N1340, N810);
nor NOR3 (N1382, N1379, N49, N7);
nor NOR2 (N1383, N1378, N1322);
xor XOR2 (N1384, N1375, N834);
and AND4 (N1385, N1374, N1187, N1153, N954);
nor NOR4 (N1386, N1385, N975, N1113, N588);
nor NOR3 (N1387, N1365, N1343, N22);
xor XOR2 (N1388, N1380, N773);
or OR2 (N1389, N1386, N1071);
nor NOR2 (N1390, N1381, N1155);
and AND4 (N1391, N1390, N549, N896, N450);
or OR3 (N1392, N1383, N376, N861);
or OR3 (N1393, N1388, N776, N593);
xor XOR2 (N1394, N1384, N107);
or OR3 (N1395, N1389, N1243, N944);
not NOT1 (N1396, N1393);
or OR3 (N1397, N1391, N839, N1264);
nand NAND3 (N1398, N1377, N925, N486);
nor NOR3 (N1399, N1396, N484, N216);
nand NAND4 (N1400, N1399, N995, N1121, N171);
nor NOR3 (N1401, N1373, N519, N952);
and AND3 (N1402, N1397, N240, N88);
xor XOR2 (N1403, N1392, N642);
nor NOR3 (N1404, N1403, N1350, N847);
nor NOR3 (N1405, N1400, N1312, N999);
not NOT1 (N1406, N1398);
buf BUF1 (N1407, N1394);
not NOT1 (N1408, N1382);
and AND3 (N1409, N1407, N107, N294);
nand NAND4 (N1410, N1404, N512, N795, N1200);
nor NOR3 (N1411, N1395, N603, N568);
buf BUF1 (N1412, N1406);
xor XOR2 (N1413, N1410, N830);
xor XOR2 (N1414, N1409, N1235);
nor NOR2 (N1415, N1414, N516);
buf BUF1 (N1416, N1408);
nor NOR4 (N1417, N1412, N596, N374, N741);
buf BUF1 (N1418, N1368);
not NOT1 (N1419, N1402);
nand NAND3 (N1420, N1415, N128, N1026);
and AND4 (N1421, N1418, N61, N1148, N141);
nand NAND3 (N1422, N1413, N1013, N44);
xor XOR2 (N1423, N1387, N1241);
or OR2 (N1424, N1417, N160);
nor NOR3 (N1425, N1416, N546, N1320);
nand NAND4 (N1426, N1424, N425, N881, N826);
buf BUF1 (N1427, N1425);
or OR3 (N1428, N1427, N831, N585);
nand NAND4 (N1429, N1423, N447, N139, N719);
or OR2 (N1430, N1405, N48);
or OR4 (N1431, N1428, N820, N1022, N174);
nand NAND2 (N1432, N1430, N570);
nor NOR3 (N1433, N1419, N133, N720);
and AND4 (N1434, N1432, N1188, N218, N1123);
not NOT1 (N1435, N1421);
nor NOR2 (N1436, N1434, N238);
nand NAND4 (N1437, N1431, N109, N483, N1076);
xor XOR2 (N1438, N1411, N968);
buf BUF1 (N1439, N1420);
or OR4 (N1440, N1426, N1098, N1375, N939);
and AND4 (N1441, N1437, N557, N761, N768);
xor XOR2 (N1442, N1441, N861);
or OR2 (N1443, N1440, N710);
nand NAND4 (N1444, N1439, N755, N128, N1023);
buf BUF1 (N1445, N1422);
nor NOR3 (N1446, N1429, N1238, N763);
or OR4 (N1447, N1435, N891, N188, N1116);
or OR3 (N1448, N1436, N740, N246);
not NOT1 (N1449, N1448);
nand NAND2 (N1450, N1443, N1309);
or OR2 (N1451, N1442, N597);
xor XOR2 (N1452, N1451, N1075);
buf BUF1 (N1453, N1401);
nand NAND2 (N1454, N1450, N1124);
xor XOR2 (N1455, N1452, N383);
xor XOR2 (N1456, N1446, N1039);
not NOT1 (N1457, N1433);
or OR2 (N1458, N1456, N1187);
buf BUF1 (N1459, N1445);
xor XOR2 (N1460, N1457, N952);
buf BUF1 (N1461, N1459);
buf BUF1 (N1462, N1453);
buf BUF1 (N1463, N1455);
nand NAND2 (N1464, N1460, N1154);
xor XOR2 (N1465, N1462, N1290);
not NOT1 (N1466, N1461);
buf BUF1 (N1467, N1466);
xor XOR2 (N1468, N1438, N526);
nor NOR3 (N1469, N1465, N1184, N207);
not NOT1 (N1470, N1444);
or OR2 (N1471, N1458, N1087);
nor NOR2 (N1472, N1468, N1407);
buf BUF1 (N1473, N1471);
not NOT1 (N1474, N1464);
nor NOR4 (N1475, N1467, N1199, N1281, N1277);
or OR4 (N1476, N1449, N835, N1249, N1128);
not NOT1 (N1477, N1454);
or OR3 (N1478, N1463, N1214, N319);
nand NAND3 (N1479, N1472, N1368, N253);
buf BUF1 (N1480, N1470);
and AND3 (N1481, N1469, N51, N659);
buf BUF1 (N1482, N1480);
not NOT1 (N1483, N1482);
xor XOR2 (N1484, N1476, N1383);
nand NAND4 (N1485, N1447, N382, N1061, N713);
not NOT1 (N1486, N1473);
not NOT1 (N1487, N1484);
buf BUF1 (N1488, N1485);
xor XOR2 (N1489, N1477, N924);
and AND2 (N1490, N1487, N794);
nor NOR3 (N1491, N1489, N350, N189);
not NOT1 (N1492, N1486);
and AND4 (N1493, N1483, N1061, N1075, N1120);
xor XOR2 (N1494, N1475, N101);
and AND3 (N1495, N1494, N785, N53);
or OR4 (N1496, N1478, N1186, N300, N1415);
xor XOR2 (N1497, N1492, N549);
nor NOR4 (N1498, N1474, N183, N950, N187);
nand NAND3 (N1499, N1488, N442, N474);
xor XOR2 (N1500, N1497, N713);
xor XOR2 (N1501, N1495, N1445);
nor NOR3 (N1502, N1493, N1292, N559);
nand NAND4 (N1503, N1479, N263, N104, N577);
or OR3 (N1504, N1498, N847, N136);
nor NOR3 (N1505, N1504, N895, N740);
buf BUF1 (N1506, N1501);
nor NOR3 (N1507, N1481, N491, N602);
not NOT1 (N1508, N1496);
or OR3 (N1509, N1506, N345, N170);
buf BUF1 (N1510, N1502);
or OR4 (N1511, N1507, N1023, N385, N1228);
xor XOR2 (N1512, N1500, N441);
xor XOR2 (N1513, N1511, N404);
or OR2 (N1514, N1508, N1479);
nor NOR3 (N1515, N1505, N1505, N8);
not NOT1 (N1516, N1515);
not NOT1 (N1517, N1510);
nand NAND4 (N1518, N1516, N1280, N798, N445);
or OR3 (N1519, N1513, N1509, N736);
nand NAND3 (N1520, N1007, N388, N1018);
or OR3 (N1521, N1517, N60, N687);
nand NAND4 (N1522, N1499, N384, N48, N1388);
or OR4 (N1523, N1514, N361, N605, N578);
nor NOR4 (N1524, N1523, N397, N1255, N1398);
nand NAND2 (N1525, N1490, N892);
nand NAND2 (N1526, N1520, N1312);
and AND2 (N1527, N1525, N461);
nand NAND2 (N1528, N1521, N65);
buf BUF1 (N1529, N1503);
or OR3 (N1530, N1519, N166, N789);
not NOT1 (N1531, N1527);
and AND4 (N1532, N1530, N954, N783, N343);
xor XOR2 (N1533, N1518, N754);
or OR2 (N1534, N1491, N694);
buf BUF1 (N1535, N1512);
or OR4 (N1536, N1529, N1007, N822, N118);
buf BUF1 (N1537, N1524);
and AND2 (N1538, N1526, N1034);
nand NAND4 (N1539, N1537, N797, N168, N1538);
nor NOR3 (N1540, N477, N763, N130);
xor XOR2 (N1541, N1535, N1307);
buf BUF1 (N1542, N1531);
nor NOR2 (N1543, N1541, N1526);
buf BUF1 (N1544, N1542);
not NOT1 (N1545, N1533);
and AND3 (N1546, N1540, N1039, N835);
xor XOR2 (N1547, N1522, N1430);
or OR2 (N1548, N1539, N647);
xor XOR2 (N1549, N1546, N1526);
or OR4 (N1550, N1549, N413, N293, N1066);
or OR2 (N1551, N1528, N1115);
not NOT1 (N1552, N1547);
xor XOR2 (N1553, N1544, N571);
and AND4 (N1554, N1532, N947, N596, N1539);
buf BUF1 (N1555, N1552);
nand NAND4 (N1556, N1545, N1455, N324, N2);
and AND4 (N1557, N1543, N774, N107, N1107);
and AND4 (N1558, N1534, N1272, N364, N1361);
or OR2 (N1559, N1551, N589);
and AND2 (N1560, N1550, N1003);
nor NOR3 (N1561, N1548, N217, N315);
nand NAND2 (N1562, N1559, N1289);
buf BUF1 (N1563, N1557);
or OR4 (N1564, N1553, N1058, N683, N1330);
buf BUF1 (N1565, N1554);
and AND2 (N1566, N1555, N37);
or OR3 (N1567, N1561, N1152, N176);
buf BUF1 (N1568, N1565);
and AND3 (N1569, N1562, N1100, N1397);
and AND4 (N1570, N1566, N747, N1307, N294);
not NOT1 (N1571, N1558);
buf BUF1 (N1572, N1560);
xor XOR2 (N1573, N1572, N604);
nand NAND3 (N1574, N1568, N520, N567);
or OR2 (N1575, N1569, N526);
xor XOR2 (N1576, N1570, N785);
buf BUF1 (N1577, N1567);
nand NAND3 (N1578, N1563, N1021, N1416);
nand NAND3 (N1579, N1556, N1316, N170);
nand NAND4 (N1580, N1577, N1548, N309, N1459);
nor NOR4 (N1581, N1579, N857, N600, N899);
buf BUF1 (N1582, N1574);
not NOT1 (N1583, N1571);
buf BUF1 (N1584, N1573);
xor XOR2 (N1585, N1584, N1123);
xor XOR2 (N1586, N1582, N318);
or OR4 (N1587, N1536, N983, N14, N166);
not NOT1 (N1588, N1564);
not NOT1 (N1589, N1587);
xor XOR2 (N1590, N1588, N568);
and AND2 (N1591, N1575, N215);
xor XOR2 (N1592, N1578, N8);
xor XOR2 (N1593, N1586, N1411);
and AND4 (N1594, N1581, N1448, N357, N493);
and AND4 (N1595, N1594, N1089, N871, N547);
xor XOR2 (N1596, N1590, N347);
xor XOR2 (N1597, N1580, N981);
buf BUF1 (N1598, N1597);
and AND4 (N1599, N1595, N646, N1158, N17);
not NOT1 (N1600, N1589);
xor XOR2 (N1601, N1592, N1008);
or OR2 (N1602, N1601, N1340);
buf BUF1 (N1603, N1583);
nor NOR3 (N1604, N1596, N1432, N1064);
buf BUF1 (N1605, N1598);
nand NAND4 (N1606, N1591, N920, N906, N745);
buf BUF1 (N1607, N1605);
xor XOR2 (N1608, N1593, N379);
or OR2 (N1609, N1606, N974);
xor XOR2 (N1610, N1603, N1345);
and AND2 (N1611, N1609, N644);
not NOT1 (N1612, N1608);
buf BUF1 (N1613, N1600);
nor NOR3 (N1614, N1585, N1407, N134);
and AND3 (N1615, N1612, N1400, N527);
xor XOR2 (N1616, N1602, N128);
nand NAND4 (N1617, N1607, N800, N865, N1032);
buf BUF1 (N1618, N1613);
or OR4 (N1619, N1599, N797, N260, N1543);
or OR2 (N1620, N1615, N1276);
buf BUF1 (N1621, N1576);
and AND2 (N1622, N1611, N660);
nor NOR3 (N1623, N1610, N1295, N342);
nand NAND4 (N1624, N1617, N106, N1037, N335);
nor NOR3 (N1625, N1616, N67, N903);
buf BUF1 (N1626, N1622);
or OR3 (N1627, N1621, N1260, N1341);
nand NAND2 (N1628, N1614, N307);
nand NAND2 (N1629, N1619, N756);
or OR2 (N1630, N1624, N304);
buf BUF1 (N1631, N1626);
or OR2 (N1632, N1618, N253);
buf BUF1 (N1633, N1632);
and AND4 (N1634, N1628, N207, N1279, N636);
nor NOR4 (N1635, N1620, N724, N859, N1094);
and AND3 (N1636, N1604, N887, N488);
not NOT1 (N1637, N1631);
and AND4 (N1638, N1633, N500, N556, N733);
xor XOR2 (N1639, N1629, N1101);
and AND2 (N1640, N1625, N1497);
xor XOR2 (N1641, N1637, N866);
or OR4 (N1642, N1627, N832, N136, N1263);
and AND2 (N1643, N1638, N1467);
not NOT1 (N1644, N1630);
or OR2 (N1645, N1636, N1634);
not NOT1 (N1646, N1609);
xor XOR2 (N1647, N1623, N532);
xor XOR2 (N1648, N1644, N558);
xor XOR2 (N1649, N1647, N1558);
buf BUF1 (N1650, N1649);
not NOT1 (N1651, N1643);
buf BUF1 (N1652, N1650);
not NOT1 (N1653, N1639);
buf BUF1 (N1654, N1652);
nor NOR2 (N1655, N1645, N1473);
nor NOR2 (N1656, N1653, N138);
buf BUF1 (N1657, N1654);
nand NAND4 (N1658, N1656, N160, N115, N922);
nand NAND4 (N1659, N1648, N1591, N979, N767);
and AND3 (N1660, N1646, N1492, N1532);
xor XOR2 (N1661, N1651, N21);
or OR3 (N1662, N1658, N1192, N170);
buf BUF1 (N1663, N1655);
nand NAND2 (N1664, N1635, N968);
or OR4 (N1665, N1662, N1594, N48, N1638);
buf BUF1 (N1666, N1641);
not NOT1 (N1667, N1665);
nand NAND2 (N1668, N1657, N1158);
nor NOR3 (N1669, N1659, N364, N379);
not NOT1 (N1670, N1666);
nor NOR2 (N1671, N1661, N487);
not NOT1 (N1672, N1640);
not NOT1 (N1673, N1668);
nand NAND2 (N1674, N1660, N417);
xor XOR2 (N1675, N1642, N449);
nand NAND3 (N1676, N1672, N185, N1445);
and AND2 (N1677, N1669, N1025);
not NOT1 (N1678, N1677);
nor NOR4 (N1679, N1678, N299, N668, N657);
nand NAND4 (N1680, N1675, N1401, N214, N1251);
or OR4 (N1681, N1670, N409, N1209, N1523);
not NOT1 (N1682, N1680);
xor XOR2 (N1683, N1664, N1044);
xor XOR2 (N1684, N1667, N1260);
and AND4 (N1685, N1679, N473, N929, N1626);
buf BUF1 (N1686, N1683);
buf BUF1 (N1687, N1684);
and AND4 (N1688, N1686, N34, N187, N1052);
or OR2 (N1689, N1663, N1674);
nor NOR2 (N1690, N209, N637);
xor XOR2 (N1691, N1681, N1226);
xor XOR2 (N1692, N1688, N313);
nor NOR4 (N1693, N1673, N1672, N1564, N1156);
or OR2 (N1694, N1676, N1593);
xor XOR2 (N1695, N1689, N971);
not NOT1 (N1696, N1695);
xor XOR2 (N1697, N1692, N1395);
nor NOR4 (N1698, N1697, N1020, N732, N1495);
not NOT1 (N1699, N1685);
not NOT1 (N1700, N1694);
nor NOR3 (N1701, N1696, N1367, N754);
buf BUF1 (N1702, N1691);
nor NOR2 (N1703, N1699, N1344);
nand NAND2 (N1704, N1687, N1306);
buf BUF1 (N1705, N1671);
xor XOR2 (N1706, N1690, N420);
nand NAND2 (N1707, N1706, N501);
and AND2 (N1708, N1701, N416);
or OR2 (N1709, N1708, N1289);
or OR4 (N1710, N1707, N977, N1217, N1619);
not NOT1 (N1711, N1700);
buf BUF1 (N1712, N1704);
not NOT1 (N1713, N1703);
not NOT1 (N1714, N1682);
xor XOR2 (N1715, N1713, N1622);
not NOT1 (N1716, N1712);
and AND2 (N1717, N1715, N617);
or OR3 (N1718, N1705, N1479, N682);
nor NOR3 (N1719, N1698, N161, N1681);
or OR4 (N1720, N1711, N1115, N1690, N648);
or OR4 (N1721, N1710, N130, N1184, N353);
xor XOR2 (N1722, N1702, N1229);
or OR3 (N1723, N1709, N584, N1382);
nand NAND2 (N1724, N1717, N1094);
and AND4 (N1725, N1723, N1712, N1156, N606);
nand NAND4 (N1726, N1693, N1612, N1286, N9);
or OR4 (N1727, N1720, N448, N1059, N837);
nand NAND3 (N1728, N1719, N1212, N497);
nand NAND3 (N1729, N1725, N353, N1420);
and AND4 (N1730, N1718, N419, N1125, N519);
or OR3 (N1731, N1721, N367, N721);
buf BUF1 (N1732, N1724);
nor NOR2 (N1733, N1714, N73);
or OR3 (N1734, N1722, N265, N383);
not NOT1 (N1735, N1734);
nor NOR2 (N1736, N1733, N1115);
xor XOR2 (N1737, N1732, N1641);
and AND3 (N1738, N1735, N1188, N923);
nor NOR2 (N1739, N1727, N1564);
or OR3 (N1740, N1729, N1708, N975);
nor NOR3 (N1741, N1737, N1425, N1120);
and AND3 (N1742, N1716, N714, N703);
not NOT1 (N1743, N1738);
nand NAND2 (N1744, N1726, N387);
nor NOR4 (N1745, N1744, N511, N820, N1312);
xor XOR2 (N1746, N1740, N1408);
buf BUF1 (N1747, N1736);
or OR2 (N1748, N1742, N1487);
buf BUF1 (N1749, N1745);
and AND3 (N1750, N1748, N41, N1155);
nor NOR2 (N1751, N1743, N1245);
nor NOR2 (N1752, N1747, N1586);
xor XOR2 (N1753, N1739, N286);
buf BUF1 (N1754, N1746);
and AND4 (N1755, N1749, N33, N581, N150);
xor XOR2 (N1756, N1752, N675);
not NOT1 (N1757, N1741);
xor XOR2 (N1758, N1731, N342);
buf BUF1 (N1759, N1754);
not NOT1 (N1760, N1753);
buf BUF1 (N1761, N1730);
nor NOR3 (N1762, N1757, N58, N1418);
xor XOR2 (N1763, N1750, N857);
xor XOR2 (N1764, N1755, N822);
and AND2 (N1765, N1728, N236);
buf BUF1 (N1766, N1758);
buf BUF1 (N1767, N1764);
and AND2 (N1768, N1760, N136);
and AND4 (N1769, N1767, N351, N1268, N634);
not NOT1 (N1770, N1751);
and AND2 (N1771, N1762, N1530);
nand NAND4 (N1772, N1766, N1155, N798, N584);
xor XOR2 (N1773, N1765, N778);
or OR2 (N1774, N1773, N791);
nor NOR2 (N1775, N1756, N973);
not NOT1 (N1776, N1759);
xor XOR2 (N1777, N1768, N1125);
nor NOR3 (N1778, N1777, N1160, N1260);
nand NAND2 (N1779, N1775, N785);
and AND3 (N1780, N1774, N714, N1077);
and AND3 (N1781, N1770, N1598, N1655);
or OR2 (N1782, N1781, N764);
not NOT1 (N1783, N1761);
not NOT1 (N1784, N1778);
or OR4 (N1785, N1779, N270, N751, N1105);
or OR3 (N1786, N1763, N612, N689);
and AND4 (N1787, N1786, N635, N611, N1736);
buf BUF1 (N1788, N1787);
nand NAND4 (N1789, N1782, N654, N985, N871);
not NOT1 (N1790, N1769);
and AND4 (N1791, N1771, N1076, N1545, N1065);
or OR3 (N1792, N1790, N1491, N1502);
buf BUF1 (N1793, N1772);
xor XOR2 (N1794, N1788, N914);
not NOT1 (N1795, N1789);
not NOT1 (N1796, N1793);
nand NAND3 (N1797, N1794, N356, N277);
buf BUF1 (N1798, N1795);
xor XOR2 (N1799, N1792, N21);
xor XOR2 (N1800, N1791, N279);
and AND3 (N1801, N1800, N174, N317);
xor XOR2 (N1802, N1797, N362);
and AND3 (N1803, N1783, N1715, N1057);
xor XOR2 (N1804, N1784, N1342);
nor NOR4 (N1805, N1802, N1275, N753, N261);
buf BUF1 (N1806, N1804);
and AND4 (N1807, N1776, N94, N335, N922);
xor XOR2 (N1808, N1801, N780);
buf BUF1 (N1809, N1803);
or OR4 (N1810, N1808, N162, N195, N1356);
or OR2 (N1811, N1806, N1196);
not NOT1 (N1812, N1798);
and AND3 (N1813, N1811, N1534, N1768);
nor NOR2 (N1814, N1805, N1090);
or OR4 (N1815, N1809, N1380, N651, N1236);
nand NAND4 (N1816, N1796, N179, N850, N84);
or OR3 (N1817, N1812, N911, N884);
buf BUF1 (N1818, N1799);
and AND3 (N1819, N1817, N1158, N1066);
not NOT1 (N1820, N1785);
buf BUF1 (N1821, N1816);
not NOT1 (N1822, N1807);
buf BUF1 (N1823, N1818);
and AND2 (N1824, N1815, N841);
not NOT1 (N1825, N1820);
buf BUF1 (N1826, N1822);
not NOT1 (N1827, N1813);
nor NOR4 (N1828, N1810, N267, N1544, N1177);
buf BUF1 (N1829, N1828);
or OR4 (N1830, N1821, N857, N1316, N979);
not NOT1 (N1831, N1819);
not NOT1 (N1832, N1830);
or OR3 (N1833, N1831, N1418, N543);
xor XOR2 (N1834, N1824, N327);
xor XOR2 (N1835, N1826, N1667);
buf BUF1 (N1836, N1780);
and AND3 (N1837, N1829, N346, N596);
xor XOR2 (N1838, N1832, N1421);
nand NAND3 (N1839, N1835, N1259, N842);
and AND2 (N1840, N1823, N738);
buf BUF1 (N1841, N1837);
not NOT1 (N1842, N1827);
nand NAND3 (N1843, N1825, N399, N378);
xor XOR2 (N1844, N1843, N296);
nor NOR4 (N1845, N1834, N943, N1072, N435);
nand NAND4 (N1846, N1838, N1637, N1446, N672);
nand NAND2 (N1847, N1839, N4);
xor XOR2 (N1848, N1846, N152);
not NOT1 (N1849, N1841);
nor NOR4 (N1850, N1847, N1707, N176, N358);
nand NAND3 (N1851, N1844, N1847, N1720);
buf BUF1 (N1852, N1850);
nand NAND2 (N1853, N1849, N1425);
xor XOR2 (N1854, N1814, N1385);
xor XOR2 (N1855, N1851, N218);
and AND4 (N1856, N1836, N857, N1418, N646);
nor NOR3 (N1857, N1855, N594, N87);
not NOT1 (N1858, N1840);
and AND4 (N1859, N1857, N1104, N292, N813);
not NOT1 (N1860, N1853);
or OR4 (N1861, N1856, N1133, N1461, N227);
nor NOR2 (N1862, N1854, N1118);
buf BUF1 (N1863, N1833);
nand NAND4 (N1864, N1842, N838, N1451, N1247);
nand NAND2 (N1865, N1863, N1394);
xor XOR2 (N1866, N1862, N1026);
and AND2 (N1867, N1852, N1121);
buf BUF1 (N1868, N1859);
not NOT1 (N1869, N1868);
nand NAND2 (N1870, N1860, N1062);
xor XOR2 (N1871, N1865, N1631);
and AND4 (N1872, N1861, N365, N1856, N327);
or OR2 (N1873, N1845, N441);
nor NOR3 (N1874, N1858, N441, N940);
xor XOR2 (N1875, N1874, N1067);
not NOT1 (N1876, N1871);
nor NOR3 (N1877, N1870, N1744, N1577);
buf BUF1 (N1878, N1877);
xor XOR2 (N1879, N1872, N255);
xor XOR2 (N1880, N1878, N1767);
nor NOR3 (N1881, N1864, N987, N967);
not NOT1 (N1882, N1848);
nor NOR2 (N1883, N1867, N1216);
or OR2 (N1884, N1880, N386);
nor NOR4 (N1885, N1884, N215, N1562, N1443);
nand NAND2 (N1886, N1885, N1531);
buf BUF1 (N1887, N1869);
buf BUF1 (N1888, N1866);
and AND4 (N1889, N1886, N506, N922, N1638);
and AND2 (N1890, N1883, N1674);
not NOT1 (N1891, N1875);
and AND3 (N1892, N1891, N390, N1695);
and AND4 (N1893, N1876, N233, N293, N1843);
nor NOR4 (N1894, N1881, N1210, N1097, N1890);
and AND2 (N1895, N1387, N1149);
buf BUF1 (N1896, N1894);
nand NAND4 (N1897, N1896, N1300, N211, N707);
buf BUF1 (N1898, N1897);
nand NAND3 (N1899, N1898, N1635, N1375);
xor XOR2 (N1900, N1892, N766);
xor XOR2 (N1901, N1889, N856);
nand NAND2 (N1902, N1901, N238);
not NOT1 (N1903, N1882);
xor XOR2 (N1904, N1879, N1416);
nand NAND2 (N1905, N1888, N676);
nor NOR4 (N1906, N1904, N1158, N394, N129);
xor XOR2 (N1907, N1902, N1134);
nor NOR3 (N1908, N1887, N821, N152);
or OR3 (N1909, N1906, N722, N658);
xor XOR2 (N1910, N1893, N1902);
buf BUF1 (N1911, N1873);
and AND4 (N1912, N1903, N895, N1680, N481);
not NOT1 (N1913, N1905);
xor XOR2 (N1914, N1913, N960);
nor NOR3 (N1915, N1912, N5, N270);
not NOT1 (N1916, N1908);
nor NOR2 (N1917, N1910, N1487);
or OR2 (N1918, N1914, N133);
xor XOR2 (N1919, N1918, N1877);
or OR2 (N1920, N1919, N1283);
not NOT1 (N1921, N1917);
nand NAND4 (N1922, N1900, N1249, N1432, N283);
not NOT1 (N1923, N1916);
and AND2 (N1924, N1921, N139);
nand NAND4 (N1925, N1924, N418, N260, N1294);
nand NAND2 (N1926, N1895, N983);
or OR3 (N1927, N1911, N649, N585);
xor XOR2 (N1928, N1899, N1589);
and AND4 (N1929, N1907, N1823, N1071, N574);
nand NAND4 (N1930, N1926, N83, N1770, N1337);
or OR4 (N1931, N1927, N55, N662, N751);
and AND2 (N1932, N1925, N355);
nand NAND2 (N1933, N1909, N837);
not NOT1 (N1934, N1933);
not NOT1 (N1935, N1923);
or OR3 (N1936, N1931, N82, N1926);
not NOT1 (N1937, N1934);
and AND4 (N1938, N1937, N559, N1877, N1215);
and AND3 (N1939, N1922, N295, N709);
not NOT1 (N1940, N1939);
xor XOR2 (N1941, N1932, N1716);
nand NAND4 (N1942, N1930, N1348, N232, N207);
buf BUF1 (N1943, N1936);
or OR3 (N1944, N1915, N1114, N790);
and AND4 (N1945, N1938, N80, N1914, N331);
or OR4 (N1946, N1935, N503, N1296, N1259);
nor NOR2 (N1947, N1942, N972);
xor XOR2 (N1948, N1928, N4);
nor NOR4 (N1949, N1946, N10, N1793, N2);
nand NAND4 (N1950, N1940, N1473, N1871, N608);
not NOT1 (N1951, N1920);
xor XOR2 (N1952, N1945, N329);
and AND2 (N1953, N1949, N1451);
buf BUF1 (N1954, N1941);
and AND2 (N1955, N1944, N266);
xor XOR2 (N1956, N1948, N1126);
nand NAND2 (N1957, N1953, N599);
buf BUF1 (N1958, N1957);
and AND2 (N1959, N1929, N1248);
and AND2 (N1960, N1959, N831);
or OR3 (N1961, N1958, N905, N1719);
xor XOR2 (N1962, N1952, N1666);
or OR2 (N1963, N1960, N1890);
xor XOR2 (N1964, N1947, N476);
nor NOR2 (N1965, N1962, N376);
buf BUF1 (N1966, N1956);
nand NAND4 (N1967, N1943, N612, N1876, N355);
buf BUF1 (N1968, N1950);
buf BUF1 (N1969, N1955);
xor XOR2 (N1970, N1954, N889);
not NOT1 (N1971, N1968);
and AND4 (N1972, N1970, N1296, N1109, N122);
and AND2 (N1973, N1972, N1459);
xor XOR2 (N1974, N1951, N1970);
and AND4 (N1975, N1969, N948, N1942, N373);
or OR4 (N1976, N1975, N59, N1347, N733);
xor XOR2 (N1977, N1963, N230);
not NOT1 (N1978, N1977);
nand NAND4 (N1979, N1961, N959, N1122, N304);
buf BUF1 (N1980, N1967);
or OR2 (N1981, N1971, N726);
buf BUF1 (N1982, N1965);
buf BUF1 (N1983, N1982);
and AND4 (N1984, N1974, N243, N1400, N1590);
and AND4 (N1985, N1984, N1676, N130, N261);
and AND4 (N1986, N1976, N42, N1783, N621);
not NOT1 (N1987, N1981);
buf BUF1 (N1988, N1979);
xor XOR2 (N1989, N1987, N476);
and AND2 (N1990, N1985, N1315);
nor NOR3 (N1991, N1986, N1089, N1282);
nand NAND3 (N1992, N1990, N1371, N1846);
or OR3 (N1993, N1980, N1822, N210);
xor XOR2 (N1994, N1983, N237);
not NOT1 (N1995, N1993);
xor XOR2 (N1996, N1978, N471);
and AND2 (N1997, N1996, N1362);
or OR4 (N1998, N1966, N1475, N110, N1955);
or OR3 (N1999, N1998, N1195, N1288);
and AND3 (N2000, N1994, N260, N1246);
or OR2 (N2001, N1992, N115);
not NOT1 (N2002, N1991);
or OR4 (N2003, N2000, N341, N1672, N1667);
buf BUF1 (N2004, N1973);
nor NOR4 (N2005, N1988, N1596, N1817, N933);
nand NAND4 (N2006, N2001, N1377, N427, N791);
and AND4 (N2007, N1995, N1731, N773, N1343);
xor XOR2 (N2008, N2007, N285);
and AND2 (N2009, N1999, N1718);
nor NOR2 (N2010, N1997, N478);
and AND4 (N2011, N1989, N1058, N186, N1727);
not NOT1 (N2012, N1964);
or OR2 (N2013, N2006, N510);
not NOT1 (N2014, N2012);
nand NAND2 (N2015, N2014, N1392);
xor XOR2 (N2016, N2015, N328);
nand NAND2 (N2017, N2003, N1637);
and AND3 (N2018, N2008, N959, N1485);
not NOT1 (N2019, N2016);
not NOT1 (N2020, N2011);
buf BUF1 (N2021, N2017);
nor NOR4 (N2022, N2005, N507, N878, N539);
nand NAND2 (N2023, N2004, N5);
or OR3 (N2024, N2013, N931, N626);
or OR2 (N2025, N2023, N678);
xor XOR2 (N2026, N2009, N199);
nand NAND4 (N2027, N2025, N830, N1716, N1422);
nand NAND3 (N2028, N2024, N486, N752);
nor NOR4 (N2029, N2026, N10, N725, N97);
nor NOR3 (N2030, N2010, N401, N766);
buf BUF1 (N2031, N2020);
nand NAND3 (N2032, N2028, N1400, N1075);
nand NAND2 (N2033, N2027, N1157);
buf BUF1 (N2034, N2021);
and AND2 (N2035, N2033, N215);
nor NOR4 (N2036, N2031, N626, N1239, N154);
or OR4 (N2037, N2035, N496, N64, N990);
nand NAND4 (N2038, N2030, N1528, N506, N298);
not NOT1 (N2039, N2032);
nand NAND4 (N2040, N2037, N454, N1470, N822);
nand NAND2 (N2041, N2029, N693);
or OR2 (N2042, N2036, N1982);
and AND3 (N2043, N2040, N1804, N1565);
or OR4 (N2044, N2042, N1262, N762, N2030);
nand NAND4 (N2045, N2002, N729, N940, N1560);
buf BUF1 (N2046, N2044);
and AND2 (N2047, N2043, N1079);
or OR2 (N2048, N2034, N379);
or OR4 (N2049, N2039, N1086, N1284, N495);
or OR3 (N2050, N2047, N138, N772);
and AND4 (N2051, N2048, N1109, N1967, N2020);
nor NOR4 (N2052, N2019, N1997, N456, N1748);
xor XOR2 (N2053, N2038, N734);
buf BUF1 (N2054, N2045);
nor NOR2 (N2055, N2022, N1078);
nand NAND2 (N2056, N2046, N258);
nand NAND3 (N2057, N2053, N1202, N193);
and AND4 (N2058, N2052, N1995, N508, N1048);
nor NOR2 (N2059, N2058, N411);
xor XOR2 (N2060, N2054, N1667);
or OR2 (N2061, N2060, N1058);
or OR3 (N2062, N2055, N1375, N2009);
buf BUF1 (N2063, N2018);
and AND2 (N2064, N2063, N1918);
or OR2 (N2065, N2041, N1708);
xor XOR2 (N2066, N2064, N992);
nand NAND2 (N2067, N2051, N540);
nand NAND3 (N2068, N2050, N1130, N87);
and AND4 (N2069, N2061, N212, N41, N268);
nand NAND3 (N2070, N2065, N1970, N1440);
and AND4 (N2071, N2057, N2038, N1930, N43);
xor XOR2 (N2072, N2066, N749);
xor XOR2 (N2073, N2067, N578);
and AND3 (N2074, N2068, N62, N1362);
and AND3 (N2075, N2071, N90, N96);
nand NAND2 (N2076, N2075, N1034);
and AND4 (N2077, N2062, N1601, N1412, N1457);
nor NOR4 (N2078, N2076, N26, N1549, N1431);
nand NAND2 (N2079, N2056, N1455);
nand NAND2 (N2080, N2073, N1331);
and AND3 (N2081, N2072, N1116, N1449);
or OR4 (N2082, N2079, N1472, N1321, N1813);
or OR3 (N2083, N2049, N471, N223);
not NOT1 (N2084, N2080);
nand NAND4 (N2085, N2069, N633, N1385, N1675);
not NOT1 (N2086, N2081);
nand NAND4 (N2087, N2074, N840, N914, N1291);
buf BUF1 (N2088, N2078);
or OR3 (N2089, N2083, N1653, N853);
buf BUF1 (N2090, N2059);
or OR4 (N2091, N2090, N1919, N789, N778);
buf BUF1 (N2092, N2088);
buf BUF1 (N2093, N2082);
nor NOR2 (N2094, N2087, N1287);
buf BUF1 (N2095, N2089);
not NOT1 (N2096, N2091);
and AND2 (N2097, N2093, N603);
buf BUF1 (N2098, N2092);
and AND4 (N2099, N2094, N1375, N1785, N582);
not NOT1 (N2100, N2070);
xor XOR2 (N2101, N2096, N113);
xor XOR2 (N2102, N2098, N1018);
nand NAND3 (N2103, N2095, N905, N1233);
nor NOR3 (N2104, N2099, N103, N74);
xor XOR2 (N2105, N2086, N465);
or OR2 (N2106, N2101, N782);
xor XOR2 (N2107, N2103, N831);
xor XOR2 (N2108, N2077, N1414);
nand NAND2 (N2109, N2107, N1703);
and AND4 (N2110, N2108, N1607, N66, N1877);
or OR4 (N2111, N2084, N410, N1907, N946);
buf BUF1 (N2112, N2100);
nor NOR4 (N2113, N2106, N158, N611, N1481);
not NOT1 (N2114, N2097);
nand NAND3 (N2115, N2085, N1659, N107);
buf BUF1 (N2116, N2115);
nand NAND3 (N2117, N2113, N1104, N1482);
and AND2 (N2118, N2116, N713);
nand NAND4 (N2119, N2114, N1471, N1573, N1832);
and AND2 (N2120, N2118, N966);
buf BUF1 (N2121, N2105);
and AND4 (N2122, N2102, N503, N966, N570);
buf BUF1 (N2123, N2122);
not NOT1 (N2124, N2104);
or OR2 (N2125, N2121, N1084);
not NOT1 (N2126, N2124);
and AND4 (N2127, N2117, N1211, N483, N765);
nand NAND2 (N2128, N2110, N1319);
nand NAND2 (N2129, N2126, N524);
or OR4 (N2130, N2112, N1034, N2123, N892);
nor NOR4 (N2131, N1320, N1782, N1752, N1992);
buf BUF1 (N2132, N2130);
and AND4 (N2133, N2131, N622, N1132, N398);
nand NAND3 (N2134, N2132, N62, N1811);
not NOT1 (N2135, N2111);
xor XOR2 (N2136, N2125, N3);
and AND4 (N2137, N2127, N821, N367, N532);
or OR4 (N2138, N2120, N1762, N625, N1450);
buf BUF1 (N2139, N2136);
nor NOR3 (N2140, N2135, N1403, N1531);
xor XOR2 (N2141, N2129, N489);
or OR2 (N2142, N2109, N992);
and AND3 (N2143, N2139, N370, N1935);
and AND4 (N2144, N2137, N1592, N325, N1007);
and AND3 (N2145, N2144, N642, N1491);
buf BUF1 (N2146, N2134);
nand NAND3 (N2147, N2138, N1024, N412);
and AND2 (N2148, N2143, N1612);
nor NOR3 (N2149, N2119, N272, N769);
and AND2 (N2150, N2148, N322);
nand NAND2 (N2151, N2142, N853);
nor NOR4 (N2152, N2141, N778, N727, N1245);
buf BUF1 (N2153, N2140);
and AND4 (N2154, N2149, N29, N1953, N496);
xor XOR2 (N2155, N2152, N548);
xor XOR2 (N2156, N2150, N1513);
or OR3 (N2157, N2147, N1508, N80);
nor NOR2 (N2158, N2146, N1053);
nor NOR2 (N2159, N2157, N156);
buf BUF1 (N2160, N2159);
nor NOR4 (N2161, N2151, N73, N2066, N282);
not NOT1 (N2162, N2153);
nand NAND2 (N2163, N2161, N1913);
not NOT1 (N2164, N2160);
or OR3 (N2165, N2133, N917, N1344);
nand NAND4 (N2166, N2156, N600, N411, N1343);
xor XOR2 (N2167, N2165, N119);
and AND3 (N2168, N2164, N1178, N1168);
buf BUF1 (N2169, N2155);
nand NAND2 (N2170, N2168, N1823);
xor XOR2 (N2171, N2166, N344);
nor NOR4 (N2172, N2154, N785, N1719, N821);
buf BUF1 (N2173, N2145);
or OR3 (N2174, N2172, N1370, N1146);
not NOT1 (N2175, N2128);
buf BUF1 (N2176, N2158);
and AND4 (N2177, N2163, N1275, N2176, N947);
not NOT1 (N2178, N745);
buf BUF1 (N2179, N2171);
nand NAND4 (N2180, N2173, N1178, N1439, N1469);
not NOT1 (N2181, N2177);
and AND4 (N2182, N2174, N1085, N2117, N1574);
nor NOR2 (N2183, N2169, N151);
nor NOR4 (N2184, N2181, N345, N884, N419);
nor NOR2 (N2185, N2167, N792);
not NOT1 (N2186, N2170);
buf BUF1 (N2187, N2185);
xor XOR2 (N2188, N2187, N1530);
or OR3 (N2189, N2162, N376, N1247);
xor XOR2 (N2190, N2178, N1317);
xor XOR2 (N2191, N2190, N2083);
nand NAND2 (N2192, N2188, N375);
xor XOR2 (N2193, N2189, N694);
nand NAND2 (N2194, N2180, N1589);
not NOT1 (N2195, N2182);
buf BUF1 (N2196, N2183);
buf BUF1 (N2197, N2195);
or OR2 (N2198, N2184, N586);
not NOT1 (N2199, N2192);
not NOT1 (N2200, N2196);
nand NAND4 (N2201, N2194, N281, N341, N634);
nand NAND3 (N2202, N2175, N1465, N952);
and AND3 (N2203, N2199, N1629, N1106);
buf BUF1 (N2204, N2186);
nand NAND4 (N2205, N2202, N695, N701, N1293);
not NOT1 (N2206, N2203);
buf BUF1 (N2207, N2179);
and AND3 (N2208, N2204, N2091, N99);
and AND4 (N2209, N2206, N308, N689, N1432);
or OR2 (N2210, N2209, N502);
and AND4 (N2211, N2208, N1697, N1962, N1999);
nand NAND4 (N2212, N2191, N1388, N1492, N84);
not NOT1 (N2213, N2198);
not NOT1 (N2214, N2211);
nor NOR4 (N2215, N2213, N474, N2188, N1782);
or OR2 (N2216, N2210, N118);
buf BUF1 (N2217, N2215);
xor XOR2 (N2218, N2214, N1227);
and AND3 (N2219, N2197, N2108, N229);
not NOT1 (N2220, N2193);
nand NAND4 (N2221, N2216, N921, N915, N273);
nor NOR3 (N2222, N2200, N2093, N188);
xor XOR2 (N2223, N2222, N1302);
xor XOR2 (N2224, N2221, N358);
xor XOR2 (N2225, N2223, N888);
not NOT1 (N2226, N2225);
buf BUF1 (N2227, N2205);
buf BUF1 (N2228, N2227);
buf BUF1 (N2229, N2218);
not NOT1 (N2230, N2207);
and AND3 (N2231, N2230, N1001, N257);
not NOT1 (N2232, N2224);
buf BUF1 (N2233, N2219);
buf BUF1 (N2234, N2212);
nand NAND2 (N2235, N2231, N542);
and AND3 (N2236, N2217, N1171, N514);
and AND2 (N2237, N2233, N794);
and AND4 (N2238, N2220, N822, N857, N532);
nor NOR4 (N2239, N2228, N1327, N486, N718);
or OR3 (N2240, N2229, N2111, N993);
not NOT1 (N2241, N2232);
nor NOR4 (N2242, N2240, N731, N1646, N1902);
not NOT1 (N2243, N2235);
xor XOR2 (N2244, N2242, N1710);
or OR4 (N2245, N2244, N263, N1000, N361);
nand NAND3 (N2246, N2238, N1300, N1173);
or OR4 (N2247, N2241, N990, N941, N970);
nor NOR4 (N2248, N2239, N584, N1152, N78);
or OR4 (N2249, N2248, N2109, N1139, N2014);
buf BUF1 (N2250, N2247);
not NOT1 (N2251, N2236);
not NOT1 (N2252, N2251);
not NOT1 (N2253, N2252);
not NOT1 (N2254, N2253);
xor XOR2 (N2255, N2245, N1875);
and AND2 (N2256, N2201, N2133);
and AND2 (N2257, N2243, N113);
or OR4 (N2258, N2256, N1271, N1679, N1471);
nand NAND2 (N2259, N2257, N598);
buf BUF1 (N2260, N2249);
or OR4 (N2261, N2258, N869, N1210, N1443);
buf BUF1 (N2262, N2250);
and AND4 (N2263, N2254, N1761, N254, N113);
and AND4 (N2264, N2237, N1967, N291, N584);
nand NAND2 (N2265, N2226, N266);
nor NOR4 (N2266, N2261, N346, N255, N1408);
buf BUF1 (N2267, N2262);
xor XOR2 (N2268, N2266, N1414);
or OR2 (N2269, N2259, N1532);
xor XOR2 (N2270, N2265, N1618);
buf BUF1 (N2271, N2268);
nand NAND3 (N2272, N2246, N1620, N981);
or OR3 (N2273, N2271, N487, N1456);
nor NOR2 (N2274, N2270, N1818);
xor XOR2 (N2275, N2263, N1509);
nand NAND3 (N2276, N2234, N1221, N1138);
and AND4 (N2277, N2276, N73, N1410, N2148);
not NOT1 (N2278, N2272);
buf BUF1 (N2279, N2277);
not NOT1 (N2280, N2255);
not NOT1 (N2281, N2274);
nor NOR4 (N2282, N2260, N119, N1459, N270);
or OR4 (N2283, N2281, N1982, N257, N365);
nand NAND4 (N2284, N2273, N178, N1616, N842);
xor XOR2 (N2285, N2283, N109);
and AND4 (N2286, N2275, N1685, N447, N659);
xor XOR2 (N2287, N2284, N933);
and AND4 (N2288, N2287, N1903, N1930, N1556);
not NOT1 (N2289, N2267);
or OR3 (N2290, N2286, N294, N2269);
xor XOR2 (N2291, N1930, N2279);
xor XOR2 (N2292, N956, N182);
nor NOR4 (N2293, N2264, N2086, N1078, N1373);
buf BUF1 (N2294, N2290);
or OR3 (N2295, N2291, N1678, N292);
xor XOR2 (N2296, N2285, N1244);
xor XOR2 (N2297, N2295, N471);
not NOT1 (N2298, N2292);
not NOT1 (N2299, N2289);
or OR3 (N2300, N2293, N1251, N933);
or OR3 (N2301, N2280, N1787, N129);
not NOT1 (N2302, N2299);
and AND2 (N2303, N2278, N219);
buf BUF1 (N2304, N2296);
nand NAND2 (N2305, N2294, N1466);
nand NAND2 (N2306, N2288, N513);
nand NAND2 (N2307, N2282, N1996);
buf BUF1 (N2308, N2305);
xor XOR2 (N2309, N2307, N1429);
xor XOR2 (N2310, N2308, N1480);
not NOT1 (N2311, N2306);
xor XOR2 (N2312, N2310, N1524);
xor XOR2 (N2313, N2300, N1169);
or OR2 (N2314, N2301, N2219);
or OR3 (N2315, N2314, N1211, N625);
or OR2 (N2316, N2312, N2047);
xor XOR2 (N2317, N2302, N418);
or OR2 (N2318, N2311, N48);
and AND2 (N2319, N2313, N2191);
and AND2 (N2320, N2316, N1685);
nand NAND2 (N2321, N2304, N965);
xor XOR2 (N2322, N2320, N582);
xor XOR2 (N2323, N2303, N793);
or OR3 (N2324, N2317, N943, N909);
or OR2 (N2325, N2318, N509);
xor XOR2 (N2326, N2325, N618);
or OR2 (N2327, N2315, N2260);
and AND2 (N2328, N2326, N1506);
not NOT1 (N2329, N2319);
nand NAND3 (N2330, N2328, N840, N1015);
buf BUF1 (N2331, N2330);
nand NAND2 (N2332, N2309, N884);
or OR3 (N2333, N2323, N444, N1280);
or OR4 (N2334, N2324, N2188, N2026, N790);
not NOT1 (N2335, N2329);
not NOT1 (N2336, N2333);
not NOT1 (N2337, N2297);
xor XOR2 (N2338, N2321, N882);
not NOT1 (N2339, N2334);
and AND3 (N2340, N2327, N1821, N1618);
or OR2 (N2341, N2331, N1771);
nor NOR3 (N2342, N2341, N2220, N800);
not NOT1 (N2343, N2338);
nand NAND3 (N2344, N2332, N1892, N1943);
or OR3 (N2345, N2322, N1280, N784);
nor NOR2 (N2346, N2336, N262);
not NOT1 (N2347, N2340);
or OR4 (N2348, N2343, N473, N846, N1370);
nand NAND3 (N2349, N2347, N1379, N1382);
xor XOR2 (N2350, N2345, N902);
and AND3 (N2351, N2337, N2138, N289);
buf BUF1 (N2352, N2335);
not NOT1 (N2353, N2352);
nand NAND2 (N2354, N2348, N1496);
buf BUF1 (N2355, N2346);
not NOT1 (N2356, N2351);
and AND4 (N2357, N2342, N457, N680, N358);
buf BUF1 (N2358, N2357);
buf BUF1 (N2359, N2353);
or OR3 (N2360, N2356, N252, N2215);
or OR2 (N2361, N2349, N2272);
nor NOR2 (N2362, N2298, N1496);
not NOT1 (N2363, N2355);
or OR2 (N2364, N2360, N1964);
buf BUF1 (N2365, N2358);
xor XOR2 (N2366, N2359, N2041);
xor XOR2 (N2367, N2362, N2269);
nand NAND3 (N2368, N2344, N1881, N282);
buf BUF1 (N2369, N2350);
buf BUF1 (N2370, N2369);
xor XOR2 (N2371, N2368, N2242);
not NOT1 (N2372, N2366);
not NOT1 (N2373, N2372);
nor NOR3 (N2374, N2365, N1478, N2023);
nor NOR3 (N2375, N2371, N1755, N1358);
xor XOR2 (N2376, N2373, N1301);
not NOT1 (N2377, N2367);
nor NOR3 (N2378, N2363, N1343, N1072);
xor XOR2 (N2379, N2374, N495);
xor XOR2 (N2380, N2379, N1737);
xor XOR2 (N2381, N2364, N948);
not NOT1 (N2382, N2377);
xor XOR2 (N2383, N2380, N2236);
xor XOR2 (N2384, N2354, N2362);
not NOT1 (N2385, N2382);
xor XOR2 (N2386, N2376, N744);
nand NAND2 (N2387, N2383, N967);
nand NAND4 (N2388, N2339, N548, N2118, N745);
nand NAND3 (N2389, N2361, N1082, N383);
nand NAND3 (N2390, N2388, N537, N1532);
not NOT1 (N2391, N2389);
and AND4 (N2392, N2387, N2013, N458, N1928);
or OR2 (N2393, N2384, N429);
or OR4 (N2394, N2378, N918, N612, N1230);
nand NAND3 (N2395, N2381, N843, N609);
and AND3 (N2396, N2393, N2258, N150);
and AND4 (N2397, N2395, N468, N1460, N2086);
and AND2 (N2398, N2397, N740);
not NOT1 (N2399, N2375);
nor NOR4 (N2400, N2399, N1556, N1103, N1645);
not NOT1 (N2401, N2396);
or OR3 (N2402, N2400, N1172, N709);
and AND4 (N2403, N2385, N123, N1497, N1770);
not NOT1 (N2404, N2394);
xor XOR2 (N2405, N2398, N2256);
xor XOR2 (N2406, N2370, N1410);
nand NAND3 (N2407, N2402, N1958, N2006);
buf BUF1 (N2408, N2390);
nand NAND3 (N2409, N2408, N2395, N540);
xor XOR2 (N2410, N2392, N1974);
not NOT1 (N2411, N2391);
or OR2 (N2412, N2404, N1131);
xor XOR2 (N2413, N2406, N1106);
and AND2 (N2414, N2410, N2124);
xor XOR2 (N2415, N2413, N1200);
nand NAND4 (N2416, N2407, N2090, N957, N1255);
xor XOR2 (N2417, N2411, N1309);
nand NAND2 (N2418, N2405, N527);
or OR3 (N2419, N2409, N1630, N2291);
buf BUF1 (N2420, N2416);
nand NAND3 (N2421, N2417, N296, N238);
xor XOR2 (N2422, N2419, N184);
or OR4 (N2423, N2421, N209, N2196, N1249);
buf BUF1 (N2424, N2412);
xor XOR2 (N2425, N2420, N442);
or OR3 (N2426, N2425, N1771, N1956);
or OR3 (N2427, N2424, N743, N1939);
xor XOR2 (N2428, N2427, N1436);
nand NAND4 (N2429, N2415, N580, N949, N924);
buf BUF1 (N2430, N2422);
and AND3 (N2431, N2414, N1006, N288);
xor XOR2 (N2432, N2386, N708);
nand NAND2 (N2433, N2429, N563);
buf BUF1 (N2434, N2426);
xor XOR2 (N2435, N2401, N39);
nand NAND4 (N2436, N2428, N851, N973, N1920);
nand NAND2 (N2437, N2433, N1838);
xor XOR2 (N2438, N2431, N2213);
xor XOR2 (N2439, N2434, N2352);
not NOT1 (N2440, N2437);
not NOT1 (N2441, N2423);
and AND3 (N2442, N2418, N2276, N805);
nor NOR4 (N2443, N2438, N2300, N2428, N1419);
nand NAND4 (N2444, N2403, N1134, N1325, N762);
or OR3 (N2445, N2432, N87, N2291);
xor XOR2 (N2446, N2445, N459);
and AND2 (N2447, N2435, N1706);
not NOT1 (N2448, N2444);
buf BUF1 (N2449, N2441);
and AND4 (N2450, N2449, N1776, N2285, N1112);
nor NOR2 (N2451, N2448, N1355);
buf BUF1 (N2452, N2442);
nand NAND4 (N2453, N2443, N1999, N28, N546);
buf BUF1 (N2454, N2430);
nand NAND4 (N2455, N2454, N2046, N1904, N267);
xor XOR2 (N2456, N2451, N142);
xor XOR2 (N2457, N2450, N1613);
buf BUF1 (N2458, N2453);
xor XOR2 (N2459, N2457, N1278);
buf BUF1 (N2460, N2459);
xor XOR2 (N2461, N2455, N1473);
buf BUF1 (N2462, N2436);
nand NAND4 (N2463, N2439, N476, N621, N385);
xor XOR2 (N2464, N2447, N455);
xor XOR2 (N2465, N2458, N884);
xor XOR2 (N2466, N2462, N570);
buf BUF1 (N2467, N2452);
not NOT1 (N2468, N2465);
not NOT1 (N2469, N2461);
xor XOR2 (N2470, N2466, N2285);
not NOT1 (N2471, N2468);
and AND3 (N2472, N2463, N1992, N1138);
nand NAND4 (N2473, N2472, N1481, N703, N2197);
xor XOR2 (N2474, N2471, N561);
and AND2 (N2475, N2464, N1019);
and AND4 (N2476, N2475, N1599, N402, N2187);
nand NAND4 (N2477, N2446, N2059, N273, N1178);
and AND2 (N2478, N2476, N264);
buf BUF1 (N2479, N2474);
and AND3 (N2480, N2470, N1300, N551);
nor NOR3 (N2481, N2473, N1136, N1255);
and AND2 (N2482, N2478, N1730);
xor XOR2 (N2483, N2460, N1741);
and AND2 (N2484, N2482, N469);
and AND2 (N2485, N2479, N1712);
nor NOR4 (N2486, N2480, N107, N265, N1571);
nand NAND4 (N2487, N2467, N1822, N1902, N1121);
buf BUF1 (N2488, N2483);
not NOT1 (N2489, N2487);
or OR4 (N2490, N2456, N2471, N1667, N1209);
buf BUF1 (N2491, N2484);
and AND3 (N2492, N2489, N2240, N1958);
and AND3 (N2493, N2490, N912, N1932);
nor NOR4 (N2494, N2485, N2, N229, N155);
not NOT1 (N2495, N2492);
nor NOR3 (N2496, N2491, N1083, N1235);
not NOT1 (N2497, N2494);
nor NOR2 (N2498, N2495, N962);
buf BUF1 (N2499, N2486);
nand NAND4 (N2500, N2469, N1576, N1987, N1270);
not NOT1 (N2501, N2498);
nor NOR2 (N2502, N2499, N2186);
xor XOR2 (N2503, N2500, N1949);
buf BUF1 (N2504, N2477);
or OR2 (N2505, N2488, N974);
nand NAND3 (N2506, N2496, N1058, N223);
nor NOR3 (N2507, N2497, N507, N1523);
nor NOR3 (N2508, N2493, N2237, N1113);
xor XOR2 (N2509, N2508, N562);
or OR4 (N2510, N2507, N2482, N362, N947);
or OR3 (N2511, N2506, N98, N1855);
nor NOR3 (N2512, N2505, N1453, N503);
not NOT1 (N2513, N2511);
xor XOR2 (N2514, N2513, N822);
not NOT1 (N2515, N2510);
nor NOR2 (N2516, N2440, N1398);
buf BUF1 (N2517, N2503);
xor XOR2 (N2518, N2501, N1768);
buf BUF1 (N2519, N2509);
buf BUF1 (N2520, N2504);
and AND3 (N2521, N2481, N427, N2474);
not NOT1 (N2522, N2514);
xor XOR2 (N2523, N2519, N1109);
or OR3 (N2524, N2520, N1477, N1569);
nand NAND2 (N2525, N2517, N621);
or OR2 (N2526, N2523, N410);
and AND3 (N2527, N2502, N1304, N1111);
not NOT1 (N2528, N2526);
not NOT1 (N2529, N2512);
nand NAND3 (N2530, N2528, N894, N1710);
nand NAND2 (N2531, N2518, N2027);
nor NOR2 (N2532, N2516, N902);
nor NOR4 (N2533, N2527, N237, N2030, N755);
nor NOR3 (N2534, N2525, N909, N2223);
buf BUF1 (N2535, N2522);
and AND2 (N2536, N2533, N681);
xor XOR2 (N2537, N2515, N793);
nand NAND2 (N2538, N2537, N1465);
xor XOR2 (N2539, N2531, N1808);
buf BUF1 (N2540, N2530);
and AND3 (N2541, N2524, N772, N244);
not NOT1 (N2542, N2538);
xor XOR2 (N2543, N2534, N823);
buf BUF1 (N2544, N2536);
or OR3 (N2545, N2532, N714, N2519);
or OR4 (N2546, N2540, N1523, N1839, N1551);
nor NOR4 (N2547, N2535, N1946, N1225, N2133);
nor NOR3 (N2548, N2541, N985, N874);
and AND3 (N2549, N2547, N1012, N164);
nor NOR4 (N2550, N2546, N1176, N1292, N209);
nand NAND2 (N2551, N2521, N1878);
not NOT1 (N2552, N2543);
nor NOR3 (N2553, N2544, N1823, N1404);
nor NOR3 (N2554, N2551, N2398, N506);
nor NOR2 (N2555, N2548, N2519);
buf BUF1 (N2556, N2554);
xor XOR2 (N2557, N2550, N800);
and AND4 (N2558, N2556, N210, N1590, N1608);
nand NAND2 (N2559, N2558, N778);
nor NOR4 (N2560, N2542, N1963, N296, N1553);
or OR2 (N2561, N2560, N2225);
nand NAND2 (N2562, N2545, N231);
or OR2 (N2563, N2559, N1240);
xor XOR2 (N2564, N2555, N406);
xor XOR2 (N2565, N2563, N2013);
or OR4 (N2566, N2539, N1380, N1989, N2170);
buf BUF1 (N2567, N2564);
nor NOR3 (N2568, N2565, N2392, N1854);
or OR3 (N2569, N2553, N741, N2148);
or OR4 (N2570, N2557, N1221, N1276, N526);
nand NAND4 (N2571, N2561, N2163, N2053, N2555);
xor XOR2 (N2572, N2569, N891);
nor NOR4 (N2573, N2549, N1826, N68, N890);
xor XOR2 (N2574, N2567, N1396);
or OR3 (N2575, N2571, N883, N2232);
nand NAND4 (N2576, N2573, N653, N490, N1897);
and AND3 (N2577, N2552, N182, N977);
and AND4 (N2578, N2576, N1623, N1250, N1817);
or OR2 (N2579, N2575, N80);
buf BUF1 (N2580, N2574);
nor NOR4 (N2581, N2568, N1425, N747, N653);
and AND3 (N2582, N2562, N413, N226);
xor XOR2 (N2583, N2579, N1030);
nor NOR4 (N2584, N2583, N1001, N1825, N2399);
nand NAND3 (N2585, N2529, N2232, N1643);
and AND3 (N2586, N2578, N1620, N766);
xor XOR2 (N2587, N2585, N2358);
and AND4 (N2588, N2572, N2374, N281, N787);
xor XOR2 (N2589, N2581, N385);
nor NOR4 (N2590, N2589, N964, N949, N283);
and AND4 (N2591, N2587, N2055, N1588, N2058);
not NOT1 (N2592, N2570);
xor XOR2 (N2593, N2592, N2205);
and AND3 (N2594, N2580, N1717, N414);
and AND3 (N2595, N2591, N1607, N2203);
nor NOR3 (N2596, N2577, N1230, N1838);
buf BUF1 (N2597, N2595);
nand NAND3 (N2598, N2566, N1131, N786);
nor NOR4 (N2599, N2593, N872, N2142, N2104);
xor XOR2 (N2600, N2590, N1267);
nor NOR2 (N2601, N2597, N1316);
buf BUF1 (N2602, N2588);
buf BUF1 (N2603, N2586);
buf BUF1 (N2604, N2599);
or OR3 (N2605, N2584, N274, N955);
or OR3 (N2606, N2600, N2513, N504);
and AND2 (N2607, N2605, N751);
xor XOR2 (N2608, N2582, N472);
or OR3 (N2609, N2601, N1245, N1354);
not NOT1 (N2610, N2598);
not NOT1 (N2611, N2603);
xor XOR2 (N2612, N2596, N2058);
nor NOR3 (N2613, N2612, N1871, N2474);
nor NOR3 (N2614, N2611, N70, N2122);
nand NAND4 (N2615, N2602, N85, N1367, N1117);
not NOT1 (N2616, N2613);
and AND2 (N2617, N2608, N598);
nand NAND4 (N2618, N2610, N511, N1917, N375);
nor NOR2 (N2619, N2594, N1611);
buf BUF1 (N2620, N2617);
xor XOR2 (N2621, N2616, N368);
and AND4 (N2622, N2607, N1504, N1858, N2452);
xor XOR2 (N2623, N2609, N1559);
and AND3 (N2624, N2619, N1991, N1300);
buf BUF1 (N2625, N2621);
buf BUF1 (N2626, N2614);
nor NOR2 (N2627, N2625, N2292);
xor XOR2 (N2628, N2624, N1147);
nand NAND4 (N2629, N2622, N900, N134, N837);
nand NAND2 (N2630, N2627, N2322);
or OR2 (N2631, N2630, N617);
xor XOR2 (N2632, N2626, N1044);
buf BUF1 (N2633, N2632);
xor XOR2 (N2634, N2633, N585);
xor XOR2 (N2635, N2606, N1654);
not NOT1 (N2636, N2631);
buf BUF1 (N2637, N2618);
or OR2 (N2638, N2604, N1259);
nand NAND3 (N2639, N2629, N949, N699);
buf BUF1 (N2640, N2634);
nor NOR2 (N2641, N2628, N618);
and AND4 (N2642, N2615, N570, N2085, N830);
buf BUF1 (N2643, N2640);
or OR4 (N2644, N2641, N816, N313, N1906);
and AND3 (N2645, N2642, N628, N643);
xor XOR2 (N2646, N2623, N2485);
nand NAND4 (N2647, N2643, N2616, N1581, N2426);
xor XOR2 (N2648, N2644, N3);
nand NAND2 (N2649, N2647, N1513);
not NOT1 (N2650, N2648);
xor XOR2 (N2651, N2650, N506);
or OR4 (N2652, N2637, N106, N2295, N1863);
nor NOR2 (N2653, N2639, N2370);
nand NAND2 (N2654, N2620, N213);
buf BUF1 (N2655, N2649);
and AND2 (N2656, N2652, N175);
and AND3 (N2657, N2635, N1513, N1465);
and AND3 (N2658, N2638, N663, N2410);
buf BUF1 (N2659, N2656);
nand NAND2 (N2660, N2654, N655);
or OR4 (N2661, N2659, N2318, N926, N1848);
nand NAND2 (N2662, N2651, N1448);
buf BUF1 (N2663, N2636);
and AND4 (N2664, N2646, N1118, N1328, N1872);
and AND4 (N2665, N2658, N1152, N101, N1977);
buf BUF1 (N2666, N2662);
and AND4 (N2667, N2661, N2130, N1896, N1206);
nand NAND4 (N2668, N2663, N1928, N912, N196);
nor NOR4 (N2669, N2664, N470, N1551, N2557);
and AND3 (N2670, N2669, N2272, N216);
nand NAND4 (N2671, N2660, N2473, N157, N259);
and AND2 (N2672, N2657, N1543);
nand NAND2 (N2673, N2665, N1034);
nand NAND3 (N2674, N2667, N2079, N463);
nand NAND3 (N2675, N2674, N169, N1076);
or OR4 (N2676, N2671, N2340, N2649, N947);
nand NAND4 (N2677, N2672, N1867, N2079, N531);
or OR4 (N2678, N2675, N412, N654, N1083);
nand NAND2 (N2679, N2668, N1456);
xor XOR2 (N2680, N2655, N82);
nand NAND3 (N2681, N2670, N900, N64);
and AND3 (N2682, N2673, N663, N2371);
not NOT1 (N2683, N2645);
not NOT1 (N2684, N2683);
nor NOR3 (N2685, N2677, N587, N965);
nand NAND2 (N2686, N2681, N815);
or OR4 (N2687, N2679, N2447, N95, N809);
nor NOR4 (N2688, N2676, N1326, N2227, N2505);
xor XOR2 (N2689, N2678, N2630);
xor XOR2 (N2690, N2689, N2462);
nor NOR2 (N2691, N2687, N1302);
or OR3 (N2692, N2690, N1219, N1929);
nor NOR4 (N2693, N2692, N542, N241, N1092);
nand NAND2 (N2694, N2685, N319);
or OR2 (N2695, N2684, N638);
buf BUF1 (N2696, N2693);
or OR3 (N2697, N2686, N802, N258);
xor XOR2 (N2698, N2697, N2460);
and AND4 (N2699, N2698, N2277, N806, N856);
nor NOR3 (N2700, N2682, N2448, N1265);
and AND3 (N2701, N2680, N2386, N474);
nand NAND4 (N2702, N2701, N893, N1019, N1152);
not NOT1 (N2703, N2700);
or OR2 (N2704, N2694, N2482);
nand NAND3 (N2705, N2691, N336, N464);
nand NAND4 (N2706, N2695, N2422, N1028, N1069);
not NOT1 (N2707, N2702);
buf BUF1 (N2708, N2704);
or OR4 (N2709, N2699, N941, N1959, N92);
and AND4 (N2710, N2666, N1256, N1268, N824);
or OR3 (N2711, N2709, N2588, N66);
or OR2 (N2712, N2711, N153);
nand NAND4 (N2713, N2706, N816, N1621, N2461);
not NOT1 (N2714, N2705);
buf BUF1 (N2715, N2707);
nand NAND2 (N2716, N2710, N2230);
and AND4 (N2717, N2696, N1126, N613, N1276);
and AND3 (N2718, N2712, N91, N1879);
and AND3 (N2719, N2715, N1171, N573);
or OR4 (N2720, N2714, N2279, N1132, N2301);
buf BUF1 (N2721, N2719);
not NOT1 (N2722, N2688);
nand NAND4 (N2723, N2717, N1570, N894, N1005);
not NOT1 (N2724, N2716);
nand NAND3 (N2725, N2713, N2698, N118);
not NOT1 (N2726, N2653);
nand NAND2 (N2727, N2718, N953);
buf BUF1 (N2728, N2721);
nor NOR4 (N2729, N2726, N853, N1004, N139);
nor NOR2 (N2730, N2728, N2481);
not NOT1 (N2731, N2708);
and AND2 (N2732, N2722, N20);
nand NAND3 (N2733, N2727, N553, N1316);
or OR2 (N2734, N2732, N625);
not NOT1 (N2735, N2730);
nor NOR3 (N2736, N2703, N726, N845);
not NOT1 (N2737, N2736);
xor XOR2 (N2738, N2723, N1784);
buf BUF1 (N2739, N2731);
and AND3 (N2740, N2739, N2235, N968);
and AND2 (N2741, N2738, N701);
nand NAND2 (N2742, N2737, N1164);
xor XOR2 (N2743, N2742, N120);
not NOT1 (N2744, N2720);
or OR3 (N2745, N2733, N457, N508);
nand NAND3 (N2746, N2744, N1555, N1328);
buf BUF1 (N2747, N2735);
nand NAND3 (N2748, N2729, N742, N1539);
buf BUF1 (N2749, N2734);
nor NOR2 (N2750, N2741, N2092);
nor NOR3 (N2751, N2743, N1206, N120);
buf BUF1 (N2752, N2740);
and AND2 (N2753, N2751, N1711);
and AND2 (N2754, N2748, N1603);
not NOT1 (N2755, N2746);
or OR2 (N2756, N2753, N2688);
not NOT1 (N2757, N2749);
buf BUF1 (N2758, N2750);
or OR4 (N2759, N2725, N114, N1313, N1560);
and AND4 (N2760, N2752, N1627, N304, N382);
buf BUF1 (N2761, N2756);
xor XOR2 (N2762, N2758, N620);
buf BUF1 (N2763, N2747);
nand NAND4 (N2764, N2757, N2036, N747, N2740);
nand NAND3 (N2765, N2761, N2075, N2662);
not NOT1 (N2766, N2755);
and AND3 (N2767, N2763, N563, N468);
not NOT1 (N2768, N2760);
buf BUF1 (N2769, N2724);
buf BUF1 (N2770, N2745);
not NOT1 (N2771, N2768);
buf BUF1 (N2772, N2759);
and AND4 (N2773, N2762, N1799, N2654, N1235);
nand NAND2 (N2774, N2754, N1052);
or OR3 (N2775, N2769, N1131, N1562);
buf BUF1 (N2776, N2772);
nor NOR4 (N2777, N2775, N466, N830, N1593);
nor NOR2 (N2778, N2774, N1783);
not NOT1 (N2779, N2773);
nor NOR4 (N2780, N2771, N2716, N2079, N935);
not NOT1 (N2781, N2766);
or OR4 (N2782, N2776, N848, N607, N18);
buf BUF1 (N2783, N2782);
buf BUF1 (N2784, N2765);
not NOT1 (N2785, N2783);
nor NOR3 (N2786, N2778, N1944, N2018);
xor XOR2 (N2787, N2777, N1096);
not NOT1 (N2788, N2764);
nor NOR3 (N2789, N2770, N1027, N543);
buf BUF1 (N2790, N2767);
not NOT1 (N2791, N2781);
and AND4 (N2792, N2789, N592, N109, N1702);
not NOT1 (N2793, N2785);
not NOT1 (N2794, N2788);
xor XOR2 (N2795, N2779, N2500);
or OR2 (N2796, N2784, N911);
nand NAND4 (N2797, N2786, N2692, N2258, N1651);
and AND2 (N2798, N2797, N872);
nor NOR3 (N2799, N2798, N2363, N2684);
and AND3 (N2800, N2791, N1883, N669);
or OR2 (N2801, N2793, N705);
buf BUF1 (N2802, N2801);
or OR2 (N2803, N2800, N459);
and AND4 (N2804, N2799, N1684, N1199, N1622);
buf BUF1 (N2805, N2796);
xor XOR2 (N2806, N2787, N99);
and AND3 (N2807, N2795, N1267, N330);
and AND2 (N2808, N2802, N182);
nor NOR2 (N2809, N2792, N2784);
or OR3 (N2810, N2803, N2008, N1254);
nor NOR4 (N2811, N2808, N2466, N1132, N1797);
or OR3 (N2812, N2805, N1, N1769);
and AND4 (N2813, N2810, N2168, N1515, N2689);
not NOT1 (N2814, N2790);
nor NOR4 (N2815, N2809, N625, N2524, N1689);
and AND2 (N2816, N2794, N748);
not NOT1 (N2817, N2812);
and AND3 (N2818, N2804, N1475, N1035);
buf BUF1 (N2819, N2780);
buf BUF1 (N2820, N2807);
not NOT1 (N2821, N2817);
and AND4 (N2822, N2813, N1568, N103, N430);
nand NAND4 (N2823, N2818, N1368, N1855, N2216);
and AND4 (N2824, N2820, N1818, N1783, N221);
buf BUF1 (N2825, N2819);
buf BUF1 (N2826, N2825);
xor XOR2 (N2827, N2826, N2747);
buf BUF1 (N2828, N2814);
and AND4 (N2829, N2816, N1664, N1018, N144);
not NOT1 (N2830, N2821);
or OR4 (N2831, N2824, N197, N772, N834);
xor XOR2 (N2832, N2815, N1942);
nand NAND3 (N2833, N2806, N890, N513);
or OR3 (N2834, N2832, N1478, N1184);
buf BUF1 (N2835, N2811);
xor XOR2 (N2836, N2823, N61);
nand NAND4 (N2837, N2828, N1598, N1146, N2421);
buf BUF1 (N2838, N2837);
not NOT1 (N2839, N2835);
or OR3 (N2840, N2829, N2169, N860);
or OR3 (N2841, N2834, N1674, N177);
or OR4 (N2842, N2830, N1927, N2243, N550);
nor NOR4 (N2843, N2827, N559, N759, N2401);
buf BUF1 (N2844, N2841);
or OR2 (N2845, N2843, N1700);
and AND3 (N2846, N2838, N1417, N1786);
and AND2 (N2847, N2845, N2820);
not NOT1 (N2848, N2822);
not NOT1 (N2849, N2844);
nand NAND2 (N2850, N2848, N2398);
nand NAND3 (N2851, N2839, N1422, N1399);
or OR4 (N2852, N2847, N924, N1444, N1604);
buf BUF1 (N2853, N2850);
buf BUF1 (N2854, N2833);
nor NOR2 (N2855, N2851, N243);
buf BUF1 (N2856, N2840);
or OR3 (N2857, N2854, N2152, N2249);
and AND3 (N2858, N2853, N1837, N2668);
not NOT1 (N2859, N2831);
buf BUF1 (N2860, N2859);
nor NOR3 (N2861, N2857, N1603, N2356);
xor XOR2 (N2862, N2849, N802);
nor NOR4 (N2863, N2858, N110, N2125, N640);
and AND2 (N2864, N2863, N344);
and AND4 (N2865, N2836, N1581, N2762, N357);
xor XOR2 (N2866, N2865, N48);
nand NAND2 (N2867, N2856, N2804);
and AND2 (N2868, N2855, N2605);
or OR4 (N2869, N2862, N579, N1777, N1151);
buf BUF1 (N2870, N2852);
nor NOR3 (N2871, N2846, N2627, N2161);
nor NOR2 (N2872, N2861, N926);
and AND3 (N2873, N2871, N294, N413);
buf BUF1 (N2874, N2864);
or OR2 (N2875, N2869, N885);
not NOT1 (N2876, N2872);
nor NOR4 (N2877, N2874, N2674, N2179, N578);
nor NOR2 (N2878, N2866, N799);
and AND2 (N2879, N2875, N2550);
and AND4 (N2880, N2842, N2473, N1336, N473);
or OR2 (N2881, N2880, N2347);
buf BUF1 (N2882, N2867);
buf BUF1 (N2883, N2877);
buf BUF1 (N2884, N2868);
not NOT1 (N2885, N2860);
buf BUF1 (N2886, N2881);
nand NAND3 (N2887, N2879, N1224, N1076);
or OR4 (N2888, N2876, N2478, N2574, N276);
xor XOR2 (N2889, N2885, N1325);
nor NOR2 (N2890, N2873, N149);
or OR2 (N2891, N2889, N1858);
xor XOR2 (N2892, N2887, N339);
not NOT1 (N2893, N2892);
not NOT1 (N2894, N2882);
or OR4 (N2895, N2886, N620, N2027, N1089);
buf BUF1 (N2896, N2893);
or OR4 (N2897, N2890, N2510, N917, N1768);
not NOT1 (N2898, N2883);
nor NOR4 (N2899, N2897, N1344, N1569, N436);
nand NAND2 (N2900, N2870, N1011);
buf BUF1 (N2901, N2894);
or OR2 (N2902, N2884, N1093);
or OR4 (N2903, N2900, N2362, N1308, N1510);
nand NAND2 (N2904, N2901, N2533);
nand NAND4 (N2905, N2895, N491, N2115, N1332);
not NOT1 (N2906, N2902);
not NOT1 (N2907, N2899);
and AND2 (N2908, N2898, N1027);
nor NOR2 (N2909, N2908, N95);
not NOT1 (N2910, N2903);
nand NAND4 (N2911, N2905, N204, N2623, N858);
or OR2 (N2912, N2907, N364);
not NOT1 (N2913, N2878);
not NOT1 (N2914, N2904);
nor NOR3 (N2915, N2914, N2090, N496);
and AND3 (N2916, N2896, N956, N1073);
nor NOR3 (N2917, N2916, N2614, N1213);
not NOT1 (N2918, N2911);
buf BUF1 (N2919, N2906);
nand NAND3 (N2920, N2918, N2673, N530);
nor NOR4 (N2921, N2909, N1111, N2473, N2393);
xor XOR2 (N2922, N2910, N776);
nor NOR3 (N2923, N2917, N2301, N197);
buf BUF1 (N2924, N2912);
nand NAND3 (N2925, N2915, N520, N351);
buf BUF1 (N2926, N2922);
nor NOR4 (N2927, N2924, N1931, N2916, N2467);
nand NAND2 (N2928, N2891, N233);
nor NOR4 (N2929, N2888, N4, N211, N335);
nand NAND4 (N2930, N2929, N1727, N1388, N180);
and AND3 (N2931, N2930, N1952, N2398);
or OR3 (N2932, N2913, N141, N2421);
nand NAND3 (N2933, N2932, N1854, N1024);
buf BUF1 (N2934, N2919);
buf BUF1 (N2935, N2927);
not NOT1 (N2936, N2926);
and AND2 (N2937, N2935, N1126);
nand NAND2 (N2938, N2933, N1366);
not NOT1 (N2939, N2921);
xor XOR2 (N2940, N2937, N562);
buf BUF1 (N2941, N2931);
or OR4 (N2942, N2936, N1961, N2063, N837);
or OR2 (N2943, N2938, N1113);
buf BUF1 (N2944, N2928);
nor NOR4 (N2945, N2944, N1021, N2778, N323);
nand NAND4 (N2946, N2920, N1686, N2798, N2496);
xor XOR2 (N2947, N2941, N2944);
xor XOR2 (N2948, N2923, N2235);
and AND3 (N2949, N2947, N1112, N2853);
or OR4 (N2950, N2942, N146, N2466, N473);
xor XOR2 (N2951, N2949, N2140);
or OR3 (N2952, N2945, N1821, N1314);
nand NAND3 (N2953, N2925, N2931, N1005);
or OR3 (N2954, N2943, N1320, N307);
or OR4 (N2955, N2934, N339, N2525, N728);
nand NAND2 (N2956, N2951, N604);
nand NAND4 (N2957, N2954, N492, N1649, N2383);
nor NOR3 (N2958, N2956, N443, N1632);
xor XOR2 (N2959, N2955, N1231);
xor XOR2 (N2960, N2948, N1869);
and AND4 (N2961, N2960, N1491, N1213, N1707);
not NOT1 (N2962, N2952);
or OR4 (N2963, N2958, N744, N1648, N946);
not NOT1 (N2964, N2946);
buf BUF1 (N2965, N2959);
buf BUF1 (N2966, N2961);
xor XOR2 (N2967, N2950, N2697);
or OR3 (N2968, N2965, N1182, N641);
nor NOR3 (N2969, N2966, N2641, N934);
nor NOR2 (N2970, N2953, N66);
and AND3 (N2971, N2967, N1852, N2429);
not NOT1 (N2972, N2963);
buf BUF1 (N2973, N2962);
buf BUF1 (N2974, N2964);
xor XOR2 (N2975, N2973, N1001);
or OR2 (N2976, N2972, N2372);
not NOT1 (N2977, N2974);
or OR2 (N2978, N2969, N476);
nand NAND3 (N2979, N2968, N1580, N1122);
buf BUF1 (N2980, N2970);
nor NOR4 (N2981, N2979, N1607, N1886, N2400);
or OR2 (N2982, N2978, N807);
xor XOR2 (N2983, N2939, N490);
nand NAND3 (N2984, N2977, N2151, N2027);
and AND4 (N2985, N2983, N839, N1699, N308);
nor NOR3 (N2986, N2940, N1333, N2397);
or OR3 (N2987, N2976, N1315, N1137);
buf BUF1 (N2988, N2975);
buf BUF1 (N2989, N2957);
not NOT1 (N2990, N2981);
not NOT1 (N2991, N2987);
nand NAND2 (N2992, N2980, N2900);
buf BUF1 (N2993, N2989);
nand NAND4 (N2994, N2988, N2967, N2438, N1156);
not NOT1 (N2995, N2991);
nand NAND3 (N2996, N2992, N2292, N1701);
nand NAND2 (N2997, N2971, N1678);
nor NOR2 (N2998, N2994, N2907);
nor NOR3 (N2999, N2995, N1421, N2114);
or OR2 (N3000, N2985, N2940);
xor XOR2 (N3001, N2986, N1407);
buf BUF1 (N3002, N2984);
buf BUF1 (N3003, N2990);
and AND4 (N3004, N2997, N795, N365, N529);
nand NAND2 (N3005, N2993, N2328);
not NOT1 (N3006, N2996);
buf BUF1 (N3007, N2998);
or OR4 (N3008, N2999, N249, N1074, N30);
not NOT1 (N3009, N3004);
nand NAND4 (N3010, N3009, N302, N1209, N2186);
not NOT1 (N3011, N3000);
or OR4 (N3012, N3008, N1834, N2418, N594);
not NOT1 (N3013, N3011);
xor XOR2 (N3014, N3001, N1232);
xor XOR2 (N3015, N3014, N793);
xor XOR2 (N3016, N3013, N2909);
not NOT1 (N3017, N3006);
nor NOR2 (N3018, N2982, N1975);
xor XOR2 (N3019, N3017, N2581);
nand NAND3 (N3020, N3016, N2759, N1369);
buf BUF1 (N3021, N3012);
nor NOR4 (N3022, N3007, N2623, N673, N99);
nand NAND3 (N3023, N3003, N1678, N12);
or OR2 (N3024, N3022, N227);
nand NAND4 (N3025, N3019, N952, N2506, N1823);
xor XOR2 (N3026, N3002, N1441);
nor NOR2 (N3027, N3010, N853);
or OR3 (N3028, N3021, N375, N2973);
not NOT1 (N3029, N3028);
xor XOR2 (N3030, N3026, N2770);
or OR3 (N3031, N3023, N2130, N2715);
nor NOR3 (N3032, N3031, N1380, N1128);
nor NOR2 (N3033, N3005, N982);
or OR3 (N3034, N3032, N2556, N1607);
or OR3 (N3035, N3020, N2286, N1255);
buf BUF1 (N3036, N3018);
nor NOR4 (N3037, N3033, N2878, N1025, N2113);
and AND4 (N3038, N3024, N1579, N1746, N2318);
nor NOR4 (N3039, N3027, N2053, N1141, N700);
not NOT1 (N3040, N3039);
nor NOR2 (N3041, N3037, N1514);
nor NOR4 (N3042, N3029, N1570, N641, N1582);
not NOT1 (N3043, N3041);
buf BUF1 (N3044, N3036);
and AND3 (N3045, N3034, N2820, N232);
xor XOR2 (N3046, N3045, N2630);
and AND4 (N3047, N3042, N1979, N1899, N1767);
not NOT1 (N3048, N3040);
xor XOR2 (N3049, N3025, N645);
and AND2 (N3050, N3035, N557);
buf BUF1 (N3051, N3038);
and AND2 (N3052, N3051, N2347);
nor NOR3 (N3053, N3047, N3037, N1538);
not NOT1 (N3054, N3050);
and AND4 (N3055, N3030, N2081, N2716, N2291);
xor XOR2 (N3056, N3044, N2601);
xor XOR2 (N3057, N3055, N2580);
not NOT1 (N3058, N3053);
buf BUF1 (N3059, N3015);
nand NAND3 (N3060, N3046, N1870, N2351);
nor NOR3 (N3061, N3048, N962, N2689);
xor XOR2 (N3062, N3056, N2829);
xor XOR2 (N3063, N3061, N1124);
nand NAND4 (N3064, N3043, N1469, N1590, N360);
buf BUF1 (N3065, N3058);
and AND4 (N3066, N3060, N2961, N2957, N1423);
and AND4 (N3067, N3065, N1685, N2277, N693);
buf BUF1 (N3068, N3049);
or OR2 (N3069, N3063, N1868);
not NOT1 (N3070, N3069);
xor XOR2 (N3071, N3066, N2797);
and AND3 (N3072, N3057, N279, N2291);
nor NOR4 (N3073, N3054, N1957, N573, N2922);
or OR4 (N3074, N3070, N102, N349, N1227);
xor XOR2 (N3075, N3071, N260);
buf BUF1 (N3076, N3059);
buf BUF1 (N3077, N3073);
and AND4 (N3078, N3076, N2515, N1362, N402);
not NOT1 (N3079, N3067);
buf BUF1 (N3080, N3068);
not NOT1 (N3081, N3080);
buf BUF1 (N3082, N3072);
buf BUF1 (N3083, N3075);
buf BUF1 (N3084, N3064);
and AND2 (N3085, N3082, N157);
xor XOR2 (N3086, N3077, N88);
or OR2 (N3087, N3079, N1168);
xor XOR2 (N3088, N3085, N1706);
xor XOR2 (N3089, N3087, N1182);
buf BUF1 (N3090, N3086);
buf BUF1 (N3091, N3052);
xor XOR2 (N3092, N3083, N1517);
nor NOR3 (N3093, N3074, N1019, N772);
nand NAND4 (N3094, N3089, N799, N2136, N1001);
nor NOR4 (N3095, N3088, N2876, N1816, N1798);
or OR3 (N3096, N3091, N16, N1056);
buf BUF1 (N3097, N3062);
or OR2 (N3098, N3078, N1618);
nor NOR3 (N3099, N3090, N1684, N1454);
and AND3 (N3100, N3096, N1658, N2545);
buf BUF1 (N3101, N3092);
nor NOR3 (N3102, N3095, N978, N2850);
xor XOR2 (N3103, N3097, N773);
nor NOR3 (N3104, N3099, N2998, N2621);
xor XOR2 (N3105, N3103, N2312);
xor XOR2 (N3106, N3102, N927);
not NOT1 (N3107, N3093);
xor XOR2 (N3108, N3081, N1462);
xor XOR2 (N3109, N3098, N199);
and AND4 (N3110, N3105, N2561, N2676, N2107);
and AND3 (N3111, N3106, N2996, N2997);
xor XOR2 (N3112, N3104, N301);
xor XOR2 (N3113, N3094, N943);
buf BUF1 (N3114, N3100);
nor NOR2 (N3115, N3112, N1248);
and AND2 (N3116, N3115, N1241);
buf BUF1 (N3117, N3113);
or OR4 (N3118, N3111, N1415, N1239, N195);
nor NOR4 (N3119, N3114, N1040, N679, N1104);
nor NOR4 (N3120, N3110, N2547, N2600, N1540);
nand NAND2 (N3121, N3118, N853);
or OR3 (N3122, N3121, N1087, N2920);
and AND2 (N3123, N3108, N2777);
not NOT1 (N3124, N3107);
not NOT1 (N3125, N3120);
and AND2 (N3126, N3084, N2805);
not NOT1 (N3127, N3126);
buf BUF1 (N3128, N3124);
and AND3 (N3129, N3127, N2417, N3029);
nand NAND4 (N3130, N3129, N2135, N1998, N1689);
or OR4 (N3131, N3123, N2432, N2374, N1530);
nand NAND3 (N3132, N3128, N1013, N1342);
xor XOR2 (N3133, N3101, N3024);
buf BUF1 (N3134, N3132);
or OR4 (N3135, N3130, N720, N2432, N389);
and AND3 (N3136, N3119, N2682, N1704);
xor XOR2 (N3137, N3109, N2593);
or OR4 (N3138, N3134, N3011, N1968, N967);
buf BUF1 (N3139, N3138);
nor NOR4 (N3140, N3133, N2543, N1356, N998);
nor NOR2 (N3141, N3125, N3076);
nand NAND3 (N3142, N3135, N2772, N2075);
not NOT1 (N3143, N3141);
nor NOR4 (N3144, N3122, N1775, N199, N1509);
and AND4 (N3145, N3139, N1779, N2218, N2508);
or OR4 (N3146, N3131, N404, N2152, N2599);
not NOT1 (N3147, N3117);
xor XOR2 (N3148, N3116, N2025);
and AND3 (N3149, N3143, N2682, N2695);
not NOT1 (N3150, N3140);
nand NAND4 (N3151, N3146, N2884, N2765, N2256);
xor XOR2 (N3152, N3148, N2941);
and AND2 (N3153, N3136, N325);
and AND4 (N3154, N3153, N1254, N2707, N1552);
buf BUF1 (N3155, N3151);
not NOT1 (N3156, N3145);
buf BUF1 (N3157, N3149);
buf BUF1 (N3158, N3144);
or OR3 (N3159, N3158, N2850, N109);
and AND4 (N3160, N3150, N1060, N414, N2506);
and AND3 (N3161, N3160, N2093, N2875);
or OR2 (N3162, N3137, N701);
buf BUF1 (N3163, N3142);
nand NAND3 (N3164, N3152, N158, N1373);
not NOT1 (N3165, N3162);
nand NAND4 (N3166, N3156, N2034, N2842, N1549);
nand NAND3 (N3167, N3155, N507, N2163);
xor XOR2 (N3168, N3157, N1306);
nand NAND4 (N3169, N3164, N1076, N1480, N104);
xor XOR2 (N3170, N3167, N1975);
buf BUF1 (N3171, N3159);
nor NOR4 (N3172, N3165, N1733, N2691, N1721);
nand NAND2 (N3173, N3147, N2414);
buf BUF1 (N3174, N3166);
buf BUF1 (N3175, N3172);
xor XOR2 (N3176, N3161, N988);
and AND4 (N3177, N3168, N391, N1280, N2639);
or OR3 (N3178, N3170, N2670, N1057);
nor NOR2 (N3179, N3178, N606);
nand NAND3 (N3180, N3179, N417, N2861);
buf BUF1 (N3181, N3154);
not NOT1 (N3182, N3169);
or OR3 (N3183, N3182, N2125, N1999);
nand NAND3 (N3184, N3163, N328, N233);
xor XOR2 (N3185, N3175, N1698);
and AND4 (N3186, N3181, N1351, N611, N3083);
and AND2 (N3187, N3171, N3045);
buf BUF1 (N3188, N3184);
nand NAND4 (N3189, N3174, N2290, N2457, N2114);
nand NAND3 (N3190, N3177, N2612, N1116);
xor XOR2 (N3191, N3190, N2540);
buf BUF1 (N3192, N3189);
not NOT1 (N3193, N3191);
nor NOR2 (N3194, N3186, N3185);
nor NOR4 (N3195, N2656, N1816, N1226, N1035);
and AND4 (N3196, N3180, N1460, N567, N1298);
buf BUF1 (N3197, N3195);
xor XOR2 (N3198, N3176, N1643);
buf BUF1 (N3199, N3187);
nor NOR2 (N3200, N3197, N211);
nor NOR4 (N3201, N3199, N2296, N2042, N2414);
buf BUF1 (N3202, N3188);
nor NOR4 (N3203, N3200, N1985, N1598, N388);
nor NOR3 (N3204, N3193, N720, N852);
nand NAND2 (N3205, N3198, N2023);
and AND3 (N3206, N3203, N1972, N3183);
not NOT1 (N3207, N3062);
not NOT1 (N3208, N3192);
or OR2 (N3209, N3201, N1229);
nor NOR3 (N3210, N3194, N2809, N3111);
not NOT1 (N3211, N3204);
or OR3 (N3212, N3208, N2722, N955);
buf BUF1 (N3213, N3196);
nand NAND4 (N3214, N3211, N215, N1570, N2834);
and AND2 (N3215, N3214, N3030);
buf BUF1 (N3216, N3215);
or OR4 (N3217, N3216, N724, N1783, N1128);
not NOT1 (N3218, N3212);
nor NOR4 (N3219, N3210, N1951, N1726, N355);
not NOT1 (N3220, N3206);
xor XOR2 (N3221, N3202, N3107);
nand NAND2 (N3222, N3173, N2341);
xor XOR2 (N3223, N3207, N3123);
nand NAND3 (N3224, N3213, N1190, N1519);
nand NAND2 (N3225, N3218, N881);
not NOT1 (N3226, N3222);
not NOT1 (N3227, N3224);
not NOT1 (N3228, N3220);
nor NOR3 (N3229, N3209, N2475, N1990);
and AND3 (N3230, N3225, N868, N1127);
and AND2 (N3231, N3226, N1331);
nor NOR2 (N3232, N3219, N1250);
nand NAND2 (N3233, N3228, N345);
or OR3 (N3234, N3221, N1382, N3077);
not NOT1 (N3235, N3230);
not NOT1 (N3236, N3231);
not NOT1 (N3237, N3234);
not NOT1 (N3238, N3217);
nor NOR4 (N3239, N3238, N1239, N461, N3229);
and AND2 (N3240, N3123, N655);
nand NAND2 (N3241, N3236, N274);
nand NAND2 (N3242, N3233, N219);
not NOT1 (N3243, N3235);
not NOT1 (N3244, N3232);
nor NOR2 (N3245, N3243, N2614);
xor XOR2 (N3246, N3245, N1826);
xor XOR2 (N3247, N3242, N3006);
not NOT1 (N3248, N3241);
nand NAND4 (N3249, N3205, N2004, N290, N2342);
xor XOR2 (N3250, N3223, N936);
and AND4 (N3251, N3239, N675, N930, N376);
not NOT1 (N3252, N3251);
or OR4 (N3253, N3240, N2656, N1540, N375);
and AND4 (N3254, N3249, N2945, N3219, N2128);
nor NOR4 (N3255, N3252, N2477, N338, N2931);
buf BUF1 (N3256, N3250);
not NOT1 (N3257, N3244);
nand NAND2 (N3258, N3227, N617);
buf BUF1 (N3259, N3257);
and AND4 (N3260, N3258, N2326, N3139, N988);
or OR3 (N3261, N3255, N2935, N3055);
not NOT1 (N3262, N3260);
and AND3 (N3263, N3262, N1842, N1389);
not NOT1 (N3264, N3263);
and AND3 (N3265, N3264, N1691, N768);
nand NAND3 (N3266, N3261, N1446, N2453);
not NOT1 (N3267, N3246);
and AND3 (N3268, N3266, N606, N439);
buf BUF1 (N3269, N3253);
and AND3 (N3270, N3237, N1850, N1833);
nand NAND2 (N3271, N3267, N652);
buf BUF1 (N3272, N3270);
buf BUF1 (N3273, N3259);
or OR4 (N3274, N3265, N1362, N105, N2376);
and AND3 (N3275, N3256, N2065, N321);
buf BUF1 (N3276, N3247);
nor NOR2 (N3277, N3269, N900);
not NOT1 (N3278, N3272);
buf BUF1 (N3279, N3268);
or OR3 (N3280, N3254, N2445, N483);
buf BUF1 (N3281, N3278);
or OR3 (N3282, N3276, N1820, N315);
and AND4 (N3283, N3279, N386, N2496, N225);
nor NOR3 (N3284, N3277, N1729, N3244);
not NOT1 (N3285, N3248);
not NOT1 (N3286, N3285);
or OR3 (N3287, N3273, N2451, N3126);
not NOT1 (N3288, N3283);
and AND3 (N3289, N3286, N1060, N1351);
nand NAND4 (N3290, N3288, N736, N2696, N878);
nand NAND3 (N3291, N3287, N185, N1910);
or OR3 (N3292, N3271, N424, N254);
xor XOR2 (N3293, N3281, N2151);
xor XOR2 (N3294, N3275, N1642);
not NOT1 (N3295, N3293);
not NOT1 (N3296, N3294);
or OR3 (N3297, N3296, N799, N1596);
xor XOR2 (N3298, N3292, N1689);
nand NAND2 (N3299, N3284, N966);
nand NAND2 (N3300, N3282, N427);
and AND4 (N3301, N3299, N1846, N2025, N2294);
nand NAND4 (N3302, N3295, N1417, N3067, N470);
and AND2 (N3303, N3301, N1843);
xor XOR2 (N3304, N3291, N2059);
not NOT1 (N3305, N3280);
not NOT1 (N3306, N3302);
not NOT1 (N3307, N3304);
nand NAND2 (N3308, N3289, N3253);
and AND2 (N3309, N3306, N348);
and AND4 (N3310, N3307, N126, N1386, N1444);
or OR2 (N3311, N3274, N1374);
not NOT1 (N3312, N3308);
not NOT1 (N3313, N3300);
and AND2 (N3314, N3305, N1217);
or OR4 (N3315, N3303, N455, N3302, N2374);
buf BUF1 (N3316, N3314);
nor NOR2 (N3317, N3298, N2593);
buf BUF1 (N3318, N3315);
nand NAND4 (N3319, N3290, N3152, N765, N1591);
nand NAND2 (N3320, N3313, N403);
nor NOR2 (N3321, N3318, N2549);
nand NAND2 (N3322, N3312, N7);
and AND4 (N3323, N3310, N495, N1167, N1794);
buf BUF1 (N3324, N3319);
or OR2 (N3325, N3317, N367);
and AND4 (N3326, N3325, N3111, N3303, N1781);
nor NOR3 (N3327, N3297, N2343, N2090);
and AND3 (N3328, N3323, N273, N31);
nor NOR2 (N3329, N3322, N2688);
and AND2 (N3330, N3328, N2865);
xor XOR2 (N3331, N3316, N2699);
buf BUF1 (N3332, N3327);
and AND4 (N3333, N3311, N2875, N1035, N839);
and AND2 (N3334, N3330, N1960);
not NOT1 (N3335, N3333);
and AND3 (N3336, N3324, N643, N1628);
and AND3 (N3337, N3326, N1159, N988);
nand NAND4 (N3338, N3329, N2643, N1615, N623);
and AND2 (N3339, N3334, N1729);
buf BUF1 (N3340, N3320);
buf BUF1 (N3341, N3340);
not NOT1 (N3342, N3321);
or OR4 (N3343, N3337, N1884, N2302, N208);
buf BUF1 (N3344, N3309);
buf BUF1 (N3345, N3344);
nand NAND2 (N3346, N3336, N332);
or OR4 (N3347, N3331, N3159, N2166, N56);
and AND3 (N3348, N3342, N3252, N569);
xor XOR2 (N3349, N3345, N3312);
buf BUF1 (N3350, N3349);
nand NAND4 (N3351, N3348, N2887, N3172, N2620);
xor XOR2 (N3352, N3341, N1101);
nand NAND4 (N3353, N3343, N647, N408, N691);
xor XOR2 (N3354, N3332, N1066);
nand NAND2 (N3355, N3354, N2634);
xor XOR2 (N3356, N3355, N2235);
buf BUF1 (N3357, N3352);
or OR3 (N3358, N3339, N3320, N318);
and AND2 (N3359, N3353, N1298);
nand NAND4 (N3360, N3346, N630, N64, N694);
and AND2 (N3361, N3356, N961);
nor NOR3 (N3362, N3351, N2047, N1905);
and AND4 (N3363, N3359, N3138, N2805, N1442);
nand NAND4 (N3364, N3350, N2260, N494, N360);
and AND4 (N3365, N3347, N1278, N2301, N1687);
buf BUF1 (N3366, N3335);
not NOT1 (N3367, N3338);
nor NOR3 (N3368, N3363, N2214, N2802);
nand NAND3 (N3369, N3365, N1717, N3169);
or OR4 (N3370, N3358, N32, N1240, N2940);
and AND2 (N3371, N3362, N2791);
not NOT1 (N3372, N3364);
nor NOR3 (N3373, N3371, N3356, N2821);
nor NOR2 (N3374, N3357, N218);
buf BUF1 (N3375, N3373);
or OR3 (N3376, N3372, N3216, N386);
nand NAND2 (N3377, N3361, N2628);
nand NAND3 (N3378, N3369, N919, N153);
xor XOR2 (N3379, N3377, N3358);
and AND4 (N3380, N3366, N3377, N182, N3211);
not NOT1 (N3381, N3370);
nor NOR4 (N3382, N3381, N1395, N3330, N955);
xor XOR2 (N3383, N3367, N605);
or OR3 (N3384, N3376, N576, N999);
or OR4 (N3385, N3382, N1661, N132, N629);
nand NAND2 (N3386, N3379, N660);
not NOT1 (N3387, N3385);
or OR2 (N3388, N3387, N3049);
or OR4 (N3389, N3368, N2647, N1709, N123);
buf BUF1 (N3390, N3389);
not NOT1 (N3391, N3388);
xor XOR2 (N3392, N3375, N3141);
not NOT1 (N3393, N3360);
xor XOR2 (N3394, N3378, N1049);
xor XOR2 (N3395, N3392, N2263);
xor XOR2 (N3396, N3374, N1423);
or OR2 (N3397, N3394, N1360);
or OR3 (N3398, N3397, N213, N2699);
xor XOR2 (N3399, N3380, N1058);
and AND4 (N3400, N3393, N883, N2859, N1828);
and AND4 (N3401, N3384, N1149, N157, N515);
nand NAND3 (N3402, N3391, N2415, N441);
xor XOR2 (N3403, N3383, N1078);
and AND3 (N3404, N3403, N423, N3193);
or OR4 (N3405, N3404, N583, N2104, N1031);
not NOT1 (N3406, N3401);
and AND4 (N3407, N3402, N1998, N92, N609);
xor XOR2 (N3408, N3396, N529);
nand NAND4 (N3409, N3408, N2253, N2364, N2289);
nand NAND4 (N3410, N3395, N2174, N3049, N826);
or OR2 (N3411, N3399, N2877);
buf BUF1 (N3412, N3398);
xor XOR2 (N3413, N3386, N1760);
xor XOR2 (N3414, N3411, N2514);
nand NAND4 (N3415, N3405, N912, N2699, N1664);
nand NAND3 (N3416, N3410, N112, N2440);
xor XOR2 (N3417, N3414, N1543);
not NOT1 (N3418, N3415);
nand NAND3 (N3419, N3416, N310, N214);
and AND3 (N3420, N3400, N2484, N585);
nand NAND3 (N3421, N3406, N308, N1157);
nand NAND3 (N3422, N3390, N784, N28);
and AND2 (N3423, N3417, N2931);
nor NOR3 (N3424, N3418, N1907, N1008);
nor NOR3 (N3425, N3424, N2461, N2792);
xor XOR2 (N3426, N3422, N415);
or OR3 (N3427, N3409, N333, N181);
and AND2 (N3428, N3419, N1357);
buf BUF1 (N3429, N3423);
not NOT1 (N3430, N3407);
or OR2 (N3431, N3429, N1475);
not NOT1 (N3432, N3430);
xor XOR2 (N3433, N3431, N1934);
and AND2 (N3434, N3413, N891);
not NOT1 (N3435, N3433);
or OR3 (N3436, N3426, N1262, N871);
and AND4 (N3437, N3421, N2721, N1898, N1964);
or OR4 (N3438, N3425, N1271, N492, N1286);
nand NAND3 (N3439, N3436, N750, N1429);
not NOT1 (N3440, N3427);
xor XOR2 (N3441, N3440, N120);
xor XOR2 (N3442, N3441, N1208);
not NOT1 (N3443, N3435);
buf BUF1 (N3444, N3434);
xor XOR2 (N3445, N3438, N1611);
nor NOR2 (N3446, N3437, N2711);
or OR3 (N3447, N3432, N360, N979);
nor NOR4 (N3448, N3446, N1229, N2256, N3088);
buf BUF1 (N3449, N3445);
nand NAND3 (N3450, N3442, N2485, N2154);
nor NOR3 (N3451, N3448, N1928, N549);
or OR3 (N3452, N3443, N2753, N2739);
and AND3 (N3453, N3449, N2885, N1815);
buf BUF1 (N3454, N3444);
nand NAND2 (N3455, N3454, N1950);
buf BUF1 (N3456, N3439);
xor XOR2 (N3457, N3412, N408);
and AND2 (N3458, N3428, N3288);
or OR3 (N3459, N3455, N720, N130);
nand NAND4 (N3460, N3459, N1103, N1185, N135);
xor XOR2 (N3461, N3456, N1408);
or OR3 (N3462, N3452, N3160, N3106);
xor XOR2 (N3463, N3462, N2738);
or OR3 (N3464, N3451, N3364, N3224);
or OR3 (N3465, N3461, N363, N2933);
buf BUF1 (N3466, N3464);
xor XOR2 (N3467, N3466, N495);
xor XOR2 (N3468, N3458, N1583);
nor NOR2 (N3469, N3463, N1617);
nor NOR4 (N3470, N3469, N2399, N1716, N20);
nand NAND2 (N3471, N3470, N628);
and AND3 (N3472, N3450, N2246, N491);
xor XOR2 (N3473, N3467, N1027);
xor XOR2 (N3474, N3471, N1785);
or OR4 (N3475, N3474, N445, N1798, N1208);
nand NAND3 (N3476, N3457, N1717, N2279);
nor NOR4 (N3477, N3473, N562, N2788, N1192);
or OR4 (N3478, N3468, N2872, N604, N2099);
nand NAND4 (N3479, N3460, N929, N1924, N20);
and AND2 (N3480, N3420, N1704);
not NOT1 (N3481, N3447);
nand NAND2 (N3482, N3465, N287);
or OR4 (N3483, N3478, N2267, N3314, N3250);
xor XOR2 (N3484, N3477, N510);
nand NAND3 (N3485, N3472, N2651, N2230);
buf BUF1 (N3486, N3476);
not NOT1 (N3487, N3485);
buf BUF1 (N3488, N3487);
xor XOR2 (N3489, N3486, N2493);
buf BUF1 (N3490, N3488);
and AND4 (N3491, N3484, N379, N2953, N821);
nor NOR2 (N3492, N3481, N2794);
buf BUF1 (N3493, N3482);
not NOT1 (N3494, N3492);
not NOT1 (N3495, N3489);
nand NAND3 (N3496, N3453, N986, N3432);
not NOT1 (N3497, N3490);
not NOT1 (N3498, N3497);
nand NAND2 (N3499, N3479, N270);
xor XOR2 (N3500, N3494, N2733);
or OR4 (N3501, N3495, N2833, N2939, N1018);
not NOT1 (N3502, N3499);
not NOT1 (N3503, N3500);
or OR2 (N3504, N3502, N1250);
not NOT1 (N3505, N3493);
or OR2 (N3506, N3475, N58);
buf BUF1 (N3507, N3501);
buf BUF1 (N3508, N3506);
xor XOR2 (N3509, N3480, N2297);
and AND3 (N3510, N3498, N262, N2650);
buf BUF1 (N3511, N3505);
or OR3 (N3512, N3511, N1333, N1898);
endmodule