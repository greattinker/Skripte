// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N8004,N8005,N7992,N8008,N7988,N8013,N8011,N8010,N8012,N8014;

nand NAND3 (N15, N1, N12, N9);
nor NOR2 (N16, N11, N12);
not NOT1 (N17, N6);
and AND2 (N18, N10, N9);
nand NAND2 (N19, N16, N6);
xor XOR2 (N20, N10, N10);
nand NAND2 (N21, N4, N14);
or OR4 (N22, N21, N3, N16, N19);
buf BUF1 (N23, N6);
not NOT1 (N24, N17);
and AND2 (N25, N10, N17);
nor NOR4 (N26, N25, N3, N15, N25);
nand NAND4 (N27, N3, N6, N18, N2);
nor NOR2 (N28, N6, N1);
nand NAND4 (N29, N16, N13, N14, N11);
buf BUF1 (N30, N6);
xor XOR2 (N31, N1, N3);
and AND4 (N32, N27, N19, N29, N21);
or OR2 (N33, N2, N10);
and AND2 (N34, N24, N32);
or OR3 (N35, N26, N17, N27);
nor NOR3 (N36, N16, N26, N20);
and AND3 (N37, N6, N24, N31);
or OR4 (N38, N23, N4, N20, N28);
nand NAND2 (N39, N16, N29);
or OR4 (N40, N1, N37, N7, N33);
buf BUF1 (N41, N39);
and AND4 (N42, N16, N25, N35, N9);
or OR4 (N43, N28, N30, N19, N6);
not NOT1 (N44, N9);
nand NAND2 (N45, N1, N19);
nor NOR3 (N46, N34, N14, N45);
or OR2 (N47, N2, N42);
nor NOR2 (N48, N36, N45);
or OR2 (N49, N7, N28);
nor NOR2 (N50, N43, N25);
or OR2 (N51, N47, N6);
nand NAND4 (N52, N38, N6, N13, N42);
and AND3 (N53, N40, N43, N3);
buf BUF1 (N54, N22);
and AND3 (N55, N48, N4, N23);
and AND3 (N56, N49, N11, N13);
or OR2 (N57, N46, N38);
nor NOR4 (N58, N50, N3, N38, N20);
or OR3 (N59, N44, N51, N45);
and AND4 (N60, N6, N37, N4, N58);
or OR2 (N61, N45, N37);
buf BUF1 (N62, N55);
or OR3 (N63, N54, N52, N40);
buf BUF1 (N64, N28);
and AND4 (N65, N59, N9, N20, N47);
xor XOR2 (N66, N61, N49);
or OR4 (N67, N41, N60, N59, N41);
xor XOR2 (N68, N29, N57);
not NOT1 (N69, N39);
nand NAND2 (N70, N69, N57);
nor NOR3 (N71, N64, N32, N46);
xor XOR2 (N72, N67, N41);
buf BUF1 (N73, N72);
or OR4 (N74, N53, N20, N63, N27);
nand NAND3 (N75, N54, N24, N3);
not NOT1 (N76, N68);
not NOT1 (N77, N70);
not NOT1 (N78, N74);
nand NAND2 (N79, N78, N2);
xor XOR2 (N80, N79, N13);
xor XOR2 (N81, N73, N43);
nor NOR3 (N82, N65, N29, N68);
or OR4 (N83, N77, N15, N3, N21);
or OR2 (N84, N56, N76);
buf BUF1 (N85, N29);
and AND4 (N86, N71, N55, N83, N82);
or OR2 (N87, N52, N45);
xor XOR2 (N88, N71, N8);
nor NOR2 (N89, N88, N23);
nor NOR3 (N90, N86, N3, N44);
and AND3 (N91, N85, N6, N77);
or OR3 (N92, N84, N19, N81);
not NOT1 (N93, N13);
nor NOR2 (N94, N75, N62);
or OR4 (N95, N32, N30, N89, N43);
buf BUF1 (N96, N93);
nand NAND3 (N97, N35, N93, N74);
nor NOR4 (N98, N91, N87, N85, N55);
xor XOR2 (N99, N10, N11);
buf BUF1 (N100, N94);
nand NAND2 (N101, N98, N11);
and AND4 (N102, N96, N87, N77, N54);
nand NAND2 (N103, N66, N18);
and AND4 (N104, N101, N53, N37, N73);
nand NAND4 (N105, N80, N10, N94, N90);
xor XOR2 (N106, N76, N82);
buf BUF1 (N107, N95);
not NOT1 (N108, N99);
buf BUF1 (N109, N105);
and AND3 (N110, N102, N81, N95);
nor NOR2 (N111, N109, N16);
and AND3 (N112, N97, N30, N81);
and AND3 (N113, N104, N11, N39);
xor XOR2 (N114, N92, N10);
nand NAND2 (N115, N103, N26);
xor XOR2 (N116, N113, N91);
not NOT1 (N117, N111);
or OR4 (N118, N108, N55, N71, N3);
xor XOR2 (N119, N115, N57);
nand NAND4 (N120, N112, N65, N108, N100);
nand NAND4 (N121, N106, N68, N117, N29);
not NOT1 (N122, N4);
and AND4 (N123, N28, N101, N9, N67);
nand NAND2 (N124, N120, N40);
not NOT1 (N125, N124);
buf BUF1 (N126, N125);
and AND3 (N127, N118, N28, N92);
or OR3 (N128, N119, N118, N77);
not NOT1 (N129, N122);
nor NOR3 (N130, N129, N35, N82);
nor NOR2 (N131, N110, N93);
and AND4 (N132, N121, N37, N64, N129);
nand NAND2 (N133, N130, N60);
and AND3 (N134, N132, N32, N57);
and AND2 (N135, N133, N53);
nor NOR4 (N136, N107, N125, N70, N66);
buf BUF1 (N137, N134);
buf BUF1 (N138, N135);
not NOT1 (N139, N137);
or OR4 (N140, N116, N17, N38, N64);
or OR2 (N141, N138, N12);
not NOT1 (N142, N127);
buf BUF1 (N143, N136);
nand NAND2 (N144, N126, N44);
xor XOR2 (N145, N141, N31);
xor XOR2 (N146, N128, N134);
or OR4 (N147, N131, N86, N109, N117);
and AND3 (N148, N114, N40, N131);
nand NAND2 (N149, N143, N121);
not NOT1 (N150, N149);
or OR4 (N151, N150, N139, N45, N60);
and AND4 (N152, N2, N29, N20, N5);
or OR4 (N153, N147, N100, N114, N77);
buf BUF1 (N154, N145);
not NOT1 (N155, N152);
buf BUF1 (N156, N142);
and AND3 (N157, N151, N74, N71);
nand NAND3 (N158, N156, N143, N39);
or OR4 (N159, N148, N17, N4, N86);
buf BUF1 (N160, N123);
nand NAND4 (N161, N157, N125, N134, N88);
buf BUF1 (N162, N144);
buf BUF1 (N163, N153);
not NOT1 (N164, N162);
or OR3 (N165, N161, N133, N20);
not NOT1 (N166, N165);
and AND2 (N167, N166, N60);
nor NOR4 (N168, N163, N22, N153, N33);
nand NAND3 (N169, N168, N109, N6);
xor XOR2 (N170, N169, N36);
xor XOR2 (N171, N146, N73);
nand NAND4 (N172, N160, N163, N138, N126);
buf BUF1 (N173, N171);
buf BUF1 (N174, N159);
or OR3 (N175, N155, N79, N131);
nand NAND3 (N176, N173, N17, N88);
and AND2 (N177, N140, N173);
buf BUF1 (N178, N158);
nand NAND3 (N179, N174, N134, N155);
nor NOR2 (N180, N172, N129);
and AND4 (N181, N176, N178, N96, N85);
buf BUF1 (N182, N151);
nand NAND2 (N183, N182, N39);
nor NOR2 (N184, N167, N94);
or OR2 (N185, N177, N11);
and AND3 (N186, N175, N93, N65);
nor NOR4 (N187, N185, N169, N140, N80);
nand NAND2 (N188, N186, N110);
nor NOR2 (N189, N181, N132);
or OR4 (N190, N180, N20, N86, N1);
buf BUF1 (N191, N187);
nand NAND2 (N192, N190, N70);
not NOT1 (N193, N170);
xor XOR2 (N194, N192, N31);
not NOT1 (N195, N154);
not NOT1 (N196, N183);
xor XOR2 (N197, N179, N108);
or OR2 (N198, N196, N74);
buf BUF1 (N199, N191);
nor NOR4 (N200, N197, N26, N133, N104);
xor XOR2 (N201, N193, N105);
not NOT1 (N202, N198);
not NOT1 (N203, N184);
buf BUF1 (N204, N164);
nor NOR4 (N205, N203, N123, N202, N155);
not NOT1 (N206, N121);
buf BUF1 (N207, N200);
buf BUF1 (N208, N207);
not NOT1 (N209, N206);
not NOT1 (N210, N205);
and AND3 (N211, N208, N151, N61);
xor XOR2 (N212, N209, N115);
or OR4 (N213, N211, N47, N166, N32);
or OR3 (N214, N204, N39, N77);
and AND3 (N215, N213, N179, N90);
or OR2 (N216, N194, N120);
xor XOR2 (N217, N189, N171);
buf BUF1 (N218, N214);
xor XOR2 (N219, N212, N36);
nor NOR3 (N220, N199, N120, N162);
nor NOR4 (N221, N220, N113, N140, N107);
nor NOR3 (N222, N218, N198, N81);
nor NOR4 (N223, N221, N132, N16, N131);
not NOT1 (N224, N195);
and AND2 (N225, N222, N138);
and AND2 (N226, N210, N60);
or OR3 (N227, N226, N219, N150);
not NOT1 (N228, N134);
xor XOR2 (N229, N227, N172);
xor XOR2 (N230, N201, N190);
buf BUF1 (N231, N216);
not NOT1 (N232, N230);
or OR3 (N233, N229, N169, N110);
buf BUF1 (N234, N228);
and AND4 (N235, N231, N121, N229, N120);
nor NOR3 (N236, N188, N234, N181);
nand NAND3 (N237, N142, N165, N167);
buf BUF1 (N238, N225);
xor XOR2 (N239, N236, N199);
nand NAND4 (N240, N223, N115, N209, N154);
not NOT1 (N241, N217);
nor NOR2 (N242, N239, N44);
xor XOR2 (N243, N235, N202);
and AND4 (N244, N238, N112, N36, N119);
or OR4 (N245, N224, N214, N16, N146);
nand NAND2 (N246, N241, N97);
nor NOR2 (N247, N232, N181);
not NOT1 (N248, N215);
nor NOR3 (N249, N246, N62, N216);
xor XOR2 (N250, N244, N234);
and AND4 (N251, N237, N242, N166, N81);
nor NOR3 (N252, N157, N157, N161);
not NOT1 (N253, N248);
or OR4 (N254, N249, N236, N150, N59);
or OR4 (N255, N245, N134, N52, N169);
buf BUF1 (N256, N253);
nor NOR3 (N257, N247, N6, N31);
and AND2 (N258, N251, N223);
nor NOR3 (N259, N243, N85, N24);
nor NOR4 (N260, N256, N209, N102, N108);
buf BUF1 (N261, N254);
nand NAND2 (N262, N252, N218);
not NOT1 (N263, N258);
and AND2 (N264, N255, N135);
and AND2 (N265, N264, N150);
and AND2 (N266, N261, N130);
nor NOR3 (N267, N266, N22, N27);
nor NOR2 (N268, N262, N90);
nor NOR2 (N269, N257, N209);
xor XOR2 (N270, N260, N39);
nor NOR4 (N271, N267, N186, N94, N81);
buf BUF1 (N272, N259);
and AND2 (N273, N263, N126);
buf BUF1 (N274, N265);
or OR3 (N275, N233, N181, N157);
nor NOR2 (N276, N250, N115);
and AND4 (N277, N270, N114, N164, N87);
xor XOR2 (N278, N268, N66);
xor XOR2 (N279, N272, N166);
and AND4 (N280, N271, N98, N12, N56);
not NOT1 (N281, N240);
nand NAND2 (N282, N273, N71);
xor XOR2 (N283, N280, N273);
nor NOR2 (N284, N282, N240);
nor NOR4 (N285, N276, N211, N137, N85);
buf BUF1 (N286, N269);
and AND4 (N287, N274, N164, N249, N130);
or OR4 (N288, N283, N134, N1, N244);
nand NAND4 (N289, N287, N91, N227, N260);
nor NOR4 (N290, N275, N266, N205, N164);
buf BUF1 (N291, N288);
nor NOR4 (N292, N281, N25, N194, N45);
or OR4 (N293, N286, N103, N86, N249);
buf BUF1 (N294, N278);
xor XOR2 (N295, N292, N38);
xor XOR2 (N296, N291, N141);
and AND2 (N297, N289, N207);
buf BUF1 (N298, N285);
nor NOR4 (N299, N295, N206, N147, N189);
buf BUF1 (N300, N293);
and AND4 (N301, N294, N94, N168, N51);
nand NAND4 (N302, N284, N93, N295, N83);
nand NAND2 (N303, N298, N82);
and AND3 (N304, N296, N8, N113);
nor NOR3 (N305, N300, N235, N199);
not NOT1 (N306, N277);
nor NOR4 (N307, N297, N184, N149, N183);
buf BUF1 (N308, N290);
buf BUF1 (N309, N305);
nand NAND4 (N310, N306, N260, N172, N284);
and AND4 (N311, N309, N79, N112, N178);
or OR3 (N312, N304, N173, N151);
not NOT1 (N313, N279);
nor NOR2 (N314, N311, N74);
not NOT1 (N315, N310);
nor NOR2 (N316, N299, N144);
nor NOR4 (N317, N307, N178, N51, N202);
or OR2 (N318, N313, N116);
buf BUF1 (N319, N314);
or OR4 (N320, N318, N226, N157, N58);
or OR3 (N321, N308, N130, N152);
nand NAND3 (N322, N301, N201, N187);
and AND3 (N323, N303, N181, N83);
or OR2 (N324, N312, N256);
nor NOR3 (N325, N319, N278, N7);
or OR3 (N326, N323, N16, N209);
or OR2 (N327, N322, N27);
and AND2 (N328, N317, N26);
xor XOR2 (N329, N328, N89);
nor NOR2 (N330, N316, N273);
not NOT1 (N331, N326);
xor XOR2 (N332, N330, N20);
nand NAND3 (N333, N329, N181, N199);
or OR2 (N334, N321, N27);
buf BUF1 (N335, N320);
or OR3 (N336, N325, N118, N181);
nand NAND3 (N337, N327, N291, N98);
or OR3 (N338, N335, N150, N305);
or OR3 (N339, N331, N5, N305);
and AND2 (N340, N332, N186);
xor XOR2 (N341, N324, N140);
not NOT1 (N342, N333);
or OR4 (N343, N337, N64, N58, N232);
or OR4 (N344, N302, N325, N290, N245);
or OR3 (N345, N342, N103, N89);
and AND3 (N346, N334, N315, N32);
buf BUF1 (N347, N57);
or OR4 (N348, N341, N91, N199, N187);
nor NOR3 (N349, N339, N303, N130);
nor NOR4 (N350, N347, N164, N207, N304);
or OR4 (N351, N350, N320, N78, N28);
not NOT1 (N352, N344);
or OR2 (N353, N351, N16);
and AND4 (N354, N343, N289, N253, N70);
xor XOR2 (N355, N345, N231);
not NOT1 (N356, N346);
not NOT1 (N357, N352);
nand NAND2 (N358, N354, N90);
and AND3 (N359, N336, N342, N1);
buf BUF1 (N360, N338);
or OR4 (N361, N360, N248, N209, N292);
not NOT1 (N362, N361);
nand NAND3 (N363, N357, N126, N192);
or OR3 (N364, N356, N214, N184);
buf BUF1 (N365, N362);
xor XOR2 (N366, N364, N252);
or OR4 (N367, N358, N225, N102, N357);
not NOT1 (N368, N348);
nand NAND2 (N369, N353, N290);
or OR3 (N370, N349, N252, N206);
not NOT1 (N371, N340);
xor XOR2 (N372, N370, N219);
buf BUF1 (N373, N365);
nand NAND3 (N374, N372, N310, N335);
xor XOR2 (N375, N371, N294);
and AND2 (N376, N374, N129);
buf BUF1 (N377, N359);
not NOT1 (N378, N355);
nor NOR4 (N379, N378, N136, N353, N117);
nor NOR3 (N380, N369, N378, N223);
buf BUF1 (N381, N379);
nor NOR4 (N382, N363, N106, N267, N343);
xor XOR2 (N383, N366, N178);
nand NAND4 (N384, N375, N142, N187, N75);
xor XOR2 (N385, N380, N51);
nor NOR3 (N386, N381, N174, N255);
not NOT1 (N387, N367);
and AND3 (N388, N384, N387, N65);
not NOT1 (N389, N325);
and AND2 (N390, N388, N178);
not NOT1 (N391, N376);
not NOT1 (N392, N390);
buf BUF1 (N393, N382);
or OR4 (N394, N393, N88, N183, N303);
nand NAND3 (N395, N386, N87, N3);
nor NOR2 (N396, N373, N119);
xor XOR2 (N397, N391, N66);
and AND4 (N398, N395, N239, N365, N20);
nor NOR4 (N399, N383, N30, N5, N305);
xor XOR2 (N400, N377, N191);
not NOT1 (N401, N398);
and AND3 (N402, N396, N99, N342);
nand NAND3 (N403, N397, N163, N84);
or OR2 (N404, N368, N64);
buf BUF1 (N405, N402);
nor NOR4 (N406, N389, N80, N117, N14);
xor XOR2 (N407, N405, N171);
and AND2 (N408, N400, N2);
buf BUF1 (N409, N407);
nand NAND4 (N410, N401, N172, N309, N318);
not NOT1 (N411, N385);
nor NOR2 (N412, N410, N88);
not NOT1 (N413, N408);
or OR2 (N414, N392, N401);
buf BUF1 (N415, N412);
or OR4 (N416, N415, N405, N22, N264);
buf BUF1 (N417, N413);
xor XOR2 (N418, N417, N12);
not NOT1 (N419, N409);
or OR3 (N420, N406, N305, N316);
buf BUF1 (N421, N394);
buf BUF1 (N422, N421);
buf BUF1 (N423, N414);
nor NOR2 (N424, N419, N347);
xor XOR2 (N425, N403, N320);
xor XOR2 (N426, N399, N350);
or OR4 (N427, N411, N193, N248, N345);
and AND3 (N428, N404, N395, N365);
not NOT1 (N429, N426);
buf BUF1 (N430, N418);
nor NOR3 (N431, N429, N87, N62);
nand NAND3 (N432, N416, N101, N377);
and AND2 (N433, N425, N319);
nand NAND2 (N434, N431, N404);
nor NOR2 (N435, N430, N318);
and AND3 (N436, N422, N14, N23);
or OR3 (N437, N433, N16, N282);
or OR4 (N438, N420, N131, N328, N293);
nor NOR3 (N439, N428, N261, N25);
nand NAND3 (N440, N435, N181, N246);
nor NOR2 (N441, N427, N332);
xor XOR2 (N442, N437, N162);
not NOT1 (N443, N424);
nor NOR2 (N444, N440, N155);
xor XOR2 (N445, N436, N292);
or OR2 (N446, N439, N22);
nand NAND4 (N447, N444, N291, N65, N80);
buf BUF1 (N448, N423);
or OR2 (N449, N445, N185);
nor NOR3 (N450, N432, N448, N74);
xor XOR2 (N451, N40, N288);
nand NAND3 (N452, N442, N71, N424);
xor XOR2 (N453, N450, N318);
or OR2 (N454, N443, N193);
nor NOR3 (N455, N451, N155, N448);
nand NAND2 (N456, N453, N40);
nor NOR2 (N457, N447, N74);
nor NOR4 (N458, N449, N233, N163, N336);
xor XOR2 (N459, N446, N106);
or OR3 (N460, N459, N148, N92);
nor NOR2 (N461, N458, N226);
and AND3 (N462, N434, N161, N361);
nand NAND2 (N463, N461, N70);
buf BUF1 (N464, N463);
xor XOR2 (N465, N456, N408);
nand NAND4 (N466, N457, N335, N333, N164);
or OR3 (N467, N438, N376, N202);
nand NAND2 (N468, N462, N28);
and AND2 (N469, N465, N318);
buf BUF1 (N470, N452);
buf BUF1 (N471, N464);
and AND3 (N472, N454, N438, N217);
nand NAND4 (N473, N466, N349, N251, N8);
or OR3 (N474, N467, N32, N291);
xor XOR2 (N475, N473, N68);
and AND2 (N476, N469, N414);
or OR2 (N477, N441, N332);
nand NAND2 (N478, N474, N172);
and AND3 (N479, N476, N218, N304);
nand NAND3 (N480, N472, N235, N364);
not NOT1 (N481, N478);
not NOT1 (N482, N475);
nor NOR3 (N483, N468, N74, N104);
or OR4 (N484, N455, N199, N76, N114);
buf BUF1 (N485, N471);
xor XOR2 (N486, N481, N279);
buf BUF1 (N487, N477);
nand NAND3 (N488, N484, N386, N14);
and AND4 (N489, N460, N194, N276, N36);
xor XOR2 (N490, N487, N116);
and AND4 (N491, N489, N368, N68, N311);
and AND3 (N492, N485, N459, N366);
and AND3 (N493, N470, N383, N141);
buf BUF1 (N494, N482);
nand NAND4 (N495, N479, N337, N55, N414);
nor NOR2 (N496, N483, N294);
nor NOR2 (N497, N480, N29);
nor NOR4 (N498, N491, N305, N394, N441);
or OR2 (N499, N486, N20);
nand NAND3 (N500, N494, N257, N407);
xor XOR2 (N501, N500, N468);
and AND4 (N502, N497, N449, N348, N200);
buf BUF1 (N503, N495);
nand NAND4 (N504, N493, N272, N77, N177);
nor NOR4 (N505, N496, N434, N328, N51);
not NOT1 (N506, N499);
nand NAND2 (N507, N498, N6);
or OR2 (N508, N503, N507);
nand NAND4 (N509, N195, N394, N493, N42);
nor NOR4 (N510, N506, N439, N382, N92);
xor XOR2 (N511, N504, N323);
nor NOR3 (N512, N505, N391, N88);
xor XOR2 (N513, N502, N240);
and AND4 (N514, N509, N347, N208, N259);
or OR4 (N515, N488, N249, N496, N27);
buf BUF1 (N516, N492);
and AND2 (N517, N514, N24);
nor NOR4 (N518, N511, N209, N25, N424);
or OR2 (N519, N515, N146);
nor NOR2 (N520, N512, N178);
buf BUF1 (N521, N510);
not NOT1 (N522, N518);
xor XOR2 (N523, N490, N513);
nand NAND3 (N524, N104, N164, N115);
xor XOR2 (N525, N521, N226);
xor XOR2 (N526, N525, N433);
and AND4 (N527, N520, N166, N25, N225);
xor XOR2 (N528, N524, N448);
buf BUF1 (N529, N508);
and AND4 (N530, N528, N466, N222, N23);
and AND3 (N531, N527, N30, N9);
or OR3 (N532, N501, N131, N514);
nor NOR4 (N533, N526, N232, N206, N508);
buf BUF1 (N534, N532);
and AND3 (N535, N533, N474, N525);
buf BUF1 (N536, N531);
buf BUF1 (N537, N535);
nand NAND2 (N538, N536, N426);
or OR3 (N539, N517, N87, N394);
and AND4 (N540, N530, N231, N519, N432);
nor NOR3 (N541, N229, N400, N66);
xor XOR2 (N542, N537, N441);
not NOT1 (N543, N523);
nand NAND3 (N544, N516, N203, N245);
and AND3 (N545, N529, N197, N98);
not NOT1 (N546, N540);
or OR3 (N547, N546, N4, N418);
nor NOR4 (N548, N544, N320, N308, N547);
not NOT1 (N549, N330);
nor NOR3 (N550, N522, N218, N235);
nor NOR4 (N551, N549, N206, N274, N336);
xor XOR2 (N552, N543, N395);
xor XOR2 (N553, N548, N471);
buf BUF1 (N554, N550);
not NOT1 (N555, N534);
or OR4 (N556, N553, N127, N154, N373);
nor NOR4 (N557, N556, N523, N554, N306);
nor NOR3 (N558, N209, N151, N49);
or OR4 (N559, N558, N463, N425, N177);
not NOT1 (N560, N538);
and AND2 (N561, N559, N443);
not NOT1 (N562, N551);
buf BUF1 (N563, N561);
or OR4 (N564, N562, N303, N376, N220);
or OR3 (N565, N560, N385, N407);
or OR4 (N566, N541, N189, N279, N397);
or OR3 (N567, N564, N433, N409);
not NOT1 (N568, N545);
xor XOR2 (N569, N563, N38);
nor NOR2 (N570, N557, N153);
and AND4 (N571, N539, N426, N116, N59);
nor NOR3 (N572, N570, N287, N67);
nor NOR3 (N573, N572, N136, N260);
buf BUF1 (N574, N555);
buf BUF1 (N575, N542);
buf BUF1 (N576, N571);
xor XOR2 (N577, N575, N543);
buf BUF1 (N578, N573);
and AND2 (N579, N577, N339);
not NOT1 (N580, N566);
and AND2 (N581, N565, N230);
nor NOR4 (N582, N581, N555, N193, N485);
buf BUF1 (N583, N567);
not NOT1 (N584, N576);
not NOT1 (N585, N552);
or OR3 (N586, N584, N217, N34);
nor NOR4 (N587, N578, N574, N402, N390);
xor XOR2 (N588, N340, N122);
or OR4 (N589, N582, N519, N44, N444);
or OR4 (N590, N569, N285, N518, N562);
nor NOR4 (N591, N568, N87, N206, N308);
xor XOR2 (N592, N583, N497);
and AND4 (N593, N586, N251, N499, N185);
xor XOR2 (N594, N580, N481);
or OR2 (N595, N588, N350);
and AND4 (N596, N587, N60, N440, N554);
not NOT1 (N597, N579);
not NOT1 (N598, N596);
or OR4 (N599, N585, N116, N223, N128);
nor NOR4 (N600, N590, N509, N326, N132);
and AND4 (N601, N594, N187, N409, N132);
not NOT1 (N602, N595);
nand NAND3 (N603, N593, N483, N244);
or OR4 (N604, N600, N583, N295, N315);
or OR4 (N605, N599, N130, N370, N244);
nand NAND2 (N606, N592, N484);
nor NOR3 (N607, N598, N410, N149);
xor XOR2 (N608, N605, N603);
not NOT1 (N609, N109);
buf BUF1 (N610, N597);
not NOT1 (N611, N609);
buf BUF1 (N612, N611);
nor NOR4 (N613, N608, N297, N389, N488);
and AND3 (N614, N589, N390, N354);
xor XOR2 (N615, N607, N125);
nand NAND3 (N616, N612, N26, N294);
xor XOR2 (N617, N604, N439);
buf BUF1 (N618, N614);
nor NOR4 (N619, N606, N509, N21, N275);
not NOT1 (N620, N613);
not NOT1 (N621, N619);
or OR2 (N622, N616, N369);
nand NAND4 (N623, N618, N599, N102, N131);
nor NOR4 (N624, N623, N202, N431, N552);
not NOT1 (N625, N624);
not NOT1 (N626, N620);
buf BUF1 (N627, N591);
nand NAND3 (N628, N625, N375, N179);
nor NOR4 (N629, N627, N350, N349, N497);
buf BUF1 (N630, N622);
and AND3 (N631, N630, N628, N120);
not NOT1 (N632, N152);
nor NOR4 (N633, N626, N15, N588, N406);
xor XOR2 (N634, N615, N133);
nand NAND4 (N635, N633, N422, N333, N426);
xor XOR2 (N636, N634, N612);
not NOT1 (N637, N610);
buf BUF1 (N638, N631);
xor XOR2 (N639, N635, N372);
or OR3 (N640, N617, N181, N44);
nand NAND3 (N641, N638, N30, N248);
buf BUF1 (N642, N637);
not NOT1 (N643, N601);
and AND4 (N644, N642, N259, N137, N597);
nand NAND4 (N645, N636, N210, N140, N629);
or OR3 (N646, N312, N512, N30);
or OR2 (N647, N646, N470);
or OR4 (N648, N647, N94, N349, N565);
nand NAND3 (N649, N648, N71, N17);
not NOT1 (N650, N632);
nor NOR4 (N651, N639, N480, N522, N305);
not NOT1 (N652, N641);
nor NOR4 (N653, N645, N134, N636, N97);
nor NOR2 (N654, N653, N566);
and AND2 (N655, N640, N132);
and AND3 (N656, N649, N308, N529);
or OR4 (N657, N654, N377, N140, N494);
or OR2 (N658, N652, N99);
not NOT1 (N659, N651);
xor XOR2 (N660, N602, N552);
nor NOR3 (N661, N643, N176, N572);
xor XOR2 (N662, N650, N537);
and AND4 (N663, N657, N541, N330, N205);
xor XOR2 (N664, N660, N236);
buf BUF1 (N665, N663);
xor XOR2 (N666, N659, N636);
not NOT1 (N667, N656);
and AND2 (N668, N664, N116);
xor XOR2 (N669, N665, N612);
or OR2 (N670, N658, N372);
not NOT1 (N671, N667);
not NOT1 (N672, N621);
nor NOR4 (N673, N655, N16, N566, N136);
or OR4 (N674, N673, N217, N642, N252);
nor NOR2 (N675, N666, N67);
not NOT1 (N676, N670);
not NOT1 (N677, N676);
not NOT1 (N678, N672);
not NOT1 (N679, N671);
buf BUF1 (N680, N674);
or OR4 (N681, N675, N482, N490, N479);
or OR2 (N682, N661, N607);
nor NOR3 (N683, N677, N128, N166);
not NOT1 (N684, N679);
xor XOR2 (N685, N684, N108);
buf BUF1 (N686, N662);
nor NOR2 (N687, N681, N487);
not NOT1 (N688, N668);
xor XOR2 (N689, N680, N22);
not NOT1 (N690, N678);
not NOT1 (N691, N683);
not NOT1 (N692, N689);
nor NOR4 (N693, N691, N491, N646, N93);
and AND3 (N694, N692, N173, N372);
not NOT1 (N695, N686);
nor NOR2 (N696, N690, N316);
nand NAND2 (N697, N644, N284);
buf BUF1 (N698, N696);
not NOT1 (N699, N687);
or OR4 (N700, N694, N275, N643, N51);
not NOT1 (N701, N693);
nand NAND3 (N702, N669, N424, N487);
and AND2 (N703, N702, N690);
xor XOR2 (N704, N703, N119);
xor XOR2 (N705, N685, N47);
xor XOR2 (N706, N682, N559);
xor XOR2 (N707, N705, N620);
not NOT1 (N708, N697);
not NOT1 (N709, N707);
not NOT1 (N710, N701);
buf BUF1 (N711, N695);
xor XOR2 (N712, N699, N159);
buf BUF1 (N713, N712);
nor NOR4 (N714, N711, N462, N468, N434);
nand NAND2 (N715, N710, N527);
and AND4 (N716, N688, N530, N160, N285);
nand NAND4 (N717, N716, N612, N477, N237);
buf BUF1 (N718, N717);
xor XOR2 (N719, N708, N539);
buf BUF1 (N720, N719);
and AND4 (N721, N709, N661, N332, N481);
and AND2 (N722, N706, N437);
nor NOR4 (N723, N721, N284, N689, N373);
and AND4 (N724, N714, N387, N650, N24);
nor NOR2 (N725, N700, N289);
not NOT1 (N726, N724);
buf BUF1 (N727, N725);
and AND3 (N728, N727, N460, N397);
nand NAND3 (N729, N726, N381, N70);
and AND4 (N730, N728, N224, N675, N658);
and AND3 (N731, N704, N561, N517);
nand NAND3 (N732, N698, N685, N204);
nor NOR3 (N733, N715, N427, N37);
buf BUF1 (N734, N722);
or OR3 (N735, N718, N661, N673);
or OR3 (N736, N723, N294, N724);
nor NOR4 (N737, N730, N601, N530, N672);
not NOT1 (N738, N734);
or OR3 (N739, N731, N651, N254);
nor NOR3 (N740, N739, N729, N587);
and AND3 (N741, N352, N333, N529);
buf BUF1 (N742, N733);
xor XOR2 (N743, N737, N26);
nand NAND2 (N744, N743, N269);
buf BUF1 (N745, N740);
or OR2 (N746, N741, N744);
and AND4 (N747, N413, N89, N72, N374);
nand NAND2 (N748, N745, N657);
not NOT1 (N749, N732);
and AND3 (N750, N746, N435, N508);
nor NOR2 (N751, N748, N48);
nand NAND2 (N752, N735, N361);
nand NAND4 (N753, N713, N24, N643, N126);
not NOT1 (N754, N747);
xor XOR2 (N755, N753, N660);
xor XOR2 (N756, N742, N561);
nand NAND4 (N757, N751, N113, N269, N88);
nand NAND2 (N758, N752, N59);
xor XOR2 (N759, N750, N164);
or OR2 (N760, N749, N603);
or OR3 (N761, N754, N233, N446);
nand NAND2 (N762, N736, N183);
xor XOR2 (N763, N738, N670);
nand NAND4 (N764, N720, N695, N750, N650);
xor XOR2 (N765, N758, N656);
or OR2 (N766, N763, N77);
buf BUF1 (N767, N761);
nor NOR4 (N768, N760, N547, N336, N662);
nor NOR4 (N769, N765, N600, N307, N571);
xor XOR2 (N770, N766, N20);
buf BUF1 (N771, N757);
and AND3 (N772, N759, N55, N660);
and AND4 (N773, N769, N546, N505, N431);
not NOT1 (N774, N770);
or OR3 (N775, N762, N172, N260);
or OR2 (N776, N767, N264);
not NOT1 (N777, N774);
nor NOR3 (N778, N775, N581, N465);
nor NOR2 (N779, N773, N252);
nand NAND4 (N780, N755, N125, N402, N158);
buf BUF1 (N781, N768);
nor NOR2 (N782, N756, N663);
buf BUF1 (N783, N764);
and AND3 (N784, N780, N674, N768);
and AND2 (N785, N777, N279);
buf BUF1 (N786, N778);
and AND3 (N787, N779, N294, N29);
xor XOR2 (N788, N772, N65);
or OR3 (N789, N788, N413, N214);
not NOT1 (N790, N776);
nor NOR3 (N791, N781, N218, N238);
and AND2 (N792, N791, N330);
or OR2 (N793, N790, N528);
and AND4 (N794, N771, N58, N47, N11);
buf BUF1 (N795, N784);
nor NOR3 (N796, N782, N88, N374);
nor NOR2 (N797, N786, N498);
nor NOR2 (N798, N785, N133);
and AND3 (N799, N789, N238, N594);
nand NAND2 (N800, N793, N390);
buf BUF1 (N801, N787);
or OR2 (N802, N796, N717);
nand NAND4 (N803, N802, N787, N14, N596);
or OR4 (N804, N798, N388, N22, N95);
nand NAND3 (N805, N783, N261, N310);
not NOT1 (N806, N800);
or OR2 (N807, N795, N43);
buf BUF1 (N808, N803);
and AND3 (N809, N805, N237, N104);
or OR4 (N810, N792, N736, N316, N368);
or OR3 (N811, N804, N423, N207);
and AND2 (N812, N808, N456);
nand NAND3 (N813, N809, N245, N334);
buf BUF1 (N814, N807);
or OR3 (N815, N811, N313, N243);
or OR4 (N816, N815, N775, N215, N693);
nand NAND4 (N817, N806, N453, N213, N201);
not NOT1 (N818, N799);
nand NAND4 (N819, N812, N806, N452, N776);
xor XOR2 (N820, N810, N728);
not NOT1 (N821, N816);
nor NOR2 (N822, N794, N102);
nor NOR2 (N823, N819, N192);
nor NOR4 (N824, N813, N180, N54, N59);
xor XOR2 (N825, N817, N95);
and AND2 (N826, N797, N690);
nor NOR2 (N827, N824, N172);
not NOT1 (N828, N825);
nor NOR2 (N829, N826, N373);
nand NAND3 (N830, N820, N541, N199);
not NOT1 (N831, N830);
or OR3 (N832, N822, N37, N779);
not NOT1 (N833, N801);
nand NAND2 (N834, N828, N632);
not NOT1 (N835, N831);
nor NOR2 (N836, N834, N456);
buf BUF1 (N837, N836);
or OR2 (N838, N823, N692);
nor NOR2 (N839, N835, N278);
nand NAND2 (N840, N832, N141);
nand NAND3 (N841, N837, N278, N225);
and AND2 (N842, N838, N528);
or OR4 (N843, N821, N284, N447, N751);
xor XOR2 (N844, N843, N694);
nand NAND4 (N845, N840, N344, N160, N521);
nor NOR2 (N846, N818, N524);
xor XOR2 (N847, N827, N47);
or OR2 (N848, N829, N290);
and AND4 (N849, N845, N495, N118, N595);
not NOT1 (N850, N848);
and AND3 (N851, N844, N25, N338);
or OR4 (N852, N841, N661, N474, N627);
or OR3 (N853, N833, N338, N244);
or OR3 (N854, N846, N812, N293);
nand NAND3 (N855, N854, N472, N25);
and AND3 (N856, N814, N511, N370);
nand NAND3 (N857, N855, N227, N98);
buf BUF1 (N858, N857);
buf BUF1 (N859, N839);
or OR2 (N860, N852, N764);
xor XOR2 (N861, N859, N451);
or OR3 (N862, N860, N77, N808);
or OR3 (N863, N856, N458, N621);
or OR2 (N864, N851, N435);
or OR2 (N865, N849, N535);
and AND2 (N866, N858, N625);
nor NOR4 (N867, N847, N50, N386, N427);
not NOT1 (N868, N861);
and AND4 (N869, N868, N52, N830, N286);
buf BUF1 (N870, N864);
or OR2 (N871, N866, N167);
nor NOR4 (N872, N863, N342, N836, N313);
buf BUF1 (N873, N850);
nand NAND4 (N874, N872, N280, N503, N606);
nand NAND3 (N875, N873, N785, N220);
and AND4 (N876, N870, N339, N490, N576);
xor XOR2 (N877, N875, N375);
buf BUF1 (N878, N869);
not NOT1 (N879, N877);
buf BUF1 (N880, N874);
and AND3 (N881, N878, N868, N283);
xor XOR2 (N882, N876, N556);
xor XOR2 (N883, N853, N213);
xor XOR2 (N884, N862, N126);
or OR2 (N885, N871, N274);
nand NAND2 (N886, N867, N118);
nor NOR4 (N887, N886, N49, N868, N535);
or OR2 (N888, N885, N277);
and AND3 (N889, N884, N594, N472);
not NOT1 (N890, N882);
xor XOR2 (N891, N881, N608);
and AND4 (N892, N879, N471, N641, N296);
xor XOR2 (N893, N842, N418);
nor NOR3 (N894, N889, N361, N148);
nor NOR4 (N895, N880, N96, N426, N19);
nand NAND3 (N896, N893, N80, N735);
buf BUF1 (N897, N888);
nor NOR2 (N898, N894, N208);
not NOT1 (N899, N895);
and AND4 (N900, N887, N318, N606, N486);
and AND3 (N901, N897, N707, N698);
or OR3 (N902, N891, N115, N184);
nor NOR2 (N903, N898, N280);
nor NOR2 (N904, N896, N667);
not NOT1 (N905, N903);
not NOT1 (N906, N902);
buf BUF1 (N907, N900);
nor NOR4 (N908, N899, N560, N321, N248);
not NOT1 (N909, N904);
nor NOR4 (N910, N909, N185, N481, N353);
xor XOR2 (N911, N892, N727);
nor NOR3 (N912, N901, N773, N854);
or OR3 (N913, N910, N32, N570);
nor NOR3 (N914, N865, N906, N289);
xor XOR2 (N915, N427, N687);
nor NOR2 (N916, N907, N257);
not NOT1 (N917, N890);
not NOT1 (N918, N911);
not NOT1 (N919, N905);
not NOT1 (N920, N914);
buf BUF1 (N921, N912);
and AND2 (N922, N915, N747);
not NOT1 (N923, N921);
or OR3 (N924, N917, N596, N436);
nor NOR3 (N925, N919, N127, N400);
buf BUF1 (N926, N922);
nor NOR4 (N927, N925, N362, N222, N490);
nor NOR3 (N928, N908, N68, N720);
and AND2 (N929, N923, N499);
or OR4 (N930, N920, N313, N777, N775);
nor NOR2 (N931, N918, N202);
or OR4 (N932, N883, N712, N901, N6);
nor NOR3 (N933, N926, N896, N393);
and AND4 (N934, N930, N131, N670, N419);
buf BUF1 (N935, N931);
nand NAND4 (N936, N928, N505, N80, N640);
not NOT1 (N937, N913);
buf BUF1 (N938, N932);
nor NOR2 (N939, N937, N603);
not NOT1 (N940, N939);
buf BUF1 (N941, N924);
nand NAND4 (N942, N938, N94, N255, N797);
nand NAND3 (N943, N941, N751, N63);
nand NAND3 (N944, N935, N445, N309);
nor NOR4 (N945, N942, N97, N455, N595);
and AND2 (N946, N933, N555);
xor XOR2 (N947, N934, N467);
and AND2 (N948, N943, N695);
not NOT1 (N949, N944);
not NOT1 (N950, N947);
xor XOR2 (N951, N916, N548);
buf BUF1 (N952, N946);
xor XOR2 (N953, N950, N937);
and AND3 (N954, N952, N476, N255);
and AND4 (N955, N951, N461, N909, N289);
xor XOR2 (N956, N936, N478);
or OR2 (N957, N953, N666);
buf BUF1 (N958, N955);
nor NOR4 (N959, N957, N695, N672, N266);
nor NOR2 (N960, N940, N459);
nor NOR3 (N961, N960, N757, N564);
and AND2 (N962, N954, N340);
nor NOR4 (N963, N929, N782, N823, N215);
not NOT1 (N964, N961);
not NOT1 (N965, N948);
buf BUF1 (N966, N927);
buf BUF1 (N967, N962);
xor XOR2 (N968, N967, N773);
nand NAND4 (N969, N945, N278, N865, N202);
nand NAND4 (N970, N965, N746, N601, N251);
nor NOR2 (N971, N969, N640);
and AND2 (N972, N966, N377);
or OR3 (N973, N971, N349, N778);
not NOT1 (N974, N973);
nand NAND3 (N975, N968, N403, N239);
and AND4 (N976, N974, N870, N181, N7);
nor NOR4 (N977, N964, N914, N463, N282);
xor XOR2 (N978, N956, N727);
nand NAND2 (N979, N975, N512);
and AND4 (N980, N978, N671, N151, N141);
buf BUF1 (N981, N963);
xor XOR2 (N982, N981, N584);
buf BUF1 (N983, N982);
buf BUF1 (N984, N959);
buf BUF1 (N985, N979);
or OR4 (N986, N980, N30, N769, N229);
xor XOR2 (N987, N977, N118);
nor NOR4 (N988, N949, N743, N886, N676);
and AND4 (N989, N972, N508, N526, N769);
nor NOR4 (N990, N987, N635, N931, N499);
buf BUF1 (N991, N988);
xor XOR2 (N992, N990, N664);
xor XOR2 (N993, N984, N699);
nor NOR2 (N994, N989, N735);
nor NOR4 (N995, N991, N194, N299, N425);
buf BUF1 (N996, N993);
or OR4 (N997, N995, N837, N132, N727);
xor XOR2 (N998, N986, N772);
nand NAND4 (N999, N994, N522, N187, N285);
nand NAND3 (N1000, N997, N929, N959);
xor XOR2 (N1001, N992, N911);
or OR2 (N1002, N998, N573);
not NOT1 (N1003, N999);
and AND2 (N1004, N983, N69);
and AND4 (N1005, N1004, N134, N671, N782);
not NOT1 (N1006, N970);
and AND2 (N1007, N1000, N730);
xor XOR2 (N1008, N1003, N694);
buf BUF1 (N1009, N1005);
buf BUF1 (N1010, N1009);
and AND4 (N1011, N1010, N554, N967, N679);
xor XOR2 (N1012, N1006, N879);
not NOT1 (N1013, N1001);
xor XOR2 (N1014, N985, N469);
nand NAND4 (N1015, N976, N307, N241, N355);
xor XOR2 (N1016, N1008, N344);
buf BUF1 (N1017, N1016);
or OR3 (N1018, N1012, N530, N885);
or OR3 (N1019, N1011, N973, N49);
buf BUF1 (N1020, N1013);
not NOT1 (N1021, N1018);
xor XOR2 (N1022, N958, N724);
buf BUF1 (N1023, N1014);
or OR4 (N1024, N1015, N252, N389, N170);
buf BUF1 (N1025, N1024);
xor XOR2 (N1026, N1021, N600);
and AND4 (N1027, N1022, N186, N468, N152);
xor XOR2 (N1028, N1020, N169);
buf BUF1 (N1029, N1026);
or OR4 (N1030, N996, N1000, N119, N297);
and AND2 (N1031, N1002, N105);
and AND4 (N1032, N1019, N565, N975, N470);
and AND3 (N1033, N1025, N397, N954);
nand NAND3 (N1034, N1007, N214, N933);
and AND2 (N1035, N1032, N49);
and AND2 (N1036, N1027, N73);
xor XOR2 (N1037, N1028, N830);
xor XOR2 (N1038, N1037, N821);
not NOT1 (N1039, N1031);
or OR2 (N1040, N1038, N443);
xor XOR2 (N1041, N1030, N344);
not NOT1 (N1042, N1041);
and AND3 (N1043, N1039, N820, N762);
not NOT1 (N1044, N1033);
nand NAND4 (N1045, N1043, N661, N347, N529);
or OR4 (N1046, N1035, N884, N356, N53);
and AND4 (N1047, N1017, N162, N266, N614);
nand NAND4 (N1048, N1047, N362, N115, N437);
buf BUF1 (N1049, N1042);
nor NOR4 (N1050, N1040, N401, N14, N621);
not NOT1 (N1051, N1036);
xor XOR2 (N1052, N1051, N298);
nand NAND3 (N1053, N1050, N590, N496);
nand NAND4 (N1054, N1029, N915, N548, N516);
buf BUF1 (N1055, N1046);
xor XOR2 (N1056, N1044, N598);
and AND4 (N1057, N1034, N520, N950, N439);
xor XOR2 (N1058, N1049, N220);
and AND2 (N1059, N1053, N402);
not NOT1 (N1060, N1045);
buf BUF1 (N1061, N1056);
and AND4 (N1062, N1054, N3, N744, N718);
nand NAND2 (N1063, N1052, N860);
nand NAND2 (N1064, N1059, N596);
buf BUF1 (N1065, N1061);
or OR2 (N1066, N1064, N909);
xor XOR2 (N1067, N1057, N603);
not NOT1 (N1068, N1066);
and AND2 (N1069, N1048, N30);
nand NAND4 (N1070, N1063, N110, N259, N731);
xor XOR2 (N1071, N1055, N1070);
and AND4 (N1072, N655, N691, N662, N220);
and AND3 (N1073, N1068, N352, N809);
buf BUF1 (N1074, N1065);
and AND3 (N1075, N1072, N42, N12);
or OR3 (N1076, N1062, N163, N513);
nand NAND3 (N1077, N1074, N155, N380);
and AND3 (N1078, N1069, N853, N271);
or OR2 (N1079, N1075, N617);
xor XOR2 (N1080, N1023, N464);
or OR3 (N1081, N1060, N697, N445);
nand NAND2 (N1082, N1067, N220);
nand NAND3 (N1083, N1081, N125, N1051);
xor XOR2 (N1084, N1073, N651);
not NOT1 (N1085, N1078);
xor XOR2 (N1086, N1082, N148);
not NOT1 (N1087, N1058);
not NOT1 (N1088, N1079);
and AND4 (N1089, N1080, N5, N864, N954);
nand NAND4 (N1090, N1088, N1037, N419, N354);
not NOT1 (N1091, N1084);
and AND2 (N1092, N1085, N389);
or OR2 (N1093, N1076, N346);
nor NOR3 (N1094, N1089, N1040, N114);
nand NAND2 (N1095, N1083, N895);
nor NOR3 (N1096, N1094, N889, N354);
xor XOR2 (N1097, N1093, N333);
nand NAND2 (N1098, N1096, N871);
and AND4 (N1099, N1091, N861, N158, N769);
nand NAND3 (N1100, N1098, N647, N134);
or OR2 (N1101, N1090, N75);
not NOT1 (N1102, N1097);
not NOT1 (N1103, N1095);
or OR2 (N1104, N1103, N126);
nor NOR2 (N1105, N1071, N502);
and AND3 (N1106, N1092, N355, N568);
or OR3 (N1107, N1087, N1043, N724);
or OR3 (N1108, N1077, N12, N867);
buf BUF1 (N1109, N1100);
and AND3 (N1110, N1109, N998, N179);
nor NOR4 (N1111, N1101, N153, N18, N213);
not NOT1 (N1112, N1107);
xor XOR2 (N1113, N1102, N353);
or OR4 (N1114, N1106, N897, N201, N385);
nor NOR2 (N1115, N1104, N1056);
nor NOR2 (N1116, N1115, N139);
not NOT1 (N1117, N1116);
xor XOR2 (N1118, N1111, N645);
nor NOR3 (N1119, N1110, N75, N992);
buf BUF1 (N1120, N1113);
xor XOR2 (N1121, N1119, N374);
and AND2 (N1122, N1108, N843);
not NOT1 (N1123, N1120);
nand NAND2 (N1124, N1122, N600);
not NOT1 (N1125, N1123);
xor XOR2 (N1126, N1112, N40);
nor NOR4 (N1127, N1118, N613, N473, N947);
xor XOR2 (N1128, N1127, N489);
nor NOR3 (N1129, N1114, N240, N940);
xor XOR2 (N1130, N1129, N928);
and AND3 (N1131, N1121, N156, N921);
nor NOR4 (N1132, N1086, N362, N70, N805);
nand NAND4 (N1133, N1124, N783, N784, N955);
nand NAND3 (N1134, N1128, N1025, N474);
xor XOR2 (N1135, N1099, N879);
not NOT1 (N1136, N1135);
and AND2 (N1137, N1134, N982);
nand NAND2 (N1138, N1117, N34);
or OR4 (N1139, N1126, N36, N398, N459);
and AND4 (N1140, N1133, N939, N701, N863);
or OR3 (N1141, N1125, N449, N1060);
buf BUF1 (N1142, N1138);
not NOT1 (N1143, N1141);
nor NOR2 (N1144, N1136, N419);
nor NOR3 (N1145, N1143, N1071, N71);
xor XOR2 (N1146, N1105, N972);
xor XOR2 (N1147, N1137, N252);
or OR3 (N1148, N1139, N1039, N718);
or OR3 (N1149, N1130, N290, N746);
and AND2 (N1150, N1142, N1096);
buf BUF1 (N1151, N1149);
nor NOR2 (N1152, N1131, N822);
nor NOR2 (N1153, N1150, N1033);
nand NAND2 (N1154, N1140, N494);
xor XOR2 (N1155, N1148, N254);
or OR2 (N1156, N1152, N106);
and AND2 (N1157, N1155, N926);
and AND2 (N1158, N1157, N308);
buf BUF1 (N1159, N1156);
or OR3 (N1160, N1154, N459, N290);
nand NAND3 (N1161, N1160, N589, N714);
not NOT1 (N1162, N1158);
xor XOR2 (N1163, N1162, N1017);
nand NAND4 (N1164, N1159, N719, N499, N146);
not NOT1 (N1165, N1161);
not NOT1 (N1166, N1151);
xor XOR2 (N1167, N1146, N52);
xor XOR2 (N1168, N1163, N941);
xor XOR2 (N1169, N1132, N79);
buf BUF1 (N1170, N1167);
xor XOR2 (N1171, N1164, N416);
or OR2 (N1172, N1145, N53);
nor NOR3 (N1173, N1144, N3, N363);
xor XOR2 (N1174, N1170, N346);
or OR4 (N1175, N1153, N495, N386, N204);
nor NOR2 (N1176, N1172, N812);
buf BUF1 (N1177, N1173);
or OR2 (N1178, N1166, N835);
or OR2 (N1179, N1168, N437);
nand NAND2 (N1180, N1169, N144);
and AND4 (N1181, N1180, N1053, N805, N90);
or OR4 (N1182, N1176, N519, N623, N833);
nand NAND2 (N1183, N1165, N1165);
buf BUF1 (N1184, N1171);
buf BUF1 (N1185, N1181);
buf BUF1 (N1186, N1175);
nand NAND2 (N1187, N1182, N852);
nor NOR3 (N1188, N1187, N101, N926);
or OR2 (N1189, N1177, N316);
xor XOR2 (N1190, N1185, N350);
not NOT1 (N1191, N1186);
nor NOR4 (N1192, N1174, N267, N558, N500);
not NOT1 (N1193, N1147);
and AND3 (N1194, N1193, N1173, N269);
or OR3 (N1195, N1190, N45, N1058);
nor NOR3 (N1196, N1189, N318, N785);
or OR4 (N1197, N1194, N457, N463, N209);
buf BUF1 (N1198, N1178);
xor XOR2 (N1199, N1184, N222);
not NOT1 (N1200, N1199);
buf BUF1 (N1201, N1200);
or OR2 (N1202, N1198, N521);
nor NOR4 (N1203, N1183, N798, N205, N263);
xor XOR2 (N1204, N1191, N1067);
buf BUF1 (N1205, N1195);
nor NOR2 (N1206, N1205, N432);
not NOT1 (N1207, N1201);
nand NAND3 (N1208, N1207, N440, N69);
nand NAND2 (N1209, N1188, N535);
buf BUF1 (N1210, N1202);
nand NAND3 (N1211, N1206, N389, N249);
and AND2 (N1212, N1179, N1081);
not NOT1 (N1213, N1196);
and AND3 (N1214, N1204, N374, N1026);
nor NOR2 (N1215, N1214, N553);
nor NOR3 (N1216, N1215, N435, N1086);
or OR2 (N1217, N1211, N147);
nand NAND4 (N1218, N1197, N422, N703, N362);
buf BUF1 (N1219, N1212);
buf BUF1 (N1220, N1213);
not NOT1 (N1221, N1208);
nor NOR3 (N1222, N1220, N423, N53);
xor XOR2 (N1223, N1222, N277);
nor NOR2 (N1224, N1218, N659);
xor XOR2 (N1225, N1216, N30);
nor NOR4 (N1226, N1219, N200, N1056, N688);
buf BUF1 (N1227, N1203);
nor NOR4 (N1228, N1209, N661, N342, N164);
not NOT1 (N1229, N1217);
nand NAND3 (N1230, N1228, N835, N316);
and AND3 (N1231, N1223, N412, N669);
xor XOR2 (N1232, N1229, N241);
nand NAND3 (N1233, N1226, N526, N220);
not NOT1 (N1234, N1231);
and AND3 (N1235, N1221, N1019, N912);
not NOT1 (N1236, N1230);
nand NAND3 (N1237, N1236, N1028, N544);
xor XOR2 (N1238, N1227, N785);
or OR4 (N1239, N1232, N1006, N1078, N832);
buf BUF1 (N1240, N1192);
not NOT1 (N1241, N1234);
not NOT1 (N1242, N1210);
and AND3 (N1243, N1238, N857, N574);
nor NOR2 (N1244, N1240, N1107);
not NOT1 (N1245, N1244);
xor XOR2 (N1246, N1233, N973);
or OR4 (N1247, N1239, N226, N701, N1161);
nor NOR2 (N1248, N1224, N10);
or OR2 (N1249, N1246, N45);
buf BUF1 (N1250, N1225);
nor NOR4 (N1251, N1248, N1072, N464, N828);
not NOT1 (N1252, N1245);
xor XOR2 (N1253, N1242, N141);
not NOT1 (N1254, N1243);
not NOT1 (N1255, N1254);
and AND4 (N1256, N1251, N1134, N553, N460);
nor NOR3 (N1257, N1252, N1025, N22);
or OR3 (N1258, N1237, N734, N717);
nor NOR2 (N1259, N1258, N333);
or OR3 (N1260, N1247, N209, N454);
and AND3 (N1261, N1253, N671, N491);
not NOT1 (N1262, N1257);
xor XOR2 (N1263, N1259, N929);
not NOT1 (N1264, N1249);
nor NOR2 (N1265, N1241, N479);
nand NAND4 (N1266, N1235, N355, N1091, N905);
nand NAND4 (N1267, N1262, N484, N1148, N390);
buf BUF1 (N1268, N1266);
and AND4 (N1269, N1263, N733, N155, N753);
not NOT1 (N1270, N1265);
nand NAND3 (N1271, N1261, N1189, N792);
or OR2 (N1272, N1256, N649);
or OR3 (N1273, N1271, N1105, N1049);
and AND3 (N1274, N1268, N215, N1132);
buf BUF1 (N1275, N1264);
and AND4 (N1276, N1267, N389, N709, N876);
nand NAND4 (N1277, N1273, N75, N241, N1056);
nand NAND2 (N1278, N1277, N920);
buf BUF1 (N1279, N1274);
xor XOR2 (N1280, N1279, N1252);
and AND2 (N1281, N1260, N550);
and AND4 (N1282, N1270, N416, N1153, N476);
nor NOR4 (N1283, N1281, N184, N1018, N594);
nand NAND4 (N1284, N1278, N489, N1156, N102);
nand NAND3 (N1285, N1282, N267, N798);
and AND4 (N1286, N1285, N959, N389, N1269);
nor NOR2 (N1287, N607, N205);
buf BUF1 (N1288, N1250);
not NOT1 (N1289, N1272);
not NOT1 (N1290, N1276);
not NOT1 (N1291, N1283);
nor NOR4 (N1292, N1289, N221, N538, N266);
buf BUF1 (N1293, N1286);
or OR4 (N1294, N1292, N1110, N1149, N63);
nor NOR3 (N1295, N1290, N171, N614);
nor NOR4 (N1296, N1287, N873, N1115, N1184);
xor XOR2 (N1297, N1296, N863);
xor XOR2 (N1298, N1297, N219);
xor XOR2 (N1299, N1275, N710);
xor XOR2 (N1300, N1294, N392);
and AND4 (N1301, N1295, N229, N503, N93);
and AND3 (N1302, N1293, N1047, N319);
and AND3 (N1303, N1291, N910, N760);
nor NOR4 (N1304, N1300, N887, N1135, N965);
buf BUF1 (N1305, N1299);
nor NOR4 (N1306, N1301, N795, N679, N331);
nand NAND4 (N1307, N1304, N552, N835, N619);
xor XOR2 (N1308, N1288, N821);
nor NOR4 (N1309, N1298, N67, N1047, N124);
nand NAND2 (N1310, N1302, N739);
nand NAND3 (N1311, N1309, N98, N1014);
buf BUF1 (N1312, N1306);
or OR4 (N1313, N1308, N738, N694, N789);
not NOT1 (N1314, N1284);
not NOT1 (N1315, N1255);
xor XOR2 (N1316, N1280, N995);
and AND2 (N1317, N1311, N277);
nor NOR3 (N1318, N1310, N315, N545);
nand NAND2 (N1319, N1307, N683);
nand NAND3 (N1320, N1313, N1056, N539);
or OR3 (N1321, N1320, N766, N289);
nand NAND2 (N1322, N1316, N124);
nor NOR4 (N1323, N1321, N1258, N99, N863);
buf BUF1 (N1324, N1315);
nand NAND3 (N1325, N1317, N423, N1138);
xor XOR2 (N1326, N1305, N1237);
or OR2 (N1327, N1322, N922);
nor NOR2 (N1328, N1323, N201);
and AND3 (N1329, N1312, N564, N299);
nor NOR2 (N1330, N1318, N689);
nand NAND3 (N1331, N1325, N1186, N608);
and AND2 (N1332, N1330, N254);
nor NOR3 (N1333, N1331, N1008, N791);
nor NOR4 (N1334, N1324, N198, N692, N1235);
or OR3 (N1335, N1303, N638, N883);
or OR4 (N1336, N1334, N1185, N823, N834);
not NOT1 (N1337, N1326);
nand NAND3 (N1338, N1335, N376, N1111);
nand NAND4 (N1339, N1336, N536, N597, N1203);
xor XOR2 (N1340, N1332, N298);
xor XOR2 (N1341, N1339, N314);
not NOT1 (N1342, N1338);
nor NOR4 (N1343, N1319, N106, N753, N85);
and AND2 (N1344, N1314, N451);
xor XOR2 (N1345, N1343, N153);
and AND3 (N1346, N1328, N544, N1214);
and AND4 (N1347, N1341, N1176, N864, N654);
nand NAND4 (N1348, N1344, N1141, N821, N34);
xor XOR2 (N1349, N1345, N1090);
not NOT1 (N1350, N1342);
nand NAND4 (N1351, N1347, N1181, N196, N944);
buf BUF1 (N1352, N1351);
buf BUF1 (N1353, N1346);
buf BUF1 (N1354, N1353);
nand NAND2 (N1355, N1354, N535);
and AND2 (N1356, N1329, N80);
nand NAND3 (N1357, N1355, N969, N246);
buf BUF1 (N1358, N1352);
and AND4 (N1359, N1333, N69, N349, N643);
xor XOR2 (N1360, N1358, N984);
not NOT1 (N1361, N1348);
or OR3 (N1362, N1340, N257, N1180);
nand NAND3 (N1363, N1360, N415, N401);
nand NAND2 (N1364, N1363, N175);
and AND4 (N1365, N1327, N855, N91, N712);
buf BUF1 (N1366, N1357);
not NOT1 (N1367, N1364);
not NOT1 (N1368, N1349);
or OR4 (N1369, N1361, N668, N528, N984);
or OR3 (N1370, N1362, N1367, N622);
nor NOR4 (N1371, N1081, N387, N1326, N1022);
xor XOR2 (N1372, N1350, N386);
not NOT1 (N1373, N1369);
nand NAND4 (N1374, N1366, N1339, N610, N115);
nor NOR3 (N1375, N1372, N486, N1266);
xor XOR2 (N1376, N1368, N40);
not NOT1 (N1377, N1376);
xor XOR2 (N1378, N1337, N854);
and AND4 (N1379, N1370, N1238, N1221, N709);
nor NOR2 (N1380, N1356, N687);
xor XOR2 (N1381, N1375, N1065);
nand NAND4 (N1382, N1379, N555, N681, N1092);
xor XOR2 (N1383, N1381, N464);
not NOT1 (N1384, N1373);
nor NOR2 (N1385, N1384, N377);
nand NAND4 (N1386, N1380, N15, N429, N1346);
xor XOR2 (N1387, N1386, N27);
nor NOR4 (N1388, N1383, N678, N1356, N325);
not NOT1 (N1389, N1377);
xor XOR2 (N1390, N1389, N1327);
not NOT1 (N1391, N1387);
nand NAND3 (N1392, N1388, N876, N1063);
not NOT1 (N1393, N1392);
or OR4 (N1394, N1385, N397, N408, N1045);
buf BUF1 (N1395, N1382);
and AND2 (N1396, N1378, N147);
xor XOR2 (N1397, N1395, N153);
nor NOR2 (N1398, N1374, N225);
buf BUF1 (N1399, N1390);
xor XOR2 (N1400, N1359, N1244);
or OR4 (N1401, N1393, N1067, N1036, N360);
or OR3 (N1402, N1398, N740, N828);
xor XOR2 (N1403, N1401, N1129);
xor XOR2 (N1404, N1400, N286);
buf BUF1 (N1405, N1403);
and AND4 (N1406, N1404, N95, N1172, N467);
or OR4 (N1407, N1371, N304, N333, N1151);
or OR4 (N1408, N1397, N1085, N220, N316);
buf BUF1 (N1409, N1365);
nand NAND4 (N1410, N1391, N1064, N177, N524);
xor XOR2 (N1411, N1396, N1184);
and AND2 (N1412, N1405, N1020);
not NOT1 (N1413, N1399);
not NOT1 (N1414, N1407);
not NOT1 (N1415, N1408);
nor NOR3 (N1416, N1414, N566, N1275);
nor NOR4 (N1417, N1413, N62, N1406, N853);
and AND3 (N1418, N740, N806, N51);
buf BUF1 (N1419, N1410);
xor XOR2 (N1420, N1415, N191);
nand NAND3 (N1421, N1416, N446, N1196);
nor NOR3 (N1422, N1420, N54, N214);
not NOT1 (N1423, N1409);
nor NOR3 (N1424, N1423, N355, N111);
nor NOR4 (N1425, N1422, N284, N1221, N809);
nand NAND2 (N1426, N1402, N1355);
nand NAND2 (N1427, N1418, N937);
nor NOR4 (N1428, N1394, N824, N117, N660);
nor NOR2 (N1429, N1421, N56);
buf BUF1 (N1430, N1429);
not NOT1 (N1431, N1412);
not NOT1 (N1432, N1419);
or OR3 (N1433, N1424, N61, N518);
nand NAND2 (N1434, N1425, N1322);
nand NAND4 (N1435, N1428, N1189, N864, N781);
xor XOR2 (N1436, N1430, N853);
and AND4 (N1437, N1431, N1344, N192, N1010);
and AND2 (N1438, N1433, N358);
nor NOR2 (N1439, N1432, N1157);
not NOT1 (N1440, N1434);
nor NOR4 (N1441, N1440, N485, N353, N1322);
and AND4 (N1442, N1426, N1378, N134, N841);
nor NOR3 (N1443, N1427, N1039, N64);
and AND3 (N1444, N1443, N1269, N1419);
xor XOR2 (N1445, N1439, N390);
and AND4 (N1446, N1437, N1341, N59, N959);
not NOT1 (N1447, N1435);
nor NOR3 (N1448, N1441, N1437, N460);
buf BUF1 (N1449, N1417);
nor NOR4 (N1450, N1436, N380, N111, N1164);
xor XOR2 (N1451, N1438, N1027);
and AND2 (N1452, N1444, N1266);
not NOT1 (N1453, N1449);
or OR4 (N1454, N1446, N823, N88, N1030);
or OR4 (N1455, N1445, N1219, N1140, N1326);
buf BUF1 (N1456, N1442);
xor XOR2 (N1457, N1454, N905);
buf BUF1 (N1458, N1455);
xor XOR2 (N1459, N1458, N7);
buf BUF1 (N1460, N1457);
nand NAND3 (N1461, N1456, N907, N1121);
not NOT1 (N1462, N1411);
not NOT1 (N1463, N1462);
nand NAND2 (N1464, N1447, N793);
xor XOR2 (N1465, N1453, N1322);
buf BUF1 (N1466, N1465);
buf BUF1 (N1467, N1450);
or OR2 (N1468, N1459, N631);
buf BUF1 (N1469, N1451);
not NOT1 (N1470, N1467);
buf BUF1 (N1471, N1461);
nand NAND3 (N1472, N1470, N141, N1439);
not NOT1 (N1473, N1469);
and AND3 (N1474, N1460, N34, N1268);
xor XOR2 (N1475, N1452, N81);
xor XOR2 (N1476, N1472, N1121);
not NOT1 (N1477, N1448);
xor XOR2 (N1478, N1477, N1417);
and AND3 (N1479, N1468, N149, N415);
nand NAND2 (N1480, N1478, N625);
buf BUF1 (N1481, N1479);
and AND3 (N1482, N1475, N1442, N688);
xor XOR2 (N1483, N1482, N317);
not NOT1 (N1484, N1471);
and AND3 (N1485, N1481, N903, N499);
nor NOR4 (N1486, N1485, N841, N71, N219);
or OR3 (N1487, N1463, N843, N1363);
or OR4 (N1488, N1474, N1467, N161, N999);
not NOT1 (N1489, N1484);
nand NAND4 (N1490, N1488, N1122, N116, N530);
or OR2 (N1491, N1490, N1410);
nand NAND3 (N1492, N1483, N503, N1478);
nor NOR3 (N1493, N1486, N844, N1378);
xor XOR2 (N1494, N1476, N173);
buf BUF1 (N1495, N1466);
nor NOR2 (N1496, N1487, N373);
xor XOR2 (N1497, N1473, N1267);
buf BUF1 (N1498, N1491);
and AND4 (N1499, N1493, N211, N619, N260);
or OR2 (N1500, N1497, N1434);
nand NAND4 (N1501, N1489, N346, N1155, N53);
nor NOR3 (N1502, N1480, N1074, N1394);
not NOT1 (N1503, N1498);
nand NAND3 (N1504, N1464, N637, N364);
xor XOR2 (N1505, N1504, N686);
buf BUF1 (N1506, N1499);
nand NAND4 (N1507, N1501, N163, N1313, N526);
buf BUF1 (N1508, N1502);
not NOT1 (N1509, N1506);
buf BUF1 (N1510, N1495);
buf BUF1 (N1511, N1509);
and AND3 (N1512, N1505, N497, N592);
buf BUF1 (N1513, N1494);
or OR3 (N1514, N1496, N52, N1068);
buf BUF1 (N1515, N1492);
and AND4 (N1516, N1514, N312, N40, N222);
or OR4 (N1517, N1511, N926, N1404, N476);
or OR4 (N1518, N1516, N98, N741, N250);
not NOT1 (N1519, N1503);
buf BUF1 (N1520, N1512);
or OR2 (N1521, N1515, N1299);
and AND3 (N1522, N1500, N1084, N398);
not NOT1 (N1523, N1520);
or OR3 (N1524, N1510, N1058, N154);
not NOT1 (N1525, N1522);
and AND2 (N1526, N1521, N1010);
nand NAND2 (N1527, N1513, N256);
nor NOR3 (N1528, N1508, N1240, N1394);
nand NAND4 (N1529, N1517, N1417, N598, N1131);
buf BUF1 (N1530, N1526);
nor NOR3 (N1531, N1507, N952, N1020);
buf BUF1 (N1532, N1531);
nand NAND3 (N1533, N1523, N926, N476);
not NOT1 (N1534, N1518);
not NOT1 (N1535, N1527);
and AND2 (N1536, N1532, N518);
nor NOR4 (N1537, N1534, N1239, N755, N416);
or OR4 (N1538, N1519, N1528, N1082, N1450);
nor NOR4 (N1539, N140, N643, N379, N717);
and AND2 (N1540, N1524, N49);
buf BUF1 (N1541, N1530);
nor NOR4 (N1542, N1540, N1507, N364, N959);
and AND4 (N1543, N1541, N808, N224, N1116);
or OR2 (N1544, N1536, N145);
not NOT1 (N1545, N1538);
xor XOR2 (N1546, N1537, N796);
nand NAND4 (N1547, N1525, N723, N849, N1227);
not NOT1 (N1548, N1542);
not NOT1 (N1549, N1539);
nor NOR2 (N1550, N1544, N992);
or OR4 (N1551, N1548, N1041, N589, N690);
xor XOR2 (N1552, N1550, N173);
nand NAND2 (N1553, N1545, N33);
not NOT1 (N1554, N1552);
xor XOR2 (N1555, N1547, N353);
not NOT1 (N1556, N1549);
or OR4 (N1557, N1551, N732, N1324, N1315);
or OR3 (N1558, N1546, N233, N1530);
or OR3 (N1559, N1543, N1186, N341);
xor XOR2 (N1560, N1535, N696);
nor NOR2 (N1561, N1553, N293);
and AND2 (N1562, N1558, N704);
nor NOR4 (N1563, N1533, N593, N1392, N469);
buf BUF1 (N1564, N1559);
or OR2 (N1565, N1529, N1090);
buf BUF1 (N1566, N1564);
buf BUF1 (N1567, N1557);
and AND2 (N1568, N1561, N463);
nor NOR2 (N1569, N1554, N52);
not NOT1 (N1570, N1555);
or OR4 (N1571, N1566, N1370, N1288, N190);
nor NOR3 (N1572, N1569, N299, N973);
xor XOR2 (N1573, N1565, N1464);
and AND2 (N1574, N1573, N865);
or OR4 (N1575, N1571, N1336, N1114, N1261);
and AND3 (N1576, N1560, N575, N1023);
xor XOR2 (N1577, N1574, N1503);
not NOT1 (N1578, N1563);
nand NAND2 (N1579, N1578, N734);
not NOT1 (N1580, N1556);
nand NAND3 (N1581, N1572, N1177, N251);
nor NOR4 (N1582, N1579, N1, N1329, N1313);
not NOT1 (N1583, N1568);
nand NAND4 (N1584, N1581, N290, N987, N1064);
buf BUF1 (N1585, N1562);
nand NAND3 (N1586, N1570, N1454, N1185);
nand NAND2 (N1587, N1583, N1227);
or OR3 (N1588, N1584, N28, N1494);
nor NOR2 (N1589, N1577, N391);
xor XOR2 (N1590, N1589, N1065);
nor NOR3 (N1591, N1575, N242, N558);
and AND3 (N1592, N1576, N47, N265);
not NOT1 (N1593, N1586);
or OR3 (N1594, N1591, N1435, N1437);
nand NAND4 (N1595, N1588, N959, N1238, N390);
nor NOR4 (N1596, N1593, N691, N337, N907);
or OR4 (N1597, N1596, N1187, N895, N328);
not NOT1 (N1598, N1592);
and AND2 (N1599, N1567, N1203);
xor XOR2 (N1600, N1582, N1335);
or OR4 (N1601, N1594, N700, N314, N587);
nand NAND4 (N1602, N1590, N3, N1238, N119);
nor NOR2 (N1603, N1598, N980);
buf BUF1 (N1604, N1587);
xor XOR2 (N1605, N1604, N204);
nand NAND4 (N1606, N1580, N167, N204, N987);
buf BUF1 (N1607, N1601);
xor XOR2 (N1608, N1600, N489);
nor NOR4 (N1609, N1606, N423, N861, N846);
buf BUF1 (N1610, N1595);
not NOT1 (N1611, N1609);
or OR4 (N1612, N1607, N1227, N393, N1078);
buf BUF1 (N1613, N1599);
buf BUF1 (N1614, N1613);
and AND4 (N1615, N1597, N249, N526, N1200);
nor NOR4 (N1616, N1612, N1561, N257, N107);
nand NAND4 (N1617, N1608, N645, N805, N1323);
buf BUF1 (N1618, N1616);
and AND2 (N1619, N1617, N742);
or OR4 (N1620, N1585, N1243, N812, N451);
or OR4 (N1621, N1614, N868, N1598, N13);
or OR4 (N1622, N1602, N516, N1070, N192);
xor XOR2 (N1623, N1622, N68);
not NOT1 (N1624, N1621);
and AND2 (N1625, N1624, N455);
and AND4 (N1626, N1611, N841, N559, N1374);
nand NAND3 (N1627, N1618, N1264, N871);
and AND4 (N1628, N1605, N1140, N697, N1209);
buf BUF1 (N1629, N1610);
or OR4 (N1630, N1603, N529, N90, N1308);
not NOT1 (N1631, N1615);
or OR3 (N1632, N1623, N1288, N785);
and AND3 (N1633, N1626, N1341, N1051);
not NOT1 (N1634, N1620);
nand NAND2 (N1635, N1631, N1618);
xor XOR2 (N1636, N1625, N1628);
nor NOR4 (N1637, N449, N1318, N170, N254);
buf BUF1 (N1638, N1634);
xor XOR2 (N1639, N1632, N1298);
nand NAND2 (N1640, N1630, N1318);
nor NOR2 (N1641, N1638, N250);
or OR4 (N1642, N1619, N960, N320, N1249);
buf BUF1 (N1643, N1635);
and AND3 (N1644, N1629, N1398, N13);
not NOT1 (N1645, N1639);
or OR2 (N1646, N1643, N1367);
nor NOR2 (N1647, N1645, N689);
and AND4 (N1648, N1647, N1627, N717, N39);
or OR4 (N1649, N510, N1165, N868, N84);
and AND3 (N1650, N1649, N1417, N1030);
buf BUF1 (N1651, N1642);
or OR4 (N1652, N1646, N1317, N172, N1310);
nor NOR2 (N1653, N1651, N910);
nand NAND2 (N1654, N1650, N210);
and AND4 (N1655, N1633, N920, N231, N1265);
nor NOR2 (N1656, N1640, N1120);
not NOT1 (N1657, N1641);
not NOT1 (N1658, N1656);
buf BUF1 (N1659, N1652);
nand NAND3 (N1660, N1654, N1426, N303);
and AND4 (N1661, N1636, N1123, N666, N60);
or OR3 (N1662, N1660, N507, N1413);
buf BUF1 (N1663, N1644);
and AND3 (N1664, N1653, N498, N212);
nand NAND2 (N1665, N1659, N46);
nor NOR2 (N1666, N1663, N687);
xor XOR2 (N1667, N1648, N997);
or OR4 (N1668, N1667, N789, N410, N1171);
not NOT1 (N1669, N1661);
nor NOR3 (N1670, N1657, N305, N255);
nor NOR2 (N1671, N1664, N1633);
nand NAND3 (N1672, N1669, N1345, N1181);
or OR4 (N1673, N1637, N1016, N214, N199);
nand NAND4 (N1674, N1666, N1627, N1138, N771);
and AND2 (N1675, N1670, N1315);
or OR3 (N1676, N1672, N1669, N1675);
or OR2 (N1677, N887, N19);
buf BUF1 (N1678, N1658);
buf BUF1 (N1679, N1655);
xor XOR2 (N1680, N1677, N880);
nor NOR3 (N1681, N1676, N1496, N751);
nand NAND2 (N1682, N1662, N958);
nand NAND4 (N1683, N1665, N1597, N675, N1359);
xor XOR2 (N1684, N1673, N448);
xor XOR2 (N1685, N1683, N276);
and AND4 (N1686, N1681, N1209, N169, N817);
and AND2 (N1687, N1685, N345);
buf BUF1 (N1688, N1684);
xor XOR2 (N1689, N1682, N391);
and AND4 (N1690, N1680, N178, N464, N1105);
or OR4 (N1691, N1668, N104, N1102, N495);
xor XOR2 (N1692, N1674, N1113);
xor XOR2 (N1693, N1692, N1350);
not NOT1 (N1694, N1671);
nand NAND3 (N1695, N1693, N589, N1063);
xor XOR2 (N1696, N1689, N1681);
buf BUF1 (N1697, N1679);
buf BUF1 (N1698, N1686);
buf BUF1 (N1699, N1697);
buf BUF1 (N1700, N1699);
and AND3 (N1701, N1700, N568, N314);
or OR2 (N1702, N1678, N1316);
nor NOR2 (N1703, N1694, N1457);
buf BUF1 (N1704, N1701);
not NOT1 (N1705, N1696);
and AND4 (N1706, N1698, N1496, N1343, N1127);
or OR2 (N1707, N1705, N847);
nand NAND3 (N1708, N1707, N107, N438);
xor XOR2 (N1709, N1703, N1655);
buf BUF1 (N1710, N1690);
and AND2 (N1711, N1691, N1444);
not NOT1 (N1712, N1708);
not NOT1 (N1713, N1695);
not NOT1 (N1714, N1687);
buf BUF1 (N1715, N1710);
nand NAND2 (N1716, N1709, N591);
not NOT1 (N1717, N1715);
nor NOR4 (N1718, N1706, N1379, N1544, N730);
not NOT1 (N1719, N1702);
nand NAND3 (N1720, N1717, N786, N125);
not NOT1 (N1721, N1688);
and AND2 (N1722, N1720, N799);
xor XOR2 (N1723, N1719, N783);
nor NOR2 (N1724, N1716, N668);
buf BUF1 (N1725, N1718);
buf BUF1 (N1726, N1721);
xor XOR2 (N1727, N1726, N275);
buf BUF1 (N1728, N1711);
or OR2 (N1729, N1723, N158);
buf BUF1 (N1730, N1704);
not NOT1 (N1731, N1714);
nand NAND3 (N1732, N1728, N1034, N70);
and AND4 (N1733, N1712, N546, N862, N1500);
buf BUF1 (N1734, N1713);
nor NOR3 (N1735, N1722, N584, N985);
and AND2 (N1736, N1734, N283);
buf BUF1 (N1737, N1725);
xor XOR2 (N1738, N1727, N413);
nor NOR2 (N1739, N1738, N627);
nand NAND3 (N1740, N1735, N848, N1688);
not NOT1 (N1741, N1737);
or OR4 (N1742, N1732, N525, N1137, N700);
xor XOR2 (N1743, N1736, N1642);
not NOT1 (N1744, N1730);
nor NOR3 (N1745, N1742, N215, N800);
nand NAND4 (N1746, N1724, N687, N1551, N249);
not NOT1 (N1747, N1729);
nand NAND2 (N1748, N1739, N506);
not NOT1 (N1749, N1746);
not NOT1 (N1750, N1745);
not NOT1 (N1751, N1747);
buf BUF1 (N1752, N1731);
and AND3 (N1753, N1750, N1571, N1032);
or OR2 (N1754, N1752, N1675);
and AND4 (N1755, N1751, N36, N457, N598);
or OR4 (N1756, N1743, N1343, N534, N1427);
xor XOR2 (N1757, N1741, N519);
not NOT1 (N1758, N1756);
xor XOR2 (N1759, N1753, N1639);
not NOT1 (N1760, N1759);
xor XOR2 (N1761, N1733, N445);
nand NAND3 (N1762, N1754, N1706, N823);
nor NOR3 (N1763, N1740, N283, N1038);
and AND2 (N1764, N1757, N1318);
xor XOR2 (N1765, N1762, N604);
buf BUF1 (N1766, N1758);
nor NOR4 (N1767, N1763, N531, N1695, N769);
nor NOR3 (N1768, N1744, N1336, N107);
nand NAND3 (N1769, N1748, N1189, N162);
xor XOR2 (N1770, N1755, N1400);
nor NOR2 (N1771, N1761, N677);
nand NAND4 (N1772, N1767, N1027, N187, N54);
not NOT1 (N1773, N1768);
and AND2 (N1774, N1772, N1504);
nor NOR3 (N1775, N1765, N1541, N1187);
xor XOR2 (N1776, N1773, N1465);
nor NOR2 (N1777, N1774, N1063);
nand NAND4 (N1778, N1769, N1658, N292, N547);
and AND4 (N1779, N1775, N503, N1217, N1269);
and AND2 (N1780, N1771, N1139);
xor XOR2 (N1781, N1770, N1283);
and AND4 (N1782, N1777, N1740, N846, N147);
or OR3 (N1783, N1782, N400, N1193);
or OR4 (N1784, N1780, N1508, N1060, N1259);
not NOT1 (N1785, N1784);
and AND2 (N1786, N1785, N606);
and AND3 (N1787, N1779, N67, N383);
xor XOR2 (N1788, N1764, N593);
and AND2 (N1789, N1783, N813);
and AND2 (N1790, N1789, N224);
buf BUF1 (N1791, N1781);
or OR4 (N1792, N1766, N408, N512, N778);
xor XOR2 (N1793, N1788, N1154);
or OR3 (N1794, N1790, N418, N951);
nor NOR2 (N1795, N1749, N749);
or OR3 (N1796, N1786, N1367, N1724);
buf BUF1 (N1797, N1792);
nor NOR2 (N1798, N1776, N482);
not NOT1 (N1799, N1787);
xor XOR2 (N1800, N1799, N176);
nor NOR4 (N1801, N1796, N1066, N62, N1799);
not NOT1 (N1802, N1791);
nor NOR4 (N1803, N1795, N759, N1140, N1456);
and AND3 (N1804, N1803, N988, N4);
not NOT1 (N1805, N1793);
not NOT1 (N1806, N1804);
or OR2 (N1807, N1800, N1678);
xor XOR2 (N1808, N1797, N185);
or OR3 (N1809, N1802, N917, N208);
and AND3 (N1810, N1807, N505, N826);
not NOT1 (N1811, N1808);
or OR3 (N1812, N1810, N555, N39);
not NOT1 (N1813, N1760);
buf BUF1 (N1814, N1809);
or OR4 (N1815, N1812, N261, N1157, N959);
and AND4 (N1816, N1805, N1026, N1300, N578);
or OR4 (N1817, N1815, N755, N213, N1290);
buf BUF1 (N1818, N1816);
not NOT1 (N1819, N1794);
xor XOR2 (N1820, N1817, N124);
buf BUF1 (N1821, N1798);
nor NOR4 (N1822, N1806, N711, N106, N57);
xor XOR2 (N1823, N1813, N1667);
not NOT1 (N1824, N1818);
xor XOR2 (N1825, N1824, N1421);
buf BUF1 (N1826, N1778);
not NOT1 (N1827, N1811);
nand NAND2 (N1828, N1826, N889);
not NOT1 (N1829, N1823);
and AND2 (N1830, N1821, N775);
and AND4 (N1831, N1829, N273, N1660, N1797);
and AND3 (N1832, N1831, N1506, N463);
not NOT1 (N1833, N1801);
or OR3 (N1834, N1832, N656, N1585);
or OR2 (N1835, N1828, N1317);
nor NOR2 (N1836, N1830, N212);
xor XOR2 (N1837, N1814, N692);
or OR3 (N1838, N1825, N1522, N82);
and AND3 (N1839, N1820, N299, N67);
buf BUF1 (N1840, N1819);
xor XOR2 (N1841, N1827, N897);
and AND4 (N1842, N1833, N1190, N1057, N294);
and AND2 (N1843, N1835, N1207);
nand NAND2 (N1844, N1841, N1377);
or OR2 (N1845, N1843, N602);
nand NAND2 (N1846, N1834, N106);
nand NAND2 (N1847, N1842, N638);
nand NAND2 (N1848, N1847, N1434);
and AND4 (N1849, N1838, N1329, N201, N393);
nand NAND3 (N1850, N1844, N1785, N845);
or OR4 (N1851, N1850, N175, N255, N1273);
nor NOR2 (N1852, N1822, N159);
or OR3 (N1853, N1836, N779, N313);
nor NOR3 (N1854, N1848, N531, N961);
or OR4 (N1855, N1839, N148, N76, N1493);
nor NOR3 (N1856, N1851, N187, N1325);
not NOT1 (N1857, N1855);
or OR4 (N1858, N1852, N1269, N1540, N1724);
xor XOR2 (N1859, N1856, N327);
or OR2 (N1860, N1849, N666);
not NOT1 (N1861, N1846);
and AND2 (N1862, N1837, N475);
or OR4 (N1863, N1857, N847, N1860, N1277);
buf BUF1 (N1864, N19);
xor XOR2 (N1865, N1863, N178);
xor XOR2 (N1866, N1864, N392);
or OR3 (N1867, N1862, N484, N127);
xor XOR2 (N1868, N1853, N737);
nor NOR4 (N1869, N1858, N832, N1178, N1001);
and AND4 (N1870, N1859, N433, N681, N1353);
nor NOR2 (N1871, N1840, N1010);
nor NOR2 (N1872, N1854, N314);
xor XOR2 (N1873, N1861, N609);
or OR4 (N1874, N1871, N1684, N1316, N235);
not NOT1 (N1875, N1872);
xor XOR2 (N1876, N1868, N1771);
xor XOR2 (N1877, N1845, N987);
xor XOR2 (N1878, N1873, N859);
nand NAND3 (N1879, N1870, N758, N609);
nand NAND4 (N1880, N1867, N1604, N1594, N1258);
not NOT1 (N1881, N1869);
not NOT1 (N1882, N1876);
nor NOR3 (N1883, N1882, N696, N257);
xor XOR2 (N1884, N1878, N551);
nand NAND2 (N1885, N1883, N93);
or OR3 (N1886, N1884, N1117, N2);
buf BUF1 (N1887, N1885);
and AND2 (N1888, N1880, N1022);
xor XOR2 (N1889, N1881, N1792);
nand NAND3 (N1890, N1886, N1532, N597);
nor NOR2 (N1891, N1889, N830);
not NOT1 (N1892, N1890);
or OR3 (N1893, N1874, N120, N803);
and AND2 (N1894, N1866, N565);
buf BUF1 (N1895, N1887);
or OR2 (N1896, N1875, N206);
nor NOR4 (N1897, N1865, N1131, N254, N1584);
xor XOR2 (N1898, N1888, N183);
not NOT1 (N1899, N1896);
nand NAND3 (N1900, N1899, N1844, N1253);
buf BUF1 (N1901, N1877);
buf BUF1 (N1902, N1897);
or OR4 (N1903, N1879, N1734, N369, N1287);
or OR4 (N1904, N1900, N1761, N919, N160);
buf BUF1 (N1905, N1891);
xor XOR2 (N1906, N1901, N102);
and AND2 (N1907, N1895, N1820);
and AND4 (N1908, N1907, N528, N1751, N1047);
nor NOR4 (N1909, N1903, N163, N403, N10);
or OR4 (N1910, N1894, N742, N1473, N1001);
nand NAND4 (N1911, N1905, N1236, N1611, N39);
nand NAND4 (N1912, N1911, N1814, N541, N1261);
nor NOR3 (N1913, N1909, N272, N1575);
buf BUF1 (N1914, N1904);
or OR4 (N1915, N1912, N1034, N697, N1180);
not NOT1 (N1916, N1913);
and AND3 (N1917, N1910, N1134, N645);
not NOT1 (N1918, N1893);
xor XOR2 (N1919, N1892, N1626);
buf BUF1 (N1920, N1908);
buf BUF1 (N1921, N1906);
nand NAND2 (N1922, N1914, N1455);
xor XOR2 (N1923, N1920, N1160);
and AND2 (N1924, N1918, N99);
buf BUF1 (N1925, N1922);
xor XOR2 (N1926, N1921, N790);
nand NAND2 (N1927, N1923, N1139);
not NOT1 (N1928, N1927);
not NOT1 (N1929, N1926);
nand NAND2 (N1930, N1902, N563);
nand NAND3 (N1931, N1929, N375, N1542);
or OR4 (N1932, N1915, N177, N1812, N109);
or OR4 (N1933, N1925, N1258, N1410, N440);
nand NAND4 (N1934, N1932, N1384, N1610, N1815);
nor NOR2 (N1935, N1916, N616);
nor NOR4 (N1936, N1917, N1417, N289, N522);
xor XOR2 (N1937, N1928, N1679);
buf BUF1 (N1938, N1934);
xor XOR2 (N1939, N1937, N1538);
nand NAND4 (N1940, N1924, N1700, N817, N471);
nor NOR2 (N1941, N1940, N1847);
nand NAND4 (N1942, N1938, N216, N239, N961);
buf BUF1 (N1943, N1935);
nor NOR3 (N1944, N1942, N1667, N633);
not NOT1 (N1945, N1944);
buf BUF1 (N1946, N1933);
not NOT1 (N1947, N1919);
xor XOR2 (N1948, N1946, N1768);
or OR3 (N1949, N1939, N1650, N1293);
nand NAND4 (N1950, N1947, N1649, N1891, N1408);
not NOT1 (N1951, N1898);
not NOT1 (N1952, N1948);
or OR2 (N1953, N1930, N1665);
and AND2 (N1954, N1941, N1519);
xor XOR2 (N1955, N1949, N1928);
and AND2 (N1956, N1954, N1328);
nor NOR4 (N1957, N1952, N493, N666, N1296);
xor XOR2 (N1958, N1936, N942);
not NOT1 (N1959, N1951);
buf BUF1 (N1960, N1959);
or OR2 (N1961, N1957, N1865);
nor NOR4 (N1962, N1943, N134, N1079, N1471);
xor XOR2 (N1963, N1961, N127);
buf BUF1 (N1964, N1956);
nor NOR3 (N1965, N1931, N1292, N871);
and AND3 (N1966, N1955, N464, N694);
nand NAND3 (N1967, N1962, N781, N1572);
not NOT1 (N1968, N1960);
and AND4 (N1969, N1964, N331, N40, N756);
not NOT1 (N1970, N1967);
xor XOR2 (N1971, N1963, N1280);
buf BUF1 (N1972, N1971);
nor NOR3 (N1973, N1968, N1452, N757);
not NOT1 (N1974, N1953);
buf BUF1 (N1975, N1973);
and AND2 (N1976, N1966, N153);
nor NOR3 (N1977, N1958, N1333, N1872);
buf BUF1 (N1978, N1950);
nor NOR3 (N1979, N1972, N1958, N1626);
nor NOR2 (N1980, N1969, N1394);
not NOT1 (N1981, N1970);
or OR2 (N1982, N1965, N672);
buf BUF1 (N1983, N1975);
not NOT1 (N1984, N1981);
or OR4 (N1985, N1974, N1268, N1882, N393);
buf BUF1 (N1986, N1976);
nand NAND2 (N1987, N1985, N224);
or OR2 (N1988, N1986, N445);
buf BUF1 (N1989, N1945);
nor NOR4 (N1990, N1978, N1932, N658, N358);
buf BUF1 (N1991, N1989);
xor XOR2 (N1992, N1984, N1725);
not NOT1 (N1993, N1979);
not NOT1 (N1994, N1982);
xor XOR2 (N1995, N1980, N404);
not NOT1 (N1996, N1977);
or OR4 (N1997, N1994, N87, N1990, N228);
xor XOR2 (N1998, N505, N1206);
buf BUF1 (N1999, N1987);
nand NAND2 (N2000, N1983, N1839);
nor NOR3 (N2001, N1988, N284, N1838);
buf BUF1 (N2002, N1996);
not NOT1 (N2003, N1998);
nor NOR3 (N2004, N2000, N346, N844);
and AND4 (N2005, N1991, N749, N347, N131);
xor XOR2 (N2006, N1992, N182);
or OR2 (N2007, N2005, N144);
nand NAND4 (N2008, N2006, N386, N370, N830);
xor XOR2 (N2009, N1993, N290);
and AND4 (N2010, N2004, N1288, N1388, N843);
nor NOR2 (N2011, N2001, N831);
nand NAND2 (N2012, N2003, N1378);
nor NOR4 (N2013, N2012, N784, N1223, N295);
or OR2 (N2014, N2011, N713);
nor NOR4 (N2015, N1997, N589, N1945, N1844);
or OR2 (N2016, N2008, N752);
buf BUF1 (N2017, N2014);
buf BUF1 (N2018, N2013);
or OR4 (N2019, N2017, N1488, N956, N222);
xor XOR2 (N2020, N1995, N551);
xor XOR2 (N2021, N2010, N1630);
buf BUF1 (N2022, N2016);
nor NOR2 (N2023, N2020, N1324);
nand NAND3 (N2024, N2019, N326, N1095);
and AND2 (N2025, N2002, N299);
or OR2 (N2026, N2025, N989);
nand NAND3 (N2027, N2024, N1078, N1571);
buf BUF1 (N2028, N2027);
or OR3 (N2029, N2026, N1434, N1387);
not NOT1 (N2030, N2022);
xor XOR2 (N2031, N2028, N1674);
not NOT1 (N2032, N2007);
not NOT1 (N2033, N2009);
nand NAND4 (N2034, N2023, N1264, N687, N1033);
or OR3 (N2035, N2034, N31, N715);
nand NAND2 (N2036, N2035, N1280);
or OR3 (N2037, N2031, N1760, N1413);
xor XOR2 (N2038, N2015, N528);
nand NAND3 (N2039, N2021, N874, N1526);
or OR3 (N2040, N2039, N767, N894);
not NOT1 (N2041, N2036);
and AND4 (N2042, N2029, N246, N171, N1927);
nor NOR2 (N2043, N2041, N247);
buf BUF1 (N2044, N2038);
xor XOR2 (N2045, N2033, N1787);
and AND3 (N2046, N2044, N2012, N95);
xor XOR2 (N2047, N2030, N766);
not NOT1 (N2048, N2042);
and AND3 (N2049, N2045, N1402, N1000);
and AND4 (N2050, N2018, N99, N294, N1141);
and AND3 (N2051, N2043, N1931, N1614);
or OR4 (N2052, N2037, N1633, N603, N1822);
nor NOR4 (N2053, N2052, N224, N1103, N318);
xor XOR2 (N2054, N2053, N65);
nand NAND2 (N2055, N2051, N1754);
nand NAND4 (N2056, N2055, N978, N1405, N1223);
not NOT1 (N2057, N2040);
nand NAND4 (N2058, N2057, N1914, N1500, N1909);
buf BUF1 (N2059, N2058);
nor NOR3 (N2060, N2047, N509, N133);
or OR4 (N2061, N2048, N1531, N1480, N660);
buf BUF1 (N2062, N2032);
or OR3 (N2063, N2060, N495, N782);
nand NAND2 (N2064, N2049, N1102);
and AND3 (N2065, N2046, N1764, N669);
xor XOR2 (N2066, N2064, N1753);
and AND4 (N2067, N2063, N1137, N1723, N1159);
and AND3 (N2068, N2056, N17, N1424);
or OR3 (N2069, N2050, N1010, N1071);
xor XOR2 (N2070, N2054, N731);
and AND2 (N2071, N2062, N713);
and AND3 (N2072, N2061, N1415, N1782);
buf BUF1 (N2073, N1999);
and AND2 (N2074, N2071, N1418);
buf BUF1 (N2075, N2073);
and AND3 (N2076, N2075, N1339, N2027);
nor NOR3 (N2077, N2067, N594, N908);
nand NAND4 (N2078, N2072, N1802, N932, N975);
or OR2 (N2079, N2069, N1659);
or OR2 (N2080, N2074, N825);
nand NAND2 (N2081, N2078, N972);
nand NAND3 (N2082, N2059, N622, N304);
xor XOR2 (N2083, N2066, N1562);
nor NOR2 (N2084, N2082, N1611);
nor NOR3 (N2085, N2080, N960, N2067);
not NOT1 (N2086, N2076);
and AND2 (N2087, N2083, N592);
and AND4 (N2088, N2065, N1593, N603, N1979);
nand NAND4 (N2089, N2081, N585, N345, N989);
xor XOR2 (N2090, N2089, N1249);
buf BUF1 (N2091, N2090);
and AND4 (N2092, N2088, N1811, N2003, N1479);
nand NAND3 (N2093, N2091, N763, N1003);
nand NAND4 (N2094, N2085, N1619, N416, N1190);
nor NOR2 (N2095, N2084, N1183);
buf BUF1 (N2096, N2087);
nand NAND4 (N2097, N2070, N1422, N560, N65);
xor XOR2 (N2098, N2079, N66);
not NOT1 (N2099, N2093);
xor XOR2 (N2100, N2096, N1453);
or OR3 (N2101, N2098, N1649, N203);
or OR2 (N2102, N2095, N454);
and AND4 (N2103, N2102, N418, N1283, N1900);
not NOT1 (N2104, N2092);
nand NAND4 (N2105, N2104, N1013, N314, N1715);
or OR4 (N2106, N2094, N1807, N657, N1186);
nor NOR3 (N2107, N2101, N2074, N1944);
nand NAND2 (N2108, N2100, N541);
and AND3 (N2109, N2068, N2088, N1899);
or OR3 (N2110, N2086, N290, N1453);
not NOT1 (N2111, N2108);
nand NAND4 (N2112, N2077, N1206, N118, N1742);
nor NOR4 (N2113, N2099, N1155, N1729, N1739);
and AND2 (N2114, N2107, N2085);
xor XOR2 (N2115, N2113, N1895);
nor NOR2 (N2116, N2106, N306);
nor NOR2 (N2117, N2110, N989);
xor XOR2 (N2118, N2112, N953);
buf BUF1 (N2119, N2117);
not NOT1 (N2120, N2103);
nor NOR4 (N2121, N2120, N392, N1988, N549);
or OR3 (N2122, N2109, N1874, N2096);
xor XOR2 (N2123, N2115, N367);
nor NOR2 (N2124, N2105, N1931);
and AND3 (N2125, N2121, N1275, N507);
not NOT1 (N2126, N2111);
xor XOR2 (N2127, N2116, N328);
or OR3 (N2128, N2126, N252, N589);
xor XOR2 (N2129, N2097, N343);
or OR4 (N2130, N2119, N373, N1166, N65);
not NOT1 (N2131, N2129);
buf BUF1 (N2132, N2124);
nor NOR3 (N2133, N2114, N173, N537);
nor NOR4 (N2134, N2118, N2030, N1071, N1550);
and AND2 (N2135, N2133, N2123);
and AND4 (N2136, N95, N355, N267, N1837);
buf BUF1 (N2137, N2127);
not NOT1 (N2138, N2137);
nand NAND2 (N2139, N2130, N1043);
or OR3 (N2140, N2135, N1315, N666);
and AND4 (N2141, N2132, N596, N1883, N1447);
xor XOR2 (N2142, N2136, N1969);
not NOT1 (N2143, N2140);
nor NOR4 (N2144, N2125, N1283, N941, N1566);
not NOT1 (N2145, N2143);
or OR4 (N2146, N2122, N81, N2074, N874);
nor NOR3 (N2147, N2134, N1295, N199);
nor NOR4 (N2148, N2144, N577, N1953, N468);
not NOT1 (N2149, N2147);
and AND2 (N2150, N2131, N456);
not NOT1 (N2151, N2142);
and AND3 (N2152, N2138, N1745, N1926);
not NOT1 (N2153, N2145);
or OR2 (N2154, N2149, N1543);
not NOT1 (N2155, N2146);
nor NOR2 (N2156, N2151, N2144);
xor XOR2 (N2157, N2128, N1455);
not NOT1 (N2158, N2141);
nand NAND2 (N2159, N2148, N603);
and AND4 (N2160, N2150, N375, N1636, N1958);
xor XOR2 (N2161, N2152, N980);
or OR2 (N2162, N2154, N85);
nor NOR3 (N2163, N2158, N1116, N912);
nand NAND3 (N2164, N2159, N39, N577);
not NOT1 (N2165, N2155);
not NOT1 (N2166, N2139);
buf BUF1 (N2167, N2166);
or OR4 (N2168, N2156, N2026, N969, N1926);
not NOT1 (N2169, N2165);
xor XOR2 (N2170, N2157, N520);
nand NAND3 (N2171, N2160, N1175, N1417);
xor XOR2 (N2172, N2171, N21);
or OR4 (N2173, N2172, N1328, N852, N544);
or OR4 (N2174, N2167, N1872, N1552, N1507);
buf BUF1 (N2175, N2153);
xor XOR2 (N2176, N2163, N1451);
xor XOR2 (N2177, N2169, N728);
nor NOR3 (N2178, N2168, N1262, N1791);
xor XOR2 (N2179, N2174, N10);
not NOT1 (N2180, N2162);
xor XOR2 (N2181, N2170, N1379);
and AND4 (N2182, N2179, N1068, N1401, N910);
or OR2 (N2183, N2175, N1090);
xor XOR2 (N2184, N2173, N1781);
xor XOR2 (N2185, N2176, N1399);
and AND3 (N2186, N2164, N900, N155);
nand NAND3 (N2187, N2184, N2183, N549);
and AND2 (N2188, N31, N160);
not NOT1 (N2189, N2161);
nor NOR4 (N2190, N2177, N895, N1820, N557);
and AND2 (N2191, N2180, N1144);
nand NAND3 (N2192, N2188, N145, N1057);
nand NAND4 (N2193, N2182, N1190, N726, N1175);
and AND3 (N2194, N2193, N87, N1157);
nand NAND2 (N2195, N2192, N737);
nand NAND3 (N2196, N2195, N1734, N1855);
xor XOR2 (N2197, N2181, N726);
not NOT1 (N2198, N2178);
and AND4 (N2199, N2186, N2077, N308, N1715);
xor XOR2 (N2200, N2187, N95);
nor NOR4 (N2201, N2189, N2077, N683, N1301);
not NOT1 (N2202, N2198);
or OR2 (N2203, N2185, N944);
or OR2 (N2204, N2196, N488);
buf BUF1 (N2205, N2191);
nor NOR4 (N2206, N2204, N1637, N741, N609);
not NOT1 (N2207, N2205);
nor NOR4 (N2208, N2202, N1467, N1169, N254);
not NOT1 (N2209, N2199);
xor XOR2 (N2210, N2208, N832);
xor XOR2 (N2211, N2197, N545);
not NOT1 (N2212, N2211);
and AND2 (N2213, N2210, N935);
and AND4 (N2214, N2206, N1310, N1679, N418);
and AND4 (N2215, N2214, N2210, N1365, N1158);
and AND3 (N2216, N2201, N722, N1160);
xor XOR2 (N2217, N2215, N639);
buf BUF1 (N2218, N2190);
not NOT1 (N2219, N2217);
and AND3 (N2220, N2213, N606, N927);
or OR2 (N2221, N2212, N2106);
nor NOR3 (N2222, N2221, N903, N1634);
or OR3 (N2223, N2216, N1588, N1731);
nand NAND3 (N2224, N2203, N119, N1306);
nor NOR2 (N2225, N2224, N639);
not NOT1 (N2226, N2207);
not NOT1 (N2227, N2219);
nor NOR3 (N2228, N2218, N1270, N1852);
not NOT1 (N2229, N2223);
not NOT1 (N2230, N2228);
nand NAND3 (N2231, N2194, N146, N1756);
nand NAND3 (N2232, N2209, N1025, N1033);
nor NOR3 (N2233, N2226, N126, N859);
xor XOR2 (N2234, N2220, N1208);
or OR2 (N2235, N2231, N1885);
or OR2 (N2236, N2233, N565);
xor XOR2 (N2237, N2225, N2223);
nor NOR4 (N2238, N2234, N1925, N1134, N1297);
not NOT1 (N2239, N2237);
nor NOR2 (N2240, N2235, N1004);
buf BUF1 (N2241, N2239);
and AND4 (N2242, N2238, N1577, N1986, N738);
xor XOR2 (N2243, N2227, N2056);
buf BUF1 (N2244, N2241);
not NOT1 (N2245, N2244);
nand NAND3 (N2246, N2243, N335, N121);
and AND3 (N2247, N2200, N537, N741);
and AND2 (N2248, N2242, N1022);
buf BUF1 (N2249, N2247);
nand NAND2 (N2250, N2248, N2243);
buf BUF1 (N2251, N2249);
buf BUF1 (N2252, N2222);
xor XOR2 (N2253, N2252, N2121);
not NOT1 (N2254, N2246);
and AND3 (N2255, N2229, N1839, N599);
not NOT1 (N2256, N2253);
not NOT1 (N2257, N2245);
and AND2 (N2258, N2257, N1516);
or OR2 (N2259, N2254, N2150);
xor XOR2 (N2260, N2251, N1850);
and AND4 (N2261, N2256, N864, N335, N942);
xor XOR2 (N2262, N2260, N1533);
nand NAND4 (N2263, N2258, N741, N328, N1417);
xor XOR2 (N2264, N2263, N530);
xor XOR2 (N2265, N2264, N869);
nor NOR2 (N2266, N2255, N180);
buf BUF1 (N2267, N2259);
xor XOR2 (N2268, N2232, N1743);
buf BUF1 (N2269, N2236);
xor XOR2 (N2270, N2250, N1445);
nor NOR3 (N2271, N2265, N1983, N2091);
not NOT1 (N2272, N2262);
nor NOR2 (N2273, N2267, N163);
nor NOR2 (N2274, N2261, N1488);
buf BUF1 (N2275, N2272);
xor XOR2 (N2276, N2266, N1425);
and AND2 (N2277, N2274, N2023);
nand NAND4 (N2278, N2270, N1227, N1370, N1890);
xor XOR2 (N2279, N2240, N634);
nor NOR3 (N2280, N2271, N314, N1650);
and AND3 (N2281, N2230, N1558, N787);
nor NOR3 (N2282, N2269, N2026, N166);
and AND4 (N2283, N2276, N2087, N1839, N591);
buf BUF1 (N2284, N2277);
not NOT1 (N2285, N2279);
buf BUF1 (N2286, N2282);
and AND2 (N2287, N2285, N1571);
buf BUF1 (N2288, N2268);
nor NOR4 (N2289, N2288, N1464, N1996, N1002);
buf BUF1 (N2290, N2280);
xor XOR2 (N2291, N2286, N1410);
xor XOR2 (N2292, N2291, N82);
or OR3 (N2293, N2290, N1432, N1354);
nor NOR4 (N2294, N2273, N274, N888, N2021);
nor NOR2 (N2295, N2289, N1108);
buf BUF1 (N2296, N2287);
not NOT1 (N2297, N2278);
and AND2 (N2298, N2275, N448);
xor XOR2 (N2299, N2284, N1373);
buf BUF1 (N2300, N2292);
and AND4 (N2301, N2298, N876, N768, N143);
xor XOR2 (N2302, N2297, N1196);
or OR2 (N2303, N2293, N906);
or OR4 (N2304, N2295, N882, N215, N1798);
and AND3 (N2305, N2294, N11, N2149);
and AND2 (N2306, N2304, N1794);
nor NOR3 (N2307, N2300, N2302, N381);
or OR3 (N2308, N1496, N1692, N89);
nand NAND3 (N2309, N2296, N1260, N2154);
not NOT1 (N2310, N2281);
xor XOR2 (N2311, N2309, N2262);
and AND3 (N2312, N2283, N1010, N36);
xor XOR2 (N2313, N2312, N1089);
buf BUF1 (N2314, N2301);
not NOT1 (N2315, N2311);
or OR3 (N2316, N2308, N715, N1079);
nor NOR3 (N2317, N2305, N297, N2032);
nor NOR2 (N2318, N2307, N1728);
not NOT1 (N2319, N2314);
nor NOR4 (N2320, N2316, N2003, N1526, N532);
buf BUF1 (N2321, N2310);
or OR4 (N2322, N2319, N1349, N2157, N1622);
nand NAND2 (N2323, N2313, N2309);
nor NOR3 (N2324, N2303, N150, N1432);
buf BUF1 (N2325, N2315);
or OR3 (N2326, N2324, N148, N1460);
not NOT1 (N2327, N2299);
buf BUF1 (N2328, N2320);
nor NOR2 (N2329, N2317, N1963);
xor XOR2 (N2330, N2306, N2281);
and AND2 (N2331, N2327, N793);
nor NOR4 (N2332, N2318, N63, N2189, N2260);
nand NAND3 (N2333, N2326, N1105, N1866);
xor XOR2 (N2334, N2330, N322);
nand NAND4 (N2335, N2322, N2055, N582, N756);
nand NAND4 (N2336, N2335, N420, N380, N325);
and AND2 (N2337, N2336, N1599);
and AND2 (N2338, N2329, N2079);
and AND3 (N2339, N2323, N138, N1910);
xor XOR2 (N2340, N2333, N1714);
and AND3 (N2341, N2334, N246, N249);
nor NOR4 (N2342, N2337, N662, N2266, N259);
buf BUF1 (N2343, N2338);
nand NAND4 (N2344, N2321, N808, N901, N1961);
or OR4 (N2345, N2344, N516, N2186, N1089);
buf BUF1 (N2346, N2343);
nor NOR2 (N2347, N2328, N1342);
xor XOR2 (N2348, N2342, N962);
or OR3 (N2349, N2340, N631, N977);
nand NAND2 (N2350, N2346, N497);
buf BUF1 (N2351, N2348);
nand NAND3 (N2352, N2349, N354, N1098);
nand NAND2 (N2353, N2347, N765);
and AND4 (N2354, N2351, N1079, N1422, N672);
not NOT1 (N2355, N2350);
nand NAND4 (N2356, N2339, N1189, N1945, N1840);
xor XOR2 (N2357, N2325, N1278);
or OR2 (N2358, N2345, N856);
buf BUF1 (N2359, N2353);
not NOT1 (N2360, N2331);
xor XOR2 (N2361, N2358, N1606);
xor XOR2 (N2362, N2341, N274);
not NOT1 (N2363, N2332);
or OR4 (N2364, N2356, N1839, N1484, N637);
nor NOR3 (N2365, N2360, N2216, N124);
buf BUF1 (N2366, N2364);
and AND3 (N2367, N2361, N821, N601);
nor NOR3 (N2368, N2367, N1503, N900);
buf BUF1 (N2369, N2365);
and AND4 (N2370, N2362, N2351, N17, N356);
nand NAND2 (N2371, N2354, N768);
nor NOR2 (N2372, N2371, N1494);
nor NOR4 (N2373, N2372, N899, N1747, N988);
not NOT1 (N2374, N2363);
nand NAND3 (N2375, N2369, N391, N2081);
nand NAND2 (N2376, N2375, N1810);
xor XOR2 (N2377, N2366, N120);
nor NOR4 (N2378, N2359, N1783, N1168, N963);
buf BUF1 (N2379, N2357);
xor XOR2 (N2380, N2352, N818);
or OR2 (N2381, N2370, N1087);
and AND4 (N2382, N2380, N511, N1052, N2097);
buf BUF1 (N2383, N2376);
nor NOR3 (N2384, N2368, N1158, N1915);
nand NAND4 (N2385, N2383, N1174, N246, N320);
nor NOR2 (N2386, N2382, N1052);
and AND3 (N2387, N2355, N1328, N1487);
buf BUF1 (N2388, N2384);
or OR3 (N2389, N2378, N2022, N524);
or OR3 (N2390, N2374, N1145, N1514);
nor NOR2 (N2391, N2389, N71);
nand NAND3 (N2392, N2377, N300, N71);
nand NAND2 (N2393, N2391, N1403);
xor XOR2 (N2394, N2373, N1570);
nand NAND4 (N2395, N2379, N905, N1950, N2280);
or OR2 (N2396, N2386, N1825);
buf BUF1 (N2397, N2387);
nand NAND4 (N2398, N2395, N1676, N2029, N1694);
nor NOR2 (N2399, N2388, N1009);
xor XOR2 (N2400, N2381, N399);
nor NOR4 (N2401, N2400, N407, N2246, N1651);
nand NAND2 (N2402, N2393, N1846);
nor NOR4 (N2403, N2385, N1935, N905, N288);
xor XOR2 (N2404, N2398, N1150);
or OR3 (N2405, N2404, N1832, N216);
nor NOR3 (N2406, N2402, N453, N12);
or OR3 (N2407, N2406, N1513, N1235);
or OR2 (N2408, N2405, N1990);
not NOT1 (N2409, N2394);
or OR2 (N2410, N2407, N2339);
and AND2 (N2411, N2397, N223);
nor NOR4 (N2412, N2410, N2311, N51, N129);
buf BUF1 (N2413, N2409);
or OR4 (N2414, N2408, N268, N1360, N639);
nor NOR3 (N2415, N2414, N14, N1320);
nor NOR4 (N2416, N2411, N1271, N1511, N2032);
nand NAND3 (N2417, N2392, N268, N1923);
buf BUF1 (N2418, N2412);
or OR4 (N2419, N2399, N1437, N985, N2120);
or OR3 (N2420, N2403, N556, N624);
buf BUF1 (N2421, N2401);
buf BUF1 (N2422, N2415);
not NOT1 (N2423, N2422);
xor XOR2 (N2424, N2423, N958);
or OR3 (N2425, N2396, N449, N1197);
and AND2 (N2426, N2418, N1176);
xor XOR2 (N2427, N2413, N313);
nor NOR4 (N2428, N2425, N1069, N256, N898);
or OR3 (N2429, N2417, N1621, N1743);
and AND3 (N2430, N2426, N2233, N1866);
xor XOR2 (N2431, N2429, N1961);
nor NOR3 (N2432, N2431, N1558, N2248);
not NOT1 (N2433, N2427);
or OR4 (N2434, N2420, N913, N1810, N1489);
buf BUF1 (N2435, N2424);
and AND3 (N2436, N2434, N362, N2204);
and AND2 (N2437, N2433, N545);
or OR4 (N2438, N2416, N1916, N689, N901);
or OR4 (N2439, N2419, N819, N1213, N2120);
not NOT1 (N2440, N2390);
buf BUF1 (N2441, N2440);
or OR3 (N2442, N2435, N2074, N2009);
nand NAND4 (N2443, N2442, N381, N2121, N1408);
buf BUF1 (N2444, N2443);
and AND3 (N2445, N2437, N1274, N9);
and AND4 (N2446, N2441, N2108, N729, N109);
xor XOR2 (N2447, N2444, N844);
nand NAND3 (N2448, N2439, N1312, N1427);
nor NOR4 (N2449, N2430, N142, N895, N849);
or OR4 (N2450, N2432, N1251, N943, N2009);
or OR2 (N2451, N2421, N1045);
xor XOR2 (N2452, N2445, N2365);
nand NAND2 (N2453, N2436, N1036);
and AND2 (N2454, N2453, N261);
nand NAND2 (N2455, N2438, N745);
nor NOR4 (N2456, N2450, N1800, N882, N122);
xor XOR2 (N2457, N2447, N264);
and AND4 (N2458, N2457, N1688, N1044, N346);
buf BUF1 (N2459, N2428);
nand NAND2 (N2460, N2449, N209);
nor NOR4 (N2461, N2456, N572, N2330, N2391);
nand NAND3 (N2462, N2452, N1769, N2381);
nor NOR3 (N2463, N2458, N1727, N2147);
buf BUF1 (N2464, N2455);
not NOT1 (N2465, N2461);
buf BUF1 (N2466, N2463);
nand NAND3 (N2467, N2451, N2093, N948);
xor XOR2 (N2468, N2467, N1963);
not NOT1 (N2469, N2454);
not NOT1 (N2470, N2448);
nor NOR2 (N2471, N2469, N824);
nor NOR3 (N2472, N2471, N851, N1422);
nor NOR2 (N2473, N2466, N1682);
xor XOR2 (N2474, N2473, N409);
buf BUF1 (N2475, N2460);
and AND3 (N2476, N2472, N520, N1985);
xor XOR2 (N2477, N2459, N935);
xor XOR2 (N2478, N2462, N2401);
not NOT1 (N2479, N2476);
xor XOR2 (N2480, N2465, N1979);
and AND4 (N2481, N2446, N1506, N1696, N96);
and AND4 (N2482, N2470, N1127, N851, N1035);
nor NOR3 (N2483, N2464, N75, N1873);
and AND4 (N2484, N2478, N1518, N1120, N71);
nand NAND2 (N2485, N2483, N1533);
or OR2 (N2486, N2485, N550);
buf BUF1 (N2487, N2477);
nand NAND4 (N2488, N2480, N609, N1138, N2063);
nand NAND3 (N2489, N2486, N1541, N193);
xor XOR2 (N2490, N2489, N1895);
nand NAND2 (N2491, N2468, N250);
nor NOR2 (N2492, N2474, N1805);
nor NOR3 (N2493, N2488, N2260, N705);
nand NAND2 (N2494, N2481, N1349);
nand NAND3 (N2495, N2487, N1627, N227);
xor XOR2 (N2496, N2484, N1701);
buf BUF1 (N2497, N2495);
not NOT1 (N2498, N2475);
nand NAND3 (N2499, N2490, N1281, N1957);
xor XOR2 (N2500, N2479, N39);
nor NOR2 (N2501, N2493, N2151);
not NOT1 (N2502, N2492);
buf BUF1 (N2503, N2497);
and AND3 (N2504, N2482, N1294, N1546);
not NOT1 (N2505, N2502);
not NOT1 (N2506, N2498);
not NOT1 (N2507, N2494);
xor XOR2 (N2508, N2505, N1740);
and AND2 (N2509, N2503, N1012);
or OR4 (N2510, N2509, N1068, N1923, N1217);
nor NOR2 (N2511, N2500, N120);
nand NAND4 (N2512, N2496, N2415, N356, N432);
not NOT1 (N2513, N2499);
and AND2 (N2514, N2513, N204);
nand NAND3 (N2515, N2506, N2083, N1961);
or OR2 (N2516, N2510, N1451);
nand NAND2 (N2517, N2512, N2386);
and AND2 (N2518, N2491, N1324);
xor XOR2 (N2519, N2507, N1997);
or OR2 (N2520, N2519, N1152);
xor XOR2 (N2521, N2516, N2044);
nand NAND2 (N2522, N2518, N841);
xor XOR2 (N2523, N2504, N908);
nor NOR3 (N2524, N2514, N677, N838);
nor NOR3 (N2525, N2501, N1797, N2026);
not NOT1 (N2526, N2520);
nand NAND2 (N2527, N2515, N1320);
nor NOR3 (N2528, N2508, N1797, N1347);
or OR2 (N2529, N2521, N282);
buf BUF1 (N2530, N2528);
buf BUF1 (N2531, N2511);
or OR4 (N2532, N2517, N133, N1463, N1838);
not NOT1 (N2533, N2523);
and AND2 (N2534, N2527, N760);
or OR2 (N2535, N2522, N395);
buf BUF1 (N2536, N2531);
nand NAND2 (N2537, N2535, N345);
nor NOR2 (N2538, N2536, N323);
nor NOR2 (N2539, N2538, N726);
xor XOR2 (N2540, N2533, N1054);
or OR4 (N2541, N2540, N1816, N1760, N1000);
nand NAND2 (N2542, N2524, N801);
buf BUF1 (N2543, N2532);
nor NOR2 (N2544, N2534, N1472);
not NOT1 (N2545, N2529);
and AND4 (N2546, N2543, N2373, N799, N317);
or OR4 (N2547, N2530, N984, N1588, N2384);
nor NOR4 (N2548, N2526, N1934, N709, N1381);
nor NOR2 (N2549, N2545, N1319);
or OR3 (N2550, N2539, N919, N402);
and AND4 (N2551, N2546, N2215, N1562, N90);
and AND2 (N2552, N2551, N2186);
nand NAND4 (N2553, N2548, N1573, N1469, N1546);
nand NAND2 (N2554, N2552, N1540);
or OR2 (N2555, N2537, N2458);
xor XOR2 (N2556, N2553, N467);
nor NOR3 (N2557, N2525, N306, N1906);
xor XOR2 (N2558, N2547, N1362);
not NOT1 (N2559, N2541);
not NOT1 (N2560, N2555);
and AND4 (N2561, N2557, N1239, N1093, N2152);
not NOT1 (N2562, N2544);
not NOT1 (N2563, N2558);
or OR2 (N2564, N2560, N2321);
and AND2 (N2565, N2554, N169);
and AND3 (N2566, N2549, N390, N2047);
nor NOR3 (N2567, N2556, N742, N2078);
xor XOR2 (N2568, N2542, N965);
nand NAND2 (N2569, N2564, N1861);
nand NAND4 (N2570, N2569, N95, N2016, N899);
nor NOR2 (N2571, N2563, N1575);
xor XOR2 (N2572, N2561, N342);
xor XOR2 (N2573, N2565, N2205);
and AND3 (N2574, N2562, N1860, N2448);
buf BUF1 (N2575, N2571);
or OR4 (N2576, N2567, N2179, N2156, N635);
xor XOR2 (N2577, N2566, N1820);
buf BUF1 (N2578, N2550);
nor NOR4 (N2579, N2573, N666, N1680, N175);
nand NAND3 (N2580, N2574, N1754, N897);
nor NOR4 (N2581, N2559, N357, N2080, N1574);
nor NOR3 (N2582, N2572, N251, N26);
nand NAND2 (N2583, N2575, N499);
nor NOR2 (N2584, N2578, N471);
not NOT1 (N2585, N2582);
or OR4 (N2586, N2580, N2460, N1568, N2468);
nor NOR2 (N2587, N2577, N1109);
and AND3 (N2588, N2579, N1801, N1326);
not NOT1 (N2589, N2584);
nor NOR2 (N2590, N2576, N258);
nand NAND3 (N2591, N2581, N847, N1787);
nor NOR2 (N2592, N2585, N1773);
buf BUF1 (N2593, N2570);
buf BUF1 (N2594, N2590);
not NOT1 (N2595, N2592);
and AND4 (N2596, N2587, N2512, N1924, N1056);
nor NOR2 (N2597, N2594, N1561);
buf BUF1 (N2598, N2591);
buf BUF1 (N2599, N2593);
xor XOR2 (N2600, N2568, N467);
or OR3 (N2601, N2586, N9, N850);
nor NOR3 (N2602, N2600, N2150, N534);
buf BUF1 (N2603, N2598);
nand NAND4 (N2604, N2596, N2246, N451, N1267);
nand NAND2 (N2605, N2602, N827);
not NOT1 (N2606, N2583);
nand NAND3 (N2607, N2597, N1775, N2130);
not NOT1 (N2608, N2603);
or OR2 (N2609, N2588, N98);
buf BUF1 (N2610, N2608);
buf BUF1 (N2611, N2604);
and AND4 (N2612, N2601, N1690, N1638, N951);
xor XOR2 (N2613, N2612, N399);
nor NOR4 (N2614, N2610, N851, N2097, N169);
buf BUF1 (N2615, N2605);
nand NAND3 (N2616, N2613, N1245, N827);
nor NOR2 (N2617, N2599, N952);
not NOT1 (N2618, N2606);
xor XOR2 (N2619, N2595, N1665);
nor NOR2 (N2620, N2611, N1768);
xor XOR2 (N2621, N2609, N2318);
and AND3 (N2622, N2617, N1932, N1146);
nand NAND2 (N2623, N2614, N2373);
nor NOR4 (N2624, N2623, N1840, N1158, N1322);
xor XOR2 (N2625, N2620, N2227);
and AND3 (N2626, N2622, N2122, N1036);
xor XOR2 (N2627, N2626, N2225);
nand NAND3 (N2628, N2624, N1552, N1939);
xor XOR2 (N2629, N2618, N2622);
buf BUF1 (N2630, N2616);
and AND2 (N2631, N2607, N1210);
or OR4 (N2632, N2619, N1311, N1358, N2086);
nand NAND4 (N2633, N2631, N1978, N1326, N1260);
xor XOR2 (N2634, N2627, N726);
nor NOR4 (N2635, N2625, N510, N1301, N1515);
xor XOR2 (N2636, N2629, N178);
not NOT1 (N2637, N2630);
buf BUF1 (N2638, N2633);
not NOT1 (N2639, N2615);
not NOT1 (N2640, N2628);
buf BUF1 (N2641, N2640);
or OR2 (N2642, N2636, N1373);
nor NOR2 (N2643, N2589, N2135);
and AND2 (N2644, N2634, N2268);
nor NOR4 (N2645, N2641, N1222, N1880, N681);
nand NAND2 (N2646, N2621, N1753);
buf BUF1 (N2647, N2639);
nand NAND4 (N2648, N2645, N2491, N2361, N1616);
or OR3 (N2649, N2643, N916, N2545);
or OR2 (N2650, N2646, N455);
buf BUF1 (N2651, N2632);
xor XOR2 (N2652, N2637, N1106);
buf BUF1 (N2653, N2652);
nor NOR4 (N2654, N2651, N947, N902, N2148);
buf BUF1 (N2655, N2648);
nor NOR2 (N2656, N2654, N1329);
xor XOR2 (N2657, N2644, N941);
buf BUF1 (N2658, N2655);
xor XOR2 (N2659, N2635, N648);
buf BUF1 (N2660, N2649);
nand NAND4 (N2661, N2658, N915, N255, N1205);
nor NOR2 (N2662, N2647, N1102);
nor NOR3 (N2663, N2650, N480, N1276);
and AND4 (N2664, N2663, N1314, N895, N1333);
xor XOR2 (N2665, N2642, N375);
not NOT1 (N2666, N2662);
xor XOR2 (N2667, N2653, N401);
and AND2 (N2668, N2666, N609);
not NOT1 (N2669, N2656);
nand NAND3 (N2670, N2668, N1726, N1962);
nor NOR3 (N2671, N2660, N2622, N856);
nor NOR2 (N2672, N2657, N1477);
or OR3 (N2673, N2669, N2032, N932);
buf BUF1 (N2674, N2661);
and AND3 (N2675, N2659, N1201, N1787);
and AND3 (N2676, N2665, N424, N2156);
nor NOR2 (N2677, N2676, N2111);
nor NOR2 (N2678, N2674, N2527);
nor NOR3 (N2679, N2677, N899, N2101);
or OR4 (N2680, N2679, N1770, N1920, N2580);
buf BUF1 (N2681, N2670);
nor NOR2 (N2682, N2672, N1093);
nor NOR4 (N2683, N2673, N1425, N948, N1727);
and AND4 (N2684, N2638, N433, N1586, N619);
not NOT1 (N2685, N2671);
nor NOR2 (N2686, N2664, N327);
or OR4 (N2687, N2686, N2365, N210, N2373);
not NOT1 (N2688, N2687);
and AND2 (N2689, N2667, N1331);
nand NAND3 (N2690, N2675, N227, N20);
nor NOR3 (N2691, N2689, N1728, N607);
nand NAND4 (N2692, N2680, N1320, N2589, N2665);
not NOT1 (N2693, N2692);
or OR3 (N2694, N2682, N2412, N1434);
nand NAND2 (N2695, N2678, N721);
buf BUF1 (N2696, N2691);
nor NOR3 (N2697, N2688, N1776, N1380);
not NOT1 (N2698, N2685);
and AND3 (N2699, N2681, N2111, N1471);
and AND4 (N2700, N2683, N1348, N516, N26);
not NOT1 (N2701, N2696);
and AND3 (N2702, N2700, N1410, N341);
nor NOR4 (N2703, N2695, N2463, N2300, N2685);
buf BUF1 (N2704, N2702);
xor XOR2 (N2705, N2699, N637);
nor NOR4 (N2706, N2705, N2423, N523, N1959);
nand NAND4 (N2707, N2701, N2385, N69, N526);
and AND3 (N2708, N2693, N1771, N482);
xor XOR2 (N2709, N2694, N1816);
xor XOR2 (N2710, N2708, N2678);
buf BUF1 (N2711, N2698);
and AND3 (N2712, N2709, N782, N556);
nand NAND2 (N2713, N2712, N2417);
not NOT1 (N2714, N2707);
or OR4 (N2715, N2690, N2383, N1325, N2486);
nand NAND3 (N2716, N2704, N1591, N452);
xor XOR2 (N2717, N2684, N48);
or OR3 (N2718, N2697, N1976, N2298);
buf BUF1 (N2719, N2711);
buf BUF1 (N2720, N2715);
xor XOR2 (N2721, N2718, N382);
or OR3 (N2722, N2710, N308, N255);
or OR3 (N2723, N2713, N415, N504);
and AND3 (N2724, N2719, N126, N18);
nor NOR3 (N2725, N2706, N1535, N145);
buf BUF1 (N2726, N2714);
xor XOR2 (N2727, N2716, N2059);
nand NAND4 (N2728, N2717, N1943, N1531, N2439);
and AND4 (N2729, N2727, N586, N2618, N2045);
and AND4 (N2730, N2723, N1392, N2360, N1585);
xor XOR2 (N2731, N2721, N24);
not NOT1 (N2732, N2720);
nor NOR3 (N2733, N2728, N1437, N922);
and AND4 (N2734, N2729, N535, N1839, N1982);
nand NAND3 (N2735, N2732, N158, N2330);
xor XOR2 (N2736, N2733, N2259);
buf BUF1 (N2737, N2735);
buf BUF1 (N2738, N2722);
nand NAND4 (N2739, N2738, N2111, N1050, N2264);
nand NAND4 (N2740, N2724, N1282, N2171, N1239);
and AND4 (N2741, N2703, N2548, N2098, N775);
nor NOR4 (N2742, N2726, N1408, N2318, N1395);
buf BUF1 (N2743, N2725);
nand NAND2 (N2744, N2736, N1366);
nor NOR3 (N2745, N2741, N303, N362);
nor NOR2 (N2746, N2740, N979);
nor NOR2 (N2747, N2744, N1556);
not NOT1 (N2748, N2739);
nor NOR2 (N2749, N2737, N2287);
xor XOR2 (N2750, N2745, N2455);
buf BUF1 (N2751, N2749);
not NOT1 (N2752, N2750);
or OR3 (N2753, N2751, N1346, N1948);
nor NOR4 (N2754, N2742, N1623, N2622, N614);
nand NAND3 (N2755, N2752, N1800, N2190);
buf BUF1 (N2756, N2755);
and AND2 (N2757, N2746, N898);
not NOT1 (N2758, N2743);
buf BUF1 (N2759, N2748);
or OR3 (N2760, N2758, N1153, N1860);
and AND2 (N2761, N2753, N2471);
nand NAND3 (N2762, N2754, N1851, N2370);
not NOT1 (N2763, N2756);
buf BUF1 (N2764, N2760);
not NOT1 (N2765, N2763);
buf BUF1 (N2766, N2762);
xor XOR2 (N2767, N2766, N134);
xor XOR2 (N2768, N2759, N1676);
not NOT1 (N2769, N2764);
not NOT1 (N2770, N2761);
nand NAND2 (N2771, N2757, N287);
and AND2 (N2772, N2765, N1487);
nand NAND2 (N2773, N2747, N2085);
and AND2 (N2774, N2731, N1967);
buf BUF1 (N2775, N2734);
nand NAND4 (N2776, N2773, N2288, N1458, N2082);
nor NOR4 (N2777, N2772, N2684, N1851, N1483);
xor XOR2 (N2778, N2770, N678);
not NOT1 (N2779, N2730);
xor XOR2 (N2780, N2777, N1155);
buf BUF1 (N2781, N2779);
buf BUF1 (N2782, N2771);
buf BUF1 (N2783, N2769);
not NOT1 (N2784, N2783);
xor XOR2 (N2785, N2780, N973);
and AND2 (N2786, N2767, N1252);
nand NAND3 (N2787, N2781, N1048, N1561);
buf BUF1 (N2788, N2776);
nor NOR4 (N2789, N2768, N769, N22, N809);
nand NAND3 (N2790, N2778, N974, N2103);
and AND4 (N2791, N2788, N1666, N392, N1621);
buf BUF1 (N2792, N2784);
not NOT1 (N2793, N2787);
not NOT1 (N2794, N2782);
nor NOR3 (N2795, N2794, N771, N2341);
and AND2 (N2796, N2792, N613);
not NOT1 (N2797, N2775);
buf BUF1 (N2798, N2785);
nor NOR2 (N2799, N2793, N506);
and AND4 (N2800, N2774, N366, N2580, N1003);
not NOT1 (N2801, N2795);
xor XOR2 (N2802, N2799, N880);
nand NAND2 (N2803, N2786, N2597);
nand NAND4 (N2804, N2789, N497, N1459, N1713);
xor XOR2 (N2805, N2803, N1122);
not NOT1 (N2806, N2800);
buf BUF1 (N2807, N2804);
not NOT1 (N2808, N2796);
nand NAND3 (N2809, N2808, N2697, N867);
nor NOR3 (N2810, N2805, N1458, N54);
and AND4 (N2811, N2810, N1457, N2473, N585);
and AND4 (N2812, N2791, N1911, N2635, N102);
or OR4 (N2813, N2798, N1001, N2281, N519);
xor XOR2 (N2814, N2807, N1979);
xor XOR2 (N2815, N2814, N2420);
xor XOR2 (N2816, N2790, N1337);
nor NOR3 (N2817, N2809, N1726, N1148);
nor NOR3 (N2818, N2811, N598, N1227);
and AND2 (N2819, N2812, N1459);
nor NOR2 (N2820, N2797, N2499);
nor NOR4 (N2821, N2818, N1455, N286, N2445);
nor NOR2 (N2822, N2817, N2798);
buf BUF1 (N2823, N2815);
and AND4 (N2824, N2813, N2793, N1240, N2582);
xor XOR2 (N2825, N2820, N2189);
xor XOR2 (N2826, N2806, N1996);
or OR4 (N2827, N2822, N2054, N1641, N1680);
xor XOR2 (N2828, N2802, N20);
nand NAND3 (N2829, N2826, N1198, N610);
nand NAND3 (N2830, N2819, N355, N878);
nand NAND2 (N2831, N2816, N1445);
not NOT1 (N2832, N2823);
and AND3 (N2833, N2825, N1091, N1724);
not NOT1 (N2834, N2833);
and AND2 (N2835, N2830, N2650);
nand NAND4 (N2836, N2835, N1975, N568, N581);
not NOT1 (N2837, N2834);
or OR2 (N2838, N2824, N80);
nand NAND3 (N2839, N2837, N1534, N1866);
not NOT1 (N2840, N2801);
xor XOR2 (N2841, N2827, N1943);
not NOT1 (N2842, N2829);
nand NAND2 (N2843, N2840, N106);
xor XOR2 (N2844, N2839, N2831);
xor XOR2 (N2845, N2602, N297);
nand NAND3 (N2846, N2828, N180, N1734);
and AND3 (N2847, N2845, N458, N1600);
and AND3 (N2848, N2846, N1794, N2180);
nor NOR2 (N2849, N2838, N1146);
xor XOR2 (N2850, N2836, N935);
xor XOR2 (N2851, N2847, N498);
nor NOR2 (N2852, N2832, N1088);
nand NAND3 (N2853, N2852, N1724, N2109);
xor XOR2 (N2854, N2821, N2317);
buf BUF1 (N2855, N2851);
nand NAND3 (N2856, N2855, N2744, N2825);
buf BUF1 (N2857, N2842);
xor XOR2 (N2858, N2844, N2630);
not NOT1 (N2859, N2853);
nand NAND2 (N2860, N2859, N1190);
or OR4 (N2861, N2848, N1013, N2415, N1862);
or OR2 (N2862, N2849, N2809);
nand NAND3 (N2863, N2843, N2114, N456);
xor XOR2 (N2864, N2850, N1773);
and AND2 (N2865, N2854, N2857);
nor NOR2 (N2866, N2554, N2346);
or OR3 (N2867, N2861, N997, N1395);
or OR2 (N2868, N2866, N247);
nand NAND4 (N2869, N2864, N1022, N553, N2268);
nand NAND4 (N2870, N2841, N1600, N51, N1280);
nand NAND3 (N2871, N2865, N1157, N1752);
buf BUF1 (N2872, N2863);
not NOT1 (N2873, N2867);
and AND2 (N2874, N2868, N1314);
and AND4 (N2875, N2862, N447, N1761, N830);
and AND4 (N2876, N2869, N2644, N2748, N418);
and AND2 (N2877, N2858, N2031);
and AND2 (N2878, N2872, N622);
or OR3 (N2879, N2870, N1812, N178);
and AND2 (N2880, N2875, N2235);
buf BUF1 (N2881, N2877);
buf BUF1 (N2882, N2876);
or OR3 (N2883, N2860, N2056, N2674);
not NOT1 (N2884, N2874);
nor NOR2 (N2885, N2856, N391);
or OR2 (N2886, N2873, N2484);
nor NOR3 (N2887, N2878, N214, N985);
nor NOR2 (N2888, N2887, N712);
xor XOR2 (N2889, N2884, N2328);
not NOT1 (N2890, N2881);
buf BUF1 (N2891, N2883);
nor NOR3 (N2892, N2891, N2747, N2685);
not NOT1 (N2893, N2892);
nand NAND3 (N2894, N2890, N1908, N1834);
nand NAND2 (N2895, N2885, N1184);
not NOT1 (N2896, N2880);
and AND2 (N2897, N2882, N2551);
nand NAND4 (N2898, N2893, N656, N609, N2245);
nor NOR3 (N2899, N2894, N1311, N2403);
not NOT1 (N2900, N2879);
not NOT1 (N2901, N2886);
xor XOR2 (N2902, N2889, N2220);
nand NAND4 (N2903, N2900, N1170, N1798, N2682);
not NOT1 (N2904, N2899);
nor NOR2 (N2905, N2895, N1103);
xor XOR2 (N2906, N2898, N1140);
nand NAND4 (N2907, N2901, N1908, N1531, N1403);
and AND4 (N2908, N2896, N1601, N2875, N142);
and AND3 (N2909, N2908, N311, N2837);
xor XOR2 (N2910, N2907, N2221);
nand NAND3 (N2911, N2897, N2409, N1933);
nand NAND4 (N2912, N2903, N2738, N18, N1187);
not NOT1 (N2913, N2902);
xor XOR2 (N2914, N2888, N288);
xor XOR2 (N2915, N2904, N2406);
nor NOR4 (N2916, N2915, N2743, N1016, N564);
and AND2 (N2917, N2911, N181);
and AND2 (N2918, N2906, N1944);
or OR4 (N2919, N2905, N2653, N2664, N1170);
buf BUF1 (N2920, N2909);
and AND4 (N2921, N2913, N490, N2791, N2222);
buf BUF1 (N2922, N2919);
xor XOR2 (N2923, N2916, N2641);
and AND3 (N2924, N2912, N2250, N689);
buf BUF1 (N2925, N2924);
and AND2 (N2926, N2918, N2229);
nand NAND4 (N2927, N2871, N1333, N199, N2857);
nand NAND4 (N2928, N2925, N2727, N2761, N2678);
xor XOR2 (N2929, N2923, N1362);
or OR4 (N2930, N2929, N1086, N2856, N1003);
not NOT1 (N2931, N2921);
nand NAND2 (N2932, N2920, N2375);
not NOT1 (N2933, N2928);
not NOT1 (N2934, N2922);
buf BUF1 (N2935, N2910);
nor NOR3 (N2936, N2917, N450, N2695);
xor XOR2 (N2937, N2934, N614);
nor NOR2 (N2938, N2931, N667);
nor NOR2 (N2939, N2926, N565);
nand NAND4 (N2940, N2938, N1601, N739, N369);
nor NOR2 (N2941, N2932, N1091);
nand NAND4 (N2942, N2941, N921, N2007, N2886);
or OR3 (N2943, N2933, N1032, N1942);
xor XOR2 (N2944, N2935, N2209);
nor NOR2 (N2945, N2943, N351);
or OR3 (N2946, N2936, N2528, N42);
or OR2 (N2947, N2940, N1757);
xor XOR2 (N2948, N2942, N1732);
buf BUF1 (N2949, N2939);
and AND4 (N2950, N2930, N2188, N864, N909);
nand NAND3 (N2951, N2947, N1342, N1315);
nor NOR2 (N2952, N2950, N452);
buf BUF1 (N2953, N2949);
or OR3 (N2954, N2944, N2319, N352);
xor XOR2 (N2955, N2945, N2339);
or OR2 (N2956, N2952, N644);
not NOT1 (N2957, N2953);
nand NAND2 (N2958, N2951, N2813);
nor NOR4 (N2959, N2948, N2474, N1021, N556);
nor NOR3 (N2960, N2957, N1723, N1356);
xor XOR2 (N2961, N2954, N2658);
not NOT1 (N2962, N2914);
and AND4 (N2963, N2946, N2422, N154, N1110);
and AND2 (N2964, N2963, N2491);
nor NOR3 (N2965, N2927, N614, N559);
nor NOR4 (N2966, N2962, N265, N2380, N1672);
or OR3 (N2967, N2937, N2141, N1233);
buf BUF1 (N2968, N2956);
nor NOR4 (N2969, N2958, N1386, N1732, N394);
nor NOR3 (N2970, N2969, N2606, N65);
xor XOR2 (N2971, N2967, N2030);
and AND3 (N2972, N2966, N1285, N1459);
nand NAND2 (N2973, N2964, N2235);
xor XOR2 (N2974, N2970, N187);
nand NAND3 (N2975, N2972, N1520, N593);
nor NOR2 (N2976, N2968, N2886);
buf BUF1 (N2977, N2959);
not NOT1 (N2978, N2961);
buf BUF1 (N2979, N2955);
not NOT1 (N2980, N2978);
nor NOR4 (N2981, N2976, N1945, N2888, N2751);
not NOT1 (N2982, N2981);
nor NOR3 (N2983, N2974, N2825, N1851);
nor NOR3 (N2984, N2960, N23, N873);
nand NAND2 (N2985, N2982, N2141);
nand NAND2 (N2986, N2965, N88);
nand NAND4 (N2987, N2979, N2323, N819, N109);
not NOT1 (N2988, N2987);
or OR2 (N2989, N2977, N1536);
and AND4 (N2990, N2988, N2458, N1511, N607);
or OR4 (N2991, N2985, N449, N1461, N2087);
buf BUF1 (N2992, N2971);
or OR4 (N2993, N2975, N2386, N2371, N1188);
buf BUF1 (N2994, N2973);
and AND2 (N2995, N2983, N2739);
or OR2 (N2996, N2995, N1125);
nand NAND2 (N2997, N2993, N2936);
buf BUF1 (N2998, N2996);
not NOT1 (N2999, N2998);
or OR4 (N3000, N2980, N255, N707, N971);
or OR3 (N3001, N2992, N1382, N1478);
buf BUF1 (N3002, N2999);
and AND2 (N3003, N2997, N1457);
or OR4 (N3004, N3000, N1659, N1629, N2635);
not NOT1 (N3005, N3003);
and AND2 (N3006, N2984, N1866);
xor XOR2 (N3007, N3004, N2692);
and AND2 (N3008, N3005, N415);
not NOT1 (N3009, N2991);
or OR4 (N3010, N3009, N624, N82, N1640);
nor NOR4 (N3011, N3008, N200, N1034, N1709);
xor XOR2 (N3012, N3001, N1205);
nor NOR4 (N3013, N3010, N1755, N2518, N2734);
xor XOR2 (N3014, N2986, N845);
nor NOR4 (N3015, N2989, N2100, N1865, N127);
xor XOR2 (N3016, N3002, N2358);
not NOT1 (N3017, N3006);
nor NOR4 (N3018, N3013, N1986, N2060, N313);
not NOT1 (N3019, N3017);
and AND2 (N3020, N2990, N191);
nor NOR2 (N3021, N3016, N1045);
or OR2 (N3022, N3015, N366);
or OR4 (N3023, N3020, N513, N2060, N890);
xor XOR2 (N3024, N3023, N2867);
not NOT1 (N3025, N3012);
nand NAND3 (N3026, N3022, N362, N96);
nor NOR3 (N3027, N3019, N1435, N2271);
xor XOR2 (N3028, N3007, N2428);
buf BUF1 (N3029, N3028);
buf BUF1 (N3030, N3018);
or OR2 (N3031, N3029, N1478);
and AND3 (N3032, N3014, N2572, N91);
and AND4 (N3033, N3030, N2747, N1241, N80);
xor XOR2 (N3034, N2994, N1412);
buf BUF1 (N3035, N3031);
xor XOR2 (N3036, N3026, N55);
nor NOR2 (N3037, N3021, N2788);
nand NAND4 (N3038, N3034, N244, N2337, N545);
nor NOR3 (N3039, N3025, N2459, N2194);
buf BUF1 (N3040, N3039);
not NOT1 (N3041, N3033);
not NOT1 (N3042, N3036);
nand NAND3 (N3043, N3037, N2521, N1358);
nor NOR3 (N3044, N3027, N43, N2480);
or OR2 (N3045, N3040, N2365);
or OR4 (N3046, N3032, N1127, N1647, N1067);
buf BUF1 (N3047, N3044);
and AND3 (N3048, N3011, N1633, N2576);
xor XOR2 (N3049, N3042, N1335);
and AND3 (N3050, N3046, N2705, N2893);
or OR3 (N3051, N3038, N1457, N22);
nor NOR4 (N3052, N3024, N1055, N786, N2757);
nand NAND2 (N3053, N3035, N1086);
nor NOR3 (N3054, N3045, N198, N2252);
xor XOR2 (N3055, N3052, N1657);
xor XOR2 (N3056, N3049, N801);
not NOT1 (N3057, N3056);
and AND3 (N3058, N3053, N2497, N2404);
nand NAND2 (N3059, N3051, N1479);
xor XOR2 (N3060, N3047, N1929);
not NOT1 (N3061, N3060);
buf BUF1 (N3062, N3041);
and AND2 (N3063, N3043, N2764);
nand NAND3 (N3064, N3063, N1708, N907);
buf BUF1 (N3065, N3059);
buf BUF1 (N3066, N3065);
and AND3 (N3067, N3058, N2309, N1001);
nor NOR2 (N3068, N3048, N118);
not NOT1 (N3069, N3062);
or OR4 (N3070, N3050, N2888, N1316, N1307);
and AND2 (N3071, N3066, N2158);
or OR2 (N3072, N3057, N714);
xor XOR2 (N3073, N3055, N2574);
not NOT1 (N3074, N3069);
nor NOR4 (N3075, N3072, N1349, N2005, N1080);
and AND4 (N3076, N3074, N1747, N1043, N1071);
buf BUF1 (N3077, N3067);
xor XOR2 (N3078, N3068, N1629);
and AND3 (N3079, N3076, N1353, N376);
nor NOR2 (N3080, N3079, N1501);
buf BUF1 (N3081, N3075);
and AND4 (N3082, N3080, N207, N1944, N2224);
and AND2 (N3083, N3070, N2275);
nor NOR2 (N3084, N3064, N1558);
and AND3 (N3085, N3083, N696, N2609);
or OR3 (N3086, N3085, N1172, N1916);
nand NAND2 (N3087, N3084, N1371);
or OR4 (N3088, N3071, N2477, N1584, N2968);
xor XOR2 (N3089, N3054, N2583);
or OR3 (N3090, N3087, N2142, N1717);
or OR2 (N3091, N3090, N467);
and AND2 (N3092, N3078, N2898);
and AND2 (N3093, N3091, N2139);
or OR4 (N3094, N3073, N1745, N1164, N274);
nor NOR2 (N3095, N3081, N2081);
nand NAND4 (N3096, N3093, N2549, N574, N2592);
buf BUF1 (N3097, N3094);
not NOT1 (N3098, N3077);
buf BUF1 (N3099, N3086);
not NOT1 (N3100, N3097);
nand NAND2 (N3101, N3099, N1593);
or OR2 (N3102, N3101, N243);
nand NAND3 (N3103, N3082, N1767, N2671);
or OR4 (N3104, N3102, N2485, N924, N2898);
or OR2 (N3105, N3092, N1324);
or OR2 (N3106, N3096, N275);
nor NOR3 (N3107, N3105, N3092, N1955);
nor NOR3 (N3108, N3106, N910, N2054);
and AND2 (N3109, N3095, N2013);
buf BUF1 (N3110, N3098);
nand NAND4 (N3111, N3110, N1377, N173, N384);
buf BUF1 (N3112, N3111);
nor NOR4 (N3113, N3103, N181, N2908, N2462);
and AND4 (N3114, N3104, N325, N10, N802);
and AND4 (N3115, N3112, N76, N1574, N1991);
or OR2 (N3116, N3109, N417);
nor NOR4 (N3117, N3116, N832, N1798, N2548);
not NOT1 (N3118, N3113);
xor XOR2 (N3119, N3118, N1001);
nor NOR2 (N3120, N3119, N1102);
xor XOR2 (N3121, N3117, N62);
nand NAND3 (N3122, N3115, N135, N1256);
xor XOR2 (N3123, N3088, N1456);
buf BUF1 (N3124, N3114);
not NOT1 (N3125, N3120);
not NOT1 (N3126, N3061);
or OR3 (N3127, N3122, N2095, N1925);
nor NOR2 (N3128, N3100, N2328);
xor XOR2 (N3129, N3128, N2937);
and AND2 (N3130, N3121, N1376);
buf BUF1 (N3131, N3124);
or OR4 (N3132, N3125, N2785, N407, N132);
xor XOR2 (N3133, N3108, N2364);
and AND4 (N3134, N3107, N1029, N125, N2804);
nand NAND4 (N3135, N3129, N2112, N516, N783);
nor NOR2 (N3136, N3123, N349);
not NOT1 (N3137, N3127);
nand NAND3 (N3138, N3134, N1749, N1560);
nor NOR3 (N3139, N3133, N2839, N2880);
or OR2 (N3140, N3136, N1994);
and AND3 (N3141, N3140, N914, N766);
and AND4 (N3142, N3130, N1958, N2592, N834);
and AND4 (N3143, N3137, N2960, N860, N2102);
not NOT1 (N3144, N3142);
buf BUF1 (N3145, N3132);
nor NOR4 (N3146, N3145, N2395, N362, N2649);
and AND2 (N3147, N3144, N1624);
nand NAND2 (N3148, N3147, N2831);
or OR2 (N3149, N3143, N422);
xor XOR2 (N3150, N3131, N2746);
and AND4 (N3151, N3141, N2356, N2183, N616);
nor NOR3 (N3152, N3151, N1115, N2822);
nand NAND4 (N3153, N3089, N2365, N842, N1711);
not NOT1 (N3154, N3150);
not NOT1 (N3155, N3138);
or OR4 (N3156, N3155, N2511, N858, N381);
nand NAND3 (N3157, N3149, N183, N329);
xor XOR2 (N3158, N3148, N1309);
nor NOR2 (N3159, N3152, N507);
nand NAND2 (N3160, N3158, N2799);
and AND2 (N3161, N3126, N2964);
xor XOR2 (N3162, N3159, N2091);
or OR2 (N3163, N3154, N1248);
buf BUF1 (N3164, N3153);
xor XOR2 (N3165, N3156, N887);
nand NAND3 (N3166, N3161, N2370, N623);
nand NAND4 (N3167, N3139, N2909, N2392, N1044);
not NOT1 (N3168, N3164);
not NOT1 (N3169, N3157);
nor NOR3 (N3170, N3163, N3009, N2921);
and AND2 (N3171, N3169, N670);
not NOT1 (N3172, N3167);
not NOT1 (N3173, N3171);
xor XOR2 (N3174, N3146, N1872);
nor NOR2 (N3175, N3160, N2774);
and AND4 (N3176, N3168, N698, N2453, N2202);
not NOT1 (N3177, N3172);
nor NOR2 (N3178, N3174, N2350);
not NOT1 (N3179, N3170);
xor XOR2 (N3180, N3178, N1575);
buf BUF1 (N3181, N3173);
nand NAND2 (N3182, N3176, N143);
nor NOR3 (N3183, N3180, N262, N1641);
nor NOR3 (N3184, N3166, N2464, N500);
nor NOR2 (N3185, N3181, N2131);
or OR4 (N3186, N3165, N2215, N1430, N2003);
xor XOR2 (N3187, N3184, N1800);
not NOT1 (N3188, N3135);
or OR2 (N3189, N3177, N1397);
nand NAND3 (N3190, N3162, N215, N2865);
buf BUF1 (N3191, N3187);
buf BUF1 (N3192, N3190);
or OR4 (N3193, N3175, N1142, N288, N2781);
or OR3 (N3194, N3183, N313, N2479);
and AND2 (N3195, N3189, N3061);
not NOT1 (N3196, N3188);
not NOT1 (N3197, N3191);
nand NAND2 (N3198, N3182, N1465);
and AND2 (N3199, N3193, N941);
nor NOR3 (N3200, N3197, N556, N2713);
buf BUF1 (N3201, N3200);
xor XOR2 (N3202, N3201, N2137);
or OR4 (N3203, N3199, N1051, N14, N130);
xor XOR2 (N3204, N3195, N789);
nand NAND3 (N3205, N3192, N1364, N3186);
nand NAND4 (N3206, N2622, N917, N181, N1697);
xor XOR2 (N3207, N3196, N2453);
xor XOR2 (N3208, N3185, N100);
buf BUF1 (N3209, N3206);
and AND3 (N3210, N3179, N1643, N2913);
and AND4 (N3211, N3209, N482, N343, N245);
or OR4 (N3212, N3204, N2298, N184, N379);
not NOT1 (N3213, N3207);
not NOT1 (N3214, N3213);
nand NAND3 (N3215, N3208, N421, N1883);
nor NOR2 (N3216, N3205, N904);
not NOT1 (N3217, N3214);
xor XOR2 (N3218, N3198, N2078);
or OR4 (N3219, N3202, N1285, N1622, N1571);
or OR4 (N3220, N3216, N485, N1584, N1544);
nor NOR4 (N3221, N3215, N3098, N1325, N2228);
not NOT1 (N3222, N3217);
not NOT1 (N3223, N3218);
xor XOR2 (N3224, N3203, N1111);
and AND3 (N3225, N3222, N3209, N178);
or OR2 (N3226, N3212, N475);
nand NAND4 (N3227, N3224, N1532, N2600, N2775);
and AND4 (N3228, N3211, N543, N2418, N2546);
buf BUF1 (N3229, N3219);
nor NOR2 (N3230, N3228, N2508);
or OR4 (N3231, N3220, N476, N1756, N1687);
xor XOR2 (N3232, N3225, N2403);
or OR2 (N3233, N3226, N1181);
buf BUF1 (N3234, N3230);
nor NOR3 (N3235, N3194, N2081, N1942);
xor XOR2 (N3236, N3231, N777);
nor NOR4 (N3237, N3229, N2003, N1575, N1972);
and AND2 (N3238, N3221, N1465);
not NOT1 (N3239, N3237);
nand NAND4 (N3240, N3232, N1283, N1337, N264);
nand NAND2 (N3241, N3223, N3046);
xor XOR2 (N3242, N3240, N1740);
or OR4 (N3243, N3234, N2511, N2026, N1287);
nand NAND4 (N3244, N3210, N3163, N2816, N3101);
buf BUF1 (N3245, N3233);
xor XOR2 (N3246, N3239, N2634);
and AND3 (N3247, N3243, N472, N3179);
and AND4 (N3248, N3235, N2601, N389, N1781);
nand NAND3 (N3249, N3244, N126, N807);
and AND3 (N3250, N3245, N1307, N433);
nor NOR4 (N3251, N3246, N2377, N1250, N2848);
not NOT1 (N3252, N3247);
nand NAND2 (N3253, N3227, N1992);
nor NOR4 (N3254, N3236, N2122, N254, N2405);
buf BUF1 (N3255, N3252);
nor NOR3 (N3256, N3250, N1345, N752);
nand NAND4 (N3257, N3255, N1337, N1442, N3038);
nand NAND4 (N3258, N3254, N869, N1015, N1293);
not NOT1 (N3259, N3257);
buf BUF1 (N3260, N3242);
and AND2 (N3261, N3260, N2907);
buf BUF1 (N3262, N3261);
and AND2 (N3263, N3262, N2908);
buf BUF1 (N3264, N3259);
and AND4 (N3265, N3251, N1309, N1727, N776);
xor XOR2 (N3266, N3238, N2471);
nor NOR4 (N3267, N3263, N3191, N29, N825);
not NOT1 (N3268, N3256);
xor XOR2 (N3269, N3268, N1827);
nand NAND4 (N3270, N3266, N1955, N1851, N1928);
nor NOR4 (N3271, N3249, N1279, N25, N884);
or OR4 (N3272, N3269, N1423, N498, N188);
or OR3 (N3273, N3253, N2352, N519);
nor NOR3 (N3274, N3270, N1121, N3239);
buf BUF1 (N3275, N3248);
not NOT1 (N3276, N3274);
or OR3 (N3277, N3271, N1083, N2321);
not NOT1 (N3278, N3275);
not NOT1 (N3279, N3258);
buf BUF1 (N3280, N3279);
not NOT1 (N3281, N3278);
nand NAND2 (N3282, N3273, N1839);
and AND3 (N3283, N3272, N1486, N1805);
or OR4 (N3284, N3276, N2445, N1972, N3175);
nor NOR3 (N3285, N3241, N2281, N979);
nand NAND3 (N3286, N3267, N1106, N3000);
or OR4 (N3287, N3280, N297, N2864, N488);
not NOT1 (N3288, N3285);
not NOT1 (N3289, N3265);
xor XOR2 (N3290, N3286, N165);
nor NOR4 (N3291, N3264, N2113, N726, N1626);
nor NOR3 (N3292, N3290, N2691, N2589);
nor NOR4 (N3293, N3282, N2443, N1332, N1101);
not NOT1 (N3294, N3287);
xor XOR2 (N3295, N3277, N2454);
or OR2 (N3296, N3283, N2991);
or OR3 (N3297, N3292, N1999, N2580);
nor NOR4 (N3298, N3288, N2406, N194, N115);
not NOT1 (N3299, N3284);
or OR3 (N3300, N3291, N1886, N2555);
nand NAND4 (N3301, N3300, N3116, N605, N1490);
buf BUF1 (N3302, N3289);
not NOT1 (N3303, N3299);
or OR4 (N3304, N3294, N1607, N695, N2716);
xor XOR2 (N3305, N3301, N1110);
nand NAND3 (N3306, N3295, N868, N946);
and AND2 (N3307, N3305, N2900);
and AND4 (N3308, N3297, N340, N1636, N307);
or OR4 (N3309, N3306, N215, N1020, N406);
not NOT1 (N3310, N3298);
not NOT1 (N3311, N3307);
buf BUF1 (N3312, N3311);
nand NAND3 (N3313, N3303, N2701, N2162);
buf BUF1 (N3314, N3304);
and AND2 (N3315, N3310, N2398);
nor NOR3 (N3316, N3302, N2107, N496);
and AND2 (N3317, N3316, N911);
xor XOR2 (N3318, N3296, N2631);
xor XOR2 (N3319, N3317, N2491);
buf BUF1 (N3320, N3308);
nand NAND3 (N3321, N3312, N1624, N1199);
nor NOR4 (N3322, N3281, N1835, N1689, N2198);
or OR4 (N3323, N3319, N2817, N2245, N1634);
buf BUF1 (N3324, N3318);
and AND2 (N3325, N3313, N1269);
xor XOR2 (N3326, N3321, N262);
nand NAND4 (N3327, N3293, N911, N1116, N342);
not NOT1 (N3328, N3323);
nand NAND3 (N3329, N3327, N630, N91);
nor NOR4 (N3330, N3324, N246, N1691, N875);
not NOT1 (N3331, N3329);
nor NOR4 (N3332, N3314, N2247, N311, N2579);
nand NAND3 (N3333, N3325, N1078, N1322);
or OR3 (N3334, N3326, N950, N2163);
or OR4 (N3335, N3332, N2947, N708, N1898);
nor NOR2 (N3336, N3309, N437);
or OR4 (N3337, N3334, N3221, N1864, N3077);
and AND4 (N3338, N3335, N2555, N810, N1978);
buf BUF1 (N3339, N3336);
nor NOR3 (N3340, N3315, N1030, N466);
or OR2 (N3341, N3320, N1828);
xor XOR2 (N3342, N3340, N1539);
and AND4 (N3343, N3339, N1997, N408, N3324);
nor NOR4 (N3344, N3322, N909, N2655, N2378);
nand NAND2 (N3345, N3342, N2169);
and AND3 (N3346, N3343, N3088, N1485);
xor XOR2 (N3347, N3328, N2281);
or OR2 (N3348, N3333, N1057);
not NOT1 (N3349, N3348);
buf BUF1 (N3350, N3337);
not NOT1 (N3351, N3345);
or OR3 (N3352, N3338, N570, N757);
buf BUF1 (N3353, N3331);
xor XOR2 (N3354, N3344, N2305);
nand NAND3 (N3355, N3353, N2257, N1716);
xor XOR2 (N3356, N3341, N1150);
nand NAND4 (N3357, N3354, N1535, N1, N391);
or OR2 (N3358, N3351, N178);
nor NOR2 (N3359, N3357, N1971);
nand NAND4 (N3360, N3352, N3132, N1864, N3023);
xor XOR2 (N3361, N3360, N1677);
or OR4 (N3362, N3355, N1920, N2243, N2276);
or OR2 (N3363, N3359, N119);
nor NOR3 (N3364, N3330, N2482, N2960);
xor XOR2 (N3365, N3347, N2394);
and AND3 (N3366, N3361, N2730, N1132);
or OR2 (N3367, N3366, N2387);
and AND3 (N3368, N3365, N549, N1325);
and AND4 (N3369, N3346, N1321, N1399, N373);
buf BUF1 (N3370, N3356);
nand NAND4 (N3371, N3363, N1116, N42, N1889);
and AND4 (N3372, N3371, N819, N1347, N919);
xor XOR2 (N3373, N3362, N814);
not NOT1 (N3374, N3358);
nand NAND2 (N3375, N3349, N3300);
xor XOR2 (N3376, N3370, N2698);
and AND4 (N3377, N3369, N2476, N376, N178);
or OR3 (N3378, N3372, N1023, N2220);
or OR4 (N3379, N3376, N1883, N399, N2864);
nor NOR2 (N3380, N3374, N1773);
not NOT1 (N3381, N3375);
buf BUF1 (N3382, N3373);
or OR2 (N3383, N3379, N72);
buf BUF1 (N3384, N3381);
buf BUF1 (N3385, N3377);
xor XOR2 (N3386, N3367, N999);
not NOT1 (N3387, N3350);
or OR4 (N3388, N3384, N949, N2108, N2220);
xor XOR2 (N3389, N3387, N490);
and AND3 (N3390, N3382, N2823, N2955);
not NOT1 (N3391, N3380);
nor NOR2 (N3392, N3383, N647);
xor XOR2 (N3393, N3389, N1785);
xor XOR2 (N3394, N3391, N630);
nor NOR2 (N3395, N3378, N2291);
and AND2 (N3396, N3390, N2641);
or OR2 (N3397, N3392, N2299);
buf BUF1 (N3398, N3394);
buf BUF1 (N3399, N3397);
nor NOR4 (N3400, N3386, N2709, N1547, N419);
or OR2 (N3401, N3396, N857);
not NOT1 (N3402, N3364);
xor XOR2 (N3403, N3402, N89);
nand NAND4 (N3404, N3385, N1413, N3175, N2675);
or OR3 (N3405, N3395, N8, N1249);
nand NAND3 (N3406, N3393, N3137, N661);
xor XOR2 (N3407, N3405, N1898);
or OR2 (N3408, N3398, N2833);
nand NAND4 (N3409, N3406, N1562, N1096, N709);
and AND2 (N3410, N3407, N2478);
nand NAND2 (N3411, N3401, N1170);
nand NAND2 (N3412, N3388, N51);
nor NOR3 (N3413, N3403, N3048, N2905);
not NOT1 (N3414, N3410);
not NOT1 (N3415, N3414);
xor XOR2 (N3416, N3412, N747);
nor NOR3 (N3417, N3413, N2456, N2431);
not NOT1 (N3418, N3415);
and AND4 (N3419, N3400, N2033, N2094, N675);
or OR2 (N3420, N3411, N1746);
nand NAND3 (N3421, N3418, N1316, N860);
nor NOR4 (N3422, N3420, N2508, N2416, N1750);
nand NAND2 (N3423, N3417, N444);
buf BUF1 (N3424, N3421);
or OR4 (N3425, N3422, N1321, N7, N2209);
buf BUF1 (N3426, N3423);
nor NOR4 (N3427, N3425, N1904, N2895, N2834);
or OR2 (N3428, N3408, N2397);
xor XOR2 (N3429, N3424, N779);
nand NAND2 (N3430, N3409, N3302);
nor NOR4 (N3431, N3416, N1332, N525, N3176);
not NOT1 (N3432, N3399);
nand NAND4 (N3433, N3432, N1939, N922, N518);
or OR4 (N3434, N3368, N2700, N2263, N1372);
or OR2 (N3435, N3427, N2047);
nand NAND4 (N3436, N3429, N2741, N216, N1449);
or OR3 (N3437, N3419, N2714, N3064);
nor NOR3 (N3438, N3431, N2349, N1627);
xor XOR2 (N3439, N3430, N1967);
xor XOR2 (N3440, N3437, N2296);
or OR4 (N3441, N3433, N318, N3015, N1613);
or OR4 (N3442, N3428, N2088, N2918, N1977);
xor XOR2 (N3443, N3438, N3168);
and AND3 (N3444, N3435, N2748, N3045);
or OR2 (N3445, N3434, N2599);
buf BUF1 (N3446, N3441);
nor NOR2 (N3447, N3442, N881);
and AND2 (N3448, N3436, N1226);
and AND3 (N3449, N3443, N1783, N1740);
buf BUF1 (N3450, N3439);
nand NAND4 (N3451, N3445, N3363, N1942, N831);
nor NOR3 (N3452, N3446, N250, N1045);
buf BUF1 (N3453, N3447);
xor XOR2 (N3454, N3451, N362);
buf BUF1 (N3455, N3448);
or OR4 (N3456, N3444, N2852, N244, N2470);
xor XOR2 (N3457, N3404, N1546);
nor NOR3 (N3458, N3449, N2052, N1966);
buf BUF1 (N3459, N3457);
or OR3 (N3460, N3458, N530, N3339);
or OR4 (N3461, N3426, N2619, N1921, N2553);
xor XOR2 (N3462, N3456, N2535);
buf BUF1 (N3463, N3455);
and AND2 (N3464, N3454, N3134);
or OR2 (N3465, N3440, N2059);
buf BUF1 (N3466, N3464);
nor NOR4 (N3467, N3466, N685, N1734, N2972);
nor NOR2 (N3468, N3450, N1460);
or OR2 (N3469, N3463, N3200);
not NOT1 (N3470, N3461);
or OR4 (N3471, N3462, N3196, N1382, N525);
or OR2 (N3472, N3468, N444);
nor NOR3 (N3473, N3452, N1009, N2219);
nor NOR4 (N3474, N3465, N2312, N1107, N991);
xor XOR2 (N3475, N3470, N1999);
and AND2 (N3476, N3475, N199);
buf BUF1 (N3477, N3476);
buf BUF1 (N3478, N3471);
buf BUF1 (N3479, N3478);
buf BUF1 (N3480, N3460);
or OR4 (N3481, N3453, N3064, N898, N199);
not NOT1 (N3482, N3480);
buf BUF1 (N3483, N3472);
xor XOR2 (N3484, N3467, N2617);
and AND2 (N3485, N3477, N1752);
nand NAND3 (N3486, N3484, N1389, N1540);
nor NOR4 (N3487, N3469, N869, N402, N778);
nand NAND2 (N3488, N3486, N768);
xor XOR2 (N3489, N3473, N898);
not NOT1 (N3490, N3485);
xor XOR2 (N3491, N3482, N2534);
or OR2 (N3492, N3474, N1219);
and AND2 (N3493, N3490, N2605);
not NOT1 (N3494, N3479);
or OR2 (N3495, N3489, N2837);
nand NAND2 (N3496, N3483, N450);
or OR2 (N3497, N3494, N353);
or OR4 (N3498, N3496, N3217, N1875, N3197);
xor XOR2 (N3499, N3498, N3093);
xor XOR2 (N3500, N3492, N3449);
nor NOR3 (N3501, N3481, N2174, N1052);
nor NOR2 (N3502, N3500, N2292);
nand NAND4 (N3503, N3459, N1665, N1223, N49);
nor NOR4 (N3504, N3497, N1045, N1299, N2712);
nand NAND2 (N3505, N3504, N3278);
buf BUF1 (N3506, N3487);
or OR3 (N3507, N3499, N1556, N1196);
buf BUF1 (N3508, N3503);
nor NOR4 (N3509, N3501, N715, N2348, N1114);
and AND4 (N3510, N3502, N2274, N3073, N1797);
buf BUF1 (N3511, N3495);
or OR2 (N3512, N3510, N1569);
not NOT1 (N3513, N3509);
or OR3 (N3514, N3507, N421, N2280);
and AND4 (N3515, N3511, N2651, N995, N486);
nand NAND4 (N3516, N3515, N1200, N935, N1261);
nor NOR3 (N3517, N3488, N586, N1382);
nor NOR3 (N3518, N3506, N3498, N3195);
nand NAND2 (N3519, N3491, N544);
or OR4 (N3520, N3516, N83, N515, N349);
nor NOR3 (N3521, N3493, N3078, N2414);
nand NAND4 (N3522, N3521, N1061, N3284, N3497);
buf BUF1 (N3523, N3517);
xor XOR2 (N3524, N3505, N239);
xor XOR2 (N3525, N3513, N57);
xor XOR2 (N3526, N3519, N1653);
nor NOR3 (N3527, N3520, N14, N184);
not NOT1 (N3528, N3508);
and AND4 (N3529, N3522, N1065, N2871, N1184);
or OR2 (N3530, N3524, N1656);
buf BUF1 (N3531, N3528);
buf BUF1 (N3532, N3518);
buf BUF1 (N3533, N3530);
and AND3 (N3534, N3533, N307, N797);
nand NAND4 (N3535, N3514, N1335, N1695, N2471);
or OR4 (N3536, N3531, N383, N1452, N1647);
or OR2 (N3537, N3534, N3259);
nor NOR2 (N3538, N3535, N1521);
not NOT1 (N3539, N3512);
and AND2 (N3540, N3536, N2751);
or OR2 (N3541, N3539, N1116);
or OR3 (N3542, N3541, N2005, N680);
nand NAND4 (N3543, N3526, N405, N580, N1921);
xor XOR2 (N3544, N3532, N465);
xor XOR2 (N3545, N3540, N3051);
nand NAND2 (N3546, N3527, N258);
or OR4 (N3547, N3543, N3362, N1629, N2715);
not NOT1 (N3548, N3544);
and AND3 (N3549, N3545, N690, N1384);
nand NAND4 (N3550, N3525, N666, N1562, N1818);
or OR2 (N3551, N3550, N1799);
not NOT1 (N3552, N3551);
and AND4 (N3553, N3529, N3340, N31, N2915);
nor NOR3 (N3554, N3548, N225, N138);
xor XOR2 (N3555, N3547, N2726);
buf BUF1 (N3556, N3537);
and AND3 (N3557, N3556, N1811, N758);
nand NAND2 (N3558, N3538, N2032);
xor XOR2 (N3559, N3549, N1696);
xor XOR2 (N3560, N3557, N1356);
nand NAND3 (N3561, N3546, N1099, N182);
nor NOR4 (N3562, N3552, N1687, N1511, N290);
xor XOR2 (N3563, N3562, N670);
nand NAND3 (N3564, N3553, N2479, N3340);
buf BUF1 (N3565, N3561);
xor XOR2 (N3566, N3560, N1192);
not NOT1 (N3567, N3523);
not NOT1 (N3568, N3558);
nand NAND2 (N3569, N3542, N1063);
nor NOR3 (N3570, N3568, N2840, N964);
not NOT1 (N3571, N3563);
and AND2 (N3572, N3559, N3047);
buf BUF1 (N3573, N3554);
and AND4 (N3574, N3555, N2482, N671, N231);
xor XOR2 (N3575, N3565, N1510);
nand NAND4 (N3576, N3572, N3363, N3433, N286);
xor XOR2 (N3577, N3576, N582);
not NOT1 (N3578, N3577);
nor NOR3 (N3579, N3574, N2649, N2941);
buf BUF1 (N3580, N3564);
or OR2 (N3581, N3567, N1306);
buf BUF1 (N3582, N3580);
or OR3 (N3583, N3579, N3515, N1135);
and AND2 (N3584, N3566, N2190);
or OR4 (N3585, N3571, N1263, N1124, N2687);
not NOT1 (N3586, N3583);
nor NOR3 (N3587, N3586, N602, N1853);
xor XOR2 (N3588, N3584, N1893);
nand NAND2 (N3589, N3578, N2293);
nor NOR3 (N3590, N3588, N1638, N2663);
xor XOR2 (N3591, N3569, N458);
buf BUF1 (N3592, N3575);
buf BUF1 (N3593, N3591);
not NOT1 (N3594, N3582);
nand NAND2 (N3595, N3587, N229);
nor NOR2 (N3596, N3570, N2128);
nor NOR3 (N3597, N3595, N2930, N3280);
xor XOR2 (N3598, N3594, N1683);
buf BUF1 (N3599, N3589);
nor NOR2 (N3600, N3597, N1073);
not NOT1 (N3601, N3596);
nand NAND2 (N3602, N3581, N70);
xor XOR2 (N3603, N3592, N3543);
or OR2 (N3604, N3603, N1803);
and AND2 (N3605, N3601, N1126);
nand NAND3 (N3606, N3604, N877, N1888);
not NOT1 (N3607, N3606);
xor XOR2 (N3608, N3573, N1641);
or OR2 (N3609, N3602, N535);
buf BUF1 (N3610, N3593);
and AND4 (N3611, N3600, N1001, N1192, N160);
nand NAND4 (N3612, N3585, N3355, N3594, N2940);
nor NOR3 (N3613, N3599, N1832, N483);
and AND2 (N3614, N3598, N2869);
nor NOR3 (N3615, N3605, N78, N2583);
and AND4 (N3616, N3590, N1940, N333, N2711);
nand NAND4 (N3617, N3613, N1468, N1413, N2038);
nor NOR4 (N3618, N3617, N886, N1269, N1858);
not NOT1 (N3619, N3610);
buf BUF1 (N3620, N3607);
buf BUF1 (N3621, N3611);
nand NAND3 (N3622, N3619, N411, N1821);
nand NAND2 (N3623, N3616, N2499);
nor NOR4 (N3624, N3621, N2204, N726, N2849);
or OR4 (N3625, N3623, N986, N1326, N1853);
nand NAND4 (N3626, N3620, N758, N487, N2562);
xor XOR2 (N3627, N3614, N389);
not NOT1 (N3628, N3625);
or OR4 (N3629, N3618, N3516, N964, N682);
or OR2 (N3630, N3622, N525);
and AND4 (N3631, N3615, N578, N1738, N3630);
nor NOR2 (N3632, N1307, N934);
xor XOR2 (N3633, N3628, N755);
xor XOR2 (N3634, N3631, N3582);
nand NAND2 (N3635, N3634, N1380);
and AND4 (N3636, N3633, N2796, N949, N2141);
or OR4 (N3637, N3612, N720, N9, N99);
not NOT1 (N3638, N3629);
nor NOR2 (N3639, N3609, N2078);
not NOT1 (N3640, N3635);
not NOT1 (N3641, N3624);
nor NOR2 (N3642, N3627, N2334);
xor XOR2 (N3643, N3632, N1493);
not NOT1 (N3644, N3626);
or OR3 (N3645, N3644, N453, N2989);
nor NOR3 (N3646, N3645, N2901, N3054);
and AND3 (N3647, N3638, N2563, N1821);
buf BUF1 (N3648, N3642);
buf BUF1 (N3649, N3639);
nor NOR3 (N3650, N3636, N2276, N1510);
and AND4 (N3651, N3637, N1162, N1426, N2532);
nand NAND4 (N3652, N3643, N357, N172, N81);
xor XOR2 (N3653, N3646, N1374);
nand NAND4 (N3654, N3652, N2130, N3118, N3593);
or OR2 (N3655, N3654, N2222);
not NOT1 (N3656, N3648);
xor XOR2 (N3657, N3650, N2296);
or OR2 (N3658, N3608, N948);
and AND4 (N3659, N3653, N682, N1171, N2118);
or OR2 (N3660, N3641, N74);
nand NAND4 (N3661, N3656, N1486, N2058, N1489);
and AND3 (N3662, N3658, N3538, N102);
and AND2 (N3663, N3660, N1425);
and AND3 (N3664, N3659, N125, N459);
or OR2 (N3665, N3663, N677);
and AND4 (N3666, N3662, N1998, N1899, N1113);
xor XOR2 (N3667, N3665, N2075);
xor XOR2 (N3668, N3640, N355);
and AND3 (N3669, N3649, N632, N557);
nor NOR4 (N3670, N3668, N3487, N1567, N760);
not NOT1 (N3671, N3664);
xor XOR2 (N3672, N3669, N2468);
nor NOR4 (N3673, N3667, N3206, N2351, N3592);
nor NOR4 (N3674, N3666, N1874, N372, N2089);
nor NOR3 (N3675, N3672, N1312, N2381);
nand NAND2 (N3676, N3651, N597);
nand NAND4 (N3677, N3670, N2396, N2133, N2421);
or OR2 (N3678, N3675, N2185);
xor XOR2 (N3679, N3655, N1353);
buf BUF1 (N3680, N3677);
nand NAND4 (N3681, N3647, N1323, N2831, N434);
not NOT1 (N3682, N3680);
nor NOR2 (N3683, N3673, N461);
buf BUF1 (N3684, N3679);
buf BUF1 (N3685, N3684);
buf BUF1 (N3686, N3661);
nand NAND2 (N3687, N3681, N3325);
nand NAND2 (N3688, N3685, N2957);
nand NAND2 (N3689, N3678, N2384);
buf BUF1 (N3690, N3689);
not NOT1 (N3691, N3674);
and AND3 (N3692, N3688, N2264, N149);
not NOT1 (N3693, N3692);
buf BUF1 (N3694, N3657);
xor XOR2 (N3695, N3671, N3001);
xor XOR2 (N3696, N3687, N3023);
or OR4 (N3697, N3695, N1756, N405, N2011);
nand NAND2 (N3698, N3693, N111);
buf BUF1 (N3699, N3697);
and AND2 (N3700, N3691, N2838);
nand NAND3 (N3701, N3694, N2020, N2247);
or OR3 (N3702, N3700, N2796, N3039);
buf BUF1 (N3703, N3701);
xor XOR2 (N3704, N3703, N1941);
not NOT1 (N3705, N3702);
xor XOR2 (N3706, N3698, N2844);
or OR4 (N3707, N3699, N1419, N1298, N441);
not NOT1 (N3708, N3706);
xor XOR2 (N3709, N3704, N3215);
buf BUF1 (N3710, N3696);
and AND2 (N3711, N3683, N2622);
and AND3 (N3712, N3710, N380, N3212);
nor NOR3 (N3713, N3686, N743, N2429);
nand NAND2 (N3714, N3708, N250);
nand NAND2 (N3715, N3705, N3288);
buf BUF1 (N3716, N3712);
not NOT1 (N3717, N3713);
nand NAND4 (N3718, N3716, N1279, N168, N3582);
or OR2 (N3719, N3707, N2554);
nor NOR2 (N3720, N3718, N3280);
not NOT1 (N3721, N3690);
and AND3 (N3722, N3714, N1899, N223);
xor XOR2 (N3723, N3719, N3041);
xor XOR2 (N3724, N3682, N235);
nor NOR3 (N3725, N3717, N3402, N3227);
nand NAND4 (N3726, N3711, N979, N3350, N65);
and AND2 (N3727, N3722, N1066);
nor NOR3 (N3728, N3721, N931, N446);
xor XOR2 (N3729, N3725, N433);
nor NOR4 (N3730, N3729, N1773, N1607, N3650);
buf BUF1 (N3731, N3724);
xor XOR2 (N3732, N3723, N3304);
or OR2 (N3733, N3727, N535);
nand NAND3 (N3734, N3676, N3721, N1036);
or OR4 (N3735, N3709, N1657, N3576, N2789);
or OR2 (N3736, N3732, N3513);
nor NOR4 (N3737, N3720, N2410, N1237, N941);
not NOT1 (N3738, N3715);
xor XOR2 (N3739, N3726, N2835);
or OR2 (N3740, N3733, N2664);
xor XOR2 (N3741, N3736, N1023);
xor XOR2 (N3742, N3731, N1774);
xor XOR2 (N3743, N3739, N2089);
nand NAND3 (N3744, N3741, N3179, N1103);
or OR3 (N3745, N3738, N389, N1353);
nor NOR3 (N3746, N3745, N2457, N919);
xor XOR2 (N3747, N3734, N1010);
buf BUF1 (N3748, N3742);
buf BUF1 (N3749, N3747);
buf BUF1 (N3750, N3728);
nor NOR4 (N3751, N3740, N2584, N585, N1713);
buf BUF1 (N3752, N3743);
not NOT1 (N3753, N3749);
buf BUF1 (N3754, N3751);
and AND4 (N3755, N3752, N322, N154, N266);
buf BUF1 (N3756, N3754);
buf BUF1 (N3757, N3737);
and AND4 (N3758, N3757, N3597, N1961, N2042);
xor XOR2 (N3759, N3755, N42);
nor NOR2 (N3760, N3759, N9);
xor XOR2 (N3761, N3760, N2027);
and AND2 (N3762, N3748, N2189);
xor XOR2 (N3763, N3753, N3668);
or OR3 (N3764, N3756, N1633, N54);
not NOT1 (N3765, N3763);
xor XOR2 (N3766, N3746, N1692);
not NOT1 (N3767, N3761);
buf BUF1 (N3768, N3765);
buf BUF1 (N3769, N3764);
not NOT1 (N3770, N3730);
nand NAND4 (N3771, N3767, N2264, N677, N3552);
buf BUF1 (N3772, N3771);
buf BUF1 (N3773, N3770);
or OR2 (N3774, N3762, N1997);
xor XOR2 (N3775, N3750, N1333);
and AND2 (N3776, N3774, N1413);
nand NAND4 (N3777, N3766, N2803, N2776, N3379);
nand NAND3 (N3778, N3758, N485, N1053);
or OR3 (N3779, N3778, N979, N226);
or OR4 (N3780, N3775, N1082, N3038, N2092);
not NOT1 (N3781, N3769);
or OR3 (N3782, N3776, N2644, N683);
nor NOR3 (N3783, N3768, N2082, N650);
xor XOR2 (N3784, N3783, N3161);
and AND3 (N3785, N3782, N135, N556);
not NOT1 (N3786, N3735);
buf BUF1 (N3787, N3785);
xor XOR2 (N3788, N3786, N1535);
nand NAND3 (N3789, N3784, N1806, N2946);
or OR2 (N3790, N3773, N2180);
nor NOR2 (N3791, N3780, N230);
buf BUF1 (N3792, N3777);
and AND3 (N3793, N3787, N871, N2477);
nand NAND2 (N3794, N3792, N3633);
and AND4 (N3795, N3744, N546, N668, N3047);
nor NOR2 (N3796, N3772, N3069);
or OR4 (N3797, N3788, N3194, N2166, N326);
or OR4 (N3798, N3779, N2811, N1465, N1506);
not NOT1 (N3799, N3796);
not NOT1 (N3800, N3799);
nand NAND3 (N3801, N3781, N336, N2810);
nor NOR2 (N3802, N3789, N14);
nor NOR2 (N3803, N3795, N3025);
not NOT1 (N3804, N3802);
buf BUF1 (N3805, N3793);
nand NAND3 (N3806, N3798, N1290, N420);
xor XOR2 (N3807, N3794, N1976);
buf BUF1 (N3808, N3803);
or OR2 (N3809, N3807, N488);
or OR4 (N3810, N3805, N2948, N611, N717);
and AND4 (N3811, N3809, N2470, N2437, N1127);
not NOT1 (N3812, N3806);
xor XOR2 (N3813, N3808, N1615);
and AND3 (N3814, N3811, N60, N203);
not NOT1 (N3815, N3800);
and AND4 (N3816, N3815, N2727, N3, N45);
buf BUF1 (N3817, N3804);
or OR4 (N3818, N3817, N788, N1458, N2130);
buf BUF1 (N3819, N3816);
and AND2 (N3820, N3797, N2800);
or OR4 (N3821, N3820, N3800, N2462, N2029);
nand NAND4 (N3822, N3812, N3229, N1616, N1713);
buf BUF1 (N3823, N3819);
nand NAND4 (N3824, N3791, N3480, N815, N2064);
nor NOR4 (N3825, N3810, N2722, N549, N951);
nor NOR2 (N3826, N3813, N287);
buf BUF1 (N3827, N3818);
not NOT1 (N3828, N3825);
not NOT1 (N3829, N3824);
buf BUF1 (N3830, N3790);
or OR3 (N3831, N3827, N2696, N1183);
or OR2 (N3832, N3814, N545);
or OR3 (N3833, N3829, N2219, N3628);
nor NOR2 (N3834, N3832, N1502);
and AND2 (N3835, N3833, N3731);
not NOT1 (N3836, N3801);
and AND4 (N3837, N3836, N673, N2105, N2784);
nor NOR3 (N3838, N3830, N610, N1558);
nor NOR3 (N3839, N3838, N48, N3559);
xor XOR2 (N3840, N3828, N3079);
nor NOR2 (N3841, N3821, N2745);
nor NOR2 (N3842, N3839, N1004);
nor NOR4 (N3843, N3840, N3048, N3778, N3595);
buf BUF1 (N3844, N3837);
buf BUF1 (N3845, N3841);
nor NOR2 (N3846, N3822, N1797);
xor XOR2 (N3847, N3843, N70);
nand NAND3 (N3848, N3842, N3219, N105);
and AND3 (N3849, N3826, N180, N969);
and AND2 (N3850, N3835, N1206);
not NOT1 (N3851, N3849);
nor NOR3 (N3852, N3851, N1899, N2238);
nor NOR2 (N3853, N3845, N836);
and AND3 (N3854, N3852, N2820, N1447);
buf BUF1 (N3855, N3823);
and AND3 (N3856, N3850, N1716, N2848);
nand NAND4 (N3857, N3854, N2922, N3852, N1476);
or OR4 (N3858, N3847, N2952, N3339, N821);
nor NOR4 (N3859, N3834, N2652, N114, N1233);
xor XOR2 (N3860, N3857, N1181);
buf BUF1 (N3861, N3844);
buf BUF1 (N3862, N3861);
nand NAND2 (N3863, N3860, N2275);
xor XOR2 (N3864, N3856, N3688);
and AND2 (N3865, N3862, N1865);
nor NOR3 (N3866, N3864, N2912, N2617);
or OR4 (N3867, N3846, N1286, N2301, N2527);
buf BUF1 (N3868, N3865);
buf BUF1 (N3869, N3848);
and AND2 (N3870, N3863, N749);
or OR3 (N3871, N3866, N325, N2680);
not NOT1 (N3872, N3869);
not NOT1 (N3873, N3872);
nand NAND3 (N3874, N3853, N67, N1555);
not NOT1 (N3875, N3858);
not NOT1 (N3876, N3873);
and AND4 (N3877, N3876, N2608, N1036, N3781);
not NOT1 (N3878, N3831);
nand NAND2 (N3879, N3878, N1780);
buf BUF1 (N3880, N3879);
nor NOR3 (N3881, N3871, N1760, N3864);
or OR2 (N3882, N3867, N2454);
nand NAND3 (N3883, N3877, N2748, N2081);
buf BUF1 (N3884, N3881);
and AND2 (N3885, N3870, N2397);
nor NOR2 (N3886, N3859, N2411);
nor NOR2 (N3887, N3855, N1985);
xor XOR2 (N3888, N3883, N3477);
xor XOR2 (N3889, N3888, N1275);
not NOT1 (N3890, N3886);
xor XOR2 (N3891, N3884, N537);
buf BUF1 (N3892, N3875);
nand NAND2 (N3893, N3887, N15);
and AND3 (N3894, N3889, N2113, N1238);
nand NAND2 (N3895, N3894, N3698);
nand NAND2 (N3896, N3892, N2226);
xor XOR2 (N3897, N3880, N480);
buf BUF1 (N3898, N3895);
or OR2 (N3899, N3897, N2654);
and AND2 (N3900, N3891, N2863);
nand NAND4 (N3901, N3898, N319, N3630, N3443);
nand NAND3 (N3902, N3868, N1463, N1027);
nor NOR4 (N3903, N3900, N2121, N303, N174);
xor XOR2 (N3904, N3890, N259);
nand NAND2 (N3905, N3882, N1709);
nand NAND4 (N3906, N3896, N2988, N595, N1096);
and AND3 (N3907, N3901, N2810, N251);
xor XOR2 (N3908, N3905, N2944);
xor XOR2 (N3909, N3908, N3674);
nand NAND3 (N3910, N3899, N482, N3733);
not NOT1 (N3911, N3903);
buf BUF1 (N3912, N3874);
xor XOR2 (N3913, N3893, N3226);
xor XOR2 (N3914, N3910, N1830);
and AND3 (N3915, N3904, N3150, N1895);
buf BUF1 (N3916, N3907);
nor NOR3 (N3917, N3913, N3404, N2787);
xor XOR2 (N3918, N3917, N3630);
xor XOR2 (N3919, N3885, N3861);
and AND2 (N3920, N3909, N2625);
buf BUF1 (N3921, N3906);
or OR3 (N3922, N3902, N2978, N2014);
and AND2 (N3923, N3916, N937);
and AND4 (N3924, N3915, N330, N1110, N3745);
nand NAND2 (N3925, N3911, N1073);
xor XOR2 (N3926, N3922, N2029);
and AND4 (N3927, N3918, N2570, N3213, N1304);
and AND3 (N3928, N3914, N2109, N1169);
buf BUF1 (N3929, N3919);
or OR3 (N3930, N3920, N1296, N3898);
or OR4 (N3931, N3925, N1143, N1831, N907);
and AND4 (N3932, N3928, N2152, N1011, N3693);
and AND2 (N3933, N3927, N3082);
and AND2 (N3934, N3933, N3559);
nor NOR3 (N3935, N3932, N1147, N1616);
and AND3 (N3936, N3930, N3676, N1546);
buf BUF1 (N3937, N3936);
and AND4 (N3938, N3931, N3330, N2637, N2766);
xor XOR2 (N3939, N3938, N467);
nand NAND2 (N3940, N3939, N1395);
not NOT1 (N3941, N3912);
buf BUF1 (N3942, N3923);
or OR3 (N3943, N3929, N2129, N1707);
not NOT1 (N3944, N3934);
nor NOR4 (N3945, N3924, N2747, N3691, N1843);
nor NOR3 (N3946, N3921, N2848, N960);
buf BUF1 (N3947, N3926);
or OR2 (N3948, N3940, N1061);
or OR4 (N3949, N3948, N448, N374, N73);
or OR4 (N3950, N3941, N774, N3513, N1664);
nor NOR4 (N3951, N3942, N894, N1814, N3687);
nand NAND3 (N3952, N3944, N1790, N538);
xor XOR2 (N3953, N3945, N2335);
not NOT1 (N3954, N3952);
nand NAND3 (N3955, N3946, N1835, N1970);
nor NOR3 (N3956, N3951, N3512, N97);
buf BUF1 (N3957, N3954);
or OR2 (N3958, N3956, N2639);
nor NOR3 (N3959, N3955, N1769, N1987);
nand NAND2 (N3960, N3947, N1153);
and AND3 (N3961, N3953, N2560, N96);
and AND2 (N3962, N3937, N573);
buf BUF1 (N3963, N3961);
xor XOR2 (N3964, N3959, N2699);
xor XOR2 (N3965, N3960, N1404);
not NOT1 (N3966, N3943);
and AND2 (N3967, N3957, N2831);
not NOT1 (N3968, N3949);
buf BUF1 (N3969, N3935);
xor XOR2 (N3970, N3966, N617);
buf BUF1 (N3971, N3950);
nand NAND2 (N3972, N3958, N1734);
or OR3 (N3973, N3965, N2679, N3639);
or OR4 (N3974, N3963, N3282, N1619, N2347);
buf BUF1 (N3975, N3964);
nor NOR4 (N3976, N3974, N1381, N2171, N3223);
nand NAND3 (N3977, N3973, N1026, N1487);
not NOT1 (N3978, N3975);
and AND2 (N3979, N3969, N810);
xor XOR2 (N3980, N3979, N3672);
xor XOR2 (N3981, N3970, N2595);
not NOT1 (N3982, N3977);
or OR3 (N3983, N3967, N1628, N3562);
buf BUF1 (N3984, N3982);
and AND4 (N3985, N3983, N182, N87, N2073);
xor XOR2 (N3986, N3976, N1967);
not NOT1 (N3987, N3978);
not NOT1 (N3988, N3971);
nor NOR3 (N3989, N3985, N1496, N3075);
and AND3 (N3990, N3984, N1490, N1004);
buf BUF1 (N3991, N3972);
or OR4 (N3992, N3987, N1783, N901, N1640);
or OR4 (N3993, N3992, N2597, N1243, N2605);
not NOT1 (N3994, N3968);
or OR3 (N3995, N3990, N1291, N2538);
buf BUF1 (N3996, N3991);
buf BUF1 (N3997, N3980);
nand NAND4 (N3998, N3986, N1016, N974, N1414);
xor XOR2 (N3999, N3981, N3192);
nand NAND4 (N4000, N3996, N465, N702, N813);
and AND4 (N4001, N3994, N2404, N4, N1804);
buf BUF1 (N4002, N3988);
or OR3 (N4003, N3995, N1737, N614);
not NOT1 (N4004, N4002);
and AND4 (N4005, N3993, N601, N2265, N1033);
xor XOR2 (N4006, N3989, N3077);
not NOT1 (N4007, N4006);
nor NOR2 (N4008, N4004, N3754);
xor XOR2 (N4009, N3962, N2369);
not NOT1 (N4010, N4008);
or OR3 (N4011, N4007, N2441, N2207);
nor NOR4 (N4012, N3999, N3694, N3946, N664);
not NOT1 (N4013, N4005);
xor XOR2 (N4014, N4011, N3216);
buf BUF1 (N4015, N3997);
and AND4 (N4016, N4015, N3055, N1243, N86);
buf BUF1 (N4017, N4012);
not NOT1 (N4018, N4000);
not NOT1 (N4019, N4003);
and AND4 (N4020, N4009, N3686, N3754, N1702);
nor NOR4 (N4021, N4001, N3473, N3669, N1082);
nor NOR4 (N4022, N4016, N3604, N622, N1491);
not NOT1 (N4023, N4020);
not NOT1 (N4024, N4014);
nand NAND4 (N4025, N4013, N23, N1930, N1176);
or OR3 (N4026, N4019, N2528, N1375);
and AND3 (N4027, N4010, N2838, N2428);
buf BUF1 (N4028, N4027);
nor NOR2 (N4029, N4023, N3068);
buf BUF1 (N4030, N4028);
not NOT1 (N4031, N4030);
buf BUF1 (N4032, N3998);
or OR2 (N4033, N4017, N733);
buf BUF1 (N4034, N4018);
xor XOR2 (N4035, N4034, N2440);
nand NAND4 (N4036, N4022, N1141, N2084, N1169);
or OR3 (N4037, N4032, N1970, N498);
nor NOR4 (N4038, N4021, N1478, N3194, N3952);
buf BUF1 (N4039, N4038);
nand NAND2 (N4040, N4035, N2154);
and AND2 (N4041, N4037, N3291);
nand NAND4 (N4042, N4040, N1873, N3339, N341);
not NOT1 (N4043, N4031);
nand NAND3 (N4044, N4042, N2922, N3004);
and AND3 (N4045, N4039, N11, N826);
nor NOR4 (N4046, N4029, N3943, N3357, N2032);
buf BUF1 (N4047, N4046);
nand NAND3 (N4048, N4036, N528, N877);
buf BUF1 (N4049, N4033);
or OR4 (N4050, N4026, N1323, N3069, N1028);
nor NOR4 (N4051, N4044, N3050, N3894, N2800);
and AND4 (N4052, N4045, N2987, N3062, N2010);
xor XOR2 (N4053, N4051, N1951);
or OR3 (N4054, N4050, N372, N2098);
and AND3 (N4055, N4052, N3036, N514);
or OR4 (N4056, N4055, N2084, N527, N882);
not NOT1 (N4057, N4047);
and AND2 (N4058, N4025, N1761);
not NOT1 (N4059, N4058);
nand NAND2 (N4060, N4024, N2599);
xor XOR2 (N4061, N4041, N683);
not NOT1 (N4062, N4054);
not NOT1 (N4063, N4059);
or OR4 (N4064, N4053, N2925, N2140, N1739);
not NOT1 (N4065, N4063);
or OR4 (N4066, N4043, N3989, N2332, N1995);
not NOT1 (N4067, N4066);
not NOT1 (N4068, N4062);
not NOT1 (N4069, N4068);
nor NOR2 (N4070, N4064, N158);
nor NOR4 (N4071, N4056, N1448, N1787, N1634);
buf BUF1 (N4072, N4069);
buf BUF1 (N4073, N4065);
xor XOR2 (N4074, N4057, N2305);
xor XOR2 (N4075, N4074, N4038);
not NOT1 (N4076, N4060);
and AND4 (N4077, N4049, N36, N3506, N2622);
xor XOR2 (N4078, N4071, N1572);
buf BUF1 (N4079, N4072);
xor XOR2 (N4080, N4079, N3665);
nand NAND3 (N4081, N4048, N2140, N2351);
or OR4 (N4082, N4080, N3130, N2252, N1543);
nor NOR2 (N4083, N4076, N228);
nor NOR4 (N4084, N4073, N3716, N3626, N1132);
and AND4 (N4085, N4075, N207, N950, N3263);
not NOT1 (N4086, N4067);
and AND2 (N4087, N4085, N3177);
and AND3 (N4088, N4078, N1923, N3398);
xor XOR2 (N4089, N4070, N1728);
xor XOR2 (N4090, N4077, N1120);
buf BUF1 (N4091, N4086);
buf BUF1 (N4092, N4088);
xor XOR2 (N4093, N4089, N285);
and AND4 (N4094, N4084, N3529, N3242, N3807);
nand NAND3 (N4095, N4091, N3681, N483);
xor XOR2 (N4096, N4090, N2640);
nand NAND4 (N4097, N4087, N851, N1177, N77);
not NOT1 (N4098, N4094);
buf BUF1 (N4099, N4061);
or OR4 (N4100, N4082, N2591, N3113, N3757);
and AND3 (N4101, N4081, N2783, N1150);
nor NOR4 (N4102, N4095, N1169, N1718, N3446);
not NOT1 (N4103, N4099);
buf BUF1 (N4104, N4092);
and AND4 (N4105, N4103, N1803, N2253, N1144);
xor XOR2 (N4106, N4102, N1071);
nor NOR2 (N4107, N4083, N1583);
not NOT1 (N4108, N4106);
buf BUF1 (N4109, N4105);
and AND2 (N4110, N4104, N1372);
not NOT1 (N4111, N4100);
and AND2 (N4112, N4111, N3949);
and AND2 (N4113, N4098, N2004);
nand NAND2 (N4114, N4097, N1201);
nor NOR4 (N4115, N4093, N2560, N1059, N1738);
buf BUF1 (N4116, N4114);
nand NAND4 (N4117, N4107, N2698, N1246, N1539);
not NOT1 (N4118, N4108);
buf BUF1 (N4119, N4109);
not NOT1 (N4120, N4115);
or OR2 (N4121, N4120, N2514);
nor NOR4 (N4122, N4118, N1271, N1826, N362);
not NOT1 (N4123, N4122);
buf BUF1 (N4124, N4121);
nor NOR4 (N4125, N4110, N585, N3843, N2769);
and AND2 (N4126, N4116, N3090);
or OR3 (N4127, N4117, N245, N2482);
not NOT1 (N4128, N4127);
xor XOR2 (N4129, N4113, N277);
xor XOR2 (N4130, N4112, N635);
and AND2 (N4131, N4126, N3674);
buf BUF1 (N4132, N4128);
or OR2 (N4133, N4130, N1823);
nor NOR3 (N4134, N4131, N1387, N3321);
xor XOR2 (N4135, N4125, N3771);
nand NAND2 (N4136, N4119, N541);
or OR4 (N4137, N4133, N1161, N870, N221);
and AND2 (N4138, N4101, N966);
or OR2 (N4139, N4096, N1669);
or OR2 (N4140, N4137, N3443);
or OR4 (N4141, N4139, N153, N352, N1713);
nand NAND2 (N4142, N4138, N1182);
or OR2 (N4143, N4136, N2596);
nor NOR2 (N4144, N4129, N3280);
xor XOR2 (N4145, N4143, N3758);
not NOT1 (N4146, N4135);
buf BUF1 (N4147, N4123);
nor NOR3 (N4148, N4146, N3692, N3541);
nand NAND2 (N4149, N4144, N513);
nand NAND4 (N4150, N4141, N1716, N3884, N3505);
or OR2 (N4151, N4148, N2889);
xor XOR2 (N4152, N4124, N2123);
nor NOR4 (N4153, N4132, N3054, N1159, N128);
nor NOR4 (N4154, N4134, N2417, N2423, N34);
not NOT1 (N4155, N4150);
nand NAND4 (N4156, N4145, N1563, N887, N3159);
or OR2 (N4157, N4149, N3167);
not NOT1 (N4158, N4142);
nand NAND4 (N4159, N4152, N3467, N2106, N1916);
xor XOR2 (N4160, N4153, N3296);
xor XOR2 (N4161, N4155, N4044);
nor NOR2 (N4162, N4161, N569);
not NOT1 (N4163, N4140);
nand NAND2 (N4164, N4154, N2615);
not NOT1 (N4165, N4163);
not NOT1 (N4166, N4165);
or OR3 (N4167, N4164, N2854, N3676);
and AND4 (N4168, N4160, N3902, N1031, N1350);
and AND2 (N4169, N4157, N3233);
not NOT1 (N4170, N4168);
buf BUF1 (N4171, N4159);
nand NAND2 (N4172, N4151, N3724);
xor XOR2 (N4173, N4166, N1283);
xor XOR2 (N4174, N4171, N1697);
nand NAND4 (N4175, N4167, N2840, N7, N214);
nand NAND2 (N4176, N4173, N1043);
buf BUF1 (N4177, N4175);
buf BUF1 (N4178, N4169);
nand NAND2 (N4179, N4158, N1235);
or OR3 (N4180, N4178, N535, N4173);
and AND2 (N4181, N4172, N3146);
buf BUF1 (N4182, N4179);
not NOT1 (N4183, N4180);
buf BUF1 (N4184, N4177);
xor XOR2 (N4185, N4162, N2786);
xor XOR2 (N4186, N4184, N3765);
nor NOR4 (N4187, N4170, N1113, N3473, N818);
xor XOR2 (N4188, N4186, N2556);
xor XOR2 (N4189, N4182, N3822);
nand NAND3 (N4190, N4188, N232, N1274);
xor XOR2 (N4191, N4185, N566);
buf BUF1 (N4192, N4190);
nand NAND3 (N4193, N4192, N1143, N30);
nor NOR3 (N4194, N4191, N2205, N1268);
nor NOR2 (N4195, N4181, N1560);
not NOT1 (N4196, N4174);
xor XOR2 (N4197, N4176, N2457);
nand NAND2 (N4198, N4197, N1388);
nand NAND4 (N4199, N4187, N1749, N2319, N1204);
or OR2 (N4200, N4194, N2008);
nand NAND4 (N4201, N4147, N955, N13, N572);
xor XOR2 (N4202, N4199, N3297);
or OR4 (N4203, N4195, N1582, N2980, N709);
buf BUF1 (N4204, N4189);
xor XOR2 (N4205, N4183, N4128);
or OR4 (N4206, N4156, N695, N3087, N4125);
not NOT1 (N4207, N4193);
not NOT1 (N4208, N4207);
and AND3 (N4209, N4206, N1041, N3383);
nor NOR4 (N4210, N4204, N3099, N422, N2051);
and AND4 (N4211, N4196, N197, N134, N4203);
nand NAND2 (N4212, N3681, N4201);
xor XOR2 (N4213, N973, N162);
nor NOR3 (N4214, N4202, N4164, N1495);
and AND3 (N4215, N4208, N3158, N975);
and AND2 (N4216, N4210, N2165);
not NOT1 (N4217, N4209);
xor XOR2 (N4218, N4214, N4132);
xor XOR2 (N4219, N4212, N606);
buf BUF1 (N4220, N4211);
nor NOR3 (N4221, N4215, N73, N2883);
not NOT1 (N4222, N4220);
nand NAND3 (N4223, N4213, N1184, N577);
and AND4 (N4224, N4200, N3410, N1702, N3071);
nand NAND3 (N4225, N4223, N2550, N329);
buf BUF1 (N4226, N4219);
buf BUF1 (N4227, N4226);
buf BUF1 (N4228, N4227);
nand NAND4 (N4229, N4218, N2543, N2342, N2303);
nor NOR4 (N4230, N4229, N629, N2319, N1077);
not NOT1 (N4231, N4198);
not NOT1 (N4232, N4225);
not NOT1 (N4233, N4222);
buf BUF1 (N4234, N4231);
not NOT1 (N4235, N4228);
xor XOR2 (N4236, N4232, N2073);
nand NAND2 (N4237, N4221, N1845);
buf BUF1 (N4238, N4237);
not NOT1 (N4239, N4230);
xor XOR2 (N4240, N4205, N7);
xor XOR2 (N4241, N4236, N3159);
nand NAND3 (N4242, N4240, N1168, N3085);
xor XOR2 (N4243, N4238, N567);
nand NAND2 (N4244, N4239, N2254);
buf BUF1 (N4245, N4224);
nor NOR3 (N4246, N4244, N1529, N1947);
buf BUF1 (N4247, N4235);
nor NOR3 (N4248, N4216, N828, N3588);
nand NAND3 (N4249, N4242, N3351, N3674);
not NOT1 (N4250, N4233);
buf BUF1 (N4251, N4250);
nor NOR3 (N4252, N4241, N2852, N4038);
buf BUF1 (N4253, N4243);
nand NAND2 (N4254, N4251, N447);
buf BUF1 (N4255, N4234);
nor NOR3 (N4256, N4217, N1021, N623);
or OR3 (N4257, N4254, N4172, N4246);
or OR2 (N4258, N2221, N2335);
and AND3 (N4259, N4252, N655, N2939);
nor NOR4 (N4260, N4258, N1048, N1135, N1414);
xor XOR2 (N4261, N4253, N1053);
or OR4 (N4262, N4257, N1654, N3578, N3700);
xor XOR2 (N4263, N4247, N1248);
and AND3 (N4264, N4261, N1266, N3402);
buf BUF1 (N4265, N4264);
and AND2 (N4266, N4248, N2300);
not NOT1 (N4267, N4266);
nand NAND4 (N4268, N4259, N285, N58, N2575);
xor XOR2 (N4269, N4267, N2906);
or OR3 (N4270, N4256, N4114, N2314);
and AND2 (N4271, N4263, N2642);
nand NAND4 (N4272, N4270, N713, N999, N1178);
buf BUF1 (N4273, N4249);
nand NAND4 (N4274, N4268, N3343, N2205, N3241);
buf BUF1 (N4275, N4269);
nand NAND3 (N4276, N4272, N882, N145);
nand NAND3 (N4277, N4274, N3041, N2684);
buf BUF1 (N4278, N4271);
or OR2 (N4279, N4265, N410);
buf BUF1 (N4280, N4260);
not NOT1 (N4281, N4273);
buf BUF1 (N4282, N4279);
not NOT1 (N4283, N4255);
xor XOR2 (N4284, N4280, N3601);
buf BUF1 (N4285, N4283);
buf BUF1 (N4286, N4277);
nand NAND3 (N4287, N4275, N3033, N1614);
nor NOR4 (N4288, N4278, N3911, N1421, N1017);
xor XOR2 (N4289, N4262, N227);
or OR3 (N4290, N4287, N1090, N936);
or OR2 (N4291, N4281, N793);
buf BUF1 (N4292, N4285);
nand NAND3 (N4293, N4292, N3415, N4155);
not NOT1 (N4294, N4293);
not NOT1 (N4295, N4294);
nor NOR3 (N4296, N4289, N2629, N4276);
buf BUF1 (N4297, N1986);
or OR2 (N4298, N4286, N3540);
buf BUF1 (N4299, N4284);
or OR2 (N4300, N4298, N1471);
or OR4 (N4301, N4296, N4089, N500, N489);
or OR4 (N4302, N4290, N290, N3590, N804);
not NOT1 (N4303, N4295);
and AND3 (N4304, N4301, N1706, N667);
nor NOR2 (N4305, N4302, N2470);
xor XOR2 (N4306, N4305, N983);
xor XOR2 (N4307, N4303, N3555);
nor NOR2 (N4308, N4306, N3504);
nand NAND2 (N4309, N4304, N4037);
not NOT1 (N4310, N4245);
xor XOR2 (N4311, N4309, N4248);
or OR3 (N4312, N4300, N1443, N1206);
nand NAND4 (N4313, N4297, N2000, N87, N1437);
buf BUF1 (N4314, N4312);
nand NAND2 (N4315, N4308, N4288);
nand NAND2 (N4316, N1961, N2754);
not NOT1 (N4317, N4282);
not NOT1 (N4318, N4315);
and AND3 (N4319, N4310, N1549, N3743);
xor XOR2 (N4320, N4299, N4120);
nor NOR4 (N4321, N4318, N3402, N3687, N3935);
xor XOR2 (N4322, N4314, N147);
buf BUF1 (N4323, N4307);
or OR3 (N4324, N4323, N1236, N911);
buf BUF1 (N4325, N4319);
or OR4 (N4326, N4291, N607, N1537, N3099);
buf BUF1 (N4327, N4322);
buf BUF1 (N4328, N4313);
and AND4 (N4329, N4326, N2679, N1474, N2991);
buf BUF1 (N4330, N4329);
nand NAND2 (N4331, N4328, N2864);
xor XOR2 (N4332, N4321, N1344);
xor XOR2 (N4333, N4320, N3913);
not NOT1 (N4334, N4316);
buf BUF1 (N4335, N4317);
not NOT1 (N4336, N4335);
nor NOR2 (N4337, N4311, N148);
not NOT1 (N4338, N4324);
xor XOR2 (N4339, N4333, N870);
buf BUF1 (N4340, N4337);
not NOT1 (N4341, N4327);
and AND4 (N4342, N4325, N3257, N4164, N3980);
buf BUF1 (N4343, N4339);
nand NAND4 (N4344, N4340, N2907, N545, N216);
nand NAND3 (N4345, N4332, N3363, N2654);
and AND4 (N4346, N4330, N4232, N251, N900);
buf BUF1 (N4347, N4346);
not NOT1 (N4348, N4338);
xor XOR2 (N4349, N4336, N3861);
not NOT1 (N4350, N4334);
nand NAND2 (N4351, N4345, N1848);
not NOT1 (N4352, N4348);
nand NAND4 (N4353, N4347, N3251, N1617, N2973);
nand NAND2 (N4354, N4351, N962);
nor NOR2 (N4355, N4342, N4288);
xor XOR2 (N4356, N4353, N1985);
nand NAND2 (N4357, N4356, N3084);
nor NOR3 (N4358, N4344, N457, N1663);
xor XOR2 (N4359, N4349, N1749);
and AND4 (N4360, N4352, N2061, N189, N1519);
nand NAND4 (N4361, N4354, N4061, N4195, N808);
and AND4 (N4362, N4355, N1877, N3131, N1195);
or OR2 (N4363, N4361, N2935);
not NOT1 (N4364, N4357);
or OR3 (N4365, N4358, N847, N1551);
nand NAND3 (N4366, N4365, N1660, N3074);
or OR4 (N4367, N4366, N1097, N1870, N3078);
not NOT1 (N4368, N4367);
and AND4 (N4369, N4331, N2905, N2117, N3709);
not NOT1 (N4370, N4359);
xor XOR2 (N4371, N4341, N3498);
buf BUF1 (N4372, N4371);
nor NOR3 (N4373, N4362, N3607, N894);
xor XOR2 (N4374, N4370, N2790);
buf BUF1 (N4375, N4369);
or OR4 (N4376, N4372, N3903, N2956, N173);
nor NOR2 (N4377, N4343, N2712);
nor NOR4 (N4378, N4376, N2257, N1321, N142);
or OR2 (N4379, N4350, N3689);
and AND2 (N4380, N4374, N1306);
xor XOR2 (N4381, N4368, N2062);
not NOT1 (N4382, N4377);
nor NOR2 (N4383, N4363, N4180);
xor XOR2 (N4384, N4360, N1424);
not NOT1 (N4385, N4378);
nor NOR4 (N4386, N4373, N2287, N3800, N2228);
buf BUF1 (N4387, N4381);
and AND3 (N4388, N4379, N887, N1202);
nand NAND2 (N4389, N4383, N4152);
or OR2 (N4390, N4382, N1887);
or OR3 (N4391, N4364, N703, N209);
not NOT1 (N4392, N4375);
or OR4 (N4393, N4390, N376, N1092, N1907);
nor NOR3 (N4394, N4380, N2668, N1447);
nor NOR2 (N4395, N4391, N2395);
not NOT1 (N4396, N4393);
and AND2 (N4397, N4395, N4288);
or OR4 (N4398, N4396, N3640, N440, N1981);
not NOT1 (N4399, N4398);
or OR4 (N4400, N4387, N2463, N4203, N163);
xor XOR2 (N4401, N4384, N1333);
xor XOR2 (N4402, N4389, N1244);
not NOT1 (N4403, N4402);
xor XOR2 (N4404, N4399, N580);
or OR4 (N4405, N4403, N2125, N2849, N1707);
nand NAND2 (N4406, N4386, N2744);
nor NOR2 (N4407, N4400, N2714);
nand NAND4 (N4408, N4405, N729, N1250, N2886);
xor XOR2 (N4409, N4397, N4378);
and AND4 (N4410, N4406, N2016, N2793, N1282);
not NOT1 (N4411, N4408);
xor XOR2 (N4412, N4401, N2751);
buf BUF1 (N4413, N4409);
not NOT1 (N4414, N4388);
or OR3 (N4415, N4411, N37, N4366);
nor NOR4 (N4416, N4407, N2024, N3359, N456);
nor NOR2 (N4417, N4394, N4284);
buf BUF1 (N4418, N4414);
or OR2 (N4419, N4410, N3056);
xor XOR2 (N4420, N4385, N3359);
xor XOR2 (N4421, N4419, N755);
not NOT1 (N4422, N4413);
or OR3 (N4423, N4404, N2685, N3473);
nor NOR4 (N4424, N4415, N2635, N3589, N4325);
xor XOR2 (N4425, N4418, N4021);
nand NAND2 (N4426, N4420, N2586);
xor XOR2 (N4427, N4416, N2755);
or OR4 (N4428, N4425, N219, N4213, N2188);
xor XOR2 (N4429, N4428, N427);
nand NAND3 (N4430, N4421, N38, N2736);
and AND2 (N4431, N4426, N1220);
nor NOR4 (N4432, N4423, N1907, N1811, N1238);
buf BUF1 (N4433, N4424);
or OR4 (N4434, N4429, N3152, N3152, N1215);
and AND3 (N4435, N4392, N4028, N3118);
not NOT1 (N4436, N4412);
xor XOR2 (N4437, N4432, N2458);
not NOT1 (N4438, N4431);
buf BUF1 (N4439, N4436);
not NOT1 (N4440, N4417);
or OR2 (N4441, N4439, N1821);
or OR4 (N4442, N4441, N713, N4407, N4142);
not NOT1 (N4443, N4437);
nor NOR3 (N4444, N4440, N3728, N4057);
or OR3 (N4445, N4438, N262, N470);
and AND3 (N4446, N4433, N4382, N3307);
not NOT1 (N4447, N4435);
or OR4 (N4448, N4434, N2656, N279, N453);
nor NOR2 (N4449, N4430, N3608);
not NOT1 (N4450, N4444);
not NOT1 (N4451, N4450);
xor XOR2 (N4452, N4448, N871);
nor NOR3 (N4453, N4452, N3387, N220);
nand NAND2 (N4454, N4443, N3553);
xor XOR2 (N4455, N4447, N63);
nor NOR3 (N4456, N4422, N4309, N3729);
or OR2 (N4457, N4451, N1574);
xor XOR2 (N4458, N4454, N2865);
or OR3 (N4459, N4427, N2795, N2079);
xor XOR2 (N4460, N4458, N1440);
xor XOR2 (N4461, N4449, N2618);
or OR4 (N4462, N4457, N1579, N208, N819);
or OR2 (N4463, N4456, N1794);
and AND3 (N4464, N4460, N1455, N3119);
and AND3 (N4465, N4455, N2705, N2967);
xor XOR2 (N4466, N4465, N3764);
not NOT1 (N4467, N4466);
xor XOR2 (N4468, N4461, N3986);
nor NOR2 (N4469, N4446, N299);
buf BUF1 (N4470, N4453);
and AND3 (N4471, N4459, N968, N459);
and AND2 (N4472, N4468, N1957);
and AND3 (N4473, N4472, N2155, N697);
or OR2 (N4474, N4467, N176);
buf BUF1 (N4475, N4442);
or OR3 (N4476, N4473, N1105, N574);
not NOT1 (N4477, N4463);
nor NOR2 (N4478, N4471, N2777);
nand NAND2 (N4479, N4462, N3678);
nand NAND4 (N4480, N4464, N2530, N882, N134);
xor XOR2 (N4481, N4470, N3046);
nor NOR2 (N4482, N4480, N1026);
nor NOR2 (N4483, N4474, N1062);
buf BUF1 (N4484, N4475);
nor NOR2 (N4485, N4482, N2757);
or OR3 (N4486, N4445, N1048, N2621);
and AND2 (N4487, N4477, N1682);
nor NOR2 (N4488, N4469, N2744);
xor XOR2 (N4489, N4487, N3706);
or OR4 (N4490, N4476, N2664, N748, N1287);
xor XOR2 (N4491, N4489, N1601);
nor NOR4 (N4492, N4491, N478, N1369, N1968);
not NOT1 (N4493, N4488);
nor NOR3 (N4494, N4483, N1405, N2618);
or OR3 (N4495, N4493, N491, N173);
buf BUF1 (N4496, N4492);
buf BUF1 (N4497, N4485);
buf BUF1 (N4498, N4479);
xor XOR2 (N4499, N4494, N2984);
not NOT1 (N4500, N4495);
buf BUF1 (N4501, N4484);
nand NAND4 (N4502, N4500, N3907, N1523, N3442);
buf BUF1 (N4503, N4502);
not NOT1 (N4504, N4496);
buf BUF1 (N4505, N4497);
buf BUF1 (N4506, N4486);
and AND3 (N4507, N4504, N484, N515);
buf BUF1 (N4508, N4498);
xor XOR2 (N4509, N4499, N2409);
buf BUF1 (N4510, N4503);
nand NAND4 (N4511, N4510, N2054, N2056, N4210);
nand NAND3 (N4512, N4505, N2773, N271);
nand NAND2 (N4513, N4506, N2400);
nand NAND4 (N4514, N4507, N1207, N1296, N1840);
nor NOR3 (N4515, N4513, N315, N1205);
not NOT1 (N4516, N4501);
buf BUF1 (N4517, N4509);
and AND2 (N4518, N4508, N2692);
and AND3 (N4519, N4481, N2848, N857);
and AND4 (N4520, N4516, N529, N4094, N2676);
or OR3 (N4521, N4520, N4024, N939);
xor XOR2 (N4522, N4519, N2259);
nand NAND4 (N4523, N4478, N2594, N3557, N1249);
buf BUF1 (N4524, N4523);
not NOT1 (N4525, N4515);
xor XOR2 (N4526, N4521, N723);
xor XOR2 (N4527, N4490, N4396);
xor XOR2 (N4528, N4524, N4309);
and AND3 (N4529, N4528, N125, N2444);
xor XOR2 (N4530, N4512, N3426);
nor NOR4 (N4531, N4511, N3593, N1994, N2694);
or OR3 (N4532, N4522, N1082, N1996);
buf BUF1 (N4533, N4532);
nand NAND2 (N4534, N4518, N1989);
nand NAND4 (N4535, N4530, N1012, N2179, N3881);
buf BUF1 (N4536, N4534);
or OR4 (N4537, N4533, N2823, N2673, N2491);
not NOT1 (N4538, N4536);
nor NOR3 (N4539, N4537, N3293, N1837);
nor NOR2 (N4540, N4538, N2092);
buf BUF1 (N4541, N4535);
buf BUF1 (N4542, N4539);
nor NOR4 (N4543, N4541, N1271, N2123, N752);
buf BUF1 (N4544, N4540);
and AND4 (N4545, N4542, N1294, N4357, N524);
and AND4 (N4546, N4514, N4365, N803, N272);
xor XOR2 (N4547, N4529, N292);
not NOT1 (N4548, N4531);
buf BUF1 (N4549, N4544);
nand NAND2 (N4550, N4545, N4504);
not NOT1 (N4551, N4548);
nand NAND2 (N4552, N4549, N3041);
not NOT1 (N4553, N4525);
not NOT1 (N4554, N4551);
and AND2 (N4555, N4547, N3023);
nor NOR4 (N4556, N4555, N1852, N2734, N1177);
nand NAND2 (N4557, N4550, N4378);
or OR2 (N4558, N4527, N1207);
not NOT1 (N4559, N4526);
not NOT1 (N4560, N4553);
and AND4 (N4561, N4557, N1296, N4420, N3237);
nor NOR3 (N4562, N4559, N4241, N1710);
buf BUF1 (N4563, N4560);
buf BUF1 (N4564, N4543);
buf BUF1 (N4565, N4517);
xor XOR2 (N4566, N4558, N3908);
buf BUF1 (N4567, N4565);
not NOT1 (N4568, N4566);
not NOT1 (N4569, N4552);
buf BUF1 (N4570, N4563);
or OR2 (N4571, N4556, N803);
nand NAND2 (N4572, N4568, N4158);
not NOT1 (N4573, N4561);
nand NAND4 (N4574, N4564, N3362, N3196, N3878);
or OR3 (N4575, N4562, N1674, N2305);
not NOT1 (N4576, N4572);
or OR2 (N4577, N4546, N2905);
xor XOR2 (N4578, N4569, N958);
and AND4 (N4579, N4573, N383, N4332, N2098);
xor XOR2 (N4580, N4571, N673);
xor XOR2 (N4581, N4579, N2679);
or OR3 (N4582, N4578, N1683, N1801);
xor XOR2 (N4583, N4580, N1774);
nor NOR4 (N4584, N4554, N3928, N4486, N3892);
nor NOR3 (N4585, N4576, N1014, N1974);
nor NOR4 (N4586, N4574, N134, N2411, N183);
nor NOR2 (N4587, N4583, N2536);
or OR2 (N4588, N4570, N2318);
buf BUF1 (N4589, N4577);
nor NOR2 (N4590, N4567, N2629);
and AND2 (N4591, N4581, N990);
xor XOR2 (N4592, N4587, N2070);
nand NAND2 (N4593, N4586, N4516);
or OR4 (N4594, N4585, N2828, N2242, N2626);
not NOT1 (N4595, N4591);
xor XOR2 (N4596, N4592, N1946);
nor NOR4 (N4597, N4595, N97, N1991, N4073);
xor XOR2 (N4598, N4593, N4288);
xor XOR2 (N4599, N4588, N1753);
or OR4 (N4600, N4594, N690, N2361, N1926);
buf BUF1 (N4601, N4598);
nor NOR4 (N4602, N4584, N4478, N3344, N1905);
or OR2 (N4603, N4602, N335);
xor XOR2 (N4604, N4599, N1548);
buf BUF1 (N4605, N4590);
xor XOR2 (N4606, N4601, N1299);
not NOT1 (N4607, N4600);
or OR3 (N4608, N4605, N707, N3804);
nor NOR4 (N4609, N4596, N1306, N1300, N1776);
or OR2 (N4610, N4604, N70);
nor NOR3 (N4611, N4607, N777, N222);
or OR2 (N4612, N4603, N1607);
not NOT1 (N4613, N4610);
buf BUF1 (N4614, N4609);
buf BUF1 (N4615, N4582);
xor XOR2 (N4616, N4608, N3437);
or OR3 (N4617, N4613, N2035, N3714);
nand NAND4 (N4618, N4575, N2259, N1786, N751);
nor NOR2 (N4619, N4589, N432);
or OR3 (N4620, N4619, N2718, N1427);
or OR4 (N4621, N4612, N2061, N2829, N4515);
and AND4 (N4622, N4615, N4020, N291, N2033);
or OR3 (N4623, N4606, N516, N1012);
not NOT1 (N4624, N4620);
and AND2 (N4625, N4614, N1281);
not NOT1 (N4626, N4623);
nand NAND3 (N4627, N4597, N6, N129);
buf BUF1 (N4628, N4624);
and AND4 (N4629, N4628, N2399, N36, N3199);
xor XOR2 (N4630, N4617, N1975);
nand NAND3 (N4631, N4622, N3413, N623);
or OR2 (N4632, N4618, N268);
or OR4 (N4633, N4611, N2160, N1956, N3793);
buf BUF1 (N4634, N4632);
buf BUF1 (N4635, N4630);
and AND2 (N4636, N4635, N2689);
and AND2 (N4637, N4629, N2861);
xor XOR2 (N4638, N4633, N4464);
and AND4 (N4639, N4636, N430, N3198, N1387);
nor NOR3 (N4640, N4631, N3269, N885);
nor NOR4 (N4641, N4621, N2299, N2183, N2715);
buf BUF1 (N4642, N4641);
or OR2 (N4643, N4642, N1483);
nor NOR4 (N4644, N4625, N1952, N2725, N335);
and AND3 (N4645, N4616, N2822, N2319);
nor NOR2 (N4646, N4626, N3452);
nor NOR4 (N4647, N4637, N307, N4306, N215);
xor XOR2 (N4648, N4644, N4110);
and AND2 (N4649, N4643, N616);
not NOT1 (N4650, N4638);
nor NOR3 (N4651, N4634, N812, N2468);
nand NAND3 (N4652, N4650, N670, N3586);
or OR2 (N4653, N4627, N833);
buf BUF1 (N4654, N4651);
nor NOR3 (N4655, N4646, N3895, N3509);
and AND3 (N4656, N4645, N25, N435);
not NOT1 (N4657, N4639);
not NOT1 (N4658, N4647);
and AND4 (N4659, N4654, N3899, N2931, N611);
xor XOR2 (N4660, N4658, N1187);
xor XOR2 (N4661, N4656, N2863);
nand NAND3 (N4662, N4657, N1789, N4292);
xor XOR2 (N4663, N4640, N1152);
buf BUF1 (N4664, N4660);
or OR2 (N4665, N4655, N3687);
not NOT1 (N4666, N4663);
nor NOR3 (N4667, N4664, N3739, N4498);
not NOT1 (N4668, N4659);
or OR4 (N4669, N4652, N2966, N2122, N3470);
buf BUF1 (N4670, N4662);
not NOT1 (N4671, N4649);
nor NOR4 (N4672, N4661, N3706, N3858, N2238);
nor NOR3 (N4673, N4671, N2103, N4502);
nor NOR4 (N4674, N4653, N784, N2211, N4354);
and AND3 (N4675, N4666, N1366, N1487);
or OR4 (N4676, N4674, N2128, N3789, N718);
nand NAND4 (N4677, N4665, N679, N1647, N2549);
buf BUF1 (N4678, N4670);
buf BUF1 (N4679, N4667);
nand NAND2 (N4680, N4669, N1785);
or OR3 (N4681, N4675, N796, N3731);
xor XOR2 (N4682, N4668, N4228);
or OR2 (N4683, N4648, N2824);
nand NAND4 (N4684, N4682, N4019, N2105, N3029);
and AND4 (N4685, N4683, N2743, N1164, N1443);
xor XOR2 (N4686, N4676, N407);
nor NOR3 (N4687, N4677, N4669, N844);
and AND3 (N4688, N4680, N3822, N1338);
and AND4 (N4689, N4684, N4340, N2625, N2403);
buf BUF1 (N4690, N4686);
xor XOR2 (N4691, N4687, N4015);
xor XOR2 (N4692, N4673, N3233);
xor XOR2 (N4693, N4681, N818);
nor NOR3 (N4694, N4689, N1996, N2685);
buf BUF1 (N4695, N4679);
not NOT1 (N4696, N4688);
not NOT1 (N4697, N4696);
nand NAND2 (N4698, N4692, N3524);
xor XOR2 (N4699, N4672, N4599);
buf BUF1 (N4700, N4690);
xor XOR2 (N4701, N4699, N3099);
buf BUF1 (N4702, N4695);
not NOT1 (N4703, N4700);
or OR2 (N4704, N4698, N3768);
nand NAND4 (N4705, N4678, N4378, N785, N3323);
nand NAND4 (N4706, N4697, N982, N1327, N3789);
buf BUF1 (N4707, N4703);
xor XOR2 (N4708, N4702, N2550);
nor NOR4 (N4709, N4694, N3409, N4274, N302);
not NOT1 (N4710, N4706);
not NOT1 (N4711, N4709);
buf BUF1 (N4712, N4705);
buf BUF1 (N4713, N4704);
nor NOR4 (N4714, N4713, N881, N1067, N1270);
buf BUF1 (N4715, N4693);
xor XOR2 (N4716, N4708, N3509);
nor NOR2 (N4717, N4701, N4611);
xor XOR2 (N4718, N4710, N297);
or OR4 (N4719, N4717, N695, N2138, N963);
buf BUF1 (N4720, N4718);
or OR2 (N4721, N4707, N4534);
or OR2 (N4722, N4719, N1130);
or OR2 (N4723, N4715, N3958);
xor XOR2 (N4724, N4712, N552);
nand NAND4 (N4725, N4714, N2019, N134, N1249);
and AND2 (N4726, N4720, N4236);
and AND2 (N4727, N4723, N3742);
nand NAND4 (N4728, N4725, N2978, N458, N1593);
xor XOR2 (N4729, N4727, N3764);
xor XOR2 (N4730, N4685, N2347);
buf BUF1 (N4731, N4721);
nor NOR4 (N4732, N4728, N3018, N4474, N4200);
xor XOR2 (N4733, N4729, N1734);
xor XOR2 (N4734, N4733, N4205);
nand NAND2 (N4735, N4726, N2914);
nand NAND3 (N4736, N4691, N2418, N682);
xor XOR2 (N4737, N4735, N2886);
and AND4 (N4738, N4730, N3412, N2935, N2304);
or OR3 (N4739, N4731, N1212, N2102);
and AND3 (N4740, N4737, N397, N1671);
and AND2 (N4741, N4734, N1912);
buf BUF1 (N4742, N4732);
nand NAND4 (N4743, N4722, N4368, N3143, N1367);
not NOT1 (N4744, N4739);
buf BUF1 (N4745, N4744);
buf BUF1 (N4746, N4743);
or OR2 (N4747, N4711, N2024);
not NOT1 (N4748, N4716);
nor NOR4 (N4749, N4742, N1484, N2012, N2350);
xor XOR2 (N4750, N4736, N752);
xor XOR2 (N4751, N4750, N4383);
and AND4 (N4752, N4740, N415, N1379, N1753);
nand NAND2 (N4753, N4752, N4144);
and AND2 (N4754, N4753, N1561);
not NOT1 (N4755, N4754);
nor NOR2 (N4756, N4746, N2212);
not NOT1 (N4757, N4755);
buf BUF1 (N4758, N4757);
or OR2 (N4759, N4738, N2470);
not NOT1 (N4760, N4751);
nor NOR2 (N4761, N4747, N2138);
buf BUF1 (N4762, N4724);
xor XOR2 (N4763, N4745, N3656);
not NOT1 (N4764, N4748);
and AND4 (N4765, N4759, N273, N209, N1310);
nand NAND4 (N4766, N4758, N2691, N1041, N4430);
not NOT1 (N4767, N4756);
xor XOR2 (N4768, N4764, N1247);
xor XOR2 (N4769, N4761, N3342);
nand NAND4 (N4770, N4767, N2326, N2527, N1717);
nand NAND3 (N4771, N4768, N570, N3190);
nand NAND3 (N4772, N4760, N90, N825);
not NOT1 (N4773, N4770);
nand NAND4 (N4774, N4771, N2431, N4464, N2522);
nor NOR3 (N4775, N4769, N3653, N556);
not NOT1 (N4776, N4772);
nand NAND3 (N4777, N4765, N2295, N2857);
buf BUF1 (N4778, N4777);
not NOT1 (N4779, N4741);
xor XOR2 (N4780, N4778, N650);
not NOT1 (N4781, N4779);
nand NAND2 (N4782, N4749, N4255);
buf BUF1 (N4783, N4773);
buf BUF1 (N4784, N4774);
nor NOR3 (N4785, N4763, N1619, N1628);
not NOT1 (N4786, N4784);
xor XOR2 (N4787, N4783, N1681);
nand NAND4 (N4788, N4785, N3317, N3318, N3797);
xor XOR2 (N4789, N4762, N4197);
nor NOR4 (N4790, N4789, N3840, N2921, N3366);
xor XOR2 (N4791, N4776, N2518);
not NOT1 (N4792, N4780);
not NOT1 (N4793, N4787);
nand NAND4 (N4794, N4786, N206, N3846, N2729);
nor NOR2 (N4795, N4775, N1776);
or OR4 (N4796, N4795, N633, N3595, N4479);
nand NAND2 (N4797, N4796, N4459);
xor XOR2 (N4798, N4791, N3910);
xor XOR2 (N4799, N4798, N2937);
not NOT1 (N4800, N4794);
xor XOR2 (N4801, N4793, N2726);
not NOT1 (N4802, N4799);
not NOT1 (N4803, N4797);
nand NAND3 (N4804, N4782, N1344, N108);
not NOT1 (N4805, N4801);
xor XOR2 (N4806, N4800, N820);
and AND4 (N4807, N4766, N3724, N3386, N702);
xor XOR2 (N4808, N4806, N692);
xor XOR2 (N4809, N4802, N1493);
and AND2 (N4810, N4805, N1277);
nand NAND2 (N4811, N4792, N1093);
nand NAND3 (N4812, N4811, N2002, N4742);
buf BUF1 (N4813, N4807);
xor XOR2 (N4814, N4790, N932);
nor NOR2 (N4815, N4804, N2844);
nor NOR3 (N4816, N4812, N1626, N4774);
xor XOR2 (N4817, N4781, N1613);
nor NOR2 (N4818, N4809, N4432);
not NOT1 (N4819, N4808);
buf BUF1 (N4820, N4816);
and AND4 (N4821, N4813, N4411, N986, N327);
and AND4 (N4822, N4820, N1658, N179, N1008);
not NOT1 (N4823, N4819);
xor XOR2 (N4824, N4817, N2712);
and AND4 (N4825, N4823, N4436, N2533, N3618);
and AND4 (N4826, N4803, N4242, N4206, N1246);
nor NOR2 (N4827, N4814, N3420);
buf BUF1 (N4828, N4788);
and AND4 (N4829, N4815, N1223, N3418, N2603);
and AND2 (N4830, N4828, N1654);
and AND2 (N4831, N4825, N1846);
not NOT1 (N4832, N4826);
buf BUF1 (N4833, N4824);
or OR3 (N4834, N4810, N2302, N1919);
or OR4 (N4835, N4829, N3120, N2667, N4115);
not NOT1 (N4836, N4821);
and AND2 (N4837, N4818, N2065);
nor NOR3 (N4838, N4830, N2240, N4415);
nor NOR2 (N4839, N4836, N2627);
nand NAND2 (N4840, N4837, N3471);
not NOT1 (N4841, N4822);
buf BUF1 (N4842, N4832);
xor XOR2 (N4843, N4841, N4156);
and AND4 (N4844, N4840, N43, N3789, N978);
xor XOR2 (N4845, N4843, N1231);
nand NAND2 (N4846, N4845, N1379);
xor XOR2 (N4847, N4838, N2037);
and AND2 (N4848, N4847, N1457);
not NOT1 (N4849, N4848);
buf BUF1 (N4850, N4844);
xor XOR2 (N4851, N4850, N1018);
not NOT1 (N4852, N4846);
and AND3 (N4853, N4827, N2753, N4311);
not NOT1 (N4854, N4851);
xor XOR2 (N4855, N4839, N3564);
nor NOR2 (N4856, N4849, N1399);
nand NAND4 (N4857, N4853, N490, N1248, N3594);
or OR4 (N4858, N4831, N3198, N3520, N426);
xor XOR2 (N4859, N4854, N2165);
buf BUF1 (N4860, N4835);
xor XOR2 (N4861, N4860, N2626);
nand NAND4 (N4862, N4834, N4327, N1599, N1222);
nand NAND4 (N4863, N4833, N4643, N4313, N1123);
and AND4 (N4864, N4842, N3770, N2226, N4141);
not NOT1 (N4865, N4852);
nand NAND2 (N4866, N4858, N2949);
nor NOR4 (N4867, N4857, N2554, N1530, N4621);
buf BUF1 (N4868, N4863);
and AND3 (N4869, N4859, N2581, N2760);
nor NOR3 (N4870, N4861, N1296, N1786);
xor XOR2 (N4871, N4856, N1502);
or OR2 (N4872, N4868, N4810);
and AND3 (N4873, N4862, N1769, N2242);
nand NAND3 (N4874, N4872, N3373, N2933);
xor XOR2 (N4875, N4870, N4013);
nand NAND2 (N4876, N4874, N1493);
not NOT1 (N4877, N4866);
nand NAND3 (N4878, N4865, N1532, N1624);
or OR2 (N4879, N4875, N4441);
or OR3 (N4880, N4864, N4035, N1269);
xor XOR2 (N4881, N4880, N3446);
not NOT1 (N4882, N4867);
xor XOR2 (N4883, N4881, N14);
nor NOR4 (N4884, N4871, N4159, N18, N2113);
not NOT1 (N4885, N4878);
nor NOR4 (N4886, N4877, N305, N3070, N941);
not NOT1 (N4887, N4879);
and AND2 (N4888, N4887, N154);
not NOT1 (N4889, N4873);
not NOT1 (N4890, N4885);
nor NOR3 (N4891, N4888, N25, N843);
not NOT1 (N4892, N4886);
xor XOR2 (N4893, N4855, N2052);
or OR3 (N4894, N4883, N4716, N2506);
not NOT1 (N4895, N4890);
buf BUF1 (N4896, N4869);
or OR2 (N4897, N4876, N877);
nand NAND2 (N4898, N4892, N2744);
not NOT1 (N4899, N4893);
buf BUF1 (N4900, N4895);
buf BUF1 (N4901, N4897);
or OR3 (N4902, N4894, N3054, N1451);
not NOT1 (N4903, N4899);
nor NOR3 (N4904, N4896, N4637, N515);
buf BUF1 (N4905, N4904);
nor NOR3 (N4906, N4902, N4558, N798);
not NOT1 (N4907, N4884);
nand NAND4 (N4908, N4900, N2085, N3729, N4332);
and AND4 (N4909, N4903, N4029, N3604, N3046);
nand NAND3 (N4910, N4909, N1529, N225);
nor NOR2 (N4911, N4907, N1619);
nor NOR3 (N4912, N4911, N3529, N4073);
or OR2 (N4913, N4910, N1689);
or OR2 (N4914, N4913, N4429);
and AND2 (N4915, N4889, N2666);
xor XOR2 (N4916, N4882, N1089);
nor NOR4 (N4917, N4898, N536, N3880, N2763);
buf BUF1 (N4918, N4905);
nor NOR4 (N4919, N4914, N4814, N4625, N583);
buf BUF1 (N4920, N4915);
nor NOR2 (N4921, N4918, N786);
nor NOR4 (N4922, N4920, N2600, N2862, N3822);
nand NAND2 (N4923, N4921, N3869);
and AND3 (N4924, N4919, N2690, N2504);
nand NAND3 (N4925, N4906, N2762, N4467);
nand NAND2 (N4926, N4912, N4344);
xor XOR2 (N4927, N4925, N844);
or OR4 (N4928, N4923, N2315, N3155, N4637);
xor XOR2 (N4929, N4891, N3308);
nor NOR3 (N4930, N4929, N2096, N1736);
or OR2 (N4931, N4927, N2263);
nor NOR2 (N4932, N4928, N2548);
buf BUF1 (N4933, N4932);
and AND2 (N4934, N4926, N3258);
not NOT1 (N4935, N4924);
not NOT1 (N4936, N4922);
and AND2 (N4937, N4901, N124);
and AND4 (N4938, N4934, N4206, N3056, N1544);
and AND4 (N4939, N4937, N3021, N3543, N2823);
nor NOR4 (N4940, N4938, N1711, N1509, N2099);
buf BUF1 (N4941, N4917);
or OR3 (N4942, N4930, N3996, N2561);
xor XOR2 (N4943, N4916, N479);
and AND4 (N4944, N4935, N2476, N769, N2966);
nor NOR4 (N4945, N4943, N4311, N1837, N2159);
nand NAND3 (N4946, N4936, N4748, N1581);
nand NAND4 (N4947, N4945, N4659, N4048, N2525);
and AND4 (N4948, N4939, N3159, N487, N4902);
not NOT1 (N4949, N4933);
not NOT1 (N4950, N4942);
not NOT1 (N4951, N4940);
and AND2 (N4952, N4941, N3976);
buf BUF1 (N4953, N4947);
nand NAND2 (N4954, N4944, N3070);
nand NAND3 (N4955, N4931, N3679, N3053);
nand NAND4 (N4956, N4949, N2183, N68, N384);
xor XOR2 (N4957, N4952, N1631);
nor NOR3 (N4958, N4951, N4193, N704);
buf BUF1 (N4959, N4948);
nand NAND4 (N4960, N4954, N1688, N92, N1480);
nor NOR2 (N4961, N4953, N4501);
or OR3 (N4962, N4960, N1056, N4657);
nand NAND3 (N4963, N4961, N1460, N4019);
xor XOR2 (N4964, N4956, N4882);
xor XOR2 (N4965, N4955, N4073);
xor XOR2 (N4966, N4964, N152);
not NOT1 (N4967, N4957);
not NOT1 (N4968, N4958);
nand NAND3 (N4969, N4968, N3333, N4567);
and AND2 (N4970, N4967, N4863);
nand NAND4 (N4971, N4963, N1553, N4945, N2231);
nor NOR3 (N4972, N4965, N3000, N2101);
buf BUF1 (N4973, N4908);
buf BUF1 (N4974, N4950);
buf BUF1 (N4975, N4959);
not NOT1 (N4976, N4970);
not NOT1 (N4977, N4973);
not NOT1 (N4978, N4962);
not NOT1 (N4979, N4976);
not NOT1 (N4980, N4966);
xor XOR2 (N4981, N4971, N4837);
buf BUF1 (N4982, N4974);
buf BUF1 (N4983, N4980);
or OR2 (N4984, N4969, N4216);
xor XOR2 (N4985, N4979, N1028);
xor XOR2 (N4986, N4972, N2770);
buf BUF1 (N4987, N4975);
and AND2 (N4988, N4977, N761);
nor NOR2 (N4989, N4946, N4442);
nand NAND3 (N4990, N4983, N2480, N1404);
and AND2 (N4991, N4988, N3426);
nor NOR3 (N4992, N4982, N4768, N1617);
not NOT1 (N4993, N4978);
nand NAND3 (N4994, N4993, N2941, N1166);
buf BUF1 (N4995, N4992);
nand NAND2 (N4996, N4990, N2398);
xor XOR2 (N4997, N4995, N3064);
buf BUF1 (N4998, N4984);
not NOT1 (N4999, N4989);
xor XOR2 (N5000, N4981, N997);
not NOT1 (N5001, N4997);
nand NAND4 (N5002, N5001, N167, N3524, N3665);
nor NOR3 (N5003, N5000, N733, N4176);
nor NOR3 (N5004, N4999, N3056, N3078);
not NOT1 (N5005, N5004);
xor XOR2 (N5006, N4994, N3812);
or OR2 (N5007, N4987, N1014);
or OR3 (N5008, N4996, N336, N1940);
xor XOR2 (N5009, N4998, N3245);
not NOT1 (N5010, N4986);
nand NAND3 (N5011, N4985, N703, N4637);
nor NOR3 (N5012, N4991, N1072, N2585);
nand NAND2 (N5013, N5010, N3548);
or OR4 (N5014, N5006, N4717, N2435, N4042);
and AND3 (N5015, N5008, N2860, N4913);
xor XOR2 (N5016, N5005, N4752);
buf BUF1 (N5017, N5002);
not NOT1 (N5018, N5014);
nand NAND2 (N5019, N5003, N3588);
buf BUF1 (N5020, N5009);
or OR2 (N5021, N5007, N4147);
nand NAND2 (N5022, N5012, N2247);
buf BUF1 (N5023, N5021);
xor XOR2 (N5024, N5016, N73);
buf BUF1 (N5025, N5024);
nand NAND3 (N5026, N5025, N116, N777);
and AND2 (N5027, N5015, N649);
and AND4 (N5028, N5023, N3021, N3171, N4624);
nor NOR2 (N5029, N5028, N2353);
nor NOR2 (N5030, N5011, N4935);
or OR3 (N5031, N5020, N30, N3482);
and AND2 (N5032, N5019, N682);
buf BUF1 (N5033, N5018);
buf BUF1 (N5034, N5026);
not NOT1 (N5035, N5033);
or OR2 (N5036, N5035, N107);
and AND3 (N5037, N5017, N1371, N3719);
xor XOR2 (N5038, N5027, N4315);
nand NAND3 (N5039, N5022, N292, N2106);
xor XOR2 (N5040, N5034, N4768);
or OR2 (N5041, N5030, N983);
and AND3 (N5042, N5032, N3595, N2527);
nor NOR3 (N5043, N5029, N972, N1037);
nand NAND3 (N5044, N5031, N1722, N2235);
buf BUF1 (N5045, N5036);
nor NOR3 (N5046, N5041, N4155, N616);
or OR2 (N5047, N5044, N3923);
nand NAND3 (N5048, N5037, N4747, N1119);
or OR2 (N5049, N5043, N4537);
nor NOR2 (N5050, N5046, N4433);
xor XOR2 (N5051, N5045, N3313);
nor NOR4 (N5052, N5039, N3078, N1794, N2776);
buf BUF1 (N5053, N5042);
nand NAND2 (N5054, N5038, N1643);
nand NAND4 (N5055, N5052, N465, N4562, N4189);
xor XOR2 (N5056, N5048, N3468);
not NOT1 (N5057, N5013);
or OR3 (N5058, N5047, N891, N845);
not NOT1 (N5059, N5055);
nor NOR2 (N5060, N5040, N3783);
nor NOR3 (N5061, N5049, N2658, N1296);
buf BUF1 (N5062, N5056);
buf BUF1 (N5063, N5050);
xor XOR2 (N5064, N5063, N876);
not NOT1 (N5065, N5057);
nand NAND2 (N5066, N5062, N4367);
xor XOR2 (N5067, N5060, N52);
nor NOR3 (N5068, N5067, N1047, N3157);
nand NAND2 (N5069, N5058, N4243);
nand NAND2 (N5070, N5066, N3782);
buf BUF1 (N5071, N5069);
xor XOR2 (N5072, N5051, N152);
or OR3 (N5073, N5072, N4977, N1164);
xor XOR2 (N5074, N5064, N2640);
xor XOR2 (N5075, N5073, N3677);
nand NAND4 (N5076, N5071, N1419, N4675, N490);
or OR3 (N5077, N5054, N1977, N448);
xor XOR2 (N5078, N5075, N5);
and AND2 (N5079, N5068, N3205);
or OR2 (N5080, N5070, N4050);
xor XOR2 (N5081, N5061, N3007);
not NOT1 (N5082, N5076);
not NOT1 (N5083, N5074);
buf BUF1 (N5084, N5083);
and AND3 (N5085, N5079, N4471, N1258);
nand NAND3 (N5086, N5081, N3224, N1573);
nand NAND4 (N5087, N5077, N815, N307, N2613);
buf BUF1 (N5088, N5085);
buf BUF1 (N5089, N5086);
nor NOR2 (N5090, N5089, N4698);
buf BUF1 (N5091, N5065);
nor NOR3 (N5092, N5082, N1840, N4072);
xor XOR2 (N5093, N5091, N2214);
or OR2 (N5094, N5088, N1798);
nor NOR3 (N5095, N5092, N1100, N4042);
nor NOR2 (N5096, N5090, N264);
or OR4 (N5097, N5053, N4714, N4640, N3750);
or OR2 (N5098, N5084, N2548);
nor NOR3 (N5099, N5093, N4974, N3112);
and AND3 (N5100, N5097, N3833, N3814);
xor XOR2 (N5101, N5098, N4813);
xor XOR2 (N5102, N5095, N3752);
buf BUF1 (N5103, N5059);
buf BUF1 (N5104, N5080);
xor XOR2 (N5105, N5099, N2395);
or OR2 (N5106, N5078, N1154);
and AND2 (N5107, N5106, N1797);
xor XOR2 (N5108, N5096, N5098);
not NOT1 (N5109, N5087);
not NOT1 (N5110, N5100);
and AND3 (N5111, N5094, N38, N376);
and AND2 (N5112, N5102, N4179);
xor XOR2 (N5113, N5101, N1440);
nor NOR4 (N5114, N5112, N2840, N3541, N485);
nand NAND2 (N5115, N5114, N2201);
and AND4 (N5116, N5109, N3025, N34, N4044);
not NOT1 (N5117, N5113);
not NOT1 (N5118, N5105);
or OR3 (N5119, N5103, N4395, N87);
xor XOR2 (N5120, N5107, N2474);
nor NOR4 (N5121, N5120, N4774, N621, N4623);
or OR2 (N5122, N5116, N4085);
nor NOR2 (N5123, N5121, N3812);
or OR4 (N5124, N5104, N5067, N194, N2558);
buf BUF1 (N5125, N5124);
buf BUF1 (N5126, N5123);
or OR2 (N5127, N5115, N3291);
nand NAND3 (N5128, N5125, N3265, N1043);
buf BUF1 (N5129, N5119);
and AND4 (N5130, N5122, N630, N4357, N4571);
nand NAND2 (N5131, N5130, N4984);
xor XOR2 (N5132, N5128, N2839);
buf BUF1 (N5133, N5108);
not NOT1 (N5134, N5118);
and AND4 (N5135, N5110, N1780, N2334, N2961);
xor XOR2 (N5136, N5111, N2401);
xor XOR2 (N5137, N5126, N4775);
xor XOR2 (N5138, N5117, N3605);
xor XOR2 (N5139, N5132, N646);
buf BUF1 (N5140, N5135);
xor XOR2 (N5141, N5129, N1293);
and AND3 (N5142, N5133, N523, N1225);
nor NOR2 (N5143, N5140, N3104);
and AND4 (N5144, N5141, N2215, N4320, N1624);
buf BUF1 (N5145, N5127);
buf BUF1 (N5146, N5134);
and AND2 (N5147, N5143, N642);
and AND4 (N5148, N5139, N3667, N3076, N1629);
nor NOR4 (N5149, N5144, N174, N3221, N1651);
buf BUF1 (N5150, N5136);
nor NOR4 (N5151, N5142, N4137, N2103, N677);
nand NAND3 (N5152, N5148, N4800, N1227);
nor NOR4 (N5153, N5152, N2451, N3750, N1465);
nor NOR4 (N5154, N5151, N3450, N219, N3350);
and AND3 (N5155, N5137, N4025, N848);
or OR3 (N5156, N5138, N5141, N2590);
xor XOR2 (N5157, N5153, N3706);
not NOT1 (N5158, N5146);
xor XOR2 (N5159, N5157, N3148);
or OR2 (N5160, N5150, N3294);
or OR4 (N5161, N5149, N4961, N760, N1957);
nand NAND4 (N5162, N5156, N1331, N1690, N2688);
nor NOR4 (N5163, N5154, N4103, N242, N616);
and AND2 (N5164, N5159, N648);
nor NOR3 (N5165, N5162, N2311, N669);
nand NAND2 (N5166, N5147, N3024);
xor XOR2 (N5167, N5155, N4080);
not NOT1 (N5168, N5161);
buf BUF1 (N5169, N5168);
not NOT1 (N5170, N5160);
not NOT1 (N5171, N5164);
xor XOR2 (N5172, N5163, N3642);
and AND3 (N5173, N5172, N2756, N3291);
xor XOR2 (N5174, N5173, N3775);
nand NAND2 (N5175, N5171, N2141);
buf BUF1 (N5176, N5167);
or OR3 (N5177, N5174, N3279, N1124);
or OR2 (N5178, N5170, N869);
nor NOR4 (N5179, N5178, N2135, N1020, N1417);
xor XOR2 (N5180, N5145, N1149);
not NOT1 (N5181, N5180);
or OR3 (N5182, N5176, N4742, N1211);
buf BUF1 (N5183, N5166);
xor XOR2 (N5184, N5177, N2418);
or OR4 (N5185, N5182, N154, N3788, N3470);
nor NOR4 (N5186, N5183, N1771, N368, N1719);
or OR2 (N5187, N5165, N112);
xor XOR2 (N5188, N5185, N3760);
nor NOR4 (N5189, N5131, N1490, N2222, N4459);
xor XOR2 (N5190, N5189, N5016);
xor XOR2 (N5191, N5179, N3326);
nand NAND3 (N5192, N5158, N1367, N3075);
nand NAND3 (N5193, N5184, N2625, N3185);
xor XOR2 (N5194, N5186, N170);
and AND3 (N5195, N5192, N1259, N355);
or OR4 (N5196, N5187, N4333, N432, N4768);
not NOT1 (N5197, N5190);
not NOT1 (N5198, N5197);
buf BUF1 (N5199, N5198);
buf BUF1 (N5200, N5196);
xor XOR2 (N5201, N5191, N2205);
nand NAND4 (N5202, N5169, N841, N2578, N1957);
buf BUF1 (N5203, N5200);
not NOT1 (N5204, N5199);
nand NAND3 (N5205, N5204, N511, N2075);
buf BUF1 (N5206, N5181);
nand NAND3 (N5207, N5203, N826, N762);
not NOT1 (N5208, N5201);
nand NAND4 (N5209, N5202, N940, N5176, N3135);
or OR3 (N5210, N5194, N4608, N1485);
nor NOR2 (N5211, N5188, N3182);
buf BUF1 (N5212, N5211);
xor XOR2 (N5213, N5210, N4358);
and AND2 (N5214, N5212, N3137);
not NOT1 (N5215, N5175);
buf BUF1 (N5216, N5208);
xor XOR2 (N5217, N5195, N4369);
or OR4 (N5218, N5216, N4991, N1380, N4583);
nor NOR4 (N5219, N5213, N1465, N2357, N3435);
or OR2 (N5220, N5207, N3397);
nor NOR4 (N5221, N5193, N1857, N1455, N386);
not NOT1 (N5222, N5206);
buf BUF1 (N5223, N5214);
xor XOR2 (N5224, N5218, N4923);
or OR4 (N5225, N5217, N4664, N2203, N2394);
nor NOR3 (N5226, N5224, N28, N1137);
buf BUF1 (N5227, N5220);
nor NOR4 (N5228, N5225, N4447, N1401, N345);
nand NAND2 (N5229, N5205, N849);
nand NAND3 (N5230, N5215, N3371, N2901);
buf BUF1 (N5231, N5229);
nand NAND2 (N5232, N5230, N3064);
or OR2 (N5233, N5221, N5039);
xor XOR2 (N5234, N5223, N4808);
buf BUF1 (N5235, N5222);
nand NAND4 (N5236, N5235, N420, N655, N460);
or OR4 (N5237, N5236, N218, N2399, N1475);
xor XOR2 (N5238, N5231, N2318);
xor XOR2 (N5239, N5233, N2955);
nand NAND3 (N5240, N5237, N2690, N4889);
and AND3 (N5241, N5227, N2613, N1166);
xor XOR2 (N5242, N5226, N2569);
not NOT1 (N5243, N5209);
nand NAND2 (N5244, N5239, N2845);
nor NOR3 (N5245, N5244, N2628, N3069);
nand NAND2 (N5246, N5228, N1761);
or OR3 (N5247, N5234, N887, N3608);
nand NAND3 (N5248, N5232, N4488, N1832);
or OR2 (N5249, N5242, N4983);
nand NAND2 (N5250, N5241, N4189);
nand NAND4 (N5251, N5219, N1061, N2669, N2267);
not NOT1 (N5252, N5243);
or OR4 (N5253, N5238, N3947, N3064, N2297);
nor NOR4 (N5254, N5246, N1387, N1573, N2728);
xor XOR2 (N5255, N5247, N4731);
or OR2 (N5256, N5254, N64);
and AND4 (N5257, N5245, N406, N785, N4912);
nor NOR3 (N5258, N5250, N4236, N3923);
buf BUF1 (N5259, N5249);
nor NOR3 (N5260, N5259, N4129, N2239);
and AND3 (N5261, N5255, N2084, N45);
nand NAND3 (N5262, N5258, N4412, N4482);
xor XOR2 (N5263, N5251, N3332);
nor NOR4 (N5264, N5256, N3406, N1868, N322);
not NOT1 (N5265, N5264);
xor XOR2 (N5266, N5263, N1881);
nand NAND2 (N5267, N5248, N27);
buf BUF1 (N5268, N5267);
xor XOR2 (N5269, N5252, N3324);
and AND3 (N5270, N5240, N582, N90);
xor XOR2 (N5271, N5268, N169);
nand NAND2 (N5272, N5262, N4678);
or OR3 (N5273, N5257, N321, N657);
not NOT1 (N5274, N5265);
or OR2 (N5275, N5266, N3783);
nor NOR3 (N5276, N5273, N2362, N783);
xor XOR2 (N5277, N5269, N2196);
nor NOR3 (N5278, N5274, N4840, N2762);
and AND3 (N5279, N5276, N313, N987);
nand NAND2 (N5280, N5279, N5056);
buf BUF1 (N5281, N5260);
xor XOR2 (N5282, N5280, N1434);
nor NOR4 (N5283, N5261, N1781, N2403, N3967);
and AND3 (N5284, N5270, N2447, N4314);
not NOT1 (N5285, N5278);
buf BUF1 (N5286, N5275);
buf BUF1 (N5287, N5286);
not NOT1 (N5288, N5253);
nand NAND4 (N5289, N5284, N861, N4252, N4392);
nand NAND4 (N5290, N5281, N1659, N3371, N4420);
and AND2 (N5291, N5283, N1392);
or OR2 (N5292, N5272, N4346);
nor NOR2 (N5293, N5285, N278);
nand NAND2 (N5294, N5287, N1214);
or OR4 (N5295, N5292, N1609, N4723, N2104);
or OR4 (N5296, N5294, N4864, N365, N1763);
not NOT1 (N5297, N5295);
nand NAND2 (N5298, N5291, N1096);
not NOT1 (N5299, N5298);
buf BUF1 (N5300, N5299);
and AND3 (N5301, N5282, N3079, N3304);
not NOT1 (N5302, N5296);
or OR3 (N5303, N5290, N4797, N1799);
and AND4 (N5304, N5297, N2357, N3132, N844);
nand NAND2 (N5305, N5271, N2770);
xor XOR2 (N5306, N5301, N974);
xor XOR2 (N5307, N5306, N2541);
xor XOR2 (N5308, N5302, N4319);
buf BUF1 (N5309, N5308);
not NOT1 (N5310, N5307);
nand NAND2 (N5311, N5288, N3527);
xor XOR2 (N5312, N5277, N2863);
and AND4 (N5313, N5305, N703, N2591, N451);
xor XOR2 (N5314, N5312, N526);
and AND2 (N5315, N5289, N1831);
nor NOR3 (N5316, N5314, N1324, N4976);
and AND3 (N5317, N5313, N1853, N1238);
nand NAND2 (N5318, N5293, N4467);
not NOT1 (N5319, N5318);
nor NOR3 (N5320, N5310, N5095, N668);
or OR4 (N5321, N5320, N7, N4114, N5);
nand NAND3 (N5322, N5316, N2939, N4296);
xor XOR2 (N5323, N5321, N4990);
xor XOR2 (N5324, N5317, N1742);
nand NAND2 (N5325, N5311, N1111);
not NOT1 (N5326, N5323);
buf BUF1 (N5327, N5315);
buf BUF1 (N5328, N5303);
and AND3 (N5329, N5309, N4271, N4094);
xor XOR2 (N5330, N5300, N5133);
and AND4 (N5331, N5324, N4633, N2595, N4649);
or OR3 (N5332, N5328, N1849, N4069);
nor NOR3 (N5333, N5330, N3368, N4042);
nor NOR2 (N5334, N5304, N1813);
nand NAND3 (N5335, N5332, N5313, N3497);
or OR4 (N5336, N5334, N1006, N2837, N5182);
xor XOR2 (N5337, N5329, N234);
nand NAND2 (N5338, N5333, N2432);
and AND2 (N5339, N5319, N4813);
nor NOR2 (N5340, N5325, N5237);
buf BUF1 (N5341, N5339);
and AND3 (N5342, N5326, N1333, N5201);
or OR3 (N5343, N5341, N3988, N2469);
and AND4 (N5344, N5337, N3581, N1099, N2156);
nand NAND2 (N5345, N5344, N4012);
not NOT1 (N5346, N5335);
or OR3 (N5347, N5345, N2902, N1702);
and AND4 (N5348, N5331, N3178, N2517, N4681);
or OR3 (N5349, N5327, N2384, N4968);
or OR4 (N5350, N5349, N2730, N3528, N5005);
xor XOR2 (N5351, N5347, N4842);
buf BUF1 (N5352, N5336);
and AND2 (N5353, N5352, N5064);
or OR4 (N5354, N5342, N4067, N2712, N4257);
nand NAND4 (N5355, N5343, N5031, N5106, N826);
buf BUF1 (N5356, N5340);
xor XOR2 (N5357, N5354, N4614);
and AND3 (N5358, N5355, N3891, N1928);
not NOT1 (N5359, N5353);
xor XOR2 (N5360, N5356, N3059);
not NOT1 (N5361, N5359);
not NOT1 (N5362, N5357);
or OR4 (N5363, N5358, N2744, N3546, N1607);
xor XOR2 (N5364, N5362, N51);
and AND2 (N5365, N5346, N4493);
nor NOR3 (N5366, N5364, N4673, N2600);
or OR3 (N5367, N5363, N4466, N2124);
xor XOR2 (N5368, N5365, N4141);
or OR3 (N5369, N5350, N2333, N270);
nor NOR4 (N5370, N5366, N4591, N261, N2654);
and AND2 (N5371, N5351, N2338);
or OR4 (N5372, N5361, N3143, N1281, N4284);
buf BUF1 (N5373, N5372);
buf BUF1 (N5374, N5369);
nand NAND2 (N5375, N5322, N3775);
and AND4 (N5376, N5367, N4611, N1120, N542);
xor XOR2 (N5377, N5373, N3950);
or OR3 (N5378, N5338, N4690, N590);
not NOT1 (N5379, N5368);
buf BUF1 (N5380, N5378);
nand NAND2 (N5381, N5348, N1623);
or OR3 (N5382, N5360, N2254, N1218);
and AND3 (N5383, N5380, N2145, N2099);
nor NOR3 (N5384, N5370, N3515, N4103);
and AND4 (N5385, N5377, N4113, N3964, N2538);
and AND4 (N5386, N5375, N2772, N4157, N3864);
not NOT1 (N5387, N5382);
buf BUF1 (N5388, N5383);
not NOT1 (N5389, N5376);
or OR3 (N5390, N5374, N2007, N4408);
buf BUF1 (N5391, N5384);
xor XOR2 (N5392, N5379, N4414);
buf BUF1 (N5393, N5390);
nand NAND2 (N5394, N5381, N4859);
or OR3 (N5395, N5391, N2147, N1016);
buf BUF1 (N5396, N5388);
and AND2 (N5397, N5389, N1188);
or OR4 (N5398, N5397, N3540, N1629, N5012);
nand NAND4 (N5399, N5385, N728, N5249, N2330);
buf BUF1 (N5400, N5386);
not NOT1 (N5401, N5393);
nand NAND4 (N5402, N5398, N5135, N3106, N4856);
nand NAND2 (N5403, N5395, N1462);
nor NOR3 (N5404, N5399, N4490, N4813);
nand NAND4 (N5405, N5403, N4130, N892, N932);
buf BUF1 (N5406, N5371);
nor NOR2 (N5407, N5404, N4228);
xor XOR2 (N5408, N5402, N5037);
xor XOR2 (N5409, N5407, N4325);
xor XOR2 (N5410, N5409, N3490);
nand NAND2 (N5411, N5394, N718);
xor XOR2 (N5412, N5408, N3430);
not NOT1 (N5413, N5405);
nand NAND4 (N5414, N5396, N5261, N2426, N2795);
nor NOR2 (N5415, N5401, N49);
nor NOR2 (N5416, N5415, N3291);
xor XOR2 (N5417, N5387, N5244);
nand NAND3 (N5418, N5400, N1117, N4521);
nand NAND3 (N5419, N5414, N882, N1645);
not NOT1 (N5420, N5392);
or OR3 (N5421, N5406, N2636, N951);
not NOT1 (N5422, N5410);
buf BUF1 (N5423, N5418);
nor NOR4 (N5424, N5420, N4773, N4287, N2624);
nand NAND3 (N5425, N5422, N1969, N5270);
buf BUF1 (N5426, N5416);
or OR3 (N5427, N5411, N3321, N5115);
xor XOR2 (N5428, N5423, N2659);
nand NAND4 (N5429, N5417, N4600, N3748, N820);
xor XOR2 (N5430, N5429, N4674);
not NOT1 (N5431, N5425);
nand NAND4 (N5432, N5419, N1814, N4392, N285);
xor XOR2 (N5433, N5426, N3652);
not NOT1 (N5434, N5430);
and AND4 (N5435, N5432, N2328, N2214, N2191);
xor XOR2 (N5436, N5412, N4666);
nand NAND2 (N5437, N5421, N2575);
buf BUF1 (N5438, N5435);
and AND4 (N5439, N5431, N4246, N3646, N1856);
not NOT1 (N5440, N5438);
buf BUF1 (N5441, N5413);
and AND2 (N5442, N5424, N3472);
and AND4 (N5443, N5434, N1286, N5278, N2320);
xor XOR2 (N5444, N5439, N3150);
not NOT1 (N5445, N5428);
buf BUF1 (N5446, N5441);
not NOT1 (N5447, N5444);
or OR2 (N5448, N5433, N2884);
nor NOR2 (N5449, N5442, N5433);
or OR2 (N5450, N5445, N2599);
buf BUF1 (N5451, N5450);
nand NAND4 (N5452, N5440, N2466, N4410, N3462);
not NOT1 (N5453, N5448);
nand NAND4 (N5454, N5453, N2463, N3857, N844);
not NOT1 (N5455, N5427);
buf BUF1 (N5456, N5447);
nor NOR4 (N5457, N5436, N3623, N1264, N1694);
or OR4 (N5458, N5452, N2726, N3851, N3955);
xor XOR2 (N5459, N5457, N1591);
and AND3 (N5460, N5449, N4627, N1903);
or OR4 (N5461, N5437, N1452, N730, N3860);
nor NOR2 (N5462, N5461, N1450);
xor XOR2 (N5463, N5454, N5175);
not NOT1 (N5464, N5451);
buf BUF1 (N5465, N5443);
nand NAND4 (N5466, N5446, N4660, N2964, N201);
nor NOR3 (N5467, N5458, N4924, N2934);
nand NAND4 (N5468, N5455, N873, N4763, N4444);
not NOT1 (N5469, N5466);
nand NAND2 (N5470, N5468, N4874);
nor NOR2 (N5471, N5469, N288);
and AND3 (N5472, N5467, N2248, N247);
not NOT1 (N5473, N5456);
nor NOR2 (N5474, N5460, N2252);
nand NAND3 (N5475, N5471, N1235, N2131);
xor XOR2 (N5476, N5462, N1260);
and AND4 (N5477, N5464, N836, N3382, N1254);
and AND2 (N5478, N5476, N4788);
not NOT1 (N5479, N5472);
not NOT1 (N5480, N5478);
or OR3 (N5481, N5479, N358, N5230);
buf BUF1 (N5482, N5480);
buf BUF1 (N5483, N5465);
xor XOR2 (N5484, N5463, N1478);
nand NAND4 (N5485, N5459, N3125, N3215, N2179);
nand NAND2 (N5486, N5475, N133);
and AND4 (N5487, N5484, N2969, N3469, N2469);
not NOT1 (N5488, N5485);
nor NOR2 (N5489, N5483, N2039);
and AND4 (N5490, N5489, N3034, N5072, N5432);
xor XOR2 (N5491, N5474, N25);
buf BUF1 (N5492, N5486);
nor NOR2 (N5493, N5482, N3940);
or OR4 (N5494, N5487, N1723, N2643, N3172);
nand NAND4 (N5495, N5470, N3146, N3137, N4124);
and AND3 (N5496, N5493, N3154, N5229);
nor NOR2 (N5497, N5491, N1337);
xor XOR2 (N5498, N5496, N3620);
nand NAND2 (N5499, N5488, N3249);
not NOT1 (N5500, N5492);
xor XOR2 (N5501, N5495, N1613);
buf BUF1 (N5502, N5497);
and AND2 (N5503, N5473, N3165);
nand NAND3 (N5504, N5481, N3504, N4580);
nor NOR3 (N5505, N5490, N2109, N106);
xor XOR2 (N5506, N5505, N162);
and AND2 (N5507, N5502, N4232);
nor NOR2 (N5508, N5507, N4825);
buf BUF1 (N5509, N5503);
and AND3 (N5510, N5477, N406, N57);
buf BUF1 (N5511, N5501);
xor XOR2 (N5512, N5500, N871);
nand NAND2 (N5513, N5510, N1332);
xor XOR2 (N5514, N5494, N5291);
not NOT1 (N5515, N5499);
nand NAND2 (N5516, N5509, N4291);
buf BUF1 (N5517, N5513);
or OR2 (N5518, N5515, N1192);
not NOT1 (N5519, N5511);
xor XOR2 (N5520, N5516, N3355);
not NOT1 (N5521, N5517);
nand NAND4 (N5522, N5514, N1027, N4079, N3669);
buf BUF1 (N5523, N5504);
and AND3 (N5524, N5508, N2478, N5377);
not NOT1 (N5525, N5506);
not NOT1 (N5526, N5518);
or OR3 (N5527, N5526, N2269, N1968);
xor XOR2 (N5528, N5525, N3027);
xor XOR2 (N5529, N5521, N5321);
nor NOR4 (N5530, N5523, N2550, N1831, N4315);
or OR2 (N5531, N5519, N386);
xor XOR2 (N5532, N5527, N899);
xor XOR2 (N5533, N5531, N1017);
not NOT1 (N5534, N5532);
nand NAND4 (N5535, N5533, N4874, N2824, N5385);
buf BUF1 (N5536, N5520);
buf BUF1 (N5537, N5534);
nand NAND4 (N5538, N5522, N4120, N2414, N5028);
nor NOR3 (N5539, N5537, N3734, N2115);
and AND4 (N5540, N5528, N1455, N4634, N775);
nor NOR4 (N5541, N5530, N2733, N1893, N3294);
nor NOR2 (N5542, N5512, N3072);
and AND3 (N5543, N5524, N1267, N1311);
not NOT1 (N5544, N5535);
xor XOR2 (N5545, N5498, N4373);
buf BUF1 (N5546, N5536);
xor XOR2 (N5547, N5545, N865);
not NOT1 (N5548, N5543);
nand NAND4 (N5549, N5541, N19, N3161, N1755);
nor NOR4 (N5550, N5547, N1097, N847, N3314);
xor XOR2 (N5551, N5546, N3794);
and AND2 (N5552, N5542, N2585);
and AND2 (N5553, N5550, N4037);
buf BUF1 (N5554, N5538);
nor NOR4 (N5555, N5548, N2613, N175, N4573);
nand NAND3 (N5556, N5540, N3071, N1300);
xor XOR2 (N5557, N5553, N2520);
nor NOR4 (N5558, N5557, N3696, N3956, N2434);
nand NAND4 (N5559, N5555, N5098, N4356, N284);
nor NOR3 (N5560, N5559, N833, N838);
xor XOR2 (N5561, N5552, N2375);
and AND3 (N5562, N5529, N2474, N1515);
buf BUF1 (N5563, N5539);
or OR4 (N5564, N5544, N3337, N5309, N1723);
and AND4 (N5565, N5561, N4384, N4778, N2732);
not NOT1 (N5566, N5562);
and AND3 (N5567, N5564, N3694, N5393);
buf BUF1 (N5568, N5554);
not NOT1 (N5569, N5556);
nand NAND3 (N5570, N5565, N290, N1898);
nor NOR3 (N5571, N5558, N5138, N4664);
xor XOR2 (N5572, N5567, N4588);
buf BUF1 (N5573, N5566);
and AND2 (N5574, N5563, N4963);
xor XOR2 (N5575, N5549, N1418);
nor NOR4 (N5576, N5572, N3137, N1752, N1839);
not NOT1 (N5577, N5571);
nand NAND4 (N5578, N5573, N2974, N1376, N353);
not NOT1 (N5579, N5577);
nand NAND2 (N5580, N5569, N5048);
buf BUF1 (N5581, N5580);
nor NOR3 (N5582, N5579, N5250, N2604);
xor XOR2 (N5583, N5576, N1659);
and AND3 (N5584, N5575, N2377, N3589);
buf BUF1 (N5585, N5584);
nor NOR3 (N5586, N5551, N4929, N1111);
xor XOR2 (N5587, N5574, N3628);
not NOT1 (N5588, N5570);
not NOT1 (N5589, N5582);
not NOT1 (N5590, N5568);
nand NAND2 (N5591, N5560, N2972);
or OR4 (N5592, N5591, N382, N2697, N4193);
buf BUF1 (N5593, N5588);
or OR3 (N5594, N5581, N2512, N3739);
buf BUF1 (N5595, N5578);
and AND2 (N5596, N5593, N1984);
or OR3 (N5597, N5594, N1628, N1119);
buf BUF1 (N5598, N5585);
nand NAND2 (N5599, N5587, N1914);
xor XOR2 (N5600, N5597, N3147);
buf BUF1 (N5601, N5592);
xor XOR2 (N5602, N5599, N928);
xor XOR2 (N5603, N5598, N2542);
xor XOR2 (N5604, N5596, N5133);
and AND2 (N5605, N5603, N995);
or OR3 (N5606, N5589, N2900, N1421);
buf BUF1 (N5607, N5601);
nand NAND2 (N5608, N5607, N701);
xor XOR2 (N5609, N5608, N5372);
or OR3 (N5610, N5590, N4485, N450);
buf BUF1 (N5611, N5595);
and AND3 (N5612, N5600, N4679, N2359);
not NOT1 (N5613, N5586);
buf BUF1 (N5614, N5609);
buf BUF1 (N5615, N5605);
xor XOR2 (N5616, N5606, N4013);
nor NOR4 (N5617, N5602, N3058, N4531, N143);
and AND4 (N5618, N5604, N5466, N3220, N4764);
buf BUF1 (N5619, N5613);
buf BUF1 (N5620, N5615);
and AND3 (N5621, N5617, N5126, N2079);
nor NOR3 (N5622, N5620, N3546, N5178);
not NOT1 (N5623, N5610);
nor NOR4 (N5624, N5611, N2952, N5534, N4005);
buf BUF1 (N5625, N5623);
xor XOR2 (N5626, N5618, N5477);
not NOT1 (N5627, N5625);
nor NOR3 (N5628, N5622, N2976, N5310);
and AND3 (N5629, N5619, N1344, N2704);
buf BUF1 (N5630, N5627);
buf BUF1 (N5631, N5628);
buf BUF1 (N5632, N5626);
and AND3 (N5633, N5631, N2653, N2465);
nor NOR3 (N5634, N5612, N3875, N4010);
buf BUF1 (N5635, N5616);
nand NAND4 (N5636, N5624, N3429, N390, N3464);
xor XOR2 (N5637, N5632, N2311);
nand NAND4 (N5638, N5630, N1771, N4386, N207);
and AND2 (N5639, N5637, N1928);
or OR2 (N5640, N5638, N89);
not NOT1 (N5641, N5640);
or OR3 (N5642, N5641, N4015, N5603);
xor XOR2 (N5643, N5642, N3059);
xor XOR2 (N5644, N5636, N1126);
and AND2 (N5645, N5614, N4698);
buf BUF1 (N5646, N5629);
nand NAND2 (N5647, N5639, N1502);
and AND4 (N5648, N5644, N110, N783, N5200);
nor NOR3 (N5649, N5645, N2768, N5535);
and AND2 (N5650, N5621, N3466);
or OR3 (N5651, N5648, N3939, N4290);
or OR4 (N5652, N5646, N491, N1001, N5412);
or OR3 (N5653, N5633, N4607, N223);
nor NOR2 (N5654, N5650, N2230);
not NOT1 (N5655, N5651);
nand NAND4 (N5656, N5583, N5394, N2451, N5248);
nor NOR3 (N5657, N5655, N4049, N970);
or OR2 (N5658, N5634, N4775);
xor XOR2 (N5659, N5652, N2788);
buf BUF1 (N5660, N5635);
nand NAND4 (N5661, N5658, N3649, N2608, N5164);
nand NAND3 (N5662, N5647, N5336, N754);
or OR3 (N5663, N5656, N1950, N1723);
or OR3 (N5664, N5643, N4359, N2021);
buf BUF1 (N5665, N5660);
buf BUF1 (N5666, N5657);
nand NAND3 (N5667, N5649, N631, N5283);
nand NAND2 (N5668, N5663, N4688);
nand NAND2 (N5669, N5662, N3705);
nand NAND4 (N5670, N5664, N3426, N3574, N1666);
or OR2 (N5671, N5669, N125);
or OR3 (N5672, N5670, N1626, N169);
nor NOR4 (N5673, N5665, N939, N3124, N4724);
xor XOR2 (N5674, N5671, N5090);
and AND3 (N5675, N5667, N5620, N1972);
or OR3 (N5676, N5659, N4724, N2920);
or OR4 (N5677, N5653, N2697, N4865, N3862);
and AND3 (N5678, N5654, N1656, N4486);
xor XOR2 (N5679, N5666, N4854);
xor XOR2 (N5680, N5661, N2524);
and AND2 (N5681, N5677, N1193);
buf BUF1 (N5682, N5673);
xor XOR2 (N5683, N5675, N4460);
nor NOR4 (N5684, N5683, N2684, N1342, N5367);
not NOT1 (N5685, N5668);
buf BUF1 (N5686, N5681);
xor XOR2 (N5687, N5682, N2779);
and AND2 (N5688, N5672, N1472);
not NOT1 (N5689, N5680);
or OR2 (N5690, N5685, N707);
not NOT1 (N5691, N5690);
or OR2 (N5692, N5688, N5198);
nor NOR3 (N5693, N5679, N294, N2067);
buf BUF1 (N5694, N5692);
buf BUF1 (N5695, N5694);
xor XOR2 (N5696, N5678, N1061);
and AND4 (N5697, N5696, N1475, N1750, N2381);
xor XOR2 (N5698, N5689, N1368);
or OR4 (N5699, N5687, N1095, N3430, N2232);
xor XOR2 (N5700, N5695, N2192);
and AND3 (N5701, N5699, N1998, N3956);
buf BUF1 (N5702, N5676);
xor XOR2 (N5703, N5697, N4773);
buf BUF1 (N5704, N5686);
not NOT1 (N5705, N5693);
not NOT1 (N5706, N5684);
xor XOR2 (N5707, N5698, N1529);
buf BUF1 (N5708, N5701);
or OR4 (N5709, N5702, N4418, N4106, N3923);
or OR4 (N5710, N5674, N2770, N3492, N1368);
nand NAND3 (N5711, N5709, N431, N2709);
or OR3 (N5712, N5711, N195, N558);
nor NOR3 (N5713, N5706, N19, N2304);
nor NOR2 (N5714, N5704, N2627);
buf BUF1 (N5715, N5714);
not NOT1 (N5716, N5712);
nand NAND3 (N5717, N5691, N5646, N2168);
not NOT1 (N5718, N5717);
and AND2 (N5719, N5710, N174);
xor XOR2 (N5720, N5713, N3237);
buf BUF1 (N5721, N5703);
buf BUF1 (N5722, N5708);
buf BUF1 (N5723, N5719);
xor XOR2 (N5724, N5720, N4132);
or OR3 (N5725, N5715, N3683, N4999);
xor XOR2 (N5726, N5700, N3927);
xor XOR2 (N5727, N5723, N2315);
xor XOR2 (N5728, N5727, N3407);
not NOT1 (N5729, N5707);
nand NAND2 (N5730, N5705, N3335);
not NOT1 (N5731, N5728);
nand NAND4 (N5732, N5725, N4361, N84, N5015);
buf BUF1 (N5733, N5721);
xor XOR2 (N5734, N5731, N620);
nand NAND4 (N5735, N5733, N2350, N4112, N3301);
nand NAND4 (N5736, N5716, N2716, N954, N3095);
buf BUF1 (N5737, N5735);
and AND2 (N5738, N5718, N584);
nor NOR3 (N5739, N5738, N3113, N969);
nor NOR3 (N5740, N5734, N2568, N3349);
not NOT1 (N5741, N5732);
not NOT1 (N5742, N5724);
nor NOR4 (N5743, N5726, N75, N4478, N5305);
nand NAND3 (N5744, N5742, N1154, N2013);
and AND3 (N5745, N5739, N3499, N1451);
and AND3 (N5746, N5741, N2972, N5548);
and AND3 (N5747, N5737, N1692, N1971);
and AND3 (N5748, N5740, N256, N4046);
nor NOR4 (N5749, N5747, N226, N2356, N3251);
or OR2 (N5750, N5729, N3336);
and AND4 (N5751, N5744, N644, N296, N3254);
buf BUF1 (N5752, N5746);
nand NAND4 (N5753, N5752, N133, N4332, N5101);
buf BUF1 (N5754, N5753);
or OR2 (N5755, N5743, N5120);
nor NOR2 (N5756, N5749, N185);
and AND4 (N5757, N5756, N1698, N2446, N559);
nor NOR2 (N5758, N5755, N1239);
nor NOR2 (N5759, N5745, N491);
not NOT1 (N5760, N5754);
and AND2 (N5761, N5758, N472);
or OR2 (N5762, N5722, N1328);
not NOT1 (N5763, N5748);
nand NAND4 (N5764, N5750, N450, N9, N4793);
nand NAND2 (N5765, N5759, N1261);
not NOT1 (N5766, N5763);
nor NOR3 (N5767, N5761, N5348, N301);
and AND4 (N5768, N5765, N1283, N2037, N978);
nand NAND4 (N5769, N5768, N76, N268, N3379);
nand NAND4 (N5770, N5769, N3756, N3759, N274);
and AND2 (N5771, N5760, N3682);
buf BUF1 (N5772, N5771);
buf BUF1 (N5773, N5751);
or OR3 (N5774, N5730, N3529, N1171);
buf BUF1 (N5775, N5736);
or OR3 (N5776, N5757, N4589, N205);
xor XOR2 (N5777, N5773, N3827);
nor NOR2 (N5778, N5777, N2895);
and AND3 (N5779, N5774, N2148, N4648);
or OR3 (N5780, N5764, N417, N5300);
or OR4 (N5781, N5762, N2525, N2580, N1696);
xor XOR2 (N5782, N5778, N554);
nand NAND4 (N5783, N5782, N3450, N327, N250);
and AND4 (N5784, N5766, N2811, N4383, N1576);
not NOT1 (N5785, N5779);
and AND2 (N5786, N5770, N2657);
buf BUF1 (N5787, N5785);
xor XOR2 (N5788, N5767, N2214);
buf BUF1 (N5789, N5776);
not NOT1 (N5790, N5781);
xor XOR2 (N5791, N5775, N4572);
nand NAND4 (N5792, N5788, N2562, N2107, N3002);
nor NOR3 (N5793, N5790, N4741, N613);
and AND3 (N5794, N5792, N3670, N2761);
buf BUF1 (N5795, N5789);
xor XOR2 (N5796, N5783, N5451);
nand NAND4 (N5797, N5787, N461, N1792, N556);
and AND4 (N5798, N5796, N888, N2977, N3661);
or OR2 (N5799, N5791, N5008);
nand NAND2 (N5800, N5784, N4952);
nand NAND2 (N5801, N5780, N4895);
nor NOR2 (N5802, N5800, N2691);
and AND3 (N5803, N5801, N845, N50);
or OR4 (N5804, N5797, N2620, N2550, N1384);
and AND2 (N5805, N5793, N3833);
or OR2 (N5806, N5798, N3301);
or OR3 (N5807, N5795, N2822, N4045);
not NOT1 (N5808, N5807);
nor NOR2 (N5809, N5802, N3943);
or OR2 (N5810, N5804, N2257);
and AND3 (N5811, N5803, N3589, N692);
xor XOR2 (N5812, N5794, N1820);
not NOT1 (N5813, N5799);
buf BUF1 (N5814, N5811);
and AND3 (N5815, N5809, N4836, N3570);
nor NOR3 (N5816, N5808, N5044, N4235);
nand NAND2 (N5817, N5812, N5271);
buf BUF1 (N5818, N5814);
nor NOR2 (N5819, N5817, N3551);
nand NAND2 (N5820, N5813, N1023);
not NOT1 (N5821, N5805);
or OR3 (N5822, N5810, N4922, N4748);
nor NOR4 (N5823, N5786, N479, N2331, N2006);
buf BUF1 (N5824, N5816);
or OR4 (N5825, N5818, N4966, N2383, N1019);
and AND4 (N5826, N5821, N4602, N4745, N1658);
not NOT1 (N5827, N5825);
buf BUF1 (N5828, N5772);
nor NOR3 (N5829, N5806, N3886, N3963);
xor XOR2 (N5830, N5815, N275);
buf BUF1 (N5831, N5824);
nor NOR3 (N5832, N5831, N4659, N212);
xor XOR2 (N5833, N5823, N3938);
or OR3 (N5834, N5833, N2944, N1967);
buf BUF1 (N5835, N5820);
buf BUF1 (N5836, N5835);
and AND3 (N5837, N5832, N3751, N5686);
and AND3 (N5838, N5836, N770, N1999);
xor XOR2 (N5839, N5827, N5019);
and AND3 (N5840, N5830, N379, N682);
and AND4 (N5841, N5837, N5823, N4818, N2324);
not NOT1 (N5842, N5822);
nor NOR4 (N5843, N5842, N3208, N3564, N1562);
xor XOR2 (N5844, N5838, N3222);
and AND3 (N5845, N5819, N3518, N2480);
nor NOR4 (N5846, N5841, N3782, N5543, N705);
not NOT1 (N5847, N5834);
and AND3 (N5848, N5845, N193, N4744);
buf BUF1 (N5849, N5829);
nor NOR3 (N5850, N5846, N1319, N1430);
buf BUF1 (N5851, N5828);
buf BUF1 (N5852, N5849);
not NOT1 (N5853, N5848);
nand NAND3 (N5854, N5843, N4690, N3375);
nand NAND3 (N5855, N5851, N795, N972);
nand NAND4 (N5856, N5854, N433, N93, N4507);
xor XOR2 (N5857, N5850, N4583);
buf BUF1 (N5858, N5839);
buf BUF1 (N5859, N5844);
nor NOR4 (N5860, N5855, N218, N4670, N1124);
nor NOR2 (N5861, N5826, N2671);
xor XOR2 (N5862, N5853, N608);
xor XOR2 (N5863, N5840, N2999);
not NOT1 (N5864, N5859);
not NOT1 (N5865, N5847);
and AND4 (N5866, N5860, N1267, N93, N2052);
not NOT1 (N5867, N5856);
buf BUF1 (N5868, N5867);
buf BUF1 (N5869, N5861);
not NOT1 (N5870, N5863);
buf BUF1 (N5871, N5864);
not NOT1 (N5872, N5857);
nor NOR4 (N5873, N5868, N610, N4349, N4357);
buf BUF1 (N5874, N5873);
nor NOR3 (N5875, N5862, N1226, N4604);
xor XOR2 (N5876, N5874, N5044);
or OR2 (N5877, N5865, N1963);
not NOT1 (N5878, N5870);
and AND2 (N5879, N5878, N1122);
nor NOR2 (N5880, N5852, N5015);
and AND2 (N5881, N5869, N3668);
nor NOR4 (N5882, N5880, N5040, N385, N3090);
buf BUF1 (N5883, N5882);
nand NAND2 (N5884, N5875, N3375);
xor XOR2 (N5885, N5858, N2137);
nor NOR3 (N5886, N5879, N3011, N894);
nand NAND4 (N5887, N5871, N1821, N3039, N5877);
buf BUF1 (N5888, N5499);
not NOT1 (N5889, N5883);
and AND4 (N5890, N5885, N3265, N2689, N702);
nand NAND2 (N5891, N5888, N2695);
or OR4 (N5892, N5891, N150, N710, N346);
or OR2 (N5893, N5890, N5682);
buf BUF1 (N5894, N5887);
xor XOR2 (N5895, N5889, N3577);
and AND4 (N5896, N5866, N1370, N4539, N5632);
xor XOR2 (N5897, N5876, N419);
not NOT1 (N5898, N5893);
or OR2 (N5899, N5895, N2299);
xor XOR2 (N5900, N5881, N3784);
and AND3 (N5901, N5897, N3189, N1384);
buf BUF1 (N5902, N5872);
not NOT1 (N5903, N5901);
xor XOR2 (N5904, N5899, N4236);
and AND4 (N5905, N5896, N1920, N5838, N2706);
and AND2 (N5906, N5905, N1308);
or OR4 (N5907, N5900, N4177, N5184, N3129);
and AND4 (N5908, N5884, N5326, N2272, N2226);
or OR3 (N5909, N5894, N5023, N1080);
not NOT1 (N5910, N5907);
not NOT1 (N5911, N5906);
buf BUF1 (N5912, N5904);
buf BUF1 (N5913, N5911);
nand NAND3 (N5914, N5903, N362, N4373);
and AND4 (N5915, N5913, N1853, N2845, N174);
nor NOR4 (N5916, N5902, N1484, N1526, N1720);
nand NAND2 (N5917, N5909, N3184);
and AND2 (N5918, N5917, N510);
nand NAND4 (N5919, N5915, N4427, N406, N4281);
not NOT1 (N5920, N5919);
nor NOR2 (N5921, N5914, N4862);
nor NOR4 (N5922, N5908, N4638, N5737, N5025);
or OR4 (N5923, N5912, N4232, N431, N5786);
and AND3 (N5924, N5923, N2756, N5912);
nand NAND4 (N5925, N5924, N3668, N4310, N4315);
and AND4 (N5926, N5922, N4330, N866, N4084);
xor XOR2 (N5927, N5918, N2507);
and AND3 (N5928, N5927, N1174, N3770);
not NOT1 (N5929, N5886);
buf BUF1 (N5930, N5926);
nor NOR2 (N5931, N5898, N5765);
nand NAND3 (N5932, N5920, N3066, N5837);
xor XOR2 (N5933, N5929, N3216);
xor XOR2 (N5934, N5932, N3758);
or OR2 (N5935, N5921, N2844);
nand NAND3 (N5936, N5916, N3318, N229);
nor NOR3 (N5937, N5928, N4741, N5548);
nand NAND2 (N5938, N5910, N5093);
and AND4 (N5939, N5934, N384, N1541, N33);
and AND3 (N5940, N5931, N2116, N4230);
xor XOR2 (N5941, N5936, N3672);
nand NAND3 (N5942, N5933, N1456, N2344);
nor NOR3 (N5943, N5937, N3208, N1696);
not NOT1 (N5944, N5892);
and AND2 (N5945, N5930, N4564);
and AND4 (N5946, N5938, N518, N3846, N704);
nor NOR3 (N5947, N5946, N449, N231);
or OR4 (N5948, N5940, N3137, N5457, N3558);
xor XOR2 (N5949, N5935, N2059);
nor NOR2 (N5950, N5939, N1375);
or OR2 (N5951, N5941, N3064);
nor NOR2 (N5952, N5942, N76);
buf BUF1 (N5953, N5947);
xor XOR2 (N5954, N5949, N4192);
nand NAND2 (N5955, N5950, N5467);
buf BUF1 (N5956, N5925);
buf BUF1 (N5957, N5943);
and AND2 (N5958, N5957, N4461);
and AND3 (N5959, N5952, N3001, N4421);
not NOT1 (N5960, N5944);
or OR4 (N5961, N5959, N1839, N3942, N3793);
xor XOR2 (N5962, N5951, N1740);
xor XOR2 (N5963, N5953, N509);
nor NOR3 (N5964, N5961, N821, N5068);
nor NOR3 (N5965, N5964, N2725, N2647);
nand NAND2 (N5966, N5956, N1134);
nor NOR2 (N5967, N5962, N4498);
and AND4 (N5968, N5966, N2483, N5210, N3937);
and AND3 (N5969, N5968, N2191, N3989);
and AND2 (N5970, N5955, N1690);
xor XOR2 (N5971, N5967, N164);
nand NAND3 (N5972, N5948, N2200, N355);
or OR3 (N5973, N5958, N4137, N2226);
nor NOR4 (N5974, N5971, N5832, N2047, N1146);
xor XOR2 (N5975, N5974, N3707);
or OR2 (N5976, N5960, N3198);
and AND2 (N5977, N5973, N5871);
nand NAND2 (N5978, N5977, N5245);
nor NOR3 (N5979, N5972, N3435, N26);
not NOT1 (N5980, N5963);
and AND2 (N5981, N5954, N4797);
or OR4 (N5982, N5975, N1811, N2484, N4555);
or OR3 (N5983, N5965, N4745, N646);
and AND4 (N5984, N5970, N2232, N714, N3551);
not NOT1 (N5985, N5980);
and AND4 (N5986, N5982, N1494, N5275, N1811);
not NOT1 (N5987, N5978);
or OR2 (N5988, N5983, N2964);
and AND3 (N5989, N5984, N1438, N5731);
or OR4 (N5990, N5988, N4141, N114, N4446);
not NOT1 (N5991, N5985);
and AND4 (N5992, N5945, N1654, N5361, N5916);
buf BUF1 (N5993, N5992);
buf BUF1 (N5994, N5993);
xor XOR2 (N5995, N5986, N5951);
and AND2 (N5996, N5981, N2339);
xor XOR2 (N5997, N5969, N1634);
nor NOR2 (N5998, N5997, N4114);
not NOT1 (N5999, N5994);
nor NOR2 (N6000, N5991, N614);
and AND3 (N6001, N6000, N5502, N2562);
not NOT1 (N6002, N5999);
buf BUF1 (N6003, N5989);
nand NAND4 (N6004, N6002, N4084, N5948, N575);
not NOT1 (N6005, N5995);
nand NAND2 (N6006, N6004, N2924);
xor XOR2 (N6007, N5998, N448);
not NOT1 (N6008, N5996);
xor XOR2 (N6009, N6001, N5720);
buf BUF1 (N6010, N6007);
or OR3 (N6011, N6008, N2866, N229);
nor NOR2 (N6012, N6010, N4450);
nor NOR4 (N6013, N5990, N5664, N4778, N5207);
nand NAND2 (N6014, N6003, N3148);
and AND3 (N6015, N5987, N5942, N413);
not NOT1 (N6016, N6014);
not NOT1 (N6017, N5976);
xor XOR2 (N6018, N6011, N3910);
and AND3 (N6019, N6006, N4737, N5905);
not NOT1 (N6020, N5979);
nand NAND3 (N6021, N6020, N4199, N4309);
and AND3 (N6022, N6019, N4604, N1841);
xor XOR2 (N6023, N6018, N4723);
nand NAND2 (N6024, N6022, N5122);
and AND4 (N6025, N6023, N5422, N3838, N3203);
and AND2 (N6026, N6012, N3565);
buf BUF1 (N6027, N6009);
nand NAND4 (N6028, N6024, N2591, N1169, N3387);
xor XOR2 (N6029, N6027, N5520);
nand NAND4 (N6030, N6025, N359, N2500, N3005);
buf BUF1 (N6031, N6026);
and AND4 (N6032, N6016, N405, N5419, N5121);
or OR3 (N6033, N6021, N1510, N2335);
and AND2 (N6034, N6028, N1013);
nand NAND2 (N6035, N6017, N2999);
nor NOR3 (N6036, N6013, N3172, N5503);
nor NOR2 (N6037, N6034, N1982);
or OR4 (N6038, N6030, N2184, N5641, N34);
not NOT1 (N6039, N6029);
nor NOR3 (N6040, N6036, N1327, N5085);
xor XOR2 (N6041, N6037, N3383);
nor NOR2 (N6042, N6041, N1156);
and AND2 (N6043, N6015, N2074);
and AND4 (N6044, N6039, N5996, N5438, N4087);
or OR3 (N6045, N6044, N3126, N2781);
or OR4 (N6046, N6035, N4190, N2726, N2608);
nand NAND2 (N6047, N6042, N4133);
buf BUF1 (N6048, N6040);
nand NAND4 (N6049, N6033, N1004, N5306, N3682);
nor NOR4 (N6050, N6005, N1385, N4844, N113);
nand NAND2 (N6051, N6045, N2551);
nor NOR3 (N6052, N6050, N2730, N3361);
xor XOR2 (N6053, N6046, N3256);
nor NOR4 (N6054, N6048, N2647, N5613, N3376);
not NOT1 (N6055, N6047);
xor XOR2 (N6056, N6051, N4132);
and AND3 (N6057, N6056, N198, N5950);
nor NOR2 (N6058, N6049, N2762);
not NOT1 (N6059, N6052);
not NOT1 (N6060, N6053);
xor XOR2 (N6061, N6060, N400);
not NOT1 (N6062, N6059);
nor NOR2 (N6063, N6038, N801);
nor NOR4 (N6064, N6057, N1019, N5997, N4264);
nand NAND3 (N6065, N6062, N3, N790);
nor NOR4 (N6066, N6063, N3009, N3185, N2375);
xor XOR2 (N6067, N6066, N5621);
xor XOR2 (N6068, N6061, N3340);
nand NAND4 (N6069, N6068, N2587, N4766, N485);
nand NAND2 (N6070, N6064, N3841);
and AND2 (N6071, N6031, N2860);
not NOT1 (N6072, N6043);
or OR4 (N6073, N6065, N5040, N5747, N3134);
buf BUF1 (N6074, N6069);
nand NAND4 (N6075, N6073, N3880, N5270, N549);
nand NAND2 (N6076, N6071, N1105);
and AND2 (N6077, N6032, N4089);
nand NAND3 (N6078, N6067, N1057, N3906);
and AND4 (N6079, N6054, N5286, N1812, N4395);
xor XOR2 (N6080, N6075, N3501);
and AND3 (N6081, N6078, N2042, N4068);
xor XOR2 (N6082, N6080, N4172);
xor XOR2 (N6083, N6076, N3500);
nand NAND4 (N6084, N6058, N4744, N4482, N3588);
not NOT1 (N6085, N6072);
not NOT1 (N6086, N6084);
not NOT1 (N6087, N6085);
buf BUF1 (N6088, N6077);
xor XOR2 (N6089, N6081, N4436);
or OR4 (N6090, N6079, N741, N3491, N78);
and AND4 (N6091, N6088, N2513, N3750, N2048);
not NOT1 (N6092, N6082);
or OR2 (N6093, N6087, N3886);
and AND3 (N6094, N6055, N996, N1583);
not NOT1 (N6095, N6074);
buf BUF1 (N6096, N6093);
not NOT1 (N6097, N6070);
nand NAND4 (N6098, N6095, N2954, N1117, N4300);
nor NOR3 (N6099, N6098, N3265, N1475);
and AND3 (N6100, N6096, N1302, N5290);
nand NAND3 (N6101, N6091, N4943, N2126);
or OR4 (N6102, N6092, N114, N4840, N1140);
or OR4 (N6103, N6097, N1961, N2395, N68);
nor NOR4 (N6104, N6090, N716, N5150, N1222);
buf BUF1 (N6105, N6083);
or OR3 (N6106, N6094, N4256, N6004);
xor XOR2 (N6107, N6100, N5917);
and AND3 (N6108, N6089, N1026, N261);
and AND3 (N6109, N6086, N2379, N2866);
buf BUF1 (N6110, N6103);
buf BUF1 (N6111, N6101);
and AND2 (N6112, N6107, N1035);
not NOT1 (N6113, N6110);
or OR4 (N6114, N6112, N5119, N5408, N2041);
nor NOR4 (N6115, N6099, N1971, N5406, N2618);
buf BUF1 (N6116, N6108);
and AND3 (N6117, N6116, N1849, N5663);
buf BUF1 (N6118, N6115);
or OR2 (N6119, N6105, N5112);
or OR2 (N6120, N6119, N5319);
xor XOR2 (N6121, N6120, N2969);
xor XOR2 (N6122, N6102, N1286);
and AND4 (N6123, N6113, N4316, N2011, N333);
not NOT1 (N6124, N6121);
not NOT1 (N6125, N6106);
nor NOR3 (N6126, N6125, N802, N4286);
not NOT1 (N6127, N6117);
nand NAND4 (N6128, N6122, N2996, N5459, N485);
not NOT1 (N6129, N6128);
or OR4 (N6130, N6129, N2727, N5284, N5768);
or OR4 (N6131, N6104, N1060, N1768, N1287);
and AND4 (N6132, N6118, N3371, N2917, N5921);
not NOT1 (N6133, N6127);
and AND2 (N6134, N6133, N2096);
or OR2 (N6135, N6134, N3198);
xor XOR2 (N6136, N6130, N5928);
or OR4 (N6137, N6111, N3113, N4432, N5108);
nand NAND3 (N6138, N6136, N3699, N2417);
nand NAND4 (N6139, N6132, N1301, N5573, N3764);
not NOT1 (N6140, N6109);
or OR2 (N6141, N6140, N5990);
buf BUF1 (N6142, N6141);
buf BUF1 (N6143, N6131);
nand NAND4 (N6144, N6137, N2063, N3535, N2309);
or OR2 (N6145, N6138, N5004);
and AND2 (N6146, N6123, N2399);
and AND2 (N6147, N6126, N5817);
buf BUF1 (N6148, N6145);
nor NOR4 (N6149, N6143, N3718, N488, N2449);
buf BUF1 (N6150, N6142);
nor NOR4 (N6151, N6147, N5476, N2699, N1655);
nand NAND2 (N6152, N6151, N1240);
xor XOR2 (N6153, N6150, N4910);
not NOT1 (N6154, N6135);
buf BUF1 (N6155, N6139);
and AND3 (N6156, N6148, N3431, N2688);
and AND3 (N6157, N6153, N882, N959);
buf BUF1 (N6158, N6124);
nor NOR3 (N6159, N6149, N4293, N3185);
not NOT1 (N6160, N6114);
or OR3 (N6161, N6159, N77, N5285);
not NOT1 (N6162, N6146);
or OR4 (N6163, N6144, N5581, N1309, N1708);
nor NOR3 (N6164, N6157, N1640, N5890);
buf BUF1 (N6165, N6152);
or OR2 (N6166, N6158, N1976);
buf BUF1 (N6167, N6165);
nand NAND2 (N6168, N6164, N1704);
nand NAND4 (N6169, N6154, N625, N1779, N6092);
buf BUF1 (N6170, N6160);
xor XOR2 (N6171, N6166, N3517);
not NOT1 (N6172, N6171);
buf BUF1 (N6173, N6161);
and AND2 (N6174, N6155, N4530);
nand NAND2 (N6175, N6162, N4438);
buf BUF1 (N6176, N6175);
not NOT1 (N6177, N6156);
and AND2 (N6178, N6172, N813);
or OR2 (N6179, N6170, N158);
not NOT1 (N6180, N6177);
nor NOR4 (N6181, N6174, N4946, N2136, N2911);
xor XOR2 (N6182, N6176, N2312);
not NOT1 (N6183, N6169);
buf BUF1 (N6184, N6180);
and AND2 (N6185, N6181, N53);
nor NOR3 (N6186, N6184, N2027, N1886);
buf BUF1 (N6187, N6186);
and AND4 (N6188, N6173, N4561, N977, N1002);
nand NAND3 (N6189, N6167, N907, N3277);
not NOT1 (N6190, N6168);
xor XOR2 (N6191, N6183, N267);
and AND2 (N6192, N6191, N4729);
nand NAND3 (N6193, N6178, N4337, N875);
and AND2 (N6194, N6179, N4752);
nand NAND2 (N6195, N6163, N4729);
nand NAND3 (N6196, N6182, N6058, N4999);
not NOT1 (N6197, N6196);
buf BUF1 (N6198, N6188);
and AND2 (N6199, N6193, N2734);
nand NAND4 (N6200, N6192, N160, N893, N473);
nor NOR2 (N6201, N6195, N887);
buf BUF1 (N6202, N6189);
and AND4 (N6203, N6200, N4679, N5231, N6028);
nand NAND3 (N6204, N6187, N6195, N2389);
nand NAND4 (N6205, N6185, N3447, N1643, N1417);
nor NOR4 (N6206, N6204, N2208, N2648, N668);
xor XOR2 (N6207, N6201, N5714);
nand NAND2 (N6208, N6206, N1256);
nand NAND3 (N6209, N6202, N801, N1411);
and AND3 (N6210, N6194, N4053, N2280);
buf BUF1 (N6211, N6205);
not NOT1 (N6212, N6203);
buf BUF1 (N6213, N6197);
nand NAND3 (N6214, N6190, N5383, N3617);
not NOT1 (N6215, N6209);
and AND4 (N6216, N6198, N4189, N2361, N3629);
and AND3 (N6217, N6207, N5651, N3222);
not NOT1 (N6218, N6216);
nor NOR4 (N6219, N6211, N6069, N266, N4630);
xor XOR2 (N6220, N6213, N2890);
and AND2 (N6221, N6208, N224);
and AND3 (N6222, N6221, N3388, N802);
xor XOR2 (N6223, N6217, N5716);
buf BUF1 (N6224, N6214);
and AND3 (N6225, N6220, N2801, N374);
and AND2 (N6226, N6210, N5752);
xor XOR2 (N6227, N6226, N6158);
or OR4 (N6228, N6224, N162, N656, N5104);
not NOT1 (N6229, N6199);
or OR3 (N6230, N6212, N4411, N5172);
not NOT1 (N6231, N6215);
or OR4 (N6232, N6230, N5225, N4127, N5259);
or OR2 (N6233, N6223, N5004);
and AND3 (N6234, N6218, N1078, N4484);
not NOT1 (N6235, N6234);
nor NOR2 (N6236, N6232, N1206);
xor XOR2 (N6237, N6225, N426);
or OR4 (N6238, N6235, N4369, N2655, N1433);
nand NAND3 (N6239, N6222, N1865, N5652);
not NOT1 (N6240, N6237);
and AND4 (N6241, N6227, N3581, N1613, N2501);
xor XOR2 (N6242, N6240, N4093);
nand NAND4 (N6243, N6242, N960, N5931, N4891);
and AND4 (N6244, N6229, N4202, N2725, N562);
nor NOR3 (N6245, N6231, N4600, N310);
buf BUF1 (N6246, N6239);
nand NAND2 (N6247, N6236, N1563);
not NOT1 (N6248, N6245);
or OR3 (N6249, N6228, N356, N635);
nor NOR3 (N6250, N6248, N1114, N1448);
not NOT1 (N6251, N6238);
buf BUF1 (N6252, N6246);
xor XOR2 (N6253, N6233, N4965);
nand NAND3 (N6254, N6252, N6025, N4453);
not NOT1 (N6255, N6244);
and AND2 (N6256, N6251, N803);
or OR4 (N6257, N6255, N3068, N5968, N1718);
or OR3 (N6258, N6257, N5520, N3996);
and AND4 (N6259, N6219, N4374, N1603, N5526);
or OR4 (N6260, N6250, N948, N5442, N6160);
not NOT1 (N6261, N6254);
buf BUF1 (N6262, N6260);
and AND3 (N6263, N6253, N4363, N278);
buf BUF1 (N6264, N6258);
nor NOR2 (N6265, N6262, N264);
nor NOR3 (N6266, N6259, N4821, N4495);
buf BUF1 (N6267, N6263);
buf BUF1 (N6268, N6267);
buf BUF1 (N6269, N6243);
not NOT1 (N6270, N6265);
buf BUF1 (N6271, N6268);
nor NOR2 (N6272, N6261, N2753);
or OR4 (N6273, N6264, N3723, N3865, N5507);
xor XOR2 (N6274, N6249, N3460);
buf BUF1 (N6275, N6256);
nand NAND3 (N6276, N6241, N1128, N3040);
nand NAND4 (N6277, N6270, N5027, N2121, N4698);
xor XOR2 (N6278, N6269, N2558);
or OR2 (N6279, N6278, N6142);
or OR4 (N6280, N6275, N407, N3604, N5206);
nor NOR4 (N6281, N6273, N2484, N5039, N1028);
not NOT1 (N6282, N6279);
buf BUF1 (N6283, N6272);
or OR4 (N6284, N6274, N3647, N2138, N3924);
xor XOR2 (N6285, N6276, N1211);
not NOT1 (N6286, N6285);
xor XOR2 (N6287, N6283, N2948);
or OR3 (N6288, N6277, N4369, N3148);
xor XOR2 (N6289, N6288, N6083);
nand NAND2 (N6290, N6280, N920);
nand NAND4 (N6291, N6247, N2391, N346, N5370);
nor NOR2 (N6292, N6266, N3715);
buf BUF1 (N6293, N6281);
nor NOR4 (N6294, N6286, N1248, N3166, N2693);
not NOT1 (N6295, N6271);
xor XOR2 (N6296, N6293, N1578);
not NOT1 (N6297, N6282);
xor XOR2 (N6298, N6291, N1599);
and AND3 (N6299, N6290, N2968, N3129);
or OR4 (N6300, N6292, N3569, N904, N5520);
or OR4 (N6301, N6284, N2063, N3877, N901);
xor XOR2 (N6302, N6299, N6154);
xor XOR2 (N6303, N6287, N1386);
nand NAND2 (N6304, N6300, N807);
and AND2 (N6305, N6289, N4341);
xor XOR2 (N6306, N6305, N5156);
xor XOR2 (N6307, N6306, N3653);
xor XOR2 (N6308, N6302, N6015);
xor XOR2 (N6309, N6296, N6258);
nand NAND4 (N6310, N6301, N3792, N2136, N2648);
and AND3 (N6311, N6298, N4294, N6131);
not NOT1 (N6312, N6295);
not NOT1 (N6313, N6304);
and AND3 (N6314, N6312, N4686, N5194);
not NOT1 (N6315, N6309);
xor XOR2 (N6316, N6308, N3329);
xor XOR2 (N6317, N6311, N5097);
nand NAND4 (N6318, N6316, N796, N5843, N2728);
not NOT1 (N6319, N6307);
xor XOR2 (N6320, N6313, N4213);
buf BUF1 (N6321, N6297);
xor XOR2 (N6322, N6310, N1457);
and AND2 (N6323, N6320, N2592);
buf BUF1 (N6324, N6318);
or OR4 (N6325, N6317, N4991, N315, N1985);
or OR4 (N6326, N6303, N2382, N290, N5241);
and AND4 (N6327, N6319, N342, N3065, N5663);
or OR2 (N6328, N6314, N2067);
buf BUF1 (N6329, N6294);
and AND2 (N6330, N6323, N2529);
buf BUF1 (N6331, N6328);
nor NOR2 (N6332, N6326, N84);
and AND2 (N6333, N6331, N6146);
xor XOR2 (N6334, N6330, N365);
or OR3 (N6335, N6329, N3026, N2236);
nor NOR3 (N6336, N6324, N5758, N5117);
xor XOR2 (N6337, N6336, N3027);
or OR4 (N6338, N6315, N6137, N631, N2020);
or OR4 (N6339, N6337, N5661, N2423, N1051);
not NOT1 (N6340, N6332);
nand NAND4 (N6341, N6335, N6098, N4933, N1429);
buf BUF1 (N6342, N6325);
nand NAND2 (N6343, N6322, N5753);
nand NAND2 (N6344, N6339, N486);
or OR4 (N6345, N6333, N1143, N3668, N40);
nand NAND3 (N6346, N6341, N774, N3238);
nor NOR4 (N6347, N6343, N4373, N622, N2305);
and AND3 (N6348, N6346, N4310, N3338);
nand NAND4 (N6349, N6344, N4158, N1708, N4158);
nand NAND4 (N6350, N6348, N6065, N1948, N613);
not NOT1 (N6351, N6347);
buf BUF1 (N6352, N6321);
or OR2 (N6353, N6342, N6078);
not NOT1 (N6354, N6345);
buf BUF1 (N6355, N6340);
not NOT1 (N6356, N6355);
xor XOR2 (N6357, N6356, N2300);
nand NAND4 (N6358, N6352, N4616, N54, N668);
and AND4 (N6359, N6350, N576, N1540, N5148);
or OR2 (N6360, N6358, N1090);
not NOT1 (N6361, N6354);
xor XOR2 (N6362, N6353, N5694);
and AND2 (N6363, N6359, N5577);
not NOT1 (N6364, N6351);
or OR2 (N6365, N6349, N4901);
and AND3 (N6366, N6361, N5460, N4830);
not NOT1 (N6367, N6363);
xor XOR2 (N6368, N6362, N2631);
or OR2 (N6369, N6357, N310);
and AND2 (N6370, N6338, N4570);
and AND3 (N6371, N6368, N4553, N766);
nor NOR2 (N6372, N6327, N5996);
nand NAND2 (N6373, N6371, N508);
not NOT1 (N6374, N6360);
xor XOR2 (N6375, N6365, N3698);
and AND3 (N6376, N6364, N6358, N6117);
not NOT1 (N6377, N6372);
buf BUF1 (N6378, N6376);
not NOT1 (N6379, N6370);
nor NOR2 (N6380, N6373, N2776);
nor NOR2 (N6381, N6375, N1684);
buf BUF1 (N6382, N6367);
buf BUF1 (N6383, N6380);
not NOT1 (N6384, N6382);
or OR4 (N6385, N6379, N1354, N2442, N2266);
nor NOR4 (N6386, N6381, N235, N3935, N3649);
buf BUF1 (N6387, N6374);
buf BUF1 (N6388, N6386);
buf BUF1 (N6389, N6388);
buf BUF1 (N6390, N6334);
xor XOR2 (N6391, N6390, N3723);
xor XOR2 (N6392, N6391, N6008);
or OR4 (N6393, N6366, N5825, N388, N1725);
not NOT1 (N6394, N6384);
not NOT1 (N6395, N6377);
nand NAND2 (N6396, N6369, N6276);
xor XOR2 (N6397, N6395, N6053);
nor NOR2 (N6398, N6387, N859);
xor XOR2 (N6399, N6383, N2620);
nor NOR4 (N6400, N6392, N4286, N1756, N5165);
xor XOR2 (N6401, N6398, N5059);
not NOT1 (N6402, N6378);
buf BUF1 (N6403, N6397);
and AND4 (N6404, N6399, N3468, N2206, N1435);
xor XOR2 (N6405, N6401, N2078);
buf BUF1 (N6406, N6403);
not NOT1 (N6407, N6393);
and AND4 (N6408, N6404, N6166, N1154, N4358);
not NOT1 (N6409, N6396);
nor NOR2 (N6410, N6409, N3846);
nor NOR2 (N6411, N6402, N5909);
nand NAND4 (N6412, N6410, N3382, N5951, N4189);
or OR3 (N6413, N6400, N2959, N5834);
buf BUF1 (N6414, N6406);
xor XOR2 (N6415, N6389, N6143);
xor XOR2 (N6416, N6405, N6341);
or OR2 (N6417, N6394, N1496);
not NOT1 (N6418, N6414);
nor NOR3 (N6419, N6416, N3915, N5582);
nor NOR3 (N6420, N6385, N5225, N6287);
buf BUF1 (N6421, N6413);
nor NOR4 (N6422, N6421, N162, N5201, N2823);
xor XOR2 (N6423, N6420, N6316);
nor NOR4 (N6424, N6407, N5618, N1229, N3805);
not NOT1 (N6425, N6418);
or OR3 (N6426, N6425, N5438, N2632);
and AND2 (N6427, N6422, N3392);
or OR4 (N6428, N6424, N2608, N3005, N4977);
nor NOR3 (N6429, N6411, N4598, N1226);
and AND4 (N6430, N6408, N4266, N4421, N754);
nor NOR4 (N6431, N6423, N4331, N3832, N6398);
not NOT1 (N6432, N6427);
xor XOR2 (N6433, N6431, N4301);
nand NAND2 (N6434, N6432, N4207);
buf BUF1 (N6435, N6415);
nor NOR2 (N6436, N6426, N5185);
and AND4 (N6437, N6435, N5135, N3070, N5952);
buf BUF1 (N6438, N6434);
xor XOR2 (N6439, N6437, N2213);
or OR3 (N6440, N6428, N4248, N4314);
not NOT1 (N6441, N6419);
not NOT1 (N6442, N6436);
and AND2 (N6443, N6429, N4574);
nor NOR3 (N6444, N6440, N4715, N4984);
xor XOR2 (N6445, N6444, N5024);
nand NAND4 (N6446, N6417, N2546, N6032, N6146);
nand NAND4 (N6447, N6439, N6054, N4599, N5874);
nor NOR3 (N6448, N6445, N4520, N754);
nor NOR3 (N6449, N6448, N4703, N5260);
not NOT1 (N6450, N6449);
nand NAND4 (N6451, N6442, N1575, N2787, N4296);
and AND2 (N6452, N6438, N4868);
nor NOR2 (N6453, N6433, N3379);
not NOT1 (N6454, N6443);
not NOT1 (N6455, N6447);
buf BUF1 (N6456, N6455);
or OR3 (N6457, N6446, N3677, N790);
or OR3 (N6458, N6457, N2368, N326);
xor XOR2 (N6459, N6456, N4689);
or OR3 (N6460, N6453, N3359, N1198);
nor NOR4 (N6461, N6452, N4778, N3149, N574);
not NOT1 (N6462, N6458);
nand NAND2 (N6463, N6451, N4993);
xor XOR2 (N6464, N6460, N3406);
nand NAND3 (N6465, N6462, N6254, N2837);
nor NOR2 (N6466, N6450, N2154);
xor XOR2 (N6467, N6412, N895);
nand NAND3 (N6468, N6461, N5852, N2850);
xor XOR2 (N6469, N6465, N3808);
not NOT1 (N6470, N6466);
not NOT1 (N6471, N6470);
or OR3 (N6472, N6430, N1365, N2778);
nor NOR3 (N6473, N6441, N3486, N6162);
nor NOR4 (N6474, N6473, N1402, N5518, N5940);
nor NOR4 (N6475, N6467, N4324, N1521, N4150);
nor NOR4 (N6476, N6468, N5816, N3219, N677);
or OR3 (N6477, N6474, N3838, N6418);
nand NAND2 (N6478, N6476, N257);
nand NAND4 (N6479, N6471, N575, N2770, N4682);
nand NAND4 (N6480, N6464, N4569, N4082, N245);
buf BUF1 (N6481, N6469);
and AND4 (N6482, N6477, N3532, N4218, N106);
nand NAND3 (N6483, N6454, N1679, N1764);
nand NAND4 (N6484, N6480, N952, N2804, N983);
not NOT1 (N6485, N6472);
and AND2 (N6486, N6459, N818);
not NOT1 (N6487, N6483);
nor NOR4 (N6488, N6478, N491, N3094, N2754);
nor NOR3 (N6489, N6475, N1171, N4359);
nand NAND4 (N6490, N6482, N4650, N3799, N1128);
or OR2 (N6491, N6463, N4076);
or OR4 (N6492, N6489, N414, N6155, N1276);
and AND3 (N6493, N6488, N719, N5234);
nand NAND3 (N6494, N6486, N617, N6055);
or OR4 (N6495, N6487, N1573, N4150, N2818);
buf BUF1 (N6496, N6479);
not NOT1 (N6497, N6493);
nand NAND3 (N6498, N6481, N5074, N6422);
or OR3 (N6499, N6492, N4221, N4121);
xor XOR2 (N6500, N6485, N30);
not NOT1 (N6501, N6484);
not NOT1 (N6502, N6497);
xor XOR2 (N6503, N6494, N2976);
not NOT1 (N6504, N6502);
and AND2 (N6505, N6499, N6358);
or OR4 (N6506, N6504, N6091, N2024, N1763);
or OR3 (N6507, N6496, N569, N4561);
and AND3 (N6508, N6500, N5976, N4406);
buf BUF1 (N6509, N6501);
xor XOR2 (N6510, N6508, N5178);
not NOT1 (N6511, N6491);
and AND3 (N6512, N6490, N1061, N810);
or OR4 (N6513, N6509, N4426, N2207, N4035);
or OR2 (N6514, N6510, N5776);
xor XOR2 (N6515, N6505, N820);
and AND2 (N6516, N6512, N3807);
buf BUF1 (N6517, N6507);
or OR2 (N6518, N6516, N2446);
buf BUF1 (N6519, N6517);
nand NAND3 (N6520, N6515, N5019, N1967);
xor XOR2 (N6521, N6506, N4730);
or OR2 (N6522, N6520, N5971);
nor NOR3 (N6523, N6498, N2584, N6355);
nand NAND2 (N6524, N6495, N6021);
not NOT1 (N6525, N6522);
nor NOR4 (N6526, N6513, N109, N5567, N333);
nor NOR4 (N6527, N6521, N4410, N6181, N648);
not NOT1 (N6528, N6527);
and AND3 (N6529, N6514, N1864, N4352);
nor NOR4 (N6530, N6524, N2047, N6089, N3028);
and AND3 (N6531, N6528, N4310, N3272);
or OR4 (N6532, N6531, N1557, N5774, N2210);
nand NAND3 (N6533, N6523, N3425, N763);
nand NAND2 (N6534, N6529, N1568);
and AND2 (N6535, N6533, N4286);
buf BUF1 (N6536, N6511);
not NOT1 (N6537, N6503);
not NOT1 (N6538, N6536);
and AND2 (N6539, N6538, N558);
and AND4 (N6540, N6518, N4714, N529, N6357);
buf BUF1 (N6541, N6526);
nor NOR4 (N6542, N6532, N6537, N4695, N1657);
and AND2 (N6543, N2770, N3068);
nor NOR3 (N6544, N6540, N6205, N412);
or OR2 (N6545, N6539, N1005);
xor XOR2 (N6546, N6530, N5917);
and AND2 (N6547, N6545, N4787);
xor XOR2 (N6548, N6535, N2962);
nor NOR3 (N6549, N6547, N1653, N4525);
nor NOR4 (N6550, N6541, N3532, N96, N4494);
buf BUF1 (N6551, N6534);
nor NOR2 (N6552, N6544, N4965);
xor XOR2 (N6553, N6551, N4146);
not NOT1 (N6554, N6525);
or OR4 (N6555, N6550, N2020, N6440, N4834);
nand NAND2 (N6556, N6543, N4706);
buf BUF1 (N6557, N6555);
nor NOR4 (N6558, N6556, N2988, N3211, N3227);
buf BUF1 (N6559, N6542);
xor XOR2 (N6560, N6559, N461);
not NOT1 (N6561, N6560);
buf BUF1 (N6562, N6554);
nand NAND3 (N6563, N6548, N4243, N1975);
nand NAND2 (N6564, N6549, N3924);
or OR2 (N6565, N6546, N2070);
xor XOR2 (N6566, N6558, N5361);
buf BUF1 (N6567, N6565);
and AND2 (N6568, N6563, N2578);
nand NAND4 (N6569, N6519, N4015, N6432, N4944);
and AND4 (N6570, N6567, N4080, N4925, N6103);
buf BUF1 (N6571, N6570);
and AND2 (N6572, N6571, N165);
or OR4 (N6573, N6552, N2341, N574, N6145);
nand NAND2 (N6574, N6572, N3938);
or OR4 (N6575, N6566, N1912, N4942, N2495);
or OR4 (N6576, N6569, N5897, N3211, N3262);
and AND3 (N6577, N6557, N5428, N5465);
xor XOR2 (N6578, N6564, N4143);
or OR4 (N6579, N6575, N1696, N1276, N4802);
or OR2 (N6580, N6573, N2063);
nor NOR4 (N6581, N6574, N794, N5668, N2349);
buf BUF1 (N6582, N6562);
not NOT1 (N6583, N6579);
xor XOR2 (N6584, N6583, N2502);
and AND3 (N6585, N6553, N2164, N3811);
xor XOR2 (N6586, N6576, N6095);
xor XOR2 (N6587, N6584, N2552);
buf BUF1 (N6588, N6561);
and AND2 (N6589, N6578, N6277);
buf BUF1 (N6590, N6585);
nand NAND3 (N6591, N6590, N4357, N1770);
xor XOR2 (N6592, N6591, N3363);
nand NAND4 (N6593, N6582, N1940, N5635, N145);
nor NOR3 (N6594, N6587, N1513, N1440);
xor XOR2 (N6595, N6581, N3240);
nand NAND4 (N6596, N6588, N407, N4149, N1643);
xor XOR2 (N6597, N6595, N6444);
nand NAND4 (N6598, N6596, N281, N5652, N3750);
nand NAND3 (N6599, N6577, N6507, N1309);
buf BUF1 (N6600, N6580);
nand NAND3 (N6601, N6568, N814, N6181);
xor XOR2 (N6602, N6586, N2746);
buf BUF1 (N6603, N6599);
nor NOR3 (N6604, N6593, N4321, N3836);
buf BUF1 (N6605, N6600);
nor NOR3 (N6606, N6605, N2210, N2407);
not NOT1 (N6607, N6601);
not NOT1 (N6608, N6592);
nor NOR4 (N6609, N6594, N2712, N1267, N2065);
and AND2 (N6610, N6604, N639);
nand NAND3 (N6611, N6603, N204, N5765);
or OR3 (N6612, N6608, N556, N1595);
nand NAND3 (N6613, N6602, N5160, N3629);
xor XOR2 (N6614, N6607, N1878);
or OR2 (N6615, N6597, N4624);
nand NAND2 (N6616, N6609, N4411);
xor XOR2 (N6617, N6612, N2759);
or OR3 (N6618, N6614, N4779, N979);
buf BUF1 (N6619, N6616);
nor NOR2 (N6620, N6617, N2469);
xor XOR2 (N6621, N6610, N5074);
not NOT1 (N6622, N6606);
or OR4 (N6623, N6618, N2281, N2551, N6126);
and AND4 (N6624, N6621, N6246, N614, N2189);
buf BUF1 (N6625, N6611);
nor NOR2 (N6626, N6615, N198);
and AND3 (N6627, N6613, N3672, N5122);
xor XOR2 (N6628, N6627, N3571);
or OR3 (N6629, N6619, N5655, N1239);
or OR3 (N6630, N6628, N3863, N5475);
or OR2 (N6631, N6598, N5658);
nor NOR2 (N6632, N6624, N4007);
xor XOR2 (N6633, N6620, N6527);
nor NOR4 (N6634, N6632, N3378, N4937, N2530);
not NOT1 (N6635, N6589);
or OR2 (N6636, N6631, N1209);
or OR3 (N6637, N6630, N2958, N5698);
not NOT1 (N6638, N6625);
nor NOR2 (N6639, N6634, N139);
buf BUF1 (N6640, N6636);
nand NAND4 (N6641, N6635, N360, N3591, N5185);
nand NAND2 (N6642, N6623, N5762);
and AND2 (N6643, N6639, N6256);
xor XOR2 (N6644, N6641, N1945);
or OR2 (N6645, N6640, N837);
nor NOR3 (N6646, N6645, N576, N4892);
and AND3 (N6647, N6642, N2130, N1134);
and AND4 (N6648, N6637, N389, N4134, N5076);
nand NAND4 (N6649, N6629, N5648, N5507, N241);
and AND2 (N6650, N6649, N375);
not NOT1 (N6651, N6626);
xor XOR2 (N6652, N6633, N2529);
or OR4 (N6653, N6622, N5931, N1388, N2049);
nand NAND4 (N6654, N6652, N2726, N3101, N4045);
or OR3 (N6655, N6654, N754, N4547);
and AND2 (N6656, N6647, N813);
nand NAND3 (N6657, N6653, N2183, N5800);
nand NAND2 (N6658, N6650, N3344);
and AND2 (N6659, N6648, N5698);
nand NAND3 (N6660, N6659, N1363, N5828);
nand NAND4 (N6661, N6638, N2201, N1380, N6150);
nor NOR4 (N6662, N6644, N2975, N434, N1543);
xor XOR2 (N6663, N6660, N2820);
nand NAND4 (N6664, N6661, N4288, N5420, N327);
xor XOR2 (N6665, N6651, N4441);
nand NAND2 (N6666, N6663, N1202);
or OR3 (N6667, N6666, N1820, N6434);
nand NAND4 (N6668, N6665, N5964, N3273, N5246);
or OR2 (N6669, N6667, N1380);
and AND4 (N6670, N6668, N3362, N5818, N4487);
or OR2 (N6671, N6655, N3695);
not NOT1 (N6672, N6657);
xor XOR2 (N6673, N6664, N2899);
buf BUF1 (N6674, N6669);
nand NAND4 (N6675, N6674, N6068, N3788, N1655);
xor XOR2 (N6676, N6670, N3586);
buf BUF1 (N6677, N6676);
not NOT1 (N6678, N6646);
or OR3 (N6679, N6656, N1249, N6352);
nand NAND2 (N6680, N6675, N881);
nand NAND4 (N6681, N6680, N328, N771, N6351);
or OR4 (N6682, N6643, N465, N4645, N5494);
or OR3 (N6683, N6658, N3987, N2872);
not NOT1 (N6684, N6683);
xor XOR2 (N6685, N6678, N1653);
xor XOR2 (N6686, N6682, N5099);
xor XOR2 (N6687, N6686, N4994);
not NOT1 (N6688, N6662);
xor XOR2 (N6689, N6688, N2318);
buf BUF1 (N6690, N6677);
buf BUF1 (N6691, N6673);
not NOT1 (N6692, N6672);
xor XOR2 (N6693, N6692, N87);
nand NAND3 (N6694, N6691, N2533, N6560);
nor NOR4 (N6695, N6681, N2822, N3508, N2465);
and AND4 (N6696, N6689, N3653, N4405, N670);
not NOT1 (N6697, N6685);
xor XOR2 (N6698, N6690, N6675);
nor NOR4 (N6699, N6684, N2528, N3901, N333);
xor XOR2 (N6700, N6695, N2491);
and AND4 (N6701, N6694, N4496, N1484, N2831);
nor NOR3 (N6702, N6698, N2935, N1620);
buf BUF1 (N6703, N6701);
xor XOR2 (N6704, N6693, N336);
buf BUF1 (N6705, N6697);
buf BUF1 (N6706, N6696);
xor XOR2 (N6707, N6706, N4050);
nor NOR3 (N6708, N6679, N825, N4712);
buf BUF1 (N6709, N6703);
xor XOR2 (N6710, N6699, N4169);
nand NAND2 (N6711, N6705, N2968);
nor NOR3 (N6712, N6687, N26, N4574);
or OR4 (N6713, N6707, N3895, N1779, N6128);
nand NAND2 (N6714, N6702, N726);
xor XOR2 (N6715, N6712, N5506);
and AND2 (N6716, N6710, N6259);
nand NAND3 (N6717, N6713, N3038, N2670);
nand NAND2 (N6718, N6709, N3305);
buf BUF1 (N6719, N6700);
not NOT1 (N6720, N6719);
nand NAND3 (N6721, N6708, N3681, N4954);
nor NOR4 (N6722, N6671, N2819, N5461, N2423);
buf BUF1 (N6723, N6722);
not NOT1 (N6724, N6721);
nand NAND4 (N6725, N6717, N3581, N3489, N2373);
nor NOR3 (N6726, N6716, N3952, N5724);
or OR3 (N6727, N6714, N2397, N3816);
nor NOR4 (N6728, N6724, N5866, N3519, N2363);
nand NAND2 (N6729, N6727, N2492);
xor XOR2 (N6730, N6729, N1059);
and AND2 (N6731, N6718, N3018);
not NOT1 (N6732, N6725);
buf BUF1 (N6733, N6723);
or OR3 (N6734, N6704, N330, N400);
nand NAND3 (N6735, N6734, N3006, N1915);
not NOT1 (N6736, N6715);
or OR2 (N6737, N6711, N4198);
buf BUF1 (N6738, N6737);
nand NAND4 (N6739, N6731, N3469, N4711, N3641);
not NOT1 (N6740, N6730);
not NOT1 (N6741, N6740);
nor NOR2 (N6742, N6733, N519);
and AND3 (N6743, N6741, N3208, N1764);
and AND4 (N6744, N6728, N4576, N3579, N2131);
nand NAND3 (N6745, N6726, N3768, N5678);
nor NOR4 (N6746, N6738, N426, N5282, N1001);
or OR4 (N6747, N6735, N3868, N4488, N6191);
or OR2 (N6748, N6746, N1688);
xor XOR2 (N6749, N6743, N3187);
nor NOR4 (N6750, N6749, N4603, N3152, N3190);
xor XOR2 (N6751, N6744, N458);
xor XOR2 (N6752, N6750, N3507);
nand NAND2 (N6753, N6739, N1813);
nor NOR4 (N6754, N6752, N2062, N6230, N3013);
not NOT1 (N6755, N6736);
xor XOR2 (N6756, N6720, N2048);
xor XOR2 (N6757, N6753, N5962);
buf BUF1 (N6758, N6747);
nor NOR2 (N6759, N6732, N2065);
not NOT1 (N6760, N6756);
buf BUF1 (N6761, N6754);
nor NOR2 (N6762, N6759, N3293);
buf BUF1 (N6763, N6742);
buf BUF1 (N6764, N6758);
and AND2 (N6765, N6748, N2568);
nor NOR2 (N6766, N6765, N187);
or OR3 (N6767, N6757, N5708, N1591);
and AND4 (N6768, N6755, N764, N3868, N3011);
nor NOR2 (N6769, N6767, N6427);
not NOT1 (N6770, N6768);
nor NOR3 (N6771, N6770, N5091, N4832);
nand NAND3 (N6772, N6761, N4395, N3857);
and AND4 (N6773, N6760, N6437, N6481, N6746);
not NOT1 (N6774, N6762);
xor XOR2 (N6775, N6745, N955);
and AND2 (N6776, N6751, N6012);
nor NOR4 (N6777, N6764, N2868, N6406, N735);
or OR2 (N6778, N6777, N3709);
nor NOR4 (N6779, N6772, N5155, N5331, N5984);
nor NOR2 (N6780, N6778, N3642);
nor NOR3 (N6781, N6779, N4637, N6473);
or OR2 (N6782, N6773, N5261);
xor XOR2 (N6783, N6776, N1594);
or OR3 (N6784, N6782, N6158, N3069);
and AND2 (N6785, N6771, N6439);
nand NAND2 (N6786, N6781, N1781);
or OR3 (N6787, N6775, N2477, N2959);
nand NAND2 (N6788, N6787, N4432);
not NOT1 (N6789, N6780);
nand NAND2 (N6790, N6784, N6453);
nor NOR2 (N6791, N6769, N1107);
buf BUF1 (N6792, N6766);
or OR2 (N6793, N6785, N843);
buf BUF1 (N6794, N6793);
or OR2 (N6795, N6794, N5495);
or OR2 (N6796, N6786, N6230);
and AND2 (N6797, N6791, N6160);
or OR3 (N6798, N6790, N2906, N1708);
and AND2 (N6799, N6774, N5721);
not NOT1 (N6800, N6789);
not NOT1 (N6801, N6795);
xor XOR2 (N6802, N6792, N3403);
or OR2 (N6803, N6763, N6198);
not NOT1 (N6804, N6797);
not NOT1 (N6805, N6803);
and AND3 (N6806, N6804, N96, N542);
or OR3 (N6807, N6788, N3916, N400);
nor NOR3 (N6808, N6798, N809, N4482);
not NOT1 (N6809, N6808);
not NOT1 (N6810, N6805);
xor XOR2 (N6811, N6801, N6791);
not NOT1 (N6812, N6809);
not NOT1 (N6813, N6807);
not NOT1 (N6814, N6799);
buf BUF1 (N6815, N6814);
and AND4 (N6816, N6811, N3469, N4496, N4241);
or OR2 (N6817, N6802, N6510);
not NOT1 (N6818, N6815);
xor XOR2 (N6819, N6783, N3011);
xor XOR2 (N6820, N6806, N1866);
nor NOR2 (N6821, N6800, N2142);
buf BUF1 (N6822, N6796);
xor XOR2 (N6823, N6820, N6389);
and AND4 (N6824, N6818, N2283, N976, N137);
buf BUF1 (N6825, N6816);
or OR3 (N6826, N6823, N4178, N2082);
not NOT1 (N6827, N6821);
not NOT1 (N6828, N6824);
and AND3 (N6829, N6827, N606, N5830);
buf BUF1 (N6830, N6817);
not NOT1 (N6831, N6828);
or OR4 (N6832, N6829, N808, N2672, N530);
not NOT1 (N6833, N6812);
xor XOR2 (N6834, N6826, N3268);
or OR4 (N6835, N6831, N5519, N5592, N6469);
nand NAND3 (N6836, N6834, N2203, N3400);
not NOT1 (N6837, N6810);
or OR2 (N6838, N6832, N5387);
buf BUF1 (N6839, N6825);
and AND4 (N6840, N6819, N6808, N1839, N6604);
or OR4 (N6841, N6822, N6339, N3218, N5912);
and AND2 (N6842, N6839, N2983);
and AND4 (N6843, N6813, N2648, N4419, N4571);
nand NAND3 (N6844, N6841, N2890, N3190);
xor XOR2 (N6845, N6835, N3248);
not NOT1 (N6846, N6830);
nand NAND3 (N6847, N6845, N1284, N656);
xor XOR2 (N6848, N6837, N352);
or OR3 (N6849, N6833, N2355, N982);
not NOT1 (N6850, N6848);
nand NAND2 (N6851, N6842, N4778);
and AND3 (N6852, N6847, N4880, N5000);
xor XOR2 (N6853, N6851, N3913);
nor NOR2 (N6854, N6852, N4363);
nor NOR3 (N6855, N6844, N4822, N2664);
or OR2 (N6856, N6849, N2650);
or OR4 (N6857, N6850, N1619, N1254, N4266);
not NOT1 (N6858, N6855);
xor XOR2 (N6859, N6838, N2057);
not NOT1 (N6860, N6859);
and AND3 (N6861, N6843, N3318, N6578);
nor NOR2 (N6862, N6861, N2566);
nand NAND2 (N6863, N6858, N4891);
not NOT1 (N6864, N6836);
nand NAND4 (N6865, N6840, N2095, N5577, N140);
and AND4 (N6866, N6854, N4195, N3426, N813);
or OR4 (N6867, N6862, N1363, N5638, N4810);
nand NAND3 (N6868, N6856, N3526, N603);
xor XOR2 (N6869, N6857, N1067);
not NOT1 (N6870, N6860);
nor NOR4 (N6871, N6864, N3122, N5919, N840);
or OR3 (N6872, N6865, N6192, N5370);
xor XOR2 (N6873, N6853, N5966);
xor XOR2 (N6874, N6867, N5624);
and AND4 (N6875, N6869, N2657, N768, N213);
or OR4 (N6876, N6868, N4948, N141, N4393);
xor XOR2 (N6877, N6871, N969);
nor NOR2 (N6878, N6846, N4655);
xor XOR2 (N6879, N6876, N623);
or OR2 (N6880, N6875, N4756);
buf BUF1 (N6881, N6870);
or OR2 (N6882, N6881, N4594);
and AND4 (N6883, N6874, N3607, N1878, N6487);
xor XOR2 (N6884, N6880, N4110);
xor XOR2 (N6885, N6878, N2477);
nand NAND3 (N6886, N6863, N637, N2250);
nand NAND3 (N6887, N6882, N2090, N6809);
nor NOR4 (N6888, N6883, N4417, N1500, N3661);
xor XOR2 (N6889, N6885, N6313);
or OR3 (N6890, N6879, N6385, N831);
nand NAND2 (N6891, N6877, N3103);
nand NAND2 (N6892, N6888, N5823);
or OR4 (N6893, N6886, N5884, N1036, N3724);
nor NOR2 (N6894, N6891, N4369);
nand NAND3 (N6895, N6872, N5599, N4310);
xor XOR2 (N6896, N6890, N5954);
nand NAND2 (N6897, N6895, N2727);
and AND4 (N6898, N6889, N125, N3795, N3319);
buf BUF1 (N6899, N6898);
or OR4 (N6900, N6873, N2611, N2552, N5861);
nor NOR3 (N6901, N6884, N3320, N5675);
nor NOR2 (N6902, N6901, N3090);
not NOT1 (N6903, N6893);
and AND2 (N6904, N6899, N450);
buf BUF1 (N6905, N6897);
nor NOR2 (N6906, N6903, N3894);
nand NAND2 (N6907, N6904, N3293);
or OR4 (N6908, N6894, N1660, N2829, N36);
and AND2 (N6909, N6896, N1435);
not NOT1 (N6910, N6909);
not NOT1 (N6911, N6907);
xor XOR2 (N6912, N6905, N1205);
and AND2 (N6913, N6912, N940);
buf BUF1 (N6914, N6902);
or OR3 (N6915, N6892, N5159, N6511);
nor NOR3 (N6916, N6914, N6574, N1007);
nand NAND2 (N6917, N6908, N2491);
xor XOR2 (N6918, N6913, N5236);
and AND2 (N6919, N6906, N5920);
nor NOR4 (N6920, N6910, N3229, N5625, N393);
not NOT1 (N6921, N6917);
not NOT1 (N6922, N6915);
or OR4 (N6923, N6916, N3741, N3959, N3263);
nor NOR4 (N6924, N6922, N6468, N2507, N4690);
not NOT1 (N6925, N6921);
or OR2 (N6926, N6923, N4217);
nor NOR3 (N6927, N6911, N4058, N5534);
nand NAND2 (N6928, N6887, N4080);
and AND3 (N6929, N6866, N6467, N4568);
xor XOR2 (N6930, N6924, N2229);
nand NAND2 (N6931, N6929, N4465);
buf BUF1 (N6932, N6920);
and AND2 (N6933, N6932, N17);
xor XOR2 (N6934, N6928, N3701);
not NOT1 (N6935, N6918);
or OR2 (N6936, N6933, N6272);
xor XOR2 (N6937, N6926, N3001);
buf BUF1 (N6938, N6936);
and AND4 (N6939, N6930, N2470, N3651, N2971);
buf BUF1 (N6940, N6931);
xor XOR2 (N6941, N6940, N632);
not NOT1 (N6942, N6937);
nor NOR2 (N6943, N6935, N2243);
nor NOR3 (N6944, N6925, N3972, N6430);
or OR4 (N6945, N6900, N292, N1498, N4806);
nand NAND4 (N6946, N6942, N3902, N6883, N2414);
or OR3 (N6947, N6927, N4562, N4221);
nor NOR3 (N6948, N6938, N5649, N815);
not NOT1 (N6949, N6939);
nor NOR3 (N6950, N6944, N3792, N2071);
or OR3 (N6951, N6941, N3493, N3443);
xor XOR2 (N6952, N6946, N2795);
buf BUF1 (N6953, N6952);
nor NOR3 (N6954, N6953, N4120, N4503);
nor NOR4 (N6955, N6954, N902, N5008, N1182);
not NOT1 (N6956, N6951);
and AND2 (N6957, N6950, N3543);
buf BUF1 (N6958, N6945);
xor XOR2 (N6959, N6943, N98);
or OR4 (N6960, N6948, N4893, N1448, N1598);
nand NAND2 (N6961, N6958, N4194);
or OR2 (N6962, N6919, N2221);
nor NOR3 (N6963, N6934, N3249, N449);
xor XOR2 (N6964, N6957, N1849);
and AND2 (N6965, N6963, N2984);
or OR3 (N6966, N6961, N5025, N4602);
nand NAND3 (N6967, N6959, N1809, N5165);
xor XOR2 (N6968, N6947, N478);
or OR3 (N6969, N6964, N4955, N2857);
not NOT1 (N6970, N6965);
nor NOR2 (N6971, N6967, N1614);
and AND4 (N6972, N6968, N1723, N4399, N3941);
or OR3 (N6973, N6966, N6216, N5389);
nor NOR4 (N6974, N6970, N3552, N1743, N3965);
xor XOR2 (N6975, N6960, N4303);
or OR2 (N6976, N6971, N3717);
and AND3 (N6977, N6969, N4936, N4198);
or OR4 (N6978, N6974, N3108, N6641, N2718);
and AND2 (N6979, N6972, N13);
or OR2 (N6980, N6979, N1929);
or OR3 (N6981, N6973, N1675, N6901);
or OR2 (N6982, N6949, N5402);
buf BUF1 (N6983, N6962);
buf BUF1 (N6984, N6980);
buf BUF1 (N6985, N6975);
nor NOR4 (N6986, N6982, N3532, N917, N6280);
xor XOR2 (N6987, N6955, N809);
nor NOR4 (N6988, N6956, N3242, N3259, N6841);
xor XOR2 (N6989, N6988, N2276);
and AND2 (N6990, N6983, N4086);
nor NOR2 (N6991, N6987, N1658);
nand NAND4 (N6992, N6985, N6728, N3602, N3213);
or OR2 (N6993, N6990, N3171);
or OR4 (N6994, N6977, N6470, N4927, N542);
not NOT1 (N6995, N6991);
or OR4 (N6996, N6992, N6790, N708, N3330);
not NOT1 (N6997, N6978);
not NOT1 (N6998, N6981);
buf BUF1 (N6999, N6976);
or OR4 (N7000, N6986, N2044, N3724, N6680);
xor XOR2 (N7001, N6995, N4463);
buf BUF1 (N7002, N6994);
nor NOR3 (N7003, N6984, N66, N324);
xor XOR2 (N7004, N6993, N2074);
and AND4 (N7005, N7003, N6, N6902, N3078);
and AND4 (N7006, N7002, N853, N1798, N1637);
or OR4 (N7007, N7000, N6709, N4739, N2475);
or OR3 (N7008, N7001, N3843, N3162);
and AND2 (N7009, N6998, N1345);
xor XOR2 (N7010, N6996, N1240);
nor NOR3 (N7011, N7005, N5623, N1798);
nor NOR4 (N7012, N7004, N5327, N6702, N1298);
and AND4 (N7013, N7006, N5655, N557, N2013);
buf BUF1 (N7014, N6989);
buf BUF1 (N7015, N7012);
not NOT1 (N7016, N7013);
nand NAND3 (N7017, N7008, N5165, N1293);
nand NAND2 (N7018, N7014, N4132);
nor NOR3 (N7019, N7011, N114, N808);
xor XOR2 (N7020, N7009, N4870);
xor XOR2 (N7021, N7010, N1191);
xor XOR2 (N7022, N6997, N2356);
nor NOR4 (N7023, N7016, N2915, N3538, N4228);
xor XOR2 (N7024, N7021, N3197);
nand NAND3 (N7025, N7018, N1613, N5942);
nand NAND2 (N7026, N7020, N5605);
nand NAND3 (N7027, N7023, N6071, N909);
and AND2 (N7028, N7025, N786);
nor NOR2 (N7029, N7022, N556);
nor NOR4 (N7030, N7029, N5462, N6391, N2350);
or OR3 (N7031, N7017, N5025, N4018);
or OR4 (N7032, N7030, N2064, N4444, N6898);
or OR4 (N7033, N7019, N2036, N2017, N4157);
buf BUF1 (N7034, N7032);
and AND4 (N7035, N6999, N1008, N878, N919);
or OR3 (N7036, N7007, N1642, N4894);
not NOT1 (N7037, N7026);
not NOT1 (N7038, N7033);
xor XOR2 (N7039, N7035, N968);
or OR3 (N7040, N7037, N878, N6515);
or OR3 (N7041, N7031, N1445, N2795);
xor XOR2 (N7042, N7038, N3879);
nand NAND3 (N7043, N7042, N1865, N4196);
nand NAND4 (N7044, N7024, N4423, N6008, N5087);
buf BUF1 (N7045, N7043);
or OR3 (N7046, N7041, N434, N4111);
nor NOR3 (N7047, N7036, N5114, N1477);
xor XOR2 (N7048, N7028, N4988);
nor NOR4 (N7049, N7039, N4352, N6927, N1342);
nor NOR4 (N7050, N7046, N979, N5364, N4937);
nor NOR3 (N7051, N7044, N621, N1764);
xor XOR2 (N7052, N7040, N3241);
xor XOR2 (N7053, N7034, N5633);
and AND2 (N7054, N7048, N2237);
xor XOR2 (N7055, N7051, N1330);
nor NOR2 (N7056, N7054, N1818);
nor NOR3 (N7057, N7056, N6107, N1672);
and AND3 (N7058, N7052, N2732, N6575);
xor XOR2 (N7059, N7053, N1469);
not NOT1 (N7060, N7059);
xor XOR2 (N7061, N7050, N6484);
nor NOR2 (N7062, N7061, N4709);
buf BUF1 (N7063, N7015);
and AND3 (N7064, N7045, N6515, N175);
nor NOR3 (N7065, N7047, N4847, N6116);
buf BUF1 (N7066, N7063);
nand NAND4 (N7067, N7066, N493, N3195, N2397);
buf BUF1 (N7068, N7027);
buf BUF1 (N7069, N7049);
or OR4 (N7070, N7065, N2088, N4010, N278);
not NOT1 (N7071, N7068);
nor NOR4 (N7072, N7071, N5894, N2856, N4825);
and AND3 (N7073, N7069, N6266, N6275);
buf BUF1 (N7074, N7073);
buf BUF1 (N7075, N7055);
xor XOR2 (N7076, N7060, N2161);
or OR4 (N7077, N7062, N98, N6932, N6096);
nand NAND2 (N7078, N7075, N6586);
nor NOR3 (N7079, N7077, N3854, N3360);
and AND3 (N7080, N7072, N2642, N6877);
or OR3 (N7081, N7074, N5295, N2600);
and AND4 (N7082, N7057, N4996, N6133, N3085);
nand NAND2 (N7083, N7067, N2092);
buf BUF1 (N7084, N7076);
nor NOR3 (N7085, N7083, N4660, N6392);
not NOT1 (N7086, N7078);
buf BUF1 (N7087, N7070);
buf BUF1 (N7088, N7081);
and AND2 (N7089, N7082, N6403);
xor XOR2 (N7090, N7080, N1901);
or OR2 (N7091, N7064, N4356);
not NOT1 (N7092, N7090);
nor NOR3 (N7093, N7087, N637, N928);
and AND4 (N7094, N7088, N1988, N6430, N3001);
buf BUF1 (N7095, N7093);
buf BUF1 (N7096, N7084);
or OR4 (N7097, N7086, N4632, N3253, N3517);
not NOT1 (N7098, N7095);
and AND2 (N7099, N7058, N2408);
xor XOR2 (N7100, N7098, N5405);
nor NOR3 (N7101, N7096, N6611, N6569);
xor XOR2 (N7102, N7100, N4746);
not NOT1 (N7103, N7102);
nor NOR3 (N7104, N7079, N1604, N2146);
or OR3 (N7105, N7101, N62, N702);
not NOT1 (N7106, N7105);
or OR2 (N7107, N7092, N1289);
xor XOR2 (N7108, N7094, N3497);
buf BUF1 (N7109, N7107);
nor NOR2 (N7110, N7103, N3792);
not NOT1 (N7111, N7109);
not NOT1 (N7112, N7085);
nand NAND2 (N7113, N7104, N925);
and AND3 (N7114, N7091, N6076, N3266);
buf BUF1 (N7115, N7114);
xor XOR2 (N7116, N7112, N5431);
buf BUF1 (N7117, N7116);
and AND3 (N7118, N7108, N1110, N4189);
buf BUF1 (N7119, N7113);
and AND4 (N7120, N7106, N3356, N670, N1578);
not NOT1 (N7121, N7120);
and AND3 (N7122, N7117, N284, N1594);
not NOT1 (N7123, N7099);
nor NOR2 (N7124, N7110, N5509);
or OR2 (N7125, N7123, N6855);
nor NOR3 (N7126, N7121, N6340, N3893);
xor XOR2 (N7127, N7126, N7112);
xor XOR2 (N7128, N7097, N274);
and AND4 (N7129, N7115, N1740, N4062, N2886);
and AND4 (N7130, N7111, N1321, N6946, N690);
nand NAND3 (N7131, N7122, N4380, N3702);
nand NAND2 (N7132, N7125, N7010);
or OR4 (N7133, N7119, N823, N3879, N2070);
nor NOR2 (N7134, N7130, N3441);
buf BUF1 (N7135, N7132);
not NOT1 (N7136, N7133);
buf BUF1 (N7137, N7131);
nor NOR2 (N7138, N7127, N1689);
or OR3 (N7139, N7128, N3073, N958);
nor NOR2 (N7140, N7137, N6794);
xor XOR2 (N7141, N7138, N3762);
nor NOR3 (N7142, N7118, N333, N4143);
xor XOR2 (N7143, N7089, N3778);
or OR4 (N7144, N7142, N6290, N1474, N356);
not NOT1 (N7145, N7141);
or OR2 (N7146, N7144, N4672);
and AND3 (N7147, N7124, N7067, N1947);
or OR4 (N7148, N7134, N1797, N160, N6503);
buf BUF1 (N7149, N7143);
xor XOR2 (N7150, N7147, N5268);
not NOT1 (N7151, N7140);
and AND4 (N7152, N7148, N441, N6728, N5500);
nand NAND4 (N7153, N7145, N5469, N1031, N2963);
xor XOR2 (N7154, N7152, N3368);
buf BUF1 (N7155, N7154);
nand NAND4 (N7156, N7139, N6611, N3321, N7113);
nor NOR3 (N7157, N7129, N1039, N1376);
or OR4 (N7158, N7151, N2929, N1753, N2651);
xor XOR2 (N7159, N7156, N5302);
not NOT1 (N7160, N7153);
nand NAND2 (N7161, N7160, N2097);
buf BUF1 (N7162, N7161);
or OR3 (N7163, N7162, N2329, N1439);
not NOT1 (N7164, N7136);
nand NAND3 (N7165, N7157, N5250, N40);
not NOT1 (N7166, N7165);
nor NOR2 (N7167, N7159, N3062);
nor NOR4 (N7168, N7163, N1883, N3492, N2417);
and AND4 (N7169, N7155, N2560, N3089, N7147);
nor NOR2 (N7170, N7146, N6283);
not NOT1 (N7171, N7170);
buf BUF1 (N7172, N7169);
or OR3 (N7173, N7158, N1118, N4676);
xor XOR2 (N7174, N7167, N5450);
nor NOR3 (N7175, N7174, N6577, N1294);
and AND4 (N7176, N7164, N5656, N4147, N4378);
or OR3 (N7177, N7176, N377, N2586);
buf BUF1 (N7178, N7175);
nand NAND4 (N7179, N7149, N796, N4724, N5841);
nor NOR4 (N7180, N7135, N1461, N3962, N885);
not NOT1 (N7181, N7177);
nor NOR4 (N7182, N7179, N83, N1097, N3486);
xor XOR2 (N7183, N7181, N1014);
nand NAND4 (N7184, N7178, N4443, N504, N4212);
not NOT1 (N7185, N7173);
xor XOR2 (N7186, N7182, N6272);
xor XOR2 (N7187, N7183, N6035);
not NOT1 (N7188, N7186);
nor NOR4 (N7189, N7171, N293, N5589, N4068);
nor NOR2 (N7190, N7184, N6480);
or OR4 (N7191, N7168, N6367, N2524, N1799);
not NOT1 (N7192, N7187);
or OR4 (N7193, N7180, N7154, N1853, N4502);
and AND3 (N7194, N7190, N1608, N2508);
xor XOR2 (N7195, N7188, N5567);
xor XOR2 (N7196, N7189, N4730);
nand NAND3 (N7197, N7195, N833, N3383);
nor NOR2 (N7198, N7193, N2916);
nor NOR4 (N7199, N7191, N1767, N2870, N5001);
or OR2 (N7200, N7166, N701);
or OR4 (N7201, N7199, N5279, N2597, N5704);
nor NOR3 (N7202, N7198, N5688, N7094);
xor XOR2 (N7203, N7172, N4454);
xor XOR2 (N7204, N7196, N318);
buf BUF1 (N7205, N7200);
nor NOR3 (N7206, N7185, N690, N6512);
or OR2 (N7207, N7201, N2724);
xor XOR2 (N7208, N7202, N3588);
not NOT1 (N7209, N7207);
not NOT1 (N7210, N7197);
buf BUF1 (N7211, N7209);
xor XOR2 (N7212, N7204, N2503);
nor NOR3 (N7213, N7194, N3641, N1943);
nor NOR2 (N7214, N7208, N6812);
not NOT1 (N7215, N7212);
nor NOR2 (N7216, N7214, N5993);
and AND2 (N7217, N7205, N4013);
nor NOR4 (N7218, N7203, N2960, N5947, N3298);
or OR2 (N7219, N7216, N6839);
nand NAND2 (N7220, N7213, N6368);
nor NOR3 (N7221, N7217, N543, N170);
or OR3 (N7222, N7192, N4200, N5170);
not NOT1 (N7223, N7206);
and AND3 (N7224, N7221, N5039, N1777);
not NOT1 (N7225, N7150);
xor XOR2 (N7226, N7222, N6201);
buf BUF1 (N7227, N7224);
xor XOR2 (N7228, N7218, N2428);
and AND4 (N7229, N7219, N1292, N1667, N1809);
not NOT1 (N7230, N7226);
nand NAND3 (N7231, N7228, N4879, N2339);
or OR2 (N7232, N7230, N6192);
nor NOR3 (N7233, N7223, N4032, N2817);
and AND3 (N7234, N7215, N354, N4126);
buf BUF1 (N7235, N7220);
or OR2 (N7236, N7235, N4005);
xor XOR2 (N7237, N7227, N676);
or OR2 (N7238, N7231, N5717);
nor NOR4 (N7239, N7210, N2247, N474, N2040);
nor NOR2 (N7240, N7232, N2458);
buf BUF1 (N7241, N7238);
xor XOR2 (N7242, N7236, N6385);
buf BUF1 (N7243, N7241);
not NOT1 (N7244, N7229);
and AND4 (N7245, N7244, N1764, N7223, N4019);
or OR2 (N7246, N7245, N923);
buf BUF1 (N7247, N7211);
xor XOR2 (N7248, N7234, N4866);
and AND3 (N7249, N7247, N1315, N6432);
xor XOR2 (N7250, N7239, N4553);
xor XOR2 (N7251, N7233, N2996);
and AND3 (N7252, N7251, N5402, N4206);
nand NAND4 (N7253, N7248, N3594, N4815, N2332);
buf BUF1 (N7254, N7242);
xor XOR2 (N7255, N7240, N231);
or OR2 (N7256, N7252, N5835);
xor XOR2 (N7257, N7250, N3168);
not NOT1 (N7258, N7256);
not NOT1 (N7259, N7253);
or OR3 (N7260, N7237, N5967, N6130);
xor XOR2 (N7261, N7249, N569);
not NOT1 (N7262, N7260);
not NOT1 (N7263, N7243);
buf BUF1 (N7264, N7259);
xor XOR2 (N7265, N7258, N1061);
or OR3 (N7266, N7246, N615, N2143);
nor NOR3 (N7267, N7263, N22, N6406);
buf BUF1 (N7268, N7265);
or OR2 (N7269, N7225, N6959);
or OR2 (N7270, N7254, N4968);
xor XOR2 (N7271, N7270, N2371);
buf BUF1 (N7272, N7267);
buf BUF1 (N7273, N7264);
xor XOR2 (N7274, N7262, N6132);
nand NAND4 (N7275, N7255, N4256, N5167, N1357);
or OR3 (N7276, N7269, N4086, N2106);
nand NAND4 (N7277, N7272, N2093, N1493, N2116);
or OR4 (N7278, N7257, N4606, N5517, N2859);
nand NAND4 (N7279, N7266, N3252, N4804, N767);
xor XOR2 (N7280, N7276, N61);
nand NAND4 (N7281, N7278, N73, N1995, N1292);
buf BUF1 (N7282, N7273);
not NOT1 (N7283, N7281);
xor XOR2 (N7284, N7277, N1329);
xor XOR2 (N7285, N7279, N5074);
nor NOR2 (N7286, N7280, N1964);
nor NOR3 (N7287, N7285, N1207, N1679);
nor NOR3 (N7288, N7271, N2704, N5835);
nand NAND2 (N7289, N7288, N6558);
xor XOR2 (N7290, N7286, N6376);
and AND2 (N7291, N7284, N1071);
and AND4 (N7292, N7287, N6222, N3550, N6538);
and AND2 (N7293, N7289, N656);
nand NAND2 (N7294, N7274, N6445);
nand NAND2 (N7295, N7292, N2795);
nand NAND4 (N7296, N7295, N2020, N2016, N4);
buf BUF1 (N7297, N7290);
or OR2 (N7298, N7297, N1567);
or OR2 (N7299, N7291, N3853);
not NOT1 (N7300, N7282);
xor XOR2 (N7301, N7294, N4045);
nor NOR3 (N7302, N7293, N2103, N1488);
and AND4 (N7303, N7268, N827, N4127, N7216);
or OR2 (N7304, N7300, N4114);
nand NAND2 (N7305, N7303, N6381);
nand NAND4 (N7306, N7299, N4994, N1603, N6111);
buf BUF1 (N7307, N7304);
buf BUF1 (N7308, N7275);
xor XOR2 (N7309, N7305, N1613);
nor NOR4 (N7310, N7283, N312, N4876, N7197);
xor XOR2 (N7311, N7298, N5293);
not NOT1 (N7312, N7307);
buf BUF1 (N7313, N7302);
buf BUF1 (N7314, N7306);
nor NOR4 (N7315, N7310, N1306, N426, N2944);
buf BUF1 (N7316, N7296);
and AND3 (N7317, N7301, N2637, N6923);
and AND4 (N7318, N7311, N1642, N1715, N3288);
buf BUF1 (N7319, N7261);
not NOT1 (N7320, N7312);
not NOT1 (N7321, N7315);
or OR3 (N7322, N7313, N424, N4936);
not NOT1 (N7323, N7319);
xor XOR2 (N7324, N7323, N3898);
and AND2 (N7325, N7322, N628);
not NOT1 (N7326, N7325);
buf BUF1 (N7327, N7317);
not NOT1 (N7328, N7308);
buf BUF1 (N7329, N7320);
xor XOR2 (N7330, N7328, N3934);
nand NAND4 (N7331, N7324, N1512, N840, N6183);
xor XOR2 (N7332, N7318, N2612);
nor NOR2 (N7333, N7331, N1028);
xor XOR2 (N7334, N7329, N1740);
not NOT1 (N7335, N7334);
or OR3 (N7336, N7332, N7053, N1465);
nor NOR2 (N7337, N7326, N2751);
buf BUF1 (N7338, N7337);
nor NOR4 (N7339, N7330, N4214, N5663, N7035);
nand NAND2 (N7340, N7327, N5955);
xor XOR2 (N7341, N7314, N2398);
not NOT1 (N7342, N7321);
xor XOR2 (N7343, N7340, N7276);
not NOT1 (N7344, N7316);
not NOT1 (N7345, N7342);
not NOT1 (N7346, N7341);
not NOT1 (N7347, N7343);
not NOT1 (N7348, N7309);
or OR4 (N7349, N7346, N6219, N1885, N2383);
and AND3 (N7350, N7335, N990, N5811);
or OR3 (N7351, N7349, N4307, N1387);
or OR2 (N7352, N7339, N4738);
nand NAND2 (N7353, N7352, N3249);
not NOT1 (N7354, N7345);
and AND3 (N7355, N7347, N3797, N3669);
xor XOR2 (N7356, N7350, N3844);
not NOT1 (N7357, N7348);
or OR4 (N7358, N7336, N7140, N1768, N2389);
xor XOR2 (N7359, N7351, N6043);
nor NOR4 (N7360, N7356, N4051, N5895, N4499);
xor XOR2 (N7361, N7360, N3103);
nand NAND4 (N7362, N7354, N2008, N4905, N2403);
or OR4 (N7363, N7355, N888, N342, N5972);
buf BUF1 (N7364, N7344);
nand NAND3 (N7365, N7353, N5839, N1289);
buf BUF1 (N7366, N7338);
xor XOR2 (N7367, N7364, N764);
xor XOR2 (N7368, N7359, N4818);
xor XOR2 (N7369, N7333, N5534);
and AND2 (N7370, N7363, N1027);
xor XOR2 (N7371, N7366, N1442);
nor NOR4 (N7372, N7357, N4186, N5687, N4961);
and AND3 (N7373, N7372, N727, N2003);
or OR4 (N7374, N7367, N1496, N7297, N6397);
nor NOR2 (N7375, N7368, N5);
or OR3 (N7376, N7361, N1643, N5631);
and AND4 (N7377, N7370, N4754, N7090, N2127);
nor NOR4 (N7378, N7369, N6421, N4973, N4148);
nor NOR2 (N7379, N7373, N4289);
nor NOR4 (N7380, N7376, N6360, N1550, N6710);
and AND3 (N7381, N7377, N5743, N5646);
nor NOR4 (N7382, N7358, N4751, N5853, N4580);
or OR4 (N7383, N7371, N6119, N4871, N6576);
or OR2 (N7384, N7374, N6938);
nor NOR4 (N7385, N7382, N351, N6523, N1567);
xor XOR2 (N7386, N7381, N6157);
or OR4 (N7387, N7385, N2944, N1463, N5161);
or OR2 (N7388, N7387, N7345);
not NOT1 (N7389, N7365);
and AND2 (N7390, N7389, N2502);
and AND3 (N7391, N7386, N3982, N6598);
buf BUF1 (N7392, N7378);
buf BUF1 (N7393, N7388);
or OR4 (N7394, N7392, N3775, N3821, N5827);
not NOT1 (N7395, N7379);
buf BUF1 (N7396, N7391);
not NOT1 (N7397, N7380);
and AND4 (N7398, N7396, N5415, N7048, N4194);
xor XOR2 (N7399, N7390, N877);
buf BUF1 (N7400, N7398);
and AND4 (N7401, N7393, N1880, N2450, N1085);
buf BUF1 (N7402, N7399);
or OR3 (N7403, N7401, N4977, N4434);
or OR2 (N7404, N7375, N288);
nand NAND2 (N7405, N7397, N4503);
not NOT1 (N7406, N7394);
or OR4 (N7407, N7406, N5117, N5072, N5833);
buf BUF1 (N7408, N7404);
not NOT1 (N7409, N7384);
and AND3 (N7410, N7402, N5579, N3172);
nand NAND2 (N7411, N7405, N6224);
nand NAND2 (N7412, N7403, N2885);
and AND2 (N7413, N7383, N5628);
or OR3 (N7414, N7408, N1910, N3286);
buf BUF1 (N7415, N7409);
and AND3 (N7416, N7411, N3147, N1974);
or OR3 (N7417, N7362, N6124, N1430);
and AND4 (N7418, N7416, N1225, N1344, N2300);
not NOT1 (N7419, N7415);
and AND2 (N7420, N7413, N7240);
not NOT1 (N7421, N7417);
nor NOR4 (N7422, N7400, N3605, N2738, N3023);
nor NOR3 (N7423, N7418, N4943, N278);
xor XOR2 (N7424, N7423, N4855);
and AND4 (N7425, N7421, N6868, N1649, N926);
or OR3 (N7426, N7395, N2206, N507);
xor XOR2 (N7427, N7425, N665);
nand NAND4 (N7428, N7420, N1531, N4572, N683);
buf BUF1 (N7429, N7422);
and AND2 (N7430, N7407, N1475);
buf BUF1 (N7431, N7429);
nor NOR2 (N7432, N7428, N5287);
nor NOR3 (N7433, N7427, N6199, N7096);
or OR3 (N7434, N7424, N2911, N3203);
or OR2 (N7435, N7434, N5024);
buf BUF1 (N7436, N7435);
buf BUF1 (N7437, N7412);
not NOT1 (N7438, N7426);
and AND4 (N7439, N7419, N3634, N1659, N3484);
not NOT1 (N7440, N7439);
xor XOR2 (N7441, N7410, N3);
nand NAND4 (N7442, N7440, N3290, N4824, N5447);
not NOT1 (N7443, N7414);
or OR2 (N7444, N7432, N6079);
not NOT1 (N7445, N7438);
or OR2 (N7446, N7431, N4482);
buf BUF1 (N7447, N7443);
not NOT1 (N7448, N7447);
not NOT1 (N7449, N7446);
buf BUF1 (N7450, N7441);
nor NOR3 (N7451, N7442, N1168, N2260);
xor XOR2 (N7452, N7445, N3571);
xor XOR2 (N7453, N7444, N3571);
not NOT1 (N7454, N7437);
nor NOR4 (N7455, N7433, N275, N1440, N5812);
not NOT1 (N7456, N7430);
buf BUF1 (N7457, N7448);
xor XOR2 (N7458, N7451, N3301);
and AND2 (N7459, N7453, N4805);
or OR2 (N7460, N7449, N2100);
or OR3 (N7461, N7457, N2895, N4576);
nand NAND3 (N7462, N7436, N3855, N7240);
nand NAND3 (N7463, N7458, N5675, N5374);
nor NOR3 (N7464, N7452, N5413, N3444);
xor XOR2 (N7465, N7460, N1995);
or OR3 (N7466, N7450, N1349, N3133);
not NOT1 (N7467, N7456);
nor NOR2 (N7468, N7454, N6375);
buf BUF1 (N7469, N7467);
buf BUF1 (N7470, N7461);
buf BUF1 (N7471, N7464);
nand NAND2 (N7472, N7465, N3626);
buf BUF1 (N7473, N7469);
xor XOR2 (N7474, N7455, N443);
or OR3 (N7475, N7459, N2942, N7342);
not NOT1 (N7476, N7468);
and AND2 (N7477, N7472, N7179);
xor XOR2 (N7478, N7470, N6674);
buf BUF1 (N7479, N7475);
buf BUF1 (N7480, N7462);
xor XOR2 (N7481, N7466, N3524);
or OR3 (N7482, N7477, N515, N3795);
not NOT1 (N7483, N7480);
nor NOR4 (N7484, N7471, N2421, N6245, N2588);
nand NAND2 (N7485, N7482, N65);
buf BUF1 (N7486, N7473);
and AND4 (N7487, N7463, N7317, N5355, N4833);
or OR3 (N7488, N7478, N6923, N3103);
and AND2 (N7489, N7484, N7347);
buf BUF1 (N7490, N7486);
xor XOR2 (N7491, N7483, N6047);
nand NAND4 (N7492, N7481, N4881, N3097, N4161);
nand NAND3 (N7493, N7485, N2121, N5378);
nor NOR3 (N7494, N7492, N1408, N1391);
not NOT1 (N7495, N7494);
not NOT1 (N7496, N7490);
buf BUF1 (N7497, N7491);
xor XOR2 (N7498, N7476, N1812);
buf BUF1 (N7499, N7488);
or OR3 (N7500, N7496, N7144, N1779);
xor XOR2 (N7501, N7479, N2922);
nor NOR4 (N7502, N7501, N4763, N5555, N4362);
or OR3 (N7503, N7500, N4923, N4372);
buf BUF1 (N7504, N7502);
and AND3 (N7505, N7503, N5937, N7466);
and AND3 (N7506, N7499, N347, N608);
xor XOR2 (N7507, N7495, N1103);
nor NOR3 (N7508, N7493, N1407, N5807);
xor XOR2 (N7509, N7498, N4685);
nand NAND4 (N7510, N7506, N4369, N762, N3186);
nand NAND3 (N7511, N7497, N2364, N1535);
and AND4 (N7512, N7504, N6868, N4234, N5934);
or OR2 (N7513, N7511, N4679);
not NOT1 (N7514, N7510);
nand NAND4 (N7515, N7487, N6706, N665, N5194);
buf BUF1 (N7516, N7474);
and AND4 (N7517, N7505, N822, N7194, N3793);
nor NOR2 (N7518, N7515, N4324);
buf BUF1 (N7519, N7507);
xor XOR2 (N7520, N7518, N1269);
nand NAND2 (N7521, N7520, N3852);
nor NOR2 (N7522, N7516, N1318);
nand NAND2 (N7523, N7517, N1412);
and AND4 (N7524, N7513, N34, N6974, N4883);
and AND2 (N7525, N7514, N3650);
and AND2 (N7526, N7524, N6131);
nand NAND4 (N7527, N7525, N499, N6581, N6472);
nand NAND4 (N7528, N7527, N5705, N2370, N5520);
nor NOR4 (N7529, N7528, N1183, N4029, N3854);
nand NAND3 (N7530, N7529, N4542, N2002);
buf BUF1 (N7531, N7521);
xor XOR2 (N7532, N7508, N1633);
nor NOR4 (N7533, N7509, N2180, N1433, N6575);
or OR2 (N7534, N7523, N6985);
nor NOR3 (N7535, N7522, N2068, N3394);
not NOT1 (N7536, N7533);
buf BUF1 (N7537, N7531);
xor XOR2 (N7538, N7489, N6650);
not NOT1 (N7539, N7536);
nand NAND2 (N7540, N7535, N806);
and AND2 (N7541, N7526, N4589);
nor NOR4 (N7542, N7541, N5931, N4484, N2127);
nand NAND4 (N7543, N7538, N3687, N905, N218);
buf BUF1 (N7544, N7512);
nand NAND4 (N7545, N7532, N6391, N6879, N6303);
nand NAND4 (N7546, N7539, N2504, N6718, N5726);
or OR2 (N7547, N7534, N393);
or OR3 (N7548, N7545, N1896, N2643);
and AND2 (N7549, N7546, N2287);
buf BUF1 (N7550, N7548);
nor NOR3 (N7551, N7550, N5669, N4857);
and AND2 (N7552, N7543, N7033);
xor XOR2 (N7553, N7537, N3980);
and AND4 (N7554, N7547, N4830, N171, N4606);
nand NAND3 (N7555, N7540, N5532, N5242);
xor XOR2 (N7556, N7552, N7228);
xor XOR2 (N7557, N7555, N6955);
or OR4 (N7558, N7551, N6498, N3488, N7340);
nand NAND4 (N7559, N7556, N2621, N789, N821);
xor XOR2 (N7560, N7554, N6742);
and AND2 (N7561, N7557, N6690);
not NOT1 (N7562, N7549);
buf BUF1 (N7563, N7559);
and AND4 (N7564, N7542, N3892, N523, N2943);
buf BUF1 (N7565, N7558);
not NOT1 (N7566, N7519);
nand NAND4 (N7567, N7565, N117, N3231, N5170);
and AND2 (N7568, N7544, N5845);
or OR3 (N7569, N7560, N4384, N4206);
xor XOR2 (N7570, N7564, N334);
buf BUF1 (N7571, N7570);
xor XOR2 (N7572, N7530, N517);
not NOT1 (N7573, N7572);
or OR3 (N7574, N7573, N3616, N4245);
xor XOR2 (N7575, N7569, N2190);
nand NAND3 (N7576, N7574, N6658, N7011);
buf BUF1 (N7577, N7563);
xor XOR2 (N7578, N7567, N1261);
not NOT1 (N7579, N7568);
nand NAND3 (N7580, N7566, N5354, N4108);
buf BUF1 (N7581, N7553);
nand NAND2 (N7582, N7577, N215);
buf BUF1 (N7583, N7578);
buf BUF1 (N7584, N7576);
and AND2 (N7585, N7581, N979);
and AND4 (N7586, N7584, N2089, N6016, N3563);
nor NOR3 (N7587, N7579, N1653, N112);
nand NAND2 (N7588, N7575, N5420);
nand NAND2 (N7589, N7580, N3964);
or OR2 (N7590, N7583, N2358);
or OR3 (N7591, N7571, N4859, N3073);
or OR4 (N7592, N7587, N3211, N5662, N2523);
nand NAND3 (N7593, N7582, N4244, N5215);
nand NAND2 (N7594, N7561, N3184);
nand NAND3 (N7595, N7591, N4526, N2079);
or OR3 (N7596, N7595, N4976, N4553);
and AND2 (N7597, N7588, N7523);
xor XOR2 (N7598, N7589, N4497);
and AND2 (N7599, N7594, N6005);
nand NAND4 (N7600, N7599, N2648, N6887, N4501);
not NOT1 (N7601, N7600);
not NOT1 (N7602, N7597);
not NOT1 (N7603, N7586);
or OR2 (N7604, N7596, N4414);
xor XOR2 (N7605, N7590, N6901);
or OR2 (N7606, N7602, N1466);
and AND2 (N7607, N7606, N216);
xor XOR2 (N7608, N7562, N3123);
nor NOR2 (N7609, N7603, N3629);
or OR3 (N7610, N7593, N5476, N4939);
and AND2 (N7611, N7585, N273);
or OR3 (N7612, N7608, N1223, N4440);
xor XOR2 (N7613, N7605, N256);
xor XOR2 (N7614, N7611, N5295);
xor XOR2 (N7615, N7604, N5664);
buf BUF1 (N7616, N7615);
and AND2 (N7617, N7609, N4090);
xor XOR2 (N7618, N7613, N901);
nand NAND2 (N7619, N7592, N6246);
and AND3 (N7620, N7617, N2043, N278);
nand NAND3 (N7621, N7598, N1250, N753);
not NOT1 (N7622, N7616);
buf BUF1 (N7623, N7610);
nand NAND2 (N7624, N7618, N5758);
and AND2 (N7625, N7620, N6678);
buf BUF1 (N7626, N7622);
nand NAND3 (N7627, N7601, N7369, N1875);
not NOT1 (N7628, N7623);
xor XOR2 (N7629, N7628, N4438);
and AND3 (N7630, N7619, N5662, N3787);
and AND3 (N7631, N7626, N1910, N6147);
buf BUF1 (N7632, N7607);
buf BUF1 (N7633, N7629);
not NOT1 (N7634, N7625);
not NOT1 (N7635, N7627);
nand NAND2 (N7636, N7631, N3378);
nand NAND4 (N7637, N7635, N4903, N7096, N1302);
nor NOR2 (N7638, N7636, N7636);
not NOT1 (N7639, N7633);
or OR3 (N7640, N7630, N4016, N176);
nor NOR3 (N7641, N7640, N6103, N5756);
not NOT1 (N7642, N7634);
xor XOR2 (N7643, N7638, N4293);
not NOT1 (N7644, N7637);
nor NOR3 (N7645, N7614, N4761, N6041);
and AND3 (N7646, N7621, N193, N1476);
nand NAND3 (N7647, N7639, N2236, N1118);
nor NOR2 (N7648, N7642, N972);
buf BUF1 (N7649, N7645);
and AND2 (N7650, N7649, N5876);
buf BUF1 (N7651, N7644);
buf BUF1 (N7652, N7641);
nor NOR2 (N7653, N7612, N1737);
buf BUF1 (N7654, N7653);
and AND4 (N7655, N7650, N2077, N1930, N6269);
xor XOR2 (N7656, N7647, N964);
xor XOR2 (N7657, N7624, N1853);
nand NAND4 (N7658, N7651, N7594, N6194, N400);
xor XOR2 (N7659, N7656, N5389);
xor XOR2 (N7660, N7657, N4387);
nor NOR2 (N7661, N7654, N1553);
not NOT1 (N7662, N7660);
not NOT1 (N7663, N7655);
not NOT1 (N7664, N7632);
buf BUF1 (N7665, N7652);
nor NOR3 (N7666, N7661, N1979, N1101);
and AND2 (N7667, N7648, N169);
and AND3 (N7668, N7667, N1487, N3369);
nor NOR3 (N7669, N7664, N4645, N2377);
buf BUF1 (N7670, N7658);
xor XOR2 (N7671, N7669, N2414);
nor NOR4 (N7672, N7646, N595, N7578, N2465);
xor XOR2 (N7673, N7668, N6514);
xor XOR2 (N7674, N7672, N1825);
not NOT1 (N7675, N7666);
nand NAND3 (N7676, N7662, N5814, N4369);
not NOT1 (N7677, N7671);
buf BUF1 (N7678, N7673);
nor NOR3 (N7679, N7675, N2770, N4833);
buf BUF1 (N7680, N7663);
nor NOR3 (N7681, N7674, N4563, N5197);
xor XOR2 (N7682, N7643, N1186);
not NOT1 (N7683, N7681);
buf BUF1 (N7684, N7680);
not NOT1 (N7685, N7665);
not NOT1 (N7686, N7659);
nor NOR4 (N7687, N7670, N1217, N2801, N5390);
xor XOR2 (N7688, N7678, N1280);
not NOT1 (N7689, N7685);
nor NOR2 (N7690, N7688, N5401);
not NOT1 (N7691, N7689);
buf BUF1 (N7692, N7684);
or OR3 (N7693, N7679, N7384, N936);
nor NOR4 (N7694, N7676, N6193, N5347, N2234);
xor XOR2 (N7695, N7691, N4486);
buf BUF1 (N7696, N7695);
not NOT1 (N7697, N7694);
or OR4 (N7698, N7683, N3554, N7013, N7060);
buf BUF1 (N7699, N7692);
xor XOR2 (N7700, N7698, N4238);
nor NOR4 (N7701, N7687, N3521, N1005, N4695);
nor NOR3 (N7702, N7677, N4958, N914);
and AND3 (N7703, N7699, N3894, N1098);
or OR4 (N7704, N7700, N288, N2726, N6033);
nand NAND4 (N7705, N7701, N4726, N265, N310);
and AND4 (N7706, N7697, N4006, N1689, N4975);
buf BUF1 (N7707, N7682);
nand NAND3 (N7708, N7693, N2344, N2383);
and AND4 (N7709, N7696, N2095, N859, N3343);
nand NAND2 (N7710, N7706, N1228);
nor NOR3 (N7711, N7710, N3025, N1446);
buf BUF1 (N7712, N7704);
not NOT1 (N7713, N7709);
nand NAND2 (N7714, N7713, N710);
nor NOR2 (N7715, N7707, N6437);
and AND4 (N7716, N7690, N1237, N3306, N5670);
buf BUF1 (N7717, N7716);
nor NOR2 (N7718, N7717, N4292);
or OR3 (N7719, N7711, N4518, N2943);
or OR2 (N7720, N7686, N7470);
and AND4 (N7721, N7705, N6614, N6381, N351);
nor NOR2 (N7722, N7719, N6413);
buf BUF1 (N7723, N7715);
or OR4 (N7724, N7720, N5472, N3876, N6120);
xor XOR2 (N7725, N7702, N2654);
xor XOR2 (N7726, N7721, N3136);
xor XOR2 (N7727, N7718, N1448);
nand NAND3 (N7728, N7703, N5510, N5806);
not NOT1 (N7729, N7723);
buf BUF1 (N7730, N7714);
not NOT1 (N7731, N7724);
and AND3 (N7732, N7708, N3292, N6350);
nor NOR4 (N7733, N7712, N5485, N4189, N2035);
xor XOR2 (N7734, N7726, N6549);
nand NAND2 (N7735, N7731, N3152);
xor XOR2 (N7736, N7730, N1624);
buf BUF1 (N7737, N7722);
xor XOR2 (N7738, N7735, N3142);
and AND3 (N7739, N7736, N1985, N96);
xor XOR2 (N7740, N7725, N3908);
xor XOR2 (N7741, N7733, N1989);
xor XOR2 (N7742, N7727, N6790);
nor NOR3 (N7743, N7739, N3072, N3873);
buf BUF1 (N7744, N7743);
not NOT1 (N7745, N7737);
buf BUF1 (N7746, N7734);
or OR3 (N7747, N7738, N6114, N7520);
or OR2 (N7748, N7745, N7340);
nand NAND2 (N7749, N7741, N368);
and AND2 (N7750, N7747, N839);
nor NOR2 (N7751, N7740, N7500);
not NOT1 (N7752, N7749);
not NOT1 (N7753, N7751);
or OR2 (N7754, N7750, N5887);
nor NOR2 (N7755, N7729, N629);
or OR4 (N7756, N7732, N1570, N5636, N3545);
nand NAND2 (N7757, N7746, N5796);
and AND3 (N7758, N7752, N669, N4499);
buf BUF1 (N7759, N7742);
buf BUF1 (N7760, N7758);
buf BUF1 (N7761, N7748);
xor XOR2 (N7762, N7754, N1848);
xor XOR2 (N7763, N7744, N6823);
nand NAND2 (N7764, N7728, N1747);
buf BUF1 (N7765, N7763);
buf BUF1 (N7766, N7757);
nor NOR3 (N7767, N7764, N352, N1785);
buf BUF1 (N7768, N7765);
nor NOR2 (N7769, N7768, N2658);
xor XOR2 (N7770, N7761, N3581);
and AND2 (N7771, N7769, N2263);
not NOT1 (N7772, N7753);
buf BUF1 (N7773, N7771);
not NOT1 (N7774, N7767);
nand NAND3 (N7775, N7774, N2734, N4973);
and AND4 (N7776, N7773, N3374, N1693, N3155);
nor NOR3 (N7777, N7755, N3149, N5823);
not NOT1 (N7778, N7775);
or OR2 (N7779, N7759, N3574);
not NOT1 (N7780, N7762);
nand NAND3 (N7781, N7778, N5623, N2254);
not NOT1 (N7782, N7766);
nor NOR2 (N7783, N7772, N7072);
nand NAND2 (N7784, N7783, N2683);
and AND4 (N7785, N7779, N4077, N1210, N6616);
and AND4 (N7786, N7782, N5293, N2861, N7189);
buf BUF1 (N7787, N7785);
and AND4 (N7788, N7780, N7150, N2733, N3460);
or OR3 (N7789, N7770, N5595, N7508);
xor XOR2 (N7790, N7787, N7644);
or OR3 (N7791, N7760, N3053, N1197);
nor NOR4 (N7792, N7776, N5375, N7159, N2191);
nand NAND2 (N7793, N7756, N4968);
and AND4 (N7794, N7777, N2168, N109, N6655);
or OR2 (N7795, N7793, N546);
nand NAND2 (N7796, N7786, N6500);
xor XOR2 (N7797, N7796, N5893);
nand NAND2 (N7798, N7788, N747);
buf BUF1 (N7799, N7784);
not NOT1 (N7800, N7789);
not NOT1 (N7801, N7792);
not NOT1 (N7802, N7781);
and AND2 (N7803, N7800, N889);
xor XOR2 (N7804, N7795, N6141);
buf BUF1 (N7805, N7803);
or OR2 (N7806, N7797, N1053);
and AND3 (N7807, N7794, N2553, N720);
nand NAND2 (N7808, N7804, N4170);
buf BUF1 (N7809, N7801);
nor NOR3 (N7810, N7798, N5055, N2067);
nor NOR2 (N7811, N7809, N1025);
xor XOR2 (N7812, N7806, N6730);
and AND3 (N7813, N7807, N4996, N5042);
buf BUF1 (N7814, N7811);
buf BUF1 (N7815, N7799);
nand NAND4 (N7816, N7814, N7599, N791, N4858);
nand NAND2 (N7817, N7808, N3321);
xor XOR2 (N7818, N7817, N5574);
buf BUF1 (N7819, N7815);
xor XOR2 (N7820, N7818, N7404);
and AND2 (N7821, N7791, N4176);
or OR3 (N7822, N7816, N6754, N826);
xor XOR2 (N7823, N7820, N5636);
and AND3 (N7824, N7822, N3064, N7582);
nand NAND4 (N7825, N7819, N555, N2096, N6408);
not NOT1 (N7826, N7810);
or OR2 (N7827, N7805, N4680);
buf BUF1 (N7828, N7802);
xor XOR2 (N7829, N7826, N7513);
nand NAND4 (N7830, N7824, N1042, N496, N7072);
not NOT1 (N7831, N7790);
not NOT1 (N7832, N7830);
not NOT1 (N7833, N7827);
nand NAND4 (N7834, N7812, N4844, N6771, N2265);
buf BUF1 (N7835, N7832);
nor NOR4 (N7836, N7831, N3268, N5556, N174);
or OR4 (N7837, N7825, N924, N7759, N5814);
or OR4 (N7838, N7813, N6609, N572, N5512);
nor NOR4 (N7839, N7821, N1477, N2708, N2244);
nor NOR2 (N7840, N7828, N1809);
buf BUF1 (N7841, N7839);
nor NOR2 (N7842, N7833, N5569);
buf BUF1 (N7843, N7840);
xor XOR2 (N7844, N7837, N2291);
not NOT1 (N7845, N7843);
buf BUF1 (N7846, N7834);
and AND3 (N7847, N7846, N5837, N2301);
buf BUF1 (N7848, N7845);
buf BUF1 (N7849, N7823);
and AND2 (N7850, N7835, N7298);
or OR2 (N7851, N7848, N698);
buf BUF1 (N7852, N7851);
buf BUF1 (N7853, N7847);
or OR3 (N7854, N7829, N7157, N1234);
buf BUF1 (N7855, N7838);
not NOT1 (N7856, N7849);
nand NAND4 (N7857, N7853, N6475, N2935, N2731);
nor NOR3 (N7858, N7842, N6712, N1924);
nor NOR4 (N7859, N7857, N7412, N1728, N7548);
xor XOR2 (N7860, N7856, N3336);
nor NOR3 (N7861, N7858, N1010, N2938);
nand NAND2 (N7862, N7850, N1359);
and AND4 (N7863, N7862, N7209, N6692, N1185);
nor NOR2 (N7864, N7855, N1958);
or OR2 (N7865, N7854, N99);
xor XOR2 (N7866, N7841, N7047);
xor XOR2 (N7867, N7859, N1982);
and AND4 (N7868, N7852, N2532, N6062, N7378);
buf BUF1 (N7869, N7868);
not NOT1 (N7870, N7863);
or OR2 (N7871, N7864, N1697);
and AND2 (N7872, N7861, N5581);
buf BUF1 (N7873, N7865);
or OR3 (N7874, N7860, N5338, N1469);
or OR2 (N7875, N7870, N1422);
xor XOR2 (N7876, N7872, N4829);
and AND4 (N7877, N7867, N6512, N2695, N7224);
buf BUF1 (N7878, N7877);
xor XOR2 (N7879, N7874, N4111);
buf BUF1 (N7880, N7844);
nor NOR3 (N7881, N7869, N4007, N1614);
buf BUF1 (N7882, N7879);
nand NAND4 (N7883, N7875, N2757, N7449, N1374);
and AND2 (N7884, N7883, N4417);
and AND3 (N7885, N7884, N6206, N3790);
buf BUF1 (N7886, N7882);
or OR2 (N7887, N7878, N2369);
or OR3 (N7888, N7886, N4745, N106);
nor NOR2 (N7889, N7836, N2671);
nor NOR4 (N7890, N7887, N1061, N7856, N2736);
nand NAND2 (N7891, N7866, N2334);
buf BUF1 (N7892, N7880);
nor NOR2 (N7893, N7871, N7791);
xor XOR2 (N7894, N7876, N4748);
xor XOR2 (N7895, N7890, N7567);
and AND4 (N7896, N7895, N3700, N4274, N416);
not NOT1 (N7897, N7894);
or OR2 (N7898, N7888, N3952);
and AND4 (N7899, N7873, N3997, N4929, N4427);
or OR4 (N7900, N7897, N4328, N4355, N5009);
nand NAND2 (N7901, N7899, N6094);
and AND2 (N7902, N7901, N2387);
nand NAND2 (N7903, N7893, N2769);
nor NOR2 (N7904, N7891, N4487);
xor XOR2 (N7905, N7904, N4289);
nand NAND4 (N7906, N7900, N4129, N944, N2140);
xor XOR2 (N7907, N7902, N6836);
nand NAND2 (N7908, N7889, N3577);
and AND3 (N7909, N7903, N4635, N724);
nand NAND4 (N7910, N7896, N2273, N191, N5397);
nor NOR2 (N7911, N7906, N93);
nor NOR4 (N7912, N7911, N4672, N3995, N367);
and AND4 (N7913, N7905, N3603, N4256, N1539);
or OR4 (N7914, N7898, N6099, N2790, N3913);
buf BUF1 (N7915, N7914);
xor XOR2 (N7916, N7910, N3320);
nor NOR2 (N7917, N7892, N5155);
buf BUF1 (N7918, N7881);
xor XOR2 (N7919, N7885, N2172);
buf BUF1 (N7920, N7919);
buf BUF1 (N7921, N7916);
and AND2 (N7922, N7907, N3978);
and AND4 (N7923, N7915, N2605, N2142, N4639);
buf BUF1 (N7924, N7912);
buf BUF1 (N7925, N7921);
and AND2 (N7926, N7925, N7123);
and AND3 (N7927, N7913, N4066, N787);
not NOT1 (N7928, N7927);
and AND3 (N7929, N7922, N771, N7156);
or OR2 (N7930, N7917, N7262);
or OR4 (N7931, N7920, N161, N2823, N5353);
xor XOR2 (N7932, N7931, N3735);
xor XOR2 (N7933, N7930, N2480);
buf BUF1 (N7934, N7924);
buf BUF1 (N7935, N7926);
nor NOR4 (N7936, N7933, N4627, N5046, N1370);
xor XOR2 (N7937, N7935, N6841);
and AND3 (N7938, N7937, N2882, N2209);
xor XOR2 (N7939, N7938, N7269);
and AND2 (N7940, N7934, N2629);
or OR4 (N7941, N7908, N2260, N3911, N7904);
buf BUF1 (N7942, N7928);
nand NAND2 (N7943, N7923, N5093);
nand NAND3 (N7944, N7936, N7333, N3091);
buf BUF1 (N7945, N7941);
not NOT1 (N7946, N7909);
buf BUF1 (N7947, N7918);
or OR2 (N7948, N7932, N6169);
and AND2 (N7949, N7939, N3866);
nand NAND3 (N7950, N7940, N3861, N7686);
buf BUF1 (N7951, N7945);
xor XOR2 (N7952, N7950, N6408);
not NOT1 (N7953, N7948);
nor NOR3 (N7954, N7949, N7003, N1937);
not NOT1 (N7955, N7946);
xor XOR2 (N7956, N7944, N3815);
nor NOR4 (N7957, N7929, N85, N5615, N5403);
buf BUF1 (N7958, N7956);
xor XOR2 (N7959, N7943, N2896);
buf BUF1 (N7960, N7952);
nor NOR3 (N7961, N7954, N1339, N6585);
and AND2 (N7962, N7959, N1838);
nand NAND4 (N7963, N7962, N445, N3387, N3889);
nand NAND4 (N7964, N7953, N6193, N2236, N7141);
buf BUF1 (N7965, N7947);
xor XOR2 (N7966, N7961, N4373);
not NOT1 (N7967, N7963);
buf BUF1 (N7968, N7964);
nor NOR4 (N7969, N7955, N2187, N1485, N2907);
nor NOR4 (N7970, N7966, N7015, N460, N1221);
and AND2 (N7971, N7957, N5207);
and AND3 (N7972, N7968, N3471, N3808);
not NOT1 (N7973, N7969);
buf BUF1 (N7974, N7972);
buf BUF1 (N7975, N7958);
buf BUF1 (N7976, N7974);
nor NOR3 (N7977, N7975, N2052, N2234);
not NOT1 (N7978, N7960);
nor NOR4 (N7979, N7967, N714, N955, N5653);
or OR4 (N7980, N7942, N6596, N61, N4077);
nand NAND3 (N7981, N7979, N3729, N4363);
nor NOR3 (N7982, N7978, N769, N783);
not NOT1 (N7983, N7976);
xor XOR2 (N7984, N7965, N6430);
nand NAND3 (N7985, N7973, N4140, N7704);
and AND2 (N7986, N7951, N1121);
or OR2 (N7987, N7983, N2310);
not NOT1 (N7988, N7987);
not NOT1 (N7989, N7977);
xor XOR2 (N7990, N7980, N7797);
and AND4 (N7991, N7971, N159, N5762, N5526);
or OR3 (N7992, N7982, N5823, N6653);
buf BUF1 (N7993, N7970);
or OR4 (N7994, N7990, N656, N6547, N145);
buf BUF1 (N7995, N7984);
and AND2 (N7996, N7993, N6889);
or OR4 (N7997, N7989, N6079, N3775, N180);
and AND3 (N7998, N7997, N1822, N1610);
not NOT1 (N7999, N7981);
buf BUF1 (N8000, N7999);
nor NOR3 (N8001, N7996, N698, N7829);
buf BUF1 (N8002, N7985);
buf BUF1 (N8003, N7994);
nor NOR4 (N8004, N8003, N3330, N5027, N2655);
buf BUF1 (N8005, N7986);
not NOT1 (N8006, N7991);
and AND3 (N8007, N8001, N6848, N4706);
xor XOR2 (N8008, N7998, N252);
or OR4 (N8009, N8000, N7583, N5844, N6897);
buf BUF1 (N8010, N7995);
xor XOR2 (N8011, N8006, N1566);
buf BUF1 (N8012, N8009);
xor XOR2 (N8013, N8007, N7942);
or OR3 (N8014, N8002, N1832, N3644);
endmodule