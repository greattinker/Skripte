// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N206,N203,N218,N196,N216,N212,N215,N208,N219;

xor XOR2 (N20, N18, N13);
buf BUF1 (N21, N16);
or OR4 (N22, N12, N20, N8, N1);
and AND4 (N23, N6, N13, N20, N19);
and AND3 (N24, N12, N7, N17);
buf BUF1 (N25, N16);
buf BUF1 (N26, N25);
nand NAND3 (N27, N2, N7, N7);
not NOT1 (N28, N22);
and AND2 (N29, N12, N23);
nor NOR4 (N30, N27, N5, N21, N10);
nand NAND2 (N31, N17, N25);
nor NOR3 (N32, N10, N6, N27);
not NOT1 (N33, N29);
and AND4 (N34, N17, N12, N14, N22);
nor NOR4 (N35, N21, N21, N17, N33);
and AND2 (N36, N33, N23);
and AND3 (N37, N32, N2, N21);
not NOT1 (N38, N24);
xor XOR2 (N39, N9, N33);
nor NOR4 (N40, N31, N27, N9, N20);
or OR2 (N41, N30, N4);
nor NOR2 (N42, N26, N21);
nor NOR2 (N43, N42, N29);
xor XOR2 (N44, N34, N23);
nor NOR2 (N45, N35, N12);
not NOT1 (N46, N41);
or OR3 (N47, N40, N32, N20);
nor NOR4 (N48, N28, N23, N35, N44);
buf BUF1 (N49, N25);
not NOT1 (N50, N48);
not NOT1 (N51, N43);
not NOT1 (N52, N38);
or OR4 (N53, N36, N8, N16, N15);
nand NAND3 (N54, N50, N4, N11);
nand NAND3 (N55, N45, N43, N10);
nand NAND2 (N56, N47, N54);
xor XOR2 (N57, N44, N33);
nand NAND3 (N58, N39, N39, N12);
nor NOR4 (N59, N52, N30, N12, N46);
nor NOR2 (N60, N8, N48);
nor NOR2 (N61, N59, N52);
nand NAND2 (N62, N49, N41);
xor XOR2 (N63, N53, N7);
or OR3 (N64, N57, N33, N1);
buf BUF1 (N65, N61);
or OR2 (N66, N58, N42);
or OR2 (N67, N56, N57);
nand NAND4 (N68, N63, N60, N60, N23);
buf BUF1 (N69, N46);
not NOT1 (N70, N67);
not NOT1 (N71, N62);
and AND4 (N72, N70, N7, N69, N55);
nand NAND2 (N73, N57, N32);
or OR2 (N74, N63, N62);
not NOT1 (N75, N66);
nand NAND3 (N76, N73, N72, N15);
or OR3 (N77, N75, N57, N25);
and AND2 (N78, N12, N4);
or OR2 (N79, N77, N5);
nor NOR3 (N80, N74, N12, N69);
and AND3 (N81, N64, N44, N80);
nor NOR3 (N82, N78, N24, N37);
xor XOR2 (N83, N8, N9);
xor XOR2 (N84, N7, N37);
and AND4 (N85, N71, N44, N71, N84);
or OR3 (N86, N69, N2, N82);
nor NOR3 (N87, N32, N79, N62);
not NOT1 (N88, N21);
xor XOR2 (N89, N85, N76);
not NOT1 (N90, N50);
nor NOR3 (N91, N86, N35, N40);
and AND4 (N92, N90, N83, N50, N40);
not NOT1 (N93, N62);
not NOT1 (N94, N93);
or OR2 (N95, N92, N65);
buf BUF1 (N96, N71);
not NOT1 (N97, N96);
buf BUF1 (N98, N68);
nand NAND2 (N99, N94, N81);
xor XOR2 (N100, N44, N96);
and AND2 (N101, N100, N67);
buf BUF1 (N102, N98);
nor NOR2 (N103, N101, N39);
nand NAND2 (N104, N103, N102);
and AND2 (N105, N29, N83);
buf BUF1 (N106, N97);
nor NOR4 (N107, N88, N106, N76, N34);
not NOT1 (N108, N52);
and AND4 (N109, N105, N31, N66, N30);
or OR3 (N110, N87, N25, N108);
nand NAND2 (N111, N74, N60);
and AND3 (N112, N51, N58, N65);
nor NOR3 (N113, N91, N86, N107);
nand NAND4 (N114, N104, N85, N6, N61);
and AND3 (N115, N30, N54, N90);
or OR3 (N116, N112, N35, N40);
nand NAND4 (N117, N99, N25, N112, N93);
not NOT1 (N118, N109);
xor XOR2 (N119, N111, N115);
and AND2 (N120, N18, N6);
not NOT1 (N121, N113);
nand NAND4 (N122, N120, N15, N43, N7);
not NOT1 (N123, N110);
xor XOR2 (N124, N114, N38);
nor NOR2 (N125, N122, N21);
buf BUF1 (N126, N118);
nand NAND4 (N127, N123, N54, N13, N4);
buf BUF1 (N128, N124);
buf BUF1 (N129, N89);
nand NAND3 (N130, N126, N66, N20);
and AND4 (N131, N125, N114, N71, N37);
nor NOR4 (N132, N121, N9, N23, N102);
and AND4 (N133, N117, N121, N120, N94);
nand NAND3 (N134, N128, N37, N108);
xor XOR2 (N135, N119, N30);
and AND4 (N136, N95, N134, N123, N128);
nor NOR2 (N137, N26, N3);
or OR2 (N138, N116, N20);
or OR4 (N139, N133, N45, N122, N33);
not NOT1 (N140, N138);
xor XOR2 (N141, N127, N57);
nor NOR2 (N142, N141, N7);
xor XOR2 (N143, N139, N49);
and AND4 (N144, N143, N22, N5, N76);
nand NAND2 (N145, N131, N41);
not NOT1 (N146, N144);
nand NAND4 (N147, N129, N103, N94, N117);
xor XOR2 (N148, N132, N71);
or OR2 (N149, N130, N61);
buf BUF1 (N150, N136);
nand NAND3 (N151, N146, N120, N117);
buf BUF1 (N152, N145);
and AND3 (N153, N135, N41, N69);
or OR4 (N154, N137, N81, N6, N76);
not NOT1 (N155, N153);
nor NOR4 (N156, N151, N34, N140, N82);
buf BUF1 (N157, N51);
xor XOR2 (N158, N156, N7);
or OR2 (N159, N152, N69);
not NOT1 (N160, N150);
or OR3 (N161, N155, N14, N32);
nor NOR2 (N162, N147, N116);
and AND2 (N163, N142, N90);
nand NAND2 (N164, N149, N22);
and AND4 (N165, N154, N61, N61, N29);
and AND2 (N166, N159, N94);
and AND3 (N167, N148, N147, N4);
nand NAND3 (N168, N158, N64, N18);
nor NOR3 (N169, N167, N56, N29);
and AND3 (N170, N166, N4, N168);
and AND2 (N171, N159, N151);
not NOT1 (N172, N160);
not NOT1 (N173, N171);
and AND2 (N174, N169, N102);
not NOT1 (N175, N163);
or OR2 (N176, N175, N22);
nor NOR2 (N177, N173, N74);
and AND3 (N178, N176, N104, N128);
not NOT1 (N179, N170);
nand NAND4 (N180, N165, N147, N160, N134);
xor XOR2 (N181, N179, N151);
nand NAND4 (N182, N180, N15, N70, N19);
or OR3 (N183, N162, N116, N62);
buf BUF1 (N184, N174);
nand NAND3 (N185, N172, N183, N115);
nand NAND4 (N186, N111, N44, N87, N45);
not NOT1 (N187, N182);
buf BUF1 (N188, N184);
xor XOR2 (N189, N164, N56);
xor XOR2 (N190, N187, N109);
xor XOR2 (N191, N186, N8);
not NOT1 (N192, N181);
nand NAND2 (N193, N185, N131);
and AND3 (N194, N157, N149, N166);
or OR4 (N195, N188, N36, N149, N128);
nor NOR3 (N196, N189, N172, N81);
nor NOR4 (N197, N190, N158, N78, N132);
not NOT1 (N198, N177);
xor XOR2 (N199, N191, N88);
and AND2 (N200, N195, N31);
nand NAND4 (N201, N194, N82, N198, N69);
and AND4 (N202, N120, N104, N60, N21);
xor XOR2 (N203, N202, N110);
or OR2 (N204, N197, N133);
nand NAND4 (N205, N193, N45, N17, N125);
or OR2 (N206, N204, N73);
nor NOR4 (N207, N178, N204, N121, N108);
nor NOR2 (N208, N199, N101);
xor XOR2 (N209, N200, N29);
or OR2 (N210, N201, N100);
buf BUF1 (N211, N161);
not NOT1 (N212, N209);
not NOT1 (N213, N207);
nor NOR3 (N214, N205, N52, N200);
not NOT1 (N215, N192);
nor NOR2 (N216, N213, N9);
buf BUF1 (N217, N210);
nand NAND2 (N218, N217, N192);
and AND4 (N219, N211, N214, N68, N173);
endmodule