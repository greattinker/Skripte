// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N6416,N6411,N6415,N6412,N6413,N6417,N6406,N6399,N6414,N6418;

and AND3 (N19, N7, N4, N3);
buf BUF1 (N20, N19);
not NOT1 (N21, N12);
xor XOR2 (N22, N8, N19);
not NOT1 (N23, N20);
nand NAND3 (N24, N15, N23, N2);
xor XOR2 (N25, N3, N7);
and AND3 (N26, N7, N6, N11);
buf BUF1 (N27, N12);
buf BUF1 (N28, N8);
not NOT1 (N29, N6);
not NOT1 (N30, N16);
or OR3 (N31, N15, N25, N8);
not NOT1 (N32, N2);
nand NAND4 (N33, N29, N19, N15, N32);
nor NOR2 (N34, N31, N24);
or OR3 (N35, N8, N26, N23);
nand NAND3 (N36, N21, N24, N25);
xor XOR2 (N37, N5, N13);
and AND3 (N38, N33, N28, N25);
xor XOR2 (N39, N9, N2);
and AND4 (N40, N5, N16, N30, N27);
and AND3 (N41, N32, N10, N25);
nor NOR3 (N42, N35, N28, N41);
nand NAND3 (N43, N1, N20, N28);
nor NOR4 (N44, N30, N40, N11, N5);
or OR2 (N45, N42, N37);
nand NAND3 (N46, N5, N1, N42);
or OR4 (N47, N12, N43, N39, N25);
and AND2 (N48, N44, N28);
or OR2 (N49, N23, N5);
and AND2 (N50, N25, N8);
or OR2 (N51, N34, N13);
not NOT1 (N52, N48);
buf BUF1 (N53, N46);
and AND2 (N54, N51, N44);
buf BUF1 (N55, N53);
and AND2 (N56, N22, N25);
and AND2 (N57, N56, N17);
nor NOR4 (N58, N38, N19, N13, N53);
not NOT1 (N59, N52);
nand NAND2 (N60, N49, N20);
nand NAND3 (N61, N54, N55, N27);
nor NOR4 (N62, N17, N19, N11, N15);
nor NOR3 (N63, N57, N10, N10);
nand NAND2 (N64, N36, N41);
nor NOR4 (N65, N62, N36, N6, N43);
and AND2 (N66, N59, N12);
buf BUF1 (N67, N64);
or OR3 (N68, N67, N61, N49);
nand NAND2 (N69, N17, N44);
xor XOR2 (N70, N69, N38);
buf BUF1 (N71, N65);
xor XOR2 (N72, N63, N21);
and AND2 (N73, N66, N33);
nor NOR3 (N74, N72, N30, N22);
not NOT1 (N75, N60);
not NOT1 (N76, N50);
not NOT1 (N77, N75);
and AND3 (N78, N58, N57, N14);
nand NAND2 (N79, N68, N76);
not NOT1 (N80, N68);
and AND2 (N81, N74, N72);
buf BUF1 (N82, N73);
not NOT1 (N83, N80);
and AND4 (N84, N83, N67, N33, N53);
and AND2 (N85, N79, N63);
buf BUF1 (N86, N70);
and AND2 (N87, N47, N73);
nand NAND3 (N88, N86, N8, N48);
xor XOR2 (N89, N85, N27);
nand NAND4 (N90, N89, N33, N49, N70);
nor NOR2 (N91, N81, N57);
and AND4 (N92, N84, N84, N24, N57);
and AND4 (N93, N88, N73, N70, N1);
not NOT1 (N94, N93);
xor XOR2 (N95, N78, N94);
not NOT1 (N96, N1);
or OR4 (N97, N95, N94, N1, N64);
and AND3 (N98, N92, N1, N39);
or OR2 (N99, N71, N91);
nor NOR2 (N100, N43, N91);
nand NAND2 (N101, N97, N67);
xor XOR2 (N102, N90, N49);
and AND4 (N103, N101, N34, N84, N76);
and AND4 (N104, N100, N49, N45, N55);
nand NAND2 (N105, N57, N9);
buf BUF1 (N106, N104);
nand NAND4 (N107, N82, N60, N64, N24);
not NOT1 (N108, N107);
not NOT1 (N109, N77);
nand NAND3 (N110, N87, N15, N42);
nor NOR3 (N111, N99, N20, N3);
not NOT1 (N112, N109);
not NOT1 (N113, N96);
nor NOR2 (N114, N113, N111);
not NOT1 (N115, N47);
or OR3 (N116, N110, N90, N39);
nor NOR3 (N117, N105, N49, N77);
buf BUF1 (N118, N106);
not NOT1 (N119, N114);
nor NOR4 (N120, N112, N40, N5, N10);
and AND2 (N121, N115, N91);
nand NAND3 (N122, N98, N59, N88);
nor NOR2 (N123, N103, N85);
nand NAND2 (N124, N108, N106);
nor NOR4 (N125, N122, N69, N35, N107);
xor XOR2 (N126, N123, N67);
buf BUF1 (N127, N118);
buf BUF1 (N128, N102);
nand NAND3 (N129, N117, N117, N61);
or OR4 (N130, N127, N115, N66, N50);
xor XOR2 (N131, N119, N48);
not NOT1 (N132, N131);
buf BUF1 (N133, N129);
or OR2 (N134, N126, N88);
nor NOR4 (N135, N130, N62, N130, N21);
and AND4 (N136, N116, N57, N10, N91);
not NOT1 (N137, N134);
or OR3 (N138, N136, N94, N61);
or OR2 (N139, N120, N136);
not NOT1 (N140, N121);
not NOT1 (N141, N140);
nand NAND4 (N142, N133, N57, N80, N93);
and AND3 (N143, N132, N23, N66);
nand NAND2 (N144, N124, N79);
xor XOR2 (N145, N128, N116);
or OR3 (N146, N135, N134, N84);
xor XOR2 (N147, N137, N3);
not NOT1 (N148, N125);
xor XOR2 (N149, N144, N42);
nand NAND2 (N150, N141, N23);
buf BUF1 (N151, N147);
xor XOR2 (N152, N139, N32);
nor NOR3 (N153, N138, N73, N27);
not NOT1 (N154, N152);
nand NAND2 (N155, N146, N138);
and AND2 (N156, N155, N129);
xor XOR2 (N157, N150, N117);
not NOT1 (N158, N154);
and AND4 (N159, N156, N66, N138, N139);
and AND2 (N160, N143, N137);
not NOT1 (N161, N142);
or OR4 (N162, N149, N144, N43, N121);
or OR2 (N163, N162, N73);
or OR3 (N164, N158, N157, N19);
nand NAND3 (N165, N119, N78, N58);
buf BUF1 (N166, N161);
nor NOR4 (N167, N163, N166, N48, N98);
nor NOR4 (N168, N110, N54, N114, N23);
or OR3 (N169, N164, N80, N120);
nor NOR3 (N170, N151, N4, N132);
buf BUF1 (N171, N148);
and AND2 (N172, N170, N112);
nor NOR4 (N173, N171, N39, N120, N107);
or OR3 (N174, N153, N123, N162);
not NOT1 (N175, N174);
or OR3 (N176, N172, N28, N2);
xor XOR2 (N177, N168, N1);
xor XOR2 (N178, N175, N118);
xor XOR2 (N179, N159, N9);
or OR4 (N180, N165, N117, N157, N140);
nand NAND3 (N181, N178, N11, N147);
xor XOR2 (N182, N167, N4);
and AND4 (N183, N176, N116, N4, N50);
xor XOR2 (N184, N145, N47);
or OR4 (N185, N180, N125, N109, N125);
xor XOR2 (N186, N177, N77);
nor NOR3 (N187, N184, N62, N87);
xor XOR2 (N188, N179, N121);
nand NAND2 (N189, N173, N128);
and AND4 (N190, N182, N47, N16, N109);
nand NAND3 (N191, N185, N21, N119);
nand NAND2 (N192, N189, N45);
xor XOR2 (N193, N192, N181);
and AND4 (N194, N89, N28, N120, N17);
or OR2 (N195, N194, N109);
xor XOR2 (N196, N183, N185);
buf BUF1 (N197, N169);
not NOT1 (N198, N196);
buf BUF1 (N199, N160);
and AND3 (N200, N186, N157, N165);
and AND3 (N201, N193, N10, N10);
nor NOR4 (N202, N191, N34, N198, N85);
xor XOR2 (N203, N13, N152);
or OR2 (N204, N197, N139);
nor NOR4 (N205, N202, N30, N95, N25);
not NOT1 (N206, N188);
and AND4 (N207, N187, N120, N179, N92);
nand NAND2 (N208, N199, N85);
nor NOR3 (N209, N206, N31, N89);
nand NAND3 (N210, N205, N124, N60);
not NOT1 (N211, N204);
not NOT1 (N212, N190);
nor NOR2 (N213, N212, N99);
xor XOR2 (N214, N207, N55);
not NOT1 (N215, N211);
nand NAND3 (N216, N208, N63, N127);
nand NAND4 (N217, N216, N156, N125, N86);
and AND2 (N218, N209, N87);
nand NAND4 (N219, N213, N65, N58, N204);
buf BUF1 (N220, N200);
xor XOR2 (N221, N218, N172);
buf BUF1 (N222, N219);
and AND4 (N223, N214, N114, N220, N114);
buf BUF1 (N224, N113);
or OR4 (N225, N201, N191, N116, N12);
buf BUF1 (N226, N217);
xor XOR2 (N227, N226, N204);
buf BUF1 (N228, N227);
nand NAND3 (N229, N195, N145, N205);
nor NOR4 (N230, N221, N112, N95, N29);
nor NOR2 (N231, N229, N13);
not NOT1 (N232, N225);
nand NAND4 (N233, N231, N150, N105, N60);
xor XOR2 (N234, N215, N230);
xor XOR2 (N235, N125, N123);
or OR4 (N236, N232, N224, N61, N2);
not NOT1 (N237, N47);
buf BUF1 (N238, N236);
xor XOR2 (N239, N234, N10);
or OR4 (N240, N238, N35, N64, N140);
or OR2 (N241, N233, N68);
not NOT1 (N242, N241);
and AND2 (N243, N242, N5);
and AND3 (N244, N240, N6, N200);
not NOT1 (N245, N223);
not NOT1 (N246, N245);
xor XOR2 (N247, N239, N135);
xor XOR2 (N248, N246, N153);
and AND4 (N249, N235, N76, N41, N231);
xor XOR2 (N250, N210, N28);
and AND4 (N251, N250, N143, N210, N241);
not NOT1 (N252, N203);
buf BUF1 (N253, N247);
buf BUF1 (N254, N237);
not NOT1 (N255, N244);
or OR3 (N256, N251, N249, N211);
or OR4 (N257, N231, N196, N111, N231);
nor NOR2 (N258, N256, N140);
not NOT1 (N259, N222);
buf BUF1 (N260, N254);
buf BUF1 (N261, N248);
buf BUF1 (N262, N261);
nand NAND2 (N263, N252, N252);
or OR3 (N264, N228, N98, N156);
or OR2 (N265, N262, N260);
and AND2 (N266, N205, N165);
buf BUF1 (N267, N255);
not NOT1 (N268, N257);
not NOT1 (N269, N259);
nor NOR3 (N270, N264, N54, N42);
and AND4 (N271, N269, N71, N87, N217);
not NOT1 (N272, N258);
and AND2 (N273, N270, N56);
xor XOR2 (N274, N268, N69);
nand NAND2 (N275, N267, N197);
not NOT1 (N276, N272);
or OR3 (N277, N271, N273, N258);
and AND3 (N278, N11, N270, N67);
nor NOR4 (N279, N263, N94, N168, N204);
nor NOR3 (N280, N278, N79, N148);
nand NAND3 (N281, N279, N99, N86);
and AND2 (N282, N280, N9);
nand NAND3 (N283, N243, N183, N7);
nand NAND4 (N284, N253, N219, N212, N163);
or OR2 (N285, N284, N95);
nor NOR2 (N286, N265, N19);
buf BUF1 (N287, N285);
xor XOR2 (N288, N287, N282);
or OR2 (N289, N71, N251);
or OR2 (N290, N266, N55);
buf BUF1 (N291, N274);
or OR2 (N292, N291, N26);
xor XOR2 (N293, N286, N259);
nor NOR4 (N294, N281, N207, N83, N8);
not NOT1 (N295, N275);
or OR2 (N296, N293, N189);
or OR3 (N297, N277, N82, N169);
buf BUF1 (N298, N283);
or OR2 (N299, N297, N270);
nand NAND4 (N300, N295, N126, N204, N108);
buf BUF1 (N301, N299);
nor NOR4 (N302, N300, N90, N222, N8);
buf BUF1 (N303, N276);
xor XOR2 (N304, N303, N120);
nor NOR2 (N305, N290, N4);
nor NOR4 (N306, N296, N270, N112, N60);
xor XOR2 (N307, N294, N61);
nand NAND4 (N308, N304, N44, N265, N261);
buf BUF1 (N309, N289);
buf BUF1 (N310, N308);
or OR3 (N311, N288, N245, N216);
buf BUF1 (N312, N311);
nand NAND2 (N313, N301, N122);
nor NOR2 (N314, N306, N102);
nand NAND3 (N315, N307, N149, N80);
xor XOR2 (N316, N314, N249);
nand NAND4 (N317, N313, N316, N34, N52);
nor NOR2 (N318, N140, N220);
nor NOR4 (N319, N310, N91, N80, N305);
buf BUF1 (N320, N179);
xor XOR2 (N321, N315, N243);
or OR4 (N322, N292, N211, N149, N136);
and AND2 (N323, N321, N37);
nor NOR4 (N324, N302, N96, N196, N154);
and AND4 (N325, N317, N185, N285, N275);
or OR3 (N326, N298, N3, N115);
nor NOR3 (N327, N323, N100, N286);
not NOT1 (N328, N312);
buf BUF1 (N329, N326);
not NOT1 (N330, N309);
and AND4 (N331, N322, N93, N94, N323);
nand NAND3 (N332, N329, N22, N101);
nor NOR2 (N333, N325, N80);
not NOT1 (N334, N333);
nand NAND3 (N335, N319, N118, N116);
buf BUF1 (N336, N331);
or OR4 (N337, N332, N152, N138, N146);
and AND4 (N338, N324, N117, N254, N328);
nand NAND4 (N339, N106, N74, N121, N1);
or OR3 (N340, N318, N59, N23);
nand NAND4 (N341, N340, N248, N226, N35);
or OR3 (N342, N330, N253, N178);
or OR4 (N343, N342, N129, N159, N269);
nor NOR4 (N344, N327, N161, N155, N67);
nor NOR4 (N345, N334, N119, N104, N235);
not NOT1 (N346, N343);
not NOT1 (N347, N336);
buf BUF1 (N348, N346);
or OR4 (N349, N345, N106, N237, N214);
nand NAND4 (N350, N320, N194, N334, N169);
xor XOR2 (N351, N349, N212);
nor NOR4 (N352, N348, N321, N93, N6);
nor NOR4 (N353, N341, N104, N10, N287);
or OR2 (N354, N338, N47);
xor XOR2 (N355, N352, N287);
and AND2 (N356, N347, N117);
or OR3 (N357, N351, N241, N111);
nand NAND2 (N358, N354, N22);
nor NOR2 (N359, N350, N158);
xor XOR2 (N360, N355, N135);
buf BUF1 (N361, N339);
buf BUF1 (N362, N337);
not NOT1 (N363, N356);
buf BUF1 (N364, N357);
nand NAND4 (N365, N360, N170, N304, N358);
not NOT1 (N366, N130);
not NOT1 (N367, N366);
xor XOR2 (N368, N364, N222);
or OR3 (N369, N359, N352, N261);
and AND3 (N370, N368, N233, N311);
or OR2 (N371, N361, N270);
and AND3 (N372, N371, N78, N309);
not NOT1 (N373, N353);
nand NAND3 (N374, N344, N285, N360);
nor NOR4 (N375, N372, N16, N114, N60);
nor NOR3 (N376, N335, N322, N227);
xor XOR2 (N377, N376, N336);
nand NAND4 (N378, N377, N266, N300, N180);
nand NAND2 (N379, N375, N85);
or OR2 (N380, N369, N121);
and AND3 (N381, N363, N107, N372);
and AND3 (N382, N373, N113, N319);
xor XOR2 (N383, N362, N11);
or OR2 (N384, N374, N221);
or OR2 (N385, N383, N219);
nor NOR2 (N386, N382, N337);
not NOT1 (N387, N386);
and AND4 (N388, N378, N270, N238, N288);
nor NOR4 (N389, N387, N371, N36, N82);
not NOT1 (N390, N380);
xor XOR2 (N391, N384, N265);
not NOT1 (N392, N389);
or OR2 (N393, N390, N135);
nor NOR2 (N394, N388, N44);
and AND2 (N395, N379, N264);
and AND2 (N396, N370, N216);
xor XOR2 (N397, N391, N72);
and AND2 (N398, N385, N232);
nand NAND4 (N399, N365, N117, N175, N297);
or OR4 (N400, N393, N150, N209, N136);
not NOT1 (N401, N394);
nand NAND4 (N402, N397, N205, N300, N150);
and AND3 (N403, N396, N163, N18);
not NOT1 (N404, N399);
or OR3 (N405, N392, N80, N250);
nand NAND2 (N406, N398, N403);
xor XOR2 (N407, N171, N109);
xor XOR2 (N408, N367, N247);
buf BUF1 (N409, N408);
nand NAND3 (N410, N405, N306, N281);
nand NAND3 (N411, N407, N22, N381);
buf BUF1 (N412, N265);
nor NOR3 (N413, N400, N52, N97);
nor NOR3 (N414, N410, N276, N104);
and AND3 (N415, N401, N101, N132);
nand NAND4 (N416, N414, N69, N318, N8);
and AND4 (N417, N413, N181, N311, N334);
buf BUF1 (N418, N411);
xor XOR2 (N419, N409, N77);
and AND4 (N420, N406, N304, N41, N250);
buf BUF1 (N421, N402);
nand NAND3 (N422, N415, N164, N27);
or OR3 (N423, N395, N198, N83);
nand NAND2 (N424, N404, N360);
nor NOR4 (N425, N412, N402, N329, N392);
and AND4 (N426, N418, N6, N58, N395);
nand NAND3 (N427, N421, N148, N251);
and AND3 (N428, N427, N347, N421);
or OR4 (N429, N417, N21, N217, N101);
and AND2 (N430, N416, N195);
nor NOR3 (N431, N425, N232, N208);
and AND2 (N432, N429, N391);
buf BUF1 (N433, N431);
and AND3 (N434, N433, N327, N217);
xor XOR2 (N435, N420, N224);
not NOT1 (N436, N422);
not NOT1 (N437, N426);
nand NAND2 (N438, N423, N390);
and AND4 (N439, N438, N406, N310, N185);
nand NAND2 (N440, N432, N348);
nor NOR4 (N441, N437, N64, N207, N246);
xor XOR2 (N442, N428, N438);
buf BUF1 (N443, N434);
buf BUF1 (N444, N435);
and AND4 (N445, N440, N252, N383, N295);
nand NAND2 (N446, N424, N325);
or OR3 (N447, N445, N299, N35);
xor XOR2 (N448, N436, N222);
nor NOR3 (N449, N444, N318, N407);
or OR3 (N450, N449, N353, N435);
nand NAND4 (N451, N443, N82, N248, N259);
or OR2 (N452, N441, N164);
or OR3 (N453, N447, N332, N137);
xor XOR2 (N454, N448, N17);
nor NOR2 (N455, N454, N309);
not NOT1 (N456, N453);
and AND3 (N457, N451, N281, N358);
nand NAND3 (N458, N430, N183, N418);
buf BUF1 (N459, N455);
and AND4 (N460, N458, N313, N39, N327);
xor XOR2 (N461, N446, N247);
buf BUF1 (N462, N439);
not NOT1 (N463, N459);
nand NAND2 (N464, N419, N372);
not NOT1 (N465, N461);
and AND3 (N466, N442, N258, N454);
nand NAND2 (N467, N462, N11);
not NOT1 (N468, N457);
buf BUF1 (N469, N463);
nor NOR3 (N470, N464, N339, N53);
xor XOR2 (N471, N460, N7);
nor NOR2 (N472, N469, N198);
buf BUF1 (N473, N452);
buf BUF1 (N474, N472);
buf BUF1 (N475, N474);
not NOT1 (N476, N475);
buf BUF1 (N477, N470);
nor NOR4 (N478, N471, N302, N153, N360);
buf BUF1 (N479, N478);
nor NOR2 (N480, N479, N442);
xor XOR2 (N481, N476, N445);
not NOT1 (N482, N456);
and AND4 (N483, N450, N458, N317, N197);
or OR3 (N484, N467, N146, N429);
nand NAND4 (N485, N473, N148, N456, N140);
xor XOR2 (N486, N483, N36);
xor XOR2 (N487, N486, N455);
buf BUF1 (N488, N465);
buf BUF1 (N489, N481);
nand NAND4 (N490, N487, N221, N300, N200);
nand NAND2 (N491, N477, N461);
or OR3 (N492, N488, N458, N402);
not NOT1 (N493, N482);
nand NAND3 (N494, N485, N241, N67);
not NOT1 (N495, N490);
not NOT1 (N496, N495);
or OR4 (N497, N494, N407, N227, N342);
nor NOR4 (N498, N496, N497, N7, N309);
not NOT1 (N499, N177);
nor NOR3 (N500, N466, N407, N422);
buf BUF1 (N501, N484);
buf BUF1 (N502, N489);
nand NAND4 (N503, N502, N74, N60, N316);
and AND4 (N504, N500, N325, N130, N121);
or OR4 (N505, N504, N394, N485, N395);
and AND4 (N506, N493, N204, N41, N489);
xor XOR2 (N507, N501, N11);
not NOT1 (N508, N468);
not NOT1 (N509, N506);
xor XOR2 (N510, N499, N24);
buf BUF1 (N511, N505);
nand NAND4 (N512, N510, N289, N220, N202);
buf BUF1 (N513, N512);
or OR4 (N514, N513, N239, N216, N248);
or OR3 (N515, N498, N457, N86);
buf BUF1 (N516, N514);
and AND2 (N517, N503, N152);
nor NOR4 (N518, N480, N412, N301, N511);
nor NOR3 (N519, N159, N517, N247);
buf BUF1 (N520, N500);
and AND4 (N521, N518, N387, N448, N99);
not NOT1 (N522, N507);
nor NOR3 (N523, N508, N258, N288);
nor NOR4 (N524, N520, N329, N312, N14);
nand NAND3 (N525, N519, N240, N74);
nand NAND4 (N526, N516, N398, N299, N338);
buf BUF1 (N527, N509);
and AND3 (N528, N521, N177, N366);
nor NOR3 (N529, N525, N76, N395);
and AND4 (N530, N524, N303, N48, N503);
nand NAND4 (N531, N522, N297, N307, N489);
nand NAND3 (N532, N529, N174, N388);
and AND3 (N533, N532, N428, N10);
not NOT1 (N534, N531);
not NOT1 (N535, N534);
xor XOR2 (N536, N535, N430);
buf BUF1 (N537, N491);
nand NAND2 (N538, N527, N268);
not NOT1 (N539, N528);
buf BUF1 (N540, N523);
nor NOR2 (N541, N533, N442);
nand NAND4 (N542, N526, N216, N478, N538);
and AND3 (N543, N302, N122, N165);
nor NOR4 (N544, N515, N204, N303, N259);
and AND4 (N545, N492, N68, N76, N290);
xor XOR2 (N546, N545, N432);
buf BUF1 (N547, N539);
xor XOR2 (N548, N544, N388);
and AND4 (N549, N536, N410, N472, N233);
and AND3 (N550, N541, N445, N11);
and AND4 (N551, N550, N54, N212, N351);
and AND4 (N552, N542, N313, N71, N292);
nor NOR2 (N553, N546, N292);
not NOT1 (N554, N549);
nand NAND2 (N555, N537, N323);
xor XOR2 (N556, N551, N217);
nand NAND3 (N557, N547, N41, N261);
and AND3 (N558, N543, N552, N80);
not NOT1 (N559, N515);
xor XOR2 (N560, N558, N470);
buf BUF1 (N561, N540);
and AND3 (N562, N554, N467, N340);
nand NAND4 (N563, N562, N375, N190, N544);
nand NAND2 (N564, N530, N26);
not NOT1 (N565, N560);
or OR3 (N566, N555, N112, N498);
and AND3 (N567, N563, N176, N508);
buf BUF1 (N568, N565);
xor XOR2 (N569, N566, N138);
nand NAND2 (N570, N567, N308);
nand NAND2 (N571, N553, N224);
xor XOR2 (N572, N564, N14);
not NOT1 (N573, N556);
buf BUF1 (N574, N569);
xor XOR2 (N575, N548, N153);
nand NAND2 (N576, N568, N31);
or OR2 (N577, N557, N112);
not NOT1 (N578, N576);
buf BUF1 (N579, N574);
buf BUF1 (N580, N577);
xor XOR2 (N581, N570, N264);
not NOT1 (N582, N581);
buf BUF1 (N583, N578);
nor NOR3 (N584, N572, N228, N108);
xor XOR2 (N585, N584, N427);
buf BUF1 (N586, N585);
xor XOR2 (N587, N579, N575);
and AND4 (N588, N383, N11, N354, N72);
not NOT1 (N589, N588);
nor NOR3 (N590, N559, N455, N109);
and AND3 (N591, N571, N127, N296);
xor XOR2 (N592, N580, N397);
nand NAND4 (N593, N583, N312, N469, N219);
nand NAND4 (N594, N593, N17, N545, N560);
not NOT1 (N595, N561);
buf BUF1 (N596, N589);
not NOT1 (N597, N591);
nor NOR3 (N598, N582, N242, N529);
not NOT1 (N599, N594);
nand NAND4 (N600, N586, N314, N185, N581);
not NOT1 (N601, N596);
and AND4 (N602, N595, N454, N310, N79);
xor XOR2 (N603, N587, N196);
not NOT1 (N604, N598);
and AND2 (N605, N602, N338);
or OR2 (N606, N573, N151);
or OR2 (N607, N605, N497);
nand NAND2 (N608, N599, N555);
xor XOR2 (N609, N601, N334);
nand NAND2 (N610, N600, N544);
xor XOR2 (N611, N604, N527);
nand NAND2 (N612, N608, N38);
or OR2 (N613, N606, N106);
buf BUF1 (N614, N607);
nor NOR2 (N615, N614, N269);
buf BUF1 (N616, N613);
not NOT1 (N617, N615);
or OR2 (N618, N611, N374);
buf BUF1 (N619, N597);
nor NOR3 (N620, N617, N584, N460);
nor NOR4 (N621, N592, N147, N588, N509);
not NOT1 (N622, N621);
and AND3 (N623, N603, N301, N326);
nand NAND3 (N624, N610, N150, N446);
and AND4 (N625, N620, N588, N217, N482);
buf BUF1 (N626, N623);
and AND4 (N627, N622, N170, N182, N452);
not NOT1 (N628, N618);
and AND4 (N629, N609, N374, N533, N208);
and AND2 (N630, N628, N55);
not NOT1 (N631, N629);
buf BUF1 (N632, N612);
not NOT1 (N633, N627);
nand NAND2 (N634, N625, N117);
buf BUF1 (N635, N632);
nor NOR3 (N636, N633, N522, N216);
not NOT1 (N637, N636);
buf BUF1 (N638, N635);
and AND2 (N639, N619, N197);
not NOT1 (N640, N624);
buf BUF1 (N641, N616);
and AND3 (N642, N631, N382, N91);
nand NAND4 (N643, N637, N563, N553, N549);
nor NOR4 (N644, N634, N271, N450, N60);
not NOT1 (N645, N640);
xor XOR2 (N646, N643, N621);
not NOT1 (N647, N630);
nand NAND2 (N648, N647, N399);
nand NAND2 (N649, N648, N590);
not NOT1 (N650, N238);
not NOT1 (N651, N650);
nor NOR2 (N652, N639, N244);
xor XOR2 (N653, N646, N636);
not NOT1 (N654, N651);
buf BUF1 (N655, N654);
not NOT1 (N656, N645);
not NOT1 (N657, N642);
and AND4 (N658, N653, N601, N37, N459);
xor XOR2 (N659, N641, N78);
nand NAND4 (N660, N658, N544, N235, N52);
not NOT1 (N661, N644);
xor XOR2 (N662, N656, N30);
not NOT1 (N663, N652);
buf BUF1 (N664, N659);
not NOT1 (N665, N655);
buf BUF1 (N666, N664);
nor NOR2 (N667, N638, N203);
nand NAND4 (N668, N657, N512, N306, N372);
nor NOR3 (N669, N665, N393, N13);
or OR2 (N670, N649, N302);
xor XOR2 (N671, N667, N592);
or OR2 (N672, N662, N492);
or OR2 (N673, N626, N76);
not NOT1 (N674, N670);
not NOT1 (N675, N661);
nor NOR2 (N676, N663, N513);
nor NOR3 (N677, N673, N267, N54);
and AND3 (N678, N677, N605, N221);
and AND2 (N679, N672, N53);
buf BUF1 (N680, N668);
or OR3 (N681, N676, N312, N247);
not NOT1 (N682, N678);
or OR2 (N683, N682, N40);
buf BUF1 (N684, N669);
xor XOR2 (N685, N684, N293);
nor NOR3 (N686, N666, N399, N228);
not NOT1 (N687, N675);
xor XOR2 (N688, N671, N338);
or OR4 (N689, N680, N456, N386, N455);
buf BUF1 (N690, N686);
not NOT1 (N691, N688);
not NOT1 (N692, N691);
xor XOR2 (N693, N681, N87);
not NOT1 (N694, N683);
or OR2 (N695, N685, N691);
and AND4 (N696, N692, N445, N430, N173);
nand NAND4 (N697, N695, N89, N63, N73);
not NOT1 (N698, N693);
and AND2 (N699, N694, N518);
buf BUF1 (N700, N687);
xor XOR2 (N701, N696, N355);
or OR4 (N702, N689, N554, N96, N285);
nand NAND2 (N703, N697, N662);
or OR2 (N704, N674, N78);
nand NAND3 (N705, N690, N198, N484);
nor NOR3 (N706, N705, N127, N413);
nand NAND4 (N707, N660, N430, N470, N668);
nand NAND4 (N708, N706, N12, N677, N153);
nor NOR3 (N709, N679, N263, N255);
and AND2 (N710, N699, N606);
xor XOR2 (N711, N710, N504);
buf BUF1 (N712, N711);
not NOT1 (N713, N704);
nor NOR3 (N714, N700, N60, N73);
nand NAND3 (N715, N703, N189, N365);
or OR2 (N716, N708, N690);
not NOT1 (N717, N716);
nor NOR4 (N718, N717, N556, N376, N596);
nor NOR4 (N719, N698, N320, N431, N487);
and AND4 (N720, N707, N270, N546, N142);
or OR2 (N721, N719, N256);
xor XOR2 (N722, N713, N446);
not NOT1 (N723, N718);
nand NAND3 (N724, N709, N500, N599);
nand NAND3 (N725, N721, N51, N158);
buf BUF1 (N726, N720);
not NOT1 (N727, N723);
not NOT1 (N728, N725);
and AND3 (N729, N715, N328, N411);
nand NAND4 (N730, N726, N11, N591, N432);
nor NOR2 (N731, N730, N587);
not NOT1 (N732, N722);
nand NAND2 (N733, N727, N91);
and AND3 (N734, N729, N546, N595);
not NOT1 (N735, N714);
nand NAND2 (N736, N732, N369);
nand NAND4 (N737, N728, N383, N583, N518);
or OR2 (N738, N734, N655);
not NOT1 (N739, N736);
xor XOR2 (N740, N724, N4);
or OR4 (N741, N740, N571, N298, N416);
nor NOR2 (N742, N733, N571);
and AND4 (N743, N735, N559, N509, N248);
buf BUF1 (N744, N742);
buf BUF1 (N745, N741);
nor NOR4 (N746, N701, N467, N104, N344);
and AND3 (N747, N739, N585, N18);
buf BUF1 (N748, N745);
and AND4 (N749, N731, N746, N186, N16);
xor XOR2 (N750, N118, N164);
not NOT1 (N751, N738);
buf BUF1 (N752, N748);
and AND4 (N753, N702, N301, N660, N460);
not NOT1 (N754, N743);
buf BUF1 (N755, N749);
buf BUF1 (N756, N753);
xor XOR2 (N757, N754, N448);
not NOT1 (N758, N744);
not NOT1 (N759, N747);
or OR2 (N760, N757, N7);
and AND3 (N761, N758, N678, N588);
or OR2 (N762, N760, N17);
nor NOR3 (N763, N712, N224, N144);
and AND4 (N764, N756, N369, N560, N426);
nand NAND4 (N765, N763, N230, N361, N106);
nor NOR2 (N766, N752, N212);
and AND3 (N767, N750, N328, N64);
xor XOR2 (N768, N737, N153);
xor XOR2 (N769, N761, N679);
nand NAND3 (N770, N759, N261, N163);
or OR2 (N771, N751, N13);
buf BUF1 (N772, N755);
nand NAND4 (N773, N764, N171, N432, N194);
nand NAND4 (N774, N767, N247, N526, N523);
or OR4 (N775, N774, N67, N244, N120);
nor NOR3 (N776, N769, N474, N603);
xor XOR2 (N777, N775, N504);
and AND3 (N778, N766, N498, N155);
nor NOR2 (N779, N778, N314);
nand NAND2 (N780, N770, N28);
xor XOR2 (N781, N777, N562);
nor NOR3 (N782, N776, N695, N112);
and AND3 (N783, N768, N523, N327);
and AND4 (N784, N771, N376, N585, N460);
not NOT1 (N785, N781);
not NOT1 (N786, N772);
not NOT1 (N787, N785);
or OR2 (N788, N784, N772);
or OR4 (N789, N788, N45, N336, N288);
not NOT1 (N790, N786);
nor NOR2 (N791, N783, N104);
buf BUF1 (N792, N762);
not NOT1 (N793, N773);
xor XOR2 (N794, N782, N394);
buf BUF1 (N795, N793);
and AND2 (N796, N789, N232);
xor XOR2 (N797, N787, N649);
buf BUF1 (N798, N779);
nand NAND3 (N799, N790, N713, N625);
nor NOR4 (N800, N797, N379, N291, N147);
buf BUF1 (N801, N765);
buf BUF1 (N802, N780);
xor XOR2 (N803, N796, N204);
not NOT1 (N804, N803);
and AND2 (N805, N792, N71);
nor NOR4 (N806, N795, N709, N757, N274);
and AND4 (N807, N802, N691, N509, N344);
buf BUF1 (N808, N794);
buf BUF1 (N809, N807);
or OR4 (N810, N809, N200, N338, N215);
or OR4 (N811, N805, N489, N532, N194);
nand NAND2 (N812, N791, N229);
not NOT1 (N813, N808);
or OR3 (N814, N813, N743, N588);
not NOT1 (N815, N801);
xor XOR2 (N816, N815, N359);
nand NAND3 (N817, N799, N392, N155);
or OR2 (N818, N817, N704);
or OR3 (N819, N814, N436, N248);
buf BUF1 (N820, N800);
nor NOR3 (N821, N812, N719, N517);
or OR4 (N822, N818, N271, N495, N294);
xor XOR2 (N823, N806, N558);
buf BUF1 (N824, N816);
xor XOR2 (N825, N821, N577);
buf BUF1 (N826, N819);
or OR4 (N827, N823, N244, N688, N643);
nand NAND4 (N828, N825, N12, N615, N683);
nor NOR2 (N829, N822, N623);
or OR2 (N830, N824, N642);
nor NOR3 (N831, N804, N790, N261);
buf BUF1 (N832, N820);
and AND4 (N833, N798, N323, N33, N759);
or OR4 (N834, N830, N756, N329, N147);
and AND2 (N835, N827, N443);
nor NOR3 (N836, N828, N602, N510);
nand NAND4 (N837, N833, N320, N103, N481);
not NOT1 (N838, N810);
xor XOR2 (N839, N837, N381);
nand NAND4 (N840, N811, N514, N252, N404);
and AND4 (N841, N838, N294, N135, N89);
or OR2 (N842, N836, N804);
buf BUF1 (N843, N839);
nand NAND4 (N844, N843, N112, N743, N63);
nand NAND2 (N845, N826, N246);
or OR4 (N846, N834, N262, N321, N618);
nand NAND3 (N847, N829, N809, N331);
nand NAND4 (N848, N847, N59, N793, N770);
xor XOR2 (N849, N832, N470);
not NOT1 (N850, N831);
buf BUF1 (N851, N846);
not NOT1 (N852, N850);
and AND4 (N853, N845, N404, N673, N442);
buf BUF1 (N854, N848);
nor NOR3 (N855, N844, N221, N542);
nor NOR4 (N856, N854, N116, N197, N52);
not NOT1 (N857, N853);
buf BUF1 (N858, N851);
or OR3 (N859, N856, N406, N439);
or OR2 (N860, N842, N220);
nor NOR2 (N861, N857, N128);
and AND3 (N862, N855, N455, N128);
nand NAND2 (N863, N852, N41);
nand NAND2 (N864, N861, N38);
buf BUF1 (N865, N858);
nand NAND2 (N866, N864, N501);
xor XOR2 (N867, N859, N418);
not NOT1 (N868, N866);
buf BUF1 (N869, N849);
and AND2 (N870, N869, N560);
not NOT1 (N871, N841);
or OR4 (N872, N835, N510, N68, N368);
nor NOR2 (N873, N870, N286);
buf BUF1 (N874, N860);
not NOT1 (N875, N872);
buf BUF1 (N876, N862);
and AND4 (N877, N840, N201, N225, N571);
nor NOR3 (N878, N874, N102, N279);
xor XOR2 (N879, N871, N723);
not NOT1 (N880, N876);
nand NAND4 (N881, N877, N631, N876, N232);
buf BUF1 (N882, N868);
xor XOR2 (N883, N875, N369);
nand NAND2 (N884, N863, N407);
nor NOR4 (N885, N865, N463, N655, N390);
nor NOR2 (N886, N873, N609);
buf BUF1 (N887, N879);
not NOT1 (N888, N867);
or OR4 (N889, N886, N451, N141, N537);
or OR3 (N890, N885, N694, N379);
not NOT1 (N891, N890);
or OR3 (N892, N880, N756, N562);
not NOT1 (N893, N887);
xor XOR2 (N894, N893, N52);
buf BUF1 (N895, N894);
xor XOR2 (N896, N888, N888);
nand NAND3 (N897, N884, N145, N93);
not NOT1 (N898, N897);
not NOT1 (N899, N883);
or OR2 (N900, N892, N722);
nor NOR2 (N901, N878, N742);
xor XOR2 (N902, N891, N80);
and AND4 (N903, N899, N399, N605, N759);
nand NAND4 (N904, N896, N369, N674, N717);
or OR2 (N905, N895, N483);
nor NOR3 (N906, N903, N755, N898);
nor NOR4 (N907, N222, N888, N801, N804);
xor XOR2 (N908, N881, N121);
nand NAND2 (N909, N906, N798);
nor NOR3 (N910, N905, N620, N662);
not NOT1 (N911, N901);
not NOT1 (N912, N909);
not NOT1 (N913, N912);
nor NOR4 (N914, N913, N870, N583, N439);
or OR2 (N915, N904, N614);
nor NOR4 (N916, N908, N857, N52, N173);
nor NOR3 (N917, N915, N827, N56);
not NOT1 (N918, N917);
nor NOR3 (N919, N900, N391, N716);
nand NAND4 (N920, N918, N179, N168, N444);
xor XOR2 (N921, N902, N643);
buf BUF1 (N922, N889);
nand NAND3 (N923, N920, N349, N815);
and AND4 (N924, N921, N645, N225, N280);
nor NOR3 (N925, N914, N805, N538);
nor NOR3 (N926, N916, N736, N188);
or OR2 (N927, N910, N727);
or OR3 (N928, N927, N339, N503);
nor NOR3 (N929, N926, N567, N663);
and AND4 (N930, N929, N1, N43, N416);
xor XOR2 (N931, N930, N495);
buf BUF1 (N932, N922);
buf BUF1 (N933, N919);
buf BUF1 (N934, N911);
or OR2 (N935, N907, N308);
or OR4 (N936, N925, N269, N548, N166);
xor XOR2 (N937, N931, N203);
xor XOR2 (N938, N935, N482);
xor XOR2 (N939, N924, N578);
and AND2 (N940, N928, N453);
xor XOR2 (N941, N923, N360);
or OR2 (N942, N939, N223);
xor XOR2 (N943, N941, N416);
nor NOR2 (N944, N932, N110);
nor NOR4 (N945, N938, N604, N701, N880);
nand NAND3 (N946, N936, N739, N452);
nor NOR3 (N947, N934, N809, N6);
not NOT1 (N948, N945);
and AND3 (N949, N946, N195, N17);
and AND2 (N950, N933, N831);
nand NAND4 (N951, N949, N348, N204, N681);
nor NOR2 (N952, N944, N538);
or OR3 (N953, N951, N684, N193);
or OR3 (N954, N948, N230, N826);
nand NAND2 (N955, N882, N847);
nor NOR4 (N956, N947, N927, N24, N302);
and AND4 (N957, N953, N606, N636, N633);
and AND2 (N958, N937, N571);
nor NOR3 (N959, N942, N236, N912);
nor NOR2 (N960, N956, N721);
and AND4 (N961, N957, N718, N375, N675);
or OR2 (N962, N959, N598);
xor XOR2 (N963, N961, N131);
xor XOR2 (N964, N963, N496);
and AND4 (N965, N943, N100, N964, N696);
buf BUF1 (N966, N961);
xor XOR2 (N967, N966, N341);
not NOT1 (N968, N960);
nor NOR4 (N969, N940, N474, N637, N492);
and AND4 (N970, N965, N249, N271, N573);
or OR3 (N971, N969, N394, N635);
nand NAND3 (N972, N955, N902, N258);
buf BUF1 (N973, N962);
nand NAND3 (N974, N958, N429, N179);
nand NAND4 (N975, N967, N654, N810, N824);
not NOT1 (N976, N950);
buf BUF1 (N977, N971);
nand NAND3 (N978, N975, N875, N792);
not NOT1 (N979, N974);
xor XOR2 (N980, N968, N585);
nand NAND4 (N981, N954, N673, N522, N940);
not NOT1 (N982, N972);
buf BUF1 (N983, N981);
not NOT1 (N984, N980);
nor NOR4 (N985, N983, N692, N426, N512);
and AND3 (N986, N984, N580, N376);
xor XOR2 (N987, N976, N798);
not NOT1 (N988, N979);
buf BUF1 (N989, N978);
and AND2 (N990, N977, N406);
not NOT1 (N991, N986);
or OR2 (N992, N982, N149);
and AND4 (N993, N990, N308, N235, N54);
nand NAND4 (N994, N952, N126, N516, N32);
and AND3 (N995, N970, N383, N759);
nand NAND3 (N996, N988, N859, N833);
xor XOR2 (N997, N996, N372);
xor XOR2 (N998, N992, N365);
buf BUF1 (N999, N985);
and AND2 (N1000, N991, N49);
and AND4 (N1001, N987, N407, N685, N620);
or OR2 (N1002, N1000, N997);
buf BUF1 (N1003, N243);
not NOT1 (N1004, N999);
and AND4 (N1005, N994, N130, N804, N219);
not NOT1 (N1006, N973);
nor NOR4 (N1007, N1004, N26, N797, N324);
and AND4 (N1008, N1002, N977, N326, N791);
xor XOR2 (N1009, N995, N229);
and AND3 (N1010, N1007, N462, N895);
or OR4 (N1011, N998, N242, N256, N980);
buf BUF1 (N1012, N1005);
buf BUF1 (N1013, N1006);
not NOT1 (N1014, N993);
or OR2 (N1015, N1001, N84);
and AND3 (N1016, N1014, N77, N495);
or OR4 (N1017, N1009, N215, N102, N51);
or OR4 (N1018, N1015, N820, N121, N447);
or OR4 (N1019, N1012, N782, N511, N461);
nand NAND4 (N1020, N1016, N45, N732, N959);
not NOT1 (N1021, N1020);
buf BUF1 (N1022, N1008);
nor NOR3 (N1023, N1017, N647, N775);
xor XOR2 (N1024, N1018, N194);
not NOT1 (N1025, N1022);
or OR3 (N1026, N1003, N382, N672);
nand NAND4 (N1027, N1011, N18, N900, N447);
nor NOR2 (N1028, N1010, N219);
buf BUF1 (N1029, N1013);
xor XOR2 (N1030, N989, N914);
and AND3 (N1031, N1028, N451, N146);
nand NAND4 (N1032, N1030, N449, N771, N239);
nor NOR2 (N1033, N1024, N838);
or OR3 (N1034, N1031, N290, N501);
not NOT1 (N1035, N1033);
or OR4 (N1036, N1021, N780, N585, N298);
nand NAND3 (N1037, N1036, N599, N6);
nor NOR2 (N1038, N1025, N810);
xor XOR2 (N1039, N1019, N545);
and AND3 (N1040, N1023, N495, N497);
and AND3 (N1041, N1040, N809, N276);
or OR2 (N1042, N1041, N178);
and AND4 (N1043, N1026, N774, N1027, N625);
nand NAND4 (N1044, N192, N839, N264, N411);
nand NAND2 (N1045, N1044, N590);
and AND2 (N1046, N1032, N921);
or OR2 (N1047, N1042, N745);
buf BUF1 (N1048, N1029);
not NOT1 (N1049, N1038);
nor NOR4 (N1050, N1048, N302, N486, N579);
and AND3 (N1051, N1050, N27, N369);
xor XOR2 (N1052, N1039, N343);
nor NOR3 (N1053, N1047, N749, N1045);
buf BUF1 (N1054, N1009);
not NOT1 (N1055, N1051);
buf BUF1 (N1056, N1055);
buf BUF1 (N1057, N1052);
xor XOR2 (N1058, N1056, N655);
buf BUF1 (N1059, N1034);
buf BUF1 (N1060, N1054);
nand NAND2 (N1061, N1058, N286);
or OR3 (N1062, N1049, N467, N990);
and AND2 (N1063, N1037, N440);
xor XOR2 (N1064, N1053, N15);
nand NAND2 (N1065, N1043, N238);
xor XOR2 (N1066, N1064, N268);
not NOT1 (N1067, N1062);
buf BUF1 (N1068, N1067);
buf BUF1 (N1069, N1035);
nand NAND2 (N1070, N1069, N927);
nand NAND2 (N1071, N1061, N241);
xor XOR2 (N1072, N1068, N43);
nor NOR2 (N1073, N1057, N85);
not NOT1 (N1074, N1063);
buf BUF1 (N1075, N1070);
or OR4 (N1076, N1075, N615, N1016, N263);
xor XOR2 (N1077, N1076, N683);
nand NAND4 (N1078, N1065, N416, N170, N139);
not NOT1 (N1079, N1074);
xor XOR2 (N1080, N1072, N261);
not NOT1 (N1081, N1073);
buf BUF1 (N1082, N1046);
nand NAND2 (N1083, N1080, N437);
xor XOR2 (N1084, N1060, N42);
and AND3 (N1085, N1077, N548, N687);
and AND4 (N1086, N1084, N955, N692, N788);
nand NAND2 (N1087, N1086, N804);
not NOT1 (N1088, N1087);
nor NOR4 (N1089, N1079, N19, N854, N872);
or OR2 (N1090, N1082, N823);
xor XOR2 (N1091, N1078, N140);
xor XOR2 (N1092, N1059, N9);
and AND4 (N1093, N1083, N34, N587, N826);
not NOT1 (N1094, N1066);
xor XOR2 (N1095, N1094, N988);
not NOT1 (N1096, N1071);
or OR2 (N1097, N1090, N176);
xor XOR2 (N1098, N1091, N125);
nor NOR4 (N1099, N1089, N524, N923, N561);
nand NAND4 (N1100, N1088, N141, N146, N474);
nand NAND4 (N1101, N1097, N927, N26, N727);
nor NOR4 (N1102, N1093, N466, N1004, N965);
and AND2 (N1103, N1081, N27);
not NOT1 (N1104, N1095);
nand NAND2 (N1105, N1092, N566);
or OR4 (N1106, N1085, N941, N342, N897);
and AND3 (N1107, N1103, N393, N896);
xor XOR2 (N1108, N1106, N881);
buf BUF1 (N1109, N1096);
buf BUF1 (N1110, N1099);
nand NAND4 (N1111, N1107, N217, N862, N791);
or OR4 (N1112, N1108, N267, N989, N608);
not NOT1 (N1113, N1109);
and AND2 (N1114, N1100, N945);
nand NAND4 (N1115, N1104, N673, N220, N660);
xor XOR2 (N1116, N1113, N1069);
nor NOR3 (N1117, N1111, N88, N1023);
and AND3 (N1118, N1105, N155, N296);
and AND3 (N1119, N1118, N766, N52);
or OR2 (N1120, N1101, N276);
not NOT1 (N1121, N1102);
nand NAND4 (N1122, N1098, N12, N1107, N7);
nor NOR2 (N1123, N1114, N698);
nor NOR2 (N1124, N1116, N764);
nor NOR2 (N1125, N1121, N274);
nand NAND3 (N1126, N1117, N651, N921);
buf BUF1 (N1127, N1125);
nor NOR4 (N1128, N1112, N533, N187, N939);
nor NOR3 (N1129, N1120, N533, N526);
or OR3 (N1130, N1126, N621, N826);
or OR2 (N1131, N1123, N635);
or OR3 (N1132, N1115, N609, N635);
nor NOR2 (N1133, N1127, N636);
or OR4 (N1134, N1130, N799, N283, N878);
or OR2 (N1135, N1128, N1079);
nand NAND3 (N1136, N1135, N913, N630);
nor NOR3 (N1137, N1129, N164, N1127);
nand NAND4 (N1138, N1131, N319, N1077, N1006);
or OR3 (N1139, N1138, N426, N350);
nand NAND3 (N1140, N1133, N235, N421);
nor NOR2 (N1141, N1134, N414);
xor XOR2 (N1142, N1141, N246);
not NOT1 (N1143, N1142);
buf BUF1 (N1144, N1139);
nor NOR4 (N1145, N1124, N1112, N668, N755);
not NOT1 (N1146, N1137);
not NOT1 (N1147, N1119);
nor NOR3 (N1148, N1146, N304, N100);
buf BUF1 (N1149, N1147);
and AND4 (N1150, N1122, N508, N476, N179);
nand NAND3 (N1151, N1143, N455, N199);
nor NOR4 (N1152, N1149, N111, N363, N703);
nand NAND3 (N1153, N1140, N1054, N767);
not NOT1 (N1154, N1110);
and AND4 (N1155, N1153, N493, N480, N707);
or OR3 (N1156, N1136, N1099, N849);
or OR3 (N1157, N1154, N304, N225);
and AND3 (N1158, N1156, N494, N75);
and AND3 (N1159, N1152, N1089, N238);
xor XOR2 (N1160, N1145, N573);
xor XOR2 (N1161, N1160, N318);
and AND2 (N1162, N1150, N575);
buf BUF1 (N1163, N1159);
not NOT1 (N1164, N1132);
nor NOR4 (N1165, N1162, N775, N473, N688);
nor NOR4 (N1166, N1155, N814, N834, N483);
not NOT1 (N1167, N1158);
buf BUF1 (N1168, N1167);
buf BUF1 (N1169, N1148);
nand NAND4 (N1170, N1157, N419, N1103, N1024);
nand NAND2 (N1171, N1164, N984);
and AND4 (N1172, N1169, N372, N427, N537);
buf BUF1 (N1173, N1166);
and AND4 (N1174, N1168, N749, N27, N820);
nor NOR3 (N1175, N1151, N232, N829);
buf BUF1 (N1176, N1170);
nand NAND4 (N1177, N1171, N956, N67, N714);
and AND4 (N1178, N1177, N619, N1031, N176);
nand NAND2 (N1179, N1174, N1106);
and AND4 (N1180, N1144, N1017, N488, N1117);
or OR2 (N1181, N1175, N844);
not NOT1 (N1182, N1161);
nand NAND2 (N1183, N1181, N260);
xor XOR2 (N1184, N1183, N346);
nor NOR2 (N1185, N1180, N639);
or OR3 (N1186, N1185, N759, N1009);
not NOT1 (N1187, N1178);
nor NOR2 (N1188, N1173, N311);
and AND2 (N1189, N1179, N198);
or OR4 (N1190, N1172, N704, N1123, N429);
nor NOR3 (N1191, N1189, N26, N333);
or OR3 (N1192, N1182, N398, N1099);
nand NAND4 (N1193, N1188, N828, N675, N1107);
nor NOR3 (N1194, N1186, N953, N398);
nor NOR4 (N1195, N1184, N1015, N396, N1141);
or OR3 (N1196, N1191, N300, N1039);
nand NAND4 (N1197, N1165, N842, N1158, N1073);
buf BUF1 (N1198, N1194);
xor XOR2 (N1199, N1187, N383);
nor NOR2 (N1200, N1198, N1108);
nand NAND3 (N1201, N1195, N1006, N335);
or OR4 (N1202, N1201, N726, N1164, N658);
buf BUF1 (N1203, N1202);
nor NOR3 (N1204, N1196, N1201, N932);
xor XOR2 (N1205, N1190, N688);
or OR2 (N1206, N1204, N36);
not NOT1 (N1207, N1203);
xor XOR2 (N1208, N1207, N1100);
buf BUF1 (N1209, N1200);
or OR2 (N1210, N1197, N389);
nor NOR2 (N1211, N1176, N534);
buf BUF1 (N1212, N1163);
or OR2 (N1213, N1212, N889);
not NOT1 (N1214, N1192);
and AND3 (N1215, N1208, N954, N1204);
xor XOR2 (N1216, N1214, N382);
nand NAND2 (N1217, N1213, N319);
buf BUF1 (N1218, N1215);
nand NAND4 (N1219, N1199, N929, N117, N303);
and AND3 (N1220, N1206, N572, N10);
and AND2 (N1221, N1217, N205);
buf BUF1 (N1222, N1193);
nor NOR2 (N1223, N1218, N409);
xor XOR2 (N1224, N1211, N909);
nor NOR2 (N1225, N1223, N768);
xor XOR2 (N1226, N1225, N1122);
xor XOR2 (N1227, N1222, N957);
or OR3 (N1228, N1227, N910, N1008);
xor XOR2 (N1229, N1221, N491);
nor NOR4 (N1230, N1216, N204, N482, N942);
xor XOR2 (N1231, N1228, N260);
xor XOR2 (N1232, N1229, N396);
buf BUF1 (N1233, N1231);
or OR4 (N1234, N1224, N441, N389, N824);
or OR2 (N1235, N1226, N70);
and AND2 (N1236, N1230, N350);
not NOT1 (N1237, N1209);
and AND4 (N1238, N1210, N1171, N927, N593);
nor NOR2 (N1239, N1234, N317);
nand NAND4 (N1240, N1239, N251, N267, N411);
xor XOR2 (N1241, N1238, N1058);
nand NAND2 (N1242, N1237, N364);
buf BUF1 (N1243, N1220);
buf BUF1 (N1244, N1232);
nand NAND2 (N1245, N1235, N13);
and AND2 (N1246, N1233, N882);
buf BUF1 (N1247, N1245);
xor XOR2 (N1248, N1246, N875);
xor XOR2 (N1249, N1248, N972);
nand NAND2 (N1250, N1242, N282);
buf BUF1 (N1251, N1236);
nor NOR4 (N1252, N1250, N207, N13, N144);
and AND4 (N1253, N1240, N116, N314, N298);
xor XOR2 (N1254, N1205, N30);
not NOT1 (N1255, N1251);
not NOT1 (N1256, N1253);
and AND2 (N1257, N1219, N826);
nand NAND2 (N1258, N1255, N296);
xor XOR2 (N1259, N1254, N707);
or OR3 (N1260, N1257, N460, N426);
nand NAND4 (N1261, N1243, N635, N903, N1013);
nand NAND2 (N1262, N1249, N495);
xor XOR2 (N1263, N1252, N93);
xor XOR2 (N1264, N1244, N1189);
not NOT1 (N1265, N1256);
or OR4 (N1266, N1262, N726, N380, N42);
nand NAND4 (N1267, N1259, N414, N233, N925);
buf BUF1 (N1268, N1247);
nand NAND2 (N1269, N1265, N751);
xor XOR2 (N1270, N1260, N403);
buf BUF1 (N1271, N1264);
not NOT1 (N1272, N1263);
xor XOR2 (N1273, N1241, N782);
xor XOR2 (N1274, N1266, N550);
nand NAND3 (N1275, N1261, N435, N682);
not NOT1 (N1276, N1271);
and AND4 (N1277, N1269, N798, N522, N339);
xor XOR2 (N1278, N1273, N856);
nor NOR2 (N1279, N1274, N180);
xor XOR2 (N1280, N1277, N496);
buf BUF1 (N1281, N1267);
or OR2 (N1282, N1270, N598);
xor XOR2 (N1283, N1282, N768);
xor XOR2 (N1284, N1276, N214);
buf BUF1 (N1285, N1268);
buf BUF1 (N1286, N1275);
not NOT1 (N1287, N1280);
buf BUF1 (N1288, N1283);
and AND3 (N1289, N1279, N1075, N516);
nor NOR3 (N1290, N1285, N179, N1139);
nand NAND3 (N1291, N1281, N1030, N1138);
and AND2 (N1292, N1272, N910);
buf BUF1 (N1293, N1292);
nor NOR3 (N1294, N1258, N738, N1278);
buf BUF1 (N1295, N1153);
xor XOR2 (N1296, N1288, N299);
nand NAND3 (N1297, N1295, N978, N1006);
not NOT1 (N1298, N1290);
and AND4 (N1299, N1284, N220, N629, N113);
and AND2 (N1300, N1294, N575);
nand NAND4 (N1301, N1291, N151, N326, N514);
not NOT1 (N1302, N1296);
xor XOR2 (N1303, N1302, N1150);
and AND2 (N1304, N1293, N1101);
xor XOR2 (N1305, N1298, N583);
not NOT1 (N1306, N1289);
or OR2 (N1307, N1297, N578);
or OR3 (N1308, N1305, N714, N518);
and AND2 (N1309, N1287, N154);
not NOT1 (N1310, N1303);
xor XOR2 (N1311, N1308, N1000);
and AND4 (N1312, N1299, N670, N73, N312);
and AND4 (N1313, N1310, N910, N1194, N478);
xor XOR2 (N1314, N1311, N811);
and AND2 (N1315, N1307, N129);
xor XOR2 (N1316, N1313, N1133);
buf BUF1 (N1317, N1315);
and AND3 (N1318, N1309, N194, N307);
buf BUF1 (N1319, N1317);
and AND3 (N1320, N1300, N1082, N305);
not NOT1 (N1321, N1286);
or OR4 (N1322, N1321, N1098, N160, N885);
not NOT1 (N1323, N1316);
or OR4 (N1324, N1323, N822, N672, N233);
buf BUF1 (N1325, N1314);
buf BUF1 (N1326, N1325);
not NOT1 (N1327, N1319);
and AND2 (N1328, N1320, N19);
or OR2 (N1329, N1312, N1110);
not NOT1 (N1330, N1306);
or OR4 (N1331, N1304, N408, N1136, N218);
nand NAND4 (N1332, N1301, N1306, N1157, N568);
not NOT1 (N1333, N1329);
nand NAND3 (N1334, N1326, N946, N703);
and AND3 (N1335, N1334, N367, N584);
not NOT1 (N1336, N1328);
or OR3 (N1337, N1331, N189, N1101);
or OR2 (N1338, N1330, N339);
not NOT1 (N1339, N1322);
nand NAND2 (N1340, N1335, N456);
nor NOR3 (N1341, N1332, N398, N443);
buf BUF1 (N1342, N1339);
xor XOR2 (N1343, N1333, N124);
or OR4 (N1344, N1340, N1241, N907, N1258);
not NOT1 (N1345, N1324);
buf BUF1 (N1346, N1345);
or OR4 (N1347, N1337, N885, N1139, N39);
nor NOR3 (N1348, N1344, N126, N455);
nor NOR4 (N1349, N1348, N962, N566, N220);
not NOT1 (N1350, N1327);
and AND3 (N1351, N1341, N184, N360);
and AND3 (N1352, N1318, N240, N282);
not NOT1 (N1353, N1352);
nor NOR2 (N1354, N1346, N1261);
nand NAND3 (N1355, N1351, N641, N625);
nor NOR3 (N1356, N1342, N1345, N201);
buf BUF1 (N1357, N1349);
or OR3 (N1358, N1347, N826, N895);
not NOT1 (N1359, N1358);
or OR2 (N1360, N1356, N451);
buf BUF1 (N1361, N1359);
buf BUF1 (N1362, N1343);
nor NOR4 (N1363, N1355, N745, N57, N451);
or OR4 (N1364, N1338, N1002, N1079, N597);
xor XOR2 (N1365, N1354, N140);
not NOT1 (N1366, N1363);
xor XOR2 (N1367, N1362, N103);
and AND3 (N1368, N1361, N631, N1206);
or OR2 (N1369, N1360, N1143);
nand NAND2 (N1370, N1336, N404);
buf BUF1 (N1371, N1370);
not NOT1 (N1372, N1368);
nand NAND2 (N1373, N1366, N1231);
and AND3 (N1374, N1353, N373, N1359);
not NOT1 (N1375, N1364);
nor NOR4 (N1376, N1372, N596, N104, N572);
nor NOR2 (N1377, N1369, N258);
not NOT1 (N1378, N1375);
nor NOR2 (N1379, N1367, N243);
nor NOR4 (N1380, N1350, N46, N710, N11);
and AND4 (N1381, N1371, N1017, N9, N373);
or OR2 (N1382, N1380, N12);
nor NOR3 (N1383, N1377, N142, N985);
and AND2 (N1384, N1357, N245);
nor NOR4 (N1385, N1365, N477, N788, N304);
nand NAND4 (N1386, N1378, N737, N972, N665);
xor XOR2 (N1387, N1381, N427);
xor XOR2 (N1388, N1384, N1045);
nand NAND3 (N1389, N1386, N636, N954);
not NOT1 (N1390, N1383);
nand NAND4 (N1391, N1388, N104, N306, N660);
not NOT1 (N1392, N1390);
nand NAND2 (N1393, N1379, N464);
nand NAND3 (N1394, N1391, N1177, N325);
nand NAND4 (N1395, N1373, N1027, N992, N975);
or OR2 (N1396, N1389, N841);
nand NAND3 (N1397, N1393, N136, N909);
not NOT1 (N1398, N1395);
nand NAND4 (N1399, N1396, N299, N253, N626);
buf BUF1 (N1400, N1399);
or OR2 (N1401, N1398, N1388);
buf BUF1 (N1402, N1394);
nand NAND4 (N1403, N1385, N532, N1071, N312);
nand NAND4 (N1404, N1382, N690, N1131, N444);
buf BUF1 (N1405, N1400);
nand NAND3 (N1406, N1374, N924, N937);
and AND3 (N1407, N1404, N14, N371);
nor NOR4 (N1408, N1401, N1132, N1143, N1387);
nand NAND4 (N1409, N413, N255, N713, N890);
and AND4 (N1410, N1407, N174, N51, N254);
nor NOR3 (N1411, N1376, N1316, N766);
buf BUF1 (N1412, N1405);
not NOT1 (N1413, N1408);
buf BUF1 (N1414, N1397);
nand NAND3 (N1415, N1403, N1224, N83);
nand NAND2 (N1416, N1409, N211);
nand NAND4 (N1417, N1402, N860, N216, N177);
and AND3 (N1418, N1406, N509, N554);
or OR4 (N1419, N1412, N478, N1254, N133);
not NOT1 (N1420, N1413);
nor NOR4 (N1421, N1415, N1262, N1016, N1020);
nand NAND4 (N1422, N1392, N1347, N708, N303);
buf BUF1 (N1423, N1422);
nor NOR3 (N1424, N1420, N592, N333);
not NOT1 (N1425, N1423);
or OR2 (N1426, N1419, N822);
or OR3 (N1427, N1418, N650, N1181);
and AND2 (N1428, N1416, N469);
not NOT1 (N1429, N1410);
nor NOR2 (N1430, N1427, N1138);
and AND4 (N1431, N1426, N204, N394, N828);
buf BUF1 (N1432, N1424);
nor NOR4 (N1433, N1428, N1386, N466, N413);
nor NOR3 (N1434, N1430, N258, N1340);
nor NOR2 (N1435, N1421, N1115);
nand NAND2 (N1436, N1431, N196);
and AND3 (N1437, N1432, N998, N1390);
nand NAND3 (N1438, N1435, N1190, N932);
and AND4 (N1439, N1436, N1127, N1271, N264);
nor NOR4 (N1440, N1433, N228, N734, N540);
nor NOR3 (N1441, N1434, N447, N462);
buf BUF1 (N1442, N1440);
nor NOR2 (N1443, N1441, N865);
nor NOR4 (N1444, N1443, N1400, N681, N609);
xor XOR2 (N1445, N1425, N1406);
and AND4 (N1446, N1444, N1048, N100, N55);
or OR3 (N1447, N1414, N744, N1164);
xor XOR2 (N1448, N1417, N786);
or OR3 (N1449, N1445, N623, N752);
xor XOR2 (N1450, N1442, N1381);
and AND4 (N1451, N1439, N349, N1251, N812);
and AND2 (N1452, N1450, N105);
nand NAND4 (N1453, N1451, N45, N416, N508);
nand NAND3 (N1454, N1429, N699, N292);
nor NOR3 (N1455, N1452, N1079, N803);
and AND4 (N1456, N1446, N1433, N491, N1169);
or OR3 (N1457, N1456, N54, N311);
and AND2 (N1458, N1411, N676);
not NOT1 (N1459, N1457);
buf BUF1 (N1460, N1455);
and AND4 (N1461, N1458, N1087, N1353, N1146);
not NOT1 (N1462, N1447);
nor NOR3 (N1463, N1459, N1431, N413);
buf BUF1 (N1464, N1448);
buf BUF1 (N1465, N1460);
buf BUF1 (N1466, N1449);
or OR2 (N1467, N1453, N752);
nand NAND2 (N1468, N1465, N89);
or OR2 (N1469, N1466, N40);
nand NAND2 (N1470, N1464, N1318);
not NOT1 (N1471, N1454);
nand NAND3 (N1472, N1462, N1408, N1355);
or OR3 (N1473, N1461, N1304, N1291);
nand NAND4 (N1474, N1471, N618, N1100, N621);
nor NOR3 (N1475, N1438, N310, N973);
xor XOR2 (N1476, N1472, N494);
xor XOR2 (N1477, N1437, N60);
buf BUF1 (N1478, N1476);
nor NOR4 (N1479, N1467, N78, N583, N1295);
not NOT1 (N1480, N1477);
not NOT1 (N1481, N1479);
buf BUF1 (N1482, N1481);
or OR2 (N1483, N1478, N1428);
nor NOR2 (N1484, N1463, N625);
nor NOR4 (N1485, N1475, N1114, N1047, N937);
xor XOR2 (N1486, N1485, N1132);
and AND4 (N1487, N1480, N118, N660, N189);
or OR4 (N1488, N1486, N1193, N759, N473);
nor NOR2 (N1489, N1487, N1267);
and AND4 (N1490, N1468, N1442, N485, N145);
nor NOR3 (N1491, N1488, N132, N1238);
and AND4 (N1492, N1484, N439, N1449, N55);
and AND3 (N1493, N1474, N814, N796);
not NOT1 (N1494, N1491);
buf BUF1 (N1495, N1482);
buf BUF1 (N1496, N1493);
nor NOR4 (N1497, N1469, N790, N956, N207);
not NOT1 (N1498, N1492);
nand NAND2 (N1499, N1496, N198);
nor NOR3 (N1500, N1483, N835, N630);
not NOT1 (N1501, N1500);
xor XOR2 (N1502, N1498, N958);
and AND2 (N1503, N1470, N742);
xor XOR2 (N1504, N1489, N856);
not NOT1 (N1505, N1473);
not NOT1 (N1506, N1505);
nor NOR4 (N1507, N1502, N520, N1495, N86);
xor XOR2 (N1508, N1152, N736);
nor NOR2 (N1509, N1503, N315);
and AND4 (N1510, N1499, N1496, N1477, N1163);
nand NAND2 (N1511, N1510, N1099);
and AND3 (N1512, N1501, N41, N215);
and AND4 (N1513, N1490, N2, N164, N296);
and AND3 (N1514, N1511, N231, N837);
or OR3 (N1515, N1514, N1184, N845);
and AND3 (N1516, N1507, N1134, N115);
buf BUF1 (N1517, N1515);
not NOT1 (N1518, N1512);
xor XOR2 (N1519, N1509, N1400);
xor XOR2 (N1520, N1519, N929);
nor NOR2 (N1521, N1513, N1134);
and AND2 (N1522, N1518, N935);
buf BUF1 (N1523, N1497);
xor XOR2 (N1524, N1506, N822);
or OR4 (N1525, N1521, N1443, N545, N838);
and AND2 (N1526, N1525, N369);
nand NAND3 (N1527, N1520, N34, N962);
nand NAND2 (N1528, N1523, N1231);
not NOT1 (N1529, N1526);
not NOT1 (N1530, N1528);
xor XOR2 (N1531, N1524, N238);
buf BUF1 (N1532, N1530);
nor NOR2 (N1533, N1529, N1366);
buf BUF1 (N1534, N1508);
nor NOR3 (N1535, N1522, N328, N92);
nand NAND2 (N1536, N1517, N1469);
xor XOR2 (N1537, N1536, N793);
not NOT1 (N1538, N1494);
buf BUF1 (N1539, N1534);
not NOT1 (N1540, N1527);
not NOT1 (N1541, N1535);
nor NOR2 (N1542, N1537, N1012);
nor NOR3 (N1543, N1516, N1419, N1343);
or OR2 (N1544, N1532, N214);
not NOT1 (N1545, N1541);
nand NAND4 (N1546, N1544, N1445, N19, N1466);
or OR4 (N1547, N1540, N152, N260, N618);
nor NOR4 (N1548, N1539, N1017, N864, N102);
nor NOR2 (N1549, N1543, N835);
and AND4 (N1550, N1546, N475, N1004, N248);
nor NOR3 (N1551, N1547, N686, N1384);
nand NAND3 (N1552, N1548, N238, N1217);
not NOT1 (N1553, N1531);
nor NOR3 (N1554, N1553, N225, N1444);
xor XOR2 (N1555, N1538, N1457);
xor XOR2 (N1556, N1554, N1399);
xor XOR2 (N1557, N1550, N1309);
nand NAND4 (N1558, N1556, N886, N492, N1460);
nor NOR4 (N1559, N1557, N937, N75, N8);
xor XOR2 (N1560, N1552, N332);
xor XOR2 (N1561, N1533, N534);
or OR2 (N1562, N1504, N158);
nor NOR4 (N1563, N1562, N578, N377, N927);
nand NAND2 (N1564, N1555, N1102);
and AND3 (N1565, N1542, N836, N284);
nand NAND2 (N1566, N1551, N157);
xor XOR2 (N1567, N1563, N413);
xor XOR2 (N1568, N1549, N975);
nor NOR3 (N1569, N1566, N1018, N1343);
buf BUF1 (N1570, N1560);
nor NOR3 (N1571, N1558, N576, N147);
buf BUF1 (N1572, N1565);
nand NAND4 (N1573, N1545, N1361, N666, N502);
and AND2 (N1574, N1568, N688);
not NOT1 (N1575, N1571);
not NOT1 (N1576, N1575);
nand NAND4 (N1577, N1559, N527, N323, N190);
and AND2 (N1578, N1567, N31);
nand NAND4 (N1579, N1561, N602, N610, N726);
not NOT1 (N1580, N1574);
xor XOR2 (N1581, N1578, N365);
buf BUF1 (N1582, N1579);
and AND4 (N1583, N1581, N216, N336, N931);
nand NAND2 (N1584, N1570, N1485);
xor XOR2 (N1585, N1576, N1101);
buf BUF1 (N1586, N1585);
xor XOR2 (N1587, N1584, N1362);
and AND3 (N1588, N1586, N238, N1014);
buf BUF1 (N1589, N1580);
nor NOR2 (N1590, N1569, N727);
not NOT1 (N1591, N1573);
and AND4 (N1592, N1590, N672, N1221, N1095);
and AND2 (N1593, N1589, N1364);
or OR2 (N1594, N1592, N197);
xor XOR2 (N1595, N1564, N1419);
and AND2 (N1596, N1594, N998);
xor XOR2 (N1597, N1588, N723);
nor NOR3 (N1598, N1582, N649, N114);
nor NOR2 (N1599, N1596, N1252);
xor XOR2 (N1600, N1577, N1428);
nand NAND3 (N1601, N1583, N625, N108);
and AND3 (N1602, N1593, N950, N1241);
or OR4 (N1603, N1597, N893, N201, N1435);
and AND3 (N1604, N1601, N1549, N1022);
xor XOR2 (N1605, N1572, N356);
nor NOR3 (N1606, N1603, N1213, N1489);
nor NOR4 (N1607, N1604, N454, N1511, N1491);
nand NAND2 (N1608, N1599, N156);
nor NOR3 (N1609, N1600, N453, N516);
and AND4 (N1610, N1609, N1058, N422, N331);
and AND3 (N1611, N1607, N594, N474);
not NOT1 (N1612, N1608);
and AND3 (N1613, N1606, N301, N1588);
xor XOR2 (N1614, N1613, N141);
nor NOR2 (N1615, N1605, N1412);
or OR4 (N1616, N1598, N1325, N51, N220);
xor XOR2 (N1617, N1614, N637);
nor NOR3 (N1618, N1602, N973, N240);
nand NAND3 (N1619, N1610, N1523, N1025);
and AND2 (N1620, N1619, N784);
not NOT1 (N1621, N1611);
xor XOR2 (N1622, N1618, N533);
nor NOR4 (N1623, N1615, N1155, N503, N1130);
xor XOR2 (N1624, N1612, N546);
and AND2 (N1625, N1623, N1074);
nand NAND2 (N1626, N1621, N1101);
buf BUF1 (N1627, N1624);
xor XOR2 (N1628, N1622, N1579);
and AND4 (N1629, N1595, N493, N1306, N1491);
or OR4 (N1630, N1629, N320, N1104, N154);
not NOT1 (N1631, N1587);
xor XOR2 (N1632, N1617, N780);
not NOT1 (N1633, N1632);
or OR2 (N1634, N1625, N547);
not NOT1 (N1635, N1627);
xor XOR2 (N1636, N1591, N978);
nand NAND2 (N1637, N1635, N400);
xor XOR2 (N1638, N1616, N1365);
or OR4 (N1639, N1631, N100, N1381, N1184);
buf BUF1 (N1640, N1633);
and AND2 (N1641, N1637, N1508);
xor XOR2 (N1642, N1628, N685);
or OR3 (N1643, N1620, N254, N1143);
buf BUF1 (N1644, N1641);
not NOT1 (N1645, N1636);
not NOT1 (N1646, N1639);
nor NOR2 (N1647, N1642, N963);
buf BUF1 (N1648, N1638);
xor XOR2 (N1649, N1644, N798);
nand NAND3 (N1650, N1626, N281, N797);
and AND2 (N1651, N1630, N862);
buf BUF1 (N1652, N1634);
or OR3 (N1653, N1650, N633, N638);
not NOT1 (N1654, N1649);
or OR2 (N1655, N1640, N277);
or OR3 (N1656, N1646, N1532, N635);
nor NOR2 (N1657, N1655, N1004);
or OR4 (N1658, N1651, N265, N1534, N736);
and AND2 (N1659, N1643, N928);
nor NOR4 (N1660, N1653, N1036, N66, N401);
xor XOR2 (N1661, N1657, N639);
and AND2 (N1662, N1656, N879);
buf BUF1 (N1663, N1647);
or OR3 (N1664, N1645, N481, N1601);
not NOT1 (N1665, N1654);
and AND3 (N1666, N1665, N303, N1110);
not NOT1 (N1667, N1663);
or OR3 (N1668, N1667, N671, N1227);
xor XOR2 (N1669, N1661, N1388);
nor NOR3 (N1670, N1668, N966, N188);
buf BUF1 (N1671, N1670);
not NOT1 (N1672, N1659);
or OR2 (N1673, N1652, N1662);
nor NOR4 (N1674, N26, N1319, N521, N1444);
nand NAND2 (N1675, N1664, N1140);
xor XOR2 (N1676, N1658, N1319);
and AND4 (N1677, N1660, N1146, N1392, N185);
buf BUF1 (N1678, N1673);
and AND4 (N1679, N1677, N1074, N449, N1470);
buf BUF1 (N1680, N1678);
xor XOR2 (N1681, N1674, N369);
and AND2 (N1682, N1679, N1158);
nand NAND4 (N1683, N1675, N21, N908, N879);
and AND3 (N1684, N1680, N518, N1389);
buf BUF1 (N1685, N1671);
or OR2 (N1686, N1682, N186);
buf BUF1 (N1687, N1676);
buf BUF1 (N1688, N1683);
nand NAND2 (N1689, N1685, N248);
nor NOR2 (N1690, N1669, N1272);
xor XOR2 (N1691, N1690, N1168);
nor NOR2 (N1692, N1684, N644);
not NOT1 (N1693, N1689);
nor NOR3 (N1694, N1692, N792, N1146);
nand NAND4 (N1695, N1694, N1256, N891, N1257);
and AND4 (N1696, N1693, N1084, N57, N1035);
xor XOR2 (N1697, N1695, N41);
nand NAND3 (N1698, N1687, N547, N586);
and AND3 (N1699, N1691, N720, N1595);
xor XOR2 (N1700, N1697, N748);
nand NAND3 (N1701, N1666, N1520, N1504);
xor XOR2 (N1702, N1701, N847);
buf BUF1 (N1703, N1700);
nand NAND3 (N1704, N1672, N1669, N533);
not NOT1 (N1705, N1688);
and AND3 (N1706, N1681, N1117, N781);
or OR3 (N1707, N1698, N881, N807);
nand NAND2 (N1708, N1702, N590);
or OR3 (N1709, N1703, N1541, N1070);
nor NOR3 (N1710, N1686, N1395, N152);
xor XOR2 (N1711, N1708, N751);
xor XOR2 (N1712, N1710, N503);
buf BUF1 (N1713, N1706);
and AND3 (N1714, N1648, N234, N1560);
and AND3 (N1715, N1704, N1705, N1290);
nand NAND2 (N1716, N1166, N1057);
nor NOR4 (N1717, N1699, N277, N71, N1129);
and AND3 (N1718, N1716, N395, N1096);
buf BUF1 (N1719, N1718);
and AND2 (N1720, N1696, N1299);
or OR3 (N1721, N1715, N49, N260);
xor XOR2 (N1722, N1714, N909);
nand NAND4 (N1723, N1717, N94, N718, N1293);
and AND3 (N1724, N1711, N594, N194);
buf BUF1 (N1725, N1721);
buf BUF1 (N1726, N1722);
not NOT1 (N1727, N1719);
xor XOR2 (N1728, N1726, N1584);
not NOT1 (N1729, N1723);
or OR3 (N1730, N1713, N96, N1367);
nand NAND3 (N1731, N1730, N835, N1199);
and AND4 (N1732, N1728, N167, N613, N239);
nor NOR2 (N1733, N1724, N1350);
not NOT1 (N1734, N1720);
nor NOR4 (N1735, N1733, N556, N362, N258);
nor NOR4 (N1736, N1732, N938, N535, N1037);
not NOT1 (N1737, N1735);
nor NOR2 (N1738, N1709, N927);
xor XOR2 (N1739, N1707, N854);
not NOT1 (N1740, N1737);
not NOT1 (N1741, N1729);
not NOT1 (N1742, N1740);
buf BUF1 (N1743, N1741);
xor XOR2 (N1744, N1743, N707);
or OR2 (N1745, N1731, N296);
buf BUF1 (N1746, N1744);
buf BUF1 (N1747, N1725);
not NOT1 (N1748, N1745);
nor NOR3 (N1749, N1748, N880, N1127);
or OR2 (N1750, N1739, N287);
or OR2 (N1751, N1742, N882);
or OR4 (N1752, N1746, N1538, N649, N340);
or OR2 (N1753, N1750, N605);
and AND2 (N1754, N1747, N267);
and AND4 (N1755, N1712, N1355, N1496, N1712);
and AND4 (N1756, N1727, N1224, N1444, N1141);
and AND2 (N1757, N1749, N461);
xor XOR2 (N1758, N1734, N819);
nor NOR3 (N1759, N1757, N309, N248);
nand NAND3 (N1760, N1756, N976, N1682);
nor NOR2 (N1761, N1738, N1053);
nor NOR2 (N1762, N1752, N869);
nand NAND2 (N1763, N1760, N30);
and AND2 (N1764, N1751, N99);
nand NAND4 (N1765, N1761, N1076, N6, N759);
xor XOR2 (N1766, N1759, N135);
xor XOR2 (N1767, N1754, N146);
xor XOR2 (N1768, N1758, N774);
not NOT1 (N1769, N1762);
nor NOR2 (N1770, N1755, N1381);
nand NAND3 (N1771, N1766, N1425, N277);
and AND3 (N1772, N1768, N1610, N1658);
not NOT1 (N1773, N1767);
nand NAND3 (N1774, N1736, N864, N169);
and AND2 (N1775, N1771, N1050);
nor NOR2 (N1776, N1769, N684);
xor XOR2 (N1777, N1764, N730);
or OR2 (N1778, N1777, N1014);
buf BUF1 (N1779, N1772);
and AND2 (N1780, N1753, N1469);
nor NOR3 (N1781, N1778, N1246, N82);
nand NAND4 (N1782, N1780, N292, N1279, N1559);
xor XOR2 (N1783, N1776, N1140);
or OR2 (N1784, N1765, N424);
buf BUF1 (N1785, N1763);
nor NOR2 (N1786, N1784, N633);
nand NAND2 (N1787, N1785, N798);
not NOT1 (N1788, N1783);
nand NAND2 (N1789, N1775, N288);
and AND3 (N1790, N1789, N637, N1221);
buf BUF1 (N1791, N1774);
or OR4 (N1792, N1779, N100, N303, N538);
nor NOR4 (N1793, N1788, N1064, N31, N1116);
not NOT1 (N1794, N1791);
not NOT1 (N1795, N1793);
or OR3 (N1796, N1782, N1729, N1085);
and AND3 (N1797, N1786, N911, N1061);
and AND2 (N1798, N1787, N568);
or OR3 (N1799, N1781, N470, N1519);
buf BUF1 (N1800, N1770);
xor XOR2 (N1801, N1792, N375);
not NOT1 (N1802, N1800);
xor XOR2 (N1803, N1796, N168);
not NOT1 (N1804, N1799);
buf BUF1 (N1805, N1797);
buf BUF1 (N1806, N1801);
xor XOR2 (N1807, N1798, N1164);
nand NAND2 (N1808, N1806, N850);
nor NOR3 (N1809, N1807, N553, N1020);
not NOT1 (N1810, N1790);
nor NOR2 (N1811, N1802, N1197);
or OR4 (N1812, N1773, N1281, N1316, N470);
and AND4 (N1813, N1808, N1267, N439, N64);
nor NOR2 (N1814, N1805, N101);
not NOT1 (N1815, N1814);
buf BUF1 (N1816, N1809);
or OR3 (N1817, N1803, N1771, N416);
or OR3 (N1818, N1811, N595, N1663);
nand NAND4 (N1819, N1815, N1692, N760, N1129);
xor XOR2 (N1820, N1818, N991);
buf BUF1 (N1821, N1819);
buf BUF1 (N1822, N1812);
not NOT1 (N1823, N1813);
not NOT1 (N1824, N1817);
and AND2 (N1825, N1823, N964);
or OR2 (N1826, N1821, N1441);
or OR3 (N1827, N1795, N424, N524);
nor NOR3 (N1828, N1827, N1231, N1416);
nor NOR3 (N1829, N1822, N597, N711);
nor NOR4 (N1830, N1824, N1538, N261, N857);
nand NAND2 (N1831, N1794, N1452);
nor NOR2 (N1832, N1828, N916);
buf BUF1 (N1833, N1829);
nand NAND3 (N1834, N1825, N739, N59);
xor XOR2 (N1835, N1832, N861);
and AND4 (N1836, N1826, N243, N1777, N41);
not NOT1 (N1837, N1820);
xor XOR2 (N1838, N1804, N1233);
buf BUF1 (N1839, N1838);
xor XOR2 (N1840, N1834, N1598);
not NOT1 (N1841, N1835);
xor XOR2 (N1842, N1810, N182);
or OR2 (N1843, N1833, N744);
nor NOR2 (N1844, N1843, N1242);
or OR4 (N1845, N1830, N1135, N1307, N1456);
buf BUF1 (N1846, N1837);
or OR3 (N1847, N1840, N1738, N791);
or OR3 (N1848, N1839, N267, N724);
xor XOR2 (N1849, N1848, N867);
xor XOR2 (N1850, N1836, N1334);
nand NAND3 (N1851, N1831, N470, N1170);
buf BUF1 (N1852, N1847);
nand NAND2 (N1853, N1849, N345);
or OR3 (N1854, N1852, N586, N205);
nand NAND2 (N1855, N1854, N4);
or OR4 (N1856, N1842, N1586, N1820, N985);
and AND4 (N1857, N1845, N566, N1097, N1338);
not NOT1 (N1858, N1816);
not NOT1 (N1859, N1841);
nand NAND4 (N1860, N1859, N1800, N499, N183);
nand NAND3 (N1861, N1858, N554, N781);
nand NAND3 (N1862, N1857, N643, N1472);
xor XOR2 (N1863, N1850, N1504);
xor XOR2 (N1864, N1856, N1008);
or OR3 (N1865, N1853, N664, N769);
nor NOR3 (N1866, N1846, N1155, N1421);
and AND4 (N1867, N1864, N1322, N689, N466);
and AND3 (N1868, N1844, N1505, N507);
nand NAND3 (N1869, N1867, N1706, N523);
xor XOR2 (N1870, N1861, N1018);
and AND3 (N1871, N1860, N368, N241);
buf BUF1 (N1872, N1863);
nor NOR3 (N1873, N1865, N1803, N356);
and AND4 (N1874, N1873, N1696, N619, N181);
and AND2 (N1875, N1868, N1656);
xor XOR2 (N1876, N1862, N1843);
or OR2 (N1877, N1855, N977);
or OR3 (N1878, N1874, N1001, N1448);
or OR2 (N1879, N1872, N831);
nand NAND2 (N1880, N1879, N1517);
or OR4 (N1881, N1875, N1457, N404, N47);
not NOT1 (N1882, N1876);
xor XOR2 (N1883, N1878, N1486);
nand NAND3 (N1884, N1869, N1323, N1259);
nor NOR4 (N1885, N1881, N812, N1349, N397);
xor XOR2 (N1886, N1884, N550);
not NOT1 (N1887, N1871);
nand NAND4 (N1888, N1883, N915, N174, N439);
xor XOR2 (N1889, N1887, N1838);
and AND2 (N1890, N1851, N1653);
or OR2 (N1891, N1880, N1242);
not NOT1 (N1892, N1870);
buf BUF1 (N1893, N1885);
not NOT1 (N1894, N1882);
nand NAND4 (N1895, N1866, N1679, N1051, N1546);
and AND2 (N1896, N1892, N1474);
buf BUF1 (N1897, N1886);
not NOT1 (N1898, N1893);
or OR4 (N1899, N1897, N490, N1266, N1334);
nand NAND4 (N1900, N1877, N396, N1293, N1090);
not NOT1 (N1901, N1895);
xor XOR2 (N1902, N1889, N1774);
xor XOR2 (N1903, N1898, N176);
xor XOR2 (N1904, N1899, N1541);
buf BUF1 (N1905, N1891);
or OR3 (N1906, N1890, N324, N559);
buf BUF1 (N1907, N1902);
and AND3 (N1908, N1901, N1472, N793);
nor NOR2 (N1909, N1905, N409);
or OR2 (N1910, N1907, N1384);
xor XOR2 (N1911, N1908, N1399);
not NOT1 (N1912, N1896);
or OR3 (N1913, N1906, N1607, N39);
and AND3 (N1914, N1911, N100, N1439);
xor XOR2 (N1915, N1904, N1819);
not NOT1 (N1916, N1894);
not NOT1 (N1917, N1915);
xor XOR2 (N1918, N1909, N1808);
or OR4 (N1919, N1910, N924, N752, N857);
nor NOR2 (N1920, N1888, N786);
or OR3 (N1921, N1912, N1174, N996);
nor NOR4 (N1922, N1920, N78, N1049, N1758);
xor XOR2 (N1923, N1919, N1473);
buf BUF1 (N1924, N1913);
nand NAND3 (N1925, N1923, N684, N330);
not NOT1 (N1926, N1924);
not NOT1 (N1927, N1914);
buf BUF1 (N1928, N1918);
buf BUF1 (N1929, N1925);
buf BUF1 (N1930, N1900);
xor XOR2 (N1931, N1903, N1308);
buf BUF1 (N1932, N1916);
and AND2 (N1933, N1929, N889);
nand NAND2 (N1934, N1931, N249);
nor NOR2 (N1935, N1930, N531);
nor NOR3 (N1936, N1921, N1570, N1339);
and AND2 (N1937, N1928, N1240);
nand NAND3 (N1938, N1917, N1898, N290);
or OR3 (N1939, N1937, N408, N959);
and AND4 (N1940, N1939, N1154, N366, N1193);
and AND3 (N1941, N1934, N819, N1462);
and AND3 (N1942, N1938, N339, N1394);
and AND3 (N1943, N1940, N1011, N1888);
not NOT1 (N1944, N1941);
not NOT1 (N1945, N1935);
or OR2 (N1946, N1945, N1524);
xor XOR2 (N1947, N1932, N1392);
xor XOR2 (N1948, N1946, N393);
and AND2 (N1949, N1942, N296);
nor NOR3 (N1950, N1936, N350, N1215);
and AND3 (N1951, N1933, N144, N64);
not NOT1 (N1952, N1944);
not NOT1 (N1953, N1947);
nand NAND4 (N1954, N1952, N720, N1490, N469);
nor NOR2 (N1955, N1949, N1848);
and AND4 (N1956, N1927, N1936, N157, N1723);
nand NAND4 (N1957, N1950, N1247, N661, N47);
nand NAND3 (N1958, N1953, N1882, N63);
or OR3 (N1959, N1956, N1117, N106);
xor XOR2 (N1960, N1926, N7);
buf BUF1 (N1961, N1954);
xor XOR2 (N1962, N1922, N35);
xor XOR2 (N1963, N1943, N482);
and AND2 (N1964, N1961, N675);
nor NOR2 (N1965, N1955, N77);
and AND2 (N1966, N1958, N760);
xor XOR2 (N1967, N1951, N1158);
or OR4 (N1968, N1962, N661, N736, N113);
nor NOR4 (N1969, N1959, N1432, N1777, N31);
buf BUF1 (N1970, N1968);
not NOT1 (N1971, N1967);
nand NAND2 (N1972, N1970, N1153);
xor XOR2 (N1973, N1948, N1690);
and AND4 (N1974, N1969, N1200, N509, N703);
buf BUF1 (N1975, N1972);
or OR2 (N1976, N1963, N1209);
or OR4 (N1977, N1965, N1604, N364, N110);
nor NOR3 (N1978, N1975, N553, N1590);
and AND4 (N1979, N1977, N1224, N1310, N381);
or OR2 (N1980, N1973, N31);
and AND2 (N1981, N1957, N1514);
and AND4 (N1982, N1979, N1783, N753, N505);
and AND3 (N1983, N1982, N899, N259);
nor NOR3 (N1984, N1983, N351, N1785);
nor NOR2 (N1985, N1978, N684);
nor NOR3 (N1986, N1984, N1213, N1623);
buf BUF1 (N1987, N1960);
and AND2 (N1988, N1980, N1561);
and AND2 (N1989, N1966, N1519);
buf BUF1 (N1990, N1986);
buf BUF1 (N1991, N1974);
nand NAND3 (N1992, N1985, N1930, N755);
nor NOR4 (N1993, N1987, N985, N1085, N1341);
or OR4 (N1994, N1971, N1282, N1660, N494);
not NOT1 (N1995, N1994);
nand NAND3 (N1996, N1991, N374, N570);
xor XOR2 (N1997, N1995, N1304);
or OR2 (N1998, N1993, N830);
buf BUF1 (N1999, N1976);
or OR3 (N2000, N1999, N1349, N1294);
and AND2 (N2001, N1992, N1189);
or OR3 (N2002, N1981, N1079, N1264);
xor XOR2 (N2003, N1996, N393);
xor XOR2 (N2004, N2001, N1244);
or OR3 (N2005, N1990, N1706, N1876);
xor XOR2 (N2006, N1997, N1242);
or OR3 (N2007, N2000, N1575, N1623);
nor NOR2 (N2008, N1998, N1130);
or OR2 (N2009, N1964, N943);
nor NOR4 (N2010, N2004, N688, N1566, N300);
nor NOR3 (N2011, N2010, N767, N437);
nand NAND3 (N2012, N1989, N256, N408);
buf BUF1 (N2013, N2008);
nor NOR3 (N2014, N2013, N1350, N1440);
nor NOR4 (N2015, N2014, N1635, N967, N1422);
nor NOR3 (N2016, N2003, N1716, N615);
and AND3 (N2017, N2012, N142, N1324);
buf BUF1 (N2018, N2017);
or OR3 (N2019, N2011, N157, N1409);
xor XOR2 (N2020, N2015, N205);
not NOT1 (N2021, N2020);
nor NOR3 (N2022, N2016, N714, N1011);
nand NAND3 (N2023, N2005, N1449, N334);
and AND4 (N2024, N2002, N1010, N787, N712);
buf BUF1 (N2025, N2018);
not NOT1 (N2026, N2009);
and AND2 (N2027, N2021, N1808);
nor NOR2 (N2028, N2006, N1434);
not NOT1 (N2029, N2026);
not NOT1 (N2030, N1988);
xor XOR2 (N2031, N2019, N1096);
nor NOR2 (N2032, N2030, N1792);
not NOT1 (N2033, N2031);
buf BUF1 (N2034, N2032);
or OR2 (N2035, N2028, N247);
buf BUF1 (N2036, N2007);
nand NAND3 (N2037, N2036, N813, N1687);
not NOT1 (N2038, N2029);
buf BUF1 (N2039, N2025);
xor XOR2 (N2040, N2039, N250);
buf BUF1 (N2041, N2034);
xor XOR2 (N2042, N2022, N1268);
or OR2 (N2043, N2038, N240);
nor NOR2 (N2044, N2027, N519);
not NOT1 (N2045, N2035);
nand NAND2 (N2046, N2045, N981);
or OR2 (N2047, N2044, N151);
and AND3 (N2048, N2037, N419, N1870);
buf BUF1 (N2049, N2043);
buf BUF1 (N2050, N2023);
nand NAND4 (N2051, N2049, N1495, N1508, N1879);
and AND3 (N2052, N2047, N445, N117);
not NOT1 (N2053, N2046);
and AND3 (N2054, N2051, N187, N193);
xor XOR2 (N2055, N2040, N837);
nand NAND3 (N2056, N2048, N393, N796);
nor NOR3 (N2057, N2054, N2037, N896);
and AND2 (N2058, N2050, N1184);
and AND4 (N2059, N2058, N1227, N1236, N1751);
and AND3 (N2060, N2052, N316, N1003);
and AND4 (N2061, N2059, N68, N2020, N1382);
or OR4 (N2062, N2056, N1782, N20, N1322);
xor XOR2 (N2063, N2041, N100);
or OR3 (N2064, N2053, N1952, N1420);
nand NAND3 (N2065, N2033, N449, N880);
buf BUF1 (N2066, N2057);
buf BUF1 (N2067, N2062);
or OR4 (N2068, N2024, N1747, N484, N125);
xor XOR2 (N2069, N2055, N3);
not NOT1 (N2070, N2060);
or OR2 (N2071, N2067, N586);
and AND4 (N2072, N2065, N1716, N1381, N1555);
xor XOR2 (N2073, N2064, N1337);
and AND3 (N2074, N2070, N1697, N1071);
or OR2 (N2075, N2073, N1331);
and AND4 (N2076, N2071, N1244, N527, N1788);
nor NOR2 (N2077, N2075, N1572);
nor NOR3 (N2078, N2066, N52, N1502);
buf BUF1 (N2079, N2069);
xor XOR2 (N2080, N2068, N616);
not NOT1 (N2081, N2061);
nand NAND3 (N2082, N2078, N1548, N426);
xor XOR2 (N2083, N2063, N1190);
and AND2 (N2084, N2080, N606);
xor XOR2 (N2085, N2084, N217);
not NOT1 (N2086, N2079);
not NOT1 (N2087, N2072);
and AND3 (N2088, N2082, N1889, N1873);
or OR3 (N2089, N2087, N407, N1817);
nor NOR3 (N2090, N2081, N1451, N1226);
and AND2 (N2091, N2090, N1219);
not NOT1 (N2092, N2091);
or OR4 (N2093, N2076, N1430, N1232, N523);
nor NOR3 (N2094, N2074, N146, N1056);
xor XOR2 (N2095, N2088, N25);
nand NAND2 (N2096, N2042, N1321);
xor XOR2 (N2097, N2092, N764);
and AND4 (N2098, N2094, N1929, N1435, N1786);
nand NAND4 (N2099, N2077, N903, N2047, N1139);
nor NOR4 (N2100, N2089, N428, N1395, N599);
nor NOR4 (N2101, N2086, N1946, N1538, N673);
buf BUF1 (N2102, N2097);
not NOT1 (N2103, N2102);
buf BUF1 (N2104, N2083);
nand NAND3 (N2105, N2096, N1741, N1639);
not NOT1 (N2106, N2095);
buf BUF1 (N2107, N2085);
buf BUF1 (N2108, N2103);
not NOT1 (N2109, N2101);
nand NAND2 (N2110, N2107, N928);
xor XOR2 (N2111, N2093, N1969);
or OR3 (N2112, N2104, N670, N2014);
xor XOR2 (N2113, N2111, N462);
and AND4 (N2114, N2108, N633, N1542, N570);
or OR2 (N2115, N2113, N1310);
buf BUF1 (N2116, N2114);
and AND2 (N2117, N2115, N1503);
xor XOR2 (N2118, N2106, N1547);
xor XOR2 (N2119, N2099, N399);
not NOT1 (N2120, N2098);
and AND2 (N2121, N2105, N300);
or OR4 (N2122, N2100, N1582, N92, N1552);
xor XOR2 (N2123, N2119, N1510);
buf BUF1 (N2124, N2109);
nand NAND3 (N2125, N2112, N509, N1465);
buf BUF1 (N2126, N2121);
buf BUF1 (N2127, N2126);
or OR4 (N2128, N2116, N1933, N1713, N832);
or OR3 (N2129, N2128, N118, N1097);
or OR3 (N2130, N2123, N1244, N2050);
nor NOR4 (N2131, N2110, N1730, N926, N1302);
buf BUF1 (N2132, N2130);
or OR3 (N2133, N2120, N1558, N1397);
not NOT1 (N2134, N2133);
or OR2 (N2135, N2124, N1961);
and AND4 (N2136, N2135, N72, N1211, N495);
not NOT1 (N2137, N2127);
or OR4 (N2138, N2131, N1067, N2086, N384);
nand NAND3 (N2139, N2136, N686, N1441);
nand NAND2 (N2140, N2132, N1683);
not NOT1 (N2141, N2139);
xor XOR2 (N2142, N2141, N51);
or OR3 (N2143, N2140, N2058, N1338);
xor XOR2 (N2144, N2117, N217);
xor XOR2 (N2145, N2138, N2049);
and AND2 (N2146, N2144, N1356);
buf BUF1 (N2147, N2134);
buf BUF1 (N2148, N2122);
not NOT1 (N2149, N2147);
not NOT1 (N2150, N2146);
or OR2 (N2151, N2125, N152);
and AND3 (N2152, N2143, N845, N835);
nor NOR2 (N2153, N2149, N1277);
not NOT1 (N2154, N2137);
nand NAND4 (N2155, N2154, N436, N1391, N219);
or OR3 (N2156, N2118, N996, N987);
or OR4 (N2157, N2152, N169, N483, N553);
or OR4 (N2158, N2148, N1502, N630, N121);
xor XOR2 (N2159, N2150, N79);
not NOT1 (N2160, N2129);
and AND2 (N2161, N2145, N1743);
nor NOR4 (N2162, N2161, N1357, N266, N641);
not NOT1 (N2163, N2155);
not NOT1 (N2164, N2158);
xor XOR2 (N2165, N2163, N995);
nor NOR4 (N2166, N2164, N967, N874, N1477);
nand NAND4 (N2167, N2159, N45, N792, N749);
buf BUF1 (N2168, N2165);
or OR3 (N2169, N2160, N1618, N1858);
buf BUF1 (N2170, N2142);
nor NOR3 (N2171, N2153, N627, N387);
or OR2 (N2172, N2169, N125);
buf BUF1 (N2173, N2151);
and AND2 (N2174, N2157, N154);
not NOT1 (N2175, N2162);
not NOT1 (N2176, N2172);
not NOT1 (N2177, N2171);
xor XOR2 (N2178, N2175, N1046);
or OR4 (N2179, N2168, N39, N1891, N1552);
nand NAND3 (N2180, N2167, N578, N2033);
nor NOR2 (N2181, N2173, N195);
xor XOR2 (N2182, N2178, N857);
xor XOR2 (N2183, N2179, N1252);
buf BUF1 (N2184, N2177);
buf BUF1 (N2185, N2184);
or OR3 (N2186, N2181, N2146, N1587);
buf BUF1 (N2187, N2166);
nor NOR3 (N2188, N2174, N1722, N263);
nand NAND4 (N2189, N2182, N1726, N1230, N933);
and AND3 (N2190, N2156, N101, N1227);
nand NAND4 (N2191, N2185, N1318, N1622, N677);
nand NAND2 (N2192, N2170, N969);
nand NAND4 (N2193, N2188, N407, N605, N642);
and AND4 (N2194, N2180, N488, N2050, N2101);
xor XOR2 (N2195, N2193, N1091);
and AND4 (N2196, N2186, N1484, N2052, N1702);
buf BUF1 (N2197, N2183);
buf BUF1 (N2198, N2197);
xor XOR2 (N2199, N2198, N1515);
not NOT1 (N2200, N2187);
nor NOR4 (N2201, N2195, N2165, N809, N2036);
nand NAND4 (N2202, N2200, N900, N1112, N1515);
xor XOR2 (N2203, N2190, N1036);
xor XOR2 (N2204, N2176, N1279);
buf BUF1 (N2205, N2196);
not NOT1 (N2206, N2204);
and AND3 (N2207, N2203, N515, N1162);
and AND2 (N2208, N2202, N1383);
xor XOR2 (N2209, N2189, N2171);
xor XOR2 (N2210, N2206, N603);
xor XOR2 (N2211, N2210, N55);
nand NAND2 (N2212, N2208, N1799);
xor XOR2 (N2213, N2199, N1588);
not NOT1 (N2214, N2212);
and AND4 (N2215, N2214, N778, N869, N578);
xor XOR2 (N2216, N2215, N890);
buf BUF1 (N2217, N2192);
nand NAND3 (N2218, N2201, N1086, N695);
nor NOR4 (N2219, N2211, N1229, N94, N331);
nor NOR2 (N2220, N2207, N1261);
not NOT1 (N2221, N2216);
nor NOR2 (N2222, N2219, N1208);
nor NOR4 (N2223, N2194, N2089, N2168, N22);
or OR3 (N2224, N2191, N452, N2055);
or OR4 (N2225, N2220, N1100, N613, N1556);
xor XOR2 (N2226, N2221, N1204);
nor NOR2 (N2227, N2205, N1463);
not NOT1 (N2228, N2218);
nand NAND3 (N2229, N2226, N27, N1264);
not NOT1 (N2230, N2227);
or OR3 (N2231, N2217, N1242, N2012);
or OR3 (N2232, N2231, N562, N1676);
nor NOR4 (N2233, N2225, N1227, N904, N1295);
not NOT1 (N2234, N2233);
xor XOR2 (N2235, N2228, N2033);
nor NOR2 (N2236, N2230, N638);
buf BUF1 (N2237, N2235);
buf BUF1 (N2238, N2209);
and AND4 (N2239, N2213, N155, N1177, N1994);
buf BUF1 (N2240, N2236);
buf BUF1 (N2241, N2224);
not NOT1 (N2242, N2223);
not NOT1 (N2243, N2222);
xor XOR2 (N2244, N2229, N1341);
and AND3 (N2245, N2232, N75, N1873);
and AND2 (N2246, N2240, N1969);
xor XOR2 (N2247, N2245, N1581);
or OR4 (N2248, N2244, N1655, N672, N2154);
or OR3 (N2249, N2239, N698, N355);
buf BUF1 (N2250, N2234);
not NOT1 (N2251, N2242);
and AND3 (N2252, N2248, N661, N647);
nor NOR3 (N2253, N2249, N2034, N654);
nand NAND3 (N2254, N2247, N800, N396);
or OR2 (N2255, N2250, N1087);
buf BUF1 (N2256, N2237);
not NOT1 (N2257, N2256);
and AND4 (N2258, N2246, N1583, N1779, N2248);
nand NAND3 (N2259, N2241, N1664, N902);
nand NAND2 (N2260, N2253, N1902);
nor NOR4 (N2261, N2243, N317, N736, N416);
and AND4 (N2262, N2259, N1979, N363, N358);
xor XOR2 (N2263, N2255, N1717);
xor XOR2 (N2264, N2257, N935);
not NOT1 (N2265, N2260);
nor NOR4 (N2266, N2264, N6, N1049, N542);
and AND3 (N2267, N2262, N1434, N2145);
or OR2 (N2268, N2238, N2190);
and AND2 (N2269, N2267, N1649);
or OR3 (N2270, N2261, N1097, N1937);
and AND4 (N2271, N2268, N1338, N318, N1810);
and AND4 (N2272, N2265, N267, N784, N2048);
xor XOR2 (N2273, N2254, N1896);
not NOT1 (N2274, N2252);
xor XOR2 (N2275, N2251, N631);
and AND4 (N2276, N2269, N516, N1528, N2);
buf BUF1 (N2277, N2270);
nor NOR4 (N2278, N2274, N802, N136, N1204);
or OR4 (N2279, N2271, N1259, N2123, N1914);
or OR2 (N2280, N2272, N997);
xor XOR2 (N2281, N2263, N1985);
and AND4 (N2282, N2266, N2258, N249, N2009);
nor NOR4 (N2283, N253, N918, N538, N89);
not NOT1 (N2284, N2282);
and AND4 (N2285, N2281, N1051, N522, N182);
xor XOR2 (N2286, N2273, N643);
not NOT1 (N2287, N2275);
nor NOR2 (N2288, N2278, N1258);
nor NOR3 (N2289, N2279, N1019, N682);
buf BUF1 (N2290, N2286);
and AND4 (N2291, N2285, N212, N1588, N695);
nor NOR3 (N2292, N2288, N2096, N1710);
buf BUF1 (N2293, N2280);
and AND4 (N2294, N2289, N1856, N2042, N469);
xor XOR2 (N2295, N2290, N115);
or OR3 (N2296, N2276, N2240, N2039);
and AND2 (N2297, N2294, N1277);
xor XOR2 (N2298, N2287, N824);
or OR3 (N2299, N2297, N1305, N1973);
or OR2 (N2300, N2291, N277);
nand NAND2 (N2301, N2300, N1533);
buf BUF1 (N2302, N2295);
or OR3 (N2303, N2298, N2042, N2264);
nand NAND3 (N2304, N2303, N813, N1577);
nor NOR4 (N2305, N2302, N2004, N1037, N1412);
nor NOR3 (N2306, N2299, N1382, N1773);
xor XOR2 (N2307, N2293, N178);
or OR2 (N2308, N2305, N1388);
nand NAND2 (N2309, N2304, N428);
or OR3 (N2310, N2284, N2247, N856);
not NOT1 (N2311, N2296);
xor XOR2 (N2312, N2292, N2203);
buf BUF1 (N2313, N2309);
buf BUF1 (N2314, N2307);
buf BUF1 (N2315, N2277);
nor NOR2 (N2316, N2301, N2273);
or OR3 (N2317, N2311, N2140, N1330);
not NOT1 (N2318, N2312);
buf BUF1 (N2319, N2317);
nand NAND4 (N2320, N2319, N2140, N912, N1708);
buf BUF1 (N2321, N2316);
or OR4 (N2322, N2283, N432, N2197, N2122);
nand NAND3 (N2323, N2320, N1469, N627);
and AND3 (N2324, N2313, N1758, N395);
not NOT1 (N2325, N2310);
or OR3 (N2326, N2318, N37, N1476);
not NOT1 (N2327, N2315);
not NOT1 (N2328, N2314);
not NOT1 (N2329, N2308);
buf BUF1 (N2330, N2321);
or OR2 (N2331, N2323, N2159);
xor XOR2 (N2332, N2327, N2035);
buf BUF1 (N2333, N2306);
xor XOR2 (N2334, N2328, N1719);
buf BUF1 (N2335, N2329);
xor XOR2 (N2336, N2325, N1267);
nor NOR3 (N2337, N2334, N1899, N1098);
nor NOR4 (N2338, N2335, N973, N1512, N2292);
and AND2 (N2339, N2326, N175);
buf BUF1 (N2340, N2324);
or OR3 (N2341, N2339, N2320, N992);
nand NAND3 (N2342, N2337, N1388, N1238);
nand NAND4 (N2343, N2336, N1909, N696, N640);
xor XOR2 (N2344, N2332, N1715);
xor XOR2 (N2345, N2331, N1478);
or OR4 (N2346, N2341, N67, N1099, N612);
nor NOR2 (N2347, N2340, N281);
nor NOR3 (N2348, N2338, N1206, N889);
xor XOR2 (N2349, N2330, N445);
not NOT1 (N2350, N2345);
nand NAND3 (N2351, N2344, N684, N1443);
nor NOR3 (N2352, N2351, N891, N930);
or OR2 (N2353, N2333, N1341);
nand NAND2 (N2354, N2353, N2136);
nand NAND3 (N2355, N2322, N570, N683);
and AND3 (N2356, N2346, N1309, N413);
buf BUF1 (N2357, N2343);
nor NOR4 (N2358, N2356, N1669, N2316, N543);
or OR2 (N2359, N2347, N1908);
nor NOR4 (N2360, N2349, N1909, N1754, N605);
and AND2 (N2361, N2355, N134);
buf BUF1 (N2362, N2357);
nor NOR2 (N2363, N2350, N748);
not NOT1 (N2364, N2363);
and AND4 (N2365, N2361, N1092, N1001, N1603);
and AND4 (N2366, N2358, N1859, N291, N1722);
xor XOR2 (N2367, N2362, N462);
xor XOR2 (N2368, N2365, N1578);
and AND4 (N2369, N2366, N1738, N2102, N796);
and AND4 (N2370, N2368, N1992, N302, N1188);
buf BUF1 (N2371, N2367);
not NOT1 (N2372, N2370);
nand NAND3 (N2373, N2359, N505, N86);
nand NAND4 (N2374, N2364, N1461, N1155, N1296);
buf BUF1 (N2375, N2342);
nand NAND4 (N2376, N2374, N1448, N484, N988);
nand NAND4 (N2377, N2376, N1556, N2342, N2118);
buf BUF1 (N2378, N2369);
and AND2 (N2379, N2360, N436);
not NOT1 (N2380, N2377);
buf BUF1 (N2381, N2372);
xor XOR2 (N2382, N2379, N997);
xor XOR2 (N2383, N2380, N1300);
nand NAND2 (N2384, N2354, N1883);
xor XOR2 (N2385, N2383, N1143);
nor NOR2 (N2386, N2373, N1522);
not NOT1 (N2387, N2381);
or OR4 (N2388, N2371, N1713, N2127, N1784);
nand NAND2 (N2389, N2378, N1472);
or OR4 (N2390, N2389, N1495, N1123, N164);
and AND3 (N2391, N2387, N1666, N1689);
not NOT1 (N2392, N2390);
nand NAND3 (N2393, N2348, N1426, N1476);
or OR3 (N2394, N2391, N1170, N982);
xor XOR2 (N2395, N2382, N958);
not NOT1 (N2396, N2384);
nor NOR3 (N2397, N2386, N1633, N1363);
or OR2 (N2398, N2395, N1363);
nand NAND4 (N2399, N2394, N1562, N2339, N606);
nand NAND2 (N2400, N2392, N562);
xor XOR2 (N2401, N2388, N522);
buf BUF1 (N2402, N2400);
or OR3 (N2403, N2393, N688, N334);
and AND4 (N2404, N2375, N83, N97, N1928);
or OR2 (N2405, N2399, N1717);
nor NOR4 (N2406, N2397, N1763, N995, N783);
buf BUF1 (N2407, N2401);
and AND2 (N2408, N2404, N1466);
and AND4 (N2409, N2407, N1190, N363, N1092);
nor NOR4 (N2410, N2352, N1561, N2398, N1742);
buf BUF1 (N2411, N1922);
nor NOR4 (N2412, N2385, N43, N862, N672);
not NOT1 (N2413, N2409);
nor NOR2 (N2414, N2406, N2226);
not NOT1 (N2415, N2412);
xor XOR2 (N2416, N2405, N1042);
nor NOR2 (N2417, N2396, N679);
nor NOR2 (N2418, N2416, N868);
or OR2 (N2419, N2411, N402);
xor XOR2 (N2420, N2408, N305);
not NOT1 (N2421, N2419);
xor XOR2 (N2422, N2402, N1116);
or OR3 (N2423, N2403, N275, N917);
nand NAND3 (N2424, N2415, N951, N929);
xor XOR2 (N2425, N2418, N1896);
nand NAND4 (N2426, N2414, N1143, N1222, N1549);
nor NOR4 (N2427, N2420, N464, N1011, N556);
nand NAND4 (N2428, N2410, N1271, N403, N1818);
buf BUF1 (N2429, N2417);
and AND4 (N2430, N2424, N930, N2407, N311);
nor NOR3 (N2431, N2427, N2092, N435);
nand NAND3 (N2432, N2429, N2224, N146);
and AND2 (N2433, N2425, N1153);
buf BUF1 (N2434, N2423);
buf BUF1 (N2435, N2434);
or OR3 (N2436, N2430, N171, N1268);
nor NOR3 (N2437, N2422, N2275, N2046);
not NOT1 (N2438, N2433);
nand NAND3 (N2439, N2426, N609, N1340);
not NOT1 (N2440, N2432);
and AND2 (N2441, N2431, N799);
nor NOR2 (N2442, N2413, N639);
nor NOR4 (N2443, N2436, N69, N462, N1618);
or OR2 (N2444, N2438, N1787);
not NOT1 (N2445, N2444);
nor NOR2 (N2446, N2441, N1325);
or OR4 (N2447, N2437, N509, N367, N242);
nand NAND3 (N2448, N2428, N2014, N989);
not NOT1 (N2449, N2443);
nor NOR2 (N2450, N2449, N2384);
not NOT1 (N2451, N2450);
not NOT1 (N2452, N2440);
or OR3 (N2453, N2439, N1300, N1007);
or OR4 (N2454, N2421, N2186, N2313, N250);
xor XOR2 (N2455, N2453, N564);
not NOT1 (N2456, N2448);
or OR4 (N2457, N2456, N2088, N1099, N557);
buf BUF1 (N2458, N2446);
not NOT1 (N2459, N2454);
and AND4 (N2460, N2435, N1624, N2417, N351);
xor XOR2 (N2461, N2459, N1295);
or OR2 (N2462, N2458, N776);
nor NOR2 (N2463, N2452, N932);
or OR2 (N2464, N2457, N1753);
nand NAND3 (N2465, N2451, N45, N1926);
nor NOR2 (N2466, N2461, N1269);
xor XOR2 (N2467, N2465, N165);
nand NAND3 (N2468, N2455, N1099, N865);
nor NOR3 (N2469, N2466, N1969, N1943);
and AND3 (N2470, N2445, N779, N1214);
and AND4 (N2471, N2467, N1154, N1707, N2289);
buf BUF1 (N2472, N2470);
nor NOR3 (N2473, N2462, N359, N263);
xor XOR2 (N2474, N2463, N1063);
nor NOR3 (N2475, N2474, N1539, N709);
not NOT1 (N2476, N2471);
not NOT1 (N2477, N2442);
nand NAND4 (N2478, N2460, N1304, N66, N1403);
or OR4 (N2479, N2475, N115, N1543, N1896);
nor NOR3 (N2480, N2476, N298, N430);
nor NOR2 (N2481, N2468, N2353);
xor XOR2 (N2482, N2481, N1356);
nand NAND2 (N2483, N2472, N2096);
nor NOR3 (N2484, N2482, N224, N882);
xor XOR2 (N2485, N2484, N1146);
nor NOR4 (N2486, N2485, N1346, N1709, N852);
buf BUF1 (N2487, N2477);
not NOT1 (N2488, N2480);
and AND4 (N2489, N2488, N93, N2301, N2342);
buf BUF1 (N2490, N2487);
or OR3 (N2491, N2489, N1492, N1113);
or OR2 (N2492, N2491, N1588);
xor XOR2 (N2493, N2483, N2387);
and AND2 (N2494, N2469, N1710);
nand NAND4 (N2495, N2490, N1870, N896, N2421);
and AND3 (N2496, N2493, N317, N1404);
not NOT1 (N2497, N2492);
and AND3 (N2498, N2478, N326, N1929);
not NOT1 (N2499, N2473);
not NOT1 (N2500, N2494);
nand NAND3 (N2501, N2479, N656, N999);
or OR3 (N2502, N2495, N1214, N1471);
nand NAND4 (N2503, N2464, N832, N2239, N2113);
not NOT1 (N2504, N2447);
nor NOR4 (N2505, N2496, N1016, N414, N1787);
buf BUF1 (N2506, N2505);
nand NAND2 (N2507, N2499, N71);
or OR3 (N2508, N2501, N1115, N867);
or OR3 (N2509, N2502, N729, N2103);
buf BUF1 (N2510, N2503);
and AND2 (N2511, N2510, N1418);
buf BUF1 (N2512, N2509);
not NOT1 (N2513, N2511);
and AND3 (N2514, N2486, N1180, N2363);
nor NOR4 (N2515, N2512, N2028, N1132, N1816);
or OR2 (N2516, N2508, N1380);
and AND3 (N2517, N2515, N2048, N2400);
nand NAND4 (N2518, N2517, N1901, N837, N800);
buf BUF1 (N2519, N2506);
or OR2 (N2520, N2498, N1085);
nand NAND3 (N2521, N2513, N2470, N2045);
nor NOR4 (N2522, N2519, N1764, N1154, N730);
not NOT1 (N2523, N2514);
nand NAND4 (N2524, N2522, N388, N230, N73);
and AND2 (N2525, N2518, N1593);
or OR4 (N2526, N2524, N706, N655, N2171);
not NOT1 (N2527, N2520);
nor NOR4 (N2528, N2526, N2396, N1553, N275);
xor XOR2 (N2529, N2528, N762);
not NOT1 (N2530, N2497);
nor NOR3 (N2531, N2516, N472, N2151);
buf BUF1 (N2532, N2529);
nand NAND2 (N2533, N2532, N344);
not NOT1 (N2534, N2531);
not NOT1 (N2535, N2527);
or OR4 (N2536, N2535, N2358, N727, N2052);
nor NOR3 (N2537, N2523, N1984, N1582);
nand NAND3 (N2538, N2537, N683, N195);
nand NAND4 (N2539, N2507, N1151, N24, N972);
nand NAND3 (N2540, N2530, N335, N34);
nand NAND3 (N2541, N2500, N480, N1273);
nor NOR4 (N2542, N2533, N379, N1883, N123);
nor NOR2 (N2543, N2525, N402);
nand NAND4 (N2544, N2536, N1149, N755, N2305);
not NOT1 (N2545, N2540);
nor NOR3 (N2546, N2539, N680, N2252);
nor NOR2 (N2547, N2538, N1505);
buf BUF1 (N2548, N2547);
nor NOR3 (N2549, N2541, N2157, N312);
buf BUF1 (N2550, N2521);
buf BUF1 (N2551, N2550);
nand NAND4 (N2552, N2551, N596, N1872, N2170);
xor XOR2 (N2553, N2546, N1136);
xor XOR2 (N2554, N2553, N675);
xor XOR2 (N2555, N2554, N1927);
not NOT1 (N2556, N2549);
buf BUF1 (N2557, N2534);
or OR2 (N2558, N2544, N1711);
and AND2 (N2559, N2545, N136);
or OR3 (N2560, N2558, N540, N1334);
not NOT1 (N2561, N2552);
and AND3 (N2562, N2556, N1732, N1790);
xor XOR2 (N2563, N2559, N949);
or OR2 (N2564, N2560, N1159);
or OR2 (N2565, N2504, N548);
or OR4 (N2566, N2564, N246, N1121, N1297);
nand NAND4 (N2567, N2562, N997, N606, N1029);
nand NAND3 (N2568, N2565, N1530, N680);
or OR2 (N2569, N2561, N1708);
buf BUF1 (N2570, N2555);
and AND2 (N2571, N2563, N2091);
buf BUF1 (N2572, N2567);
nand NAND3 (N2573, N2571, N734, N1043);
nand NAND4 (N2574, N2557, N648, N56, N1298);
nand NAND2 (N2575, N2568, N1077);
and AND4 (N2576, N2542, N747, N2542, N1574);
not NOT1 (N2577, N2570);
or OR2 (N2578, N2543, N1900);
nor NOR4 (N2579, N2575, N84, N128, N1552);
nor NOR2 (N2580, N2573, N1211);
xor XOR2 (N2581, N2579, N469);
xor XOR2 (N2582, N2580, N1347);
or OR4 (N2583, N2578, N1517, N1985, N1989);
buf BUF1 (N2584, N2569);
or OR3 (N2585, N2566, N484, N630);
xor XOR2 (N2586, N2585, N1354);
nand NAND3 (N2587, N2584, N1576, N2517);
nand NAND2 (N2588, N2572, N1609);
and AND2 (N2589, N2577, N1357);
not NOT1 (N2590, N2589);
not NOT1 (N2591, N2583);
xor XOR2 (N2592, N2548, N268);
nor NOR3 (N2593, N2582, N1909, N972);
not NOT1 (N2594, N2591);
or OR3 (N2595, N2590, N2040, N377);
nand NAND3 (N2596, N2588, N2459, N1288);
not NOT1 (N2597, N2594);
xor XOR2 (N2598, N2587, N187);
or OR2 (N2599, N2581, N2225);
and AND3 (N2600, N2586, N795, N2597);
nor NOR3 (N2601, N355, N1487, N77);
not NOT1 (N2602, N2599);
buf BUF1 (N2603, N2576);
or OR2 (N2604, N2595, N2006);
xor XOR2 (N2605, N2598, N1366);
buf BUF1 (N2606, N2603);
xor XOR2 (N2607, N2574, N497);
or OR4 (N2608, N2596, N1876, N1339, N871);
nand NAND2 (N2609, N2593, N492);
or OR4 (N2610, N2606, N1199, N88, N1830);
and AND2 (N2611, N2604, N814);
xor XOR2 (N2612, N2610, N2283);
or OR3 (N2613, N2605, N1668, N1706);
and AND2 (N2614, N2612, N1143);
or OR3 (N2615, N2600, N1878, N1127);
nor NOR4 (N2616, N2607, N1981, N1251, N1951);
not NOT1 (N2617, N2602);
or OR3 (N2618, N2614, N593, N142);
or OR2 (N2619, N2592, N1390);
not NOT1 (N2620, N2618);
not NOT1 (N2621, N2601);
buf BUF1 (N2622, N2611);
nor NOR3 (N2623, N2609, N1720, N719);
nor NOR4 (N2624, N2622, N2327, N2234, N253);
xor XOR2 (N2625, N2608, N1710);
and AND4 (N2626, N2625, N1702, N241, N1019);
not NOT1 (N2627, N2619);
not NOT1 (N2628, N2620);
not NOT1 (N2629, N2617);
nor NOR4 (N2630, N2615, N1984, N1399, N337);
buf BUF1 (N2631, N2627);
nand NAND2 (N2632, N2629, N446);
nand NAND2 (N2633, N2632, N877);
xor XOR2 (N2634, N2616, N2483);
xor XOR2 (N2635, N2624, N2057);
nand NAND3 (N2636, N2623, N360, N1569);
or OR2 (N2637, N2626, N510);
or OR2 (N2638, N2634, N2061);
nor NOR2 (N2639, N2636, N1131);
nor NOR4 (N2640, N2639, N2143, N2005, N48);
and AND3 (N2641, N2631, N466, N1518);
buf BUF1 (N2642, N2635);
or OR2 (N2643, N2640, N199);
xor XOR2 (N2644, N2638, N1738);
buf BUF1 (N2645, N2637);
and AND3 (N2646, N2642, N1867, N52);
nor NOR3 (N2647, N2613, N1875, N1679);
and AND3 (N2648, N2630, N1224, N1741);
buf BUF1 (N2649, N2643);
buf BUF1 (N2650, N2646);
or OR2 (N2651, N2644, N2189);
and AND3 (N2652, N2633, N1168, N1426);
not NOT1 (N2653, N2641);
buf BUF1 (N2654, N2645);
nor NOR4 (N2655, N2647, N343, N2235, N964);
nand NAND2 (N2656, N2628, N966);
and AND4 (N2657, N2649, N963, N1061, N1204);
or OR4 (N2658, N2651, N2158, N243, N532);
buf BUF1 (N2659, N2657);
and AND4 (N2660, N2658, N697, N2202, N540);
not NOT1 (N2661, N2650);
buf BUF1 (N2662, N2621);
xor XOR2 (N2663, N2653, N1387);
xor XOR2 (N2664, N2660, N690);
nor NOR2 (N2665, N2661, N1963);
xor XOR2 (N2666, N2656, N1538);
xor XOR2 (N2667, N2648, N859);
and AND3 (N2668, N2665, N421, N1014);
or OR2 (N2669, N2654, N1680);
nand NAND4 (N2670, N2659, N2226, N378, N1838);
not NOT1 (N2671, N2664);
xor XOR2 (N2672, N2666, N32);
or OR3 (N2673, N2662, N1368, N1019);
and AND4 (N2674, N2652, N2135, N1512, N2307);
not NOT1 (N2675, N2655);
not NOT1 (N2676, N2669);
and AND3 (N2677, N2670, N1409, N2527);
nand NAND3 (N2678, N2675, N516, N546);
or OR4 (N2679, N2663, N1588, N823, N730);
buf BUF1 (N2680, N2671);
nand NAND4 (N2681, N2677, N2418, N1450, N2183);
not NOT1 (N2682, N2672);
not NOT1 (N2683, N2680);
not NOT1 (N2684, N2667);
and AND3 (N2685, N2683, N948, N870);
nand NAND3 (N2686, N2685, N2391, N1557);
or OR2 (N2687, N2676, N139);
not NOT1 (N2688, N2668);
xor XOR2 (N2689, N2674, N83);
or OR3 (N2690, N2682, N2022, N334);
and AND2 (N2691, N2688, N38);
nand NAND4 (N2692, N2687, N1912, N2231, N1805);
not NOT1 (N2693, N2692);
and AND3 (N2694, N2689, N369, N2428);
nor NOR3 (N2695, N2679, N999, N31);
nand NAND2 (N2696, N2690, N1309);
and AND2 (N2697, N2681, N1569);
nor NOR2 (N2698, N2691, N2575);
nor NOR3 (N2699, N2695, N374, N1272);
nand NAND2 (N2700, N2686, N1296);
and AND2 (N2701, N2697, N1713);
xor XOR2 (N2702, N2700, N1409);
nand NAND2 (N2703, N2698, N2457);
nand NAND4 (N2704, N2696, N2401, N312, N507);
or OR2 (N2705, N2684, N2089);
and AND4 (N2706, N2673, N1903, N2312, N1481);
or OR3 (N2707, N2699, N1551, N2379);
or OR4 (N2708, N2705, N1445, N1395, N995);
not NOT1 (N2709, N2693);
buf BUF1 (N2710, N2703);
nand NAND3 (N2711, N2678, N708, N1972);
not NOT1 (N2712, N2708);
or OR4 (N2713, N2704, N2628, N462, N2099);
and AND3 (N2714, N2702, N1187, N1525);
nor NOR2 (N2715, N2714, N1389);
xor XOR2 (N2716, N2711, N35);
xor XOR2 (N2717, N2709, N1316);
nor NOR4 (N2718, N2716, N1703, N1278, N1262);
buf BUF1 (N2719, N2710);
buf BUF1 (N2720, N2712);
buf BUF1 (N2721, N2694);
not NOT1 (N2722, N2701);
and AND3 (N2723, N2718, N646, N401);
and AND2 (N2724, N2706, N74);
xor XOR2 (N2725, N2713, N424);
buf BUF1 (N2726, N2725);
not NOT1 (N2727, N2717);
nand NAND3 (N2728, N2724, N1146, N1162);
xor XOR2 (N2729, N2728, N2437);
xor XOR2 (N2730, N2715, N2376);
or OR4 (N2731, N2720, N733, N1584, N2340);
xor XOR2 (N2732, N2730, N1497);
or OR2 (N2733, N2723, N1622);
not NOT1 (N2734, N2707);
nor NOR3 (N2735, N2719, N2275, N1967);
buf BUF1 (N2736, N2722);
xor XOR2 (N2737, N2734, N2680);
nor NOR3 (N2738, N2726, N1221, N1989);
nand NAND2 (N2739, N2733, N1699);
not NOT1 (N2740, N2736);
nand NAND4 (N2741, N2739, N2675, N1137, N15);
and AND2 (N2742, N2735, N2448);
or OR4 (N2743, N2731, N1003, N996, N2491);
nor NOR3 (N2744, N2740, N2480, N2095);
xor XOR2 (N2745, N2744, N208);
and AND4 (N2746, N2741, N2170, N1101, N1000);
not NOT1 (N2747, N2743);
nand NAND3 (N2748, N2732, N948, N2329);
or OR2 (N2749, N2729, N1050);
xor XOR2 (N2750, N2747, N1359);
not NOT1 (N2751, N2748);
nand NAND4 (N2752, N2742, N1553, N2019, N1764);
nor NOR4 (N2753, N2737, N1998, N915, N898);
or OR3 (N2754, N2752, N1830, N941);
and AND4 (N2755, N2753, N412, N1688, N800);
or OR4 (N2756, N2746, N2653, N1036, N1031);
and AND3 (N2757, N2755, N300, N690);
nor NOR3 (N2758, N2754, N2565, N1954);
and AND3 (N2759, N2758, N2620, N103);
and AND3 (N2760, N2749, N507, N466);
buf BUF1 (N2761, N2738);
nand NAND4 (N2762, N2750, N533, N1291, N1056);
not NOT1 (N2763, N2751);
buf BUF1 (N2764, N2745);
xor XOR2 (N2765, N2759, N2691);
or OR3 (N2766, N2761, N1744, N490);
xor XOR2 (N2767, N2760, N2457);
not NOT1 (N2768, N2721);
nor NOR3 (N2769, N2768, N2603, N268);
nand NAND2 (N2770, N2766, N2362);
not NOT1 (N2771, N2762);
not NOT1 (N2772, N2770);
nor NOR2 (N2773, N2756, N2450);
nand NAND4 (N2774, N2767, N1201, N1743, N1053);
nand NAND2 (N2775, N2769, N1031);
not NOT1 (N2776, N2775);
xor XOR2 (N2777, N2765, N2464);
nor NOR2 (N2778, N2772, N2165);
buf BUF1 (N2779, N2771);
or OR4 (N2780, N2773, N674, N731, N1660);
nor NOR2 (N2781, N2780, N2179);
nand NAND2 (N2782, N2779, N1598);
or OR2 (N2783, N2763, N853);
or OR4 (N2784, N2757, N1254, N2599, N1067);
xor XOR2 (N2785, N2776, N815);
nand NAND4 (N2786, N2764, N1076, N14, N880);
buf BUF1 (N2787, N2777);
and AND4 (N2788, N2784, N1227, N776, N1369);
nor NOR4 (N2789, N2786, N1656, N1283, N2699);
not NOT1 (N2790, N2788);
buf BUF1 (N2791, N2783);
nand NAND2 (N2792, N2789, N1205);
or OR2 (N2793, N2792, N911);
not NOT1 (N2794, N2791);
buf BUF1 (N2795, N2785);
and AND3 (N2796, N2781, N741, N2345);
buf BUF1 (N2797, N2790);
nor NOR3 (N2798, N2774, N689, N1250);
nor NOR2 (N2799, N2796, N2318);
buf BUF1 (N2800, N2727);
nor NOR3 (N2801, N2795, N2246, N1061);
nand NAND3 (N2802, N2798, N1128, N1323);
xor XOR2 (N2803, N2778, N282);
and AND3 (N2804, N2794, N2617, N65);
buf BUF1 (N2805, N2787);
and AND4 (N2806, N2804, N2543, N245, N1764);
buf BUF1 (N2807, N2803);
buf BUF1 (N2808, N2807);
nand NAND2 (N2809, N2793, N1267);
nor NOR3 (N2810, N2799, N282, N661);
nor NOR2 (N2811, N2805, N1913);
nor NOR3 (N2812, N2782, N7, N2173);
or OR3 (N2813, N2812, N776, N129);
xor XOR2 (N2814, N2808, N1606);
xor XOR2 (N2815, N2813, N1328);
nor NOR2 (N2816, N2811, N2714);
xor XOR2 (N2817, N2809, N1179);
buf BUF1 (N2818, N2800);
and AND3 (N2819, N2801, N2172, N2143);
buf BUF1 (N2820, N2797);
and AND2 (N2821, N2814, N479);
xor XOR2 (N2822, N2817, N2680);
nor NOR4 (N2823, N2822, N2236, N1203, N791);
buf BUF1 (N2824, N2818);
nand NAND2 (N2825, N2802, N1562);
buf BUF1 (N2826, N2816);
xor XOR2 (N2827, N2823, N930);
or OR3 (N2828, N2820, N2564, N2257);
buf BUF1 (N2829, N2815);
nor NOR3 (N2830, N2824, N1509, N667);
xor XOR2 (N2831, N2819, N1303);
nand NAND4 (N2832, N2825, N1154, N1509, N785);
xor XOR2 (N2833, N2827, N729);
not NOT1 (N2834, N2832);
nor NOR4 (N2835, N2828, N121, N2038, N1920);
not NOT1 (N2836, N2829);
nand NAND3 (N2837, N2834, N115, N28);
nand NAND4 (N2838, N2836, N482, N2192, N942);
and AND4 (N2839, N2838, N655, N2333, N342);
nor NOR2 (N2840, N2821, N2234);
and AND3 (N2841, N2835, N806, N941);
and AND3 (N2842, N2810, N657, N1947);
nand NAND4 (N2843, N2831, N1399, N816, N768);
not NOT1 (N2844, N2833);
xor XOR2 (N2845, N2843, N936);
and AND4 (N2846, N2840, N1163, N105, N502);
and AND2 (N2847, N2830, N616);
not NOT1 (N2848, N2837);
nand NAND3 (N2849, N2806, N2204, N985);
or OR4 (N2850, N2839, N427, N1947, N1410);
not NOT1 (N2851, N2826);
not NOT1 (N2852, N2842);
buf BUF1 (N2853, N2845);
or OR4 (N2854, N2847, N1608, N2332, N1528);
buf BUF1 (N2855, N2850);
not NOT1 (N2856, N2851);
not NOT1 (N2857, N2846);
nand NAND2 (N2858, N2856, N2188);
xor XOR2 (N2859, N2844, N2083);
or OR4 (N2860, N2849, N2169, N461, N2280);
and AND4 (N2861, N2852, N78, N745, N2632);
and AND2 (N2862, N2861, N2017);
nand NAND4 (N2863, N2855, N401, N2319, N454);
or OR2 (N2864, N2858, N1820);
buf BUF1 (N2865, N2864);
not NOT1 (N2866, N2865);
nor NOR3 (N2867, N2860, N2818, N111);
buf BUF1 (N2868, N2862);
xor XOR2 (N2869, N2866, N749);
not NOT1 (N2870, N2869);
xor XOR2 (N2871, N2857, N368);
not NOT1 (N2872, N2871);
and AND4 (N2873, N2859, N533, N282, N554);
xor XOR2 (N2874, N2868, N2364);
not NOT1 (N2875, N2854);
nand NAND3 (N2876, N2867, N163, N2269);
or OR3 (N2877, N2841, N302, N64);
and AND4 (N2878, N2853, N667, N2043, N760);
or OR4 (N2879, N2870, N1198, N1592, N1222);
and AND4 (N2880, N2879, N1264, N2417, N1921);
or OR3 (N2881, N2863, N1819, N1282);
nand NAND2 (N2882, N2872, N2216);
nand NAND4 (N2883, N2880, N2583, N324, N2387);
not NOT1 (N2884, N2875);
xor XOR2 (N2885, N2873, N2841);
nor NOR3 (N2886, N2882, N2821, N1664);
or OR2 (N2887, N2881, N2667);
buf BUF1 (N2888, N2885);
not NOT1 (N2889, N2886);
nor NOR2 (N2890, N2876, N1942);
nor NOR2 (N2891, N2888, N2027);
not NOT1 (N2892, N2889);
not NOT1 (N2893, N2883);
xor XOR2 (N2894, N2878, N1060);
not NOT1 (N2895, N2890);
xor XOR2 (N2896, N2874, N625);
buf BUF1 (N2897, N2893);
buf BUF1 (N2898, N2892);
nor NOR3 (N2899, N2898, N2405, N2566);
nor NOR4 (N2900, N2894, N2622, N1624, N410);
buf BUF1 (N2901, N2900);
nand NAND4 (N2902, N2896, N2421, N2818, N520);
buf BUF1 (N2903, N2897);
not NOT1 (N2904, N2877);
and AND3 (N2905, N2904, N1798, N2790);
buf BUF1 (N2906, N2899);
or OR4 (N2907, N2891, N2031, N949, N2413);
nand NAND3 (N2908, N2903, N336, N1468);
or OR2 (N2909, N2848, N2576);
xor XOR2 (N2910, N2884, N2462);
buf BUF1 (N2911, N2902);
xor XOR2 (N2912, N2911, N1499);
buf BUF1 (N2913, N2901);
not NOT1 (N2914, N2910);
nor NOR2 (N2915, N2905, N690);
or OR2 (N2916, N2912, N2088);
not NOT1 (N2917, N2907);
or OR4 (N2918, N2908, N1913, N900, N1135);
nor NOR3 (N2919, N2895, N2476, N256);
not NOT1 (N2920, N2909);
not NOT1 (N2921, N2887);
nor NOR3 (N2922, N2915, N91, N2649);
nand NAND4 (N2923, N2919, N2567, N1402, N158);
and AND4 (N2924, N2923, N2057, N1996, N512);
nor NOR2 (N2925, N2906, N2481);
nor NOR2 (N2926, N2914, N1607);
not NOT1 (N2927, N2922);
nor NOR4 (N2928, N2916, N1778, N2533, N2489);
nand NAND4 (N2929, N2924, N1778, N591, N2441);
xor XOR2 (N2930, N2929, N340);
buf BUF1 (N2931, N2925);
or OR4 (N2932, N2918, N1964, N884, N1657);
or OR2 (N2933, N2928, N1652);
buf BUF1 (N2934, N2932);
nand NAND2 (N2935, N2927, N2768);
nor NOR4 (N2936, N2934, N439, N2620, N2695);
nand NAND3 (N2937, N2931, N1278, N567);
and AND4 (N2938, N2913, N2250, N2785, N1030);
and AND2 (N2939, N2937, N1120);
and AND4 (N2940, N2935, N2640, N2928, N1554);
or OR3 (N2941, N2930, N312, N1496);
not NOT1 (N2942, N2940);
or OR4 (N2943, N2933, N711, N477, N2199);
nand NAND2 (N2944, N2942, N1636);
nand NAND4 (N2945, N2921, N438, N2426, N14);
nor NOR2 (N2946, N2938, N753);
nand NAND2 (N2947, N2939, N1644);
nand NAND4 (N2948, N2943, N1282, N1995, N1418);
nand NAND2 (N2949, N2936, N347);
not NOT1 (N2950, N2941);
or OR3 (N2951, N2949, N2757, N366);
and AND3 (N2952, N2917, N2896, N590);
buf BUF1 (N2953, N2926);
not NOT1 (N2954, N2920);
nor NOR4 (N2955, N2948, N2126, N2127, N2006);
xor XOR2 (N2956, N2947, N1370);
buf BUF1 (N2957, N2954);
or OR3 (N2958, N2956, N1043, N1975);
buf BUF1 (N2959, N2952);
or OR2 (N2960, N2957, N2180);
buf BUF1 (N2961, N2958);
and AND2 (N2962, N2959, N938);
or OR4 (N2963, N2960, N83, N1931, N1964);
and AND3 (N2964, N2955, N2253, N1837);
nor NOR4 (N2965, N2964, N2702, N2286, N363);
buf BUF1 (N2966, N2965);
buf BUF1 (N2967, N2963);
or OR4 (N2968, N2946, N1954, N805, N1274);
or OR3 (N2969, N2966, N1375, N1337);
nor NOR2 (N2970, N2944, N484);
or OR2 (N2971, N2969, N1054);
xor XOR2 (N2972, N2968, N439);
buf BUF1 (N2973, N2971);
xor XOR2 (N2974, N2951, N2808);
xor XOR2 (N2975, N2961, N1890);
or OR2 (N2976, N2967, N969);
not NOT1 (N2977, N2953);
buf BUF1 (N2978, N2976);
not NOT1 (N2979, N2973);
and AND2 (N2980, N2972, N2664);
buf BUF1 (N2981, N2978);
nor NOR4 (N2982, N2980, N469, N2729, N1074);
nand NAND4 (N2983, N2977, N618, N1196, N1599);
xor XOR2 (N2984, N2981, N1324);
and AND4 (N2985, N2982, N1438, N1762, N1386);
nor NOR4 (N2986, N2974, N2374, N2281, N2413);
or OR2 (N2987, N2975, N2672);
nand NAND2 (N2988, N2970, N189);
or OR4 (N2989, N2987, N2526, N1115, N1678);
and AND2 (N2990, N2945, N810);
or OR4 (N2991, N2962, N2959, N1123, N2160);
nand NAND4 (N2992, N2990, N2801, N1940, N1580);
nand NAND4 (N2993, N2991, N395, N440, N2747);
and AND4 (N2994, N2988, N729, N2702, N2445);
not NOT1 (N2995, N2992);
not NOT1 (N2996, N2986);
and AND2 (N2997, N2984, N2206);
or OR3 (N2998, N2995, N123, N2547);
nor NOR4 (N2999, N2998, N21, N504, N2079);
buf BUF1 (N3000, N2950);
and AND4 (N3001, N2993, N1334, N642, N668);
xor XOR2 (N3002, N2999, N1688);
buf BUF1 (N3003, N3000);
buf BUF1 (N3004, N2989);
nor NOR4 (N3005, N3003, N483, N262, N2845);
not NOT1 (N3006, N3001);
xor XOR2 (N3007, N3002, N2742);
nand NAND4 (N3008, N2996, N2337, N2690, N1518);
xor XOR2 (N3009, N3007, N2198);
not NOT1 (N3010, N2983);
and AND4 (N3011, N2985, N1515, N1756, N425);
not NOT1 (N3012, N3004);
xor XOR2 (N3013, N3009, N2209);
buf BUF1 (N3014, N2997);
nand NAND2 (N3015, N3005, N377);
and AND4 (N3016, N3012, N722, N2998, N1270);
or OR4 (N3017, N3015, N2090, N39, N1671);
nand NAND3 (N3018, N3017, N1728, N2878);
buf BUF1 (N3019, N3016);
and AND4 (N3020, N3006, N896, N568, N2967);
and AND2 (N3021, N3019, N578);
nand NAND3 (N3022, N3013, N1712, N141);
not NOT1 (N3023, N3014);
not NOT1 (N3024, N3018);
nor NOR4 (N3025, N3008, N340, N1036, N144);
and AND2 (N3026, N2979, N1487);
nor NOR2 (N3027, N3025, N2252);
nor NOR4 (N3028, N3027, N2678, N1877, N1133);
buf BUF1 (N3029, N2994);
or OR2 (N3030, N3011, N1315);
buf BUF1 (N3031, N3030);
nor NOR3 (N3032, N3023, N1482, N1832);
or OR3 (N3033, N3021, N598, N2202);
and AND3 (N3034, N3010, N1035, N51);
buf BUF1 (N3035, N3020);
xor XOR2 (N3036, N3029, N2380);
nor NOR2 (N3037, N3024, N35);
buf BUF1 (N3038, N3033);
or OR4 (N3039, N3026, N1804, N1266, N1283);
buf BUF1 (N3040, N3022);
and AND3 (N3041, N3036, N534, N3009);
not NOT1 (N3042, N3034);
nor NOR3 (N3043, N3038, N694, N3011);
nand NAND3 (N3044, N3042, N368, N365);
or OR2 (N3045, N3031, N1146);
buf BUF1 (N3046, N3040);
xor XOR2 (N3047, N3037, N2894);
not NOT1 (N3048, N3032);
xor XOR2 (N3049, N3047, N1606);
nand NAND4 (N3050, N3043, N587, N414, N2955);
and AND3 (N3051, N3028, N2805, N137);
nor NOR4 (N3052, N3044, N1569, N319, N2759);
not NOT1 (N3053, N3049);
not NOT1 (N3054, N3052);
or OR4 (N3055, N3050, N1164, N2286, N3030);
xor XOR2 (N3056, N3045, N283);
xor XOR2 (N3057, N3046, N1044);
nor NOR4 (N3058, N3053, N316, N2077, N1148);
and AND4 (N3059, N3058, N488, N115, N2369);
and AND3 (N3060, N3055, N2514, N698);
not NOT1 (N3061, N3035);
xor XOR2 (N3062, N3051, N2778);
and AND2 (N3063, N3048, N2758);
buf BUF1 (N3064, N3062);
buf BUF1 (N3065, N3041);
nand NAND2 (N3066, N3064, N2029);
buf BUF1 (N3067, N3056);
not NOT1 (N3068, N3065);
not NOT1 (N3069, N3061);
not NOT1 (N3070, N3054);
nor NOR3 (N3071, N3057, N3011, N1321);
xor XOR2 (N3072, N3063, N41);
not NOT1 (N3073, N3059);
nand NAND4 (N3074, N3069, N689, N545, N942);
and AND3 (N3075, N3072, N2957, N291);
not NOT1 (N3076, N3070);
nand NAND4 (N3077, N3074, N1570, N1532, N2797);
nor NOR2 (N3078, N3071, N2133);
nor NOR2 (N3079, N3075, N240);
and AND2 (N3080, N3077, N803);
or OR3 (N3081, N3073, N2080, N355);
or OR2 (N3082, N3060, N1214);
nand NAND4 (N3083, N3082, N1805, N2855, N907);
not NOT1 (N3084, N3066);
nand NAND2 (N3085, N3067, N2562);
xor XOR2 (N3086, N3085, N649);
and AND3 (N3087, N3079, N2979, N1405);
and AND3 (N3088, N3076, N2334, N485);
xor XOR2 (N3089, N3086, N721);
not NOT1 (N3090, N3084);
not NOT1 (N3091, N3080);
and AND3 (N3092, N3083, N2930, N1800);
not NOT1 (N3093, N3089);
not NOT1 (N3094, N3068);
not NOT1 (N3095, N3088);
buf BUF1 (N3096, N3094);
nor NOR4 (N3097, N3096, N720, N221, N2374);
xor XOR2 (N3098, N3090, N2791);
nand NAND3 (N3099, N3095, N1293, N2175);
buf BUF1 (N3100, N3087);
xor XOR2 (N3101, N3091, N2907);
not NOT1 (N3102, N3099);
nor NOR2 (N3103, N3098, N1254);
xor XOR2 (N3104, N3100, N2255);
not NOT1 (N3105, N3101);
not NOT1 (N3106, N3081);
and AND4 (N3107, N3039, N1577, N1661, N15);
and AND2 (N3108, N3107, N118);
xor XOR2 (N3109, N3092, N1920);
nor NOR4 (N3110, N3078, N1328, N1822, N1445);
xor XOR2 (N3111, N3104, N1471);
nor NOR3 (N3112, N3110, N150, N896);
buf BUF1 (N3113, N3108);
nor NOR2 (N3114, N3097, N2847);
or OR2 (N3115, N3109, N1929);
not NOT1 (N3116, N3115);
xor XOR2 (N3117, N3112, N2706);
nor NOR2 (N3118, N3116, N565);
xor XOR2 (N3119, N3114, N2474);
nor NOR4 (N3120, N3111, N1370, N2210, N743);
or OR4 (N3121, N3120, N3120, N1556, N972);
nand NAND4 (N3122, N3106, N2017, N995, N2244);
xor XOR2 (N3123, N3102, N73);
and AND2 (N3124, N3119, N32);
or OR4 (N3125, N3122, N1076, N2720, N1156);
nand NAND3 (N3126, N3105, N2645, N317);
buf BUF1 (N3127, N3124);
nand NAND4 (N3128, N3093, N2553, N2731, N1859);
nor NOR3 (N3129, N3123, N2822, N440);
not NOT1 (N3130, N3121);
nand NAND4 (N3131, N3118, N424, N2850, N2429);
nand NAND3 (N3132, N3103, N1031, N236);
not NOT1 (N3133, N3127);
nor NOR2 (N3134, N3128, N2874);
nand NAND2 (N3135, N3117, N1276);
buf BUF1 (N3136, N3125);
and AND2 (N3137, N3134, N2917);
nand NAND2 (N3138, N3137, N238);
nand NAND2 (N3139, N3129, N2118);
buf BUF1 (N3140, N3126);
or OR3 (N3141, N3113, N1901, N2175);
nor NOR2 (N3142, N3130, N71);
and AND2 (N3143, N3135, N2257);
or OR4 (N3144, N3139, N3111, N38, N1380);
and AND3 (N3145, N3141, N49, N1453);
and AND3 (N3146, N3133, N3037, N1313);
and AND2 (N3147, N3138, N1394);
and AND2 (N3148, N3140, N202);
or OR2 (N3149, N3146, N2077);
not NOT1 (N3150, N3136);
xor XOR2 (N3151, N3145, N2218);
not NOT1 (N3152, N3132);
buf BUF1 (N3153, N3131);
nor NOR4 (N3154, N3147, N367, N1872, N1680);
and AND2 (N3155, N3154, N2414);
nor NOR3 (N3156, N3155, N1911, N2466);
not NOT1 (N3157, N3144);
or OR2 (N3158, N3142, N2802);
nand NAND3 (N3159, N3149, N2722, N2700);
and AND2 (N3160, N3148, N1778);
buf BUF1 (N3161, N3157);
buf BUF1 (N3162, N3156);
xor XOR2 (N3163, N3143, N2705);
nand NAND3 (N3164, N3152, N249, N1308);
xor XOR2 (N3165, N3159, N970);
nor NOR4 (N3166, N3160, N411, N3, N3107);
nor NOR2 (N3167, N3166, N2928);
not NOT1 (N3168, N3150);
buf BUF1 (N3169, N3158);
not NOT1 (N3170, N3164);
nand NAND4 (N3171, N3161, N2594, N2736, N1932);
and AND2 (N3172, N3168, N1406);
not NOT1 (N3173, N3171);
nor NOR4 (N3174, N3167, N7, N611, N579);
or OR4 (N3175, N3162, N2624, N730, N2956);
xor XOR2 (N3176, N3172, N3118);
buf BUF1 (N3177, N3170);
not NOT1 (N3178, N3165);
nand NAND4 (N3179, N3177, N2411, N1700, N2327);
nand NAND4 (N3180, N3169, N3134, N2536, N671);
nand NAND3 (N3181, N3179, N18, N1862);
xor XOR2 (N3182, N3173, N2887);
xor XOR2 (N3183, N3153, N439);
nand NAND3 (N3184, N3182, N1568, N8);
nor NOR2 (N3185, N3181, N2086);
not NOT1 (N3186, N3185);
nand NAND2 (N3187, N3184, N599);
buf BUF1 (N3188, N3186);
and AND4 (N3189, N3187, N719, N2718, N1191);
buf BUF1 (N3190, N3174);
nor NOR4 (N3191, N3175, N2116, N646, N1056);
not NOT1 (N3192, N3163);
not NOT1 (N3193, N3191);
buf BUF1 (N3194, N3183);
nor NOR3 (N3195, N3188, N1128, N1150);
buf BUF1 (N3196, N3180);
nand NAND3 (N3197, N3189, N2317, N1448);
nand NAND2 (N3198, N3190, N530);
nor NOR4 (N3199, N3194, N830, N240, N2525);
and AND4 (N3200, N3197, N961, N345, N2620);
nand NAND3 (N3201, N3199, N2470, N2586);
buf BUF1 (N3202, N3193);
nor NOR2 (N3203, N3196, N3086);
buf BUF1 (N3204, N3201);
and AND4 (N3205, N3204, N865, N1559, N1199);
or OR4 (N3206, N3200, N89, N2223, N1803);
or OR2 (N3207, N3195, N296);
or OR4 (N3208, N3207, N65, N233, N1123);
nor NOR3 (N3209, N3176, N1397, N1193);
nor NOR4 (N3210, N3208, N414, N2446, N322);
nand NAND3 (N3211, N3210, N2869, N2320);
not NOT1 (N3212, N3151);
nor NOR3 (N3213, N3211, N2334, N1002);
not NOT1 (N3214, N3198);
and AND4 (N3215, N3205, N2856, N1420, N583);
buf BUF1 (N3216, N3192);
not NOT1 (N3217, N3203);
nor NOR2 (N3218, N3217, N2056);
nor NOR4 (N3219, N3216, N42, N2985, N457);
or OR3 (N3220, N3202, N1588, N819);
nor NOR2 (N3221, N3219, N2615);
buf BUF1 (N3222, N3215);
not NOT1 (N3223, N3206);
and AND4 (N3224, N3223, N514, N3158, N1624);
or OR3 (N3225, N3212, N2111, N576);
not NOT1 (N3226, N3224);
nand NAND2 (N3227, N3218, N332);
nand NAND4 (N3228, N3222, N1372, N3141, N2812);
nand NAND2 (N3229, N3214, N1208);
not NOT1 (N3230, N3225);
nand NAND3 (N3231, N3213, N657, N977);
nand NAND4 (N3232, N3226, N718, N959, N652);
buf BUF1 (N3233, N3231);
nor NOR3 (N3234, N3233, N1125, N2012);
nor NOR3 (N3235, N3230, N1438, N76);
nor NOR2 (N3236, N3221, N588);
and AND3 (N3237, N3227, N1031, N1531);
or OR3 (N3238, N3228, N2397, N2084);
and AND4 (N3239, N3236, N2248, N2352, N357);
nor NOR4 (N3240, N3232, N1345, N726, N432);
nor NOR3 (N3241, N3220, N1039, N2367);
nor NOR4 (N3242, N3239, N22, N1246, N1182);
or OR3 (N3243, N3241, N1048, N1446);
xor XOR2 (N3244, N3229, N88);
nand NAND3 (N3245, N3244, N2356, N716);
not NOT1 (N3246, N3178);
nand NAND4 (N3247, N3245, N2236, N2722, N1698);
nor NOR4 (N3248, N3242, N3199, N1848, N2044);
nand NAND2 (N3249, N3209, N578);
not NOT1 (N3250, N3249);
or OR3 (N3251, N3250, N152, N1267);
not NOT1 (N3252, N3240);
buf BUF1 (N3253, N3251);
xor XOR2 (N3254, N3235, N1313);
nor NOR4 (N3255, N3252, N2779, N3017, N66);
not NOT1 (N3256, N3246);
and AND4 (N3257, N3256, N2511, N1848, N1503);
or OR2 (N3258, N3248, N1162);
nor NOR4 (N3259, N3257, N3082, N1475, N2072);
not NOT1 (N3260, N3258);
nor NOR2 (N3261, N3260, N960);
and AND3 (N3262, N3243, N378, N78);
xor XOR2 (N3263, N3261, N3231);
nor NOR2 (N3264, N3262, N3256);
not NOT1 (N3265, N3255);
nand NAND2 (N3266, N3265, N1008);
and AND2 (N3267, N3263, N1330);
nand NAND4 (N3268, N3254, N2470, N2356, N195);
nor NOR4 (N3269, N3253, N2920, N2665, N497);
and AND2 (N3270, N3237, N996);
xor XOR2 (N3271, N3259, N3046);
nor NOR3 (N3272, N3264, N791, N416);
or OR4 (N3273, N3266, N2843, N945, N94);
nand NAND3 (N3274, N3268, N1933, N1850);
buf BUF1 (N3275, N3273);
not NOT1 (N3276, N3270);
xor XOR2 (N3277, N3267, N1280);
not NOT1 (N3278, N3269);
and AND2 (N3279, N3277, N583);
nand NAND3 (N3280, N3274, N2006, N1362);
not NOT1 (N3281, N3272);
not NOT1 (N3282, N3234);
buf BUF1 (N3283, N3280);
xor XOR2 (N3284, N3278, N434);
not NOT1 (N3285, N3247);
buf BUF1 (N3286, N3284);
or OR3 (N3287, N3279, N3140, N1071);
buf BUF1 (N3288, N3283);
nand NAND2 (N3289, N3276, N2415);
not NOT1 (N3290, N3275);
or OR4 (N3291, N3290, N889, N1922, N2324);
buf BUF1 (N3292, N3287);
nor NOR3 (N3293, N3285, N1638, N2761);
or OR4 (N3294, N3282, N758, N2697, N1286);
buf BUF1 (N3295, N3292);
nor NOR4 (N3296, N3238, N1055, N852, N2623);
nand NAND2 (N3297, N3288, N2455);
not NOT1 (N3298, N3281);
or OR3 (N3299, N3298, N2718, N2358);
or OR3 (N3300, N3299, N2091, N2215);
and AND4 (N3301, N3271, N2902, N259, N1292);
and AND2 (N3302, N3291, N2366);
xor XOR2 (N3303, N3286, N1816);
buf BUF1 (N3304, N3296);
and AND2 (N3305, N3301, N2297);
and AND3 (N3306, N3289, N2261, N3253);
nor NOR2 (N3307, N3305, N1198);
nand NAND4 (N3308, N3303, N2683, N791, N1389);
not NOT1 (N3309, N3297);
xor XOR2 (N3310, N3295, N2193);
nor NOR3 (N3311, N3307, N1012, N257);
buf BUF1 (N3312, N3304);
xor XOR2 (N3313, N3294, N2906);
and AND4 (N3314, N3309, N859, N2101, N489);
not NOT1 (N3315, N3293);
buf BUF1 (N3316, N3306);
and AND3 (N3317, N3300, N3107, N2192);
not NOT1 (N3318, N3308);
nor NOR4 (N3319, N3302, N274, N141, N759);
or OR2 (N3320, N3311, N159);
nor NOR3 (N3321, N3310, N1414, N289);
xor XOR2 (N3322, N3314, N1968);
nor NOR2 (N3323, N3322, N117);
or OR2 (N3324, N3316, N1435);
buf BUF1 (N3325, N3313);
not NOT1 (N3326, N3324);
and AND4 (N3327, N3319, N3275, N954, N2888);
buf BUF1 (N3328, N3327);
and AND3 (N3329, N3318, N3143, N2351);
xor XOR2 (N3330, N3329, N487);
nor NOR3 (N3331, N3321, N2317, N2260);
and AND4 (N3332, N3326, N472, N3280, N703);
or OR2 (N3333, N3325, N772);
not NOT1 (N3334, N3312);
nand NAND4 (N3335, N3331, N2212, N2181, N1551);
not NOT1 (N3336, N3335);
xor XOR2 (N3337, N3328, N3127);
xor XOR2 (N3338, N3332, N708);
buf BUF1 (N3339, N3336);
nor NOR3 (N3340, N3330, N899, N2965);
nand NAND2 (N3341, N3315, N885);
or OR3 (N3342, N3320, N1135, N1625);
xor XOR2 (N3343, N3334, N1807);
and AND4 (N3344, N3337, N641, N1177, N601);
or OR3 (N3345, N3341, N639, N1113);
nand NAND4 (N3346, N3340, N3213, N2416, N644);
xor XOR2 (N3347, N3317, N714);
or OR2 (N3348, N3342, N2738);
nand NAND2 (N3349, N3347, N462);
nand NAND3 (N3350, N3339, N2025, N2759);
nand NAND2 (N3351, N3323, N392);
or OR3 (N3352, N3338, N1954, N3199);
buf BUF1 (N3353, N3344);
buf BUF1 (N3354, N3333);
xor XOR2 (N3355, N3352, N1008);
nor NOR2 (N3356, N3345, N2685);
and AND4 (N3357, N3350, N1355, N1443, N1411);
or OR4 (N3358, N3357, N1275, N1048, N1719);
buf BUF1 (N3359, N3349);
xor XOR2 (N3360, N3346, N2092);
nor NOR3 (N3361, N3354, N2722, N458);
buf BUF1 (N3362, N3356);
and AND4 (N3363, N3362, N1315, N2204, N1361);
or OR2 (N3364, N3361, N2067);
and AND3 (N3365, N3348, N1407, N1594);
buf BUF1 (N3366, N3355);
nor NOR3 (N3367, N3364, N1004, N464);
buf BUF1 (N3368, N3353);
nand NAND4 (N3369, N3368, N6, N2541, N3185);
nand NAND4 (N3370, N3365, N1871, N2786, N1858);
not NOT1 (N3371, N3351);
not NOT1 (N3372, N3367);
buf BUF1 (N3373, N3370);
xor XOR2 (N3374, N3372, N3353);
or OR2 (N3375, N3343, N1062);
buf BUF1 (N3376, N3358);
or OR2 (N3377, N3359, N1691);
not NOT1 (N3378, N3369);
not NOT1 (N3379, N3377);
or OR2 (N3380, N3360, N1233);
buf BUF1 (N3381, N3378);
buf BUF1 (N3382, N3376);
nand NAND3 (N3383, N3363, N2417, N2614);
and AND2 (N3384, N3380, N1056);
and AND4 (N3385, N3381, N328, N1113, N3247);
not NOT1 (N3386, N3385);
and AND2 (N3387, N3386, N221);
xor XOR2 (N3388, N3384, N1818);
nand NAND4 (N3389, N3382, N3340, N2749, N2177);
and AND3 (N3390, N3388, N966, N2911);
or OR2 (N3391, N3366, N3358);
or OR3 (N3392, N3390, N1133, N2558);
nand NAND2 (N3393, N3371, N1055);
not NOT1 (N3394, N3374);
or OR3 (N3395, N3375, N2894, N2687);
xor XOR2 (N3396, N3391, N2759);
and AND4 (N3397, N3387, N213, N198, N2934);
and AND3 (N3398, N3394, N1028, N2998);
or OR3 (N3399, N3373, N1603, N1530);
nand NAND2 (N3400, N3396, N2751);
buf BUF1 (N3401, N3383);
nor NOR2 (N3402, N3389, N2250);
and AND3 (N3403, N3392, N2450, N2508);
xor XOR2 (N3404, N3395, N307);
nor NOR4 (N3405, N3400, N1164, N2523, N2435);
or OR3 (N3406, N3404, N2655, N3095);
xor XOR2 (N3407, N3379, N1639);
xor XOR2 (N3408, N3397, N2505);
nand NAND3 (N3409, N3405, N3349, N1838);
buf BUF1 (N3410, N3406);
nor NOR2 (N3411, N3401, N1064);
nand NAND3 (N3412, N3398, N3177, N2941);
nor NOR2 (N3413, N3399, N1626);
nor NOR3 (N3414, N3407, N1884, N1914);
nor NOR4 (N3415, N3414, N1437, N2845, N2543);
xor XOR2 (N3416, N3412, N1499);
buf BUF1 (N3417, N3402);
buf BUF1 (N3418, N3411);
xor XOR2 (N3419, N3413, N961);
xor XOR2 (N3420, N3417, N3414);
and AND2 (N3421, N3410, N1204);
not NOT1 (N3422, N3419);
buf BUF1 (N3423, N3420);
xor XOR2 (N3424, N3393, N514);
xor XOR2 (N3425, N3408, N10);
or OR4 (N3426, N3422, N694, N480, N155);
or OR3 (N3427, N3416, N2209, N1272);
xor XOR2 (N3428, N3418, N2785);
nor NOR3 (N3429, N3424, N111, N1728);
buf BUF1 (N3430, N3421);
or OR2 (N3431, N3425, N1270);
and AND2 (N3432, N3429, N3047);
not NOT1 (N3433, N3423);
nand NAND4 (N3434, N3431, N3416, N2745, N3070);
xor XOR2 (N3435, N3432, N2700);
and AND2 (N3436, N3430, N582);
buf BUF1 (N3437, N3433);
xor XOR2 (N3438, N3435, N128);
buf BUF1 (N3439, N3409);
or OR2 (N3440, N3439, N2693);
xor XOR2 (N3441, N3427, N1583);
or OR4 (N3442, N3403, N759, N968, N922);
buf BUF1 (N3443, N3438);
nand NAND4 (N3444, N3415, N1778, N445, N2321);
and AND3 (N3445, N3426, N1128, N1808);
nor NOR2 (N3446, N3443, N2161);
or OR2 (N3447, N3445, N260);
nor NOR3 (N3448, N3442, N2822, N2003);
and AND3 (N3449, N3434, N2424, N1150);
xor XOR2 (N3450, N3437, N2102);
buf BUF1 (N3451, N3436);
and AND3 (N3452, N3448, N3143, N2232);
nor NOR4 (N3453, N3446, N3015, N2824, N985);
nor NOR3 (N3454, N3428, N1876, N528);
nor NOR2 (N3455, N3440, N266);
buf BUF1 (N3456, N3449);
or OR3 (N3457, N3441, N173, N2808);
or OR2 (N3458, N3450, N2978);
buf BUF1 (N3459, N3453);
or OR4 (N3460, N3451, N1603, N2918, N1733);
buf BUF1 (N3461, N3457);
and AND3 (N3462, N3458, N2016, N332);
xor XOR2 (N3463, N3455, N552);
xor XOR2 (N3464, N3454, N2174);
or OR3 (N3465, N3461, N2352, N985);
xor XOR2 (N3466, N3444, N3086);
or OR4 (N3467, N3452, N2224, N1536, N3460);
xor XOR2 (N3468, N1443, N389);
nand NAND4 (N3469, N3447, N1451, N123, N3000);
xor XOR2 (N3470, N3468, N265);
nand NAND3 (N3471, N3466, N494, N274);
not NOT1 (N3472, N3470);
or OR2 (N3473, N3465, N2919);
xor XOR2 (N3474, N3459, N897);
or OR4 (N3475, N3462, N1790, N1592, N3407);
nand NAND4 (N3476, N3474, N284, N504, N1992);
nand NAND4 (N3477, N3475, N2428, N690, N2751);
nor NOR4 (N3478, N3472, N1834, N2273, N738);
xor XOR2 (N3479, N3476, N31);
xor XOR2 (N3480, N3477, N197);
buf BUF1 (N3481, N3471);
nand NAND4 (N3482, N3464, N62, N2926, N3226);
or OR2 (N3483, N3456, N2735);
not NOT1 (N3484, N3479);
buf BUF1 (N3485, N3483);
and AND2 (N3486, N3484, N2137);
xor XOR2 (N3487, N3480, N3396);
xor XOR2 (N3488, N3487, N2731);
buf BUF1 (N3489, N3486);
xor XOR2 (N3490, N3469, N1567);
or OR4 (N3491, N3478, N3132, N2916, N70);
xor XOR2 (N3492, N3463, N2847);
not NOT1 (N3493, N3490);
xor XOR2 (N3494, N3485, N1649);
nand NAND4 (N3495, N3473, N268, N2771, N341);
and AND3 (N3496, N3494, N1068, N1308);
nand NAND2 (N3497, N3493, N3255);
or OR2 (N3498, N3491, N3212);
buf BUF1 (N3499, N3498);
nor NOR2 (N3500, N3492, N1215);
buf BUF1 (N3501, N3495);
xor XOR2 (N3502, N3467, N1776);
or OR2 (N3503, N3488, N1129);
buf BUF1 (N3504, N3481);
nor NOR3 (N3505, N3489, N2105, N1926);
nand NAND3 (N3506, N3497, N2438, N3218);
xor XOR2 (N3507, N3496, N547);
buf BUF1 (N3508, N3505);
or OR4 (N3509, N3482, N2461, N550, N3089);
nand NAND4 (N3510, N3509, N704, N2918, N1044);
or OR4 (N3511, N3503, N261, N1589, N3115);
buf BUF1 (N3512, N3500);
buf BUF1 (N3513, N3507);
not NOT1 (N3514, N3502);
nand NAND2 (N3515, N3510, N2230);
or OR3 (N3516, N3504, N1125, N87);
nor NOR3 (N3517, N3514, N179, N958);
nand NAND3 (N3518, N3499, N2147, N675);
not NOT1 (N3519, N3512);
not NOT1 (N3520, N3501);
buf BUF1 (N3521, N3517);
or OR3 (N3522, N3516, N1089, N752);
nand NAND2 (N3523, N3521, N2281);
nand NAND4 (N3524, N3518, N2693, N2669, N3061);
nor NOR2 (N3525, N3513, N2496);
and AND4 (N3526, N3520, N2503, N2409, N1003);
nor NOR4 (N3527, N3511, N1794, N770, N3476);
or OR3 (N3528, N3527, N2631, N1070);
nand NAND4 (N3529, N3523, N1062, N2579, N1598);
and AND2 (N3530, N3515, N3492);
or OR3 (N3531, N3529, N85, N1680);
or OR2 (N3532, N3525, N703);
buf BUF1 (N3533, N3508);
and AND3 (N3534, N3531, N3273, N3112);
nor NOR2 (N3535, N3532, N705);
not NOT1 (N3536, N3535);
nand NAND2 (N3537, N3524, N1234);
and AND2 (N3538, N3506, N3070);
buf BUF1 (N3539, N3534);
or OR2 (N3540, N3536, N802);
or OR3 (N3541, N3540, N289, N1675);
nand NAND2 (N3542, N3522, N1125);
not NOT1 (N3543, N3538);
and AND2 (N3544, N3541, N1327);
or OR4 (N3545, N3539, N3338, N1840, N551);
not NOT1 (N3546, N3542);
xor XOR2 (N3547, N3544, N2735);
and AND2 (N3548, N3537, N931);
buf BUF1 (N3549, N3548);
nand NAND3 (N3550, N3547, N213, N594);
nand NAND4 (N3551, N3526, N2187, N2042, N727);
not NOT1 (N3552, N3528);
or OR3 (N3553, N3519, N205, N3134);
nand NAND3 (N3554, N3552, N678, N2800);
nor NOR2 (N3555, N3546, N3289);
buf BUF1 (N3556, N3554);
not NOT1 (N3557, N3533);
buf BUF1 (N3558, N3555);
nand NAND3 (N3559, N3550, N568, N2370);
or OR4 (N3560, N3530, N2350, N1265, N1482);
and AND2 (N3561, N3556, N2162);
xor XOR2 (N3562, N3559, N36);
buf BUF1 (N3563, N3558);
buf BUF1 (N3564, N3543);
buf BUF1 (N3565, N3564);
xor XOR2 (N3566, N3553, N3526);
buf BUF1 (N3567, N3560);
or OR4 (N3568, N3566, N1319, N2246, N785);
nand NAND4 (N3569, N3562, N3087, N1330, N1734);
nor NOR4 (N3570, N3569, N2749, N1380, N613);
xor XOR2 (N3571, N3563, N2626);
not NOT1 (N3572, N3551);
xor XOR2 (N3573, N3565, N2649);
or OR4 (N3574, N3568, N2541, N2404, N2433);
and AND3 (N3575, N3561, N3022, N2646);
nor NOR2 (N3576, N3567, N788);
nand NAND4 (N3577, N3570, N3473, N1397, N2250);
nand NAND4 (N3578, N3571, N2631, N3436, N874);
nor NOR4 (N3579, N3557, N516, N1245, N990);
nor NOR2 (N3580, N3577, N2977);
nor NOR4 (N3581, N3580, N2239, N1073, N362);
and AND2 (N3582, N3545, N2754);
nand NAND4 (N3583, N3573, N3529, N499, N2776);
nor NOR4 (N3584, N3575, N1971, N514, N386);
buf BUF1 (N3585, N3572);
or OR2 (N3586, N3579, N2275);
nor NOR3 (N3587, N3549, N3559, N1043);
or OR2 (N3588, N3582, N2051);
nand NAND4 (N3589, N3583, N1200, N1483, N568);
and AND2 (N3590, N3576, N588);
not NOT1 (N3591, N3589);
not NOT1 (N3592, N3586);
nand NAND4 (N3593, N3581, N2350, N2171, N190);
or OR2 (N3594, N3588, N1105);
or OR3 (N3595, N3578, N2964, N119);
not NOT1 (N3596, N3585);
or OR3 (N3597, N3595, N920, N1627);
or OR3 (N3598, N3596, N2712, N2288);
nor NOR4 (N3599, N3574, N1935, N3342, N1636);
nand NAND2 (N3600, N3599, N134);
nand NAND3 (N3601, N3598, N199, N1094);
and AND4 (N3602, N3592, N1292, N3495, N1415);
nand NAND3 (N3603, N3584, N3241, N2302);
xor XOR2 (N3604, N3603, N2157);
buf BUF1 (N3605, N3590);
xor XOR2 (N3606, N3594, N1299);
and AND4 (N3607, N3606, N685, N2810, N2938);
or OR4 (N3608, N3597, N3348, N308, N962);
not NOT1 (N3609, N3587);
or OR4 (N3610, N3605, N1905, N1650, N1393);
not NOT1 (N3611, N3607);
buf BUF1 (N3612, N3602);
nand NAND2 (N3613, N3611, N96);
xor XOR2 (N3614, N3609, N797);
nor NOR4 (N3615, N3593, N2110, N2145, N417);
nor NOR4 (N3616, N3613, N580, N620, N2504);
nor NOR2 (N3617, N3610, N3028);
nand NAND2 (N3618, N3615, N2317);
nor NOR3 (N3619, N3614, N411, N561);
not NOT1 (N3620, N3619);
buf BUF1 (N3621, N3601);
buf BUF1 (N3622, N3608);
nor NOR4 (N3623, N3604, N542, N1454, N1476);
nand NAND3 (N3624, N3621, N3085, N3380);
buf BUF1 (N3625, N3617);
buf BUF1 (N3626, N3623);
xor XOR2 (N3627, N3618, N3545);
or OR4 (N3628, N3626, N528, N1642, N354);
or OR2 (N3629, N3622, N1196);
nand NAND4 (N3630, N3629, N3437, N865, N2768);
buf BUF1 (N3631, N3612);
xor XOR2 (N3632, N3616, N1888);
or OR2 (N3633, N3600, N1058);
buf BUF1 (N3634, N3632);
and AND2 (N3635, N3630, N1205);
and AND4 (N3636, N3627, N1030, N2477, N1898);
buf BUF1 (N3637, N3634);
not NOT1 (N3638, N3637);
buf BUF1 (N3639, N3628);
nand NAND2 (N3640, N3636, N3530);
buf BUF1 (N3641, N3631);
buf BUF1 (N3642, N3625);
buf BUF1 (N3643, N3642);
or OR3 (N3644, N3633, N2129, N3187);
buf BUF1 (N3645, N3620);
and AND3 (N3646, N3645, N340, N1133);
nor NOR2 (N3647, N3639, N1406);
and AND2 (N3648, N3646, N3422);
and AND2 (N3649, N3638, N2053);
xor XOR2 (N3650, N3640, N1410);
and AND2 (N3651, N3643, N172);
and AND4 (N3652, N3648, N748, N709, N3569);
nand NAND2 (N3653, N3591, N986);
or OR3 (N3654, N3644, N1040, N2213);
or OR3 (N3655, N3635, N361, N888);
not NOT1 (N3656, N3649);
and AND2 (N3657, N3654, N2245);
or OR2 (N3658, N3647, N2598);
and AND2 (N3659, N3651, N1428);
not NOT1 (N3660, N3656);
nand NAND3 (N3661, N3657, N589, N188);
xor XOR2 (N3662, N3652, N1906);
or OR3 (N3663, N3661, N1560, N2465);
nor NOR4 (N3664, N3624, N2350, N897, N3294);
not NOT1 (N3665, N3658);
nand NAND2 (N3666, N3665, N778);
xor XOR2 (N3667, N3666, N3222);
and AND3 (N3668, N3667, N999, N3625);
nor NOR2 (N3669, N3660, N1486);
nand NAND2 (N3670, N3664, N1138);
nor NOR2 (N3671, N3662, N2004);
nand NAND4 (N3672, N3668, N434, N2867, N169);
xor XOR2 (N3673, N3672, N3145);
buf BUF1 (N3674, N3669);
and AND3 (N3675, N3663, N344, N2342);
and AND3 (N3676, N3653, N3378, N186);
nand NAND2 (N3677, N3641, N649);
buf BUF1 (N3678, N3650);
nor NOR2 (N3679, N3659, N2208);
nand NAND4 (N3680, N3670, N1424, N2252, N506);
nor NOR2 (N3681, N3676, N1150);
not NOT1 (N3682, N3675);
buf BUF1 (N3683, N3677);
nand NAND3 (N3684, N3655, N2220, N647);
not NOT1 (N3685, N3684);
and AND2 (N3686, N3682, N2718);
not NOT1 (N3687, N3681);
nand NAND4 (N3688, N3680, N388, N2534, N1416);
nand NAND4 (N3689, N3685, N89, N2519, N3646);
and AND4 (N3690, N3683, N3102, N186, N2572);
xor XOR2 (N3691, N3671, N2630);
nand NAND2 (N3692, N3690, N2399);
nand NAND4 (N3693, N3691, N901, N203, N2525);
nand NAND2 (N3694, N3692, N1194);
nor NOR3 (N3695, N3674, N1095, N3591);
xor XOR2 (N3696, N3673, N1573);
or OR3 (N3697, N3686, N2744, N912);
nand NAND4 (N3698, N3678, N1325, N1329, N2329);
buf BUF1 (N3699, N3698);
and AND4 (N3700, N3679, N3405, N1923, N1444);
and AND4 (N3701, N3696, N297, N2679, N2806);
buf BUF1 (N3702, N3694);
nor NOR3 (N3703, N3700, N834, N2255);
nor NOR2 (N3704, N3697, N1093);
nor NOR2 (N3705, N3699, N2981);
nand NAND4 (N3706, N3693, N113, N246, N2364);
xor XOR2 (N3707, N3689, N1300);
not NOT1 (N3708, N3695);
xor XOR2 (N3709, N3703, N2696);
nand NAND4 (N3710, N3705, N922, N167, N1949);
or OR3 (N3711, N3688, N2310, N1913);
nor NOR3 (N3712, N3701, N1209, N2831);
not NOT1 (N3713, N3706);
not NOT1 (N3714, N3710);
nor NOR4 (N3715, N3709, N3535, N829, N2226);
nor NOR4 (N3716, N3702, N2276, N1432, N3630);
xor XOR2 (N3717, N3704, N1534);
buf BUF1 (N3718, N3716);
and AND3 (N3719, N3715, N38, N2282);
not NOT1 (N3720, N3719);
not NOT1 (N3721, N3707);
buf BUF1 (N3722, N3721);
not NOT1 (N3723, N3712);
nor NOR4 (N3724, N3722, N79, N1663, N2835);
and AND3 (N3725, N3718, N3275, N3611);
or OR4 (N3726, N3723, N637, N3582, N385);
xor XOR2 (N3727, N3713, N513);
nand NAND2 (N3728, N3726, N3421);
nor NOR3 (N3729, N3728, N1094, N3600);
and AND3 (N3730, N3724, N1773, N1431);
nand NAND3 (N3731, N3729, N1639, N3419);
nand NAND3 (N3732, N3708, N311, N3546);
xor XOR2 (N3733, N3717, N3342);
not NOT1 (N3734, N3731);
nand NAND3 (N3735, N3732, N500, N1443);
and AND2 (N3736, N3733, N3663);
nor NOR3 (N3737, N3725, N1769, N240);
xor XOR2 (N3738, N3720, N291);
and AND4 (N3739, N3738, N3165, N774, N884);
buf BUF1 (N3740, N3735);
nand NAND3 (N3741, N3711, N254, N1471);
buf BUF1 (N3742, N3739);
nor NOR4 (N3743, N3687, N335, N3528, N2583);
nor NOR2 (N3744, N3740, N773);
not NOT1 (N3745, N3743);
nor NOR3 (N3746, N3736, N2449, N1041);
not NOT1 (N3747, N3741);
and AND3 (N3748, N3734, N3204, N2828);
and AND3 (N3749, N3714, N2481, N367);
xor XOR2 (N3750, N3737, N2422);
nor NOR3 (N3751, N3745, N3696, N3434);
or OR2 (N3752, N3751, N3287);
not NOT1 (N3753, N3748);
nand NAND2 (N3754, N3730, N3389);
and AND3 (N3755, N3753, N2732, N842);
not NOT1 (N3756, N3747);
buf BUF1 (N3757, N3744);
nand NAND2 (N3758, N3749, N1380);
buf BUF1 (N3759, N3757);
buf BUF1 (N3760, N3750);
nor NOR4 (N3761, N3756, N554, N2898, N1017);
or OR2 (N3762, N3760, N266);
xor XOR2 (N3763, N3758, N1067);
or OR3 (N3764, N3754, N1806, N954);
and AND2 (N3765, N3762, N3406);
and AND4 (N3766, N3764, N1688, N107, N579);
buf BUF1 (N3767, N3755);
nand NAND2 (N3768, N3742, N2488);
buf BUF1 (N3769, N3766);
nand NAND4 (N3770, N3759, N1694, N447, N2144);
or OR2 (N3771, N3727, N2281);
xor XOR2 (N3772, N3763, N521);
xor XOR2 (N3773, N3770, N2113);
not NOT1 (N3774, N3746);
not NOT1 (N3775, N3774);
not NOT1 (N3776, N3768);
or OR4 (N3777, N3775, N1373, N1010, N2564);
nand NAND2 (N3778, N3765, N2774);
or OR2 (N3779, N3777, N3451);
nand NAND4 (N3780, N3761, N2371, N615, N2517);
nor NOR2 (N3781, N3767, N2715);
not NOT1 (N3782, N3780);
buf BUF1 (N3783, N3773);
nor NOR3 (N3784, N3781, N1239, N2831);
and AND3 (N3785, N3769, N936, N2913);
nand NAND2 (N3786, N3779, N1507);
or OR4 (N3787, N3776, N3612, N3413, N3519);
nand NAND2 (N3788, N3772, N3548);
and AND2 (N3789, N3783, N692);
and AND4 (N3790, N3752, N588, N1406, N295);
buf BUF1 (N3791, N3789);
nand NAND3 (N3792, N3790, N488, N1881);
or OR3 (N3793, N3786, N1146, N373);
and AND4 (N3794, N3788, N2507, N79, N3199);
xor XOR2 (N3795, N3791, N2588);
and AND3 (N3796, N3771, N1809, N1180);
nor NOR2 (N3797, N3796, N379);
or OR3 (N3798, N3795, N2223, N2092);
xor XOR2 (N3799, N3793, N451);
not NOT1 (N3800, N3794);
xor XOR2 (N3801, N3800, N2680);
or OR3 (N3802, N3797, N3465, N3331);
not NOT1 (N3803, N3799);
nand NAND2 (N3804, N3798, N3083);
buf BUF1 (N3805, N3804);
nand NAND3 (N3806, N3785, N3705, N3139);
buf BUF1 (N3807, N3802);
nor NOR2 (N3808, N3801, N2362);
not NOT1 (N3809, N3792);
or OR4 (N3810, N3784, N1972, N165, N433);
nor NOR4 (N3811, N3809, N1799, N2677, N467);
and AND3 (N3812, N3782, N3253, N2902);
buf BUF1 (N3813, N3787);
not NOT1 (N3814, N3807);
and AND3 (N3815, N3803, N3283, N3227);
not NOT1 (N3816, N3805);
or OR4 (N3817, N3814, N2823, N2534, N3288);
and AND4 (N3818, N3778, N1946, N716, N1129);
nor NOR3 (N3819, N3806, N3594, N2769);
nand NAND3 (N3820, N3810, N1325, N975);
nand NAND3 (N3821, N3819, N2207, N3158);
nor NOR3 (N3822, N3812, N3761, N3454);
buf BUF1 (N3823, N3818);
not NOT1 (N3824, N3817);
buf BUF1 (N3825, N3820);
xor XOR2 (N3826, N3816, N1886);
not NOT1 (N3827, N3826);
nor NOR2 (N3828, N3825, N2023);
not NOT1 (N3829, N3823);
or OR4 (N3830, N3811, N2583, N867, N1440);
not NOT1 (N3831, N3827);
nand NAND2 (N3832, N3822, N2667);
or OR2 (N3833, N3831, N3016);
or OR4 (N3834, N3821, N633, N3400, N861);
or OR4 (N3835, N3830, N1148, N2480, N3371);
and AND2 (N3836, N3824, N199);
nand NAND4 (N3837, N3836, N2238, N2860, N2585);
not NOT1 (N3838, N3813);
and AND4 (N3839, N3833, N3218, N2662, N1150);
xor XOR2 (N3840, N3838, N3483);
or OR4 (N3841, N3828, N2969, N2237, N1092);
xor XOR2 (N3842, N3839, N1072);
buf BUF1 (N3843, N3829);
xor XOR2 (N3844, N3835, N1784);
buf BUF1 (N3845, N3815);
nor NOR4 (N3846, N3832, N1207, N1393, N3247);
buf BUF1 (N3847, N3808);
nor NOR4 (N3848, N3847, N3516, N636, N651);
xor XOR2 (N3849, N3834, N3823);
or OR3 (N3850, N3840, N2634, N2359);
or OR2 (N3851, N3844, N231);
and AND2 (N3852, N3843, N1680);
not NOT1 (N3853, N3845);
or OR2 (N3854, N3852, N2939);
nand NAND4 (N3855, N3850, N1074, N3554, N945);
not NOT1 (N3856, N3848);
or OR2 (N3857, N3854, N2320);
nor NOR2 (N3858, N3851, N1747);
and AND4 (N3859, N3841, N3513, N155, N713);
not NOT1 (N3860, N3859);
not NOT1 (N3861, N3858);
not NOT1 (N3862, N3855);
xor XOR2 (N3863, N3857, N2055);
nand NAND2 (N3864, N3862, N2396);
not NOT1 (N3865, N3853);
not NOT1 (N3866, N3846);
or OR3 (N3867, N3865, N2864, N1109);
and AND2 (N3868, N3856, N538);
not NOT1 (N3869, N3842);
or OR3 (N3870, N3837, N443, N1913);
nor NOR4 (N3871, N3849, N905, N1462, N2283);
buf BUF1 (N3872, N3864);
nand NAND3 (N3873, N3869, N3183, N2126);
buf BUF1 (N3874, N3863);
not NOT1 (N3875, N3861);
or OR3 (N3876, N3873, N709, N2854);
buf BUF1 (N3877, N3872);
buf BUF1 (N3878, N3874);
or OR2 (N3879, N3866, N801);
nor NOR3 (N3880, N3879, N2890, N3867);
and AND3 (N3881, N1172, N1036, N1335);
buf BUF1 (N3882, N3878);
buf BUF1 (N3883, N3868);
nand NAND4 (N3884, N3880, N2189, N492, N1713);
and AND4 (N3885, N3884, N2172, N990, N1205);
buf BUF1 (N3886, N3885);
xor XOR2 (N3887, N3860, N2490);
nand NAND3 (N3888, N3883, N1471, N3364);
nand NAND4 (N3889, N3875, N660, N116, N2305);
and AND2 (N3890, N3889, N1149);
not NOT1 (N3891, N3888);
nand NAND3 (N3892, N3876, N1798, N1603);
not NOT1 (N3893, N3882);
and AND2 (N3894, N3887, N544);
and AND2 (N3895, N3871, N259);
or OR3 (N3896, N3881, N2398, N1111);
buf BUF1 (N3897, N3886);
nor NOR3 (N3898, N3892, N3457, N1572);
nand NAND4 (N3899, N3891, N1515, N474, N1442);
buf BUF1 (N3900, N3899);
buf BUF1 (N3901, N3893);
and AND4 (N3902, N3897, N1591, N551, N2638);
buf BUF1 (N3903, N3877);
xor XOR2 (N3904, N3896, N412);
nor NOR2 (N3905, N3904, N1353);
and AND2 (N3906, N3900, N604);
and AND2 (N3907, N3870, N3151);
xor XOR2 (N3908, N3907, N2373);
not NOT1 (N3909, N3894);
xor XOR2 (N3910, N3902, N1551);
xor XOR2 (N3911, N3909, N2154);
buf BUF1 (N3912, N3910);
nand NAND4 (N3913, N3908, N3200, N1706, N2690);
nand NAND3 (N3914, N3898, N3332, N1694);
not NOT1 (N3915, N3905);
nor NOR3 (N3916, N3903, N2544, N1475);
nand NAND4 (N3917, N3914, N1633, N3481, N1162);
buf BUF1 (N3918, N3917);
nand NAND3 (N3919, N3915, N2120, N1862);
nor NOR4 (N3920, N3913, N1472, N2583, N1823);
xor XOR2 (N3921, N3916, N871);
not NOT1 (N3922, N3890);
nor NOR3 (N3923, N3920, N2969, N2649);
nor NOR4 (N3924, N3919, N1308, N825, N1174);
and AND3 (N3925, N3901, N1662, N1670);
xor XOR2 (N3926, N3924, N659);
or OR4 (N3927, N3921, N285, N2559, N1268);
xor XOR2 (N3928, N3918, N1236);
and AND2 (N3929, N3912, N2770);
or OR2 (N3930, N3927, N2862);
or OR4 (N3931, N3911, N577, N184, N3524);
and AND4 (N3932, N3925, N2891, N958, N174);
not NOT1 (N3933, N3923);
or OR4 (N3934, N3931, N32, N1455, N1634);
nand NAND4 (N3935, N3934, N162, N514, N2783);
nor NOR3 (N3936, N3930, N3397, N581);
not NOT1 (N3937, N3926);
nor NOR4 (N3938, N3932, N3080, N148, N3137);
not NOT1 (N3939, N3938);
buf BUF1 (N3940, N3928);
buf BUF1 (N3941, N3929);
and AND4 (N3942, N3937, N1102, N798, N2255);
and AND2 (N3943, N3941, N1406);
xor XOR2 (N3944, N3935, N184);
and AND2 (N3945, N3939, N3631);
not NOT1 (N3946, N3942);
and AND4 (N3947, N3946, N2720, N1872, N1097);
or OR4 (N3948, N3945, N3115, N70, N373);
xor XOR2 (N3949, N3906, N1882);
buf BUF1 (N3950, N3949);
not NOT1 (N3951, N3948);
and AND4 (N3952, N3940, N206, N622, N1169);
nor NOR2 (N3953, N3947, N2381);
nor NOR3 (N3954, N3895, N404, N1385);
and AND2 (N3955, N3953, N834);
not NOT1 (N3956, N3955);
buf BUF1 (N3957, N3951);
or OR2 (N3958, N3944, N1899);
xor XOR2 (N3959, N3958, N450);
not NOT1 (N3960, N3956);
or OR2 (N3961, N3922, N268);
nand NAND2 (N3962, N3960, N1790);
xor XOR2 (N3963, N3959, N3623);
not NOT1 (N3964, N3961);
or OR2 (N3965, N3936, N2313);
xor XOR2 (N3966, N3957, N107);
or OR2 (N3967, N3952, N3947);
nand NAND3 (N3968, N3933, N34, N2617);
nor NOR4 (N3969, N3966, N3922, N3869, N3864);
not NOT1 (N3970, N3968);
xor XOR2 (N3971, N3967, N3282);
buf BUF1 (N3972, N3965);
or OR4 (N3973, N3962, N1998, N2176, N1534);
xor XOR2 (N3974, N3950, N2363);
nand NAND3 (N3975, N3973, N2276, N2801);
or OR3 (N3976, N3969, N402, N2566);
or OR3 (N3977, N3964, N733, N1981);
not NOT1 (N3978, N3976);
xor XOR2 (N3979, N3963, N3576);
xor XOR2 (N3980, N3975, N90);
xor XOR2 (N3981, N3974, N2786);
and AND4 (N3982, N3954, N2071, N2452, N2562);
buf BUF1 (N3983, N3980);
nor NOR3 (N3984, N3983, N2337, N4);
not NOT1 (N3985, N3970);
nor NOR3 (N3986, N3982, N3665, N2306);
xor XOR2 (N3987, N3978, N91);
nor NOR2 (N3988, N3972, N3517);
not NOT1 (N3989, N3979);
not NOT1 (N3990, N3989);
buf BUF1 (N3991, N3987);
or OR2 (N3992, N3943, N436);
or OR4 (N3993, N3988, N1200, N1279, N952);
and AND4 (N3994, N3985, N1425, N3319, N52);
xor XOR2 (N3995, N3971, N711);
xor XOR2 (N3996, N3981, N988);
or OR2 (N3997, N3984, N2203);
buf BUF1 (N3998, N3995);
buf BUF1 (N3999, N3977);
not NOT1 (N4000, N3998);
or OR4 (N4001, N4000, N1724, N1364, N1067);
not NOT1 (N4002, N3993);
buf BUF1 (N4003, N3994);
buf BUF1 (N4004, N3997);
buf BUF1 (N4005, N3991);
or OR2 (N4006, N4001, N3447);
not NOT1 (N4007, N4006);
not NOT1 (N4008, N4003);
and AND2 (N4009, N3992, N1306);
xor XOR2 (N4010, N4002, N2639);
and AND2 (N4011, N4009, N2545);
not NOT1 (N4012, N4008);
nand NAND4 (N4013, N4012, N1624, N1995, N1638);
or OR3 (N4014, N4010, N141, N2924);
buf BUF1 (N4015, N4014);
xor XOR2 (N4016, N4015, N1920);
buf BUF1 (N4017, N4007);
buf BUF1 (N4018, N3999);
and AND3 (N4019, N4013, N1838, N767);
or OR3 (N4020, N4017, N2547, N2543);
buf BUF1 (N4021, N4005);
nor NOR4 (N4022, N4018, N4013, N1918, N3558);
nand NAND3 (N4023, N4020, N164, N2846);
and AND3 (N4024, N4004, N2820, N1471);
and AND4 (N4025, N4023, N3594, N2621, N1119);
xor XOR2 (N4026, N4011, N3232);
xor XOR2 (N4027, N4024, N2276);
not NOT1 (N4028, N4027);
or OR3 (N4029, N3990, N3948, N2567);
nand NAND3 (N4030, N4025, N1041, N2931);
xor XOR2 (N4031, N4028, N342);
nor NOR2 (N4032, N4022, N866);
or OR4 (N4033, N4019, N2520, N3440, N1050);
nor NOR2 (N4034, N4033, N3291);
buf BUF1 (N4035, N4016);
nor NOR3 (N4036, N4029, N3383, N1118);
buf BUF1 (N4037, N4031);
nor NOR3 (N4038, N4035, N2466, N1469);
not NOT1 (N4039, N4036);
and AND3 (N4040, N4032, N3976, N3163);
buf BUF1 (N4041, N4038);
and AND2 (N4042, N4040, N3573);
xor XOR2 (N4043, N4041, N310);
nand NAND2 (N4044, N3986, N1071);
not NOT1 (N4045, N4034);
nand NAND3 (N4046, N3996, N121, N612);
nor NOR3 (N4047, N4045, N1671, N2436);
buf BUF1 (N4048, N4044);
nand NAND2 (N4049, N4048, N1887);
nand NAND4 (N4050, N4021, N2863, N3943, N3611);
not NOT1 (N4051, N4047);
or OR2 (N4052, N4030, N3309);
buf BUF1 (N4053, N4046);
buf BUF1 (N4054, N4042);
nand NAND3 (N4055, N4054, N3735, N1572);
and AND3 (N4056, N4050, N3140, N324);
and AND2 (N4057, N4055, N2598);
nor NOR2 (N4058, N4039, N1155);
xor XOR2 (N4059, N4053, N1854);
buf BUF1 (N4060, N4049);
nor NOR2 (N4061, N4026, N125);
nor NOR3 (N4062, N4052, N3727, N767);
buf BUF1 (N4063, N4057);
and AND3 (N4064, N4043, N2552, N438);
and AND4 (N4065, N4059, N947, N631, N2460);
or OR3 (N4066, N4058, N774, N3722);
xor XOR2 (N4067, N4056, N1098);
and AND2 (N4068, N4060, N2388);
buf BUF1 (N4069, N4061);
buf BUF1 (N4070, N4069);
not NOT1 (N4071, N4051);
not NOT1 (N4072, N4066);
not NOT1 (N4073, N4065);
or OR3 (N4074, N4063, N1163, N2224);
not NOT1 (N4075, N4068);
and AND4 (N4076, N4075, N2716, N1133, N867);
xor XOR2 (N4077, N4070, N1053);
nor NOR3 (N4078, N4072, N1541, N2659);
nor NOR4 (N4079, N4071, N1518, N948, N1654);
and AND4 (N4080, N4073, N1637, N2354, N3785);
nand NAND3 (N4081, N4077, N3828, N1731);
not NOT1 (N4082, N4064);
nand NAND2 (N4083, N4078, N2731);
nor NOR3 (N4084, N4079, N3712, N3445);
or OR2 (N4085, N4082, N2419);
xor XOR2 (N4086, N4081, N1779);
xor XOR2 (N4087, N4084, N214);
nand NAND3 (N4088, N4074, N51, N355);
xor XOR2 (N4089, N4067, N3232);
not NOT1 (N4090, N4062);
buf BUF1 (N4091, N4090);
not NOT1 (N4092, N4083);
nor NOR4 (N4093, N4091, N2127, N3243, N3939);
nand NAND3 (N4094, N4093, N1230, N3732);
buf BUF1 (N4095, N4089);
and AND3 (N4096, N4094, N3809, N2863);
nand NAND4 (N4097, N4095, N1597, N1490, N1042);
not NOT1 (N4098, N4097);
not NOT1 (N4099, N4085);
buf BUF1 (N4100, N4092);
xor XOR2 (N4101, N4087, N3289);
nand NAND4 (N4102, N4096, N1340, N483, N377);
and AND3 (N4103, N4086, N2565, N3708);
nor NOR4 (N4104, N4088, N1772, N2658, N60);
xor XOR2 (N4105, N4099, N2617);
or OR2 (N4106, N4037, N2769);
nor NOR3 (N4107, N4106, N484, N1771);
buf BUF1 (N4108, N4103);
xor XOR2 (N4109, N4107, N1725);
not NOT1 (N4110, N4102);
nor NOR3 (N4111, N4104, N3290, N143);
buf BUF1 (N4112, N4100);
not NOT1 (N4113, N4076);
nand NAND4 (N4114, N4109, N2551, N2184, N2801);
xor XOR2 (N4115, N4113, N344);
nand NAND2 (N4116, N4112, N3397);
or OR3 (N4117, N4105, N363, N3235);
nor NOR4 (N4118, N4108, N2423, N3945, N3717);
nor NOR4 (N4119, N4098, N3048, N2156, N718);
xor XOR2 (N4120, N4114, N3654);
nand NAND4 (N4121, N4118, N3184, N1631, N943);
xor XOR2 (N4122, N4115, N352);
not NOT1 (N4123, N4119);
nor NOR2 (N4124, N4116, N2401);
nor NOR4 (N4125, N4111, N3401, N3830, N3909);
nor NOR3 (N4126, N4117, N1393, N1595);
nand NAND3 (N4127, N4123, N811, N2706);
nor NOR2 (N4128, N4110, N2282);
nor NOR2 (N4129, N4124, N3187);
not NOT1 (N4130, N4121);
and AND2 (N4131, N4126, N2074);
xor XOR2 (N4132, N4122, N3040);
and AND3 (N4133, N4132, N166, N2199);
nor NOR2 (N4134, N4080, N3376);
nor NOR4 (N4135, N4134, N2075, N2532, N3853);
buf BUF1 (N4136, N4125);
and AND3 (N4137, N4127, N2588, N2122);
not NOT1 (N4138, N4120);
nor NOR2 (N4139, N4101, N2904);
not NOT1 (N4140, N4136);
not NOT1 (N4141, N4131);
and AND2 (N4142, N4128, N2560);
nor NOR2 (N4143, N4141, N3170);
and AND4 (N4144, N4143, N314, N1029, N3685);
nor NOR2 (N4145, N4135, N1165);
nand NAND4 (N4146, N4133, N3910, N3689, N670);
not NOT1 (N4147, N4146);
not NOT1 (N4148, N4130);
buf BUF1 (N4149, N4145);
buf BUF1 (N4150, N4140);
xor XOR2 (N4151, N4150, N287);
nor NOR2 (N4152, N4138, N4010);
not NOT1 (N4153, N4148);
not NOT1 (N4154, N4153);
or OR3 (N4155, N4137, N265, N1566);
and AND4 (N4156, N4142, N1890, N2182, N3967);
nor NOR2 (N4157, N4154, N2011);
or OR4 (N4158, N4139, N3403, N2498, N2106);
and AND4 (N4159, N4129, N1154, N3461, N4011);
not NOT1 (N4160, N4144);
and AND4 (N4161, N4149, N542, N2190, N108);
and AND4 (N4162, N4157, N2140, N2423, N24);
xor XOR2 (N4163, N4151, N815);
nand NAND4 (N4164, N4155, N1930, N3143, N2617);
nand NAND4 (N4165, N4161, N1289, N3871, N1467);
or OR4 (N4166, N4162, N3315, N2888, N1266);
not NOT1 (N4167, N4152);
buf BUF1 (N4168, N4160);
xor XOR2 (N4169, N4168, N4113);
nor NOR2 (N4170, N4147, N3285);
buf BUF1 (N4171, N4164);
and AND4 (N4172, N4159, N148, N3094, N1791);
nor NOR3 (N4173, N4172, N387, N2850);
not NOT1 (N4174, N4166);
nand NAND4 (N4175, N4170, N520, N1785, N76);
and AND4 (N4176, N4163, N2303, N195, N1996);
or OR2 (N4177, N4171, N2675);
nor NOR3 (N4178, N4174, N677, N2081);
xor XOR2 (N4179, N4178, N2582);
nor NOR4 (N4180, N4177, N76, N1197, N100);
xor XOR2 (N4181, N4158, N3551);
not NOT1 (N4182, N4180);
xor XOR2 (N4183, N4169, N3683);
xor XOR2 (N4184, N4182, N2295);
nor NOR4 (N4185, N4167, N1499, N3749, N2556);
xor XOR2 (N4186, N4176, N1191);
buf BUF1 (N4187, N4184);
or OR4 (N4188, N4181, N1637, N2947, N3667);
buf BUF1 (N4189, N4186);
and AND2 (N4190, N4188, N3745);
and AND3 (N4191, N4187, N1178, N3527);
nand NAND2 (N4192, N4183, N3044);
or OR3 (N4193, N4190, N1805, N1863);
nor NOR2 (N4194, N4189, N4146);
not NOT1 (N4195, N4179);
nor NOR4 (N4196, N4173, N512, N2506, N1770);
or OR3 (N4197, N4196, N1225, N2387);
not NOT1 (N4198, N4175);
nor NOR2 (N4199, N4193, N3731);
nor NOR2 (N4200, N4191, N52);
or OR4 (N4201, N4199, N1770, N2717, N1215);
and AND2 (N4202, N4200, N3957);
and AND2 (N4203, N4201, N574);
not NOT1 (N4204, N4198);
not NOT1 (N4205, N4195);
not NOT1 (N4206, N4185);
xor XOR2 (N4207, N4205, N3080);
nand NAND3 (N4208, N4197, N2597, N2340);
or OR4 (N4209, N4207, N437, N3774, N3294);
nand NAND4 (N4210, N4206, N648, N1129, N785);
not NOT1 (N4211, N4156);
nand NAND3 (N4212, N4208, N2827, N4098);
not NOT1 (N4213, N4194);
nand NAND2 (N4214, N4192, N977);
buf BUF1 (N4215, N4209);
nand NAND3 (N4216, N4210, N3115, N2548);
xor XOR2 (N4217, N4165, N475);
xor XOR2 (N4218, N4216, N1524);
nand NAND3 (N4219, N4214, N1785, N703);
not NOT1 (N4220, N4217);
buf BUF1 (N4221, N4215);
buf BUF1 (N4222, N4204);
not NOT1 (N4223, N4218);
or OR3 (N4224, N4222, N3976, N496);
nor NOR4 (N4225, N4213, N667, N1208, N2376);
buf BUF1 (N4226, N4220);
nand NAND2 (N4227, N4202, N3047);
nand NAND2 (N4228, N4224, N627);
buf BUF1 (N4229, N4212);
xor XOR2 (N4230, N4228, N3485);
and AND2 (N4231, N4203, N3532);
not NOT1 (N4232, N4211);
buf BUF1 (N4233, N4223);
not NOT1 (N4234, N4229);
and AND2 (N4235, N4234, N2991);
or OR2 (N4236, N4231, N3456);
not NOT1 (N4237, N4232);
xor XOR2 (N4238, N4225, N443);
buf BUF1 (N4239, N4233);
nand NAND3 (N4240, N4238, N1976, N2586);
not NOT1 (N4241, N4240);
not NOT1 (N4242, N4227);
xor XOR2 (N4243, N4239, N4002);
and AND4 (N4244, N4237, N1892, N1443, N2123);
or OR3 (N4245, N4230, N3273, N2965);
nand NAND4 (N4246, N4221, N2178, N253, N1539);
and AND2 (N4247, N4243, N2900);
nor NOR2 (N4248, N4235, N1477);
buf BUF1 (N4249, N4219);
and AND4 (N4250, N4236, N2075, N253, N568);
nor NOR3 (N4251, N4242, N3799, N3078);
or OR4 (N4252, N4226, N2601, N3422, N2783);
nor NOR3 (N4253, N4247, N519, N120);
and AND4 (N4254, N4252, N3088, N1899, N1772);
not NOT1 (N4255, N4244);
nor NOR3 (N4256, N4250, N3425, N922);
not NOT1 (N4257, N4251);
xor XOR2 (N4258, N4241, N3484);
nor NOR4 (N4259, N4258, N2070, N340, N258);
xor XOR2 (N4260, N4245, N3551);
not NOT1 (N4261, N4249);
and AND4 (N4262, N4257, N3782, N2351, N4210);
not NOT1 (N4263, N4256);
nand NAND3 (N4264, N4262, N2507, N1213);
not NOT1 (N4265, N4261);
or OR4 (N4266, N4259, N1589, N133, N3501);
or OR3 (N4267, N4260, N3290, N4082);
buf BUF1 (N4268, N4246);
and AND4 (N4269, N4253, N669, N1819, N3535);
xor XOR2 (N4270, N4264, N1816);
nand NAND4 (N4271, N4248, N2191, N3872, N52);
xor XOR2 (N4272, N4267, N2531);
nand NAND2 (N4273, N4269, N377);
or OR4 (N4274, N4272, N4244, N270, N3869);
buf BUF1 (N4275, N4254);
xor XOR2 (N4276, N4274, N683);
buf BUF1 (N4277, N4271);
and AND3 (N4278, N4265, N485, N2013);
not NOT1 (N4279, N4278);
not NOT1 (N4280, N4277);
or OR2 (N4281, N4255, N2165);
not NOT1 (N4282, N4279);
nor NOR3 (N4283, N4276, N3853, N3196);
nor NOR2 (N4284, N4268, N3120);
not NOT1 (N4285, N4282);
xor XOR2 (N4286, N4285, N3795);
and AND2 (N4287, N4284, N1925);
nor NOR3 (N4288, N4280, N2468, N982);
nand NAND4 (N4289, N4263, N1734, N2948, N2271);
not NOT1 (N4290, N4283);
or OR4 (N4291, N4281, N278, N1885, N3008);
xor XOR2 (N4292, N4291, N2398);
nor NOR4 (N4293, N4290, N67, N2007, N3448);
nor NOR4 (N4294, N4288, N554, N3799, N2353);
nand NAND2 (N4295, N4294, N2308);
and AND4 (N4296, N4273, N4065, N1070, N3018);
and AND4 (N4297, N4295, N526, N2975, N3957);
or OR4 (N4298, N4287, N3412, N2818, N3392);
and AND2 (N4299, N4293, N808);
nor NOR4 (N4300, N4299, N3955, N1304, N313);
buf BUF1 (N4301, N4270);
xor XOR2 (N4302, N4301, N943);
or OR2 (N4303, N4289, N2369);
not NOT1 (N4304, N4302);
xor XOR2 (N4305, N4292, N1708);
xor XOR2 (N4306, N4305, N3337);
buf BUF1 (N4307, N4304);
or OR4 (N4308, N4307, N3872, N2912, N141);
nor NOR2 (N4309, N4303, N2659);
xor XOR2 (N4310, N4308, N3218);
buf BUF1 (N4311, N4286);
buf BUF1 (N4312, N4266);
or OR2 (N4313, N4300, N1145);
nor NOR4 (N4314, N4297, N633, N2593, N2304);
or OR3 (N4315, N4310, N1329, N3828);
and AND3 (N4316, N4296, N876, N2817);
and AND4 (N4317, N4298, N3118, N1286, N521);
buf BUF1 (N4318, N4311);
xor XOR2 (N4319, N4275, N4251);
xor XOR2 (N4320, N4318, N2874);
xor XOR2 (N4321, N4313, N163);
and AND4 (N4322, N4312, N1593, N2310, N233);
or OR3 (N4323, N4314, N1320, N1033);
xor XOR2 (N4324, N4316, N1804);
nor NOR4 (N4325, N4322, N2308, N164, N1582);
or OR2 (N4326, N4325, N711);
and AND2 (N4327, N4306, N3584);
buf BUF1 (N4328, N4320);
buf BUF1 (N4329, N4319);
or OR2 (N4330, N4327, N155);
and AND4 (N4331, N4329, N2632, N3673, N1950);
nand NAND2 (N4332, N4321, N2119);
xor XOR2 (N4333, N4317, N546);
buf BUF1 (N4334, N4330);
not NOT1 (N4335, N4331);
or OR2 (N4336, N4335, N4032);
xor XOR2 (N4337, N4324, N4134);
or OR2 (N4338, N4332, N2434);
or OR2 (N4339, N4326, N3687);
not NOT1 (N4340, N4336);
xor XOR2 (N4341, N4338, N820);
nand NAND4 (N4342, N4323, N607, N672, N3871);
not NOT1 (N4343, N4333);
nand NAND4 (N4344, N4339, N2557, N1454, N1666);
buf BUF1 (N4345, N4337);
not NOT1 (N4346, N4345);
buf BUF1 (N4347, N4341);
nor NOR3 (N4348, N4340, N2778, N3007);
not NOT1 (N4349, N4315);
buf BUF1 (N4350, N4347);
xor XOR2 (N4351, N4350, N2073);
or OR4 (N4352, N4351, N1823, N1238, N2533);
not NOT1 (N4353, N4352);
nor NOR4 (N4354, N4334, N591, N1791, N1054);
xor XOR2 (N4355, N4309, N3437);
nor NOR4 (N4356, N4344, N3808, N307, N1037);
and AND3 (N4357, N4354, N764, N2603);
not NOT1 (N4358, N4343);
and AND2 (N4359, N4357, N3499);
xor XOR2 (N4360, N4346, N1160);
buf BUF1 (N4361, N4360);
nand NAND3 (N4362, N4361, N4115, N2652);
nor NOR4 (N4363, N4348, N987, N2483, N1146);
xor XOR2 (N4364, N4353, N3650);
buf BUF1 (N4365, N4364);
and AND4 (N4366, N4363, N3354, N2851, N3700);
or OR3 (N4367, N4359, N2961, N2686);
xor XOR2 (N4368, N4342, N2849);
xor XOR2 (N4369, N4365, N4024);
buf BUF1 (N4370, N4366);
nor NOR4 (N4371, N4369, N1457, N417, N2902);
nor NOR3 (N4372, N4368, N1556, N3477);
or OR3 (N4373, N4362, N2903, N36);
or OR2 (N4374, N4372, N3180);
or OR2 (N4375, N4355, N3566);
nand NAND4 (N4376, N4371, N3768, N2012, N1653);
not NOT1 (N4377, N4374);
nand NAND4 (N4378, N4375, N2327, N3195, N1493);
xor XOR2 (N4379, N4378, N1936);
nand NAND4 (N4380, N4376, N1754, N926, N3298);
or OR4 (N4381, N4328, N2240, N950, N1763);
nand NAND2 (N4382, N4373, N989);
nor NOR3 (N4383, N4379, N713, N3147);
or OR2 (N4384, N4356, N3088);
xor XOR2 (N4385, N4381, N379);
xor XOR2 (N4386, N4370, N1961);
xor XOR2 (N4387, N4386, N1761);
nand NAND2 (N4388, N4358, N1401);
or OR3 (N4389, N4388, N1508, N1021);
or OR4 (N4390, N4385, N3149, N360, N2217);
not NOT1 (N4391, N4367);
nand NAND3 (N4392, N4390, N3316, N781);
not NOT1 (N4393, N4349);
not NOT1 (N4394, N4377);
or OR2 (N4395, N4383, N3503);
or OR3 (N4396, N4391, N3016, N1352);
or OR3 (N4397, N4380, N3135, N4093);
xor XOR2 (N4398, N4384, N1322);
nand NAND2 (N4399, N4387, N2542);
xor XOR2 (N4400, N4395, N868);
and AND2 (N4401, N4396, N2270);
or OR2 (N4402, N4392, N3316);
buf BUF1 (N4403, N4398);
xor XOR2 (N4404, N4397, N3141);
nand NAND2 (N4405, N4393, N3189);
or OR4 (N4406, N4404, N879, N575, N3439);
nor NOR2 (N4407, N4402, N1852);
and AND4 (N4408, N4401, N688, N3319, N3932);
nor NOR2 (N4409, N4406, N393);
nand NAND4 (N4410, N4389, N1382, N2635, N2139);
or OR2 (N4411, N4394, N1298);
buf BUF1 (N4412, N4403);
nand NAND3 (N4413, N4410, N252, N1434);
and AND2 (N4414, N4382, N3589);
or OR2 (N4415, N4399, N475);
nor NOR4 (N4416, N4414, N1225, N919, N3358);
buf BUF1 (N4417, N4405);
xor XOR2 (N4418, N4400, N1754);
nor NOR3 (N4419, N4415, N840, N3338);
not NOT1 (N4420, N4407);
nor NOR2 (N4421, N4416, N1724);
xor XOR2 (N4422, N4417, N2942);
or OR3 (N4423, N4420, N1626, N4239);
and AND4 (N4424, N4409, N4351, N492, N1618);
xor XOR2 (N4425, N4419, N3601);
nor NOR3 (N4426, N4411, N715, N219);
not NOT1 (N4427, N4418);
or OR4 (N4428, N4423, N47, N4123, N869);
nor NOR4 (N4429, N4427, N4043, N2293, N2483);
xor XOR2 (N4430, N4426, N3269);
nor NOR2 (N4431, N4429, N1793);
buf BUF1 (N4432, N4430);
nand NAND3 (N4433, N4421, N550, N3804);
nor NOR3 (N4434, N4428, N1095, N4309);
or OR4 (N4435, N4431, N2806, N1263, N2222);
xor XOR2 (N4436, N4432, N133);
xor XOR2 (N4437, N4435, N2816);
or OR4 (N4438, N4434, N3014, N996, N1381);
nand NAND2 (N4439, N4433, N3463);
xor XOR2 (N4440, N4438, N3427);
nand NAND4 (N4441, N4436, N663, N1216, N1605);
not NOT1 (N4442, N4425);
buf BUF1 (N4443, N4422);
xor XOR2 (N4444, N4408, N3858);
nor NOR3 (N4445, N4412, N2857, N4011);
not NOT1 (N4446, N4441);
or OR3 (N4447, N4442, N4361, N480);
nor NOR4 (N4448, N4447, N567, N2519, N886);
buf BUF1 (N4449, N4448);
xor XOR2 (N4450, N4445, N4424);
and AND3 (N4451, N1548, N2246, N1959);
and AND2 (N4452, N4437, N3955);
or OR4 (N4453, N4439, N146, N2847, N724);
xor XOR2 (N4454, N4446, N4296);
buf BUF1 (N4455, N4454);
nor NOR3 (N4456, N4453, N175, N2495);
buf BUF1 (N4457, N4413);
or OR2 (N4458, N4457, N541);
not NOT1 (N4459, N4444);
nand NAND4 (N4460, N4451, N837, N1475, N150);
or OR2 (N4461, N4452, N1307);
buf BUF1 (N4462, N4443);
or OR2 (N4463, N4450, N1440);
and AND4 (N4464, N4458, N2393, N3764, N2720);
or OR2 (N4465, N4440, N1732);
xor XOR2 (N4466, N4455, N166);
nand NAND4 (N4467, N4460, N3874, N1966, N1163);
and AND3 (N4468, N4465, N175, N3828);
or OR2 (N4469, N4461, N435);
or OR3 (N4470, N4467, N1302, N856);
xor XOR2 (N4471, N4449, N3897);
or OR2 (N4472, N4463, N3740);
and AND4 (N4473, N4456, N1443, N4263, N346);
xor XOR2 (N4474, N4459, N1327);
or OR2 (N4475, N4462, N4319);
and AND2 (N4476, N4473, N730);
nor NOR4 (N4477, N4472, N3113, N941, N1821);
and AND4 (N4478, N4470, N4469, N2880, N3541);
nor NOR2 (N4479, N906, N2669);
xor XOR2 (N4480, N4468, N4372);
nor NOR3 (N4481, N4464, N3145, N1470);
and AND3 (N4482, N4474, N1132, N1763);
and AND4 (N4483, N4466, N1037, N3272, N3649);
not NOT1 (N4484, N4477);
and AND2 (N4485, N4471, N1424);
or OR3 (N4486, N4479, N2071, N254);
xor XOR2 (N4487, N4481, N2661);
buf BUF1 (N4488, N4485);
or OR3 (N4489, N4487, N451, N1070);
buf BUF1 (N4490, N4484);
nor NOR2 (N4491, N4476, N2668);
buf BUF1 (N4492, N4483);
buf BUF1 (N4493, N4488);
not NOT1 (N4494, N4475);
buf BUF1 (N4495, N4482);
and AND4 (N4496, N4490, N4289, N3210, N173);
buf BUF1 (N4497, N4494);
and AND4 (N4498, N4495, N2768, N722, N2367);
buf BUF1 (N4499, N4498);
or OR4 (N4500, N4496, N2282, N3496, N67);
nand NAND3 (N4501, N4499, N2977, N4293);
not NOT1 (N4502, N4500);
buf BUF1 (N4503, N4491);
or OR4 (N4504, N4486, N2222, N1747, N72);
nor NOR4 (N4505, N4480, N358, N630, N2329);
xor XOR2 (N4506, N4478, N3831);
not NOT1 (N4507, N4493);
nand NAND2 (N4508, N4503, N3444);
or OR2 (N4509, N4492, N3054);
xor XOR2 (N4510, N4497, N4017);
or OR3 (N4511, N4501, N2769, N4170);
nand NAND3 (N4512, N4510, N4361, N2099);
nor NOR3 (N4513, N4505, N2372, N1345);
not NOT1 (N4514, N4513);
buf BUF1 (N4515, N4489);
not NOT1 (N4516, N4507);
and AND2 (N4517, N4516, N3970);
nor NOR4 (N4518, N4511, N2456, N2687, N3250);
buf BUF1 (N4519, N4512);
buf BUF1 (N4520, N4506);
not NOT1 (N4521, N4520);
and AND3 (N4522, N4517, N1704, N3768);
nand NAND2 (N4523, N4504, N4113);
or OR3 (N4524, N4522, N1794, N2702);
or OR2 (N4525, N4502, N3333);
nand NAND4 (N4526, N4523, N2548, N3326, N2282);
and AND3 (N4527, N4514, N2495, N4239);
or OR3 (N4528, N4521, N1374, N2869);
not NOT1 (N4529, N4518);
nor NOR3 (N4530, N4524, N281, N2920);
xor XOR2 (N4531, N4509, N1167);
buf BUF1 (N4532, N4519);
or OR4 (N4533, N4527, N2682, N1210, N2031);
buf BUF1 (N4534, N4526);
buf BUF1 (N4535, N4533);
buf BUF1 (N4536, N4535);
or OR3 (N4537, N4530, N1148, N3336);
not NOT1 (N4538, N4532);
xor XOR2 (N4539, N4508, N1493);
and AND4 (N4540, N4538, N3059, N4445, N3978);
or OR2 (N4541, N4534, N3395);
and AND3 (N4542, N4537, N3802, N4377);
and AND3 (N4543, N4539, N3965, N1009);
and AND2 (N4544, N4540, N2338);
or OR3 (N4545, N4525, N781, N3749);
nand NAND3 (N4546, N4542, N227, N4123);
and AND3 (N4547, N4536, N667, N4223);
buf BUF1 (N4548, N4544);
nor NOR4 (N4549, N4546, N2772, N1690, N2624);
xor XOR2 (N4550, N4531, N4272);
buf BUF1 (N4551, N4543);
or OR2 (N4552, N4528, N2656);
buf BUF1 (N4553, N4515);
and AND3 (N4554, N4553, N2231, N336);
or OR2 (N4555, N4551, N1984);
not NOT1 (N4556, N4549);
xor XOR2 (N4557, N4548, N1140);
nand NAND3 (N4558, N4541, N4119, N709);
not NOT1 (N4559, N4554);
nor NOR2 (N4560, N4557, N826);
buf BUF1 (N4561, N4529);
and AND3 (N4562, N4559, N3576, N3244);
or OR4 (N4563, N4561, N253, N1144, N2829);
nor NOR3 (N4564, N4556, N1685, N3646);
or OR4 (N4565, N4547, N2475, N782, N1931);
xor XOR2 (N4566, N4558, N1751);
nand NAND4 (N4567, N4560, N2210, N421, N2047);
nor NOR2 (N4568, N4567, N2114);
nor NOR4 (N4569, N4552, N3975, N3785, N3585);
not NOT1 (N4570, N4564);
xor XOR2 (N4571, N4566, N1693);
or OR3 (N4572, N4563, N2085, N919);
xor XOR2 (N4573, N4562, N955);
xor XOR2 (N4574, N4571, N1773);
nor NOR4 (N4575, N4555, N2710, N2818, N623);
buf BUF1 (N4576, N4573);
xor XOR2 (N4577, N4565, N3345);
and AND4 (N4578, N4575, N1900, N4290, N2817);
buf BUF1 (N4579, N4568);
not NOT1 (N4580, N4579);
xor XOR2 (N4581, N4580, N90);
not NOT1 (N4582, N4550);
nand NAND4 (N4583, N4569, N3933, N4514, N1016);
nor NOR4 (N4584, N4581, N4283, N3669, N2008);
and AND4 (N4585, N4578, N332, N1688, N1091);
not NOT1 (N4586, N4572);
xor XOR2 (N4587, N4585, N460);
or OR4 (N4588, N4574, N749, N3501, N77);
buf BUF1 (N4589, N4583);
or OR3 (N4590, N4545, N519, N1818);
not NOT1 (N4591, N4577);
and AND2 (N4592, N4589, N2463);
and AND3 (N4593, N4590, N573, N2416);
not NOT1 (N4594, N4576);
not NOT1 (N4595, N4591);
buf BUF1 (N4596, N4584);
nor NOR3 (N4597, N4588, N1828, N3392);
buf BUF1 (N4598, N4570);
or OR2 (N4599, N4582, N1739);
not NOT1 (N4600, N4599);
and AND4 (N4601, N4594, N1076, N2581, N2000);
not NOT1 (N4602, N4596);
nand NAND4 (N4603, N4593, N1456, N1120, N155);
nor NOR2 (N4604, N4595, N284);
buf BUF1 (N4605, N4587);
nor NOR3 (N4606, N4601, N4081, N1877);
buf BUF1 (N4607, N4598);
buf BUF1 (N4608, N4603);
buf BUF1 (N4609, N4586);
xor XOR2 (N4610, N4592, N1116);
buf BUF1 (N4611, N4605);
not NOT1 (N4612, N4597);
buf BUF1 (N4613, N4610);
or OR3 (N4614, N4613, N4351, N187);
or OR2 (N4615, N4609, N1366);
nor NOR2 (N4616, N4608, N1484);
nand NAND3 (N4617, N4604, N164, N1942);
and AND2 (N4618, N4606, N3388);
not NOT1 (N4619, N4611);
nand NAND3 (N4620, N4617, N149, N4054);
xor XOR2 (N4621, N4620, N4415);
xor XOR2 (N4622, N4602, N2064);
and AND2 (N4623, N4600, N131);
not NOT1 (N4624, N4619);
and AND2 (N4625, N4624, N2594);
and AND2 (N4626, N4614, N1415);
not NOT1 (N4627, N4607);
not NOT1 (N4628, N4627);
and AND2 (N4629, N4621, N1963);
nand NAND4 (N4630, N4618, N2937, N4469, N2308);
or OR3 (N4631, N4616, N3418, N2549);
or OR3 (N4632, N4630, N594, N30);
buf BUF1 (N4633, N4631);
xor XOR2 (N4634, N4628, N953);
buf BUF1 (N4635, N4625);
or OR3 (N4636, N4635, N4024, N182);
or OR4 (N4637, N4622, N1700, N675, N4231);
and AND2 (N4638, N4637, N4112);
nand NAND2 (N4639, N4638, N3421);
nor NOR3 (N4640, N4615, N2951, N1932);
nand NAND2 (N4641, N4629, N4314);
not NOT1 (N4642, N4639);
nand NAND4 (N4643, N4612, N2053, N3159, N4545);
buf BUF1 (N4644, N4623);
nand NAND4 (N4645, N4643, N3756, N3990, N1473);
and AND3 (N4646, N4645, N982, N3116);
xor XOR2 (N4647, N4632, N3995);
xor XOR2 (N4648, N4633, N2155);
nor NOR4 (N4649, N4648, N2547, N3277, N903);
nor NOR4 (N4650, N4626, N3591, N3866, N4480);
nand NAND3 (N4651, N4634, N1065, N3963);
buf BUF1 (N4652, N4647);
nor NOR4 (N4653, N4646, N1495, N266, N3305);
buf BUF1 (N4654, N4651);
xor XOR2 (N4655, N4642, N1212);
xor XOR2 (N4656, N4640, N21);
xor XOR2 (N4657, N4644, N742);
nor NOR2 (N4658, N4653, N977);
and AND3 (N4659, N4658, N1192, N1761);
xor XOR2 (N4660, N4650, N1827);
buf BUF1 (N4661, N4652);
not NOT1 (N4662, N4654);
or OR3 (N4663, N4659, N1811, N3398);
nor NOR3 (N4664, N4649, N1419, N3992);
not NOT1 (N4665, N4660);
or OR2 (N4666, N4655, N534);
nand NAND2 (N4667, N4641, N3238);
nand NAND4 (N4668, N4661, N575, N260, N2588);
buf BUF1 (N4669, N4663);
nand NAND2 (N4670, N4667, N3768);
or OR4 (N4671, N4662, N1445, N518, N2187);
xor XOR2 (N4672, N4669, N810);
or OR4 (N4673, N4656, N2890, N4329, N2474);
or OR4 (N4674, N4673, N671, N4203, N1625);
not NOT1 (N4675, N4664);
and AND3 (N4676, N4636, N3028, N1923);
xor XOR2 (N4677, N4676, N1539);
or OR2 (N4678, N4675, N1899);
not NOT1 (N4679, N4678);
nand NAND3 (N4680, N4672, N203, N458);
not NOT1 (N4681, N4666);
nand NAND4 (N4682, N4677, N1842, N4322, N1116);
nand NAND3 (N4683, N4674, N3126, N3261);
or OR4 (N4684, N4682, N634, N2097, N1192);
and AND3 (N4685, N4670, N2867, N763);
and AND3 (N4686, N4668, N2882, N1268);
or OR3 (N4687, N4679, N2722, N4523);
nor NOR2 (N4688, N4685, N1673);
nand NAND2 (N4689, N4687, N2302);
nor NOR2 (N4690, N4686, N2157);
nand NAND4 (N4691, N4690, N3539, N371, N1681);
nand NAND2 (N4692, N4657, N4115);
nand NAND2 (N4693, N4692, N172);
not NOT1 (N4694, N4680);
and AND3 (N4695, N4665, N110, N1076);
not NOT1 (N4696, N4684);
not NOT1 (N4697, N4683);
buf BUF1 (N4698, N4696);
buf BUF1 (N4699, N4695);
and AND4 (N4700, N4689, N3490, N696, N613);
buf BUF1 (N4701, N4698);
xor XOR2 (N4702, N4671, N590);
not NOT1 (N4703, N4697);
and AND3 (N4704, N4688, N1172, N3380);
and AND2 (N4705, N4699, N2105);
nor NOR2 (N4706, N4705, N1316);
nand NAND4 (N4707, N4694, N4085, N3023, N132);
or OR2 (N4708, N4707, N3363);
and AND3 (N4709, N4700, N170, N4320);
buf BUF1 (N4710, N4693);
nor NOR2 (N4711, N4708, N3754);
xor XOR2 (N4712, N4701, N1983);
and AND4 (N4713, N4691, N1566, N629, N4353);
or OR3 (N4714, N4704, N1027, N132);
nor NOR2 (N4715, N4681, N1836);
nand NAND2 (N4716, N4703, N3314);
nand NAND3 (N4717, N4712, N3627, N2649);
and AND2 (N4718, N4717, N2088);
and AND3 (N4719, N4706, N2935, N3865);
buf BUF1 (N4720, N4718);
nand NAND4 (N4721, N4720, N3431, N1451, N2335);
nor NOR2 (N4722, N4702, N2932);
nor NOR2 (N4723, N4721, N1420);
not NOT1 (N4724, N4719);
buf BUF1 (N4725, N4709);
buf BUF1 (N4726, N4713);
not NOT1 (N4727, N4714);
not NOT1 (N4728, N4715);
or OR4 (N4729, N4726, N3065, N4540, N2160);
nor NOR4 (N4730, N4716, N1259, N1028, N3946);
nand NAND2 (N4731, N4730, N996);
and AND4 (N4732, N4727, N1112, N3533, N3277);
xor XOR2 (N4733, N4728, N3482);
xor XOR2 (N4734, N4722, N149);
or OR3 (N4735, N4731, N1012, N4216);
and AND4 (N4736, N4734, N2797, N2825, N4635);
buf BUF1 (N4737, N4736);
buf BUF1 (N4738, N4737);
buf BUF1 (N4739, N4732);
nand NAND3 (N4740, N4725, N3600, N3353);
and AND4 (N4741, N4729, N2317, N4028, N3432);
buf BUF1 (N4742, N4740);
nand NAND4 (N4743, N4710, N533, N3058, N1574);
nor NOR3 (N4744, N4739, N717, N2687);
buf BUF1 (N4745, N4744);
not NOT1 (N4746, N4735);
not NOT1 (N4747, N4741);
not NOT1 (N4748, N4724);
or OR4 (N4749, N4745, N281, N4246, N3362);
or OR3 (N4750, N4746, N3540, N2795);
or OR3 (N4751, N4747, N1009, N3837);
nor NOR3 (N4752, N4743, N3126, N3121);
nand NAND3 (N4753, N4748, N1107, N1232);
buf BUF1 (N4754, N4751);
nand NAND3 (N4755, N4738, N3489, N3920);
buf BUF1 (N4756, N4733);
or OR4 (N4757, N4755, N3208, N435, N4737);
nand NAND2 (N4758, N4757, N135);
or OR3 (N4759, N4750, N788, N54);
not NOT1 (N4760, N4711);
nand NAND3 (N4761, N4756, N3832, N3214);
or OR3 (N4762, N4742, N232, N654);
xor XOR2 (N4763, N4753, N3865);
and AND3 (N4764, N4762, N4154, N4539);
nand NAND3 (N4765, N4759, N255, N1755);
and AND3 (N4766, N4760, N4762, N148);
nor NOR3 (N4767, N4758, N2552, N341);
nand NAND3 (N4768, N4723, N1363, N2054);
buf BUF1 (N4769, N4765);
not NOT1 (N4770, N4768);
or OR4 (N4771, N4763, N135, N3511, N3413);
not NOT1 (N4772, N4766);
buf BUF1 (N4773, N4749);
and AND2 (N4774, N4772, N3431);
xor XOR2 (N4775, N4767, N2347);
nor NOR4 (N4776, N4764, N4275, N1524, N584);
or OR4 (N4777, N4775, N102, N3385, N4607);
and AND2 (N4778, N4777, N3228);
nor NOR3 (N4779, N4774, N4744, N1179);
or OR2 (N4780, N4761, N1100);
nand NAND4 (N4781, N4778, N1842, N2376, N909);
buf BUF1 (N4782, N4771);
xor XOR2 (N4783, N4780, N1216);
nand NAND3 (N4784, N4773, N713, N4251);
buf BUF1 (N4785, N4769);
not NOT1 (N4786, N4784);
xor XOR2 (N4787, N4781, N346);
not NOT1 (N4788, N4783);
xor XOR2 (N4789, N4754, N2236);
or OR4 (N4790, N4779, N171, N111, N2144);
and AND2 (N4791, N4790, N751);
nor NOR2 (N4792, N4770, N4017);
and AND4 (N4793, N4788, N3813, N303, N2541);
nand NAND4 (N4794, N4752, N2023, N819, N840);
nor NOR3 (N4795, N4792, N1636, N1321);
nand NAND4 (N4796, N4776, N3371, N2699, N1465);
xor XOR2 (N4797, N4785, N4388);
nand NAND3 (N4798, N4797, N4732, N1515);
nor NOR4 (N4799, N4787, N2947, N2604, N3507);
buf BUF1 (N4800, N4798);
nand NAND4 (N4801, N4786, N644, N571, N4446);
and AND4 (N4802, N4793, N3124, N2354, N213);
or OR3 (N4803, N4794, N281, N3460);
and AND3 (N4804, N4782, N3562, N2450);
nor NOR2 (N4805, N4800, N3897);
xor XOR2 (N4806, N4801, N1423);
or OR4 (N4807, N4803, N229, N1303, N707);
nand NAND4 (N4808, N4806, N720, N4595, N194);
or OR2 (N4809, N4799, N1947);
or OR4 (N4810, N4802, N1561, N4804, N1201);
nand NAND3 (N4811, N1473, N1553, N1858);
xor XOR2 (N4812, N4809, N2768);
or OR2 (N4813, N4805, N3872);
nand NAND4 (N4814, N4812, N646, N4304, N2937);
nand NAND2 (N4815, N4813, N3266);
xor XOR2 (N4816, N4796, N1161);
or OR2 (N4817, N4810, N2515);
xor XOR2 (N4818, N4814, N2555);
not NOT1 (N4819, N4816);
xor XOR2 (N4820, N4789, N1734);
nand NAND2 (N4821, N4817, N876);
or OR4 (N4822, N4795, N1970, N4464, N3963);
not NOT1 (N4823, N4791);
xor XOR2 (N4824, N4820, N4616);
buf BUF1 (N4825, N4822);
or OR3 (N4826, N4811, N3850, N3048);
nand NAND4 (N4827, N4823, N3213, N1193, N891);
buf BUF1 (N4828, N4818);
and AND3 (N4829, N4808, N99, N4492);
xor XOR2 (N4830, N4821, N4475);
nor NOR3 (N4831, N4819, N2392, N2136);
not NOT1 (N4832, N4828);
xor XOR2 (N4833, N4825, N875);
buf BUF1 (N4834, N4831);
xor XOR2 (N4835, N4833, N1152);
buf BUF1 (N4836, N4826);
nand NAND3 (N4837, N4807, N575, N3382);
and AND3 (N4838, N4834, N1422, N4672);
buf BUF1 (N4839, N4837);
nand NAND4 (N4840, N4815, N33, N4281, N1467);
nor NOR4 (N4841, N4830, N4414, N4212, N2797);
and AND2 (N4842, N4841, N3481);
nand NAND3 (N4843, N4840, N2935, N3370);
or OR3 (N4844, N4824, N4301, N2942);
buf BUF1 (N4845, N4843);
xor XOR2 (N4846, N4827, N3829);
not NOT1 (N4847, N4835);
buf BUF1 (N4848, N4839);
nand NAND3 (N4849, N4844, N3352, N4002);
and AND4 (N4850, N4849, N661, N892, N2797);
or OR3 (N4851, N4829, N1469, N3264);
nor NOR3 (N4852, N4848, N1897, N1149);
not NOT1 (N4853, N4842);
nor NOR2 (N4854, N4832, N2446);
and AND3 (N4855, N4852, N3063, N2513);
nor NOR2 (N4856, N4845, N292);
nand NAND2 (N4857, N4850, N4051);
buf BUF1 (N4858, N4854);
buf BUF1 (N4859, N4855);
nand NAND3 (N4860, N4838, N2832, N3102);
and AND3 (N4861, N4836, N175, N3593);
and AND2 (N4862, N4857, N1678);
and AND3 (N4863, N4862, N67, N2656);
not NOT1 (N4864, N4846);
or OR2 (N4865, N4863, N2878);
buf BUF1 (N4866, N4853);
or OR3 (N4867, N4864, N3586, N254);
not NOT1 (N4868, N4867);
not NOT1 (N4869, N4856);
nand NAND4 (N4870, N4861, N2293, N1672, N2870);
and AND3 (N4871, N4858, N4335, N1463);
xor XOR2 (N4872, N4865, N571);
not NOT1 (N4873, N4847);
xor XOR2 (N4874, N4871, N929);
and AND3 (N4875, N4859, N3250, N502);
nand NAND2 (N4876, N4860, N4734);
nand NAND3 (N4877, N4874, N4677, N4679);
and AND2 (N4878, N4875, N1984);
buf BUF1 (N4879, N4873);
nor NOR2 (N4880, N4869, N2496);
nand NAND3 (N4881, N4877, N2028, N182);
or OR4 (N4882, N4876, N743, N1138, N3573);
nor NOR2 (N4883, N4868, N4664);
or OR3 (N4884, N4879, N4760, N2931);
or OR2 (N4885, N4884, N2229);
not NOT1 (N4886, N4883);
nand NAND2 (N4887, N4878, N2141);
and AND4 (N4888, N4870, N3930, N1562, N2740);
buf BUF1 (N4889, N4866);
nand NAND3 (N4890, N4886, N3094, N1706);
nand NAND4 (N4891, N4880, N2373, N3665, N3987);
and AND2 (N4892, N4882, N1738);
nand NAND3 (N4893, N4892, N2259, N1191);
nor NOR4 (N4894, N4851, N1087, N4757, N466);
not NOT1 (N4895, N4889);
nand NAND2 (N4896, N4890, N3583);
buf BUF1 (N4897, N4893);
xor XOR2 (N4898, N4891, N4602);
not NOT1 (N4899, N4895);
not NOT1 (N4900, N4885);
not NOT1 (N4901, N4897);
nand NAND2 (N4902, N4894, N4546);
or OR3 (N4903, N4887, N1382, N4367);
and AND4 (N4904, N4888, N3058, N2148, N2489);
or OR2 (N4905, N4901, N4370);
nand NAND4 (N4906, N4902, N4051, N4748, N915);
and AND2 (N4907, N4905, N88);
buf BUF1 (N4908, N4899);
nor NOR4 (N4909, N4896, N342, N740, N3461);
buf BUF1 (N4910, N4881);
buf BUF1 (N4911, N4903);
nand NAND3 (N4912, N4910, N4209, N2342);
not NOT1 (N4913, N4872);
not NOT1 (N4914, N4912);
nor NOR3 (N4915, N4913, N2229, N946);
nand NAND3 (N4916, N4909, N3226, N2153);
not NOT1 (N4917, N4907);
or OR3 (N4918, N4916, N692, N3987);
xor XOR2 (N4919, N4906, N94);
xor XOR2 (N4920, N4898, N4658);
buf BUF1 (N4921, N4920);
and AND4 (N4922, N4921, N1915, N3375, N4269);
not NOT1 (N4923, N4908);
not NOT1 (N4924, N4917);
xor XOR2 (N4925, N4904, N3056);
nand NAND2 (N4926, N4911, N3102);
xor XOR2 (N4927, N4923, N2069);
and AND2 (N4928, N4925, N2744);
and AND2 (N4929, N4928, N1213);
buf BUF1 (N4930, N4924);
xor XOR2 (N4931, N4919, N546);
nand NAND2 (N4932, N4929, N4225);
xor XOR2 (N4933, N4931, N3349);
and AND2 (N4934, N4926, N337);
not NOT1 (N4935, N4927);
or OR3 (N4936, N4914, N735, N4613);
and AND3 (N4937, N4936, N3462, N4017);
nor NOR2 (N4938, N4933, N302);
xor XOR2 (N4939, N4915, N117);
nand NAND4 (N4940, N4935, N1745, N2520, N2613);
nand NAND2 (N4941, N4918, N4171);
nand NAND2 (N4942, N4934, N137);
xor XOR2 (N4943, N4941, N770);
xor XOR2 (N4944, N4939, N4674);
xor XOR2 (N4945, N4943, N613);
or OR4 (N4946, N4942, N1521, N2931, N1296);
nand NAND2 (N4947, N4944, N2090);
buf BUF1 (N4948, N4932);
and AND2 (N4949, N4945, N1759);
nor NOR3 (N4950, N4900, N301, N3003);
or OR3 (N4951, N4946, N3142, N4676);
and AND4 (N4952, N4937, N2657, N4914, N1854);
xor XOR2 (N4953, N4947, N3000);
nand NAND4 (N4954, N4930, N3407, N3620, N781);
xor XOR2 (N4955, N4950, N591);
not NOT1 (N4956, N4951);
nor NOR4 (N4957, N4938, N4861, N1010, N1577);
nand NAND4 (N4958, N4954, N4883, N2256, N1483);
buf BUF1 (N4959, N4957);
nand NAND2 (N4960, N4952, N4203);
and AND3 (N4961, N4949, N2989, N4066);
and AND3 (N4962, N4922, N363, N3745);
nand NAND4 (N4963, N4953, N4605, N956, N2151);
or OR3 (N4964, N4958, N1185, N509);
xor XOR2 (N4965, N4940, N4596);
xor XOR2 (N4966, N4959, N1241);
nand NAND3 (N4967, N4960, N1194, N4346);
xor XOR2 (N4968, N4961, N4359);
buf BUF1 (N4969, N4968);
or OR2 (N4970, N4963, N2365);
or OR2 (N4971, N4948, N2074);
buf BUF1 (N4972, N4970);
xor XOR2 (N4973, N4969, N3753);
not NOT1 (N4974, N4967);
or OR3 (N4975, N4955, N1972, N3702);
xor XOR2 (N4976, N4956, N2076);
and AND3 (N4977, N4972, N2643, N1511);
nand NAND4 (N4978, N4975, N2342, N860, N2021);
nand NAND3 (N4979, N4973, N410, N347);
nand NAND4 (N4980, N4965, N51, N2602, N4900);
or OR3 (N4981, N4980, N1982, N4655);
xor XOR2 (N4982, N4981, N3357);
xor XOR2 (N4983, N4964, N645);
buf BUF1 (N4984, N4983);
buf BUF1 (N4985, N4984);
nand NAND2 (N4986, N4962, N3481);
nor NOR4 (N4987, N4978, N613, N3464, N4124);
buf BUF1 (N4988, N4985);
not NOT1 (N4989, N4977);
or OR4 (N4990, N4989, N4003, N3720, N2135);
buf BUF1 (N4991, N4974);
nor NOR2 (N4992, N4979, N4172);
xor XOR2 (N4993, N4976, N2636);
buf BUF1 (N4994, N4988);
or OR3 (N4995, N4993, N763, N2536);
and AND4 (N4996, N4982, N3373, N4612, N4973);
xor XOR2 (N4997, N4990, N770);
nand NAND3 (N4998, N4971, N102, N906);
and AND2 (N4999, N4986, N4174);
or OR4 (N5000, N4991, N4276, N1716, N3427);
and AND3 (N5001, N4966, N1352, N1099);
or OR2 (N5002, N4998, N4000);
buf BUF1 (N5003, N5000);
not NOT1 (N5004, N5003);
xor XOR2 (N5005, N4997, N2416);
not NOT1 (N5006, N4987);
and AND3 (N5007, N5006, N2902, N4966);
and AND3 (N5008, N4995, N1355, N4060);
or OR3 (N5009, N5001, N3946, N2625);
nand NAND4 (N5010, N5009, N956, N3258, N302);
or OR2 (N5011, N5002, N1283);
not NOT1 (N5012, N5011);
not NOT1 (N5013, N5007);
not NOT1 (N5014, N4994);
and AND4 (N5015, N5012, N3398, N4937, N3869);
buf BUF1 (N5016, N5004);
buf BUF1 (N5017, N5013);
xor XOR2 (N5018, N4992, N221);
xor XOR2 (N5019, N5014, N447);
not NOT1 (N5020, N5018);
and AND4 (N5021, N5005, N3649, N676, N1845);
not NOT1 (N5022, N4996);
or OR3 (N5023, N5020, N824, N4375);
not NOT1 (N5024, N5017);
not NOT1 (N5025, N5019);
buf BUF1 (N5026, N5015);
nand NAND4 (N5027, N5016, N3966, N92, N3488);
nor NOR3 (N5028, N5024, N2301, N1841);
nor NOR2 (N5029, N5026, N1123);
nor NOR4 (N5030, N5029, N72, N2389, N2559);
and AND3 (N5031, N5008, N4590, N1797);
buf BUF1 (N5032, N4999);
buf BUF1 (N5033, N5025);
and AND2 (N5034, N5023, N4627);
buf BUF1 (N5035, N5021);
nor NOR4 (N5036, N5028, N2306, N4585, N1910);
nor NOR3 (N5037, N5033, N2931, N2614);
and AND3 (N5038, N5027, N2482, N2206);
nand NAND2 (N5039, N5022, N2699);
buf BUF1 (N5040, N5034);
buf BUF1 (N5041, N5040);
or OR4 (N5042, N5035, N4500, N560, N4789);
nand NAND2 (N5043, N5031, N965);
nand NAND3 (N5044, N5010, N2420, N4017);
xor XOR2 (N5045, N5041, N4123);
xor XOR2 (N5046, N5042, N1832);
not NOT1 (N5047, N5044);
not NOT1 (N5048, N5043);
nor NOR2 (N5049, N5038, N844);
not NOT1 (N5050, N5037);
nor NOR2 (N5051, N5050, N3785);
nor NOR4 (N5052, N5039, N3329, N180, N1026);
nor NOR2 (N5053, N5048, N2825);
nor NOR3 (N5054, N5046, N3066, N1165);
and AND2 (N5055, N5030, N2805);
nor NOR3 (N5056, N5045, N1213, N4861);
buf BUF1 (N5057, N5054);
nor NOR4 (N5058, N5032, N2693, N379, N827);
or OR3 (N5059, N5057, N3612, N898);
xor XOR2 (N5060, N5049, N4052);
or OR3 (N5061, N5052, N1829, N1340);
buf BUF1 (N5062, N5053);
not NOT1 (N5063, N5060);
and AND3 (N5064, N5063, N3049, N991);
nand NAND2 (N5065, N5058, N3717);
nand NAND2 (N5066, N5056, N4471);
not NOT1 (N5067, N5055);
not NOT1 (N5068, N5064);
or OR2 (N5069, N5068, N3759);
nand NAND2 (N5070, N5047, N3733);
buf BUF1 (N5071, N5067);
and AND2 (N5072, N5061, N1577);
not NOT1 (N5073, N5059);
buf BUF1 (N5074, N5051);
or OR3 (N5075, N5066, N2576, N1081);
and AND3 (N5076, N5070, N1053, N4241);
and AND3 (N5077, N5065, N4211, N1865);
nand NAND3 (N5078, N5071, N2400, N3462);
or OR2 (N5079, N5073, N1249);
or OR4 (N5080, N5076, N448, N542, N693);
nand NAND2 (N5081, N5074, N1113);
nor NOR2 (N5082, N5079, N683);
and AND3 (N5083, N5081, N543, N3121);
not NOT1 (N5084, N5069);
nand NAND2 (N5085, N5078, N4495);
nand NAND2 (N5086, N5083, N1594);
nand NAND3 (N5087, N5072, N628, N2737);
or OR3 (N5088, N5062, N3496, N2415);
or OR2 (N5089, N5080, N4089);
or OR2 (N5090, N5086, N2803);
nand NAND2 (N5091, N5036, N4878);
not NOT1 (N5092, N5085);
and AND4 (N5093, N5089, N442, N2453, N44);
nor NOR3 (N5094, N5082, N938, N1524);
and AND2 (N5095, N5093, N4908);
xor XOR2 (N5096, N5090, N1838);
nand NAND4 (N5097, N5091, N233, N3355, N998);
buf BUF1 (N5098, N5097);
and AND4 (N5099, N5075, N3740, N209, N3753);
nand NAND2 (N5100, N5092, N3178);
nand NAND3 (N5101, N5100, N5003, N2101);
nor NOR4 (N5102, N5088, N4750, N2511, N2761);
not NOT1 (N5103, N5096);
and AND2 (N5104, N5087, N1690);
or OR3 (N5105, N5084, N706, N1505);
not NOT1 (N5106, N5099);
or OR4 (N5107, N5103, N3628, N2195, N1556);
nand NAND2 (N5108, N5106, N1577);
xor XOR2 (N5109, N5102, N3262);
and AND4 (N5110, N5104, N4386, N3961, N3810);
nor NOR2 (N5111, N5105, N4952);
not NOT1 (N5112, N5077);
not NOT1 (N5113, N5107);
and AND2 (N5114, N5098, N1528);
buf BUF1 (N5115, N5108);
buf BUF1 (N5116, N5109);
xor XOR2 (N5117, N5111, N1068);
buf BUF1 (N5118, N5110);
xor XOR2 (N5119, N5101, N4351);
nor NOR4 (N5120, N5113, N3775, N847, N2849);
or OR3 (N5121, N5120, N1889, N3723);
nor NOR3 (N5122, N5094, N3932, N388);
or OR2 (N5123, N5115, N1053);
xor XOR2 (N5124, N5122, N3766);
xor XOR2 (N5125, N5121, N260);
nor NOR4 (N5126, N5125, N4407, N3153, N3379);
not NOT1 (N5127, N5114);
buf BUF1 (N5128, N5124);
buf BUF1 (N5129, N5116);
xor XOR2 (N5130, N5095, N2945);
and AND4 (N5131, N5123, N3700, N81, N4563);
not NOT1 (N5132, N5128);
and AND2 (N5133, N5130, N1894);
or OR2 (N5134, N5129, N4803);
or OR3 (N5135, N5126, N688, N2721);
nand NAND3 (N5136, N5117, N3590, N2566);
xor XOR2 (N5137, N5131, N2268);
not NOT1 (N5138, N5118);
or OR2 (N5139, N5112, N3240);
xor XOR2 (N5140, N5138, N2043);
and AND4 (N5141, N5140, N2921, N4231, N688);
or OR4 (N5142, N5119, N224, N5124, N2787);
nor NOR4 (N5143, N5135, N3718, N4142, N3710);
xor XOR2 (N5144, N5142, N4131);
nand NAND2 (N5145, N5143, N5097);
and AND3 (N5146, N5144, N2898, N2925);
not NOT1 (N5147, N5139);
nor NOR3 (N5148, N5137, N4044, N873);
or OR2 (N5149, N5146, N1263);
buf BUF1 (N5150, N5147);
and AND4 (N5151, N5150, N1936, N1862, N3281);
nand NAND4 (N5152, N5133, N1983, N1813, N5090);
not NOT1 (N5153, N5151);
buf BUF1 (N5154, N5149);
or OR3 (N5155, N5132, N483, N2468);
nand NAND3 (N5156, N5148, N3022, N1245);
not NOT1 (N5157, N5153);
and AND3 (N5158, N5157, N1500, N2175);
xor XOR2 (N5159, N5158, N3665);
nor NOR2 (N5160, N5152, N1031);
xor XOR2 (N5161, N5136, N855);
and AND2 (N5162, N5161, N1119);
nand NAND2 (N5163, N5155, N3256);
nor NOR3 (N5164, N5127, N1128, N3308);
and AND4 (N5165, N5145, N2050, N3392, N4018);
xor XOR2 (N5166, N5134, N1303);
and AND3 (N5167, N5164, N4133, N795);
nor NOR4 (N5168, N5163, N1160, N3144, N4798);
xor XOR2 (N5169, N5168, N5024);
not NOT1 (N5170, N5165);
buf BUF1 (N5171, N5156);
nor NOR3 (N5172, N5160, N1289, N2172);
and AND3 (N5173, N5166, N2985, N841);
and AND2 (N5174, N5171, N3531);
not NOT1 (N5175, N5167);
nor NOR2 (N5176, N5172, N3946);
not NOT1 (N5177, N5175);
buf BUF1 (N5178, N5173);
and AND4 (N5179, N5159, N308, N3777, N3971);
xor XOR2 (N5180, N5179, N4597);
and AND4 (N5181, N5178, N4724, N1548, N1771);
not NOT1 (N5182, N5169);
or OR3 (N5183, N5182, N1547, N1754);
or OR3 (N5184, N5176, N649, N3409);
not NOT1 (N5185, N5141);
and AND2 (N5186, N5184, N4494);
not NOT1 (N5187, N5180);
or OR4 (N5188, N5187, N152, N1110, N131);
buf BUF1 (N5189, N5162);
and AND3 (N5190, N5174, N3285, N3192);
xor XOR2 (N5191, N5185, N1672);
not NOT1 (N5192, N5170);
buf BUF1 (N5193, N5183);
not NOT1 (N5194, N5189);
and AND2 (N5195, N5186, N4790);
not NOT1 (N5196, N5154);
or OR4 (N5197, N5177, N4698, N567, N1948);
nand NAND4 (N5198, N5181, N3621, N2453, N3342);
nor NOR4 (N5199, N5195, N3247, N2681, N41);
nor NOR3 (N5200, N5197, N4773, N4543);
or OR2 (N5201, N5191, N128);
xor XOR2 (N5202, N5201, N4689);
and AND3 (N5203, N5192, N1487, N3292);
and AND4 (N5204, N5196, N3765, N2737, N2687);
or OR2 (N5205, N5203, N674);
xor XOR2 (N5206, N5198, N2657);
nand NAND2 (N5207, N5194, N1839);
buf BUF1 (N5208, N5200);
or OR4 (N5209, N5202, N2836, N662, N2262);
nor NOR4 (N5210, N5190, N3335, N4695, N952);
or OR2 (N5211, N5210, N985);
or OR4 (N5212, N5205, N3430, N1490, N389);
xor XOR2 (N5213, N5193, N3581);
buf BUF1 (N5214, N5212);
xor XOR2 (N5215, N5188, N1965);
nor NOR2 (N5216, N5206, N3774);
buf BUF1 (N5217, N5214);
buf BUF1 (N5218, N5209);
xor XOR2 (N5219, N5213, N5085);
buf BUF1 (N5220, N5211);
xor XOR2 (N5221, N5219, N1038);
nor NOR4 (N5222, N5208, N1307, N3308, N2579);
nor NOR2 (N5223, N5215, N3587);
nor NOR3 (N5224, N5199, N268, N474);
buf BUF1 (N5225, N5222);
nand NAND4 (N5226, N5225, N787, N4542, N2105);
nor NOR2 (N5227, N5226, N4240);
and AND4 (N5228, N5220, N4189, N538, N1015);
xor XOR2 (N5229, N5207, N469);
buf BUF1 (N5230, N5216);
nand NAND4 (N5231, N5227, N1174, N2568, N675);
xor XOR2 (N5232, N5218, N789);
not NOT1 (N5233, N5228);
nand NAND2 (N5234, N5229, N511);
nor NOR3 (N5235, N5223, N3660, N289);
not NOT1 (N5236, N5232);
or OR4 (N5237, N5234, N1293, N2757, N4700);
not NOT1 (N5238, N5231);
nand NAND3 (N5239, N5236, N4519, N1858);
xor XOR2 (N5240, N5221, N1104);
nor NOR4 (N5241, N5238, N570, N1699, N790);
buf BUF1 (N5242, N5217);
not NOT1 (N5243, N5240);
nor NOR4 (N5244, N5242, N1433, N577, N340);
nand NAND4 (N5245, N5244, N4607, N738, N3059);
and AND4 (N5246, N5245, N2838, N3751, N4994);
xor XOR2 (N5247, N5204, N3390);
and AND4 (N5248, N5246, N777, N3849, N1319);
buf BUF1 (N5249, N5241);
and AND3 (N5250, N5224, N905, N2319);
xor XOR2 (N5251, N5230, N282);
nor NOR3 (N5252, N5237, N4039, N3598);
xor XOR2 (N5253, N5239, N862);
buf BUF1 (N5254, N5247);
nor NOR3 (N5255, N5250, N2792, N208);
buf BUF1 (N5256, N5253);
nor NOR4 (N5257, N5252, N4291, N150, N4176);
buf BUF1 (N5258, N5254);
not NOT1 (N5259, N5256);
nor NOR2 (N5260, N5255, N4792);
xor XOR2 (N5261, N5249, N3166);
and AND4 (N5262, N5248, N3327, N3063, N532);
nand NAND2 (N5263, N5235, N144);
nand NAND3 (N5264, N5258, N1272, N2242);
xor XOR2 (N5265, N5257, N1546);
nor NOR4 (N5266, N5251, N50, N1834, N3266);
xor XOR2 (N5267, N5265, N1982);
not NOT1 (N5268, N5233);
and AND3 (N5269, N5267, N4093, N595);
not NOT1 (N5270, N5261);
buf BUF1 (N5271, N5268);
and AND3 (N5272, N5260, N241, N1082);
or OR3 (N5273, N5270, N54, N3319);
not NOT1 (N5274, N5272);
xor XOR2 (N5275, N5262, N1694);
buf BUF1 (N5276, N5271);
xor XOR2 (N5277, N5266, N4268);
not NOT1 (N5278, N5275);
nand NAND3 (N5279, N5269, N3029, N432);
nand NAND2 (N5280, N5279, N490);
xor XOR2 (N5281, N5277, N2490);
xor XOR2 (N5282, N5276, N4926);
xor XOR2 (N5283, N5273, N2302);
or OR3 (N5284, N5283, N1550, N2373);
not NOT1 (N5285, N5281);
xor XOR2 (N5286, N5274, N1256);
buf BUF1 (N5287, N5280);
buf BUF1 (N5288, N5264);
nand NAND3 (N5289, N5285, N4378, N4064);
nand NAND2 (N5290, N5289, N1332);
not NOT1 (N5291, N5286);
nand NAND2 (N5292, N5291, N3208);
or OR4 (N5293, N5284, N2230, N592, N3585);
or OR3 (N5294, N5293, N5009, N3471);
not NOT1 (N5295, N5294);
nor NOR2 (N5296, N5292, N772);
nor NOR2 (N5297, N5288, N585);
or OR4 (N5298, N5295, N4396, N928, N2059);
nand NAND3 (N5299, N5243, N5151, N5289);
or OR2 (N5300, N5282, N4708);
not NOT1 (N5301, N5298);
nand NAND4 (N5302, N5290, N3831, N107, N3615);
buf BUF1 (N5303, N5296);
buf BUF1 (N5304, N5299);
and AND2 (N5305, N5304, N2338);
nor NOR3 (N5306, N5302, N2836, N3511);
nand NAND4 (N5307, N5306, N4425, N4565, N1590);
xor XOR2 (N5308, N5300, N1709);
nor NOR4 (N5309, N5305, N2318, N10, N1987);
buf BUF1 (N5310, N5263);
or OR2 (N5311, N5259, N2530);
nor NOR4 (N5312, N5303, N821, N2725, N901);
buf BUF1 (N5313, N5307);
not NOT1 (N5314, N5309);
buf BUF1 (N5315, N5313);
nand NAND3 (N5316, N5311, N3997, N3448);
nor NOR2 (N5317, N5315, N2090);
buf BUF1 (N5318, N5278);
nand NAND2 (N5319, N5316, N5159);
buf BUF1 (N5320, N5312);
or OR3 (N5321, N5287, N4547, N850);
and AND3 (N5322, N5297, N5074, N3048);
buf BUF1 (N5323, N5317);
xor XOR2 (N5324, N5310, N3676);
buf BUF1 (N5325, N5324);
or OR2 (N5326, N5319, N2362);
xor XOR2 (N5327, N5322, N4240);
not NOT1 (N5328, N5321);
not NOT1 (N5329, N5325);
or OR2 (N5330, N5327, N1130);
nand NAND3 (N5331, N5323, N613, N2274);
or OR2 (N5332, N5329, N3352);
and AND3 (N5333, N5326, N4390, N379);
nand NAND4 (N5334, N5332, N1057, N1297, N3142);
nand NAND4 (N5335, N5331, N3790, N5258, N3920);
and AND3 (N5336, N5320, N360, N1146);
or OR4 (N5337, N5301, N1457, N2948, N2851);
xor XOR2 (N5338, N5335, N2169);
xor XOR2 (N5339, N5330, N3993);
nand NAND2 (N5340, N5334, N4561);
nand NAND3 (N5341, N5314, N2858, N2868);
or OR3 (N5342, N5339, N3479, N972);
nand NAND4 (N5343, N5342, N4690, N1241, N667);
or OR2 (N5344, N5337, N4922);
xor XOR2 (N5345, N5318, N5061);
not NOT1 (N5346, N5340);
or OR4 (N5347, N5343, N2712, N3766, N2526);
or OR4 (N5348, N5344, N1809, N1163, N3828);
nand NAND4 (N5349, N5345, N384, N2194, N704);
xor XOR2 (N5350, N5328, N1747);
buf BUF1 (N5351, N5348);
nand NAND4 (N5352, N5336, N4546, N4677, N1549);
or OR2 (N5353, N5352, N1333);
and AND2 (N5354, N5341, N4137);
or OR4 (N5355, N5350, N1148, N4191, N1303);
nand NAND2 (N5356, N5338, N3602);
buf BUF1 (N5357, N5347);
buf BUF1 (N5358, N5353);
xor XOR2 (N5359, N5357, N782);
buf BUF1 (N5360, N5354);
buf BUF1 (N5361, N5360);
nand NAND4 (N5362, N5333, N5085, N25, N571);
not NOT1 (N5363, N5361);
nand NAND4 (N5364, N5308, N481, N3994, N2932);
not NOT1 (N5365, N5346);
buf BUF1 (N5366, N5356);
or OR4 (N5367, N5359, N1332, N2121, N4301);
and AND2 (N5368, N5362, N4088);
not NOT1 (N5369, N5364);
nand NAND4 (N5370, N5349, N1800, N578, N1316);
xor XOR2 (N5371, N5365, N602);
nand NAND4 (N5372, N5368, N2805, N4676, N797);
nand NAND4 (N5373, N5369, N1554, N803, N1173);
nand NAND4 (N5374, N5371, N3737, N3562, N2976);
buf BUF1 (N5375, N5372);
and AND2 (N5376, N5366, N2331);
xor XOR2 (N5377, N5376, N1152);
xor XOR2 (N5378, N5375, N3537);
buf BUF1 (N5379, N5378);
not NOT1 (N5380, N5358);
and AND2 (N5381, N5355, N1878);
or OR3 (N5382, N5370, N1982, N1219);
and AND4 (N5383, N5381, N1279, N5109, N5101);
nand NAND4 (N5384, N5383, N2741, N2330, N4296);
or OR4 (N5385, N5382, N74, N1294, N2602);
nor NOR2 (N5386, N5374, N1077);
buf BUF1 (N5387, N5351);
nor NOR2 (N5388, N5379, N4720);
and AND3 (N5389, N5387, N296, N2020);
not NOT1 (N5390, N5373);
buf BUF1 (N5391, N5384);
and AND3 (N5392, N5388, N4268, N5124);
not NOT1 (N5393, N5377);
xor XOR2 (N5394, N5367, N1134);
or OR4 (N5395, N5394, N3993, N1963, N1509);
xor XOR2 (N5396, N5386, N1857);
buf BUF1 (N5397, N5380);
and AND2 (N5398, N5389, N4986);
xor XOR2 (N5399, N5395, N3400);
nand NAND4 (N5400, N5391, N3707, N16, N3907);
not NOT1 (N5401, N5385);
or OR2 (N5402, N5400, N864);
not NOT1 (N5403, N5402);
nor NOR3 (N5404, N5399, N1829, N4705);
nor NOR3 (N5405, N5392, N4436, N645);
xor XOR2 (N5406, N5390, N4383);
or OR4 (N5407, N5363, N1138, N3793, N1322);
or OR3 (N5408, N5403, N3614, N1757);
nand NAND4 (N5409, N5396, N2795, N4347, N1780);
buf BUF1 (N5410, N5393);
not NOT1 (N5411, N5398);
not NOT1 (N5412, N5406);
nand NAND3 (N5413, N5404, N2561, N1626);
nand NAND4 (N5414, N5401, N3426, N3819, N3273);
xor XOR2 (N5415, N5413, N5316);
xor XOR2 (N5416, N5411, N1466);
xor XOR2 (N5417, N5415, N2519);
xor XOR2 (N5418, N5416, N1100);
and AND4 (N5419, N5414, N2550, N2759, N2854);
buf BUF1 (N5420, N5419);
or OR2 (N5421, N5408, N280);
or OR2 (N5422, N5418, N2271);
xor XOR2 (N5423, N5422, N669);
nand NAND4 (N5424, N5407, N600, N3789, N3382);
buf BUF1 (N5425, N5410);
xor XOR2 (N5426, N5405, N329);
nand NAND4 (N5427, N5424, N268, N2113, N3233);
nor NOR4 (N5428, N5423, N4725, N4670, N2047);
and AND4 (N5429, N5412, N966, N358, N2468);
buf BUF1 (N5430, N5425);
or OR3 (N5431, N5421, N4382, N438);
nand NAND4 (N5432, N5431, N818, N234, N5366);
nor NOR4 (N5433, N5426, N2462, N474, N2642);
buf BUF1 (N5434, N5427);
or OR4 (N5435, N5429, N277, N63, N4845);
or OR3 (N5436, N5420, N1777, N1466);
or OR4 (N5437, N5417, N2177, N3730, N2086);
and AND4 (N5438, N5432, N1383, N1075, N852);
xor XOR2 (N5439, N5433, N778);
or OR2 (N5440, N5428, N2657);
nor NOR2 (N5441, N5435, N1265);
nand NAND2 (N5442, N5430, N1136);
buf BUF1 (N5443, N5434);
or OR3 (N5444, N5409, N2542, N1671);
not NOT1 (N5445, N5441);
xor XOR2 (N5446, N5444, N3100);
not NOT1 (N5447, N5439);
nand NAND4 (N5448, N5437, N2232, N4784, N2350);
nand NAND2 (N5449, N5445, N2759);
not NOT1 (N5450, N5442);
buf BUF1 (N5451, N5448);
xor XOR2 (N5452, N5447, N878);
xor XOR2 (N5453, N5452, N2609);
nand NAND2 (N5454, N5440, N2127);
and AND4 (N5455, N5450, N4107, N4863, N2218);
xor XOR2 (N5456, N5436, N3227);
nor NOR3 (N5457, N5446, N4956, N2102);
buf BUF1 (N5458, N5443);
buf BUF1 (N5459, N5453);
buf BUF1 (N5460, N5438);
not NOT1 (N5461, N5458);
and AND4 (N5462, N5455, N1439, N2602, N4819);
not NOT1 (N5463, N5457);
xor XOR2 (N5464, N5449, N1885);
or OR4 (N5465, N5463, N2858, N964, N5037);
nor NOR4 (N5466, N5451, N715, N3130, N5337);
buf BUF1 (N5467, N5462);
xor XOR2 (N5468, N5461, N2023);
not NOT1 (N5469, N5460);
xor XOR2 (N5470, N5468, N2613);
xor XOR2 (N5471, N5466, N1522);
nor NOR2 (N5472, N5464, N2787);
buf BUF1 (N5473, N5456);
not NOT1 (N5474, N5467);
nand NAND4 (N5475, N5469, N3126, N4808, N2686);
and AND2 (N5476, N5475, N2572);
xor XOR2 (N5477, N5471, N300);
not NOT1 (N5478, N5472);
not NOT1 (N5479, N5476);
nand NAND4 (N5480, N5397, N5433, N1168, N2094);
nand NAND2 (N5481, N5465, N1159);
nor NOR2 (N5482, N5478, N1737);
or OR3 (N5483, N5474, N5240, N4977);
not NOT1 (N5484, N5454);
xor XOR2 (N5485, N5477, N5027);
and AND2 (N5486, N5483, N4847);
nand NAND2 (N5487, N5485, N4688);
buf BUF1 (N5488, N5484);
or OR3 (N5489, N5479, N3827, N2036);
nor NOR2 (N5490, N5482, N3906);
not NOT1 (N5491, N5490);
buf BUF1 (N5492, N5480);
nor NOR4 (N5493, N5492, N2795, N13, N3547);
nor NOR4 (N5494, N5473, N488, N3361, N429);
and AND4 (N5495, N5493, N1021, N1756, N1239);
or OR4 (N5496, N5488, N4946, N5111, N2041);
and AND4 (N5497, N5486, N4528, N4390, N1479);
nor NOR3 (N5498, N5496, N937, N1595);
nand NAND4 (N5499, N5497, N3500, N2502, N2537);
and AND4 (N5500, N5459, N3127, N2904, N2928);
nand NAND4 (N5501, N5494, N2832, N4076, N5141);
buf BUF1 (N5502, N5489);
nor NOR3 (N5503, N5500, N1020, N1419);
xor XOR2 (N5504, N5491, N3156);
nor NOR4 (N5505, N5481, N999, N4288, N4382);
nor NOR4 (N5506, N5503, N1804, N2067, N5404);
nor NOR4 (N5507, N5498, N5361, N3024, N182);
nor NOR4 (N5508, N5487, N3026, N1606, N4034);
xor XOR2 (N5509, N5499, N3265);
and AND3 (N5510, N5501, N3809, N3852);
buf BUF1 (N5511, N5495);
nor NOR4 (N5512, N5510, N5497, N1914, N3488);
and AND3 (N5513, N5502, N2225, N2172);
or OR4 (N5514, N5512, N3323, N1878, N2102);
nor NOR2 (N5515, N5511, N4462);
buf BUF1 (N5516, N5513);
xor XOR2 (N5517, N5507, N955);
nor NOR3 (N5518, N5516, N836, N2237);
or OR3 (N5519, N5505, N1925, N53);
or OR2 (N5520, N5518, N2023);
or OR2 (N5521, N5519, N1335);
xor XOR2 (N5522, N5508, N1027);
nand NAND3 (N5523, N5514, N2102, N3585);
xor XOR2 (N5524, N5515, N2156);
nor NOR3 (N5525, N5509, N477, N3994);
nor NOR3 (N5526, N5517, N2378, N1094);
xor XOR2 (N5527, N5526, N4647);
and AND3 (N5528, N5527, N4157, N2134);
and AND3 (N5529, N5524, N2067, N4010);
not NOT1 (N5530, N5528);
buf BUF1 (N5531, N5530);
not NOT1 (N5532, N5506);
not NOT1 (N5533, N5521);
xor XOR2 (N5534, N5531, N551);
or OR3 (N5535, N5520, N4374, N383);
nand NAND3 (N5536, N5523, N2880, N2784);
xor XOR2 (N5537, N5533, N358);
buf BUF1 (N5538, N5529);
nor NOR2 (N5539, N5536, N853);
nor NOR4 (N5540, N5470, N809, N2883, N126);
and AND2 (N5541, N5537, N4307);
nor NOR4 (N5542, N5538, N2832, N4178, N742);
buf BUF1 (N5543, N5541);
not NOT1 (N5544, N5522);
buf BUF1 (N5545, N5540);
nand NAND4 (N5546, N5535, N3970, N4552, N5392);
or OR4 (N5547, N5525, N1965, N423, N5508);
buf BUF1 (N5548, N5543);
xor XOR2 (N5549, N5544, N1467);
nor NOR4 (N5550, N5542, N4428, N1393, N1944);
nand NAND2 (N5551, N5546, N3231);
and AND2 (N5552, N5548, N4967);
xor XOR2 (N5553, N5550, N2714);
nor NOR2 (N5554, N5534, N4142);
nor NOR2 (N5555, N5545, N2796);
buf BUF1 (N5556, N5552);
buf BUF1 (N5557, N5539);
not NOT1 (N5558, N5532);
not NOT1 (N5559, N5547);
xor XOR2 (N5560, N5559, N267);
xor XOR2 (N5561, N5554, N5255);
and AND4 (N5562, N5555, N513, N4829, N2444);
xor XOR2 (N5563, N5561, N5272);
or OR3 (N5564, N5557, N4998, N2223);
not NOT1 (N5565, N5504);
nand NAND2 (N5566, N5565, N3738);
not NOT1 (N5567, N5556);
and AND4 (N5568, N5564, N3024, N4712, N668);
and AND2 (N5569, N5553, N272);
nor NOR2 (N5570, N5568, N2599);
nor NOR4 (N5571, N5569, N643, N3177, N872);
or OR2 (N5572, N5563, N5413);
nor NOR4 (N5573, N5570, N4496, N1887, N83);
nand NAND2 (N5574, N5573, N1713);
xor XOR2 (N5575, N5566, N97);
not NOT1 (N5576, N5558);
and AND4 (N5577, N5562, N562, N2045, N4101);
and AND2 (N5578, N5572, N5555);
and AND4 (N5579, N5567, N2600, N548, N5575);
not NOT1 (N5580, N3320);
xor XOR2 (N5581, N5578, N1414);
and AND2 (N5582, N5549, N4730);
or OR4 (N5583, N5580, N477, N2286, N2692);
xor XOR2 (N5584, N5582, N2835);
or OR4 (N5585, N5579, N4596, N3547, N5121);
nor NOR4 (N5586, N5571, N1838, N132, N4731);
and AND3 (N5587, N5577, N5403, N3097);
xor XOR2 (N5588, N5583, N1860);
or OR3 (N5589, N5560, N1871, N4062);
xor XOR2 (N5590, N5576, N1132);
or OR4 (N5591, N5590, N5440, N5293, N2243);
and AND3 (N5592, N5589, N4770, N1243);
buf BUF1 (N5593, N5585);
buf BUF1 (N5594, N5593);
nand NAND4 (N5595, N5587, N1756, N2437, N2711);
buf BUF1 (N5596, N5581);
not NOT1 (N5597, N5591);
not NOT1 (N5598, N5574);
or OR4 (N5599, N5592, N540, N1588, N829);
and AND2 (N5600, N5597, N2262);
xor XOR2 (N5601, N5596, N4589);
xor XOR2 (N5602, N5598, N4769);
nor NOR3 (N5603, N5602, N545, N2757);
buf BUF1 (N5604, N5601);
and AND4 (N5605, N5604, N2233, N1065, N4934);
not NOT1 (N5606, N5595);
not NOT1 (N5607, N5551);
and AND2 (N5608, N5584, N3343);
xor XOR2 (N5609, N5603, N4965);
or OR2 (N5610, N5607, N1443);
xor XOR2 (N5611, N5594, N4154);
nand NAND4 (N5612, N5606, N5515, N2242, N5062);
not NOT1 (N5613, N5611);
not NOT1 (N5614, N5586);
nor NOR2 (N5615, N5608, N5371);
xor XOR2 (N5616, N5614, N3341);
buf BUF1 (N5617, N5588);
xor XOR2 (N5618, N5612, N1386);
not NOT1 (N5619, N5617);
nand NAND3 (N5620, N5619, N4069, N3365);
xor XOR2 (N5621, N5620, N1703);
buf BUF1 (N5622, N5600);
buf BUF1 (N5623, N5609);
or OR4 (N5624, N5599, N4087, N5456, N695);
and AND3 (N5625, N5622, N3621, N2104);
nor NOR4 (N5626, N5623, N2956, N2790, N3921);
xor XOR2 (N5627, N5613, N4083);
nand NAND3 (N5628, N5610, N3994, N3291);
or OR4 (N5629, N5616, N3902, N136, N4796);
not NOT1 (N5630, N5628);
and AND2 (N5631, N5615, N3027);
xor XOR2 (N5632, N5605, N3831);
xor XOR2 (N5633, N5625, N4016);
buf BUF1 (N5634, N5627);
and AND4 (N5635, N5630, N1744, N1459, N2694);
or OR2 (N5636, N5631, N4698);
or OR3 (N5637, N5618, N387, N3399);
xor XOR2 (N5638, N5635, N3536);
not NOT1 (N5639, N5637);
nor NOR3 (N5640, N5636, N2895, N328);
not NOT1 (N5641, N5621);
and AND4 (N5642, N5633, N4333, N5296, N2995);
and AND4 (N5643, N5641, N758, N3025, N4854);
buf BUF1 (N5644, N5640);
or OR2 (N5645, N5644, N2052);
xor XOR2 (N5646, N5626, N2588);
and AND2 (N5647, N5645, N3733);
buf BUF1 (N5648, N5642);
or OR4 (N5649, N5632, N5134, N2816, N3759);
not NOT1 (N5650, N5643);
not NOT1 (N5651, N5649);
xor XOR2 (N5652, N5634, N3474);
not NOT1 (N5653, N5624);
or OR2 (N5654, N5638, N4895);
nor NOR2 (N5655, N5654, N3431);
not NOT1 (N5656, N5647);
or OR4 (N5657, N5648, N4709, N4865, N3575);
nand NAND2 (N5658, N5639, N4110);
buf BUF1 (N5659, N5658);
not NOT1 (N5660, N5653);
nor NOR2 (N5661, N5659, N1335);
not NOT1 (N5662, N5655);
not NOT1 (N5663, N5662);
nand NAND3 (N5664, N5656, N1070, N5394);
not NOT1 (N5665, N5657);
not NOT1 (N5666, N5646);
buf BUF1 (N5667, N5660);
xor XOR2 (N5668, N5665, N5593);
xor XOR2 (N5669, N5668, N393);
or OR3 (N5670, N5661, N1955, N1572);
and AND3 (N5671, N5650, N3591, N3246);
and AND3 (N5672, N5670, N1905, N4645);
nand NAND2 (N5673, N5651, N3460);
buf BUF1 (N5674, N5672);
not NOT1 (N5675, N5671);
not NOT1 (N5676, N5652);
nand NAND2 (N5677, N5629, N1310);
or OR4 (N5678, N5673, N2985, N4429, N2643);
not NOT1 (N5679, N5675);
nor NOR2 (N5680, N5678, N2568);
not NOT1 (N5681, N5674);
or OR2 (N5682, N5677, N4469);
nor NOR2 (N5683, N5679, N1671);
or OR3 (N5684, N5666, N1822, N1383);
and AND4 (N5685, N5663, N3073, N5335, N3858);
nor NOR3 (N5686, N5683, N4350, N2513);
nor NOR4 (N5687, N5667, N4342, N3819, N4302);
nor NOR3 (N5688, N5669, N2012, N2900);
nand NAND2 (N5689, N5685, N567);
nand NAND3 (N5690, N5680, N2348, N3965);
nand NAND3 (N5691, N5689, N4620, N3675);
nand NAND4 (N5692, N5664, N3183, N3758, N1345);
nand NAND2 (N5693, N5687, N5496);
and AND4 (N5694, N5686, N1082, N2188, N5581);
or OR3 (N5695, N5684, N2827, N1165);
xor XOR2 (N5696, N5688, N515);
or OR4 (N5697, N5682, N3184, N4780, N208);
or OR2 (N5698, N5690, N3194);
not NOT1 (N5699, N5693);
nand NAND2 (N5700, N5696, N3762);
nand NAND4 (N5701, N5692, N2665, N2702, N540);
not NOT1 (N5702, N5676);
nor NOR3 (N5703, N5691, N2076, N2008);
and AND4 (N5704, N5703, N2632, N2477, N3551);
buf BUF1 (N5705, N5702);
buf BUF1 (N5706, N5695);
or OR2 (N5707, N5681, N1518);
and AND2 (N5708, N5694, N2546);
or OR3 (N5709, N5701, N5339, N2945);
or OR2 (N5710, N5706, N2112);
nand NAND2 (N5711, N5704, N1363);
and AND4 (N5712, N5700, N99, N1958, N2036);
buf BUF1 (N5713, N5699);
xor XOR2 (N5714, N5711, N3186);
not NOT1 (N5715, N5707);
not NOT1 (N5716, N5697);
xor XOR2 (N5717, N5709, N4689);
and AND3 (N5718, N5714, N5016, N1270);
xor XOR2 (N5719, N5717, N4998);
nand NAND4 (N5720, N5718, N1786, N306, N4633);
nand NAND2 (N5721, N5710, N1233);
nand NAND2 (N5722, N5698, N5602);
buf BUF1 (N5723, N5713);
buf BUF1 (N5724, N5720);
nor NOR3 (N5725, N5722, N5283, N3143);
not NOT1 (N5726, N5721);
xor XOR2 (N5727, N5705, N2946);
or OR3 (N5728, N5715, N724, N4702);
xor XOR2 (N5729, N5724, N326);
not NOT1 (N5730, N5708);
xor XOR2 (N5731, N5719, N4008);
and AND4 (N5732, N5727, N83, N5228, N5429);
and AND4 (N5733, N5729, N3429, N2469, N3700);
buf BUF1 (N5734, N5733);
xor XOR2 (N5735, N5734, N2090);
buf BUF1 (N5736, N5728);
nand NAND3 (N5737, N5730, N2361, N330);
or OR2 (N5738, N5712, N5305);
nand NAND4 (N5739, N5736, N2130, N5576, N61);
nand NAND3 (N5740, N5731, N1983, N134);
buf BUF1 (N5741, N5716);
or OR2 (N5742, N5740, N772);
or OR4 (N5743, N5738, N4984, N1378, N5041);
and AND3 (N5744, N5743, N4610, N5108);
nand NAND2 (N5745, N5744, N2721);
nand NAND4 (N5746, N5737, N2123, N4398, N134);
not NOT1 (N5747, N5725);
not NOT1 (N5748, N5741);
xor XOR2 (N5749, N5735, N2703);
buf BUF1 (N5750, N5742);
or OR3 (N5751, N5723, N2891, N5649);
and AND3 (N5752, N5748, N5530, N4695);
or OR3 (N5753, N5752, N2771, N4916);
not NOT1 (N5754, N5739);
not NOT1 (N5755, N5749);
and AND4 (N5756, N5754, N344, N125, N3090);
and AND4 (N5757, N5751, N2567, N3829, N5050);
xor XOR2 (N5758, N5746, N1623);
nor NOR3 (N5759, N5758, N4766, N3112);
nand NAND4 (N5760, N5756, N1750, N1511, N2605);
or OR3 (N5761, N5732, N973, N1856);
nand NAND4 (N5762, N5745, N741, N1116, N217);
and AND3 (N5763, N5747, N3942, N2080);
xor XOR2 (N5764, N5759, N2160);
xor XOR2 (N5765, N5764, N2252);
xor XOR2 (N5766, N5726, N5550);
and AND3 (N5767, N5755, N1700, N981);
xor XOR2 (N5768, N5760, N3722);
nor NOR2 (N5769, N5766, N4205);
buf BUF1 (N5770, N5765);
buf BUF1 (N5771, N5757);
or OR3 (N5772, N5762, N4998, N1719);
not NOT1 (N5773, N5763);
or OR4 (N5774, N5761, N4205, N818, N5716);
nor NOR4 (N5775, N5770, N5589, N1522, N1138);
buf BUF1 (N5776, N5773);
nand NAND2 (N5777, N5768, N4251);
and AND4 (N5778, N5772, N1358, N4666, N4067);
or OR4 (N5779, N5778, N2847, N5675, N4624);
and AND4 (N5780, N5774, N2654, N3264, N885);
or OR4 (N5781, N5775, N4149, N2696, N2578);
not NOT1 (N5782, N5781);
nand NAND2 (N5783, N5750, N637);
or OR2 (N5784, N5780, N5120);
nand NAND2 (N5785, N5779, N3252);
not NOT1 (N5786, N5785);
xor XOR2 (N5787, N5784, N5133);
xor XOR2 (N5788, N5782, N3717);
xor XOR2 (N5789, N5753, N3563);
and AND3 (N5790, N5769, N2937, N5560);
xor XOR2 (N5791, N5777, N597);
nor NOR4 (N5792, N5776, N2540, N4996, N5422);
buf BUF1 (N5793, N5788);
buf BUF1 (N5794, N5790);
buf BUF1 (N5795, N5792);
or OR2 (N5796, N5787, N4735);
and AND4 (N5797, N5791, N2691, N1894, N4789);
and AND3 (N5798, N5796, N5588, N4130);
not NOT1 (N5799, N5794);
or OR3 (N5800, N5797, N3154, N4573);
xor XOR2 (N5801, N5798, N2284);
or OR2 (N5802, N5800, N2399);
or OR2 (N5803, N5793, N2741);
buf BUF1 (N5804, N5783);
not NOT1 (N5805, N5767);
buf BUF1 (N5806, N5799);
not NOT1 (N5807, N5789);
and AND2 (N5808, N5802, N2418);
not NOT1 (N5809, N5808);
not NOT1 (N5810, N5771);
nor NOR3 (N5811, N5806, N5515, N3209);
nand NAND3 (N5812, N5809, N960, N2594);
and AND3 (N5813, N5812, N3871, N4717);
not NOT1 (N5814, N5807);
not NOT1 (N5815, N5811);
or OR4 (N5816, N5803, N3127, N4621, N1381);
and AND3 (N5817, N5801, N2242, N4916);
nand NAND3 (N5818, N5814, N2746, N3501);
buf BUF1 (N5819, N5816);
or OR3 (N5820, N5813, N24, N623);
nand NAND2 (N5821, N5786, N1348);
nor NOR3 (N5822, N5804, N2493, N1456);
nand NAND3 (N5823, N5805, N690, N3441);
nor NOR2 (N5824, N5820, N4878);
or OR3 (N5825, N5818, N3098, N1147);
nand NAND2 (N5826, N5825, N2105);
nor NOR2 (N5827, N5822, N425);
or OR4 (N5828, N5817, N3254, N2086, N5739);
nand NAND3 (N5829, N5821, N2036, N404);
or OR4 (N5830, N5828, N4012, N3908, N2411);
xor XOR2 (N5831, N5823, N3532);
not NOT1 (N5832, N5827);
xor XOR2 (N5833, N5829, N1222);
and AND3 (N5834, N5830, N3897, N2856);
nor NOR3 (N5835, N5810, N4896, N378);
nor NOR4 (N5836, N5831, N5231, N5600, N5444);
nor NOR3 (N5837, N5835, N4582, N5461);
buf BUF1 (N5838, N5826);
nand NAND2 (N5839, N5832, N3139);
not NOT1 (N5840, N5819);
buf BUF1 (N5841, N5839);
xor XOR2 (N5842, N5837, N2233);
xor XOR2 (N5843, N5815, N3921);
buf BUF1 (N5844, N5833);
not NOT1 (N5845, N5840);
xor XOR2 (N5846, N5845, N2662);
nand NAND3 (N5847, N5843, N4751, N1260);
nor NOR4 (N5848, N5836, N3724, N660, N1201);
buf BUF1 (N5849, N5824);
or OR4 (N5850, N5841, N68, N5247, N5415);
and AND3 (N5851, N5838, N4826, N2414);
nor NOR2 (N5852, N5795, N4731);
nor NOR3 (N5853, N5847, N5715, N835);
buf BUF1 (N5854, N5844);
and AND4 (N5855, N5842, N3750, N1469, N1867);
and AND2 (N5856, N5846, N1229);
buf BUF1 (N5857, N5848);
nor NOR3 (N5858, N5834, N2461, N4534);
or OR2 (N5859, N5856, N3712);
not NOT1 (N5860, N5859);
not NOT1 (N5861, N5855);
not NOT1 (N5862, N5849);
nor NOR2 (N5863, N5857, N932);
nor NOR3 (N5864, N5861, N3169, N469);
nor NOR4 (N5865, N5852, N1025, N2660, N675);
buf BUF1 (N5866, N5865);
buf BUF1 (N5867, N5863);
nand NAND2 (N5868, N5858, N196);
nor NOR3 (N5869, N5867, N4655, N4905);
xor XOR2 (N5870, N5854, N3492);
nor NOR4 (N5871, N5866, N2697, N3347, N4136);
buf BUF1 (N5872, N5850);
not NOT1 (N5873, N5871);
nand NAND2 (N5874, N5864, N1457);
buf BUF1 (N5875, N5853);
xor XOR2 (N5876, N5868, N3133);
nor NOR4 (N5877, N5874, N372, N38, N2710);
nand NAND4 (N5878, N5862, N4749, N4711, N1638);
buf BUF1 (N5879, N5875);
and AND2 (N5880, N5877, N5756);
or OR4 (N5881, N5870, N2741, N5498, N4533);
and AND4 (N5882, N5881, N705, N3150, N3776);
or OR2 (N5883, N5873, N612);
or OR4 (N5884, N5869, N4772, N2637, N3443);
buf BUF1 (N5885, N5884);
not NOT1 (N5886, N5880);
nand NAND2 (N5887, N5879, N3773);
xor XOR2 (N5888, N5882, N1136);
not NOT1 (N5889, N5872);
or OR3 (N5890, N5878, N142, N5062);
buf BUF1 (N5891, N5860);
xor XOR2 (N5892, N5889, N2887);
xor XOR2 (N5893, N5887, N929);
xor XOR2 (N5894, N5893, N4045);
or OR2 (N5895, N5883, N1411);
and AND3 (N5896, N5885, N5688, N2865);
nand NAND4 (N5897, N5890, N2689, N5164, N1051);
or OR2 (N5898, N5888, N3987);
nand NAND4 (N5899, N5897, N5106, N1576, N356);
not NOT1 (N5900, N5899);
nor NOR2 (N5901, N5894, N2163);
nand NAND3 (N5902, N5876, N713, N4005);
nor NOR4 (N5903, N5895, N3209, N4976, N1552);
xor XOR2 (N5904, N5902, N3165);
and AND4 (N5905, N5898, N5892, N2116, N922);
nand NAND4 (N5906, N4316, N2159, N848, N4631);
xor XOR2 (N5907, N5904, N2475);
nand NAND2 (N5908, N5851, N401);
xor XOR2 (N5909, N5891, N2584);
xor XOR2 (N5910, N5906, N660);
xor XOR2 (N5911, N5896, N5566);
nand NAND4 (N5912, N5911, N2587, N4700, N3036);
xor XOR2 (N5913, N5909, N1127);
nor NOR4 (N5914, N5912, N4045, N2493, N4713);
or OR4 (N5915, N5886, N1980, N2776, N4373);
or OR3 (N5916, N5901, N5064, N3393);
nor NOR2 (N5917, N5900, N5808);
and AND3 (N5918, N5908, N4151, N152);
or OR4 (N5919, N5907, N3075, N2977, N3668);
xor XOR2 (N5920, N5916, N1206);
or OR4 (N5921, N5917, N1902, N640, N2617);
or OR3 (N5922, N5910, N4988, N4138);
xor XOR2 (N5923, N5905, N1236);
and AND2 (N5924, N5922, N2380);
nand NAND4 (N5925, N5918, N92, N1878, N1187);
and AND4 (N5926, N5924, N3714, N3155, N4715);
nor NOR2 (N5927, N5913, N2239);
not NOT1 (N5928, N5914);
nand NAND3 (N5929, N5915, N2491, N2925);
or OR3 (N5930, N5920, N3596, N4981);
and AND3 (N5931, N5926, N53, N5186);
nand NAND2 (N5932, N5929, N5775);
buf BUF1 (N5933, N5928);
not NOT1 (N5934, N5930);
or OR3 (N5935, N5927, N3633, N1092);
not NOT1 (N5936, N5933);
xor XOR2 (N5937, N5935, N563);
buf BUF1 (N5938, N5921);
nand NAND2 (N5939, N5931, N2642);
not NOT1 (N5940, N5919);
xor XOR2 (N5941, N5903, N5590);
xor XOR2 (N5942, N5923, N3895);
buf BUF1 (N5943, N5938);
buf BUF1 (N5944, N5941);
or OR2 (N5945, N5925, N4029);
nor NOR4 (N5946, N5937, N4920, N670, N1669);
xor XOR2 (N5947, N5934, N4002);
or OR2 (N5948, N5940, N3530);
nand NAND4 (N5949, N5939, N66, N5783, N4102);
buf BUF1 (N5950, N5947);
buf BUF1 (N5951, N5945);
nor NOR3 (N5952, N5942, N722, N5182);
nand NAND2 (N5953, N5946, N285);
or OR3 (N5954, N5944, N1534, N3374);
not NOT1 (N5955, N5948);
or OR2 (N5956, N5932, N3503);
nor NOR4 (N5957, N5949, N531, N2469, N772);
nor NOR4 (N5958, N5957, N1153, N461, N3354);
nand NAND3 (N5959, N5943, N3557, N5953);
nor NOR4 (N5960, N2415, N1240, N1268, N621);
nor NOR2 (N5961, N5956, N5854);
buf BUF1 (N5962, N5936);
xor XOR2 (N5963, N5951, N4780);
nor NOR3 (N5964, N5958, N2709, N4438);
buf BUF1 (N5965, N5954);
xor XOR2 (N5966, N5959, N1287);
nand NAND3 (N5967, N5964, N1825, N3409);
xor XOR2 (N5968, N5965, N240);
nor NOR4 (N5969, N5952, N1341, N3116, N442);
nand NAND4 (N5970, N5969, N4330, N2185, N3181);
buf BUF1 (N5971, N5966);
not NOT1 (N5972, N5961);
xor XOR2 (N5973, N5970, N1818);
or OR4 (N5974, N5972, N3508, N1142, N4964);
or OR4 (N5975, N5960, N2307, N1519, N2847);
nor NOR4 (N5976, N5974, N3328, N2858, N3111);
nor NOR2 (N5977, N5975, N1369);
and AND2 (N5978, N5962, N2959);
and AND3 (N5979, N5973, N1668, N2726);
xor XOR2 (N5980, N5978, N2578);
nand NAND2 (N5981, N5977, N1447);
not NOT1 (N5982, N5980);
xor XOR2 (N5983, N5982, N5914);
xor XOR2 (N5984, N5979, N900);
buf BUF1 (N5985, N5955);
not NOT1 (N5986, N5967);
xor XOR2 (N5987, N5968, N898);
nor NOR2 (N5988, N5984, N3116);
nand NAND2 (N5989, N5971, N3721);
buf BUF1 (N5990, N5963);
buf BUF1 (N5991, N5987);
nor NOR4 (N5992, N5986, N2669, N963, N2650);
buf BUF1 (N5993, N5989);
or OR2 (N5994, N5991, N243);
not NOT1 (N5995, N5976);
and AND3 (N5996, N5950, N3929, N1452);
not NOT1 (N5997, N5995);
not NOT1 (N5998, N5985);
not NOT1 (N5999, N5990);
xor XOR2 (N6000, N5983, N2657);
buf BUF1 (N6001, N5994);
and AND3 (N6002, N5988, N3450, N2419);
buf BUF1 (N6003, N6000);
not NOT1 (N6004, N5981);
nor NOR4 (N6005, N6001, N667, N1807, N1041);
not NOT1 (N6006, N6004);
nor NOR4 (N6007, N6002, N883, N2445, N5590);
and AND3 (N6008, N5999, N1271, N5763);
buf BUF1 (N6009, N6008);
nor NOR2 (N6010, N6003, N2500);
nand NAND4 (N6011, N5997, N951, N4858, N1011);
xor XOR2 (N6012, N6010, N518);
and AND3 (N6013, N5996, N58, N4119);
nor NOR2 (N6014, N6011, N3654);
and AND3 (N6015, N5992, N351, N1201);
and AND4 (N6016, N6015, N4589, N2330, N2298);
nand NAND2 (N6017, N5998, N1330);
buf BUF1 (N6018, N6009);
not NOT1 (N6019, N6018);
and AND4 (N6020, N6005, N4695, N295, N3780);
not NOT1 (N6021, N6020);
buf BUF1 (N6022, N6017);
or OR4 (N6023, N6022, N2754, N457, N1767);
or OR3 (N6024, N6012, N85, N281);
and AND2 (N6025, N6024, N4657);
nor NOR3 (N6026, N6021, N4677, N5248);
nor NOR4 (N6027, N6014, N5337, N691, N3139);
nand NAND3 (N6028, N6025, N1779, N5685);
buf BUF1 (N6029, N6019);
nor NOR3 (N6030, N6028, N167, N1597);
nand NAND3 (N6031, N6013, N2341, N1694);
or OR4 (N6032, N6029, N5906, N2705, N5566);
nor NOR3 (N6033, N6023, N3891, N2177);
not NOT1 (N6034, N6026);
or OR2 (N6035, N6034, N3492);
nor NOR2 (N6036, N6007, N3771);
xor XOR2 (N6037, N6032, N515);
and AND3 (N6038, N6006, N3249, N535);
xor XOR2 (N6039, N6036, N2508);
or OR3 (N6040, N6016, N3043, N3661);
or OR3 (N6041, N6027, N1800, N5708);
xor XOR2 (N6042, N6040, N2308);
xor XOR2 (N6043, N6038, N1953);
buf BUF1 (N6044, N6031);
xor XOR2 (N6045, N6043, N4244);
or OR3 (N6046, N5993, N1842, N1132);
or OR4 (N6047, N6035, N2345, N1270, N503);
nand NAND4 (N6048, N6046, N711, N5704, N3597);
and AND2 (N6049, N6048, N3387);
not NOT1 (N6050, N6042);
xor XOR2 (N6051, N6045, N2269);
buf BUF1 (N6052, N6041);
xor XOR2 (N6053, N6037, N4370);
nand NAND2 (N6054, N6049, N3491);
or OR2 (N6055, N6051, N4419);
xor XOR2 (N6056, N6052, N3125);
and AND4 (N6057, N6033, N3494, N5735, N4867);
not NOT1 (N6058, N6056);
buf BUF1 (N6059, N6039);
and AND4 (N6060, N6044, N3241, N1758, N1722);
and AND3 (N6061, N6057, N5602, N1720);
not NOT1 (N6062, N6059);
buf BUF1 (N6063, N6050);
not NOT1 (N6064, N6062);
not NOT1 (N6065, N6061);
and AND4 (N6066, N6030, N5713, N67, N70);
and AND4 (N6067, N6063, N4433, N1176, N5431);
nand NAND4 (N6068, N6064, N1154, N832, N1153);
buf BUF1 (N6069, N6066);
xor XOR2 (N6070, N6069, N2072);
and AND3 (N6071, N6065, N1650, N890);
xor XOR2 (N6072, N6060, N81);
nand NAND2 (N6073, N6058, N4703);
xor XOR2 (N6074, N6068, N4706);
and AND2 (N6075, N6054, N1042);
nand NAND2 (N6076, N6075, N1704);
nor NOR3 (N6077, N6055, N461, N414);
nor NOR4 (N6078, N6070, N2481, N1283, N4187);
nor NOR4 (N6079, N6076, N1421, N4721, N3335);
buf BUF1 (N6080, N6078);
nor NOR2 (N6081, N6073, N3784);
or OR4 (N6082, N6067, N1144, N4315, N2201);
or OR4 (N6083, N6071, N5885, N2455, N4637);
not NOT1 (N6084, N6077);
buf BUF1 (N6085, N6079);
and AND4 (N6086, N6082, N1892, N512, N16);
nand NAND3 (N6087, N6080, N1501, N2990);
or OR4 (N6088, N6072, N4018, N5259, N5412);
buf BUF1 (N6089, N6085);
nand NAND4 (N6090, N6083, N5551, N4268, N5009);
nand NAND4 (N6091, N6087, N1389, N3256, N2675);
nor NOR3 (N6092, N6074, N3498, N3900);
nand NAND4 (N6093, N6047, N5538, N1881, N534);
and AND3 (N6094, N6084, N2722, N5382);
xor XOR2 (N6095, N6053, N870);
nor NOR3 (N6096, N6090, N3641, N4027);
nand NAND2 (N6097, N6094, N2343);
or OR4 (N6098, N6093, N645, N5675, N4797);
not NOT1 (N6099, N6088);
xor XOR2 (N6100, N6096, N4464);
buf BUF1 (N6101, N6092);
buf BUF1 (N6102, N6101);
not NOT1 (N6103, N6098);
or OR2 (N6104, N6100, N5627);
nand NAND4 (N6105, N6091, N5165, N4680, N4147);
nand NAND3 (N6106, N6099, N2267, N3034);
nor NOR3 (N6107, N6102, N4706, N2176);
xor XOR2 (N6108, N6106, N4511);
buf BUF1 (N6109, N6089);
xor XOR2 (N6110, N6095, N5448);
xor XOR2 (N6111, N6108, N2466);
and AND3 (N6112, N6110, N2080, N5062);
buf BUF1 (N6113, N6107);
buf BUF1 (N6114, N6103);
xor XOR2 (N6115, N6114, N1759);
xor XOR2 (N6116, N6115, N1760);
or OR3 (N6117, N6081, N138, N1508);
xor XOR2 (N6118, N6112, N5505);
buf BUF1 (N6119, N6118);
nor NOR2 (N6120, N6105, N3414);
buf BUF1 (N6121, N6104);
xor XOR2 (N6122, N6116, N1713);
nand NAND2 (N6123, N6119, N2249);
nor NOR2 (N6124, N6121, N2581);
buf BUF1 (N6125, N6111);
nor NOR4 (N6126, N6086, N3862, N5261, N3892);
not NOT1 (N6127, N6097);
nand NAND4 (N6128, N6123, N4742, N2792, N5310);
buf BUF1 (N6129, N6128);
xor XOR2 (N6130, N6129, N1290);
or OR3 (N6131, N6120, N902, N578);
buf BUF1 (N6132, N6109);
nor NOR3 (N6133, N6124, N5837, N4905);
buf BUF1 (N6134, N6125);
not NOT1 (N6135, N6122);
not NOT1 (N6136, N6135);
xor XOR2 (N6137, N6130, N4222);
nor NOR3 (N6138, N6133, N638, N5336);
nand NAND3 (N6139, N6127, N2703, N940);
and AND2 (N6140, N6117, N4319);
buf BUF1 (N6141, N6132);
or OR4 (N6142, N6126, N976, N3947, N3280);
or OR3 (N6143, N6140, N4556, N5853);
buf BUF1 (N6144, N6141);
nor NOR4 (N6145, N6144, N1395, N5197, N4125);
and AND2 (N6146, N6134, N2312);
nor NOR2 (N6147, N6137, N4975);
buf BUF1 (N6148, N6136);
buf BUF1 (N6149, N6145);
nor NOR2 (N6150, N6146, N4302);
and AND2 (N6151, N6131, N5425);
and AND4 (N6152, N6139, N5409, N4086, N178);
not NOT1 (N6153, N6113);
not NOT1 (N6154, N6148);
buf BUF1 (N6155, N6143);
buf BUF1 (N6156, N6147);
nand NAND3 (N6157, N6149, N4447, N3820);
nor NOR2 (N6158, N6155, N474);
xor XOR2 (N6159, N6142, N3871);
buf BUF1 (N6160, N6138);
buf BUF1 (N6161, N6153);
or OR4 (N6162, N6154, N2919, N66, N3516);
and AND3 (N6163, N6162, N3948, N2380);
xor XOR2 (N6164, N6157, N2902);
xor XOR2 (N6165, N6151, N1604);
not NOT1 (N6166, N6159);
nor NOR4 (N6167, N6160, N2160, N4659, N4103);
nor NOR4 (N6168, N6164, N4771, N1970, N2778);
xor XOR2 (N6169, N6161, N2455);
buf BUF1 (N6170, N6163);
xor XOR2 (N6171, N6165, N494);
nand NAND2 (N6172, N6166, N2507);
and AND2 (N6173, N6150, N2115);
or OR3 (N6174, N6152, N4248, N935);
buf BUF1 (N6175, N6174);
buf BUF1 (N6176, N6156);
or OR4 (N6177, N6171, N3080, N3519, N432);
xor XOR2 (N6178, N6169, N612);
nor NOR3 (N6179, N6173, N4371, N2074);
not NOT1 (N6180, N6167);
not NOT1 (N6181, N6178);
and AND2 (N6182, N6180, N6046);
or OR4 (N6183, N6177, N3363, N1280, N4153);
and AND2 (N6184, N6182, N5451);
nor NOR2 (N6185, N6181, N5834);
xor XOR2 (N6186, N6184, N2090);
nor NOR3 (N6187, N6168, N5068, N4637);
and AND3 (N6188, N6187, N4078, N3420);
or OR3 (N6189, N6170, N6187, N2676);
and AND4 (N6190, N6188, N4108, N1891, N3148);
not NOT1 (N6191, N6158);
nor NOR2 (N6192, N6191, N2232);
not NOT1 (N6193, N6175);
xor XOR2 (N6194, N6190, N3209);
xor XOR2 (N6195, N6186, N1034);
and AND2 (N6196, N6189, N5595);
nor NOR4 (N6197, N6195, N3413, N3374, N1628);
buf BUF1 (N6198, N6179);
or OR4 (N6199, N6193, N4938, N3875, N3150);
nor NOR4 (N6200, N6185, N273, N4734, N1124);
or OR3 (N6201, N6176, N4222, N5197);
nand NAND2 (N6202, N6197, N2127);
buf BUF1 (N6203, N6198);
nor NOR3 (N6204, N6196, N2678, N1925);
nor NOR4 (N6205, N6204, N5717, N271, N1897);
buf BUF1 (N6206, N6202);
nor NOR2 (N6207, N6183, N3462);
not NOT1 (N6208, N6203);
buf BUF1 (N6209, N6172);
nand NAND3 (N6210, N6207, N5348, N100);
buf BUF1 (N6211, N6210);
buf BUF1 (N6212, N6201);
nand NAND2 (N6213, N6200, N6154);
buf BUF1 (N6214, N6206);
and AND4 (N6215, N6199, N2564, N5881, N3469);
xor XOR2 (N6216, N6205, N4757);
buf BUF1 (N6217, N6209);
or OR3 (N6218, N6213, N4679, N5271);
nor NOR2 (N6219, N6215, N351);
not NOT1 (N6220, N6192);
nor NOR3 (N6221, N6214, N486, N3354);
or OR2 (N6222, N6212, N3560);
xor XOR2 (N6223, N6216, N4579);
and AND4 (N6224, N6218, N3039, N90, N5174);
nand NAND3 (N6225, N6220, N1498, N5325);
or OR3 (N6226, N6221, N3491, N1549);
and AND4 (N6227, N6225, N15, N2201, N721);
buf BUF1 (N6228, N6208);
buf BUF1 (N6229, N6228);
and AND4 (N6230, N6194, N689, N2689, N237);
and AND3 (N6231, N6226, N3159, N5775);
buf BUF1 (N6232, N6211);
xor XOR2 (N6233, N6223, N2624);
not NOT1 (N6234, N6229);
xor XOR2 (N6235, N6227, N1813);
or OR3 (N6236, N6235, N2269, N3690);
and AND3 (N6237, N6222, N36, N519);
nand NAND2 (N6238, N6233, N1986);
and AND3 (N6239, N6232, N1915, N5112);
or OR3 (N6240, N6217, N858, N5643);
and AND4 (N6241, N6239, N2201, N1196, N1548);
nor NOR3 (N6242, N6224, N2991, N4871);
xor XOR2 (N6243, N6242, N2576);
and AND4 (N6244, N6241, N3143, N1039, N886);
nand NAND2 (N6245, N6236, N744);
nand NAND4 (N6246, N6234, N1793, N6202, N3439);
xor XOR2 (N6247, N6238, N2068);
nor NOR4 (N6248, N6230, N1165, N3770, N112);
nor NOR3 (N6249, N6243, N2807, N459);
and AND4 (N6250, N6246, N2842, N4198, N4291);
nor NOR2 (N6251, N6244, N3124);
or OR4 (N6252, N6248, N3784, N5248, N3643);
and AND3 (N6253, N6219, N2444, N5999);
xor XOR2 (N6254, N6251, N5076);
nand NAND4 (N6255, N6247, N1500, N5547, N1114);
and AND2 (N6256, N6253, N5607);
nand NAND4 (N6257, N6250, N1545, N882, N215);
xor XOR2 (N6258, N6255, N2487);
nor NOR3 (N6259, N6254, N560, N2977);
not NOT1 (N6260, N6252);
xor XOR2 (N6261, N6259, N3925);
xor XOR2 (N6262, N6260, N857);
xor XOR2 (N6263, N6261, N2603);
or OR2 (N6264, N6256, N3497);
nand NAND4 (N6265, N6249, N3519, N3738, N1981);
xor XOR2 (N6266, N6264, N1376);
nor NOR4 (N6267, N6265, N3698, N6235, N2868);
nor NOR3 (N6268, N6267, N4018, N2687);
and AND2 (N6269, N6262, N1406);
and AND3 (N6270, N6237, N1555, N4935);
buf BUF1 (N6271, N6268);
not NOT1 (N6272, N6266);
or OR4 (N6273, N6257, N6088, N5533, N2432);
buf BUF1 (N6274, N6273);
and AND4 (N6275, N6274, N4579, N971, N5539);
or OR4 (N6276, N6269, N1290, N299, N2900);
nand NAND2 (N6277, N6245, N1423);
nor NOR2 (N6278, N6231, N5014);
and AND2 (N6279, N6270, N1094);
not NOT1 (N6280, N6275);
nand NAND3 (N6281, N6280, N5447, N1592);
not NOT1 (N6282, N6258);
nor NOR4 (N6283, N6271, N3645, N3035, N1248);
or OR2 (N6284, N6240, N2772);
not NOT1 (N6285, N6279);
nor NOR3 (N6286, N6282, N1896, N3713);
buf BUF1 (N6287, N6276);
not NOT1 (N6288, N6284);
and AND3 (N6289, N6277, N5245, N3764);
and AND3 (N6290, N6289, N872, N5436);
xor XOR2 (N6291, N6281, N208);
not NOT1 (N6292, N6278);
not NOT1 (N6293, N6285);
nand NAND4 (N6294, N6288, N3740, N989, N393);
nor NOR4 (N6295, N6283, N1173, N681, N296);
buf BUF1 (N6296, N6263);
buf BUF1 (N6297, N6295);
xor XOR2 (N6298, N6286, N465);
buf BUF1 (N6299, N6294);
not NOT1 (N6300, N6299);
xor XOR2 (N6301, N6272, N5681);
or OR4 (N6302, N6291, N3928, N4408, N4662);
not NOT1 (N6303, N6290);
nand NAND3 (N6304, N6302, N1667, N2019);
not NOT1 (N6305, N6292);
xor XOR2 (N6306, N6296, N3922);
not NOT1 (N6307, N6306);
nor NOR4 (N6308, N6298, N1558, N4206, N3701);
buf BUF1 (N6309, N6307);
xor XOR2 (N6310, N6287, N2506);
or OR3 (N6311, N6303, N5075, N976);
nor NOR4 (N6312, N6304, N5126, N3204, N1047);
and AND3 (N6313, N6293, N5345, N3875);
xor XOR2 (N6314, N6313, N2723);
and AND3 (N6315, N6308, N3385, N3001);
nand NAND2 (N6316, N6311, N108);
not NOT1 (N6317, N6301);
xor XOR2 (N6318, N6300, N304);
nand NAND4 (N6319, N6317, N1009, N1956, N6009);
or OR2 (N6320, N6319, N6130);
or OR2 (N6321, N6312, N5346);
xor XOR2 (N6322, N6321, N4876);
not NOT1 (N6323, N6320);
nor NOR2 (N6324, N6297, N5232);
nand NAND3 (N6325, N6309, N737, N5907);
buf BUF1 (N6326, N6314);
nor NOR4 (N6327, N6310, N4530, N723, N6046);
xor XOR2 (N6328, N6325, N518);
buf BUF1 (N6329, N6327);
xor XOR2 (N6330, N6324, N5731);
or OR2 (N6331, N6318, N5595);
nand NAND2 (N6332, N6305, N6110);
buf BUF1 (N6333, N6322);
nor NOR3 (N6334, N6323, N3472, N451);
and AND3 (N6335, N6326, N833, N5808);
or OR4 (N6336, N6335, N1929, N6091, N3718);
xor XOR2 (N6337, N6334, N4665);
xor XOR2 (N6338, N6330, N4466);
xor XOR2 (N6339, N6328, N1257);
not NOT1 (N6340, N6332);
nor NOR3 (N6341, N6331, N5730, N104);
nand NAND4 (N6342, N6329, N5758, N376, N4563);
or OR4 (N6343, N6341, N1725, N4597, N1067);
and AND3 (N6344, N6338, N2489, N435);
xor XOR2 (N6345, N6343, N1597);
nor NOR3 (N6346, N6316, N1496, N4004);
not NOT1 (N6347, N6336);
nor NOR4 (N6348, N6315, N3786, N2494, N506);
nor NOR3 (N6349, N6339, N4205, N1150);
and AND2 (N6350, N6347, N5391);
not NOT1 (N6351, N6337);
xor XOR2 (N6352, N6340, N4649);
nand NAND4 (N6353, N6344, N5507, N6196, N3621);
and AND2 (N6354, N6345, N4896);
nor NOR4 (N6355, N6346, N3988, N2773, N1217);
buf BUF1 (N6356, N6352);
or OR2 (N6357, N6354, N170);
or OR3 (N6358, N6342, N1401, N2752);
and AND2 (N6359, N6355, N3674);
or OR2 (N6360, N6333, N510);
buf BUF1 (N6361, N6356);
nand NAND4 (N6362, N6348, N5712, N6285, N3022);
xor XOR2 (N6363, N6351, N3767);
or OR3 (N6364, N6362, N4079, N772);
not NOT1 (N6365, N6358);
buf BUF1 (N6366, N6353);
or OR3 (N6367, N6366, N4290, N4449);
xor XOR2 (N6368, N6364, N587);
xor XOR2 (N6369, N6367, N4845);
not NOT1 (N6370, N6359);
xor XOR2 (N6371, N6360, N4951);
not NOT1 (N6372, N6363);
or OR4 (N6373, N6371, N2293, N4200, N2728);
not NOT1 (N6374, N6369);
nor NOR3 (N6375, N6370, N5310, N1684);
nor NOR3 (N6376, N6368, N702, N4293);
buf BUF1 (N6377, N6373);
or OR4 (N6378, N6349, N6316, N1940, N4776);
and AND4 (N6379, N6378, N5474, N2241, N5227);
and AND2 (N6380, N6357, N1057);
not NOT1 (N6381, N6374);
buf BUF1 (N6382, N6376);
and AND4 (N6383, N6350, N2762, N3819, N4605);
or OR2 (N6384, N6382, N3241);
nand NAND3 (N6385, N6377, N1721, N3766);
and AND3 (N6386, N6384, N2535, N905);
or OR2 (N6387, N6379, N5949);
not NOT1 (N6388, N6383);
and AND3 (N6389, N6365, N798, N5445);
nor NOR4 (N6390, N6385, N690, N246, N4750);
xor XOR2 (N6391, N6375, N901);
nand NAND4 (N6392, N6372, N2924, N5578, N3887);
xor XOR2 (N6393, N6361, N2118);
or OR3 (N6394, N6387, N723, N6030);
or OR4 (N6395, N6392, N652, N440, N6071);
buf BUF1 (N6396, N6389);
nand NAND2 (N6397, N6386, N1039);
or OR4 (N6398, N6395, N4252, N4039, N5191);
buf BUF1 (N6399, N6393);
or OR2 (N6400, N6388, N2749);
buf BUF1 (N6401, N6390);
buf BUF1 (N6402, N6380);
and AND4 (N6403, N6400, N2201, N3537, N6231);
nor NOR3 (N6404, N6394, N739, N6356);
nand NAND3 (N6405, N6398, N3217, N4639);
or OR2 (N6406, N6401, N359);
or OR4 (N6407, N6396, N3366, N4194, N2300);
xor XOR2 (N6408, N6402, N5773);
nand NAND4 (N6409, N6407, N120, N1332, N4169);
and AND3 (N6410, N6403, N1685, N4542);
xor XOR2 (N6411, N6408, N4194);
not NOT1 (N6412, N6405);
nand NAND3 (N6413, N6391, N5088, N1142);
and AND4 (N6414, N6410, N468, N5155, N2413);
and AND3 (N6415, N6409, N5622, N2986);
and AND4 (N6416, N6381, N4473, N1524, N1210);
buf BUF1 (N6417, N6404);
or OR3 (N6418, N6397, N4793, N1725);
endmodule