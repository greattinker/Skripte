// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N811,N814,N820,N818,N809,N812,N822,N806,N821,N823;

nor NOR3 (N24, N2, N11, N9);
xor XOR2 (N25, N18, N10);
buf BUF1 (N26, N24);
or OR4 (N27, N25, N15, N11, N13);
buf BUF1 (N28, N27);
not NOT1 (N29, N22);
and AND3 (N30, N23, N27, N25);
buf BUF1 (N31, N1);
buf BUF1 (N32, N19);
nand NAND4 (N33, N4, N27, N29, N17);
nor NOR2 (N34, N23, N12);
and AND3 (N35, N15, N20, N12);
nor NOR2 (N36, N16, N6);
not NOT1 (N37, N26);
or OR4 (N38, N19, N30, N16, N35);
not NOT1 (N39, N35);
not NOT1 (N40, N12);
or OR3 (N41, N38, N13, N12);
or OR3 (N42, N28, N40, N32);
xor XOR2 (N43, N14, N34);
buf BUF1 (N44, N28);
buf BUF1 (N45, N40);
nor NOR2 (N46, N42, N45);
nand NAND2 (N47, N16, N8);
buf BUF1 (N48, N31);
nor NOR2 (N49, N44, N14);
xor XOR2 (N50, N46, N7);
not NOT1 (N51, N37);
nand NAND2 (N52, N47, N41);
and AND2 (N53, N43, N48);
or OR2 (N54, N23, N49);
xor XOR2 (N55, N51, N37);
xor XOR2 (N56, N35, N51);
or OR2 (N57, N13, N20);
or OR2 (N58, N54, N47);
or OR2 (N59, N56, N29);
buf BUF1 (N60, N36);
or OR4 (N61, N53, N2, N60, N4);
nor NOR4 (N62, N61, N58, N8, N18);
or OR4 (N63, N12, N25, N5, N32);
xor XOR2 (N64, N61, N22);
and AND2 (N65, N50, N27);
nand NAND3 (N66, N59, N20, N47);
and AND3 (N67, N62, N58, N66);
or OR4 (N68, N35, N36, N50, N21);
buf BUF1 (N69, N63);
nand NAND3 (N70, N65, N22, N25);
buf BUF1 (N71, N52);
xor XOR2 (N72, N71, N54);
xor XOR2 (N73, N67, N14);
and AND3 (N74, N64, N18, N4);
or OR4 (N75, N73, N22, N43, N22);
xor XOR2 (N76, N68, N53);
not NOT1 (N77, N74);
not NOT1 (N78, N70);
xor XOR2 (N79, N78, N4);
nor NOR2 (N80, N76, N65);
and AND3 (N81, N80, N55, N46);
not NOT1 (N82, N5);
and AND2 (N83, N79, N13);
or OR2 (N84, N82, N65);
or OR2 (N85, N84, N20);
buf BUF1 (N86, N85);
and AND2 (N87, N81, N57);
buf BUF1 (N88, N11);
nand NAND3 (N89, N88, N85, N24);
nand NAND3 (N90, N83, N2, N73);
nor NOR2 (N91, N75, N78);
not NOT1 (N92, N87);
or OR3 (N93, N39, N6, N70);
or OR3 (N94, N72, N26, N81);
nor NOR3 (N95, N90, N19, N22);
nor NOR3 (N96, N91, N76, N90);
and AND4 (N97, N93, N65, N94, N28);
nor NOR3 (N98, N23, N29, N92);
nand NAND2 (N99, N91, N26);
nand NAND2 (N100, N96, N87);
and AND4 (N101, N97, N66, N81, N85);
nor NOR4 (N102, N33, N26, N88, N61);
and AND2 (N103, N99, N26);
xor XOR2 (N104, N101, N28);
or OR4 (N105, N69, N63, N16, N62);
and AND3 (N106, N104, N57, N98);
nor NOR4 (N107, N9, N70, N92, N64);
nor NOR4 (N108, N100, N99, N21, N63);
and AND3 (N109, N89, N3, N78);
buf BUF1 (N110, N105);
nand NAND4 (N111, N86, N46, N28, N3);
nor NOR4 (N112, N77, N50, N87, N18);
or OR2 (N113, N103, N58);
nor NOR3 (N114, N110, N102, N6);
xor XOR2 (N115, N50, N88);
nand NAND4 (N116, N111, N32, N63, N106);
not NOT1 (N117, N56);
nand NAND2 (N118, N115, N76);
xor XOR2 (N119, N112, N39);
buf BUF1 (N120, N118);
not NOT1 (N121, N116);
xor XOR2 (N122, N109, N96);
buf BUF1 (N123, N120);
nand NAND3 (N124, N113, N99, N123);
nor NOR2 (N125, N112, N97);
and AND2 (N126, N108, N17);
nand NAND2 (N127, N126, N4);
not NOT1 (N128, N114);
buf BUF1 (N129, N95);
xor XOR2 (N130, N124, N18);
buf BUF1 (N131, N107);
nand NAND4 (N132, N119, N25, N125, N126);
xor XOR2 (N133, N69, N130);
and AND4 (N134, N100, N92, N19, N106);
nor NOR2 (N135, N117, N7);
xor XOR2 (N136, N132, N113);
xor XOR2 (N137, N129, N52);
nand NAND2 (N138, N131, N94);
and AND2 (N139, N121, N43);
xor XOR2 (N140, N136, N53);
buf BUF1 (N141, N128);
buf BUF1 (N142, N140);
and AND4 (N143, N122, N121, N5, N100);
xor XOR2 (N144, N138, N18);
nor NOR3 (N145, N143, N89, N137);
not NOT1 (N146, N21);
nand NAND4 (N147, N141, N129, N17, N116);
nor NOR2 (N148, N145, N129);
and AND2 (N149, N144, N133);
nor NOR2 (N150, N95, N131);
buf BUF1 (N151, N146);
nand NAND3 (N152, N127, N90, N141);
buf BUF1 (N153, N134);
not NOT1 (N154, N153);
not NOT1 (N155, N139);
xor XOR2 (N156, N148, N106);
or OR3 (N157, N150, N61, N5);
and AND2 (N158, N149, N37);
nand NAND2 (N159, N157, N16);
buf BUF1 (N160, N152);
nand NAND2 (N161, N154, N144);
nor NOR3 (N162, N142, N158, N130);
xor XOR2 (N163, N41, N33);
and AND3 (N164, N161, N64, N125);
not NOT1 (N165, N147);
not NOT1 (N166, N135);
and AND3 (N167, N163, N73, N80);
not NOT1 (N168, N155);
nor NOR3 (N169, N156, N54, N133);
and AND2 (N170, N167, N128);
and AND4 (N171, N159, N17, N36, N79);
nor NOR2 (N172, N162, N161);
and AND3 (N173, N165, N122, N35);
and AND2 (N174, N172, N6);
or OR2 (N175, N173, N73);
xor XOR2 (N176, N175, N6);
xor XOR2 (N177, N151, N152);
xor XOR2 (N178, N169, N71);
and AND2 (N179, N160, N19);
nor NOR2 (N180, N171, N47);
nand NAND4 (N181, N166, N108, N100, N4);
or OR2 (N182, N178, N22);
xor XOR2 (N183, N182, N58);
buf BUF1 (N184, N180);
xor XOR2 (N185, N164, N47);
not NOT1 (N186, N168);
nand NAND2 (N187, N176, N98);
buf BUF1 (N188, N186);
not NOT1 (N189, N170);
xor XOR2 (N190, N181, N99);
nor NOR3 (N191, N189, N11, N127);
buf BUF1 (N192, N188);
or OR3 (N193, N187, N86, N141);
nor NOR4 (N194, N190, N144, N138, N77);
and AND4 (N195, N192, N35, N139, N157);
buf BUF1 (N196, N177);
xor XOR2 (N197, N195, N66);
nand NAND4 (N198, N196, N175, N19, N71);
and AND3 (N199, N194, N72, N123);
nand NAND2 (N200, N174, N138);
not NOT1 (N201, N184);
buf BUF1 (N202, N199);
not NOT1 (N203, N185);
or OR2 (N204, N179, N159);
nor NOR2 (N205, N193, N123);
nand NAND3 (N206, N205, N16, N66);
xor XOR2 (N207, N201, N206);
buf BUF1 (N208, N128);
nand NAND4 (N209, N200, N84, N145, N173);
not NOT1 (N210, N203);
xor XOR2 (N211, N191, N11);
or OR3 (N212, N210, N173, N9);
and AND4 (N213, N204, N9, N108, N203);
buf BUF1 (N214, N183);
xor XOR2 (N215, N197, N38);
or OR3 (N216, N209, N92, N12);
and AND4 (N217, N208, N119, N141, N54);
or OR2 (N218, N217, N53);
nor NOR3 (N219, N212, N174, N116);
and AND4 (N220, N219, N64, N43, N56);
not NOT1 (N221, N214);
and AND4 (N222, N211, N130, N59, N80);
xor XOR2 (N223, N218, N110);
xor XOR2 (N224, N198, N54);
nor NOR3 (N225, N220, N58, N200);
or OR4 (N226, N215, N85, N150, N222);
buf BUF1 (N227, N167);
not NOT1 (N228, N221);
nand NAND3 (N229, N227, N160, N73);
nor NOR2 (N230, N223, N174);
xor XOR2 (N231, N228, N41);
or OR4 (N232, N231, N127, N189, N185);
not NOT1 (N233, N229);
not NOT1 (N234, N230);
or OR4 (N235, N213, N102, N2, N115);
nand NAND3 (N236, N232, N130, N120);
buf BUF1 (N237, N225);
nor NOR3 (N238, N216, N113, N171);
and AND2 (N239, N226, N188);
not NOT1 (N240, N237);
nor NOR2 (N241, N207, N8);
and AND3 (N242, N234, N77, N96);
xor XOR2 (N243, N240, N92);
xor XOR2 (N244, N239, N218);
or OR3 (N245, N202, N91, N86);
nand NAND2 (N246, N243, N76);
nand NAND2 (N247, N241, N207);
nor NOR3 (N248, N242, N11, N49);
nor NOR3 (N249, N246, N68, N40);
xor XOR2 (N250, N248, N136);
and AND3 (N251, N238, N221, N126);
or OR4 (N252, N247, N14, N201, N171);
and AND3 (N253, N250, N86, N136);
and AND4 (N254, N233, N121, N79, N180);
and AND3 (N255, N245, N116, N135);
not NOT1 (N256, N244);
buf BUF1 (N257, N251);
nand NAND4 (N258, N255, N199, N23, N226);
not NOT1 (N259, N252);
or OR4 (N260, N259, N41, N181, N150);
not NOT1 (N261, N249);
and AND3 (N262, N224, N64, N257);
xor XOR2 (N263, N128, N123);
buf BUF1 (N264, N254);
or OR3 (N265, N261, N233, N23);
or OR2 (N266, N265, N202);
or OR3 (N267, N266, N8, N197);
and AND2 (N268, N264, N111);
and AND2 (N269, N258, N49);
nor NOR3 (N270, N235, N37, N128);
and AND3 (N271, N262, N105, N141);
or OR3 (N272, N236, N134, N225);
buf BUF1 (N273, N272);
and AND3 (N274, N269, N272, N34);
nor NOR3 (N275, N268, N47, N197);
and AND2 (N276, N267, N148);
buf BUF1 (N277, N260);
not NOT1 (N278, N263);
xor XOR2 (N279, N256, N140);
buf BUF1 (N280, N276);
nor NOR3 (N281, N280, N152, N100);
not NOT1 (N282, N253);
and AND3 (N283, N274, N282, N257);
buf BUF1 (N284, N185);
and AND3 (N285, N271, N6, N121);
nand NAND4 (N286, N281, N48, N70, N264);
not NOT1 (N287, N270);
or OR3 (N288, N278, N189, N94);
and AND4 (N289, N285, N19, N97, N215);
not NOT1 (N290, N275);
buf BUF1 (N291, N279);
nor NOR4 (N292, N283, N124, N186, N142);
nand NAND4 (N293, N290, N55, N172, N224);
buf BUF1 (N294, N277);
xor XOR2 (N295, N273, N262);
nor NOR2 (N296, N289, N87);
buf BUF1 (N297, N294);
xor XOR2 (N298, N295, N297);
xor XOR2 (N299, N256, N188);
and AND3 (N300, N287, N214, N253);
nor NOR2 (N301, N299, N170);
or OR3 (N302, N298, N139, N217);
buf BUF1 (N303, N301);
not NOT1 (N304, N291);
xor XOR2 (N305, N296, N274);
nand NAND4 (N306, N304, N295, N201, N189);
xor XOR2 (N307, N300, N68);
not NOT1 (N308, N286);
and AND2 (N309, N288, N179);
buf BUF1 (N310, N306);
buf BUF1 (N311, N293);
nor NOR4 (N312, N302, N89, N47, N301);
and AND4 (N313, N311, N209, N259, N232);
nand NAND3 (N314, N284, N249, N308);
buf BUF1 (N315, N210);
nor NOR4 (N316, N310, N168, N241, N296);
nor NOR4 (N317, N303, N234, N64, N159);
and AND2 (N318, N292, N74);
xor XOR2 (N319, N305, N200);
nor NOR3 (N320, N312, N55, N256);
xor XOR2 (N321, N315, N84);
or OR4 (N322, N314, N276, N305, N281);
or OR2 (N323, N317, N160);
nand NAND2 (N324, N316, N52);
xor XOR2 (N325, N320, N33);
or OR2 (N326, N321, N305);
not NOT1 (N327, N319);
nand NAND4 (N328, N324, N193, N40, N230);
buf BUF1 (N329, N307);
nor NOR3 (N330, N329, N49, N292);
nor NOR2 (N331, N318, N311);
and AND4 (N332, N323, N78, N142, N323);
buf BUF1 (N333, N332);
nand NAND2 (N334, N326, N110);
not NOT1 (N335, N309);
nand NAND4 (N336, N333, N6, N317, N125);
nor NOR3 (N337, N328, N216, N196);
and AND2 (N338, N337, N224);
nor NOR2 (N339, N338, N4);
not NOT1 (N340, N313);
or OR4 (N341, N339, N156, N215, N108);
xor XOR2 (N342, N330, N213);
and AND2 (N343, N322, N2);
and AND2 (N344, N340, N306);
or OR2 (N345, N336, N253);
nor NOR2 (N346, N344, N302);
xor XOR2 (N347, N343, N240);
nor NOR4 (N348, N346, N65, N289, N300);
nor NOR2 (N349, N347, N53);
xor XOR2 (N350, N331, N179);
buf BUF1 (N351, N334);
buf BUF1 (N352, N335);
nand NAND3 (N353, N342, N157, N159);
not NOT1 (N354, N349);
xor XOR2 (N355, N353, N260);
not NOT1 (N356, N354);
nand NAND3 (N357, N356, N164, N165);
buf BUF1 (N358, N355);
and AND4 (N359, N327, N35, N169, N142);
nor NOR4 (N360, N351, N71, N323, N31);
xor XOR2 (N361, N352, N347);
buf BUF1 (N362, N341);
not NOT1 (N363, N345);
nand NAND2 (N364, N360, N261);
buf BUF1 (N365, N363);
nor NOR4 (N366, N325, N308, N138, N353);
nand NAND4 (N367, N362, N152, N279, N249);
or OR4 (N368, N357, N82, N223, N263);
buf BUF1 (N369, N350);
or OR2 (N370, N359, N109);
and AND3 (N371, N370, N331, N258);
nand NAND4 (N372, N348, N367, N140, N340);
xor XOR2 (N373, N230, N156);
buf BUF1 (N374, N366);
not NOT1 (N375, N372);
xor XOR2 (N376, N361, N127);
buf BUF1 (N377, N369);
buf BUF1 (N378, N377);
buf BUF1 (N379, N373);
or OR4 (N380, N368, N57, N319, N94);
not NOT1 (N381, N374);
buf BUF1 (N382, N364);
and AND4 (N383, N375, N23, N223, N22);
not NOT1 (N384, N379);
buf BUF1 (N385, N380);
buf BUF1 (N386, N378);
or OR4 (N387, N381, N129, N20, N107);
buf BUF1 (N388, N365);
nand NAND2 (N389, N376, N74);
xor XOR2 (N390, N389, N353);
not NOT1 (N391, N388);
nand NAND4 (N392, N386, N46, N156, N129);
nor NOR3 (N393, N391, N261, N132);
buf BUF1 (N394, N382);
xor XOR2 (N395, N387, N339);
and AND4 (N396, N392, N120, N221, N107);
not NOT1 (N397, N394);
buf BUF1 (N398, N397);
and AND4 (N399, N371, N243, N340, N32);
nor NOR4 (N400, N396, N50, N339, N219);
and AND2 (N401, N399, N297);
buf BUF1 (N402, N400);
buf BUF1 (N403, N390);
buf BUF1 (N404, N383);
buf BUF1 (N405, N404);
buf BUF1 (N406, N384);
nand NAND4 (N407, N395, N123, N199, N205);
or OR4 (N408, N385, N404, N319, N74);
nand NAND2 (N409, N408, N329);
not NOT1 (N410, N398);
xor XOR2 (N411, N407, N25);
buf BUF1 (N412, N405);
nor NOR2 (N413, N358, N145);
nor NOR3 (N414, N412, N40, N125);
and AND2 (N415, N403, N362);
not NOT1 (N416, N406);
nand NAND3 (N417, N409, N406, N186);
nor NOR3 (N418, N415, N167, N80);
nand NAND2 (N419, N417, N117);
or OR3 (N420, N414, N51, N240);
and AND3 (N421, N402, N375, N196);
and AND4 (N422, N401, N34, N191, N321);
nor NOR2 (N423, N422, N87);
buf BUF1 (N424, N420);
and AND3 (N425, N411, N132, N273);
buf BUF1 (N426, N421);
and AND3 (N427, N426, N184, N300);
xor XOR2 (N428, N423, N238);
xor XOR2 (N429, N428, N99);
xor XOR2 (N430, N424, N425);
buf BUF1 (N431, N278);
or OR3 (N432, N413, N118, N180);
buf BUF1 (N433, N416);
or OR4 (N434, N410, N98, N210, N258);
buf BUF1 (N435, N431);
xor XOR2 (N436, N418, N112);
or OR2 (N437, N429, N159);
not NOT1 (N438, N435);
buf BUF1 (N439, N437);
buf BUF1 (N440, N419);
xor XOR2 (N441, N439, N78);
buf BUF1 (N442, N441);
buf BUF1 (N443, N430);
or OR4 (N444, N436, N348, N416, N367);
xor XOR2 (N445, N393, N15);
nor NOR3 (N446, N434, N278, N338);
nor NOR3 (N447, N442, N444, N52);
buf BUF1 (N448, N284);
buf BUF1 (N449, N446);
nand NAND3 (N450, N427, N154, N389);
or OR4 (N451, N445, N142, N323, N371);
and AND3 (N452, N448, N248, N208);
not NOT1 (N453, N451);
xor XOR2 (N454, N452, N194);
or OR2 (N455, N443, N125);
or OR3 (N456, N447, N186, N154);
nor NOR3 (N457, N433, N190, N413);
and AND2 (N458, N450, N170);
xor XOR2 (N459, N457, N191);
buf BUF1 (N460, N453);
or OR3 (N461, N440, N413, N454);
not NOT1 (N462, N132);
xor XOR2 (N463, N461, N430);
nand NAND2 (N464, N456, N272);
and AND3 (N465, N432, N295, N81);
buf BUF1 (N466, N459);
xor XOR2 (N467, N462, N96);
or OR4 (N468, N464, N66, N369, N125);
buf BUF1 (N469, N449);
not NOT1 (N470, N466);
or OR3 (N471, N455, N372, N437);
nor NOR2 (N472, N438, N190);
xor XOR2 (N473, N468, N123);
nor NOR4 (N474, N470, N114, N36, N390);
and AND3 (N475, N473, N452, N151);
and AND2 (N476, N460, N327);
or OR3 (N477, N465, N72, N183);
and AND2 (N478, N469, N257);
and AND4 (N479, N458, N87, N125, N447);
xor XOR2 (N480, N478, N444);
not NOT1 (N481, N471);
nand NAND3 (N482, N477, N59, N419);
nor NOR4 (N483, N479, N266, N155, N455);
xor XOR2 (N484, N476, N418);
not NOT1 (N485, N481);
buf BUF1 (N486, N467);
and AND4 (N487, N482, N14, N403, N486);
nor NOR4 (N488, N431, N347, N104, N279);
not NOT1 (N489, N488);
nor NOR2 (N490, N484, N463);
nand NAND3 (N491, N358, N70, N224);
xor XOR2 (N492, N475, N61);
and AND2 (N493, N491, N279);
nor NOR2 (N494, N493, N378);
and AND2 (N495, N492, N342);
nand NAND2 (N496, N474, N452);
not NOT1 (N497, N495);
and AND3 (N498, N490, N216, N217);
and AND4 (N499, N489, N95, N268, N405);
nor NOR3 (N500, N497, N401, N260);
and AND3 (N501, N500, N115, N194);
buf BUF1 (N502, N480);
nand NAND2 (N503, N485, N467);
buf BUF1 (N504, N498);
and AND2 (N505, N503, N3);
nor NOR4 (N506, N499, N230, N449, N38);
or OR3 (N507, N496, N441, N382);
or OR4 (N508, N504, N212, N64, N249);
nor NOR3 (N509, N502, N85, N316);
nor NOR3 (N510, N505, N324, N76);
buf BUF1 (N511, N508);
and AND2 (N512, N509, N173);
or OR2 (N513, N510, N274);
buf BUF1 (N514, N501);
buf BUF1 (N515, N472);
nor NOR4 (N516, N513, N419, N104, N387);
xor XOR2 (N517, N506, N84);
nor NOR3 (N518, N512, N11, N362);
and AND2 (N519, N483, N32);
xor XOR2 (N520, N514, N136);
xor XOR2 (N521, N515, N240);
xor XOR2 (N522, N521, N108);
not NOT1 (N523, N517);
nor NOR4 (N524, N487, N124, N225, N31);
xor XOR2 (N525, N511, N494);
xor XOR2 (N526, N319, N127);
and AND2 (N527, N526, N89);
buf BUF1 (N528, N527);
xor XOR2 (N529, N523, N402);
not NOT1 (N530, N516);
buf BUF1 (N531, N518);
nor NOR4 (N532, N524, N299, N338, N471);
buf BUF1 (N533, N520);
buf BUF1 (N534, N529);
not NOT1 (N535, N531);
xor XOR2 (N536, N534, N306);
and AND2 (N537, N535, N154);
not NOT1 (N538, N533);
xor XOR2 (N539, N507, N160);
and AND4 (N540, N536, N172, N228, N120);
or OR2 (N541, N540, N516);
and AND2 (N542, N541, N109);
nor NOR2 (N543, N525, N524);
xor XOR2 (N544, N539, N150);
nor NOR3 (N545, N544, N94, N308);
nor NOR4 (N546, N532, N369, N130, N237);
nand NAND3 (N547, N528, N365, N230);
xor XOR2 (N548, N538, N268);
nor NOR2 (N549, N530, N85);
not NOT1 (N550, N543);
or OR4 (N551, N547, N494, N471, N49);
nor NOR2 (N552, N522, N426);
and AND3 (N553, N545, N485, N235);
buf BUF1 (N554, N519);
and AND3 (N555, N552, N334, N550);
nor NOR2 (N556, N493, N353);
not NOT1 (N557, N556);
or OR3 (N558, N553, N557, N417);
or OR4 (N559, N303, N22, N237, N211);
nor NOR2 (N560, N551, N193);
not NOT1 (N561, N537);
and AND2 (N562, N555, N323);
not NOT1 (N563, N558);
nor NOR4 (N564, N546, N332, N435, N507);
nor NOR3 (N565, N542, N393, N561);
or OR2 (N566, N457, N224);
and AND4 (N567, N565, N360, N413, N460);
nor NOR4 (N568, N548, N68, N111, N136);
xor XOR2 (N569, N549, N317);
buf BUF1 (N570, N567);
not NOT1 (N571, N570);
nor NOR4 (N572, N564, N281, N145, N478);
and AND3 (N573, N566, N336, N408);
nor NOR2 (N574, N572, N37);
not NOT1 (N575, N569);
nor NOR4 (N576, N563, N158, N340, N160);
xor XOR2 (N577, N574, N487);
buf BUF1 (N578, N575);
xor XOR2 (N579, N560, N339);
nand NAND2 (N580, N577, N446);
buf BUF1 (N581, N571);
not NOT1 (N582, N573);
not NOT1 (N583, N582);
or OR2 (N584, N578, N86);
and AND2 (N585, N576, N14);
and AND3 (N586, N585, N447, N427);
nor NOR2 (N587, N568, N97);
nor NOR2 (N588, N559, N314);
not NOT1 (N589, N584);
nand NAND2 (N590, N588, N38);
or OR2 (N591, N583, N491);
or OR4 (N592, N580, N391, N140, N483);
nor NOR3 (N593, N586, N501, N478);
not NOT1 (N594, N562);
nor NOR4 (N595, N581, N299, N44, N77);
nor NOR4 (N596, N591, N424, N267, N439);
xor XOR2 (N597, N595, N530);
not NOT1 (N598, N594);
buf BUF1 (N599, N596);
xor XOR2 (N600, N554, N476);
buf BUF1 (N601, N587);
xor XOR2 (N602, N597, N583);
xor XOR2 (N603, N579, N266);
or OR3 (N604, N599, N534, N233);
not NOT1 (N605, N598);
nor NOR4 (N606, N603, N159, N139, N503);
and AND2 (N607, N592, N578);
or OR4 (N608, N590, N56, N506, N478);
and AND4 (N609, N607, N16, N34, N276);
xor XOR2 (N610, N602, N313);
buf BUF1 (N611, N589);
nor NOR2 (N612, N593, N118);
or OR3 (N613, N609, N53, N417);
xor XOR2 (N614, N610, N185);
buf BUF1 (N615, N612);
and AND4 (N616, N606, N563, N419, N553);
or OR3 (N617, N601, N420, N69);
nand NAND2 (N618, N604, N548);
and AND2 (N619, N605, N479);
nand NAND3 (N620, N616, N15, N355);
and AND3 (N621, N608, N102, N361);
and AND2 (N622, N611, N163);
or OR2 (N623, N618, N105);
xor XOR2 (N624, N621, N332);
nor NOR2 (N625, N623, N396);
nand NAND3 (N626, N615, N316, N317);
not NOT1 (N627, N619);
xor XOR2 (N628, N620, N350);
nor NOR2 (N629, N625, N424);
or OR4 (N630, N628, N521, N166, N629);
or OR2 (N631, N212, N139);
and AND3 (N632, N624, N232, N341);
nand NAND2 (N633, N632, N238);
buf BUF1 (N634, N600);
not NOT1 (N635, N626);
and AND2 (N636, N634, N379);
nand NAND3 (N637, N630, N452, N207);
not NOT1 (N638, N614);
xor XOR2 (N639, N635, N53);
nand NAND3 (N640, N617, N506, N210);
xor XOR2 (N641, N622, N158);
buf BUF1 (N642, N640);
or OR4 (N643, N613, N577, N589, N82);
or OR4 (N644, N627, N24, N541, N91);
nor NOR3 (N645, N631, N306, N589);
buf BUF1 (N646, N639);
and AND2 (N647, N642, N191);
or OR4 (N648, N646, N615, N160, N91);
nor NOR2 (N649, N648, N296);
nor NOR4 (N650, N647, N110, N592, N360);
xor XOR2 (N651, N645, N615);
buf BUF1 (N652, N651);
nor NOR3 (N653, N649, N291, N292);
not NOT1 (N654, N653);
or OR4 (N655, N643, N236, N43, N335);
nor NOR2 (N656, N636, N330);
not NOT1 (N657, N652);
nor NOR2 (N658, N644, N381);
not NOT1 (N659, N657);
xor XOR2 (N660, N659, N337);
not NOT1 (N661, N660);
nor NOR3 (N662, N633, N632, N254);
not NOT1 (N663, N658);
and AND2 (N664, N655, N176);
and AND2 (N665, N637, N39);
nor NOR2 (N666, N661, N87);
not NOT1 (N667, N662);
xor XOR2 (N668, N656, N509);
or OR4 (N669, N666, N402, N148, N449);
xor XOR2 (N670, N668, N630);
xor XOR2 (N671, N654, N207);
not NOT1 (N672, N663);
nand NAND4 (N673, N664, N608, N562, N406);
nor NOR3 (N674, N669, N586, N64);
nor NOR2 (N675, N641, N274);
nand NAND4 (N676, N673, N147, N542, N383);
nand NAND2 (N677, N674, N511);
or OR3 (N678, N638, N47, N142);
buf BUF1 (N679, N665);
xor XOR2 (N680, N670, N263);
or OR2 (N681, N680, N276);
xor XOR2 (N682, N671, N350);
nand NAND3 (N683, N678, N7, N157);
nand NAND2 (N684, N679, N583);
and AND2 (N685, N672, N359);
nand NAND4 (N686, N667, N139, N46, N394);
not NOT1 (N687, N685);
or OR4 (N688, N687, N448, N452, N50);
not NOT1 (N689, N682);
nor NOR3 (N690, N677, N380, N534);
xor XOR2 (N691, N675, N290);
and AND3 (N692, N689, N214, N458);
nand NAND2 (N693, N691, N307);
not NOT1 (N694, N681);
nor NOR3 (N695, N683, N403, N659);
nand NAND3 (N696, N695, N15, N572);
or OR2 (N697, N694, N679);
buf BUF1 (N698, N686);
and AND4 (N699, N688, N216, N153, N334);
or OR4 (N700, N690, N572, N414, N484);
or OR2 (N701, N698, N207);
or OR3 (N702, N696, N431, N40);
nand NAND3 (N703, N697, N152, N557);
buf BUF1 (N704, N701);
xor XOR2 (N705, N700, N338);
nand NAND4 (N706, N676, N200, N653, N33);
or OR3 (N707, N705, N620, N400);
xor XOR2 (N708, N684, N307);
xor XOR2 (N709, N706, N466);
nand NAND3 (N710, N702, N223, N580);
xor XOR2 (N711, N707, N601);
nand NAND3 (N712, N650, N687, N50);
buf BUF1 (N713, N703);
or OR3 (N714, N692, N322, N387);
buf BUF1 (N715, N704);
xor XOR2 (N716, N693, N157);
nor NOR3 (N717, N713, N391, N274);
and AND4 (N718, N714, N642, N84, N553);
nand NAND4 (N719, N715, N604, N73, N538);
buf BUF1 (N720, N699);
xor XOR2 (N721, N708, N562);
or OR3 (N722, N718, N395, N242);
and AND4 (N723, N719, N420, N337, N149);
not NOT1 (N724, N710);
not NOT1 (N725, N724);
nand NAND3 (N726, N721, N706, N593);
nand NAND3 (N727, N711, N151, N430);
and AND2 (N728, N720, N590);
xor XOR2 (N729, N726, N686);
nand NAND3 (N730, N727, N530, N567);
or OR4 (N731, N722, N179, N146, N379);
nand NAND2 (N732, N728, N317);
and AND4 (N733, N717, N724, N100, N429);
not NOT1 (N734, N716);
or OR3 (N735, N712, N15, N319);
not NOT1 (N736, N709);
xor XOR2 (N737, N734, N242);
xor XOR2 (N738, N729, N111);
or OR2 (N739, N738, N382);
buf BUF1 (N740, N737);
nor NOR2 (N741, N730, N28);
nand NAND3 (N742, N732, N637, N284);
or OR4 (N743, N735, N24, N527, N658);
nor NOR4 (N744, N723, N741, N584, N706);
not NOT1 (N745, N617);
nor NOR4 (N746, N743, N525, N206, N361);
not NOT1 (N747, N740);
xor XOR2 (N748, N725, N192);
and AND4 (N749, N736, N363, N602, N323);
not NOT1 (N750, N739);
or OR3 (N751, N747, N538, N673);
nor NOR3 (N752, N744, N512, N144);
or OR2 (N753, N733, N208);
xor XOR2 (N754, N746, N342);
buf BUF1 (N755, N752);
and AND4 (N756, N745, N613, N347, N584);
not NOT1 (N757, N731);
or OR2 (N758, N754, N660);
nor NOR3 (N759, N748, N505, N10);
and AND4 (N760, N757, N280, N392, N590);
nand NAND4 (N761, N742, N201, N459, N207);
nor NOR2 (N762, N749, N139);
buf BUF1 (N763, N758);
nand NAND4 (N764, N750, N614, N203, N239);
nand NAND4 (N765, N763, N295, N52, N500);
or OR4 (N766, N759, N82, N1, N277);
nor NOR4 (N767, N760, N287, N109, N439);
or OR2 (N768, N753, N8);
nand NAND2 (N769, N751, N514);
not NOT1 (N770, N764);
nand NAND3 (N771, N769, N540, N367);
not NOT1 (N772, N770);
buf BUF1 (N773, N756);
not NOT1 (N774, N773);
nand NAND2 (N775, N772, N592);
xor XOR2 (N776, N775, N496);
not NOT1 (N777, N774);
xor XOR2 (N778, N766, N607);
xor XOR2 (N779, N765, N142);
nand NAND2 (N780, N779, N174);
buf BUF1 (N781, N755);
and AND4 (N782, N762, N649, N631, N147);
not NOT1 (N783, N771);
and AND3 (N784, N767, N767, N310);
or OR4 (N785, N768, N656, N693, N419);
nor NOR2 (N786, N785, N334);
nand NAND2 (N787, N780, N623);
xor XOR2 (N788, N761, N704);
buf BUF1 (N789, N778);
nand NAND4 (N790, N789, N606, N651, N482);
nor NOR2 (N791, N788, N296);
or OR3 (N792, N777, N708, N415);
nand NAND3 (N793, N783, N623, N757);
nor NOR4 (N794, N790, N637, N324, N211);
or OR3 (N795, N776, N702, N361);
or OR2 (N796, N784, N791);
not NOT1 (N797, N212);
xor XOR2 (N798, N792, N253);
or OR4 (N799, N795, N105, N793, N431);
or OR4 (N800, N605, N372, N296, N36);
xor XOR2 (N801, N787, N82);
or OR4 (N802, N798, N464, N682, N166);
or OR3 (N803, N781, N111, N506);
nand NAND2 (N804, N782, N155);
or OR3 (N805, N802, N488, N45);
nand NAND3 (N806, N800, N94, N465);
not NOT1 (N807, N797);
buf BUF1 (N808, N799);
nor NOR2 (N809, N794, N120);
and AND3 (N810, N807, N667, N543);
or OR2 (N811, N810, N296);
xor XOR2 (N812, N808, N18);
buf BUF1 (N813, N805);
buf BUF1 (N814, N803);
and AND2 (N815, N801, N654);
xor XOR2 (N816, N786, N786);
nand NAND2 (N817, N815, N147);
xor XOR2 (N818, N817, N37);
or OR3 (N819, N796, N718, N128);
nor NOR2 (N820, N804, N558);
nand NAND4 (N821, N819, N652, N813, N535);
nand NAND2 (N822, N607, N450);
nand NAND3 (N823, N816, N57, N372);
endmodule