// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N717,N708,N722,N687,N712,N720,N707,N716,N718,N724;

xor XOR2 (N25, N22, N3);
nor NOR4 (N26, N20, N11, N19, N20);
nand NAND4 (N27, N15, N13, N3, N9);
or OR4 (N28, N19, N23, N1, N11);
nand NAND2 (N29, N8, N19);
not NOT1 (N30, N4);
or OR4 (N31, N12, N12, N27, N10);
nand NAND2 (N32, N7, N18);
or OR3 (N33, N20, N16, N18);
buf BUF1 (N34, N10);
nor NOR4 (N35, N26, N30, N30, N14);
xor XOR2 (N36, N20, N1);
not NOT1 (N37, N25);
not NOT1 (N38, N8);
not NOT1 (N39, N33);
xor XOR2 (N40, N28, N20);
nand NAND4 (N41, N32, N28, N29, N14);
buf BUF1 (N42, N27);
not NOT1 (N43, N39);
nor NOR3 (N44, N40, N15, N27);
xor XOR2 (N45, N38, N14);
not NOT1 (N46, N45);
or OR4 (N47, N46, N5, N5, N10);
or OR4 (N48, N37, N8, N34, N8);
or OR2 (N49, N7, N24);
or OR4 (N50, N48, N39, N15, N39);
and AND2 (N51, N49, N17);
buf BUF1 (N52, N50);
nand NAND2 (N53, N41, N40);
buf BUF1 (N54, N51);
buf BUF1 (N55, N43);
and AND3 (N56, N31, N28, N7);
nand NAND2 (N57, N36, N2);
or OR2 (N58, N54, N6);
or OR4 (N59, N42, N7, N20, N20);
xor XOR2 (N60, N57, N22);
or OR3 (N61, N47, N37, N35);
nor NOR4 (N62, N29, N2, N17, N19);
xor XOR2 (N63, N61, N39);
nor NOR4 (N64, N53, N50, N60, N57);
xor XOR2 (N65, N61, N33);
or OR3 (N66, N62, N16, N17);
or OR3 (N67, N55, N9, N33);
nor NOR2 (N68, N52, N54);
nor NOR3 (N69, N67, N25, N25);
xor XOR2 (N70, N59, N16);
and AND3 (N71, N70, N5, N12);
nor NOR4 (N72, N64, N52, N19, N61);
and AND3 (N73, N58, N9, N16);
or OR4 (N74, N66, N54, N45, N12);
not NOT1 (N75, N74);
nand NAND4 (N76, N72, N1, N12, N4);
and AND3 (N77, N63, N63, N73);
or OR4 (N78, N12, N16, N34, N37);
not NOT1 (N79, N71);
nor NOR3 (N80, N76, N29, N29);
nand NAND3 (N81, N77, N25, N32);
or OR3 (N82, N75, N36, N62);
xor XOR2 (N83, N79, N73);
nor NOR3 (N84, N78, N81, N14);
nor NOR4 (N85, N41, N10, N13, N43);
nor NOR4 (N86, N82, N82, N79, N65);
or OR3 (N87, N85, N56, N26);
nand NAND4 (N88, N53, N44, N33, N44);
nand NAND2 (N89, N45, N73);
nand NAND4 (N90, N42, N7, N9, N67);
and AND2 (N91, N68, N46);
nand NAND3 (N92, N69, N82, N18);
xor XOR2 (N93, N87, N44);
xor XOR2 (N94, N90, N77);
xor XOR2 (N95, N94, N90);
and AND4 (N96, N84, N77, N83, N24);
xor XOR2 (N97, N33, N44);
or OR2 (N98, N96, N5);
buf BUF1 (N99, N89);
xor XOR2 (N100, N92, N63);
nand NAND3 (N101, N98, N44, N34);
and AND3 (N102, N91, N13, N84);
not NOT1 (N103, N86);
or OR4 (N104, N88, N73, N68, N81);
xor XOR2 (N105, N104, N43);
nor NOR2 (N106, N97, N105);
not NOT1 (N107, N47);
nand NAND2 (N108, N95, N40);
buf BUF1 (N109, N102);
nand NAND4 (N110, N103, N74, N18, N24);
xor XOR2 (N111, N109, N50);
buf BUF1 (N112, N106);
or OR4 (N113, N110, N35, N7, N78);
or OR2 (N114, N80, N52);
not NOT1 (N115, N107);
nand NAND3 (N116, N112, N62, N60);
not NOT1 (N117, N100);
buf BUF1 (N118, N116);
or OR3 (N119, N108, N61, N39);
xor XOR2 (N120, N118, N89);
buf BUF1 (N121, N119);
and AND3 (N122, N120, N121, N87);
nor NOR2 (N123, N80, N81);
not NOT1 (N124, N115);
or OR2 (N125, N101, N14);
and AND4 (N126, N111, N101, N32, N9);
nor NOR4 (N127, N113, N115, N117, N52);
xor XOR2 (N128, N100, N72);
or OR2 (N129, N127, N34);
or OR2 (N130, N99, N108);
or OR2 (N131, N129, N26);
xor XOR2 (N132, N131, N130);
nand NAND3 (N133, N19, N82, N8);
xor XOR2 (N134, N123, N33);
or OR3 (N135, N128, N46, N107);
xor XOR2 (N136, N125, N72);
nand NAND3 (N137, N126, N129, N17);
xor XOR2 (N138, N136, N136);
not NOT1 (N139, N122);
xor XOR2 (N140, N138, N43);
nor NOR4 (N141, N114, N116, N25, N37);
and AND4 (N142, N134, N46, N19, N118);
xor XOR2 (N143, N135, N85);
not NOT1 (N144, N141);
buf BUF1 (N145, N133);
or OR3 (N146, N140, N32, N8);
nor NOR4 (N147, N142, N115, N67, N145);
or OR2 (N148, N112, N142);
buf BUF1 (N149, N124);
nor NOR4 (N150, N148, N104, N70, N87);
buf BUF1 (N151, N149);
nand NAND4 (N152, N139, N106, N115, N79);
nand NAND2 (N153, N144, N50);
and AND4 (N154, N146, N66, N86, N1);
and AND2 (N155, N93, N108);
nand NAND2 (N156, N147, N117);
or OR3 (N157, N150, N149, N67);
and AND4 (N158, N154, N88, N10, N126);
or OR4 (N159, N151, N24, N110, N36);
and AND3 (N160, N155, N53, N132);
nand NAND2 (N161, N18, N34);
buf BUF1 (N162, N153);
not NOT1 (N163, N156);
buf BUF1 (N164, N157);
or OR3 (N165, N143, N15, N42);
nand NAND2 (N166, N165, N85);
nor NOR3 (N167, N164, N70, N28);
nand NAND4 (N168, N162, N94, N126, N40);
or OR3 (N169, N166, N142, N54);
xor XOR2 (N170, N152, N117);
nand NAND4 (N171, N137, N143, N19, N73);
or OR2 (N172, N170, N166);
nand NAND4 (N173, N159, N127, N100, N98);
and AND2 (N174, N167, N123);
buf BUF1 (N175, N174);
and AND2 (N176, N158, N135);
not NOT1 (N177, N175);
and AND2 (N178, N177, N130);
nand NAND2 (N179, N169, N38);
nor NOR3 (N180, N171, N121, N15);
nand NAND3 (N181, N178, N125, N1);
or OR4 (N182, N168, N87, N165, N12);
nor NOR4 (N183, N172, N129, N80, N87);
nor NOR3 (N184, N181, N168, N126);
nor NOR4 (N185, N179, N8, N134, N103);
nor NOR2 (N186, N160, N12);
buf BUF1 (N187, N184);
and AND2 (N188, N186, N105);
not NOT1 (N189, N180);
xor XOR2 (N190, N183, N33);
nand NAND4 (N191, N187, N59, N53, N125);
nor NOR2 (N192, N189, N42);
and AND3 (N193, N163, N173, N120);
or OR4 (N194, N74, N26, N25, N186);
nand NAND3 (N195, N192, N67, N108);
or OR4 (N196, N188, N15, N22, N32);
xor XOR2 (N197, N161, N156);
nor NOR4 (N198, N190, N167, N9, N141);
or OR3 (N199, N191, N19, N119);
nor NOR3 (N200, N193, N127, N20);
xor XOR2 (N201, N194, N148);
nand NAND2 (N202, N199, N49);
not NOT1 (N203, N182);
not NOT1 (N204, N185);
xor XOR2 (N205, N197, N138);
buf BUF1 (N206, N196);
and AND2 (N207, N195, N132);
and AND3 (N208, N205, N105, N108);
not NOT1 (N209, N208);
buf BUF1 (N210, N207);
and AND4 (N211, N204, N12, N47, N65);
and AND2 (N212, N200, N103);
not NOT1 (N213, N176);
nor NOR4 (N214, N210, N197, N111, N21);
not NOT1 (N215, N213);
not NOT1 (N216, N201);
xor XOR2 (N217, N203, N88);
not NOT1 (N218, N212);
nor NOR2 (N219, N211, N185);
buf BUF1 (N220, N206);
nor NOR4 (N221, N219, N133, N49, N10);
or OR3 (N222, N198, N139, N103);
or OR4 (N223, N215, N169, N146, N6);
or OR3 (N224, N221, N187, N120);
nor NOR4 (N225, N223, N97, N131, N191);
buf BUF1 (N226, N216);
nor NOR3 (N227, N222, N196, N24);
nand NAND2 (N228, N218, N94);
nand NAND2 (N229, N227, N167);
buf BUF1 (N230, N226);
xor XOR2 (N231, N220, N224);
not NOT1 (N232, N106);
and AND3 (N233, N231, N157, N89);
and AND4 (N234, N232, N154, N19, N89);
xor XOR2 (N235, N233, N226);
nand NAND2 (N236, N225, N98);
and AND3 (N237, N217, N183, N13);
not NOT1 (N238, N237);
xor XOR2 (N239, N235, N8);
or OR3 (N240, N214, N28, N128);
buf BUF1 (N241, N234);
not NOT1 (N242, N239);
nor NOR4 (N243, N230, N26, N158, N70);
xor XOR2 (N244, N228, N192);
nor NOR4 (N245, N236, N134, N216, N77);
or OR3 (N246, N244, N84, N33);
nor NOR4 (N247, N229, N125, N9, N102);
nand NAND3 (N248, N209, N208, N138);
or OR3 (N249, N246, N167, N176);
xor XOR2 (N250, N245, N219);
buf BUF1 (N251, N243);
or OR4 (N252, N248, N131, N161, N222);
or OR3 (N253, N247, N65, N106);
buf BUF1 (N254, N251);
or OR2 (N255, N202, N235);
xor XOR2 (N256, N240, N158);
and AND4 (N257, N238, N44, N221, N35);
and AND4 (N258, N249, N106, N181, N187);
or OR4 (N259, N256, N68, N26, N26);
nor NOR2 (N260, N252, N25);
xor XOR2 (N261, N255, N224);
or OR4 (N262, N258, N118, N196, N124);
not NOT1 (N263, N241);
not NOT1 (N264, N254);
and AND2 (N265, N261, N35);
nand NAND4 (N266, N262, N210, N44, N85);
xor XOR2 (N267, N259, N214);
not NOT1 (N268, N264);
xor XOR2 (N269, N242, N56);
buf BUF1 (N270, N260);
nand NAND2 (N271, N266, N83);
or OR4 (N272, N257, N159, N32, N250);
buf BUF1 (N273, N178);
buf BUF1 (N274, N273);
buf BUF1 (N275, N267);
not NOT1 (N276, N271);
nor NOR3 (N277, N253, N198, N79);
buf BUF1 (N278, N274);
xor XOR2 (N279, N278, N131);
nand NAND2 (N280, N265, N43);
and AND4 (N281, N280, N78, N259, N112);
not NOT1 (N282, N277);
nor NOR2 (N283, N282, N135);
nor NOR2 (N284, N270, N32);
and AND4 (N285, N272, N112, N58, N89);
not NOT1 (N286, N276);
nand NAND4 (N287, N279, N126, N219, N81);
buf BUF1 (N288, N283);
nand NAND3 (N289, N288, N210, N196);
xor XOR2 (N290, N287, N262);
and AND4 (N291, N263, N282, N33, N119);
nor NOR2 (N292, N284, N95);
or OR4 (N293, N291, N116, N183, N32);
buf BUF1 (N294, N285);
not NOT1 (N295, N293);
nand NAND2 (N296, N269, N174);
nand NAND2 (N297, N290, N255);
and AND3 (N298, N295, N66, N74);
and AND2 (N299, N292, N31);
xor XOR2 (N300, N294, N193);
nand NAND4 (N301, N300, N184, N129, N67);
nor NOR3 (N302, N286, N95, N239);
or OR3 (N303, N301, N129, N39);
xor XOR2 (N304, N302, N81);
buf BUF1 (N305, N297);
not NOT1 (N306, N275);
nand NAND4 (N307, N281, N203, N112, N57);
or OR3 (N308, N307, N251, N100);
xor XOR2 (N309, N303, N307);
buf BUF1 (N310, N299);
and AND4 (N311, N289, N142, N187, N232);
nor NOR4 (N312, N298, N259, N64, N32);
xor XOR2 (N313, N311, N280);
and AND2 (N314, N313, N25);
nor NOR2 (N315, N304, N6);
or OR4 (N316, N309, N279, N29, N27);
not NOT1 (N317, N268);
nor NOR4 (N318, N296, N47, N132, N85);
or OR2 (N319, N310, N232);
xor XOR2 (N320, N315, N185);
not NOT1 (N321, N312);
xor XOR2 (N322, N316, N287);
xor XOR2 (N323, N319, N211);
not NOT1 (N324, N317);
or OR2 (N325, N305, N309);
and AND2 (N326, N323, N77);
buf BUF1 (N327, N308);
xor XOR2 (N328, N322, N267);
not NOT1 (N329, N324);
nor NOR3 (N330, N321, N234, N59);
and AND3 (N331, N327, N176, N32);
nand NAND4 (N332, N331, N313, N128, N253);
nor NOR3 (N333, N328, N22, N297);
xor XOR2 (N334, N314, N260);
nor NOR3 (N335, N332, N99, N175);
not NOT1 (N336, N320);
or OR2 (N337, N336, N236);
buf BUF1 (N338, N330);
xor XOR2 (N339, N337, N311);
and AND4 (N340, N318, N30, N12, N114);
or OR2 (N341, N333, N56);
nor NOR4 (N342, N306, N171, N319, N101);
or OR4 (N343, N341, N130, N198, N267);
nor NOR3 (N344, N326, N116, N15);
or OR2 (N345, N334, N63);
and AND2 (N346, N329, N31);
buf BUF1 (N347, N342);
buf BUF1 (N348, N339);
nor NOR4 (N349, N338, N74, N192, N58);
nor NOR4 (N350, N348, N277, N271, N172);
not NOT1 (N351, N325);
nand NAND4 (N352, N349, N117, N186, N267);
and AND4 (N353, N352, N46, N173, N186);
nand NAND2 (N354, N345, N158);
nand NAND4 (N355, N346, N42, N344, N41);
buf BUF1 (N356, N208);
buf BUF1 (N357, N356);
not NOT1 (N358, N343);
xor XOR2 (N359, N340, N170);
nand NAND2 (N360, N354, N181);
and AND3 (N361, N351, N320, N131);
buf BUF1 (N362, N359);
buf BUF1 (N363, N347);
or OR4 (N364, N335, N153, N80, N18);
not NOT1 (N365, N361);
not NOT1 (N366, N355);
buf BUF1 (N367, N350);
and AND4 (N368, N358, N129, N361, N56);
nand NAND3 (N369, N357, N227, N112);
not NOT1 (N370, N365);
or OR3 (N371, N370, N266, N262);
or OR3 (N372, N371, N104, N30);
or OR2 (N373, N366, N333);
or OR3 (N374, N363, N253, N343);
nor NOR4 (N375, N362, N280, N356, N205);
nand NAND4 (N376, N369, N260, N373, N370);
and AND2 (N377, N46, N23);
nor NOR3 (N378, N360, N373, N322);
nor NOR4 (N379, N375, N292, N27, N263);
not NOT1 (N380, N374);
xor XOR2 (N381, N364, N220);
nor NOR4 (N382, N376, N20, N31, N187);
buf BUF1 (N383, N367);
and AND3 (N384, N379, N165, N21);
nand NAND4 (N385, N372, N267, N97, N197);
xor XOR2 (N386, N383, N144);
and AND2 (N387, N353, N164);
or OR2 (N388, N380, N196);
nor NOR2 (N389, N382, N85);
xor XOR2 (N390, N389, N57);
buf BUF1 (N391, N378);
not NOT1 (N392, N377);
and AND3 (N393, N390, N2, N173);
nand NAND4 (N394, N387, N99, N178, N294);
nand NAND3 (N395, N385, N25, N202);
nor NOR4 (N396, N391, N389, N395, N187);
nand NAND4 (N397, N151, N360, N7, N89);
and AND3 (N398, N392, N270, N363);
xor XOR2 (N399, N396, N127);
nand NAND2 (N400, N368, N384);
nand NAND3 (N401, N250, N10, N25);
nand NAND4 (N402, N398, N26, N191, N328);
buf BUF1 (N403, N401);
nand NAND2 (N404, N381, N16);
nand NAND2 (N405, N394, N68);
xor XOR2 (N406, N403, N130);
nor NOR4 (N407, N399, N391, N256, N110);
xor XOR2 (N408, N406, N367);
xor XOR2 (N409, N402, N89);
or OR4 (N410, N386, N127, N33, N362);
buf BUF1 (N411, N407);
nor NOR2 (N412, N400, N256);
buf BUF1 (N413, N393);
not NOT1 (N414, N411);
or OR3 (N415, N410, N275, N200);
and AND3 (N416, N412, N27, N55);
nand NAND4 (N417, N397, N62, N250, N184);
not NOT1 (N418, N408);
not NOT1 (N419, N388);
buf BUF1 (N420, N409);
buf BUF1 (N421, N415);
nand NAND4 (N422, N420, N103, N14, N301);
xor XOR2 (N423, N418, N362);
buf BUF1 (N424, N423);
and AND4 (N425, N417, N1, N293, N124);
xor XOR2 (N426, N404, N110);
buf BUF1 (N427, N414);
not NOT1 (N428, N421);
nor NOR4 (N429, N416, N381, N217, N120);
and AND3 (N430, N419, N180, N149);
nand NAND2 (N431, N425, N155);
buf BUF1 (N432, N429);
xor XOR2 (N433, N432, N270);
and AND2 (N434, N433, N6);
nand NAND2 (N435, N422, N358);
or OR4 (N436, N405, N195, N29, N255);
xor XOR2 (N437, N436, N95);
buf BUF1 (N438, N431);
nor NOR2 (N439, N413, N325);
nand NAND4 (N440, N437, N105, N315, N127);
buf BUF1 (N441, N434);
nand NAND2 (N442, N439, N145);
or OR3 (N443, N440, N72, N330);
nand NAND4 (N444, N438, N115, N192, N246);
and AND4 (N445, N444, N6, N6, N81);
not NOT1 (N446, N424);
and AND4 (N447, N435, N73, N302, N318);
or OR2 (N448, N442, N342);
nand NAND2 (N449, N428, N425);
not NOT1 (N450, N447);
and AND4 (N451, N427, N398, N99, N374);
and AND2 (N452, N441, N289);
nand NAND3 (N453, N446, N436, N65);
and AND2 (N454, N430, N159);
and AND3 (N455, N445, N380, N139);
buf BUF1 (N456, N450);
not NOT1 (N457, N448);
not NOT1 (N458, N455);
or OR2 (N459, N457, N417);
nand NAND3 (N460, N453, N373, N361);
xor XOR2 (N461, N458, N107);
not NOT1 (N462, N460);
and AND3 (N463, N426, N51, N279);
xor XOR2 (N464, N456, N291);
not NOT1 (N465, N459);
nand NAND3 (N466, N463, N10, N123);
nand NAND3 (N467, N465, N237, N149);
xor XOR2 (N468, N443, N373);
and AND4 (N469, N461, N285, N456, N79);
xor XOR2 (N470, N449, N161);
nor NOR3 (N471, N469, N400, N365);
and AND3 (N472, N470, N54, N415);
or OR3 (N473, N462, N164, N288);
or OR2 (N474, N466, N57);
buf BUF1 (N475, N452);
nor NOR4 (N476, N454, N298, N97, N359);
and AND4 (N477, N451, N220, N340, N363);
nor NOR4 (N478, N471, N8, N296, N229);
nor NOR2 (N479, N472, N440);
buf BUF1 (N480, N473);
not NOT1 (N481, N467);
not NOT1 (N482, N479);
xor XOR2 (N483, N468, N455);
nor NOR4 (N484, N480, N190, N464, N41);
buf BUF1 (N485, N18);
nand NAND2 (N486, N474, N125);
buf BUF1 (N487, N478);
not NOT1 (N488, N476);
or OR4 (N489, N483, N205, N287, N255);
nor NOR4 (N490, N489, N378, N116, N386);
or OR4 (N491, N485, N274, N74, N98);
and AND3 (N492, N486, N210, N184);
buf BUF1 (N493, N477);
not NOT1 (N494, N488);
xor XOR2 (N495, N475, N461);
buf BUF1 (N496, N491);
nand NAND2 (N497, N493, N99);
buf BUF1 (N498, N496);
and AND4 (N499, N482, N360, N73, N103);
or OR3 (N500, N499, N166, N486);
and AND3 (N501, N492, N403, N120);
buf BUF1 (N502, N500);
or OR3 (N503, N501, N69, N336);
or OR3 (N504, N497, N274, N352);
or OR3 (N505, N484, N9, N56);
xor XOR2 (N506, N498, N359);
nand NAND4 (N507, N504, N316, N221, N202);
nand NAND3 (N508, N502, N153, N493);
xor XOR2 (N509, N487, N74);
not NOT1 (N510, N509);
nor NOR4 (N511, N490, N495, N134, N41);
not NOT1 (N512, N113);
nand NAND3 (N513, N512, N89, N365);
not NOT1 (N514, N506);
and AND2 (N515, N481, N333);
xor XOR2 (N516, N494, N233);
buf BUF1 (N517, N515);
buf BUF1 (N518, N508);
not NOT1 (N519, N510);
nand NAND3 (N520, N517, N3, N279);
or OR2 (N521, N518, N445);
xor XOR2 (N522, N507, N355);
xor XOR2 (N523, N516, N104);
and AND3 (N524, N505, N484, N384);
not NOT1 (N525, N513);
buf BUF1 (N526, N519);
buf BUF1 (N527, N522);
buf BUF1 (N528, N514);
not NOT1 (N529, N526);
nor NOR3 (N530, N503, N217, N462);
nor NOR2 (N531, N529, N96);
nor NOR4 (N532, N521, N490, N397, N399);
xor XOR2 (N533, N511, N151);
buf BUF1 (N534, N532);
xor XOR2 (N535, N530, N128);
buf BUF1 (N536, N524);
xor XOR2 (N537, N527, N65);
xor XOR2 (N538, N536, N242);
not NOT1 (N539, N523);
not NOT1 (N540, N531);
nand NAND3 (N541, N528, N87, N203);
and AND4 (N542, N538, N389, N265, N77);
nor NOR4 (N543, N540, N469, N10, N109);
and AND4 (N544, N539, N202, N328, N298);
buf BUF1 (N545, N535);
not NOT1 (N546, N543);
and AND3 (N547, N545, N44, N91);
buf BUF1 (N548, N542);
nor NOR4 (N549, N544, N301, N132, N199);
or OR4 (N550, N547, N27, N213, N31);
and AND3 (N551, N533, N401, N205);
nand NAND4 (N552, N550, N280, N98, N520);
nor NOR2 (N553, N17, N112);
nand NAND3 (N554, N549, N450, N423);
nor NOR4 (N555, N525, N275, N356, N497);
and AND2 (N556, N541, N84);
not NOT1 (N557, N537);
nand NAND2 (N558, N551, N245);
or OR3 (N559, N552, N362, N280);
and AND3 (N560, N548, N473, N181);
not NOT1 (N561, N558);
xor XOR2 (N562, N556, N423);
buf BUF1 (N563, N554);
or OR2 (N564, N563, N247);
buf BUF1 (N565, N557);
xor XOR2 (N566, N561, N130);
or OR2 (N567, N566, N146);
or OR4 (N568, N546, N440, N182, N40);
nand NAND3 (N569, N560, N513, N165);
or OR3 (N570, N567, N396, N538);
nand NAND3 (N571, N559, N76, N221);
nor NOR3 (N572, N534, N110, N13);
and AND4 (N573, N569, N52, N530, N99);
and AND4 (N574, N572, N569, N545, N118);
and AND2 (N575, N565, N103);
or OR2 (N576, N571, N118);
not NOT1 (N577, N555);
and AND4 (N578, N577, N360, N410, N223);
nor NOR2 (N579, N562, N457);
buf BUF1 (N580, N568);
nor NOR4 (N581, N579, N250, N162, N338);
buf BUF1 (N582, N564);
buf BUF1 (N583, N580);
buf BUF1 (N584, N581);
not NOT1 (N585, N570);
and AND2 (N586, N585, N180);
buf BUF1 (N587, N586);
xor XOR2 (N588, N582, N30);
buf BUF1 (N589, N553);
nand NAND3 (N590, N573, N269, N341);
and AND2 (N591, N575, N141);
xor XOR2 (N592, N590, N174);
and AND2 (N593, N588, N464);
or OR2 (N594, N589, N4);
buf BUF1 (N595, N576);
xor XOR2 (N596, N595, N236);
not NOT1 (N597, N591);
nand NAND3 (N598, N594, N331, N34);
xor XOR2 (N599, N592, N96);
xor XOR2 (N600, N598, N547);
xor XOR2 (N601, N596, N111);
buf BUF1 (N602, N599);
or OR4 (N603, N601, N186, N219, N2);
not NOT1 (N604, N584);
nand NAND4 (N605, N602, N40, N462, N450);
xor XOR2 (N606, N603, N579);
nand NAND2 (N607, N606, N540);
and AND2 (N608, N578, N50);
buf BUF1 (N609, N593);
xor XOR2 (N610, N605, N446);
or OR2 (N611, N600, N512);
xor XOR2 (N612, N611, N17);
xor XOR2 (N613, N604, N340);
or OR3 (N614, N612, N577, N399);
nand NAND4 (N615, N610, N362, N21, N568);
nor NOR2 (N616, N597, N321);
not NOT1 (N617, N587);
xor XOR2 (N618, N583, N323);
nand NAND2 (N619, N613, N102);
nand NAND4 (N620, N617, N318, N413, N250);
buf BUF1 (N621, N620);
xor XOR2 (N622, N574, N165);
nor NOR2 (N623, N618, N422);
and AND3 (N624, N607, N158, N24);
nor NOR3 (N625, N619, N302, N542);
nor NOR4 (N626, N624, N299, N255, N126);
or OR2 (N627, N615, N593);
xor XOR2 (N628, N623, N558);
nor NOR2 (N629, N621, N283);
not NOT1 (N630, N628);
xor XOR2 (N631, N608, N416);
xor XOR2 (N632, N614, N318);
nand NAND3 (N633, N625, N445, N533);
not NOT1 (N634, N631);
not NOT1 (N635, N630);
buf BUF1 (N636, N622);
buf BUF1 (N637, N609);
not NOT1 (N638, N627);
not NOT1 (N639, N633);
not NOT1 (N640, N629);
nand NAND3 (N641, N637, N157, N461);
nor NOR3 (N642, N632, N558, N324);
buf BUF1 (N643, N636);
or OR2 (N644, N616, N20);
or OR4 (N645, N642, N560, N259, N27);
not NOT1 (N646, N634);
nand NAND2 (N647, N626, N267);
nor NOR4 (N648, N638, N254, N305, N641);
buf BUF1 (N649, N340);
not NOT1 (N650, N647);
nand NAND2 (N651, N645, N511);
buf BUF1 (N652, N649);
nand NAND4 (N653, N652, N509, N572, N487);
or OR2 (N654, N646, N617);
buf BUF1 (N655, N635);
not NOT1 (N656, N655);
and AND4 (N657, N648, N227, N91, N175);
xor XOR2 (N658, N640, N8);
xor XOR2 (N659, N644, N287);
nor NOR4 (N660, N651, N473, N342, N109);
xor XOR2 (N661, N653, N516);
xor XOR2 (N662, N650, N46);
xor XOR2 (N663, N660, N293);
nand NAND4 (N664, N662, N139, N467, N572);
or OR4 (N665, N657, N567, N288, N440);
or OR2 (N666, N663, N634);
or OR2 (N667, N639, N104);
nand NAND3 (N668, N659, N561, N233);
not NOT1 (N669, N664);
or OR3 (N670, N667, N112, N227);
xor XOR2 (N671, N669, N629);
nor NOR3 (N672, N665, N510, N346);
xor XOR2 (N673, N656, N91);
xor XOR2 (N674, N670, N601);
or OR4 (N675, N672, N158, N445, N36);
not NOT1 (N676, N675);
xor XOR2 (N677, N658, N5);
not NOT1 (N678, N668);
xor XOR2 (N679, N673, N12);
and AND2 (N680, N674, N80);
xor XOR2 (N681, N643, N497);
or OR2 (N682, N680, N505);
xor XOR2 (N683, N676, N31);
and AND3 (N684, N679, N157, N96);
nand NAND4 (N685, N654, N592, N232, N325);
xor XOR2 (N686, N666, N229);
nand NAND2 (N687, N683, N29);
or OR3 (N688, N684, N520, N42);
or OR3 (N689, N681, N322, N322);
xor XOR2 (N690, N682, N573);
nor NOR3 (N691, N677, N634, N194);
nor NOR4 (N692, N689, N557, N594, N558);
xor XOR2 (N693, N692, N663);
nand NAND4 (N694, N661, N202, N113, N43);
xor XOR2 (N695, N691, N141);
buf BUF1 (N696, N695);
xor XOR2 (N697, N690, N87);
buf BUF1 (N698, N678);
and AND3 (N699, N686, N399, N601);
not NOT1 (N700, N693);
nor NOR2 (N701, N685, N186);
nand NAND4 (N702, N698, N14, N560, N638);
and AND4 (N703, N694, N695, N518, N424);
buf BUF1 (N704, N688);
or OR4 (N705, N701, N437, N683, N388);
nand NAND3 (N706, N700, N99, N559);
nand NAND2 (N707, N703, N369);
or OR3 (N708, N704, N665, N573);
not NOT1 (N709, N696);
xor XOR2 (N710, N671, N459);
xor XOR2 (N711, N697, N132);
and AND4 (N712, N709, N162, N305, N331);
and AND3 (N713, N705, N355, N665);
or OR2 (N714, N710, N690);
nor NOR3 (N715, N713, N434, N673);
xor XOR2 (N716, N699, N163);
not NOT1 (N717, N711);
nor NOR4 (N718, N702, N249, N242, N556);
or OR2 (N719, N706, N235);
and AND2 (N720, N719, N388);
not NOT1 (N721, N714);
or OR2 (N722, N715, N468);
and AND3 (N723, N721, N602, N418);
or OR2 (N724, N723, N39);
endmodule