// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N491,N501,N509,N504,N495,N508,N502,N507,N485,N510;

and AND2 (N11, N1, N4);
or OR3 (N12, N2, N8, N9);
xor XOR2 (N13, N10, N9);
buf BUF1 (N14, N5);
nand NAND4 (N15, N1, N10, N14, N7);
xor XOR2 (N16, N10, N9);
nor NOR4 (N17, N5, N6, N11, N9);
nor NOR3 (N18, N2, N15, N7);
or OR3 (N19, N15, N18, N13);
not NOT1 (N20, N7);
not NOT1 (N21, N7);
buf BUF1 (N22, N1);
or OR4 (N23, N21, N17, N6, N5);
not NOT1 (N24, N10);
buf BUF1 (N25, N13);
not NOT1 (N26, N18);
xor XOR2 (N27, N18, N5);
or OR2 (N28, N23, N11);
not NOT1 (N29, N27);
nand NAND4 (N30, N26, N12, N23, N15);
nor NOR2 (N31, N11, N5);
and AND4 (N32, N25, N29, N20, N20);
nand NAND2 (N33, N30, N10);
buf BUF1 (N34, N8);
nand NAND2 (N35, N19, N14);
buf BUF1 (N36, N14);
buf BUF1 (N37, N28);
or OR3 (N38, N31, N8, N7);
nor NOR3 (N39, N36, N24, N33);
or OR4 (N40, N17, N9, N33, N22);
nor NOR4 (N41, N33, N1, N6, N4);
or OR2 (N42, N10, N28);
nor NOR3 (N43, N35, N33, N9);
xor XOR2 (N44, N32, N26);
not NOT1 (N45, N43);
buf BUF1 (N46, N38);
and AND2 (N47, N45, N17);
or OR4 (N48, N42, N35, N20, N1);
xor XOR2 (N49, N41, N34);
buf BUF1 (N50, N48);
nor NOR2 (N51, N17, N44);
xor XOR2 (N52, N26, N45);
nor NOR2 (N53, N49, N8);
nand NAND2 (N54, N51, N2);
xor XOR2 (N55, N16, N39);
nor NOR4 (N56, N21, N27, N29, N22);
buf BUF1 (N57, N46);
xor XOR2 (N58, N56, N29);
not NOT1 (N59, N50);
nor NOR2 (N60, N59, N24);
not NOT1 (N61, N47);
xor XOR2 (N62, N54, N33);
not NOT1 (N63, N40);
nand NAND4 (N64, N37, N50, N1, N29);
and AND3 (N65, N64, N47, N34);
xor XOR2 (N66, N65, N62);
xor XOR2 (N67, N24, N24);
xor XOR2 (N68, N60, N51);
and AND2 (N69, N63, N61);
buf BUF1 (N70, N25);
or OR3 (N71, N68, N5, N61);
nand NAND2 (N72, N67, N52);
or OR4 (N73, N31, N37, N3, N41);
not NOT1 (N74, N71);
nor NOR3 (N75, N55, N25, N70);
and AND3 (N76, N61, N67, N14);
nor NOR3 (N77, N69, N74, N40);
buf BUF1 (N78, N28);
or OR3 (N79, N53, N1, N9);
buf BUF1 (N80, N76);
nand NAND4 (N81, N73, N33, N30, N78);
xor XOR2 (N82, N74, N51);
or OR4 (N83, N81, N15, N37, N45);
or OR2 (N84, N77, N69);
nand NAND2 (N85, N84, N49);
nand NAND2 (N86, N82, N2);
nand NAND2 (N87, N80, N25);
not NOT1 (N88, N86);
not NOT1 (N89, N75);
not NOT1 (N90, N85);
buf BUF1 (N91, N66);
and AND2 (N92, N87, N77);
nand NAND3 (N93, N57, N83, N80);
and AND4 (N94, N45, N27, N64, N15);
or OR3 (N95, N91, N70, N7);
buf BUF1 (N96, N95);
or OR2 (N97, N90, N51);
nor NOR4 (N98, N79, N37, N21, N18);
buf BUF1 (N99, N98);
or OR2 (N100, N72, N93);
and AND2 (N101, N67, N16);
not NOT1 (N102, N92);
and AND2 (N103, N89, N44);
buf BUF1 (N104, N99);
nand NAND2 (N105, N97, N51);
buf BUF1 (N106, N104);
and AND3 (N107, N58, N104, N1);
or OR4 (N108, N103, N56, N30, N64);
or OR3 (N109, N108, N83, N58);
xor XOR2 (N110, N94, N24);
buf BUF1 (N111, N106);
nand NAND4 (N112, N88, N62, N74, N95);
or OR2 (N113, N102, N78);
xor XOR2 (N114, N101, N112);
and AND3 (N115, N68, N71, N53);
or OR2 (N116, N110, N84);
and AND3 (N117, N113, N26, N94);
xor XOR2 (N118, N116, N93);
or OR2 (N119, N96, N82);
and AND4 (N120, N109, N105, N44, N62);
buf BUF1 (N121, N35);
nand NAND2 (N122, N107, N8);
and AND4 (N123, N119, N89, N28, N56);
not NOT1 (N124, N120);
xor XOR2 (N125, N114, N57);
xor XOR2 (N126, N125, N25);
buf BUF1 (N127, N111);
nor NOR4 (N128, N123, N111, N25, N60);
and AND2 (N129, N100, N34);
nand NAND3 (N130, N115, N94, N102);
not NOT1 (N131, N117);
nand NAND3 (N132, N121, N120, N2);
nand NAND3 (N133, N131, N41, N130);
nor NOR2 (N134, N12, N124);
xor XOR2 (N135, N3, N5);
or OR4 (N136, N134, N84, N130, N41);
nor NOR4 (N137, N127, N76, N95, N23);
buf BUF1 (N138, N126);
buf BUF1 (N139, N138);
or OR4 (N140, N133, N110, N121, N41);
nor NOR4 (N141, N122, N16, N70, N67);
nand NAND3 (N142, N137, N35, N94);
nand NAND3 (N143, N142, N76, N37);
and AND2 (N144, N132, N63);
or OR3 (N145, N140, N27, N78);
or OR4 (N146, N141, N45, N82, N96);
nand NAND2 (N147, N143, N74);
xor XOR2 (N148, N139, N75);
or OR3 (N149, N146, N106, N22);
not NOT1 (N150, N149);
nor NOR2 (N151, N135, N29);
nor NOR3 (N152, N136, N62, N85);
not NOT1 (N153, N152);
and AND4 (N154, N147, N35, N86, N73);
nand NAND3 (N155, N151, N133, N130);
nor NOR4 (N156, N145, N23, N141, N100);
not NOT1 (N157, N144);
not NOT1 (N158, N118);
buf BUF1 (N159, N150);
nor NOR3 (N160, N155, N64, N25);
and AND4 (N161, N158, N153, N70, N63);
nand NAND2 (N162, N121, N26);
buf BUF1 (N163, N156);
nand NAND3 (N164, N148, N84, N79);
not NOT1 (N165, N162);
xor XOR2 (N166, N165, N118);
nand NAND3 (N167, N164, N136, N29);
buf BUF1 (N168, N157);
and AND2 (N169, N160, N97);
not NOT1 (N170, N154);
xor XOR2 (N171, N163, N108);
nor NOR4 (N172, N171, N70, N31, N50);
not NOT1 (N173, N168);
xor XOR2 (N174, N167, N12);
not NOT1 (N175, N161);
or OR2 (N176, N173, N31);
and AND3 (N177, N128, N10, N141);
or OR2 (N178, N174, N104);
xor XOR2 (N179, N178, N46);
nand NAND2 (N180, N129, N58);
nor NOR4 (N181, N159, N85, N158, N140);
and AND4 (N182, N179, N38, N101, N110);
nor NOR3 (N183, N172, N61, N106);
nor NOR3 (N184, N166, N173, N154);
xor XOR2 (N185, N175, N150);
not NOT1 (N186, N185);
or OR2 (N187, N183, N110);
buf BUF1 (N188, N177);
or OR4 (N189, N170, N153, N4, N52);
buf BUF1 (N190, N180);
and AND3 (N191, N184, N54, N71);
nand NAND4 (N192, N182, N146, N116, N96);
nand NAND4 (N193, N189, N144, N22, N70);
xor XOR2 (N194, N192, N41);
nand NAND4 (N195, N169, N51, N169, N166);
nor NOR4 (N196, N191, N8, N123, N86);
and AND3 (N197, N181, N14, N154);
nor NOR2 (N198, N195, N196);
and AND2 (N199, N33, N62);
or OR3 (N200, N197, N80, N113);
nand NAND2 (N201, N176, N91);
buf BUF1 (N202, N194);
or OR2 (N203, N201, N148);
buf BUF1 (N204, N187);
nor NOR3 (N205, N198, N85, N55);
not NOT1 (N206, N199);
or OR4 (N207, N186, N72, N16, N89);
xor XOR2 (N208, N200, N191);
and AND3 (N209, N207, N166, N67);
and AND2 (N210, N203, N24);
nor NOR2 (N211, N208, N67);
not NOT1 (N212, N210);
nand NAND4 (N213, N211, N33, N155, N197);
nand NAND4 (N214, N190, N204, N160, N28);
nand NAND4 (N215, N127, N81, N104, N58);
nand NAND2 (N216, N202, N37);
or OR2 (N217, N213, N88);
nand NAND4 (N218, N209, N74, N110, N81);
buf BUF1 (N219, N217);
nand NAND4 (N220, N215, N8, N101, N70);
nand NAND2 (N221, N188, N84);
nor NOR2 (N222, N193, N137);
and AND4 (N223, N216, N171, N169, N188);
nand NAND4 (N224, N218, N145, N159, N10);
or OR3 (N225, N222, N43, N30);
not NOT1 (N226, N225);
and AND2 (N227, N205, N128);
or OR4 (N228, N220, N30, N90, N170);
buf BUF1 (N229, N221);
or OR3 (N230, N219, N98, N191);
or OR2 (N231, N206, N150);
or OR3 (N232, N226, N226, N13);
buf BUF1 (N233, N228);
buf BUF1 (N234, N231);
not NOT1 (N235, N227);
and AND2 (N236, N223, N19);
not NOT1 (N237, N236);
buf BUF1 (N238, N232);
and AND4 (N239, N235, N129, N235, N121);
xor XOR2 (N240, N237, N60);
and AND3 (N241, N214, N198, N3);
buf BUF1 (N242, N241);
or OR4 (N243, N224, N27, N164, N74);
xor XOR2 (N244, N240, N132);
xor XOR2 (N245, N233, N109);
buf BUF1 (N246, N238);
nand NAND4 (N247, N246, N155, N242, N94);
nand NAND3 (N248, N41, N196, N92);
nor NOR4 (N249, N245, N172, N202, N208);
not NOT1 (N250, N239);
nand NAND3 (N251, N248, N56, N181);
buf BUF1 (N252, N212);
or OR4 (N253, N251, N246, N62, N227);
nor NOR4 (N254, N229, N22, N168, N72);
xor XOR2 (N255, N234, N41);
and AND2 (N256, N254, N163);
buf BUF1 (N257, N230);
and AND3 (N258, N250, N201, N101);
nor NOR2 (N259, N255, N227);
xor XOR2 (N260, N256, N39);
buf BUF1 (N261, N249);
xor XOR2 (N262, N252, N111);
or OR2 (N263, N253, N51);
not NOT1 (N264, N243);
not NOT1 (N265, N264);
not NOT1 (N266, N262);
and AND4 (N267, N261, N263, N113, N82);
nor NOR2 (N268, N257, N73);
nor NOR2 (N269, N235, N181);
not NOT1 (N270, N244);
buf BUF1 (N271, N268);
xor XOR2 (N272, N247, N134);
nor NOR4 (N273, N267, N162, N28, N223);
xor XOR2 (N274, N258, N163);
and AND3 (N275, N265, N180, N143);
or OR3 (N276, N272, N222, N82);
nand NAND4 (N277, N274, N263, N53, N144);
xor XOR2 (N278, N276, N232);
not NOT1 (N279, N271);
and AND2 (N280, N275, N31);
nor NOR3 (N281, N270, N155, N111);
nor NOR3 (N282, N279, N50, N48);
buf BUF1 (N283, N282);
nand NAND3 (N284, N281, N44, N36);
xor XOR2 (N285, N273, N63);
buf BUF1 (N286, N260);
and AND2 (N287, N285, N68);
nand NAND2 (N288, N266, N146);
nor NOR3 (N289, N288, N252, N133);
and AND3 (N290, N286, N18, N86);
and AND3 (N291, N278, N7, N19);
nor NOR4 (N292, N259, N43, N70, N4);
buf BUF1 (N293, N287);
not NOT1 (N294, N290);
buf BUF1 (N295, N294);
buf BUF1 (N296, N277);
or OR2 (N297, N284, N109);
xor XOR2 (N298, N269, N176);
xor XOR2 (N299, N291, N22);
nor NOR4 (N300, N292, N118, N108, N118);
or OR2 (N301, N296, N77);
and AND2 (N302, N300, N140);
or OR2 (N303, N299, N55);
not NOT1 (N304, N289);
buf BUF1 (N305, N304);
not NOT1 (N306, N298);
not NOT1 (N307, N306);
nor NOR4 (N308, N303, N131, N31, N165);
nor NOR4 (N309, N295, N116, N290, N141);
not NOT1 (N310, N302);
buf BUF1 (N311, N310);
not NOT1 (N312, N307);
or OR2 (N313, N280, N193);
or OR2 (N314, N313, N267);
nor NOR3 (N315, N309, N236, N289);
nor NOR4 (N316, N297, N21, N229, N244);
xor XOR2 (N317, N312, N119);
nor NOR4 (N318, N317, N20, N41, N113);
nand NAND4 (N319, N305, N179, N273, N63);
nor NOR2 (N320, N318, N82);
nor NOR2 (N321, N283, N121);
nor NOR3 (N322, N314, N247, N55);
and AND2 (N323, N308, N57);
buf BUF1 (N324, N293);
nor NOR2 (N325, N311, N228);
not NOT1 (N326, N324);
or OR4 (N327, N315, N153, N27, N9);
or OR3 (N328, N316, N163, N175);
or OR3 (N329, N319, N39, N280);
buf BUF1 (N330, N322);
or OR2 (N331, N321, N70);
xor XOR2 (N332, N330, N94);
buf BUF1 (N333, N328);
xor XOR2 (N334, N331, N254);
nor NOR3 (N335, N327, N65, N241);
nor NOR4 (N336, N334, N267, N26, N66);
and AND2 (N337, N333, N27);
not NOT1 (N338, N301);
and AND2 (N339, N323, N196);
not NOT1 (N340, N325);
nand NAND3 (N341, N339, N274, N271);
nand NAND4 (N342, N320, N306, N59, N102);
buf BUF1 (N343, N335);
or OR4 (N344, N340, N98, N327, N2);
and AND3 (N345, N342, N128, N343);
not NOT1 (N346, N328);
nor NOR3 (N347, N337, N150, N12);
nor NOR3 (N348, N326, N15, N104);
or OR2 (N349, N347, N305);
not NOT1 (N350, N341);
and AND4 (N351, N338, N127, N93, N188);
nor NOR3 (N352, N349, N170, N83);
or OR2 (N353, N348, N289);
buf BUF1 (N354, N353);
not NOT1 (N355, N345);
nor NOR4 (N356, N329, N169, N75, N169);
and AND2 (N357, N352, N326);
nor NOR2 (N358, N356, N333);
xor XOR2 (N359, N351, N274);
nor NOR3 (N360, N359, N133, N87);
and AND3 (N361, N336, N39, N337);
not NOT1 (N362, N350);
nor NOR2 (N363, N346, N119);
xor XOR2 (N364, N360, N44);
nor NOR4 (N365, N363, N19, N296, N88);
or OR4 (N366, N362, N152, N176, N346);
not NOT1 (N367, N358);
and AND3 (N368, N354, N183, N174);
xor XOR2 (N369, N357, N231);
nor NOR3 (N370, N367, N40, N352);
buf BUF1 (N371, N361);
not NOT1 (N372, N355);
buf BUF1 (N373, N372);
nand NAND3 (N374, N344, N293, N289);
nor NOR4 (N375, N371, N28, N18, N58);
not NOT1 (N376, N332);
xor XOR2 (N377, N369, N123);
nand NAND2 (N378, N365, N3);
nand NAND2 (N379, N368, N66);
nand NAND2 (N380, N375, N161);
xor XOR2 (N381, N380, N297);
xor XOR2 (N382, N374, N29);
and AND4 (N383, N382, N214, N350, N352);
nand NAND2 (N384, N378, N368);
and AND2 (N385, N373, N298);
nand NAND4 (N386, N364, N101, N173, N282);
xor XOR2 (N387, N366, N173);
xor XOR2 (N388, N385, N275);
nand NAND2 (N389, N383, N279);
buf BUF1 (N390, N377);
nor NOR3 (N391, N389, N272, N22);
xor XOR2 (N392, N386, N304);
buf BUF1 (N393, N370);
nand NAND3 (N394, N387, N93, N9);
buf BUF1 (N395, N381);
and AND2 (N396, N393, N40);
xor XOR2 (N397, N395, N62);
and AND4 (N398, N391, N73, N137, N42);
and AND3 (N399, N396, N47, N71);
nor NOR4 (N400, N399, N366, N198, N288);
nand NAND2 (N401, N392, N232);
and AND3 (N402, N390, N337, N25);
or OR3 (N403, N402, N100, N320);
nor NOR3 (N404, N401, N48, N376);
nand NAND2 (N405, N226, N234);
nand NAND4 (N406, N394, N284, N44, N328);
nor NOR2 (N407, N400, N209);
and AND3 (N408, N403, N228, N365);
nor NOR3 (N409, N407, N28, N381);
not NOT1 (N410, N408);
and AND3 (N411, N384, N33, N49);
buf BUF1 (N412, N398);
buf BUF1 (N413, N406);
buf BUF1 (N414, N388);
and AND3 (N415, N379, N49, N114);
and AND2 (N416, N411, N380);
nand NAND4 (N417, N404, N383, N234, N124);
and AND3 (N418, N414, N242, N131);
buf BUF1 (N419, N413);
buf BUF1 (N420, N410);
nor NOR3 (N421, N397, N182, N101);
not NOT1 (N422, N420);
and AND3 (N423, N421, N201, N112);
not NOT1 (N424, N416);
nand NAND2 (N425, N418, N368);
nor NOR2 (N426, N425, N367);
nor NOR4 (N427, N405, N89, N242, N254);
and AND3 (N428, N419, N249, N409);
or OR4 (N429, N232, N134, N224, N328);
xor XOR2 (N430, N423, N180);
nor NOR3 (N431, N426, N219, N311);
buf BUF1 (N432, N417);
buf BUF1 (N433, N427);
nor NOR2 (N434, N415, N85);
and AND2 (N435, N429, N100);
nor NOR4 (N436, N430, N334, N366, N1);
and AND2 (N437, N432, N340);
nor NOR4 (N438, N436, N51, N184, N282);
buf BUF1 (N439, N422);
or OR3 (N440, N412, N352, N109);
xor XOR2 (N441, N431, N193);
xor XOR2 (N442, N437, N71);
not NOT1 (N443, N433);
and AND2 (N444, N440, N337);
buf BUF1 (N445, N434);
buf BUF1 (N446, N439);
nor NOR3 (N447, N438, N135, N419);
or OR2 (N448, N445, N122);
buf BUF1 (N449, N435);
nand NAND2 (N450, N441, N152);
nand NAND3 (N451, N450, N213, N228);
nor NOR3 (N452, N444, N312, N394);
xor XOR2 (N453, N448, N197);
buf BUF1 (N454, N424);
nor NOR3 (N455, N446, N99, N357);
nor NOR2 (N456, N447, N198);
and AND3 (N457, N443, N246, N253);
and AND2 (N458, N428, N287);
nor NOR4 (N459, N455, N223, N271, N406);
buf BUF1 (N460, N457);
or OR4 (N461, N452, N142, N349, N125);
not NOT1 (N462, N451);
or OR2 (N463, N442, N99);
or OR3 (N464, N461, N398, N228);
not NOT1 (N465, N454);
or OR2 (N466, N462, N366);
not NOT1 (N467, N459);
buf BUF1 (N468, N460);
not NOT1 (N469, N453);
nor NOR4 (N470, N464, N427, N397, N251);
or OR3 (N471, N466, N117, N64);
nand NAND3 (N472, N463, N463, N288);
and AND2 (N473, N469, N238);
nor NOR2 (N474, N471, N164);
not NOT1 (N475, N470);
xor XOR2 (N476, N449, N288);
xor XOR2 (N477, N467, N451);
nor NOR2 (N478, N475, N40);
and AND4 (N479, N476, N133, N19, N400);
or OR3 (N480, N456, N193, N358);
or OR4 (N481, N478, N218, N14, N336);
or OR3 (N482, N481, N193, N391);
buf BUF1 (N483, N479);
or OR2 (N484, N474, N433);
not NOT1 (N485, N458);
buf BUF1 (N486, N473);
buf BUF1 (N487, N480);
nand NAND3 (N488, N487, N29, N378);
and AND2 (N489, N482, N144);
nor NOR3 (N490, N483, N40, N181);
xor XOR2 (N491, N490, N392);
buf BUF1 (N492, N484);
buf BUF1 (N493, N492);
not NOT1 (N494, N472);
not NOT1 (N495, N494);
nor NOR3 (N496, N465, N407, N145);
not NOT1 (N497, N488);
and AND2 (N498, N477, N355);
and AND3 (N499, N497, N403, N299);
nor NOR3 (N500, N489, N387, N379);
xor XOR2 (N501, N486, N34);
or OR2 (N502, N496, N34);
buf BUF1 (N503, N493);
nor NOR4 (N504, N503, N302, N497, N180);
or OR3 (N505, N499, N280, N371);
or OR2 (N506, N500, N73);
buf BUF1 (N507, N506);
nor NOR4 (N508, N505, N450, N344, N478);
buf BUF1 (N509, N498);
buf BUF1 (N510, N468);
endmodule