// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N3014,N3013,N3002,N3016,N3012,N3008,N3015,N3017,N3011,N3018;

xor XOR2 (N19, N3, N17);
nand NAND4 (N20, N9, N17, N13, N3);
and AND2 (N21, N11, N9);
not NOT1 (N22, N1);
and AND2 (N23, N22, N10);
nand NAND3 (N24, N22, N20, N8);
xor XOR2 (N25, N19, N24);
and AND4 (N26, N1, N12, N24, N1);
xor XOR2 (N27, N21, N24);
nor NOR4 (N28, N18, N20, N26, N1);
nor NOR4 (N29, N15, N14, N26, N12);
nand NAND4 (N30, N2, N7, N15, N4);
not NOT1 (N31, N7);
xor XOR2 (N32, N24, N15);
xor XOR2 (N33, N2, N18);
nor NOR3 (N34, N32, N13, N18);
and AND4 (N35, N2, N31, N24, N25);
and AND2 (N36, N28, N18);
or OR4 (N37, N12, N36, N20, N18);
or OR4 (N38, N23, N20, N24, N36);
nand NAND4 (N39, N8, N37, N33, N21);
buf BUF1 (N40, N19);
xor XOR2 (N41, N7, N28);
buf BUF1 (N42, N34);
nor NOR2 (N43, N23, N25);
and AND4 (N44, N29, N8, N37, N9);
xor XOR2 (N45, N43, N36);
or OR4 (N46, N27, N5, N45, N28);
not NOT1 (N47, N46);
nand NAND2 (N48, N19, N27);
and AND2 (N49, N47, N27);
xor XOR2 (N50, N38, N43);
xor XOR2 (N51, N50, N31);
xor XOR2 (N52, N39, N16);
xor XOR2 (N53, N35, N9);
buf BUF1 (N54, N52);
xor XOR2 (N55, N42, N27);
buf BUF1 (N56, N49);
and AND3 (N57, N54, N9, N44);
nand NAND3 (N58, N8, N7, N25);
not NOT1 (N59, N41);
buf BUF1 (N60, N51);
nor NOR2 (N61, N60, N15);
xor XOR2 (N62, N56, N61);
buf BUF1 (N63, N12);
nor NOR4 (N64, N57, N59, N32, N8);
buf BUF1 (N65, N26);
buf BUF1 (N66, N30);
buf BUF1 (N67, N64);
or OR2 (N68, N67, N3);
not NOT1 (N69, N65);
not NOT1 (N70, N55);
nor NOR4 (N71, N68, N47, N40, N68);
not NOT1 (N72, N24);
and AND2 (N73, N63, N2);
nand NAND3 (N74, N66, N64, N16);
xor XOR2 (N75, N72, N4);
xor XOR2 (N76, N48, N2);
not NOT1 (N77, N58);
nand NAND2 (N78, N71, N41);
or OR4 (N79, N76, N69, N60, N38);
xor XOR2 (N80, N50, N9);
not NOT1 (N81, N70);
xor XOR2 (N82, N74, N75);
xor XOR2 (N83, N78, N35);
xor XOR2 (N84, N48, N9);
buf BUF1 (N85, N82);
not NOT1 (N86, N84);
or OR2 (N87, N86, N72);
xor XOR2 (N88, N79, N49);
not NOT1 (N89, N62);
or OR2 (N90, N85, N36);
xor XOR2 (N91, N87, N30);
and AND4 (N92, N73, N88, N29, N19);
xor XOR2 (N93, N65, N46);
xor XOR2 (N94, N81, N46);
nor NOR3 (N95, N77, N85, N49);
or OR3 (N96, N90, N72, N67);
not NOT1 (N97, N95);
not NOT1 (N98, N91);
buf BUF1 (N99, N53);
not NOT1 (N100, N98);
buf BUF1 (N101, N97);
xor XOR2 (N102, N89, N48);
xor XOR2 (N103, N101, N49);
xor XOR2 (N104, N93, N14);
nor NOR4 (N105, N94, N21, N52, N52);
or OR3 (N106, N103, N3, N49);
and AND3 (N107, N99, N91, N36);
xor XOR2 (N108, N106, N28);
not NOT1 (N109, N102);
xor XOR2 (N110, N109, N72);
nor NOR2 (N111, N83, N70);
or OR3 (N112, N100, N73, N97);
or OR4 (N113, N110, N74, N98, N94);
nand NAND4 (N114, N107, N104, N5, N99);
not NOT1 (N115, N24);
not NOT1 (N116, N105);
nor NOR2 (N117, N113, N34);
not NOT1 (N118, N115);
nor NOR4 (N119, N114, N61, N29, N25);
buf BUF1 (N120, N112);
xor XOR2 (N121, N111, N41);
nand NAND3 (N122, N96, N4, N30);
or OR4 (N123, N117, N1, N85, N92);
nor NOR3 (N124, N70, N94, N31);
nand NAND4 (N125, N118, N107, N21, N29);
buf BUF1 (N126, N80);
and AND2 (N127, N120, N50);
nand NAND2 (N128, N126, N99);
xor XOR2 (N129, N123, N6);
xor XOR2 (N130, N125, N65);
or OR4 (N131, N119, N19, N46, N22);
or OR2 (N132, N122, N88);
and AND4 (N133, N127, N72, N67, N123);
and AND4 (N134, N124, N84, N21, N67);
xor XOR2 (N135, N108, N43);
or OR4 (N136, N129, N12, N55, N61);
buf BUF1 (N137, N132);
and AND3 (N138, N133, N112, N40);
and AND2 (N139, N138, N33);
nor NOR4 (N140, N116, N39, N10, N11);
buf BUF1 (N141, N131);
or OR4 (N142, N135, N4, N67, N6);
and AND3 (N143, N140, N23, N91);
and AND4 (N144, N134, N70, N26, N120);
xor XOR2 (N145, N136, N13);
nor NOR4 (N146, N130, N109, N49, N140);
nor NOR4 (N147, N142, N15, N4, N36);
nand NAND2 (N148, N145, N25);
nor NOR3 (N149, N146, N70, N141);
nand NAND2 (N150, N112, N95);
or OR2 (N151, N128, N4);
not NOT1 (N152, N144);
and AND2 (N153, N121, N3);
nand NAND4 (N154, N150, N142, N140, N35);
xor XOR2 (N155, N154, N50);
not NOT1 (N156, N137);
nand NAND3 (N157, N155, N73, N109);
not NOT1 (N158, N139);
or OR4 (N159, N149, N39, N118, N136);
nand NAND2 (N160, N159, N146);
nand NAND2 (N161, N158, N9);
xor XOR2 (N162, N156, N18);
buf BUF1 (N163, N162);
nor NOR3 (N164, N143, N142, N6);
xor XOR2 (N165, N147, N57);
nor NOR3 (N166, N164, N104, N86);
and AND3 (N167, N151, N94, N166);
nor NOR4 (N168, N134, N131, N45, N99);
xor XOR2 (N169, N153, N10);
not NOT1 (N170, N160);
not NOT1 (N171, N157);
not NOT1 (N172, N171);
nor NOR4 (N173, N169, N74, N37, N99);
buf BUF1 (N174, N168);
nor NOR4 (N175, N173, N40, N128, N158);
and AND2 (N176, N175, N84);
nor NOR3 (N177, N176, N32, N101);
or OR4 (N178, N174, N99, N120, N117);
or OR4 (N179, N165, N46, N87, N136);
not NOT1 (N180, N161);
nor NOR3 (N181, N167, N171, N37);
nand NAND2 (N182, N148, N180);
not NOT1 (N183, N171);
xor XOR2 (N184, N170, N159);
and AND3 (N185, N179, N176, N115);
buf BUF1 (N186, N185);
nor NOR3 (N187, N182, N145, N10);
and AND2 (N188, N181, N68);
not NOT1 (N189, N163);
buf BUF1 (N190, N184);
and AND2 (N191, N172, N113);
nor NOR4 (N192, N152, N21, N13, N16);
and AND4 (N193, N191, N28, N91, N145);
or OR2 (N194, N186, N43);
not NOT1 (N195, N192);
or OR3 (N196, N178, N1, N139);
nand NAND3 (N197, N183, N98, N42);
and AND3 (N198, N196, N197, N15);
or OR3 (N199, N14, N144, N60);
or OR4 (N200, N199, N61, N194, N14);
nand NAND3 (N201, N47, N148, N17);
nand NAND4 (N202, N193, N71, N112, N152);
xor XOR2 (N203, N201, N38);
and AND2 (N204, N195, N151);
nand NAND4 (N205, N203, N132, N130, N204);
buf BUF1 (N206, N190);
or OR3 (N207, N201, N44, N132);
xor XOR2 (N208, N202, N89);
nor NOR2 (N209, N198, N119);
nand NAND2 (N210, N209, N52);
or OR3 (N211, N206, N34, N180);
buf BUF1 (N212, N208);
buf BUF1 (N213, N188);
and AND4 (N214, N177, N201, N86, N58);
buf BUF1 (N215, N214);
not NOT1 (N216, N187);
xor XOR2 (N217, N213, N203);
nand NAND3 (N218, N217, N192, N106);
nor NOR4 (N219, N200, N88, N17, N132);
buf BUF1 (N220, N189);
buf BUF1 (N221, N212);
or OR4 (N222, N221, N120, N52, N19);
nand NAND2 (N223, N220, N151);
or OR2 (N224, N205, N67);
not NOT1 (N225, N223);
buf BUF1 (N226, N215);
buf BUF1 (N227, N219);
xor XOR2 (N228, N210, N117);
and AND2 (N229, N228, N168);
not NOT1 (N230, N207);
not NOT1 (N231, N216);
xor XOR2 (N232, N218, N51);
not NOT1 (N233, N211);
nand NAND3 (N234, N229, N87, N201);
not NOT1 (N235, N225);
not NOT1 (N236, N224);
buf BUF1 (N237, N232);
nor NOR3 (N238, N222, N93, N162);
xor XOR2 (N239, N236, N12);
xor XOR2 (N240, N230, N192);
nand NAND2 (N241, N233, N27);
not NOT1 (N242, N238);
xor XOR2 (N243, N226, N200);
nand NAND2 (N244, N242, N186);
xor XOR2 (N245, N231, N36);
nand NAND4 (N246, N239, N218, N101, N21);
not NOT1 (N247, N234);
and AND2 (N248, N235, N68);
not NOT1 (N249, N246);
and AND3 (N250, N227, N13, N222);
nor NOR2 (N251, N240, N71);
not NOT1 (N252, N237);
nor NOR2 (N253, N248, N81);
and AND3 (N254, N253, N54, N11);
nand NAND3 (N255, N245, N148, N120);
nor NOR3 (N256, N250, N35, N72);
nor NOR2 (N257, N256, N225);
xor XOR2 (N258, N252, N14);
not NOT1 (N259, N244);
and AND4 (N260, N254, N39, N243, N109);
nand NAND4 (N261, N65, N87, N50, N41);
nand NAND3 (N262, N251, N10, N62);
buf BUF1 (N263, N260);
and AND2 (N264, N241, N171);
nor NOR4 (N265, N247, N136, N231, N204);
nor NOR3 (N266, N258, N66, N112);
nand NAND2 (N267, N261, N117);
nor NOR4 (N268, N267, N51, N118, N168);
and AND3 (N269, N266, N109, N73);
or OR3 (N270, N269, N131, N255);
not NOT1 (N271, N115);
buf BUF1 (N272, N268);
not NOT1 (N273, N271);
or OR4 (N274, N264, N115, N131, N136);
not NOT1 (N275, N259);
and AND3 (N276, N274, N31, N252);
xor XOR2 (N277, N275, N132);
nor NOR4 (N278, N277, N187, N94, N60);
or OR3 (N279, N262, N50, N159);
buf BUF1 (N280, N265);
or OR3 (N281, N280, N229, N112);
or OR3 (N282, N278, N271, N57);
or OR4 (N283, N273, N231, N98, N281);
buf BUF1 (N284, N42);
xor XOR2 (N285, N282, N136);
buf BUF1 (N286, N263);
and AND4 (N287, N270, N121, N91, N127);
xor XOR2 (N288, N286, N238);
nor NOR4 (N289, N276, N198, N266, N58);
not NOT1 (N290, N279);
nor NOR2 (N291, N284, N199);
buf BUF1 (N292, N288);
xor XOR2 (N293, N283, N30);
xor XOR2 (N294, N257, N210);
buf BUF1 (N295, N292);
buf BUF1 (N296, N295);
nor NOR2 (N297, N287, N69);
and AND2 (N298, N294, N257);
nand NAND3 (N299, N289, N139, N207);
or OR4 (N300, N249, N221, N132, N49);
buf BUF1 (N301, N293);
and AND2 (N302, N298, N52);
xor XOR2 (N303, N297, N131);
not NOT1 (N304, N303);
nand NAND3 (N305, N300, N20, N137);
nor NOR2 (N306, N272, N61);
and AND3 (N307, N296, N72, N155);
nor NOR3 (N308, N290, N141, N248);
or OR4 (N309, N285, N256, N177, N308);
nor NOR3 (N310, N261, N225, N55);
nor NOR2 (N311, N302, N48);
nand NAND3 (N312, N311, N182, N193);
not NOT1 (N313, N306);
nand NAND2 (N314, N305, N61);
xor XOR2 (N315, N291, N96);
or OR4 (N316, N310, N37, N30, N196);
and AND4 (N317, N301, N139, N136, N56);
or OR3 (N318, N312, N280, N88);
xor XOR2 (N319, N309, N121);
and AND4 (N320, N317, N276, N151, N32);
nand NAND2 (N321, N315, N220);
buf BUF1 (N322, N313);
nand NAND4 (N323, N322, N72, N151, N272);
nand NAND2 (N324, N320, N48);
nor NOR3 (N325, N304, N144, N130);
xor XOR2 (N326, N318, N294);
or OR4 (N327, N324, N309, N261, N275);
or OR2 (N328, N319, N87);
buf BUF1 (N329, N327);
not NOT1 (N330, N328);
nand NAND3 (N331, N323, N164, N259);
xor XOR2 (N332, N329, N40);
nand NAND4 (N333, N314, N258, N332, N84);
and AND3 (N334, N36, N251, N154);
or OR3 (N335, N331, N51, N58);
or OR2 (N336, N316, N273);
and AND3 (N337, N307, N232, N138);
xor XOR2 (N338, N336, N89);
nor NOR2 (N339, N330, N151);
not NOT1 (N340, N321);
not NOT1 (N341, N326);
xor XOR2 (N342, N299, N45);
nor NOR4 (N343, N337, N162, N33, N235);
not NOT1 (N344, N335);
buf BUF1 (N345, N338);
nor NOR4 (N346, N333, N313, N290, N311);
not NOT1 (N347, N339);
nor NOR4 (N348, N344, N257, N66, N94);
nand NAND2 (N349, N347, N291);
and AND3 (N350, N346, N309, N226);
or OR2 (N351, N348, N50);
buf BUF1 (N352, N325);
buf BUF1 (N353, N341);
or OR4 (N354, N342, N227, N269, N66);
xor XOR2 (N355, N345, N230);
nand NAND4 (N356, N351, N10, N125, N180);
nand NAND4 (N357, N354, N338, N344, N247);
nand NAND2 (N358, N356, N133);
nor NOR4 (N359, N353, N138, N51, N245);
buf BUF1 (N360, N343);
nand NAND4 (N361, N359, N253, N46, N285);
not NOT1 (N362, N352);
nor NOR3 (N363, N334, N112, N112);
xor XOR2 (N364, N363, N99);
or OR2 (N365, N350, N42);
not NOT1 (N366, N360);
or OR4 (N367, N358, N239, N225, N236);
xor XOR2 (N368, N349, N285);
nand NAND2 (N369, N340, N340);
xor XOR2 (N370, N368, N169);
xor XOR2 (N371, N365, N128);
and AND4 (N372, N355, N343, N235, N259);
and AND3 (N373, N364, N3, N310);
and AND4 (N374, N369, N147, N61, N335);
and AND2 (N375, N374, N134);
or OR3 (N376, N371, N321, N239);
not NOT1 (N377, N367);
buf BUF1 (N378, N375);
buf BUF1 (N379, N366);
or OR4 (N380, N377, N325, N105, N46);
buf BUF1 (N381, N370);
or OR3 (N382, N373, N135, N240);
nand NAND4 (N383, N379, N172, N273, N4);
or OR4 (N384, N362, N222, N5, N142);
not NOT1 (N385, N361);
nor NOR3 (N386, N376, N331, N19);
xor XOR2 (N387, N357, N318);
nor NOR2 (N388, N384, N30);
buf BUF1 (N389, N386);
or OR3 (N390, N387, N159, N13);
not NOT1 (N391, N382);
not NOT1 (N392, N385);
nand NAND4 (N393, N390, N101, N137, N274);
nand NAND3 (N394, N389, N341, N214);
buf BUF1 (N395, N388);
and AND2 (N396, N380, N297);
nand NAND4 (N397, N396, N136, N223, N89);
xor XOR2 (N398, N372, N105);
nor NOR4 (N399, N394, N273, N51, N253);
nand NAND2 (N400, N383, N383);
nor NOR2 (N401, N393, N320);
xor XOR2 (N402, N392, N209);
nor NOR4 (N403, N401, N243, N58, N126);
nor NOR2 (N404, N381, N371);
xor XOR2 (N405, N398, N320);
nand NAND4 (N406, N400, N196, N285, N225);
nor NOR2 (N407, N399, N273);
nand NAND4 (N408, N405, N24, N272, N159);
nor NOR2 (N409, N378, N389);
buf BUF1 (N410, N402);
xor XOR2 (N411, N397, N325);
nand NAND2 (N412, N406, N270);
nor NOR4 (N413, N408, N287, N34, N350);
or OR4 (N414, N404, N194, N279, N69);
or OR2 (N415, N409, N8);
xor XOR2 (N416, N411, N210);
nor NOR2 (N417, N391, N192);
and AND2 (N418, N417, N146);
nor NOR4 (N419, N395, N333, N328, N145);
not NOT1 (N420, N412);
not NOT1 (N421, N413);
buf BUF1 (N422, N419);
or OR4 (N423, N416, N285, N348, N51);
not NOT1 (N424, N418);
or OR3 (N425, N422, N194, N12);
or OR2 (N426, N407, N137);
xor XOR2 (N427, N425, N133);
and AND2 (N428, N410, N179);
or OR2 (N429, N414, N82);
or OR4 (N430, N428, N429, N423, N167);
xor XOR2 (N431, N195, N63);
nor NOR4 (N432, N255, N66, N176, N115);
not NOT1 (N433, N432);
nand NAND4 (N434, N403, N233, N163, N354);
and AND2 (N435, N420, N423);
and AND3 (N436, N426, N45, N431);
xor XOR2 (N437, N381, N21);
buf BUF1 (N438, N433);
not NOT1 (N439, N434);
nor NOR2 (N440, N424, N392);
not NOT1 (N441, N435);
buf BUF1 (N442, N421);
or OR4 (N443, N438, N320, N227, N123);
xor XOR2 (N444, N442, N259);
not NOT1 (N445, N440);
nor NOR4 (N446, N439, N20, N239, N166);
and AND3 (N447, N436, N335, N47);
not NOT1 (N448, N441);
nand NAND3 (N449, N415, N36, N112);
or OR2 (N450, N444, N253);
nor NOR2 (N451, N427, N168);
buf BUF1 (N452, N449);
and AND3 (N453, N446, N347, N423);
not NOT1 (N454, N452);
nand NAND3 (N455, N445, N294, N295);
nor NOR2 (N456, N450, N237);
buf BUF1 (N457, N453);
or OR3 (N458, N437, N52, N171);
not NOT1 (N459, N443);
xor XOR2 (N460, N448, N6);
buf BUF1 (N461, N460);
nor NOR2 (N462, N461, N109);
xor XOR2 (N463, N459, N450);
nand NAND4 (N464, N457, N358, N291, N243);
and AND2 (N465, N455, N385);
and AND2 (N466, N454, N120);
and AND2 (N467, N465, N328);
and AND3 (N468, N430, N47, N75);
not NOT1 (N469, N468);
or OR2 (N470, N447, N365);
and AND3 (N471, N462, N171, N44);
or OR3 (N472, N470, N267, N469);
nand NAND2 (N473, N391, N102);
not NOT1 (N474, N472);
not NOT1 (N475, N471);
buf BUF1 (N476, N458);
nor NOR3 (N477, N473, N325, N435);
not NOT1 (N478, N467);
or OR4 (N479, N456, N102, N151, N401);
or OR3 (N480, N479, N96, N393);
xor XOR2 (N481, N451, N266);
or OR3 (N482, N480, N1, N324);
not NOT1 (N483, N463);
nand NAND3 (N484, N466, N101, N380);
xor XOR2 (N485, N474, N93);
and AND2 (N486, N482, N134);
nor NOR3 (N487, N478, N260, N115);
or OR2 (N488, N477, N19);
or OR4 (N489, N476, N243, N133, N449);
and AND4 (N490, N487, N233, N440, N157);
and AND2 (N491, N483, N11);
xor XOR2 (N492, N491, N225);
buf BUF1 (N493, N481);
buf BUF1 (N494, N492);
nand NAND4 (N495, N490, N464, N280, N46);
or OR4 (N496, N138, N149, N263, N235);
xor XOR2 (N497, N493, N75);
or OR2 (N498, N485, N36);
not NOT1 (N499, N489);
buf BUF1 (N500, N496);
and AND2 (N501, N497, N413);
or OR3 (N502, N499, N237, N32);
nand NAND2 (N503, N500, N465);
not NOT1 (N504, N503);
buf BUF1 (N505, N498);
or OR4 (N506, N505, N49, N424, N458);
buf BUF1 (N507, N502);
nor NOR3 (N508, N475, N414, N239);
nor NOR3 (N509, N488, N16, N16);
not NOT1 (N510, N501);
nand NAND3 (N511, N509, N85, N135);
buf BUF1 (N512, N508);
xor XOR2 (N513, N512, N359);
not NOT1 (N514, N504);
nand NAND4 (N515, N495, N421, N119, N480);
not NOT1 (N516, N511);
not NOT1 (N517, N515);
nor NOR4 (N518, N486, N301, N382, N102);
nor NOR2 (N519, N514, N495);
not NOT1 (N520, N513);
and AND4 (N521, N510, N74, N238, N221);
buf BUF1 (N522, N519);
nor NOR3 (N523, N520, N374, N112);
buf BUF1 (N524, N522);
nand NAND4 (N525, N506, N433, N309, N369);
nor NOR4 (N526, N517, N508, N124, N7);
and AND4 (N527, N526, N113, N233, N103);
nor NOR4 (N528, N507, N455, N153, N52);
and AND3 (N529, N516, N217, N371);
not NOT1 (N530, N518);
nand NAND3 (N531, N521, N449, N344);
nor NOR3 (N532, N524, N372, N170);
or OR2 (N533, N527, N513);
nand NAND2 (N534, N533, N130);
buf BUF1 (N535, N525);
nor NOR4 (N536, N531, N511, N261, N501);
buf BUF1 (N537, N535);
not NOT1 (N538, N529);
xor XOR2 (N539, N532, N3);
and AND4 (N540, N523, N202, N276, N390);
and AND3 (N541, N540, N378, N209);
buf BUF1 (N542, N530);
and AND4 (N543, N537, N210, N128, N542);
xor XOR2 (N544, N227, N375);
or OR2 (N545, N534, N356);
buf BUF1 (N546, N544);
not NOT1 (N547, N528);
or OR2 (N548, N543, N325);
nand NAND4 (N549, N546, N148, N332, N486);
buf BUF1 (N550, N541);
not NOT1 (N551, N536);
not NOT1 (N552, N539);
not NOT1 (N553, N551);
and AND4 (N554, N548, N118, N327, N33);
nand NAND2 (N555, N547, N80);
nand NAND2 (N556, N554, N408);
not NOT1 (N557, N545);
and AND3 (N558, N484, N42, N83);
not NOT1 (N559, N552);
buf BUF1 (N560, N556);
buf BUF1 (N561, N557);
xor XOR2 (N562, N538, N44);
nor NOR4 (N563, N553, N334, N322, N493);
buf BUF1 (N564, N555);
or OR4 (N565, N549, N170, N121, N214);
nand NAND4 (N566, N560, N85, N293, N368);
nor NOR4 (N567, N561, N106, N187, N239);
or OR3 (N568, N558, N556, N498);
xor XOR2 (N569, N494, N92);
nand NAND2 (N570, N563, N277);
and AND3 (N571, N568, N383, N182);
nor NOR4 (N572, N570, N2, N273, N284);
and AND3 (N573, N571, N55, N135);
nor NOR4 (N574, N550, N567, N265, N197);
nor NOR4 (N575, N371, N382, N155, N136);
nand NAND2 (N576, N565, N161);
nor NOR2 (N577, N559, N558);
not NOT1 (N578, N574);
or OR2 (N579, N572, N3);
nor NOR4 (N580, N576, N345, N37, N133);
xor XOR2 (N581, N564, N237);
not NOT1 (N582, N579);
not NOT1 (N583, N577);
not NOT1 (N584, N581);
and AND2 (N585, N578, N237);
buf BUF1 (N586, N569);
buf BUF1 (N587, N580);
or OR2 (N588, N562, N243);
buf BUF1 (N589, N575);
or OR2 (N590, N588, N293);
buf BUF1 (N591, N582);
nand NAND2 (N592, N590, N165);
xor XOR2 (N593, N591, N455);
or OR4 (N594, N587, N437, N416, N378);
not NOT1 (N595, N573);
nand NAND2 (N596, N585, N274);
nand NAND2 (N597, N595, N162);
buf BUF1 (N598, N596);
nand NAND4 (N599, N598, N545, N475, N485);
xor XOR2 (N600, N586, N126);
buf BUF1 (N601, N600);
nor NOR3 (N602, N597, N105, N90);
buf BUF1 (N603, N602);
nand NAND3 (N604, N593, N51, N191);
and AND3 (N605, N592, N421, N503);
xor XOR2 (N606, N566, N331);
xor XOR2 (N607, N603, N528);
buf BUF1 (N608, N599);
and AND2 (N609, N594, N336);
nand NAND3 (N610, N583, N3, N252);
buf BUF1 (N611, N607);
xor XOR2 (N612, N584, N340);
or OR3 (N613, N589, N93, N505);
nor NOR3 (N614, N608, N100, N600);
or OR2 (N615, N609, N439);
nor NOR2 (N616, N610, N376);
and AND4 (N617, N612, N146, N533, N161);
nand NAND4 (N618, N611, N29, N188, N424);
or OR4 (N619, N614, N102, N145, N384);
or OR3 (N620, N604, N553, N239);
nand NAND3 (N621, N601, N565, N272);
nand NAND3 (N622, N619, N427, N334);
nor NOR4 (N623, N617, N269, N290, N585);
or OR4 (N624, N616, N71, N172, N496);
or OR3 (N625, N623, N121, N25);
buf BUF1 (N626, N625);
or OR4 (N627, N613, N241, N373, N210);
nor NOR4 (N628, N627, N80, N483, N463);
not NOT1 (N629, N626);
nor NOR3 (N630, N605, N490, N462);
not NOT1 (N631, N630);
xor XOR2 (N632, N629, N222);
and AND4 (N633, N615, N418, N335, N105);
nor NOR3 (N634, N621, N530, N63);
or OR3 (N635, N628, N347, N270);
nand NAND3 (N636, N632, N281, N375);
xor XOR2 (N637, N635, N630);
buf BUF1 (N638, N633);
or OR3 (N639, N620, N547, N381);
nor NOR2 (N640, N624, N134);
or OR3 (N641, N618, N555, N344);
and AND3 (N642, N606, N284, N491);
buf BUF1 (N643, N634);
nand NAND3 (N644, N642, N354, N379);
or OR3 (N645, N640, N396, N97);
not NOT1 (N646, N622);
buf BUF1 (N647, N641);
buf BUF1 (N648, N631);
or OR4 (N649, N643, N524, N358, N611);
and AND2 (N650, N636, N322);
nor NOR3 (N651, N645, N511, N152);
nand NAND3 (N652, N646, N340, N403);
and AND2 (N653, N650, N628);
and AND4 (N654, N651, N442, N239, N209);
and AND2 (N655, N652, N524);
nor NOR3 (N656, N648, N203, N102);
nor NOR4 (N657, N649, N64, N412, N133);
nor NOR2 (N658, N638, N498);
buf BUF1 (N659, N656);
or OR4 (N660, N637, N238, N652, N99);
xor XOR2 (N661, N654, N621);
buf BUF1 (N662, N660);
not NOT1 (N663, N661);
or OR3 (N664, N662, N253, N90);
xor XOR2 (N665, N663, N324);
not NOT1 (N666, N644);
not NOT1 (N667, N659);
or OR2 (N668, N647, N597);
buf BUF1 (N669, N655);
buf BUF1 (N670, N664);
xor XOR2 (N671, N653, N485);
nor NOR2 (N672, N657, N428);
and AND3 (N673, N670, N427, N367);
xor XOR2 (N674, N671, N492);
and AND2 (N675, N674, N558);
not NOT1 (N676, N675);
and AND3 (N677, N639, N22, N556);
and AND3 (N678, N676, N414, N499);
not NOT1 (N679, N673);
nor NOR3 (N680, N672, N37, N252);
nor NOR4 (N681, N667, N123, N572, N241);
or OR4 (N682, N665, N578, N475, N474);
nand NAND4 (N683, N658, N652, N606, N58);
not NOT1 (N684, N669);
and AND2 (N685, N680, N43);
nor NOR2 (N686, N679, N493);
buf BUF1 (N687, N682);
nor NOR4 (N688, N668, N610, N373, N260);
xor XOR2 (N689, N666, N507);
xor XOR2 (N690, N683, N533);
not NOT1 (N691, N678);
or OR2 (N692, N677, N418);
xor XOR2 (N693, N681, N145);
not NOT1 (N694, N689);
buf BUF1 (N695, N694);
nand NAND3 (N696, N685, N606, N130);
and AND3 (N697, N684, N59, N421);
buf BUF1 (N698, N697);
or OR3 (N699, N696, N682, N689);
and AND4 (N700, N690, N209, N106, N504);
xor XOR2 (N701, N686, N692);
buf BUF1 (N702, N636);
nor NOR2 (N703, N702, N211);
buf BUF1 (N704, N698);
or OR3 (N705, N701, N173, N110);
not NOT1 (N706, N705);
nand NAND2 (N707, N699, N108);
or OR2 (N708, N706, N27);
nor NOR4 (N709, N708, N54, N378, N685);
and AND3 (N710, N687, N624, N687);
nor NOR3 (N711, N695, N58, N42);
nand NAND2 (N712, N700, N698);
buf BUF1 (N713, N710);
and AND3 (N714, N709, N384, N238);
not NOT1 (N715, N713);
and AND4 (N716, N714, N605, N47, N244);
xor XOR2 (N717, N712, N291);
nor NOR2 (N718, N717, N490);
nand NAND2 (N719, N693, N470);
nand NAND4 (N720, N691, N124, N413, N81);
and AND2 (N721, N711, N335);
nor NOR4 (N722, N721, N697, N460, N464);
nor NOR4 (N723, N718, N163, N586, N427);
nor NOR3 (N724, N719, N429, N652);
xor XOR2 (N725, N723, N629);
nand NAND4 (N726, N722, N538, N418, N393);
and AND2 (N727, N704, N8);
nor NOR3 (N728, N724, N614, N22);
nand NAND4 (N729, N688, N556, N518, N718);
buf BUF1 (N730, N728);
nor NOR3 (N731, N729, N16, N57);
nand NAND4 (N732, N730, N438, N78, N341);
not NOT1 (N733, N725);
buf BUF1 (N734, N707);
and AND2 (N735, N727, N304);
nand NAND3 (N736, N734, N640, N256);
not NOT1 (N737, N715);
xor XOR2 (N738, N726, N255);
or OR3 (N739, N716, N705, N679);
not NOT1 (N740, N736);
nor NOR4 (N741, N703, N604, N735, N267);
and AND2 (N742, N636, N591);
and AND2 (N743, N732, N686);
nand NAND3 (N744, N731, N713, N496);
nor NOR3 (N745, N740, N249, N620);
nand NAND2 (N746, N720, N423);
nor NOR2 (N747, N743, N325);
nand NAND4 (N748, N733, N64, N236, N346);
or OR2 (N749, N741, N471);
nand NAND2 (N750, N749, N415);
buf BUF1 (N751, N738);
or OR3 (N752, N747, N401, N51);
nand NAND4 (N753, N739, N532, N216, N641);
or OR2 (N754, N746, N554);
or OR2 (N755, N742, N58);
and AND2 (N756, N748, N465);
or OR2 (N757, N753, N544);
buf BUF1 (N758, N755);
or OR2 (N759, N750, N545);
not NOT1 (N760, N745);
buf BUF1 (N761, N752);
not NOT1 (N762, N761);
or OR3 (N763, N756, N621, N471);
xor XOR2 (N764, N757, N142);
or OR2 (N765, N764, N440);
not NOT1 (N766, N758);
xor XOR2 (N767, N744, N699);
xor XOR2 (N768, N767, N474);
and AND3 (N769, N765, N731, N330);
buf BUF1 (N770, N768);
xor XOR2 (N771, N737, N589);
xor XOR2 (N772, N763, N210);
nor NOR3 (N773, N754, N34, N463);
xor XOR2 (N774, N771, N35);
buf BUF1 (N775, N774);
not NOT1 (N776, N769);
or OR2 (N777, N775, N445);
or OR4 (N778, N759, N166, N36, N588);
buf BUF1 (N779, N778);
xor XOR2 (N780, N751, N192);
buf BUF1 (N781, N780);
xor XOR2 (N782, N773, N310);
not NOT1 (N783, N770);
xor XOR2 (N784, N760, N763);
and AND2 (N785, N784, N382);
xor XOR2 (N786, N785, N109);
or OR3 (N787, N781, N208, N166);
xor XOR2 (N788, N787, N763);
not NOT1 (N789, N786);
not NOT1 (N790, N762);
not NOT1 (N791, N766);
nor NOR2 (N792, N791, N41);
and AND3 (N793, N782, N303, N536);
nor NOR4 (N794, N789, N299, N168, N533);
buf BUF1 (N795, N779);
and AND2 (N796, N794, N665);
not NOT1 (N797, N777);
nor NOR4 (N798, N790, N388, N256, N399);
nand NAND2 (N799, N795, N367);
and AND2 (N800, N798, N771);
not NOT1 (N801, N796);
not NOT1 (N802, N788);
nor NOR2 (N803, N802, N794);
buf BUF1 (N804, N792);
not NOT1 (N805, N797);
nand NAND4 (N806, N800, N219, N359, N581);
buf BUF1 (N807, N783);
buf BUF1 (N808, N801);
and AND2 (N809, N793, N257);
and AND4 (N810, N805, N715, N309, N426);
xor XOR2 (N811, N810, N354);
buf BUF1 (N812, N799);
nand NAND2 (N813, N812, N75);
or OR2 (N814, N803, N262);
buf BUF1 (N815, N814);
nor NOR4 (N816, N806, N156, N211, N20);
or OR2 (N817, N808, N807);
and AND2 (N818, N216, N61);
nand NAND4 (N819, N772, N171, N586, N729);
nand NAND2 (N820, N818, N187);
or OR2 (N821, N816, N814);
and AND4 (N822, N820, N427, N782, N8);
and AND3 (N823, N809, N449, N565);
buf BUF1 (N824, N821);
not NOT1 (N825, N813);
nor NOR3 (N826, N824, N707, N384);
and AND2 (N827, N811, N170);
xor XOR2 (N828, N817, N738);
nor NOR3 (N829, N823, N283, N761);
not NOT1 (N830, N819);
or OR3 (N831, N804, N37, N310);
not NOT1 (N832, N822);
and AND3 (N833, N827, N13, N481);
xor XOR2 (N834, N830, N315);
xor XOR2 (N835, N834, N711);
buf BUF1 (N836, N833);
buf BUF1 (N837, N835);
buf BUF1 (N838, N826);
and AND2 (N839, N836, N718);
xor XOR2 (N840, N825, N779);
not NOT1 (N841, N828);
not NOT1 (N842, N832);
not NOT1 (N843, N841);
or OR2 (N844, N831, N600);
or OR3 (N845, N776, N291, N430);
nand NAND2 (N846, N837, N430);
buf BUF1 (N847, N815);
xor XOR2 (N848, N844, N381);
nand NAND2 (N849, N848, N735);
or OR3 (N850, N829, N810, N492);
buf BUF1 (N851, N847);
nand NAND4 (N852, N843, N56, N557, N44);
and AND3 (N853, N838, N617, N645);
not NOT1 (N854, N853);
or OR4 (N855, N851, N634, N737, N695);
or OR4 (N856, N839, N764, N853, N502);
buf BUF1 (N857, N842);
not NOT1 (N858, N849);
buf BUF1 (N859, N857);
xor XOR2 (N860, N852, N363);
buf BUF1 (N861, N858);
and AND2 (N862, N845, N315);
not NOT1 (N863, N860);
and AND4 (N864, N854, N198, N353, N238);
buf BUF1 (N865, N859);
buf BUF1 (N866, N850);
xor XOR2 (N867, N865, N244);
and AND2 (N868, N864, N75);
not NOT1 (N869, N868);
or OR4 (N870, N846, N26, N327, N561);
nand NAND2 (N871, N870, N713);
buf BUF1 (N872, N856);
nand NAND2 (N873, N862, N441);
buf BUF1 (N874, N869);
or OR2 (N875, N867, N790);
nor NOR4 (N876, N840, N383, N136, N601);
not NOT1 (N877, N875);
nor NOR2 (N878, N866, N615);
xor XOR2 (N879, N878, N398);
xor XOR2 (N880, N877, N34);
nand NAND4 (N881, N863, N679, N26, N250);
and AND3 (N882, N874, N840, N167);
nand NAND3 (N883, N855, N264, N560);
not NOT1 (N884, N879);
and AND2 (N885, N880, N560);
xor XOR2 (N886, N882, N225);
xor XOR2 (N887, N885, N711);
nor NOR2 (N888, N876, N754);
nor NOR3 (N889, N873, N791, N21);
nand NAND3 (N890, N861, N501, N232);
nor NOR3 (N891, N884, N231, N156);
buf BUF1 (N892, N889);
and AND4 (N893, N890, N316, N655, N461);
not NOT1 (N894, N881);
nor NOR4 (N895, N888, N590, N211, N143);
nand NAND4 (N896, N872, N891, N286, N799);
nand NAND3 (N897, N189, N320, N56);
buf BUF1 (N898, N892);
buf BUF1 (N899, N893);
nor NOR3 (N900, N894, N651, N743);
not NOT1 (N901, N886);
xor XOR2 (N902, N900, N882);
and AND4 (N903, N871, N714, N27, N360);
nand NAND4 (N904, N899, N269, N142, N68);
xor XOR2 (N905, N883, N426);
xor XOR2 (N906, N905, N326);
xor XOR2 (N907, N904, N735);
nor NOR4 (N908, N895, N600, N156, N607);
not NOT1 (N909, N901);
nor NOR2 (N910, N896, N539);
xor XOR2 (N911, N910, N327);
and AND3 (N912, N908, N869, N491);
and AND2 (N913, N902, N288);
buf BUF1 (N914, N898);
and AND3 (N915, N913, N663, N95);
and AND4 (N916, N912, N422, N172, N853);
not NOT1 (N917, N903);
not NOT1 (N918, N915);
not NOT1 (N919, N887);
or OR2 (N920, N916, N653);
nor NOR2 (N921, N917, N554);
nand NAND3 (N922, N911, N752, N256);
or OR3 (N923, N909, N861, N779);
xor XOR2 (N924, N918, N577);
and AND3 (N925, N914, N495, N37);
buf BUF1 (N926, N920);
nand NAND4 (N927, N924, N553, N681, N182);
nand NAND4 (N928, N926, N826, N417, N912);
buf BUF1 (N929, N907);
buf BUF1 (N930, N897);
and AND2 (N931, N906, N877);
and AND3 (N932, N930, N77, N283);
nor NOR4 (N933, N922, N431, N618, N223);
nand NAND4 (N934, N927, N420, N500, N921);
not NOT1 (N935, N852);
nor NOR3 (N936, N935, N404, N900);
nand NAND4 (N937, N933, N468, N628, N407);
and AND4 (N938, N937, N799, N601, N465);
buf BUF1 (N939, N938);
not NOT1 (N940, N925);
nor NOR3 (N941, N931, N368, N225);
or OR2 (N942, N932, N387);
and AND4 (N943, N928, N532, N493, N734);
nor NOR3 (N944, N942, N518, N366);
nand NAND2 (N945, N923, N192);
not NOT1 (N946, N940);
nor NOR4 (N947, N936, N539, N104, N620);
nand NAND2 (N948, N947, N707);
nor NOR2 (N949, N943, N65);
or OR2 (N950, N919, N534);
nand NAND2 (N951, N949, N443);
xor XOR2 (N952, N950, N17);
and AND3 (N953, N929, N92, N782);
buf BUF1 (N954, N948);
xor XOR2 (N955, N934, N27);
xor XOR2 (N956, N945, N29);
and AND3 (N957, N941, N713, N855);
xor XOR2 (N958, N944, N170);
xor XOR2 (N959, N953, N563);
buf BUF1 (N960, N952);
xor XOR2 (N961, N958, N232);
or OR4 (N962, N957, N523, N343, N595);
nand NAND3 (N963, N951, N682, N596);
nor NOR3 (N964, N962, N792, N955);
xor XOR2 (N965, N125, N628);
or OR4 (N966, N963, N791, N929, N188);
or OR4 (N967, N939, N467, N726, N419);
xor XOR2 (N968, N965, N684);
nand NAND3 (N969, N964, N172, N686);
not NOT1 (N970, N967);
buf BUF1 (N971, N959);
or OR3 (N972, N960, N677, N651);
nand NAND2 (N973, N966, N76);
and AND2 (N974, N970, N610);
xor XOR2 (N975, N974, N459);
nand NAND2 (N976, N956, N834);
nor NOR3 (N977, N976, N145, N400);
nand NAND3 (N978, N971, N149, N608);
xor XOR2 (N979, N975, N432);
not NOT1 (N980, N946);
not NOT1 (N981, N977);
not NOT1 (N982, N954);
buf BUF1 (N983, N980);
nor NOR3 (N984, N969, N414, N546);
buf BUF1 (N985, N978);
buf BUF1 (N986, N983);
nand NAND2 (N987, N961, N709);
nor NOR3 (N988, N984, N755, N215);
xor XOR2 (N989, N988, N203);
and AND4 (N990, N987, N95, N434, N687);
or OR4 (N991, N979, N764, N534, N69);
or OR4 (N992, N982, N398, N406, N405);
xor XOR2 (N993, N986, N760);
not NOT1 (N994, N992);
nor NOR4 (N995, N973, N863, N647, N597);
not NOT1 (N996, N994);
not NOT1 (N997, N991);
nand NAND2 (N998, N981, N748);
xor XOR2 (N999, N995, N871);
xor XOR2 (N1000, N997, N547);
xor XOR2 (N1001, N985, N920);
nand NAND2 (N1002, N972, N920);
and AND4 (N1003, N990, N18, N467, N630);
xor XOR2 (N1004, N1002, N95);
and AND3 (N1005, N989, N571, N266);
buf BUF1 (N1006, N1001);
not NOT1 (N1007, N998);
not NOT1 (N1008, N999);
xor XOR2 (N1009, N1007, N1004);
xor XOR2 (N1010, N664, N825);
xor XOR2 (N1011, N996, N684);
nor NOR3 (N1012, N1010, N480, N624);
not NOT1 (N1013, N1009);
xor XOR2 (N1014, N1000, N793);
buf BUF1 (N1015, N1014);
or OR4 (N1016, N1003, N825, N74, N423);
not NOT1 (N1017, N1011);
nor NOR2 (N1018, N1012, N484);
and AND4 (N1019, N1005, N354, N422, N693);
or OR4 (N1020, N1016, N768, N553, N947);
buf BUF1 (N1021, N1006);
and AND2 (N1022, N1020, N352);
nor NOR4 (N1023, N1019, N637, N846, N950);
or OR3 (N1024, N1021, N461, N304);
nor NOR4 (N1025, N993, N345, N906, N906);
or OR2 (N1026, N1024, N455);
nor NOR4 (N1027, N1023, N261, N539, N228);
and AND4 (N1028, N1013, N223, N406, N898);
nand NAND3 (N1029, N1017, N31, N150);
nor NOR4 (N1030, N1025, N591, N758, N727);
or OR3 (N1031, N1026, N793, N678);
nor NOR2 (N1032, N968, N646);
not NOT1 (N1033, N1015);
xor XOR2 (N1034, N1008, N140);
or OR2 (N1035, N1032, N653);
buf BUF1 (N1036, N1035);
buf BUF1 (N1037, N1029);
or OR3 (N1038, N1031, N345, N774);
or OR2 (N1039, N1037, N976);
xor XOR2 (N1040, N1033, N1003);
nor NOR3 (N1041, N1039, N781, N687);
buf BUF1 (N1042, N1036);
buf BUF1 (N1043, N1040);
or OR3 (N1044, N1038, N54, N580);
and AND4 (N1045, N1030, N229, N719, N746);
xor XOR2 (N1046, N1041, N765);
nand NAND3 (N1047, N1044, N130, N456);
not NOT1 (N1048, N1022);
nor NOR4 (N1049, N1048, N316, N817, N384);
not NOT1 (N1050, N1028);
or OR4 (N1051, N1027, N430, N333, N9);
nand NAND3 (N1052, N1043, N631, N913);
not NOT1 (N1053, N1034);
and AND2 (N1054, N1045, N651);
buf BUF1 (N1055, N1042);
or OR2 (N1056, N1052, N1050);
and AND3 (N1057, N800, N394, N574);
xor XOR2 (N1058, N1057, N417);
nor NOR2 (N1059, N1054, N1026);
buf BUF1 (N1060, N1049);
and AND2 (N1061, N1056, N163);
and AND3 (N1062, N1055, N388, N434);
or OR3 (N1063, N1060, N799, N291);
buf BUF1 (N1064, N1053);
or OR2 (N1065, N1062, N744);
xor XOR2 (N1066, N1046, N888);
nand NAND2 (N1067, N1051, N751);
nor NOR4 (N1068, N1047, N240, N59, N818);
nand NAND3 (N1069, N1018, N426, N440);
or OR2 (N1070, N1058, N3);
and AND3 (N1071, N1059, N127, N612);
and AND3 (N1072, N1068, N343, N1047);
xor XOR2 (N1073, N1067, N305);
nand NAND2 (N1074, N1066, N1008);
and AND3 (N1075, N1070, N554, N502);
nor NOR3 (N1076, N1074, N866, N674);
buf BUF1 (N1077, N1069);
not NOT1 (N1078, N1063);
nor NOR4 (N1079, N1076, N449, N164, N783);
not NOT1 (N1080, N1072);
or OR4 (N1081, N1065, N178, N941, N695);
buf BUF1 (N1082, N1078);
and AND4 (N1083, N1082, N529, N421, N58);
buf BUF1 (N1084, N1073);
buf BUF1 (N1085, N1081);
buf BUF1 (N1086, N1080);
xor XOR2 (N1087, N1075, N188);
buf BUF1 (N1088, N1085);
nand NAND2 (N1089, N1079, N455);
or OR2 (N1090, N1089, N191);
nor NOR3 (N1091, N1083, N723, N532);
not NOT1 (N1092, N1091);
xor XOR2 (N1093, N1086, N136);
nand NAND2 (N1094, N1090, N440);
xor XOR2 (N1095, N1084, N745);
not NOT1 (N1096, N1088);
nand NAND2 (N1097, N1061, N910);
buf BUF1 (N1098, N1071);
nor NOR2 (N1099, N1077, N1093);
xor XOR2 (N1100, N840, N1068);
not NOT1 (N1101, N1098);
nand NAND2 (N1102, N1099, N1028);
not NOT1 (N1103, N1102);
xor XOR2 (N1104, N1087, N368);
and AND3 (N1105, N1097, N560, N258);
or OR4 (N1106, N1096, N623, N256, N736);
buf BUF1 (N1107, N1094);
or OR3 (N1108, N1103, N318, N970);
nor NOR3 (N1109, N1105, N827, N555);
and AND4 (N1110, N1106, N531, N385, N1071);
and AND3 (N1111, N1108, N544, N637);
or OR2 (N1112, N1095, N638);
xor XOR2 (N1113, N1111, N576);
or OR2 (N1114, N1107, N1051);
not NOT1 (N1115, N1064);
nor NOR3 (N1116, N1110, N204, N19);
nor NOR2 (N1117, N1104, N1063);
and AND2 (N1118, N1115, N453);
not NOT1 (N1119, N1117);
not NOT1 (N1120, N1109);
or OR3 (N1121, N1100, N413, N521);
buf BUF1 (N1122, N1120);
buf BUF1 (N1123, N1092);
nand NAND2 (N1124, N1119, N37);
nor NOR2 (N1125, N1116, N273);
or OR2 (N1126, N1123, N540);
buf BUF1 (N1127, N1121);
not NOT1 (N1128, N1114);
or OR4 (N1129, N1127, N434, N710, N102);
not NOT1 (N1130, N1129);
and AND4 (N1131, N1130, N316, N1024, N182);
nand NAND3 (N1132, N1124, N410, N950);
nand NAND3 (N1133, N1112, N739, N1021);
or OR3 (N1134, N1101, N638, N1082);
nand NAND3 (N1135, N1125, N946, N845);
nor NOR2 (N1136, N1118, N1126);
nand NAND3 (N1137, N103, N561, N1075);
nor NOR4 (N1138, N1122, N1029, N1093, N265);
nand NAND4 (N1139, N1135, N540, N480, N137);
xor XOR2 (N1140, N1133, N240);
nand NAND4 (N1141, N1139, N328, N106, N805);
or OR3 (N1142, N1134, N249, N205);
or OR4 (N1143, N1136, N15, N424, N343);
xor XOR2 (N1144, N1138, N841);
nand NAND3 (N1145, N1143, N592, N871);
buf BUF1 (N1146, N1142);
or OR3 (N1147, N1113, N57, N1052);
xor XOR2 (N1148, N1132, N759);
buf BUF1 (N1149, N1144);
nor NOR3 (N1150, N1146, N340, N877);
and AND4 (N1151, N1131, N674, N290, N349);
xor XOR2 (N1152, N1140, N152);
or OR3 (N1153, N1147, N516, N378);
and AND4 (N1154, N1137, N1025, N214, N867);
and AND4 (N1155, N1149, N801, N837, N694);
or OR3 (N1156, N1150, N1003, N409);
nor NOR2 (N1157, N1155, N981);
and AND2 (N1158, N1156, N240);
not NOT1 (N1159, N1158);
xor XOR2 (N1160, N1154, N338);
or OR4 (N1161, N1159, N104, N460, N352);
nor NOR3 (N1162, N1148, N47, N192);
or OR2 (N1163, N1141, N677);
not NOT1 (N1164, N1163);
buf BUF1 (N1165, N1160);
buf BUF1 (N1166, N1153);
nand NAND3 (N1167, N1164, N1165, N419);
and AND3 (N1168, N717, N830, N1035);
nand NAND2 (N1169, N1151, N246);
xor XOR2 (N1170, N1161, N331);
and AND4 (N1171, N1170, N784, N201, N286);
and AND4 (N1172, N1145, N524, N473, N1141);
nand NAND3 (N1173, N1168, N20, N755);
nand NAND3 (N1174, N1128, N1089, N339);
and AND3 (N1175, N1171, N16, N1147);
and AND3 (N1176, N1167, N408, N213);
nor NOR2 (N1177, N1166, N240);
or OR4 (N1178, N1177, N546, N1018, N364);
nor NOR2 (N1179, N1178, N1121);
xor XOR2 (N1180, N1176, N246);
and AND4 (N1181, N1152, N603, N1163, N1086);
and AND4 (N1182, N1172, N89, N1025, N136);
nand NAND3 (N1183, N1157, N1045, N329);
nand NAND4 (N1184, N1182, N376, N1125, N1066);
buf BUF1 (N1185, N1183);
not NOT1 (N1186, N1179);
not NOT1 (N1187, N1169);
not NOT1 (N1188, N1181);
nand NAND3 (N1189, N1186, N28, N2);
nand NAND2 (N1190, N1187, N577);
or OR3 (N1191, N1184, N408, N41);
not NOT1 (N1192, N1185);
or OR2 (N1193, N1173, N593);
not NOT1 (N1194, N1191);
xor XOR2 (N1195, N1194, N1027);
buf BUF1 (N1196, N1162);
nand NAND2 (N1197, N1195, N385);
nand NAND4 (N1198, N1180, N841, N585, N895);
and AND4 (N1199, N1189, N536, N272, N4);
nor NOR2 (N1200, N1192, N830);
nor NOR2 (N1201, N1200, N1138);
buf BUF1 (N1202, N1174);
buf BUF1 (N1203, N1201);
not NOT1 (N1204, N1203);
not NOT1 (N1205, N1188);
xor XOR2 (N1206, N1190, N824);
nand NAND2 (N1207, N1175, N1017);
buf BUF1 (N1208, N1207);
not NOT1 (N1209, N1202);
nor NOR2 (N1210, N1209, N593);
or OR2 (N1211, N1199, N16);
and AND3 (N1212, N1211, N453, N987);
not NOT1 (N1213, N1206);
and AND4 (N1214, N1196, N729, N72, N1201);
and AND4 (N1215, N1213, N162, N292, N468);
nor NOR2 (N1216, N1212, N707);
and AND2 (N1217, N1198, N515);
xor XOR2 (N1218, N1216, N1107);
nand NAND2 (N1219, N1218, N72);
nand NAND2 (N1220, N1208, N1159);
not NOT1 (N1221, N1210);
buf BUF1 (N1222, N1220);
and AND2 (N1223, N1217, N1021);
buf BUF1 (N1224, N1223);
xor XOR2 (N1225, N1205, N730);
and AND2 (N1226, N1221, N733);
nand NAND3 (N1227, N1197, N744, N651);
or OR2 (N1228, N1224, N1088);
buf BUF1 (N1229, N1214);
xor XOR2 (N1230, N1227, N6);
xor XOR2 (N1231, N1193, N253);
or OR4 (N1232, N1229, N389, N279, N71);
nand NAND2 (N1233, N1225, N1095);
nand NAND3 (N1234, N1215, N492, N246);
and AND4 (N1235, N1231, N454, N653, N1173);
and AND2 (N1236, N1234, N1183);
or OR4 (N1237, N1230, N491, N776, N115);
nor NOR2 (N1238, N1237, N1183);
not NOT1 (N1239, N1235);
nand NAND4 (N1240, N1236, N761, N1008, N125);
buf BUF1 (N1241, N1228);
nand NAND3 (N1242, N1222, N92, N750);
xor XOR2 (N1243, N1204, N105);
xor XOR2 (N1244, N1219, N775);
not NOT1 (N1245, N1244);
not NOT1 (N1246, N1226);
and AND3 (N1247, N1232, N233, N1131);
nor NOR4 (N1248, N1238, N828, N1180, N1196);
nand NAND4 (N1249, N1233, N188, N710, N587);
buf BUF1 (N1250, N1249);
nor NOR2 (N1251, N1250, N490);
nor NOR2 (N1252, N1242, N337);
or OR2 (N1253, N1246, N1200);
nand NAND2 (N1254, N1248, N451);
nor NOR3 (N1255, N1243, N73, N228);
buf BUF1 (N1256, N1239);
buf BUF1 (N1257, N1241);
and AND4 (N1258, N1251, N309, N559, N654);
xor XOR2 (N1259, N1254, N767);
nor NOR4 (N1260, N1247, N305, N481, N1108);
not NOT1 (N1261, N1245);
or OR4 (N1262, N1259, N926, N1164, N608);
xor XOR2 (N1263, N1253, N751);
buf BUF1 (N1264, N1256);
and AND3 (N1265, N1262, N1215, N34);
and AND2 (N1266, N1261, N554);
buf BUF1 (N1267, N1260);
xor XOR2 (N1268, N1255, N272);
nor NOR2 (N1269, N1240, N206);
xor XOR2 (N1270, N1266, N1161);
buf BUF1 (N1271, N1269);
or OR3 (N1272, N1263, N1189, N486);
or OR4 (N1273, N1268, N12, N220, N57);
xor XOR2 (N1274, N1271, N106);
buf BUF1 (N1275, N1274);
or OR2 (N1276, N1270, N1093);
buf BUF1 (N1277, N1272);
nand NAND3 (N1278, N1275, N685, N1150);
nor NOR3 (N1279, N1264, N616, N873);
nand NAND4 (N1280, N1277, N188, N1147, N1062);
and AND3 (N1281, N1280, N213, N1192);
nand NAND3 (N1282, N1279, N1156, N355);
xor XOR2 (N1283, N1273, N496);
or OR3 (N1284, N1283, N625, N1203);
buf BUF1 (N1285, N1278);
not NOT1 (N1286, N1281);
nor NOR4 (N1287, N1257, N173, N1201, N412);
buf BUF1 (N1288, N1258);
xor XOR2 (N1289, N1276, N668);
not NOT1 (N1290, N1287);
nand NAND2 (N1291, N1282, N863);
and AND2 (N1292, N1286, N973);
or OR2 (N1293, N1289, N655);
nor NOR2 (N1294, N1285, N810);
buf BUF1 (N1295, N1288);
xor XOR2 (N1296, N1284, N508);
or OR3 (N1297, N1290, N134, N1077);
buf BUF1 (N1298, N1294);
and AND3 (N1299, N1292, N1208, N216);
xor XOR2 (N1300, N1265, N877);
or OR4 (N1301, N1296, N328, N333, N866);
buf BUF1 (N1302, N1299);
xor XOR2 (N1303, N1267, N1280);
nor NOR2 (N1304, N1297, N576);
nand NAND4 (N1305, N1295, N689, N1126, N1236);
xor XOR2 (N1306, N1300, N142);
xor XOR2 (N1307, N1298, N871);
nor NOR4 (N1308, N1252, N1144, N191, N133);
not NOT1 (N1309, N1308);
buf BUF1 (N1310, N1293);
xor XOR2 (N1311, N1310, N581);
nor NOR3 (N1312, N1305, N803, N705);
buf BUF1 (N1313, N1312);
buf BUF1 (N1314, N1301);
and AND3 (N1315, N1313, N47, N207);
and AND4 (N1316, N1307, N208, N393, N854);
buf BUF1 (N1317, N1291);
xor XOR2 (N1318, N1309, N747);
or OR2 (N1319, N1311, N1250);
xor XOR2 (N1320, N1317, N838);
xor XOR2 (N1321, N1304, N374);
not NOT1 (N1322, N1314);
nor NOR3 (N1323, N1316, N64, N138);
and AND4 (N1324, N1323, N924, N417, N310);
not NOT1 (N1325, N1321);
xor XOR2 (N1326, N1322, N203);
nor NOR3 (N1327, N1318, N1161, N607);
nand NAND4 (N1328, N1320, N508, N1129, N1169);
buf BUF1 (N1329, N1328);
or OR4 (N1330, N1324, N1084, N460, N919);
buf BUF1 (N1331, N1319);
nand NAND3 (N1332, N1303, N240, N68);
buf BUF1 (N1333, N1329);
buf BUF1 (N1334, N1327);
buf BUF1 (N1335, N1332);
nand NAND4 (N1336, N1315, N700, N744, N7);
buf BUF1 (N1337, N1302);
nand NAND4 (N1338, N1325, N352, N1226, N1172);
buf BUF1 (N1339, N1331);
and AND3 (N1340, N1326, N491, N594);
nor NOR2 (N1341, N1338, N1203);
nor NOR2 (N1342, N1335, N1193);
nor NOR4 (N1343, N1330, N202, N1026, N104);
nor NOR4 (N1344, N1336, N1138, N1248, N1104);
xor XOR2 (N1345, N1340, N847);
and AND2 (N1346, N1339, N799);
nor NOR4 (N1347, N1341, N441, N663, N1104);
buf BUF1 (N1348, N1344);
nand NAND4 (N1349, N1346, N902, N740, N234);
nand NAND3 (N1350, N1345, N1128, N1189);
xor XOR2 (N1351, N1347, N798);
nand NAND3 (N1352, N1306, N255, N596);
and AND4 (N1353, N1343, N677, N525, N463);
and AND3 (N1354, N1334, N768, N156);
and AND4 (N1355, N1351, N218, N816, N1329);
buf BUF1 (N1356, N1353);
or OR3 (N1357, N1348, N1064, N866);
nand NAND4 (N1358, N1349, N685, N1333, N1148);
buf BUF1 (N1359, N1016);
or OR3 (N1360, N1342, N434, N1174);
xor XOR2 (N1361, N1352, N943);
or OR4 (N1362, N1350, N950, N610, N779);
and AND4 (N1363, N1362, N431, N1278, N1272);
and AND2 (N1364, N1361, N133);
not NOT1 (N1365, N1358);
nand NAND3 (N1366, N1354, N561, N1335);
or OR2 (N1367, N1360, N387);
and AND4 (N1368, N1337, N142, N1018, N209);
and AND2 (N1369, N1357, N694);
or OR2 (N1370, N1355, N83);
or OR4 (N1371, N1369, N476, N452, N675);
nor NOR4 (N1372, N1364, N880, N298, N1324);
and AND3 (N1373, N1356, N576, N470);
buf BUF1 (N1374, N1371);
xor XOR2 (N1375, N1373, N1020);
nor NOR3 (N1376, N1359, N550, N307);
xor XOR2 (N1377, N1376, N119);
not NOT1 (N1378, N1372);
nor NOR2 (N1379, N1374, N1111);
not NOT1 (N1380, N1365);
or OR4 (N1381, N1370, N1180, N826, N676);
not NOT1 (N1382, N1367);
not NOT1 (N1383, N1363);
not NOT1 (N1384, N1368);
xor XOR2 (N1385, N1383, N587);
nor NOR2 (N1386, N1378, N913);
nand NAND4 (N1387, N1385, N1295, N357, N1092);
buf BUF1 (N1388, N1366);
buf BUF1 (N1389, N1375);
and AND2 (N1390, N1388, N936);
xor XOR2 (N1391, N1390, N1229);
buf BUF1 (N1392, N1389);
and AND3 (N1393, N1379, N335, N593);
nor NOR2 (N1394, N1386, N293);
nor NOR4 (N1395, N1387, N798, N1052, N845);
buf BUF1 (N1396, N1394);
nor NOR3 (N1397, N1392, N624, N1123);
buf BUF1 (N1398, N1381);
xor XOR2 (N1399, N1382, N742);
not NOT1 (N1400, N1384);
buf BUF1 (N1401, N1398);
and AND4 (N1402, N1391, N184, N939, N900);
not NOT1 (N1403, N1401);
xor XOR2 (N1404, N1397, N957);
or OR2 (N1405, N1404, N680);
buf BUF1 (N1406, N1402);
and AND4 (N1407, N1395, N960, N256, N747);
and AND4 (N1408, N1406, N117, N165, N694);
or OR4 (N1409, N1400, N329, N701, N123);
buf BUF1 (N1410, N1399);
or OR2 (N1411, N1396, N910);
not NOT1 (N1412, N1393);
or OR4 (N1413, N1411, N754, N1070, N20);
xor XOR2 (N1414, N1403, N113);
or OR3 (N1415, N1408, N50, N180);
xor XOR2 (N1416, N1412, N1295);
and AND2 (N1417, N1377, N1317);
or OR3 (N1418, N1416, N237, N48);
or OR2 (N1419, N1405, N909);
and AND2 (N1420, N1414, N852);
and AND2 (N1421, N1418, N500);
not NOT1 (N1422, N1419);
and AND2 (N1423, N1421, N1346);
xor XOR2 (N1424, N1409, N394);
xor XOR2 (N1425, N1423, N1366);
nand NAND4 (N1426, N1415, N1223, N1354, N1412);
xor XOR2 (N1427, N1413, N648);
xor XOR2 (N1428, N1380, N1249);
nand NAND4 (N1429, N1424, N386, N731, N1345);
not NOT1 (N1430, N1427);
nor NOR4 (N1431, N1420, N503, N1039, N146);
nand NAND4 (N1432, N1417, N224, N390, N703);
not NOT1 (N1433, N1430);
nor NOR3 (N1434, N1422, N1380, N286);
nor NOR4 (N1435, N1431, N532, N1085, N624);
xor XOR2 (N1436, N1435, N162);
not NOT1 (N1437, N1433);
buf BUF1 (N1438, N1429);
buf BUF1 (N1439, N1434);
not NOT1 (N1440, N1425);
xor XOR2 (N1441, N1439, N165);
buf BUF1 (N1442, N1440);
buf BUF1 (N1443, N1432);
or OR4 (N1444, N1426, N209, N745, N1207);
nor NOR3 (N1445, N1441, N20, N1156);
nor NOR3 (N1446, N1438, N326, N1261);
nor NOR2 (N1447, N1410, N769);
xor XOR2 (N1448, N1445, N1157);
nor NOR3 (N1449, N1436, N1012, N1329);
buf BUF1 (N1450, N1446);
xor XOR2 (N1451, N1448, N385);
or OR4 (N1452, N1437, N803, N84, N257);
xor XOR2 (N1453, N1452, N1346);
nand NAND2 (N1454, N1453, N1167);
nor NOR3 (N1455, N1428, N648, N1297);
nand NAND3 (N1456, N1443, N709, N784);
nand NAND3 (N1457, N1444, N1049, N427);
nand NAND3 (N1458, N1456, N496, N66);
xor XOR2 (N1459, N1450, N732);
nor NOR4 (N1460, N1459, N227, N924, N775);
xor XOR2 (N1461, N1442, N1051);
and AND4 (N1462, N1460, N742, N941, N805);
or OR2 (N1463, N1461, N1452);
xor XOR2 (N1464, N1449, N972);
nor NOR4 (N1465, N1457, N915, N1322, N896);
nand NAND2 (N1466, N1455, N1105);
not NOT1 (N1467, N1465);
not NOT1 (N1468, N1454);
xor XOR2 (N1469, N1407, N1444);
nand NAND3 (N1470, N1463, N903, N1181);
not NOT1 (N1471, N1464);
not NOT1 (N1472, N1468);
not NOT1 (N1473, N1466);
not NOT1 (N1474, N1469);
nand NAND4 (N1475, N1472, N167, N1098, N1264);
and AND3 (N1476, N1451, N679, N1170);
or OR4 (N1477, N1467, N1152, N670, N967);
not NOT1 (N1478, N1473);
not NOT1 (N1479, N1470);
or OR4 (N1480, N1475, N176, N1079, N660);
and AND2 (N1481, N1474, N134);
nand NAND3 (N1482, N1447, N188, N930);
buf BUF1 (N1483, N1479);
nand NAND3 (N1484, N1471, N1057, N1286);
and AND4 (N1485, N1484, N723, N1111, N849);
or OR3 (N1486, N1478, N147, N235);
buf BUF1 (N1487, N1480);
or OR3 (N1488, N1485, N669, N1274);
buf BUF1 (N1489, N1483);
xor XOR2 (N1490, N1458, N505);
nor NOR4 (N1491, N1477, N868, N1056, N324);
buf BUF1 (N1492, N1486);
xor XOR2 (N1493, N1489, N319);
nand NAND3 (N1494, N1488, N988, N386);
buf BUF1 (N1495, N1493);
nand NAND4 (N1496, N1490, N1071, N879, N374);
not NOT1 (N1497, N1482);
and AND3 (N1498, N1476, N667, N530);
not NOT1 (N1499, N1496);
nand NAND3 (N1500, N1487, N837, N939);
nand NAND4 (N1501, N1491, N1015, N502, N716);
and AND3 (N1502, N1492, N684, N561);
buf BUF1 (N1503, N1499);
or OR2 (N1504, N1500, N1221);
or OR3 (N1505, N1497, N1296, N1416);
xor XOR2 (N1506, N1481, N558);
not NOT1 (N1507, N1503);
not NOT1 (N1508, N1504);
or OR2 (N1509, N1462, N454);
not NOT1 (N1510, N1495);
xor XOR2 (N1511, N1506, N885);
nand NAND4 (N1512, N1498, N1119, N411, N708);
xor XOR2 (N1513, N1509, N1311);
and AND3 (N1514, N1505, N1156, N1246);
or OR3 (N1515, N1501, N1231, N858);
and AND3 (N1516, N1513, N897, N442);
nand NAND2 (N1517, N1511, N196);
nor NOR4 (N1518, N1510, N162, N1419, N775);
or OR2 (N1519, N1514, N556);
nor NOR2 (N1520, N1519, N464);
and AND3 (N1521, N1520, N711, N219);
and AND2 (N1522, N1507, N1113);
nor NOR3 (N1523, N1518, N862, N1369);
nor NOR2 (N1524, N1517, N302);
not NOT1 (N1525, N1522);
buf BUF1 (N1526, N1516);
or OR4 (N1527, N1521, N876, N1060, N1146);
not NOT1 (N1528, N1512);
xor XOR2 (N1529, N1523, N82);
and AND3 (N1530, N1526, N1501, N91);
nand NAND2 (N1531, N1502, N226);
buf BUF1 (N1532, N1525);
buf BUF1 (N1533, N1515);
or OR3 (N1534, N1529, N1105, N1365);
nand NAND3 (N1535, N1528, N49, N1067);
not NOT1 (N1536, N1534);
not NOT1 (N1537, N1508);
buf BUF1 (N1538, N1533);
nand NAND2 (N1539, N1532, N669);
and AND3 (N1540, N1535, N1171, N1085);
not NOT1 (N1541, N1539);
xor XOR2 (N1542, N1527, N174);
xor XOR2 (N1543, N1537, N676);
xor XOR2 (N1544, N1524, N1426);
nor NOR3 (N1545, N1542, N1398, N1302);
and AND3 (N1546, N1494, N1210, N562);
and AND4 (N1547, N1538, N199, N281, N1393);
buf BUF1 (N1548, N1544);
nand NAND3 (N1549, N1545, N290, N1057);
not NOT1 (N1550, N1549);
nand NAND2 (N1551, N1550, N1362);
and AND3 (N1552, N1531, N1305, N1200);
or OR2 (N1553, N1552, N748);
nand NAND2 (N1554, N1546, N427);
xor XOR2 (N1555, N1543, N897);
nor NOR2 (N1556, N1547, N855);
or OR3 (N1557, N1548, N1422, N1306);
and AND3 (N1558, N1541, N1020, N641);
not NOT1 (N1559, N1551);
not NOT1 (N1560, N1557);
nand NAND3 (N1561, N1560, N1268, N1014);
and AND3 (N1562, N1540, N649, N569);
and AND3 (N1563, N1530, N1357, N92);
xor XOR2 (N1564, N1562, N1384);
xor XOR2 (N1565, N1536, N878);
nand NAND4 (N1566, N1556, N1295, N1035, N528);
nor NOR4 (N1567, N1566, N630, N171, N736);
xor XOR2 (N1568, N1567, N655);
xor XOR2 (N1569, N1568, N568);
nor NOR4 (N1570, N1554, N1469, N404, N1033);
not NOT1 (N1571, N1553);
xor XOR2 (N1572, N1570, N1016);
and AND3 (N1573, N1564, N1156, N1096);
nor NOR3 (N1574, N1571, N495, N908);
and AND3 (N1575, N1572, N458, N949);
xor XOR2 (N1576, N1558, N303);
buf BUF1 (N1577, N1555);
not NOT1 (N1578, N1559);
not NOT1 (N1579, N1573);
and AND2 (N1580, N1575, N1117);
not NOT1 (N1581, N1577);
or OR4 (N1582, N1565, N688, N1025, N452);
nor NOR3 (N1583, N1576, N773, N259);
not NOT1 (N1584, N1582);
and AND3 (N1585, N1574, N61, N42);
nor NOR2 (N1586, N1580, N902);
not NOT1 (N1587, N1561);
nor NOR4 (N1588, N1587, N916, N1511, N216);
xor XOR2 (N1589, N1579, N573);
or OR2 (N1590, N1589, N1269);
buf BUF1 (N1591, N1583);
not NOT1 (N1592, N1591);
and AND4 (N1593, N1592, N355, N1540, N1156);
or OR2 (N1594, N1581, N191);
xor XOR2 (N1595, N1590, N1389);
nand NAND2 (N1596, N1586, N1389);
nand NAND3 (N1597, N1596, N1282, N2);
not NOT1 (N1598, N1588);
or OR2 (N1599, N1584, N397);
buf BUF1 (N1600, N1563);
buf BUF1 (N1601, N1600);
xor XOR2 (N1602, N1569, N395);
or OR4 (N1603, N1593, N192, N1081, N884);
and AND4 (N1604, N1601, N940, N67, N831);
xor XOR2 (N1605, N1597, N1248);
buf BUF1 (N1606, N1578);
or OR2 (N1607, N1598, N238);
not NOT1 (N1608, N1607);
not NOT1 (N1609, N1608);
and AND3 (N1610, N1594, N886, N153);
or OR3 (N1611, N1603, N242, N357);
not NOT1 (N1612, N1606);
and AND3 (N1613, N1611, N818, N131);
and AND4 (N1614, N1612, N808, N1072, N1336);
not NOT1 (N1615, N1595);
buf BUF1 (N1616, N1614);
nand NAND3 (N1617, N1613, N945, N806);
not NOT1 (N1618, N1616);
and AND2 (N1619, N1605, N941);
nand NAND3 (N1620, N1617, N1553, N1320);
buf BUF1 (N1621, N1619);
and AND3 (N1622, N1610, N1075, N992);
nor NOR4 (N1623, N1585, N836, N620, N14);
buf BUF1 (N1624, N1621);
not NOT1 (N1625, N1604);
xor XOR2 (N1626, N1615, N246);
buf BUF1 (N1627, N1623);
nand NAND4 (N1628, N1627, N674, N120, N1303);
or OR4 (N1629, N1602, N969, N1265, N1579);
not NOT1 (N1630, N1609);
and AND3 (N1631, N1618, N176, N357);
xor XOR2 (N1632, N1622, N1206);
or OR3 (N1633, N1628, N457, N895);
buf BUF1 (N1634, N1620);
buf BUF1 (N1635, N1625);
and AND4 (N1636, N1630, N481, N465, N820);
buf BUF1 (N1637, N1626);
not NOT1 (N1638, N1632);
and AND4 (N1639, N1637, N645, N397, N1586);
or OR4 (N1640, N1624, N819, N152, N836);
buf BUF1 (N1641, N1631);
and AND4 (N1642, N1629, N1137, N1083, N211);
nor NOR3 (N1643, N1638, N571, N701);
nand NAND2 (N1644, N1643, N1103);
nor NOR4 (N1645, N1599, N1624, N627, N24);
or OR2 (N1646, N1642, N1219);
not NOT1 (N1647, N1641);
not NOT1 (N1648, N1640);
nor NOR3 (N1649, N1639, N1596, N935);
and AND2 (N1650, N1647, N54);
and AND3 (N1651, N1634, N1048, N752);
nor NOR3 (N1652, N1651, N296, N1463);
or OR2 (N1653, N1635, N1378);
and AND2 (N1654, N1649, N457);
and AND2 (N1655, N1653, N997);
and AND2 (N1656, N1636, N120);
nand NAND2 (N1657, N1655, N1013);
xor XOR2 (N1658, N1644, N778);
xor XOR2 (N1659, N1656, N736);
or OR2 (N1660, N1658, N1552);
xor XOR2 (N1661, N1652, N775);
xor XOR2 (N1662, N1661, N757);
nor NOR2 (N1663, N1657, N952);
xor XOR2 (N1664, N1646, N21);
xor XOR2 (N1665, N1663, N1165);
xor XOR2 (N1666, N1664, N315);
or OR3 (N1667, N1645, N1510, N1665);
nand NAND3 (N1668, N345, N709, N1531);
nand NAND3 (N1669, N1650, N991, N235);
nand NAND2 (N1670, N1633, N1113);
not NOT1 (N1671, N1670);
nand NAND3 (N1672, N1666, N419, N1654);
nand NAND4 (N1673, N364, N826, N615, N1241);
xor XOR2 (N1674, N1662, N1656);
nor NOR2 (N1675, N1671, N335);
buf BUF1 (N1676, N1659);
or OR2 (N1677, N1676, N848);
not NOT1 (N1678, N1669);
buf BUF1 (N1679, N1648);
and AND2 (N1680, N1667, N112);
and AND3 (N1681, N1674, N363, N819);
or OR4 (N1682, N1668, N1186, N201, N1215);
not NOT1 (N1683, N1677);
nor NOR4 (N1684, N1682, N554, N1086, N60);
nand NAND2 (N1685, N1680, N51);
or OR2 (N1686, N1660, N657);
and AND3 (N1687, N1678, N74, N918);
nand NAND4 (N1688, N1681, N1105, N1221, N878);
nor NOR4 (N1689, N1685, N772, N545, N762);
buf BUF1 (N1690, N1683);
or OR4 (N1691, N1673, N771, N496, N515);
nand NAND4 (N1692, N1689, N380, N924, N711);
and AND4 (N1693, N1692, N1521, N1283, N1130);
xor XOR2 (N1694, N1687, N1339);
and AND3 (N1695, N1690, N313, N1256);
xor XOR2 (N1696, N1691, N818);
not NOT1 (N1697, N1696);
nand NAND2 (N1698, N1694, N330);
not NOT1 (N1699, N1695);
and AND4 (N1700, N1688, N910, N1450, N742);
xor XOR2 (N1701, N1679, N1167);
and AND2 (N1702, N1697, N191);
or OR2 (N1703, N1672, N1119);
nand NAND3 (N1704, N1701, N882, N1643);
buf BUF1 (N1705, N1702);
nor NOR4 (N1706, N1705, N1645, N943, N1271);
nand NAND4 (N1707, N1686, N890, N863, N1643);
or OR4 (N1708, N1693, N41, N212, N113);
not NOT1 (N1709, N1704);
not NOT1 (N1710, N1708);
not NOT1 (N1711, N1707);
or OR2 (N1712, N1700, N1637);
nor NOR4 (N1713, N1699, N1115, N20, N626);
xor XOR2 (N1714, N1712, N463);
nand NAND4 (N1715, N1710, N792, N223, N967);
nor NOR4 (N1716, N1709, N1310, N1708, N303);
and AND2 (N1717, N1711, N1619);
xor XOR2 (N1718, N1716, N1468);
or OR4 (N1719, N1703, N995, N1551, N481);
and AND4 (N1720, N1713, N371, N583, N1159);
nor NOR2 (N1721, N1718, N211);
not NOT1 (N1722, N1675);
or OR3 (N1723, N1722, N312, N1307);
buf BUF1 (N1724, N1684);
xor XOR2 (N1725, N1714, N1328);
or OR2 (N1726, N1721, N340);
nor NOR2 (N1727, N1720, N196);
nand NAND3 (N1728, N1717, N421, N1365);
and AND4 (N1729, N1719, N1398, N1033, N172);
xor XOR2 (N1730, N1724, N1697);
nor NOR2 (N1731, N1698, N491);
not NOT1 (N1732, N1723);
xor XOR2 (N1733, N1715, N86);
nand NAND3 (N1734, N1726, N1574, N1377);
buf BUF1 (N1735, N1725);
xor XOR2 (N1736, N1734, N234);
buf BUF1 (N1737, N1736);
nand NAND2 (N1738, N1728, N772);
not NOT1 (N1739, N1706);
and AND4 (N1740, N1738, N1066, N1577, N513);
xor XOR2 (N1741, N1730, N1481);
not NOT1 (N1742, N1729);
and AND3 (N1743, N1739, N868, N494);
or OR3 (N1744, N1735, N123, N365);
nor NOR4 (N1745, N1731, N1450, N1183, N576);
or OR3 (N1746, N1745, N277, N568);
and AND3 (N1747, N1746, N975, N311);
buf BUF1 (N1748, N1737);
buf BUF1 (N1749, N1748);
xor XOR2 (N1750, N1732, N929);
not NOT1 (N1751, N1744);
nand NAND4 (N1752, N1749, N1669, N158, N822);
xor XOR2 (N1753, N1751, N1744);
nand NAND4 (N1754, N1741, N1232, N916, N1485);
or OR2 (N1755, N1727, N450);
xor XOR2 (N1756, N1752, N1689);
xor XOR2 (N1757, N1753, N211);
and AND3 (N1758, N1755, N1282, N222);
nand NAND3 (N1759, N1758, N464, N353);
nand NAND4 (N1760, N1757, N240, N1107, N13);
buf BUF1 (N1761, N1733);
buf BUF1 (N1762, N1756);
buf BUF1 (N1763, N1759);
and AND2 (N1764, N1743, N1661);
nor NOR3 (N1765, N1754, N236, N705);
nor NOR4 (N1766, N1762, N1365, N645, N389);
nor NOR2 (N1767, N1750, N54);
nand NAND3 (N1768, N1765, N1550, N1758);
and AND4 (N1769, N1767, N1519, N1332, N547);
not NOT1 (N1770, N1763);
and AND3 (N1771, N1742, N1240, N1669);
xor XOR2 (N1772, N1747, N869);
buf BUF1 (N1773, N1764);
xor XOR2 (N1774, N1770, N209);
nor NOR2 (N1775, N1773, N631);
not NOT1 (N1776, N1771);
xor XOR2 (N1777, N1740, N1296);
or OR4 (N1778, N1775, N790, N1747, N1668);
buf BUF1 (N1779, N1768);
buf BUF1 (N1780, N1776);
buf BUF1 (N1781, N1760);
buf BUF1 (N1782, N1778);
or OR3 (N1783, N1779, N136, N74);
not NOT1 (N1784, N1777);
nor NOR4 (N1785, N1766, N1673, N888, N897);
not NOT1 (N1786, N1782);
and AND4 (N1787, N1761, N1281, N235, N1257);
or OR3 (N1788, N1785, N1180, N738);
nand NAND3 (N1789, N1781, N128, N728);
nor NOR2 (N1790, N1784, N522);
or OR2 (N1791, N1786, N83);
xor XOR2 (N1792, N1788, N1343);
xor XOR2 (N1793, N1780, N803);
or OR3 (N1794, N1769, N660, N677);
nor NOR4 (N1795, N1787, N236, N1710, N1384);
and AND4 (N1796, N1789, N486, N505, N1343);
not NOT1 (N1797, N1783);
or OR3 (N1798, N1794, N1687, N1718);
nand NAND4 (N1799, N1790, N1467, N1638, N795);
and AND3 (N1800, N1791, N802, N214);
nor NOR4 (N1801, N1774, N740, N1695, N1490);
nand NAND4 (N1802, N1792, N1463, N905, N1650);
xor XOR2 (N1803, N1797, N1123);
not NOT1 (N1804, N1798);
xor XOR2 (N1805, N1801, N1243);
and AND3 (N1806, N1796, N1708, N449);
not NOT1 (N1807, N1800);
and AND2 (N1808, N1804, N1224);
nor NOR3 (N1809, N1799, N1493, N1575);
not NOT1 (N1810, N1802);
nand NAND4 (N1811, N1809, N53, N585, N1116);
nand NAND2 (N1812, N1808, N1035);
xor XOR2 (N1813, N1811, N1602);
nand NAND2 (N1814, N1772, N197);
not NOT1 (N1815, N1805);
not NOT1 (N1816, N1812);
buf BUF1 (N1817, N1807);
buf BUF1 (N1818, N1793);
nor NOR3 (N1819, N1817, N1073, N1449);
xor XOR2 (N1820, N1806, N1688);
not NOT1 (N1821, N1819);
not NOT1 (N1822, N1813);
not NOT1 (N1823, N1818);
nor NOR4 (N1824, N1821, N469, N1551, N1136);
and AND4 (N1825, N1803, N353, N1811, N32);
or OR2 (N1826, N1824, N1054);
nand NAND3 (N1827, N1815, N217, N399);
not NOT1 (N1828, N1810);
buf BUF1 (N1829, N1827);
nor NOR3 (N1830, N1826, N308, N1123);
xor XOR2 (N1831, N1822, N1822);
not NOT1 (N1832, N1795);
nand NAND2 (N1833, N1814, N1147);
xor XOR2 (N1834, N1832, N476);
and AND3 (N1835, N1825, N694, N1260);
and AND2 (N1836, N1835, N1273);
nor NOR4 (N1837, N1831, N1564, N1775, N647);
and AND2 (N1838, N1829, N1336);
xor XOR2 (N1839, N1837, N508);
nand NAND2 (N1840, N1816, N721);
and AND2 (N1841, N1839, N397);
nand NAND2 (N1842, N1834, N311);
nor NOR4 (N1843, N1842, N1415, N375, N1332);
or OR3 (N1844, N1833, N1351, N912);
not NOT1 (N1845, N1841);
not NOT1 (N1846, N1838);
buf BUF1 (N1847, N1843);
xor XOR2 (N1848, N1840, N909);
nor NOR4 (N1849, N1846, N330, N1832, N61);
nor NOR4 (N1850, N1823, N1265, N1057, N123);
xor XOR2 (N1851, N1848, N873);
and AND2 (N1852, N1830, N487);
nand NAND3 (N1853, N1849, N744, N1138);
not NOT1 (N1854, N1828);
not NOT1 (N1855, N1851);
nor NOR3 (N1856, N1845, N1779, N536);
nand NAND4 (N1857, N1820, N330, N1478, N1494);
xor XOR2 (N1858, N1853, N679);
or OR3 (N1859, N1858, N1461, N641);
nand NAND2 (N1860, N1852, N1356);
and AND2 (N1861, N1857, N700);
or OR3 (N1862, N1860, N496, N935);
buf BUF1 (N1863, N1856);
buf BUF1 (N1864, N1854);
xor XOR2 (N1865, N1863, N1741);
and AND2 (N1866, N1865, N1393);
not NOT1 (N1867, N1850);
nand NAND3 (N1868, N1864, N1554, N1481);
buf BUF1 (N1869, N1867);
buf BUF1 (N1870, N1859);
or OR4 (N1871, N1844, N134, N526, N759);
and AND2 (N1872, N1861, N661);
buf BUF1 (N1873, N1869);
nand NAND3 (N1874, N1871, N542, N496);
xor XOR2 (N1875, N1868, N1202);
or OR4 (N1876, N1870, N825, N399, N876);
or OR4 (N1877, N1874, N1241, N467, N52);
buf BUF1 (N1878, N1836);
buf BUF1 (N1879, N1875);
or OR3 (N1880, N1878, N66, N617);
buf BUF1 (N1881, N1872);
xor XOR2 (N1882, N1880, N845);
nor NOR4 (N1883, N1862, N1467, N288, N276);
nor NOR2 (N1884, N1847, N1237);
nor NOR4 (N1885, N1877, N1652, N1067, N532);
nor NOR2 (N1886, N1885, N982);
or OR2 (N1887, N1855, N1155);
nor NOR2 (N1888, N1879, N1505);
or OR3 (N1889, N1883, N135, N524);
nor NOR2 (N1890, N1884, N103);
buf BUF1 (N1891, N1873);
nand NAND3 (N1892, N1891, N72, N1408);
and AND2 (N1893, N1892, N806);
buf BUF1 (N1894, N1882);
buf BUF1 (N1895, N1893);
not NOT1 (N1896, N1889);
nand NAND2 (N1897, N1876, N1412);
buf BUF1 (N1898, N1890);
and AND4 (N1899, N1887, N527, N1361, N1035);
nand NAND4 (N1900, N1895, N1837, N275, N818);
nand NAND4 (N1901, N1897, N1846, N965, N477);
and AND4 (N1902, N1894, N256, N618, N1476);
nor NOR2 (N1903, N1866, N713);
buf BUF1 (N1904, N1903);
xor XOR2 (N1905, N1886, N1533);
xor XOR2 (N1906, N1888, N530);
nor NOR4 (N1907, N1906, N317, N1473, N138);
xor XOR2 (N1908, N1901, N1344);
or OR2 (N1909, N1896, N1739);
and AND3 (N1910, N1909, N1239, N1840);
nand NAND3 (N1911, N1900, N180, N347);
nor NOR2 (N1912, N1902, N1338);
buf BUF1 (N1913, N1908);
or OR2 (N1914, N1905, N1252);
buf BUF1 (N1915, N1899);
buf BUF1 (N1916, N1907);
xor XOR2 (N1917, N1904, N1373);
xor XOR2 (N1918, N1915, N1195);
and AND2 (N1919, N1913, N888);
not NOT1 (N1920, N1911);
nand NAND4 (N1921, N1898, N388, N1453, N1717);
nor NOR2 (N1922, N1921, N1348);
or OR2 (N1923, N1920, N433);
and AND4 (N1924, N1922, N1834, N946, N1051);
nand NAND3 (N1925, N1910, N519, N923);
not NOT1 (N1926, N1924);
buf BUF1 (N1927, N1919);
and AND3 (N1928, N1881, N770, N1672);
not NOT1 (N1929, N1914);
buf BUF1 (N1930, N1927);
xor XOR2 (N1931, N1929, N16);
buf BUF1 (N1932, N1926);
and AND3 (N1933, N1923, N1424, N1684);
not NOT1 (N1934, N1931);
or OR2 (N1935, N1918, N62);
and AND2 (N1936, N1912, N644);
not NOT1 (N1937, N1925);
not NOT1 (N1938, N1930);
xor XOR2 (N1939, N1916, N784);
nor NOR2 (N1940, N1934, N16);
or OR3 (N1941, N1932, N1559, N1777);
nand NAND2 (N1942, N1917, N1144);
nand NAND3 (N1943, N1936, N1693, N1852);
buf BUF1 (N1944, N1935);
buf BUF1 (N1945, N1939);
or OR4 (N1946, N1937, N1043, N1788, N1793);
and AND2 (N1947, N1933, N1714);
nor NOR4 (N1948, N1941, N305, N1403, N322);
and AND2 (N1949, N1943, N672);
and AND2 (N1950, N1948, N185);
and AND3 (N1951, N1945, N238, N401);
buf BUF1 (N1952, N1949);
or OR3 (N1953, N1952, N1030, N636);
and AND2 (N1954, N1940, N534);
buf BUF1 (N1955, N1954);
buf BUF1 (N1956, N1947);
buf BUF1 (N1957, N1951);
or OR2 (N1958, N1956, N1692);
and AND4 (N1959, N1946, N883, N647, N429);
buf BUF1 (N1960, N1944);
and AND3 (N1961, N1938, N1686, N1085);
or OR2 (N1962, N1958, N170);
not NOT1 (N1963, N1955);
and AND4 (N1964, N1961, N634, N409, N784);
xor XOR2 (N1965, N1963, N882);
and AND2 (N1966, N1962, N1271);
buf BUF1 (N1967, N1928);
xor XOR2 (N1968, N1964, N434);
nand NAND4 (N1969, N1965, N174, N497, N374);
nor NOR2 (N1970, N1966, N62);
or OR2 (N1971, N1950, N585);
xor XOR2 (N1972, N1959, N1731);
buf BUF1 (N1973, N1971);
not NOT1 (N1974, N1942);
buf BUF1 (N1975, N1972);
nor NOR3 (N1976, N1967, N807, N1330);
and AND3 (N1977, N1974, N542, N1944);
and AND2 (N1978, N1969, N1413);
and AND3 (N1979, N1976, N669, N1052);
nand NAND4 (N1980, N1979, N1308, N1105, N426);
nand NAND3 (N1981, N1968, N655, N1783);
nor NOR4 (N1982, N1957, N1531, N801, N962);
and AND2 (N1983, N1981, N1472);
and AND3 (N1984, N1953, N1557, N868);
not NOT1 (N1985, N1970);
or OR4 (N1986, N1960, N117, N1785, N131);
and AND4 (N1987, N1983, N566, N152, N15);
or OR4 (N1988, N1987, N1314, N1603, N1144);
xor XOR2 (N1989, N1988, N1952);
buf BUF1 (N1990, N1977);
or OR2 (N1991, N1980, N44);
buf BUF1 (N1992, N1990);
nor NOR3 (N1993, N1989, N1225, N340);
or OR4 (N1994, N1986, N864, N1644, N505);
xor XOR2 (N1995, N1978, N1312);
nand NAND2 (N1996, N1995, N1903);
and AND3 (N1997, N1985, N739, N1938);
xor XOR2 (N1998, N1994, N1207);
or OR3 (N1999, N1993, N662, N1815);
not NOT1 (N2000, N1998);
buf BUF1 (N2001, N1991);
nand NAND4 (N2002, N1999, N1369, N1688, N448);
not NOT1 (N2003, N2002);
xor XOR2 (N2004, N2000, N915);
not NOT1 (N2005, N1992);
and AND4 (N2006, N1984, N986, N1355, N1142);
xor XOR2 (N2007, N1997, N959);
not NOT1 (N2008, N1975);
buf BUF1 (N2009, N2006);
buf BUF1 (N2010, N1996);
and AND2 (N2011, N2010, N538);
nor NOR4 (N2012, N2009, N809, N429, N1589);
nor NOR3 (N2013, N1982, N247, N1724);
nand NAND3 (N2014, N2011, N1238, N282);
xor XOR2 (N2015, N1973, N1472);
xor XOR2 (N2016, N2012, N1708);
or OR2 (N2017, N2013, N1849);
nand NAND4 (N2018, N2004, N562, N1844, N510);
nand NAND4 (N2019, N2017, N1624, N1467, N649);
buf BUF1 (N2020, N2015);
nand NAND2 (N2021, N2008, N834);
xor XOR2 (N2022, N2007, N655);
xor XOR2 (N2023, N2019, N169);
or OR4 (N2024, N2020, N1701, N1744, N709);
not NOT1 (N2025, N2014);
nor NOR4 (N2026, N2021, N1052, N1238, N1699);
xor XOR2 (N2027, N2005, N724);
nor NOR3 (N2028, N2018, N981, N1369);
not NOT1 (N2029, N2023);
buf BUF1 (N2030, N2001);
or OR2 (N2031, N2016, N411);
xor XOR2 (N2032, N2025, N61);
buf BUF1 (N2033, N2028);
not NOT1 (N2034, N2030);
not NOT1 (N2035, N2022);
or OR2 (N2036, N2035, N1838);
buf BUF1 (N2037, N2036);
and AND3 (N2038, N2026, N347, N1182);
xor XOR2 (N2039, N2038, N1712);
or OR2 (N2040, N2032, N1227);
not NOT1 (N2041, N2024);
nand NAND3 (N2042, N2041, N1356, N853);
nor NOR2 (N2043, N2029, N227);
nand NAND2 (N2044, N2042, N1951);
nor NOR2 (N2045, N2044, N265);
not NOT1 (N2046, N2033);
nor NOR3 (N2047, N2027, N1925, N1265);
nor NOR3 (N2048, N2040, N829, N429);
nor NOR3 (N2049, N2003, N1610, N1676);
and AND4 (N2050, N2045, N1475, N1849, N147);
and AND3 (N2051, N2050, N635, N1526);
buf BUF1 (N2052, N2043);
buf BUF1 (N2053, N2031);
and AND4 (N2054, N2039, N867, N162, N296);
nand NAND2 (N2055, N2054, N1316);
not NOT1 (N2056, N2034);
or OR3 (N2057, N2055, N683, N1102);
not NOT1 (N2058, N2052);
and AND4 (N2059, N2053, N1396, N606, N1842);
xor XOR2 (N2060, N2049, N1024);
buf BUF1 (N2061, N2046);
nand NAND2 (N2062, N2051, N1825);
nor NOR2 (N2063, N2057, N258);
buf BUF1 (N2064, N2048);
xor XOR2 (N2065, N2037, N1941);
or OR4 (N2066, N2063, N565, N1331, N592);
and AND2 (N2067, N2065, N1691);
xor XOR2 (N2068, N2061, N466);
nand NAND2 (N2069, N2064, N2004);
nor NOR2 (N2070, N2066, N1852);
buf BUF1 (N2071, N2062);
and AND3 (N2072, N2059, N1834, N1818);
and AND2 (N2073, N2067, N96);
buf BUF1 (N2074, N2072);
not NOT1 (N2075, N2070);
nand NAND2 (N2076, N2073, N1313);
xor XOR2 (N2077, N2056, N686);
buf BUF1 (N2078, N2075);
xor XOR2 (N2079, N2074, N1870);
nand NAND4 (N2080, N2058, N967, N1454, N1207);
or OR2 (N2081, N2078, N1315);
and AND3 (N2082, N2076, N1813, N300);
nor NOR4 (N2083, N2068, N1404, N969, N627);
and AND4 (N2084, N2080, N772, N1577, N1928);
and AND3 (N2085, N2069, N904, N916);
or OR3 (N2086, N2082, N286, N1630);
nand NAND4 (N2087, N2085, N483, N1172, N1419);
nor NOR2 (N2088, N2047, N1635);
nand NAND4 (N2089, N2083, N1671, N989, N1074);
xor XOR2 (N2090, N2081, N297);
or OR4 (N2091, N2084, N91, N338, N784);
buf BUF1 (N2092, N2090);
and AND2 (N2093, N2060, N213);
not NOT1 (N2094, N2086);
or OR4 (N2095, N2089, N334, N2088, N1991);
or OR3 (N2096, N488, N1303, N96);
and AND4 (N2097, N2087, N1270, N781, N1285);
not NOT1 (N2098, N2071);
xor XOR2 (N2099, N2095, N1385);
xor XOR2 (N2100, N2094, N1815);
or OR3 (N2101, N2091, N2024, N668);
nor NOR2 (N2102, N2097, N1402);
and AND2 (N2103, N2100, N1765);
nand NAND3 (N2104, N2099, N2007, N1442);
xor XOR2 (N2105, N2098, N966);
buf BUF1 (N2106, N2102);
nand NAND2 (N2107, N2092, N816);
nand NAND3 (N2108, N2107, N718, N794);
nor NOR4 (N2109, N2077, N240, N1521, N1039);
nor NOR4 (N2110, N2101, N383, N636, N1189);
not NOT1 (N2111, N2079);
buf BUF1 (N2112, N2106);
and AND3 (N2113, N2105, N1414, N428);
buf BUF1 (N2114, N2108);
and AND2 (N2115, N2111, N316);
or OR2 (N2116, N2103, N1910);
nor NOR4 (N2117, N2109, N1071, N2063, N1846);
and AND3 (N2118, N2093, N1163, N992);
xor XOR2 (N2119, N2110, N1238);
not NOT1 (N2120, N2115);
nand NAND4 (N2121, N2104, N100, N1987, N920);
buf BUF1 (N2122, N2116);
xor XOR2 (N2123, N2096, N1762);
buf BUF1 (N2124, N2122);
and AND2 (N2125, N2119, N1199);
xor XOR2 (N2126, N2124, N381);
not NOT1 (N2127, N2125);
and AND4 (N2128, N2123, N1052, N719, N101);
nand NAND2 (N2129, N2112, N292);
and AND4 (N2130, N2120, N1204, N710, N32);
buf BUF1 (N2131, N2121);
xor XOR2 (N2132, N2129, N742);
and AND4 (N2133, N2128, N1684, N2027, N119);
or OR3 (N2134, N2133, N1200, N1612);
nand NAND4 (N2135, N2126, N87, N974, N1596);
nand NAND4 (N2136, N2134, N707, N1873, N1132);
xor XOR2 (N2137, N2127, N874);
nor NOR3 (N2138, N2131, N1855, N384);
nor NOR4 (N2139, N2138, N1094, N1103, N432);
xor XOR2 (N2140, N2136, N1525);
and AND4 (N2141, N2139, N2078, N1553, N835);
xor XOR2 (N2142, N2113, N1618);
or OR3 (N2143, N2135, N1518, N1815);
nor NOR4 (N2144, N2137, N860, N1544, N1228);
nor NOR4 (N2145, N2130, N52, N651, N1644);
and AND2 (N2146, N2142, N1638);
not NOT1 (N2147, N2146);
not NOT1 (N2148, N2132);
xor XOR2 (N2149, N2145, N879);
nor NOR4 (N2150, N2147, N1244, N2027, N130);
buf BUF1 (N2151, N2140);
not NOT1 (N2152, N2118);
or OR4 (N2153, N2144, N745, N1572, N782);
nand NAND2 (N2154, N2150, N973);
buf BUF1 (N2155, N2153);
not NOT1 (N2156, N2152);
or OR4 (N2157, N2155, N895, N2149, N1641);
and AND2 (N2158, N1638, N425);
nor NOR2 (N2159, N2158, N648);
or OR2 (N2160, N2154, N789);
nor NOR2 (N2161, N2156, N1979);
and AND4 (N2162, N2161, N1807, N1117, N1238);
not NOT1 (N2163, N2114);
nand NAND4 (N2164, N2141, N1186, N57, N1209);
and AND3 (N2165, N2164, N210, N24);
buf BUF1 (N2166, N2148);
nand NAND3 (N2167, N2162, N1140, N1634);
and AND2 (N2168, N2117, N863);
buf BUF1 (N2169, N2159);
and AND4 (N2170, N2163, N1550, N1708, N1959);
buf BUF1 (N2171, N2143);
or OR3 (N2172, N2166, N874, N1121);
or OR3 (N2173, N2165, N347, N917);
or OR4 (N2174, N2167, N1949, N1153, N1284);
and AND4 (N2175, N2174, N1800, N918, N927);
nand NAND4 (N2176, N2171, N675, N1483, N1169);
not NOT1 (N2177, N2172);
nand NAND4 (N2178, N2160, N131, N873, N938);
not NOT1 (N2179, N2151);
xor XOR2 (N2180, N2157, N148);
xor XOR2 (N2181, N2178, N1072);
not NOT1 (N2182, N2175);
xor XOR2 (N2183, N2173, N1962);
or OR2 (N2184, N2179, N86);
xor XOR2 (N2185, N2168, N1637);
nor NOR4 (N2186, N2183, N418, N545, N1916);
xor XOR2 (N2187, N2169, N1897);
nand NAND4 (N2188, N2181, N2064, N1929, N1939);
or OR2 (N2189, N2180, N1085);
buf BUF1 (N2190, N2189);
nand NAND4 (N2191, N2186, N540, N1658, N1043);
nand NAND4 (N2192, N2191, N125, N1071, N571);
and AND2 (N2193, N2187, N1916);
nand NAND4 (N2194, N2185, N1183, N313, N734);
or OR4 (N2195, N2194, N1776, N594, N222);
xor XOR2 (N2196, N2193, N1397);
nand NAND4 (N2197, N2192, N294, N1573, N87);
or OR3 (N2198, N2182, N1914, N1076);
xor XOR2 (N2199, N2188, N1610);
xor XOR2 (N2200, N2198, N1700);
nand NAND3 (N2201, N2195, N224, N1190);
and AND3 (N2202, N2200, N1846, N1260);
xor XOR2 (N2203, N2176, N1870);
xor XOR2 (N2204, N2184, N1551);
or OR3 (N2205, N2202, N895, N264);
not NOT1 (N2206, N2190);
xor XOR2 (N2207, N2177, N147);
not NOT1 (N2208, N2170);
xor XOR2 (N2209, N2203, N2138);
xor XOR2 (N2210, N2208, N197);
or OR3 (N2211, N2201, N797, N1057);
xor XOR2 (N2212, N2204, N727);
or OR3 (N2213, N2212, N13, N437);
or OR3 (N2214, N2213, N139, N490);
xor XOR2 (N2215, N2211, N2121);
nand NAND2 (N2216, N2214, N1929);
not NOT1 (N2217, N2205);
nand NAND2 (N2218, N2207, N1826);
xor XOR2 (N2219, N2215, N1358);
nand NAND3 (N2220, N2216, N1986, N828);
not NOT1 (N2221, N2209);
nand NAND2 (N2222, N2206, N370);
buf BUF1 (N2223, N2219);
xor XOR2 (N2224, N2217, N673);
not NOT1 (N2225, N2222);
and AND4 (N2226, N2220, N948, N1064, N1288);
not NOT1 (N2227, N2225);
and AND4 (N2228, N2218, N1051, N362, N690);
or OR4 (N2229, N2221, N2228, N1124, N1711);
and AND2 (N2230, N1908, N166);
and AND4 (N2231, N2223, N1046, N495, N2075);
buf BUF1 (N2232, N2199);
not NOT1 (N2233, N2224);
and AND4 (N2234, N2230, N1852, N543, N1044);
not NOT1 (N2235, N2196);
not NOT1 (N2236, N2197);
not NOT1 (N2237, N2229);
nand NAND4 (N2238, N2232, N1011, N1351, N758);
nand NAND3 (N2239, N2226, N560, N1672);
nor NOR2 (N2240, N2210, N1285);
nand NAND4 (N2241, N2227, N209, N1526, N1419);
nand NAND4 (N2242, N2241, N1900, N1475, N1039);
buf BUF1 (N2243, N2235);
and AND3 (N2244, N2242, N1243, N2014);
nor NOR3 (N2245, N2243, N1433, N1270);
and AND2 (N2246, N2233, N702);
buf BUF1 (N2247, N2244);
nand NAND3 (N2248, N2234, N1976, N564);
xor XOR2 (N2249, N2238, N644);
and AND4 (N2250, N2246, N116, N2140, N759);
not NOT1 (N2251, N2245);
nand NAND3 (N2252, N2247, N2156, N687);
and AND4 (N2253, N2240, N457, N498, N1026);
not NOT1 (N2254, N2237);
not NOT1 (N2255, N2249);
xor XOR2 (N2256, N2250, N1947);
or OR3 (N2257, N2239, N1625, N1541);
buf BUF1 (N2258, N2255);
or OR3 (N2259, N2258, N865, N314);
nor NOR2 (N2260, N2256, N1617);
or OR3 (N2261, N2254, N922, N132);
or OR3 (N2262, N2252, N2171, N86);
buf BUF1 (N2263, N2253);
not NOT1 (N2264, N2248);
or OR4 (N2265, N2260, N311, N372, N676);
nor NOR3 (N2266, N2263, N149, N192);
buf BUF1 (N2267, N2257);
xor XOR2 (N2268, N2265, N1280);
nor NOR2 (N2269, N2267, N177);
or OR2 (N2270, N2251, N1211);
nand NAND4 (N2271, N2261, N1314, N2154, N1123);
buf BUF1 (N2272, N2264);
buf BUF1 (N2273, N2269);
nand NAND4 (N2274, N2231, N654, N1587, N805);
and AND4 (N2275, N2270, N1038, N1499, N922);
nand NAND3 (N2276, N2262, N817, N477);
nor NOR3 (N2277, N2236, N1570, N217);
and AND2 (N2278, N2271, N1810);
or OR3 (N2279, N2259, N1052, N1079);
not NOT1 (N2280, N2268);
not NOT1 (N2281, N2275);
not NOT1 (N2282, N2278);
xor XOR2 (N2283, N2272, N1734);
not NOT1 (N2284, N2276);
nor NOR4 (N2285, N2273, N1226, N663, N2193);
xor XOR2 (N2286, N2266, N581);
xor XOR2 (N2287, N2284, N983);
buf BUF1 (N2288, N2282);
or OR2 (N2289, N2288, N2096);
nand NAND4 (N2290, N2281, N65, N1699, N961);
or OR2 (N2291, N2277, N161);
not NOT1 (N2292, N2291);
and AND3 (N2293, N2292, N2051, N783);
xor XOR2 (N2294, N2279, N2020);
nand NAND4 (N2295, N2285, N1457, N813, N1196);
and AND3 (N2296, N2287, N2036, N1716);
nor NOR2 (N2297, N2290, N164);
xor XOR2 (N2298, N2274, N994);
nor NOR3 (N2299, N2297, N2209, N1844);
buf BUF1 (N2300, N2289);
buf BUF1 (N2301, N2296);
buf BUF1 (N2302, N2280);
and AND3 (N2303, N2299, N1889, N1029);
or OR2 (N2304, N2294, N389);
and AND4 (N2305, N2300, N479, N677, N2224);
xor XOR2 (N2306, N2301, N1672);
or OR4 (N2307, N2302, N12, N1627, N1746);
and AND2 (N2308, N2283, N1);
xor XOR2 (N2309, N2307, N1403);
not NOT1 (N2310, N2304);
and AND3 (N2311, N2309, N590, N851);
and AND2 (N2312, N2305, N2278);
nand NAND4 (N2313, N2295, N48, N1210, N818);
or OR4 (N2314, N2306, N1323, N205, N273);
and AND4 (N2315, N2303, N1915, N1451, N631);
not NOT1 (N2316, N2313);
not NOT1 (N2317, N2314);
and AND4 (N2318, N2316, N1193, N1071, N112);
nand NAND3 (N2319, N2318, N674, N1273);
nor NOR4 (N2320, N2293, N2150, N1067, N808);
not NOT1 (N2321, N2298);
nand NAND4 (N2322, N2317, N306, N155, N2194);
and AND3 (N2323, N2320, N1028, N1364);
and AND4 (N2324, N2311, N2240, N257, N1964);
nor NOR4 (N2325, N2323, N1508, N1394, N1788);
xor XOR2 (N2326, N2308, N1821);
xor XOR2 (N2327, N2326, N653);
not NOT1 (N2328, N2322);
nand NAND3 (N2329, N2328, N545, N1644);
buf BUF1 (N2330, N2312);
nand NAND3 (N2331, N2310, N1551, N1933);
nand NAND3 (N2332, N2330, N1429, N1634);
or OR3 (N2333, N2315, N149, N1349);
nor NOR3 (N2334, N2327, N1403, N671);
buf BUF1 (N2335, N2286);
buf BUF1 (N2336, N2333);
not NOT1 (N2337, N2321);
nand NAND2 (N2338, N2329, N1670);
or OR3 (N2339, N2334, N760, N1310);
xor XOR2 (N2340, N2337, N1584);
buf BUF1 (N2341, N2319);
nand NAND2 (N2342, N2325, N543);
nand NAND2 (N2343, N2332, N959);
not NOT1 (N2344, N2342);
nor NOR3 (N2345, N2338, N1482, N2032);
not NOT1 (N2346, N2341);
nand NAND3 (N2347, N2344, N881, N393);
buf BUF1 (N2348, N2347);
nand NAND3 (N2349, N2335, N2205, N1595);
buf BUF1 (N2350, N2348);
buf BUF1 (N2351, N2340);
not NOT1 (N2352, N2349);
buf BUF1 (N2353, N2346);
not NOT1 (N2354, N2345);
xor XOR2 (N2355, N2354, N800);
nand NAND2 (N2356, N2324, N1319);
nand NAND4 (N2357, N2353, N1655, N424, N1919);
and AND2 (N2358, N2343, N641);
and AND2 (N2359, N2339, N1608);
and AND3 (N2360, N2351, N2327, N2011);
xor XOR2 (N2361, N2360, N1142);
nand NAND3 (N2362, N2356, N22, N1579);
not NOT1 (N2363, N2361);
and AND4 (N2364, N2331, N645, N1482, N888);
and AND3 (N2365, N2352, N793, N1609);
buf BUF1 (N2366, N2364);
nand NAND3 (N2367, N2358, N2169, N2254);
xor XOR2 (N2368, N2359, N1082);
nor NOR3 (N2369, N2363, N630, N1742);
nor NOR2 (N2370, N2369, N1217);
xor XOR2 (N2371, N2336, N1122);
and AND2 (N2372, N2367, N2067);
buf BUF1 (N2373, N2372);
buf BUF1 (N2374, N2373);
or OR3 (N2375, N2350, N507, N2295);
and AND3 (N2376, N2355, N311, N94);
and AND4 (N2377, N2375, N2245, N352, N837);
and AND4 (N2378, N2368, N907, N647, N34);
and AND2 (N2379, N2376, N1971);
or OR2 (N2380, N2362, N2079);
not NOT1 (N2381, N2379);
nor NOR3 (N2382, N2380, N702, N40);
nor NOR2 (N2383, N2377, N843);
nand NAND2 (N2384, N2374, N1418);
nor NOR3 (N2385, N2370, N258, N975);
not NOT1 (N2386, N2365);
nand NAND3 (N2387, N2381, N1998, N105);
and AND2 (N2388, N2384, N2333);
buf BUF1 (N2389, N2387);
nand NAND3 (N2390, N2382, N1553, N719);
nand NAND2 (N2391, N2357, N935);
or OR4 (N2392, N2388, N2206, N1067, N1145);
not NOT1 (N2393, N2383);
buf BUF1 (N2394, N2386);
nor NOR2 (N2395, N2392, N309);
or OR4 (N2396, N2391, N2024, N1435, N748);
and AND2 (N2397, N2390, N1676);
not NOT1 (N2398, N2396);
xor XOR2 (N2399, N2395, N1430);
buf BUF1 (N2400, N2389);
xor XOR2 (N2401, N2394, N2180);
nand NAND4 (N2402, N2397, N2, N1660, N1424);
nand NAND3 (N2403, N2366, N1022, N107);
not NOT1 (N2404, N2399);
nor NOR2 (N2405, N2371, N481);
and AND4 (N2406, N2401, N2096, N1478, N961);
nand NAND4 (N2407, N2400, N2218, N224, N451);
nor NOR4 (N2408, N2403, N474, N1641, N295);
not NOT1 (N2409, N2404);
nand NAND4 (N2410, N2407, N611, N1436, N2011);
not NOT1 (N2411, N2378);
not NOT1 (N2412, N2385);
xor XOR2 (N2413, N2406, N1033);
nor NOR4 (N2414, N2410, N795, N1253, N422);
or OR2 (N2415, N2409, N814);
not NOT1 (N2416, N2408);
buf BUF1 (N2417, N2411);
nand NAND3 (N2418, N2415, N1493, N1476);
nor NOR3 (N2419, N2417, N262, N132);
not NOT1 (N2420, N2412);
buf BUF1 (N2421, N2416);
nand NAND3 (N2422, N2393, N2263, N2127);
xor XOR2 (N2423, N2422, N665);
nor NOR4 (N2424, N2419, N1378, N2421, N835);
not NOT1 (N2425, N2058);
or OR4 (N2426, N2398, N137, N955, N1798);
and AND4 (N2427, N2414, N388, N1512, N1492);
not NOT1 (N2428, N2425);
and AND2 (N2429, N2413, N1812);
nor NOR3 (N2430, N2418, N1939, N874);
not NOT1 (N2431, N2405);
buf BUF1 (N2432, N2430);
nor NOR3 (N2433, N2426, N1860, N1410);
xor XOR2 (N2434, N2423, N1186);
or OR4 (N2435, N2432, N229, N1703, N1041);
nor NOR4 (N2436, N2428, N1596, N610, N1350);
nor NOR3 (N2437, N2434, N755, N102);
nor NOR2 (N2438, N2424, N813);
xor XOR2 (N2439, N2429, N361);
nor NOR4 (N2440, N2433, N591, N907, N2414);
nand NAND3 (N2441, N2440, N1786, N493);
not NOT1 (N2442, N2436);
not NOT1 (N2443, N2439);
nand NAND4 (N2444, N2441, N1430, N1777, N892);
or OR4 (N2445, N2427, N264, N1610, N230);
not NOT1 (N2446, N2438);
not NOT1 (N2447, N2446);
or OR4 (N2448, N2443, N390, N1062, N1641);
not NOT1 (N2449, N2420);
nand NAND4 (N2450, N2445, N314, N2385, N2298);
buf BUF1 (N2451, N2449);
xor XOR2 (N2452, N2447, N1172);
nand NAND4 (N2453, N2448, N898, N1135, N871);
buf BUF1 (N2454, N2431);
nor NOR4 (N2455, N2442, N163, N1797, N493);
nand NAND2 (N2456, N2451, N1442);
not NOT1 (N2457, N2453);
xor XOR2 (N2458, N2450, N162);
xor XOR2 (N2459, N2455, N665);
or OR2 (N2460, N2444, N313);
nand NAND4 (N2461, N2458, N1804, N1703, N455);
and AND4 (N2462, N2459, N1169, N168, N1733);
or OR2 (N2463, N2452, N1538);
buf BUF1 (N2464, N2437);
nand NAND2 (N2465, N2454, N774);
or OR4 (N2466, N2456, N871, N161, N1414);
nand NAND3 (N2467, N2466, N260, N468);
nand NAND3 (N2468, N2435, N257, N2259);
and AND4 (N2469, N2457, N1505, N2133, N1597);
not NOT1 (N2470, N2464);
xor XOR2 (N2471, N2461, N2326);
and AND3 (N2472, N2467, N270, N779);
nand NAND3 (N2473, N2460, N1768, N1354);
or OR3 (N2474, N2462, N2303, N1827);
nand NAND4 (N2475, N2402, N1082, N1197, N1290);
buf BUF1 (N2476, N2474);
nand NAND2 (N2477, N2469, N604);
buf BUF1 (N2478, N2468);
and AND2 (N2479, N2473, N1252);
nor NOR2 (N2480, N2463, N757);
xor XOR2 (N2481, N2470, N231);
buf BUF1 (N2482, N2479);
or OR3 (N2483, N2471, N2398, N797);
not NOT1 (N2484, N2472);
or OR2 (N2485, N2480, N1706);
and AND3 (N2486, N2478, N2087, N66);
or OR3 (N2487, N2482, N708, N1322);
nand NAND3 (N2488, N2483, N316, N857);
or OR4 (N2489, N2488, N1592, N1854, N1171);
or OR2 (N2490, N2476, N1381);
xor XOR2 (N2491, N2485, N1685);
and AND3 (N2492, N2484, N1935, N1712);
nand NAND4 (N2493, N2487, N1614, N1551, N2128);
buf BUF1 (N2494, N2481);
nand NAND4 (N2495, N2489, N112, N1988, N2319);
nor NOR2 (N2496, N2465, N1549);
nand NAND2 (N2497, N2493, N294);
buf BUF1 (N2498, N2477);
nand NAND3 (N2499, N2495, N2483, N1968);
not NOT1 (N2500, N2494);
nor NOR2 (N2501, N2500, N1752);
buf BUF1 (N2502, N2491);
nand NAND3 (N2503, N2498, N2001, N1438);
or OR3 (N2504, N2492, N1559, N1165);
nor NOR3 (N2505, N2499, N1230, N881);
buf BUF1 (N2506, N2497);
xor XOR2 (N2507, N2505, N2275);
and AND3 (N2508, N2504, N1575, N2501);
buf BUF1 (N2509, N39);
nor NOR2 (N2510, N2508, N2288);
xor XOR2 (N2511, N2503, N515);
or OR4 (N2512, N2486, N862, N2094, N942);
nor NOR2 (N2513, N2490, N62);
or OR2 (N2514, N2511, N1085);
nand NAND4 (N2515, N2510, N1747, N281, N1249);
or OR4 (N2516, N2502, N2331, N2025, N852);
buf BUF1 (N2517, N2513);
xor XOR2 (N2518, N2517, N1588);
nor NOR3 (N2519, N2515, N26, N2280);
xor XOR2 (N2520, N2516, N1500);
and AND4 (N2521, N2509, N968, N474, N1928);
and AND4 (N2522, N2519, N18, N2048, N506);
and AND4 (N2523, N2518, N24, N442, N1823);
nand NAND2 (N2524, N2512, N1192);
xor XOR2 (N2525, N2507, N1021);
and AND4 (N2526, N2496, N1607, N2007, N688);
or OR4 (N2527, N2520, N1585, N1896, N1444);
or OR4 (N2528, N2514, N1293, N450, N1324);
nand NAND2 (N2529, N2475, N306);
nand NAND2 (N2530, N2524, N1612);
nor NOR2 (N2531, N2522, N1172);
nor NOR4 (N2532, N2521, N373, N1034, N1166);
or OR4 (N2533, N2529, N1012, N327, N1193);
buf BUF1 (N2534, N2528);
nor NOR4 (N2535, N2530, N701, N393, N682);
nand NAND4 (N2536, N2523, N335, N1275, N903);
buf BUF1 (N2537, N2532);
and AND4 (N2538, N2527, N722, N2136, N1724);
xor XOR2 (N2539, N2526, N1552);
nor NOR4 (N2540, N2534, N507, N2145, N1908);
and AND3 (N2541, N2538, N1130, N477);
not NOT1 (N2542, N2525);
or OR3 (N2543, N2536, N561, N464);
xor XOR2 (N2544, N2541, N410);
buf BUF1 (N2545, N2542);
or OR4 (N2546, N2535, N495, N622, N2387);
and AND3 (N2547, N2545, N894, N1873);
buf BUF1 (N2548, N2533);
and AND4 (N2549, N2537, N1596, N1588, N14);
nor NOR2 (N2550, N2547, N427);
not NOT1 (N2551, N2550);
xor XOR2 (N2552, N2549, N755);
nand NAND2 (N2553, N2543, N2168);
and AND2 (N2554, N2546, N1207);
buf BUF1 (N2555, N2540);
and AND4 (N2556, N2506, N1710, N2486, N240);
nor NOR3 (N2557, N2548, N724, N180);
not NOT1 (N2558, N2553);
not NOT1 (N2559, N2531);
xor XOR2 (N2560, N2559, N973);
buf BUF1 (N2561, N2552);
buf BUF1 (N2562, N2544);
or OR3 (N2563, N2558, N1386, N762);
and AND4 (N2564, N2563, N1235, N882, N1108);
nor NOR4 (N2565, N2551, N2283, N2295, N1945);
xor XOR2 (N2566, N2554, N371);
nand NAND2 (N2567, N2555, N886);
not NOT1 (N2568, N2556);
or OR2 (N2569, N2565, N1728);
xor XOR2 (N2570, N2567, N2387);
xor XOR2 (N2571, N2570, N597);
nor NOR2 (N2572, N2561, N1197);
and AND4 (N2573, N2571, N1468, N1354, N411);
not NOT1 (N2574, N2557);
not NOT1 (N2575, N2539);
and AND3 (N2576, N2572, N2564, N2541);
not NOT1 (N2577, N192);
nand NAND2 (N2578, N2574, N50);
or OR4 (N2579, N2578, N331, N2419, N1240);
nor NOR2 (N2580, N2562, N2398);
buf BUF1 (N2581, N2568);
and AND4 (N2582, N2580, N2387, N181, N2497);
buf BUF1 (N2583, N2582);
xor XOR2 (N2584, N2560, N2118);
not NOT1 (N2585, N2577);
not NOT1 (N2586, N2573);
nor NOR2 (N2587, N2585, N930);
nand NAND4 (N2588, N2584, N1157, N901, N1102);
and AND4 (N2589, N2587, N1664, N1017, N1862);
nor NOR2 (N2590, N2566, N1564);
nor NOR4 (N2591, N2583, N338, N153, N168);
nand NAND2 (N2592, N2581, N2105);
xor XOR2 (N2593, N2586, N138);
not NOT1 (N2594, N2576);
xor XOR2 (N2595, N2590, N1986);
not NOT1 (N2596, N2569);
buf BUF1 (N2597, N2594);
buf BUF1 (N2598, N2579);
nor NOR3 (N2599, N2592, N2597, N1353);
buf BUF1 (N2600, N1923);
buf BUF1 (N2601, N2595);
xor XOR2 (N2602, N2598, N2458);
or OR4 (N2603, N2602, N1544, N1254, N942);
and AND2 (N2604, N2588, N2454);
xor XOR2 (N2605, N2600, N971);
or OR3 (N2606, N2599, N194, N701);
or OR4 (N2607, N2606, N628, N432, N2195);
and AND3 (N2608, N2605, N1013, N1118);
or OR3 (N2609, N2575, N1725, N1535);
nor NOR2 (N2610, N2601, N66);
nor NOR4 (N2611, N2604, N2216, N1856, N1240);
xor XOR2 (N2612, N2608, N1349);
nor NOR3 (N2613, N2591, N858, N2136);
nand NAND3 (N2614, N2593, N1100, N2125);
and AND3 (N2615, N2610, N1830, N441);
nor NOR2 (N2616, N2607, N2189);
and AND2 (N2617, N2603, N1184);
or OR2 (N2618, N2612, N1054);
and AND3 (N2619, N2589, N1301, N162);
nand NAND2 (N2620, N2619, N547);
and AND4 (N2621, N2618, N386, N177, N1002);
and AND4 (N2622, N2611, N2284, N2341, N74);
not NOT1 (N2623, N2613);
or OR3 (N2624, N2617, N1160, N2052);
xor XOR2 (N2625, N2616, N694);
nand NAND3 (N2626, N2622, N728, N118);
nand NAND4 (N2627, N2615, N1092, N2436, N879);
xor XOR2 (N2628, N2620, N654);
xor XOR2 (N2629, N2609, N2589);
not NOT1 (N2630, N2624);
nand NAND3 (N2631, N2623, N2001, N365);
and AND4 (N2632, N2630, N951, N1810, N776);
nand NAND3 (N2633, N2614, N2531, N2334);
xor XOR2 (N2634, N2631, N2096);
nor NOR4 (N2635, N2596, N992, N267, N1182);
not NOT1 (N2636, N2627);
not NOT1 (N2637, N2629);
xor XOR2 (N2638, N2626, N1179);
and AND4 (N2639, N2625, N1485, N923, N2167);
and AND3 (N2640, N2636, N962, N81);
and AND3 (N2641, N2628, N1653, N2186);
nand NAND2 (N2642, N2637, N1371);
nor NOR3 (N2643, N2641, N2306, N297);
and AND4 (N2644, N2640, N616, N635, N2108);
nor NOR2 (N2645, N2634, N2133);
or OR3 (N2646, N2645, N467, N203);
not NOT1 (N2647, N2638);
xor XOR2 (N2648, N2633, N2426);
or OR2 (N2649, N2642, N1083);
nor NOR4 (N2650, N2649, N789, N1013, N2292);
not NOT1 (N2651, N2644);
and AND4 (N2652, N2621, N1912, N1850, N123);
and AND3 (N2653, N2651, N570, N2090);
nand NAND4 (N2654, N2643, N2172, N1963, N837);
buf BUF1 (N2655, N2650);
not NOT1 (N2656, N2648);
nor NOR2 (N2657, N2639, N705);
not NOT1 (N2658, N2635);
not NOT1 (N2659, N2647);
xor XOR2 (N2660, N2632, N2358);
or OR3 (N2661, N2659, N225, N1977);
not NOT1 (N2662, N2656);
xor XOR2 (N2663, N2661, N898);
buf BUF1 (N2664, N2663);
nor NOR3 (N2665, N2662, N2113, N1199);
xor XOR2 (N2666, N2646, N1333);
buf BUF1 (N2667, N2653);
xor XOR2 (N2668, N2658, N1933);
not NOT1 (N2669, N2660);
buf BUF1 (N2670, N2669);
nand NAND2 (N2671, N2652, N674);
or OR2 (N2672, N2655, N2055);
and AND3 (N2673, N2664, N2185, N36);
or OR4 (N2674, N2668, N286, N1214, N931);
xor XOR2 (N2675, N2657, N2125);
or OR3 (N2676, N2671, N1287, N2428);
nand NAND2 (N2677, N2673, N2438);
nor NOR2 (N2678, N2674, N309);
nand NAND4 (N2679, N2667, N1016, N1890, N1003);
or OR4 (N2680, N2670, N2574, N2120, N399);
buf BUF1 (N2681, N2672);
not NOT1 (N2682, N2681);
nand NAND3 (N2683, N2654, N709, N282);
not NOT1 (N2684, N2678);
nor NOR3 (N2685, N2684, N1, N2085);
not NOT1 (N2686, N2677);
not NOT1 (N2687, N2685);
nand NAND2 (N2688, N2666, N1062);
xor XOR2 (N2689, N2688, N2344);
nand NAND3 (N2690, N2676, N995, N1522);
buf BUF1 (N2691, N2680);
nor NOR4 (N2692, N2683, N1603, N1606, N1791);
not NOT1 (N2693, N2665);
buf BUF1 (N2694, N2693);
not NOT1 (N2695, N2682);
or OR4 (N2696, N2691, N1280, N2464, N1336);
nor NOR3 (N2697, N2675, N581, N1628);
xor XOR2 (N2698, N2696, N670);
not NOT1 (N2699, N2692);
nor NOR2 (N2700, N2690, N2006);
or OR4 (N2701, N2689, N2541, N2574, N1929);
not NOT1 (N2702, N2698);
nor NOR3 (N2703, N2699, N733, N1302);
nor NOR4 (N2704, N2701, N223, N1758, N1836);
and AND3 (N2705, N2700, N1274, N779);
buf BUF1 (N2706, N2702);
or OR2 (N2707, N2705, N633);
nand NAND2 (N2708, N2687, N1387);
buf BUF1 (N2709, N2707);
buf BUF1 (N2710, N2679);
nand NAND2 (N2711, N2686, N2383);
and AND4 (N2712, N2704, N2155, N277, N1480);
not NOT1 (N2713, N2694);
or OR4 (N2714, N2697, N2103, N1550, N986);
xor XOR2 (N2715, N2711, N975);
and AND3 (N2716, N2708, N1943, N1667);
nor NOR4 (N2717, N2713, N1095, N2127, N1829);
or OR4 (N2718, N2695, N2653, N1305, N936);
buf BUF1 (N2719, N2706);
nor NOR2 (N2720, N2714, N1782);
not NOT1 (N2721, N2717);
not NOT1 (N2722, N2703);
nor NOR4 (N2723, N2709, N698, N2416, N1610);
nor NOR4 (N2724, N2722, N187, N2179, N1185);
xor XOR2 (N2725, N2719, N2034);
and AND2 (N2726, N2724, N769);
and AND3 (N2727, N2712, N582, N2152);
and AND3 (N2728, N2723, N574, N1430);
nand NAND2 (N2729, N2726, N2411);
xor XOR2 (N2730, N2716, N2578);
or OR4 (N2731, N2729, N687, N2683, N1113);
buf BUF1 (N2732, N2728);
nand NAND3 (N2733, N2731, N376, N765);
and AND2 (N2734, N2721, N1262);
or OR3 (N2735, N2710, N1388, N867);
nand NAND3 (N2736, N2727, N1559, N433);
not NOT1 (N2737, N2720);
buf BUF1 (N2738, N2737);
or OR2 (N2739, N2735, N626);
nor NOR3 (N2740, N2736, N1196, N273);
nand NAND3 (N2741, N2734, N2391, N643);
nand NAND2 (N2742, N2718, N106);
not NOT1 (N2743, N2715);
nor NOR4 (N2744, N2733, N66, N1876, N201);
nor NOR4 (N2745, N2742, N115, N2279, N1277);
and AND3 (N2746, N2741, N66, N1390);
or OR4 (N2747, N2732, N661, N79, N1522);
and AND4 (N2748, N2738, N1974, N2608, N2259);
buf BUF1 (N2749, N2739);
xor XOR2 (N2750, N2744, N1006);
or OR4 (N2751, N2746, N62, N1175, N982);
nor NOR2 (N2752, N2730, N1988);
xor XOR2 (N2753, N2747, N472);
xor XOR2 (N2754, N2745, N2306);
xor XOR2 (N2755, N2740, N530);
or OR2 (N2756, N2749, N181);
nand NAND4 (N2757, N2754, N2590, N1965, N503);
xor XOR2 (N2758, N2748, N2704);
or OR4 (N2759, N2756, N873, N1049, N2595);
xor XOR2 (N2760, N2750, N163);
buf BUF1 (N2761, N2760);
or OR3 (N2762, N2759, N137, N900);
and AND2 (N2763, N2725, N2146);
and AND4 (N2764, N2758, N2720, N2190, N1719);
not NOT1 (N2765, N2752);
nor NOR4 (N2766, N2753, N1361, N550, N2489);
or OR3 (N2767, N2765, N2480, N2693);
nor NOR2 (N2768, N2763, N1463);
nor NOR4 (N2769, N2743, N1418, N1886, N2455);
and AND2 (N2770, N2761, N1068);
buf BUF1 (N2771, N2755);
buf BUF1 (N2772, N2751);
nor NOR3 (N2773, N2762, N2525, N1495);
nand NAND2 (N2774, N2757, N343);
xor XOR2 (N2775, N2769, N952);
and AND2 (N2776, N2771, N1552);
and AND3 (N2777, N2767, N1517, N2046);
xor XOR2 (N2778, N2777, N2483);
or OR4 (N2779, N2778, N1517, N1700, N1963);
xor XOR2 (N2780, N2768, N2137);
nor NOR2 (N2781, N2764, N120);
not NOT1 (N2782, N2780);
xor XOR2 (N2783, N2766, N315);
xor XOR2 (N2784, N2775, N347);
and AND3 (N2785, N2772, N275, N664);
nand NAND2 (N2786, N2776, N2426);
nor NOR4 (N2787, N2786, N1831, N1979, N1965);
nor NOR2 (N2788, N2781, N1381);
nand NAND2 (N2789, N2785, N1105);
and AND4 (N2790, N2774, N516, N756, N1506);
xor XOR2 (N2791, N2779, N1429);
nor NOR3 (N2792, N2789, N303, N636);
buf BUF1 (N2793, N2787);
xor XOR2 (N2794, N2773, N2756);
or OR3 (N2795, N2793, N2637, N1669);
buf BUF1 (N2796, N2792);
nand NAND4 (N2797, N2784, N1994, N2380, N38);
not NOT1 (N2798, N2770);
or OR2 (N2799, N2797, N2029);
not NOT1 (N2800, N2783);
or OR3 (N2801, N2800, N1365, N194);
and AND2 (N2802, N2796, N1624);
not NOT1 (N2803, N2802);
buf BUF1 (N2804, N2799);
or OR2 (N2805, N2794, N1032);
buf BUF1 (N2806, N2801);
nor NOR4 (N2807, N2788, N2458, N710, N2081);
buf BUF1 (N2808, N2791);
nand NAND4 (N2809, N2798, N1301, N519, N802);
and AND3 (N2810, N2803, N1144, N229);
nand NAND2 (N2811, N2804, N1691);
or OR4 (N2812, N2805, N1672, N422, N1295);
and AND3 (N2813, N2812, N269, N980);
buf BUF1 (N2814, N2807);
buf BUF1 (N2815, N2806);
or OR2 (N2816, N2814, N2563);
nor NOR2 (N2817, N2810, N2167);
nor NOR3 (N2818, N2813, N1888, N2384);
nor NOR4 (N2819, N2811, N379, N167, N2058);
and AND3 (N2820, N2816, N2080, N2175);
not NOT1 (N2821, N2795);
xor XOR2 (N2822, N2819, N1313);
and AND4 (N2823, N2817, N1499, N837, N504);
nand NAND2 (N2824, N2820, N37);
nand NAND3 (N2825, N2823, N1665, N1154);
nand NAND3 (N2826, N2824, N382, N2291);
not NOT1 (N2827, N2818);
or OR4 (N2828, N2815, N2548, N1437, N255);
and AND3 (N2829, N2808, N103, N580);
xor XOR2 (N2830, N2828, N936);
not NOT1 (N2831, N2826);
not NOT1 (N2832, N2782);
nor NOR2 (N2833, N2827, N128);
nand NAND3 (N2834, N2821, N177, N577);
xor XOR2 (N2835, N2790, N529);
nand NAND3 (N2836, N2825, N669, N1939);
not NOT1 (N2837, N2809);
not NOT1 (N2838, N2832);
not NOT1 (N2839, N2822);
nor NOR3 (N2840, N2831, N522, N1294);
or OR3 (N2841, N2829, N1662, N2453);
xor XOR2 (N2842, N2840, N1364);
and AND2 (N2843, N2833, N1832);
not NOT1 (N2844, N2834);
buf BUF1 (N2845, N2838);
nand NAND4 (N2846, N2843, N2573, N1910, N143);
xor XOR2 (N2847, N2835, N703);
xor XOR2 (N2848, N2847, N1252);
or OR3 (N2849, N2839, N2154, N1310);
xor XOR2 (N2850, N2837, N2552);
xor XOR2 (N2851, N2841, N2311);
and AND4 (N2852, N2842, N656, N1483, N781);
and AND3 (N2853, N2846, N2371, N486);
nand NAND3 (N2854, N2845, N560, N2161);
not NOT1 (N2855, N2850);
and AND2 (N2856, N2849, N2849);
nor NOR4 (N2857, N2836, N1804, N2330, N1862);
nand NAND3 (N2858, N2851, N2253, N1472);
nand NAND3 (N2859, N2854, N843, N2616);
nor NOR3 (N2860, N2844, N873, N1712);
not NOT1 (N2861, N2859);
not NOT1 (N2862, N2852);
not NOT1 (N2863, N2855);
and AND3 (N2864, N2862, N729, N2512);
nor NOR3 (N2865, N2864, N1594, N2701);
not NOT1 (N2866, N2857);
not NOT1 (N2867, N2865);
xor XOR2 (N2868, N2863, N2140);
not NOT1 (N2869, N2848);
or OR3 (N2870, N2856, N1358, N2225);
not NOT1 (N2871, N2869);
and AND4 (N2872, N2860, N1937, N898, N2486);
and AND3 (N2873, N2871, N2731, N864);
nor NOR4 (N2874, N2853, N2157, N1683, N1587);
buf BUF1 (N2875, N2858);
buf BUF1 (N2876, N2875);
nand NAND4 (N2877, N2867, N2552, N2341, N2130);
buf BUF1 (N2878, N2868);
buf BUF1 (N2879, N2866);
not NOT1 (N2880, N2876);
buf BUF1 (N2881, N2880);
or OR4 (N2882, N2870, N1476, N1230, N1237);
nor NOR2 (N2883, N2873, N2824);
not NOT1 (N2884, N2883);
xor XOR2 (N2885, N2882, N1003);
or OR2 (N2886, N2861, N2264);
or OR4 (N2887, N2874, N2129, N2581, N2579);
nand NAND3 (N2888, N2885, N2224, N1227);
nor NOR2 (N2889, N2887, N169);
xor XOR2 (N2890, N2881, N2608);
or OR4 (N2891, N2889, N1741, N2219, N1784);
nand NAND2 (N2892, N2890, N1290);
and AND2 (N2893, N2877, N1705);
not NOT1 (N2894, N2893);
nand NAND3 (N2895, N2886, N2339, N2455);
xor XOR2 (N2896, N2892, N157);
and AND3 (N2897, N2894, N1983, N758);
nor NOR4 (N2898, N2830, N2471, N2292, N1799);
not NOT1 (N2899, N2884);
nor NOR4 (N2900, N2896, N2666, N453, N995);
not NOT1 (N2901, N2900);
buf BUF1 (N2902, N2878);
nor NOR3 (N2903, N2888, N2886, N558);
not NOT1 (N2904, N2901);
xor XOR2 (N2905, N2891, N2228);
nor NOR2 (N2906, N2879, N1457);
and AND3 (N2907, N2898, N2408, N2247);
xor XOR2 (N2908, N2897, N2468);
xor XOR2 (N2909, N2899, N443);
buf BUF1 (N2910, N2908);
or OR3 (N2911, N2872, N2713, N2383);
xor XOR2 (N2912, N2906, N2899);
and AND2 (N2913, N2895, N2283);
nor NOR2 (N2914, N2912, N2629);
and AND2 (N2915, N2902, N885);
buf BUF1 (N2916, N2905);
not NOT1 (N2917, N2907);
or OR4 (N2918, N2917, N2571, N1139, N211);
not NOT1 (N2919, N2904);
and AND3 (N2920, N2909, N1848, N886);
nand NAND3 (N2921, N2918, N2039, N2425);
nor NOR3 (N2922, N2903, N1017, N2009);
and AND3 (N2923, N2921, N1064, N382);
nor NOR4 (N2924, N2923, N2244, N2221, N2413);
or OR2 (N2925, N2915, N2124);
nor NOR4 (N2926, N2913, N1253, N2866, N2617);
xor XOR2 (N2927, N2920, N1395);
nor NOR4 (N2928, N2925, N917, N1139, N2470);
or OR4 (N2929, N2916, N280, N605, N1636);
buf BUF1 (N2930, N2927);
nand NAND2 (N2931, N2930, N2423);
or OR4 (N2932, N2910, N1639, N2494, N2005);
or OR4 (N2933, N2911, N1548, N1402, N1466);
xor XOR2 (N2934, N2924, N2018);
xor XOR2 (N2935, N2914, N1430);
nor NOR4 (N2936, N2932, N835, N412, N595);
not NOT1 (N2937, N2935);
not NOT1 (N2938, N2931);
and AND3 (N2939, N2934, N273, N1118);
xor XOR2 (N2940, N2937, N1578);
nor NOR4 (N2941, N2939, N2734, N2834, N1819);
not NOT1 (N2942, N2922);
or OR3 (N2943, N2928, N2036, N2830);
not NOT1 (N2944, N2941);
xor XOR2 (N2945, N2926, N729);
nor NOR4 (N2946, N2919, N844, N1960, N2404);
nor NOR4 (N2947, N2929, N2579, N1384, N167);
nand NAND4 (N2948, N2933, N1304, N645, N94);
nor NOR2 (N2949, N2945, N530);
and AND4 (N2950, N2944, N1839, N1115, N1672);
nand NAND4 (N2951, N2940, N1170, N1464, N2901);
and AND4 (N2952, N2942, N366, N967, N1843);
xor XOR2 (N2953, N2952, N275);
nand NAND3 (N2954, N2950, N1393, N1881);
nand NAND3 (N2955, N2946, N275, N1031);
buf BUF1 (N2956, N2948);
nand NAND4 (N2957, N2956, N2038, N2163, N2692);
and AND4 (N2958, N2954, N1816, N92, N2595);
xor XOR2 (N2959, N2943, N1599);
buf BUF1 (N2960, N2953);
xor XOR2 (N2961, N2960, N1863);
nand NAND4 (N2962, N2961, N1441, N460, N417);
buf BUF1 (N2963, N2938);
and AND3 (N2964, N2951, N879, N2775);
and AND4 (N2965, N2936, N2759, N2344, N2811);
or OR4 (N2966, N2959, N2783, N722, N2837);
nand NAND3 (N2967, N2962, N1505, N1311);
xor XOR2 (N2968, N2957, N1141);
not NOT1 (N2969, N2958);
buf BUF1 (N2970, N2955);
nor NOR3 (N2971, N2970, N2703, N1947);
not NOT1 (N2972, N2947);
and AND2 (N2973, N2965, N1035);
nor NOR3 (N2974, N2972, N1239, N2186);
xor XOR2 (N2975, N2973, N2317);
not NOT1 (N2976, N2949);
nand NAND3 (N2977, N2974, N2650, N151);
and AND4 (N2978, N2967, N1599, N855, N947);
nand NAND2 (N2979, N2975, N1029);
buf BUF1 (N2980, N2964);
or OR4 (N2981, N2977, N2359, N1609, N954);
and AND4 (N2982, N2969, N139, N2935, N1100);
nor NOR3 (N2983, N2980, N803, N1121);
and AND3 (N2984, N2963, N72, N2222);
and AND2 (N2985, N2976, N246);
xor XOR2 (N2986, N2983, N766);
not NOT1 (N2987, N2986);
or OR4 (N2988, N2978, N1260, N2194, N2504);
not NOT1 (N2989, N2981);
buf BUF1 (N2990, N2971);
and AND3 (N2991, N2968, N347, N977);
nand NAND4 (N2992, N2989, N2923, N1393, N2224);
nor NOR3 (N2993, N2991, N525, N987);
or OR2 (N2994, N2987, N98);
nand NAND3 (N2995, N2994, N1903, N2322);
nor NOR4 (N2996, N2985, N311, N2006, N560);
and AND2 (N2997, N2990, N1456);
buf BUF1 (N2998, N2988);
nor NOR3 (N2999, N2996, N97, N1008);
not NOT1 (N3000, N2984);
and AND4 (N3001, N2966, N2560, N576, N2378);
not NOT1 (N3002, N2998);
nand NAND4 (N3003, N2979, N1821, N2964, N2956);
xor XOR2 (N3004, N2992, N1323);
nand NAND2 (N3005, N3001, N2915);
or OR3 (N3006, N2993, N1536, N2029);
xor XOR2 (N3007, N3005, N37);
and AND2 (N3008, N3006, N1267);
nor NOR3 (N3009, N3007, N2232, N1883);
not NOT1 (N3010, N3000);
nor NOR4 (N3011, N2997, N1527, N768, N2452);
not NOT1 (N3012, N2982);
not NOT1 (N3013, N3009);
nor NOR4 (N3014, N3003, N1347, N2597, N1134);
nand NAND3 (N3015, N3004, N1504, N699);
xor XOR2 (N3016, N2999, N2381);
nor NOR4 (N3017, N2995, N1980, N2061, N1979);
or OR4 (N3018, N3010, N749, N1347, N2172);
endmodule