// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;

output N6396,N6409,N6413,N6405,N6411,N6404,N6407,N6408,N6397,N6415;

not NOT1 (N16, N10);
or OR4 (N17, N15, N16, N8, N10);
nor NOR3 (N18, N16, N11, N10);
nand NAND2 (N19, N8, N4);
or OR4 (N20, N11, N10, N1, N15);
buf BUF1 (N21, N7);
not NOT1 (N22, N5);
and AND4 (N23, N9, N2, N19, N10);
nor NOR4 (N24, N13, N9, N3, N21);
or OR2 (N25, N22, N20);
not NOT1 (N26, N8);
or OR3 (N27, N19, N25, N6);
nor NOR4 (N28, N25, N11, N22, N14);
nand NAND4 (N29, N21, N19, N1, N26);
nand NAND2 (N30, N6, N28);
buf BUF1 (N31, N15);
not NOT1 (N32, N26);
or OR3 (N33, N1, N17, N14);
nand NAND2 (N34, N2, N29);
nor NOR2 (N35, N29, N18);
nor NOR3 (N36, N29, N21, N3);
nor NOR2 (N37, N35, N11);
nor NOR3 (N38, N37, N32, N36);
and AND3 (N39, N3, N35, N21);
nor NOR3 (N40, N4, N25, N4);
nor NOR2 (N41, N34, N40);
buf BUF1 (N42, N23);
nand NAND3 (N43, N26, N13, N22);
not NOT1 (N44, N33);
buf BUF1 (N45, N42);
and AND4 (N46, N30, N6, N33, N34);
and AND2 (N47, N38, N43);
xor XOR2 (N48, N45, N1);
nor NOR2 (N49, N35, N30);
not NOT1 (N50, N49);
and AND2 (N51, N41, N32);
xor XOR2 (N52, N48, N8);
buf BUF1 (N53, N47);
nand NAND2 (N54, N51, N39);
nor NOR3 (N55, N47, N23, N48);
or OR3 (N56, N27, N36, N3);
not NOT1 (N57, N46);
buf BUF1 (N58, N57);
xor XOR2 (N59, N53, N7);
nor NOR2 (N60, N58, N17);
nor NOR4 (N61, N54, N34, N40, N32);
and AND2 (N62, N55, N30);
nor NOR2 (N63, N31, N15);
or OR2 (N64, N44, N35);
buf BUF1 (N65, N24);
xor XOR2 (N66, N64, N27);
nand NAND3 (N67, N65, N44, N10);
buf BUF1 (N68, N66);
not NOT1 (N69, N59);
xor XOR2 (N70, N56, N31);
nor NOR3 (N71, N50, N48, N20);
or OR2 (N72, N63, N13);
nand NAND2 (N73, N72, N4);
xor XOR2 (N74, N60, N14);
nor NOR4 (N75, N71, N48, N69, N28);
xor XOR2 (N76, N38, N63);
and AND2 (N77, N61, N28);
xor XOR2 (N78, N74, N40);
nor NOR2 (N79, N78, N35);
and AND3 (N80, N76, N72, N73);
nor NOR4 (N81, N52, N69, N19, N32);
not NOT1 (N82, N70);
and AND3 (N83, N56, N69, N27);
not NOT1 (N84, N81);
not NOT1 (N85, N84);
not NOT1 (N86, N77);
xor XOR2 (N87, N67, N51);
buf BUF1 (N88, N80);
not NOT1 (N89, N87);
not NOT1 (N90, N79);
or OR4 (N91, N68, N21, N30, N45);
and AND4 (N92, N90, N89, N13, N30);
xor XOR2 (N93, N54, N64);
nand NAND2 (N94, N85, N51);
nand NAND4 (N95, N91, N77, N58, N49);
not NOT1 (N96, N95);
nor NOR2 (N97, N94, N3);
not NOT1 (N98, N62);
not NOT1 (N99, N92);
or OR3 (N100, N75, N83, N82);
buf BUF1 (N101, N39);
not NOT1 (N102, N56);
nand NAND3 (N103, N96, N27, N79);
not NOT1 (N104, N98);
buf BUF1 (N105, N93);
buf BUF1 (N106, N102);
xor XOR2 (N107, N97, N13);
not NOT1 (N108, N99);
or OR3 (N109, N100, N2, N32);
and AND4 (N110, N108, N30, N95, N48);
nand NAND4 (N111, N105, N48, N20, N27);
and AND3 (N112, N107, N52, N75);
buf BUF1 (N113, N106);
buf BUF1 (N114, N101);
not NOT1 (N115, N110);
xor XOR2 (N116, N115, N20);
or OR2 (N117, N116, N97);
not NOT1 (N118, N113);
nor NOR3 (N119, N114, N20, N79);
or OR3 (N120, N104, N19, N61);
buf BUF1 (N121, N120);
or OR2 (N122, N119, N82);
nor NOR2 (N123, N109, N84);
and AND4 (N124, N122, N75, N24, N62);
nand NAND3 (N125, N103, N100, N73);
or OR4 (N126, N121, N112, N68, N73);
buf BUF1 (N127, N46);
nor NOR4 (N128, N123, N51, N49, N95);
not NOT1 (N129, N117);
not NOT1 (N130, N111);
not NOT1 (N131, N126);
nor NOR3 (N132, N125, N111, N4);
xor XOR2 (N133, N127, N132);
and AND4 (N134, N90, N52, N116, N76);
or OR2 (N135, N128, N15);
xor XOR2 (N136, N88, N91);
not NOT1 (N137, N135);
nand NAND3 (N138, N134, N17, N3);
nor NOR2 (N139, N136, N8);
buf BUF1 (N140, N139);
buf BUF1 (N141, N140);
not NOT1 (N142, N141);
buf BUF1 (N143, N118);
nor NOR2 (N144, N142, N37);
nand NAND3 (N145, N143, N30, N118);
or OR4 (N146, N133, N117, N63, N83);
nand NAND4 (N147, N129, N52, N63, N122);
nor NOR4 (N148, N146, N106, N9, N75);
nand NAND2 (N149, N138, N36);
nand NAND4 (N150, N124, N146, N87, N111);
or OR4 (N151, N144, N141, N100, N29);
xor XOR2 (N152, N137, N58);
xor XOR2 (N153, N147, N94);
or OR3 (N154, N86, N7, N57);
or OR3 (N155, N152, N152, N123);
xor XOR2 (N156, N153, N149);
buf BUF1 (N157, N105);
or OR2 (N158, N156, N12);
xor XOR2 (N159, N154, N79);
or OR4 (N160, N148, N26, N47, N93);
not NOT1 (N161, N157);
and AND4 (N162, N160, N32, N150, N50);
buf BUF1 (N163, N94);
or OR3 (N164, N131, N107, N81);
xor XOR2 (N165, N151, N156);
and AND3 (N166, N155, N63, N155);
not NOT1 (N167, N159);
nor NOR4 (N168, N145, N158, N124, N75);
or OR4 (N169, N17, N122, N130, N81);
not NOT1 (N170, N147);
and AND3 (N171, N168, N97, N3);
nand NAND3 (N172, N161, N50, N28);
buf BUF1 (N173, N166);
buf BUF1 (N174, N171);
nor NOR4 (N175, N167, N174, N7, N90);
or OR4 (N176, N144, N79, N100, N49);
nand NAND2 (N177, N162, N11);
nor NOR2 (N178, N165, N78);
nand NAND2 (N179, N172, N87);
nor NOR3 (N180, N175, N85, N72);
and AND3 (N181, N173, N130, N131);
nand NAND2 (N182, N170, N72);
nor NOR4 (N183, N169, N73, N16, N104);
xor XOR2 (N184, N163, N168);
and AND4 (N185, N178, N110, N72, N174);
buf BUF1 (N186, N180);
or OR2 (N187, N179, N124);
not NOT1 (N188, N181);
or OR3 (N189, N177, N21, N93);
and AND4 (N190, N184, N31, N35, N153);
nor NOR3 (N191, N176, N19, N168);
buf BUF1 (N192, N164);
and AND2 (N193, N191, N71);
and AND3 (N194, N193, N60, N62);
nand NAND4 (N195, N194, N154, N121, N19);
or OR3 (N196, N183, N34, N168);
not NOT1 (N197, N187);
not NOT1 (N198, N190);
buf BUF1 (N199, N185);
buf BUF1 (N200, N186);
xor XOR2 (N201, N189, N81);
or OR2 (N202, N201, N37);
and AND4 (N203, N202, N201, N74, N197);
nand NAND3 (N204, N173, N75, N193);
and AND4 (N205, N196, N149, N37, N27);
or OR3 (N206, N205, N41, N111);
or OR3 (N207, N198, N190, N72);
xor XOR2 (N208, N207, N78);
nand NAND4 (N209, N195, N75, N9, N5);
not NOT1 (N210, N182);
and AND2 (N211, N209, N151);
buf BUF1 (N212, N208);
nand NAND2 (N213, N200, N4);
or OR3 (N214, N211, N160, N79);
nand NAND4 (N215, N192, N96, N28, N24);
nor NOR2 (N216, N213, N24);
not NOT1 (N217, N215);
not NOT1 (N218, N206);
and AND2 (N219, N218, N168);
or OR2 (N220, N214, N97);
nor NOR3 (N221, N204, N17, N143);
not NOT1 (N222, N219);
nand NAND3 (N223, N216, N214, N214);
or OR3 (N224, N210, N118, N31);
or OR3 (N225, N221, N94, N194);
not NOT1 (N226, N199);
nand NAND2 (N227, N224, N216);
nor NOR2 (N228, N222, N101);
not NOT1 (N229, N226);
and AND2 (N230, N203, N94);
buf BUF1 (N231, N223);
xor XOR2 (N232, N228, N120);
or OR4 (N233, N231, N25, N67, N73);
nand NAND3 (N234, N188, N183, N10);
or OR3 (N235, N230, N156, N111);
xor XOR2 (N236, N212, N187);
not NOT1 (N237, N236);
xor XOR2 (N238, N217, N32);
nor NOR3 (N239, N225, N195, N90);
buf BUF1 (N240, N229);
nand NAND3 (N241, N239, N123, N138);
nor NOR4 (N242, N238, N84, N55, N218);
nand NAND3 (N243, N234, N193, N87);
not NOT1 (N244, N220);
not NOT1 (N245, N233);
nor NOR2 (N246, N241, N162);
and AND4 (N247, N242, N144, N114, N228);
or OR4 (N248, N227, N221, N211, N121);
xor XOR2 (N249, N246, N236);
nor NOR3 (N250, N232, N232, N126);
or OR2 (N251, N243, N135);
and AND2 (N252, N248, N242);
xor XOR2 (N253, N245, N163);
or OR2 (N254, N252, N76);
not NOT1 (N255, N237);
xor XOR2 (N256, N244, N159);
xor XOR2 (N257, N255, N21);
nor NOR4 (N258, N256, N212, N98, N248);
and AND3 (N259, N249, N251, N5);
not NOT1 (N260, N35);
nor NOR3 (N261, N260, N81, N209);
or OR4 (N262, N235, N59, N174, N208);
nor NOR4 (N263, N261, N49, N139, N196);
buf BUF1 (N264, N254);
xor XOR2 (N265, N250, N135);
or OR2 (N266, N264, N260);
or OR2 (N267, N263, N144);
nor NOR3 (N268, N259, N94, N138);
not NOT1 (N269, N266);
xor XOR2 (N270, N253, N216);
or OR2 (N271, N257, N237);
nor NOR3 (N272, N268, N105, N77);
or OR2 (N273, N269, N99);
nor NOR3 (N274, N272, N59, N182);
xor XOR2 (N275, N240, N130);
buf BUF1 (N276, N275);
buf BUF1 (N277, N274);
not NOT1 (N278, N277);
or OR2 (N279, N270, N79);
nor NOR2 (N280, N265, N198);
and AND3 (N281, N276, N90, N11);
buf BUF1 (N282, N267);
nor NOR2 (N283, N280, N256);
buf BUF1 (N284, N262);
nand NAND2 (N285, N247, N122);
buf BUF1 (N286, N279);
and AND4 (N287, N271, N187, N71, N155);
buf BUF1 (N288, N281);
buf BUF1 (N289, N278);
or OR4 (N290, N289, N275, N70, N50);
nor NOR2 (N291, N285, N175);
nand NAND3 (N292, N284, N225, N58);
or OR4 (N293, N287, N99, N182, N19);
or OR2 (N294, N293, N138);
nor NOR3 (N295, N273, N193, N22);
and AND2 (N296, N294, N205);
nor NOR4 (N297, N292, N167, N185, N294);
nor NOR2 (N298, N295, N104);
buf BUF1 (N299, N290);
not NOT1 (N300, N296);
xor XOR2 (N301, N300, N181);
xor XOR2 (N302, N258, N128);
nor NOR3 (N303, N297, N53, N94);
xor XOR2 (N304, N301, N270);
xor XOR2 (N305, N302, N294);
nor NOR2 (N306, N305, N45);
nor NOR2 (N307, N306, N4);
or OR3 (N308, N307, N58, N227);
or OR3 (N309, N286, N113, N285);
and AND2 (N310, N299, N45);
nand NAND3 (N311, N282, N281, N262);
not NOT1 (N312, N288);
not NOT1 (N313, N311);
not NOT1 (N314, N310);
xor XOR2 (N315, N298, N178);
nand NAND4 (N316, N315, N197, N52, N19);
or OR4 (N317, N304, N196, N193, N292);
and AND2 (N318, N309, N5);
not NOT1 (N319, N283);
nand NAND2 (N320, N314, N30);
nor NOR2 (N321, N320, N106);
not NOT1 (N322, N318);
and AND3 (N323, N312, N284, N150);
buf BUF1 (N324, N313);
buf BUF1 (N325, N303);
not NOT1 (N326, N323);
and AND3 (N327, N322, N8, N173);
nor NOR3 (N328, N327, N5, N273);
nand NAND3 (N329, N291, N308, N280);
buf BUF1 (N330, N18);
not NOT1 (N331, N329);
buf BUF1 (N332, N316);
and AND3 (N333, N328, N6, N167);
buf BUF1 (N334, N319);
xor XOR2 (N335, N324, N73);
not NOT1 (N336, N330);
not NOT1 (N337, N331);
nand NAND2 (N338, N326, N231);
nor NOR3 (N339, N317, N317, N242);
and AND2 (N340, N338, N15);
not NOT1 (N341, N337);
buf BUF1 (N342, N334);
not NOT1 (N343, N325);
nor NOR3 (N344, N335, N224, N48);
nor NOR3 (N345, N332, N32, N71);
nor NOR3 (N346, N333, N235, N292);
and AND4 (N347, N346, N10, N71, N233);
buf BUF1 (N348, N347);
xor XOR2 (N349, N336, N184);
and AND3 (N350, N345, N123, N215);
or OR2 (N351, N343, N3);
and AND2 (N352, N344, N290);
not NOT1 (N353, N349);
and AND3 (N354, N321, N303, N60);
and AND2 (N355, N340, N226);
not NOT1 (N356, N348);
nor NOR3 (N357, N342, N245, N295);
nor NOR4 (N358, N350, N215, N137, N239);
nand NAND2 (N359, N352, N15);
buf BUF1 (N360, N358);
and AND2 (N361, N359, N70);
or OR2 (N362, N353, N138);
not NOT1 (N363, N360);
or OR2 (N364, N339, N258);
and AND4 (N365, N361, N338, N311, N150);
nand NAND4 (N366, N356, N84, N297, N269);
nand NAND3 (N367, N351, N164, N341);
or OR4 (N368, N185, N113, N358, N164);
and AND2 (N369, N367, N107);
and AND3 (N370, N362, N302, N13);
buf BUF1 (N371, N370);
not NOT1 (N372, N368);
xor XOR2 (N373, N364, N132);
buf BUF1 (N374, N369);
or OR4 (N375, N365, N55, N25, N198);
xor XOR2 (N376, N354, N12);
and AND3 (N377, N375, N362, N177);
and AND2 (N378, N357, N239);
and AND4 (N379, N372, N374, N275, N363);
nand NAND2 (N380, N173, N27);
not NOT1 (N381, N3);
not NOT1 (N382, N373);
not NOT1 (N383, N381);
and AND4 (N384, N355, N142, N118, N179);
buf BUF1 (N385, N382);
and AND2 (N386, N371, N340);
not NOT1 (N387, N366);
not NOT1 (N388, N376);
and AND2 (N389, N380, N221);
nor NOR2 (N390, N377, N388);
buf BUF1 (N391, N46);
nor NOR2 (N392, N378, N118);
or OR4 (N393, N391, N41, N236, N186);
buf BUF1 (N394, N389);
nor NOR4 (N395, N390, N341, N340, N62);
xor XOR2 (N396, N394, N124);
not NOT1 (N397, N393);
xor XOR2 (N398, N397, N74);
xor XOR2 (N399, N385, N111);
buf BUF1 (N400, N386);
not NOT1 (N401, N383);
or OR4 (N402, N398, N183, N258, N206);
xor XOR2 (N403, N401, N297);
and AND4 (N404, N396, N151, N277, N354);
and AND4 (N405, N400, N126, N169, N270);
and AND3 (N406, N402, N331, N80);
not NOT1 (N407, N399);
buf BUF1 (N408, N407);
xor XOR2 (N409, N392, N145);
or OR2 (N410, N387, N208);
nand NAND3 (N411, N403, N62, N283);
nor NOR4 (N412, N409, N381, N95, N201);
nand NAND4 (N413, N406, N412, N357, N2);
nand NAND2 (N414, N72, N280);
buf BUF1 (N415, N414);
nand NAND2 (N416, N415, N402);
nand NAND3 (N417, N384, N49, N387);
buf BUF1 (N418, N404);
not NOT1 (N419, N416);
or OR2 (N420, N405, N122);
and AND3 (N421, N410, N30, N214);
nand NAND4 (N422, N411, N300, N170, N377);
xor XOR2 (N423, N395, N135);
not NOT1 (N424, N420);
nor NOR2 (N425, N408, N246);
nor NOR3 (N426, N417, N22, N121);
not NOT1 (N427, N422);
nor NOR4 (N428, N421, N129, N394, N290);
not NOT1 (N429, N424);
not NOT1 (N430, N426);
or OR4 (N431, N413, N14, N301, N322);
and AND3 (N432, N430, N420, N179);
not NOT1 (N433, N425);
or OR2 (N434, N379, N19);
or OR4 (N435, N431, N367, N303, N34);
not NOT1 (N436, N419);
buf BUF1 (N437, N418);
nor NOR4 (N438, N434, N411, N314, N8);
nand NAND4 (N439, N438, N86, N171, N264);
xor XOR2 (N440, N436, N253);
or OR3 (N441, N439, N165, N397);
nor NOR4 (N442, N432, N345, N255, N54);
buf BUF1 (N443, N435);
or OR2 (N444, N437, N352);
xor XOR2 (N445, N444, N259);
nand NAND3 (N446, N440, N85, N139);
not NOT1 (N447, N423);
and AND4 (N448, N445, N429, N147, N343);
nor NOR2 (N449, N339, N141);
nand NAND3 (N450, N442, N319, N339);
xor XOR2 (N451, N441, N203);
xor XOR2 (N452, N448, N426);
nor NOR3 (N453, N447, N280, N271);
nor NOR3 (N454, N427, N398, N11);
not NOT1 (N455, N446);
and AND3 (N456, N428, N32, N352);
or OR3 (N457, N452, N17, N26);
nor NOR3 (N458, N454, N181, N151);
buf BUF1 (N459, N457);
nand NAND3 (N460, N450, N450, N244);
buf BUF1 (N461, N451);
nand NAND3 (N462, N459, N444, N145);
and AND2 (N463, N460, N204);
or OR3 (N464, N456, N354, N124);
and AND3 (N465, N462, N349, N163);
xor XOR2 (N466, N463, N222);
xor XOR2 (N467, N443, N270);
and AND2 (N468, N449, N324);
and AND2 (N469, N453, N245);
not NOT1 (N470, N458);
or OR2 (N471, N467, N289);
nor NOR4 (N472, N471, N446, N147, N362);
buf BUF1 (N473, N469);
or OR3 (N474, N473, N136, N17);
and AND4 (N475, N465, N155, N212, N406);
not NOT1 (N476, N464);
nor NOR4 (N477, N455, N316, N392, N79);
nand NAND3 (N478, N433, N256, N74);
nor NOR2 (N479, N477, N157);
not NOT1 (N480, N466);
buf BUF1 (N481, N480);
nor NOR2 (N482, N478, N2);
xor XOR2 (N483, N474, N376);
not NOT1 (N484, N479);
nand NAND2 (N485, N468, N475);
buf BUF1 (N486, N345);
not NOT1 (N487, N486);
xor XOR2 (N488, N470, N330);
or OR4 (N489, N476, N184, N356, N117);
not NOT1 (N490, N481);
nor NOR3 (N491, N483, N417, N138);
buf BUF1 (N492, N491);
xor XOR2 (N493, N488, N344);
or OR2 (N494, N461, N264);
or OR3 (N495, N490, N296, N349);
xor XOR2 (N496, N493, N300);
and AND3 (N497, N484, N407, N13);
or OR2 (N498, N497, N137);
nor NOR2 (N499, N472, N378);
buf BUF1 (N500, N495);
nand NAND4 (N501, N498, N284, N372, N259);
not NOT1 (N502, N496);
or OR3 (N503, N492, N194, N91);
and AND2 (N504, N485, N342);
xor XOR2 (N505, N500, N118);
and AND4 (N506, N499, N259, N172, N367);
xor XOR2 (N507, N494, N356);
or OR2 (N508, N505, N237);
nor NOR3 (N509, N502, N201, N480);
not NOT1 (N510, N506);
not NOT1 (N511, N501);
not NOT1 (N512, N482);
xor XOR2 (N513, N487, N236);
or OR3 (N514, N504, N492, N321);
nor NOR2 (N515, N509, N481);
nand NAND3 (N516, N503, N103, N285);
nand NAND3 (N517, N512, N494, N442);
not NOT1 (N518, N516);
not NOT1 (N519, N517);
xor XOR2 (N520, N508, N65);
buf BUF1 (N521, N519);
not NOT1 (N522, N510);
buf BUF1 (N523, N520);
xor XOR2 (N524, N514, N263);
or OR4 (N525, N524, N10, N187, N356);
or OR4 (N526, N513, N308, N400, N407);
buf BUF1 (N527, N526);
buf BUF1 (N528, N521);
not NOT1 (N529, N515);
nor NOR2 (N530, N523, N86);
nand NAND3 (N531, N525, N155, N195);
nor NOR2 (N532, N507, N41);
not NOT1 (N533, N511);
xor XOR2 (N534, N533, N82);
nor NOR3 (N535, N518, N81, N21);
nand NAND3 (N536, N522, N326, N196);
or OR2 (N537, N530, N172);
nor NOR3 (N538, N537, N228, N363);
xor XOR2 (N539, N529, N405);
not NOT1 (N540, N528);
nor NOR3 (N541, N538, N12, N30);
not NOT1 (N542, N536);
buf BUF1 (N543, N541);
nor NOR4 (N544, N535, N303, N205, N153);
not NOT1 (N545, N539);
buf BUF1 (N546, N527);
nor NOR3 (N547, N489, N196, N480);
not NOT1 (N548, N532);
nor NOR4 (N549, N548, N4, N520, N394);
xor XOR2 (N550, N534, N359);
not NOT1 (N551, N546);
and AND4 (N552, N531, N483, N442, N175);
buf BUF1 (N553, N540);
nor NOR3 (N554, N543, N525, N520);
and AND3 (N555, N554, N177, N531);
nor NOR4 (N556, N549, N312, N47, N311);
nor NOR2 (N557, N556, N373);
xor XOR2 (N558, N545, N223);
and AND3 (N559, N542, N438, N227);
nand NAND4 (N560, N553, N121, N461, N377);
or OR4 (N561, N551, N17, N87, N376);
or OR3 (N562, N552, N480, N351);
or OR3 (N563, N557, N176, N489);
nand NAND4 (N564, N563, N467, N396, N448);
nand NAND3 (N565, N564, N286, N496);
buf BUF1 (N566, N565);
or OR4 (N567, N555, N224, N88, N396);
not NOT1 (N568, N550);
and AND3 (N569, N561, N172, N66);
nand NAND2 (N570, N566, N298);
and AND2 (N571, N558, N116);
not NOT1 (N572, N559);
xor XOR2 (N573, N544, N323);
or OR2 (N574, N570, N493);
not NOT1 (N575, N547);
not NOT1 (N576, N562);
nand NAND4 (N577, N575, N196, N568, N238);
not NOT1 (N578, N360);
or OR4 (N579, N574, N106, N43, N369);
or OR2 (N580, N579, N186);
buf BUF1 (N581, N580);
or OR3 (N582, N571, N169, N483);
and AND4 (N583, N572, N322, N323, N73);
nand NAND2 (N584, N567, N415);
nand NAND4 (N585, N578, N25, N583, N135);
and AND4 (N586, N570, N375, N27, N450);
buf BUF1 (N587, N584);
not NOT1 (N588, N587);
nor NOR2 (N589, N569, N539);
buf BUF1 (N590, N588);
xor XOR2 (N591, N590, N120);
xor XOR2 (N592, N577, N546);
not NOT1 (N593, N560);
and AND2 (N594, N582, N334);
not NOT1 (N595, N592);
xor XOR2 (N596, N595, N345);
not NOT1 (N597, N591);
buf BUF1 (N598, N585);
nor NOR2 (N599, N573, N253);
buf BUF1 (N600, N596);
nand NAND3 (N601, N600, N241, N447);
and AND3 (N602, N581, N22, N152);
nand NAND3 (N603, N594, N343, N431);
buf BUF1 (N604, N601);
xor XOR2 (N605, N589, N204);
or OR3 (N606, N599, N584, N451);
not NOT1 (N607, N606);
buf BUF1 (N608, N607);
not NOT1 (N609, N576);
not NOT1 (N610, N586);
xor XOR2 (N611, N603, N92);
and AND3 (N612, N610, N571, N272);
xor XOR2 (N613, N598, N332);
or OR3 (N614, N593, N376, N194);
and AND4 (N615, N609, N332, N376, N330);
xor XOR2 (N616, N612, N135);
and AND4 (N617, N615, N401, N482, N266);
nand NAND4 (N618, N613, N478, N49, N106);
and AND3 (N619, N608, N494, N184);
or OR3 (N620, N605, N492, N579);
not NOT1 (N621, N604);
nand NAND2 (N622, N621, N344);
xor XOR2 (N623, N618, N257);
or OR2 (N624, N622, N283);
xor XOR2 (N625, N623, N286);
nand NAND3 (N626, N611, N571, N104);
or OR4 (N627, N625, N32, N582, N394);
xor XOR2 (N628, N626, N102);
or OR4 (N629, N620, N177, N240, N119);
and AND4 (N630, N617, N391, N434, N359);
not NOT1 (N631, N629);
or OR4 (N632, N619, N298, N359, N565);
and AND2 (N633, N614, N321);
xor XOR2 (N634, N616, N37);
nor NOR2 (N635, N628, N249);
buf BUF1 (N636, N632);
nand NAND4 (N637, N635, N133, N409, N253);
nand NAND4 (N638, N636, N617, N607, N500);
buf BUF1 (N639, N637);
xor XOR2 (N640, N627, N495);
nor NOR3 (N641, N634, N539, N624);
buf BUF1 (N642, N492);
buf BUF1 (N643, N597);
nand NAND3 (N644, N633, N267, N289);
nor NOR2 (N645, N639, N233);
buf BUF1 (N646, N631);
nand NAND4 (N647, N643, N422, N295, N463);
nor NOR3 (N648, N641, N431, N267);
or OR4 (N649, N602, N179, N471, N155);
nor NOR2 (N650, N638, N625);
xor XOR2 (N651, N647, N127);
nand NAND3 (N652, N645, N117, N552);
or OR4 (N653, N644, N494, N413, N535);
or OR4 (N654, N649, N354, N650, N311);
nand NAND3 (N655, N558, N372, N44);
nor NOR2 (N656, N651, N525);
nand NAND2 (N657, N654, N602);
nor NOR2 (N658, N657, N481);
nor NOR2 (N659, N640, N567);
and AND2 (N660, N656, N155);
or OR2 (N661, N648, N462);
nor NOR2 (N662, N658, N526);
not NOT1 (N663, N646);
nor NOR3 (N664, N652, N24, N648);
nor NOR4 (N665, N660, N260, N417, N453);
and AND4 (N666, N665, N76, N652, N300);
xor XOR2 (N667, N661, N629);
nand NAND3 (N668, N667, N498, N550);
not NOT1 (N669, N642);
and AND3 (N670, N655, N276, N88);
nand NAND3 (N671, N668, N413, N661);
xor XOR2 (N672, N662, N264);
nor NOR4 (N673, N630, N136, N593, N76);
not NOT1 (N674, N669);
buf BUF1 (N675, N666);
buf BUF1 (N676, N673);
buf BUF1 (N677, N676);
and AND3 (N678, N670, N99, N53);
and AND4 (N679, N671, N430, N121, N322);
and AND4 (N680, N653, N189, N362, N246);
or OR4 (N681, N674, N291, N187, N332);
nor NOR2 (N682, N672, N1);
nand NAND3 (N683, N681, N645, N458);
buf BUF1 (N684, N680);
or OR4 (N685, N683, N92, N163, N54);
and AND3 (N686, N663, N300, N494);
xor XOR2 (N687, N679, N417);
and AND2 (N688, N684, N213);
nor NOR3 (N689, N664, N93, N479);
nor NOR4 (N690, N659, N632, N653, N484);
or OR2 (N691, N682, N293);
or OR2 (N692, N689, N441);
buf BUF1 (N693, N687);
nor NOR3 (N694, N693, N175, N70);
or OR3 (N695, N686, N402, N428);
nor NOR2 (N696, N688, N148);
or OR3 (N697, N685, N183, N271);
not NOT1 (N698, N678);
nand NAND3 (N699, N691, N481, N337);
nor NOR2 (N700, N695, N65);
or OR2 (N701, N699, N269);
buf BUF1 (N702, N692);
xor XOR2 (N703, N702, N129);
nand NAND4 (N704, N698, N117, N30, N391);
buf BUF1 (N705, N696);
nand NAND3 (N706, N704, N437, N208);
or OR2 (N707, N697, N165);
buf BUF1 (N708, N706);
not NOT1 (N709, N708);
xor XOR2 (N710, N694, N164);
nor NOR3 (N711, N677, N604, N587);
not NOT1 (N712, N710);
and AND3 (N713, N712, N601, N121);
nor NOR4 (N714, N711, N176, N490, N418);
nor NOR3 (N715, N709, N238, N196);
or OR2 (N716, N700, N145);
and AND3 (N717, N703, N294, N506);
nand NAND2 (N718, N714, N208);
xor XOR2 (N719, N716, N523);
nand NAND2 (N720, N705, N604);
nor NOR4 (N721, N713, N717, N369, N472);
or OR4 (N722, N135, N382, N452, N114);
nor NOR3 (N723, N715, N251, N647);
and AND2 (N724, N701, N459);
buf BUF1 (N725, N720);
buf BUF1 (N726, N690);
and AND3 (N727, N719, N78, N571);
or OR3 (N728, N722, N280, N489);
or OR4 (N729, N718, N641, N83, N530);
not NOT1 (N730, N721);
and AND4 (N731, N727, N58, N294, N195);
or OR2 (N732, N725, N449);
nor NOR4 (N733, N730, N441, N556, N376);
buf BUF1 (N734, N733);
or OR3 (N735, N732, N7, N149);
or OR2 (N736, N675, N547);
and AND2 (N737, N734, N112);
not NOT1 (N738, N728);
nor NOR4 (N739, N726, N324, N220, N31);
nor NOR2 (N740, N707, N149);
or OR2 (N741, N738, N90);
not NOT1 (N742, N731);
buf BUF1 (N743, N741);
buf BUF1 (N744, N729);
xor XOR2 (N745, N743, N735);
xor XOR2 (N746, N285, N54);
buf BUF1 (N747, N736);
or OR4 (N748, N746, N490, N54, N614);
xor XOR2 (N749, N745, N62);
or OR2 (N750, N748, N515);
not NOT1 (N751, N742);
nor NOR3 (N752, N747, N53, N279);
nand NAND3 (N753, N724, N524, N433);
not NOT1 (N754, N739);
buf BUF1 (N755, N751);
or OR3 (N756, N753, N329, N281);
and AND4 (N757, N744, N691, N141, N225);
buf BUF1 (N758, N723);
nor NOR4 (N759, N755, N596, N748, N376);
buf BUF1 (N760, N758);
buf BUF1 (N761, N759);
not NOT1 (N762, N737);
xor XOR2 (N763, N762, N219);
nand NAND2 (N764, N757, N384);
or OR3 (N765, N756, N646, N320);
and AND4 (N766, N749, N519, N672, N302);
xor XOR2 (N767, N760, N499);
not NOT1 (N768, N761);
nand NAND4 (N769, N763, N249, N508, N146);
or OR4 (N770, N766, N364, N302, N581);
buf BUF1 (N771, N740);
or OR3 (N772, N769, N35, N448);
nand NAND3 (N773, N754, N346, N597);
nand NAND2 (N774, N773, N229);
and AND4 (N775, N765, N279, N398, N663);
or OR2 (N776, N750, N53);
xor XOR2 (N777, N768, N711);
xor XOR2 (N778, N764, N692);
not NOT1 (N779, N775);
buf BUF1 (N780, N778);
xor XOR2 (N781, N770, N206);
or OR3 (N782, N777, N336, N26);
or OR3 (N783, N774, N425, N584);
and AND2 (N784, N772, N24);
not NOT1 (N785, N779);
and AND4 (N786, N782, N459, N592, N325);
buf BUF1 (N787, N776);
nor NOR4 (N788, N784, N353, N155, N583);
nand NAND3 (N789, N771, N221, N570);
buf BUF1 (N790, N767);
buf BUF1 (N791, N786);
xor XOR2 (N792, N791, N705);
nor NOR4 (N793, N781, N327, N544, N485);
buf BUF1 (N794, N780);
not NOT1 (N795, N792);
and AND4 (N796, N788, N563, N73, N157);
and AND4 (N797, N794, N360, N84, N571);
xor XOR2 (N798, N796, N278);
nor NOR2 (N799, N789, N247);
nor NOR4 (N800, N798, N645, N718, N796);
nand NAND2 (N801, N795, N588);
and AND2 (N802, N793, N257);
buf BUF1 (N803, N790);
buf BUF1 (N804, N797);
or OR2 (N805, N800, N672);
not NOT1 (N806, N803);
not NOT1 (N807, N752);
and AND2 (N808, N785, N186);
nor NOR4 (N809, N807, N258, N523, N233);
nand NAND4 (N810, N802, N92, N625, N420);
and AND3 (N811, N805, N789, N157);
nand NAND4 (N812, N787, N54, N192, N691);
not NOT1 (N813, N799);
buf BUF1 (N814, N808);
nor NOR4 (N815, N814, N766, N685, N795);
nor NOR3 (N816, N804, N726, N230);
nand NAND4 (N817, N809, N167, N480, N82);
nor NOR2 (N818, N815, N502);
buf BUF1 (N819, N801);
buf BUF1 (N820, N783);
buf BUF1 (N821, N818);
nand NAND3 (N822, N812, N601, N744);
and AND2 (N823, N813, N732);
buf BUF1 (N824, N806);
buf BUF1 (N825, N823);
nand NAND2 (N826, N821, N54);
nand NAND2 (N827, N811, N820);
buf BUF1 (N828, N672);
nand NAND4 (N829, N824, N313, N10, N605);
xor XOR2 (N830, N825, N811);
buf BUF1 (N831, N816);
not NOT1 (N832, N831);
xor XOR2 (N833, N827, N129);
buf BUF1 (N834, N830);
nor NOR4 (N835, N832, N514, N70, N182);
not NOT1 (N836, N835);
nand NAND3 (N837, N826, N383, N57);
not NOT1 (N838, N817);
or OR3 (N839, N828, N443, N297);
or OR2 (N840, N839, N251);
buf BUF1 (N841, N829);
not NOT1 (N842, N838);
and AND4 (N843, N822, N749, N627, N627);
nand NAND3 (N844, N840, N772, N518);
xor XOR2 (N845, N834, N732);
or OR2 (N846, N842, N464);
buf BUF1 (N847, N810);
or OR2 (N848, N845, N662);
xor XOR2 (N849, N819, N240);
not NOT1 (N850, N849);
and AND2 (N851, N837, N309);
buf BUF1 (N852, N846);
xor XOR2 (N853, N843, N410);
not NOT1 (N854, N850);
xor XOR2 (N855, N854, N628);
and AND3 (N856, N852, N343, N245);
not NOT1 (N857, N848);
nor NOR3 (N858, N836, N6, N13);
or OR2 (N859, N858, N641);
buf BUF1 (N860, N856);
xor XOR2 (N861, N855, N765);
and AND3 (N862, N857, N615, N465);
nor NOR3 (N863, N860, N307, N793);
and AND3 (N864, N861, N850, N432);
not NOT1 (N865, N853);
buf BUF1 (N866, N865);
buf BUF1 (N867, N859);
nor NOR2 (N868, N866, N338);
not NOT1 (N869, N862);
xor XOR2 (N870, N864, N863);
nand NAND3 (N871, N507, N165, N387);
and AND4 (N872, N851, N393, N588, N814);
xor XOR2 (N873, N871, N222);
not NOT1 (N874, N872);
not NOT1 (N875, N868);
not NOT1 (N876, N873);
and AND3 (N877, N847, N422, N721);
nor NOR3 (N878, N874, N798, N99);
and AND4 (N879, N841, N349, N230, N469);
nor NOR3 (N880, N879, N513, N757);
xor XOR2 (N881, N869, N550);
nand NAND4 (N882, N880, N72, N717, N454);
and AND4 (N883, N876, N739, N193, N43);
not NOT1 (N884, N882);
nand NAND3 (N885, N867, N392, N111);
xor XOR2 (N886, N881, N164);
nor NOR2 (N887, N833, N464);
xor XOR2 (N888, N885, N878);
nor NOR4 (N889, N191, N847, N613, N25);
buf BUF1 (N890, N884);
nor NOR2 (N891, N870, N601);
and AND4 (N892, N887, N185, N666, N712);
xor XOR2 (N893, N883, N335);
not NOT1 (N894, N888);
and AND2 (N895, N892, N275);
nand NAND3 (N896, N893, N282, N274);
xor XOR2 (N897, N877, N746);
xor XOR2 (N898, N894, N67);
xor XOR2 (N899, N890, N432);
xor XOR2 (N900, N886, N455);
and AND2 (N901, N898, N115);
or OR3 (N902, N897, N28, N239);
not NOT1 (N903, N891);
not NOT1 (N904, N896);
not NOT1 (N905, N901);
xor XOR2 (N906, N904, N786);
or OR2 (N907, N875, N525);
nand NAND2 (N908, N844, N211);
or OR4 (N909, N899, N42, N702, N653);
nor NOR4 (N910, N906, N853, N488, N29);
nand NAND2 (N911, N902, N525);
xor XOR2 (N912, N911, N873);
buf BUF1 (N913, N903);
nand NAND2 (N914, N889, N821);
and AND4 (N915, N895, N721, N33, N828);
xor XOR2 (N916, N907, N785);
not NOT1 (N917, N916);
nand NAND2 (N918, N910, N880);
and AND2 (N919, N915, N642);
buf BUF1 (N920, N919);
xor XOR2 (N921, N914, N164);
not NOT1 (N922, N908);
xor XOR2 (N923, N912, N200);
nor NOR4 (N924, N922, N623, N486, N51);
or OR2 (N925, N921, N275);
xor XOR2 (N926, N918, N34);
not NOT1 (N927, N923);
nand NAND3 (N928, N926, N467, N927);
buf BUF1 (N929, N909);
xor XOR2 (N930, N218, N312);
nand NAND2 (N931, N900, N758);
xor XOR2 (N932, N920, N193);
xor XOR2 (N933, N905, N644);
not NOT1 (N934, N924);
nand NAND4 (N935, N930, N468, N237, N166);
xor XOR2 (N936, N933, N894);
nand NAND3 (N937, N932, N163, N711);
not NOT1 (N938, N925);
nor NOR4 (N939, N929, N904, N882, N425);
buf BUF1 (N940, N931);
buf BUF1 (N941, N936);
not NOT1 (N942, N928);
nor NOR2 (N943, N934, N683);
or OR3 (N944, N917, N487, N224);
not NOT1 (N945, N937);
nor NOR2 (N946, N942, N191);
nand NAND3 (N947, N946, N565, N192);
and AND3 (N948, N940, N235, N400);
xor XOR2 (N949, N935, N372);
xor XOR2 (N950, N939, N302);
nand NAND3 (N951, N949, N195, N528);
nand NAND2 (N952, N948, N282);
and AND2 (N953, N950, N241);
nand NAND4 (N954, N938, N270, N549, N772);
nand NAND2 (N955, N951, N230);
buf BUF1 (N956, N954);
nand NAND3 (N957, N955, N865, N502);
or OR2 (N958, N913, N429);
nor NOR2 (N959, N945, N620);
buf BUF1 (N960, N941);
nand NAND4 (N961, N947, N576, N726, N313);
not NOT1 (N962, N960);
or OR4 (N963, N956, N236, N300, N536);
not NOT1 (N964, N958);
buf BUF1 (N965, N952);
nor NOR3 (N966, N944, N482, N695);
or OR3 (N967, N964, N923, N124);
xor XOR2 (N968, N966, N409);
not NOT1 (N969, N961);
not NOT1 (N970, N953);
or OR2 (N971, N943, N157);
xor XOR2 (N972, N963, N382);
nand NAND3 (N973, N972, N386, N628);
xor XOR2 (N974, N965, N318);
nor NOR4 (N975, N974, N939, N773, N50);
xor XOR2 (N976, N968, N611);
nor NOR3 (N977, N957, N42, N840);
or OR3 (N978, N967, N976, N731);
nor NOR3 (N979, N877, N698, N396);
buf BUF1 (N980, N969);
and AND4 (N981, N973, N127, N621, N638);
or OR4 (N982, N979, N165, N96, N548);
nor NOR4 (N983, N971, N142, N966, N50);
and AND3 (N984, N959, N469, N741);
or OR2 (N985, N980, N805);
buf BUF1 (N986, N962);
nor NOR4 (N987, N977, N97, N922, N451);
or OR2 (N988, N983, N715);
buf BUF1 (N989, N987);
buf BUF1 (N990, N986);
buf BUF1 (N991, N981);
not NOT1 (N992, N975);
not NOT1 (N993, N982);
nand NAND2 (N994, N991, N631);
buf BUF1 (N995, N989);
or OR4 (N996, N993, N382, N355, N101);
and AND3 (N997, N996, N326, N588);
nand NAND2 (N998, N990, N886);
or OR4 (N999, N992, N658, N865, N833);
xor XOR2 (N1000, N998, N281);
buf BUF1 (N1001, N985);
nor NOR3 (N1002, N1001, N459, N620);
nor NOR2 (N1003, N978, N338);
or OR2 (N1004, N997, N111);
buf BUF1 (N1005, N1004);
buf BUF1 (N1006, N999);
nor NOR4 (N1007, N984, N637, N14, N163);
and AND2 (N1008, N1005, N920);
nand NAND2 (N1009, N1003, N395);
nor NOR4 (N1010, N970, N234, N584, N45);
not NOT1 (N1011, N1006);
nand NAND3 (N1012, N1011, N41, N753);
buf BUF1 (N1013, N1008);
nand NAND3 (N1014, N994, N769, N787);
nand NAND3 (N1015, N1014, N262, N582);
nand NAND3 (N1016, N995, N67, N88);
xor XOR2 (N1017, N988, N967);
xor XOR2 (N1018, N1007, N183);
or OR2 (N1019, N1009, N175);
or OR2 (N1020, N1017, N909);
or OR3 (N1021, N1002, N28, N797);
and AND3 (N1022, N1020, N131, N790);
and AND4 (N1023, N1019, N599, N314, N742);
nand NAND2 (N1024, N1022, N917);
xor XOR2 (N1025, N1015, N766);
not NOT1 (N1026, N1000);
nand NAND4 (N1027, N1013, N1025, N223, N801);
and AND2 (N1028, N215, N316);
nand NAND3 (N1029, N1026, N636, N787);
or OR2 (N1030, N1016, N61);
nor NOR2 (N1031, N1030, N719);
nand NAND2 (N1032, N1028, N780);
nand NAND4 (N1033, N1012, N873, N175, N727);
xor XOR2 (N1034, N1021, N999);
xor XOR2 (N1035, N1034, N265);
not NOT1 (N1036, N1031);
nand NAND4 (N1037, N1032, N1003, N942, N556);
xor XOR2 (N1038, N1027, N3);
buf BUF1 (N1039, N1037);
not NOT1 (N1040, N1024);
nor NOR4 (N1041, N1023, N136, N661, N456);
nand NAND2 (N1042, N1041, N934);
nor NOR3 (N1043, N1029, N100, N842);
or OR2 (N1044, N1039, N79);
and AND4 (N1045, N1035, N948, N139, N508);
not NOT1 (N1046, N1040);
and AND4 (N1047, N1038, N633, N38, N660);
nand NAND2 (N1048, N1047, N1019);
nand NAND4 (N1049, N1033, N414, N679, N939);
and AND3 (N1050, N1043, N238, N613);
nand NAND3 (N1051, N1050, N651, N265);
nand NAND2 (N1052, N1044, N170);
xor XOR2 (N1053, N1018, N901);
or OR3 (N1054, N1045, N924, N514);
buf BUF1 (N1055, N1036);
nor NOR3 (N1056, N1053, N380, N964);
not NOT1 (N1057, N1010);
or OR3 (N1058, N1052, N197, N145);
and AND3 (N1059, N1042, N240, N118);
nand NAND3 (N1060, N1055, N867, N856);
or OR2 (N1061, N1059, N671);
xor XOR2 (N1062, N1049, N682);
nor NOR4 (N1063, N1058, N78, N169, N624);
xor XOR2 (N1064, N1048, N708);
nor NOR3 (N1065, N1054, N819, N688);
not NOT1 (N1066, N1065);
not NOT1 (N1067, N1057);
xor XOR2 (N1068, N1060, N1062);
xor XOR2 (N1069, N667, N675);
buf BUF1 (N1070, N1061);
nand NAND4 (N1071, N1069, N115, N532, N970);
not NOT1 (N1072, N1063);
nor NOR4 (N1073, N1071, N564, N586, N354);
or OR4 (N1074, N1068, N890, N888, N1026);
and AND2 (N1075, N1056, N523);
not NOT1 (N1076, N1075);
xor XOR2 (N1077, N1072, N909);
not NOT1 (N1078, N1070);
nor NOR4 (N1079, N1064, N440, N939, N539);
nand NAND4 (N1080, N1046, N439, N651, N366);
nor NOR3 (N1081, N1078, N59, N318);
buf BUF1 (N1082, N1073);
xor XOR2 (N1083, N1076, N297);
not NOT1 (N1084, N1083);
xor XOR2 (N1085, N1081, N231);
or OR4 (N1086, N1077, N150, N793, N653);
not NOT1 (N1087, N1067);
nand NAND3 (N1088, N1082, N506, N160);
or OR2 (N1089, N1074, N926);
not NOT1 (N1090, N1051);
or OR3 (N1091, N1086, N924, N139);
nand NAND2 (N1092, N1088, N514);
not NOT1 (N1093, N1066);
not NOT1 (N1094, N1092);
xor XOR2 (N1095, N1085, N1077);
nand NAND3 (N1096, N1094, N740, N754);
nor NOR2 (N1097, N1079, N1031);
nand NAND2 (N1098, N1084, N242);
or OR4 (N1099, N1097, N390, N327, N683);
or OR2 (N1100, N1093, N19);
nand NAND3 (N1101, N1095, N744, N980);
and AND2 (N1102, N1087, N394);
not NOT1 (N1103, N1102);
xor XOR2 (N1104, N1098, N597);
buf BUF1 (N1105, N1103);
xor XOR2 (N1106, N1089, N862);
buf BUF1 (N1107, N1090);
nor NOR3 (N1108, N1096, N326, N970);
xor XOR2 (N1109, N1108, N749);
and AND3 (N1110, N1100, N474, N190);
nor NOR3 (N1111, N1101, N190, N75);
nor NOR4 (N1112, N1091, N66, N612, N146);
and AND2 (N1113, N1105, N86);
buf BUF1 (N1114, N1080);
xor XOR2 (N1115, N1114, N133);
or OR2 (N1116, N1113, N701);
nand NAND4 (N1117, N1110, N1013, N512, N220);
nand NAND4 (N1118, N1117, N430, N52, N443);
or OR4 (N1119, N1104, N446, N1115, N258);
or OR2 (N1120, N149, N824);
or OR3 (N1121, N1116, N17, N889);
or OR4 (N1122, N1109, N166, N211, N5);
or OR3 (N1123, N1122, N151, N193);
not NOT1 (N1124, N1120);
nor NOR4 (N1125, N1107, N324, N418, N17);
and AND4 (N1126, N1121, N426, N33, N100);
xor XOR2 (N1127, N1123, N587);
or OR3 (N1128, N1125, N583, N507);
and AND4 (N1129, N1106, N1053, N551, N431);
or OR2 (N1130, N1124, N974);
or OR3 (N1131, N1130, N88, N201);
buf BUF1 (N1132, N1127);
and AND4 (N1133, N1129, N416, N355, N361);
xor XOR2 (N1134, N1132, N948);
not NOT1 (N1135, N1111);
nor NOR4 (N1136, N1126, N917, N468, N303);
not NOT1 (N1137, N1119);
nor NOR3 (N1138, N1136, N586, N1047);
or OR2 (N1139, N1133, N1003);
or OR2 (N1140, N1131, N390);
xor XOR2 (N1141, N1112, N861);
or OR3 (N1142, N1141, N37, N879);
not NOT1 (N1143, N1139);
or OR4 (N1144, N1128, N1001, N1027, N660);
nor NOR4 (N1145, N1140, N901, N982, N816);
and AND3 (N1146, N1145, N840, N922);
nand NAND4 (N1147, N1146, N395, N1111, N399);
xor XOR2 (N1148, N1144, N639);
not NOT1 (N1149, N1118);
nor NOR3 (N1150, N1137, N981, N220);
and AND4 (N1151, N1149, N782, N71, N1102);
xor XOR2 (N1152, N1147, N574);
buf BUF1 (N1153, N1134);
buf BUF1 (N1154, N1138);
not NOT1 (N1155, N1148);
nand NAND4 (N1156, N1153, N951, N1110, N919);
nor NOR3 (N1157, N1152, N409, N528);
not NOT1 (N1158, N1157);
and AND2 (N1159, N1142, N506);
and AND4 (N1160, N1150, N332, N534, N981);
or OR2 (N1161, N1155, N206);
buf BUF1 (N1162, N1158);
xor XOR2 (N1163, N1160, N1023);
nand NAND3 (N1164, N1143, N804, N173);
or OR2 (N1165, N1151, N666);
buf BUF1 (N1166, N1162);
and AND4 (N1167, N1154, N514, N548, N921);
xor XOR2 (N1168, N1165, N681);
nand NAND4 (N1169, N1166, N643, N256, N440);
buf BUF1 (N1170, N1135);
xor XOR2 (N1171, N1167, N228);
nand NAND3 (N1172, N1099, N429, N256);
not NOT1 (N1173, N1172);
xor XOR2 (N1174, N1173, N310);
xor XOR2 (N1175, N1159, N947);
not NOT1 (N1176, N1171);
nand NAND2 (N1177, N1168, N1051);
or OR3 (N1178, N1156, N557, N1159);
nand NAND2 (N1179, N1169, N434);
or OR2 (N1180, N1178, N306);
nor NOR3 (N1181, N1177, N388, N376);
and AND2 (N1182, N1176, N132);
nor NOR4 (N1183, N1161, N175, N591, N1089);
nand NAND3 (N1184, N1180, N164, N41);
xor XOR2 (N1185, N1163, N332);
nand NAND2 (N1186, N1164, N233);
not NOT1 (N1187, N1179);
or OR2 (N1188, N1170, N1067);
and AND3 (N1189, N1185, N548, N820);
nor NOR3 (N1190, N1187, N862, N91);
nor NOR2 (N1191, N1175, N663);
nand NAND2 (N1192, N1183, N532);
buf BUF1 (N1193, N1188);
buf BUF1 (N1194, N1184);
or OR2 (N1195, N1190, N374);
and AND4 (N1196, N1194, N867, N1090, N216);
xor XOR2 (N1197, N1193, N273);
not NOT1 (N1198, N1186);
nand NAND3 (N1199, N1191, N467, N62);
or OR2 (N1200, N1199, N69);
nand NAND3 (N1201, N1181, N1126, N1082);
and AND2 (N1202, N1201, N270);
buf BUF1 (N1203, N1195);
xor XOR2 (N1204, N1198, N830);
buf BUF1 (N1205, N1189);
not NOT1 (N1206, N1182);
nand NAND2 (N1207, N1192, N169);
and AND4 (N1208, N1197, N35, N481, N1169);
and AND3 (N1209, N1174, N1118, N691);
buf BUF1 (N1210, N1208);
nand NAND3 (N1211, N1207, N136, N425);
buf BUF1 (N1212, N1210);
xor XOR2 (N1213, N1206, N755);
buf BUF1 (N1214, N1203);
xor XOR2 (N1215, N1205, N745);
not NOT1 (N1216, N1202);
buf BUF1 (N1217, N1204);
xor XOR2 (N1218, N1214, N1147);
and AND4 (N1219, N1211, N978, N754, N456);
nand NAND4 (N1220, N1218, N666, N403, N340);
nor NOR2 (N1221, N1215, N187);
nor NOR4 (N1222, N1216, N1204, N577, N3);
or OR2 (N1223, N1217, N941);
xor XOR2 (N1224, N1213, N838);
buf BUF1 (N1225, N1223);
nand NAND2 (N1226, N1224, N411);
or OR3 (N1227, N1212, N200, N746);
nand NAND3 (N1228, N1225, N949, N56);
and AND4 (N1229, N1227, N1035, N498, N421);
xor XOR2 (N1230, N1221, N446);
nand NAND4 (N1231, N1222, N645, N306, N246);
nand NAND2 (N1232, N1231, N113);
or OR3 (N1233, N1232, N510, N427);
buf BUF1 (N1234, N1220);
nor NOR2 (N1235, N1228, N1045);
and AND3 (N1236, N1234, N551, N1088);
not NOT1 (N1237, N1209);
or OR4 (N1238, N1219, N470, N1013, N328);
buf BUF1 (N1239, N1226);
and AND2 (N1240, N1235, N1031);
nand NAND2 (N1241, N1238, N934);
not NOT1 (N1242, N1230);
or OR3 (N1243, N1196, N515, N1054);
buf BUF1 (N1244, N1229);
xor XOR2 (N1245, N1241, N136);
xor XOR2 (N1246, N1200, N656);
nand NAND2 (N1247, N1233, N772);
and AND2 (N1248, N1246, N919);
or OR2 (N1249, N1243, N481);
nand NAND3 (N1250, N1247, N516, N474);
nand NAND3 (N1251, N1244, N764, N561);
xor XOR2 (N1252, N1236, N849);
buf BUF1 (N1253, N1240);
nand NAND2 (N1254, N1253, N127);
nor NOR2 (N1255, N1237, N194);
xor XOR2 (N1256, N1254, N681);
nand NAND4 (N1257, N1255, N1075, N184, N1191);
and AND3 (N1258, N1249, N751, N944);
buf BUF1 (N1259, N1242);
buf BUF1 (N1260, N1256);
xor XOR2 (N1261, N1250, N293);
nand NAND4 (N1262, N1259, N156, N913, N365);
nor NOR3 (N1263, N1239, N270, N423);
nand NAND3 (N1264, N1260, N164, N58);
and AND2 (N1265, N1257, N824);
or OR2 (N1266, N1248, N1090);
buf BUF1 (N1267, N1245);
xor XOR2 (N1268, N1251, N145);
nor NOR2 (N1269, N1266, N1232);
buf BUF1 (N1270, N1268);
nand NAND2 (N1271, N1267, N159);
not NOT1 (N1272, N1252);
buf BUF1 (N1273, N1272);
nand NAND3 (N1274, N1264, N619, N167);
xor XOR2 (N1275, N1274, N298);
nor NOR2 (N1276, N1273, N987);
not NOT1 (N1277, N1263);
not NOT1 (N1278, N1258);
nand NAND2 (N1279, N1275, N128);
and AND2 (N1280, N1261, N113);
nand NAND3 (N1281, N1280, N359, N1110);
and AND2 (N1282, N1278, N681);
nor NOR3 (N1283, N1282, N1214, N1231);
and AND4 (N1284, N1265, N966, N432, N1225);
and AND3 (N1285, N1262, N57, N95);
xor XOR2 (N1286, N1285, N377);
and AND4 (N1287, N1276, N1059, N952, N1176);
buf BUF1 (N1288, N1269);
or OR2 (N1289, N1284, N1030);
or OR4 (N1290, N1288, N1158, N1192, N56);
xor XOR2 (N1291, N1287, N110);
not NOT1 (N1292, N1277);
nor NOR3 (N1293, N1270, N1121, N345);
nor NOR4 (N1294, N1290, N1007, N339, N771);
or OR4 (N1295, N1294, N997, N1266, N937);
and AND4 (N1296, N1289, N877, N770, N467);
and AND2 (N1297, N1291, N1052);
not NOT1 (N1298, N1279);
or OR2 (N1299, N1297, N1095);
not NOT1 (N1300, N1295);
not NOT1 (N1301, N1292);
nand NAND4 (N1302, N1296, N1121, N143, N24);
xor XOR2 (N1303, N1283, N571);
nand NAND4 (N1304, N1299, N49, N233, N107);
not NOT1 (N1305, N1293);
not NOT1 (N1306, N1300);
buf BUF1 (N1307, N1305);
xor XOR2 (N1308, N1303, N1223);
xor XOR2 (N1309, N1304, N287);
or OR3 (N1310, N1302, N159, N735);
nor NOR4 (N1311, N1307, N297, N897, N258);
nor NOR4 (N1312, N1306, N886, N389, N1058);
nor NOR2 (N1313, N1308, N351);
nand NAND2 (N1314, N1298, N775);
or OR2 (N1315, N1312, N425);
not NOT1 (N1316, N1315);
buf BUF1 (N1317, N1316);
or OR2 (N1318, N1317, N197);
not NOT1 (N1319, N1313);
nand NAND2 (N1320, N1319, N546);
not NOT1 (N1321, N1320);
nor NOR3 (N1322, N1321, N1243, N647);
buf BUF1 (N1323, N1286);
buf BUF1 (N1324, N1310);
nand NAND3 (N1325, N1314, N1088, N917);
nand NAND2 (N1326, N1281, N296);
not NOT1 (N1327, N1318);
buf BUF1 (N1328, N1327);
and AND4 (N1329, N1326, N768, N432, N1311);
nand NAND2 (N1330, N360, N1323);
or OR3 (N1331, N438, N218, N320);
nand NAND4 (N1332, N1329, N869, N1021, N805);
xor XOR2 (N1333, N1271, N1050);
or OR4 (N1334, N1331, N1284, N591, N1190);
xor XOR2 (N1335, N1322, N529);
buf BUF1 (N1336, N1332);
nand NAND4 (N1337, N1334, N373, N454, N293);
nor NOR4 (N1338, N1324, N679, N1296, N767);
xor XOR2 (N1339, N1325, N1142);
buf BUF1 (N1340, N1301);
or OR2 (N1341, N1340, N1227);
nor NOR3 (N1342, N1328, N1023, N1003);
not NOT1 (N1343, N1335);
or OR4 (N1344, N1336, N32, N1125, N485);
nor NOR2 (N1345, N1341, N540);
and AND3 (N1346, N1345, N670, N475);
and AND4 (N1347, N1346, N109, N550, N83);
not NOT1 (N1348, N1339);
not NOT1 (N1349, N1338);
or OR3 (N1350, N1349, N1120, N82);
buf BUF1 (N1351, N1347);
or OR4 (N1352, N1344, N86, N1310, N682);
not NOT1 (N1353, N1348);
nor NOR3 (N1354, N1352, N322, N121);
xor XOR2 (N1355, N1350, N285);
nand NAND3 (N1356, N1333, N127, N752);
and AND4 (N1357, N1355, N567, N582, N242);
or OR3 (N1358, N1354, N1070, N781);
nand NAND2 (N1359, N1337, N585);
or OR2 (N1360, N1353, N1015);
and AND4 (N1361, N1343, N1111, N1113, N463);
nor NOR2 (N1362, N1356, N1173);
nand NAND4 (N1363, N1330, N742, N725, N1007);
nand NAND3 (N1364, N1363, N850, N1323);
not NOT1 (N1365, N1351);
and AND4 (N1366, N1342, N241, N1042, N854);
nand NAND3 (N1367, N1360, N87, N855);
buf BUF1 (N1368, N1366);
not NOT1 (N1369, N1364);
nor NOR4 (N1370, N1361, N927, N902, N675);
nor NOR4 (N1371, N1362, N416, N250, N1151);
not NOT1 (N1372, N1309);
xor XOR2 (N1373, N1367, N1293);
not NOT1 (N1374, N1365);
or OR4 (N1375, N1368, N1126, N474, N118);
not NOT1 (N1376, N1357);
and AND3 (N1377, N1375, N746, N508);
not NOT1 (N1378, N1376);
or OR3 (N1379, N1359, N795, N1333);
buf BUF1 (N1380, N1358);
xor XOR2 (N1381, N1370, N1357);
nor NOR4 (N1382, N1371, N962, N546, N598);
and AND2 (N1383, N1378, N695);
not NOT1 (N1384, N1369);
not NOT1 (N1385, N1380);
buf BUF1 (N1386, N1381);
xor XOR2 (N1387, N1374, N1011);
not NOT1 (N1388, N1387);
or OR3 (N1389, N1388, N683, N292);
or OR3 (N1390, N1382, N487, N889);
nor NOR2 (N1391, N1386, N1028);
nand NAND3 (N1392, N1390, N204, N1219);
or OR2 (N1393, N1385, N524);
buf BUF1 (N1394, N1377);
and AND4 (N1395, N1373, N1372, N1340, N481);
buf BUF1 (N1396, N975);
not NOT1 (N1397, N1383);
buf BUF1 (N1398, N1379);
and AND3 (N1399, N1396, N1319, N114);
not NOT1 (N1400, N1389);
nor NOR2 (N1401, N1397, N1133);
nor NOR3 (N1402, N1400, N281, N55);
buf BUF1 (N1403, N1394);
xor XOR2 (N1404, N1402, N311);
nand NAND2 (N1405, N1398, N676);
nor NOR4 (N1406, N1401, N1113, N1107, N474);
not NOT1 (N1407, N1405);
nor NOR4 (N1408, N1395, N693, N321, N1028);
not NOT1 (N1409, N1391);
buf BUF1 (N1410, N1408);
buf BUF1 (N1411, N1410);
nor NOR3 (N1412, N1392, N607, N521);
buf BUF1 (N1413, N1404);
nor NOR4 (N1414, N1411, N1302, N476, N202);
and AND3 (N1415, N1393, N1069, N210);
nand NAND4 (N1416, N1412, N1100, N160, N986);
not NOT1 (N1417, N1399);
nor NOR2 (N1418, N1384, N311);
or OR3 (N1419, N1417, N464, N122);
not NOT1 (N1420, N1415);
not NOT1 (N1421, N1419);
nor NOR3 (N1422, N1407, N801, N1084);
buf BUF1 (N1423, N1420);
and AND4 (N1424, N1416, N1131, N809, N147);
xor XOR2 (N1425, N1413, N249);
xor XOR2 (N1426, N1425, N494);
not NOT1 (N1427, N1406);
or OR3 (N1428, N1424, N454, N1359);
or OR3 (N1429, N1409, N1262, N151);
buf BUF1 (N1430, N1418);
or OR4 (N1431, N1422, N395, N837, N76);
nand NAND4 (N1432, N1429, N975, N915, N564);
buf BUF1 (N1433, N1421);
nand NAND3 (N1434, N1430, N357, N889);
not NOT1 (N1435, N1431);
or OR4 (N1436, N1414, N1067, N523, N220);
xor XOR2 (N1437, N1423, N818);
nand NAND2 (N1438, N1433, N1277);
and AND2 (N1439, N1434, N424);
xor XOR2 (N1440, N1426, N846);
nor NOR2 (N1441, N1435, N784);
buf BUF1 (N1442, N1427);
xor XOR2 (N1443, N1441, N800);
and AND2 (N1444, N1436, N346);
or OR2 (N1445, N1403, N472);
and AND2 (N1446, N1443, N52);
xor XOR2 (N1447, N1442, N944);
buf BUF1 (N1448, N1437);
not NOT1 (N1449, N1447);
nor NOR2 (N1450, N1449, N1395);
nor NOR2 (N1451, N1444, N1308);
nor NOR4 (N1452, N1450, N459, N110, N56);
or OR2 (N1453, N1445, N998);
nor NOR2 (N1454, N1440, N106);
nor NOR3 (N1455, N1453, N288, N1156);
or OR4 (N1456, N1439, N402, N1397, N590);
not NOT1 (N1457, N1448);
or OR4 (N1458, N1432, N587, N1411, N229);
or OR3 (N1459, N1455, N841, N1442);
not NOT1 (N1460, N1456);
nor NOR3 (N1461, N1460, N792, N973);
and AND4 (N1462, N1458, N373, N1015, N920);
and AND3 (N1463, N1446, N400, N1149);
not NOT1 (N1464, N1438);
buf BUF1 (N1465, N1454);
or OR3 (N1466, N1465, N970, N300);
buf BUF1 (N1467, N1464);
xor XOR2 (N1468, N1467, N770);
xor XOR2 (N1469, N1463, N1419);
or OR4 (N1470, N1451, N1214, N229, N1085);
not NOT1 (N1471, N1461);
nand NAND4 (N1472, N1466, N65, N578, N303);
not NOT1 (N1473, N1428);
and AND3 (N1474, N1459, N1136, N480);
nand NAND2 (N1475, N1452, N313);
xor XOR2 (N1476, N1468, N116);
not NOT1 (N1477, N1462);
not NOT1 (N1478, N1475);
and AND2 (N1479, N1469, N1274);
or OR2 (N1480, N1457, N534);
or OR2 (N1481, N1479, N1414);
or OR3 (N1482, N1472, N2, N441);
and AND4 (N1483, N1474, N336, N790, N1031);
or OR3 (N1484, N1481, N654, N1242);
or OR2 (N1485, N1483, N1470);
nand NAND2 (N1486, N652, N545);
buf BUF1 (N1487, N1482);
nor NOR3 (N1488, N1478, N459, N460);
xor XOR2 (N1489, N1480, N44);
nor NOR3 (N1490, N1484, N18, N783);
nand NAND2 (N1491, N1487, N1415);
and AND3 (N1492, N1488, N1130, N706);
xor XOR2 (N1493, N1486, N1389);
nand NAND4 (N1494, N1492, N1154, N50, N1034);
buf BUF1 (N1495, N1493);
not NOT1 (N1496, N1494);
xor XOR2 (N1497, N1489, N534);
nand NAND4 (N1498, N1497, N503, N1246, N1196);
nand NAND2 (N1499, N1490, N393);
and AND3 (N1500, N1495, N710, N539);
nor NOR3 (N1501, N1498, N928, N588);
nor NOR4 (N1502, N1477, N193, N1330, N963);
buf BUF1 (N1503, N1500);
or OR2 (N1504, N1485, N478);
and AND4 (N1505, N1476, N512, N415, N351);
buf BUF1 (N1506, N1502);
nand NAND3 (N1507, N1503, N782, N1414);
buf BUF1 (N1508, N1505);
and AND2 (N1509, N1507, N885);
not NOT1 (N1510, N1506);
xor XOR2 (N1511, N1491, N631);
xor XOR2 (N1512, N1510, N1431);
buf BUF1 (N1513, N1499);
nor NOR3 (N1514, N1471, N1193, N1248);
nor NOR4 (N1515, N1504, N471, N569, N958);
xor XOR2 (N1516, N1508, N663);
and AND3 (N1517, N1514, N357, N325);
nand NAND4 (N1518, N1496, N209, N722, N759);
nand NAND3 (N1519, N1517, N457, N892);
or OR4 (N1520, N1519, N804, N237, N1300);
and AND4 (N1521, N1512, N758, N1341, N552);
nand NAND3 (N1522, N1515, N734, N1233);
buf BUF1 (N1523, N1509);
xor XOR2 (N1524, N1523, N507);
buf BUF1 (N1525, N1501);
nand NAND4 (N1526, N1518, N986, N581, N150);
xor XOR2 (N1527, N1526, N840);
and AND4 (N1528, N1522, N453, N1059, N1520);
or OR4 (N1529, N1378, N271, N202, N1094);
not NOT1 (N1530, N1525);
buf BUF1 (N1531, N1528);
xor XOR2 (N1532, N1473, N892);
or OR4 (N1533, N1524, N912, N9, N1099);
and AND3 (N1534, N1532, N901, N808);
xor XOR2 (N1535, N1533, N1455);
or OR4 (N1536, N1535, N1252, N1117, N1010);
not NOT1 (N1537, N1511);
nand NAND3 (N1538, N1530, N7, N1382);
nand NAND4 (N1539, N1531, N1422, N483, N1276);
xor XOR2 (N1540, N1537, N101);
not NOT1 (N1541, N1538);
or OR3 (N1542, N1521, N1015, N494);
nor NOR3 (N1543, N1541, N1389, N1502);
or OR3 (N1544, N1539, N892, N748);
not NOT1 (N1545, N1543);
nand NAND2 (N1546, N1544, N182);
nand NAND3 (N1547, N1536, N64, N433);
buf BUF1 (N1548, N1534);
buf BUF1 (N1549, N1546);
or OR4 (N1550, N1545, N1540, N363, N140);
nand NAND2 (N1551, N755, N930);
and AND3 (N1552, N1542, N79, N1490);
xor XOR2 (N1553, N1529, N1083);
or OR3 (N1554, N1551, N62, N95);
or OR2 (N1555, N1552, N1357);
and AND4 (N1556, N1549, N1218, N369, N273);
nor NOR4 (N1557, N1547, N23, N105, N84);
xor XOR2 (N1558, N1554, N1254);
xor XOR2 (N1559, N1527, N1452);
xor XOR2 (N1560, N1513, N56);
or OR4 (N1561, N1550, N1238, N1186, N471);
nand NAND2 (N1562, N1560, N1277);
or OR4 (N1563, N1557, N1336, N1377, N314);
buf BUF1 (N1564, N1558);
or OR2 (N1565, N1564, N662);
and AND4 (N1566, N1548, N1212, N1547, N1565);
or OR2 (N1567, N1060, N134);
xor XOR2 (N1568, N1553, N220);
not NOT1 (N1569, N1559);
or OR2 (N1570, N1561, N142);
nand NAND4 (N1571, N1568, N80, N688, N1363);
or OR4 (N1572, N1569, N318, N856, N198);
nor NOR4 (N1573, N1566, N403, N1380, N554);
and AND3 (N1574, N1562, N1521, N946);
nor NOR4 (N1575, N1572, N555, N866, N316);
not NOT1 (N1576, N1573);
nor NOR2 (N1577, N1575, N690);
or OR2 (N1578, N1576, N1496);
xor XOR2 (N1579, N1567, N267);
or OR3 (N1580, N1574, N1552, N41);
not NOT1 (N1581, N1555);
xor XOR2 (N1582, N1580, N1324);
buf BUF1 (N1583, N1571);
and AND2 (N1584, N1563, N465);
or OR4 (N1585, N1579, N671, N277, N1224);
nand NAND2 (N1586, N1583, N653);
not NOT1 (N1587, N1586);
buf BUF1 (N1588, N1587);
buf BUF1 (N1589, N1584);
xor XOR2 (N1590, N1570, N933);
not NOT1 (N1591, N1590);
buf BUF1 (N1592, N1588);
or OR2 (N1593, N1582, N701);
not NOT1 (N1594, N1577);
not NOT1 (N1595, N1591);
buf BUF1 (N1596, N1594);
nand NAND3 (N1597, N1593, N531, N1030);
nor NOR4 (N1598, N1516, N458, N67, N1327);
not NOT1 (N1599, N1597);
or OR3 (N1600, N1596, N270, N580);
nor NOR3 (N1601, N1556, N103, N435);
not NOT1 (N1602, N1578);
xor XOR2 (N1603, N1600, N1501);
nor NOR2 (N1604, N1599, N1574);
xor XOR2 (N1605, N1592, N1002);
not NOT1 (N1606, N1602);
and AND4 (N1607, N1603, N1447, N432, N161);
not NOT1 (N1608, N1598);
xor XOR2 (N1609, N1581, N453);
and AND2 (N1610, N1607, N1301);
xor XOR2 (N1611, N1608, N690);
xor XOR2 (N1612, N1606, N168);
xor XOR2 (N1613, N1589, N664);
xor XOR2 (N1614, N1595, N137);
and AND4 (N1615, N1614, N865, N1190, N1146);
and AND2 (N1616, N1605, N754);
nand NAND3 (N1617, N1609, N1492, N1309);
or OR3 (N1618, N1604, N1089, N1371);
xor XOR2 (N1619, N1618, N256);
buf BUF1 (N1620, N1613);
and AND3 (N1621, N1601, N629, N1069);
and AND3 (N1622, N1611, N809, N1131);
and AND4 (N1623, N1621, N1012, N794, N1503);
buf BUF1 (N1624, N1615);
and AND4 (N1625, N1622, N944, N1386, N779);
not NOT1 (N1626, N1610);
buf BUF1 (N1627, N1616);
or OR4 (N1628, N1617, N369, N496, N803);
buf BUF1 (N1629, N1624);
and AND3 (N1630, N1585, N59, N826);
nand NAND2 (N1631, N1626, N652);
and AND3 (N1632, N1625, N116, N360);
nor NOR4 (N1633, N1630, N23, N94, N420);
or OR2 (N1634, N1629, N442);
not NOT1 (N1635, N1623);
or OR3 (N1636, N1634, N555, N1627);
xor XOR2 (N1637, N501, N264);
and AND3 (N1638, N1628, N832, N625);
or OR3 (N1639, N1636, N969, N934);
nor NOR3 (N1640, N1635, N1391, N119);
buf BUF1 (N1641, N1638);
not NOT1 (N1642, N1637);
nand NAND2 (N1643, N1640, N1596);
or OR4 (N1644, N1633, N1093, N368, N494);
nor NOR3 (N1645, N1620, N537, N814);
not NOT1 (N1646, N1641);
nand NAND3 (N1647, N1643, N1251, N1441);
or OR2 (N1648, N1647, N39);
or OR3 (N1649, N1646, N1266, N912);
or OR3 (N1650, N1639, N1213, N1174);
nor NOR2 (N1651, N1644, N1049);
xor XOR2 (N1652, N1651, N1517);
nand NAND3 (N1653, N1649, N975, N754);
or OR4 (N1654, N1645, N1605, N1635, N373);
nand NAND4 (N1655, N1642, N1235, N1510, N1519);
nor NOR4 (N1656, N1631, N1572, N1329, N309);
nand NAND4 (N1657, N1654, N825, N959, N1294);
nor NOR2 (N1658, N1652, N673);
or OR2 (N1659, N1632, N1341);
not NOT1 (N1660, N1653);
xor XOR2 (N1661, N1612, N440);
not NOT1 (N1662, N1650);
and AND4 (N1663, N1662, N1066, N1074, N1247);
nor NOR4 (N1664, N1648, N481, N1610, N313);
xor XOR2 (N1665, N1619, N64);
nand NAND4 (N1666, N1655, N1283, N1628, N1519);
and AND3 (N1667, N1657, N980, N1377);
xor XOR2 (N1668, N1666, N1446);
nand NAND2 (N1669, N1668, N785);
buf BUF1 (N1670, N1659);
and AND2 (N1671, N1656, N1300);
not NOT1 (N1672, N1663);
buf BUF1 (N1673, N1670);
xor XOR2 (N1674, N1664, N1131);
xor XOR2 (N1675, N1669, N257);
nor NOR4 (N1676, N1665, N1620, N209, N1116);
not NOT1 (N1677, N1671);
buf BUF1 (N1678, N1676);
nor NOR4 (N1679, N1672, N1600, N93, N458);
not NOT1 (N1680, N1661);
xor XOR2 (N1681, N1679, N402);
xor XOR2 (N1682, N1673, N730);
or OR2 (N1683, N1681, N357);
nor NOR3 (N1684, N1658, N1170, N110);
buf BUF1 (N1685, N1660);
buf BUF1 (N1686, N1677);
and AND3 (N1687, N1683, N788, N1377);
and AND3 (N1688, N1678, N1141, N1058);
and AND4 (N1689, N1675, N1620, N1465, N797);
or OR4 (N1690, N1687, N1109, N986, N485);
nand NAND2 (N1691, N1688, N68);
nand NAND4 (N1692, N1684, N439, N334, N62);
and AND4 (N1693, N1690, N18, N1170, N832);
buf BUF1 (N1694, N1667);
nor NOR3 (N1695, N1674, N915, N243);
nand NAND3 (N1696, N1692, N562, N345);
not NOT1 (N1697, N1682);
nand NAND3 (N1698, N1696, N294, N292);
nor NOR3 (N1699, N1689, N844, N1145);
not NOT1 (N1700, N1694);
nor NOR3 (N1701, N1691, N659, N222);
or OR3 (N1702, N1680, N772, N1633);
xor XOR2 (N1703, N1698, N1258);
nand NAND2 (N1704, N1693, N325);
or OR2 (N1705, N1702, N392);
buf BUF1 (N1706, N1686);
buf BUF1 (N1707, N1699);
buf BUF1 (N1708, N1706);
and AND2 (N1709, N1700, N1488);
xor XOR2 (N1710, N1708, N253);
xor XOR2 (N1711, N1703, N1586);
buf BUF1 (N1712, N1711);
or OR3 (N1713, N1707, N288, N553);
or OR2 (N1714, N1685, N552);
xor XOR2 (N1715, N1713, N1345);
nand NAND4 (N1716, N1710, N1594, N1463, N350);
and AND2 (N1717, N1715, N1394);
buf BUF1 (N1718, N1717);
xor XOR2 (N1719, N1714, N325);
nand NAND4 (N1720, N1716, N899, N1440, N975);
nand NAND3 (N1721, N1712, N1191, N404);
nor NOR2 (N1722, N1709, N542);
nor NOR4 (N1723, N1722, N58, N1274, N426);
and AND2 (N1724, N1701, N429);
not NOT1 (N1725, N1704);
xor XOR2 (N1726, N1697, N1179);
buf BUF1 (N1727, N1719);
nand NAND3 (N1728, N1725, N938, N408);
nand NAND3 (N1729, N1705, N840, N1676);
buf BUF1 (N1730, N1728);
or OR2 (N1731, N1720, N1248);
nand NAND3 (N1732, N1723, N1676, N1077);
nand NAND3 (N1733, N1727, N1381, N762);
xor XOR2 (N1734, N1730, N741);
or OR3 (N1735, N1721, N1072, N77);
nand NAND3 (N1736, N1695, N1328, N851);
or OR2 (N1737, N1735, N193);
nor NOR3 (N1738, N1726, N460, N623);
or OR4 (N1739, N1724, N758, N1263, N47);
not NOT1 (N1740, N1738);
nand NAND3 (N1741, N1729, N539, N1537);
not NOT1 (N1742, N1734);
nor NOR3 (N1743, N1732, N1446, N1025);
buf BUF1 (N1744, N1733);
buf BUF1 (N1745, N1731);
or OR3 (N1746, N1740, N78, N1354);
nand NAND4 (N1747, N1741, N1112, N210, N1604);
nor NOR3 (N1748, N1747, N542, N728);
nand NAND2 (N1749, N1748, N206);
and AND3 (N1750, N1718, N701, N786);
not NOT1 (N1751, N1739);
xor XOR2 (N1752, N1751, N793);
nor NOR4 (N1753, N1742, N779, N314, N40);
not NOT1 (N1754, N1744);
buf BUF1 (N1755, N1749);
nor NOR4 (N1756, N1753, N1397, N1565, N696);
buf BUF1 (N1757, N1743);
buf BUF1 (N1758, N1745);
xor XOR2 (N1759, N1756, N1314);
not NOT1 (N1760, N1754);
nand NAND2 (N1761, N1760, N1160);
or OR2 (N1762, N1755, N320);
buf BUF1 (N1763, N1759);
nand NAND3 (N1764, N1752, N1115, N985);
and AND3 (N1765, N1758, N202, N556);
or OR2 (N1766, N1765, N1576);
nand NAND3 (N1767, N1746, N319, N20);
xor XOR2 (N1768, N1767, N11);
buf BUF1 (N1769, N1764);
nand NAND3 (N1770, N1761, N103, N250);
xor XOR2 (N1771, N1770, N393);
nand NAND2 (N1772, N1737, N1367);
nand NAND4 (N1773, N1736, N851, N349, N178);
buf BUF1 (N1774, N1750);
not NOT1 (N1775, N1774);
buf BUF1 (N1776, N1763);
nand NAND4 (N1777, N1775, N278, N1435, N654);
nor NOR4 (N1778, N1772, N1218, N619, N369);
not NOT1 (N1779, N1762);
or OR4 (N1780, N1768, N1133, N742, N1584);
xor XOR2 (N1781, N1776, N489);
not NOT1 (N1782, N1757);
and AND3 (N1783, N1769, N1087, N203);
not NOT1 (N1784, N1778);
nor NOR4 (N1785, N1773, N46, N493, N782);
not NOT1 (N1786, N1777);
not NOT1 (N1787, N1786);
or OR3 (N1788, N1783, N962, N1218);
or OR3 (N1789, N1771, N600, N1372);
nor NOR4 (N1790, N1788, N240, N1223, N273);
not NOT1 (N1791, N1789);
not NOT1 (N1792, N1779);
buf BUF1 (N1793, N1787);
not NOT1 (N1794, N1766);
nand NAND3 (N1795, N1785, N744, N102);
nand NAND2 (N1796, N1790, N1058);
nand NAND4 (N1797, N1784, N926, N1697, N778);
and AND4 (N1798, N1780, N191, N1248, N550);
or OR4 (N1799, N1795, N299, N1481, N973);
xor XOR2 (N1800, N1797, N1324);
xor XOR2 (N1801, N1791, N1712);
buf BUF1 (N1802, N1796);
nor NOR4 (N1803, N1793, N354, N532, N59);
and AND2 (N1804, N1782, N1309);
not NOT1 (N1805, N1799);
nand NAND2 (N1806, N1781, N1007);
not NOT1 (N1807, N1803);
nand NAND3 (N1808, N1805, N673, N1500);
and AND2 (N1809, N1794, N991);
and AND2 (N1810, N1792, N1575);
buf BUF1 (N1811, N1801);
buf BUF1 (N1812, N1811);
buf BUF1 (N1813, N1800);
xor XOR2 (N1814, N1806, N1309);
buf BUF1 (N1815, N1804);
not NOT1 (N1816, N1807);
or OR3 (N1817, N1813, N1496, N1037);
or OR2 (N1818, N1808, N1394);
xor XOR2 (N1819, N1812, N1479);
nor NOR4 (N1820, N1818, N762, N1789, N1337);
and AND4 (N1821, N1817, N1087, N576, N1234);
nand NAND4 (N1822, N1819, N1111, N1412, N666);
not NOT1 (N1823, N1802);
not NOT1 (N1824, N1815);
buf BUF1 (N1825, N1810);
and AND3 (N1826, N1814, N582, N331);
nor NOR4 (N1827, N1822, N959, N1265, N1551);
nand NAND2 (N1828, N1827, N732);
not NOT1 (N1829, N1820);
nand NAND3 (N1830, N1825, N1503, N1440);
or OR2 (N1831, N1826, N1815);
nor NOR3 (N1832, N1831, N217, N679);
buf BUF1 (N1833, N1823);
nor NOR2 (N1834, N1830, N903);
not NOT1 (N1835, N1829);
not NOT1 (N1836, N1832);
nor NOR2 (N1837, N1833, N540);
nand NAND2 (N1838, N1828, N255);
nor NOR3 (N1839, N1836, N480, N1586);
nor NOR3 (N1840, N1809, N718, N1379);
buf BUF1 (N1841, N1840);
nand NAND2 (N1842, N1816, N755);
not NOT1 (N1843, N1837);
not NOT1 (N1844, N1824);
and AND4 (N1845, N1844, N1778, N1293, N787);
nor NOR4 (N1846, N1834, N875, N243, N952);
and AND3 (N1847, N1841, N1250, N558);
xor XOR2 (N1848, N1821, N422);
xor XOR2 (N1849, N1843, N617);
and AND4 (N1850, N1835, N1628, N1639, N1052);
and AND2 (N1851, N1850, N692);
or OR4 (N1852, N1842, N1, N1814, N1447);
nor NOR2 (N1853, N1798, N816);
nand NAND4 (N1854, N1852, N360, N1780, N1140);
nor NOR4 (N1855, N1849, N1116, N1600, N990);
xor XOR2 (N1856, N1853, N1609);
not NOT1 (N1857, N1845);
buf BUF1 (N1858, N1855);
or OR4 (N1859, N1858, N570, N50, N1457);
not NOT1 (N1860, N1857);
nor NOR3 (N1861, N1851, N408, N380);
xor XOR2 (N1862, N1856, N1554);
not NOT1 (N1863, N1859);
nor NOR2 (N1864, N1861, N1501);
buf BUF1 (N1865, N1848);
or OR4 (N1866, N1860, N1571, N1049, N675);
or OR3 (N1867, N1839, N605, N1456);
nand NAND2 (N1868, N1865, N1066);
or OR4 (N1869, N1866, N1048, N25, N148);
xor XOR2 (N1870, N1846, N1378);
nor NOR4 (N1871, N1838, N665, N1574, N618);
xor XOR2 (N1872, N1867, N350);
not NOT1 (N1873, N1863);
nor NOR4 (N1874, N1868, N1101, N816, N271);
nand NAND4 (N1875, N1871, N743, N78, N1396);
xor XOR2 (N1876, N1870, N777);
nand NAND3 (N1877, N1862, N1648, N1482);
buf BUF1 (N1878, N1869);
not NOT1 (N1879, N1864);
nor NOR3 (N1880, N1847, N1853, N1483);
buf BUF1 (N1881, N1874);
nor NOR4 (N1882, N1872, N454, N547, N1461);
buf BUF1 (N1883, N1881);
xor XOR2 (N1884, N1877, N889);
nor NOR4 (N1885, N1884, N1574, N1747, N15);
or OR4 (N1886, N1879, N253, N36, N104);
nand NAND4 (N1887, N1883, N97, N998, N1750);
nor NOR3 (N1888, N1882, N511, N1334);
xor XOR2 (N1889, N1885, N1153);
and AND2 (N1890, N1873, N1238);
not NOT1 (N1891, N1887);
nand NAND4 (N1892, N1880, N1365, N1587, N1247);
nor NOR4 (N1893, N1892, N1376, N425, N1859);
not NOT1 (N1894, N1878);
buf BUF1 (N1895, N1894);
nor NOR3 (N1896, N1876, N107, N1389);
and AND3 (N1897, N1888, N601, N1769);
not NOT1 (N1898, N1893);
xor XOR2 (N1899, N1897, N1369);
and AND2 (N1900, N1854, N1413);
or OR4 (N1901, N1886, N594, N1352, N670);
not NOT1 (N1902, N1900);
xor XOR2 (N1903, N1895, N550);
nor NOR3 (N1904, N1896, N1701, N1177);
not NOT1 (N1905, N1891);
buf BUF1 (N1906, N1904);
xor XOR2 (N1907, N1898, N875);
xor XOR2 (N1908, N1899, N335);
and AND3 (N1909, N1875, N1255, N411);
or OR4 (N1910, N1907, N1619, N1800, N1759);
nor NOR3 (N1911, N1902, N559, N1850);
or OR2 (N1912, N1901, N1857);
nand NAND2 (N1913, N1905, N231);
nor NOR2 (N1914, N1911, N611);
xor XOR2 (N1915, N1909, N1151);
not NOT1 (N1916, N1889);
buf BUF1 (N1917, N1908);
buf BUF1 (N1918, N1906);
buf BUF1 (N1919, N1903);
buf BUF1 (N1920, N1918);
buf BUF1 (N1921, N1917);
and AND3 (N1922, N1890, N696, N1699);
nand NAND4 (N1923, N1916, N685, N1072, N1567);
not NOT1 (N1924, N1910);
nor NOR2 (N1925, N1924, N168);
or OR2 (N1926, N1912, N1793);
xor XOR2 (N1927, N1919, N1751);
or OR2 (N1928, N1922, N171);
and AND3 (N1929, N1914, N1540, N1166);
or OR4 (N1930, N1925, N48, N1823, N626);
buf BUF1 (N1931, N1928);
buf BUF1 (N1932, N1930);
xor XOR2 (N1933, N1927, N407);
not NOT1 (N1934, N1933);
and AND3 (N1935, N1923, N236, N624);
not NOT1 (N1936, N1915);
nor NOR3 (N1937, N1936, N440, N1297);
nand NAND2 (N1938, N1932, N817);
buf BUF1 (N1939, N1921);
xor XOR2 (N1940, N1937, N1600);
xor XOR2 (N1941, N1935, N310);
buf BUF1 (N1942, N1938);
not NOT1 (N1943, N1929);
nand NAND3 (N1944, N1931, N965, N103);
not NOT1 (N1945, N1943);
buf BUF1 (N1946, N1944);
xor XOR2 (N1947, N1941, N1416);
not NOT1 (N1948, N1934);
buf BUF1 (N1949, N1948);
or OR3 (N1950, N1939, N1145, N900);
or OR4 (N1951, N1940, N525, N1221, N1575);
nor NOR2 (N1952, N1949, N375);
nor NOR3 (N1953, N1950, N536, N1321);
and AND2 (N1954, N1913, N671);
or OR3 (N1955, N1920, N1931, N877);
and AND4 (N1956, N1946, N36, N117, N1001);
and AND4 (N1957, N1954, N441, N1214, N47);
nand NAND3 (N1958, N1926, N379, N79);
nand NAND4 (N1959, N1942, N529, N91, N1655);
or OR4 (N1960, N1955, N1326, N137, N1009);
or OR3 (N1961, N1956, N1660, N866);
nor NOR3 (N1962, N1952, N814, N933);
not NOT1 (N1963, N1953);
nor NOR4 (N1964, N1945, N1249, N479, N1522);
or OR3 (N1965, N1957, N510, N245);
not NOT1 (N1966, N1960);
or OR2 (N1967, N1966, N1889);
nand NAND3 (N1968, N1951, N1678, N1578);
and AND2 (N1969, N1964, N998);
nand NAND4 (N1970, N1963, N1617, N1240, N737);
nand NAND3 (N1971, N1969, N1355, N850);
and AND3 (N1972, N1970, N1054, N775);
buf BUF1 (N1973, N1971);
xor XOR2 (N1974, N1968, N316);
xor XOR2 (N1975, N1965, N1559);
nor NOR3 (N1976, N1973, N503, N1484);
not NOT1 (N1977, N1975);
or OR4 (N1978, N1967, N155, N474, N1007);
nand NAND2 (N1979, N1977, N565);
nand NAND2 (N1980, N1978, N1636);
not NOT1 (N1981, N1961);
buf BUF1 (N1982, N1980);
and AND4 (N1983, N1972, N299, N1612, N1146);
or OR2 (N1984, N1982, N831);
or OR4 (N1985, N1962, N383, N7, N1066);
nor NOR2 (N1986, N1979, N1640);
buf BUF1 (N1987, N1986);
xor XOR2 (N1988, N1987, N1390);
nor NOR4 (N1989, N1988, N948, N1553, N143);
and AND4 (N1990, N1989, N1638, N599, N479);
buf BUF1 (N1991, N1976);
or OR4 (N1992, N1990, N1020, N1339, N1823);
nor NOR2 (N1993, N1991, N1753);
buf BUF1 (N1994, N1947);
and AND4 (N1995, N1981, N338, N1241, N335);
or OR4 (N1996, N1983, N29, N1301, N1613);
not NOT1 (N1997, N1985);
or OR4 (N1998, N1958, N415, N321, N1127);
nor NOR2 (N1999, N1998, N1870);
and AND3 (N2000, N1974, N1692, N1724);
buf BUF1 (N2001, N1995);
or OR2 (N2002, N2001, N1966);
not NOT1 (N2003, N2002);
or OR3 (N2004, N1993, N797, N1887);
nand NAND2 (N2005, N1994, N1287);
nor NOR3 (N2006, N1959, N534, N1832);
buf BUF1 (N2007, N2005);
and AND2 (N2008, N1997, N387);
nand NAND3 (N2009, N1992, N1010, N1085);
nor NOR2 (N2010, N2009, N564);
buf BUF1 (N2011, N1999);
nand NAND3 (N2012, N2008, N643, N160);
buf BUF1 (N2013, N1996);
not NOT1 (N2014, N2007);
xor XOR2 (N2015, N2012, N1269);
or OR2 (N2016, N2000, N994);
nor NOR4 (N2017, N2013, N1533, N459, N1417);
nor NOR2 (N2018, N2003, N1751);
xor XOR2 (N2019, N2017, N1198);
buf BUF1 (N2020, N1984);
not NOT1 (N2021, N2014);
nor NOR4 (N2022, N2010, N1142, N1066, N1102);
nand NAND4 (N2023, N2015, N1543, N1229, N876);
or OR3 (N2024, N2016, N1254, N1279);
or OR4 (N2025, N2019, N592, N1303, N679);
and AND3 (N2026, N2020, N144, N416);
or OR4 (N2027, N2006, N377, N2008, N259);
xor XOR2 (N2028, N2027, N221);
or OR2 (N2029, N2024, N763);
xor XOR2 (N2030, N2022, N391);
not NOT1 (N2031, N2025);
nand NAND4 (N2032, N2011, N749, N1907, N343);
and AND4 (N2033, N2021, N391, N1584, N839);
nand NAND2 (N2034, N2032, N301);
nor NOR4 (N2035, N2030, N463, N1094, N944);
not NOT1 (N2036, N2028);
nor NOR2 (N2037, N2031, N1631);
xor XOR2 (N2038, N2023, N1715);
nand NAND2 (N2039, N2033, N707);
buf BUF1 (N2040, N2035);
buf BUF1 (N2041, N2036);
nand NAND2 (N2042, N2018, N1288);
and AND3 (N2043, N2041, N1525, N1394);
nor NOR2 (N2044, N2034, N872);
xor XOR2 (N2045, N2040, N681);
nand NAND3 (N2046, N2026, N251, N1257);
xor XOR2 (N2047, N2044, N893);
or OR2 (N2048, N2039, N1405);
not NOT1 (N2049, N2046);
xor XOR2 (N2050, N2038, N561);
buf BUF1 (N2051, N2049);
and AND2 (N2052, N2050, N1785);
not NOT1 (N2053, N2045);
or OR3 (N2054, N2042, N1277, N1930);
nand NAND3 (N2055, N2054, N1664, N1098);
and AND2 (N2056, N2047, N481);
and AND4 (N2057, N2004, N217, N2024, N42);
not NOT1 (N2058, N2057);
not NOT1 (N2059, N2052);
and AND3 (N2060, N2055, N465, N1118);
nand NAND4 (N2061, N2056, N1422, N690, N273);
and AND3 (N2062, N2060, N1950, N1900);
not NOT1 (N2063, N2051);
nand NAND2 (N2064, N2029, N376);
xor XOR2 (N2065, N2043, N862);
and AND4 (N2066, N2064, N1455, N1892, N2027);
xor XOR2 (N2067, N2037, N1077);
nand NAND2 (N2068, N2063, N1398);
or OR4 (N2069, N2061, N240, N3, N1368);
buf BUF1 (N2070, N2068);
not NOT1 (N2071, N2058);
or OR3 (N2072, N2053, N853, N467);
buf BUF1 (N2073, N2062);
nand NAND2 (N2074, N2073, N1945);
nor NOR3 (N2075, N2059, N1962, N245);
nand NAND4 (N2076, N2048, N1818, N1454, N1979);
xor XOR2 (N2077, N2066, N2021);
not NOT1 (N2078, N2077);
nor NOR4 (N2079, N2075, N1127, N1277, N137);
and AND3 (N2080, N2071, N1416, N1395);
xor XOR2 (N2081, N2070, N44);
and AND3 (N2082, N2079, N2059, N2041);
nand NAND4 (N2083, N2082, N1721, N1521, N838);
not NOT1 (N2084, N2076);
nor NOR3 (N2085, N2067, N341, N1378);
buf BUF1 (N2086, N2083);
not NOT1 (N2087, N2072);
and AND2 (N2088, N2084, N361);
buf BUF1 (N2089, N2078);
or OR2 (N2090, N2065, N618);
not NOT1 (N2091, N2074);
buf BUF1 (N2092, N2089);
not NOT1 (N2093, N2069);
nand NAND4 (N2094, N2080, N425, N681, N1820);
not NOT1 (N2095, N2091);
or OR4 (N2096, N2095, N1475, N208, N1239);
or OR2 (N2097, N2081, N1079);
nor NOR3 (N2098, N2087, N419, N1701);
or OR3 (N2099, N2097, N469, N1562);
xor XOR2 (N2100, N2096, N1960);
not NOT1 (N2101, N2099);
buf BUF1 (N2102, N2085);
and AND4 (N2103, N2092, N633, N1663, N1865);
buf BUF1 (N2104, N2088);
nand NAND2 (N2105, N2090, N2065);
nand NAND4 (N2106, N2103, N682, N2013, N2045);
xor XOR2 (N2107, N2100, N1032);
or OR4 (N2108, N2101, N1344, N1383, N1473);
xor XOR2 (N2109, N2102, N17);
buf BUF1 (N2110, N2108);
nand NAND4 (N2111, N2107, N1879, N1350, N1693);
xor XOR2 (N2112, N2105, N621);
xor XOR2 (N2113, N2093, N1959);
or OR4 (N2114, N2094, N2113, N775, N1151);
not NOT1 (N2115, N1367);
buf BUF1 (N2116, N2111);
or OR4 (N2117, N2114, N372, N572, N466);
or OR2 (N2118, N2106, N1996);
not NOT1 (N2119, N2110);
not NOT1 (N2120, N2104);
or OR2 (N2121, N2118, N1047);
or OR2 (N2122, N2109, N1696);
nor NOR3 (N2123, N2120, N480, N793);
not NOT1 (N2124, N2086);
and AND2 (N2125, N2124, N882);
xor XOR2 (N2126, N2112, N64);
buf BUF1 (N2127, N2126);
and AND3 (N2128, N2115, N1310, N937);
nor NOR4 (N2129, N2119, N1506, N1610, N1313);
buf BUF1 (N2130, N2123);
and AND3 (N2131, N2116, N908, N1987);
not NOT1 (N2132, N2125);
nand NAND3 (N2133, N2130, N1263, N1231);
nor NOR3 (N2134, N2128, N555, N1928);
and AND2 (N2135, N2122, N1271);
and AND4 (N2136, N2135, N1522, N114, N1845);
or OR4 (N2137, N2134, N1242, N1851, N1282);
not NOT1 (N2138, N2098);
and AND4 (N2139, N2136, N817, N967, N1539);
or OR2 (N2140, N2129, N974);
buf BUF1 (N2141, N2117);
or OR3 (N2142, N2141, N1834, N281);
and AND3 (N2143, N2139, N994, N524);
xor XOR2 (N2144, N2121, N620);
buf BUF1 (N2145, N2137);
nor NOR4 (N2146, N2142, N474, N648, N88);
not NOT1 (N2147, N2131);
and AND3 (N2148, N2133, N443, N1773);
buf BUF1 (N2149, N2143);
and AND4 (N2150, N2145, N1579, N652, N1731);
or OR3 (N2151, N2148, N1883, N37);
or OR2 (N2152, N2150, N36);
buf BUF1 (N2153, N2132);
buf BUF1 (N2154, N2127);
buf BUF1 (N2155, N2140);
or OR4 (N2156, N2153, N238, N314, N1833);
and AND3 (N2157, N2156, N1604, N1847);
nand NAND2 (N2158, N2151, N2136);
xor XOR2 (N2159, N2158, N476);
or OR3 (N2160, N2146, N1459, N1023);
nand NAND3 (N2161, N2155, N510, N927);
nor NOR2 (N2162, N2161, N1965);
nor NOR4 (N2163, N2149, N1047, N1365, N912);
and AND2 (N2164, N2147, N351);
and AND3 (N2165, N2159, N1524, N1531);
and AND2 (N2166, N2162, N1639);
buf BUF1 (N2167, N2164);
buf BUF1 (N2168, N2152);
and AND4 (N2169, N2165, N518, N1973, N1309);
xor XOR2 (N2170, N2157, N2159);
nor NOR2 (N2171, N2154, N1800);
xor XOR2 (N2172, N2163, N117);
nor NOR2 (N2173, N2166, N551);
and AND3 (N2174, N2144, N1772, N1803);
buf BUF1 (N2175, N2173);
not NOT1 (N2176, N2174);
or OR2 (N2177, N2169, N91);
and AND3 (N2178, N2170, N118, N36);
nor NOR2 (N2179, N2167, N19);
nor NOR4 (N2180, N2178, N707, N654, N926);
or OR3 (N2181, N2138, N271, N534);
or OR3 (N2182, N2172, N61, N1268);
xor XOR2 (N2183, N2177, N1234);
nand NAND2 (N2184, N2182, N1560);
not NOT1 (N2185, N2183);
and AND2 (N2186, N2160, N723);
not NOT1 (N2187, N2181);
and AND3 (N2188, N2176, N473, N639);
nand NAND4 (N2189, N2171, N772, N1980, N900);
nor NOR3 (N2190, N2186, N1519, N543);
nor NOR4 (N2191, N2188, N713, N1356, N1289);
not NOT1 (N2192, N2184);
or OR2 (N2193, N2190, N945);
xor XOR2 (N2194, N2189, N210);
xor XOR2 (N2195, N2175, N1361);
xor XOR2 (N2196, N2179, N1330);
and AND2 (N2197, N2194, N590);
nor NOR2 (N2198, N2195, N57);
and AND4 (N2199, N2198, N1173, N1808, N2026);
and AND2 (N2200, N2185, N646);
xor XOR2 (N2201, N2196, N580);
nand NAND2 (N2202, N2187, N1397);
or OR3 (N2203, N2201, N1884, N1292);
not NOT1 (N2204, N2180);
buf BUF1 (N2205, N2168);
or OR4 (N2206, N2203, N1046, N66, N1140);
and AND4 (N2207, N2202, N1864, N1287, N1694);
or OR3 (N2208, N2205, N2107, N2088);
and AND2 (N2209, N2192, N2014);
buf BUF1 (N2210, N2204);
and AND4 (N2211, N2206, N531, N2100, N308);
and AND3 (N2212, N2211, N1129, N2157);
and AND3 (N2213, N2209, N566, N1549);
xor XOR2 (N2214, N2213, N1182);
not NOT1 (N2215, N2208);
not NOT1 (N2216, N2210);
nor NOR2 (N2217, N2200, N1378);
or OR3 (N2218, N2212, N1879, N461);
and AND4 (N2219, N2217, N1293, N1614, N1671);
and AND3 (N2220, N2207, N1848, N789);
not NOT1 (N2221, N2193);
nor NOR3 (N2222, N2219, N503, N570);
not NOT1 (N2223, N2197);
and AND4 (N2224, N2199, N754, N222, N291);
and AND3 (N2225, N2215, N345, N2146);
buf BUF1 (N2226, N2218);
or OR4 (N2227, N2220, N354, N1647, N844);
or OR3 (N2228, N2226, N2081, N281);
xor XOR2 (N2229, N2216, N1324);
xor XOR2 (N2230, N2222, N317);
xor XOR2 (N2231, N2221, N524);
or OR2 (N2232, N2230, N1107);
nand NAND2 (N2233, N2225, N1250);
not NOT1 (N2234, N2233);
xor XOR2 (N2235, N2191, N1420);
not NOT1 (N2236, N2224);
xor XOR2 (N2237, N2236, N592);
nand NAND3 (N2238, N2229, N1829, N583);
nand NAND2 (N2239, N2234, N955);
nand NAND4 (N2240, N2237, N1552, N1727, N1210);
nor NOR2 (N2241, N2235, N1675);
or OR4 (N2242, N2232, N1026, N1697, N1337);
and AND4 (N2243, N2239, N2235, N1339, N312);
xor XOR2 (N2244, N2231, N2012);
xor XOR2 (N2245, N2238, N751);
and AND2 (N2246, N2243, N1789);
not NOT1 (N2247, N2214);
xor XOR2 (N2248, N2223, N664);
or OR3 (N2249, N2246, N528, N1833);
nand NAND4 (N2250, N2242, N1099, N942, N1435);
nand NAND4 (N2251, N2250, N1744, N1486, N1058);
nand NAND4 (N2252, N2244, N560, N904, N712);
nor NOR4 (N2253, N2241, N134, N197, N823);
xor XOR2 (N2254, N2253, N2150);
and AND2 (N2255, N2249, N1946);
nor NOR4 (N2256, N2240, N830, N90, N700);
or OR3 (N2257, N2248, N752, N1954);
xor XOR2 (N2258, N2256, N709);
xor XOR2 (N2259, N2228, N693);
and AND2 (N2260, N2255, N2143);
nand NAND2 (N2261, N2245, N498);
nor NOR3 (N2262, N2261, N37, N1615);
xor XOR2 (N2263, N2251, N1839);
and AND4 (N2264, N2254, N1045, N1632, N1335);
nand NAND4 (N2265, N2264, N1145, N713, N2064);
nand NAND4 (N2266, N2258, N503, N457, N1888);
and AND4 (N2267, N2266, N2179, N945, N175);
buf BUF1 (N2268, N2267);
buf BUF1 (N2269, N2257);
xor XOR2 (N2270, N2260, N2155);
xor XOR2 (N2271, N2268, N1281);
not NOT1 (N2272, N2252);
or OR2 (N2273, N2269, N882);
buf BUF1 (N2274, N2273);
nor NOR3 (N2275, N2263, N1471, N1040);
buf BUF1 (N2276, N2270);
not NOT1 (N2277, N2262);
and AND4 (N2278, N2274, N594, N389, N555);
buf BUF1 (N2279, N2271);
not NOT1 (N2280, N2247);
buf BUF1 (N2281, N2259);
and AND2 (N2282, N2275, N1176);
nor NOR3 (N2283, N2265, N1314, N558);
and AND3 (N2284, N2279, N671, N224);
buf BUF1 (N2285, N2282);
and AND4 (N2286, N2276, N497, N772, N424);
and AND2 (N2287, N2277, N1018);
nand NAND3 (N2288, N2281, N1701, N1539);
nor NOR3 (N2289, N2283, N1281, N1391);
buf BUF1 (N2290, N2285);
xor XOR2 (N2291, N2272, N1157);
or OR4 (N2292, N2278, N1192, N696, N1116);
or OR3 (N2293, N2292, N2032, N440);
nor NOR4 (N2294, N2291, N2067, N1712, N1130);
nand NAND3 (N2295, N2227, N714, N130);
and AND4 (N2296, N2287, N1459, N607, N250);
xor XOR2 (N2297, N2293, N1627);
and AND3 (N2298, N2297, N637, N2093);
nand NAND2 (N2299, N2295, N2181);
nor NOR2 (N2300, N2284, N1914);
and AND2 (N2301, N2298, N994);
nor NOR3 (N2302, N2288, N692, N1344);
buf BUF1 (N2303, N2290);
or OR3 (N2304, N2299, N736, N333);
buf BUF1 (N2305, N2303);
nor NOR4 (N2306, N2300, N2072, N1584, N196);
buf BUF1 (N2307, N2289);
nand NAND3 (N2308, N2304, N1252, N618);
not NOT1 (N2309, N2305);
not NOT1 (N2310, N2286);
buf BUF1 (N2311, N2310);
nor NOR2 (N2312, N2307, N1175);
or OR2 (N2313, N2312, N817);
not NOT1 (N2314, N2302);
not NOT1 (N2315, N2308);
and AND2 (N2316, N2315, N174);
and AND3 (N2317, N2301, N1215, N1735);
xor XOR2 (N2318, N2314, N836);
and AND3 (N2319, N2311, N176, N6);
buf BUF1 (N2320, N2309);
or OR2 (N2321, N2320, N854);
nand NAND2 (N2322, N2321, N802);
not NOT1 (N2323, N2316);
or OR4 (N2324, N2318, N2128, N654, N1399);
buf BUF1 (N2325, N2296);
xor XOR2 (N2326, N2323, N119);
nor NOR3 (N2327, N2306, N811, N1260);
xor XOR2 (N2328, N2317, N1735);
not NOT1 (N2329, N2280);
not NOT1 (N2330, N2322);
nor NOR4 (N2331, N2325, N2166, N1932, N2178);
nor NOR4 (N2332, N2327, N1357, N2176, N986);
nand NAND2 (N2333, N2332, N1047);
xor XOR2 (N2334, N2326, N2085);
or OR2 (N2335, N2333, N670);
xor XOR2 (N2336, N2313, N1407);
or OR4 (N2337, N2330, N1746, N191, N1448);
nand NAND3 (N2338, N2337, N1817, N1456);
not NOT1 (N2339, N2334);
xor XOR2 (N2340, N2336, N2304);
nand NAND2 (N2341, N2331, N1346);
buf BUF1 (N2342, N2329);
nor NOR4 (N2343, N2294, N1748, N1812, N2319);
not NOT1 (N2344, N840);
not NOT1 (N2345, N2339);
and AND3 (N2346, N2338, N926, N680);
xor XOR2 (N2347, N2342, N2092);
or OR4 (N2348, N2345, N1377, N1027, N1985);
nor NOR4 (N2349, N2347, N968, N1716, N1169);
nand NAND2 (N2350, N2349, N1986);
xor XOR2 (N2351, N2343, N907);
or OR4 (N2352, N2346, N261, N1460, N984);
buf BUF1 (N2353, N2341);
nor NOR4 (N2354, N2350, N1048, N1423, N1338);
buf BUF1 (N2355, N2352);
not NOT1 (N2356, N2324);
xor XOR2 (N2357, N2335, N2264);
or OR2 (N2358, N2351, N2263);
nand NAND4 (N2359, N2358, N1838, N1169, N629);
buf BUF1 (N2360, N2359);
or OR2 (N2361, N2354, N2188);
not NOT1 (N2362, N2348);
nand NAND2 (N2363, N2362, N2144);
or OR2 (N2364, N2360, N2146);
xor XOR2 (N2365, N2340, N613);
nor NOR4 (N2366, N2353, N1179, N1747, N1270);
not NOT1 (N2367, N2361);
buf BUF1 (N2368, N2363);
not NOT1 (N2369, N2368);
xor XOR2 (N2370, N2364, N1007);
buf BUF1 (N2371, N2365);
buf BUF1 (N2372, N2369);
and AND3 (N2373, N2328, N2207, N483);
nor NOR3 (N2374, N2357, N1618, N1859);
or OR2 (N2375, N2356, N600);
and AND2 (N2376, N2367, N402);
and AND2 (N2377, N2371, N1869);
buf BUF1 (N2378, N2366);
not NOT1 (N2379, N2344);
buf BUF1 (N2380, N2372);
and AND2 (N2381, N2374, N406);
xor XOR2 (N2382, N2381, N1663);
or OR4 (N2383, N2355, N1037, N1, N389);
xor XOR2 (N2384, N2370, N780);
nand NAND2 (N2385, N2373, N2140);
nand NAND2 (N2386, N2375, N2277);
nand NAND3 (N2387, N2380, N2092, N558);
and AND2 (N2388, N2384, N148);
buf BUF1 (N2389, N2376);
buf BUF1 (N2390, N2388);
not NOT1 (N2391, N2389);
buf BUF1 (N2392, N2391);
and AND4 (N2393, N2392, N2176, N1821, N1842);
buf BUF1 (N2394, N2383);
nor NOR2 (N2395, N2386, N2167);
not NOT1 (N2396, N2378);
not NOT1 (N2397, N2396);
nand NAND3 (N2398, N2394, N952, N1136);
buf BUF1 (N2399, N2390);
nand NAND2 (N2400, N2385, N1872);
not NOT1 (N2401, N2398);
or OR3 (N2402, N2387, N2114, N2339);
nand NAND2 (N2403, N2401, N342);
buf BUF1 (N2404, N2395);
nor NOR4 (N2405, N2404, N1851, N1624, N1749);
nor NOR2 (N2406, N2379, N438);
nand NAND4 (N2407, N2406, N753, N914, N1195);
buf BUF1 (N2408, N2403);
or OR3 (N2409, N2407, N1839, N2019);
buf BUF1 (N2410, N2382);
buf BUF1 (N2411, N2393);
buf BUF1 (N2412, N2400);
buf BUF1 (N2413, N2409);
or OR3 (N2414, N2410, N1933, N613);
or OR3 (N2415, N2399, N1201, N1317);
xor XOR2 (N2416, N2408, N1685);
and AND3 (N2417, N2415, N696, N1354);
or OR4 (N2418, N2414, N2052, N1678, N989);
and AND2 (N2419, N2412, N736);
or OR2 (N2420, N2411, N210);
nand NAND3 (N2421, N2418, N1343, N2193);
nand NAND2 (N2422, N2402, N1851);
xor XOR2 (N2423, N2416, N136);
or OR4 (N2424, N2420, N349, N1296, N2330);
xor XOR2 (N2425, N2421, N441);
nand NAND4 (N2426, N2424, N1964, N71, N1291);
xor XOR2 (N2427, N2397, N512);
nand NAND2 (N2428, N2426, N869);
nand NAND2 (N2429, N2425, N134);
not NOT1 (N2430, N2417);
not NOT1 (N2431, N2430);
buf BUF1 (N2432, N2431);
nand NAND2 (N2433, N2427, N1344);
and AND4 (N2434, N2432, N1653, N133, N29);
buf BUF1 (N2435, N2429);
or OR2 (N2436, N2434, N1884);
nand NAND4 (N2437, N2433, N1275, N335, N146);
nor NOR3 (N2438, N2428, N500, N2076);
and AND2 (N2439, N2405, N919);
buf BUF1 (N2440, N2423);
and AND3 (N2441, N2436, N207, N1147);
buf BUF1 (N2442, N2377);
and AND2 (N2443, N2441, N2010);
nor NOR4 (N2444, N2442, N1024, N440, N1363);
and AND3 (N2445, N2444, N27, N2029);
buf BUF1 (N2446, N2440);
and AND3 (N2447, N2446, N348, N1336);
buf BUF1 (N2448, N2413);
xor XOR2 (N2449, N2437, N1121);
buf BUF1 (N2450, N2449);
nor NOR3 (N2451, N2443, N1436, N36);
buf BUF1 (N2452, N2447);
and AND3 (N2453, N2452, N2086, N274);
buf BUF1 (N2454, N2450);
nand NAND3 (N2455, N2454, N405, N1222);
xor XOR2 (N2456, N2455, N266);
xor XOR2 (N2457, N2435, N1865);
or OR3 (N2458, N2453, N1770, N267);
buf BUF1 (N2459, N2445);
xor XOR2 (N2460, N2448, N466);
and AND4 (N2461, N2439, N1383, N668, N1092);
buf BUF1 (N2462, N2458);
not NOT1 (N2463, N2459);
nor NOR2 (N2464, N2461, N944);
nor NOR2 (N2465, N2422, N1592);
xor XOR2 (N2466, N2438, N624);
xor XOR2 (N2467, N2462, N514);
nor NOR2 (N2468, N2464, N1890);
xor XOR2 (N2469, N2465, N927);
or OR3 (N2470, N2469, N1271, N2418);
nand NAND3 (N2471, N2468, N263, N2456);
not NOT1 (N2472, N1791);
buf BUF1 (N2473, N2419);
nand NAND2 (N2474, N2473, N904);
not NOT1 (N2475, N2467);
nand NAND4 (N2476, N2451, N535, N2249, N981);
nor NOR4 (N2477, N2460, N2328, N2144, N1003);
or OR2 (N2478, N2470, N1290);
and AND2 (N2479, N2477, N2288);
xor XOR2 (N2480, N2474, N1977);
nand NAND3 (N2481, N2478, N2468, N1970);
xor XOR2 (N2482, N2480, N234);
and AND3 (N2483, N2471, N2219, N717);
buf BUF1 (N2484, N2472);
xor XOR2 (N2485, N2466, N2116);
nand NAND2 (N2486, N2479, N1654);
buf BUF1 (N2487, N2475);
nor NOR3 (N2488, N2487, N463, N1156);
not NOT1 (N2489, N2482);
nor NOR4 (N2490, N2463, N1112, N1411, N1350);
buf BUF1 (N2491, N2484);
and AND3 (N2492, N2488, N699, N1355);
nand NAND3 (N2493, N2490, N1427, N2027);
xor XOR2 (N2494, N2481, N737);
xor XOR2 (N2495, N2457, N477);
buf BUF1 (N2496, N2491);
or OR4 (N2497, N2492, N2383, N1741, N1535);
not NOT1 (N2498, N2495);
buf BUF1 (N2499, N2485);
not NOT1 (N2500, N2496);
xor XOR2 (N2501, N2498, N2257);
or OR3 (N2502, N2501, N1406, N485);
nor NOR3 (N2503, N2497, N2110, N2322);
buf BUF1 (N2504, N2489);
xor XOR2 (N2505, N2503, N2263);
not NOT1 (N2506, N2476);
or OR3 (N2507, N2506, N2298, N2080);
buf BUF1 (N2508, N2486);
nor NOR2 (N2509, N2502, N272);
nand NAND3 (N2510, N2483, N221, N1318);
or OR2 (N2511, N2505, N1296);
or OR3 (N2512, N2511, N4, N1907);
nor NOR4 (N2513, N2499, N277, N2195, N1887);
not NOT1 (N2514, N2504);
nand NAND4 (N2515, N2500, N1655, N307, N2311);
and AND2 (N2516, N2515, N2205);
xor XOR2 (N2517, N2494, N2415);
buf BUF1 (N2518, N2510);
nor NOR3 (N2519, N2513, N1899, N413);
buf BUF1 (N2520, N2507);
not NOT1 (N2521, N2509);
xor XOR2 (N2522, N2493, N313);
buf BUF1 (N2523, N2517);
nand NAND2 (N2524, N2512, N266);
and AND4 (N2525, N2524, N858, N1841, N999);
nor NOR4 (N2526, N2508, N1415, N766, N1234);
xor XOR2 (N2527, N2518, N1190);
buf BUF1 (N2528, N2526);
or OR3 (N2529, N2521, N1502, N372);
or OR2 (N2530, N2522, N2136);
and AND4 (N2531, N2523, N2362, N2411, N1956);
not NOT1 (N2532, N2528);
and AND4 (N2533, N2529, N2367, N1010, N366);
xor XOR2 (N2534, N2519, N546);
not NOT1 (N2535, N2516);
and AND4 (N2536, N2534, N1887, N2501, N1709);
nand NAND4 (N2537, N2530, N1522, N1761, N710);
buf BUF1 (N2538, N2525);
and AND2 (N2539, N2527, N1217);
nor NOR4 (N2540, N2535, N2389, N2441, N951);
and AND4 (N2541, N2539, N2305, N1149, N2514);
buf BUF1 (N2542, N693);
not NOT1 (N2543, N2520);
nand NAND3 (N2544, N2543, N1696, N177);
or OR4 (N2545, N2544, N294, N1608, N2354);
xor XOR2 (N2546, N2540, N1132);
buf BUF1 (N2547, N2533);
nand NAND4 (N2548, N2547, N409, N1522, N646);
nor NOR2 (N2549, N2541, N1610);
or OR4 (N2550, N2538, N1853, N1756, N127);
nor NOR4 (N2551, N2546, N320, N667, N301);
and AND4 (N2552, N2548, N352, N292, N2339);
xor XOR2 (N2553, N2536, N2340);
and AND4 (N2554, N2553, N954, N1665, N2043);
nand NAND3 (N2555, N2554, N2498, N842);
buf BUF1 (N2556, N2552);
or OR4 (N2557, N2556, N1853, N1820, N1131);
not NOT1 (N2558, N2555);
not NOT1 (N2559, N2531);
xor XOR2 (N2560, N2550, N2550);
and AND2 (N2561, N2558, N1028);
and AND3 (N2562, N2545, N1471, N194);
not NOT1 (N2563, N2542);
or OR2 (N2564, N2537, N1893);
nor NOR2 (N2565, N2560, N2421);
or OR2 (N2566, N2564, N1977);
nand NAND3 (N2567, N2562, N1301, N1998);
not NOT1 (N2568, N2567);
or OR2 (N2569, N2549, N50);
and AND4 (N2570, N2569, N1038, N1783, N1297);
nand NAND4 (N2571, N2559, N2042, N423, N220);
and AND2 (N2572, N2557, N1445);
nor NOR2 (N2573, N2565, N302);
and AND4 (N2574, N2561, N1466, N2537, N2232);
nor NOR2 (N2575, N2571, N816);
buf BUF1 (N2576, N2532);
xor XOR2 (N2577, N2563, N709);
or OR4 (N2578, N2572, N644, N1112, N376);
buf BUF1 (N2579, N2573);
and AND4 (N2580, N2574, N891, N2177, N282);
nor NOR2 (N2581, N2578, N693);
not NOT1 (N2582, N2581);
buf BUF1 (N2583, N2566);
nor NOR2 (N2584, N2570, N2441);
xor XOR2 (N2585, N2583, N574);
or OR2 (N2586, N2579, N104);
buf BUF1 (N2587, N2575);
or OR3 (N2588, N2582, N1343, N877);
xor XOR2 (N2589, N2584, N735);
nor NOR3 (N2590, N2586, N1108, N2077);
xor XOR2 (N2591, N2576, N546);
not NOT1 (N2592, N2590);
not NOT1 (N2593, N2589);
nor NOR2 (N2594, N2592, N49);
nand NAND4 (N2595, N2587, N2141, N1656, N2004);
and AND4 (N2596, N2551, N1830, N593, N2500);
and AND2 (N2597, N2593, N1087);
and AND2 (N2598, N2577, N1269);
xor XOR2 (N2599, N2580, N1198);
not NOT1 (N2600, N2594);
not NOT1 (N2601, N2599);
and AND4 (N2602, N2588, N1633, N1656, N2409);
not NOT1 (N2603, N2585);
nor NOR3 (N2604, N2597, N1207, N794);
not NOT1 (N2605, N2568);
nand NAND3 (N2606, N2591, N576, N137);
nor NOR3 (N2607, N2604, N995, N384);
buf BUF1 (N2608, N2606);
xor XOR2 (N2609, N2601, N1280);
nand NAND3 (N2610, N2596, N1890, N1952);
nor NOR2 (N2611, N2598, N2257);
buf BUF1 (N2612, N2609);
xor XOR2 (N2613, N2602, N1392);
buf BUF1 (N2614, N2607);
xor XOR2 (N2615, N2605, N978);
buf BUF1 (N2616, N2600);
and AND2 (N2617, N2614, N1767);
or OR4 (N2618, N2613, N2373, N896, N573);
not NOT1 (N2619, N2611);
or OR2 (N2620, N2618, N293);
and AND2 (N2621, N2620, N1476);
xor XOR2 (N2622, N2616, N105);
not NOT1 (N2623, N2608);
and AND4 (N2624, N2617, N97, N1439, N623);
and AND4 (N2625, N2615, N2548, N191, N323);
buf BUF1 (N2626, N2603);
nand NAND4 (N2627, N2624, N453, N2191, N488);
xor XOR2 (N2628, N2623, N850);
nand NAND3 (N2629, N2628, N1938, N1619);
not NOT1 (N2630, N2621);
not NOT1 (N2631, N2625);
xor XOR2 (N2632, N2626, N501);
and AND3 (N2633, N2622, N1595, N862);
buf BUF1 (N2634, N2627);
xor XOR2 (N2635, N2631, N148);
buf BUF1 (N2636, N2610);
nor NOR4 (N2637, N2619, N597, N1849, N1972);
and AND3 (N2638, N2634, N1965, N1205);
not NOT1 (N2639, N2636);
nor NOR3 (N2640, N2633, N634, N108);
or OR2 (N2641, N2630, N552);
xor XOR2 (N2642, N2641, N599);
or OR2 (N2643, N2632, N364);
nand NAND3 (N2644, N2638, N1851, N560);
or OR4 (N2645, N2644, N2104, N2438, N1016);
xor XOR2 (N2646, N2645, N2110);
buf BUF1 (N2647, N2640);
buf BUF1 (N2648, N2595);
or OR3 (N2649, N2637, N2200, N1945);
or OR2 (N2650, N2646, N875);
xor XOR2 (N2651, N2650, N1281);
buf BUF1 (N2652, N2643);
buf BUF1 (N2653, N2647);
and AND2 (N2654, N2642, N865);
buf BUF1 (N2655, N2648);
buf BUF1 (N2656, N2655);
and AND2 (N2657, N2629, N2385);
or OR3 (N2658, N2639, N2242, N494);
and AND2 (N2659, N2651, N785);
buf BUF1 (N2660, N2635);
xor XOR2 (N2661, N2659, N173);
not NOT1 (N2662, N2612);
or OR2 (N2663, N2662, N2018);
and AND3 (N2664, N2654, N1544, N2226);
nand NAND4 (N2665, N2661, N2399, N235, N1632);
nand NAND3 (N2666, N2656, N2451, N1031);
buf BUF1 (N2667, N2652);
or OR2 (N2668, N2657, N2513);
or OR4 (N2669, N2668, N2481, N2262, N2211);
nor NOR2 (N2670, N2649, N1674);
nor NOR4 (N2671, N2665, N2311, N343, N2309);
not NOT1 (N2672, N2667);
or OR4 (N2673, N2653, N2633, N1039, N1920);
or OR3 (N2674, N2663, N2152, N2384);
and AND4 (N2675, N2671, N713, N621, N157);
xor XOR2 (N2676, N2658, N847);
buf BUF1 (N2677, N2670);
xor XOR2 (N2678, N2672, N397);
and AND4 (N2679, N2675, N783, N861, N1464);
or OR3 (N2680, N2669, N1889, N2146);
nor NOR4 (N2681, N2664, N698, N1074, N1354);
not NOT1 (N2682, N2681);
or OR4 (N2683, N2674, N1418, N2414, N949);
xor XOR2 (N2684, N2660, N1162);
not NOT1 (N2685, N2677);
nand NAND2 (N2686, N2685, N242);
xor XOR2 (N2687, N2676, N2381);
buf BUF1 (N2688, N2684);
nand NAND4 (N2689, N2686, N1711, N2468, N559);
or OR4 (N2690, N2688, N445, N2225, N2519);
nand NAND4 (N2691, N2680, N2280, N1151, N1434);
or OR4 (N2692, N2673, N1580, N792, N2594);
nand NAND3 (N2693, N2683, N2275, N431);
buf BUF1 (N2694, N2678);
or OR2 (N2695, N2690, N1800);
or OR3 (N2696, N2689, N2136, N1754);
not NOT1 (N2697, N2666);
xor XOR2 (N2698, N2697, N1024);
xor XOR2 (N2699, N2682, N2450);
and AND3 (N2700, N2687, N2062, N1034);
buf BUF1 (N2701, N2679);
nor NOR3 (N2702, N2695, N2006, N471);
buf BUF1 (N2703, N2691);
nand NAND4 (N2704, N2699, N1694, N1448, N919);
xor XOR2 (N2705, N2704, N1800);
or OR3 (N2706, N2696, N217, N1812);
xor XOR2 (N2707, N2701, N1578);
buf BUF1 (N2708, N2702);
xor XOR2 (N2709, N2707, N2258);
xor XOR2 (N2710, N2700, N483);
nor NOR2 (N2711, N2703, N1965);
buf BUF1 (N2712, N2705);
nor NOR2 (N2713, N2710, N356);
nor NOR2 (N2714, N2693, N916);
nor NOR2 (N2715, N2694, N207);
or OR2 (N2716, N2715, N1515);
nor NOR3 (N2717, N2711, N2394, N2615);
nand NAND3 (N2718, N2698, N1724, N1167);
and AND3 (N2719, N2706, N922, N181);
buf BUF1 (N2720, N2719);
nor NOR3 (N2721, N2720, N2312, N202);
or OR3 (N2722, N2708, N1501, N754);
buf BUF1 (N2723, N2692);
and AND4 (N2724, N2723, N897, N958, N481);
xor XOR2 (N2725, N2724, N868);
or OR3 (N2726, N2721, N2676, N285);
buf BUF1 (N2727, N2726);
xor XOR2 (N2728, N2718, N254);
xor XOR2 (N2729, N2722, N1521);
xor XOR2 (N2730, N2713, N1637);
and AND4 (N2731, N2728, N1262, N254, N1275);
xor XOR2 (N2732, N2731, N1796);
buf BUF1 (N2733, N2714);
nand NAND3 (N2734, N2716, N225, N763);
buf BUF1 (N2735, N2730);
not NOT1 (N2736, N2727);
buf BUF1 (N2737, N2736);
not NOT1 (N2738, N2717);
buf BUF1 (N2739, N2725);
nand NAND2 (N2740, N2735, N747);
xor XOR2 (N2741, N2729, N1801);
buf BUF1 (N2742, N2741);
or OR3 (N2743, N2709, N1838, N1997);
not NOT1 (N2744, N2742);
not NOT1 (N2745, N2740);
buf BUF1 (N2746, N2737);
buf BUF1 (N2747, N2744);
nor NOR2 (N2748, N2738, N2600);
or OR4 (N2749, N2743, N1746, N279, N2097);
or OR3 (N2750, N2746, N2180, N690);
not NOT1 (N2751, N2748);
not NOT1 (N2752, N2732);
nor NOR4 (N2753, N2733, N1810, N2087, N2525);
buf BUF1 (N2754, N2739);
or OR3 (N2755, N2752, N2109, N2650);
nand NAND2 (N2756, N2712, N2091);
not NOT1 (N2757, N2751);
or OR3 (N2758, N2753, N1434, N617);
and AND3 (N2759, N2758, N2525, N2560);
xor XOR2 (N2760, N2749, N446);
nand NAND2 (N2761, N2755, N1776);
or OR3 (N2762, N2745, N584, N86);
or OR2 (N2763, N2762, N33);
and AND2 (N2764, N2763, N957);
xor XOR2 (N2765, N2764, N2316);
not NOT1 (N2766, N2765);
not NOT1 (N2767, N2760);
buf BUF1 (N2768, N2747);
buf BUF1 (N2769, N2750);
not NOT1 (N2770, N2734);
nor NOR2 (N2771, N2767, N1655);
xor XOR2 (N2772, N2757, N2684);
nand NAND2 (N2773, N2769, N500);
xor XOR2 (N2774, N2754, N653);
or OR4 (N2775, N2761, N411, N706, N2095);
xor XOR2 (N2776, N2756, N2501);
not NOT1 (N2777, N2759);
nor NOR3 (N2778, N2776, N1790, N2588);
xor XOR2 (N2779, N2775, N1852);
xor XOR2 (N2780, N2771, N1206);
and AND4 (N2781, N2780, N337, N1521, N2275);
and AND2 (N2782, N2778, N1015);
nor NOR2 (N2783, N2781, N1804);
and AND4 (N2784, N2768, N1433, N2236, N1080);
nand NAND3 (N2785, N2766, N1353, N2582);
or OR2 (N2786, N2773, N103);
xor XOR2 (N2787, N2786, N1552);
nand NAND3 (N2788, N2787, N1128, N1148);
nor NOR3 (N2789, N2777, N1621, N41);
not NOT1 (N2790, N2785);
nor NOR3 (N2791, N2784, N2323, N2213);
or OR4 (N2792, N2788, N1730, N1681, N2575);
xor XOR2 (N2793, N2790, N876);
buf BUF1 (N2794, N2789);
nor NOR2 (N2795, N2772, N1228);
not NOT1 (N2796, N2770);
and AND2 (N2797, N2782, N952);
nor NOR4 (N2798, N2783, N2570, N2097, N2131);
nor NOR2 (N2799, N2794, N2544);
not NOT1 (N2800, N2791);
buf BUF1 (N2801, N2797);
and AND4 (N2802, N2796, N973, N776, N159);
not NOT1 (N2803, N2799);
xor XOR2 (N2804, N2779, N170);
xor XOR2 (N2805, N2795, N372);
not NOT1 (N2806, N2804);
buf BUF1 (N2807, N2806);
buf BUF1 (N2808, N2800);
nand NAND3 (N2809, N2803, N2801, N2221);
or OR2 (N2810, N413, N2488);
nand NAND3 (N2811, N2809, N937, N1410);
not NOT1 (N2812, N2802);
xor XOR2 (N2813, N2798, N800);
nand NAND4 (N2814, N2813, N2232, N1448, N1236);
buf BUF1 (N2815, N2812);
and AND2 (N2816, N2792, N619);
or OR2 (N2817, N2815, N1647);
xor XOR2 (N2818, N2774, N1122);
or OR3 (N2819, N2817, N74, N347);
and AND4 (N2820, N2818, N183, N1760, N1082);
not NOT1 (N2821, N2807);
nor NOR3 (N2822, N2811, N1639, N1263);
nand NAND4 (N2823, N2814, N2195, N1399, N574);
buf BUF1 (N2824, N2821);
nor NOR4 (N2825, N2808, N824, N1942, N498);
not NOT1 (N2826, N2810);
nor NOR4 (N2827, N2805, N2246, N1192, N1746);
buf BUF1 (N2828, N2827);
and AND4 (N2829, N2825, N2143, N1291, N1182);
nor NOR4 (N2830, N2816, N1970, N1598, N1086);
or OR2 (N2831, N2828, N732);
not NOT1 (N2832, N2822);
buf BUF1 (N2833, N2830);
and AND4 (N2834, N2820, N1309, N2294, N1067);
and AND4 (N2835, N2831, N2423, N906, N838);
and AND2 (N2836, N2826, N2366);
xor XOR2 (N2837, N2829, N1013);
buf BUF1 (N2838, N2836);
and AND2 (N2839, N2834, N1949);
nor NOR3 (N2840, N2819, N1215, N978);
xor XOR2 (N2841, N2837, N1389);
not NOT1 (N2842, N2833);
not NOT1 (N2843, N2839);
buf BUF1 (N2844, N2841);
xor XOR2 (N2845, N2843, N1739);
and AND3 (N2846, N2793, N998, N1286);
nor NOR3 (N2847, N2835, N2014, N306);
nor NOR4 (N2848, N2824, N1653, N852, N262);
xor XOR2 (N2849, N2845, N1129);
and AND4 (N2850, N2849, N2008, N233, N1641);
not NOT1 (N2851, N2846);
buf BUF1 (N2852, N2823);
nor NOR3 (N2853, N2840, N1120, N300);
and AND4 (N2854, N2850, N1179, N1164, N2099);
xor XOR2 (N2855, N2854, N2265);
nand NAND3 (N2856, N2847, N2038, N1038);
not NOT1 (N2857, N2852);
nor NOR4 (N2858, N2844, N482, N2530, N1745);
buf BUF1 (N2859, N2848);
nand NAND3 (N2860, N2838, N2, N2415);
nand NAND2 (N2861, N2859, N272);
buf BUF1 (N2862, N2842);
nor NOR4 (N2863, N2861, N665, N1551, N1840);
buf BUF1 (N2864, N2856);
and AND3 (N2865, N2855, N486, N2366);
or OR2 (N2866, N2860, N2398);
buf BUF1 (N2867, N2858);
nor NOR3 (N2868, N2865, N1463, N1602);
not NOT1 (N2869, N2866);
buf BUF1 (N2870, N2863);
not NOT1 (N2871, N2868);
not NOT1 (N2872, N2864);
nor NOR2 (N2873, N2867, N1881);
or OR4 (N2874, N2869, N1231, N339, N1354);
or OR4 (N2875, N2874, N1279, N847, N288);
or OR4 (N2876, N2871, N305, N1765, N457);
buf BUF1 (N2877, N2857);
nand NAND4 (N2878, N2875, N587, N2611, N1272);
xor XOR2 (N2879, N2873, N1348);
and AND3 (N2880, N2851, N2350, N491);
nor NOR2 (N2881, N2880, N1866);
nor NOR3 (N2882, N2870, N1151, N1449);
nand NAND3 (N2883, N2853, N1835, N2645);
or OR2 (N2884, N2879, N1530);
nand NAND4 (N2885, N2876, N110, N2663, N153);
nor NOR3 (N2886, N2881, N1232, N2100);
not NOT1 (N2887, N2877);
and AND2 (N2888, N2886, N235);
xor XOR2 (N2889, N2862, N838);
buf BUF1 (N2890, N2872);
nand NAND3 (N2891, N2888, N1332, N2429);
xor XOR2 (N2892, N2878, N2677);
not NOT1 (N2893, N2883);
and AND3 (N2894, N2890, N2327, N1408);
xor XOR2 (N2895, N2893, N2293);
or OR4 (N2896, N2889, N2154, N413, N2252);
nand NAND2 (N2897, N2885, N20);
and AND3 (N2898, N2894, N124, N14);
and AND3 (N2899, N2882, N2395, N535);
and AND3 (N2900, N2896, N2797, N1318);
not NOT1 (N2901, N2832);
nor NOR3 (N2902, N2892, N947, N2133);
buf BUF1 (N2903, N2899);
buf BUF1 (N2904, N2900);
nor NOR2 (N2905, N2898, N849);
buf BUF1 (N2906, N2902);
nand NAND2 (N2907, N2903, N867);
nor NOR4 (N2908, N2904, N1611, N2232, N2387);
nor NOR4 (N2909, N2901, N2047, N2906, N2731);
and AND3 (N2910, N1837, N1087, N2103);
nand NAND3 (N2911, N2909, N355, N244);
and AND2 (N2912, N2884, N83);
buf BUF1 (N2913, N2887);
xor XOR2 (N2914, N2908, N612);
nand NAND3 (N2915, N2891, N1118, N1885);
and AND4 (N2916, N2907, N1667, N1284, N2002);
nand NAND2 (N2917, N2916, N2773);
xor XOR2 (N2918, N2895, N827);
and AND4 (N2919, N2917, N2241, N2531, N148);
or OR2 (N2920, N2914, N2594);
xor XOR2 (N2921, N2915, N817);
not NOT1 (N2922, N2919);
xor XOR2 (N2923, N2921, N1030);
nand NAND2 (N2924, N2912, N725);
nor NOR4 (N2925, N2897, N2533, N1731, N2390);
and AND3 (N2926, N2913, N859, N1803);
nand NAND4 (N2927, N2918, N1438, N661, N16);
and AND3 (N2928, N2910, N667, N247);
buf BUF1 (N2929, N2920);
nand NAND4 (N2930, N2924, N2642, N703, N773);
xor XOR2 (N2931, N2925, N2856);
buf BUF1 (N2932, N2930);
not NOT1 (N2933, N2931);
nand NAND4 (N2934, N2905, N563, N2839, N1801);
or OR4 (N2935, N2932, N2226, N2205, N1846);
xor XOR2 (N2936, N2928, N2101);
and AND4 (N2937, N2923, N814, N2657, N308);
nor NOR4 (N2938, N2935, N2077, N2517, N2069);
buf BUF1 (N2939, N2936);
nand NAND2 (N2940, N2926, N609);
not NOT1 (N2941, N2937);
not NOT1 (N2942, N2922);
nor NOR4 (N2943, N2942, N2835, N2523, N2419);
nand NAND4 (N2944, N2929, N282, N635, N788);
and AND3 (N2945, N2939, N635, N2071);
nand NAND3 (N2946, N2944, N2871, N2369);
xor XOR2 (N2947, N2940, N2403);
nor NOR3 (N2948, N2945, N1787, N364);
or OR4 (N2949, N2946, N1478, N434, N2077);
not NOT1 (N2950, N2911);
buf BUF1 (N2951, N2933);
buf BUF1 (N2952, N2943);
buf BUF1 (N2953, N2927);
and AND3 (N2954, N2938, N2659, N1220);
and AND2 (N2955, N2954, N2727);
nand NAND3 (N2956, N2951, N2312, N1667);
or OR4 (N2957, N2949, N122, N1494, N1196);
or OR3 (N2958, N2953, N2214, N2169);
and AND3 (N2959, N2948, N1802, N1888);
or OR3 (N2960, N2941, N527, N1961);
not NOT1 (N2961, N2950);
not NOT1 (N2962, N2958);
nand NAND4 (N2963, N2934, N2414, N2112, N1969);
xor XOR2 (N2964, N2957, N1973);
nor NOR3 (N2965, N2947, N1498, N2711);
nand NAND4 (N2966, N2961, N2705, N272, N2225);
not NOT1 (N2967, N2965);
nor NOR4 (N2968, N2966, N2155, N395, N2310);
buf BUF1 (N2969, N2956);
or OR2 (N2970, N2962, N2329);
not NOT1 (N2971, N2964);
or OR2 (N2972, N2969, N2490);
buf BUF1 (N2973, N2968);
nor NOR2 (N2974, N2963, N1352);
and AND4 (N2975, N2972, N1286, N1369, N1517);
not NOT1 (N2976, N2970);
xor XOR2 (N2977, N2952, N1581);
or OR4 (N2978, N2971, N1371, N171, N1751);
nand NAND2 (N2979, N2959, N1905);
and AND2 (N2980, N2973, N1157);
nand NAND2 (N2981, N2960, N1205);
and AND3 (N2982, N2974, N579, N70);
or OR4 (N2983, N2982, N1901, N2490, N1994);
or OR3 (N2984, N2980, N2230, N839);
xor XOR2 (N2985, N2978, N1391);
nand NAND2 (N2986, N2979, N161);
nor NOR3 (N2987, N2955, N1493, N2979);
buf BUF1 (N2988, N2975);
and AND3 (N2989, N2977, N2902, N2565);
or OR3 (N2990, N2983, N1196, N942);
nor NOR2 (N2991, N2985, N2310);
xor XOR2 (N2992, N2981, N558);
buf BUF1 (N2993, N2976);
nor NOR4 (N2994, N2989, N382, N2548, N1093);
nand NAND4 (N2995, N2986, N1294, N1069, N1001);
or OR4 (N2996, N2993, N1552, N640, N709);
not NOT1 (N2997, N2967);
nor NOR3 (N2998, N2992, N711, N2324);
nand NAND3 (N2999, N2984, N2218, N116);
and AND4 (N3000, N2990, N1148, N2363, N1934);
not NOT1 (N3001, N3000);
buf BUF1 (N3002, N3001);
and AND2 (N3003, N3002, N470);
or OR4 (N3004, N2999, N2979, N285, N2892);
xor XOR2 (N3005, N3003, N928);
and AND4 (N3006, N2994, N2630, N1719, N1009);
and AND3 (N3007, N3006, N2982, N682);
or OR3 (N3008, N2996, N2090, N817);
not NOT1 (N3009, N3008);
not NOT1 (N3010, N2998);
nand NAND4 (N3011, N2987, N1195, N937, N2465);
or OR2 (N3012, N3005, N2822);
buf BUF1 (N3013, N3007);
or OR4 (N3014, N3011, N995, N1808, N1824);
not NOT1 (N3015, N3004);
not NOT1 (N3016, N3015);
nor NOR4 (N3017, N3013, N2088, N201, N743);
and AND2 (N3018, N3012, N510);
not NOT1 (N3019, N3016);
nand NAND2 (N3020, N3014, N2216);
xor XOR2 (N3021, N3019, N535);
buf BUF1 (N3022, N2997);
not NOT1 (N3023, N3020);
nand NAND2 (N3024, N2988, N114);
not NOT1 (N3025, N3022);
and AND4 (N3026, N2991, N2886, N172, N2193);
nor NOR2 (N3027, N3023, N1212);
nor NOR4 (N3028, N3018, N1063, N24, N2616);
not NOT1 (N3029, N2995);
and AND2 (N3030, N3010, N1583);
nor NOR4 (N3031, N3027, N1090, N1962, N1041);
nand NAND4 (N3032, N3009, N1789, N1778, N585);
not NOT1 (N3033, N3021);
or OR3 (N3034, N3028, N1771, N1662);
and AND3 (N3035, N3017, N639, N1302);
and AND2 (N3036, N3032, N2466);
or OR2 (N3037, N3035, N2894);
nand NAND3 (N3038, N3025, N2591, N1748);
xor XOR2 (N3039, N3029, N1354);
nand NAND3 (N3040, N3030, N1742, N883);
xor XOR2 (N3041, N3026, N1382);
and AND3 (N3042, N3033, N2303, N1846);
buf BUF1 (N3043, N3034);
or OR2 (N3044, N3041, N2101);
nor NOR2 (N3045, N3044, N295);
nand NAND2 (N3046, N3031, N2030);
or OR3 (N3047, N3024, N2499, N2915);
buf BUF1 (N3048, N3043);
or OR4 (N3049, N3036, N3030, N386, N2361);
or OR2 (N3050, N3046, N1075);
not NOT1 (N3051, N3045);
nor NOR2 (N3052, N3042, N1091);
not NOT1 (N3053, N3039);
and AND2 (N3054, N3052, N1354);
nand NAND4 (N3055, N3038, N1010, N166, N3038);
and AND4 (N3056, N3051, N1579, N979, N2407);
or OR4 (N3057, N3047, N1555, N420, N3037);
buf BUF1 (N3058, N2041);
and AND2 (N3059, N3049, N431);
xor XOR2 (N3060, N3057, N259);
or OR4 (N3061, N3056, N1868, N2185, N246);
xor XOR2 (N3062, N3054, N944);
not NOT1 (N3063, N3061);
nor NOR4 (N3064, N3055, N2233, N2598, N1318);
and AND4 (N3065, N3048, N2965, N2058, N2678);
buf BUF1 (N3066, N3040);
and AND2 (N3067, N3062, N1477);
buf BUF1 (N3068, N3050);
not NOT1 (N3069, N3068);
nor NOR4 (N3070, N3065, N2417, N39, N2942);
not NOT1 (N3071, N3069);
not NOT1 (N3072, N3070);
nand NAND3 (N3073, N3063, N688, N396);
buf BUF1 (N3074, N3067);
nor NOR2 (N3075, N3071, N829);
buf BUF1 (N3076, N3059);
not NOT1 (N3077, N3060);
nand NAND3 (N3078, N3076, N473, N2712);
nand NAND2 (N3079, N3074, N1030);
and AND4 (N3080, N3058, N663, N1795, N2997);
not NOT1 (N3081, N3053);
nor NOR2 (N3082, N3081, N1509);
buf BUF1 (N3083, N3077);
and AND4 (N3084, N3064, N563, N1275, N1748);
and AND4 (N3085, N3084, N663, N2367, N2738);
and AND3 (N3086, N3075, N1683, N1780);
nor NOR3 (N3087, N3082, N3031, N2519);
not NOT1 (N3088, N3087);
xor XOR2 (N3089, N3079, N1361);
and AND3 (N3090, N3083, N1987, N3062);
not NOT1 (N3091, N3090);
buf BUF1 (N3092, N3073);
or OR2 (N3093, N3089, N360);
and AND3 (N3094, N3088, N1802, N2930);
xor XOR2 (N3095, N3086, N144);
nor NOR4 (N3096, N3093, N1486, N70, N2442);
nand NAND3 (N3097, N3096, N1202, N615);
and AND2 (N3098, N3080, N1630);
or OR2 (N3099, N3097, N702);
not NOT1 (N3100, N3092);
buf BUF1 (N3101, N3066);
and AND3 (N3102, N3091, N859, N1031);
or OR3 (N3103, N3100, N501, N728);
nand NAND4 (N3104, N3101, N1407, N2499, N2810);
and AND3 (N3105, N3078, N1278, N1387);
or OR3 (N3106, N3094, N2119, N893);
or OR4 (N3107, N3099, N1420, N1279, N1017);
xor XOR2 (N3108, N3104, N2330);
not NOT1 (N3109, N3108);
or OR4 (N3110, N3106, N128, N1552, N1490);
nor NOR2 (N3111, N3102, N1050);
and AND3 (N3112, N3105, N565, N783);
nand NAND4 (N3113, N3098, N1765, N860, N1992);
nand NAND3 (N3114, N3103, N2550, N746);
buf BUF1 (N3115, N3111);
nand NAND2 (N3116, N3110, N1181);
or OR3 (N3117, N3113, N45, N234);
and AND4 (N3118, N3112, N741, N1253, N1651);
xor XOR2 (N3119, N3115, N1250);
xor XOR2 (N3120, N3109, N2066);
buf BUF1 (N3121, N3120);
nor NOR2 (N3122, N3118, N1219);
and AND3 (N3123, N3116, N2435, N795);
and AND2 (N3124, N3122, N102);
not NOT1 (N3125, N3124);
buf BUF1 (N3126, N3114);
and AND3 (N3127, N3117, N405, N3101);
xor XOR2 (N3128, N3127, N676);
nor NOR3 (N3129, N3125, N1157, N2927);
and AND4 (N3130, N3119, N2501, N2281, N295);
not NOT1 (N3131, N3126);
and AND3 (N3132, N3107, N3025, N1160);
not NOT1 (N3133, N3085);
xor XOR2 (N3134, N3133, N386);
nor NOR3 (N3135, N3129, N1246, N2904);
or OR4 (N3136, N3134, N1857, N895, N1693);
not NOT1 (N3137, N3130);
nand NAND2 (N3138, N3137, N2);
nand NAND2 (N3139, N3131, N1775);
nand NAND2 (N3140, N3139, N404);
or OR2 (N3141, N3095, N1205);
and AND3 (N3142, N3141, N2913, N2394);
not NOT1 (N3143, N3138);
nor NOR3 (N3144, N3140, N2518, N1763);
buf BUF1 (N3145, N3123);
nor NOR4 (N3146, N3072, N1939, N1356, N505);
xor XOR2 (N3147, N3128, N1259);
nand NAND3 (N3148, N3145, N1015, N2169);
not NOT1 (N3149, N3135);
nand NAND4 (N3150, N3121, N3075, N113, N124);
not NOT1 (N3151, N3142);
xor XOR2 (N3152, N3132, N3137);
or OR3 (N3153, N3144, N460, N1125);
not NOT1 (N3154, N3148);
xor XOR2 (N3155, N3136, N1659);
nor NOR4 (N3156, N3150, N1317, N2087, N904);
and AND3 (N3157, N3147, N21, N2316);
buf BUF1 (N3158, N3151);
nor NOR2 (N3159, N3152, N481);
not NOT1 (N3160, N3149);
and AND4 (N3161, N3157, N1693, N2163, N468);
or OR4 (N3162, N3155, N2930, N2961, N2463);
buf BUF1 (N3163, N3156);
nor NOR3 (N3164, N3153, N840, N2334);
buf BUF1 (N3165, N3164);
nand NAND4 (N3166, N3143, N2678, N480, N163);
not NOT1 (N3167, N3158);
buf BUF1 (N3168, N3146);
and AND2 (N3169, N3168, N1058);
buf BUF1 (N3170, N3162);
xor XOR2 (N3171, N3165, N2025);
nand NAND2 (N3172, N3163, N3137);
nand NAND3 (N3173, N3167, N1667, N2495);
nand NAND3 (N3174, N3171, N686, N2984);
nand NAND3 (N3175, N3169, N1253, N2771);
and AND2 (N3176, N3170, N2006);
buf BUF1 (N3177, N3160);
buf BUF1 (N3178, N3174);
not NOT1 (N3179, N3178);
not NOT1 (N3180, N3166);
and AND3 (N3181, N3161, N172, N775);
buf BUF1 (N3182, N3181);
xor XOR2 (N3183, N3159, N1632);
nand NAND2 (N3184, N3177, N1089);
not NOT1 (N3185, N3180);
nor NOR4 (N3186, N3179, N121, N1389, N3076);
buf BUF1 (N3187, N3173);
nand NAND3 (N3188, N3185, N722, N2795);
nand NAND2 (N3189, N3175, N1825);
buf BUF1 (N3190, N3188);
xor XOR2 (N3191, N3189, N759);
xor XOR2 (N3192, N3172, N358);
xor XOR2 (N3193, N3190, N1544);
and AND3 (N3194, N3176, N236, N1454);
and AND2 (N3195, N3193, N418);
or OR4 (N3196, N3194, N331, N2880, N649);
buf BUF1 (N3197, N3187);
buf BUF1 (N3198, N3184);
nand NAND2 (N3199, N3186, N1336);
nor NOR3 (N3200, N3192, N1072, N1040);
xor XOR2 (N3201, N3197, N2333);
or OR3 (N3202, N3201, N1651, N1602);
xor XOR2 (N3203, N3195, N1990);
not NOT1 (N3204, N3196);
xor XOR2 (N3205, N3154, N615);
nor NOR4 (N3206, N3202, N384, N2391, N145);
nor NOR4 (N3207, N3183, N53, N1083, N58);
buf BUF1 (N3208, N3207);
not NOT1 (N3209, N3205);
not NOT1 (N3210, N3191);
nand NAND3 (N3211, N3206, N2414, N3127);
buf BUF1 (N3212, N3200);
or OR2 (N3213, N3210, N1511);
or OR4 (N3214, N3209, N3157, N647, N836);
buf BUF1 (N3215, N3208);
or OR2 (N3216, N3213, N1899);
nor NOR4 (N3217, N3211, N509, N2002, N897);
and AND4 (N3218, N3215, N2598, N2210, N1177);
xor XOR2 (N3219, N3218, N2945);
nand NAND2 (N3220, N3199, N2497);
not NOT1 (N3221, N3217);
buf BUF1 (N3222, N3182);
not NOT1 (N3223, N3212);
buf BUF1 (N3224, N3219);
nor NOR4 (N3225, N3198, N1572, N2727, N2056);
nor NOR2 (N3226, N3204, N731);
not NOT1 (N3227, N3220);
xor XOR2 (N3228, N3227, N533);
nor NOR3 (N3229, N3222, N388, N1471);
nand NAND2 (N3230, N3228, N965);
nor NOR3 (N3231, N3224, N678, N471);
nor NOR2 (N3232, N3225, N916);
buf BUF1 (N3233, N3229);
and AND2 (N3234, N3216, N2447);
or OR4 (N3235, N3221, N1533, N2741, N1928);
and AND3 (N3236, N3235, N625, N3101);
not NOT1 (N3237, N3203);
not NOT1 (N3238, N3226);
nor NOR2 (N3239, N3231, N1431);
not NOT1 (N3240, N3230);
buf BUF1 (N3241, N3234);
nor NOR2 (N3242, N3239, N1350);
not NOT1 (N3243, N3223);
buf BUF1 (N3244, N3233);
and AND4 (N3245, N3241, N639, N708, N2428);
or OR4 (N3246, N3238, N2655, N263, N2527);
or OR3 (N3247, N3242, N1507, N2917);
buf BUF1 (N3248, N3236);
xor XOR2 (N3249, N3248, N1372);
not NOT1 (N3250, N3247);
xor XOR2 (N3251, N3243, N2275);
nor NOR4 (N3252, N3245, N1112, N2444, N1804);
and AND2 (N3253, N3249, N3128);
buf BUF1 (N3254, N3251);
nor NOR3 (N3255, N3253, N1068, N1327);
and AND4 (N3256, N3250, N1158, N2940, N351);
buf BUF1 (N3257, N3255);
xor XOR2 (N3258, N3237, N2828);
and AND2 (N3259, N3246, N271);
not NOT1 (N3260, N3256);
buf BUF1 (N3261, N3257);
or OR4 (N3262, N3232, N962, N1586, N2562);
not NOT1 (N3263, N3262);
nor NOR4 (N3264, N3258, N406, N2716, N1996);
or OR4 (N3265, N3244, N268, N109, N2862);
not NOT1 (N3266, N3254);
nor NOR3 (N3267, N3266, N596, N2185);
not NOT1 (N3268, N3263);
not NOT1 (N3269, N3259);
buf BUF1 (N3270, N3265);
nand NAND3 (N3271, N3264, N1385, N1746);
not NOT1 (N3272, N3271);
or OR2 (N3273, N3261, N2095);
nor NOR2 (N3274, N3240, N63);
buf BUF1 (N3275, N3268);
and AND4 (N3276, N3269, N786, N453, N2887);
buf BUF1 (N3277, N3272);
and AND2 (N3278, N3260, N539);
and AND4 (N3279, N3267, N1423, N2786, N208);
xor XOR2 (N3280, N3214, N2608);
or OR3 (N3281, N3270, N2405, N699);
and AND4 (N3282, N3279, N2668, N2400, N3130);
xor XOR2 (N3283, N3252, N1339);
or OR4 (N3284, N3283, N1290, N1563, N2434);
or OR2 (N3285, N3276, N2218);
or OR2 (N3286, N3277, N2961);
buf BUF1 (N3287, N3281);
or OR2 (N3288, N3275, N2759);
nand NAND3 (N3289, N3287, N2415, N890);
nor NOR2 (N3290, N3282, N2592);
xor XOR2 (N3291, N3289, N2922);
and AND2 (N3292, N3285, N1789);
and AND3 (N3293, N3292, N1713, N56);
or OR2 (N3294, N3278, N682);
nor NOR4 (N3295, N3274, N1215, N3112, N241);
not NOT1 (N3296, N3280);
buf BUF1 (N3297, N3273);
and AND3 (N3298, N3286, N1722, N3034);
not NOT1 (N3299, N3290);
nand NAND2 (N3300, N3293, N3174);
buf BUF1 (N3301, N3296);
or OR4 (N3302, N3294, N2025, N3218, N2967);
or OR2 (N3303, N3300, N2618);
not NOT1 (N3304, N3299);
nand NAND3 (N3305, N3291, N199, N2572);
nor NOR2 (N3306, N3288, N1184);
nand NAND3 (N3307, N3303, N1140, N2165);
and AND2 (N3308, N3307, N726);
nor NOR2 (N3309, N3295, N674);
not NOT1 (N3310, N3306);
or OR4 (N3311, N3284, N1016, N1483, N853);
nand NAND4 (N3312, N3301, N217, N501, N3097);
not NOT1 (N3313, N3311);
nor NOR4 (N3314, N3310, N3311, N2219, N105);
nand NAND4 (N3315, N3302, N1197, N1740, N2777);
xor XOR2 (N3316, N3308, N2805);
not NOT1 (N3317, N3309);
nor NOR4 (N3318, N3314, N1526, N2034, N1367);
xor XOR2 (N3319, N3304, N291);
and AND2 (N3320, N3305, N1043);
nor NOR3 (N3321, N3318, N1232, N404);
xor XOR2 (N3322, N3298, N66);
not NOT1 (N3323, N3297);
nand NAND4 (N3324, N3320, N8, N2857, N419);
buf BUF1 (N3325, N3323);
nand NAND2 (N3326, N3321, N2618);
buf BUF1 (N3327, N3322);
or OR3 (N3328, N3327, N501, N2214);
nand NAND4 (N3329, N3312, N2226, N1358, N3180);
buf BUF1 (N3330, N3317);
and AND2 (N3331, N3319, N1209);
or OR4 (N3332, N3325, N781, N3206, N2286);
not NOT1 (N3333, N3331);
nor NOR2 (N3334, N3316, N2746);
nor NOR3 (N3335, N3313, N1971, N2046);
nand NAND3 (N3336, N3330, N1580, N1167);
not NOT1 (N3337, N3333);
and AND4 (N3338, N3315, N808, N1026, N2185);
or OR4 (N3339, N3324, N1927, N2476, N3050);
xor XOR2 (N3340, N3335, N2277);
xor XOR2 (N3341, N3326, N2627);
not NOT1 (N3342, N3329);
or OR3 (N3343, N3338, N1306, N1271);
xor XOR2 (N3344, N3343, N3055);
not NOT1 (N3345, N3336);
buf BUF1 (N3346, N3340);
and AND4 (N3347, N3337, N281, N375, N76);
xor XOR2 (N3348, N3347, N1535);
buf BUF1 (N3349, N3348);
buf BUF1 (N3350, N3345);
not NOT1 (N3351, N3350);
buf BUF1 (N3352, N3351);
nor NOR2 (N3353, N3341, N975);
nand NAND3 (N3354, N3352, N468, N79);
not NOT1 (N3355, N3332);
nor NOR3 (N3356, N3342, N1903, N2068);
or OR2 (N3357, N3344, N471);
and AND4 (N3358, N3356, N2150, N165, N2939);
or OR4 (N3359, N3354, N869, N2596, N176);
not NOT1 (N3360, N3328);
buf BUF1 (N3361, N3349);
not NOT1 (N3362, N3357);
nand NAND3 (N3363, N3359, N2130, N1444);
xor XOR2 (N3364, N3334, N1618);
nand NAND2 (N3365, N3358, N861);
nand NAND4 (N3366, N3363, N1633, N3074, N188);
nand NAND3 (N3367, N3355, N2316, N2800);
buf BUF1 (N3368, N3367);
xor XOR2 (N3369, N3368, N2843);
nand NAND3 (N3370, N3366, N3237, N682);
or OR3 (N3371, N3361, N986, N2874);
or OR4 (N3372, N3364, N409, N86, N1926);
xor XOR2 (N3373, N3369, N428);
xor XOR2 (N3374, N3373, N501);
nand NAND2 (N3375, N3371, N346);
nand NAND2 (N3376, N3375, N1936);
xor XOR2 (N3377, N3346, N2327);
nor NOR3 (N3378, N3377, N106, N1191);
buf BUF1 (N3379, N3376);
nor NOR2 (N3380, N3353, N1290);
nand NAND3 (N3381, N3378, N2962, N1983);
nor NOR3 (N3382, N3374, N211, N2313);
nor NOR2 (N3383, N3360, N269);
xor XOR2 (N3384, N3365, N1512);
and AND4 (N3385, N3383, N1865, N2428, N113);
nand NAND4 (N3386, N3380, N2322, N1238, N3195);
buf BUF1 (N3387, N3381);
not NOT1 (N3388, N3384);
and AND4 (N3389, N3382, N2399, N1709, N807);
not NOT1 (N3390, N3389);
xor XOR2 (N3391, N3388, N621);
nor NOR4 (N3392, N3362, N2461, N2856, N3300);
not NOT1 (N3393, N3392);
nor NOR2 (N3394, N3372, N2463);
nand NAND4 (N3395, N3386, N1391, N793, N2939);
xor XOR2 (N3396, N3379, N961);
or OR2 (N3397, N3339, N662);
nand NAND2 (N3398, N3387, N784);
nand NAND4 (N3399, N3385, N2667, N1781, N334);
xor XOR2 (N3400, N3390, N2227);
nand NAND2 (N3401, N3370, N2694);
not NOT1 (N3402, N3401);
not NOT1 (N3403, N3393);
buf BUF1 (N3404, N3394);
and AND2 (N3405, N3404, N2836);
buf BUF1 (N3406, N3402);
or OR4 (N3407, N3400, N2274, N2720, N1741);
or OR2 (N3408, N3397, N1636);
or OR3 (N3409, N3403, N3254, N3195);
or OR4 (N3410, N3409, N1981, N1707, N2388);
not NOT1 (N3411, N3405);
nand NAND2 (N3412, N3396, N2529);
or OR2 (N3413, N3410, N2184);
nor NOR3 (N3414, N3408, N542, N1519);
buf BUF1 (N3415, N3406);
buf BUF1 (N3416, N3395);
and AND4 (N3417, N3399, N986, N3103, N3193);
not NOT1 (N3418, N3411);
or OR4 (N3419, N3412, N441, N603, N2628);
buf BUF1 (N3420, N3418);
or OR4 (N3421, N3398, N1160, N1637, N1279);
not NOT1 (N3422, N3413);
or OR2 (N3423, N3419, N1049);
buf BUF1 (N3424, N3414);
buf BUF1 (N3425, N3424);
not NOT1 (N3426, N3423);
and AND4 (N3427, N3391, N163, N3160, N1056);
nor NOR4 (N3428, N3421, N3073, N1959, N1131);
and AND2 (N3429, N3426, N2104);
and AND2 (N3430, N3429, N2002);
or OR4 (N3431, N3430, N2545, N1746, N88);
buf BUF1 (N3432, N3416);
xor XOR2 (N3433, N3417, N171);
buf BUF1 (N3434, N3432);
nand NAND2 (N3435, N3422, N177);
buf BUF1 (N3436, N3427);
and AND4 (N3437, N3415, N2755, N2317, N2733);
not NOT1 (N3438, N3435);
buf BUF1 (N3439, N3428);
xor XOR2 (N3440, N3437, N2316);
nand NAND3 (N3441, N3434, N977, N598);
nor NOR3 (N3442, N3407, N3430, N740);
or OR3 (N3443, N3440, N2067, N2907);
not NOT1 (N3444, N3425);
xor XOR2 (N3445, N3436, N2949);
and AND3 (N3446, N3441, N600, N109);
nand NAND3 (N3447, N3445, N1356, N2866);
and AND3 (N3448, N3433, N2641, N1764);
or OR3 (N3449, N3448, N1420, N2302);
not NOT1 (N3450, N3447);
not NOT1 (N3451, N3431);
nand NAND2 (N3452, N3443, N669);
nand NAND2 (N3453, N3451, N3318);
nand NAND3 (N3454, N3453, N1474, N330);
buf BUF1 (N3455, N3449);
nand NAND2 (N3456, N3446, N2078);
buf BUF1 (N3457, N3455);
xor XOR2 (N3458, N3454, N306);
or OR4 (N3459, N3458, N1651, N2265, N585);
nor NOR3 (N3460, N3438, N3297, N1668);
and AND4 (N3461, N3452, N361, N2381, N80);
nand NAND4 (N3462, N3457, N2086, N354, N343);
not NOT1 (N3463, N3450);
nor NOR2 (N3464, N3444, N1890);
nor NOR2 (N3465, N3439, N2066);
nand NAND2 (N3466, N3464, N1079);
xor XOR2 (N3467, N3459, N3366);
nor NOR3 (N3468, N3461, N2971, N2763);
buf BUF1 (N3469, N3420);
nor NOR4 (N3470, N3460, N2454, N699, N3160);
or OR4 (N3471, N3467, N2038, N128, N965);
buf BUF1 (N3472, N3465);
xor XOR2 (N3473, N3468, N1619);
xor XOR2 (N3474, N3469, N1023);
nor NOR3 (N3475, N3474, N1101, N789);
nand NAND3 (N3476, N3442, N778, N2320);
or OR2 (N3477, N3466, N2381);
nand NAND4 (N3478, N3472, N931, N689, N1367);
xor XOR2 (N3479, N3456, N1077);
or OR3 (N3480, N3463, N2887, N2377);
not NOT1 (N3481, N3476);
or OR4 (N3482, N3462, N1592, N2745, N3446);
not NOT1 (N3483, N3477);
nor NOR2 (N3484, N3471, N2232);
or OR2 (N3485, N3484, N1997);
not NOT1 (N3486, N3481);
nor NOR3 (N3487, N3485, N920, N2919);
nor NOR3 (N3488, N3479, N1959, N444);
or OR4 (N3489, N3478, N1464, N2652, N1356);
not NOT1 (N3490, N3487);
buf BUF1 (N3491, N3490);
buf BUF1 (N3492, N3475);
nor NOR2 (N3493, N3482, N1407);
or OR4 (N3494, N3491, N1286, N1332, N1709);
not NOT1 (N3495, N3473);
buf BUF1 (N3496, N3494);
buf BUF1 (N3497, N3489);
and AND2 (N3498, N3493, N568);
and AND3 (N3499, N3480, N2163, N2935);
or OR2 (N3500, N3497, N3339);
or OR4 (N3501, N3483, N417, N1185, N1390);
buf BUF1 (N3502, N3501);
buf BUF1 (N3503, N3488);
buf BUF1 (N3504, N3496);
and AND2 (N3505, N3498, N2804);
and AND2 (N3506, N3504, N3375);
or OR3 (N3507, N3486, N2366, N2468);
nor NOR2 (N3508, N3492, N1842);
xor XOR2 (N3509, N3495, N2053);
nor NOR4 (N3510, N3503, N1274, N3034, N2807);
nand NAND2 (N3511, N3508, N2335);
xor XOR2 (N3512, N3502, N2381);
not NOT1 (N3513, N3507);
nand NAND3 (N3514, N3506, N2087, N592);
and AND2 (N3515, N3499, N2776);
or OR3 (N3516, N3512, N69, N3358);
xor XOR2 (N3517, N3516, N3432);
nand NAND2 (N3518, N3513, N887);
or OR4 (N3519, N3515, N567, N1087, N2126);
or OR2 (N3520, N3500, N275);
buf BUF1 (N3521, N3511);
or OR4 (N3522, N3510, N159, N2730, N485);
nand NAND4 (N3523, N3518, N776, N1420, N1355);
nand NAND4 (N3524, N3517, N682, N2530, N311);
xor XOR2 (N3525, N3524, N1193);
nand NAND4 (N3526, N3525, N1153, N1434, N227);
nand NAND2 (N3527, N3521, N2057);
xor XOR2 (N3528, N3527, N2953);
not NOT1 (N3529, N3505);
and AND2 (N3530, N3529, N1682);
xor XOR2 (N3531, N3528, N3007);
and AND3 (N3532, N3522, N1942, N1863);
buf BUF1 (N3533, N3514);
or OR2 (N3534, N3530, N1163);
xor XOR2 (N3535, N3519, N797);
and AND4 (N3536, N3535, N299, N3094, N1994);
not NOT1 (N3537, N3520);
nand NAND2 (N3538, N3534, N650);
nand NAND3 (N3539, N3536, N1435, N172);
nor NOR3 (N3540, N3532, N658, N2766);
not NOT1 (N3541, N3533);
and AND2 (N3542, N3470, N2953);
or OR2 (N3543, N3542, N3251);
and AND4 (N3544, N3526, N446, N2599, N3365);
xor XOR2 (N3545, N3543, N573);
or OR3 (N3546, N3538, N1561, N1879);
nor NOR4 (N3547, N3537, N3069, N2076, N3463);
or OR4 (N3548, N3509, N2228, N1584, N3061);
buf BUF1 (N3549, N3539);
not NOT1 (N3550, N3531);
and AND3 (N3551, N3544, N699, N1167);
not NOT1 (N3552, N3548);
or OR4 (N3553, N3523, N724, N2612, N533);
buf BUF1 (N3554, N3547);
not NOT1 (N3555, N3549);
nand NAND4 (N3556, N3540, N1270, N1763, N2222);
or OR3 (N3557, N3546, N2521, N1025);
and AND3 (N3558, N3551, N3439, N969);
nor NOR4 (N3559, N3541, N1493, N3262, N968);
or OR2 (N3560, N3552, N101);
and AND4 (N3561, N3560, N2217, N3198, N2418);
xor XOR2 (N3562, N3557, N2097);
and AND4 (N3563, N3556, N2636, N100, N1969);
nor NOR3 (N3564, N3563, N1475, N2417);
nor NOR4 (N3565, N3554, N2526, N404, N3311);
buf BUF1 (N3566, N3545);
and AND4 (N3567, N3558, N877, N2223, N138);
nand NAND4 (N3568, N3550, N3341, N939, N1415);
not NOT1 (N3569, N3561);
or OR3 (N3570, N3555, N1317, N3458);
and AND3 (N3571, N3569, N772, N2858);
and AND3 (N3572, N3562, N526, N2630);
or OR3 (N3573, N3568, N3327, N3106);
not NOT1 (N3574, N3570);
buf BUF1 (N3575, N3572);
buf BUF1 (N3576, N3565);
not NOT1 (N3577, N3564);
buf BUF1 (N3578, N3559);
nand NAND2 (N3579, N3553, N352);
and AND3 (N3580, N3578, N459, N3243);
xor XOR2 (N3581, N3567, N3387);
or OR2 (N3582, N3579, N154);
nand NAND2 (N3583, N3577, N2842);
buf BUF1 (N3584, N3571);
not NOT1 (N3585, N3580);
not NOT1 (N3586, N3574);
nor NOR3 (N3587, N3576, N1292, N1267);
and AND4 (N3588, N3585, N349, N2497, N2826);
buf BUF1 (N3589, N3575);
not NOT1 (N3590, N3583);
nand NAND2 (N3591, N3587, N2631);
nor NOR4 (N3592, N3586, N663, N2202, N1893);
or OR4 (N3593, N3590, N1429, N1297, N3187);
nor NOR2 (N3594, N3566, N108);
nor NOR4 (N3595, N3589, N1686, N1124, N1737);
xor XOR2 (N3596, N3595, N2244);
buf BUF1 (N3597, N3581);
buf BUF1 (N3598, N3596);
buf BUF1 (N3599, N3582);
nand NAND3 (N3600, N3592, N971, N3226);
and AND3 (N3601, N3597, N1041, N2623);
or OR4 (N3602, N3573, N2651, N1054, N560);
or OR3 (N3603, N3599, N2606, N2041);
nor NOR3 (N3604, N3584, N1285, N2518);
and AND4 (N3605, N3588, N2801, N3199, N1812);
not NOT1 (N3606, N3605);
xor XOR2 (N3607, N3598, N2424);
nor NOR2 (N3608, N3602, N2982);
nor NOR2 (N3609, N3600, N2096);
not NOT1 (N3610, N3609);
and AND4 (N3611, N3591, N923, N3569, N1181);
nand NAND4 (N3612, N3601, N2563, N165, N1152);
xor XOR2 (N3613, N3608, N2454);
or OR3 (N3614, N3594, N1958, N160);
nor NOR2 (N3615, N3613, N1886);
nand NAND4 (N3616, N3615, N3182, N24, N505);
or OR2 (N3617, N3607, N1582);
nand NAND4 (N3618, N3606, N1891, N2028, N3262);
xor XOR2 (N3619, N3618, N1964);
and AND2 (N3620, N3610, N2717);
nor NOR3 (N3621, N3593, N2180, N988);
buf BUF1 (N3622, N3620);
not NOT1 (N3623, N3619);
not NOT1 (N3624, N3611);
and AND3 (N3625, N3604, N508, N3435);
buf BUF1 (N3626, N3617);
xor XOR2 (N3627, N3626, N3272);
or OR3 (N3628, N3603, N1572, N1567);
nor NOR3 (N3629, N3622, N130, N604);
nand NAND3 (N3630, N3627, N1229, N596);
nand NAND3 (N3631, N3625, N1005, N2639);
or OR4 (N3632, N3614, N3300, N1876, N1103);
buf BUF1 (N3633, N3612);
nor NOR3 (N3634, N3623, N2479, N3181);
buf BUF1 (N3635, N3628);
and AND4 (N3636, N3632, N1792, N1643, N3486);
not NOT1 (N3637, N3633);
nand NAND2 (N3638, N3634, N1652);
and AND4 (N3639, N3636, N1545, N1043, N3210);
nand NAND3 (N3640, N3621, N2945, N995);
xor XOR2 (N3641, N3640, N2626);
nor NOR4 (N3642, N3630, N515, N1329, N117);
or OR4 (N3643, N3641, N2115, N1738, N1967);
and AND3 (N3644, N3642, N970, N2955);
nand NAND4 (N3645, N3624, N1801, N3291, N2663);
buf BUF1 (N3646, N3629);
nor NOR4 (N3647, N3646, N382, N686, N59);
buf BUF1 (N3648, N3616);
nor NOR3 (N3649, N3638, N885, N1210);
nand NAND3 (N3650, N3647, N3247, N2361);
not NOT1 (N3651, N3644);
nor NOR4 (N3652, N3649, N2247, N1594, N527);
not NOT1 (N3653, N3648);
xor XOR2 (N3654, N3653, N2590);
buf BUF1 (N3655, N3654);
or OR3 (N3656, N3637, N1180, N341);
and AND3 (N3657, N3643, N934, N2105);
not NOT1 (N3658, N3655);
nand NAND4 (N3659, N3656, N2638, N1723, N1377);
nand NAND2 (N3660, N3635, N501);
or OR2 (N3661, N3657, N531);
or OR4 (N3662, N3659, N317, N799, N1876);
nand NAND4 (N3663, N3645, N3627, N1434, N3407);
or OR3 (N3664, N3651, N1948, N2612);
or OR3 (N3665, N3661, N1263, N2033);
buf BUF1 (N3666, N3650);
nand NAND4 (N3667, N3660, N1573, N3551, N2544);
or OR4 (N3668, N3667, N2648, N2675, N2690);
buf BUF1 (N3669, N3666);
and AND3 (N3670, N3664, N1543, N1679);
or OR3 (N3671, N3658, N924, N3051);
buf BUF1 (N3672, N3665);
and AND4 (N3673, N3631, N1897, N1100, N2830);
and AND4 (N3674, N3669, N476, N1210, N3373);
nand NAND2 (N3675, N3639, N214);
xor XOR2 (N3676, N3673, N2711);
or OR3 (N3677, N3662, N2892, N2706);
not NOT1 (N3678, N3652);
nand NAND4 (N3679, N3671, N718, N2170, N1554);
and AND2 (N3680, N3679, N3538);
xor XOR2 (N3681, N3680, N182);
nor NOR4 (N3682, N3678, N2588, N945, N3307);
buf BUF1 (N3683, N3672);
not NOT1 (N3684, N3682);
xor XOR2 (N3685, N3674, N252);
nor NOR2 (N3686, N3685, N2728);
nor NOR2 (N3687, N3677, N1444);
nand NAND3 (N3688, N3676, N940, N2547);
nor NOR4 (N3689, N3684, N3613, N2827, N334);
xor XOR2 (N3690, N3687, N2628);
nor NOR2 (N3691, N3675, N3552);
xor XOR2 (N3692, N3686, N790);
nor NOR3 (N3693, N3690, N2438, N957);
xor XOR2 (N3694, N3688, N1267);
or OR2 (N3695, N3668, N463);
buf BUF1 (N3696, N3683);
or OR4 (N3697, N3696, N1641, N2037, N3528);
buf BUF1 (N3698, N3693);
xor XOR2 (N3699, N3670, N1348);
xor XOR2 (N3700, N3694, N1922);
xor XOR2 (N3701, N3698, N1321);
nand NAND4 (N3702, N3689, N1485, N2052, N3071);
and AND4 (N3703, N3695, N24, N3614, N3446);
nand NAND3 (N3704, N3681, N1407, N3410);
or OR4 (N3705, N3692, N3305, N2921, N582);
buf BUF1 (N3706, N3702);
buf BUF1 (N3707, N3699);
or OR3 (N3708, N3701, N3685, N717);
not NOT1 (N3709, N3707);
nand NAND3 (N3710, N3708, N2894, N1572);
xor XOR2 (N3711, N3709, N2721);
nor NOR3 (N3712, N3705, N1556, N307);
nand NAND2 (N3713, N3706, N2821);
or OR2 (N3714, N3704, N562);
not NOT1 (N3715, N3714);
nor NOR2 (N3716, N3700, N1854);
not NOT1 (N3717, N3697);
and AND3 (N3718, N3710, N499, N428);
or OR4 (N3719, N3691, N671, N601, N994);
buf BUF1 (N3720, N3718);
nor NOR2 (N3721, N3715, N429);
not NOT1 (N3722, N3703);
and AND3 (N3723, N3722, N263, N355);
and AND2 (N3724, N3720, N710);
nor NOR3 (N3725, N3719, N775, N3264);
not NOT1 (N3726, N3713);
buf BUF1 (N3727, N3711);
or OR3 (N3728, N3727, N2533, N335);
nor NOR4 (N3729, N3725, N2634, N155, N1560);
or OR2 (N3730, N3712, N623);
or OR4 (N3731, N3729, N1097, N792, N794);
nor NOR4 (N3732, N3717, N860, N1918, N3390);
nand NAND3 (N3733, N3724, N791, N1879);
and AND2 (N3734, N3726, N1555);
nand NAND4 (N3735, N3734, N3093, N3574, N794);
xor XOR2 (N3736, N3663, N2881);
xor XOR2 (N3737, N3735, N2909);
and AND3 (N3738, N3736, N3454, N331);
and AND3 (N3739, N3716, N3190, N865);
and AND3 (N3740, N3738, N1431, N1980);
and AND2 (N3741, N3733, N917);
not NOT1 (N3742, N3721);
not NOT1 (N3743, N3737);
buf BUF1 (N3744, N3743);
not NOT1 (N3745, N3744);
nand NAND3 (N3746, N3742, N145, N1424);
or OR2 (N3747, N3739, N2564);
buf BUF1 (N3748, N3745);
nor NOR3 (N3749, N3731, N787, N1790);
nand NAND2 (N3750, N3730, N1939);
nor NOR3 (N3751, N3748, N582, N1924);
nor NOR2 (N3752, N3741, N3671);
nand NAND2 (N3753, N3750, N2896);
nor NOR3 (N3754, N3747, N75, N1293);
xor XOR2 (N3755, N3754, N2865);
nand NAND3 (N3756, N3732, N1867, N1879);
or OR4 (N3757, N3755, N1071, N2877, N3577);
nand NAND4 (N3758, N3751, N2897, N3077, N896);
and AND3 (N3759, N3758, N852, N2247);
buf BUF1 (N3760, N3753);
or OR3 (N3761, N3759, N1018, N1123);
nand NAND4 (N3762, N3761, N2031, N1444, N2847);
nand NAND4 (N3763, N3723, N3583, N2967, N569);
buf BUF1 (N3764, N3749);
or OR2 (N3765, N3760, N269);
or OR2 (N3766, N3765, N894);
nor NOR2 (N3767, N3756, N2751);
nand NAND2 (N3768, N3762, N3595);
not NOT1 (N3769, N3763);
nand NAND2 (N3770, N3767, N65);
nor NOR3 (N3771, N3740, N2756, N107);
nand NAND4 (N3772, N3768, N2055, N1304, N934);
buf BUF1 (N3773, N3771);
nand NAND2 (N3774, N3728, N1472);
not NOT1 (N3775, N3757);
not NOT1 (N3776, N3752);
or OR2 (N3777, N3773, N2745);
not NOT1 (N3778, N3746);
xor XOR2 (N3779, N3778, N2666);
not NOT1 (N3780, N3775);
not NOT1 (N3781, N3770);
and AND3 (N3782, N3779, N3453, N1237);
or OR3 (N3783, N3781, N1098, N136);
buf BUF1 (N3784, N3782);
or OR4 (N3785, N3772, N3089, N1648, N1623);
buf BUF1 (N3786, N3766);
xor XOR2 (N3787, N3774, N1761);
nor NOR4 (N3788, N3786, N3047, N958, N173);
buf BUF1 (N3789, N3764);
xor XOR2 (N3790, N3788, N1055);
nand NAND4 (N3791, N3783, N2900, N147, N3168);
and AND2 (N3792, N3769, N2288);
buf BUF1 (N3793, N3776);
nand NAND4 (N3794, N3784, N473, N651, N2989);
or OR2 (N3795, N3789, N1305);
and AND3 (N3796, N3785, N1932, N917);
and AND3 (N3797, N3787, N528, N1346);
buf BUF1 (N3798, N3791);
xor XOR2 (N3799, N3790, N3444);
buf BUF1 (N3800, N3795);
buf BUF1 (N3801, N3798);
xor XOR2 (N3802, N3780, N2769);
or OR4 (N3803, N3796, N327, N1650, N173);
nand NAND2 (N3804, N3801, N3114);
not NOT1 (N3805, N3800);
not NOT1 (N3806, N3793);
or OR4 (N3807, N3806, N149, N3095, N3262);
nand NAND4 (N3808, N3792, N419, N186, N52);
not NOT1 (N3809, N3803);
or OR3 (N3810, N3802, N679, N1166);
and AND4 (N3811, N3777, N538, N2893, N352);
buf BUF1 (N3812, N3809);
xor XOR2 (N3813, N3811, N714);
xor XOR2 (N3814, N3799, N2365);
xor XOR2 (N3815, N3805, N2292);
buf BUF1 (N3816, N3810);
and AND3 (N3817, N3812, N2867, N3566);
not NOT1 (N3818, N3814);
and AND2 (N3819, N3807, N3459);
nand NAND4 (N3820, N3794, N2572, N2073, N1879);
nand NAND2 (N3821, N3820, N1846);
buf BUF1 (N3822, N3813);
nand NAND3 (N3823, N3797, N1669, N2039);
and AND4 (N3824, N3822, N1744, N3263, N506);
xor XOR2 (N3825, N3816, N3438);
buf BUF1 (N3826, N3817);
nor NOR3 (N3827, N3804, N3224, N541);
buf BUF1 (N3828, N3819);
or OR3 (N3829, N3824, N1190, N194);
xor XOR2 (N3830, N3815, N510);
nand NAND3 (N3831, N3823, N1823, N1896);
nand NAND3 (N3832, N3830, N3207, N224);
nand NAND4 (N3833, N3827, N1886, N915, N1468);
nor NOR4 (N3834, N3826, N3350, N471, N3825);
or OR2 (N3835, N1707, N2517);
not NOT1 (N3836, N3828);
buf BUF1 (N3837, N3808);
and AND4 (N3838, N3829, N3152, N2357, N2204);
and AND2 (N3839, N3818, N1106);
not NOT1 (N3840, N3838);
nor NOR3 (N3841, N3834, N3689, N548);
or OR2 (N3842, N3821, N1529);
buf BUF1 (N3843, N3831);
buf BUF1 (N3844, N3842);
xor XOR2 (N3845, N3840, N977);
or OR3 (N3846, N3836, N980, N1456);
nor NOR3 (N3847, N3835, N1515, N3806);
xor XOR2 (N3848, N3845, N1367);
and AND4 (N3849, N3843, N556, N2175, N2838);
nand NAND4 (N3850, N3848, N3757, N650, N3278);
nor NOR4 (N3851, N3846, N1791, N2733, N3780);
buf BUF1 (N3852, N3841);
and AND3 (N3853, N3839, N712, N3824);
xor XOR2 (N3854, N3853, N3347);
and AND3 (N3855, N3850, N1767, N1561);
or OR4 (N3856, N3854, N3595, N1765, N1654);
not NOT1 (N3857, N3851);
or OR4 (N3858, N3849, N2251, N3313, N316);
not NOT1 (N3859, N3856);
or OR3 (N3860, N3832, N2290, N1280);
buf BUF1 (N3861, N3855);
not NOT1 (N3862, N3837);
nor NOR4 (N3863, N3858, N3345, N3428, N1541);
not NOT1 (N3864, N3847);
buf BUF1 (N3865, N3852);
buf BUF1 (N3866, N3863);
and AND3 (N3867, N3857, N1880, N551);
or OR2 (N3868, N3859, N748);
or OR4 (N3869, N3860, N2053, N970, N2127);
or OR4 (N3870, N3868, N3763, N2512, N1571);
nor NOR4 (N3871, N3862, N207, N943, N528);
xor XOR2 (N3872, N3869, N2340);
xor XOR2 (N3873, N3866, N1895);
not NOT1 (N3874, N3833);
or OR4 (N3875, N3864, N3253, N1156, N1270);
nor NOR2 (N3876, N3867, N2249);
nand NAND3 (N3877, N3876, N2108, N1392);
and AND4 (N3878, N3874, N3397, N128, N1144);
buf BUF1 (N3879, N3878);
or OR3 (N3880, N3875, N3335, N1804);
buf BUF1 (N3881, N3872);
not NOT1 (N3882, N3870);
or OR2 (N3883, N3881, N2114);
buf BUF1 (N3884, N3871);
buf BUF1 (N3885, N3873);
and AND2 (N3886, N3861, N2224);
nor NOR2 (N3887, N3886, N2550);
buf BUF1 (N3888, N3865);
or OR2 (N3889, N3885, N170);
not NOT1 (N3890, N3883);
xor XOR2 (N3891, N3882, N2048);
and AND4 (N3892, N3877, N19, N1629, N3152);
not NOT1 (N3893, N3889);
not NOT1 (N3894, N3879);
and AND2 (N3895, N3888, N3004);
xor XOR2 (N3896, N3880, N3808);
nor NOR2 (N3897, N3891, N449);
and AND3 (N3898, N3894, N1305, N2578);
and AND4 (N3899, N3898, N1039, N1910, N1129);
or OR4 (N3900, N3896, N2917, N3721, N2220);
buf BUF1 (N3901, N3899);
buf BUF1 (N3902, N3897);
nand NAND4 (N3903, N3893, N3287, N956, N707);
or OR4 (N3904, N3902, N1022, N1145, N676);
nor NOR4 (N3905, N3887, N3009, N2692, N728);
or OR3 (N3906, N3901, N2735, N661);
and AND4 (N3907, N3900, N2298, N1094, N1824);
buf BUF1 (N3908, N3844);
buf BUF1 (N3909, N3905);
nand NAND2 (N3910, N3908, N3021);
xor XOR2 (N3911, N3909, N223);
nand NAND4 (N3912, N3884, N1751, N2994, N1370);
or OR2 (N3913, N3906, N3802);
not NOT1 (N3914, N3904);
or OR3 (N3915, N3890, N3274, N2235);
xor XOR2 (N3916, N3912, N3481);
nor NOR3 (N3917, N3914, N1660, N994);
nand NAND2 (N3918, N3903, N3862);
nand NAND3 (N3919, N3895, N3761, N2044);
nor NOR4 (N3920, N3917, N2614, N987, N881);
nor NOR3 (N3921, N3919, N2013, N891);
buf BUF1 (N3922, N3921);
xor XOR2 (N3923, N3892, N2203);
not NOT1 (N3924, N3910);
not NOT1 (N3925, N3924);
not NOT1 (N3926, N3913);
xor XOR2 (N3927, N3918, N1101);
or OR3 (N3928, N3925, N2704, N76);
or OR4 (N3929, N3926, N2560, N3883, N1368);
or OR4 (N3930, N3907, N1634, N1814, N182);
buf BUF1 (N3931, N3929);
and AND3 (N3932, N3930, N2187, N3378);
buf BUF1 (N3933, N3916);
and AND2 (N3934, N3911, N2193);
not NOT1 (N3935, N3933);
and AND3 (N3936, N3935, N1927, N2923);
xor XOR2 (N3937, N3915, N3821);
xor XOR2 (N3938, N3923, N241);
nor NOR2 (N3939, N3928, N3075);
xor XOR2 (N3940, N3927, N3632);
nand NAND2 (N3941, N3934, N436);
nand NAND4 (N3942, N3941, N3031, N1409, N3538);
xor XOR2 (N3943, N3932, N1260);
xor XOR2 (N3944, N3937, N1589);
and AND4 (N3945, N3944, N1841, N1476, N1792);
or OR4 (N3946, N3938, N532, N3325, N1450);
buf BUF1 (N3947, N3946);
and AND3 (N3948, N3939, N1268, N2353);
or OR4 (N3949, N3945, N2219, N2684, N747);
xor XOR2 (N3950, N3947, N3092);
not NOT1 (N3951, N3920);
or OR2 (N3952, N3950, N2221);
and AND3 (N3953, N3931, N2238, N441);
nand NAND2 (N3954, N3922, N2746);
and AND3 (N3955, N3943, N140, N2762);
and AND2 (N3956, N3951, N1875);
xor XOR2 (N3957, N3949, N888);
and AND2 (N3958, N3948, N3700);
buf BUF1 (N3959, N3955);
not NOT1 (N3960, N3958);
not NOT1 (N3961, N3953);
or OR3 (N3962, N3936, N2382, N1665);
nand NAND2 (N3963, N3959, N1588);
not NOT1 (N3964, N3961);
nor NOR4 (N3965, N3957, N2446, N533, N3060);
buf BUF1 (N3966, N3942);
nand NAND3 (N3967, N3962, N621, N1572);
buf BUF1 (N3968, N3963);
not NOT1 (N3969, N3967);
not NOT1 (N3970, N3968);
and AND2 (N3971, N3940, N2054);
or OR2 (N3972, N3966, N640);
not NOT1 (N3973, N3965);
or OR3 (N3974, N3969, N1106, N1080);
nor NOR3 (N3975, N3964, N3422, N3379);
buf BUF1 (N3976, N3973);
or OR3 (N3977, N3974, N2192, N3639);
and AND3 (N3978, N3975, N3518, N3311);
not NOT1 (N3979, N3954);
or OR4 (N3980, N3978, N878, N3870, N1390);
and AND3 (N3981, N3970, N3831, N650);
not NOT1 (N3982, N3971);
or OR2 (N3983, N3982, N2751);
or OR4 (N3984, N3977, N1978, N2085, N1537);
buf BUF1 (N3985, N3956);
not NOT1 (N3986, N3960);
and AND2 (N3987, N3983, N3308);
xor XOR2 (N3988, N3985, N953);
nand NAND4 (N3989, N3980, N747, N2508, N2967);
buf BUF1 (N3990, N3972);
xor XOR2 (N3991, N3984, N1135);
buf BUF1 (N3992, N3989);
not NOT1 (N3993, N3988);
xor XOR2 (N3994, N3991, N2403);
nand NAND2 (N3995, N3979, N3000);
xor XOR2 (N3996, N3990, N332);
or OR4 (N3997, N3996, N2600, N2670, N2153);
nand NAND4 (N3998, N3976, N2104, N2517, N2095);
and AND3 (N3999, N3952, N3934, N3626);
buf BUF1 (N4000, N3997);
or OR4 (N4001, N3999, N1707, N2285, N3820);
not NOT1 (N4002, N3998);
nor NOR3 (N4003, N4000, N1323, N2418);
not NOT1 (N4004, N3994);
nor NOR4 (N4005, N4002, N89, N76, N943);
buf BUF1 (N4006, N4001);
buf BUF1 (N4007, N3981);
nand NAND2 (N4008, N4007, N3280);
nand NAND3 (N4009, N4008, N326, N2844);
xor XOR2 (N4010, N3986, N651);
not NOT1 (N4011, N4005);
nand NAND2 (N4012, N4011, N3991);
xor XOR2 (N4013, N3993, N2177);
not NOT1 (N4014, N4003);
not NOT1 (N4015, N4014);
xor XOR2 (N4016, N4006, N1324);
and AND4 (N4017, N4004, N2022, N1830, N926);
buf BUF1 (N4018, N4017);
nor NOR3 (N4019, N3987, N1533, N4016);
xor XOR2 (N4020, N1732, N800);
and AND2 (N4021, N4012, N3497);
buf BUF1 (N4022, N4013);
buf BUF1 (N4023, N4021);
nor NOR3 (N4024, N4009, N2933, N592);
not NOT1 (N4025, N4015);
buf BUF1 (N4026, N4023);
or OR2 (N4027, N4018, N3427);
buf BUF1 (N4028, N4010);
and AND3 (N4029, N4024, N2873, N74);
or OR2 (N4030, N4026, N3828);
buf BUF1 (N4031, N4019);
nor NOR2 (N4032, N4020, N808);
not NOT1 (N4033, N4027);
nor NOR2 (N4034, N4030, N1190);
or OR3 (N4035, N4025, N3455, N1195);
buf BUF1 (N4036, N4028);
xor XOR2 (N4037, N4022, N3382);
and AND3 (N4038, N4036, N430, N955);
buf BUF1 (N4039, N4035);
nor NOR2 (N4040, N4034, N112);
buf BUF1 (N4041, N4037);
not NOT1 (N4042, N4041);
xor XOR2 (N4043, N4029, N2056);
xor XOR2 (N4044, N4032, N3944);
nand NAND4 (N4045, N4043, N3667, N37, N372);
nor NOR3 (N4046, N4044, N518, N511);
and AND3 (N4047, N4031, N3741, N2297);
and AND4 (N4048, N4033, N2749, N4020, N165);
xor XOR2 (N4049, N4045, N2793);
nand NAND2 (N4050, N4040, N3631);
or OR2 (N4051, N4042, N3618);
nand NAND2 (N4052, N3995, N4004);
and AND3 (N4053, N4046, N1151, N338);
not NOT1 (N4054, N4050);
xor XOR2 (N4055, N4038, N1107);
nand NAND3 (N4056, N4052, N2011, N950);
xor XOR2 (N4057, N4055, N3381);
not NOT1 (N4058, N4053);
buf BUF1 (N4059, N4048);
buf BUF1 (N4060, N4058);
xor XOR2 (N4061, N4039, N3319);
not NOT1 (N4062, N4061);
and AND2 (N4063, N4054, N874);
nor NOR3 (N4064, N3992, N1493, N3206);
nand NAND3 (N4065, N4062, N1410, N201);
buf BUF1 (N4066, N4049);
and AND4 (N4067, N4057, N3687, N2862, N2873);
and AND3 (N4068, N4060, N2843, N883);
not NOT1 (N4069, N4066);
nand NAND2 (N4070, N4065, N2836);
and AND4 (N4071, N4070, N1452, N3693, N3744);
or OR4 (N4072, N4064, N1778, N1704, N981);
or OR4 (N4073, N4072, N103, N313, N2063);
and AND2 (N4074, N4063, N2036);
not NOT1 (N4075, N4067);
nor NOR3 (N4076, N4074, N133, N1992);
buf BUF1 (N4077, N4069);
and AND3 (N4078, N4059, N3233, N3433);
buf BUF1 (N4079, N4077);
xor XOR2 (N4080, N4047, N3594);
xor XOR2 (N4081, N4078, N3084);
and AND2 (N4082, N4081, N559);
and AND2 (N4083, N4068, N3870);
and AND4 (N4084, N4071, N1250, N2145, N506);
buf BUF1 (N4085, N4082);
xor XOR2 (N4086, N4076, N2238);
xor XOR2 (N4087, N4085, N215);
xor XOR2 (N4088, N4080, N1675);
xor XOR2 (N4089, N4079, N1633);
not NOT1 (N4090, N4089);
nand NAND3 (N4091, N4073, N1181, N103);
or OR4 (N4092, N4090, N2972, N1296, N4008);
or OR2 (N4093, N4051, N772);
buf BUF1 (N4094, N4092);
nand NAND4 (N4095, N4088, N2794, N1106, N3153);
buf BUF1 (N4096, N4056);
xor XOR2 (N4097, N4087, N1028);
nand NAND4 (N4098, N4097, N2038, N1099, N3512);
nor NOR2 (N4099, N4093, N2073);
nor NOR3 (N4100, N4098, N3253, N3402);
xor XOR2 (N4101, N4094, N3095);
nand NAND2 (N4102, N4075, N354);
nor NOR4 (N4103, N4086, N2819, N3907, N843);
and AND4 (N4104, N4101, N1328, N1740, N2136);
not NOT1 (N4105, N4103);
xor XOR2 (N4106, N4095, N16);
or OR2 (N4107, N4100, N3916);
and AND2 (N4108, N4083, N1155);
nand NAND2 (N4109, N4096, N760);
nor NOR4 (N4110, N4104, N2648, N3210, N515);
nand NAND3 (N4111, N4105, N3841, N3132);
nor NOR3 (N4112, N4108, N3021, N3269);
or OR2 (N4113, N4091, N761);
not NOT1 (N4114, N4107);
nor NOR3 (N4115, N4112, N3680, N2959);
nor NOR2 (N4116, N4102, N3030);
nand NAND3 (N4117, N4110, N1412, N437);
not NOT1 (N4118, N4084);
and AND2 (N4119, N4109, N1970);
not NOT1 (N4120, N4111);
and AND4 (N4121, N4118, N626, N4044, N3945);
not NOT1 (N4122, N4106);
nor NOR3 (N4123, N4120, N3077, N1209);
buf BUF1 (N4124, N4116);
or OR2 (N4125, N4115, N3554);
xor XOR2 (N4126, N4125, N776);
xor XOR2 (N4127, N4113, N5);
buf BUF1 (N4128, N4117);
not NOT1 (N4129, N4122);
nand NAND2 (N4130, N4114, N3301);
and AND2 (N4131, N4130, N1558);
nor NOR3 (N4132, N4121, N2360, N3752);
or OR4 (N4133, N4127, N880, N3531, N339);
nand NAND4 (N4134, N4099, N1497, N2128, N715);
or OR4 (N4135, N4124, N1870, N4037, N3717);
and AND2 (N4136, N4134, N3254);
and AND4 (N4137, N4136, N3992, N1345, N3046);
buf BUF1 (N4138, N4132);
nand NAND4 (N4139, N4126, N1055, N581, N2921);
nand NAND4 (N4140, N4133, N1084, N822, N2392);
not NOT1 (N4141, N4137);
buf BUF1 (N4142, N4138);
buf BUF1 (N4143, N4131);
and AND4 (N4144, N4119, N1288, N3353, N2939);
xor XOR2 (N4145, N4143, N1231);
buf BUF1 (N4146, N4141);
buf BUF1 (N4147, N4128);
buf BUF1 (N4148, N4147);
not NOT1 (N4149, N4129);
buf BUF1 (N4150, N4139);
buf BUF1 (N4151, N4150);
buf BUF1 (N4152, N4149);
nor NOR4 (N4153, N4123, N1158, N3509, N693);
buf BUF1 (N4154, N4146);
nor NOR4 (N4155, N4145, N3772, N1976, N193);
buf BUF1 (N4156, N4153);
not NOT1 (N4157, N4144);
not NOT1 (N4158, N4155);
not NOT1 (N4159, N4152);
nand NAND3 (N4160, N4151, N1841, N3093);
or OR2 (N4161, N4158, N247);
and AND3 (N4162, N4159, N1195, N1880);
or OR2 (N4163, N4161, N2329);
nand NAND3 (N4164, N4135, N1444, N3738);
nand NAND4 (N4165, N4162, N3481, N56, N1047);
not NOT1 (N4166, N4142);
and AND3 (N4167, N4165, N954, N359);
not NOT1 (N4168, N4160);
xor XOR2 (N4169, N4167, N1336);
nand NAND2 (N4170, N4168, N2385);
nor NOR3 (N4171, N4140, N2814, N3203);
not NOT1 (N4172, N4164);
xor XOR2 (N4173, N4163, N452);
not NOT1 (N4174, N4169);
nand NAND2 (N4175, N4173, N378);
nand NAND3 (N4176, N4175, N2075, N3815);
buf BUF1 (N4177, N4176);
nor NOR3 (N4178, N4174, N2707, N604);
or OR4 (N4179, N4156, N1349, N827, N845);
buf BUF1 (N4180, N4177);
buf BUF1 (N4181, N4148);
nand NAND4 (N4182, N4181, N4049, N2948, N609);
and AND3 (N4183, N4180, N3377, N3462);
nor NOR2 (N4184, N4154, N1853);
or OR4 (N4185, N4157, N1228, N1786, N3179);
buf BUF1 (N4186, N4184);
xor XOR2 (N4187, N4179, N244);
nand NAND4 (N4188, N4171, N493, N1199, N3571);
nor NOR3 (N4189, N4178, N2077, N3934);
nand NAND2 (N4190, N4189, N4006);
not NOT1 (N4191, N4166);
and AND3 (N4192, N4172, N2279, N3099);
and AND2 (N4193, N4190, N3802);
nand NAND2 (N4194, N4186, N2165);
not NOT1 (N4195, N4170);
nor NOR4 (N4196, N4193, N1766, N2135, N1543);
buf BUF1 (N4197, N4187);
buf BUF1 (N4198, N4197);
or OR2 (N4199, N4194, N284);
not NOT1 (N4200, N4188);
xor XOR2 (N4201, N4191, N42);
nor NOR2 (N4202, N4199, N3747);
nor NOR3 (N4203, N4200, N2993, N2704);
buf BUF1 (N4204, N4201);
buf BUF1 (N4205, N4195);
nand NAND2 (N4206, N4204, N3522);
or OR2 (N4207, N4205, N1382);
buf BUF1 (N4208, N4203);
and AND4 (N4209, N4183, N305, N2919, N2);
nand NAND2 (N4210, N4206, N3879);
not NOT1 (N4211, N4198);
xor XOR2 (N4212, N4211, N3404);
or OR4 (N4213, N4210, N2180, N751, N721);
nor NOR3 (N4214, N4185, N1717, N2266);
xor XOR2 (N4215, N4214, N4178);
nor NOR3 (N4216, N4212, N1319, N2281);
not NOT1 (N4217, N4215);
or OR3 (N4218, N4216, N1805, N1547);
xor XOR2 (N4219, N4196, N1749);
xor XOR2 (N4220, N4213, N2069);
xor XOR2 (N4221, N4217, N311);
or OR3 (N4222, N4220, N2943, N2214);
buf BUF1 (N4223, N4222);
and AND3 (N4224, N4209, N3188, N88);
and AND3 (N4225, N4192, N2816, N1806);
xor XOR2 (N4226, N4223, N223);
not NOT1 (N4227, N4202);
not NOT1 (N4228, N4225);
nand NAND3 (N4229, N4221, N2120, N1166);
buf BUF1 (N4230, N4208);
nand NAND4 (N4231, N4207, N3233, N4053, N122);
nor NOR2 (N4232, N4219, N2496);
or OR4 (N4233, N4228, N3849, N316, N3855);
and AND4 (N4234, N4229, N2045, N1849, N3286);
and AND2 (N4235, N4182, N1952);
nand NAND4 (N4236, N4233, N3779, N2436, N1145);
and AND3 (N4237, N4231, N2169, N2463);
xor XOR2 (N4238, N4237, N2713);
nor NOR2 (N4239, N4227, N3073);
buf BUF1 (N4240, N4234);
xor XOR2 (N4241, N4226, N166);
not NOT1 (N4242, N4240);
and AND3 (N4243, N4224, N289, N708);
buf BUF1 (N4244, N4241);
nor NOR2 (N4245, N4242, N2414);
xor XOR2 (N4246, N4230, N2385);
or OR3 (N4247, N4238, N2143, N3754);
or OR3 (N4248, N4218, N292, N2965);
or OR4 (N4249, N4239, N673, N1023, N2782);
and AND2 (N4250, N4247, N4019);
not NOT1 (N4251, N4245);
nand NAND3 (N4252, N4244, N705, N4013);
buf BUF1 (N4253, N4248);
nand NAND2 (N4254, N4252, N4163);
buf BUF1 (N4255, N4243);
and AND4 (N4256, N4253, N1649, N1266, N924);
xor XOR2 (N4257, N4236, N409);
nand NAND4 (N4258, N4257, N3922, N692, N1696);
xor XOR2 (N4259, N4255, N61);
buf BUF1 (N4260, N4254);
not NOT1 (N4261, N4256);
not NOT1 (N4262, N4246);
and AND2 (N4263, N4249, N3865);
and AND4 (N4264, N4263, N3343, N1206, N2777);
xor XOR2 (N4265, N4258, N2101);
or OR2 (N4266, N4262, N3954);
and AND4 (N4267, N4261, N3763, N1564, N4167);
nand NAND4 (N4268, N4266, N2906, N2506, N82);
and AND3 (N4269, N4260, N45, N3741);
buf BUF1 (N4270, N4264);
not NOT1 (N4271, N4235);
nand NAND2 (N4272, N4259, N3943);
not NOT1 (N4273, N4270);
or OR2 (N4274, N4269, N2737);
or OR2 (N4275, N4274, N2248);
nor NOR3 (N4276, N4251, N3053, N703);
and AND2 (N4277, N4232, N452);
xor XOR2 (N4278, N4275, N2787);
and AND2 (N4279, N4271, N3964);
or OR2 (N4280, N4250, N1122);
buf BUF1 (N4281, N4267);
nor NOR4 (N4282, N4276, N3072, N1681, N2547);
xor XOR2 (N4283, N4277, N4187);
buf BUF1 (N4284, N4272);
and AND2 (N4285, N4279, N3413);
buf BUF1 (N4286, N4265);
or OR2 (N4287, N4283, N47);
nor NOR4 (N4288, N4278, N2092, N2542, N3399);
nand NAND4 (N4289, N4286, N1129, N4144, N865);
and AND2 (N4290, N4268, N1658);
and AND2 (N4291, N4280, N2526);
xor XOR2 (N4292, N4290, N3190);
or OR3 (N4293, N4287, N827, N918);
or OR2 (N4294, N4281, N2401);
xor XOR2 (N4295, N4291, N1634);
or OR3 (N4296, N4285, N3679, N3403);
buf BUF1 (N4297, N4284);
not NOT1 (N4298, N4295);
xor XOR2 (N4299, N4296, N2409);
and AND2 (N4300, N4292, N3363);
buf BUF1 (N4301, N4299);
xor XOR2 (N4302, N4282, N565);
or OR3 (N4303, N4273, N335, N2537);
and AND2 (N4304, N4288, N2474);
not NOT1 (N4305, N4293);
nor NOR2 (N4306, N4302, N2849);
nor NOR3 (N4307, N4300, N2851, N2850);
or OR2 (N4308, N4289, N1886);
and AND4 (N4309, N4297, N3493, N1568, N4230);
xor XOR2 (N4310, N4309, N3698);
xor XOR2 (N4311, N4304, N1333);
and AND2 (N4312, N4294, N457);
nand NAND4 (N4313, N4305, N176, N2213, N3377);
buf BUF1 (N4314, N4303);
xor XOR2 (N4315, N4308, N71);
nand NAND4 (N4316, N4301, N3920, N2779, N1249);
not NOT1 (N4317, N4306);
nand NAND2 (N4318, N4317, N1419);
nor NOR3 (N4319, N4318, N1220, N1687);
not NOT1 (N4320, N4316);
and AND2 (N4321, N4313, N581);
buf BUF1 (N4322, N4321);
or OR3 (N4323, N4312, N2065, N4029);
and AND3 (N4324, N4310, N958, N2394);
or OR2 (N4325, N4320, N2941);
buf BUF1 (N4326, N4314);
buf BUF1 (N4327, N4323);
buf BUF1 (N4328, N4326);
or OR3 (N4329, N4328, N3803, N1874);
nor NOR2 (N4330, N4329, N1828);
nor NOR2 (N4331, N4307, N1250);
buf BUF1 (N4332, N4322);
nand NAND4 (N4333, N4332, N1328, N3040, N3042);
nand NAND2 (N4334, N4327, N4063);
nand NAND4 (N4335, N4330, N2711, N3459, N1856);
not NOT1 (N4336, N4319);
nor NOR3 (N4337, N4324, N2515, N1484);
buf BUF1 (N4338, N4337);
buf BUF1 (N4339, N4334);
buf BUF1 (N4340, N4311);
nor NOR3 (N4341, N4336, N4269, N3528);
nor NOR4 (N4342, N4333, N809, N1233, N782);
and AND2 (N4343, N4325, N1090);
buf BUF1 (N4344, N4338);
not NOT1 (N4345, N4343);
or OR3 (N4346, N4339, N939, N1144);
not NOT1 (N4347, N4344);
not NOT1 (N4348, N4345);
buf BUF1 (N4349, N4335);
buf BUF1 (N4350, N4342);
or OR3 (N4351, N4340, N3447, N111);
xor XOR2 (N4352, N4350, N3558);
xor XOR2 (N4353, N4331, N3768);
xor XOR2 (N4354, N4347, N1538);
or OR2 (N4355, N4351, N2191);
nor NOR3 (N4356, N4346, N779, N2248);
nand NAND2 (N4357, N4341, N134);
buf BUF1 (N4358, N4357);
and AND4 (N4359, N4315, N3873, N2246, N4276);
nor NOR4 (N4360, N4354, N4139, N493, N729);
nor NOR2 (N4361, N4298, N3644);
xor XOR2 (N4362, N4355, N3483);
not NOT1 (N4363, N4358);
nand NAND2 (N4364, N4356, N3227);
or OR2 (N4365, N4359, N1439);
nor NOR4 (N4366, N4348, N2454, N1346, N733);
or OR4 (N4367, N4349, N3033, N3587, N2154);
buf BUF1 (N4368, N4363);
buf BUF1 (N4369, N4352);
nand NAND2 (N4370, N4361, N2559);
not NOT1 (N4371, N4362);
or OR4 (N4372, N4353, N966, N1233, N4069);
buf BUF1 (N4373, N4370);
buf BUF1 (N4374, N4366);
or OR4 (N4375, N4374, N139, N2112, N1610);
nand NAND3 (N4376, N4372, N3619, N1575);
xor XOR2 (N4377, N4368, N874);
not NOT1 (N4378, N4377);
buf BUF1 (N4379, N4376);
not NOT1 (N4380, N4379);
nand NAND4 (N4381, N4380, N1115, N2964, N1580);
nand NAND2 (N4382, N4371, N129);
xor XOR2 (N4383, N4381, N2033);
xor XOR2 (N4384, N4360, N3508);
nand NAND3 (N4385, N4365, N3433, N1533);
buf BUF1 (N4386, N4378);
nand NAND4 (N4387, N4385, N1113, N1990, N2343);
nor NOR4 (N4388, N4384, N2740, N368, N3633);
buf BUF1 (N4389, N4383);
nor NOR3 (N4390, N4369, N1112, N1451);
and AND2 (N4391, N4375, N1208);
not NOT1 (N4392, N4373);
and AND4 (N4393, N4387, N4152, N3056, N1363);
or OR2 (N4394, N4390, N737);
nor NOR4 (N4395, N4393, N3322, N3877, N1414);
not NOT1 (N4396, N4394);
nand NAND2 (N4397, N4388, N2221);
nor NOR4 (N4398, N4396, N1553, N952, N1454);
buf BUF1 (N4399, N4386);
buf BUF1 (N4400, N4364);
not NOT1 (N4401, N4400);
nand NAND4 (N4402, N4367, N3585, N2606, N3050);
not NOT1 (N4403, N4397);
or OR3 (N4404, N4382, N2190, N2118);
xor XOR2 (N4405, N4395, N2471);
buf BUF1 (N4406, N4399);
xor XOR2 (N4407, N4405, N4380);
and AND2 (N4408, N4392, N3333);
nor NOR2 (N4409, N4406, N3411);
and AND4 (N4410, N4402, N3537, N466, N3964);
nand NAND2 (N4411, N4409, N1098);
and AND3 (N4412, N4403, N2301, N1126);
not NOT1 (N4413, N4401);
buf BUF1 (N4414, N4389);
buf BUF1 (N4415, N4398);
buf BUF1 (N4416, N4407);
and AND4 (N4417, N4414, N1235, N8, N3269);
xor XOR2 (N4418, N4410, N2917);
or OR3 (N4419, N4416, N272, N2717);
or OR4 (N4420, N4419, N2277, N86, N1594);
not NOT1 (N4421, N4417);
or OR4 (N4422, N4412, N3158, N3775, N2786);
buf BUF1 (N4423, N4411);
nand NAND4 (N4424, N4418, N1266, N2607, N400);
buf BUF1 (N4425, N4415);
nand NAND4 (N4426, N4423, N163, N2414, N4318);
and AND4 (N4427, N4426, N3892, N4078, N234);
xor XOR2 (N4428, N4420, N1314);
or OR4 (N4429, N4427, N1629, N1544, N4018);
and AND3 (N4430, N4413, N1812, N4303);
or OR3 (N4431, N4422, N771, N1892);
xor XOR2 (N4432, N4428, N3274);
or OR3 (N4433, N4431, N1659, N3122);
nand NAND4 (N4434, N4424, N3131, N3106, N3517);
buf BUF1 (N4435, N4425);
buf BUF1 (N4436, N4408);
not NOT1 (N4437, N4433);
nand NAND2 (N4438, N4434, N3536);
buf BUF1 (N4439, N4432);
nor NOR4 (N4440, N4439, N10, N2305, N3554);
buf BUF1 (N4441, N4440);
buf BUF1 (N4442, N4430);
xor XOR2 (N4443, N4429, N71);
xor XOR2 (N4444, N4438, N3988);
or OR4 (N4445, N4444, N3070, N2204, N835);
xor XOR2 (N4446, N4421, N772);
buf BUF1 (N4447, N4443);
xor XOR2 (N4448, N4447, N4249);
not NOT1 (N4449, N4446);
not NOT1 (N4450, N4435);
xor XOR2 (N4451, N4391, N1022);
or OR4 (N4452, N4437, N4211, N1885, N3522);
and AND3 (N4453, N4450, N2037, N4225);
and AND2 (N4454, N4442, N1249);
or OR4 (N4455, N4445, N4062, N4000, N1039);
buf BUF1 (N4456, N4441);
xor XOR2 (N4457, N4452, N2296);
and AND2 (N4458, N4451, N4130);
buf BUF1 (N4459, N4455);
or OR4 (N4460, N4456, N30, N11, N468);
xor XOR2 (N4461, N4436, N999);
or OR2 (N4462, N4454, N1014);
xor XOR2 (N4463, N4448, N752);
xor XOR2 (N4464, N4449, N1920);
or OR4 (N4465, N4453, N973, N3763, N1874);
xor XOR2 (N4466, N4457, N4395);
buf BUF1 (N4467, N4465);
xor XOR2 (N4468, N4461, N402);
nand NAND2 (N4469, N4458, N2352);
nand NAND4 (N4470, N4404, N1947, N222, N3015);
and AND4 (N4471, N4459, N457, N3234, N2205);
and AND3 (N4472, N4470, N1820, N4053);
xor XOR2 (N4473, N4471, N3813);
nand NAND2 (N4474, N4472, N3422);
not NOT1 (N4475, N4466);
xor XOR2 (N4476, N4473, N2935);
not NOT1 (N4477, N4474);
xor XOR2 (N4478, N4476, N2896);
not NOT1 (N4479, N4462);
or OR2 (N4480, N4463, N3377);
nand NAND4 (N4481, N4469, N1733, N1325, N147);
not NOT1 (N4482, N4477);
xor XOR2 (N4483, N4468, N3458);
nand NAND4 (N4484, N4483, N1301, N319, N1605);
nand NAND4 (N4485, N4478, N164, N2735, N1197);
nand NAND2 (N4486, N4475, N4033);
not NOT1 (N4487, N4480);
buf BUF1 (N4488, N4487);
buf BUF1 (N4489, N4460);
or OR3 (N4490, N4482, N4188, N774);
xor XOR2 (N4491, N4485, N577);
xor XOR2 (N4492, N4464, N3107);
buf BUF1 (N4493, N4479);
or OR4 (N4494, N4493, N2046, N3188, N3734);
buf BUF1 (N4495, N4494);
not NOT1 (N4496, N4486);
nand NAND3 (N4497, N4491, N182, N62);
buf BUF1 (N4498, N4467);
or OR2 (N4499, N4488, N299);
nor NOR4 (N4500, N4497, N561, N3513, N1687);
buf BUF1 (N4501, N4495);
nor NOR4 (N4502, N4499, N2248, N1601, N2759);
not NOT1 (N4503, N4484);
not NOT1 (N4504, N4502);
nand NAND3 (N4505, N4498, N1462, N2390);
not NOT1 (N4506, N4500);
xor XOR2 (N4507, N4501, N3834);
nor NOR3 (N4508, N4489, N1924, N4087);
xor XOR2 (N4509, N4505, N3127);
nand NAND4 (N4510, N4509, N3959, N998, N1525);
or OR2 (N4511, N4481, N3502);
or OR4 (N4512, N4503, N3250, N3491, N3748);
and AND3 (N4513, N4504, N802, N3397);
xor XOR2 (N4514, N4492, N1161);
not NOT1 (N4515, N4508);
buf BUF1 (N4516, N4511);
and AND4 (N4517, N4513, N1492, N770, N4178);
or OR2 (N4518, N4517, N1194);
not NOT1 (N4519, N4518);
or OR4 (N4520, N4506, N2233, N3218, N1901);
xor XOR2 (N4521, N4514, N1269);
or OR2 (N4522, N4520, N1607);
buf BUF1 (N4523, N4516);
not NOT1 (N4524, N4519);
and AND3 (N4525, N4512, N3284, N2332);
buf BUF1 (N4526, N4524);
nand NAND2 (N4527, N4522, N1136);
or OR2 (N4528, N4496, N1823);
not NOT1 (N4529, N4521);
buf BUF1 (N4530, N4527);
or OR3 (N4531, N4528, N2522, N2324);
xor XOR2 (N4532, N4490, N1341);
not NOT1 (N4533, N4531);
and AND2 (N4534, N4529, N1234);
xor XOR2 (N4535, N4534, N2488);
and AND4 (N4536, N4526, N2121, N3510, N1410);
and AND4 (N4537, N4535, N285, N3008, N2831);
buf BUF1 (N4538, N4537);
buf BUF1 (N4539, N4536);
nor NOR4 (N4540, N4525, N2790, N2064, N3634);
not NOT1 (N4541, N4538);
buf BUF1 (N4542, N4530);
xor XOR2 (N4543, N4533, N42);
and AND3 (N4544, N4532, N1193, N4245);
or OR4 (N4545, N4515, N3726, N3364, N3255);
not NOT1 (N4546, N4542);
nand NAND4 (N4547, N4546, N3207, N1703, N3344);
xor XOR2 (N4548, N4545, N709);
xor XOR2 (N4549, N4547, N2485);
or OR4 (N4550, N4548, N1263, N2774, N2962);
and AND2 (N4551, N4510, N349);
or OR4 (N4552, N4540, N1200, N776, N905);
and AND3 (N4553, N4551, N3291, N1852);
and AND2 (N4554, N4553, N2961);
not NOT1 (N4555, N4554);
nor NOR3 (N4556, N4539, N2536, N2448);
or OR4 (N4557, N4556, N2355, N3643, N152);
nor NOR4 (N4558, N4552, N374, N4130, N1173);
not NOT1 (N4559, N4523);
xor XOR2 (N4560, N4543, N812);
and AND3 (N4561, N4557, N3474, N3075);
or OR3 (N4562, N4541, N3203, N3210);
and AND4 (N4563, N4544, N1093, N788, N1527);
or OR4 (N4564, N4560, N4294, N2296, N3292);
and AND3 (N4565, N4555, N958, N1204);
nor NOR2 (N4566, N4563, N4001);
buf BUF1 (N4567, N4549);
nor NOR2 (N4568, N4550, N3655);
not NOT1 (N4569, N4562);
not NOT1 (N4570, N4561);
or OR3 (N4571, N4567, N4115, N3782);
xor XOR2 (N4572, N4571, N1454);
xor XOR2 (N4573, N4570, N1907);
nor NOR2 (N4574, N4569, N1596);
xor XOR2 (N4575, N4565, N2377);
nand NAND3 (N4576, N4507, N3865, N2153);
or OR4 (N4577, N4576, N4267, N1629, N2257);
buf BUF1 (N4578, N4566);
or OR2 (N4579, N4575, N844);
nor NOR4 (N4580, N4574, N1662, N892, N4382);
xor XOR2 (N4581, N4572, N521);
and AND4 (N4582, N4580, N3516, N4477, N339);
or OR2 (N4583, N4578, N409);
xor XOR2 (N4584, N4582, N4339);
nand NAND4 (N4585, N4581, N2113, N861, N162);
buf BUF1 (N4586, N4583);
nor NOR4 (N4587, N4558, N3121, N1589, N3869);
buf BUF1 (N4588, N4568);
and AND4 (N4589, N4579, N3096, N2747, N864);
not NOT1 (N4590, N4564);
and AND4 (N4591, N4588, N2676, N2703, N921);
nand NAND3 (N4592, N4590, N1236, N2112);
nor NOR4 (N4593, N4592, N4292, N3293, N935);
buf BUF1 (N4594, N4587);
nor NOR4 (N4595, N4589, N916, N3346, N2425);
nand NAND2 (N4596, N4584, N4385);
not NOT1 (N4597, N4596);
xor XOR2 (N4598, N4594, N1428);
xor XOR2 (N4599, N4597, N843);
nor NOR4 (N4600, N4593, N1756, N220, N2317);
or OR3 (N4601, N4598, N67, N1181);
nor NOR3 (N4602, N4585, N1664, N1699);
buf BUF1 (N4603, N4601);
nand NAND2 (N4604, N4577, N2071);
and AND3 (N4605, N4586, N1190, N990);
and AND3 (N4606, N4600, N1266, N1530);
or OR3 (N4607, N4599, N3652, N2149);
and AND3 (N4608, N4607, N1956, N804);
xor XOR2 (N4609, N4605, N2340);
xor XOR2 (N4610, N4573, N3585);
nor NOR2 (N4611, N4591, N1969);
and AND3 (N4612, N4604, N135, N3087);
buf BUF1 (N4613, N4611);
nor NOR4 (N4614, N4602, N1715, N3315, N2884);
xor XOR2 (N4615, N4613, N577);
or OR2 (N4616, N4612, N1142);
or OR3 (N4617, N4609, N1323, N3293);
not NOT1 (N4618, N4559);
nor NOR2 (N4619, N4608, N3044);
nor NOR4 (N4620, N4615, N4475, N3229, N1182);
and AND2 (N4621, N4603, N2529);
not NOT1 (N4622, N4618);
and AND4 (N4623, N4595, N2619, N2646, N3978);
not NOT1 (N4624, N4620);
and AND3 (N4625, N4619, N2914, N409);
not NOT1 (N4626, N4621);
nand NAND4 (N4627, N4614, N1941, N474, N4168);
nand NAND4 (N4628, N4606, N1102, N435, N1331);
buf BUF1 (N4629, N4622);
or OR3 (N4630, N4623, N4573, N1275);
or OR3 (N4631, N4626, N4453, N4491);
xor XOR2 (N4632, N4630, N4143);
or OR2 (N4633, N4616, N900);
or OR4 (N4634, N4628, N3548, N212, N3394);
and AND2 (N4635, N4627, N2308);
buf BUF1 (N4636, N4624);
nand NAND3 (N4637, N4632, N4499, N3321);
xor XOR2 (N4638, N4631, N525);
and AND2 (N4639, N4634, N2517);
nand NAND2 (N4640, N4638, N4002);
and AND3 (N4641, N4625, N2190, N3784);
xor XOR2 (N4642, N4635, N904);
nand NAND4 (N4643, N4636, N4418, N917, N4170);
or OR3 (N4644, N4640, N4316, N866);
buf BUF1 (N4645, N4617);
nor NOR3 (N4646, N4643, N37, N1621);
nand NAND2 (N4647, N4645, N2400);
nand NAND4 (N4648, N4637, N2962, N4379, N1200);
nand NAND4 (N4649, N4647, N4231, N729, N437);
or OR2 (N4650, N4649, N1134);
and AND4 (N4651, N4644, N4473, N1740, N3341);
xor XOR2 (N4652, N4650, N2941);
buf BUF1 (N4653, N4652);
not NOT1 (N4654, N4642);
and AND3 (N4655, N4641, N4264, N2830);
nor NOR4 (N4656, N4610, N3268, N667, N2224);
or OR3 (N4657, N4629, N4048, N1642);
nand NAND4 (N4658, N4657, N3463, N495, N4201);
not NOT1 (N4659, N4633);
xor XOR2 (N4660, N4656, N4526);
buf BUF1 (N4661, N4660);
and AND3 (N4662, N4658, N2863, N2574);
nand NAND4 (N4663, N4653, N4073, N4646, N3366);
buf BUF1 (N4664, N3272);
nor NOR4 (N4665, N4639, N1266, N2650, N685);
xor XOR2 (N4666, N4663, N1251);
or OR4 (N4667, N4654, N300, N4536, N3772);
xor XOR2 (N4668, N4662, N2658);
or OR4 (N4669, N4668, N1371, N2650, N1927);
nand NAND4 (N4670, N4661, N4325, N2256, N3763);
nand NAND2 (N4671, N4655, N2057);
and AND3 (N4672, N4665, N609, N3188);
not NOT1 (N4673, N4672);
nor NOR3 (N4674, N4670, N704, N1243);
xor XOR2 (N4675, N4673, N2414);
buf BUF1 (N4676, N4674);
xor XOR2 (N4677, N4676, N2712);
buf BUF1 (N4678, N4671);
buf BUF1 (N4679, N4669);
buf BUF1 (N4680, N4659);
nor NOR2 (N4681, N4675, N704);
nor NOR3 (N4682, N4677, N4555, N929);
xor XOR2 (N4683, N4681, N4356);
and AND4 (N4684, N4682, N1179, N4334, N3284);
not NOT1 (N4685, N4679);
buf BUF1 (N4686, N4666);
nand NAND2 (N4687, N4680, N2620);
xor XOR2 (N4688, N4651, N3043);
nor NOR4 (N4689, N4667, N2266, N868, N4507);
or OR2 (N4690, N4683, N2145);
nand NAND2 (N4691, N4690, N1674);
nand NAND2 (N4692, N4687, N3980);
and AND4 (N4693, N4691, N709, N4440, N4121);
or OR4 (N4694, N4686, N4324, N515, N1908);
or OR2 (N4695, N4678, N4088);
or OR4 (N4696, N4689, N858, N4692, N4054);
nand NAND4 (N4697, N4399, N2834, N140, N4296);
nor NOR2 (N4698, N4697, N2375);
xor XOR2 (N4699, N4685, N4325);
and AND4 (N4700, N4696, N1553, N630, N86);
nand NAND2 (N4701, N4664, N4568);
not NOT1 (N4702, N4693);
not NOT1 (N4703, N4702);
xor XOR2 (N4704, N4648, N964);
nand NAND4 (N4705, N4698, N2343, N3862, N633);
nor NOR2 (N4706, N4700, N789);
not NOT1 (N4707, N4684);
xor XOR2 (N4708, N4699, N452);
nand NAND4 (N4709, N4701, N814, N2351, N1814);
nand NAND2 (N4710, N4688, N922);
xor XOR2 (N4711, N4708, N4527);
or OR2 (N4712, N4704, N2081);
buf BUF1 (N4713, N4694);
and AND3 (N4714, N4710, N2224, N4536);
and AND3 (N4715, N4709, N4396, N882);
nand NAND4 (N4716, N4705, N2619, N2501, N241);
and AND4 (N4717, N4703, N1557, N2349, N1463);
buf BUF1 (N4718, N4716);
or OR2 (N4719, N4714, N1773);
and AND2 (N4720, N4717, N3668);
or OR3 (N4721, N4715, N1640, N2512);
buf BUF1 (N4722, N4720);
buf BUF1 (N4723, N4712);
nand NAND2 (N4724, N4723, N4699);
not NOT1 (N4725, N4711);
xor XOR2 (N4726, N4706, N1804);
or OR2 (N4727, N4721, N2437);
xor XOR2 (N4728, N4707, N4459);
or OR2 (N4729, N4722, N2563);
not NOT1 (N4730, N4713);
nand NAND3 (N4731, N4729, N3839, N2747);
xor XOR2 (N4732, N4730, N1520);
or OR4 (N4733, N4726, N4538, N4481, N3827);
nand NAND4 (N4734, N4731, N4071, N2755, N1447);
xor XOR2 (N4735, N4695, N2906);
or OR4 (N4736, N4725, N2545, N3848, N2428);
or OR4 (N4737, N4736, N861, N1952, N3272);
not NOT1 (N4738, N4727);
and AND2 (N4739, N4724, N4010);
nor NOR4 (N4740, N4734, N1860, N4172, N4098);
not NOT1 (N4741, N4719);
xor XOR2 (N4742, N4738, N3656);
or OR3 (N4743, N4737, N3517, N2601);
nand NAND2 (N4744, N4742, N1380);
or OR2 (N4745, N4739, N2314);
or OR3 (N4746, N4740, N4036, N3312);
and AND4 (N4747, N4728, N3729, N1311, N1872);
nand NAND4 (N4748, N4746, N179, N2908, N4405);
xor XOR2 (N4749, N4733, N1698);
nor NOR2 (N4750, N4744, N560);
or OR4 (N4751, N4743, N3254, N3800, N3603);
xor XOR2 (N4752, N4745, N392);
and AND4 (N4753, N4748, N2081, N83, N1433);
nand NAND2 (N4754, N4752, N237);
buf BUF1 (N4755, N4732);
not NOT1 (N4756, N4750);
buf BUF1 (N4757, N4753);
or OR2 (N4758, N4757, N3588);
or OR4 (N4759, N4741, N1729, N2053, N2235);
and AND2 (N4760, N4759, N2258);
nand NAND2 (N4761, N4758, N3598);
nor NOR2 (N4762, N4751, N4426);
not NOT1 (N4763, N4760);
xor XOR2 (N4764, N4755, N2091);
nand NAND2 (N4765, N4763, N1635);
and AND4 (N4766, N4749, N4457, N1552, N3877);
not NOT1 (N4767, N4764);
not NOT1 (N4768, N4765);
not NOT1 (N4769, N4756);
or OR3 (N4770, N4762, N1669, N3315);
xor XOR2 (N4771, N4766, N2097);
not NOT1 (N4772, N4769);
buf BUF1 (N4773, N4747);
and AND3 (N4774, N4767, N1276, N2517);
nand NAND4 (N4775, N4772, N3526, N3432, N2858);
nor NOR3 (N4776, N4768, N4538, N3075);
buf BUF1 (N4777, N4774);
not NOT1 (N4778, N4754);
nor NOR4 (N4779, N4775, N588, N82, N1502);
buf BUF1 (N4780, N4718);
xor XOR2 (N4781, N4779, N2590);
buf BUF1 (N4782, N4780);
and AND2 (N4783, N4776, N945);
xor XOR2 (N4784, N4783, N4106);
and AND4 (N4785, N4782, N2192, N4039, N1883);
and AND4 (N4786, N4785, N4292, N1248, N4471);
not NOT1 (N4787, N4735);
xor XOR2 (N4788, N4777, N2965);
nor NOR2 (N4789, N4773, N2454);
xor XOR2 (N4790, N4771, N2494);
or OR3 (N4791, N4784, N1625, N2066);
nand NAND3 (N4792, N4786, N4219, N1649);
nand NAND2 (N4793, N4791, N3959);
xor XOR2 (N4794, N4793, N2372);
or OR2 (N4795, N4781, N332);
and AND3 (N4796, N4787, N1298, N500);
and AND3 (N4797, N4761, N5, N2619);
nand NAND2 (N4798, N4797, N1777);
nand NAND2 (N4799, N4798, N3884);
nand NAND4 (N4800, N4789, N3992, N2066, N4720);
buf BUF1 (N4801, N4796);
or OR4 (N4802, N4801, N1834, N197, N3494);
nor NOR2 (N4803, N4795, N3030);
or OR2 (N4804, N4794, N3019);
buf BUF1 (N4805, N4802);
buf BUF1 (N4806, N4800);
buf BUF1 (N4807, N4770);
not NOT1 (N4808, N4807);
not NOT1 (N4809, N4806);
nor NOR3 (N4810, N4809, N2372, N3113);
xor XOR2 (N4811, N4790, N611);
or OR2 (N4812, N4778, N1992);
and AND4 (N4813, N4792, N3794, N145, N3543);
not NOT1 (N4814, N4812);
nand NAND3 (N4815, N4799, N4427, N316);
nand NAND3 (N4816, N4810, N3270, N1419);
not NOT1 (N4817, N4788);
not NOT1 (N4818, N4808);
and AND4 (N4819, N4804, N2806, N4444, N1066);
and AND2 (N4820, N4815, N4573);
xor XOR2 (N4821, N4816, N3366);
nand NAND4 (N4822, N4818, N4067, N3221, N1153);
nand NAND4 (N4823, N4805, N2592, N1789, N1890);
or OR2 (N4824, N4817, N2729);
and AND4 (N4825, N4813, N3791, N106, N2945);
not NOT1 (N4826, N4824);
nor NOR3 (N4827, N4803, N1542, N326);
xor XOR2 (N4828, N4822, N1999);
or OR4 (N4829, N4826, N3264, N3738, N3100);
buf BUF1 (N4830, N4819);
not NOT1 (N4831, N4821);
xor XOR2 (N4832, N4825, N125);
xor XOR2 (N4833, N4830, N2289);
xor XOR2 (N4834, N4828, N2656);
buf BUF1 (N4835, N4814);
and AND3 (N4836, N4831, N2390, N1266);
or OR2 (N4837, N4833, N2980);
xor XOR2 (N4838, N4834, N677);
not NOT1 (N4839, N4829);
xor XOR2 (N4840, N4823, N4081);
or OR2 (N4841, N4832, N1977);
or OR2 (N4842, N4835, N580);
or OR3 (N4843, N4842, N3337, N840);
not NOT1 (N4844, N4827);
nand NAND3 (N4845, N4836, N99, N1493);
buf BUF1 (N4846, N4844);
nor NOR3 (N4847, N4845, N4604, N4191);
and AND4 (N4848, N4846, N3051, N3766, N2954);
buf BUF1 (N4849, N4840);
nor NOR3 (N4850, N4820, N2070, N565);
not NOT1 (N4851, N4838);
and AND2 (N4852, N4841, N1197);
nor NOR3 (N4853, N4839, N3433, N493);
or OR2 (N4854, N4851, N2156);
xor XOR2 (N4855, N4843, N4781);
xor XOR2 (N4856, N4847, N4700);
buf BUF1 (N4857, N4811);
not NOT1 (N4858, N4837);
and AND2 (N4859, N4855, N4726);
xor XOR2 (N4860, N4849, N2113);
not NOT1 (N4861, N4857);
buf BUF1 (N4862, N4853);
nor NOR3 (N4863, N4858, N4672, N4565);
or OR4 (N4864, N4859, N4691, N3432, N2786);
buf BUF1 (N4865, N4852);
and AND2 (N4866, N4850, N2882);
nor NOR4 (N4867, N4861, N679, N1683, N2989);
buf BUF1 (N4868, N4866);
and AND3 (N4869, N4856, N2665, N2277);
nand NAND4 (N4870, N4867, N2574, N101, N1247);
and AND2 (N4871, N4848, N1297);
not NOT1 (N4872, N4860);
and AND4 (N4873, N4862, N751, N2876, N709);
or OR2 (N4874, N4870, N3166);
or OR2 (N4875, N4864, N4395);
or OR3 (N4876, N4854, N1496, N2537);
nor NOR4 (N4877, N4863, N4341, N2183, N2950);
and AND4 (N4878, N4874, N3102, N916, N4048);
nor NOR4 (N4879, N4875, N3040, N3951, N2526);
nor NOR2 (N4880, N4877, N332);
not NOT1 (N4881, N4873);
buf BUF1 (N4882, N4872);
and AND4 (N4883, N4868, N2835, N3233, N489);
buf BUF1 (N4884, N4871);
not NOT1 (N4885, N4876);
or OR3 (N4886, N4869, N36, N3755);
not NOT1 (N4887, N4884);
or OR3 (N4888, N4885, N554, N2383);
xor XOR2 (N4889, N4880, N2487);
and AND4 (N4890, N4881, N2563, N2899, N3493);
nand NAND2 (N4891, N4883, N158);
and AND2 (N4892, N4886, N3918);
xor XOR2 (N4893, N4878, N4350);
nand NAND4 (N4894, N4887, N4048, N4345, N3178);
nand NAND4 (N4895, N4890, N3186, N1117, N3361);
or OR2 (N4896, N4892, N2290);
xor XOR2 (N4897, N4865, N4468);
xor XOR2 (N4898, N4895, N643);
nor NOR4 (N4899, N4889, N3016, N3199, N212);
xor XOR2 (N4900, N4882, N1095);
or OR3 (N4901, N4897, N4723, N4858);
nor NOR3 (N4902, N4888, N1073, N3887);
nand NAND2 (N4903, N4902, N452);
nand NAND4 (N4904, N4903, N3235, N1103, N3192);
xor XOR2 (N4905, N4896, N4742);
or OR3 (N4906, N4894, N872, N736);
nand NAND4 (N4907, N4893, N1060, N2232, N2039);
buf BUF1 (N4908, N4899);
nand NAND2 (N4909, N4898, N856);
nand NAND3 (N4910, N4907, N46, N4017);
not NOT1 (N4911, N4906);
or OR2 (N4912, N4904, N4503);
nand NAND4 (N4913, N4911, N203, N2768, N3500);
buf BUF1 (N4914, N4891);
nand NAND3 (N4915, N4909, N2243, N455);
not NOT1 (N4916, N4900);
xor XOR2 (N4917, N4914, N1444);
xor XOR2 (N4918, N4908, N4159);
xor XOR2 (N4919, N4905, N3514);
nand NAND2 (N4920, N4910, N1322);
buf BUF1 (N4921, N4916);
not NOT1 (N4922, N4913);
xor XOR2 (N4923, N4918, N1256);
xor XOR2 (N4924, N4912, N4025);
nor NOR2 (N4925, N4922, N1879);
or OR2 (N4926, N4921, N3049);
buf BUF1 (N4927, N4879);
xor XOR2 (N4928, N4901, N50);
xor XOR2 (N4929, N4919, N1833);
nand NAND2 (N4930, N4920, N1432);
buf BUF1 (N4931, N4930);
and AND2 (N4932, N4925, N4742);
nor NOR2 (N4933, N4928, N893);
buf BUF1 (N4934, N4929);
buf BUF1 (N4935, N4932);
xor XOR2 (N4936, N4923, N353);
and AND3 (N4937, N4934, N1531, N4405);
and AND3 (N4938, N4936, N246, N2967);
nor NOR3 (N4939, N4926, N3934, N4524);
and AND4 (N4940, N4924, N4830, N2863, N4289);
not NOT1 (N4941, N4937);
buf BUF1 (N4942, N4939);
nand NAND2 (N4943, N4940, N3327);
nand NAND3 (N4944, N4938, N3673, N285);
nand NAND3 (N4945, N4941, N4471, N409);
and AND4 (N4946, N4927, N3074, N3961, N4305);
nand NAND2 (N4947, N4946, N822);
and AND4 (N4948, N4917, N4565, N3606, N3398);
buf BUF1 (N4949, N4942);
and AND3 (N4950, N4944, N4052, N160);
and AND2 (N4951, N4949, N3816);
or OR3 (N4952, N4915, N3620, N4790);
buf BUF1 (N4953, N4948);
nand NAND2 (N4954, N4945, N2721);
nand NAND2 (N4955, N4952, N3210);
nor NOR2 (N4956, N4947, N1059);
nor NOR2 (N4957, N4955, N95);
xor XOR2 (N4958, N4933, N3344);
buf BUF1 (N4959, N4931);
nand NAND4 (N4960, N4958, N3148, N1631, N4936);
buf BUF1 (N4961, N4959);
and AND2 (N4962, N4956, N43);
buf BUF1 (N4963, N4943);
xor XOR2 (N4964, N4962, N3238);
nor NOR4 (N4965, N4964, N4514, N1040, N4206);
nand NAND2 (N4966, N4950, N2597);
not NOT1 (N4967, N4935);
not NOT1 (N4968, N4953);
or OR2 (N4969, N4954, N3438);
or OR3 (N4970, N4968, N1716, N1025);
not NOT1 (N4971, N4970);
nand NAND3 (N4972, N4951, N766, N1581);
nor NOR4 (N4973, N4957, N4644, N3341, N136);
buf BUF1 (N4974, N4966);
and AND4 (N4975, N4972, N354, N1002, N759);
nor NOR4 (N4976, N4967, N2840, N4403, N3201);
xor XOR2 (N4977, N4960, N2765);
nand NAND4 (N4978, N4963, N4259, N2297, N1940);
or OR2 (N4979, N4977, N3783);
nand NAND2 (N4980, N4979, N3447);
nor NOR2 (N4981, N4976, N1062);
not NOT1 (N4982, N4980);
not NOT1 (N4983, N4978);
not NOT1 (N4984, N4974);
buf BUF1 (N4985, N4961);
nor NOR3 (N4986, N4981, N2011, N4408);
nor NOR2 (N4987, N4975, N2689);
not NOT1 (N4988, N4982);
xor XOR2 (N4989, N4973, N4185);
nand NAND3 (N4990, N4983, N1392, N2899);
buf BUF1 (N4991, N4985);
nor NOR3 (N4992, N4986, N1724, N3492);
and AND2 (N4993, N4992, N4590);
or OR2 (N4994, N4969, N2021);
buf BUF1 (N4995, N4984);
nand NAND4 (N4996, N4971, N3917, N3182, N387);
xor XOR2 (N4997, N4989, N561);
nor NOR3 (N4998, N4997, N4670, N4231);
nand NAND2 (N4999, N4993, N4925);
nand NAND2 (N5000, N4995, N1474);
and AND3 (N5001, N5000, N2042, N3460);
buf BUF1 (N5002, N4998);
not NOT1 (N5003, N4994);
buf BUF1 (N5004, N5003);
nor NOR4 (N5005, N4990, N3780, N4005, N4408);
or OR2 (N5006, N5004, N4329);
not NOT1 (N5007, N5005);
buf BUF1 (N5008, N5002);
nand NAND4 (N5009, N4988, N1341, N294, N4312);
or OR4 (N5010, N4991, N3033, N4764, N4053);
nor NOR3 (N5011, N4987, N2768, N2001);
buf BUF1 (N5012, N5011);
nand NAND2 (N5013, N5008, N4870);
not NOT1 (N5014, N5007);
not NOT1 (N5015, N5001);
nor NOR2 (N5016, N5010, N193);
xor XOR2 (N5017, N5016, N4532);
or OR4 (N5018, N5012, N3677, N2948, N2631);
or OR2 (N5019, N4965, N1235);
or OR3 (N5020, N4999, N581, N2825);
buf BUF1 (N5021, N5015);
or OR2 (N5022, N5021, N3635);
not NOT1 (N5023, N5013);
or OR4 (N5024, N5017, N4647, N2005, N2551);
or OR3 (N5025, N5022, N3494, N2098);
nor NOR2 (N5026, N5018, N3272);
buf BUF1 (N5027, N5020);
buf BUF1 (N5028, N5024);
and AND2 (N5029, N5023, N2630);
buf BUF1 (N5030, N5027);
or OR4 (N5031, N5019, N4755, N4648, N51);
nor NOR4 (N5032, N5026, N3474, N1358, N4753);
not NOT1 (N5033, N5032);
and AND4 (N5034, N5028, N3298, N3321, N2688);
xor XOR2 (N5035, N5025, N325);
xor XOR2 (N5036, N5030, N4777);
not NOT1 (N5037, N5035);
xor XOR2 (N5038, N5009, N439);
nor NOR3 (N5039, N5029, N2334, N408);
xor XOR2 (N5040, N5006, N4149);
nor NOR2 (N5041, N5031, N3825);
nand NAND3 (N5042, N4996, N1900, N4391);
not NOT1 (N5043, N5034);
not NOT1 (N5044, N5036);
and AND4 (N5045, N5043, N185, N707, N2193);
buf BUF1 (N5046, N5042);
nand NAND3 (N5047, N5033, N3421, N2637);
and AND2 (N5048, N5040, N2463);
buf BUF1 (N5049, N5039);
not NOT1 (N5050, N5044);
xor XOR2 (N5051, N5047, N4481);
or OR2 (N5052, N5038, N314);
not NOT1 (N5053, N5045);
not NOT1 (N5054, N5052);
or OR3 (N5055, N5051, N2315, N2209);
not NOT1 (N5056, N5055);
not NOT1 (N5057, N5046);
and AND3 (N5058, N5049, N2152, N358);
nor NOR3 (N5059, N5014, N2199, N1958);
xor XOR2 (N5060, N5059, N3771);
nor NOR4 (N5061, N5054, N4419, N3951, N3410);
and AND3 (N5062, N5048, N1565, N504);
buf BUF1 (N5063, N5061);
or OR4 (N5064, N5056, N2181, N495, N2897);
and AND2 (N5065, N5053, N2113);
nor NOR4 (N5066, N5063, N327, N1349, N2816);
or OR2 (N5067, N5058, N1717);
xor XOR2 (N5068, N5062, N3738);
and AND4 (N5069, N5037, N5031, N2305, N2729);
not NOT1 (N5070, N5050);
nor NOR3 (N5071, N5060, N314, N4373);
or OR4 (N5072, N5065, N1758, N2168, N583);
xor XOR2 (N5073, N5069, N1248);
not NOT1 (N5074, N5068);
not NOT1 (N5075, N5074);
and AND3 (N5076, N5073, N3103, N3259);
nand NAND3 (N5077, N5072, N1300, N1867);
nand NAND4 (N5078, N5066, N3472, N2004, N2952);
nor NOR4 (N5079, N5067, N3685, N558, N3847);
and AND3 (N5080, N5071, N4711, N2330);
and AND3 (N5081, N5075, N3803, N1566);
and AND2 (N5082, N5079, N828);
and AND3 (N5083, N5064, N2426, N3592);
and AND3 (N5084, N5076, N3476, N3624);
nand NAND4 (N5085, N5041, N345, N4265, N1048);
nor NOR3 (N5086, N5082, N1050, N3477);
not NOT1 (N5087, N5070);
or OR4 (N5088, N5077, N4610, N4111, N3116);
nand NAND4 (N5089, N5086, N1115, N4172, N1818);
xor XOR2 (N5090, N5057, N3930);
nor NOR3 (N5091, N5089, N1626, N657);
xor XOR2 (N5092, N5080, N2869);
nor NOR2 (N5093, N5088, N2924);
nand NAND4 (N5094, N5090, N4230, N1404, N501);
not NOT1 (N5095, N5094);
nand NAND4 (N5096, N5083, N2023, N4387, N1351);
nand NAND2 (N5097, N5092, N2308);
not NOT1 (N5098, N5084);
buf BUF1 (N5099, N5096);
buf BUF1 (N5100, N5085);
buf BUF1 (N5101, N5100);
nor NOR3 (N5102, N5078, N2820, N2905);
xor XOR2 (N5103, N5102, N699);
xor XOR2 (N5104, N5101, N3983);
nor NOR2 (N5105, N5104, N2914);
xor XOR2 (N5106, N5095, N1075);
or OR2 (N5107, N5093, N4674);
or OR4 (N5108, N5091, N4455, N2027, N1296);
xor XOR2 (N5109, N5106, N1606);
nand NAND4 (N5110, N5107, N2300, N4098, N825);
nor NOR3 (N5111, N5099, N748, N6);
xor XOR2 (N5112, N5109, N4649);
nor NOR3 (N5113, N5105, N2177, N3622);
and AND3 (N5114, N5097, N4699, N4364);
nor NOR3 (N5115, N5112, N4225, N317);
not NOT1 (N5116, N5113);
nor NOR4 (N5117, N5087, N2239, N5034, N1512);
nand NAND4 (N5118, N5098, N871, N3067, N2725);
xor XOR2 (N5119, N5114, N87);
nor NOR3 (N5120, N5108, N3496, N2635);
not NOT1 (N5121, N5081);
buf BUF1 (N5122, N5118);
xor XOR2 (N5123, N5115, N1036);
not NOT1 (N5124, N5121);
nor NOR4 (N5125, N5124, N4539, N4120, N2763);
nand NAND3 (N5126, N5116, N3004, N764);
xor XOR2 (N5127, N5120, N381);
or OR3 (N5128, N5111, N3077, N4928);
not NOT1 (N5129, N5103);
not NOT1 (N5130, N5119);
not NOT1 (N5131, N5125);
not NOT1 (N5132, N5110);
or OR4 (N5133, N5117, N709, N2986, N2449);
buf BUF1 (N5134, N5130);
not NOT1 (N5135, N5129);
not NOT1 (N5136, N5126);
not NOT1 (N5137, N5135);
buf BUF1 (N5138, N5128);
and AND4 (N5139, N5131, N3001, N4892, N4355);
xor XOR2 (N5140, N5127, N1691);
and AND4 (N5141, N5134, N648, N1455, N2155);
xor XOR2 (N5142, N5139, N1164);
xor XOR2 (N5143, N5138, N4505);
xor XOR2 (N5144, N5140, N4098);
nand NAND4 (N5145, N5137, N2401, N3992, N427);
not NOT1 (N5146, N5136);
buf BUF1 (N5147, N5123);
and AND4 (N5148, N5122, N1037, N3360, N1034);
buf BUF1 (N5149, N5133);
xor XOR2 (N5150, N5141, N3575);
nand NAND3 (N5151, N5132, N4372, N4689);
nor NOR2 (N5152, N5145, N3476);
nor NOR4 (N5153, N5150, N5089, N2720, N2860);
nand NAND3 (N5154, N5143, N5119, N3020);
or OR4 (N5155, N5151, N3105, N4023, N2871);
nor NOR3 (N5156, N5155, N947, N1834);
nand NAND4 (N5157, N5148, N2035, N316, N3721);
nand NAND4 (N5158, N5147, N1154, N4605, N4256);
or OR3 (N5159, N5152, N2536, N3193);
nand NAND2 (N5160, N5153, N2556);
not NOT1 (N5161, N5142);
or OR2 (N5162, N5144, N3354);
nand NAND3 (N5163, N5157, N678, N3556);
or OR2 (N5164, N5154, N2870);
buf BUF1 (N5165, N5161);
or OR2 (N5166, N5163, N3842);
and AND4 (N5167, N5156, N4104, N4611, N2074);
and AND4 (N5168, N5158, N3776, N707, N4313);
and AND3 (N5169, N5149, N866, N4765);
buf BUF1 (N5170, N5160);
buf BUF1 (N5171, N5168);
nand NAND3 (N5172, N5165, N4415, N1508);
not NOT1 (N5173, N5164);
not NOT1 (N5174, N5169);
xor XOR2 (N5175, N5162, N2013);
not NOT1 (N5176, N5172);
buf BUF1 (N5177, N5170);
nor NOR4 (N5178, N5171, N3933, N5123, N3318);
nor NOR4 (N5179, N5176, N5019, N640, N3107);
xor XOR2 (N5180, N5178, N3955);
buf BUF1 (N5181, N5175);
and AND2 (N5182, N5174, N4411);
and AND4 (N5183, N5173, N4719, N755, N1733);
xor XOR2 (N5184, N5177, N681);
xor XOR2 (N5185, N5159, N1716);
not NOT1 (N5186, N5184);
nand NAND2 (N5187, N5185, N2969);
and AND3 (N5188, N5181, N1454, N958);
xor XOR2 (N5189, N5166, N2813);
nor NOR2 (N5190, N5146, N2156);
not NOT1 (N5191, N5188);
and AND3 (N5192, N5190, N4831, N960);
xor XOR2 (N5193, N5179, N1957);
xor XOR2 (N5194, N5193, N3974);
nor NOR2 (N5195, N5180, N4338);
and AND4 (N5196, N5187, N1120, N2457, N1114);
and AND3 (N5197, N5167, N431, N4730);
nor NOR4 (N5198, N5192, N1464, N4083, N4762);
not NOT1 (N5199, N5196);
or OR2 (N5200, N5194, N2277);
and AND3 (N5201, N5200, N2552, N935);
and AND3 (N5202, N5186, N1658, N703);
nor NOR3 (N5203, N5198, N1641, N372);
buf BUF1 (N5204, N5191);
nor NOR3 (N5205, N5202, N4155, N491);
nor NOR2 (N5206, N5182, N580);
nor NOR2 (N5207, N5201, N2902);
not NOT1 (N5208, N5203);
buf BUF1 (N5209, N5206);
nor NOR2 (N5210, N5189, N3573);
buf BUF1 (N5211, N5210);
nor NOR3 (N5212, N5195, N3233, N2030);
buf BUF1 (N5213, N5207);
nor NOR2 (N5214, N5213, N314);
nand NAND2 (N5215, N5199, N1310);
not NOT1 (N5216, N5208);
and AND2 (N5217, N5209, N628);
and AND2 (N5218, N5215, N3540);
nand NAND2 (N5219, N5216, N3779);
or OR4 (N5220, N5217, N1623, N2225, N591);
not NOT1 (N5221, N5204);
not NOT1 (N5222, N5219);
xor XOR2 (N5223, N5211, N2423);
xor XOR2 (N5224, N5223, N3093);
not NOT1 (N5225, N5212);
xor XOR2 (N5226, N5205, N3741);
buf BUF1 (N5227, N5224);
or OR3 (N5228, N5222, N1376, N749);
buf BUF1 (N5229, N5226);
buf BUF1 (N5230, N5227);
not NOT1 (N5231, N5225);
nand NAND2 (N5232, N5220, N4573);
and AND3 (N5233, N5197, N1061, N1365);
nand NAND2 (N5234, N5221, N1395);
buf BUF1 (N5235, N5218);
buf BUF1 (N5236, N5183);
nand NAND4 (N5237, N5236, N5224, N1182, N1038);
buf BUF1 (N5238, N5233);
nand NAND3 (N5239, N5214, N3757, N2757);
nand NAND4 (N5240, N5231, N4388, N765, N2837);
not NOT1 (N5241, N5239);
not NOT1 (N5242, N5238);
nand NAND4 (N5243, N5240, N2929, N1479, N3782);
or OR3 (N5244, N5243, N5091, N1891);
buf BUF1 (N5245, N5234);
or OR2 (N5246, N5237, N1686);
or OR4 (N5247, N5246, N700, N4171, N5042);
and AND4 (N5248, N5244, N4793, N705, N136);
not NOT1 (N5249, N5228);
buf BUF1 (N5250, N5235);
and AND4 (N5251, N5250, N2662, N3443, N1756);
and AND2 (N5252, N5245, N628);
not NOT1 (N5253, N5232);
xor XOR2 (N5254, N5252, N2373);
or OR2 (N5255, N5249, N547);
or OR4 (N5256, N5241, N3732, N2091, N2214);
not NOT1 (N5257, N5247);
nand NAND4 (N5258, N5256, N659, N4265, N112);
xor XOR2 (N5259, N5257, N1127);
buf BUF1 (N5260, N5254);
buf BUF1 (N5261, N5248);
and AND3 (N5262, N5260, N5062, N695);
and AND4 (N5263, N5253, N4847, N4638, N1476);
xor XOR2 (N5264, N5259, N2769);
and AND2 (N5265, N5263, N2414);
not NOT1 (N5266, N5255);
xor XOR2 (N5267, N5229, N2416);
xor XOR2 (N5268, N5265, N1492);
or OR4 (N5269, N5266, N5095, N2770, N786);
or OR2 (N5270, N5267, N3521);
xor XOR2 (N5271, N5262, N2667);
nor NOR2 (N5272, N5251, N4567);
xor XOR2 (N5273, N5272, N1127);
nor NOR2 (N5274, N5242, N2856);
nor NOR2 (N5275, N5271, N4534);
nor NOR2 (N5276, N5258, N3567);
or OR4 (N5277, N5274, N2625, N300, N4357);
not NOT1 (N5278, N5275);
not NOT1 (N5279, N5268);
and AND3 (N5280, N5269, N5041, N2254);
buf BUF1 (N5281, N5270);
xor XOR2 (N5282, N5230, N4817);
or OR3 (N5283, N5281, N3191, N1145);
or OR4 (N5284, N5277, N4129, N3009, N4647);
and AND2 (N5285, N5273, N1444);
and AND3 (N5286, N5278, N298, N3709);
xor XOR2 (N5287, N5286, N3906);
or OR4 (N5288, N5280, N2100, N1551, N4573);
xor XOR2 (N5289, N5284, N3523);
xor XOR2 (N5290, N5276, N629);
and AND4 (N5291, N5285, N1905, N1957, N2822);
not NOT1 (N5292, N5289);
not NOT1 (N5293, N5282);
not NOT1 (N5294, N5283);
nand NAND4 (N5295, N5288, N4240, N775, N4245);
xor XOR2 (N5296, N5290, N2416);
or OR4 (N5297, N5291, N4572, N4351, N3684);
not NOT1 (N5298, N5287);
not NOT1 (N5299, N5264);
or OR2 (N5300, N5297, N5079);
not NOT1 (N5301, N5300);
xor XOR2 (N5302, N5296, N1829);
and AND3 (N5303, N5279, N1816, N3605);
or OR2 (N5304, N5295, N1667);
buf BUF1 (N5305, N5301);
buf BUF1 (N5306, N5298);
nand NAND3 (N5307, N5293, N4031, N5284);
nor NOR2 (N5308, N5294, N3470);
xor XOR2 (N5309, N5292, N2499);
not NOT1 (N5310, N5308);
or OR3 (N5311, N5303, N1737, N4365);
nand NAND3 (N5312, N5304, N1201, N4854);
nand NAND4 (N5313, N5302, N4647, N5280, N1036);
buf BUF1 (N5314, N5313);
not NOT1 (N5315, N5310);
nor NOR3 (N5316, N5261, N2694, N259);
nor NOR3 (N5317, N5311, N4135, N2728);
xor XOR2 (N5318, N5312, N1558);
nor NOR3 (N5319, N5316, N2298, N4932);
or OR4 (N5320, N5318, N749, N3754, N1950);
not NOT1 (N5321, N5305);
not NOT1 (N5322, N5321);
buf BUF1 (N5323, N5320);
and AND4 (N5324, N5323, N4452, N624, N561);
not NOT1 (N5325, N5324);
and AND2 (N5326, N5315, N1529);
xor XOR2 (N5327, N5319, N4257);
not NOT1 (N5328, N5314);
nor NOR2 (N5329, N5325, N668);
nand NAND4 (N5330, N5328, N5094, N1270, N762);
or OR4 (N5331, N5329, N3338, N3639, N2960);
nand NAND3 (N5332, N5307, N1776, N4090);
xor XOR2 (N5333, N5332, N5023);
xor XOR2 (N5334, N5326, N405);
xor XOR2 (N5335, N5317, N2614);
buf BUF1 (N5336, N5327);
buf BUF1 (N5337, N5330);
nand NAND3 (N5338, N5333, N2476, N4146);
nor NOR4 (N5339, N5322, N1609, N1378, N686);
xor XOR2 (N5340, N5331, N1614);
and AND4 (N5341, N5309, N3256, N2995, N4);
not NOT1 (N5342, N5337);
not NOT1 (N5343, N5335);
or OR3 (N5344, N5334, N4847, N3497);
xor XOR2 (N5345, N5339, N310);
buf BUF1 (N5346, N5345);
or OR3 (N5347, N5343, N3127, N2455);
or OR2 (N5348, N5306, N1621);
and AND4 (N5349, N5342, N1728, N3908, N795);
xor XOR2 (N5350, N5341, N1248);
nor NOR2 (N5351, N5346, N23);
nor NOR2 (N5352, N5338, N4524);
buf BUF1 (N5353, N5350);
not NOT1 (N5354, N5336);
buf BUF1 (N5355, N5353);
xor XOR2 (N5356, N5351, N5223);
and AND2 (N5357, N5352, N3042);
buf BUF1 (N5358, N5355);
nand NAND3 (N5359, N5344, N416, N1742);
buf BUF1 (N5360, N5340);
or OR4 (N5361, N5299, N960, N1491, N856);
not NOT1 (N5362, N5356);
xor XOR2 (N5363, N5348, N3561);
xor XOR2 (N5364, N5361, N3823);
or OR2 (N5365, N5357, N4970);
or OR2 (N5366, N5362, N4644);
or OR3 (N5367, N5358, N309, N3476);
nor NOR4 (N5368, N5363, N69, N4445, N3383);
nand NAND3 (N5369, N5365, N2987, N4370);
or OR2 (N5370, N5349, N3582);
xor XOR2 (N5371, N5354, N5097);
and AND2 (N5372, N5371, N3660);
xor XOR2 (N5373, N5364, N4037);
not NOT1 (N5374, N5366);
nand NAND3 (N5375, N5359, N2605, N2592);
and AND2 (N5376, N5374, N768);
nor NOR4 (N5377, N5367, N4340, N2354, N4897);
nor NOR2 (N5378, N5347, N1547);
or OR2 (N5379, N5372, N495);
xor XOR2 (N5380, N5376, N5228);
xor XOR2 (N5381, N5378, N2242);
and AND4 (N5382, N5370, N4386, N767, N3863);
and AND3 (N5383, N5380, N4770, N2324);
and AND3 (N5384, N5373, N935, N4462);
nor NOR4 (N5385, N5377, N1790, N3290, N385);
not NOT1 (N5386, N5369);
nor NOR4 (N5387, N5360, N4937, N4058, N3066);
and AND4 (N5388, N5385, N3926, N4719, N4671);
and AND2 (N5389, N5382, N2194);
or OR4 (N5390, N5379, N3604, N790, N358);
nor NOR3 (N5391, N5388, N1345, N1894);
not NOT1 (N5392, N5381);
nor NOR2 (N5393, N5386, N1058);
nor NOR3 (N5394, N5393, N2349, N2006);
not NOT1 (N5395, N5387);
and AND4 (N5396, N5389, N1255, N2294, N2039);
not NOT1 (N5397, N5396);
nand NAND2 (N5398, N5390, N1);
xor XOR2 (N5399, N5368, N1402);
and AND2 (N5400, N5395, N2459);
buf BUF1 (N5401, N5384);
nor NOR3 (N5402, N5394, N5128, N3817);
not NOT1 (N5403, N5401);
buf BUF1 (N5404, N5400);
and AND3 (N5405, N5398, N3435, N4919);
or OR2 (N5406, N5375, N3369);
and AND4 (N5407, N5404, N1388, N2685, N1891);
or OR2 (N5408, N5391, N573);
nor NOR4 (N5409, N5399, N4715, N2627, N722);
and AND4 (N5410, N5383, N239, N765, N1818);
and AND3 (N5411, N5392, N2907, N326);
and AND3 (N5412, N5402, N5289, N519);
xor XOR2 (N5413, N5410, N149);
or OR3 (N5414, N5411, N3989, N4455);
nor NOR3 (N5415, N5414, N3283, N2875);
or OR3 (N5416, N5412, N1934, N4347);
buf BUF1 (N5417, N5403);
or OR2 (N5418, N5397, N3808);
nor NOR3 (N5419, N5418, N3702, N1177);
buf BUF1 (N5420, N5417);
nor NOR4 (N5421, N5405, N5272, N2616, N53);
or OR3 (N5422, N5419, N4300, N1056);
nor NOR4 (N5423, N5413, N3776, N4919, N2296);
buf BUF1 (N5424, N5408);
buf BUF1 (N5425, N5422);
buf BUF1 (N5426, N5423);
nand NAND2 (N5427, N5420, N4536);
nand NAND3 (N5428, N5425, N2823, N828);
or OR4 (N5429, N5407, N2795, N388, N410);
or OR4 (N5430, N5406, N4768, N2566, N2076);
xor XOR2 (N5431, N5430, N3562);
and AND2 (N5432, N5427, N4500);
buf BUF1 (N5433, N5429);
xor XOR2 (N5434, N5426, N745);
buf BUF1 (N5435, N5433);
or OR4 (N5436, N5416, N2160, N4616, N716);
or OR3 (N5437, N5436, N4201, N1673);
or OR2 (N5438, N5424, N869);
nor NOR3 (N5439, N5434, N247, N4984);
buf BUF1 (N5440, N5437);
not NOT1 (N5441, N5409);
nor NOR3 (N5442, N5441, N4875, N2847);
xor XOR2 (N5443, N5435, N4051);
xor XOR2 (N5444, N5438, N2616);
or OR3 (N5445, N5440, N5270, N2743);
buf BUF1 (N5446, N5444);
nor NOR4 (N5447, N5432, N4705, N241, N2916);
xor XOR2 (N5448, N5431, N4183);
and AND4 (N5449, N5443, N2615, N1415, N65);
and AND2 (N5450, N5442, N4401);
or OR2 (N5451, N5415, N1111);
or OR2 (N5452, N5446, N1044);
and AND3 (N5453, N5445, N4255, N843);
or OR3 (N5454, N5449, N4195, N235);
nor NOR3 (N5455, N5428, N2916, N923);
or OR4 (N5456, N5451, N2310, N2179, N3984);
nand NAND2 (N5457, N5439, N479);
not NOT1 (N5458, N5447);
nor NOR4 (N5459, N5448, N1248, N619, N1613);
or OR2 (N5460, N5455, N3858);
and AND2 (N5461, N5421, N4981);
and AND2 (N5462, N5459, N3163);
not NOT1 (N5463, N5453);
not NOT1 (N5464, N5452);
not NOT1 (N5465, N5464);
buf BUF1 (N5466, N5465);
nor NOR2 (N5467, N5466, N1136);
and AND4 (N5468, N5458, N4797, N3967, N3185);
buf BUF1 (N5469, N5457);
buf BUF1 (N5470, N5460);
and AND2 (N5471, N5462, N456);
buf BUF1 (N5472, N5461);
xor XOR2 (N5473, N5469, N2213);
not NOT1 (N5474, N5450);
xor XOR2 (N5475, N5471, N3361);
or OR3 (N5476, N5456, N1862, N4932);
buf BUF1 (N5477, N5470);
not NOT1 (N5478, N5472);
buf BUF1 (N5479, N5474);
and AND4 (N5480, N5476, N482, N2957, N3978);
and AND3 (N5481, N5473, N1222, N3212);
and AND2 (N5482, N5463, N1917);
xor XOR2 (N5483, N5481, N3586);
and AND2 (N5484, N5468, N4402);
or OR4 (N5485, N5475, N3326, N1450, N3993);
xor XOR2 (N5486, N5480, N2918);
buf BUF1 (N5487, N5467);
xor XOR2 (N5488, N5479, N550);
not NOT1 (N5489, N5454);
xor XOR2 (N5490, N5486, N749);
nor NOR4 (N5491, N5490, N3526, N4505, N2500);
not NOT1 (N5492, N5485);
or OR4 (N5493, N5491, N2935, N4068, N2828);
buf BUF1 (N5494, N5493);
nand NAND3 (N5495, N5492, N3928, N17);
or OR3 (N5496, N5494, N2637, N1701);
xor XOR2 (N5497, N5487, N1898);
not NOT1 (N5498, N5495);
xor XOR2 (N5499, N5483, N4110);
nand NAND2 (N5500, N5499, N2991);
and AND2 (N5501, N5477, N1368);
and AND3 (N5502, N5488, N1464, N2732);
nor NOR3 (N5503, N5501, N4166, N1188);
and AND4 (N5504, N5500, N261, N1908, N3819);
or OR3 (N5505, N5498, N5264, N5455);
nand NAND3 (N5506, N5504, N4287, N2013);
or OR2 (N5507, N5484, N4521);
nor NOR4 (N5508, N5502, N2512, N675, N1812);
nand NAND2 (N5509, N5489, N4238);
nand NAND2 (N5510, N5503, N167);
buf BUF1 (N5511, N5507);
nor NOR4 (N5512, N5482, N92, N4793, N2646);
buf BUF1 (N5513, N5512);
not NOT1 (N5514, N5506);
nand NAND2 (N5515, N5509, N2905);
buf BUF1 (N5516, N5508);
nor NOR3 (N5517, N5514, N2768, N3520);
or OR2 (N5518, N5510, N3980);
or OR2 (N5519, N5511, N1705);
nor NOR3 (N5520, N5497, N4858, N4684);
buf BUF1 (N5521, N5518);
not NOT1 (N5522, N5496);
and AND2 (N5523, N5513, N3480);
nand NAND3 (N5524, N5478, N3393, N2587);
not NOT1 (N5525, N5520);
and AND3 (N5526, N5505, N3578, N2187);
or OR4 (N5527, N5515, N3097, N1279, N5486);
xor XOR2 (N5528, N5522, N5352);
buf BUF1 (N5529, N5516);
not NOT1 (N5530, N5528);
or OR2 (N5531, N5529, N2916);
xor XOR2 (N5532, N5521, N2961);
or OR4 (N5533, N5530, N1890, N1125, N5119);
nor NOR2 (N5534, N5523, N3680);
not NOT1 (N5535, N5525);
or OR3 (N5536, N5532, N334, N2981);
nand NAND3 (N5537, N5531, N2677, N4834);
nor NOR4 (N5538, N5533, N990, N1756, N532);
buf BUF1 (N5539, N5517);
nor NOR3 (N5540, N5537, N3725, N3690);
buf BUF1 (N5541, N5536);
nand NAND2 (N5542, N5524, N4625);
xor XOR2 (N5543, N5526, N3755);
not NOT1 (N5544, N5539);
and AND4 (N5545, N5527, N3145, N3847, N3866);
or OR3 (N5546, N5543, N1189, N983);
nand NAND3 (N5547, N5534, N4210, N3500);
nand NAND4 (N5548, N5538, N112, N2269, N106);
nand NAND4 (N5549, N5547, N215, N761, N997);
not NOT1 (N5550, N5548);
or OR2 (N5551, N5550, N1131);
nand NAND4 (N5552, N5546, N3428, N972, N1015);
not NOT1 (N5553, N5552);
xor XOR2 (N5554, N5540, N2383);
or OR4 (N5555, N5553, N2019, N4258, N4890);
nand NAND4 (N5556, N5535, N3661, N102, N3489);
xor XOR2 (N5557, N5544, N4329);
and AND3 (N5558, N5549, N1594, N155);
not NOT1 (N5559, N5541);
xor XOR2 (N5560, N5519, N3365);
or OR2 (N5561, N5556, N1768);
or OR2 (N5562, N5557, N4153);
nor NOR3 (N5563, N5554, N1095, N2824);
xor XOR2 (N5564, N5563, N1175);
nor NOR3 (N5565, N5545, N5, N2712);
xor XOR2 (N5566, N5542, N410);
and AND3 (N5567, N5565, N1914, N4681);
buf BUF1 (N5568, N5555);
nor NOR3 (N5569, N5559, N2409, N4094);
nand NAND3 (N5570, N5568, N3675, N603);
nand NAND2 (N5571, N5564, N2787);
nand NAND2 (N5572, N5551, N2372);
not NOT1 (N5573, N5571);
nor NOR4 (N5574, N5572, N1073, N5011, N1040);
nand NAND4 (N5575, N5562, N1720, N1506, N2653);
not NOT1 (N5576, N5567);
or OR3 (N5577, N5560, N4079, N3883);
xor XOR2 (N5578, N5573, N2982);
nand NAND4 (N5579, N5569, N1168, N3750, N4380);
nor NOR2 (N5580, N5575, N1905);
and AND4 (N5581, N5566, N4444, N238, N4094);
and AND2 (N5582, N5558, N4275);
nor NOR2 (N5583, N5582, N3718);
not NOT1 (N5584, N5583);
and AND2 (N5585, N5579, N128);
buf BUF1 (N5586, N5578);
and AND3 (N5587, N5581, N3480, N396);
or OR3 (N5588, N5577, N709, N4651);
nand NAND3 (N5589, N5586, N3666, N4082);
nand NAND3 (N5590, N5576, N4210, N2223);
xor XOR2 (N5591, N5580, N829);
xor XOR2 (N5592, N5589, N1315);
nand NAND2 (N5593, N5574, N677);
xor XOR2 (N5594, N5584, N4676);
and AND3 (N5595, N5593, N3471, N1123);
buf BUF1 (N5596, N5587);
nand NAND3 (N5597, N5588, N251, N5343);
buf BUF1 (N5598, N5596);
xor XOR2 (N5599, N5595, N389);
nor NOR4 (N5600, N5590, N1047, N5508, N4565);
and AND3 (N5601, N5570, N1486, N1263);
not NOT1 (N5602, N5598);
and AND2 (N5603, N5594, N1346);
nor NOR4 (N5604, N5603, N5132, N5386, N272);
not NOT1 (N5605, N5561);
nor NOR2 (N5606, N5597, N5133);
nand NAND4 (N5607, N5585, N303, N1767, N2230);
nand NAND4 (N5608, N5604, N2187, N5552, N4879);
buf BUF1 (N5609, N5600);
or OR4 (N5610, N5599, N2522, N4866, N71);
xor XOR2 (N5611, N5602, N720);
buf BUF1 (N5612, N5610);
nor NOR4 (N5613, N5612, N449, N4506, N3643);
not NOT1 (N5614, N5611);
not NOT1 (N5615, N5613);
and AND2 (N5616, N5592, N4869);
or OR4 (N5617, N5607, N5167, N2169, N1726);
and AND3 (N5618, N5608, N4391, N1593);
xor XOR2 (N5619, N5618, N144);
not NOT1 (N5620, N5617);
nand NAND2 (N5621, N5606, N3780);
not NOT1 (N5622, N5619);
not NOT1 (N5623, N5620);
or OR4 (N5624, N5605, N2843, N2123, N5068);
or OR3 (N5625, N5621, N232, N3155);
or OR2 (N5626, N5615, N4184);
xor XOR2 (N5627, N5614, N1963);
nand NAND3 (N5628, N5627, N5227, N3752);
nor NOR4 (N5629, N5622, N1992, N2675, N3854);
not NOT1 (N5630, N5609);
nand NAND3 (N5631, N5629, N3579, N4625);
xor XOR2 (N5632, N5626, N2209);
xor XOR2 (N5633, N5628, N28);
nand NAND2 (N5634, N5591, N3135);
not NOT1 (N5635, N5631);
xor XOR2 (N5636, N5601, N1099);
and AND3 (N5637, N5632, N3568, N1326);
nand NAND2 (N5638, N5637, N5563);
and AND4 (N5639, N5634, N5541, N4198, N525);
buf BUF1 (N5640, N5625);
or OR4 (N5641, N5638, N5337, N4679, N1242);
xor XOR2 (N5642, N5639, N1445);
nor NOR3 (N5643, N5616, N2827, N5500);
nor NOR3 (N5644, N5643, N2265, N1994);
nand NAND3 (N5645, N5636, N1680, N4181);
xor XOR2 (N5646, N5624, N3894);
nand NAND4 (N5647, N5644, N1156, N3868, N4662);
nor NOR3 (N5648, N5633, N3632, N481);
or OR4 (N5649, N5645, N2833, N3247, N1866);
and AND3 (N5650, N5630, N810, N2346);
buf BUF1 (N5651, N5648);
nand NAND3 (N5652, N5640, N1980, N3376);
not NOT1 (N5653, N5651);
xor XOR2 (N5654, N5653, N4234);
nor NOR3 (N5655, N5642, N806, N1279);
or OR3 (N5656, N5649, N2662, N4959);
xor XOR2 (N5657, N5650, N1367);
not NOT1 (N5658, N5646);
and AND3 (N5659, N5656, N5612, N5621);
and AND4 (N5660, N5641, N5463, N1216, N200);
nor NOR2 (N5661, N5654, N1376);
buf BUF1 (N5662, N5623);
nand NAND4 (N5663, N5660, N3110, N2136, N4003);
nor NOR4 (N5664, N5647, N785, N3629, N4788);
or OR3 (N5665, N5664, N4594, N4995);
nand NAND4 (N5666, N5661, N3431, N1425, N2724);
and AND2 (N5667, N5655, N5542);
buf BUF1 (N5668, N5663);
nand NAND3 (N5669, N5658, N5605, N736);
buf BUF1 (N5670, N5666);
nand NAND2 (N5671, N5652, N1534);
not NOT1 (N5672, N5635);
or OR3 (N5673, N5659, N2393, N4898);
xor XOR2 (N5674, N5673, N2796);
or OR2 (N5675, N5672, N5150);
and AND2 (N5676, N5670, N5075);
nor NOR4 (N5677, N5669, N3097, N3878, N5383);
not NOT1 (N5678, N5667);
buf BUF1 (N5679, N5676);
not NOT1 (N5680, N5662);
not NOT1 (N5681, N5680);
or OR4 (N5682, N5671, N589, N1703, N3351);
nand NAND3 (N5683, N5675, N994, N386);
not NOT1 (N5684, N5682);
nand NAND4 (N5685, N5678, N2753, N3913, N5162);
buf BUF1 (N5686, N5685);
xor XOR2 (N5687, N5683, N4050);
xor XOR2 (N5688, N5677, N5587);
not NOT1 (N5689, N5684);
not NOT1 (N5690, N5657);
not NOT1 (N5691, N5668);
buf BUF1 (N5692, N5681);
nand NAND4 (N5693, N5679, N1992, N4494, N5153);
not NOT1 (N5694, N5686);
or OR4 (N5695, N5665, N1386, N3284, N4301);
nand NAND2 (N5696, N5689, N3368);
and AND4 (N5697, N5688, N299, N2061, N819);
xor XOR2 (N5698, N5697, N474);
buf BUF1 (N5699, N5694);
buf BUF1 (N5700, N5696);
or OR3 (N5701, N5674, N3587, N4462);
buf BUF1 (N5702, N5699);
not NOT1 (N5703, N5695);
not NOT1 (N5704, N5687);
buf BUF1 (N5705, N5700);
not NOT1 (N5706, N5701);
xor XOR2 (N5707, N5704, N4879);
xor XOR2 (N5708, N5691, N4830);
and AND3 (N5709, N5706, N4265, N2238);
xor XOR2 (N5710, N5698, N1850);
buf BUF1 (N5711, N5707);
not NOT1 (N5712, N5702);
and AND4 (N5713, N5690, N3883, N1532, N2672);
nor NOR2 (N5714, N5711, N629);
and AND2 (N5715, N5712, N3507);
nand NAND4 (N5716, N5709, N1894, N380, N5711);
or OR3 (N5717, N5713, N4805, N5101);
or OR4 (N5718, N5705, N216, N2302, N2390);
not NOT1 (N5719, N5718);
buf BUF1 (N5720, N5708);
not NOT1 (N5721, N5693);
nor NOR2 (N5722, N5710, N2293);
xor XOR2 (N5723, N5716, N1174);
or OR3 (N5724, N5720, N1120, N5572);
not NOT1 (N5725, N5714);
nor NOR4 (N5726, N5724, N4690, N2206, N2068);
not NOT1 (N5727, N5717);
nand NAND4 (N5728, N5715, N2202, N193, N1811);
xor XOR2 (N5729, N5728, N5143);
nand NAND4 (N5730, N5703, N4449, N2331, N4188);
nor NOR4 (N5731, N5719, N3704, N1173, N3219);
buf BUF1 (N5732, N5727);
or OR3 (N5733, N5726, N1094, N3454);
xor XOR2 (N5734, N5725, N2818);
xor XOR2 (N5735, N5730, N2392);
or OR3 (N5736, N5731, N1108, N3322);
or OR4 (N5737, N5692, N5032, N2267, N3378);
nand NAND2 (N5738, N5722, N3272);
nor NOR4 (N5739, N5736, N2333, N3714, N4420);
nor NOR3 (N5740, N5737, N5003, N5183);
nand NAND3 (N5741, N5734, N4187, N123);
nand NAND3 (N5742, N5740, N73, N5254);
xor XOR2 (N5743, N5733, N2825);
not NOT1 (N5744, N5723);
nand NAND2 (N5745, N5721, N3005);
buf BUF1 (N5746, N5738);
or OR4 (N5747, N5745, N4552, N720, N1836);
and AND3 (N5748, N5739, N203, N2004);
not NOT1 (N5749, N5744);
buf BUF1 (N5750, N5732);
nor NOR4 (N5751, N5743, N3175, N732, N1738);
not NOT1 (N5752, N5747);
xor XOR2 (N5753, N5735, N1359);
not NOT1 (N5754, N5750);
not NOT1 (N5755, N5752);
xor XOR2 (N5756, N5751, N971);
not NOT1 (N5757, N5755);
xor XOR2 (N5758, N5756, N439);
not NOT1 (N5759, N5729);
nor NOR2 (N5760, N5748, N1193);
xor XOR2 (N5761, N5746, N1400);
xor XOR2 (N5762, N5753, N791);
nand NAND4 (N5763, N5759, N3705, N2787, N2270);
and AND3 (N5764, N5763, N1825, N2473);
xor XOR2 (N5765, N5757, N5443);
not NOT1 (N5766, N5758);
or OR2 (N5767, N5764, N3642);
nor NOR2 (N5768, N5754, N696);
and AND3 (N5769, N5765, N1197, N3310);
or OR3 (N5770, N5760, N2969, N3127);
and AND2 (N5771, N5741, N5127);
or OR4 (N5772, N5761, N1745, N1881, N1971);
xor XOR2 (N5773, N5771, N2425);
xor XOR2 (N5774, N5770, N1378);
nor NOR4 (N5775, N5742, N256, N3592, N2093);
nor NOR4 (N5776, N5775, N2410, N1637, N1680);
nand NAND3 (N5777, N5776, N5583, N2874);
nand NAND2 (N5778, N5774, N3310);
and AND2 (N5779, N5769, N4497);
buf BUF1 (N5780, N5779);
not NOT1 (N5781, N5766);
nor NOR3 (N5782, N5749, N4266, N5101);
xor XOR2 (N5783, N5777, N3980);
and AND4 (N5784, N5778, N825, N4569, N4172);
and AND2 (N5785, N5783, N5254);
and AND3 (N5786, N5782, N3790, N5153);
nand NAND2 (N5787, N5784, N338);
and AND2 (N5788, N5772, N4842);
not NOT1 (N5789, N5788);
not NOT1 (N5790, N5785);
xor XOR2 (N5791, N5790, N4866);
and AND3 (N5792, N5789, N18, N3724);
nor NOR3 (N5793, N5767, N972, N1874);
nor NOR4 (N5794, N5793, N2013, N185, N615);
xor XOR2 (N5795, N5794, N5005);
nor NOR4 (N5796, N5762, N4126, N2557, N29);
not NOT1 (N5797, N5768);
and AND2 (N5798, N5796, N780);
buf BUF1 (N5799, N5795);
not NOT1 (N5800, N5786);
nor NOR3 (N5801, N5780, N592, N3287);
and AND4 (N5802, N5773, N529, N65, N5582);
xor XOR2 (N5803, N5802, N4322);
or OR4 (N5804, N5791, N4894, N2238, N4326);
xor XOR2 (N5805, N5799, N2726);
or OR4 (N5806, N5801, N1851, N218, N5776);
buf BUF1 (N5807, N5787);
xor XOR2 (N5808, N5804, N1849);
and AND2 (N5809, N5806, N3241);
not NOT1 (N5810, N5809);
or OR2 (N5811, N5797, N815);
not NOT1 (N5812, N5781);
buf BUF1 (N5813, N5812);
nor NOR4 (N5814, N5813, N4860, N4244, N5120);
nand NAND4 (N5815, N5805, N3586, N2948, N3489);
and AND3 (N5816, N5814, N5580, N4098);
not NOT1 (N5817, N5816);
nor NOR4 (N5818, N5810, N3055, N1574, N5345);
and AND3 (N5819, N5792, N1747, N1783);
nor NOR4 (N5820, N5808, N2793, N1660, N4236);
buf BUF1 (N5821, N5819);
nor NOR3 (N5822, N5803, N1095, N3136);
and AND3 (N5823, N5798, N3281, N1758);
or OR4 (N5824, N5823, N1085, N4663, N4660);
not NOT1 (N5825, N5807);
buf BUF1 (N5826, N5815);
nand NAND2 (N5827, N5800, N4813);
not NOT1 (N5828, N5821);
buf BUF1 (N5829, N5828);
buf BUF1 (N5830, N5824);
or OR3 (N5831, N5820, N5073, N1789);
nand NAND3 (N5832, N5826, N3900, N3247);
nand NAND4 (N5833, N5817, N5312, N3880, N5492);
or OR2 (N5834, N5822, N408);
buf BUF1 (N5835, N5831);
and AND2 (N5836, N5818, N858);
nand NAND3 (N5837, N5825, N1434, N4436);
and AND3 (N5838, N5836, N3457, N1805);
and AND4 (N5839, N5835, N3711, N401, N2689);
and AND2 (N5840, N5839, N3923);
nand NAND4 (N5841, N5811, N4994, N620, N275);
buf BUF1 (N5842, N5830);
xor XOR2 (N5843, N5834, N2418);
buf BUF1 (N5844, N5827);
nor NOR3 (N5845, N5843, N2661, N3146);
or OR4 (N5846, N5838, N3177, N2135, N1753);
xor XOR2 (N5847, N5833, N3131);
nand NAND4 (N5848, N5845, N1527, N3857, N1704);
nand NAND2 (N5849, N5841, N902);
xor XOR2 (N5850, N5829, N412);
and AND3 (N5851, N5832, N3921, N887);
or OR4 (N5852, N5846, N3759, N1115, N1826);
xor XOR2 (N5853, N5844, N2127);
not NOT1 (N5854, N5853);
and AND2 (N5855, N5852, N1760);
and AND3 (N5856, N5837, N1039, N4029);
nor NOR4 (N5857, N5849, N176, N1442, N1042);
nor NOR2 (N5858, N5840, N3711);
xor XOR2 (N5859, N5851, N97);
nand NAND2 (N5860, N5842, N5519);
or OR3 (N5861, N5848, N3372, N4304);
and AND2 (N5862, N5859, N2996);
xor XOR2 (N5863, N5857, N492);
not NOT1 (N5864, N5863);
nor NOR4 (N5865, N5858, N1116, N5383, N3284);
not NOT1 (N5866, N5855);
nand NAND3 (N5867, N5862, N179, N4679);
and AND3 (N5868, N5854, N2559, N5426);
and AND2 (N5869, N5856, N1335);
nand NAND4 (N5870, N5869, N885, N3542, N131);
not NOT1 (N5871, N5866);
or OR2 (N5872, N5867, N3459);
buf BUF1 (N5873, N5872);
not NOT1 (N5874, N5860);
buf BUF1 (N5875, N5870);
nor NOR2 (N5876, N5865, N3823);
not NOT1 (N5877, N5876);
buf BUF1 (N5878, N5873);
nand NAND3 (N5879, N5861, N3965, N5030);
xor XOR2 (N5880, N5864, N1467);
xor XOR2 (N5881, N5880, N1631);
buf BUF1 (N5882, N5875);
nor NOR4 (N5883, N5874, N5707, N778, N1223);
or OR4 (N5884, N5847, N3276, N3749, N289);
and AND2 (N5885, N5868, N3588);
nor NOR2 (N5886, N5879, N5536);
buf BUF1 (N5887, N5886);
nand NAND4 (N5888, N5885, N2454, N3401, N3362);
not NOT1 (N5889, N5888);
nor NOR4 (N5890, N5877, N1579, N4434, N439);
or OR3 (N5891, N5890, N3350, N1661);
and AND4 (N5892, N5889, N5240, N5595, N4276);
nand NAND2 (N5893, N5882, N2088);
and AND3 (N5894, N5881, N5570, N3083);
nor NOR2 (N5895, N5893, N2484);
xor XOR2 (N5896, N5850, N3954);
xor XOR2 (N5897, N5895, N3274);
nand NAND4 (N5898, N5871, N4429, N5337, N1054);
or OR3 (N5899, N5891, N498, N4238);
not NOT1 (N5900, N5899);
nor NOR3 (N5901, N5896, N2333, N2567);
buf BUF1 (N5902, N5883);
nor NOR2 (N5903, N5898, N1910);
nand NAND3 (N5904, N5892, N3337, N612);
nand NAND4 (N5905, N5903, N2655, N4524, N2347);
or OR3 (N5906, N5894, N2773, N1194);
nand NAND2 (N5907, N5902, N4366);
buf BUF1 (N5908, N5878);
or OR4 (N5909, N5900, N2733, N5840, N1021);
nor NOR4 (N5910, N5906, N3156, N3874, N4718);
nand NAND3 (N5911, N5901, N4862, N5666);
not NOT1 (N5912, N5911);
xor XOR2 (N5913, N5887, N4122);
and AND2 (N5914, N5912, N4420);
and AND2 (N5915, N5908, N5033);
or OR4 (N5916, N5909, N2741, N2532, N74);
not NOT1 (N5917, N5910);
not NOT1 (N5918, N5897);
buf BUF1 (N5919, N5917);
or OR2 (N5920, N5913, N5052);
or OR3 (N5921, N5884, N117, N2192);
or OR4 (N5922, N5904, N1012, N2520, N1464);
not NOT1 (N5923, N5916);
xor XOR2 (N5924, N5919, N5084);
buf BUF1 (N5925, N5907);
and AND4 (N5926, N5905, N1345, N5228, N12);
nand NAND4 (N5927, N5922, N4142, N1081, N3189);
or OR3 (N5928, N5924, N1540, N972);
or OR2 (N5929, N5926, N2922);
xor XOR2 (N5930, N5920, N1229);
buf BUF1 (N5931, N5923);
and AND2 (N5932, N5930, N5284);
buf BUF1 (N5933, N5929);
nand NAND3 (N5934, N5931, N1522, N3141);
nand NAND4 (N5935, N5914, N5645, N262, N2393);
or OR3 (N5936, N5918, N3524, N1605);
or OR4 (N5937, N5935, N3757, N5296, N2811);
xor XOR2 (N5938, N5921, N1155);
or OR3 (N5939, N5934, N4657, N2409);
xor XOR2 (N5940, N5915, N3801);
nand NAND4 (N5941, N5928, N1848, N1327, N189);
and AND4 (N5942, N5938, N310, N5531, N5233);
not NOT1 (N5943, N5940);
or OR4 (N5944, N5925, N4178, N1138, N835);
nand NAND3 (N5945, N5932, N597, N5087);
or OR2 (N5946, N5936, N3505);
xor XOR2 (N5947, N5942, N5356);
xor XOR2 (N5948, N5945, N3258);
nor NOR3 (N5949, N5939, N2148, N194);
xor XOR2 (N5950, N5949, N501);
and AND3 (N5951, N5950, N4805, N3429);
nor NOR3 (N5952, N5933, N3308, N2158);
or OR3 (N5953, N5948, N3210, N711);
buf BUF1 (N5954, N5953);
buf BUF1 (N5955, N5954);
xor XOR2 (N5956, N5946, N431);
buf BUF1 (N5957, N5943);
and AND2 (N5958, N5956, N76);
buf BUF1 (N5959, N5958);
nand NAND4 (N5960, N5937, N2565, N3986, N1351);
or OR4 (N5961, N5957, N2943, N2810, N60);
not NOT1 (N5962, N5944);
or OR4 (N5963, N5947, N604, N4885, N4411);
nand NAND4 (N5964, N5962, N4089, N4978, N4145);
xor XOR2 (N5965, N5960, N4852);
and AND3 (N5966, N5964, N3095, N4662);
buf BUF1 (N5967, N5951);
or OR4 (N5968, N5927, N2692, N3964, N3909);
buf BUF1 (N5969, N5965);
not NOT1 (N5970, N5967);
not NOT1 (N5971, N5966);
nand NAND3 (N5972, N5963, N1369, N251);
xor XOR2 (N5973, N5941, N1480);
or OR4 (N5974, N5961, N2134, N4925, N5640);
or OR2 (N5975, N5955, N3098);
nor NOR4 (N5976, N5971, N4524, N4905, N1858);
xor XOR2 (N5977, N5973, N1817);
buf BUF1 (N5978, N5975);
and AND4 (N5979, N5970, N3018, N5867, N2479);
not NOT1 (N5980, N5972);
or OR4 (N5981, N5969, N2634, N5733, N592);
buf BUF1 (N5982, N5976);
nor NOR4 (N5983, N5980, N1501, N5163, N5023);
or OR2 (N5984, N5959, N1962);
buf BUF1 (N5985, N5968);
xor XOR2 (N5986, N5977, N109);
or OR3 (N5987, N5978, N1297, N3466);
xor XOR2 (N5988, N5983, N900);
or OR2 (N5989, N5952, N1268);
xor XOR2 (N5990, N5989, N1106);
buf BUF1 (N5991, N5979);
or OR4 (N5992, N5988, N3559, N1128, N4376);
not NOT1 (N5993, N5981);
buf BUF1 (N5994, N5992);
not NOT1 (N5995, N5990);
xor XOR2 (N5996, N5974, N4361);
and AND4 (N5997, N5987, N5416, N3121, N2509);
xor XOR2 (N5998, N5994, N5975);
nor NOR3 (N5999, N5998, N2839, N2795);
or OR2 (N6000, N5984, N4588);
not NOT1 (N6001, N5985);
nor NOR2 (N6002, N5997, N67);
buf BUF1 (N6003, N6002);
and AND3 (N6004, N6000, N1916, N4950);
and AND2 (N6005, N5986, N738);
buf BUF1 (N6006, N5995);
not NOT1 (N6007, N5996);
nor NOR4 (N6008, N6003, N5910, N2794, N123);
and AND4 (N6009, N6001, N5322, N1707, N2539);
or OR3 (N6010, N6006, N3151, N1566);
and AND3 (N6011, N6005, N5047, N1396);
and AND3 (N6012, N5999, N5294, N2221);
nor NOR2 (N6013, N6008, N1388);
nand NAND4 (N6014, N5993, N3405, N1128, N3376);
xor XOR2 (N6015, N5982, N141);
or OR2 (N6016, N6012, N105);
not NOT1 (N6017, N6014);
nor NOR2 (N6018, N6013, N3934);
xor XOR2 (N6019, N6011, N3716);
not NOT1 (N6020, N6017);
xor XOR2 (N6021, N6009, N2356);
or OR2 (N6022, N6019, N1424);
buf BUF1 (N6023, N6022);
not NOT1 (N6024, N6015);
buf BUF1 (N6025, N6004);
nor NOR2 (N6026, N6018, N5488);
xor XOR2 (N6027, N5991, N3646);
and AND4 (N6028, N6026, N4865, N3174, N3232);
and AND4 (N6029, N6024, N5619, N2219, N4230);
and AND2 (N6030, N6007, N703);
not NOT1 (N6031, N6016);
nor NOR3 (N6032, N6028, N9, N3064);
buf BUF1 (N6033, N6023);
buf BUF1 (N6034, N6021);
and AND3 (N6035, N6025, N1074, N2424);
and AND2 (N6036, N6027, N2774);
not NOT1 (N6037, N6010);
nor NOR2 (N6038, N6034, N977);
xor XOR2 (N6039, N6038, N424);
buf BUF1 (N6040, N6037);
xor XOR2 (N6041, N6040, N3716);
or OR2 (N6042, N6041, N5621);
buf BUF1 (N6043, N6031);
xor XOR2 (N6044, N6039, N5726);
xor XOR2 (N6045, N6043, N5946);
xor XOR2 (N6046, N6042, N4758);
or OR4 (N6047, N6036, N4072, N4457, N3507);
buf BUF1 (N6048, N6033);
nor NOR3 (N6049, N6030, N4305, N2065);
not NOT1 (N6050, N6044);
nor NOR3 (N6051, N6032, N27, N4408);
xor XOR2 (N6052, N6048, N1953);
nor NOR4 (N6053, N6035, N1422, N1929, N1026);
buf BUF1 (N6054, N6020);
nand NAND4 (N6055, N6046, N3177, N3264, N5662);
nand NAND3 (N6056, N6045, N2889, N3971);
nor NOR2 (N6057, N6051, N5572);
nor NOR2 (N6058, N6057, N414);
buf BUF1 (N6059, N6054);
xor XOR2 (N6060, N6053, N428);
buf BUF1 (N6061, N6047);
and AND2 (N6062, N6052, N4628);
nor NOR3 (N6063, N6059, N5953, N3215);
not NOT1 (N6064, N6050);
not NOT1 (N6065, N6061);
not NOT1 (N6066, N6056);
xor XOR2 (N6067, N6058, N5644);
nand NAND3 (N6068, N6060, N4399, N4212);
or OR2 (N6069, N6066, N5619);
buf BUF1 (N6070, N6055);
and AND4 (N6071, N6068, N3361, N3382, N681);
and AND4 (N6072, N6029, N3970, N3705, N1744);
nor NOR3 (N6073, N6072, N247, N1957);
xor XOR2 (N6074, N6073, N5053);
nand NAND4 (N6075, N6069, N5, N1900, N5062);
nor NOR3 (N6076, N6049, N378, N548);
or OR2 (N6077, N6064, N4257);
xor XOR2 (N6078, N6067, N4556);
xor XOR2 (N6079, N6070, N5749);
nor NOR4 (N6080, N6062, N5338, N2490, N424);
and AND4 (N6081, N6079, N4437, N5465, N1547);
not NOT1 (N6082, N6074);
nand NAND4 (N6083, N6063, N1679, N4903, N3100);
and AND3 (N6084, N6080, N1208, N3495);
and AND4 (N6085, N6071, N3426, N4718, N4459);
nand NAND2 (N6086, N6083, N5185);
buf BUF1 (N6087, N6075);
buf BUF1 (N6088, N6077);
and AND2 (N6089, N6085, N5656);
buf BUF1 (N6090, N6076);
not NOT1 (N6091, N6086);
or OR3 (N6092, N6065, N5643, N3416);
or OR3 (N6093, N6092, N370, N3550);
not NOT1 (N6094, N6089);
xor XOR2 (N6095, N6087, N3465);
nand NAND2 (N6096, N6091, N973);
nand NAND3 (N6097, N6078, N131, N2032);
or OR3 (N6098, N6097, N3453, N3356);
and AND2 (N6099, N6082, N5059);
buf BUF1 (N6100, N6090);
nand NAND2 (N6101, N6100, N1893);
buf BUF1 (N6102, N6093);
and AND2 (N6103, N6081, N5021);
and AND4 (N6104, N6084, N5546, N5763, N5565);
nor NOR4 (N6105, N6102, N4979, N542, N5794);
or OR2 (N6106, N6104, N3917);
and AND2 (N6107, N6094, N5082);
nand NAND2 (N6108, N6095, N4541);
not NOT1 (N6109, N6099);
xor XOR2 (N6110, N6096, N4721);
buf BUF1 (N6111, N6108);
not NOT1 (N6112, N6106);
xor XOR2 (N6113, N6098, N87);
or OR4 (N6114, N6113, N1577, N246, N5460);
or OR3 (N6115, N6112, N250, N2200);
nor NOR2 (N6116, N6114, N1359);
or OR3 (N6117, N6116, N2997, N1298);
xor XOR2 (N6118, N6103, N2347);
nand NAND3 (N6119, N6115, N4899, N3396);
buf BUF1 (N6120, N6109);
xor XOR2 (N6121, N6110, N1486);
nor NOR3 (N6122, N6088, N4333, N3003);
not NOT1 (N6123, N6120);
or OR4 (N6124, N6123, N2681, N635, N1036);
nor NOR4 (N6125, N6118, N3211, N3317, N5907);
nand NAND4 (N6126, N6101, N4380, N4511, N608);
buf BUF1 (N6127, N6117);
xor XOR2 (N6128, N6125, N700);
or OR4 (N6129, N6126, N4490, N1612, N4311);
and AND2 (N6130, N6127, N5541);
and AND2 (N6131, N6128, N5483);
nand NAND2 (N6132, N6124, N5208);
not NOT1 (N6133, N6119);
and AND2 (N6134, N6107, N813);
buf BUF1 (N6135, N6122);
nand NAND2 (N6136, N6111, N2799);
and AND3 (N6137, N6121, N983, N1103);
nand NAND2 (N6138, N6132, N1586);
xor XOR2 (N6139, N6133, N5733);
nor NOR3 (N6140, N6130, N3895, N4022);
not NOT1 (N6141, N6129);
not NOT1 (N6142, N6138);
buf BUF1 (N6143, N6136);
not NOT1 (N6144, N6137);
not NOT1 (N6145, N6131);
and AND2 (N6146, N6144, N1109);
and AND4 (N6147, N6139, N254, N4114, N4044);
xor XOR2 (N6148, N6105, N4293);
buf BUF1 (N6149, N6140);
nor NOR4 (N6150, N6134, N2679, N5003, N4214);
or OR4 (N6151, N6143, N2754, N5457, N619);
nand NAND3 (N6152, N6141, N3420, N3160);
not NOT1 (N6153, N6135);
xor XOR2 (N6154, N6151, N2027);
buf BUF1 (N6155, N6152);
nor NOR3 (N6156, N6149, N2273, N4736);
xor XOR2 (N6157, N6148, N1619);
nor NOR3 (N6158, N6153, N4467, N2134);
or OR3 (N6159, N6142, N4816, N4554);
xor XOR2 (N6160, N6146, N4040);
xor XOR2 (N6161, N6154, N142);
nand NAND3 (N6162, N6159, N3837, N3816);
nand NAND2 (N6163, N6155, N3373);
and AND3 (N6164, N6157, N5315, N4455);
buf BUF1 (N6165, N6150);
and AND2 (N6166, N6162, N5400);
or OR4 (N6167, N6160, N4240, N806, N5757);
not NOT1 (N6168, N6164);
nand NAND4 (N6169, N6167, N1288, N2632, N976);
nor NOR3 (N6170, N6156, N3427, N4653);
buf BUF1 (N6171, N6161);
or OR4 (N6172, N6171, N3668, N3134, N1827);
nor NOR2 (N6173, N6158, N337);
or OR3 (N6174, N6165, N3390, N5263);
not NOT1 (N6175, N6169);
not NOT1 (N6176, N6170);
buf BUF1 (N6177, N6145);
nand NAND3 (N6178, N6147, N4848, N3789);
xor XOR2 (N6179, N6172, N3662);
not NOT1 (N6180, N6168);
nand NAND3 (N6181, N6163, N811, N4011);
and AND2 (N6182, N6181, N1129);
nor NOR2 (N6183, N6178, N863);
nor NOR4 (N6184, N6174, N3868, N1421, N208);
nand NAND4 (N6185, N6173, N607, N563, N4735);
or OR4 (N6186, N6166, N2295, N2851, N5867);
xor XOR2 (N6187, N6182, N2152);
not NOT1 (N6188, N6185);
buf BUF1 (N6189, N6187);
and AND2 (N6190, N6189, N3634);
not NOT1 (N6191, N6190);
xor XOR2 (N6192, N6191, N2675);
nor NOR4 (N6193, N6175, N3440, N795, N2359);
or OR3 (N6194, N6183, N1165, N5180);
nor NOR3 (N6195, N6192, N1178, N531);
xor XOR2 (N6196, N6194, N1615);
and AND3 (N6197, N6177, N3928, N3407);
or OR4 (N6198, N6186, N5254, N4824, N195);
not NOT1 (N6199, N6198);
buf BUF1 (N6200, N6179);
nor NOR3 (N6201, N6193, N2979, N1238);
and AND2 (N6202, N6180, N2983);
nand NAND4 (N6203, N6199, N3225, N2495, N3827);
and AND2 (N6204, N6201, N3781);
not NOT1 (N6205, N6184);
not NOT1 (N6206, N6203);
nand NAND2 (N6207, N6204, N2228);
not NOT1 (N6208, N6195);
nor NOR2 (N6209, N6196, N3992);
xor XOR2 (N6210, N6209, N5696);
nand NAND2 (N6211, N6208, N1314);
nand NAND4 (N6212, N6211, N3444, N4234, N931);
xor XOR2 (N6213, N6176, N2995);
not NOT1 (N6214, N6188);
buf BUF1 (N6215, N6206);
nor NOR3 (N6216, N6197, N3028, N94);
nand NAND4 (N6217, N6205, N2093, N2561, N6198);
nand NAND3 (N6218, N6207, N4146, N5900);
nor NOR3 (N6219, N6218, N6012, N3933);
xor XOR2 (N6220, N6213, N3008);
xor XOR2 (N6221, N6200, N5414);
buf BUF1 (N6222, N6214);
buf BUF1 (N6223, N6220);
or OR2 (N6224, N6217, N2058);
not NOT1 (N6225, N6210);
nor NOR2 (N6226, N6212, N2214);
not NOT1 (N6227, N6216);
and AND4 (N6228, N6223, N1943, N1492, N1241);
and AND2 (N6229, N6215, N2249);
buf BUF1 (N6230, N6202);
nand NAND4 (N6231, N6225, N4076, N5327, N293);
or OR3 (N6232, N6231, N3030, N5306);
xor XOR2 (N6233, N6229, N2861);
not NOT1 (N6234, N6219);
xor XOR2 (N6235, N6228, N1069);
xor XOR2 (N6236, N6222, N2720);
nand NAND3 (N6237, N6221, N1151, N162);
and AND2 (N6238, N6224, N4117);
buf BUF1 (N6239, N6236);
and AND4 (N6240, N6237, N4398, N1891, N507);
nand NAND4 (N6241, N6226, N5738, N634, N4170);
or OR2 (N6242, N6234, N1270);
and AND3 (N6243, N6238, N5918, N6197);
nor NOR4 (N6244, N6239, N1634, N3733, N2903);
and AND2 (N6245, N6244, N28);
and AND2 (N6246, N6233, N5901);
not NOT1 (N6247, N6230);
and AND4 (N6248, N6247, N3096, N5901, N253);
not NOT1 (N6249, N6243);
not NOT1 (N6250, N6246);
buf BUF1 (N6251, N6227);
buf BUF1 (N6252, N6251);
not NOT1 (N6253, N6242);
not NOT1 (N6254, N6245);
xor XOR2 (N6255, N6249, N5882);
not NOT1 (N6256, N6241);
not NOT1 (N6257, N6248);
nand NAND2 (N6258, N6257, N6196);
not NOT1 (N6259, N6240);
and AND3 (N6260, N6258, N2159, N565);
xor XOR2 (N6261, N6254, N4704);
not NOT1 (N6262, N6261);
xor XOR2 (N6263, N6253, N4717);
buf BUF1 (N6264, N6262);
and AND4 (N6265, N6263, N4569, N4606, N582);
buf BUF1 (N6266, N6232);
not NOT1 (N6267, N6252);
or OR2 (N6268, N6260, N3748);
buf BUF1 (N6269, N6256);
or OR4 (N6270, N6250, N4068, N3462, N6009);
not NOT1 (N6271, N6255);
nand NAND4 (N6272, N6269, N4343, N330, N4556);
not NOT1 (N6273, N6271);
or OR3 (N6274, N6273, N5937, N1085);
xor XOR2 (N6275, N6235, N1914);
nor NOR4 (N6276, N6265, N5931, N6166, N143);
buf BUF1 (N6277, N6266);
and AND4 (N6278, N6267, N5128, N2612, N360);
xor XOR2 (N6279, N6259, N1333);
xor XOR2 (N6280, N6274, N2028);
nor NOR4 (N6281, N6280, N3924, N5359, N3221);
xor XOR2 (N6282, N6270, N4761);
not NOT1 (N6283, N6268);
or OR4 (N6284, N6282, N1253, N3882, N4764);
buf BUF1 (N6285, N6275);
nor NOR4 (N6286, N6272, N5895, N4421, N4986);
buf BUF1 (N6287, N6285);
and AND4 (N6288, N6287, N1375, N3973, N5029);
or OR2 (N6289, N6288, N2695);
nand NAND4 (N6290, N6289, N1604, N3792, N886);
xor XOR2 (N6291, N6281, N1033);
nand NAND4 (N6292, N6290, N2255, N995, N4890);
and AND2 (N6293, N6264, N2070);
nand NAND3 (N6294, N6276, N4619, N4487);
or OR4 (N6295, N6294, N2594, N5276, N4550);
xor XOR2 (N6296, N6292, N1367);
nand NAND2 (N6297, N6278, N2139);
or OR4 (N6298, N6297, N1461, N5916, N5142);
not NOT1 (N6299, N6277);
nor NOR3 (N6300, N6298, N764, N3973);
buf BUF1 (N6301, N6299);
or OR4 (N6302, N6286, N3067, N1499, N5586);
not NOT1 (N6303, N6296);
not NOT1 (N6304, N6283);
xor XOR2 (N6305, N6291, N5990);
and AND3 (N6306, N6301, N1654, N5164);
and AND4 (N6307, N6279, N5092, N4158, N211);
nor NOR3 (N6308, N6284, N5012, N1058);
xor XOR2 (N6309, N6304, N3721);
nor NOR2 (N6310, N6293, N5962);
nand NAND3 (N6311, N6310, N4528, N1641);
or OR2 (N6312, N6303, N4381);
and AND3 (N6313, N6300, N1361, N4050);
xor XOR2 (N6314, N6311, N5702);
nor NOR2 (N6315, N6302, N3669);
nor NOR4 (N6316, N6305, N2150, N1590, N2290);
not NOT1 (N6317, N6307);
xor XOR2 (N6318, N6309, N4181);
or OR3 (N6319, N6314, N6042, N700);
nor NOR4 (N6320, N6308, N3471, N1478, N5854);
and AND2 (N6321, N6306, N2366);
or OR4 (N6322, N6318, N841, N1393, N3002);
or OR4 (N6323, N6319, N2763, N5636, N3582);
and AND4 (N6324, N6295, N467, N3419, N3457);
not NOT1 (N6325, N6315);
and AND4 (N6326, N6322, N2969, N1131, N6049);
buf BUF1 (N6327, N6320);
xor XOR2 (N6328, N6316, N499);
not NOT1 (N6329, N6323);
nor NOR2 (N6330, N6325, N4243);
nor NOR2 (N6331, N6327, N4494);
and AND4 (N6332, N6330, N3676, N5929, N5502);
xor XOR2 (N6333, N6326, N2773);
xor XOR2 (N6334, N6312, N1157);
or OR2 (N6335, N6332, N185);
not NOT1 (N6336, N6331);
not NOT1 (N6337, N6313);
xor XOR2 (N6338, N6324, N4342);
nor NOR3 (N6339, N6337, N3807, N3513);
xor XOR2 (N6340, N6336, N5791);
nor NOR4 (N6341, N6321, N4973, N1357, N2854);
nor NOR3 (N6342, N6334, N3417, N3222);
or OR4 (N6343, N6329, N2626, N5468, N4212);
or OR2 (N6344, N6342, N3452);
or OR2 (N6345, N6341, N1613);
or OR2 (N6346, N6339, N5486);
and AND4 (N6347, N6345, N3928, N2517, N3481);
or OR3 (N6348, N6344, N6060, N723);
nand NAND2 (N6349, N6348, N4338);
nand NAND2 (N6350, N6340, N675);
buf BUF1 (N6351, N6346);
not NOT1 (N6352, N6328);
buf BUF1 (N6353, N6333);
buf BUF1 (N6354, N6343);
not NOT1 (N6355, N6353);
nor NOR3 (N6356, N6347, N1548, N918);
xor XOR2 (N6357, N6352, N351);
nand NAND2 (N6358, N6357, N5861);
xor XOR2 (N6359, N6355, N5427);
buf BUF1 (N6360, N6359);
xor XOR2 (N6361, N6354, N2563);
xor XOR2 (N6362, N6360, N1265);
not NOT1 (N6363, N6349);
not NOT1 (N6364, N6350);
and AND3 (N6365, N6362, N3182, N3155);
nand NAND3 (N6366, N6335, N3539, N5318);
not NOT1 (N6367, N6363);
buf BUF1 (N6368, N6356);
not NOT1 (N6369, N6364);
nand NAND2 (N6370, N6367, N4480);
or OR2 (N6371, N6370, N4305);
xor XOR2 (N6372, N6365, N6224);
not NOT1 (N6373, N6361);
nand NAND3 (N6374, N6351, N1231, N5768);
buf BUF1 (N6375, N6358);
buf BUF1 (N6376, N6371);
nor NOR4 (N6377, N6375, N5402, N3917, N1130);
and AND4 (N6378, N6376, N1347, N1125, N4963);
buf BUF1 (N6379, N6317);
or OR3 (N6380, N6372, N3455, N3854);
buf BUF1 (N6381, N6374);
nor NOR4 (N6382, N6338, N5804, N1808, N3927);
and AND2 (N6383, N6380, N3405);
or OR3 (N6384, N6378, N118, N3132);
or OR3 (N6385, N6384, N2990, N4674);
not NOT1 (N6386, N6369);
nand NAND4 (N6387, N6386, N517, N1651, N5972);
nand NAND3 (N6388, N6381, N2369, N242);
xor XOR2 (N6389, N6385, N72);
or OR3 (N6390, N6387, N4325, N3267);
nor NOR2 (N6391, N6389, N3204);
and AND3 (N6392, N6383, N5352, N5869);
xor XOR2 (N6393, N6388, N2277);
and AND4 (N6394, N6391, N5671, N4318, N2813);
xor XOR2 (N6395, N6393, N5583);
or OR3 (N6396, N6392, N1068, N1685);
or OR3 (N6397, N6377, N2000, N5913);
nand NAND3 (N6398, N6382, N3500, N6012);
or OR3 (N6399, N6398, N3170, N3007);
xor XOR2 (N6400, N6390, N4877);
and AND4 (N6401, N6399, N3697, N6388, N600);
nand NAND4 (N6402, N6368, N3050, N2452, N2339);
or OR4 (N6403, N6402, N3404, N4295, N1189);
and AND4 (N6404, N6400, N4844, N1560, N428);
or OR4 (N6405, N6373, N829, N4721, N2811);
not NOT1 (N6406, N6394);
and AND4 (N6407, N6366, N2064, N6153, N3011);
nor NOR2 (N6408, N6395, N870);
nor NOR3 (N6409, N6401, N2890, N253);
nor NOR4 (N6410, N6379, N4135, N3136, N3235);
nor NOR2 (N6411, N6403, N1141);
nand NAND4 (N6412, N6410, N1506, N982, N5389);
buf BUF1 (N6413, N6406);
or OR4 (N6414, N6412, N332, N3925, N5254);
or OR4 (N6415, N6414, N3299, N5878, N607);
endmodule