// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;

output N911,N894,N910,N909,N896,N876,N905,N908,N883,N912;

nor NOR3 (N13, N6, N9, N9);
nand NAND2 (N14, N8, N5);
or OR2 (N15, N3, N1);
xor XOR2 (N16, N14, N11);
xor XOR2 (N17, N8, N10);
buf BUF1 (N18, N3);
and AND3 (N19, N8, N9, N6);
and AND2 (N20, N8, N17);
nor NOR3 (N21, N18, N13, N8);
nor NOR2 (N22, N13, N17);
or OR3 (N23, N9, N22, N4);
nand NAND2 (N24, N13, N3);
nand NAND4 (N25, N10, N13, N12, N18);
buf BUF1 (N26, N23);
buf BUF1 (N27, N1);
buf BUF1 (N28, N13);
or OR3 (N29, N27, N25, N21);
buf BUF1 (N30, N6);
xor XOR2 (N31, N10, N3);
buf BUF1 (N32, N28);
nand NAND4 (N33, N30, N32, N25, N28);
nor NOR4 (N34, N11, N9, N13, N8);
and AND2 (N35, N31, N3);
or OR3 (N36, N33, N6, N10);
and AND4 (N37, N34, N12, N6, N33);
nor NOR3 (N38, N20, N1, N2);
not NOT1 (N39, N29);
xor XOR2 (N40, N15, N22);
nand NAND4 (N41, N26, N6, N32, N10);
not NOT1 (N42, N38);
or OR4 (N43, N16, N38, N1, N7);
or OR4 (N44, N40, N11, N37, N32);
buf BUF1 (N45, N32);
buf BUF1 (N46, N24);
not NOT1 (N47, N43);
not NOT1 (N48, N45);
nand NAND2 (N49, N44, N41);
nor NOR3 (N50, N16, N22, N40);
buf BUF1 (N51, N35);
not NOT1 (N52, N50);
buf BUF1 (N53, N52);
or OR4 (N54, N47, N28, N28, N12);
xor XOR2 (N55, N53, N14);
not NOT1 (N56, N55);
nand NAND3 (N57, N56, N16, N46);
nand NAND3 (N58, N39, N28, N52);
nand NAND2 (N59, N28, N36);
nand NAND3 (N60, N32, N58, N50);
and AND3 (N61, N26, N43, N4);
nor NOR3 (N62, N54, N8, N16);
buf BUF1 (N63, N57);
or OR2 (N64, N51, N58);
nand NAND4 (N65, N61, N6, N15, N5);
nand NAND4 (N66, N19, N29, N55, N54);
not NOT1 (N67, N49);
not NOT1 (N68, N59);
and AND4 (N69, N62, N28, N51, N9);
nor NOR2 (N70, N42, N37);
buf BUF1 (N71, N70);
nand NAND3 (N72, N71, N35, N12);
nor NOR2 (N73, N63, N39);
not NOT1 (N74, N72);
and AND2 (N75, N64, N7);
xor XOR2 (N76, N65, N42);
xor XOR2 (N77, N74, N25);
nor NOR3 (N78, N77, N27, N19);
not NOT1 (N79, N67);
nor NOR2 (N80, N78, N8);
xor XOR2 (N81, N69, N74);
buf BUF1 (N82, N73);
xor XOR2 (N83, N82, N76);
xor XOR2 (N84, N67, N49);
xor XOR2 (N85, N84, N76);
or OR3 (N86, N48, N46, N33);
or OR4 (N87, N68, N3, N19, N83);
xor XOR2 (N88, N43, N53);
buf BUF1 (N89, N81);
xor XOR2 (N90, N80, N34);
xor XOR2 (N91, N87, N1);
or OR4 (N92, N79, N31, N70, N21);
nand NAND2 (N93, N92, N64);
xor XOR2 (N94, N91, N47);
nand NAND4 (N95, N85, N28, N23, N10);
nand NAND3 (N96, N60, N28, N66);
not NOT1 (N97, N82);
or OR4 (N98, N95, N83, N39, N64);
buf BUF1 (N99, N90);
and AND2 (N100, N99, N45);
nor NOR4 (N101, N97, N26, N99, N93);
xor XOR2 (N102, N56, N12);
not NOT1 (N103, N98);
nand NAND4 (N104, N94, N85, N35, N14);
xor XOR2 (N105, N102, N64);
nand NAND3 (N106, N100, N97, N100);
nand NAND2 (N107, N104, N69);
and AND3 (N108, N107, N80, N88);
nor NOR3 (N109, N91, N85, N78);
xor XOR2 (N110, N108, N56);
nand NAND3 (N111, N103, N89, N38);
or OR4 (N112, N55, N81, N97, N57);
and AND2 (N113, N109, N54);
and AND4 (N114, N111, N106, N68, N74);
nor NOR3 (N115, N36, N35, N102);
and AND3 (N116, N115, N30, N92);
xor XOR2 (N117, N101, N108);
not NOT1 (N118, N112);
nor NOR3 (N119, N116, N7, N111);
not NOT1 (N120, N113);
or OR3 (N121, N96, N28, N72);
nand NAND2 (N122, N121, N10);
xor XOR2 (N123, N122, N88);
not NOT1 (N124, N123);
xor XOR2 (N125, N75, N34);
and AND4 (N126, N117, N47, N64, N122);
not NOT1 (N127, N110);
nand NAND4 (N128, N114, N70, N8, N19);
not NOT1 (N129, N124);
not NOT1 (N130, N119);
buf BUF1 (N131, N126);
buf BUF1 (N132, N86);
not NOT1 (N133, N131);
and AND3 (N134, N120, N93, N101);
xor XOR2 (N135, N118, N93);
not NOT1 (N136, N129);
buf BUF1 (N137, N130);
not NOT1 (N138, N132);
nand NAND3 (N139, N128, N92, N60);
and AND2 (N140, N137, N24);
xor XOR2 (N141, N138, N10);
buf BUF1 (N142, N127);
and AND4 (N143, N133, N34, N26, N117);
and AND3 (N144, N105, N29, N119);
nor NOR2 (N145, N141, N103);
xor XOR2 (N146, N144, N126);
buf BUF1 (N147, N134);
nor NOR4 (N148, N140, N24, N38, N91);
or OR3 (N149, N125, N51, N22);
or OR4 (N150, N145, N33, N80, N40);
buf BUF1 (N151, N136);
or OR3 (N152, N151, N25, N17);
nand NAND4 (N153, N139, N148, N22, N134);
nor NOR3 (N154, N133, N96, N31);
buf BUF1 (N155, N143);
buf BUF1 (N156, N152);
xor XOR2 (N157, N142, N90);
nand NAND2 (N158, N157, N42);
nand NAND2 (N159, N135, N131);
or OR4 (N160, N146, N30, N64, N95);
nand NAND3 (N161, N154, N137, N111);
and AND2 (N162, N160, N143);
xor XOR2 (N163, N161, N51);
and AND4 (N164, N147, N47, N88, N22);
or OR2 (N165, N158, N11);
buf BUF1 (N166, N159);
nand NAND4 (N167, N162, N81, N147, N104);
or OR4 (N168, N167, N98, N165, N68);
and AND4 (N169, N81, N6, N96, N93);
or OR3 (N170, N168, N135, N22);
not NOT1 (N171, N156);
not NOT1 (N172, N150);
or OR3 (N173, N164, N30, N158);
and AND3 (N174, N173, N14, N33);
buf BUF1 (N175, N171);
not NOT1 (N176, N155);
nor NOR2 (N177, N169, N92);
or OR2 (N178, N149, N143);
buf BUF1 (N179, N175);
xor XOR2 (N180, N172, N40);
buf BUF1 (N181, N174);
nand NAND2 (N182, N153, N153);
not NOT1 (N183, N179);
xor XOR2 (N184, N181, N103);
and AND2 (N185, N176, N36);
not NOT1 (N186, N178);
nand NAND3 (N187, N184, N123, N22);
nand NAND4 (N188, N170, N186, N134, N46);
not NOT1 (N189, N168);
not NOT1 (N190, N189);
xor XOR2 (N191, N182, N131);
nand NAND4 (N192, N187, N169, N9, N160);
buf BUF1 (N193, N163);
or OR3 (N194, N183, N114, N48);
nand NAND4 (N195, N194, N111, N96, N35);
nor NOR4 (N196, N188, N9, N164, N192);
buf BUF1 (N197, N1);
buf BUF1 (N198, N197);
not NOT1 (N199, N180);
nand NAND2 (N200, N196, N84);
xor XOR2 (N201, N166, N23);
not NOT1 (N202, N185);
nor NOR2 (N203, N199, N23);
nand NAND4 (N204, N191, N93, N55, N150);
buf BUF1 (N205, N201);
or OR4 (N206, N204, N107, N3, N22);
not NOT1 (N207, N190);
buf BUF1 (N208, N195);
and AND4 (N209, N206, N146, N121, N165);
or OR2 (N210, N202, N170);
buf BUF1 (N211, N209);
nand NAND4 (N212, N208, N81, N31, N152);
xor XOR2 (N213, N207, N93);
nor NOR3 (N214, N198, N77, N85);
not NOT1 (N215, N203);
nor NOR3 (N216, N193, N130, N43);
nand NAND4 (N217, N211, N157, N140, N33);
nand NAND4 (N218, N215, N130, N169, N63);
buf BUF1 (N219, N212);
or OR3 (N220, N210, N213, N47);
xor XOR2 (N221, N146, N18);
not NOT1 (N222, N220);
or OR3 (N223, N218, N116, N17);
buf BUF1 (N224, N222);
not NOT1 (N225, N224);
and AND4 (N226, N177, N128, N112, N58);
buf BUF1 (N227, N221);
nor NOR2 (N228, N200, N108);
buf BUF1 (N229, N225);
buf BUF1 (N230, N216);
nor NOR3 (N231, N230, N201, N167);
nor NOR3 (N232, N226, N222, N140);
nor NOR2 (N233, N223, N34);
not NOT1 (N234, N228);
nand NAND4 (N235, N205, N107, N12, N34);
nand NAND2 (N236, N235, N192);
not NOT1 (N237, N234);
or OR2 (N238, N233, N189);
buf BUF1 (N239, N214);
xor XOR2 (N240, N219, N173);
and AND4 (N241, N232, N58, N223, N18);
xor XOR2 (N242, N238, N165);
nand NAND3 (N243, N237, N11, N59);
buf BUF1 (N244, N242);
buf BUF1 (N245, N227);
buf BUF1 (N246, N239);
or OR4 (N247, N245, N15, N41, N100);
buf BUF1 (N248, N236);
or OR3 (N249, N244, N100, N177);
or OR2 (N250, N248, N205);
and AND2 (N251, N243, N138);
and AND4 (N252, N250, N71, N244, N218);
nand NAND2 (N253, N240, N55);
nor NOR4 (N254, N249, N68, N168, N184);
or OR4 (N255, N246, N100, N81, N20);
nor NOR4 (N256, N253, N22, N199, N10);
xor XOR2 (N257, N256, N67);
xor XOR2 (N258, N217, N154);
nor NOR4 (N259, N254, N123, N71, N44);
nor NOR3 (N260, N229, N182, N34);
buf BUF1 (N261, N252);
not NOT1 (N262, N259);
nand NAND2 (N263, N241, N117);
buf BUF1 (N264, N260);
buf BUF1 (N265, N258);
not NOT1 (N266, N264);
xor XOR2 (N267, N247, N97);
and AND2 (N268, N261, N10);
or OR2 (N269, N251, N34);
xor XOR2 (N270, N267, N140);
or OR4 (N271, N255, N215, N137, N151);
buf BUF1 (N272, N266);
or OR2 (N273, N263, N140);
nand NAND3 (N274, N265, N163, N272);
and AND2 (N275, N237, N267);
nor NOR3 (N276, N274, N124, N242);
nor NOR3 (N277, N271, N141, N72);
xor XOR2 (N278, N273, N163);
not NOT1 (N279, N270);
and AND4 (N280, N268, N126, N196, N218);
xor XOR2 (N281, N257, N204);
xor XOR2 (N282, N279, N187);
or OR2 (N283, N269, N105);
nor NOR4 (N284, N277, N76, N195, N2);
nor NOR3 (N285, N283, N272, N123);
buf BUF1 (N286, N262);
xor XOR2 (N287, N231, N177);
and AND2 (N288, N284, N221);
not NOT1 (N289, N275);
and AND2 (N290, N281, N69);
and AND3 (N291, N287, N125, N140);
not NOT1 (N292, N288);
xor XOR2 (N293, N278, N201);
nand NAND4 (N294, N282, N87, N18, N200);
not NOT1 (N295, N294);
not NOT1 (N296, N293);
nor NOR4 (N297, N296, N132, N32, N20);
buf BUF1 (N298, N292);
and AND3 (N299, N291, N223, N252);
nand NAND4 (N300, N297, N295, N121, N102);
nor NOR4 (N301, N270, N5, N191, N18);
xor XOR2 (N302, N298, N125);
buf BUF1 (N303, N301);
not NOT1 (N304, N280);
buf BUF1 (N305, N286);
nand NAND2 (N306, N302, N301);
xor XOR2 (N307, N299, N128);
buf BUF1 (N308, N290);
buf BUF1 (N309, N285);
or OR3 (N310, N289, N35, N266);
or OR4 (N311, N307, N110, N102, N163);
xor XOR2 (N312, N304, N111);
or OR4 (N313, N309, N191, N72, N290);
buf BUF1 (N314, N300);
xor XOR2 (N315, N310, N231);
and AND3 (N316, N311, N281, N112);
and AND2 (N317, N312, N150);
and AND3 (N318, N303, N255, N129);
buf BUF1 (N319, N306);
xor XOR2 (N320, N305, N87);
nand NAND3 (N321, N319, N244, N300);
nand NAND3 (N322, N317, N86, N240);
nand NAND2 (N323, N308, N219);
nor NOR4 (N324, N313, N167, N122, N312);
or OR4 (N325, N318, N116, N43, N308);
not NOT1 (N326, N320);
buf BUF1 (N327, N314);
nor NOR2 (N328, N276, N322);
or OR4 (N329, N14, N134, N314, N275);
not NOT1 (N330, N315);
nor NOR2 (N331, N327, N325);
not NOT1 (N332, N185);
xor XOR2 (N333, N321, N228);
xor XOR2 (N334, N323, N72);
nor NOR2 (N335, N332, N204);
buf BUF1 (N336, N331);
and AND2 (N337, N324, N270);
buf BUF1 (N338, N335);
not NOT1 (N339, N316);
nand NAND2 (N340, N337, N143);
and AND4 (N341, N333, N151, N147, N281);
and AND2 (N342, N339, N111);
nor NOR4 (N343, N338, N232, N144, N187);
buf BUF1 (N344, N341);
not NOT1 (N345, N328);
or OR2 (N346, N340, N62);
and AND4 (N347, N330, N61, N121, N114);
not NOT1 (N348, N344);
not NOT1 (N349, N342);
and AND3 (N350, N334, N332, N88);
or OR2 (N351, N350, N304);
buf BUF1 (N352, N351);
nand NAND4 (N353, N349, N242, N333, N254);
and AND4 (N354, N346, N176, N116, N270);
nand NAND4 (N355, N354, N302, N13, N181);
nor NOR2 (N356, N352, N135);
buf BUF1 (N357, N336);
not NOT1 (N358, N329);
not NOT1 (N359, N345);
or OR2 (N360, N353, N48);
xor XOR2 (N361, N326, N124);
and AND2 (N362, N356, N237);
buf BUF1 (N363, N361);
and AND3 (N364, N347, N228, N299);
nor NOR2 (N365, N348, N191);
nor NOR3 (N366, N357, N161, N280);
nand NAND3 (N367, N365, N243, N298);
xor XOR2 (N368, N358, N196);
xor XOR2 (N369, N366, N333);
or OR3 (N370, N360, N104, N210);
not NOT1 (N371, N370);
nor NOR2 (N372, N362, N232);
nor NOR3 (N373, N364, N72, N151);
nand NAND3 (N374, N343, N207, N132);
nor NOR2 (N375, N368, N116);
buf BUF1 (N376, N372);
and AND3 (N377, N371, N33, N351);
nand NAND3 (N378, N374, N136, N175);
or OR3 (N379, N375, N353, N351);
and AND4 (N380, N373, N43, N237, N368);
nand NAND2 (N381, N369, N207);
or OR4 (N382, N380, N210, N366, N6);
nand NAND4 (N383, N359, N105, N126, N87);
buf BUF1 (N384, N379);
and AND4 (N385, N377, N66, N122, N277);
and AND4 (N386, N385, N78, N82, N255);
nand NAND2 (N387, N355, N365);
or OR3 (N388, N381, N350, N275);
nor NOR4 (N389, N384, N328, N258, N247);
or OR3 (N390, N363, N280, N13);
and AND3 (N391, N378, N257, N311);
nand NAND3 (N392, N387, N272, N72);
buf BUF1 (N393, N383);
and AND4 (N394, N393, N350, N240, N119);
not NOT1 (N395, N390);
xor XOR2 (N396, N382, N241);
and AND4 (N397, N367, N322, N184, N171);
not NOT1 (N398, N389);
nand NAND2 (N399, N394, N89);
and AND3 (N400, N396, N378, N22);
buf BUF1 (N401, N399);
nor NOR4 (N402, N388, N25, N244, N337);
xor XOR2 (N403, N386, N352);
nor NOR4 (N404, N398, N334, N84, N332);
nand NAND3 (N405, N392, N390, N234);
xor XOR2 (N406, N404, N11);
xor XOR2 (N407, N405, N35);
and AND2 (N408, N403, N73);
nand NAND4 (N409, N408, N319, N34, N106);
not NOT1 (N410, N401);
nor NOR3 (N411, N400, N293, N240);
or OR2 (N412, N395, N321);
nor NOR3 (N413, N406, N145, N145);
not NOT1 (N414, N409);
nor NOR4 (N415, N376, N358, N126, N44);
nor NOR3 (N416, N411, N63, N313);
not NOT1 (N417, N415);
nand NAND2 (N418, N397, N253);
xor XOR2 (N419, N407, N281);
xor XOR2 (N420, N416, N237);
nor NOR2 (N421, N419, N261);
and AND3 (N422, N414, N40, N352);
nor NOR3 (N423, N420, N44, N366);
and AND3 (N424, N423, N61, N364);
not NOT1 (N425, N424);
not NOT1 (N426, N421);
not NOT1 (N427, N413);
buf BUF1 (N428, N422);
not NOT1 (N429, N418);
nand NAND2 (N430, N429, N231);
xor XOR2 (N431, N402, N256);
nor NOR2 (N432, N426, N137);
not NOT1 (N433, N427);
buf BUF1 (N434, N410);
nor NOR4 (N435, N428, N415, N83, N204);
buf BUF1 (N436, N412);
or OR4 (N437, N435, N347, N405, N121);
or OR2 (N438, N432, N135);
and AND4 (N439, N417, N271, N32, N110);
buf BUF1 (N440, N437);
not NOT1 (N441, N436);
xor XOR2 (N442, N439, N371);
nand NAND3 (N443, N441, N411, N318);
xor XOR2 (N444, N430, N222);
nor NOR3 (N445, N440, N176, N99);
xor XOR2 (N446, N431, N338);
xor XOR2 (N447, N434, N350);
nor NOR2 (N448, N442, N404);
nand NAND2 (N449, N425, N417);
and AND3 (N450, N446, N81, N37);
or OR4 (N451, N443, N136, N4, N198);
xor XOR2 (N452, N449, N212);
nand NAND2 (N453, N444, N446);
or OR4 (N454, N447, N398, N226, N296);
buf BUF1 (N455, N433);
nand NAND2 (N456, N455, N409);
buf BUF1 (N457, N456);
nor NOR2 (N458, N457, N315);
not NOT1 (N459, N448);
and AND2 (N460, N451, N276);
nor NOR2 (N461, N454, N256);
buf BUF1 (N462, N452);
nor NOR2 (N463, N438, N309);
buf BUF1 (N464, N461);
nor NOR2 (N465, N445, N67);
or OR2 (N466, N450, N232);
not NOT1 (N467, N460);
nor NOR3 (N468, N462, N352, N453);
buf BUF1 (N469, N275);
not NOT1 (N470, N464);
nor NOR2 (N471, N391, N37);
and AND4 (N472, N463, N170, N332, N236);
not NOT1 (N473, N459);
xor XOR2 (N474, N469, N178);
xor XOR2 (N475, N458, N145);
or OR3 (N476, N468, N175, N233);
xor XOR2 (N477, N467, N36);
or OR3 (N478, N473, N431, N41);
and AND3 (N479, N472, N311, N247);
not NOT1 (N480, N471);
nor NOR3 (N481, N479, N19, N17);
not NOT1 (N482, N465);
buf BUF1 (N483, N477);
buf BUF1 (N484, N466);
or OR3 (N485, N478, N28, N174);
nor NOR3 (N486, N480, N343, N264);
or OR2 (N487, N474, N425);
not NOT1 (N488, N487);
nand NAND2 (N489, N483, N486);
xor XOR2 (N490, N153, N79);
nor NOR3 (N491, N470, N361, N169);
or OR4 (N492, N481, N124, N27, N246);
nand NAND4 (N493, N485, N284, N327, N143);
nand NAND4 (N494, N492, N44, N138, N459);
buf BUF1 (N495, N482);
nor NOR2 (N496, N484, N409);
nand NAND2 (N497, N493, N279);
xor XOR2 (N498, N476, N257);
or OR2 (N499, N494, N19);
xor XOR2 (N500, N491, N11);
buf BUF1 (N501, N500);
xor XOR2 (N502, N499, N124);
not NOT1 (N503, N496);
buf BUF1 (N504, N503);
not NOT1 (N505, N498);
or OR2 (N506, N495, N319);
and AND2 (N507, N502, N392);
nand NAND3 (N508, N507, N25, N3);
buf BUF1 (N509, N504);
or OR2 (N510, N508, N182);
nand NAND2 (N511, N506, N208);
nor NOR3 (N512, N488, N229, N199);
not NOT1 (N513, N475);
nor NOR2 (N514, N510, N323);
not NOT1 (N515, N511);
nor NOR2 (N516, N489, N348);
xor XOR2 (N517, N497, N510);
or OR4 (N518, N490, N382, N402, N283);
and AND4 (N519, N517, N314, N488, N278);
nor NOR2 (N520, N513, N277);
nor NOR3 (N521, N518, N508, N160);
and AND3 (N522, N509, N365, N226);
nand NAND4 (N523, N514, N290, N160, N448);
and AND2 (N524, N522, N418);
or OR2 (N525, N524, N12);
not NOT1 (N526, N525);
nand NAND3 (N527, N515, N201, N132);
buf BUF1 (N528, N512);
xor XOR2 (N529, N519, N347);
not NOT1 (N530, N523);
buf BUF1 (N531, N527);
nor NOR2 (N532, N530, N203);
xor XOR2 (N533, N531, N134);
and AND3 (N534, N520, N265, N278);
xor XOR2 (N535, N532, N194);
nor NOR4 (N536, N516, N404, N513, N254);
nor NOR4 (N537, N535, N205, N22, N312);
not NOT1 (N538, N528);
nand NAND3 (N539, N538, N313, N95);
or OR4 (N540, N505, N535, N76, N43);
xor XOR2 (N541, N521, N339);
not NOT1 (N542, N501);
nand NAND2 (N543, N539, N496);
or OR2 (N544, N540, N350);
not NOT1 (N545, N533);
nor NOR3 (N546, N542, N62, N444);
nor NOR2 (N547, N534, N518);
and AND2 (N548, N546, N243);
nand NAND2 (N549, N537, N67);
and AND3 (N550, N547, N384, N466);
xor XOR2 (N551, N549, N185);
nand NAND3 (N552, N526, N376, N122);
buf BUF1 (N553, N541);
and AND2 (N554, N545, N111);
or OR2 (N555, N551, N439);
or OR4 (N556, N552, N235, N190, N265);
buf BUF1 (N557, N543);
not NOT1 (N558, N550);
nand NAND4 (N559, N555, N496, N45, N184);
or OR3 (N560, N548, N415, N117);
or OR3 (N561, N553, N263, N85);
nor NOR3 (N562, N561, N234, N60);
nand NAND3 (N563, N529, N517, N189);
and AND4 (N564, N560, N173, N357, N159);
and AND4 (N565, N554, N103, N541, N76);
not NOT1 (N566, N564);
buf BUF1 (N567, N559);
not NOT1 (N568, N536);
and AND4 (N569, N556, N276, N20, N429);
nand NAND4 (N570, N558, N297, N263, N38);
not NOT1 (N571, N568);
xor XOR2 (N572, N557, N510);
xor XOR2 (N573, N569, N377);
xor XOR2 (N574, N566, N473);
buf BUF1 (N575, N565);
buf BUF1 (N576, N571);
not NOT1 (N577, N563);
nand NAND2 (N578, N572, N464);
and AND3 (N579, N570, N25, N239);
or OR3 (N580, N576, N215, N301);
not NOT1 (N581, N573);
xor XOR2 (N582, N574, N191);
nand NAND2 (N583, N562, N525);
not NOT1 (N584, N579);
buf BUF1 (N585, N584);
xor XOR2 (N586, N567, N288);
and AND3 (N587, N586, N298, N287);
xor XOR2 (N588, N587, N95);
or OR2 (N589, N585, N226);
nor NOR3 (N590, N589, N537, N314);
and AND3 (N591, N580, N373, N214);
and AND4 (N592, N583, N439, N522, N267);
and AND2 (N593, N582, N77);
xor XOR2 (N594, N578, N24);
or OR4 (N595, N591, N343, N112, N137);
or OR3 (N596, N581, N548, N264);
nor NOR2 (N597, N588, N558);
xor XOR2 (N598, N544, N301);
buf BUF1 (N599, N598);
nand NAND2 (N600, N575, N370);
nand NAND3 (N601, N590, N402, N526);
not NOT1 (N602, N577);
nand NAND2 (N603, N596, N66);
and AND4 (N604, N601, N258, N371, N69);
nor NOR4 (N605, N597, N33, N331, N583);
not NOT1 (N606, N600);
nand NAND2 (N607, N594, N204);
buf BUF1 (N608, N602);
xor XOR2 (N609, N605, N244);
xor XOR2 (N610, N606, N51);
nand NAND4 (N611, N603, N188, N285, N604);
not NOT1 (N612, N363);
nor NOR3 (N613, N608, N304, N448);
xor XOR2 (N614, N599, N153);
buf BUF1 (N615, N610);
or OR4 (N616, N595, N26, N145, N44);
xor XOR2 (N617, N613, N240);
nand NAND4 (N618, N616, N347, N262, N115);
nand NAND2 (N619, N607, N376);
or OR4 (N620, N611, N484, N314, N320);
buf BUF1 (N621, N593);
not NOT1 (N622, N592);
nor NOR2 (N623, N618, N471);
and AND3 (N624, N617, N40, N129);
nor NOR3 (N625, N619, N502, N274);
buf BUF1 (N626, N609);
xor XOR2 (N627, N625, N360);
buf BUF1 (N628, N615);
and AND2 (N629, N623, N41);
nand NAND4 (N630, N628, N591, N379, N446);
nand NAND2 (N631, N629, N369);
not NOT1 (N632, N612);
nor NOR2 (N633, N622, N149);
buf BUF1 (N634, N621);
nand NAND3 (N635, N626, N25, N316);
xor XOR2 (N636, N630, N124);
and AND3 (N637, N632, N222, N188);
and AND4 (N638, N633, N72, N27, N454);
not NOT1 (N639, N636);
buf BUF1 (N640, N639);
buf BUF1 (N641, N614);
and AND3 (N642, N627, N327, N22);
nand NAND3 (N643, N635, N75, N449);
and AND4 (N644, N641, N568, N204, N416);
or OR3 (N645, N634, N377, N188);
xor XOR2 (N646, N637, N238);
not NOT1 (N647, N643);
nand NAND3 (N648, N642, N372, N321);
and AND3 (N649, N646, N239, N23);
xor XOR2 (N650, N624, N68);
buf BUF1 (N651, N650);
and AND4 (N652, N638, N195, N589, N257);
or OR3 (N653, N620, N167, N611);
xor XOR2 (N654, N652, N76);
not NOT1 (N655, N651);
nor NOR3 (N656, N645, N620, N423);
xor XOR2 (N657, N644, N475);
nand NAND2 (N658, N657, N390);
buf BUF1 (N659, N649);
buf BUF1 (N660, N653);
nor NOR4 (N661, N654, N474, N179, N271);
or OR2 (N662, N661, N199);
or OR3 (N663, N660, N155, N58);
not NOT1 (N664, N663);
or OR2 (N665, N648, N277);
xor XOR2 (N666, N659, N220);
nor NOR3 (N667, N664, N513, N272);
and AND3 (N668, N640, N229, N170);
xor XOR2 (N669, N631, N327);
nand NAND4 (N670, N662, N141, N523, N21);
buf BUF1 (N671, N658);
buf BUF1 (N672, N666);
nor NOR3 (N673, N647, N345, N492);
not NOT1 (N674, N668);
buf BUF1 (N675, N670);
buf BUF1 (N676, N665);
nor NOR4 (N677, N656, N373, N39, N116);
not NOT1 (N678, N675);
or OR2 (N679, N674, N486);
nand NAND2 (N680, N679, N631);
buf BUF1 (N681, N678);
buf BUF1 (N682, N681);
nor NOR4 (N683, N667, N620, N24, N266);
xor XOR2 (N684, N655, N288);
buf BUF1 (N685, N683);
not NOT1 (N686, N685);
and AND3 (N687, N672, N283, N75);
not NOT1 (N688, N676);
and AND3 (N689, N677, N40, N560);
nand NAND4 (N690, N687, N280, N218, N91);
buf BUF1 (N691, N689);
nand NAND4 (N692, N669, N64, N156, N494);
xor XOR2 (N693, N688, N493);
xor XOR2 (N694, N692, N561);
buf BUF1 (N695, N686);
buf BUF1 (N696, N694);
or OR2 (N697, N680, N70);
buf BUF1 (N698, N691);
buf BUF1 (N699, N690);
nand NAND2 (N700, N693, N569);
nand NAND4 (N701, N700, N272, N217, N342);
not NOT1 (N702, N695);
xor XOR2 (N703, N699, N149);
xor XOR2 (N704, N701, N516);
xor XOR2 (N705, N698, N58);
or OR3 (N706, N684, N622, N139);
xor XOR2 (N707, N671, N32);
and AND2 (N708, N707, N169);
not NOT1 (N709, N708);
nor NOR2 (N710, N704, N316);
or OR4 (N711, N710, N18, N436, N73);
not NOT1 (N712, N696);
nand NAND3 (N713, N697, N560, N75);
and AND4 (N714, N712, N300, N387, N445);
nor NOR2 (N715, N703, N321);
nor NOR4 (N716, N706, N21, N537, N88);
xor XOR2 (N717, N715, N418);
and AND4 (N718, N682, N281, N139, N287);
nand NAND4 (N719, N709, N164, N97, N373);
not NOT1 (N720, N714);
nor NOR3 (N721, N711, N576, N430);
buf BUF1 (N722, N705);
nor NOR4 (N723, N720, N124, N631, N598);
xor XOR2 (N724, N702, N462);
buf BUF1 (N725, N673);
xor XOR2 (N726, N713, N162);
or OR3 (N727, N717, N549, N567);
and AND3 (N728, N723, N43, N721);
and AND2 (N729, N397, N157);
not NOT1 (N730, N728);
nor NOR3 (N731, N730, N107, N698);
nor NOR2 (N732, N726, N430);
or OR3 (N733, N727, N361, N70);
nor NOR3 (N734, N729, N156, N132);
and AND2 (N735, N722, N547);
buf BUF1 (N736, N716);
not NOT1 (N737, N736);
not NOT1 (N738, N735);
nand NAND3 (N739, N734, N656, N672);
nor NOR2 (N740, N719, N197);
xor XOR2 (N741, N724, N693);
not NOT1 (N742, N718);
not NOT1 (N743, N731);
xor XOR2 (N744, N733, N165);
buf BUF1 (N745, N739);
not NOT1 (N746, N740);
xor XOR2 (N747, N742, N465);
nand NAND2 (N748, N725, N727);
and AND2 (N749, N738, N60);
nor NOR2 (N750, N743, N697);
nand NAND2 (N751, N737, N227);
not NOT1 (N752, N751);
buf BUF1 (N753, N741);
or OR4 (N754, N746, N733, N595, N282);
xor XOR2 (N755, N744, N476);
nand NAND4 (N756, N755, N322, N426, N200);
buf BUF1 (N757, N749);
or OR3 (N758, N745, N172, N526);
nor NOR3 (N759, N747, N83, N353);
or OR2 (N760, N754, N498);
and AND2 (N761, N732, N397);
buf BUF1 (N762, N757);
and AND2 (N763, N750, N10);
xor XOR2 (N764, N756, N234);
nor NOR2 (N765, N759, N286);
buf BUF1 (N766, N764);
xor XOR2 (N767, N765, N382);
or OR4 (N768, N763, N520, N268, N662);
nor NOR2 (N769, N761, N473);
not NOT1 (N770, N752);
or OR4 (N771, N769, N493, N37, N747);
xor XOR2 (N772, N753, N165);
xor XOR2 (N773, N768, N7);
nand NAND3 (N774, N762, N701, N49);
or OR3 (N775, N773, N627, N463);
not NOT1 (N776, N767);
and AND4 (N777, N766, N327, N519, N54);
or OR4 (N778, N774, N19, N269, N339);
nor NOR2 (N779, N770, N528);
and AND4 (N780, N778, N173, N553, N322);
or OR3 (N781, N777, N695, N233);
and AND4 (N782, N780, N18, N769, N381);
not NOT1 (N783, N771);
not NOT1 (N784, N748);
buf BUF1 (N785, N784);
xor XOR2 (N786, N772, N414);
or OR2 (N787, N781, N315);
and AND4 (N788, N760, N260, N320, N549);
or OR3 (N789, N779, N467, N320);
not NOT1 (N790, N782);
buf BUF1 (N791, N758);
nor NOR2 (N792, N776, N590);
buf BUF1 (N793, N775);
nor NOR2 (N794, N783, N337);
nand NAND2 (N795, N786, N760);
or OR3 (N796, N793, N101, N658);
and AND2 (N797, N787, N568);
and AND3 (N798, N796, N333, N42);
buf BUF1 (N799, N788);
xor XOR2 (N800, N791, N626);
and AND2 (N801, N794, N156);
nor NOR3 (N802, N799, N666, N90);
xor XOR2 (N803, N792, N767);
or OR2 (N804, N785, N104);
nor NOR4 (N805, N790, N491, N177, N140);
nor NOR3 (N806, N797, N761, N4);
buf BUF1 (N807, N798);
buf BUF1 (N808, N801);
or OR3 (N809, N805, N32, N756);
and AND3 (N810, N809, N154, N67);
buf BUF1 (N811, N807);
nand NAND3 (N812, N804, N186, N499);
nand NAND2 (N813, N810, N344);
nand NAND4 (N814, N800, N46, N72, N254);
nand NAND4 (N815, N802, N581, N247, N149);
buf BUF1 (N816, N815);
nor NOR4 (N817, N808, N600, N172, N390);
xor XOR2 (N818, N789, N223);
or OR3 (N819, N812, N622, N130);
or OR3 (N820, N813, N27, N652);
buf BUF1 (N821, N818);
nor NOR4 (N822, N817, N591, N778, N54);
and AND3 (N823, N795, N732, N588);
and AND4 (N824, N820, N664, N429, N765);
nand NAND4 (N825, N814, N58, N34, N366);
xor XOR2 (N826, N811, N679);
or OR2 (N827, N819, N556);
buf BUF1 (N828, N824);
buf BUF1 (N829, N823);
xor XOR2 (N830, N826, N361);
and AND2 (N831, N825, N352);
and AND4 (N832, N816, N409, N590, N645);
nor NOR3 (N833, N829, N292, N157);
nor NOR3 (N834, N803, N288, N481);
xor XOR2 (N835, N831, N282);
nor NOR2 (N836, N833, N667);
nand NAND2 (N837, N832, N572);
or OR3 (N838, N806, N156, N491);
nor NOR2 (N839, N821, N72);
or OR2 (N840, N837, N458);
nor NOR4 (N841, N834, N51, N100, N705);
nor NOR4 (N842, N838, N595, N781, N632);
or OR4 (N843, N827, N27, N433, N823);
buf BUF1 (N844, N840);
nor NOR3 (N845, N822, N289, N536);
xor XOR2 (N846, N844, N551);
xor XOR2 (N847, N830, N305);
or OR4 (N848, N847, N226, N23, N797);
not NOT1 (N849, N846);
not NOT1 (N850, N839);
not NOT1 (N851, N843);
or OR2 (N852, N828, N267);
and AND4 (N853, N835, N308, N134, N254);
not NOT1 (N854, N848);
nor NOR3 (N855, N850, N519, N630);
not NOT1 (N856, N853);
nor NOR2 (N857, N836, N477);
and AND3 (N858, N851, N230, N723);
not NOT1 (N859, N857);
nand NAND4 (N860, N842, N349, N89, N742);
or OR2 (N861, N841, N68);
or OR3 (N862, N852, N178, N807);
xor XOR2 (N863, N849, N762);
buf BUF1 (N864, N859);
and AND3 (N865, N862, N160, N704);
xor XOR2 (N866, N856, N751);
buf BUF1 (N867, N863);
not NOT1 (N868, N864);
and AND3 (N869, N845, N184, N800);
nand NAND4 (N870, N866, N672, N30, N75);
nand NAND4 (N871, N867, N208, N803, N504);
or OR2 (N872, N855, N86);
and AND3 (N873, N865, N569, N417);
xor XOR2 (N874, N868, N518);
and AND2 (N875, N872, N363);
buf BUF1 (N876, N858);
and AND3 (N877, N875, N314, N571);
nand NAND3 (N878, N869, N507, N485);
buf BUF1 (N879, N870);
or OR4 (N880, N878, N820, N773, N361);
buf BUF1 (N881, N874);
or OR4 (N882, N881, N515, N79, N250);
or OR3 (N883, N860, N25, N290);
or OR2 (N884, N882, N559);
buf BUF1 (N885, N884);
or OR3 (N886, N861, N832, N664);
nor NOR2 (N887, N880, N736);
buf BUF1 (N888, N877);
xor XOR2 (N889, N879, N646);
and AND2 (N890, N887, N7);
buf BUF1 (N891, N871);
and AND2 (N892, N889, N270);
nand NAND4 (N893, N885, N643, N728, N678);
nor NOR2 (N894, N873, N457);
nor NOR2 (N895, N854, N409);
nand NAND2 (N896, N892, N284);
or OR2 (N897, N888, N887);
and AND4 (N898, N893, N220, N739, N880);
not NOT1 (N899, N891);
nor NOR3 (N900, N886, N449, N549);
buf BUF1 (N901, N898);
xor XOR2 (N902, N900, N826);
nand NAND4 (N903, N899, N543, N414, N118);
buf BUF1 (N904, N895);
and AND4 (N905, N903, N179, N253, N677);
and AND2 (N906, N897, N858);
nand NAND3 (N907, N906, N378, N253);
and AND4 (N908, N890, N567, N862, N276);
buf BUF1 (N909, N904);
nand NAND4 (N910, N901, N354, N265, N246);
xor XOR2 (N911, N902, N517);
or OR3 (N912, N907, N630, N258);
endmodule