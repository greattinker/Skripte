// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N611,N604,N610,N607,N616,N615,N613,N609,N594,N617;

or OR4 (N18, N7, N1, N10, N13);
buf BUF1 (N19, N6);
nor NOR3 (N20, N1, N13, N14);
buf BUF1 (N21, N17);
not NOT1 (N22, N1);
and AND3 (N23, N18, N12, N22);
xor XOR2 (N24, N13, N13);
and AND3 (N25, N9, N23, N20);
xor XOR2 (N26, N1, N25);
or OR4 (N27, N20, N13, N12, N8);
or OR2 (N28, N1, N13);
and AND2 (N29, N14, N7);
not NOT1 (N30, N15);
not NOT1 (N31, N12);
xor XOR2 (N32, N28, N22);
buf BUF1 (N33, N19);
xor XOR2 (N34, N13, N7);
and AND3 (N35, N21, N29, N32);
not NOT1 (N36, N32);
xor XOR2 (N37, N35, N19);
not NOT1 (N38, N31);
nand NAND2 (N39, N19, N4);
and AND2 (N40, N38, N1);
or OR3 (N41, N39, N36, N38);
buf BUF1 (N42, N17);
not NOT1 (N43, N42);
not NOT1 (N44, N37);
or OR4 (N45, N30, N27, N16, N21);
nand NAND2 (N46, N22, N17);
and AND3 (N47, N34, N32, N8);
xor XOR2 (N48, N40, N5);
nor NOR4 (N49, N48, N6, N12, N17);
nand NAND3 (N50, N45, N31, N11);
nor NOR2 (N51, N44, N33);
nor NOR3 (N52, N51, N27, N50);
or OR3 (N53, N24, N14, N1);
nand NAND3 (N54, N25, N15, N7);
buf BUF1 (N55, N52);
buf BUF1 (N56, N34);
or OR4 (N57, N46, N1, N22, N47);
buf BUF1 (N58, N22);
buf BUF1 (N59, N26);
xor XOR2 (N60, N53, N52);
nand NAND2 (N61, N43, N37);
nand NAND2 (N62, N54, N8);
buf BUF1 (N63, N49);
or OR3 (N64, N55, N28, N5);
nor NOR4 (N65, N41, N1, N21, N3);
nor NOR4 (N66, N63, N48, N4, N40);
and AND3 (N67, N57, N53, N24);
xor XOR2 (N68, N58, N10);
buf BUF1 (N69, N64);
xor XOR2 (N70, N59, N21);
and AND4 (N71, N66, N8, N8, N43);
nand NAND2 (N72, N60, N49);
xor XOR2 (N73, N65, N69);
or OR3 (N74, N40, N73, N42);
nand NAND4 (N75, N51, N3, N28, N2);
nand NAND3 (N76, N62, N61, N37);
not NOT1 (N77, N54);
xor XOR2 (N78, N76, N29);
or OR2 (N79, N68, N55);
and AND4 (N80, N56, N79, N42, N43);
buf BUF1 (N81, N55);
nand NAND2 (N82, N75, N38);
xor XOR2 (N83, N67, N51);
and AND4 (N84, N81, N46, N29, N63);
or OR4 (N85, N72, N51, N36, N52);
not NOT1 (N86, N82);
nand NAND3 (N87, N83, N60, N34);
nand NAND4 (N88, N85, N46, N59, N23);
and AND2 (N89, N86, N5);
and AND4 (N90, N70, N84, N23, N58);
xor XOR2 (N91, N2, N84);
buf BUF1 (N92, N89);
and AND4 (N93, N74, N8, N73, N37);
nor NOR2 (N94, N92, N21);
or OR4 (N95, N90, N12, N40, N40);
nor NOR3 (N96, N77, N62, N63);
nor NOR3 (N97, N80, N2, N7);
or OR3 (N98, N78, N81, N16);
nor NOR2 (N99, N91, N68);
and AND4 (N100, N71, N8, N37, N8);
xor XOR2 (N101, N96, N6);
buf BUF1 (N102, N97);
buf BUF1 (N103, N101);
not NOT1 (N104, N102);
or OR4 (N105, N94, N13, N52, N104);
not NOT1 (N106, N86);
not NOT1 (N107, N103);
or OR2 (N108, N100, N28);
buf BUF1 (N109, N98);
xor XOR2 (N110, N107, N26);
and AND3 (N111, N106, N105, N69);
not NOT1 (N112, N11);
and AND2 (N113, N95, N55);
nand NAND2 (N114, N110, N21);
or OR3 (N115, N99, N77, N33);
not NOT1 (N116, N108);
nor NOR3 (N117, N113, N37, N83);
nand NAND2 (N118, N115, N65);
not NOT1 (N119, N109);
nor NOR3 (N120, N87, N80, N13);
xor XOR2 (N121, N119, N113);
buf BUF1 (N122, N114);
nand NAND4 (N123, N121, N95, N45, N21);
buf BUF1 (N124, N120);
or OR4 (N125, N122, N54, N56, N90);
or OR4 (N126, N118, N8, N6, N10);
buf BUF1 (N127, N124);
xor XOR2 (N128, N123, N95);
buf BUF1 (N129, N111);
buf BUF1 (N130, N88);
nand NAND3 (N131, N125, N5, N15);
or OR3 (N132, N128, N120, N84);
nand NAND3 (N133, N117, N102, N25);
nor NOR2 (N134, N93, N131);
xor XOR2 (N135, N113, N85);
nor NOR4 (N136, N129, N113, N78, N14);
nand NAND4 (N137, N133, N80, N73, N108);
buf BUF1 (N138, N126);
not NOT1 (N139, N135);
not NOT1 (N140, N139);
buf BUF1 (N141, N140);
and AND3 (N142, N132, N107, N125);
or OR4 (N143, N134, N85, N120, N133);
or OR4 (N144, N142, N60, N74, N11);
or OR2 (N145, N127, N100);
nand NAND4 (N146, N145, N9, N2, N138);
nor NOR2 (N147, N57, N70);
buf BUF1 (N148, N147);
or OR4 (N149, N144, N70, N138, N52);
buf BUF1 (N150, N136);
and AND3 (N151, N149, N84, N121);
nor NOR3 (N152, N148, N61, N77);
xor XOR2 (N153, N116, N68);
or OR2 (N154, N150, N111);
xor XOR2 (N155, N152, N75);
buf BUF1 (N156, N154);
buf BUF1 (N157, N141);
xor XOR2 (N158, N157, N76);
xor XOR2 (N159, N155, N147);
not NOT1 (N160, N143);
nand NAND3 (N161, N112, N60, N28);
nand NAND3 (N162, N158, N114, N97);
buf BUF1 (N163, N160);
or OR4 (N164, N151, N93, N40, N157);
nand NAND4 (N165, N156, N154, N144, N128);
buf BUF1 (N166, N161);
and AND4 (N167, N146, N89, N73, N75);
or OR4 (N168, N164, N106, N107, N154);
not NOT1 (N169, N159);
or OR3 (N170, N165, N163, N67);
not NOT1 (N171, N10);
nand NAND3 (N172, N170, N71, N12);
xor XOR2 (N173, N153, N67);
xor XOR2 (N174, N167, N1);
xor XOR2 (N175, N172, N15);
or OR2 (N176, N168, N44);
and AND4 (N177, N174, N104, N60, N173);
buf BUF1 (N178, N149);
nor NOR4 (N179, N175, N30, N82, N89);
xor XOR2 (N180, N162, N63);
not NOT1 (N181, N176);
xor XOR2 (N182, N137, N39);
xor XOR2 (N183, N178, N93);
or OR3 (N184, N181, N139, N88);
not NOT1 (N185, N130);
and AND2 (N186, N183, N24);
or OR3 (N187, N186, N185, N32);
or OR2 (N188, N59, N112);
not NOT1 (N189, N179);
buf BUF1 (N190, N171);
nor NOR2 (N191, N166, N134);
not NOT1 (N192, N188);
buf BUF1 (N193, N190);
buf BUF1 (N194, N169);
or OR3 (N195, N194, N32, N129);
or OR2 (N196, N191, N50);
buf BUF1 (N197, N182);
buf BUF1 (N198, N177);
buf BUF1 (N199, N192);
or OR3 (N200, N196, N108, N144);
nand NAND3 (N201, N199, N100, N63);
xor XOR2 (N202, N200, N40);
not NOT1 (N203, N184);
nand NAND3 (N204, N203, N101, N13);
buf BUF1 (N205, N193);
or OR3 (N206, N198, N13, N41);
not NOT1 (N207, N197);
xor XOR2 (N208, N207, N54);
xor XOR2 (N209, N204, N99);
buf BUF1 (N210, N189);
or OR4 (N211, N208, N56, N33, N90);
and AND3 (N212, N201, N5, N86);
and AND2 (N213, N205, N89);
nor NOR3 (N214, N187, N52, N178);
or OR2 (N215, N213, N14);
not NOT1 (N216, N195);
nor NOR2 (N217, N215, N12);
not NOT1 (N218, N216);
nor NOR3 (N219, N210, N150, N173);
not NOT1 (N220, N212);
or OR4 (N221, N218, N145, N116, N7);
nor NOR2 (N222, N221, N111);
nor NOR2 (N223, N206, N133);
not NOT1 (N224, N222);
buf BUF1 (N225, N217);
not NOT1 (N226, N211);
nor NOR4 (N227, N202, N31, N50, N41);
buf BUF1 (N228, N224);
and AND2 (N229, N223, N87);
xor XOR2 (N230, N220, N180);
xor XOR2 (N231, N106, N71);
xor XOR2 (N232, N209, N37);
or OR3 (N233, N229, N224, N167);
not NOT1 (N234, N226);
or OR3 (N235, N214, N7, N207);
nor NOR4 (N236, N227, N135, N148, N221);
not NOT1 (N237, N225);
buf BUF1 (N238, N235);
or OR2 (N239, N232, N215);
xor XOR2 (N240, N219, N89);
and AND3 (N241, N231, N93, N103);
nand NAND4 (N242, N238, N116, N149, N30);
nand NAND3 (N243, N234, N133, N85);
nand NAND4 (N244, N230, N172, N18, N167);
or OR4 (N245, N233, N111, N91, N99);
nor NOR2 (N246, N239, N60);
not NOT1 (N247, N245);
nand NAND3 (N248, N228, N5, N149);
nor NOR4 (N249, N236, N85, N46, N89);
buf BUF1 (N250, N247);
nand NAND2 (N251, N249, N8);
nand NAND4 (N252, N242, N235, N225, N244);
xor XOR2 (N253, N219, N245);
or OR2 (N254, N250, N152);
buf BUF1 (N255, N248);
nor NOR3 (N256, N253, N27, N214);
nand NAND2 (N257, N251, N127);
nand NAND3 (N258, N246, N193, N160);
and AND2 (N259, N254, N11);
nor NOR3 (N260, N256, N53, N61);
xor XOR2 (N261, N243, N114);
xor XOR2 (N262, N241, N200);
nand NAND2 (N263, N259, N215);
xor XOR2 (N264, N252, N109);
buf BUF1 (N265, N262);
and AND4 (N266, N255, N127, N188, N131);
and AND3 (N267, N258, N110, N171);
xor XOR2 (N268, N260, N215);
and AND4 (N269, N265, N163, N19, N88);
nand NAND2 (N270, N264, N63);
nand NAND4 (N271, N266, N227, N42, N2);
xor XOR2 (N272, N268, N175);
and AND2 (N273, N240, N145);
nor NOR2 (N274, N257, N54);
nor NOR3 (N275, N237, N219, N179);
xor XOR2 (N276, N261, N45);
buf BUF1 (N277, N269);
or OR3 (N278, N267, N223, N229);
xor XOR2 (N279, N263, N235);
nand NAND3 (N280, N276, N205, N243);
not NOT1 (N281, N274);
buf BUF1 (N282, N273);
xor XOR2 (N283, N277, N19);
not NOT1 (N284, N282);
xor XOR2 (N285, N283, N239);
xor XOR2 (N286, N279, N191);
not NOT1 (N287, N271);
nor NOR2 (N288, N270, N218);
not NOT1 (N289, N272);
nor NOR3 (N290, N281, N23, N72);
and AND2 (N291, N278, N165);
nor NOR3 (N292, N284, N234, N175);
or OR2 (N293, N280, N194);
xor XOR2 (N294, N292, N212);
not NOT1 (N295, N285);
xor XOR2 (N296, N287, N120);
nor NOR2 (N297, N275, N268);
not NOT1 (N298, N297);
buf BUF1 (N299, N288);
xor XOR2 (N300, N296, N112);
buf BUF1 (N301, N298);
xor XOR2 (N302, N294, N2);
not NOT1 (N303, N301);
nor NOR2 (N304, N295, N71);
or OR4 (N305, N303, N175, N191, N11);
nand NAND3 (N306, N305, N289, N11);
or OR2 (N307, N240, N75);
or OR2 (N308, N306, N200);
nor NOR3 (N309, N299, N34, N13);
nand NAND4 (N310, N291, N92, N209, N212);
or OR2 (N311, N300, N106);
buf BUF1 (N312, N310);
nand NAND4 (N313, N308, N68, N70, N117);
and AND3 (N314, N313, N302, N303);
and AND4 (N315, N35, N195, N313, N140);
not NOT1 (N316, N286);
nor NOR4 (N317, N290, N249, N277, N148);
xor XOR2 (N318, N311, N191);
nand NAND3 (N319, N293, N246, N173);
not NOT1 (N320, N307);
nor NOR3 (N321, N319, N31, N98);
xor XOR2 (N322, N315, N163);
not NOT1 (N323, N317);
buf BUF1 (N324, N314);
xor XOR2 (N325, N320, N290);
nor NOR4 (N326, N312, N12, N271, N303);
nor NOR3 (N327, N316, N97, N305);
buf BUF1 (N328, N321);
nor NOR2 (N329, N325, N193);
or OR4 (N330, N323, N210, N265, N250);
or OR4 (N331, N304, N99, N244, N161);
xor XOR2 (N332, N331, N2);
nor NOR3 (N333, N332, N309, N133);
or OR2 (N334, N91, N301);
not NOT1 (N335, N329);
xor XOR2 (N336, N328, N46);
nand NAND2 (N337, N335, N132);
and AND4 (N338, N326, N148, N207, N128);
not NOT1 (N339, N336);
nand NAND4 (N340, N322, N80, N205, N308);
or OR4 (N341, N324, N251, N332, N23);
and AND2 (N342, N318, N9);
or OR4 (N343, N342, N2, N80, N3);
nor NOR2 (N344, N343, N203);
and AND4 (N345, N337, N172, N39, N112);
and AND4 (N346, N340, N85, N292, N285);
not NOT1 (N347, N334);
and AND4 (N348, N344, N309, N335, N275);
nor NOR3 (N349, N327, N61, N118);
not NOT1 (N350, N330);
buf BUF1 (N351, N348);
nand NAND3 (N352, N339, N2, N185);
and AND4 (N353, N351, N17, N138, N5);
and AND4 (N354, N347, N178, N101, N339);
or OR2 (N355, N353, N324);
not NOT1 (N356, N346);
buf BUF1 (N357, N338);
nand NAND2 (N358, N356, N145);
not NOT1 (N359, N345);
not NOT1 (N360, N355);
nand NAND3 (N361, N352, N282, N303);
buf BUF1 (N362, N349);
and AND2 (N363, N358, N294);
not NOT1 (N364, N354);
not NOT1 (N365, N363);
buf BUF1 (N366, N360);
or OR3 (N367, N365, N118, N148);
nand NAND2 (N368, N341, N88);
or OR2 (N369, N357, N82);
not NOT1 (N370, N359);
xor XOR2 (N371, N333, N73);
xor XOR2 (N372, N369, N224);
nor NOR2 (N373, N350, N85);
buf BUF1 (N374, N362);
not NOT1 (N375, N361);
xor XOR2 (N376, N366, N339);
or OR2 (N377, N368, N10);
and AND4 (N378, N374, N307, N296, N197);
xor XOR2 (N379, N378, N323);
and AND4 (N380, N372, N364, N165, N193);
or OR4 (N381, N169, N78, N77, N61);
or OR2 (N382, N371, N81);
xor XOR2 (N383, N381, N98);
and AND2 (N384, N379, N203);
nand NAND2 (N385, N370, N284);
buf BUF1 (N386, N367);
not NOT1 (N387, N375);
nand NAND2 (N388, N377, N376);
not NOT1 (N389, N122);
nor NOR3 (N390, N386, N64, N259);
buf BUF1 (N391, N384);
and AND2 (N392, N380, N265);
nand NAND2 (N393, N382, N346);
nand NAND4 (N394, N392, N206, N319, N105);
not NOT1 (N395, N393);
buf BUF1 (N396, N388);
and AND4 (N397, N385, N128, N24, N2);
and AND2 (N398, N390, N231);
buf BUF1 (N399, N397);
buf BUF1 (N400, N389);
nand NAND3 (N401, N400, N102, N324);
or OR3 (N402, N373, N274, N32);
nand NAND2 (N403, N391, N219);
or OR2 (N404, N398, N158);
or OR3 (N405, N404, N308, N268);
nand NAND3 (N406, N403, N78, N125);
not NOT1 (N407, N394);
and AND2 (N408, N387, N73);
not NOT1 (N409, N408);
and AND4 (N410, N405, N42, N4, N295);
or OR3 (N411, N401, N212, N398);
nand NAND3 (N412, N407, N350, N37);
buf BUF1 (N413, N383);
not NOT1 (N414, N411);
nor NOR3 (N415, N409, N157, N173);
not NOT1 (N416, N414);
nand NAND4 (N417, N396, N166, N49, N250);
not NOT1 (N418, N415);
nand NAND4 (N419, N395, N329, N84, N385);
and AND2 (N420, N406, N207);
or OR3 (N421, N402, N283, N45);
or OR3 (N422, N417, N15, N383);
buf BUF1 (N423, N421);
and AND2 (N424, N416, N275);
not NOT1 (N425, N413);
or OR2 (N426, N412, N210);
xor XOR2 (N427, N423, N373);
buf BUF1 (N428, N424);
nand NAND4 (N429, N410, N82, N279, N94);
nand NAND3 (N430, N418, N268, N401);
buf BUF1 (N431, N422);
nand NAND3 (N432, N420, N137, N205);
not NOT1 (N433, N428);
xor XOR2 (N434, N399, N134);
or OR3 (N435, N430, N285, N104);
not NOT1 (N436, N432);
buf BUF1 (N437, N425);
nor NOR2 (N438, N427, N92);
not NOT1 (N439, N419);
not NOT1 (N440, N439);
buf BUF1 (N441, N440);
nand NAND2 (N442, N429, N316);
or OR3 (N443, N436, N69, N201);
nand NAND2 (N444, N438, N391);
xor XOR2 (N445, N444, N137);
nor NOR2 (N446, N445, N206);
nand NAND4 (N447, N433, N238, N64, N170);
or OR4 (N448, N431, N429, N324, N192);
buf BUF1 (N449, N434);
not NOT1 (N450, N448);
nor NOR3 (N451, N443, N397, N196);
and AND3 (N452, N426, N333, N397);
xor XOR2 (N453, N441, N338);
not NOT1 (N454, N453);
nor NOR4 (N455, N446, N153, N235, N400);
or OR4 (N456, N455, N76, N53, N222);
nor NOR2 (N457, N456, N221);
nor NOR2 (N458, N447, N396);
or OR3 (N459, N454, N445, N197);
nand NAND3 (N460, N450, N177, N337);
nand NAND2 (N461, N458, N313);
not NOT1 (N462, N435);
not NOT1 (N463, N459);
nand NAND2 (N464, N451, N439);
or OR3 (N465, N442, N147, N63);
xor XOR2 (N466, N464, N249);
xor XOR2 (N467, N452, N138);
or OR4 (N468, N449, N139, N348, N300);
and AND3 (N469, N465, N1, N134);
buf BUF1 (N470, N463);
nand NAND4 (N471, N468, N81, N325, N62);
and AND2 (N472, N469, N446);
not NOT1 (N473, N457);
nor NOR4 (N474, N470, N253, N356, N88);
buf BUF1 (N475, N461);
not NOT1 (N476, N472);
xor XOR2 (N477, N460, N231);
and AND3 (N478, N476, N61, N279);
or OR3 (N479, N473, N49, N260);
xor XOR2 (N480, N477, N155);
buf BUF1 (N481, N471);
not NOT1 (N482, N466);
xor XOR2 (N483, N474, N264);
xor XOR2 (N484, N478, N55);
nor NOR2 (N485, N467, N132);
nor NOR4 (N486, N485, N165, N3, N292);
or OR3 (N487, N475, N423, N436);
not NOT1 (N488, N482);
and AND2 (N489, N481, N64);
buf BUF1 (N490, N462);
buf BUF1 (N491, N483);
or OR4 (N492, N480, N38, N219, N153);
xor XOR2 (N493, N437, N480);
nor NOR3 (N494, N489, N102, N59);
buf BUF1 (N495, N494);
not NOT1 (N496, N484);
xor XOR2 (N497, N486, N472);
buf BUF1 (N498, N487);
xor XOR2 (N499, N479, N318);
xor XOR2 (N500, N497, N462);
xor XOR2 (N501, N491, N168);
or OR2 (N502, N500, N30);
xor XOR2 (N503, N492, N501);
nand NAND3 (N504, N407, N434, N274);
buf BUF1 (N505, N495);
xor XOR2 (N506, N499, N179);
nand NAND4 (N507, N493, N370, N363, N356);
xor XOR2 (N508, N496, N394);
xor XOR2 (N509, N502, N461);
xor XOR2 (N510, N503, N33);
nor NOR2 (N511, N507, N132);
nand NAND4 (N512, N511, N24, N69, N415);
not NOT1 (N513, N498);
or OR2 (N514, N509, N356);
xor XOR2 (N515, N490, N161);
buf BUF1 (N516, N506);
not NOT1 (N517, N513);
not NOT1 (N518, N517);
or OR3 (N519, N505, N325, N117);
buf BUF1 (N520, N508);
nand NAND3 (N521, N488, N373, N351);
or OR4 (N522, N521, N163, N223, N258);
xor XOR2 (N523, N519, N427);
xor XOR2 (N524, N523, N45);
not NOT1 (N525, N510);
xor XOR2 (N526, N504, N232);
nor NOR2 (N527, N518, N156);
xor XOR2 (N528, N514, N94);
not NOT1 (N529, N516);
buf BUF1 (N530, N528);
buf BUF1 (N531, N525);
nand NAND2 (N532, N530, N484);
and AND3 (N533, N527, N44, N414);
not NOT1 (N534, N522);
and AND4 (N535, N533, N392, N440, N38);
or OR4 (N536, N512, N339, N54, N367);
nand NAND3 (N537, N526, N219, N202);
buf BUF1 (N538, N536);
not NOT1 (N539, N535);
xor XOR2 (N540, N524, N141);
nor NOR2 (N541, N529, N242);
nand NAND4 (N542, N540, N370, N185, N32);
nor NOR4 (N543, N520, N344, N88, N203);
nand NAND4 (N544, N542, N112, N520, N80);
nor NOR4 (N545, N544, N4, N57, N510);
nand NAND2 (N546, N515, N99);
or OR3 (N547, N537, N201, N333);
and AND3 (N548, N546, N307, N132);
xor XOR2 (N549, N531, N442);
nor NOR4 (N550, N545, N266, N492, N379);
not NOT1 (N551, N534);
xor XOR2 (N552, N548, N371);
or OR2 (N553, N547, N425);
xor XOR2 (N554, N538, N472);
not NOT1 (N555, N553);
xor XOR2 (N556, N539, N496);
xor XOR2 (N557, N532, N361);
nor NOR2 (N558, N541, N199);
and AND3 (N559, N555, N117, N179);
buf BUF1 (N560, N559);
nand NAND2 (N561, N557, N503);
nor NOR3 (N562, N549, N125, N554);
xor XOR2 (N563, N66, N155);
or OR3 (N564, N550, N461, N299);
buf BUF1 (N565, N564);
not NOT1 (N566, N563);
nand NAND4 (N567, N552, N412, N18, N379);
nand NAND2 (N568, N565, N289);
not NOT1 (N569, N560);
nor NOR4 (N570, N568, N30, N269, N560);
nand NAND3 (N571, N566, N315, N256);
or OR3 (N572, N562, N273, N455);
nand NAND4 (N573, N571, N215, N450, N348);
not NOT1 (N574, N556);
and AND3 (N575, N572, N495, N221);
nand NAND4 (N576, N575, N437, N204, N232);
xor XOR2 (N577, N570, N383);
xor XOR2 (N578, N561, N46);
xor XOR2 (N579, N558, N105);
not NOT1 (N580, N576);
xor XOR2 (N581, N573, N123);
and AND3 (N582, N577, N66, N224);
xor XOR2 (N583, N551, N529);
and AND3 (N584, N579, N120, N377);
and AND2 (N585, N569, N287);
xor XOR2 (N586, N580, N45);
nand NAND4 (N587, N567, N329, N451, N159);
nor NOR3 (N588, N586, N586, N92);
buf BUF1 (N589, N582);
nand NAND3 (N590, N584, N24, N39);
and AND2 (N591, N588, N148);
xor XOR2 (N592, N583, N268);
not NOT1 (N593, N543);
nand NAND4 (N594, N585, N32, N408, N313);
nand NAND4 (N595, N593, N215, N590, N180);
xor XOR2 (N596, N388, N122);
buf BUF1 (N597, N592);
xor XOR2 (N598, N587, N542);
nor NOR2 (N599, N596, N284);
buf BUF1 (N600, N598);
nor NOR3 (N601, N591, N242, N425);
nor NOR4 (N602, N597, N305, N258, N449);
buf BUF1 (N603, N600);
not NOT1 (N604, N589);
nor NOR2 (N605, N599, N221);
and AND2 (N606, N601, N186);
and AND4 (N607, N606, N163, N176, N286);
and AND4 (N608, N581, N243, N317, N150);
or OR3 (N609, N578, N152, N453);
or OR3 (N610, N595, N489, N353);
buf BUF1 (N611, N574);
buf BUF1 (N612, N605);
and AND2 (N613, N608, N520);
xor XOR2 (N614, N612, N225);
xor XOR2 (N615, N602, N556);
not NOT1 (N616, N614);
nor NOR3 (N617, N603, N603, N118);
endmodule