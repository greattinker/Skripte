// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N907,N916,N919,N885,N917,N920,N914,N909,N911,N921;

nor NOR2 (N22, N1, N13);
buf BUF1 (N23, N20);
nor NOR3 (N24, N2, N1, N3);
or OR2 (N25, N22, N24);
or OR3 (N26, N1, N22, N19);
and AND2 (N27, N22, N5);
and AND2 (N28, N14, N14);
not NOT1 (N29, N14);
and AND4 (N30, N2, N7, N18, N6);
nor NOR3 (N31, N12, N12, N22);
xor XOR2 (N32, N15, N3);
and AND2 (N33, N8, N13);
nand NAND3 (N34, N30, N14, N8);
xor XOR2 (N35, N29, N23);
not NOT1 (N36, N9);
nand NAND3 (N37, N32, N24, N23);
not NOT1 (N38, N28);
and AND3 (N39, N36, N10, N31);
buf BUF1 (N40, N24);
or OR3 (N41, N25, N36, N33);
buf BUF1 (N42, N25);
buf BUF1 (N43, N42);
nand NAND3 (N44, N43, N20, N15);
nor NOR4 (N45, N37, N18, N37, N18);
and AND2 (N46, N35, N21);
nand NAND2 (N47, N26, N24);
nand NAND4 (N48, N27, N7, N30, N1);
buf BUF1 (N49, N40);
and AND3 (N50, N48, N49, N26);
xor XOR2 (N51, N35, N39);
and AND4 (N52, N25, N33, N2, N18);
xor XOR2 (N53, N52, N52);
xor XOR2 (N54, N41, N37);
or OR3 (N55, N53, N12, N49);
or OR2 (N56, N50, N16);
or OR2 (N57, N51, N20);
and AND3 (N58, N54, N53, N39);
nand NAND3 (N59, N57, N38, N19);
buf BUF1 (N60, N31);
or OR4 (N61, N46, N1, N10, N10);
nor NOR4 (N62, N61, N23, N29, N45);
or OR3 (N63, N26, N18, N34);
and AND4 (N64, N15, N42, N8, N12);
buf BUF1 (N65, N63);
and AND3 (N66, N47, N57, N25);
or OR4 (N67, N58, N47, N57, N20);
and AND4 (N68, N64, N51, N8, N53);
xor XOR2 (N69, N60, N22);
or OR3 (N70, N69, N27, N53);
xor XOR2 (N71, N55, N4);
not NOT1 (N72, N62);
xor XOR2 (N73, N65, N39);
buf BUF1 (N74, N70);
nor NOR4 (N75, N74, N70, N49, N47);
buf BUF1 (N76, N71);
xor XOR2 (N77, N56, N49);
nand NAND2 (N78, N72, N47);
nand NAND3 (N79, N73, N46, N69);
not NOT1 (N80, N44);
xor XOR2 (N81, N68, N19);
nand NAND3 (N82, N80, N45, N59);
xor XOR2 (N83, N58, N51);
and AND3 (N84, N77, N60, N14);
xor XOR2 (N85, N81, N55);
not NOT1 (N86, N83);
xor XOR2 (N87, N66, N55);
or OR3 (N88, N85, N76, N75);
buf BUF1 (N89, N46);
xor XOR2 (N90, N1, N21);
nand NAND2 (N91, N86, N22);
or OR4 (N92, N79, N50, N15, N89);
and AND4 (N93, N26, N58, N39, N20);
nand NAND4 (N94, N92, N84, N34, N26);
buf BUF1 (N95, N75);
nor NOR2 (N96, N94, N59);
nand NAND2 (N97, N67, N96);
xor XOR2 (N98, N45, N41);
nor NOR3 (N99, N91, N98, N51);
and AND2 (N100, N5, N16);
xor XOR2 (N101, N97, N7);
or OR2 (N102, N93, N19);
xor XOR2 (N103, N101, N14);
and AND2 (N104, N78, N2);
or OR4 (N105, N82, N27, N34, N63);
nor NOR2 (N106, N104, N4);
nand NAND3 (N107, N102, N87, N58);
nor NOR4 (N108, N58, N92, N69, N43);
nand NAND2 (N109, N107, N16);
or OR4 (N110, N99, N77, N89, N93);
buf BUF1 (N111, N110);
nand NAND2 (N112, N111, N10);
and AND4 (N113, N109, N66, N64, N109);
and AND4 (N114, N100, N35, N27, N85);
xor XOR2 (N115, N103, N106);
buf BUF1 (N116, N23);
xor XOR2 (N117, N113, N74);
not NOT1 (N118, N117);
or OR2 (N119, N95, N90);
buf BUF1 (N120, N93);
and AND2 (N121, N88, N79);
nor NOR2 (N122, N120, N79);
or OR4 (N123, N119, N90, N115, N17);
buf BUF1 (N124, N105);
not NOT1 (N125, N80);
buf BUF1 (N126, N121);
not NOT1 (N127, N125);
and AND4 (N128, N122, N47, N77, N90);
or OR4 (N129, N126, N60, N14, N116);
not NOT1 (N130, N104);
nor NOR4 (N131, N130, N114, N107, N12);
buf BUF1 (N132, N23);
or OR3 (N133, N128, N91, N104);
nor NOR2 (N134, N127, N23);
or OR2 (N135, N124, N61);
or OR4 (N136, N135, N84, N110, N121);
and AND2 (N137, N118, N108);
buf BUF1 (N138, N20);
xor XOR2 (N139, N134, N33);
not NOT1 (N140, N112);
nor NOR3 (N141, N137, N72, N6);
xor XOR2 (N142, N129, N97);
xor XOR2 (N143, N138, N55);
buf BUF1 (N144, N142);
and AND4 (N145, N140, N13, N58, N108);
nor NOR3 (N146, N139, N76, N109);
buf BUF1 (N147, N123);
and AND3 (N148, N144, N129, N78);
nand NAND3 (N149, N148, N26, N147);
not NOT1 (N150, N40);
xor XOR2 (N151, N145, N127);
xor XOR2 (N152, N146, N71);
or OR3 (N153, N141, N32, N74);
and AND2 (N154, N132, N114);
xor XOR2 (N155, N152, N137);
or OR2 (N156, N154, N139);
nor NOR3 (N157, N150, N151, N39);
xor XOR2 (N158, N10, N111);
or OR3 (N159, N156, N97, N12);
not NOT1 (N160, N136);
xor XOR2 (N161, N157, N126);
and AND2 (N162, N133, N73);
xor XOR2 (N163, N131, N108);
nand NAND4 (N164, N149, N28, N105, N145);
nor NOR4 (N165, N158, N133, N55, N134);
or OR3 (N166, N159, N77, N158);
nor NOR3 (N167, N165, N164, N42);
and AND2 (N168, N38, N118);
buf BUF1 (N169, N168);
nor NOR2 (N170, N155, N154);
or OR4 (N171, N170, N5, N83, N142);
xor XOR2 (N172, N167, N36);
nor NOR3 (N173, N163, N43, N137);
not NOT1 (N174, N169);
nor NOR2 (N175, N166, N27);
or OR3 (N176, N153, N5, N41);
and AND4 (N177, N171, N19, N98, N153);
nand NAND4 (N178, N172, N57, N4, N65);
or OR4 (N179, N177, N144, N164, N148);
nand NAND4 (N180, N161, N31, N74, N6);
not NOT1 (N181, N178);
and AND4 (N182, N174, N143, N46, N37);
nor NOR2 (N183, N5, N6);
xor XOR2 (N184, N162, N71);
not NOT1 (N185, N182);
xor XOR2 (N186, N181, N174);
or OR3 (N187, N184, N41, N94);
not NOT1 (N188, N160);
or OR3 (N189, N176, N27, N97);
nor NOR3 (N190, N173, N75, N140);
and AND4 (N191, N189, N112, N121, N185);
or OR4 (N192, N69, N172, N20, N150);
xor XOR2 (N193, N183, N182);
nor NOR2 (N194, N186, N16);
xor XOR2 (N195, N190, N175);
buf BUF1 (N196, N1);
nor NOR3 (N197, N194, N118, N71);
nand NAND4 (N198, N196, N43, N173, N107);
nand NAND2 (N199, N187, N78);
nand NAND3 (N200, N192, N93, N62);
nor NOR3 (N201, N180, N77, N76);
or OR2 (N202, N201, N15);
and AND4 (N203, N193, N132, N31, N181);
and AND4 (N204, N200, N110, N199, N138);
xor XOR2 (N205, N11, N187);
nor NOR3 (N206, N188, N13, N176);
xor XOR2 (N207, N205, N145);
or OR4 (N208, N195, N132, N167, N85);
buf BUF1 (N209, N204);
buf BUF1 (N210, N209);
nand NAND2 (N211, N202, N139);
and AND4 (N212, N207, N20, N133, N58);
nor NOR2 (N213, N191, N79);
and AND2 (N214, N212, N22);
not NOT1 (N215, N197);
buf BUF1 (N216, N215);
and AND4 (N217, N198, N47, N108, N136);
buf BUF1 (N218, N214);
or OR3 (N219, N211, N98, N118);
nand NAND4 (N220, N218, N173, N95, N40);
nor NOR3 (N221, N217, N175, N108);
nor NOR4 (N222, N210, N105, N169, N174);
not NOT1 (N223, N203);
and AND3 (N224, N223, N24, N15);
not NOT1 (N225, N219);
and AND2 (N226, N179, N161);
buf BUF1 (N227, N226);
nor NOR4 (N228, N206, N215, N84, N166);
xor XOR2 (N229, N222, N106);
nand NAND2 (N230, N213, N11);
nor NOR2 (N231, N229, N195);
not NOT1 (N232, N208);
not NOT1 (N233, N216);
not NOT1 (N234, N221);
or OR2 (N235, N232, N79);
xor XOR2 (N236, N230, N185);
xor XOR2 (N237, N220, N110);
nor NOR2 (N238, N236, N18);
nand NAND2 (N239, N231, N228);
buf BUF1 (N240, N102);
buf BUF1 (N241, N225);
nand NAND2 (N242, N238, N236);
xor XOR2 (N243, N241, N93);
buf BUF1 (N244, N233);
nand NAND4 (N245, N224, N82, N48, N244);
not NOT1 (N246, N93);
or OR4 (N247, N234, N97, N144, N203);
xor XOR2 (N248, N245, N241);
buf BUF1 (N249, N247);
not NOT1 (N250, N227);
buf BUF1 (N251, N249);
or OR3 (N252, N250, N177, N243);
or OR4 (N253, N252, N140, N6, N5);
not NOT1 (N254, N67);
buf BUF1 (N255, N248);
nand NAND2 (N256, N254, N20);
xor XOR2 (N257, N251, N140);
xor XOR2 (N258, N253, N133);
not NOT1 (N259, N242);
nor NOR4 (N260, N237, N163, N37, N116);
xor XOR2 (N261, N258, N92);
nor NOR4 (N262, N261, N147, N6, N58);
xor XOR2 (N263, N262, N214);
and AND2 (N264, N239, N54);
not NOT1 (N265, N256);
xor XOR2 (N266, N265, N204);
not NOT1 (N267, N264);
not NOT1 (N268, N266);
nor NOR3 (N269, N235, N183, N225);
buf BUF1 (N270, N269);
xor XOR2 (N271, N259, N212);
buf BUF1 (N272, N255);
or OR4 (N273, N270, N118, N35, N11);
nor NOR2 (N274, N272, N182);
xor XOR2 (N275, N240, N176);
buf BUF1 (N276, N275);
nand NAND2 (N277, N271, N27);
xor XOR2 (N278, N274, N92);
buf BUF1 (N279, N260);
xor XOR2 (N280, N279, N152);
nand NAND3 (N281, N277, N269, N167);
buf BUF1 (N282, N276);
and AND3 (N283, N263, N125, N59);
buf BUF1 (N284, N281);
nand NAND2 (N285, N283, N92);
nor NOR2 (N286, N246, N126);
xor XOR2 (N287, N273, N268);
nor NOR4 (N288, N207, N99, N209, N72);
not NOT1 (N289, N285);
or OR2 (N290, N257, N154);
and AND3 (N291, N282, N205, N123);
nor NOR4 (N292, N291, N117, N285, N168);
nand NAND4 (N293, N289, N142, N175, N214);
not NOT1 (N294, N278);
and AND2 (N295, N290, N117);
nand NAND3 (N296, N280, N86, N240);
nand NAND4 (N297, N286, N16, N21, N212);
xor XOR2 (N298, N293, N97);
and AND3 (N299, N295, N107, N71);
nor NOR3 (N300, N288, N159, N220);
and AND3 (N301, N296, N77, N133);
xor XOR2 (N302, N292, N134);
and AND4 (N303, N298, N254, N84, N32);
buf BUF1 (N304, N267);
and AND4 (N305, N302, N199, N174, N113);
and AND3 (N306, N284, N198, N12);
nand NAND2 (N307, N304, N30);
not NOT1 (N308, N294);
xor XOR2 (N309, N308, N188);
nand NAND3 (N310, N300, N68, N27);
not NOT1 (N311, N306);
or OR3 (N312, N299, N67, N123);
nor NOR4 (N313, N310, N159, N218, N101);
nand NAND4 (N314, N313, N201, N133, N138);
and AND3 (N315, N305, N62, N206);
buf BUF1 (N316, N315);
not NOT1 (N317, N311);
buf BUF1 (N318, N297);
buf BUF1 (N319, N314);
or OR4 (N320, N317, N28, N168, N256);
nand NAND3 (N321, N318, N275, N262);
xor XOR2 (N322, N309, N112);
nor NOR4 (N323, N319, N232, N65, N72);
nand NAND4 (N324, N287, N208, N145, N295);
nand NAND3 (N325, N301, N59, N162);
and AND3 (N326, N312, N15, N297);
or OR4 (N327, N303, N162, N6, N6);
and AND4 (N328, N320, N322, N194, N214);
or OR2 (N329, N197, N111);
nand NAND4 (N330, N327, N302, N136, N110);
or OR3 (N331, N330, N74, N66);
and AND4 (N332, N328, N231, N330, N319);
buf BUF1 (N333, N324);
nand NAND4 (N334, N323, N92, N303, N88);
nor NOR3 (N335, N326, N119, N14);
or OR2 (N336, N325, N314);
nand NAND4 (N337, N335, N285, N244, N277);
and AND4 (N338, N336, N227, N62, N58);
or OR2 (N339, N337, N153);
or OR3 (N340, N307, N229, N246);
buf BUF1 (N341, N339);
nor NOR4 (N342, N331, N61, N175, N27);
and AND4 (N343, N316, N182, N292, N83);
nand NAND4 (N344, N332, N259, N227, N185);
nor NOR4 (N345, N333, N3, N209, N234);
not NOT1 (N346, N340);
and AND2 (N347, N344, N77);
buf BUF1 (N348, N343);
and AND2 (N349, N345, N127);
buf BUF1 (N350, N347);
and AND4 (N351, N329, N49, N195, N234);
buf BUF1 (N352, N341);
nor NOR2 (N353, N352, N273);
buf BUF1 (N354, N348);
nor NOR4 (N355, N321, N120, N273, N194);
not NOT1 (N356, N342);
not NOT1 (N357, N338);
and AND2 (N358, N349, N312);
buf BUF1 (N359, N354);
nor NOR4 (N360, N346, N33, N287, N295);
xor XOR2 (N361, N351, N313);
not NOT1 (N362, N334);
not NOT1 (N363, N353);
xor XOR2 (N364, N360, N300);
not NOT1 (N365, N362);
nand NAND4 (N366, N364, N223, N331, N174);
or OR4 (N367, N357, N82, N26, N105);
buf BUF1 (N368, N361);
or OR4 (N369, N368, N29, N168, N365);
nand NAND4 (N370, N368, N71, N259, N178);
nand NAND4 (N371, N356, N162, N75, N163);
and AND3 (N372, N370, N365, N229);
not NOT1 (N373, N355);
buf BUF1 (N374, N359);
xor XOR2 (N375, N373, N95);
nand NAND3 (N376, N374, N331, N37);
nand NAND2 (N377, N367, N148);
buf BUF1 (N378, N376);
nor NOR4 (N379, N378, N37, N274, N21);
nor NOR2 (N380, N358, N371);
not NOT1 (N381, N75);
xor XOR2 (N382, N363, N259);
or OR2 (N383, N380, N260);
xor XOR2 (N384, N369, N199);
and AND2 (N385, N375, N292);
nand NAND2 (N386, N385, N154);
nor NOR3 (N387, N381, N225, N192);
buf BUF1 (N388, N372);
xor XOR2 (N389, N387, N118);
and AND3 (N390, N386, N208, N362);
and AND3 (N391, N366, N213, N44);
xor XOR2 (N392, N389, N5);
buf BUF1 (N393, N379);
and AND4 (N394, N382, N298, N24, N337);
or OR4 (N395, N390, N392, N332, N64);
nand NAND2 (N396, N392, N300);
buf BUF1 (N397, N393);
nor NOR2 (N398, N397, N178);
and AND4 (N399, N394, N350, N207, N89);
nor NOR4 (N400, N240, N369, N149, N42);
xor XOR2 (N401, N400, N383);
not NOT1 (N402, N244);
nand NAND4 (N403, N391, N255, N362, N344);
buf BUF1 (N404, N388);
not NOT1 (N405, N395);
nand NAND4 (N406, N403, N114, N348, N369);
buf BUF1 (N407, N405);
nor NOR2 (N408, N404, N336);
nand NAND2 (N409, N402, N13);
and AND3 (N410, N399, N356, N242);
not NOT1 (N411, N409);
nor NOR3 (N412, N384, N60, N224);
xor XOR2 (N413, N410, N322);
buf BUF1 (N414, N377);
nand NAND3 (N415, N411, N322, N98);
not NOT1 (N416, N406);
and AND2 (N417, N401, N117);
nand NAND2 (N418, N417, N21);
and AND4 (N419, N416, N252, N195, N148);
nand NAND4 (N420, N418, N372, N381, N214);
xor XOR2 (N421, N408, N289);
nand NAND2 (N422, N415, N383);
not NOT1 (N423, N419);
not NOT1 (N424, N414);
buf BUF1 (N425, N422);
nand NAND3 (N426, N412, N258, N183);
not NOT1 (N427, N424);
nor NOR2 (N428, N396, N49);
not NOT1 (N429, N398);
nor NOR3 (N430, N427, N335, N261);
buf BUF1 (N431, N420);
and AND3 (N432, N426, N148, N241);
and AND3 (N433, N423, N326, N42);
and AND2 (N434, N425, N319);
nor NOR2 (N435, N413, N145);
nor NOR3 (N436, N434, N292, N110);
buf BUF1 (N437, N432);
not NOT1 (N438, N431);
or OR3 (N439, N407, N208, N365);
not NOT1 (N440, N433);
xor XOR2 (N441, N430, N382);
buf BUF1 (N442, N428);
and AND2 (N443, N435, N181);
nor NOR2 (N444, N437, N27);
not NOT1 (N445, N442);
and AND4 (N446, N445, N279, N127, N394);
and AND3 (N447, N443, N97, N51);
and AND2 (N448, N436, N91);
and AND3 (N449, N438, N323, N383);
nand NAND2 (N450, N429, N317);
nand NAND4 (N451, N440, N446, N344, N442);
and AND3 (N452, N255, N203, N273);
buf BUF1 (N453, N439);
or OR3 (N454, N453, N61, N342);
not NOT1 (N455, N454);
xor XOR2 (N456, N447, N288);
xor XOR2 (N457, N449, N367);
nor NOR2 (N458, N452, N178);
not NOT1 (N459, N444);
xor XOR2 (N460, N441, N257);
xor XOR2 (N461, N459, N32);
nor NOR4 (N462, N461, N398, N395, N91);
nor NOR4 (N463, N460, N132, N255, N386);
not NOT1 (N464, N451);
nor NOR3 (N465, N462, N167, N341);
or OR4 (N466, N450, N153, N260, N61);
nand NAND3 (N467, N456, N103, N38);
nand NAND3 (N468, N455, N23, N333);
or OR2 (N469, N421, N131);
not NOT1 (N470, N458);
not NOT1 (N471, N469);
nor NOR2 (N472, N465, N83);
and AND4 (N473, N468, N309, N77, N308);
nand NAND2 (N474, N472, N297);
not NOT1 (N475, N466);
xor XOR2 (N476, N470, N358);
nor NOR3 (N477, N474, N204, N347);
nor NOR4 (N478, N476, N347, N200, N261);
nand NAND3 (N479, N471, N95, N140);
or OR2 (N480, N448, N325);
or OR2 (N481, N478, N471);
nand NAND3 (N482, N480, N309, N404);
and AND2 (N483, N463, N278);
and AND2 (N484, N475, N418);
or OR4 (N485, N483, N376, N37, N37);
nor NOR3 (N486, N481, N48, N124);
nand NAND3 (N487, N467, N46, N220);
or OR2 (N488, N473, N152);
buf BUF1 (N489, N479);
nand NAND4 (N490, N477, N384, N71, N94);
and AND4 (N491, N485, N448, N412, N43);
or OR3 (N492, N484, N426, N242);
or OR3 (N493, N487, N318, N447);
or OR3 (N494, N488, N323, N311);
and AND3 (N495, N464, N236, N94);
xor XOR2 (N496, N495, N104);
and AND2 (N497, N489, N90);
and AND3 (N498, N497, N228, N6);
nand NAND2 (N499, N491, N190);
and AND4 (N500, N457, N396, N456, N63);
and AND4 (N501, N492, N381, N425, N133);
and AND3 (N502, N493, N294, N254);
xor XOR2 (N503, N501, N117);
xor XOR2 (N504, N498, N471);
not NOT1 (N505, N504);
xor XOR2 (N506, N496, N157);
buf BUF1 (N507, N506);
nand NAND4 (N508, N482, N100, N156, N179);
not NOT1 (N509, N500);
nand NAND3 (N510, N499, N223, N51);
xor XOR2 (N511, N507, N198);
or OR2 (N512, N511, N152);
or OR3 (N513, N505, N447, N46);
and AND4 (N514, N512, N242, N225, N225);
and AND3 (N515, N486, N20, N84);
buf BUF1 (N516, N494);
or OR4 (N517, N508, N207, N309, N182);
nand NAND4 (N518, N502, N428, N142, N227);
nor NOR4 (N519, N509, N470, N492, N368);
and AND3 (N520, N517, N182, N370);
or OR3 (N521, N513, N229, N199);
not NOT1 (N522, N490);
nor NOR4 (N523, N521, N479, N183, N30);
not NOT1 (N524, N514);
buf BUF1 (N525, N518);
buf BUF1 (N526, N516);
xor XOR2 (N527, N515, N475);
not NOT1 (N528, N526);
not NOT1 (N529, N523);
not NOT1 (N530, N510);
and AND2 (N531, N525, N385);
or OR3 (N532, N531, N407, N79);
nand NAND3 (N533, N530, N335, N258);
and AND3 (N534, N528, N94, N254);
nor NOR3 (N535, N524, N367, N423);
nand NAND4 (N536, N503, N318, N209, N247);
nor NOR3 (N537, N522, N125, N167);
not NOT1 (N538, N534);
xor XOR2 (N539, N520, N149);
or OR3 (N540, N539, N228, N480);
nor NOR2 (N541, N533, N506);
not NOT1 (N542, N538);
not NOT1 (N543, N537);
nand NAND4 (N544, N543, N38, N485, N166);
buf BUF1 (N545, N541);
xor XOR2 (N546, N536, N230);
and AND3 (N547, N544, N329, N372);
not NOT1 (N548, N546);
buf BUF1 (N549, N535);
nand NAND3 (N550, N549, N126, N81);
and AND2 (N551, N527, N514);
and AND2 (N552, N519, N391);
and AND2 (N553, N529, N466);
not NOT1 (N554, N548);
nor NOR2 (N555, N547, N132);
nand NAND2 (N556, N540, N398);
and AND4 (N557, N555, N207, N318, N388);
buf BUF1 (N558, N553);
nor NOR4 (N559, N552, N125, N92, N220);
nor NOR2 (N560, N532, N237);
buf BUF1 (N561, N545);
nor NOR3 (N562, N559, N76, N42);
xor XOR2 (N563, N557, N263);
nor NOR2 (N564, N542, N435);
and AND3 (N565, N562, N50, N364);
and AND4 (N566, N550, N87, N59, N479);
or OR4 (N567, N558, N470, N508, N475);
nor NOR4 (N568, N567, N493, N331, N476);
or OR2 (N569, N565, N66);
not NOT1 (N570, N556);
xor XOR2 (N571, N551, N480);
and AND2 (N572, N569, N219);
and AND2 (N573, N564, N420);
nor NOR3 (N574, N570, N287, N31);
and AND3 (N575, N566, N196, N368);
nor NOR4 (N576, N575, N201, N442, N556);
nand NAND3 (N577, N554, N541, N183);
or OR2 (N578, N576, N463);
nor NOR2 (N579, N577, N443);
buf BUF1 (N580, N568);
not NOT1 (N581, N572);
buf BUF1 (N582, N571);
buf BUF1 (N583, N579);
or OR3 (N584, N578, N513, N265);
xor XOR2 (N585, N563, N139);
or OR4 (N586, N561, N281, N46, N35);
xor XOR2 (N587, N582, N407);
nand NAND2 (N588, N574, N535);
xor XOR2 (N589, N584, N526);
buf BUF1 (N590, N588);
xor XOR2 (N591, N590, N130);
not NOT1 (N592, N587);
not NOT1 (N593, N581);
buf BUF1 (N594, N586);
and AND3 (N595, N585, N22, N278);
nand NAND2 (N596, N591, N507);
or OR4 (N597, N592, N369, N79, N562);
or OR4 (N598, N589, N234, N461, N543);
xor XOR2 (N599, N596, N264);
buf BUF1 (N600, N599);
nor NOR4 (N601, N580, N298, N141, N561);
and AND2 (N602, N573, N404);
nand NAND4 (N603, N600, N368, N544, N249);
nand NAND3 (N604, N593, N396, N21);
nor NOR4 (N605, N604, N183, N13, N222);
nor NOR4 (N606, N560, N321, N123, N445);
or OR4 (N607, N598, N445, N395, N479);
and AND2 (N608, N597, N285);
not NOT1 (N609, N605);
nand NAND3 (N610, N583, N250, N345);
not NOT1 (N611, N601);
buf BUF1 (N612, N602);
not NOT1 (N613, N611);
or OR4 (N614, N613, N60, N412, N162);
nor NOR4 (N615, N610, N611, N266, N434);
or OR3 (N616, N606, N522, N473);
xor XOR2 (N617, N616, N199);
and AND2 (N618, N612, N60);
not NOT1 (N619, N607);
buf BUF1 (N620, N595);
and AND2 (N621, N615, N194);
nor NOR2 (N622, N594, N23);
or OR3 (N623, N620, N86, N468);
or OR3 (N624, N614, N161, N434);
buf BUF1 (N625, N617);
nor NOR2 (N626, N623, N303);
xor XOR2 (N627, N608, N180);
or OR2 (N628, N619, N60);
not NOT1 (N629, N626);
nand NAND3 (N630, N627, N294, N348);
or OR3 (N631, N628, N90, N163);
and AND4 (N632, N618, N175, N70, N574);
xor XOR2 (N633, N622, N419);
xor XOR2 (N634, N621, N90);
and AND2 (N635, N632, N307);
and AND4 (N636, N625, N305, N339, N158);
buf BUF1 (N637, N631);
buf BUF1 (N638, N603);
xor XOR2 (N639, N630, N552);
nor NOR2 (N640, N639, N213);
or OR2 (N641, N629, N365);
nor NOR3 (N642, N641, N78, N270);
buf BUF1 (N643, N634);
not NOT1 (N644, N638);
not NOT1 (N645, N636);
nand NAND2 (N646, N635, N219);
and AND4 (N647, N642, N287, N157, N414);
not NOT1 (N648, N637);
nand NAND3 (N649, N609, N415, N523);
and AND4 (N650, N644, N324, N179, N89);
nand NAND3 (N651, N640, N390, N589);
and AND3 (N652, N648, N603, N649);
not NOT1 (N653, N379);
buf BUF1 (N654, N652);
nor NOR3 (N655, N633, N444, N128);
nor NOR3 (N656, N653, N4, N642);
or OR4 (N657, N646, N393, N305, N118);
buf BUF1 (N658, N651);
nand NAND2 (N659, N654, N633);
nand NAND3 (N660, N647, N343, N247);
buf BUF1 (N661, N655);
nand NAND4 (N662, N661, N273, N420, N580);
or OR3 (N663, N658, N125, N229);
buf BUF1 (N664, N662);
not NOT1 (N665, N643);
buf BUF1 (N666, N664);
buf BUF1 (N667, N659);
not NOT1 (N668, N657);
buf BUF1 (N669, N645);
and AND2 (N670, N663, N57);
or OR4 (N671, N624, N34, N472, N649);
nor NOR2 (N672, N650, N347);
not NOT1 (N673, N672);
xor XOR2 (N674, N656, N477);
xor XOR2 (N675, N666, N326);
nor NOR4 (N676, N668, N604, N264, N458);
or OR2 (N677, N665, N570);
buf BUF1 (N678, N670);
buf BUF1 (N679, N674);
nand NAND4 (N680, N660, N564, N629, N13);
or OR4 (N681, N671, N633, N70, N190);
buf BUF1 (N682, N681);
not NOT1 (N683, N679);
not NOT1 (N684, N677);
not NOT1 (N685, N683);
nand NAND2 (N686, N673, N577);
nand NAND2 (N687, N682, N10);
not NOT1 (N688, N686);
nand NAND3 (N689, N678, N576, N197);
buf BUF1 (N690, N680);
buf BUF1 (N691, N676);
not NOT1 (N692, N687);
or OR2 (N693, N669, N513);
nand NAND2 (N694, N688, N565);
nor NOR2 (N695, N685, N352);
not NOT1 (N696, N693);
and AND3 (N697, N690, N522, N473);
not NOT1 (N698, N695);
or OR4 (N699, N691, N625, N155, N7);
not NOT1 (N700, N692);
nor NOR3 (N701, N696, N495, N106);
buf BUF1 (N702, N667);
nor NOR3 (N703, N700, N298, N537);
or OR4 (N704, N702, N382, N65, N650);
or OR3 (N705, N698, N677, N277);
nor NOR2 (N706, N703, N184);
or OR4 (N707, N706, N67, N465, N370);
xor XOR2 (N708, N675, N566);
and AND2 (N709, N704, N430);
buf BUF1 (N710, N689);
nand NAND4 (N711, N705, N313, N521, N23);
and AND2 (N712, N684, N479);
and AND2 (N713, N711, N61);
xor XOR2 (N714, N712, N56);
buf BUF1 (N715, N697);
xor XOR2 (N716, N699, N137);
and AND2 (N717, N710, N452);
not NOT1 (N718, N717);
nand NAND4 (N719, N716, N99, N297, N688);
buf BUF1 (N720, N707);
xor XOR2 (N721, N701, N594);
nor NOR2 (N722, N694, N142);
not NOT1 (N723, N708);
nor NOR3 (N724, N709, N378, N504);
nand NAND3 (N725, N723, N581, N195);
xor XOR2 (N726, N714, N624);
xor XOR2 (N727, N725, N86);
nand NAND2 (N728, N721, N471);
nor NOR3 (N729, N715, N52, N648);
not NOT1 (N730, N729);
and AND2 (N731, N730, N377);
nor NOR4 (N732, N713, N243, N472, N584);
nor NOR2 (N733, N728, N82);
or OR4 (N734, N732, N203, N172, N541);
and AND2 (N735, N731, N358);
not NOT1 (N736, N718);
or OR4 (N737, N724, N467, N310, N335);
nand NAND2 (N738, N722, N673);
buf BUF1 (N739, N727);
xor XOR2 (N740, N733, N164);
not NOT1 (N741, N737);
or OR2 (N742, N739, N63);
nand NAND2 (N743, N720, N556);
nor NOR4 (N744, N719, N324, N182, N124);
and AND4 (N745, N734, N731, N316, N3);
and AND2 (N746, N736, N191);
buf BUF1 (N747, N746);
nor NOR3 (N748, N741, N153, N431);
and AND2 (N749, N744, N9);
nor NOR2 (N750, N738, N147);
xor XOR2 (N751, N740, N218);
nor NOR2 (N752, N748, N10);
and AND3 (N753, N751, N196, N30);
buf BUF1 (N754, N726);
and AND4 (N755, N743, N293, N107, N706);
nand NAND4 (N756, N742, N51, N268, N424);
xor XOR2 (N757, N754, N276);
and AND4 (N758, N747, N85, N708, N163);
nand NAND3 (N759, N758, N503, N463);
nand NAND4 (N760, N749, N703, N558, N230);
buf BUF1 (N761, N756);
buf BUF1 (N762, N745);
nor NOR2 (N763, N753, N202);
buf BUF1 (N764, N735);
buf BUF1 (N765, N761);
nor NOR4 (N766, N763, N220, N590, N403);
and AND3 (N767, N762, N525, N222);
nand NAND3 (N768, N765, N81, N590);
buf BUF1 (N769, N759);
not NOT1 (N770, N760);
and AND2 (N771, N770, N116);
nor NOR4 (N772, N755, N566, N574, N620);
buf BUF1 (N773, N767);
and AND3 (N774, N752, N735, N513);
buf BUF1 (N775, N750);
nand NAND3 (N776, N769, N547, N260);
nor NOR4 (N777, N775, N322, N78, N611);
or OR3 (N778, N771, N651, N88);
buf BUF1 (N779, N773);
and AND2 (N780, N777, N733);
xor XOR2 (N781, N778, N155);
xor XOR2 (N782, N774, N138);
not NOT1 (N783, N776);
not NOT1 (N784, N772);
not NOT1 (N785, N782);
not NOT1 (N786, N784);
nor NOR2 (N787, N780, N27);
buf BUF1 (N788, N779);
nor NOR3 (N789, N785, N289, N540);
and AND3 (N790, N786, N787, N425);
and AND4 (N791, N417, N636, N769, N751);
xor XOR2 (N792, N783, N309);
and AND2 (N793, N781, N257);
nand NAND4 (N794, N790, N732, N131, N764);
buf BUF1 (N795, N135);
not NOT1 (N796, N795);
xor XOR2 (N797, N793, N175);
nand NAND2 (N798, N791, N637);
buf BUF1 (N799, N796);
xor XOR2 (N800, N797, N298);
xor XOR2 (N801, N766, N147);
and AND4 (N802, N801, N772, N750, N525);
or OR4 (N803, N789, N169, N666, N480);
or OR4 (N804, N802, N137, N683, N157);
or OR4 (N805, N804, N398, N391, N687);
or OR2 (N806, N792, N358);
nor NOR2 (N807, N805, N604);
nor NOR4 (N808, N788, N5, N6, N72);
and AND2 (N809, N768, N799);
nand NAND4 (N810, N314, N676, N393, N514);
nand NAND2 (N811, N757, N365);
buf BUF1 (N812, N803);
xor XOR2 (N813, N800, N633);
buf BUF1 (N814, N811);
nand NAND4 (N815, N813, N352, N734, N663);
not NOT1 (N816, N815);
xor XOR2 (N817, N816, N661);
xor XOR2 (N818, N810, N796);
nor NOR3 (N819, N818, N482, N455);
not NOT1 (N820, N819);
nand NAND4 (N821, N809, N476, N587, N603);
or OR3 (N822, N807, N343, N571);
and AND4 (N823, N822, N509, N99, N420);
buf BUF1 (N824, N817);
not NOT1 (N825, N794);
and AND2 (N826, N814, N509);
xor XOR2 (N827, N824, N588);
and AND4 (N828, N806, N389, N796, N88);
nand NAND2 (N829, N812, N529);
not NOT1 (N830, N829);
not NOT1 (N831, N798);
buf BUF1 (N832, N826);
nand NAND3 (N833, N830, N764, N624);
xor XOR2 (N834, N820, N757);
nor NOR4 (N835, N834, N709, N217, N520);
or OR2 (N836, N808, N414);
not NOT1 (N837, N828);
and AND3 (N838, N827, N662, N124);
and AND3 (N839, N832, N338, N205);
or OR4 (N840, N839, N306, N511, N777);
and AND4 (N841, N840, N559, N301, N417);
nand NAND2 (N842, N836, N557);
nor NOR4 (N843, N837, N629, N319, N461);
buf BUF1 (N844, N821);
and AND2 (N845, N844, N733);
nor NOR2 (N846, N841, N268);
buf BUF1 (N847, N845);
buf BUF1 (N848, N825);
and AND2 (N849, N838, N155);
not NOT1 (N850, N849);
nand NAND3 (N851, N835, N517, N287);
not NOT1 (N852, N823);
and AND4 (N853, N831, N479, N647, N697);
not NOT1 (N854, N850);
buf BUF1 (N855, N853);
xor XOR2 (N856, N855, N398);
buf BUF1 (N857, N852);
xor XOR2 (N858, N842, N148);
buf BUF1 (N859, N846);
and AND3 (N860, N854, N459, N111);
buf BUF1 (N861, N847);
and AND2 (N862, N860, N845);
nand NAND4 (N863, N848, N177, N215, N670);
xor XOR2 (N864, N862, N455);
buf BUF1 (N865, N858);
not NOT1 (N866, N864);
nand NAND2 (N867, N866, N478);
nor NOR2 (N868, N861, N657);
buf BUF1 (N869, N857);
xor XOR2 (N870, N833, N760);
xor XOR2 (N871, N869, N725);
and AND2 (N872, N865, N302);
not NOT1 (N873, N851);
and AND4 (N874, N859, N70, N339, N194);
and AND3 (N875, N871, N219, N129);
buf BUF1 (N876, N868);
and AND4 (N877, N874, N174, N417, N775);
and AND2 (N878, N843, N134);
or OR2 (N879, N872, N14);
or OR3 (N880, N867, N299, N357);
not NOT1 (N881, N876);
nor NOR3 (N882, N879, N843, N628);
or OR2 (N883, N882, N58);
xor XOR2 (N884, N873, N700);
or OR4 (N885, N875, N560, N183, N535);
and AND2 (N886, N883, N5);
and AND4 (N887, N884, N725, N521, N254);
nor NOR3 (N888, N878, N286, N464);
nor NOR4 (N889, N863, N36, N657, N292);
and AND4 (N890, N881, N840, N150, N153);
or OR2 (N891, N877, N359);
buf BUF1 (N892, N887);
and AND4 (N893, N892, N473, N516, N413);
buf BUF1 (N894, N870);
or OR4 (N895, N891, N651, N438, N206);
xor XOR2 (N896, N893, N260);
not NOT1 (N897, N888);
nor NOR4 (N898, N886, N199, N582, N828);
and AND3 (N899, N897, N853, N562);
buf BUF1 (N900, N896);
not NOT1 (N901, N880);
nor NOR3 (N902, N900, N739, N129);
buf BUF1 (N903, N899);
nand NAND2 (N904, N894, N416);
or OR3 (N905, N898, N901, N596);
nor NOR4 (N906, N879, N549, N877, N873);
or OR3 (N907, N903, N58, N878);
and AND3 (N908, N902, N390, N133);
and AND4 (N909, N904, N127, N113, N351);
or OR2 (N910, N856, N330);
nor NOR3 (N911, N889, N213, N241);
nand NAND4 (N912, N890, N581, N709, N478);
nor NOR2 (N913, N912, N397);
nor NOR2 (N914, N913, N865);
buf BUF1 (N915, N906);
xor XOR2 (N916, N895, N802);
xor XOR2 (N917, N905, N30);
xor XOR2 (N918, N908, N861);
xor XOR2 (N919, N918, N20);
buf BUF1 (N920, N915);
and AND3 (N921, N910, N651, N600);
endmodule