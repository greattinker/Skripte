// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N195,N219,N204,N220,N215,N216,N217,N213,N205,N221;

nand NAND3 (N22, N11, N2, N19);
nor NOR3 (N23, N8, N7, N5);
not NOT1 (N24, N3);
xor XOR2 (N25, N8, N11);
nand NAND4 (N26, N17, N17, N11, N24);
buf BUF1 (N27, N19);
xor XOR2 (N28, N2, N20);
or OR4 (N29, N3, N21, N11, N10);
xor XOR2 (N30, N25, N2);
and AND3 (N31, N4, N21, N25);
not NOT1 (N32, N11);
nand NAND3 (N33, N26, N7, N4);
nand NAND3 (N34, N7, N1, N25);
xor XOR2 (N35, N27, N9);
xor XOR2 (N36, N33, N31);
nand NAND3 (N37, N27, N9, N17);
or OR2 (N38, N29, N7);
xor XOR2 (N39, N23, N12);
buf BUF1 (N40, N34);
not NOT1 (N41, N40);
xor XOR2 (N42, N32, N8);
buf BUF1 (N43, N35);
xor XOR2 (N44, N37, N43);
xor XOR2 (N45, N40, N23);
or OR2 (N46, N39, N14);
not NOT1 (N47, N38);
not NOT1 (N48, N47);
not NOT1 (N49, N48);
buf BUF1 (N50, N28);
not NOT1 (N51, N42);
xor XOR2 (N52, N30, N39);
buf BUF1 (N53, N44);
xor XOR2 (N54, N51, N43);
xor XOR2 (N55, N41, N21);
or OR2 (N56, N54, N11);
nor NOR3 (N57, N56, N48, N1);
buf BUF1 (N58, N49);
xor XOR2 (N59, N53, N10);
and AND4 (N60, N55, N33, N21, N40);
not NOT1 (N61, N57);
buf BUF1 (N62, N36);
nand NAND3 (N63, N59, N29, N26);
buf BUF1 (N64, N58);
xor XOR2 (N65, N22, N3);
buf BUF1 (N66, N45);
and AND4 (N67, N62, N28, N60, N53);
nand NAND4 (N68, N48, N15, N29, N23);
xor XOR2 (N69, N66, N9);
and AND4 (N70, N46, N5, N9, N57);
nand NAND3 (N71, N65, N39, N36);
not NOT1 (N72, N71);
not NOT1 (N73, N69);
not NOT1 (N74, N72);
and AND3 (N75, N68, N18, N44);
not NOT1 (N76, N75);
xor XOR2 (N77, N61, N65);
or OR2 (N78, N63, N23);
not NOT1 (N79, N64);
xor XOR2 (N80, N52, N48);
nor NOR2 (N81, N80, N20);
buf BUF1 (N82, N79);
nor NOR2 (N83, N67, N55);
nand NAND2 (N84, N50, N49);
nor NOR3 (N85, N70, N13, N68);
nor NOR2 (N86, N76, N24);
buf BUF1 (N87, N85);
nor NOR3 (N88, N77, N32, N29);
xor XOR2 (N89, N87, N44);
nor NOR4 (N90, N73, N4, N33, N57);
buf BUF1 (N91, N84);
xor XOR2 (N92, N86, N71);
buf BUF1 (N93, N74);
not NOT1 (N94, N81);
and AND3 (N95, N91, N8, N8);
nor NOR3 (N96, N92, N6, N20);
nor NOR3 (N97, N89, N9, N62);
xor XOR2 (N98, N94, N48);
buf BUF1 (N99, N95);
and AND2 (N100, N88, N13);
nor NOR2 (N101, N97, N91);
buf BUF1 (N102, N101);
or OR3 (N103, N78, N51, N65);
nand NAND2 (N104, N102, N42);
xor XOR2 (N105, N93, N33);
buf BUF1 (N106, N83);
nor NOR2 (N107, N99, N86);
not NOT1 (N108, N90);
nor NOR3 (N109, N104, N92, N99);
and AND3 (N110, N100, N69, N63);
xor XOR2 (N111, N109, N106);
and AND2 (N112, N40, N61);
nand NAND4 (N113, N105, N68, N3, N25);
not NOT1 (N114, N82);
and AND4 (N115, N113, N71, N73, N45);
or OR2 (N116, N112, N61);
or OR3 (N117, N114, N88, N51);
nor NOR2 (N118, N98, N13);
buf BUF1 (N119, N96);
and AND2 (N120, N119, N50);
or OR3 (N121, N120, N87, N88);
not NOT1 (N122, N121);
or OR4 (N123, N117, N90, N8, N56);
or OR4 (N124, N123, N34, N6, N14);
nand NAND3 (N125, N103, N50, N21);
nor NOR2 (N126, N107, N110);
nand NAND3 (N127, N29, N105, N80);
or OR2 (N128, N116, N108);
nand NAND4 (N129, N115, N102, N40, N42);
xor XOR2 (N130, N24, N88);
buf BUF1 (N131, N130);
and AND4 (N132, N124, N51, N92, N19);
or OR4 (N133, N118, N59, N70, N42);
nor NOR2 (N134, N127, N78);
xor XOR2 (N135, N133, N73);
xor XOR2 (N136, N126, N41);
or OR4 (N137, N132, N25, N98, N21);
and AND4 (N138, N129, N15, N123, N37);
nor NOR4 (N139, N111, N4, N41, N11);
buf BUF1 (N140, N138);
or OR4 (N141, N131, N64, N58, N103);
xor XOR2 (N142, N141, N27);
nand NAND3 (N143, N128, N2, N47);
buf BUF1 (N144, N137);
nand NAND3 (N145, N136, N32, N117);
nor NOR2 (N146, N125, N125);
xor XOR2 (N147, N146, N3);
xor XOR2 (N148, N144, N12);
or OR4 (N149, N143, N97, N147, N92);
nand NAND3 (N150, N17, N59, N10);
xor XOR2 (N151, N142, N78);
and AND4 (N152, N134, N136, N78, N90);
xor XOR2 (N153, N145, N43);
and AND3 (N154, N135, N127, N91);
and AND2 (N155, N150, N154);
nand NAND4 (N156, N36, N26, N71, N108);
and AND3 (N157, N122, N36, N133);
nor NOR3 (N158, N157, N103, N59);
not NOT1 (N159, N153);
xor XOR2 (N160, N155, N105);
not NOT1 (N161, N159);
or OR2 (N162, N139, N44);
and AND4 (N163, N140, N125, N68, N129);
and AND3 (N164, N151, N105, N132);
nand NAND3 (N165, N152, N4, N4);
nand NAND3 (N166, N158, N61, N75);
or OR3 (N167, N162, N132, N21);
nand NAND4 (N168, N167, N1, N37, N23);
nand NAND2 (N169, N148, N117);
not NOT1 (N170, N160);
buf BUF1 (N171, N163);
xor XOR2 (N172, N156, N157);
nor NOR2 (N173, N171, N5);
or OR4 (N174, N170, N11, N164, N3);
nor NOR2 (N175, N94, N156);
and AND2 (N176, N169, N12);
or OR4 (N177, N176, N79, N141, N65);
xor XOR2 (N178, N166, N133);
or OR2 (N179, N165, N45);
or OR2 (N180, N172, N142);
nor NOR2 (N181, N179, N10);
not NOT1 (N182, N168);
and AND3 (N183, N178, N107, N75);
or OR4 (N184, N180, N157, N10, N125);
not NOT1 (N185, N149);
not NOT1 (N186, N183);
and AND3 (N187, N161, N139, N100);
xor XOR2 (N188, N181, N36);
and AND2 (N189, N186, N169);
nor NOR4 (N190, N189, N106, N139, N66);
and AND4 (N191, N187, N120, N93, N95);
buf BUF1 (N192, N191);
nand NAND2 (N193, N182, N88);
buf BUF1 (N194, N184);
buf BUF1 (N195, N193);
nand NAND2 (N196, N188, N173);
xor XOR2 (N197, N56, N155);
and AND4 (N198, N197, N25, N92, N148);
nor NOR3 (N199, N175, N24, N57);
and AND2 (N200, N190, N90);
xor XOR2 (N201, N192, N145);
not NOT1 (N202, N174);
xor XOR2 (N203, N194, N45);
xor XOR2 (N204, N199, N187);
or OR3 (N205, N200, N73, N185);
nand NAND4 (N206, N162, N144, N142, N58);
xor XOR2 (N207, N206, N62);
xor XOR2 (N208, N207, N41);
xor XOR2 (N209, N202, N96);
nand NAND3 (N210, N198, N16, N130);
nand NAND2 (N211, N208, N123);
or OR3 (N212, N203, N62, N128);
nand NAND3 (N213, N177, N47, N3);
and AND3 (N214, N201, N143, N185);
not NOT1 (N215, N214);
nor NOR3 (N216, N209, N159, N9);
nand NAND3 (N217, N211, N37, N97);
nand NAND2 (N218, N212, N62);
not NOT1 (N219, N218);
not NOT1 (N220, N196);
not NOT1 (N221, N210);
endmodule