// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N119,N118,N110,N108,N116,N120,N95,N114,N113,N121;

or OR4 (N22, N12, N1, N13, N20);
xor XOR2 (N23, N9, N17);
and AND3 (N24, N4, N7, N14);
nand NAND4 (N25, N20, N18, N9, N17);
and AND4 (N26, N15, N10, N19, N11);
buf BUF1 (N27, N4);
not NOT1 (N28, N13);
not NOT1 (N29, N10);
xor XOR2 (N30, N14, N22);
or OR2 (N31, N18, N7);
xor XOR2 (N32, N28, N14);
nor NOR4 (N33, N1, N3, N4, N18);
nor NOR3 (N34, N31, N24, N22);
and AND3 (N35, N5, N30, N20);
not NOT1 (N36, N34);
xor XOR2 (N37, N11, N29);
buf BUF1 (N38, N1);
or OR4 (N39, N32, N12, N29, N13);
not NOT1 (N40, N39);
xor XOR2 (N41, N27, N1);
nand NAND3 (N42, N23, N19, N24);
xor XOR2 (N43, N37, N24);
and AND4 (N44, N36, N21, N41, N28);
nor NOR4 (N45, N22, N15, N11, N44);
not NOT1 (N46, N21);
or OR2 (N47, N35, N33);
buf BUF1 (N48, N2);
or OR3 (N49, N43, N1, N48);
xor XOR2 (N50, N29, N43);
buf BUF1 (N51, N42);
or OR3 (N52, N26, N7, N41);
buf BUF1 (N53, N50);
or OR4 (N54, N51, N31, N38, N7);
nor NOR2 (N55, N38, N12);
nand NAND3 (N56, N54, N33, N30);
nand NAND4 (N57, N45, N6, N29, N23);
not NOT1 (N58, N25);
or OR2 (N59, N58, N4);
xor XOR2 (N60, N52, N18);
xor XOR2 (N61, N40, N2);
and AND3 (N62, N60, N41, N48);
or OR2 (N63, N55, N21);
or OR4 (N64, N59, N41, N63, N59);
nand NAND4 (N65, N29, N48, N60, N21);
nor NOR2 (N66, N64, N36);
not NOT1 (N67, N49);
or OR4 (N68, N65, N32, N14, N23);
and AND4 (N69, N57, N44, N17, N30);
buf BUF1 (N70, N61);
not NOT1 (N71, N67);
and AND3 (N72, N68, N53, N56);
not NOT1 (N73, N54);
buf BUF1 (N74, N36);
and AND4 (N75, N70, N36, N70, N6);
and AND2 (N76, N71, N27);
xor XOR2 (N77, N46, N26);
not NOT1 (N78, N76);
and AND4 (N79, N62, N57, N45, N57);
nand NAND2 (N80, N75, N38);
nand NAND4 (N81, N80, N60, N20, N41);
not NOT1 (N82, N72);
buf BUF1 (N83, N82);
and AND2 (N84, N77, N41);
or OR2 (N85, N83, N35);
or OR4 (N86, N47, N33, N67, N53);
buf BUF1 (N87, N74);
buf BUF1 (N88, N87);
nor NOR3 (N89, N69, N63, N1);
not NOT1 (N90, N86);
and AND2 (N91, N89, N64);
nor NOR2 (N92, N78, N82);
buf BUF1 (N93, N73);
nor NOR2 (N94, N84, N8);
and AND2 (N95, N81, N78);
not NOT1 (N96, N93);
xor XOR2 (N97, N79, N48);
buf BUF1 (N98, N94);
nor NOR4 (N99, N92, N64, N85, N65);
buf BUF1 (N100, N52);
and AND2 (N101, N99, N71);
nand NAND3 (N102, N90, N73, N59);
xor XOR2 (N103, N66, N62);
or OR2 (N104, N102, N3);
nor NOR2 (N105, N97, N100);
nand NAND4 (N106, N63, N4, N46, N81);
not NOT1 (N107, N96);
buf BUF1 (N108, N88);
buf BUF1 (N109, N98);
nand NAND4 (N110, N103, N105, N31, N32);
or OR4 (N111, N97, N76, N25, N40);
and AND4 (N112, N109, N96, N84, N87);
and AND2 (N113, N111, N103);
or OR3 (N114, N104, N8, N39);
xor XOR2 (N115, N112, N101);
or OR4 (N116, N76, N58, N106, N98);
buf BUF1 (N117, N103);
nor NOR2 (N118, N107, N55);
not NOT1 (N119, N115);
or OR4 (N120, N117, N4, N89, N54);
buf BUF1 (N121, N91);
endmodule