// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;

output N812,N802,N808,N801,N810,N811,N807,N780,N813,N814;

nand NAND4 (N15, N3, N5, N7, N10);
or OR4 (N16, N7, N15, N9, N5);
buf BUF1 (N17, N12);
xor XOR2 (N18, N15, N12);
or OR4 (N19, N5, N17, N15, N1);
or OR2 (N20, N11, N13);
and AND3 (N21, N5, N11, N13);
xor XOR2 (N22, N14, N1);
not NOT1 (N23, N18);
or OR3 (N24, N14, N14, N12);
not NOT1 (N25, N23);
xor XOR2 (N26, N5, N17);
or OR4 (N27, N25, N5, N3, N6);
not NOT1 (N28, N7);
buf BUF1 (N29, N11);
nor NOR2 (N30, N26, N26);
nand NAND2 (N31, N30, N6);
nor NOR2 (N32, N20, N29);
xor XOR2 (N33, N28, N6);
and AND2 (N34, N2, N4);
or OR2 (N35, N31, N20);
buf BUF1 (N36, N35);
or OR2 (N37, N36, N24);
buf BUF1 (N38, N30);
or OR2 (N39, N16, N2);
and AND2 (N40, N27, N33);
buf BUF1 (N41, N17);
not NOT1 (N42, N21);
nand NAND2 (N43, N37, N13);
nand NAND4 (N44, N32, N8, N2, N6);
nand NAND2 (N45, N44, N14);
and AND2 (N46, N45, N31);
nand NAND3 (N47, N39, N34, N41);
or OR2 (N48, N44, N33);
nor NOR2 (N49, N21, N13);
buf BUF1 (N50, N40);
not NOT1 (N51, N42);
not NOT1 (N52, N46);
buf BUF1 (N53, N38);
nand NAND4 (N54, N47, N6, N6, N48);
buf BUF1 (N55, N4);
not NOT1 (N56, N53);
and AND4 (N57, N19, N42, N12, N10);
nor NOR2 (N58, N54, N19);
not NOT1 (N59, N56);
nor NOR2 (N60, N58, N44);
nand NAND4 (N61, N49, N13, N25, N31);
and AND3 (N62, N55, N56, N11);
or OR3 (N63, N61, N44, N6);
xor XOR2 (N64, N60, N34);
nor NOR2 (N65, N57, N47);
nand NAND2 (N66, N63, N2);
or OR4 (N67, N65, N59, N7, N12);
nand NAND2 (N68, N62, N20);
xor XOR2 (N69, N10, N9);
xor XOR2 (N70, N52, N31);
or OR2 (N71, N43, N26);
nand NAND2 (N72, N64, N69);
and AND3 (N73, N30, N72, N20);
and AND3 (N74, N57, N47, N66);
nand NAND3 (N75, N29, N2, N58);
not NOT1 (N76, N50);
not NOT1 (N77, N76);
buf BUF1 (N78, N75);
nand NAND2 (N79, N67, N3);
nand NAND4 (N80, N78, N27, N44, N50);
or OR4 (N81, N70, N56, N63, N16);
and AND3 (N82, N73, N65, N78);
or OR2 (N83, N81, N58);
or OR3 (N84, N79, N64, N63);
not NOT1 (N85, N22);
nand NAND4 (N86, N51, N19, N26, N64);
nand NAND4 (N87, N71, N24, N38, N76);
nand NAND3 (N88, N83, N56, N38);
nand NAND2 (N89, N74, N71);
or OR2 (N90, N84, N59);
nor NOR3 (N91, N89, N47, N18);
or OR2 (N92, N68, N45);
xor XOR2 (N93, N82, N54);
and AND2 (N94, N92, N90);
xor XOR2 (N95, N37, N19);
nor NOR3 (N96, N95, N17, N51);
and AND2 (N97, N87, N18);
xor XOR2 (N98, N80, N52);
or OR3 (N99, N86, N94, N46);
not NOT1 (N100, N59);
or OR3 (N101, N98, N92, N80);
nand NAND2 (N102, N88, N14);
xor XOR2 (N103, N77, N99);
nand NAND2 (N104, N30, N44);
and AND4 (N105, N85, N78, N70, N54);
xor XOR2 (N106, N102, N13);
xor XOR2 (N107, N103, N12);
buf BUF1 (N108, N96);
nor NOR2 (N109, N107, N73);
not NOT1 (N110, N108);
buf BUF1 (N111, N100);
or OR4 (N112, N91, N41, N70, N23);
xor XOR2 (N113, N101, N57);
nor NOR2 (N114, N93, N15);
nor NOR3 (N115, N114, N41, N13);
xor XOR2 (N116, N106, N41);
or OR4 (N117, N109, N48, N44, N84);
or OR4 (N118, N112, N116, N32, N18);
nand NAND4 (N119, N69, N35, N75, N53);
nand NAND3 (N120, N117, N86, N52);
and AND3 (N121, N118, N2, N68);
xor XOR2 (N122, N113, N101);
or OR3 (N123, N122, N87, N48);
nor NOR2 (N124, N120, N86);
not NOT1 (N125, N105);
nand NAND3 (N126, N119, N46, N7);
and AND2 (N127, N110, N32);
or OR4 (N128, N115, N122, N38, N101);
nand NAND3 (N129, N127, N66, N60);
not NOT1 (N130, N97);
not NOT1 (N131, N121);
nand NAND2 (N132, N111, N50);
buf BUF1 (N133, N123);
or OR2 (N134, N128, N116);
nand NAND2 (N135, N134, N23);
nor NOR2 (N136, N126, N58);
nor NOR2 (N137, N136, N135);
not NOT1 (N138, N101);
buf BUF1 (N139, N131);
and AND4 (N140, N129, N119, N10, N109);
not NOT1 (N141, N132);
and AND3 (N142, N138, N96, N141);
nor NOR2 (N143, N6, N127);
and AND4 (N144, N124, N132, N67, N109);
buf BUF1 (N145, N130);
nand NAND2 (N146, N144, N63);
nand NAND4 (N147, N140, N83, N29, N29);
or OR4 (N148, N146, N35, N119, N126);
xor XOR2 (N149, N147, N52);
not NOT1 (N150, N133);
buf BUF1 (N151, N148);
not NOT1 (N152, N145);
not NOT1 (N153, N143);
not NOT1 (N154, N149);
nor NOR4 (N155, N139, N28, N38, N91);
and AND3 (N156, N155, N143, N112);
nor NOR2 (N157, N150, N125);
nor NOR3 (N158, N86, N82, N108);
or OR3 (N159, N142, N143, N146);
buf BUF1 (N160, N156);
nor NOR3 (N161, N137, N21, N52);
nor NOR4 (N162, N161, N158, N20, N136);
nand NAND2 (N163, N142, N61);
xor XOR2 (N164, N157, N36);
or OR3 (N165, N162, N140, N94);
and AND4 (N166, N163, N148, N60, N112);
nor NOR2 (N167, N152, N89);
or OR2 (N168, N151, N63);
not NOT1 (N169, N164);
xor XOR2 (N170, N104, N75);
buf BUF1 (N171, N165);
buf BUF1 (N172, N154);
xor XOR2 (N173, N159, N79);
nor NOR2 (N174, N168, N39);
buf BUF1 (N175, N153);
not NOT1 (N176, N174);
xor XOR2 (N177, N170, N100);
nor NOR4 (N178, N171, N13, N137, N85);
nand NAND2 (N179, N175, N110);
nand NAND3 (N180, N167, N37, N175);
not NOT1 (N181, N178);
nand NAND3 (N182, N177, N111, N52);
or OR4 (N183, N180, N121, N39, N85);
nor NOR4 (N184, N173, N169, N115, N94);
nor NOR4 (N185, N172, N68, N146, N31);
xor XOR2 (N186, N127, N151);
nor NOR2 (N187, N184, N10);
not NOT1 (N188, N160);
nand NAND4 (N189, N186, N140, N51, N133);
nor NOR3 (N190, N185, N109, N189);
or OR3 (N191, N141, N6, N1);
nor NOR3 (N192, N166, N69, N152);
not NOT1 (N193, N191);
xor XOR2 (N194, N187, N70);
xor XOR2 (N195, N181, N65);
nand NAND3 (N196, N192, N179, N152);
nand NAND4 (N197, N157, N4, N149, N152);
buf BUF1 (N198, N190);
nor NOR2 (N199, N195, N54);
nand NAND4 (N200, N193, N30, N1, N7);
nor NOR4 (N201, N196, N122, N200, N121);
not NOT1 (N202, N73);
not NOT1 (N203, N194);
nand NAND4 (N204, N182, N108, N176, N167);
not NOT1 (N205, N86);
or OR3 (N206, N203, N198, N125);
not NOT1 (N207, N1);
xor XOR2 (N208, N199, N13);
nand NAND2 (N209, N206, N99);
buf BUF1 (N210, N201);
nor NOR3 (N211, N188, N80, N93);
nand NAND3 (N212, N209, N23, N198);
and AND2 (N213, N208, N98);
nor NOR3 (N214, N197, N33, N128);
not NOT1 (N215, N210);
xor XOR2 (N216, N213, N141);
not NOT1 (N217, N215);
xor XOR2 (N218, N217, N65);
not NOT1 (N219, N212);
xor XOR2 (N220, N205, N56);
not NOT1 (N221, N207);
or OR2 (N222, N219, N134);
xor XOR2 (N223, N221, N62);
buf BUF1 (N224, N220);
buf BUF1 (N225, N223);
buf BUF1 (N226, N204);
and AND3 (N227, N222, N107, N195);
nor NOR2 (N228, N211, N101);
nand NAND2 (N229, N214, N20);
nand NAND4 (N230, N218, N46, N144, N7);
and AND2 (N231, N216, N28);
and AND2 (N232, N202, N88);
not NOT1 (N233, N228);
xor XOR2 (N234, N224, N101);
nand NAND2 (N235, N183, N142);
nand NAND2 (N236, N231, N166);
and AND2 (N237, N236, N126);
nand NAND3 (N238, N235, N80, N200);
xor XOR2 (N239, N229, N139);
and AND4 (N240, N233, N199, N78, N53);
nand NAND3 (N241, N239, N45, N47);
nand NAND4 (N242, N230, N189, N10, N150);
nand NAND4 (N243, N240, N219, N202, N16);
or OR3 (N244, N241, N20, N232);
nand NAND3 (N245, N241, N152, N187);
nand NAND4 (N246, N237, N34, N159, N112);
and AND3 (N247, N242, N43, N11);
xor XOR2 (N248, N247, N121);
not NOT1 (N249, N243);
nand NAND4 (N250, N226, N91, N61, N140);
buf BUF1 (N251, N234);
nand NAND2 (N252, N251, N27);
xor XOR2 (N253, N227, N223);
buf BUF1 (N254, N250);
or OR2 (N255, N254, N9);
buf BUF1 (N256, N253);
and AND2 (N257, N249, N59);
buf BUF1 (N258, N252);
buf BUF1 (N259, N245);
buf BUF1 (N260, N257);
and AND4 (N261, N246, N212, N40, N216);
buf BUF1 (N262, N258);
buf BUF1 (N263, N256);
buf BUF1 (N264, N262);
xor XOR2 (N265, N261, N213);
xor XOR2 (N266, N238, N29);
buf BUF1 (N267, N265);
nor NOR3 (N268, N259, N83, N161);
xor XOR2 (N269, N268, N200);
xor XOR2 (N270, N264, N208);
xor XOR2 (N271, N270, N173);
not NOT1 (N272, N271);
nand NAND3 (N273, N260, N37, N119);
buf BUF1 (N274, N244);
nand NAND3 (N275, N263, N85, N100);
nand NAND4 (N276, N275, N127, N60, N275);
buf BUF1 (N277, N267);
and AND2 (N278, N274, N174);
xor XOR2 (N279, N276, N152);
buf BUF1 (N280, N273);
not NOT1 (N281, N279);
nand NAND2 (N282, N255, N164);
not NOT1 (N283, N281);
or OR2 (N284, N272, N25);
and AND4 (N285, N277, N224, N146, N280);
and AND4 (N286, N56, N140, N22, N30);
or OR3 (N287, N248, N164, N138);
and AND2 (N288, N266, N81);
buf BUF1 (N289, N282);
xor XOR2 (N290, N285, N286);
nand NAND2 (N291, N146, N104);
and AND2 (N292, N290, N69);
nand NAND3 (N293, N288, N35, N260);
buf BUF1 (N294, N291);
and AND4 (N295, N278, N95, N62, N24);
xor XOR2 (N296, N287, N81);
xor XOR2 (N297, N296, N131);
nor NOR4 (N298, N292, N46, N51, N178);
nor NOR4 (N299, N289, N203, N160, N278);
buf BUF1 (N300, N283);
xor XOR2 (N301, N295, N124);
buf BUF1 (N302, N297);
not NOT1 (N303, N302);
and AND2 (N304, N299, N239);
not NOT1 (N305, N300);
not NOT1 (N306, N284);
xor XOR2 (N307, N303, N130);
not NOT1 (N308, N307);
or OR4 (N309, N305, N79, N308, N27);
xor XOR2 (N310, N73, N41);
buf BUF1 (N311, N298);
and AND3 (N312, N304, N188, N267);
nand NAND4 (N313, N301, N75, N5, N309);
or OR3 (N314, N17, N295, N56);
buf BUF1 (N315, N314);
nor NOR2 (N316, N312, N43);
buf BUF1 (N317, N293);
or OR2 (N318, N225, N147);
buf BUF1 (N319, N313);
not NOT1 (N320, N316);
xor XOR2 (N321, N269, N121);
nand NAND3 (N322, N310, N138, N166);
not NOT1 (N323, N322);
or OR2 (N324, N294, N260);
and AND4 (N325, N318, N263, N160, N276);
or OR2 (N326, N317, N26);
nor NOR3 (N327, N311, N136, N232);
not NOT1 (N328, N320);
buf BUF1 (N329, N326);
or OR2 (N330, N306, N127);
nand NAND3 (N331, N328, N193, N325);
xor XOR2 (N332, N136, N284);
or OR3 (N333, N324, N146, N214);
not NOT1 (N334, N315);
and AND3 (N335, N323, N54, N209);
and AND3 (N336, N334, N190, N325);
buf BUF1 (N337, N329);
or OR4 (N338, N333, N6, N107, N96);
xor XOR2 (N339, N337, N41);
buf BUF1 (N340, N331);
and AND3 (N341, N340, N111, N320);
xor XOR2 (N342, N339, N212);
and AND2 (N343, N335, N182);
nor NOR2 (N344, N319, N37);
and AND3 (N345, N341, N195, N207);
and AND2 (N346, N332, N1);
nand NAND3 (N347, N327, N256, N127);
or OR3 (N348, N343, N111, N105);
nand NAND3 (N349, N348, N216, N41);
xor XOR2 (N350, N338, N165);
not NOT1 (N351, N330);
nand NAND2 (N352, N351, N141);
buf BUF1 (N353, N347);
not NOT1 (N354, N344);
xor XOR2 (N355, N353, N111);
not NOT1 (N356, N336);
buf BUF1 (N357, N355);
not NOT1 (N358, N321);
xor XOR2 (N359, N350, N64);
nor NOR2 (N360, N346, N270);
and AND4 (N361, N358, N194, N213, N193);
xor XOR2 (N362, N345, N265);
and AND3 (N363, N359, N348, N342);
xor XOR2 (N364, N107, N182);
not NOT1 (N365, N354);
or OR3 (N366, N361, N202, N210);
or OR2 (N367, N362, N108);
and AND2 (N368, N363, N244);
and AND2 (N369, N360, N295);
xor XOR2 (N370, N369, N17);
and AND2 (N371, N365, N114);
buf BUF1 (N372, N371);
not NOT1 (N373, N364);
nand NAND3 (N374, N357, N24, N92);
xor XOR2 (N375, N352, N86);
or OR3 (N376, N356, N273, N93);
or OR3 (N377, N372, N308, N52);
and AND4 (N378, N366, N77, N276, N286);
not NOT1 (N379, N378);
xor XOR2 (N380, N374, N361);
and AND2 (N381, N373, N311);
not NOT1 (N382, N349);
not NOT1 (N383, N381);
nand NAND3 (N384, N376, N301, N338);
buf BUF1 (N385, N383);
xor XOR2 (N386, N379, N128);
nand NAND3 (N387, N370, N339, N45);
and AND4 (N388, N377, N119, N300, N108);
or OR4 (N389, N380, N41, N342, N188);
not NOT1 (N390, N384);
xor XOR2 (N391, N386, N358);
nor NOR3 (N392, N368, N324, N96);
and AND4 (N393, N367, N66, N194, N304);
nor NOR2 (N394, N392, N367);
or OR4 (N395, N387, N229, N125, N32);
nor NOR4 (N396, N389, N141, N81, N324);
and AND3 (N397, N396, N168, N67);
xor XOR2 (N398, N394, N294);
not NOT1 (N399, N393);
buf BUF1 (N400, N382);
or OR2 (N401, N390, N391);
nand NAND4 (N402, N292, N200, N165, N86);
not NOT1 (N403, N388);
xor XOR2 (N404, N399, N297);
nor NOR3 (N405, N402, N357, N392);
nor NOR3 (N406, N403, N332, N60);
not NOT1 (N407, N375);
and AND3 (N408, N395, N104, N269);
not NOT1 (N409, N398);
not NOT1 (N410, N404);
xor XOR2 (N411, N406, N385);
or OR3 (N412, N378, N144, N406);
nand NAND3 (N413, N397, N186, N398);
nor NOR2 (N414, N401, N378);
and AND2 (N415, N413, N147);
and AND3 (N416, N412, N154, N337);
nor NOR2 (N417, N407, N80);
or OR4 (N418, N405, N60, N16, N243);
or OR3 (N419, N400, N166, N11);
nor NOR2 (N420, N414, N315);
xor XOR2 (N421, N419, N315);
or OR3 (N422, N418, N281, N5);
nor NOR3 (N423, N422, N79, N187);
buf BUF1 (N424, N416);
xor XOR2 (N425, N408, N403);
nand NAND4 (N426, N421, N252, N243, N141);
or OR2 (N427, N417, N377);
not NOT1 (N428, N411);
xor XOR2 (N429, N423, N321);
xor XOR2 (N430, N428, N385);
xor XOR2 (N431, N415, N205);
nor NOR2 (N432, N424, N129);
nand NAND3 (N433, N425, N157, N321);
nand NAND2 (N434, N433, N17);
nand NAND4 (N435, N431, N47, N295, N31);
not NOT1 (N436, N427);
xor XOR2 (N437, N410, N6);
buf BUF1 (N438, N409);
xor XOR2 (N439, N420, N72);
nor NOR4 (N440, N429, N273, N166, N379);
xor XOR2 (N441, N437, N303);
nand NAND3 (N442, N430, N298, N141);
nor NOR2 (N443, N432, N421);
nor NOR3 (N444, N440, N168, N142);
nand NAND3 (N445, N439, N128, N249);
or OR2 (N446, N442, N29);
nor NOR2 (N447, N441, N179);
nor NOR2 (N448, N447, N350);
and AND4 (N449, N445, N422, N112, N340);
nand NAND2 (N450, N446, N107);
and AND3 (N451, N443, N203, N253);
buf BUF1 (N452, N450);
nor NOR3 (N453, N436, N63, N87);
xor XOR2 (N454, N438, N84);
xor XOR2 (N455, N454, N229);
and AND3 (N456, N444, N383, N115);
or OR2 (N457, N426, N64);
nor NOR2 (N458, N448, N270);
nand NAND3 (N459, N451, N432, N260);
nor NOR4 (N460, N435, N155, N380, N96);
not NOT1 (N461, N452);
xor XOR2 (N462, N457, N90);
xor XOR2 (N463, N462, N105);
or OR3 (N464, N461, N358, N428);
and AND4 (N465, N434, N353, N347, N425);
xor XOR2 (N466, N460, N7);
nand NAND2 (N467, N463, N310);
and AND4 (N468, N467, N116, N261, N267);
nand NAND4 (N469, N456, N363, N267, N13);
nor NOR2 (N470, N464, N70);
not NOT1 (N471, N449);
buf BUF1 (N472, N458);
xor XOR2 (N473, N455, N438);
and AND3 (N474, N471, N449, N72);
xor XOR2 (N475, N474, N201);
xor XOR2 (N476, N472, N99);
nand NAND2 (N477, N468, N60);
xor XOR2 (N478, N476, N388);
nor NOR3 (N479, N478, N397, N94);
xor XOR2 (N480, N477, N194);
xor XOR2 (N481, N480, N69);
and AND4 (N482, N466, N413, N275, N373);
not NOT1 (N483, N482);
buf BUF1 (N484, N470);
and AND3 (N485, N469, N274, N259);
and AND3 (N486, N473, N50, N194);
nor NOR4 (N487, N453, N399, N447, N200);
nor NOR4 (N488, N484, N154, N191, N30);
not NOT1 (N489, N459);
buf BUF1 (N490, N488);
or OR3 (N491, N486, N259, N437);
nand NAND4 (N492, N479, N479, N478, N363);
buf BUF1 (N493, N487);
nor NOR3 (N494, N492, N142, N237);
xor XOR2 (N495, N489, N289);
xor XOR2 (N496, N491, N234);
buf BUF1 (N497, N490);
nor NOR4 (N498, N481, N12, N6, N254);
or OR2 (N499, N475, N275);
not NOT1 (N500, N498);
not NOT1 (N501, N499);
xor XOR2 (N502, N494, N250);
buf BUF1 (N503, N483);
or OR3 (N504, N496, N210, N239);
and AND2 (N505, N501, N69);
or OR4 (N506, N500, N304, N181, N48);
xor XOR2 (N507, N495, N114);
buf BUF1 (N508, N465);
nor NOR2 (N509, N503, N330);
xor XOR2 (N510, N509, N105);
and AND3 (N511, N505, N480, N161);
buf BUF1 (N512, N507);
buf BUF1 (N513, N504);
or OR2 (N514, N511, N478);
nand NAND2 (N515, N508, N413);
buf BUF1 (N516, N512);
not NOT1 (N517, N513);
or OR2 (N518, N493, N488);
not NOT1 (N519, N518);
xor XOR2 (N520, N502, N394);
xor XOR2 (N521, N506, N380);
not NOT1 (N522, N516);
nand NAND2 (N523, N497, N460);
not NOT1 (N524, N520);
nor NOR4 (N525, N485, N307, N210, N384);
nand NAND2 (N526, N510, N30);
buf BUF1 (N527, N519);
nor NOR2 (N528, N526, N143);
or OR2 (N529, N525, N376);
and AND4 (N530, N517, N156, N224, N479);
not NOT1 (N531, N523);
or OR4 (N532, N515, N142, N443, N521);
xor XOR2 (N533, N480, N468);
buf BUF1 (N534, N529);
buf BUF1 (N535, N524);
and AND2 (N536, N531, N217);
or OR3 (N537, N536, N455, N161);
xor XOR2 (N538, N534, N353);
xor XOR2 (N539, N532, N125);
nand NAND2 (N540, N533, N370);
nor NOR4 (N541, N527, N293, N209, N469);
not NOT1 (N542, N522);
not NOT1 (N543, N514);
nand NAND3 (N544, N530, N353, N395);
nor NOR2 (N545, N541, N304);
nand NAND2 (N546, N542, N163);
xor XOR2 (N547, N543, N398);
and AND2 (N548, N535, N334);
xor XOR2 (N549, N547, N89);
or OR3 (N550, N539, N263, N46);
or OR2 (N551, N544, N453);
nor NOR3 (N552, N551, N218, N303);
nand NAND2 (N553, N538, N74);
not NOT1 (N554, N537);
nand NAND2 (N555, N553, N535);
nand NAND2 (N556, N549, N490);
buf BUF1 (N557, N540);
nor NOR4 (N558, N528, N233, N258, N92);
or OR4 (N559, N550, N208, N340, N12);
not NOT1 (N560, N554);
or OR2 (N561, N557, N407);
nor NOR3 (N562, N561, N26, N51);
not NOT1 (N563, N562);
or OR3 (N564, N558, N64, N267);
nor NOR3 (N565, N564, N1, N245);
nor NOR2 (N566, N560, N504);
not NOT1 (N567, N552);
and AND3 (N568, N545, N349, N171);
nand NAND3 (N569, N556, N256, N398);
buf BUF1 (N570, N555);
and AND4 (N571, N546, N281, N389, N391);
not NOT1 (N572, N570);
or OR3 (N573, N565, N108, N182);
and AND3 (N574, N548, N315, N364);
xor XOR2 (N575, N567, N73);
xor XOR2 (N576, N563, N553);
xor XOR2 (N577, N566, N177);
nand NAND4 (N578, N574, N549, N252, N95);
nand NAND3 (N579, N573, N559, N331);
nor NOR4 (N580, N454, N11, N274, N145);
and AND3 (N581, N580, N426, N10);
not NOT1 (N582, N571);
nor NOR4 (N583, N576, N454, N172, N103);
buf BUF1 (N584, N582);
not NOT1 (N585, N579);
xor XOR2 (N586, N585, N156);
buf BUF1 (N587, N568);
nand NAND2 (N588, N577, N80);
buf BUF1 (N589, N569);
xor XOR2 (N590, N588, N563);
not NOT1 (N591, N575);
xor XOR2 (N592, N581, N459);
nand NAND2 (N593, N589, N565);
nor NOR2 (N594, N586, N58);
nand NAND4 (N595, N594, N340, N123, N468);
not NOT1 (N596, N587);
nor NOR3 (N597, N584, N503, N53);
nor NOR3 (N598, N591, N204, N213);
buf BUF1 (N599, N597);
nand NAND2 (N600, N572, N372);
and AND4 (N601, N583, N323, N436, N399);
xor XOR2 (N602, N596, N204);
or OR4 (N603, N593, N474, N439, N502);
xor XOR2 (N604, N598, N66);
and AND3 (N605, N601, N47, N569);
not NOT1 (N606, N595);
nor NOR3 (N607, N578, N349, N64);
buf BUF1 (N608, N603);
and AND2 (N609, N599, N474);
and AND3 (N610, N592, N305, N313);
xor XOR2 (N611, N590, N207);
or OR3 (N612, N609, N268, N579);
and AND4 (N613, N604, N384, N111, N321);
buf BUF1 (N614, N612);
xor XOR2 (N615, N600, N494);
not NOT1 (N616, N607);
buf BUF1 (N617, N615);
buf BUF1 (N618, N602);
xor XOR2 (N619, N611, N27);
not NOT1 (N620, N610);
xor XOR2 (N621, N613, N204);
xor XOR2 (N622, N617, N415);
nand NAND3 (N623, N606, N435, N360);
or OR4 (N624, N621, N393, N310, N352);
or OR3 (N625, N624, N486, N314);
nand NAND2 (N626, N619, N122);
and AND4 (N627, N620, N617, N78, N337);
or OR4 (N628, N625, N162, N435, N327);
and AND3 (N629, N628, N332, N607);
xor XOR2 (N630, N626, N264);
nor NOR4 (N631, N608, N586, N259, N536);
nor NOR3 (N632, N614, N206, N461);
nand NAND2 (N633, N618, N606);
nor NOR4 (N634, N629, N461, N327, N119);
xor XOR2 (N635, N634, N465);
buf BUF1 (N636, N623);
buf BUF1 (N637, N632);
nor NOR4 (N638, N631, N314, N277, N239);
not NOT1 (N639, N630);
nor NOR3 (N640, N633, N104, N495);
nor NOR4 (N641, N622, N574, N618, N186);
buf BUF1 (N642, N641);
nand NAND4 (N643, N638, N144, N610, N197);
buf BUF1 (N644, N637);
buf BUF1 (N645, N640);
and AND4 (N646, N642, N274, N252, N337);
not NOT1 (N647, N644);
buf BUF1 (N648, N639);
and AND3 (N649, N648, N434, N239);
xor XOR2 (N650, N646, N10);
buf BUF1 (N651, N645);
not NOT1 (N652, N605);
xor XOR2 (N653, N635, N109);
nand NAND4 (N654, N647, N127, N488, N403);
or OR4 (N655, N653, N435, N485, N415);
and AND4 (N656, N616, N279, N115, N21);
or OR2 (N657, N643, N628);
xor XOR2 (N658, N655, N366);
and AND2 (N659, N650, N311);
nor NOR4 (N660, N654, N24, N334, N380);
or OR2 (N661, N652, N654);
xor XOR2 (N662, N651, N660);
xor XOR2 (N663, N459, N24);
or OR4 (N664, N657, N84, N542, N77);
buf BUF1 (N665, N659);
buf BUF1 (N666, N664);
not NOT1 (N667, N661);
buf BUF1 (N668, N658);
buf BUF1 (N669, N663);
not NOT1 (N670, N662);
or OR4 (N671, N665, N40, N237, N159);
xor XOR2 (N672, N670, N520);
xor XOR2 (N673, N668, N238);
or OR2 (N674, N649, N116);
buf BUF1 (N675, N671);
nand NAND4 (N676, N669, N205, N455, N48);
not NOT1 (N677, N673);
not NOT1 (N678, N672);
not NOT1 (N679, N677);
not NOT1 (N680, N674);
nand NAND4 (N681, N636, N556, N463, N537);
nor NOR2 (N682, N676, N463);
or OR3 (N683, N681, N243, N318);
not NOT1 (N684, N627);
or OR4 (N685, N667, N43, N344, N502);
and AND3 (N686, N682, N367, N380);
not NOT1 (N687, N666);
nand NAND4 (N688, N680, N494, N62, N8);
nor NOR3 (N689, N686, N138, N160);
xor XOR2 (N690, N679, N167);
buf BUF1 (N691, N688);
nor NOR3 (N692, N656, N10, N8);
buf BUF1 (N693, N690);
nor NOR3 (N694, N678, N38, N505);
not NOT1 (N695, N685);
buf BUF1 (N696, N691);
not NOT1 (N697, N675);
or OR3 (N698, N687, N617, N412);
buf BUF1 (N699, N698);
nand NAND4 (N700, N697, N629, N459, N24);
or OR3 (N701, N700, N253, N517);
nand NAND3 (N702, N696, N29, N62);
or OR4 (N703, N701, N363, N685, N481);
or OR4 (N704, N703, N102, N672, N508);
nor NOR3 (N705, N684, N579, N360);
nand NAND4 (N706, N693, N375, N425, N421);
nor NOR2 (N707, N706, N372);
buf BUF1 (N708, N699);
buf BUF1 (N709, N692);
buf BUF1 (N710, N704);
xor XOR2 (N711, N689, N498);
buf BUF1 (N712, N705);
buf BUF1 (N713, N711);
nor NOR3 (N714, N695, N434, N3);
or OR3 (N715, N712, N387, N583);
and AND3 (N716, N694, N481, N242);
or OR3 (N717, N707, N133, N34);
buf BUF1 (N718, N715);
and AND4 (N719, N714, N438, N146, N254);
xor XOR2 (N720, N683, N485);
xor XOR2 (N721, N708, N497);
or OR4 (N722, N710, N132, N355, N109);
not NOT1 (N723, N702);
xor XOR2 (N724, N722, N467);
buf BUF1 (N725, N709);
buf BUF1 (N726, N719);
or OR2 (N727, N713, N574);
buf BUF1 (N728, N721);
not NOT1 (N729, N718);
nor NOR3 (N730, N726, N544, N546);
or OR4 (N731, N720, N660, N182, N72);
nand NAND4 (N732, N731, N475, N606, N352);
and AND2 (N733, N724, N646);
or OR4 (N734, N730, N294, N732, N639);
not NOT1 (N735, N248);
and AND2 (N736, N733, N156);
not NOT1 (N737, N716);
or OR4 (N738, N727, N651, N600, N28);
not NOT1 (N739, N728);
and AND4 (N740, N736, N487, N88, N529);
buf BUF1 (N741, N717);
and AND2 (N742, N741, N367);
nor NOR2 (N743, N742, N157);
or OR3 (N744, N729, N143, N192);
buf BUF1 (N745, N735);
nand NAND2 (N746, N740, N337);
xor XOR2 (N747, N737, N660);
not NOT1 (N748, N747);
not NOT1 (N749, N738);
and AND4 (N750, N748, N480, N273, N548);
and AND4 (N751, N749, N443, N689, N427);
nor NOR2 (N752, N750, N387);
and AND3 (N753, N734, N524, N368);
and AND4 (N754, N725, N253, N721, N429);
buf BUF1 (N755, N743);
xor XOR2 (N756, N752, N317);
xor XOR2 (N757, N739, N662);
nor NOR3 (N758, N754, N152, N399);
and AND2 (N759, N757, N47);
nand NAND3 (N760, N759, N683, N310);
xor XOR2 (N761, N723, N602);
or OR4 (N762, N761, N164, N321, N165);
not NOT1 (N763, N753);
nand NAND2 (N764, N763, N539);
buf BUF1 (N765, N764);
nand NAND2 (N766, N758, N551);
buf BUF1 (N767, N751);
xor XOR2 (N768, N767, N487);
and AND2 (N769, N766, N605);
and AND3 (N770, N755, N551, N566);
and AND3 (N771, N770, N157, N642);
buf BUF1 (N772, N771);
nand NAND3 (N773, N769, N175, N471);
nor NOR3 (N774, N745, N256, N742);
and AND3 (N775, N760, N533, N451);
not NOT1 (N776, N762);
nor NOR2 (N777, N775, N383);
not NOT1 (N778, N744);
xor XOR2 (N779, N778, N31);
and AND3 (N780, N774, N484, N560);
buf BUF1 (N781, N773);
xor XOR2 (N782, N772, N355);
nand NAND4 (N783, N768, N776, N591, N726);
or OR4 (N784, N91, N343, N298, N432);
buf BUF1 (N785, N779);
nor NOR3 (N786, N765, N687, N645);
xor XOR2 (N787, N746, N703);
and AND2 (N788, N785, N57);
buf BUF1 (N789, N788);
not NOT1 (N790, N777);
nor NOR4 (N791, N784, N33, N656, N344);
nor NOR4 (N792, N781, N414, N76, N130);
buf BUF1 (N793, N756);
and AND2 (N794, N789, N424);
or OR2 (N795, N794, N750);
nand NAND3 (N796, N791, N246, N309);
nor NOR2 (N797, N796, N598);
and AND4 (N798, N792, N294, N353, N566);
xor XOR2 (N799, N790, N303);
xor XOR2 (N800, N787, N750);
xor XOR2 (N801, N800, N253);
nand NAND2 (N802, N797, N337);
buf BUF1 (N803, N798);
xor XOR2 (N804, N782, N695);
buf BUF1 (N805, N786);
or OR2 (N806, N803, N65);
or OR2 (N807, N806, N631);
and AND2 (N808, N804, N254);
and AND2 (N809, N793, N675);
or OR2 (N810, N805, N771);
and AND3 (N811, N809, N239, N599);
nand NAND2 (N812, N783, N614);
nand NAND3 (N813, N795, N11, N764);
xor XOR2 (N814, N799, N411);
endmodule