// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N3004,N3009,N3008,N3001,N3000,N3007,N3002,N2991,N2992,N3010;

buf BUF1 (N11, N1);
or OR2 (N12, N6, N6);
nand NAND3 (N13, N2, N7, N6);
xor XOR2 (N14, N11, N9);
buf BUF1 (N15, N4);
xor XOR2 (N16, N8, N4);
nor NOR2 (N17, N9, N1);
nor NOR3 (N18, N2, N3, N1);
xor XOR2 (N19, N12, N13);
not NOT1 (N20, N8);
or OR2 (N21, N20, N7);
buf BUF1 (N22, N6);
nor NOR3 (N23, N3, N12, N20);
not NOT1 (N24, N5);
nor NOR2 (N25, N22, N15);
or OR2 (N26, N14, N24);
nand NAND3 (N27, N19, N19, N15);
xor XOR2 (N28, N6, N21);
or OR2 (N29, N13, N28);
and AND4 (N30, N1, N9, N24, N20);
or OR2 (N31, N21, N19);
not NOT1 (N32, N17);
nor NOR2 (N33, N26, N21);
nor NOR3 (N34, N23, N12, N28);
not NOT1 (N35, N32);
nor NOR2 (N36, N33, N19);
or OR2 (N37, N16, N6);
and AND2 (N38, N35, N23);
xor XOR2 (N39, N36, N13);
not NOT1 (N40, N31);
or OR4 (N41, N39, N15, N7, N14);
xor XOR2 (N42, N38, N2);
buf BUF1 (N43, N30);
nor NOR3 (N44, N27, N9, N22);
xor XOR2 (N45, N18, N9);
not NOT1 (N46, N41);
xor XOR2 (N47, N34, N13);
or OR3 (N48, N40, N45, N13);
xor XOR2 (N49, N24, N23);
nand NAND4 (N50, N46, N33, N43, N44);
nor NOR3 (N51, N44, N46, N10);
xor XOR2 (N52, N45, N43);
or OR2 (N53, N52, N40);
not NOT1 (N54, N25);
or OR3 (N55, N37, N2, N52);
not NOT1 (N56, N50);
buf BUF1 (N57, N56);
buf BUF1 (N58, N55);
or OR2 (N59, N53, N35);
and AND2 (N60, N57, N27);
buf BUF1 (N61, N29);
nand NAND3 (N62, N58, N61, N37);
xor XOR2 (N63, N24, N58);
nand NAND2 (N64, N48, N21);
buf BUF1 (N65, N60);
and AND4 (N66, N51, N24, N34, N52);
or OR3 (N67, N65, N44, N41);
xor XOR2 (N68, N49, N3);
not NOT1 (N69, N42);
nand NAND3 (N70, N59, N41, N17);
not NOT1 (N71, N54);
nor NOR3 (N72, N67, N40, N50);
nor NOR3 (N73, N70, N19, N19);
not NOT1 (N74, N68);
xor XOR2 (N75, N72, N34);
nor NOR2 (N76, N64, N42);
xor XOR2 (N77, N66, N52);
nor NOR4 (N78, N63, N42, N46, N69);
buf BUF1 (N79, N34);
nor NOR3 (N80, N62, N36, N75);
nor NOR2 (N81, N63, N24);
nor NOR3 (N82, N47, N43, N30);
not NOT1 (N83, N76);
and AND3 (N84, N80, N73, N71);
not NOT1 (N85, N73);
and AND4 (N86, N23, N42, N63, N22);
or OR4 (N87, N77, N73, N37, N50);
buf BUF1 (N88, N87);
xor XOR2 (N89, N82, N50);
buf BUF1 (N90, N81);
and AND3 (N91, N83, N81, N90);
buf BUF1 (N92, N39);
buf BUF1 (N93, N91);
nor NOR4 (N94, N74, N42, N53, N13);
xor XOR2 (N95, N79, N62);
buf BUF1 (N96, N78);
nand NAND2 (N97, N88, N62);
and AND2 (N98, N95, N66);
not NOT1 (N99, N84);
nand NAND4 (N100, N94, N79, N66, N16);
and AND4 (N101, N86, N14, N74, N8);
buf BUF1 (N102, N96);
nor NOR2 (N103, N101, N99);
and AND3 (N104, N87, N4, N48);
xor XOR2 (N105, N102, N18);
not NOT1 (N106, N100);
or OR2 (N107, N89, N7);
nand NAND3 (N108, N104, N103, N64);
buf BUF1 (N109, N93);
nand NAND4 (N110, N71, N2, N93, N109);
or OR2 (N111, N52, N12);
nand NAND2 (N112, N107, N92);
nand NAND3 (N113, N1, N16, N42);
and AND2 (N114, N105, N67);
buf BUF1 (N115, N111);
buf BUF1 (N116, N108);
buf BUF1 (N117, N98);
or OR3 (N118, N112, N8, N97);
and AND4 (N119, N73, N42, N20, N75);
or OR4 (N120, N113, N98, N91, N25);
nor NOR4 (N121, N118, N100, N113, N102);
not NOT1 (N122, N120);
buf BUF1 (N123, N114);
and AND2 (N124, N122, N81);
buf BUF1 (N125, N119);
buf BUF1 (N126, N106);
nor NOR2 (N127, N116, N92);
nand NAND4 (N128, N121, N124, N60, N62);
and AND3 (N129, N51, N108, N120);
nor NOR2 (N130, N110, N116);
nand NAND4 (N131, N85, N87, N84, N66);
xor XOR2 (N132, N130, N70);
nor NOR2 (N133, N126, N100);
xor XOR2 (N134, N129, N86);
buf BUF1 (N135, N131);
nor NOR3 (N136, N132, N65, N3);
buf BUF1 (N137, N133);
buf BUF1 (N138, N127);
or OR2 (N139, N117, N93);
nand NAND4 (N140, N136, N122, N106, N32);
nor NOR3 (N141, N134, N48, N80);
nor NOR4 (N142, N123, N41, N80, N138);
buf BUF1 (N143, N69);
xor XOR2 (N144, N135, N44);
not NOT1 (N145, N143);
not NOT1 (N146, N139);
and AND4 (N147, N142, N14, N76, N35);
or OR4 (N148, N137, N126, N25, N108);
nand NAND3 (N149, N144, N40, N101);
not NOT1 (N150, N146);
xor XOR2 (N151, N148, N43);
not NOT1 (N152, N145);
xor XOR2 (N153, N141, N132);
not NOT1 (N154, N151);
xor XOR2 (N155, N150, N137);
not NOT1 (N156, N153);
not NOT1 (N157, N115);
buf BUF1 (N158, N125);
nor NOR4 (N159, N152, N141, N23, N107);
nor NOR2 (N160, N159, N144);
not NOT1 (N161, N154);
nor NOR2 (N162, N140, N106);
and AND2 (N163, N149, N91);
nor NOR4 (N164, N155, N38, N88, N23);
xor XOR2 (N165, N163, N112);
nor NOR4 (N166, N147, N155, N107, N128);
nor NOR3 (N167, N14, N139, N94);
nor NOR2 (N168, N160, N34);
or OR4 (N169, N168, N124, N109, N112);
nand NAND3 (N170, N161, N61, N111);
nor NOR4 (N171, N162, N6, N68, N32);
nor NOR3 (N172, N167, N115, N46);
nand NAND3 (N173, N170, N59, N56);
not NOT1 (N174, N169);
nor NOR3 (N175, N172, N73, N59);
xor XOR2 (N176, N164, N146);
or OR3 (N177, N173, N22, N140);
nor NOR2 (N178, N157, N42);
nand NAND3 (N179, N174, N140, N144);
and AND2 (N180, N179, N53);
and AND4 (N181, N158, N87, N116, N155);
or OR2 (N182, N175, N174);
buf BUF1 (N183, N180);
xor XOR2 (N184, N176, N162);
buf BUF1 (N185, N181);
and AND4 (N186, N165, N160, N66, N28);
nor NOR3 (N187, N177, N150, N104);
xor XOR2 (N188, N171, N56);
or OR3 (N189, N182, N28, N26);
nand NAND2 (N190, N188, N111);
xor XOR2 (N191, N178, N88);
not NOT1 (N192, N185);
buf BUF1 (N193, N192);
and AND2 (N194, N156, N120);
or OR3 (N195, N184, N193, N110);
and AND3 (N196, N150, N166, N116);
xor XOR2 (N197, N8, N144);
nand NAND3 (N198, N186, N105, N14);
nor NOR3 (N199, N189, N18, N11);
not NOT1 (N200, N191);
nor NOR4 (N201, N197, N199, N33, N157);
not NOT1 (N202, N47);
not NOT1 (N203, N196);
nand NAND2 (N204, N183, N94);
nand NAND3 (N205, N201, N70, N111);
nor NOR3 (N206, N203, N137, N49);
buf BUF1 (N207, N200);
nand NAND3 (N208, N204, N23, N183);
not NOT1 (N209, N206);
and AND4 (N210, N194, N65, N196, N129);
and AND2 (N211, N195, N29);
nand NAND2 (N212, N207, N156);
not NOT1 (N213, N190);
not NOT1 (N214, N212);
not NOT1 (N215, N209);
and AND4 (N216, N211, N60, N13, N41);
and AND4 (N217, N210, N34, N34, N36);
not NOT1 (N218, N215);
and AND3 (N219, N202, N142, N85);
buf BUF1 (N220, N213);
and AND3 (N221, N208, N143, N141);
or OR3 (N222, N216, N38, N31);
or OR2 (N223, N222, N87);
or OR4 (N224, N198, N71, N20, N7);
and AND2 (N225, N219, N33);
nand NAND3 (N226, N221, N52, N99);
nor NOR2 (N227, N187, N91);
or OR4 (N228, N220, N83, N144, N135);
xor XOR2 (N229, N228, N119);
or OR3 (N230, N218, N105, N123);
and AND2 (N231, N230, N38);
or OR3 (N232, N229, N188, N150);
not NOT1 (N233, N227);
and AND2 (N234, N233, N81);
buf BUF1 (N235, N231);
nor NOR3 (N236, N234, N129, N32);
nor NOR4 (N237, N224, N200, N121, N101);
and AND3 (N238, N237, N204, N89);
buf BUF1 (N239, N214);
xor XOR2 (N240, N239, N19);
nor NOR4 (N241, N205, N22, N74, N158);
or OR3 (N242, N235, N40, N31);
not NOT1 (N243, N236);
nor NOR2 (N244, N223, N230);
nor NOR4 (N245, N238, N203, N202, N193);
nand NAND3 (N246, N241, N46, N76);
xor XOR2 (N247, N245, N175);
buf BUF1 (N248, N246);
nor NOR2 (N249, N242, N193);
or OR2 (N250, N225, N233);
and AND3 (N251, N250, N193, N30);
xor XOR2 (N252, N217, N105);
xor XOR2 (N253, N244, N186);
buf BUF1 (N254, N248);
not NOT1 (N255, N249);
xor XOR2 (N256, N240, N156);
xor XOR2 (N257, N251, N205);
nor NOR4 (N258, N232, N92, N241, N42);
buf BUF1 (N259, N253);
buf BUF1 (N260, N247);
nand NAND3 (N261, N252, N20, N27);
or OR4 (N262, N258, N103, N237, N181);
nor NOR4 (N263, N226, N116, N8, N244);
and AND3 (N264, N254, N56, N127);
and AND4 (N265, N260, N91, N111, N96);
not NOT1 (N266, N243);
xor XOR2 (N267, N261, N204);
nor NOR3 (N268, N264, N14, N250);
xor XOR2 (N269, N262, N255);
xor XOR2 (N270, N167, N82);
not NOT1 (N271, N267);
xor XOR2 (N272, N259, N137);
or OR4 (N273, N272, N112, N107, N114);
or OR2 (N274, N263, N260);
and AND2 (N275, N273, N183);
xor XOR2 (N276, N257, N207);
buf BUF1 (N277, N271);
xor XOR2 (N278, N268, N116);
nand NAND4 (N279, N276, N21, N60, N148);
buf BUF1 (N280, N277);
buf BUF1 (N281, N275);
or OR4 (N282, N274, N96, N120, N122);
not NOT1 (N283, N282);
nand NAND4 (N284, N283, N172, N235, N156);
and AND2 (N285, N265, N6);
xor XOR2 (N286, N281, N192);
buf BUF1 (N287, N284);
xor XOR2 (N288, N256, N48);
nand NAND2 (N289, N285, N245);
buf BUF1 (N290, N280);
nor NOR4 (N291, N289, N269, N106, N185);
and AND3 (N292, N179, N149, N39);
buf BUF1 (N293, N291);
nand NAND4 (N294, N293, N84, N229, N172);
xor XOR2 (N295, N286, N255);
nand NAND4 (N296, N278, N35, N14, N149);
nor NOR3 (N297, N295, N292, N165);
nand NAND3 (N298, N283, N174, N28);
and AND3 (N299, N279, N132, N170);
and AND3 (N300, N297, N65, N17);
nand NAND4 (N301, N287, N141, N142, N2);
xor XOR2 (N302, N296, N71);
nand NAND3 (N303, N298, N162, N49);
and AND4 (N304, N288, N270, N120, N3);
nor NOR4 (N305, N268, N52, N48, N163);
xor XOR2 (N306, N304, N117);
xor XOR2 (N307, N302, N291);
nor NOR2 (N308, N301, N127);
nand NAND3 (N309, N305, N21, N229);
and AND4 (N310, N308, N86, N95, N75);
or OR3 (N311, N309, N274, N69);
or OR4 (N312, N299, N184, N130, N223);
not NOT1 (N313, N310);
and AND4 (N314, N294, N104, N69, N120);
or OR4 (N315, N313, N79, N37, N277);
and AND3 (N316, N307, N129, N65);
nand NAND2 (N317, N290, N9);
nand NAND3 (N318, N315, N158, N146);
buf BUF1 (N319, N314);
buf BUF1 (N320, N300);
nand NAND2 (N321, N303, N249);
xor XOR2 (N322, N316, N82);
nor NOR4 (N323, N266, N136, N42, N62);
buf BUF1 (N324, N318);
xor XOR2 (N325, N317, N54);
xor XOR2 (N326, N322, N161);
xor XOR2 (N327, N320, N268);
xor XOR2 (N328, N326, N20);
not NOT1 (N329, N323);
not NOT1 (N330, N319);
or OR4 (N331, N327, N188, N90, N297);
nand NAND2 (N332, N331, N57);
and AND4 (N333, N324, N13, N101, N82);
nor NOR3 (N334, N312, N259, N165);
buf BUF1 (N335, N311);
not NOT1 (N336, N321);
or OR2 (N337, N336, N15);
nor NOR3 (N338, N335, N85, N120);
nand NAND4 (N339, N337, N82, N164, N255);
nand NAND4 (N340, N325, N3, N228, N286);
or OR2 (N341, N332, N167);
and AND2 (N342, N328, N272);
nor NOR2 (N343, N342, N206);
not NOT1 (N344, N341);
not NOT1 (N345, N339);
and AND2 (N346, N338, N47);
xor XOR2 (N347, N329, N73);
xor XOR2 (N348, N333, N212);
and AND4 (N349, N340, N326, N50, N12);
nand NAND3 (N350, N345, N246, N195);
or OR4 (N351, N350, N348, N34, N217);
or OR3 (N352, N329, N220, N315);
not NOT1 (N353, N346);
or OR4 (N354, N353, N165, N52, N32);
and AND3 (N355, N351, N318, N295);
buf BUF1 (N356, N334);
buf BUF1 (N357, N330);
nand NAND3 (N358, N355, N239, N74);
nand NAND3 (N359, N306, N1, N233);
xor XOR2 (N360, N343, N43);
or OR4 (N361, N356, N344, N151, N2);
not NOT1 (N362, N276);
nand NAND3 (N363, N360, N266, N177);
buf BUF1 (N364, N354);
buf BUF1 (N365, N361);
and AND2 (N366, N365, N298);
or OR3 (N367, N352, N229, N82);
and AND3 (N368, N364, N217, N211);
nor NOR4 (N369, N349, N315, N287, N153);
xor XOR2 (N370, N347, N340);
nand NAND4 (N371, N362, N144, N179, N37);
not NOT1 (N372, N368);
and AND3 (N373, N370, N261, N125);
buf BUF1 (N374, N363);
nand NAND4 (N375, N358, N177, N213, N209);
or OR2 (N376, N372, N346);
buf BUF1 (N377, N371);
nand NAND4 (N378, N376, N57, N256, N310);
buf BUF1 (N379, N366);
nand NAND3 (N380, N379, N134, N362);
nor NOR2 (N381, N377, N200);
nor NOR2 (N382, N375, N247);
or OR4 (N383, N382, N150, N137, N303);
nand NAND3 (N384, N380, N343, N206);
buf BUF1 (N385, N381);
not NOT1 (N386, N373);
and AND2 (N387, N367, N211);
and AND3 (N388, N374, N94, N279);
xor XOR2 (N389, N385, N201);
nor NOR2 (N390, N387, N327);
xor XOR2 (N391, N369, N224);
and AND4 (N392, N378, N193, N27, N73);
xor XOR2 (N393, N357, N194);
xor XOR2 (N394, N384, N263);
or OR4 (N395, N393, N38, N99, N210);
nand NAND2 (N396, N394, N271);
or OR2 (N397, N391, N248);
not NOT1 (N398, N386);
not NOT1 (N399, N359);
or OR4 (N400, N392, N4, N230, N146);
and AND3 (N401, N390, N221, N120);
or OR2 (N402, N395, N334);
nor NOR3 (N403, N397, N395, N45);
not NOT1 (N404, N399);
and AND3 (N405, N402, N122, N132);
not NOT1 (N406, N388);
nor NOR2 (N407, N403, N217);
xor XOR2 (N408, N406, N122);
buf BUF1 (N409, N404);
nand NAND2 (N410, N383, N189);
not NOT1 (N411, N409);
nor NOR4 (N412, N389, N291, N189, N93);
xor XOR2 (N413, N396, N322);
xor XOR2 (N414, N412, N314);
xor XOR2 (N415, N398, N133);
nand NAND2 (N416, N415, N354);
not NOT1 (N417, N414);
nor NOR3 (N418, N413, N24, N172);
and AND3 (N419, N407, N57, N25);
and AND4 (N420, N418, N305, N30, N161);
buf BUF1 (N421, N420);
and AND3 (N422, N419, N140, N409);
nor NOR2 (N423, N400, N352);
not NOT1 (N424, N411);
buf BUF1 (N425, N416);
not NOT1 (N426, N401);
or OR3 (N427, N424, N198, N258);
xor XOR2 (N428, N421, N178);
nand NAND4 (N429, N422, N96, N29, N312);
and AND3 (N430, N417, N328, N105);
not NOT1 (N431, N423);
not NOT1 (N432, N430);
nand NAND3 (N433, N431, N353, N62);
not NOT1 (N434, N408);
xor XOR2 (N435, N427, N117);
or OR3 (N436, N410, N310, N213);
xor XOR2 (N437, N428, N415);
xor XOR2 (N438, N405, N358);
and AND3 (N439, N435, N135, N169);
xor XOR2 (N440, N439, N62);
nor NOR3 (N441, N426, N253, N76);
nor NOR2 (N442, N433, N343);
or OR3 (N443, N442, N401, N422);
and AND2 (N444, N438, N74);
xor XOR2 (N445, N425, N179);
xor XOR2 (N446, N443, N27);
and AND2 (N447, N436, N174);
and AND2 (N448, N446, N67);
xor XOR2 (N449, N434, N205);
nand NAND2 (N450, N440, N418);
buf BUF1 (N451, N447);
and AND3 (N452, N429, N414, N187);
nand NAND4 (N453, N437, N28, N38, N8);
not NOT1 (N454, N441);
buf BUF1 (N455, N450);
or OR4 (N456, N449, N148, N329, N309);
not NOT1 (N457, N454);
buf BUF1 (N458, N452);
or OR2 (N459, N457, N224);
buf BUF1 (N460, N448);
xor XOR2 (N461, N432, N260);
and AND4 (N462, N451, N442, N331, N363);
not NOT1 (N463, N456);
nor NOR3 (N464, N459, N446, N447);
or OR4 (N465, N464, N239, N284, N86);
buf BUF1 (N466, N453);
not NOT1 (N467, N461);
or OR4 (N468, N465, N450, N358, N187);
buf BUF1 (N469, N462);
buf BUF1 (N470, N444);
and AND4 (N471, N470, N190, N289, N168);
not NOT1 (N472, N471);
nor NOR3 (N473, N445, N373, N395);
and AND2 (N474, N463, N153);
nand NAND3 (N475, N458, N302, N19);
buf BUF1 (N476, N472);
nor NOR3 (N477, N455, N142, N444);
nand NAND3 (N478, N469, N444, N225);
buf BUF1 (N479, N473);
not NOT1 (N480, N476);
nor NOR3 (N481, N460, N93, N14);
or OR4 (N482, N477, N377, N393, N336);
nand NAND2 (N483, N474, N30);
buf BUF1 (N484, N483);
xor XOR2 (N485, N475, N64);
buf BUF1 (N486, N479);
nand NAND2 (N487, N480, N123);
buf BUF1 (N488, N466);
buf BUF1 (N489, N487);
not NOT1 (N490, N485);
nand NAND4 (N491, N481, N95, N7, N385);
and AND3 (N492, N484, N435, N149);
nor NOR4 (N493, N467, N417, N4, N9);
nor NOR2 (N494, N493, N410);
nor NOR2 (N495, N494, N110);
buf BUF1 (N496, N486);
nor NOR4 (N497, N482, N474, N465, N282);
buf BUF1 (N498, N491);
nor NOR2 (N499, N495, N339);
nand NAND2 (N500, N498, N284);
and AND4 (N501, N497, N75, N16, N479);
nor NOR3 (N502, N501, N274, N456);
not NOT1 (N503, N488);
or OR2 (N504, N490, N217);
xor XOR2 (N505, N504, N370);
xor XOR2 (N506, N502, N349);
and AND3 (N507, N489, N364, N285);
not NOT1 (N508, N496);
nor NOR2 (N509, N503, N294);
nand NAND4 (N510, N492, N132, N390, N129);
not NOT1 (N511, N499);
xor XOR2 (N512, N478, N200);
not NOT1 (N513, N507);
or OR4 (N514, N500, N78, N173, N310);
and AND3 (N515, N509, N108, N279);
nor NOR4 (N516, N513, N493, N334, N120);
not NOT1 (N517, N468);
or OR3 (N518, N508, N482, N233);
not NOT1 (N519, N510);
nor NOR2 (N520, N514, N159);
xor XOR2 (N521, N519, N2);
buf BUF1 (N522, N512);
nand NAND2 (N523, N506, N418);
not NOT1 (N524, N518);
and AND2 (N525, N524, N388);
nand NAND4 (N526, N516, N98, N331, N489);
nor NOR4 (N527, N517, N356, N346, N362);
and AND4 (N528, N523, N475, N209, N473);
and AND3 (N529, N521, N75, N176);
and AND3 (N530, N528, N154, N171);
buf BUF1 (N531, N522);
nand NAND3 (N532, N515, N161, N505);
nor NOR3 (N533, N153, N493, N113);
nand NAND4 (N534, N532, N392, N93, N318);
and AND3 (N535, N531, N68, N180);
or OR3 (N536, N529, N95, N340);
not NOT1 (N537, N526);
not NOT1 (N538, N511);
buf BUF1 (N539, N538);
and AND3 (N540, N535, N143, N472);
or OR3 (N541, N527, N45, N260);
xor XOR2 (N542, N525, N239);
and AND3 (N543, N539, N327, N71);
or OR4 (N544, N543, N126, N51, N156);
or OR4 (N545, N541, N110, N246, N411);
nand NAND4 (N546, N540, N277, N420, N73);
xor XOR2 (N547, N520, N310);
and AND4 (N548, N545, N446, N123, N413);
nor NOR3 (N549, N546, N102, N285);
nor NOR3 (N550, N533, N203, N180);
not NOT1 (N551, N534);
or OR4 (N552, N536, N55, N479, N512);
or OR2 (N553, N542, N34);
and AND4 (N554, N548, N39, N212, N400);
and AND3 (N555, N553, N229, N224);
buf BUF1 (N556, N537);
buf BUF1 (N557, N530);
nand NAND2 (N558, N556, N399);
nand NAND2 (N559, N555, N397);
not NOT1 (N560, N552);
and AND2 (N561, N549, N320);
and AND2 (N562, N560, N413);
and AND3 (N563, N559, N493, N51);
and AND2 (N564, N557, N545);
buf BUF1 (N565, N544);
and AND4 (N566, N550, N334, N252, N311);
or OR2 (N567, N564, N180);
not NOT1 (N568, N562);
xor XOR2 (N569, N568, N340);
and AND3 (N570, N563, N267, N317);
nor NOR4 (N571, N554, N540, N183, N136);
xor XOR2 (N572, N570, N422);
nand NAND3 (N573, N572, N515, N393);
nor NOR4 (N574, N569, N480, N77, N115);
buf BUF1 (N575, N566);
buf BUF1 (N576, N575);
or OR2 (N577, N567, N313);
or OR4 (N578, N551, N10, N163, N362);
nand NAND3 (N579, N576, N487, N562);
nor NOR3 (N580, N578, N54, N32);
or OR3 (N581, N577, N482, N454);
or OR4 (N582, N574, N199, N44, N393);
nor NOR2 (N583, N580, N259);
and AND4 (N584, N565, N538, N141, N40);
or OR2 (N585, N579, N455);
and AND2 (N586, N558, N544);
or OR4 (N587, N561, N516, N556, N268);
xor XOR2 (N588, N571, N314);
and AND4 (N589, N587, N318, N277, N454);
or OR2 (N590, N585, N37);
not NOT1 (N591, N583);
buf BUF1 (N592, N547);
nand NAND4 (N593, N581, N34, N166, N213);
nand NAND3 (N594, N589, N499, N581);
xor XOR2 (N595, N582, N301);
nand NAND3 (N596, N592, N223, N310);
nor NOR3 (N597, N586, N126, N1);
nand NAND3 (N598, N596, N200, N551);
buf BUF1 (N599, N588);
not NOT1 (N600, N594);
nor NOR3 (N601, N595, N1, N127);
nand NAND3 (N602, N598, N145, N449);
nor NOR2 (N603, N602, N531);
and AND4 (N604, N573, N387, N193, N416);
buf BUF1 (N605, N597);
nor NOR4 (N606, N599, N285, N264, N412);
buf BUF1 (N607, N591);
and AND2 (N608, N605, N338);
nand NAND3 (N609, N601, N305, N405);
xor XOR2 (N610, N600, N16);
not NOT1 (N611, N590);
xor XOR2 (N612, N608, N545);
buf BUF1 (N613, N593);
nand NAND4 (N614, N584, N208, N142, N298);
nand NAND2 (N615, N613, N31);
or OR2 (N616, N604, N287);
nand NAND2 (N617, N612, N172);
nand NAND2 (N618, N616, N317);
or OR4 (N619, N615, N447, N236, N106);
nand NAND2 (N620, N606, N111);
or OR2 (N621, N611, N545);
xor XOR2 (N622, N609, N587);
nor NOR3 (N623, N619, N130, N440);
or OR2 (N624, N618, N77);
and AND2 (N625, N621, N306);
not NOT1 (N626, N622);
nand NAND3 (N627, N603, N315, N626);
and AND4 (N628, N280, N111, N617, N269);
xor XOR2 (N629, N153, N22);
xor XOR2 (N630, N628, N533);
or OR4 (N631, N607, N571, N298, N192);
buf BUF1 (N632, N627);
nor NOR2 (N633, N632, N595);
nor NOR4 (N634, N624, N1, N620, N58);
or OR2 (N635, N344, N141);
buf BUF1 (N636, N625);
or OR2 (N637, N630, N465);
not NOT1 (N638, N629);
nor NOR2 (N639, N633, N313);
not NOT1 (N640, N631);
xor XOR2 (N641, N639, N367);
buf BUF1 (N642, N641);
nand NAND2 (N643, N637, N322);
and AND2 (N644, N638, N571);
buf BUF1 (N645, N635);
not NOT1 (N646, N640);
not NOT1 (N647, N636);
and AND2 (N648, N645, N9);
not NOT1 (N649, N642);
or OR4 (N650, N643, N285, N244, N100);
nor NOR3 (N651, N649, N150, N32);
not NOT1 (N652, N610);
xor XOR2 (N653, N648, N184);
not NOT1 (N654, N646);
not NOT1 (N655, N644);
buf BUF1 (N656, N653);
and AND3 (N657, N656, N67, N538);
buf BUF1 (N658, N651);
buf BUF1 (N659, N652);
or OR4 (N660, N659, N4, N300, N358);
xor XOR2 (N661, N658, N319);
buf BUF1 (N662, N654);
xor XOR2 (N663, N634, N378);
buf BUF1 (N664, N662);
xor XOR2 (N665, N664, N355);
xor XOR2 (N666, N660, N213);
xor XOR2 (N667, N647, N646);
or OR3 (N668, N661, N27, N658);
nor NOR4 (N669, N650, N127, N509, N111);
buf BUF1 (N670, N623);
xor XOR2 (N671, N665, N13);
xor XOR2 (N672, N663, N242);
xor XOR2 (N673, N672, N608);
nor NOR3 (N674, N671, N564, N175);
xor XOR2 (N675, N670, N277);
buf BUF1 (N676, N668);
nor NOR2 (N677, N667, N409);
buf BUF1 (N678, N666);
xor XOR2 (N679, N676, N106);
or OR4 (N680, N677, N25, N312, N88);
or OR3 (N681, N669, N207, N465);
not NOT1 (N682, N681);
not NOT1 (N683, N655);
nor NOR4 (N684, N678, N171, N630, N337);
or OR4 (N685, N673, N670, N86, N78);
or OR2 (N686, N674, N197);
xor XOR2 (N687, N680, N67);
nand NAND4 (N688, N687, N179, N149, N641);
not NOT1 (N689, N675);
and AND2 (N690, N686, N441);
or OR2 (N691, N614, N104);
xor XOR2 (N692, N689, N67);
xor XOR2 (N693, N682, N14);
xor XOR2 (N694, N690, N521);
xor XOR2 (N695, N684, N158);
or OR4 (N696, N691, N674, N249, N490);
buf BUF1 (N697, N694);
and AND2 (N698, N685, N679);
nand NAND3 (N699, N489, N228, N591);
or OR3 (N700, N698, N501, N661);
not NOT1 (N701, N697);
nand NAND2 (N702, N695, N23);
nor NOR4 (N703, N699, N16, N578, N293);
and AND3 (N704, N702, N28, N612);
nor NOR3 (N705, N688, N298, N103);
or OR2 (N706, N701, N476);
or OR3 (N707, N706, N124, N297);
nand NAND2 (N708, N657, N177);
not NOT1 (N709, N692);
xor XOR2 (N710, N683, N594);
or OR4 (N711, N700, N188, N569, N433);
not NOT1 (N712, N711);
nor NOR4 (N713, N703, N413, N544, N393);
nor NOR4 (N714, N712, N429, N408, N104);
or OR2 (N715, N704, N129);
buf BUF1 (N716, N705);
not NOT1 (N717, N693);
and AND4 (N718, N714, N60, N183, N166);
and AND4 (N719, N710, N660, N593, N671);
xor XOR2 (N720, N709, N179);
or OR4 (N721, N713, N691, N447, N684);
buf BUF1 (N722, N717);
not NOT1 (N723, N707);
xor XOR2 (N724, N708, N54);
xor XOR2 (N725, N715, N282);
or OR4 (N726, N718, N1, N451, N550);
not NOT1 (N727, N719);
buf BUF1 (N728, N716);
buf BUF1 (N729, N723);
not NOT1 (N730, N727);
buf BUF1 (N731, N728);
xor XOR2 (N732, N721, N98);
not NOT1 (N733, N726);
xor XOR2 (N734, N730, N366);
not NOT1 (N735, N725);
not NOT1 (N736, N696);
nand NAND2 (N737, N735, N108);
and AND2 (N738, N732, N128);
buf BUF1 (N739, N737);
not NOT1 (N740, N734);
and AND4 (N741, N731, N466, N442, N725);
and AND4 (N742, N720, N716, N112, N155);
buf BUF1 (N743, N741);
not NOT1 (N744, N740);
and AND2 (N745, N733, N618);
nand NAND3 (N746, N736, N623, N601);
buf BUF1 (N747, N745);
nor NOR3 (N748, N743, N559, N111);
nand NAND3 (N749, N747, N174, N581);
nor NOR3 (N750, N724, N77, N626);
xor XOR2 (N751, N722, N470);
or OR2 (N752, N738, N578);
nand NAND2 (N753, N751, N13);
not NOT1 (N754, N746);
nand NAND4 (N755, N748, N353, N752, N567);
and AND4 (N756, N491, N301, N604, N656);
or OR3 (N757, N753, N652, N419);
buf BUF1 (N758, N755);
not NOT1 (N759, N758);
nor NOR2 (N760, N759, N237);
nor NOR4 (N761, N760, N90, N250, N408);
or OR2 (N762, N742, N516);
xor XOR2 (N763, N754, N545);
nor NOR3 (N764, N744, N324, N26);
nor NOR4 (N765, N749, N523, N574, N178);
not NOT1 (N766, N765);
nor NOR4 (N767, N764, N693, N118, N460);
buf BUF1 (N768, N761);
buf BUF1 (N769, N767);
nand NAND2 (N770, N769, N703);
not NOT1 (N771, N739);
xor XOR2 (N772, N771, N590);
or OR3 (N773, N762, N154, N749);
buf BUF1 (N774, N756);
xor XOR2 (N775, N766, N610);
buf BUF1 (N776, N770);
nand NAND3 (N777, N773, N97, N1);
nor NOR3 (N778, N775, N385, N524);
or OR4 (N779, N768, N413, N112, N209);
or OR3 (N780, N774, N603, N189);
and AND2 (N781, N729, N3);
xor XOR2 (N782, N772, N665);
nor NOR2 (N783, N778, N243);
nand NAND3 (N784, N763, N719, N305);
nand NAND3 (N785, N780, N287, N748);
and AND3 (N786, N785, N766, N739);
nor NOR2 (N787, N783, N591);
or OR4 (N788, N782, N157, N403, N161);
buf BUF1 (N789, N757);
and AND4 (N790, N789, N276, N590, N617);
or OR4 (N791, N787, N699, N46, N464);
nor NOR3 (N792, N790, N701, N543);
and AND3 (N793, N788, N226, N680);
or OR4 (N794, N779, N255, N387, N15);
not NOT1 (N795, N793);
xor XOR2 (N796, N791, N331);
xor XOR2 (N797, N784, N316);
and AND4 (N798, N797, N589, N596, N405);
or OR2 (N799, N777, N636);
xor XOR2 (N800, N796, N50);
not NOT1 (N801, N792);
nand NAND3 (N802, N786, N213, N348);
nand NAND4 (N803, N750, N678, N726, N659);
or OR4 (N804, N794, N260, N313, N229);
xor XOR2 (N805, N802, N141);
buf BUF1 (N806, N799);
xor XOR2 (N807, N781, N473);
buf BUF1 (N808, N803);
nand NAND4 (N809, N801, N542, N458, N176);
and AND3 (N810, N808, N397, N547);
buf BUF1 (N811, N800);
xor XOR2 (N812, N804, N157);
nand NAND4 (N813, N776, N665, N51, N734);
and AND3 (N814, N795, N720, N94);
or OR3 (N815, N807, N581, N183);
xor XOR2 (N816, N810, N112);
not NOT1 (N817, N815);
and AND2 (N818, N811, N224);
nand NAND2 (N819, N816, N217);
or OR4 (N820, N806, N96, N796, N31);
nand NAND3 (N821, N819, N209, N475);
nor NOR3 (N822, N805, N820, N60);
and AND3 (N823, N334, N686, N267);
nor NOR2 (N824, N809, N281);
and AND4 (N825, N824, N145, N726, N366);
buf BUF1 (N826, N798);
nand NAND2 (N827, N823, N491);
or OR3 (N828, N813, N782, N628);
nor NOR2 (N829, N814, N751);
not NOT1 (N830, N821);
and AND3 (N831, N822, N720, N687);
nor NOR4 (N832, N817, N485, N649, N698);
not NOT1 (N833, N818);
xor XOR2 (N834, N826, N746);
xor XOR2 (N835, N831, N31);
buf BUF1 (N836, N825);
not NOT1 (N837, N836);
buf BUF1 (N838, N812);
or OR2 (N839, N838, N387);
buf BUF1 (N840, N839);
xor XOR2 (N841, N840, N282);
buf BUF1 (N842, N833);
and AND3 (N843, N827, N565, N759);
xor XOR2 (N844, N835, N373);
nor NOR3 (N845, N834, N230, N168);
buf BUF1 (N846, N842);
nand NAND4 (N847, N843, N189, N823, N501);
buf BUF1 (N848, N832);
or OR2 (N849, N837, N432);
or OR2 (N850, N846, N60);
not NOT1 (N851, N845);
nor NOR2 (N852, N829, N84);
nand NAND2 (N853, N847, N400);
and AND2 (N854, N841, N559);
buf BUF1 (N855, N848);
buf BUF1 (N856, N851);
nor NOR3 (N857, N852, N119, N484);
not NOT1 (N858, N853);
nor NOR4 (N859, N854, N472, N18, N74);
not NOT1 (N860, N830);
and AND4 (N861, N849, N546, N812, N322);
and AND4 (N862, N844, N625, N736, N287);
or OR3 (N863, N855, N415, N549);
buf BUF1 (N864, N850);
not NOT1 (N865, N860);
not NOT1 (N866, N862);
and AND2 (N867, N864, N496);
xor XOR2 (N868, N863, N474);
nand NAND3 (N869, N865, N18, N548);
not NOT1 (N870, N858);
nor NOR4 (N871, N869, N692, N148, N696);
and AND3 (N872, N857, N596, N695);
xor XOR2 (N873, N868, N865);
not NOT1 (N874, N867);
or OR3 (N875, N861, N184, N71);
and AND4 (N876, N828, N682, N589, N519);
nand NAND2 (N877, N859, N574);
not NOT1 (N878, N876);
xor XOR2 (N879, N872, N828);
xor XOR2 (N880, N877, N457);
not NOT1 (N881, N878);
xor XOR2 (N882, N881, N510);
nor NOR3 (N883, N874, N287, N702);
or OR3 (N884, N879, N610, N883);
nand NAND3 (N885, N702, N873, N486);
or OR2 (N886, N275, N582);
nand NAND3 (N887, N856, N156, N819);
not NOT1 (N888, N875);
nor NOR4 (N889, N871, N30, N43, N209);
nand NAND4 (N890, N888, N17, N838, N163);
or OR4 (N891, N889, N330, N27, N437);
nand NAND4 (N892, N891, N80, N224, N113);
buf BUF1 (N893, N870);
not NOT1 (N894, N886);
buf BUF1 (N895, N894);
nor NOR4 (N896, N884, N602, N364, N851);
not NOT1 (N897, N893);
xor XOR2 (N898, N880, N589);
xor XOR2 (N899, N898, N761);
nand NAND4 (N900, N895, N341, N829, N404);
nor NOR2 (N901, N896, N900);
buf BUF1 (N902, N146);
buf BUF1 (N903, N887);
xor XOR2 (N904, N903, N723);
or OR4 (N905, N902, N11, N172, N396);
or OR2 (N906, N905, N823);
xor XOR2 (N907, N904, N517);
buf BUF1 (N908, N906);
xor XOR2 (N909, N897, N493);
nand NAND2 (N910, N892, N198);
xor XOR2 (N911, N882, N731);
and AND3 (N912, N890, N249, N898);
or OR4 (N913, N912, N55, N428, N764);
buf BUF1 (N914, N866);
nand NAND4 (N915, N885, N260, N4, N228);
and AND4 (N916, N908, N524, N329, N194);
nor NOR4 (N917, N911, N840, N878, N548);
xor XOR2 (N918, N915, N291);
not NOT1 (N919, N918);
not NOT1 (N920, N916);
or OR2 (N921, N914, N797);
or OR2 (N922, N920, N761);
xor XOR2 (N923, N901, N528);
and AND2 (N924, N917, N701);
not NOT1 (N925, N923);
nor NOR4 (N926, N909, N360, N44, N150);
nor NOR2 (N927, N899, N179);
nor NOR2 (N928, N925, N761);
buf BUF1 (N929, N910);
or OR4 (N930, N913, N700, N28, N397);
xor XOR2 (N931, N922, N712);
and AND2 (N932, N928, N582);
xor XOR2 (N933, N932, N301);
buf BUF1 (N934, N930);
or OR2 (N935, N933, N746);
buf BUF1 (N936, N924);
or OR4 (N937, N921, N848, N137, N409);
xor XOR2 (N938, N936, N36);
nor NOR3 (N939, N929, N527, N348);
not NOT1 (N940, N937);
nand NAND2 (N941, N940, N106);
and AND2 (N942, N941, N744);
buf BUF1 (N943, N942);
xor XOR2 (N944, N931, N308);
buf BUF1 (N945, N943);
or OR2 (N946, N919, N280);
not NOT1 (N947, N907);
nand NAND2 (N948, N945, N328);
nor NOR2 (N949, N939, N876);
nand NAND2 (N950, N935, N697);
and AND4 (N951, N926, N572, N661, N637);
xor XOR2 (N952, N944, N372);
and AND4 (N953, N952, N863, N852, N251);
xor XOR2 (N954, N950, N123);
buf BUF1 (N955, N949);
or OR2 (N956, N934, N205);
nor NOR2 (N957, N927, N784);
nand NAND3 (N958, N951, N158, N927);
and AND2 (N959, N955, N86);
xor XOR2 (N960, N938, N924);
not NOT1 (N961, N957);
nor NOR2 (N962, N961, N829);
or OR2 (N963, N956, N353);
buf BUF1 (N964, N946);
and AND4 (N965, N953, N53, N589, N204);
nor NOR2 (N966, N959, N633);
not NOT1 (N967, N958);
or OR3 (N968, N963, N724, N725);
buf BUF1 (N969, N948);
or OR4 (N970, N967, N216, N810, N259);
nand NAND3 (N971, N969, N613, N175);
nand NAND3 (N972, N970, N27, N898);
xor XOR2 (N973, N960, N644);
buf BUF1 (N974, N968);
xor XOR2 (N975, N965, N744);
or OR2 (N976, N962, N690);
not NOT1 (N977, N973);
nand NAND4 (N978, N964, N939, N208, N331);
nand NAND2 (N979, N947, N256);
xor XOR2 (N980, N974, N895);
nor NOR4 (N981, N977, N804, N543, N841);
buf BUF1 (N982, N976);
nor NOR3 (N983, N972, N166, N116);
nor NOR3 (N984, N971, N9, N178);
or OR3 (N985, N978, N119, N637);
or OR3 (N986, N982, N324, N462);
nand NAND4 (N987, N954, N739, N740, N285);
not NOT1 (N988, N979);
and AND3 (N989, N983, N108, N406);
nor NOR3 (N990, N987, N47, N785);
nand NAND2 (N991, N986, N90);
nand NAND2 (N992, N966, N908);
and AND2 (N993, N992, N77);
buf BUF1 (N994, N990);
and AND4 (N995, N991, N605, N409, N234);
or OR2 (N996, N975, N523);
xor XOR2 (N997, N989, N429);
not NOT1 (N998, N985);
and AND2 (N999, N995, N82);
nand NAND3 (N1000, N984, N279, N372);
not NOT1 (N1001, N999);
buf BUF1 (N1002, N1000);
nand NAND3 (N1003, N994, N728, N207);
not NOT1 (N1004, N993);
or OR2 (N1005, N998, N674);
not NOT1 (N1006, N1003);
xor XOR2 (N1007, N1002, N289);
buf BUF1 (N1008, N988);
not NOT1 (N1009, N997);
not NOT1 (N1010, N996);
not NOT1 (N1011, N1010);
and AND3 (N1012, N1005, N992, N857);
xor XOR2 (N1013, N1001, N701);
xor XOR2 (N1014, N980, N281);
and AND3 (N1015, N1012, N388, N615);
not NOT1 (N1016, N1011);
or OR4 (N1017, N1008, N230, N35, N877);
nand NAND3 (N1018, N1007, N897, N944);
or OR4 (N1019, N1016, N1015, N690, N755);
buf BUF1 (N1020, N216);
xor XOR2 (N1021, N1006, N439);
xor XOR2 (N1022, N1014, N679);
xor XOR2 (N1023, N1004, N318);
xor XOR2 (N1024, N1020, N950);
and AND2 (N1025, N1021, N629);
nand NAND2 (N1026, N1025, N809);
nor NOR4 (N1027, N1022, N667, N506, N693);
nor NOR4 (N1028, N1023, N211, N31, N625);
not NOT1 (N1029, N1013);
nand NAND2 (N1030, N1029, N45);
and AND4 (N1031, N1018, N1024, N768, N867);
and AND4 (N1032, N273, N186, N983, N167);
nor NOR2 (N1033, N1028, N744);
and AND4 (N1034, N1033, N271, N514, N983);
buf BUF1 (N1035, N1026);
or OR2 (N1036, N1009, N823);
not NOT1 (N1037, N1034);
and AND2 (N1038, N1037, N518);
not NOT1 (N1039, N1017);
not NOT1 (N1040, N1035);
buf BUF1 (N1041, N1038);
xor XOR2 (N1042, N1036, N900);
not NOT1 (N1043, N1031);
buf BUF1 (N1044, N1039);
xor XOR2 (N1045, N1030, N792);
buf BUF1 (N1046, N981);
nand NAND3 (N1047, N1040, N500, N730);
buf BUF1 (N1048, N1041);
buf BUF1 (N1049, N1032);
buf BUF1 (N1050, N1046);
and AND2 (N1051, N1047, N49);
xor XOR2 (N1052, N1049, N1014);
and AND3 (N1053, N1043, N165, N69);
or OR3 (N1054, N1027, N951, N34);
nand NAND4 (N1055, N1045, N460, N419, N391);
or OR2 (N1056, N1055, N157);
and AND3 (N1057, N1050, N959, N524);
nand NAND4 (N1058, N1054, N604, N252, N609);
xor XOR2 (N1059, N1019, N72);
buf BUF1 (N1060, N1058);
and AND2 (N1061, N1052, N308);
nand NAND3 (N1062, N1057, N531, N816);
not NOT1 (N1063, N1062);
or OR2 (N1064, N1059, N1056);
xor XOR2 (N1065, N433, N826);
and AND3 (N1066, N1048, N535, N1016);
nor NOR2 (N1067, N1061, N626);
or OR4 (N1068, N1042, N622, N476, N14);
nand NAND2 (N1069, N1051, N659);
nor NOR2 (N1070, N1069, N520);
xor XOR2 (N1071, N1060, N344);
or OR2 (N1072, N1070, N275);
buf BUF1 (N1073, N1066);
and AND3 (N1074, N1053, N917, N218);
and AND3 (N1075, N1065, N143, N407);
buf BUF1 (N1076, N1074);
nand NAND2 (N1077, N1044, N948);
buf BUF1 (N1078, N1075);
nand NAND3 (N1079, N1073, N616, N801);
nand NAND2 (N1080, N1068, N3);
or OR2 (N1081, N1080, N60);
xor XOR2 (N1082, N1063, N130);
xor XOR2 (N1083, N1072, N488);
not NOT1 (N1084, N1071);
or OR3 (N1085, N1082, N763, N13);
buf BUF1 (N1086, N1076);
buf BUF1 (N1087, N1079);
and AND3 (N1088, N1085, N619, N187);
nand NAND4 (N1089, N1078, N620, N19, N3);
and AND3 (N1090, N1089, N833, N352);
nand NAND3 (N1091, N1067, N965, N678);
or OR2 (N1092, N1064, N60);
not NOT1 (N1093, N1084);
or OR3 (N1094, N1081, N871, N760);
or OR2 (N1095, N1092, N217);
not NOT1 (N1096, N1095);
buf BUF1 (N1097, N1083);
buf BUF1 (N1098, N1090);
buf BUF1 (N1099, N1088);
or OR2 (N1100, N1091, N458);
nand NAND4 (N1101, N1086, N463, N1037, N264);
and AND2 (N1102, N1093, N675);
nand NAND2 (N1103, N1077, N971);
and AND4 (N1104, N1100, N1040, N217, N315);
nand NAND2 (N1105, N1101, N516);
buf BUF1 (N1106, N1087);
not NOT1 (N1107, N1102);
nand NAND4 (N1108, N1105, N1103, N688, N930);
or OR2 (N1109, N968, N251);
and AND4 (N1110, N1106, N338, N1101, N966);
and AND4 (N1111, N1097, N26, N752, N280);
buf BUF1 (N1112, N1107);
or OR4 (N1113, N1111, N529, N497, N178);
buf BUF1 (N1114, N1099);
and AND4 (N1115, N1113, N390, N760, N647);
nor NOR3 (N1116, N1094, N969, N55);
buf BUF1 (N1117, N1104);
and AND2 (N1118, N1098, N145);
not NOT1 (N1119, N1116);
or OR4 (N1120, N1118, N243, N266, N963);
nand NAND4 (N1121, N1117, N786, N921, N759);
buf BUF1 (N1122, N1096);
or OR4 (N1123, N1110, N1053, N318, N733);
xor XOR2 (N1124, N1121, N975);
and AND4 (N1125, N1123, N174, N224, N732);
xor XOR2 (N1126, N1125, N353);
xor XOR2 (N1127, N1115, N631);
not NOT1 (N1128, N1124);
not NOT1 (N1129, N1114);
or OR3 (N1130, N1126, N655, N114);
nand NAND4 (N1131, N1119, N545, N474, N811);
and AND4 (N1132, N1122, N1121, N605, N1104);
buf BUF1 (N1133, N1130);
nand NAND4 (N1134, N1108, N492, N479, N996);
or OR4 (N1135, N1128, N21, N775, N203);
buf BUF1 (N1136, N1129);
or OR3 (N1137, N1109, N411, N480);
xor XOR2 (N1138, N1112, N834);
nor NOR3 (N1139, N1136, N752, N43);
nor NOR2 (N1140, N1139, N875);
nand NAND3 (N1141, N1131, N681, N1026);
nor NOR3 (N1142, N1133, N177, N403);
xor XOR2 (N1143, N1142, N205);
xor XOR2 (N1144, N1134, N940);
buf BUF1 (N1145, N1144);
nor NOR3 (N1146, N1138, N506, N1049);
xor XOR2 (N1147, N1140, N165);
nor NOR2 (N1148, N1135, N662);
buf BUF1 (N1149, N1145);
nand NAND2 (N1150, N1137, N216);
not NOT1 (N1151, N1132);
or OR4 (N1152, N1120, N1079, N288, N895);
nand NAND4 (N1153, N1150, N80, N879, N514);
nor NOR3 (N1154, N1127, N99, N46);
nor NOR3 (N1155, N1152, N1012, N1007);
nand NAND2 (N1156, N1153, N142);
and AND2 (N1157, N1149, N968);
or OR4 (N1158, N1157, N1059, N1044, N550);
xor XOR2 (N1159, N1141, N263);
and AND4 (N1160, N1159, N441, N354, N1142);
nor NOR4 (N1161, N1154, N185, N979, N895);
xor XOR2 (N1162, N1143, N1133);
nand NAND2 (N1163, N1148, N670);
buf BUF1 (N1164, N1162);
nor NOR2 (N1165, N1146, N695);
xor XOR2 (N1166, N1165, N286);
xor XOR2 (N1167, N1163, N393);
xor XOR2 (N1168, N1158, N369);
nor NOR2 (N1169, N1166, N807);
nand NAND4 (N1170, N1151, N426, N1034, N1042);
or OR3 (N1171, N1147, N56, N425);
xor XOR2 (N1172, N1164, N122);
and AND3 (N1173, N1172, N843, N888);
nor NOR4 (N1174, N1156, N764, N881, N922);
xor XOR2 (N1175, N1168, N358);
nor NOR3 (N1176, N1174, N876, N136);
or OR4 (N1177, N1161, N962, N613, N88);
nand NAND4 (N1178, N1169, N229, N1024, N83);
nor NOR3 (N1179, N1155, N652, N1088);
not NOT1 (N1180, N1173);
or OR3 (N1181, N1177, N1158, N286);
nand NAND4 (N1182, N1175, N440, N99, N2);
nor NOR2 (N1183, N1160, N757);
xor XOR2 (N1184, N1170, N878);
nand NAND3 (N1185, N1182, N150, N494);
buf BUF1 (N1186, N1167);
nand NAND4 (N1187, N1183, N72, N587, N1185);
not NOT1 (N1188, N203);
not NOT1 (N1189, N1186);
and AND2 (N1190, N1179, N1122);
nand NAND4 (N1191, N1184, N676, N477, N381);
buf BUF1 (N1192, N1176);
and AND2 (N1193, N1189, N1029);
nor NOR4 (N1194, N1188, N367, N383, N192);
or OR3 (N1195, N1193, N787, N481);
buf BUF1 (N1196, N1195);
nand NAND3 (N1197, N1178, N682, N354);
or OR3 (N1198, N1197, N564, N67);
not NOT1 (N1199, N1180);
not NOT1 (N1200, N1199);
buf BUF1 (N1201, N1200);
xor XOR2 (N1202, N1191, N664);
nor NOR2 (N1203, N1190, N1178);
not NOT1 (N1204, N1171);
buf BUF1 (N1205, N1201);
nor NOR2 (N1206, N1196, N764);
not NOT1 (N1207, N1192);
nor NOR4 (N1208, N1198, N689, N275, N851);
or OR2 (N1209, N1207, N36);
and AND4 (N1210, N1205, N707, N954, N291);
not NOT1 (N1211, N1204);
xor XOR2 (N1212, N1206, N16);
or OR4 (N1213, N1211, N707, N409, N14);
nand NAND2 (N1214, N1187, N195);
buf BUF1 (N1215, N1181);
buf BUF1 (N1216, N1194);
and AND2 (N1217, N1210, N237);
not NOT1 (N1218, N1209);
not NOT1 (N1219, N1208);
not NOT1 (N1220, N1212);
or OR4 (N1221, N1202, N1161, N1009, N549);
not NOT1 (N1222, N1216);
buf BUF1 (N1223, N1217);
nand NAND4 (N1224, N1203, N639, N13, N262);
and AND2 (N1225, N1219, N279);
nor NOR4 (N1226, N1223, N85, N929, N683);
or OR3 (N1227, N1226, N719, N607);
or OR2 (N1228, N1227, N388);
not NOT1 (N1229, N1218);
and AND3 (N1230, N1229, N812, N515);
or OR3 (N1231, N1214, N775, N760);
nand NAND4 (N1232, N1215, N286, N431, N177);
nand NAND4 (N1233, N1232, N885, N644, N246);
buf BUF1 (N1234, N1230);
or OR3 (N1235, N1224, N366, N714);
nand NAND3 (N1236, N1222, N3, N310);
and AND4 (N1237, N1234, N496, N992, N752);
nand NAND2 (N1238, N1221, N735);
xor XOR2 (N1239, N1220, N216);
xor XOR2 (N1240, N1225, N435);
or OR4 (N1241, N1238, N812, N754, N51);
buf BUF1 (N1242, N1241);
xor XOR2 (N1243, N1213, N684);
buf BUF1 (N1244, N1231);
or OR4 (N1245, N1240, N291, N513, N635);
nand NAND4 (N1246, N1228, N176, N521, N1206);
buf BUF1 (N1247, N1236);
buf BUF1 (N1248, N1235);
nand NAND2 (N1249, N1245, N738);
xor XOR2 (N1250, N1248, N1164);
buf BUF1 (N1251, N1242);
nor NOR4 (N1252, N1251, N620, N392, N520);
and AND2 (N1253, N1250, N1123);
or OR4 (N1254, N1252, N1180, N427, N275);
nor NOR2 (N1255, N1237, N307);
or OR4 (N1256, N1249, N1051, N1203, N17);
and AND3 (N1257, N1233, N247, N143);
nor NOR2 (N1258, N1246, N1038);
nor NOR2 (N1259, N1253, N530);
not NOT1 (N1260, N1256);
nand NAND2 (N1261, N1254, N40);
not NOT1 (N1262, N1247);
nand NAND3 (N1263, N1255, N558, N411);
nor NOR3 (N1264, N1239, N241, N1040);
buf BUF1 (N1265, N1259);
and AND3 (N1266, N1262, N1005, N945);
nor NOR2 (N1267, N1243, N1012);
or OR2 (N1268, N1258, N663);
nor NOR2 (N1269, N1261, N164);
nand NAND4 (N1270, N1268, N1223, N35, N1162);
or OR2 (N1271, N1263, N490);
and AND2 (N1272, N1264, N833);
xor XOR2 (N1273, N1269, N449);
nand NAND2 (N1274, N1257, N669);
buf BUF1 (N1275, N1265);
or OR3 (N1276, N1260, N668, N111);
not NOT1 (N1277, N1273);
or OR4 (N1278, N1276, N692, N733, N21);
and AND2 (N1279, N1267, N1164);
buf BUF1 (N1280, N1272);
and AND4 (N1281, N1244, N465, N79, N126);
nand NAND4 (N1282, N1271, N963, N118, N1125);
not NOT1 (N1283, N1279);
xor XOR2 (N1284, N1274, N376);
nand NAND2 (N1285, N1282, N472);
and AND3 (N1286, N1277, N751, N78);
or OR3 (N1287, N1281, N642, N765);
nor NOR3 (N1288, N1286, N1186, N1163);
nand NAND2 (N1289, N1283, N1275);
xor XOR2 (N1290, N1164, N1144);
nand NAND4 (N1291, N1290, N916, N81, N965);
and AND4 (N1292, N1284, N754, N82, N156);
xor XOR2 (N1293, N1280, N1240);
nor NOR3 (N1294, N1293, N1133, N588);
nor NOR4 (N1295, N1287, N495, N13, N474);
or OR3 (N1296, N1292, N634, N523);
nand NAND2 (N1297, N1296, N290);
not NOT1 (N1298, N1291);
nand NAND2 (N1299, N1278, N623);
nor NOR2 (N1300, N1298, N1103);
or OR2 (N1301, N1288, N288);
and AND3 (N1302, N1300, N609, N264);
xor XOR2 (N1303, N1297, N1200);
not NOT1 (N1304, N1301);
nand NAND3 (N1305, N1294, N922, N570);
xor XOR2 (N1306, N1305, N265);
buf BUF1 (N1307, N1289);
nand NAND3 (N1308, N1266, N1186, N118);
nor NOR4 (N1309, N1270, N79, N641, N1285);
nor NOR2 (N1310, N990, N1234);
xor XOR2 (N1311, N1299, N800);
or OR3 (N1312, N1309, N321, N430);
and AND3 (N1313, N1306, N240, N721);
not NOT1 (N1314, N1310);
nand NAND4 (N1315, N1302, N756, N985, N1221);
buf BUF1 (N1316, N1304);
buf BUF1 (N1317, N1314);
xor XOR2 (N1318, N1316, N642);
xor XOR2 (N1319, N1315, N182);
and AND2 (N1320, N1319, N1066);
and AND3 (N1321, N1307, N520, N241);
or OR3 (N1322, N1311, N559, N738);
nand NAND4 (N1323, N1312, N1143, N256, N95);
buf BUF1 (N1324, N1321);
or OR3 (N1325, N1313, N807, N372);
or OR4 (N1326, N1317, N1309, N633, N1206);
xor XOR2 (N1327, N1318, N142);
buf BUF1 (N1328, N1327);
or OR3 (N1329, N1324, N801, N1108);
or OR3 (N1330, N1322, N616, N1027);
nor NOR4 (N1331, N1303, N186, N437, N539);
or OR2 (N1332, N1328, N23);
nand NAND2 (N1333, N1326, N1308);
xor XOR2 (N1334, N310, N1267);
nand NAND4 (N1335, N1331, N736, N414, N386);
nor NOR4 (N1336, N1295, N1017, N964, N82);
nor NOR2 (N1337, N1332, N286);
nand NAND2 (N1338, N1335, N905);
not NOT1 (N1339, N1323);
xor XOR2 (N1340, N1334, N433);
and AND2 (N1341, N1337, N769);
buf BUF1 (N1342, N1339);
nor NOR2 (N1343, N1325, N1120);
buf BUF1 (N1344, N1342);
nor NOR2 (N1345, N1336, N1343);
buf BUF1 (N1346, N1099);
not NOT1 (N1347, N1346);
nand NAND3 (N1348, N1330, N1085, N676);
nand NAND4 (N1349, N1340, N1338, N791, N874);
not NOT1 (N1350, N1266);
or OR3 (N1351, N1333, N483, N877);
nor NOR4 (N1352, N1320, N654, N15, N990);
buf BUF1 (N1353, N1344);
or OR3 (N1354, N1347, N1107, N580);
nor NOR4 (N1355, N1349, N1108, N415, N485);
buf BUF1 (N1356, N1350);
or OR4 (N1357, N1352, N261, N1194, N1314);
nand NAND2 (N1358, N1354, N1083);
not NOT1 (N1359, N1329);
buf BUF1 (N1360, N1358);
nand NAND4 (N1361, N1360, N1268, N318, N655);
buf BUF1 (N1362, N1357);
xor XOR2 (N1363, N1345, N230);
xor XOR2 (N1364, N1353, N273);
or OR4 (N1365, N1363, N613, N736, N1059);
or OR3 (N1366, N1365, N300, N1024);
or OR4 (N1367, N1355, N12, N593, N479);
xor XOR2 (N1368, N1356, N208);
or OR4 (N1369, N1367, N867, N107, N831);
nor NOR3 (N1370, N1341, N534, N286);
nor NOR4 (N1371, N1366, N438, N609, N1163);
xor XOR2 (N1372, N1361, N1104);
nor NOR3 (N1373, N1370, N967, N957);
or OR3 (N1374, N1351, N973, N775);
buf BUF1 (N1375, N1348);
and AND3 (N1376, N1374, N499, N649);
nand NAND2 (N1377, N1375, N1290);
xor XOR2 (N1378, N1371, N1204);
or OR4 (N1379, N1362, N338, N626, N949);
not NOT1 (N1380, N1378);
xor XOR2 (N1381, N1379, N4);
xor XOR2 (N1382, N1380, N713);
or OR3 (N1383, N1372, N1109, N550);
not NOT1 (N1384, N1383);
xor XOR2 (N1385, N1376, N70);
nand NAND4 (N1386, N1369, N239, N1081, N472);
nor NOR2 (N1387, N1364, N66);
nand NAND4 (N1388, N1359, N1246, N221, N432);
and AND3 (N1389, N1388, N644, N139);
buf BUF1 (N1390, N1368);
or OR4 (N1391, N1387, N365, N54, N849);
and AND3 (N1392, N1386, N694, N580);
nand NAND4 (N1393, N1381, N1183, N307, N140);
not NOT1 (N1394, N1373);
nand NAND4 (N1395, N1377, N534, N713, N789);
or OR4 (N1396, N1384, N480, N1379, N312);
or OR4 (N1397, N1389, N1009, N793, N154);
nand NAND2 (N1398, N1393, N935);
not NOT1 (N1399, N1396);
not NOT1 (N1400, N1382);
nor NOR2 (N1401, N1397, N372);
or OR4 (N1402, N1385, N826, N1246, N570);
and AND3 (N1403, N1391, N564, N821);
buf BUF1 (N1404, N1394);
xor XOR2 (N1405, N1400, N537);
not NOT1 (N1406, N1392);
not NOT1 (N1407, N1402);
or OR4 (N1408, N1403, N943, N911, N670);
not NOT1 (N1409, N1395);
and AND4 (N1410, N1408, N1317, N1071, N296);
and AND4 (N1411, N1407, N1160, N276, N765);
buf BUF1 (N1412, N1399);
not NOT1 (N1413, N1410);
not NOT1 (N1414, N1406);
buf BUF1 (N1415, N1405);
not NOT1 (N1416, N1412);
nand NAND3 (N1417, N1416, N699, N55);
and AND2 (N1418, N1390, N895);
xor XOR2 (N1419, N1415, N126);
and AND2 (N1420, N1409, N687);
buf BUF1 (N1421, N1420);
nor NOR2 (N1422, N1421, N334);
nand NAND3 (N1423, N1413, N1346, N924);
xor XOR2 (N1424, N1414, N382);
not NOT1 (N1425, N1404);
xor XOR2 (N1426, N1422, N1266);
buf BUF1 (N1427, N1425);
or OR2 (N1428, N1418, N1110);
nand NAND2 (N1429, N1426, N852);
nand NAND4 (N1430, N1429, N129, N1359, N569);
not NOT1 (N1431, N1398);
nor NOR3 (N1432, N1428, N1193, N120);
nand NAND2 (N1433, N1423, N612);
not NOT1 (N1434, N1419);
nand NAND2 (N1435, N1401, N155);
and AND4 (N1436, N1433, N86, N645, N474);
buf BUF1 (N1437, N1432);
not NOT1 (N1438, N1437);
and AND3 (N1439, N1434, N850, N1067);
xor XOR2 (N1440, N1427, N471);
buf BUF1 (N1441, N1431);
xor XOR2 (N1442, N1436, N1188);
nand NAND4 (N1443, N1417, N724, N441, N954);
nor NOR3 (N1444, N1441, N776, N210);
and AND3 (N1445, N1439, N1041, N745);
buf BUF1 (N1446, N1435);
or OR2 (N1447, N1438, N441);
nor NOR4 (N1448, N1444, N1034, N888, N1362);
nor NOR3 (N1449, N1445, N834, N5);
or OR3 (N1450, N1448, N1223, N301);
or OR4 (N1451, N1446, N126, N802, N772);
not NOT1 (N1452, N1451);
not NOT1 (N1453, N1411);
and AND4 (N1454, N1450, N874, N820, N1264);
or OR4 (N1455, N1443, N1395, N46, N367);
nor NOR2 (N1456, N1453, N955);
not NOT1 (N1457, N1456);
and AND3 (N1458, N1457, N467, N841);
nor NOR2 (N1459, N1442, N417);
nor NOR4 (N1460, N1458, N116, N1079, N500);
not NOT1 (N1461, N1430);
buf BUF1 (N1462, N1449);
xor XOR2 (N1463, N1454, N865);
nor NOR3 (N1464, N1452, N168, N505);
and AND2 (N1465, N1455, N1043);
nand NAND4 (N1466, N1459, N1054, N1340, N587);
or OR2 (N1467, N1462, N415);
not NOT1 (N1468, N1447);
xor XOR2 (N1469, N1464, N247);
xor XOR2 (N1470, N1460, N1404);
xor XOR2 (N1471, N1465, N833);
nand NAND4 (N1472, N1461, N479, N206, N602);
nand NAND2 (N1473, N1466, N707);
not NOT1 (N1474, N1440);
nand NAND3 (N1475, N1473, N1314, N479);
nand NAND2 (N1476, N1463, N371);
nand NAND2 (N1477, N1467, N796);
xor XOR2 (N1478, N1469, N829);
nand NAND4 (N1479, N1474, N808, N1349, N1232);
nand NAND2 (N1480, N1424, N580);
not NOT1 (N1481, N1479);
or OR4 (N1482, N1470, N733, N222, N1089);
or OR2 (N1483, N1477, N217);
or OR4 (N1484, N1471, N353, N164, N141);
or OR4 (N1485, N1475, N157, N602, N42);
and AND3 (N1486, N1484, N180, N820);
xor XOR2 (N1487, N1468, N1100);
xor XOR2 (N1488, N1486, N749);
xor XOR2 (N1489, N1481, N1404);
not NOT1 (N1490, N1482);
and AND4 (N1491, N1472, N601, N373, N336);
or OR3 (N1492, N1488, N1087, N141);
nand NAND2 (N1493, N1476, N220);
buf BUF1 (N1494, N1493);
and AND3 (N1495, N1478, N787, N256);
xor XOR2 (N1496, N1487, N1210);
buf BUF1 (N1497, N1491);
buf BUF1 (N1498, N1480);
buf BUF1 (N1499, N1490);
or OR2 (N1500, N1485, N702);
nor NOR4 (N1501, N1499, N77, N1451, N50);
buf BUF1 (N1502, N1498);
xor XOR2 (N1503, N1501, N1220);
or OR4 (N1504, N1496, N295, N469, N132);
nor NOR4 (N1505, N1495, N334, N1485, N992);
buf BUF1 (N1506, N1492);
xor XOR2 (N1507, N1494, N1240);
nand NAND4 (N1508, N1505, N72, N343, N498);
xor XOR2 (N1509, N1489, N794);
nor NOR4 (N1510, N1508, N1190, N1035, N1145);
xor XOR2 (N1511, N1502, N44);
and AND2 (N1512, N1504, N818);
nor NOR4 (N1513, N1509, N796, N1003, N578);
and AND2 (N1514, N1512, N1094);
not NOT1 (N1515, N1507);
or OR2 (N1516, N1511, N617);
or OR2 (N1517, N1514, N408);
not NOT1 (N1518, N1515);
nor NOR4 (N1519, N1518, N1099, N152, N1422);
not NOT1 (N1520, N1503);
or OR2 (N1521, N1510, N245);
nor NOR4 (N1522, N1483, N14, N1105, N1274);
or OR4 (N1523, N1522, N131, N1437, N830);
or OR2 (N1524, N1519, N1317);
xor XOR2 (N1525, N1506, N681);
or OR4 (N1526, N1520, N449, N820, N496);
nand NAND4 (N1527, N1521, N998, N823, N1341);
nor NOR3 (N1528, N1527, N597, N96);
or OR4 (N1529, N1524, N29, N1287, N666);
buf BUF1 (N1530, N1497);
and AND2 (N1531, N1523, N909);
and AND3 (N1532, N1500, N650, N1171);
not NOT1 (N1533, N1516);
nor NOR2 (N1534, N1533, N919);
xor XOR2 (N1535, N1513, N1103);
buf BUF1 (N1536, N1529);
buf BUF1 (N1537, N1526);
or OR4 (N1538, N1528, N230, N782, N487);
nand NAND4 (N1539, N1534, N63, N580, N421);
nor NOR2 (N1540, N1539, N149);
or OR4 (N1541, N1540, N1486, N1366, N998);
nor NOR3 (N1542, N1532, N981, N346);
and AND3 (N1543, N1541, N833, N521);
xor XOR2 (N1544, N1525, N725);
buf BUF1 (N1545, N1530);
or OR4 (N1546, N1545, N789, N461, N725);
xor XOR2 (N1547, N1538, N655);
nand NAND2 (N1548, N1531, N1403);
buf BUF1 (N1549, N1548);
buf BUF1 (N1550, N1537);
or OR3 (N1551, N1542, N36, N1007);
or OR4 (N1552, N1546, N864, N36, N1504);
buf BUF1 (N1553, N1536);
or OR2 (N1554, N1543, N160);
or OR4 (N1555, N1552, N98, N1295, N281);
buf BUF1 (N1556, N1547);
or OR4 (N1557, N1553, N1418, N1290, N793);
nand NAND3 (N1558, N1550, N1543, N1178);
buf BUF1 (N1559, N1554);
nand NAND3 (N1560, N1558, N1119, N1231);
nor NOR3 (N1561, N1544, N501, N1098);
xor XOR2 (N1562, N1559, N235);
nor NOR2 (N1563, N1561, N27);
not NOT1 (N1564, N1560);
buf BUF1 (N1565, N1549);
or OR2 (N1566, N1535, N580);
or OR2 (N1567, N1565, N1174);
nand NAND3 (N1568, N1555, N509, N766);
xor XOR2 (N1569, N1556, N1374);
and AND4 (N1570, N1562, N920, N1438, N1129);
or OR3 (N1571, N1567, N233, N671);
not NOT1 (N1572, N1571);
not NOT1 (N1573, N1566);
nor NOR2 (N1574, N1568, N80);
nand NAND3 (N1575, N1573, N1049, N531);
xor XOR2 (N1576, N1563, N868);
nand NAND3 (N1577, N1570, N353, N1235);
buf BUF1 (N1578, N1574);
buf BUF1 (N1579, N1557);
and AND2 (N1580, N1578, N1072);
nand NAND2 (N1581, N1572, N469);
nor NOR4 (N1582, N1581, N1251, N1052, N643);
nor NOR4 (N1583, N1517, N1438, N921, N1280);
nor NOR3 (N1584, N1569, N1384, N1236);
xor XOR2 (N1585, N1584, N171);
buf BUF1 (N1586, N1551);
buf BUF1 (N1587, N1575);
xor XOR2 (N1588, N1580, N1229);
nand NAND3 (N1589, N1564, N608, N338);
or OR3 (N1590, N1586, N1333, N1278);
buf BUF1 (N1591, N1576);
nor NOR3 (N1592, N1589, N1179, N964);
nor NOR3 (N1593, N1577, N993, N1050);
nor NOR4 (N1594, N1582, N879, N795, N792);
and AND2 (N1595, N1583, N431);
and AND2 (N1596, N1592, N1187);
buf BUF1 (N1597, N1596);
nand NAND3 (N1598, N1594, N628, N577);
and AND2 (N1599, N1597, N169);
xor XOR2 (N1600, N1598, N781);
nor NOR4 (N1601, N1588, N1169, N1405, N723);
buf BUF1 (N1602, N1595);
or OR4 (N1603, N1602, N105, N1529, N427);
xor XOR2 (N1604, N1579, N191);
nand NAND4 (N1605, N1590, N233, N59, N986);
not NOT1 (N1606, N1587);
and AND4 (N1607, N1605, N1026, N709, N1103);
buf BUF1 (N1608, N1607);
buf BUF1 (N1609, N1591);
or OR2 (N1610, N1599, N139);
nor NOR3 (N1611, N1603, N383, N1403);
nor NOR2 (N1612, N1606, N679);
or OR4 (N1613, N1612, N1510, N517, N776);
nand NAND2 (N1614, N1611, N131);
or OR3 (N1615, N1610, N856, N627);
buf BUF1 (N1616, N1585);
nand NAND3 (N1617, N1600, N336, N1439);
buf BUF1 (N1618, N1616);
or OR2 (N1619, N1601, N667);
buf BUF1 (N1620, N1613);
nor NOR4 (N1621, N1604, N1046, N813, N981);
or OR2 (N1622, N1608, N930);
nand NAND2 (N1623, N1617, N808);
or OR2 (N1624, N1618, N594);
xor XOR2 (N1625, N1614, N1068);
and AND3 (N1626, N1623, N1067, N1544);
not NOT1 (N1627, N1626);
not NOT1 (N1628, N1593);
xor XOR2 (N1629, N1615, N353);
and AND2 (N1630, N1619, N90);
nand NAND4 (N1631, N1629, N107, N1257, N1061);
and AND4 (N1632, N1630, N182, N1343, N876);
xor XOR2 (N1633, N1627, N831);
and AND4 (N1634, N1625, N1624, N1499, N1220);
buf BUF1 (N1635, N1192);
or OR3 (N1636, N1633, N1330, N740);
buf BUF1 (N1637, N1622);
buf BUF1 (N1638, N1631);
nand NAND3 (N1639, N1638, N70, N1241);
or OR2 (N1640, N1628, N771);
buf BUF1 (N1641, N1640);
buf BUF1 (N1642, N1632);
nor NOR3 (N1643, N1642, N358, N801);
nand NAND3 (N1644, N1637, N704, N1161);
not NOT1 (N1645, N1644);
nor NOR2 (N1646, N1639, N742);
and AND2 (N1647, N1635, N868);
not NOT1 (N1648, N1643);
not NOT1 (N1649, N1634);
and AND3 (N1650, N1649, N102, N146);
not NOT1 (N1651, N1621);
xor XOR2 (N1652, N1609, N536);
or OR2 (N1653, N1645, N1595);
nor NOR2 (N1654, N1650, N897);
buf BUF1 (N1655, N1641);
nand NAND3 (N1656, N1647, N1024, N187);
buf BUF1 (N1657, N1653);
nand NAND2 (N1658, N1648, N1054);
xor XOR2 (N1659, N1656, N264);
not NOT1 (N1660, N1659);
nand NAND4 (N1661, N1651, N491, N1025, N779);
nand NAND4 (N1662, N1646, N1020, N487, N267);
nand NAND3 (N1663, N1661, N1302, N636);
xor XOR2 (N1664, N1658, N1033);
not NOT1 (N1665, N1655);
or OR2 (N1666, N1657, N1404);
and AND3 (N1667, N1662, N261, N509);
or OR4 (N1668, N1666, N740, N937, N80);
or OR2 (N1669, N1652, N284);
not NOT1 (N1670, N1636);
or OR3 (N1671, N1660, N164, N20);
and AND3 (N1672, N1664, N861, N1167);
nand NAND4 (N1673, N1620, N1365, N1452, N23);
not NOT1 (N1674, N1665);
nor NOR3 (N1675, N1673, N1595, N1650);
or OR4 (N1676, N1674, N971, N1444, N1571);
xor XOR2 (N1677, N1668, N68);
not NOT1 (N1678, N1670);
and AND4 (N1679, N1676, N1651, N1545, N1275);
xor XOR2 (N1680, N1679, N1645);
nor NOR3 (N1681, N1671, N1102, N1580);
or OR2 (N1682, N1680, N1476);
buf BUF1 (N1683, N1654);
nand NAND3 (N1684, N1683, N292, N986);
nand NAND3 (N1685, N1677, N1410, N941);
or OR2 (N1686, N1681, N610);
not NOT1 (N1687, N1682);
nand NAND4 (N1688, N1675, N1446, N1315, N485);
nor NOR3 (N1689, N1663, N1473, N1036);
and AND3 (N1690, N1688, N781, N1314);
nor NOR2 (N1691, N1669, N505);
buf BUF1 (N1692, N1686);
nor NOR4 (N1693, N1687, N778, N1471, N1078);
not NOT1 (N1694, N1691);
buf BUF1 (N1695, N1667);
nor NOR4 (N1696, N1695, N1460, N460, N1409);
xor XOR2 (N1697, N1678, N1472);
and AND2 (N1698, N1692, N1585);
not NOT1 (N1699, N1696);
nand NAND2 (N1700, N1672, N445);
and AND3 (N1701, N1685, N876, N577);
not NOT1 (N1702, N1700);
xor XOR2 (N1703, N1699, N1581);
not NOT1 (N1704, N1698);
nor NOR2 (N1705, N1704, N443);
nand NAND4 (N1706, N1684, N514, N811, N24);
xor XOR2 (N1707, N1694, N201);
not NOT1 (N1708, N1701);
or OR4 (N1709, N1693, N44, N418, N764);
and AND3 (N1710, N1709, N941, N756);
or OR2 (N1711, N1703, N1132);
or OR3 (N1712, N1705, N348, N931);
nand NAND2 (N1713, N1712, N1261);
nand NAND3 (N1714, N1690, N1263, N303);
xor XOR2 (N1715, N1711, N65);
nand NAND4 (N1716, N1710, N656, N84, N836);
xor XOR2 (N1717, N1715, N1025);
and AND3 (N1718, N1707, N1476, N1620);
not NOT1 (N1719, N1689);
buf BUF1 (N1720, N1717);
nor NOR2 (N1721, N1706, N916);
buf BUF1 (N1722, N1708);
nor NOR3 (N1723, N1721, N507, N1456);
buf BUF1 (N1724, N1722);
xor XOR2 (N1725, N1719, N1446);
not NOT1 (N1726, N1724);
nand NAND3 (N1727, N1713, N1666, N752);
not NOT1 (N1728, N1697);
nor NOR2 (N1729, N1728, N650);
nor NOR2 (N1730, N1716, N1338);
and AND4 (N1731, N1720, N1453, N509, N526);
nor NOR2 (N1732, N1718, N407);
not NOT1 (N1733, N1726);
nand NAND2 (N1734, N1729, N382);
not NOT1 (N1735, N1727);
nor NOR3 (N1736, N1735, N664, N84);
not NOT1 (N1737, N1714);
nand NAND3 (N1738, N1736, N391, N539);
and AND4 (N1739, N1723, N1728, N136, N1187);
and AND2 (N1740, N1725, N1093);
nor NOR4 (N1741, N1732, N829, N39, N1563);
not NOT1 (N1742, N1733);
nand NAND4 (N1743, N1741, N648, N384, N971);
xor XOR2 (N1744, N1742, N1290);
nand NAND4 (N1745, N1738, N1517, N100, N539);
xor XOR2 (N1746, N1702, N308);
not NOT1 (N1747, N1739);
not NOT1 (N1748, N1734);
nor NOR3 (N1749, N1744, N644, N99);
nand NAND4 (N1750, N1731, N393, N737, N17);
nor NOR4 (N1751, N1750, N677, N1030, N248);
xor XOR2 (N1752, N1740, N996);
nor NOR3 (N1753, N1737, N79, N724);
and AND2 (N1754, N1753, N316);
buf BUF1 (N1755, N1751);
and AND2 (N1756, N1755, N595);
and AND2 (N1757, N1749, N1557);
or OR3 (N1758, N1756, N118, N1652);
and AND3 (N1759, N1748, N1014, N405);
or OR3 (N1760, N1758, N825, N1294);
nand NAND2 (N1761, N1752, N473);
nor NOR3 (N1762, N1760, N1646, N272);
nand NAND4 (N1763, N1762, N1114, N206, N1696);
buf BUF1 (N1764, N1757);
or OR3 (N1765, N1764, N1336, N332);
or OR3 (N1766, N1747, N840, N1440);
or OR3 (N1767, N1745, N1735, N757);
and AND3 (N1768, N1730, N11, N1620);
xor XOR2 (N1769, N1759, N1578);
buf BUF1 (N1770, N1763);
xor XOR2 (N1771, N1770, N1660);
buf BUF1 (N1772, N1768);
buf BUF1 (N1773, N1766);
buf BUF1 (N1774, N1772);
and AND3 (N1775, N1767, N939, N531);
or OR4 (N1776, N1774, N710, N1661, N50);
or OR3 (N1777, N1771, N870, N1121);
not NOT1 (N1778, N1775);
not NOT1 (N1779, N1773);
buf BUF1 (N1780, N1765);
xor XOR2 (N1781, N1778, N498);
and AND2 (N1782, N1781, N1101);
not NOT1 (N1783, N1743);
nand NAND4 (N1784, N1761, N731, N1085, N1574);
buf BUF1 (N1785, N1784);
nor NOR2 (N1786, N1776, N1435);
xor XOR2 (N1787, N1782, N186);
xor XOR2 (N1788, N1777, N261);
xor XOR2 (N1789, N1785, N864);
xor XOR2 (N1790, N1787, N567);
not NOT1 (N1791, N1769);
or OR3 (N1792, N1791, N1698, N175);
buf BUF1 (N1793, N1783);
not NOT1 (N1794, N1789);
or OR4 (N1795, N1794, N991, N1513, N1354);
not NOT1 (N1796, N1792);
or OR4 (N1797, N1779, N1184, N407, N492);
nand NAND2 (N1798, N1746, N1118);
and AND4 (N1799, N1790, N1617, N1502, N1087);
and AND3 (N1800, N1799, N104, N1406);
not NOT1 (N1801, N1796);
and AND3 (N1802, N1800, N1044, N1575);
not NOT1 (N1803, N1801);
not NOT1 (N1804, N1780);
buf BUF1 (N1805, N1803);
buf BUF1 (N1806, N1804);
or OR3 (N1807, N1754, N42, N234);
nor NOR3 (N1808, N1793, N969, N452);
or OR4 (N1809, N1806, N1385, N1128, N720);
or OR2 (N1810, N1802, N235);
or OR3 (N1811, N1788, N899, N780);
or OR3 (N1812, N1810, N862, N502);
xor XOR2 (N1813, N1812, N256);
not NOT1 (N1814, N1808);
not NOT1 (N1815, N1814);
nand NAND2 (N1816, N1797, N1479);
xor XOR2 (N1817, N1815, N429);
buf BUF1 (N1818, N1807);
not NOT1 (N1819, N1805);
nand NAND4 (N1820, N1809, N441, N483, N20);
buf BUF1 (N1821, N1819);
nand NAND3 (N1822, N1813, N1130, N1686);
nand NAND2 (N1823, N1786, N1168);
nand NAND4 (N1824, N1822, N1753, N782, N318);
buf BUF1 (N1825, N1820);
buf BUF1 (N1826, N1816);
and AND3 (N1827, N1817, N1036, N904);
and AND4 (N1828, N1818, N661, N1073, N824);
nor NOR3 (N1829, N1811, N956, N1794);
nand NAND4 (N1830, N1825, N1603, N305, N1208);
xor XOR2 (N1831, N1830, N889);
nor NOR4 (N1832, N1831, N1268, N629, N1);
nand NAND3 (N1833, N1828, N1694, N1670);
not NOT1 (N1834, N1823);
buf BUF1 (N1835, N1795);
and AND2 (N1836, N1821, N735);
nand NAND2 (N1837, N1836, N1733);
and AND2 (N1838, N1833, N1254);
nand NAND3 (N1839, N1838, N162, N356);
or OR4 (N1840, N1827, N1, N891, N162);
nor NOR3 (N1841, N1832, N867, N303);
xor XOR2 (N1842, N1840, N110);
not NOT1 (N1843, N1842);
nand NAND3 (N1844, N1834, N399, N598);
buf BUF1 (N1845, N1835);
buf BUF1 (N1846, N1845);
and AND3 (N1847, N1824, N490, N1821);
nor NOR2 (N1848, N1826, N904);
nor NOR2 (N1849, N1839, N1452);
nor NOR2 (N1850, N1848, N611);
or OR2 (N1851, N1829, N348);
buf BUF1 (N1852, N1849);
not NOT1 (N1853, N1843);
buf BUF1 (N1854, N1844);
or OR2 (N1855, N1853, N1185);
and AND2 (N1856, N1837, N270);
buf BUF1 (N1857, N1852);
xor XOR2 (N1858, N1856, N1773);
xor XOR2 (N1859, N1798, N122);
nand NAND3 (N1860, N1841, N633, N1409);
not NOT1 (N1861, N1847);
nand NAND2 (N1862, N1846, N1213);
nand NAND4 (N1863, N1861, N218, N840, N1844);
nand NAND3 (N1864, N1859, N693, N574);
nand NAND2 (N1865, N1858, N1522);
xor XOR2 (N1866, N1851, N1643);
nor NOR2 (N1867, N1860, N77);
buf BUF1 (N1868, N1855);
and AND2 (N1869, N1850, N1643);
nand NAND4 (N1870, N1867, N240, N358, N1514);
or OR4 (N1871, N1868, N1489, N374, N1832);
buf BUF1 (N1872, N1863);
nor NOR2 (N1873, N1857, N1402);
not NOT1 (N1874, N1864);
or OR2 (N1875, N1862, N506);
buf BUF1 (N1876, N1875);
xor XOR2 (N1877, N1854, N1209);
and AND3 (N1878, N1877, N267, N28);
and AND2 (N1879, N1865, N1455);
xor XOR2 (N1880, N1871, N431);
nor NOR3 (N1881, N1876, N1772, N425);
nor NOR3 (N1882, N1869, N140, N275);
or OR3 (N1883, N1881, N572, N64);
buf BUF1 (N1884, N1873);
xor XOR2 (N1885, N1872, N1337);
buf BUF1 (N1886, N1884);
and AND2 (N1887, N1883, N105);
not NOT1 (N1888, N1874);
or OR3 (N1889, N1882, N771, N1502);
nand NAND3 (N1890, N1887, N777, N1301);
xor XOR2 (N1891, N1879, N1699);
and AND3 (N1892, N1866, N1506, N1680);
not NOT1 (N1893, N1885);
or OR2 (N1894, N1891, N1653);
and AND2 (N1895, N1892, N9);
nand NAND4 (N1896, N1894, N1563, N1452, N281);
nand NAND3 (N1897, N1886, N956, N1785);
xor XOR2 (N1898, N1890, N856);
and AND3 (N1899, N1893, N410, N462);
nor NOR2 (N1900, N1898, N1447);
nand NAND4 (N1901, N1896, N1842, N1602, N1235);
xor XOR2 (N1902, N1889, N362);
nor NOR4 (N1903, N1888, N1464, N1166, N508);
or OR2 (N1904, N1900, N101);
not NOT1 (N1905, N1878);
or OR2 (N1906, N1902, N865);
nand NAND2 (N1907, N1904, N705);
buf BUF1 (N1908, N1880);
and AND3 (N1909, N1905, N1265, N578);
and AND2 (N1910, N1908, N174);
nor NOR4 (N1911, N1901, N782, N951, N227);
nor NOR4 (N1912, N1903, N856, N1870, N1654);
or OR4 (N1913, N768, N530, N807, N1454);
and AND2 (N1914, N1911, N1778);
and AND4 (N1915, N1912, N1330, N1364, N276);
buf BUF1 (N1916, N1910);
nand NAND3 (N1917, N1895, N551, N1442);
not NOT1 (N1918, N1907);
buf BUF1 (N1919, N1897);
buf BUF1 (N1920, N1916);
or OR4 (N1921, N1906, N955, N1332, N1821);
buf BUF1 (N1922, N1918);
and AND4 (N1923, N1922, N927, N333, N885);
nand NAND3 (N1924, N1919, N1439, N975);
nor NOR3 (N1925, N1921, N1364, N1775);
buf BUF1 (N1926, N1899);
not NOT1 (N1927, N1913);
not NOT1 (N1928, N1920);
or OR2 (N1929, N1909, N367);
nor NOR2 (N1930, N1926, N1164);
nor NOR3 (N1931, N1930, N170, N49);
xor XOR2 (N1932, N1924, N715);
or OR4 (N1933, N1932, N1353, N243, N194);
nor NOR2 (N1934, N1929, N737);
and AND3 (N1935, N1914, N571, N965);
and AND3 (N1936, N1935, N1813, N145);
nand NAND3 (N1937, N1923, N1247, N1249);
xor XOR2 (N1938, N1931, N943);
xor XOR2 (N1939, N1927, N1600);
buf BUF1 (N1940, N1937);
not NOT1 (N1941, N1917);
and AND2 (N1942, N1933, N521);
and AND3 (N1943, N1928, N1578, N1327);
nor NOR2 (N1944, N1943, N844);
and AND3 (N1945, N1925, N478, N421);
xor XOR2 (N1946, N1934, N979);
not NOT1 (N1947, N1946);
xor XOR2 (N1948, N1947, N1060);
xor XOR2 (N1949, N1939, N1602);
not NOT1 (N1950, N1948);
buf BUF1 (N1951, N1942);
and AND4 (N1952, N1949, N1499, N831, N1916);
or OR2 (N1953, N1941, N1819);
nand NAND3 (N1954, N1944, N1505, N932);
and AND2 (N1955, N1915, N258);
and AND3 (N1956, N1952, N731, N1825);
and AND2 (N1957, N1956, N1147);
and AND2 (N1958, N1954, N1951);
nand NAND2 (N1959, N859, N1387);
nor NOR2 (N1960, N1940, N1366);
xor XOR2 (N1961, N1953, N1347);
and AND3 (N1962, N1950, N1194, N1017);
xor XOR2 (N1963, N1957, N309);
xor XOR2 (N1964, N1960, N157);
xor XOR2 (N1965, N1958, N1287);
xor XOR2 (N1966, N1964, N596);
buf BUF1 (N1967, N1966);
nand NAND4 (N1968, N1963, N29, N1650, N1692);
or OR2 (N1969, N1945, N11);
nor NOR3 (N1970, N1959, N1352, N316);
not NOT1 (N1971, N1961);
and AND3 (N1972, N1971, N792, N1588);
and AND2 (N1973, N1938, N258);
nand NAND4 (N1974, N1955, N949, N318, N729);
not NOT1 (N1975, N1972);
and AND4 (N1976, N1968, N293, N1350, N521);
nand NAND3 (N1977, N1969, N900, N1585);
xor XOR2 (N1978, N1974, N1139);
buf BUF1 (N1979, N1965);
not NOT1 (N1980, N1970);
and AND4 (N1981, N1979, N1933, N1473, N1367);
nand NAND4 (N1982, N1975, N704, N910, N1442);
not NOT1 (N1983, N1977);
not NOT1 (N1984, N1980);
nand NAND3 (N1985, N1981, N1330, N1683);
or OR2 (N1986, N1976, N69);
or OR2 (N1987, N1984, N820);
buf BUF1 (N1988, N1985);
buf BUF1 (N1989, N1978);
and AND4 (N1990, N1936, N401, N1549, N935);
xor XOR2 (N1991, N1986, N710);
nor NOR2 (N1992, N1991, N1341);
or OR3 (N1993, N1987, N595, N1106);
nor NOR4 (N1994, N1982, N1800, N544, N1672);
or OR4 (N1995, N1990, N1677, N1687, N154);
not NOT1 (N1996, N1962);
or OR2 (N1997, N1996, N1408);
and AND2 (N1998, N1989, N1365);
or OR2 (N1999, N1973, N271);
or OR2 (N2000, N1995, N260);
nor NOR4 (N2001, N1967, N1986, N1381, N522);
xor XOR2 (N2002, N1997, N1836);
and AND4 (N2003, N1993, N651, N1536, N1599);
and AND2 (N2004, N1999, N1319);
and AND4 (N2005, N1983, N588, N519, N1554);
and AND4 (N2006, N2003, N1435, N1657, N1009);
xor XOR2 (N2007, N2000, N1332);
and AND4 (N2008, N1998, N1295, N1523, N764);
not NOT1 (N2009, N1994);
buf BUF1 (N2010, N2007);
nand NAND3 (N2011, N2005, N1855, N1247);
and AND3 (N2012, N2006, N656, N539);
xor XOR2 (N2013, N1988, N1247);
xor XOR2 (N2014, N2012, N1591);
buf BUF1 (N2015, N2014);
and AND2 (N2016, N1992, N1538);
buf BUF1 (N2017, N2002);
buf BUF1 (N2018, N2010);
nor NOR2 (N2019, N2011, N1223);
and AND4 (N2020, N2013, N1302, N1134, N862);
or OR3 (N2021, N2009, N81, N1876);
not NOT1 (N2022, N2019);
nor NOR2 (N2023, N2016, N253);
buf BUF1 (N2024, N2008);
xor XOR2 (N2025, N2018, N558);
and AND3 (N2026, N2015, N1764, N1471);
or OR3 (N2027, N2024, N756, N1957);
buf BUF1 (N2028, N2004);
nor NOR2 (N2029, N2022, N1603);
xor XOR2 (N2030, N2025, N1077);
nand NAND3 (N2031, N2028, N685, N1025);
nand NAND2 (N2032, N2031, N1165);
nor NOR3 (N2033, N2023, N939, N1446);
buf BUF1 (N2034, N2026);
buf BUF1 (N2035, N2020);
nor NOR3 (N2036, N2034, N1722, N1622);
xor XOR2 (N2037, N2035, N1947);
or OR2 (N2038, N2029, N1711);
xor XOR2 (N2039, N2001, N681);
buf BUF1 (N2040, N2027);
xor XOR2 (N2041, N2038, N1457);
nand NAND2 (N2042, N2033, N881);
or OR3 (N2043, N2039, N671, N332);
xor XOR2 (N2044, N2042, N600);
nand NAND2 (N2045, N2043, N371);
nor NOR3 (N2046, N2044, N1613, N169);
not NOT1 (N2047, N2017);
and AND3 (N2048, N2021, N457, N1630);
buf BUF1 (N2049, N2036);
not NOT1 (N2050, N2040);
or OR2 (N2051, N2045, N2014);
xor XOR2 (N2052, N2051, N57);
xor XOR2 (N2053, N2049, N892);
buf BUF1 (N2054, N2041);
nand NAND3 (N2055, N2053, N379, N1973);
nor NOR4 (N2056, N2047, N815, N1769, N292);
or OR4 (N2057, N2030, N1341, N1187, N1041);
xor XOR2 (N2058, N2032, N1303);
or OR3 (N2059, N2050, N1654, N441);
not NOT1 (N2060, N2046);
and AND3 (N2061, N2052, N1960, N568);
nand NAND4 (N2062, N2058, N496, N1598, N506);
or OR4 (N2063, N2055, N2032, N1479, N1169);
buf BUF1 (N2064, N2062);
not NOT1 (N2065, N2048);
nand NAND2 (N2066, N2065, N843);
and AND3 (N2067, N2064, N667, N1186);
nand NAND3 (N2068, N2066, N656, N1706);
buf BUF1 (N2069, N2067);
nor NOR2 (N2070, N2054, N465);
xor XOR2 (N2071, N2063, N2031);
xor XOR2 (N2072, N2059, N1023);
or OR3 (N2073, N2071, N1245, N999);
nor NOR2 (N2074, N2069, N1829);
or OR3 (N2075, N2037, N1421, N2019);
and AND4 (N2076, N2057, N1218, N813, N761);
xor XOR2 (N2077, N2060, N187);
buf BUF1 (N2078, N2075);
nor NOR3 (N2079, N2078, N1748, N681);
xor XOR2 (N2080, N2056, N1088);
buf BUF1 (N2081, N2072);
xor XOR2 (N2082, N2073, N746);
not NOT1 (N2083, N2080);
nor NOR3 (N2084, N2082, N1895, N565);
not NOT1 (N2085, N2076);
buf BUF1 (N2086, N2085);
not NOT1 (N2087, N2068);
nor NOR4 (N2088, N2084, N1689, N2001, N313);
not NOT1 (N2089, N2077);
buf BUF1 (N2090, N2088);
xor XOR2 (N2091, N2090, N213);
nor NOR3 (N2092, N2086, N1300, N1516);
and AND4 (N2093, N2092, N644, N1785, N1470);
nand NAND2 (N2094, N2070, N1149);
and AND3 (N2095, N2074, N1041, N1654);
and AND4 (N2096, N2079, N1889, N1439, N727);
nor NOR3 (N2097, N2093, N1684, N1529);
nand NAND2 (N2098, N2096, N1473);
or OR4 (N2099, N2083, N1147, N150, N684);
and AND2 (N2100, N2094, N91);
nand NAND4 (N2101, N2081, N2023, N868, N746);
or OR4 (N2102, N2101, N1897, N513, N229);
not NOT1 (N2103, N2097);
buf BUF1 (N2104, N2061);
nand NAND4 (N2105, N2103, N1939, N1573, N335);
or OR2 (N2106, N2095, N807);
or OR3 (N2107, N2099, N659, N955);
nand NAND2 (N2108, N2102, N1700);
nand NAND4 (N2109, N2089, N1839, N434, N1692);
buf BUF1 (N2110, N2087);
or OR4 (N2111, N2104, N1301, N1073, N428);
xor XOR2 (N2112, N2098, N54);
and AND4 (N2113, N2107, N23, N411, N2100);
buf BUF1 (N2114, N942);
or OR2 (N2115, N2113, N790);
and AND4 (N2116, N2114, N995, N88, N1029);
and AND4 (N2117, N2105, N1887, N862, N619);
nor NOR3 (N2118, N2112, N1088, N2031);
and AND4 (N2119, N2117, N46, N1663, N982);
and AND4 (N2120, N2111, N1639, N954, N456);
not NOT1 (N2121, N2118);
not NOT1 (N2122, N2110);
or OR3 (N2123, N2108, N345, N1564);
nor NOR4 (N2124, N2120, N190, N1119, N233);
or OR2 (N2125, N2116, N565);
and AND2 (N2126, N2121, N975);
xor XOR2 (N2127, N2126, N228);
buf BUF1 (N2128, N2127);
or OR3 (N2129, N2115, N216, N1566);
and AND2 (N2130, N2119, N106);
buf BUF1 (N2131, N2109);
and AND3 (N2132, N2129, N1938, N434);
xor XOR2 (N2133, N2091, N1549);
not NOT1 (N2134, N2122);
not NOT1 (N2135, N2125);
and AND2 (N2136, N2133, N1075);
or OR4 (N2137, N2123, N1849, N1761, N663);
or OR2 (N2138, N2124, N644);
and AND3 (N2139, N2131, N365, N1909);
buf BUF1 (N2140, N2136);
nor NOR4 (N2141, N2132, N358, N879, N712);
nor NOR2 (N2142, N2141, N365);
nor NOR4 (N2143, N2106, N930, N1001, N2141);
and AND2 (N2144, N2137, N2002);
buf BUF1 (N2145, N2128);
and AND2 (N2146, N2142, N1294);
buf BUF1 (N2147, N2140);
nor NOR2 (N2148, N2147, N113);
xor XOR2 (N2149, N2130, N1395);
nor NOR2 (N2150, N2139, N215);
buf BUF1 (N2151, N2148);
nand NAND2 (N2152, N2143, N1172);
xor XOR2 (N2153, N2152, N1998);
and AND3 (N2154, N2150, N1913, N191);
buf BUF1 (N2155, N2144);
buf BUF1 (N2156, N2138);
xor XOR2 (N2157, N2155, N268);
and AND3 (N2158, N2151, N1816, N697);
and AND3 (N2159, N2157, N1614, N1911);
buf BUF1 (N2160, N2154);
nand NAND4 (N2161, N2146, N2125, N842, N286);
buf BUF1 (N2162, N2153);
and AND4 (N2163, N2161, N2118, N221, N380);
nor NOR4 (N2164, N2160, N575, N1530, N1846);
and AND3 (N2165, N2134, N732, N1555);
and AND3 (N2166, N2149, N2015, N1724);
xor XOR2 (N2167, N2159, N1771);
nand NAND3 (N2168, N2135, N2066, N1298);
or OR3 (N2169, N2166, N362, N1737);
and AND2 (N2170, N2162, N2017);
buf BUF1 (N2171, N2167);
or OR2 (N2172, N2165, N265);
and AND4 (N2173, N2172, N262, N131, N1239);
nor NOR4 (N2174, N2170, N792, N1996, N664);
not NOT1 (N2175, N2158);
xor XOR2 (N2176, N2168, N2035);
not NOT1 (N2177, N2164);
and AND4 (N2178, N2176, N553, N2106, N1822);
buf BUF1 (N2179, N2156);
nand NAND4 (N2180, N2177, N472, N1689, N827);
buf BUF1 (N2181, N2171);
buf BUF1 (N2182, N2169);
nand NAND4 (N2183, N2178, N211, N1793, N623);
and AND4 (N2184, N2145, N1513, N683, N51);
xor XOR2 (N2185, N2179, N2017);
buf BUF1 (N2186, N2180);
not NOT1 (N2187, N2173);
nand NAND3 (N2188, N2182, N1909, N1029);
buf BUF1 (N2189, N2175);
nand NAND4 (N2190, N2188, N318, N1595, N498);
nor NOR2 (N2191, N2187, N1347);
buf BUF1 (N2192, N2189);
nor NOR3 (N2193, N2174, N554, N1432);
nor NOR3 (N2194, N2185, N1079, N221);
and AND3 (N2195, N2194, N2012, N608);
nor NOR2 (N2196, N2192, N570);
xor XOR2 (N2197, N2196, N1878);
nor NOR4 (N2198, N2163, N1231, N1188, N1957);
and AND3 (N2199, N2195, N1390, N325);
not NOT1 (N2200, N2197);
xor XOR2 (N2201, N2199, N773);
or OR4 (N2202, N2198, N553, N1236, N833);
nor NOR2 (N2203, N2186, N641);
and AND3 (N2204, N2181, N2157, N1863);
xor XOR2 (N2205, N2190, N401);
and AND2 (N2206, N2184, N578);
not NOT1 (N2207, N2191);
nand NAND2 (N2208, N2206, N919);
not NOT1 (N2209, N2203);
buf BUF1 (N2210, N2208);
nand NAND4 (N2211, N2202, N947, N113, N936);
buf BUF1 (N2212, N2204);
not NOT1 (N2213, N2205);
buf BUF1 (N2214, N2207);
xor XOR2 (N2215, N2213, N565);
nand NAND2 (N2216, N2200, N2024);
or OR3 (N2217, N2210, N702, N1692);
and AND3 (N2218, N2183, N1397, N1171);
or OR3 (N2219, N2211, N1926, N1324);
buf BUF1 (N2220, N2201);
not NOT1 (N2221, N2193);
xor XOR2 (N2222, N2219, N942);
and AND3 (N2223, N2221, N853, N573);
xor XOR2 (N2224, N2212, N1312);
nand NAND4 (N2225, N2220, N999, N2222, N37);
xor XOR2 (N2226, N714, N2222);
nand NAND3 (N2227, N2224, N476, N1405);
or OR2 (N2228, N2215, N1205);
buf BUF1 (N2229, N2209);
or OR3 (N2230, N2223, N301, N2066);
buf BUF1 (N2231, N2228);
xor XOR2 (N2232, N2230, N1423);
or OR3 (N2233, N2232, N550, N95);
nand NAND3 (N2234, N2227, N909, N1412);
and AND2 (N2235, N2217, N1518);
nand NAND3 (N2236, N2229, N702, N1668);
not NOT1 (N2237, N2226);
and AND3 (N2238, N2214, N436, N1250);
or OR4 (N2239, N2238, N375, N979, N56);
nor NOR2 (N2240, N2234, N1559);
and AND3 (N2241, N2218, N302, N1977);
not NOT1 (N2242, N2225);
nand NAND3 (N2243, N2237, N2174, N1200);
or OR4 (N2244, N2240, N1529, N461, N119);
xor XOR2 (N2245, N2216, N1833);
and AND2 (N2246, N2241, N1354);
xor XOR2 (N2247, N2245, N2157);
xor XOR2 (N2248, N2246, N1316);
nor NOR3 (N2249, N2247, N2154, N190);
or OR3 (N2250, N2239, N1229, N704);
nor NOR3 (N2251, N2250, N2132, N797);
or OR2 (N2252, N2236, N1915);
and AND2 (N2253, N2235, N479);
or OR3 (N2254, N2242, N197, N1865);
buf BUF1 (N2255, N2231);
buf BUF1 (N2256, N2249);
xor XOR2 (N2257, N2256, N1752);
and AND2 (N2258, N2248, N2191);
or OR2 (N2259, N2258, N380);
nor NOR4 (N2260, N2255, N105, N447, N1474);
not NOT1 (N2261, N2253);
or OR4 (N2262, N2254, N1836, N852, N507);
xor XOR2 (N2263, N2243, N1868);
not NOT1 (N2264, N2259);
or OR4 (N2265, N2233, N2190, N1166, N1454);
buf BUF1 (N2266, N2261);
or OR2 (N2267, N2265, N2165);
nor NOR3 (N2268, N2257, N1366, N2084);
nand NAND4 (N2269, N2266, N573, N1351, N2238);
and AND2 (N2270, N2251, N676);
xor XOR2 (N2271, N2267, N753);
not NOT1 (N2272, N2271);
xor XOR2 (N2273, N2268, N1287);
not NOT1 (N2274, N2262);
and AND4 (N2275, N2269, N1865, N1402, N1138);
and AND3 (N2276, N2264, N1284, N1734);
or OR3 (N2277, N2273, N743, N852);
xor XOR2 (N2278, N2274, N507);
nor NOR3 (N2279, N2244, N571, N1695);
nand NAND2 (N2280, N2270, N1761);
nor NOR2 (N2281, N2263, N301);
or OR3 (N2282, N2277, N680, N490);
not NOT1 (N2283, N2278);
nor NOR4 (N2284, N2283, N344, N833, N495);
nor NOR3 (N2285, N2282, N1670, N1565);
not NOT1 (N2286, N2279);
nand NAND2 (N2287, N2252, N1873);
buf BUF1 (N2288, N2260);
nand NAND4 (N2289, N2276, N812, N1350, N1105);
or OR2 (N2290, N2272, N87);
or OR3 (N2291, N2275, N1235, N979);
or OR3 (N2292, N2289, N1544, N1440);
nand NAND4 (N2293, N2292, N1798, N106, N632);
buf BUF1 (N2294, N2290);
and AND4 (N2295, N2287, N1452, N692, N1845);
xor XOR2 (N2296, N2280, N1525);
buf BUF1 (N2297, N2296);
nor NOR4 (N2298, N2281, N2143, N641, N2160);
nor NOR3 (N2299, N2297, N1398, N539);
nand NAND2 (N2300, N2293, N2100);
not NOT1 (N2301, N2299);
nand NAND4 (N2302, N2294, N739, N68, N227);
xor XOR2 (N2303, N2295, N1092);
nor NOR2 (N2304, N2286, N334);
and AND2 (N2305, N2288, N1432);
not NOT1 (N2306, N2291);
nor NOR2 (N2307, N2305, N194);
nor NOR4 (N2308, N2298, N346, N1871, N196);
xor XOR2 (N2309, N2304, N2019);
nand NAND2 (N2310, N2306, N1463);
nor NOR4 (N2311, N2301, N2183, N1349, N1849);
or OR4 (N2312, N2302, N1320, N1034, N1838);
and AND2 (N2313, N2285, N244);
not NOT1 (N2314, N2311);
xor XOR2 (N2315, N2312, N2183);
or OR4 (N2316, N2315, N2258, N597, N681);
and AND3 (N2317, N2307, N2226, N610);
nor NOR4 (N2318, N2284, N1418, N2078, N1850);
nand NAND2 (N2319, N2303, N1899);
buf BUF1 (N2320, N2319);
buf BUF1 (N2321, N2310);
xor XOR2 (N2322, N2309, N1637);
buf BUF1 (N2323, N2308);
and AND4 (N2324, N2322, N1028, N1824, N2025);
nor NOR3 (N2325, N2313, N1519, N927);
nand NAND3 (N2326, N2318, N2011, N240);
nor NOR2 (N2327, N2321, N1982);
buf BUF1 (N2328, N2320);
xor XOR2 (N2329, N2316, N2318);
xor XOR2 (N2330, N2329, N1501);
buf BUF1 (N2331, N2317);
not NOT1 (N2332, N2324);
buf BUF1 (N2333, N2314);
or OR3 (N2334, N2325, N290, N2181);
nor NOR3 (N2335, N2326, N519, N477);
xor XOR2 (N2336, N2330, N1671);
and AND3 (N2337, N2323, N20, N33);
and AND2 (N2338, N2327, N1604);
nand NAND3 (N2339, N2337, N1673, N1081);
nand NAND2 (N2340, N2328, N680);
nand NAND4 (N2341, N2340, N2178, N623, N386);
buf BUF1 (N2342, N2341);
buf BUF1 (N2343, N2334);
nor NOR3 (N2344, N2338, N1062, N341);
and AND3 (N2345, N2332, N736, N1391);
xor XOR2 (N2346, N2343, N989);
xor XOR2 (N2347, N2345, N288);
or OR2 (N2348, N2336, N693);
or OR3 (N2349, N2346, N477, N2309);
buf BUF1 (N2350, N2331);
or OR3 (N2351, N2350, N1716, N731);
and AND2 (N2352, N2348, N1776);
buf BUF1 (N2353, N2351);
buf BUF1 (N2354, N2344);
and AND3 (N2355, N2352, N2189, N2059);
or OR2 (N2356, N2349, N369);
and AND2 (N2357, N2339, N1382);
not NOT1 (N2358, N2347);
not NOT1 (N2359, N2300);
xor XOR2 (N2360, N2333, N2017);
or OR3 (N2361, N2360, N555, N1809);
buf BUF1 (N2362, N2358);
and AND4 (N2363, N2359, N1437, N304, N1032);
buf BUF1 (N2364, N2361);
nand NAND4 (N2365, N2356, N665, N1644, N270);
and AND2 (N2366, N2342, N2323);
and AND3 (N2367, N2362, N553, N1396);
buf BUF1 (N2368, N2367);
not NOT1 (N2369, N2368);
xor XOR2 (N2370, N2355, N1490);
or OR4 (N2371, N2354, N679, N987, N982);
buf BUF1 (N2372, N2335);
buf BUF1 (N2373, N2364);
xor XOR2 (N2374, N2372, N773);
buf BUF1 (N2375, N2374);
nand NAND2 (N2376, N2369, N655);
buf BUF1 (N2377, N2357);
nor NOR4 (N2378, N2363, N375, N427, N2051);
buf BUF1 (N2379, N2375);
or OR2 (N2380, N2353, N2148);
nor NOR2 (N2381, N2380, N617);
nand NAND3 (N2382, N2377, N1080, N1724);
buf BUF1 (N2383, N2381);
xor XOR2 (N2384, N2376, N1943);
or OR2 (N2385, N2373, N80);
nand NAND2 (N2386, N2383, N1770);
xor XOR2 (N2387, N2386, N10);
buf BUF1 (N2388, N2365);
buf BUF1 (N2389, N2379);
and AND3 (N2390, N2389, N2295, N1027);
not NOT1 (N2391, N2384);
not NOT1 (N2392, N2371);
xor XOR2 (N2393, N2370, N541);
or OR4 (N2394, N2391, N665, N1990, N1440);
buf BUF1 (N2395, N2387);
not NOT1 (N2396, N2378);
xor XOR2 (N2397, N2395, N329);
xor XOR2 (N2398, N2397, N2179);
xor XOR2 (N2399, N2393, N1449);
or OR4 (N2400, N2385, N1678, N1356, N1774);
nor NOR4 (N2401, N2400, N2131, N1425, N1834);
xor XOR2 (N2402, N2399, N457);
nand NAND4 (N2403, N2402, N857, N1891, N1484);
or OR3 (N2404, N2396, N631, N186);
and AND4 (N2405, N2382, N453, N555, N2400);
xor XOR2 (N2406, N2404, N2015);
nand NAND2 (N2407, N2403, N1720);
and AND4 (N2408, N2405, N1611, N1179, N1733);
nand NAND3 (N2409, N2388, N629, N902);
not NOT1 (N2410, N2409);
not NOT1 (N2411, N2410);
and AND3 (N2412, N2366, N2306, N1746);
or OR3 (N2413, N2406, N2321, N415);
buf BUF1 (N2414, N2401);
and AND2 (N2415, N2398, N517);
nand NAND2 (N2416, N2411, N139);
and AND4 (N2417, N2392, N1594, N2118, N290);
xor XOR2 (N2418, N2417, N1906);
xor XOR2 (N2419, N2414, N846);
buf BUF1 (N2420, N2419);
buf BUF1 (N2421, N2413);
buf BUF1 (N2422, N2394);
or OR4 (N2423, N2415, N872, N1623, N496);
xor XOR2 (N2424, N2407, N819);
nand NAND4 (N2425, N2423, N2, N2020, N686);
and AND3 (N2426, N2418, N394, N742);
nor NOR4 (N2427, N2426, N921, N1502, N2158);
nor NOR2 (N2428, N2421, N2310);
nand NAND4 (N2429, N2416, N183, N330, N419);
xor XOR2 (N2430, N2422, N1915);
xor XOR2 (N2431, N2390, N2212);
nor NOR3 (N2432, N2412, N1402, N1578);
buf BUF1 (N2433, N2408);
or OR4 (N2434, N2430, N2237, N805, N764);
buf BUF1 (N2435, N2433);
or OR3 (N2436, N2432, N242, N325);
not NOT1 (N2437, N2436);
or OR3 (N2438, N2437, N187, N91);
xor XOR2 (N2439, N2427, N1379);
buf BUF1 (N2440, N2425);
and AND2 (N2441, N2431, N446);
not NOT1 (N2442, N2434);
xor XOR2 (N2443, N2441, N1956);
not NOT1 (N2444, N2428);
not NOT1 (N2445, N2442);
buf BUF1 (N2446, N2435);
nor NOR4 (N2447, N2443, N1036, N925, N80);
or OR2 (N2448, N2429, N936);
xor XOR2 (N2449, N2444, N502);
xor XOR2 (N2450, N2447, N747);
not NOT1 (N2451, N2450);
and AND3 (N2452, N2449, N829, N914);
nand NAND3 (N2453, N2420, N2177, N329);
nand NAND3 (N2454, N2439, N1246, N2401);
xor XOR2 (N2455, N2424, N295);
nor NOR4 (N2456, N2453, N982, N963, N161);
or OR4 (N2457, N2451, N2346, N2029, N2308);
buf BUF1 (N2458, N2452);
nand NAND2 (N2459, N2445, N1852);
xor XOR2 (N2460, N2448, N504);
or OR2 (N2461, N2455, N2414);
buf BUF1 (N2462, N2458);
and AND2 (N2463, N2460, N1979);
buf BUF1 (N2464, N2454);
xor XOR2 (N2465, N2440, N2189);
xor XOR2 (N2466, N2462, N33);
xor XOR2 (N2467, N2464, N1539);
not NOT1 (N2468, N2467);
not NOT1 (N2469, N2468);
nand NAND2 (N2470, N2469, N261);
nand NAND4 (N2471, N2456, N597, N1792, N1922);
nor NOR2 (N2472, N2465, N1521);
nand NAND2 (N2473, N2461, N1220);
not NOT1 (N2474, N2463);
nor NOR4 (N2475, N2472, N2242, N1358, N1978);
nand NAND4 (N2476, N2457, N1604, N2352, N2041);
xor XOR2 (N2477, N2474, N1217);
xor XOR2 (N2478, N2471, N1114);
not NOT1 (N2479, N2477);
xor XOR2 (N2480, N2459, N2179);
not NOT1 (N2481, N2466);
buf BUF1 (N2482, N2446);
xor XOR2 (N2483, N2438, N753);
not NOT1 (N2484, N2470);
or OR3 (N2485, N2482, N2297, N45);
or OR4 (N2486, N2484, N2048, N800, N2184);
and AND3 (N2487, N2480, N1428, N1436);
not NOT1 (N2488, N2481);
or OR2 (N2489, N2486, N1294);
buf BUF1 (N2490, N2487);
and AND2 (N2491, N2479, N1265);
nor NOR4 (N2492, N2489, N156, N885, N380);
xor XOR2 (N2493, N2490, N2453);
and AND3 (N2494, N2473, N678, N2265);
not NOT1 (N2495, N2494);
xor XOR2 (N2496, N2492, N2024);
buf BUF1 (N2497, N2476);
nor NOR4 (N2498, N2478, N134, N867, N693);
or OR2 (N2499, N2485, N2487);
or OR3 (N2500, N2491, N170, N2199);
or OR2 (N2501, N2495, N883);
nand NAND2 (N2502, N2500, N1524);
nand NAND3 (N2503, N2497, N120, N2419);
not NOT1 (N2504, N2496);
nor NOR4 (N2505, N2499, N2218, N508, N324);
not NOT1 (N2506, N2503);
and AND4 (N2507, N2505, N1427, N2395, N2430);
not NOT1 (N2508, N2483);
not NOT1 (N2509, N2501);
buf BUF1 (N2510, N2498);
xor XOR2 (N2511, N2504, N2030);
not NOT1 (N2512, N2493);
nand NAND4 (N2513, N2508, N842, N1673, N400);
nor NOR3 (N2514, N2488, N1640, N792);
nor NOR3 (N2515, N2512, N3, N2099);
buf BUF1 (N2516, N2506);
xor XOR2 (N2517, N2513, N1587);
and AND3 (N2518, N2514, N1555, N1363);
and AND3 (N2519, N2475, N1985, N2187);
not NOT1 (N2520, N2510);
nor NOR3 (N2521, N2520, N1687, N1961);
not NOT1 (N2522, N2518);
xor XOR2 (N2523, N2517, N2230);
not NOT1 (N2524, N2516);
or OR2 (N2525, N2522, N1413);
and AND3 (N2526, N2519, N1965, N1973);
and AND2 (N2527, N2509, N1760);
xor XOR2 (N2528, N2521, N2232);
xor XOR2 (N2529, N2523, N1387);
nor NOR2 (N2530, N2527, N1600);
not NOT1 (N2531, N2526);
xor XOR2 (N2532, N2502, N505);
xor XOR2 (N2533, N2515, N1356);
and AND2 (N2534, N2511, N492);
not NOT1 (N2535, N2532);
or OR2 (N2536, N2533, N1078);
buf BUF1 (N2537, N2535);
nor NOR4 (N2538, N2536, N490, N2004, N266);
or OR2 (N2539, N2530, N298);
not NOT1 (N2540, N2525);
xor XOR2 (N2541, N2538, N1205);
nor NOR3 (N2542, N2507, N1892, N2041);
or OR3 (N2543, N2541, N394, N1069);
buf BUF1 (N2544, N2537);
nand NAND3 (N2545, N2540, N1516, N2350);
nand NAND3 (N2546, N2539, N1069, N1865);
buf BUF1 (N2547, N2543);
xor XOR2 (N2548, N2546, N2164);
and AND4 (N2549, N2524, N1582, N137, N214);
and AND3 (N2550, N2549, N1667, N645);
buf BUF1 (N2551, N2529);
or OR4 (N2552, N2534, N241, N774, N1975);
xor XOR2 (N2553, N2545, N1981);
nor NOR2 (N2554, N2552, N2245);
buf BUF1 (N2555, N2554);
nor NOR4 (N2556, N2550, N1815, N732, N2019);
or OR4 (N2557, N2528, N756, N2338, N480);
not NOT1 (N2558, N2547);
buf BUF1 (N2559, N2548);
and AND3 (N2560, N2542, N2359, N127);
or OR2 (N2561, N2551, N2100);
nor NOR2 (N2562, N2544, N2359);
xor XOR2 (N2563, N2561, N1540);
nand NAND3 (N2564, N2557, N2074, N771);
and AND3 (N2565, N2562, N899, N650);
not NOT1 (N2566, N2556);
buf BUF1 (N2567, N2555);
buf BUF1 (N2568, N2559);
nor NOR3 (N2569, N2558, N952, N2359);
nand NAND2 (N2570, N2560, N1324);
buf BUF1 (N2571, N2565);
nor NOR3 (N2572, N2568, N493, N1790);
xor XOR2 (N2573, N2571, N2468);
not NOT1 (N2574, N2569);
xor XOR2 (N2575, N2573, N1285);
nor NOR3 (N2576, N2563, N774, N189);
xor XOR2 (N2577, N2566, N543);
not NOT1 (N2578, N2575);
nand NAND4 (N2579, N2570, N1020, N1190, N1361);
buf BUF1 (N2580, N2572);
xor XOR2 (N2581, N2580, N1164);
not NOT1 (N2582, N2553);
not NOT1 (N2583, N2567);
nand NAND4 (N2584, N2564, N2180, N1439, N982);
buf BUF1 (N2585, N2577);
nand NAND4 (N2586, N2579, N708, N1143, N209);
not NOT1 (N2587, N2586);
nor NOR3 (N2588, N2531, N1570, N479);
nand NAND4 (N2589, N2574, N348, N759, N1312);
not NOT1 (N2590, N2584);
nor NOR2 (N2591, N2590, N159);
xor XOR2 (N2592, N2587, N1652);
buf BUF1 (N2593, N2591);
or OR2 (N2594, N2593, N1733);
buf BUF1 (N2595, N2585);
not NOT1 (N2596, N2588);
buf BUF1 (N2597, N2595);
not NOT1 (N2598, N2594);
xor XOR2 (N2599, N2581, N2060);
nor NOR4 (N2600, N2589, N1592, N1676, N1119);
nor NOR4 (N2601, N2592, N1744, N98, N1123);
nand NAND3 (N2602, N2578, N685, N120);
and AND3 (N2603, N2597, N997, N496);
buf BUF1 (N2604, N2599);
not NOT1 (N2605, N2602);
and AND2 (N2606, N2601, N2513);
or OR3 (N2607, N2583, N2229, N2321);
xor XOR2 (N2608, N2604, N563);
or OR3 (N2609, N2607, N2252, N2344);
not NOT1 (N2610, N2609);
nand NAND3 (N2611, N2600, N54, N1818);
xor XOR2 (N2612, N2598, N1891);
buf BUF1 (N2613, N2576);
not NOT1 (N2614, N2605);
not NOT1 (N2615, N2596);
and AND2 (N2616, N2612, N516);
and AND4 (N2617, N2616, N1895, N2233, N1625);
xor XOR2 (N2618, N2614, N1815);
and AND3 (N2619, N2617, N2360, N484);
nand NAND4 (N2620, N2603, N120, N1949, N2443);
and AND4 (N2621, N2618, N2390, N2403, N1035);
not NOT1 (N2622, N2611);
nor NOR4 (N2623, N2615, N2531, N73, N21);
buf BUF1 (N2624, N2622);
or OR4 (N2625, N2582, N170, N2028, N1923);
buf BUF1 (N2626, N2610);
nor NOR4 (N2627, N2608, N1728, N2093, N2592);
nand NAND4 (N2628, N2625, N985, N1657, N867);
buf BUF1 (N2629, N2606);
not NOT1 (N2630, N2626);
nand NAND3 (N2631, N2630, N2146, N229);
not NOT1 (N2632, N2624);
xor XOR2 (N2633, N2632, N1489);
and AND2 (N2634, N2619, N2229);
nand NAND2 (N2635, N2634, N678);
and AND2 (N2636, N2620, N1216);
and AND2 (N2637, N2613, N154);
nor NOR2 (N2638, N2627, N2294);
xor XOR2 (N2639, N2621, N1565);
nor NOR2 (N2640, N2639, N694);
buf BUF1 (N2641, N2637);
not NOT1 (N2642, N2629);
not NOT1 (N2643, N2642);
xor XOR2 (N2644, N2636, N1682);
and AND4 (N2645, N2631, N1091, N930, N548);
nor NOR3 (N2646, N2643, N520, N1134);
and AND4 (N2647, N2623, N372, N191, N1782);
not NOT1 (N2648, N2635);
or OR2 (N2649, N2640, N907);
nand NAND2 (N2650, N2648, N1176);
nand NAND4 (N2651, N2646, N723, N1953, N1222);
nor NOR2 (N2652, N2650, N1029);
buf BUF1 (N2653, N2638);
and AND4 (N2654, N2641, N1549, N102, N174);
nand NAND4 (N2655, N2654, N1571, N2641, N2123);
xor XOR2 (N2656, N2628, N1298);
and AND4 (N2657, N2644, N1284, N221, N2642);
buf BUF1 (N2658, N2633);
nand NAND3 (N2659, N2657, N800, N1218);
nor NOR4 (N2660, N2645, N1371, N557, N1475);
nor NOR2 (N2661, N2651, N146);
or OR3 (N2662, N2653, N1294, N1028);
xor XOR2 (N2663, N2656, N1297);
or OR4 (N2664, N2655, N217, N1116, N2173);
buf BUF1 (N2665, N2649);
and AND3 (N2666, N2664, N68, N1479);
buf BUF1 (N2667, N2663);
xor XOR2 (N2668, N2659, N84);
not NOT1 (N2669, N2668);
not NOT1 (N2670, N2647);
or OR2 (N2671, N2665, N586);
and AND3 (N2672, N2669, N879, N445);
nand NAND4 (N2673, N2666, N2070, N913, N203);
or OR3 (N2674, N2670, N2093, N2470);
xor XOR2 (N2675, N2658, N1056);
nand NAND4 (N2676, N2671, N649, N1469, N1446);
nor NOR3 (N2677, N2660, N2240, N1653);
xor XOR2 (N2678, N2661, N41);
and AND2 (N2679, N2676, N1012);
not NOT1 (N2680, N2675);
not NOT1 (N2681, N2673);
or OR2 (N2682, N2672, N1812);
xor XOR2 (N2683, N2678, N484);
buf BUF1 (N2684, N2667);
xor XOR2 (N2685, N2681, N1805);
or OR4 (N2686, N2662, N981, N216, N961);
or OR4 (N2687, N2682, N1432, N737, N1735);
xor XOR2 (N2688, N2652, N2022);
nor NOR4 (N2689, N2686, N1445, N1870, N1807);
xor XOR2 (N2690, N2680, N1898);
or OR3 (N2691, N2689, N923, N698);
and AND4 (N2692, N2674, N1009, N1192, N851);
and AND4 (N2693, N2692, N1637, N1644, N386);
and AND3 (N2694, N2690, N1152, N1710);
buf BUF1 (N2695, N2684);
and AND2 (N2696, N2679, N1154);
or OR2 (N2697, N2677, N825);
xor XOR2 (N2698, N2685, N1180);
nand NAND3 (N2699, N2698, N403, N499);
not NOT1 (N2700, N2695);
nand NAND3 (N2701, N2683, N1836, N2540);
and AND2 (N2702, N2691, N2277);
buf BUF1 (N2703, N2688);
nor NOR3 (N2704, N2687, N1832, N178);
or OR3 (N2705, N2703, N627, N556);
nand NAND4 (N2706, N2699, N1532, N2036, N781);
or OR4 (N2707, N2693, N66, N1671, N863);
and AND4 (N2708, N2706, N423, N1354, N408);
nor NOR2 (N2709, N2696, N1735);
xor XOR2 (N2710, N2700, N1130);
and AND2 (N2711, N2701, N2458);
and AND4 (N2712, N2694, N1502, N923, N1373);
nand NAND4 (N2713, N2711, N46, N1009, N2396);
nor NOR4 (N2714, N2713, N2, N601, N306);
not NOT1 (N2715, N2712);
buf BUF1 (N2716, N2708);
and AND4 (N2717, N2702, N2667, N1626, N933);
not NOT1 (N2718, N2704);
not NOT1 (N2719, N2707);
buf BUF1 (N2720, N2697);
buf BUF1 (N2721, N2710);
or OR4 (N2722, N2705, N605, N2583, N592);
or OR4 (N2723, N2715, N1436, N2465, N1121);
or OR3 (N2724, N2723, N1333, N1590);
nand NAND4 (N2725, N2709, N1741, N575, N1351);
nand NAND3 (N2726, N2716, N43, N704);
nor NOR4 (N2727, N2724, N250, N2432, N591);
buf BUF1 (N2728, N2720);
buf BUF1 (N2729, N2714);
xor XOR2 (N2730, N2718, N866);
and AND3 (N2731, N2721, N107, N1084);
nor NOR4 (N2732, N2730, N2671, N499, N2360);
not NOT1 (N2733, N2731);
and AND4 (N2734, N2725, N2462, N2402, N415);
or OR2 (N2735, N2719, N209);
buf BUF1 (N2736, N2735);
not NOT1 (N2737, N2727);
buf BUF1 (N2738, N2728);
and AND2 (N2739, N2729, N2351);
nand NAND2 (N2740, N2739, N2607);
buf BUF1 (N2741, N2722);
not NOT1 (N2742, N2726);
not NOT1 (N2743, N2742);
and AND3 (N2744, N2741, N298, N1335);
xor XOR2 (N2745, N2740, N2184);
and AND2 (N2746, N2737, N613);
xor XOR2 (N2747, N2744, N2365);
not NOT1 (N2748, N2746);
buf BUF1 (N2749, N2732);
buf BUF1 (N2750, N2733);
nand NAND4 (N2751, N2738, N2486, N1460, N164);
nor NOR3 (N2752, N2745, N646, N53);
or OR2 (N2753, N2736, N281);
and AND4 (N2754, N2751, N1372, N2616, N934);
nor NOR4 (N2755, N2748, N1977, N150, N2584);
nor NOR2 (N2756, N2750, N1237);
nor NOR4 (N2757, N2756, N2130, N2602, N1562);
and AND3 (N2758, N2757, N1825, N848);
buf BUF1 (N2759, N2754);
xor XOR2 (N2760, N2753, N1076);
nand NAND2 (N2761, N2759, N184);
xor XOR2 (N2762, N2743, N1234);
nor NOR2 (N2763, N2717, N2550);
nand NAND4 (N2764, N2762, N2543, N1963, N445);
xor XOR2 (N2765, N2761, N1095);
xor XOR2 (N2766, N2764, N1953);
buf BUF1 (N2767, N2734);
or OR4 (N2768, N2758, N1627, N1072, N1005);
buf BUF1 (N2769, N2752);
xor XOR2 (N2770, N2766, N2221);
and AND4 (N2771, N2763, N288, N2288, N2047);
not NOT1 (N2772, N2749);
nand NAND3 (N2773, N2755, N395, N2687);
nor NOR4 (N2774, N2769, N2588, N351, N2307);
nor NOR2 (N2775, N2771, N38);
nor NOR2 (N2776, N2774, N1562);
buf BUF1 (N2777, N2773);
not NOT1 (N2778, N2776);
or OR3 (N2779, N2775, N1328, N1691);
not NOT1 (N2780, N2770);
not NOT1 (N2781, N2765);
buf BUF1 (N2782, N2760);
nand NAND4 (N2783, N2781, N2503, N282, N2103);
or OR2 (N2784, N2768, N37);
not NOT1 (N2785, N2780);
not NOT1 (N2786, N2772);
or OR3 (N2787, N2778, N1025, N2607);
or OR2 (N2788, N2777, N2051);
buf BUF1 (N2789, N2779);
and AND2 (N2790, N2784, N918);
nand NAND3 (N2791, N2783, N772, N684);
buf BUF1 (N2792, N2767);
buf BUF1 (N2793, N2785);
nor NOR3 (N2794, N2788, N263, N395);
nor NOR3 (N2795, N2782, N1670, N2733);
and AND3 (N2796, N2786, N1540, N58);
buf BUF1 (N2797, N2793);
and AND4 (N2798, N2787, N978, N2479, N98);
xor XOR2 (N2799, N2796, N1912);
and AND2 (N2800, N2747, N2298);
nor NOR3 (N2801, N2797, N2261, N2288);
and AND3 (N2802, N2790, N2686, N1023);
not NOT1 (N2803, N2789);
or OR2 (N2804, N2799, N151);
and AND4 (N2805, N2791, N1835, N1305, N1981);
nor NOR4 (N2806, N2804, N2505, N2341, N854);
xor XOR2 (N2807, N2800, N241);
xor XOR2 (N2808, N2798, N2180);
buf BUF1 (N2809, N2803);
nand NAND4 (N2810, N2795, N1451, N2798, N2318);
or OR3 (N2811, N2809, N2047, N1294);
nand NAND2 (N2812, N2810, N1345);
or OR4 (N2813, N2802, N2728, N336, N1789);
xor XOR2 (N2814, N2805, N2422);
nor NOR2 (N2815, N2812, N2093);
or OR2 (N2816, N2792, N1951);
or OR4 (N2817, N2806, N566, N422, N1720);
nor NOR4 (N2818, N2813, N1416, N2604, N1075);
buf BUF1 (N2819, N2811);
not NOT1 (N2820, N2794);
buf BUF1 (N2821, N2818);
nor NOR4 (N2822, N2815, N943, N256, N178);
or OR3 (N2823, N2814, N2314, N1715);
not NOT1 (N2824, N2819);
buf BUF1 (N2825, N2821);
or OR2 (N2826, N2822, N1669);
buf BUF1 (N2827, N2825);
and AND3 (N2828, N2808, N1992, N2615);
xor XOR2 (N2829, N2824, N69);
and AND4 (N2830, N2826, N1211, N2685, N506);
nand NAND2 (N2831, N2830, N2598);
or OR2 (N2832, N2801, N2262);
and AND3 (N2833, N2816, N592, N455);
buf BUF1 (N2834, N2833);
xor XOR2 (N2835, N2834, N1295);
xor XOR2 (N2836, N2807, N1170);
nand NAND3 (N2837, N2827, N2096, N2538);
or OR4 (N2838, N2837, N2537, N2386, N460);
not NOT1 (N2839, N2832);
xor XOR2 (N2840, N2820, N1237);
nor NOR3 (N2841, N2829, N1167, N811);
buf BUF1 (N2842, N2835);
and AND2 (N2843, N2838, N2608);
not NOT1 (N2844, N2840);
buf BUF1 (N2845, N2841);
not NOT1 (N2846, N2844);
buf BUF1 (N2847, N2836);
and AND3 (N2848, N2823, N2324, N2360);
buf BUF1 (N2849, N2839);
nor NOR3 (N2850, N2848, N700, N1189);
xor XOR2 (N2851, N2846, N29);
not NOT1 (N2852, N2847);
nor NOR4 (N2853, N2828, N1482, N517, N428);
buf BUF1 (N2854, N2852);
and AND2 (N2855, N2853, N2699);
nand NAND2 (N2856, N2842, N402);
nand NAND2 (N2857, N2849, N1043);
xor XOR2 (N2858, N2845, N1914);
xor XOR2 (N2859, N2858, N2496);
nand NAND2 (N2860, N2856, N2270);
xor XOR2 (N2861, N2855, N663);
xor XOR2 (N2862, N2854, N2525);
nand NAND2 (N2863, N2850, N423);
nor NOR4 (N2864, N2861, N476, N2711, N746);
or OR3 (N2865, N2857, N2160, N791);
buf BUF1 (N2866, N2860);
nand NAND2 (N2867, N2843, N825);
nand NAND3 (N2868, N2817, N2068, N9);
nor NOR3 (N2869, N2863, N2643, N2632);
buf BUF1 (N2870, N2851);
not NOT1 (N2871, N2864);
not NOT1 (N2872, N2866);
not NOT1 (N2873, N2831);
nor NOR3 (N2874, N2871, N2605, N2097);
xor XOR2 (N2875, N2865, N2676);
not NOT1 (N2876, N2872);
xor XOR2 (N2877, N2862, N2178);
and AND4 (N2878, N2870, N2754, N2786, N2248);
or OR3 (N2879, N2873, N1767, N2020);
and AND3 (N2880, N2869, N101, N2831);
or OR2 (N2881, N2880, N2228);
nand NAND4 (N2882, N2876, N1810, N4, N1982);
or OR4 (N2883, N2879, N2460, N1029, N2703);
nand NAND4 (N2884, N2878, N1368, N170, N2642);
or OR2 (N2885, N2874, N572);
nor NOR4 (N2886, N2882, N2832, N2620, N2574);
xor XOR2 (N2887, N2881, N1288);
not NOT1 (N2888, N2886);
buf BUF1 (N2889, N2885);
nor NOR2 (N2890, N2867, N1376);
xor XOR2 (N2891, N2868, N1248);
nand NAND3 (N2892, N2877, N38, N1597);
nand NAND3 (N2893, N2875, N281, N422);
nor NOR4 (N2894, N2890, N831, N1138, N2036);
xor XOR2 (N2895, N2892, N1166);
not NOT1 (N2896, N2884);
not NOT1 (N2897, N2859);
nor NOR4 (N2898, N2895, N402, N1317, N1937);
nor NOR3 (N2899, N2896, N2823, N847);
xor XOR2 (N2900, N2897, N2507);
not NOT1 (N2901, N2887);
buf BUF1 (N2902, N2891);
buf BUF1 (N2903, N2888);
or OR2 (N2904, N2893, N1789);
or OR3 (N2905, N2894, N1818, N1034);
nor NOR2 (N2906, N2901, N2621);
or OR4 (N2907, N2906, N2900, N1919, N115);
nand NAND3 (N2908, N2440, N1328, N1301);
or OR3 (N2909, N2883, N2342, N2731);
not NOT1 (N2910, N2905);
or OR4 (N2911, N2904, N2783, N428, N165);
xor XOR2 (N2912, N2907, N589);
xor XOR2 (N2913, N2909, N1541);
buf BUF1 (N2914, N2899);
and AND2 (N2915, N2889, N861);
xor XOR2 (N2916, N2902, N1397);
buf BUF1 (N2917, N2916);
not NOT1 (N2918, N2912);
not NOT1 (N2919, N2908);
xor XOR2 (N2920, N2910, N1780);
and AND2 (N2921, N2911, N2776);
buf BUF1 (N2922, N2914);
buf BUF1 (N2923, N2903);
or OR3 (N2924, N2898, N1484, N2276);
not NOT1 (N2925, N2920);
or OR2 (N2926, N2913, N2755);
not NOT1 (N2927, N2924);
and AND2 (N2928, N2921, N494);
and AND4 (N2929, N2918, N2702, N2420, N2255);
xor XOR2 (N2930, N2925, N1167);
not NOT1 (N2931, N2917);
and AND4 (N2932, N2929, N828, N2398, N2754);
and AND2 (N2933, N2931, N652);
xor XOR2 (N2934, N2933, N2090);
and AND3 (N2935, N2927, N2084, N2736);
xor XOR2 (N2936, N2928, N1323);
xor XOR2 (N2937, N2919, N2358);
xor XOR2 (N2938, N2915, N753);
buf BUF1 (N2939, N2935);
nor NOR3 (N2940, N2938, N2241, N2167);
or OR3 (N2941, N2926, N1721, N1031);
buf BUF1 (N2942, N2939);
or OR4 (N2943, N2940, N109, N2383, N2109);
buf BUF1 (N2944, N2923);
and AND3 (N2945, N2934, N2865, N314);
nand NAND2 (N2946, N2944, N1943);
xor XOR2 (N2947, N2930, N1844);
buf BUF1 (N2948, N2932);
nand NAND4 (N2949, N2948, N2735, N2046, N439);
and AND3 (N2950, N2947, N376, N2105);
and AND3 (N2951, N2936, N2356, N44);
buf BUF1 (N2952, N2945);
or OR2 (N2953, N2922, N1578);
not NOT1 (N2954, N2949);
or OR3 (N2955, N2946, N334, N2177);
xor XOR2 (N2956, N2943, N1295);
or OR2 (N2957, N2951, N827);
and AND4 (N2958, N2937, N700, N2752, N1802);
nor NOR2 (N2959, N2958, N1209);
xor XOR2 (N2960, N2950, N1372);
or OR4 (N2961, N2956, N771, N450, N2381);
nand NAND2 (N2962, N2960, N1065);
or OR3 (N2963, N2959, N691, N581);
or OR4 (N2964, N2961, N658, N586, N1975);
nand NAND2 (N2965, N2942, N1638);
not NOT1 (N2966, N2952);
nand NAND2 (N2967, N2954, N2667);
nor NOR4 (N2968, N2963, N2326, N1263, N2681);
nor NOR4 (N2969, N2964, N2627, N1590, N2192);
nand NAND3 (N2970, N2941, N2620, N2550);
nor NOR2 (N2971, N2967, N718);
not NOT1 (N2972, N2965);
nor NOR2 (N2973, N2962, N2604);
nor NOR3 (N2974, N2953, N98, N198);
or OR3 (N2975, N2969, N999, N103);
nor NOR4 (N2976, N2973, N1019, N253, N804);
xor XOR2 (N2977, N2970, N2285);
not NOT1 (N2978, N2974);
buf BUF1 (N2979, N2977);
xor XOR2 (N2980, N2971, N97);
xor XOR2 (N2981, N2968, N450);
or OR4 (N2982, N2980, N1310, N111, N785);
nor NOR2 (N2983, N2982, N2855);
nor NOR2 (N2984, N2978, N1584);
nand NAND2 (N2985, N2984, N243);
nor NOR4 (N2986, N2985, N2240, N1238, N2604);
xor XOR2 (N2987, N2955, N2827);
xor XOR2 (N2988, N2972, N394);
and AND2 (N2989, N2987, N1067);
nor NOR3 (N2990, N2988, N2054, N2193);
xor XOR2 (N2991, N2989, N1139);
buf BUF1 (N2992, N2983);
not NOT1 (N2993, N2976);
or OR2 (N2994, N2986, N2961);
not NOT1 (N2995, N2966);
nor NOR3 (N2996, N2957, N459, N2911);
or OR2 (N2997, N2994, N2214);
nand NAND2 (N2998, N2979, N1925);
not NOT1 (N2999, N2990);
not NOT1 (N3000, N2996);
not NOT1 (N3001, N2993);
xor XOR2 (N3002, N2981, N549);
buf BUF1 (N3003, N2997);
nand NAND4 (N3004, N2995, N2107, N1002, N814);
nand NAND2 (N3005, N2999, N1241);
xor XOR2 (N3006, N3005, N2516);
buf BUF1 (N3007, N3003);
or OR4 (N3008, N2998, N2341, N984, N282);
not NOT1 (N3009, N2975);
nand NAND3 (N3010, N3006, N1692, N482);
endmodule