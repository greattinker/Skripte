// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N1617,N1602,N1609,N1612,N1615,N1607,N1618,N1584,N1603,N1619;

not NOT1 (N20, N9);
not NOT1 (N21, N7);
buf BUF1 (N22, N21);
buf BUF1 (N23, N16);
buf BUF1 (N24, N18);
not NOT1 (N25, N7);
or OR2 (N26, N10, N16);
and AND4 (N27, N13, N26, N26, N16);
and AND4 (N28, N20, N9, N14, N3);
nor NOR4 (N29, N11, N24, N17, N2);
nand NAND4 (N30, N11, N28, N25, N19);
nand NAND4 (N31, N12, N22, N13, N3);
nor NOR4 (N32, N16, N4, N6, N22);
nand NAND2 (N33, N25, N9);
not NOT1 (N34, N24);
not NOT1 (N35, N30);
nand NAND4 (N36, N25, N10, N6, N27);
buf BUF1 (N37, N25);
not NOT1 (N38, N33);
xor XOR2 (N39, N24, N5);
buf BUF1 (N40, N23);
nor NOR2 (N41, N31, N6);
or OR3 (N42, N37, N27, N4);
nand NAND3 (N43, N42, N15, N35);
nand NAND3 (N44, N40, N3, N16);
nor NOR4 (N45, N24, N15, N37, N38);
xor XOR2 (N46, N4, N37);
buf BUF1 (N47, N32);
and AND4 (N48, N45, N9, N23, N10);
buf BUF1 (N49, N43);
and AND2 (N50, N36, N2);
nand NAND4 (N51, N44, N11, N15, N43);
nor NOR3 (N52, N50, N16, N24);
buf BUF1 (N53, N52);
nand NAND2 (N54, N48, N23);
xor XOR2 (N55, N49, N35);
nor NOR3 (N56, N55, N40, N5);
xor XOR2 (N57, N54, N29);
not NOT1 (N58, N49);
not NOT1 (N59, N46);
nor NOR2 (N60, N39, N13);
nor NOR4 (N61, N51, N33, N35, N19);
or OR4 (N62, N56, N43, N17, N37);
xor XOR2 (N63, N57, N13);
buf BUF1 (N64, N60);
not NOT1 (N65, N41);
or OR2 (N66, N62, N40);
not NOT1 (N67, N59);
nand NAND2 (N68, N63, N48);
and AND3 (N69, N65, N7, N53);
not NOT1 (N70, N19);
buf BUF1 (N71, N61);
xor XOR2 (N72, N69, N57);
buf BUF1 (N73, N67);
nand NAND4 (N74, N64, N15, N65, N58);
and AND3 (N75, N40, N43, N12);
nor NOR2 (N76, N71, N20);
not NOT1 (N77, N34);
xor XOR2 (N78, N77, N18);
and AND2 (N79, N66, N14);
not NOT1 (N80, N75);
and AND4 (N81, N79, N39, N74, N15);
nor NOR3 (N82, N5, N3, N20);
nand NAND4 (N83, N72, N68, N64, N33);
nor NOR2 (N84, N35, N3);
not NOT1 (N85, N76);
buf BUF1 (N86, N85);
not NOT1 (N87, N70);
or OR3 (N88, N84, N46, N45);
xor XOR2 (N89, N88, N52);
nand NAND4 (N90, N78, N71, N63, N2);
not NOT1 (N91, N90);
not NOT1 (N92, N86);
nand NAND2 (N93, N89, N50);
not NOT1 (N94, N80);
and AND4 (N95, N87, N8, N60, N92);
or OR2 (N96, N54, N14);
or OR2 (N97, N96, N92);
nand NAND3 (N98, N83, N53, N71);
and AND3 (N99, N93, N86, N28);
and AND4 (N100, N81, N60, N3, N78);
or OR4 (N101, N91, N65, N92, N24);
nand NAND2 (N102, N98, N94);
nor NOR3 (N103, N79, N54, N87);
and AND4 (N104, N95, N53, N91, N70);
and AND4 (N105, N100, N50, N8, N46);
nand NAND4 (N106, N73, N58, N51, N43);
and AND2 (N107, N106, N17);
or OR3 (N108, N97, N46, N50);
and AND2 (N109, N107, N13);
and AND4 (N110, N104, N60, N107, N64);
nor NOR4 (N111, N102, N74, N15, N110);
nand NAND4 (N112, N23, N45, N100, N82);
nand NAND2 (N113, N7, N8);
nand NAND4 (N114, N105, N76, N58, N106);
not NOT1 (N115, N112);
buf BUF1 (N116, N101);
xor XOR2 (N117, N113, N29);
nand NAND2 (N118, N108, N50);
and AND2 (N119, N116, N63);
nand NAND2 (N120, N115, N13);
or OR2 (N121, N111, N46);
buf BUF1 (N122, N109);
nand NAND3 (N123, N47, N31, N35);
buf BUF1 (N124, N99);
xor XOR2 (N125, N123, N96);
buf BUF1 (N126, N125);
buf BUF1 (N127, N126);
buf BUF1 (N128, N121);
buf BUF1 (N129, N119);
xor XOR2 (N130, N128, N58);
and AND2 (N131, N103, N74);
and AND4 (N132, N118, N84, N36, N85);
and AND3 (N133, N131, N30, N67);
xor XOR2 (N134, N124, N84);
buf BUF1 (N135, N134);
buf BUF1 (N136, N120);
buf BUF1 (N137, N127);
xor XOR2 (N138, N129, N4);
xor XOR2 (N139, N137, N121);
not NOT1 (N140, N133);
xor XOR2 (N141, N135, N52);
or OR2 (N142, N139, N1);
not NOT1 (N143, N141);
or OR4 (N144, N138, N59, N33, N19);
xor XOR2 (N145, N142, N20);
xor XOR2 (N146, N122, N27);
xor XOR2 (N147, N140, N65);
xor XOR2 (N148, N136, N55);
buf BUF1 (N149, N148);
nand NAND3 (N150, N130, N3, N10);
xor XOR2 (N151, N143, N44);
xor XOR2 (N152, N132, N124);
not NOT1 (N153, N149);
nor NOR2 (N154, N153, N112);
not NOT1 (N155, N150);
or OR2 (N156, N151, N2);
and AND3 (N157, N154, N49, N78);
not NOT1 (N158, N157);
xor XOR2 (N159, N145, N145);
xor XOR2 (N160, N152, N52);
buf BUF1 (N161, N160);
xor XOR2 (N162, N159, N154);
or OR4 (N163, N146, N100, N58, N161);
xor XOR2 (N164, N112, N128);
nor NOR4 (N165, N163, N150, N53, N15);
or OR3 (N166, N117, N70, N45);
and AND4 (N167, N156, N151, N163, N55);
and AND2 (N168, N166, N11);
nand NAND3 (N169, N114, N126, N63);
buf BUF1 (N170, N155);
or OR3 (N171, N167, N139, N59);
not NOT1 (N172, N147);
nor NOR3 (N173, N158, N116, N56);
nor NOR3 (N174, N170, N13, N20);
and AND4 (N175, N169, N96, N5, N95);
nor NOR4 (N176, N172, N122, N151, N102);
nor NOR2 (N177, N175, N71);
not NOT1 (N178, N162);
not NOT1 (N179, N144);
nand NAND2 (N180, N176, N91);
nor NOR2 (N181, N178, N27);
not NOT1 (N182, N174);
or OR4 (N183, N179, N49, N151, N129);
and AND2 (N184, N164, N125);
not NOT1 (N185, N173);
buf BUF1 (N186, N168);
and AND2 (N187, N184, N166);
nand NAND2 (N188, N182, N41);
nand NAND3 (N189, N187, N100, N131);
or OR4 (N190, N181, N119, N57, N70);
buf BUF1 (N191, N186);
nor NOR3 (N192, N191, N113, N79);
xor XOR2 (N193, N192, N152);
nand NAND2 (N194, N183, N137);
not NOT1 (N195, N194);
nand NAND2 (N196, N189, N111);
not NOT1 (N197, N180);
not NOT1 (N198, N165);
not NOT1 (N199, N197);
nand NAND4 (N200, N190, N174, N22, N124);
nor NOR3 (N201, N195, N184, N156);
buf BUF1 (N202, N200);
not NOT1 (N203, N185);
nor NOR2 (N204, N201, N107);
nand NAND2 (N205, N171, N19);
buf BUF1 (N206, N205);
xor XOR2 (N207, N196, N65);
nor NOR2 (N208, N177, N85);
not NOT1 (N209, N193);
nand NAND4 (N210, N207, N96, N173, N163);
xor XOR2 (N211, N188, N71);
nor NOR3 (N212, N199, N92, N56);
not NOT1 (N213, N202);
nand NAND4 (N214, N198, N87, N51, N18);
and AND2 (N215, N212, N159);
buf BUF1 (N216, N204);
not NOT1 (N217, N210);
and AND2 (N218, N211, N123);
and AND2 (N219, N206, N35);
not NOT1 (N220, N203);
nor NOR3 (N221, N216, N111, N40);
xor XOR2 (N222, N213, N161);
or OR2 (N223, N215, N174);
xor XOR2 (N224, N218, N22);
nor NOR2 (N225, N217, N155);
nand NAND2 (N226, N221, N211);
nand NAND3 (N227, N225, N26, N60);
xor XOR2 (N228, N223, N78);
buf BUF1 (N229, N226);
buf BUF1 (N230, N208);
nor NOR3 (N231, N228, N50, N68);
or OR3 (N232, N214, N170, N130);
nand NAND4 (N233, N231, N79, N205, N188);
nand NAND2 (N234, N227, N222);
and AND3 (N235, N153, N40, N106);
nand NAND3 (N236, N232, N158, N73);
nor NOR3 (N237, N234, N181, N200);
buf BUF1 (N238, N235);
not NOT1 (N239, N219);
or OR3 (N240, N237, N107, N36);
and AND3 (N241, N220, N25, N99);
xor XOR2 (N242, N240, N52);
not NOT1 (N243, N233);
nor NOR2 (N244, N209, N49);
buf BUF1 (N245, N230);
nor NOR3 (N246, N243, N107, N185);
and AND3 (N247, N242, N5, N136);
and AND2 (N248, N238, N109);
nor NOR4 (N249, N248, N49, N201, N114);
and AND2 (N250, N247, N33);
xor XOR2 (N251, N224, N250);
xor XOR2 (N252, N38, N10);
buf BUF1 (N253, N236);
nor NOR4 (N254, N246, N38, N169, N104);
xor XOR2 (N255, N245, N249);
or OR4 (N256, N158, N209, N33, N42);
buf BUF1 (N257, N251);
nor NOR3 (N258, N229, N89, N59);
not NOT1 (N259, N255);
or OR3 (N260, N256, N112, N184);
not NOT1 (N261, N260);
and AND4 (N262, N239, N192, N69, N65);
nor NOR3 (N263, N258, N76, N161);
buf BUF1 (N264, N254);
not NOT1 (N265, N257);
nor NOR4 (N266, N261, N6, N68, N122);
not NOT1 (N267, N264);
not NOT1 (N268, N244);
and AND2 (N269, N267, N206);
buf BUF1 (N270, N252);
not NOT1 (N271, N241);
buf BUF1 (N272, N262);
nand NAND3 (N273, N268, N153, N227);
not NOT1 (N274, N272);
buf BUF1 (N275, N270);
or OR2 (N276, N266, N67);
and AND3 (N277, N276, N264, N170);
and AND2 (N278, N275, N83);
nor NOR2 (N279, N277, N99);
nor NOR4 (N280, N273, N102, N8, N189);
not NOT1 (N281, N280);
and AND2 (N282, N253, N133);
xor XOR2 (N283, N265, N218);
and AND2 (N284, N274, N247);
nand NAND3 (N285, N284, N68, N269);
or OR3 (N286, N77, N142, N44);
xor XOR2 (N287, N279, N126);
and AND4 (N288, N283, N222, N9, N70);
xor XOR2 (N289, N282, N45);
and AND2 (N290, N278, N279);
and AND2 (N291, N288, N184);
nor NOR4 (N292, N263, N40, N96, N105);
nor NOR4 (N293, N259, N3, N31, N36);
xor XOR2 (N294, N287, N160);
nor NOR3 (N295, N289, N198, N173);
nor NOR2 (N296, N293, N292);
nand NAND2 (N297, N8, N34);
nor NOR4 (N298, N285, N53, N255, N149);
xor XOR2 (N299, N286, N60);
and AND2 (N300, N296, N145);
xor XOR2 (N301, N298, N29);
buf BUF1 (N302, N281);
nand NAND4 (N303, N291, N281, N212, N175);
nor NOR4 (N304, N290, N141, N129, N131);
and AND4 (N305, N302, N59, N249, N143);
not NOT1 (N306, N294);
and AND2 (N307, N303, N110);
nand NAND3 (N308, N271, N160, N239);
or OR4 (N309, N305, N134, N300, N106);
nand NAND2 (N310, N136, N201);
buf BUF1 (N311, N304);
not NOT1 (N312, N311);
nor NOR4 (N313, N309, N244, N15, N72);
not NOT1 (N314, N297);
or OR2 (N315, N299, N7);
buf BUF1 (N316, N295);
buf BUF1 (N317, N314);
or OR4 (N318, N317, N160, N191, N55);
buf BUF1 (N319, N307);
and AND3 (N320, N310, N297, N271);
and AND3 (N321, N320, N229, N197);
buf BUF1 (N322, N316);
nor NOR2 (N323, N318, N41);
or OR3 (N324, N319, N303, N243);
and AND2 (N325, N301, N256);
nor NOR4 (N326, N312, N106, N39, N322);
and AND2 (N327, N284, N302);
or OR3 (N328, N326, N273, N221);
not NOT1 (N329, N308);
buf BUF1 (N330, N306);
or OR4 (N331, N325, N189, N249, N264);
or OR3 (N332, N315, N330, N78);
nand NAND2 (N333, N293, N132);
nor NOR2 (N334, N324, N249);
not NOT1 (N335, N327);
not NOT1 (N336, N331);
and AND3 (N337, N335, N253, N238);
nand NAND2 (N338, N329, N70);
not NOT1 (N339, N333);
and AND3 (N340, N332, N338, N262);
xor XOR2 (N341, N216, N320);
or OR3 (N342, N323, N178, N230);
buf BUF1 (N343, N340);
nor NOR2 (N344, N341, N174);
xor XOR2 (N345, N328, N313);
nor NOR3 (N346, N39, N258, N264);
xor XOR2 (N347, N337, N274);
and AND3 (N348, N321, N270, N273);
nor NOR2 (N349, N346, N269);
xor XOR2 (N350, N344, N151);
and AND2 (N351, N343, N217);
nand NAND3 (N352, N351, N41, N136);
nor NOR4 (N353, N350, N8, N322, N309);
or OR3 (N354, N336, N130, N25);
xor XOR2 (N355, N352, N305);
and AND4 (N356, N339, N56, N116, N19);
not NOT1 (N357, N354);
buf BUF1 (N358, N348);
xor XOR2 (N359, N358, N342);
nor NOR4 (N360, N330, N154, N122, N73);
xor XOR2 (N361, N357, N290);
buf BUF1 (N362, N349);
buf BUF1 (N363, N345);
not NOT1 (N364, N353);
nand NAND4 (N365, N363, N269, N127, N35);
buf BUF1 (N366, N362);
xor XOR2 (N367, N356, N157);
xor XOR2 (N368, N364, N189);
and AND3 (N369, N334, N315, N54);
buf BUF1 (N370, N369);
xor XOR2 (N371, N360, N127);
nor NOR3 (N372, N370, N26, N353);
buf BUF1 (N373, N355);
and AND4 (N374, N347, N103, N173, N74);
or OR2 (N375, N374, N236);
and AND4 (N376, N375, N59, N280, N360);
or OR4 (N377, N367, N358, N339, N37);
buf BUF1 (N378, N376);
nor NOR4 (N379, N366, N110, N151, N209);
or OR3 (N380, N371, N106, N356);
and AND2 (N381, N372, N285);
or OR3 (N382, N365, N141, N187);
xor XOR2 (N383, N382, N251);
not NOT1 (N384, N379);
or OR4 (N385, N380, N288, N229, N112);
or OR4 (N386, N385, N307, N87, N247);
or OR3 (N387, N381, N280, N172);
nor NOR2 (N388, N368, N61);
and AND3 (N389, N388, N31, N93);
buf BUF1 (N390, N373);
xor XOR2 (N391, N359, N237);
nand NAND4 (N392, N386, N105, N378, N226);
not NOT1 (N393, N144);
buf BUF1 (N394, N390);
xor XOR2 (N395, N391, N195);
xor XOR2 (N396, N392, N37);
xor XOR2 (N397, N389, N391);
nor NOR3 (N398, N397, N238, N157);
buf BUF1 (N399, N393);
buf BUF1 (N400, N395);
nor NOR2 (N401, N394, N129);
nor NOR4 (N402, N387, N275, N131, N320);
and AND4 (N403, N384, N285, N337, N358);
xor XOR2 (N404, N361, N272);
and AND2 (N405, N396, N190);
or OR3 (N406, N398, N344, N1);
or OR4 (N407, N383, N406, N139, N387);
not NOT1 (N408, N233);
and AND4 (N409, N408, N199, N136, N336);
buf BUF1 (N410, N400);
or OR4 (N411, N405, N6, N385, N369);
or OR3 (N412, N377, N84, N56);
nor NOR2 (N413, N401, N140);
buf BUF1 (N414, N407);
not NOT1 (N415, N413);
not NOT1 (N416, N410);
and AND2 (N417, N399, N320);
nand NAND4 (N418, N409, N326, N322, N67);
not NOT1 (N419, N412);
buf BUF1 (N420, N415);
and AND2 (N421, N418, N17);
not NOT1 (N422, N419);
nand NAND3 (N423, N417, N189, N341);
nor NOR2 (N424, N423, N322);
buf BUF1 (N425, N420);
buf BUF1 (N426, N424);
or OR3 (N427, N416, N97, N106);
not NOT1 (N428, N402);
nor NOR2 (N429, N422, N262);
and AND3 (N430, N421, N382, N408);
nand NAND4 (N431, N426, N347, N54, N164);
or OR3 (N432, N427, N51, N126);
nor NOR4 (N433, N425, N417, N101, N327);
nor NOR2 (N434, N414, N71);
xor XOR2 (N435, N434, N219);
and AND4 (N436, N411, N151, N359, N233);
or OR2 (N437, N431, N171);
or OR3 (N438, N435, N313, N342);
xor XOR2 (N439, N403, N32);
buf BUF1 (N440, N433);
xor XOR2 (N441, N432, N428);
nand NAND2 (N442, N79, N6);
nor NOR4 (N443, N436, N272, N242, N406);
and AND3 (N444, N439, N181, N156);
nor NOR3 (N445, N430, N5, N103);
buf BUF1 (N446, N443);
and AND3 (N447, N444, N217, N41);
not NOT1 (N448, N440);
xor XOR2 (N449, N446, N186);
nand NAND4 (N450, N441, N212, N98, N331);
nand NAND2 (N451, N429, N187);
and AND4 (N452, N448, N299, N132, N348);
buf BUF1 (N453, N452);
or OR4 (N454, N404, N3, N263, N305);
nand NAND2 (N455, N447, N84);
nor NOR3 (N456, N449, N15, N318);
nor NOR2 (N457, N453, N24);
not NOT1 (N458, N451);
and AND2 (N459, N445, N364);
nor NOR2 (N460, N456, N338);
not NOT1 (N461, N455);
nand NAND4 (N462, N454, N325, N326, N104);
and AND3 (N463, N462, N323, N23);
or OR3 (N464, N457, N398, N53);
not NOT1 (N465, N442);
nand NAND4 (N466, N465, N386, N196, N440);
nor NOR3 (N467, N437, N290, N70);
or OR3 (N468, N450, N422, N148);
nor NOR2 (N469, N459, N99);
xor XOR2 (N470, N463, N23);
nand NAND3 (N471, N467, N414, N227);
not NOT1 (N472, N458);
not NOT1 (N473, N472);
not NOT1 (N474, N461);
nor NOR3 (N475, N466, N454, N439);
xor XOR2 (N476, N464, N416);
or OR4 (N477, N460, N350, N23, N439);
not NOT1 (N478, N473);
nor NOR4 (N479, N470, N191, N164, N171);
nand NAND3 (N480, N474, N65, N68);
buf BUF1 (N481, N468);
not NOT1 (N482, N476);
nand NAND4 (N483, N477, N98, N250, N12);
xor XOR2 (N484, N471, N420);
xor XOR2 (N485, N480, N94);
nor NOR2 (N486, N438, N23);
buf BUF1 (N487, N481);
xor XOR2 (N488, N483, N423);
nand NAND4 (N489, N487, N279, N200, N292);
and AND4 (N490, N482, N118, N390, N217);
nand NAND4 (N491, N484, N35, N400, N131);
and AND2 (N492, N488, N221);
nand NAND3 (N493, N489, N400, N77);
and AND3 (N494, N485, N390, N172);
and AND3 (N495, N478, N419, N25);
and AND4 (N496, N469, N27, N232, N16);
and AND3 (N497, N492, N33, N428);
xor XOR2 (N498, N491, N437);
nor NOR3 (N499, N495, N163, N333);
buf BUF1 (N500, N494);
buf BUF1 (N501, N500);
xor XOR2 (N502, N496, N135);
or OR3 (N503, N499, N432, N408);
xor XOR2 (N504, N498, N458);
not NOT1 (N505, N497);
xor XOR2 (N506, N502, N282);
nand NAND2 (N507, N493, N454);
and AND4 (N508, N507, N75, N87, N428);
or OR2 (N509, N501, N127);
not NOT1 (N510, N509);
nor NOR4 (N511, N508, N303, N17, N49);
or OR4 (N512, N490, N293, N306, N265);
nand NAND2 (N513, N510, N45);
not NOT1 (N514, N512);
and AND3 (N515, N511, N173, N212);
nand NAND3 (N516, N503, N402, N225);
and AND2 (N517, N516, N395);
or OR3 (N518, N513, N472, N94);
and AND3 (N519, N506, N359, N206);
and AND4 (N520, N514, N62, N72, N40);
not NOT1 (N521, N519);
buf BUF1 (N522, N486);
nand NAND3 (N523, N479, N163, N94);
buf BUF1 (N524, N504);
nor NOR2 (N525, N524, N292);
or OR4 (N526, N523, N4, N521, N241);
xor XOR2 (N527, N384, N470);
or OR3 (N528, N522, N380, N526);
buf BUF1 (N529, N115);
nor NOR4 (N530, N520, N74, N42, N262);
xor XOR2 (N531, N525, N463);
nand NAND3 (N532, N475, N230, N525);
nand NAND3 (N533, N529, N271, N243);
or OR3 (N534, N527, N178, N415);
nand NAND3 (N535, N532, N128, N160);
nor NOR3 (N536, N535, N419, N506);
and AND4 (N537, N528, N185, N215, N253);
nor NOR4 (N538, N530, N506, N46, N319);
nor NOR3 (N539, N537, N533, N112);
not NOT1 (N540, N269);
xor XOR2 (N541, N540, N514);
and AND3 (N542, N515, N199, N88);
not NOT1 (N543, N538);
nor NOR2 (N544, N542, N482);
nor NOR4 (N545, N544, N375, N352, N147);
and AND4 (N546, N534, N279, N217, N141);
or OR2 (N547, N539, N141);
and AND4 (N548, N545, N73, N140, N356);
and AND2 (N549, N543, N348);
or OR4 (N550, N505, N235, N367, N195);
nand NAND3 (N551, N549, N349, N391);
or OR2 (N552, N536, N124);
or OR3 (N553, N518, N220, N480);
xor XOR2 (N554, N517, N12);
not NOT1 (N555, N546);
not NOT1 (N556, N554);
not NOT1 (N557, N552);
buf BUF1 (N558, N541);
nor NOR4 (N559, N551, N380, N291, N62);
nor NOR3 (N560, N548, N425, N56);
buf BUF1 (N561, N556);
and AND4 (N562, N559, N172, N57, N305);
nor NOR3 (N563, N562, N8, N476);
buf BUF1 (N564, N531);
nand NAND4 (N565, N553, N507, N73, N12);
nor NOR2 (N566, N565, N523);
nand NAND4 (N567, N547, N306, N341, N555);
buf BUF1 (N568, N552);
or OR4 (N569, N566, N340, N365, N391);
or OR2 (N570, N568, N233);
buf BUF1 (N571, N550);
or OR3 (N572, N569, N37, N232);
and AND3 (N573, N571, N299, N24);
nand NAND4 (N574, N570, N434, N233, N329);
nor NOR2 (N575, N573, N333);
xor XOR2 (N576, N567, N360);
and AND2 (N577, N558, N496);
buf BUF1 (N578, N574);
buf BUF1 (N579, N578);
nand NAND2 (N580, N564, N176);
buf BUF1 (N581, N561);
nand NAND3 (N582, N581, N249, N275);
and AND3 (N583, N563, N564, N307);
nor NOR2 (N584, N572, N544);
not NOT1 (N585, N583);
or OR4 (N586, N580, N54, N317, N113);
xor XOR2 (N587, N584, N12);
nor NOR3 (N588, N560, N551, N221);
nor NOR4 (N589, N585, N107, N437, N582);
nand NAND4 (N590, N586, N557, N118, N57);
buf BUF1 (N591, N5);
buf BUF1 (N592, N13);
nor NOR3 (N593, N587, N14, N361);
buf BUF1 (N594, N591);
or OR4 (N595, N588, N544, N379, N92);
not NOT1 (N596, N577);
or OR3 (N597, N592, N42, N203);
xor XOR2 (N598, N593, N262);
and AND2 (N599, N576, N394);
nor NOR3 (N600, N575, N94, N47);
or OR3 (N601, N594, N553, N429);
nor NOR2 (N602, N589, N234);
nand NAND2 (N603, N598, N4);
not NOT1 (N604, N600);
or OR2 (N605, N602, N143);
xor XOR2 (N606, N605, N398);
and AND4 (N607, N601, N342, N273, N250);
or OR2 (N608, N606, N225);
xor XOR2 (N609, N608, N343);
not NOT1 (N610, N599);
not NOT1 (N611, N607);
xor XOR2 (N612, N596, N240);
xor XOR2 (N613, N590, N478);
buf BUF1 (N614, N603);
buf BUF1 (N615, N604);
xor XOR2 (N616, N610, N179);
xor XOR2 (N617, N616, N310);
xor XOR2 (N618, N609, N415);
or OR4 (N619, N614, N339, N564, N388);
and AND3 (N620, N611, N192, N108);
buf BUF1 (N621, N620);
buf BUF1 (N622, N618);
nor NOR3 (N623, N617, N356, N406);
buf BUF1 (N624, N615);
buf BUF1 (N625, N624);
nor NOR3 (N626, N612, N575, N36);
buf BUF1 (N627, N623);
nand NAND4 (N628, N579, N15, N497, N328);
and AND4 (N629, N622, N411, N179, N445);
and AND4 (N630, N628, N326, N65, N195);
not NOT1 (N631, N595);
not NOT1 (N632, N629);
not NOT1 (N633, N627);
nand NAND3 (N634, N625, N565, N345);
or OR4 (N635, N597, N52, N235, N34);
not NOT1 (N636, N634);
not NOT1 (N637, N630);
nand NAND3 (N638, N621, N63, N335);
nand NAND3 (N639, N638, N348, N276);
xor XOR2 (N640, N637, N390);
not NOT1 (N641, N619);
not NOT1 (N642, N640);
nor NOR2 (N643, N635, N147);
and AND3 (N644, N626, N107, N450);
or OR3 (N645, N632, N131, N425);
nand NAND2 (N646, N639, N121);
buf BUF1 (N647, N633);
xor XOR2 (N648, N641, N458);
nor NOR2 (N649, N648, N314);
buf BUF1 (N650, N636);
nand NAND4 (N651, N631, N297, N504, N390);
or OR3 (N652, N613, N302, N282);
nor NOR3 (N653, N643, N290, N418);
nor NOR2 (N654, N642, N485);
buf BUF1 (N655, N649);
or OR4 (N656, N650, N626, N104, N288);
buf BUF1 (N657, N645);
nor NOR2 (N658, N644, N2);
buf BUF1 (N659, N657);
nand NAND3 (N660, N653, N317, N298);
nand NAND4 (N661, N655, N286, N69, N113);
and AND3 (N662, N654, N160, N105);
nor NOR3 (N663, N652, N418, N363);
nor NOR2 (N664, N659, N113);
nand NAND2 (N665, N647, N215);
buf BUF1 (N666, N664);
buf BUF1 (N667, N656);
nor NOR4 (N668, N662, N309, N529, N531);
xor XOR2 (N669, N646, N613);
xor XOR2 (N670, N661, N305);
or OR4 (N671, N658, N637, N404, N15);
not NOT1 (N672, N651);
or OR2 (N673, N671, N478);
nand NAND3 (N674, N670, N631, N71);
nor NOR4 (N675, N665, N532, N250, N526);
nor NOR3 (N676, N666, N349, N9);
xor XOR2 (N677, N669, N429);
nor NOR2 (N678, N660, N359);
buf BUF1 (N679, N677);
nand NAND2 (N680, N678, N549);
nor NOR3 (N681, N673, N64, N57);
nand NAND2 (N682, N668, N418);
xor XOR2 (N683, N680, N209);
nand NAND2 (N684, N681, N495);
and AND4 (N685, N679, N315, N504, N175);
nor NOR2 (N686, N674, N225);
and AND3 (N687, N672, N537, N485);
not NOT1 (N688, N685);
nor NOR3 (N689, N676, N53, N365);
not NOT1 (N690, N688);
xor XOR2 (N691, N667, N544);
or OR3 (N692, N687, N110, N220);
and AND2 (N693, N684, N663);
nor NOR4 (N694, N413, N122, N139, N109);
nand NAND4 (N695, N689, N355, N139, N609);
or OR3 (N696, N694, N433, N22);
not NOT1 (N697, N682);
buf BUF1 (N698, N692);
not NOT1 (N699, N695);
not NOT1 (N700, N696);
and AND3 (N701, N693, N650, N654);
or OR3 (N702, N675, N97, N48);
and AND3 (N703, N699, N443, N72);
buf BUF1 (N704, N701);
buf BUF1 (N705, N698);
not NOT1 (N706, N704);
nor NOR3 (N707, N706, N212, N508);
or OR3 (N708, N707, N680, N529);
nand NAND2 (N709, N691, N683);
not NOT1 (N710, N617);
nor NOR2 (N711, N703, N139);
not NOT1 (N712, N690);
not NOT1 (N713, N700);
xor XOR2 (N714, N697, N616);
and AND2 (N715, N713, N131);
not NOT1 (N716, N709);
and AND3 (N717, N686, N161, N25);
and AND4 (N718, N717, N419, N615, N200);
nand NAND3 (N719, N711, N572, N248);
nor NOR2 (N720, N708, N12);
and AND2 (N721, N716, N644);
nand NAND2 (N722, N720, N378);
nor NOR2 (N723, N710, N446);
and AND2 (N724, N712, N23);
not NOT1 (N725, N723);
nand NAND4 (N726, N725, N690, N426, N129);
not NOT1 (N727, N719);
nand NAND3 (N728, N718, N277, N707);
nor NOR4 (N729, N705, N306, N612, N683);
nor NOR2 (N730, N727, N119);
nor NOR4 (N731, N726, N178, N43, N395);
or OR2 (N732, N715, N660);
nand NAND2 (N733, N724, N86);
not NOT1 (N734, N729);
nand NAND4 (N735, N702, N183, N198, N83);
and AND3 (N736, N734, N297, N272);
buf BUF1 (N737, N730);
not NOT1 (N738, N728);
not NOT1 (N739, N733);
xor XOR2 (N740, N731, N63);
nor NOR2 (N741, N735, N33);
and AND3 (N742, N714, N406, N6);
and AND4 (N743, N737, N265, N400, N426);
buf BUF1 (N744, N740);
nor NOR3 (N745, N739, N27, N528);
and AND2 (N746, N736, N197);
nand NAND3 (N747, N732, N495, N389);
nand NAND2 (N748, N745, N270);
nor NOR2 (N749, N721, N296);
nor NOR3 (N750, N747, N560, N25);
or OR4 (N751, N738, N241, N522, N90);
not NOT1 (N752, N741);
and AND2 (N753, N748, N521);
and AND3 (N754, N744, N477, N232);
and AND2 (N755, N751, N381);
buf BUF1 (N756, N749);
and AND2 (N757, N743, N529);
or OR4 (N758, N755, N320, N186, N463);
nor NOR4 (N759, N742, N225, N495, N708);
nand NAND2 (N760, N752, N577);
and AND4 (N761, N758, N636, N594, N746);
or OR3 (N762, N256, N606, N355);
not NOT1 (N763, N756);
nand NAND4 (N764, N754, N163, N44, N418);
xor XOR2 (N765, N759, N259);
and AND4 (N766, N761, N534, N620, N23);
xor XOR2 (N767, N762, N284);
or OR2 (N768, N766, N380);
xor XOR2 (N769, N765, N172);
or OR3 (N770, N750, N549, N720);
nand NAND4 (N771, N753, N602, N382, N639);
and AND2 (N772, N722, N533);
or OR3 (N773, N763, N562, N65);
nor NOR4 (N774, N760, N658, N235, N183);
nor NOR2 (N775, N774, N313);
not NOT1 (N776, N772);
not NOT1 (N777, N764);
and AND4 (N778, N776, N14, N6, N414);
nand NAND3 (N779, N757, N348, N703);
not NOT1 (N780, N770);
buf BUF1 (N781, N777);
and AND4 (N782, N780, N94, N197, N299);
not NOT1 (N783, N769);
and AND3 (N784, N778, N145, N398);
nand NAND3 (N785, N768, N424, N331);
buf BUF1 (N786, N784);
and AND2 (N787, N781, N591);
not NOT1 (N788, N767);
or OR2 (N789, N771, N33);
or OR4 (N790, N789, N372, N524, N440);
xor XOR2 (N791, N773, N234);
buf BUF1 (N792, N779);
not NOT1 (N793, N791);
not NOT1 (N794, N783);
nand NAND2 (N795, N787, N175);
nand NAND2 (N796, N795, N505);
and AND4 (N797, N785, N312, N516, N407);
not NOT1 (N798, N797);
buf BUF1 (N799, N782);
not NOT1 (N800, N796);
buf BUF1 (N801, N775);
nand NAND4 (N802, N788, N561, N425, N410);
nand NAND4 (N803, N794, N438, N761, N300);
nor NOR4 (N804, N799, N330, N277, N337);
nor NOR4 (N805, N801, N740, N115, N679);
buf BUF1 (N806, N792);
nand NAND2 (N807, N790, N337);
nor NOR3 (N808, N798, N506, N516);
or OR2 (N809, N807, N466);
nand NAND2 (N810, N800, N316);
and AND4 (N811, N810, N27, N185, N628);
or OR4 (N812, N809, N807, N362, N312);
buf BUF1 (N813, N793);
nor NOR2 (N814, N786, N746);
nand NAND3 (N815, N812, N77, N477);
not NOT1 (N816, N813);
nor NOR3 (N817, N814, N141, N144);
and AND2 (N818, N808, N256);
nand NAND4 (N819, N803, N808, N646, N284);
nor NOR3 (N820, N815, N180, N58);
not NOT1 (N821, N811);
not NOT1 (N822, N816);
nor NOR4 (N823, N817, N666, N584, N818);
not NOT1 (N824, N662);
buf BUF1 (N825, N823);
buf BUF1 (N826, N825);
xor XOR2 (N827, N824, N760);
nand NAND2 (N828, N822, N734);
buf BUF1 (N829, N804);
xor XOR2 (N830, N826, N580);
nor NOR2 (N831, N819, N360);
or OR3 (N832, N830, N79, N330);
xor XOR2 (N833, N805, N442);
or OR2 (N834, N821, N759);
buf BUF1 (N835, N827);
not NOT1 (N836, N828);
and AND4 (N837, N820, N440, N359, N426);
or OR3 (N838, N806, N209, N574);
and AND4 (N839, N802, N490, N759, N498);
buf BUF1 (N840, N829);
nand NAND3 (N841, N834, N317, N80);
or OR2 (N842, N841, N786);
nand NAND4 (N843, N838, N275, N446, N825);
nor NOR3 (N844, N831, N746, N386);
not NOT1 (N845, N839);
xor XOR2 (N846, N843, N730);
or OR2 (N847, N837, N588);
nand NAND4 (N848, N833, N1, N115, N371);
nand NAND3 (N849, N847, N716, N124);
nand NAND4 (N850, N835, N333, N840, N478);
nand NAND2 (N851, N50, N817);
and AND4 (N852, N845, N734, N53, N452);
or OR2 (N853, N832, N235);
and AND2 (N854, N844, N436);
nand NAND3 (N855, N850, N651, N632);
and AND2 (N856, N849, N174);
buf BUF1 (N857, N846);
nor NOR2 (N858, N857, N362);
buf BUF1 (N859, N852);
not NOT1 (N860, N836);
buf BUF1 (N861, N859);
nor NOR4 (N862, N848, N833, N169, N816);
not NOT1 (N863, N861);
xor XOR2 (N864, N860, N99);
nand NAND3 (N865, N853, N372, N758);
or OR2 (N866, N864, N344);
xor XOR2 (N867, N858, N721);
buf BUF1 (N868, N862);
and AND4 (N869, N856, N227, N397, N784);
nand NAND3 (N870, N854, N7, N14);
nand NAND2 (N871, N855, N603);
or OR3 (N872, N866, N279, N305);
nand NAND4 (N873, N851, N131, N327, N604);
or OR3 (N874, N842, N185, N500);
and AND3 (N875, N872, N655, N382);
buf BUF1 (N876, N865);
xor XOR2 (N877, N869, N492);
buf BUF1 (N878, N875);
buf BUF1 (N879, N871);
xor XOR2 (N880, N877, N878);
and AND4 (N881, N176, N345, N113, N166);
and AND2 (N882, N880, N502);
nor NOR2 (N883, N874, N681);
not NOT1 (N884, N873);
not NOT1 (N885, N870);
buf BUF1 (N886, N881);
xor XOR2 (N887, N879, N678);
buf BUF1 (N888, N868);
xor XOR2 (N889, N887, N827);
not NOT1 (N890, N883);
and AND3 (N891, N882, N777, N318);
and AND4 (N892, N867, N841, N484, N880);
buf BUF1 (N893, N891);
xor XOR2 (N894, N892, N676);
and AND2 (N895, N890, N521);
nor NOR4 (N896, N863, N482, N400, N585);
xor XOR2 (N897, N884, N176);
buf BUF1 (N898, N893);
xor XOR2 (N899, N889, N310);
or OR3 (N900, N886, N694, N221);
and AND3 (N901, N894, N879, N716);
not NOT1 (N902, N898);
or OR2 (N903, N901, N397);
xor XOR2 (N904, N885, N868);
nand NAND2 (N905, N896, N378);
nand NAND2 (N906, N900, N803);
nor NOR2 (N907, N899, N482);
and AND2 (N908, N876, N371);
nand NAND3 (N909, N903, N359, N274);
or OR2 (N910, N904, N88);
or OR3 (N911, N895, N273, N45);
or OR2 (N912, N906, N677);
buf BUF1 (N913, N909);
nor NOR3 (N914, N907, N848, N394);
buf BUF1 (N915, N911);
or OR3 (N916, N915, N610, N896);
xor XOR2 (N917, N902, N571);
nand NAND2 (N918, N914, N181);
xor XOR2 (N919, N916, N422);
nand NAND4 (N920, N905, N699, N829, N793);
and AND3 (N921, N917, N403, N584);
nor NOR2 (N922, N908, N619);
nand NAND2 (N923, N888, N457);
and AND2 (N924, N922, N5);
nand NAND2 (N925, N918, N881);
nand NAND4 (N926, N923, N925, N380, N712);
and AND4 (N927, N260, N258, N199, N807);
nand NAND4 (N928, N912, N21, N850, N888);
nor NOR2 (N929, N913, N510);
nor NOR4 (N930, N920, N830, N127, N166);
and AND2 (N931, N928, N111);
xor XOR2 (N932, N897, N470);
nor NOR2 (N933, N929, N794);
nand NAND2 (N934, N932, N796);
nand NAND4 (N935, N921, N627, N564, N21);
xor XOR2 (N936, N910, N54);
or OR4 (N937, N933, N63, N65, N595);
nor NOR2 (N938, N930, N867);
nand NAND4 (N939, N938, N434, N558, N733);
nand NAND2 (N940, N936, N864);
nor NOR2 (N941, N924, N899);
nand NAND2 (N942, N937, N213);
not NOT1 (N943, N927);
and AND2 (N944, N943, N177);
and AND3 (N945, N944, N271, N610);
nand NAND2 (N946, N940, N23);
xor XOR2 (N947, N945, N59);
not NOT1 (N948, N934);
xor XOR2 (N949, N947, N294);
xor XOR2 (N950, N941, N19);
nor NOR3 (N951, N942, N540, N547);
and AND3 (N952, N926, N896, N115);
xor XOR2 (N953, N950, N760);
not NOT1 (N954, N949);
xor XOR2 (N955, N952, N805);
not NOT1 (N956, N954);
buf BUF1 (N957, N931);
nand NAND2 (N958, N939, N671);
buf BUF1 (N959, N957);
nand NAND4 (N960, N959, N450, N955, N820);
and AND2 (N961, N372, N477);
xor XOR2 (N962, N961, N354);
nor NOR4 (N963, N956, N235, N186, N703);
buf BUF1 (N964, N935);
nor NOR4 (N965, N951, N845, N510, N803);
and AND3 (N966, N958, N860, N308);
or OR3 (N967, N948, N316, N507);
nand NAND3 (N968, N953, N35, N194);
or OR3 (N969, N968, N186, N364);
or OR4 (N970, N967, N714, N73, N182);
nand NAND2 (N971, N919, N183);
and AND4 (N972, N946, N885, N366, N293);
nor NOR2 (N973, N966, N828);
nor NOR3 (N974, N972, N424, N676);
nand NAND2 (N975, N974, N570);
xor XOR2 (N976, N960, N161);
xor XOR2 (N977, N963, N207);
buf BUF1 (N978, N965);
or OR3 (N979, N970, N691, N427);
or OR3 (N980, N978, N199, N65);
nand NAND2 (N981, N973, N629);
nand NAND4 (N982, N962, N736, N839, N6);
nor NOR2 (N983, N969, N146);
or OR4 (N984, N980, N911, N302, N225);
not NOT1 (N985, N981);
nand NAND2 (N986, N964, N190);
buf BUF1 (N987, N983);
nor NOR3 (N988, N986, N984, N103);
not NOT1 (N989, N396);
xor XOR2 (N990, N975, N138);
not NOT1 (N991, N971);
and AND2 (N992, N982, N68);
buf BUF1 (N993, N988);
nand NAND3 (N994, N979, N457, N157);
and AND3 (N995, N992, N94, N793);
xor XOR2 (N996, N995, N611);
xor XOR2 (N997, N990, N292);
and AND3 (N998, N994, N950, N164);
buf BUF1 (N999, N993);
or OR3 (N1000, N998, N762, N507);
and AND4 (N1001, N999, N170, N961, N610);
xor XOR2 (N1002, N996, N353);
and AND3 (N1003, N991, N633, N400);
and AND4 (N1004, N1000, N55, N222, N177);
or OR3 (N1005, N1002, N546, N659);
nand NAND3 (N1006, N977, N745, N282);
nand NAND2 (N1007, N1004, N205);
or OR2 (N1008, N976, N848);
buf BUF1 (N1009, N997);
xor XOR2 (N1010, N985, N740);
xor XOR2 (N1011, N1009, N190);
nor NOR4 (N1012, N1007, N370, N302, N447);
nor NOR2 (N1013, N989, N257);
or OR4 (N1014, N1006, N122, N341, N934);
and AND3 (N1015, N1003, N440, N526);
nand NAND2 (N1016, N1015, N764);
nand NAND3 (N1017, N1013, N772, N554);
xor XOR2 (N1018, N1017, N698);
or OR3 (N1019, N1011, N770, N645);
and AND2 (N1020, N1014, N689);
or OR2 (N1021, N1020, N184);
nor NOR2 (N1022, N1001, N444);
nand NAND3 (N1023, N1022, N73, N971);
nand NAND2 (N1024, N987, N71);
not NOT1 (N1025, N1019);
xor XOR2 (N1026, N1018, N1015);
nor NOR2 (N1027, N1008, N210);
nand NAND2 (N1028, N1026, N704);
buf BUF1 (N1029, N1021);
not NOT1 (N1030, N1025);
not NOT1 (N1031, N1027);
buf BUF1 (N1032, N1024);
buf BUF1 (N1033, N1023);
xor XOR2 (N1034, N1010, N733);
not NOT1 (N1035, N1028);
nand NAND2 (N1036, N1034, N489);
xor XOR2 (N1037, N1036, N345);
or OR4 (N1038, N1032, N406, N868, N70);
nor NOR3 (N1039, N1012, N263, N995);
or OR3 (N1040, N1030, N443, N74);
or OR2 (N1041, N1029, N675);
or OR3 (N1042, N1037, N540, N1040);
or OR3 (N1043, N52, N324, N535);
buf BUF1 (N1044, N1005);
nor NOR2 (N1045, N1031, N822);
buf BUF1 (N1046, N1038);
nand NAND4 (N1047, N1039, N326, N542, N56);
not NOT1 (N1048, N1044);
xor XOR2 (N1049, N1041, N467);
xor XOR2 (N1050, N1045, N843);
and AND2 (N1051, N1046, N138);
nor NOR2 (N1052, N1033, N957);
xor XOR2 (N1053, N1049, N319);
nand NAND3 (N1054, N1051, N1019, N813);
nand NAND4 (N1055, N1043, N1010, N530, N755);
not NOT1 (N1056, N1047);
nor NOR2 (N1057, N1042, N1032);
not NOT1 (N1058, N1054);
buf BUF1 (N1059, N1055);
and AND3 (N1060, N1057, N722, N605);
not NOT1 (N1061, N1058);
nor NOR2 (N1062, N1035, N64);
not NOT1 (N1063, N1048);
buf BUF1 (N1064, N1061);
xor XOR2 (N1065, N1050, N904);
buf BUF1 (N1066, N1052);
nand NAND4 (N1067, N1059, N897, N355, N757);
nor NOR2 (N1068, N1053, N327);
not NOT1 (N1069, N1056);
nor NOR2 (N1070, N1067, N492);
buf BUF1 (N1071, N1060);
nand NAND3 (N1072, N1062, N465, N391);
xor XOR2 (N1073, N1071, N453);
not NOT1 (N1074, N1072);
not NOT1 (N1075, N1073);
or OR3 (N1076, N1065, N106, N907);
or OR2 (N1077, N1069, N629);
nand NAND2 (N1078, N1074, N414);
and AND4 (N1079, N1070, N605, N939, N242);
not NOT1 (N1080, N1075);
and AND2 (N1081, N1077, N709);
and AND2 (N1082, N1078, N695);
nor NOR3 (N1083, N1080, N519, N218);
not NOT1 (N1084, N1081);
and AND2 (N1085, N1084, N557);
or OR4 (N1086, N1016, N644, N75, N764);
or OR4 (N1087, N1083, N114, N1012, N372);
buf BUF1 (N1088, N1076);
nand NAND4 (N1089, N1066, N554, N449, N1);
or OR2 (N1090, N1086, N51);
or OR2 (N1091, N1090, N602);
xor XOR2 (N1092, N1082, N961);
not NOT1 (N1093, N1087);
buf BUF1 (N1094, N1093);
or OR4 (N1095, N1092, N216, N776, N317);
or OR2 (N1096, N1091, N545);
nor NOR2 (N1097, N1095, N258);
buf BUF1 (N1098, N1063);
buf BUF1 (N1099, N1097);
buf BUF1 (N1100, N1079);
not NOT1 (N1101, N1089);
nand NAND3 (N1102, N1096, N1063, N1025);
nand NAND3 (N1103, N1101, N1, N301);
nand NAND3 (N1104, N1098, N487, N869);
or OR2 (N1105, N1103, N807);
or OR3 (N1106, N1105, N285, N254);
nor NOR3 (N1107, N1094, N985, N961);
nand NAND2 (N1108, N1099, N759);
buf BUF1 (N1109, N1102);
or OR2 (N1110, N1107, N666);
not NOT1 (N1111, N1085);
or OR2 (N1112, N1100, N969);
and AND4 (N1113, N1088, N1037, N243, N49);
nor NOR4 (N1114, N1108, N59, N402, N937);
and AND2 (N1115, N1112, N1039);
buf BUF1 (N1116, N1111);
xor XOR2 (N1117, N1114, N600);
buf BUF1 (N1118, N1109);
xor XOR2 (N1119, N1118, N744);
nand NAND2 (N1120, N1113, N256);
or OR3 (N1121, N1116, N812, N102);
buf BUF1 (N1122, N1120);
or OR2 (N1123, N1068, N170);
and AND4 (N1124, N1119, N177, N784, N667);
nor NOR2 (N1125, N1104, N206);
and AND2 (N1126, N1125, N763);
or OR4 (N1127, N1121, N601, N459, N21);
buf BUF1 (N1128, N1106);
xor XOR2 (N1129, N1064, N1027);
nor NOR4 (N1130, N1122, N873, N924, N363);
or OR4 (N1131, N1127, N32, N910, N172);
xor XOR2 (N1132, N1126, N147);
nor NOR3 (N1133, N1131, N86, N787);
buf BUF1 (N1134, N1130);
and AND2 (N1135, N1132, N1009);
xor XOR2 (N1136, N1123, N584);
not NOT1 (N1137, N1128);
buf BUF1 (N1138, N1124);
not NOT1 (N1139, N1133);
and AND3 (N1140, N1139, N228, N644);
nand NAND3 (N1141, N1138, N146, N582);
xor XOR2 (N1142, N1135, N615);
buf BUF1 (N1143, N1137);
nor NOR2 (N1144, N1141, N1013);
nor NOR2 (N1145, N1142, N495);
and AND4 (N1146, N1144, N916, N569, N939);
xor XOR2 (N1147, N1136, N144);
or OR4 (N1148, N1115, N215, N439, N454);
buf BUF1 (N1149, N1143);
nor NOR4 (N1150, N1117, N826, N311, N975);
or OR4 (N1151, N1110, N577, N93, N301);
or OR2 (N1152, N1151, N818);
xor XOR2 (N1153, N1145, N733);
not NOT1 (N1154, N1148);
nand NAND2 (N1155, N1146, N15);
nand NAND3 (N1156, N1152, N554, N41);
buf BUF1 (N1157, N1134);
not NOT1 (N1158, N1150);
not NOT1 (N1159, N1140);
and AND3 (N1160, N1158, N1032, N820);
not NOT1 (N1161, N1153);
nor NOR4 (N1162, N1155, N1057, N107, N785);
buf BUF1 (N1163, N1147);
not NOT1 (N1164, N1159);
not NOT1 (N1165, N1157);
buf BUF1 (N1166, N1156);
xor XOR2 (N1167, N1129, N91);
xor XOR2 (N1168, N1149, N632);
or OR2 (N1169, N1160, N698);
nor NOR4 (N1170, N1162, N92, N951, N335);
not NOT1 (N1171, N1154);
not NOT1 (N1172, N1167);
nand NAND4 (N1173, N1165, N591, N278, N189);
nor NOR3 (N1174, N1169, N39, N433);
or OR3 (N1175, N1161, N895, N901);
and AND4 (N1176, N1171, N957, N618, N747);
nor NOR3 (N1177, N1168, N774, N260);
nand NAND3 (N1178, N1175, N155, N308);
nor NOR4 (N1179, N1163, N164, N544, N1076);
not NOT1 (N1180, N1176);
not NOT1 (N1181, N1166);
nor NOR3 (N1182, N1173, N892, N738);
buf BUF1 (N1183, N1164);
nor NOR4 (N1184, N1172, N359, N630, N1070);
or OR4 (N1185, N1170, N510, N148, N1019);
and AND4 (N1186, N1185, N619, N1053, N779);
buf BUF1 (N1187, N1186);
or OR2 (N1188, N1179, N312);
buf BUF1 (N1189, N1183);
and AND2 (N1190, N1182, N940);
and AND2 (N1191, N1187, N285);
and AND3 (N1192, N1188, N90, N323);
nor NOR2 (N1193, N1180, N1091);
nand NAND3 (N1194, N1190, N473, N888);
or OR2 (N1195, N1177, N968);
buf BUF1 (N1196, N1192);
nand NAND4 (N1197, N1194, N385, N851, N1110);
or OR2 (N1198, N1189, N1012);
not NOT1 (N1199, N1178);
and AND3 (N1200, N1174, N770, N398);
nand NAND3 (N1201, N1196, N313, N361);
or OR3 (N1202, N1184, N412, N321);
and AND4 (N1203, N1199, N370, N1070, N848);
nor NOR3 (N1204, N1197, N926, N63);
xor XOR2 (N1205, N1204, N518);
buf BUF1 (N1206, N1181);
or OR4 (N1207, N1205, N686, N1073, N1134);
and AND4 (N1208, N1195, N983, N936, N506);
not NOT1 (N1209, N1208);
or OR3 (N1210, N1201, N31, N520);
buf BUF1 (N1211, N1191);
nand NAND4 (N1212, N1202, N53, N1086, N209);
not NOT1 (N1213, N1211);
and AND3 (N1214, N1198, N83, N60);
buf BUF1 (N1215, N1209);
not NOT1 (N1216, N1210);
nor NOR3 (N1217, N1212, N1104, N501);
xor XOR2 (N1218, N1213, N430);
nor NOR2 (N1219, N1206, N1015);
nor NOR4 (N1220, N1216, N832, N250, N1144);
nand NAND3 (N1221, N1200, N429, N984);
nor NOR4 (N1222, N1215, N1018, N375, N829);
buf BUF1 (N1223, N1222);
and AND4 (N1224, N1221, N124, N504, N1081);
buf BUF1 (N1225, N1217);
nor NOR4 (N1226, N1220, N345, N530, N41);
xor XOR2 (N1227, N1224, N926);
nand NAND2 (N1228, N1227, N452);
nand NAND3 (N1229, N1228, N905, N976);
xor XOR2 (N1230, N1214, N15);
or OR2 (N1231, N1223, N657);
nand NAND2 (N1232, N1229, N677);
not NOT1 (N1233, N1225);
nor NOR4 (N1234, N1232, N463, N955, N652);
nand NAND3 (N1235, N1230, N955, N498);
nand NAND3 (N1236, N1231, N521, N443);
or OR3 (N1237, N1203, N95, N202);
xor XOR2 (N1238, N1207, N879);
nor NOR4 (N1239, N1193, N1045, N894, N868);
not NOT1 (N1240, N1234);
nor NOR4 (N1241, N1239, N916, N919, N576);
nor NOR3 (N1242, N1226, N898, N511);
nor NOR4 (N1243, N1235, N121, N1029, N283);
nand NAND2 (N1244, N1236, N907);
nor NOR3 (N1245, N1238, N792, N364);
buf BUF1 (N1246, N1237);
and AND4 (N1247, N1233, N1126, N379, N44);
xor XOR2 (N1248, N1243, N403);
and AND4 (N1249, N1218, N996, N593, N554);
buf BUF1 (N1250, N1242);
nor NOR3 (N1251, N1219, N246, N39);
and AND2 (N1252, N1251, N371);
nand NAND4 (N1253, N1241, N79, N1115, N859);
buf BUF1 (N1254, N1247);
buf BUF1 (N1255, N1244);
or OR2 (N1256, N1255, N11);
nand NAND3 (N1257, N1253, N670, N213);
xor XOR2 (N1258, N1252, N28);
not NOT1 (N1259, N1256);
or OR3 (N1260, N1257, N943, N769);
or OR2 (N1261, N1248, N899);
or OR3 (N1262, N1260, N984, N366);
not NOT1 (N1263, N1259);
and AND2 (N1264, N1250, N165);
and AND2 (N1265, N1249, N549);
nor NOR2 (N1266, N1265, N447);
nand NAND3 (N1267, N1262, N582, N733);
and AND3 (N1268, N1266, N45, N915);
nor NOR3 (N1269, N1246, N730, N1012);
not NOT1 (N1270, N1267);
nand NAND3 (N1271, N1245, N897, N1247);
xor XOR2 (N1272, N1240, N204);
nand NAND3 (N1273, N1268, N292, N1262);
nor NOR4 (N1274, N1261, N1031, N1028, N14);
xor XOR2 (N1275, N1263, N754);
not NOT1 (N1276, N1269);
buf BUF1 (N1277, N1276);
nor NOR3 (N1278, N1273, N24, N505);
or OR3 (N1279, N1274, N222, N848);
not NOT1 (N1280, N1277);
nor NOR2 (N1281, N1280, N262);
nor NOR4 (N1282, N1258, N624, N236, N376);
or OR3 (N1283, N1254, N164, N1189);
or OR4 (N1284, N1282, N257, N768, N63);
xor XOR2 (N1285, N1264, N164);
not NOT1 (N1286, N1279);
nand NAND2 (N1287, N1275, N1073);
nand NAND3 (N1288, N1272, N1260, N1259);
nand NAND4 (N1289, N1288, N144, N589, N188);
and AND3 (N1290, N1271, N1125, N608);
nor NOR3 (N1291, N1284, N284, N842);
or OR2 (N1292, N1278, N637);
not NOT1 (N1293, N1270);
buf BUF1 (N1294, N1287);
nand NAND2 (N1295, N1290, N167);
not NOT1 (N1296, N1292);
xor XOR2 (N1297, N1293, N50);
nor NOR4 (N1298, N1285, N1144, N4, N652);
or OR2 (N1299, N1294, N30);
xor XOR2 (N1300, N1291, N1019);
nor NOR4 (N1301, N1296, N851, N903, N394);
nand NAND3 (N1302, N1298, N663, N403);
buf BUF1 (N1303, N1301);
buf BUF1 (N1304, N1297);
nor NOR3 (N1305, N1286, N117, N965);
and AND4 (N1306, N1303, N1078, N1038, N65);
and AND2 (N1307, N1302, N899);
nor NOR3 (N1308, N1281, N785, N773);
xor XOR2 (N1309, N1307, N70);
not NOT1 (N1310, N1306);
nor NOR3 (N1311, N1299, N76, N693);
and AND2 (N1312, N1311, N847);
or OR3 (N1313, N1305, N1100, N1115);
and AND4 (N1314, N1295, N1282, N968, N158);
not NOT1 (N1315, N1314);
xor XOR2 (N1316, N1304, N811);
xor XOR2 (N1317, N1315, N171);
nor NOR3 (N1318, N1312, N289, N430);
not NOT1 (N1319, N1310);
buf BUF1 (N1320, N1308);
nor NOR4 (N1321, N1320, N657, N957, N3);
buf BUF1 (N1322, N1319);
nand NAND2 (N1323, N1317, N1127);
not NOT1 (N1324, N1321);
xor XOR2 (N1325, N1323, N1085);
buf BUF1 (N1326, N1313);
buf BUF1 (N1327, N1283);
and AND3 (N1328, N1327, N915, N859);
nand NAND3 (N1329, N1326, N446, N152);
nor NOR4 (N1330, N1324, N963, N736, N642);
nor NOR2 (N1331, N1329, N912);
buf BUF1 (N1332, N1300);
not NOT1 (N1333, N1322);
or OR3 (N1334, N1309, N1019, N346);
not NOT1 (N1335, N1325);
or OR2 (N1336, N1334, N972);
nand NAND4 (N1337, N1331, N441, N377, N955);
or OR4 (N1338, N1336, N1331, N428, N353);
or OR4 (N1339, N1289, N14, N346, N1131);
xor XOR2 (N1340, N1337, N842);
not NOT1 (N1341, N1328);
and AND2 (N1342, N1340, N355);
or OR3 (N1343, N1339, N212, N155);
and AND2 (N1344, N1316, N1302);
and AND3 (N1345, N1344, N354, N950);
or OR2 (N1346, N1318, N1299);
not NOT1 (N1347, N1330);
xor XOR2 (N1348, N1346, N142);
nor NOR2 (N1349, N1348, N1074);
not NOT1 (N1350, N1347);
or OR2 (N1351, N1343, N653);
nor NOR4 (N1352, N1350, N460, N1316, N1029);
and AND3 (N1353, N1338, N430, N694);
not NOT1 (N1354, N1345);
buf BUF1 (N1355, N1354);
nand NAND3 (N1356, N1342, N1202, N556);
nor NOR2 (N1357, N1341, N537);
and AND4 (N1358, N1356, N1318, N854, N876);
nand NAND2 (N1359, N1333, N182);
xor XOR2 (N1360, N1359, N1216);
or OR2 (N1361, N1352, N1292);
nand NAND3 (N1362, N1332, N875, N794);
or OR3 (N1363, N1361, N515, N1052);
not NOT1 (N1364, N1351);
and AND2 (N1365, N1363, N1058);
nand NAND2 (N1366, N1360, N110);
or OR2 (N1367, N1365, N961);
xor XOR2 (N1368, N1362, N459);
nor NOR4 (N1369, N1353, N1111, N494, N1158);
buf BUF1 (N1370, N1364);
not NOT1 (N1371, N1357);
or OR3 (N1372, N1335, N936, N594);
xor XOR2 (N1373, N1358, N441);
nor NOR4 (N1374, N1372, N929, N633, N318);
nand NAND2 (N1375, N1366, N523);
buf BUF1 (N1376, N1355);
not NOT1 (N1377, N1368);
buf BUF1 (N1378, N1369);
xor XOR2 (N1379, N1376, N1286);
and AND3 (N1380, N1379, N1323, N918);
or OR3 (N1381, N1374, N1014, N674);
or OR2 (N1382, N1380, N190);
and AND2 (N1383, N1367, N999);
xor XOR2 (N1384, N1373, N555);
and AND4 (N1385, N1371, N1218, N191, N999);
nand NAND2 (N1386, N1377, N767);
and AND3 (N1387, N1382, N968, N1266);
buf BUF1 (N1388, N1385);
nand NAND3 (N1389, N1387, N886, N108);
xor XOR2 (N1390, N1388, N840);
or OR2 (N1391, N1375, N1156);
xor XOR2 (N1392, N1386, N732);
nor NOR4 (N1393, N1392, N1186, N299, N823);
or OR3 (N1394, N1389, N393, N690);
xor XOR2 (N1395, N1349, N1021);
and AND2 (N1396, N1383, N266);
nor NOR4 (N1397, N1381, N1110, N382, N1248);
xor XOR2 (N1398, N1397, N846);
nor NOR4 (N1399, N1391, N123, N167, N654);
or OR3 (N1400, N1399, N1119, N1384);
nor NOR4 (N1401, N212, N900, N508, N177);
xor XOR2 (N1402, N1393, N436);
not NOT1 (N1403, N1401);
nor NOR3 (N1404, N1370, N852, N516);
nand NAND3 (N1405, N1396, N498, N884);
not NOT1 (N1406, N1402);
nand NAND4 (N1407, N1378, N790, N11, N300);
and AND3 (N1408, N1394, N626, N310);
xor XOR2 (N1409, N1398, N206);
and AND2 (N1410, N1409, N1162);
xor XOR2 (N1411, N1407, N1148);
not NOT1 (N1412, N1395);
nand NAND3 (N1413, N1404, N1243, N209);
not NOT1 (N1414, N1406);
and AND2 (N1415, N1390, N1171);
nor NOR3 (N1416, N1414, N959, N810);
and AND4 (N1417, N1416, N241, N798, N125);
nand NAND3 (N1418, N1408, N1040, N1069);
nand NAND4 (N1419, N1413, N1173, N1125, N562);
xor XOR2 (N1420, N1415, N1318);
and AND2 (N1421, N1412, N1205);
xor XOR2 (N1422, N1420, N166);
and AND2 (N1423, N1417, N32);
nor NOR3 (N1424, N1411, N1086, N560);
buf BUF1 (N1425, N1421);
nor NOR2 (N1426, N1418, N255);
and AND4 (N1427, N1426, N348, N781, N460);
buf BUF1 (N1428, N1419);
nor NOR4 (N1429, N1424, N1310, N637, N1033);
and AND3 (N1430, N1427, N938, N977);
nand NAND2 (N1431, N1405, N576);
or OR2 (N1432, N1423, N449);
and AND4 (N1433, N1422, N304, N670, N881);
buf BUF1 (N1434, N1431);
and AND3 (N1435, N1428, N596, N13);
buf BUF1 (N1436, N1430);
buf BUF1 (N1437, N1434);
xor XOR2 (N1438, N1432, N1030);
and AND3 (N1439, N1437, N448, N8);
nand NAND4 (N1440, N1436, N192, N657, N1209);
not NOT1 (N1441, N1440);
buf BUF1 (N1442, N1403);
or OR4 (N1443, N1433, N265, N360, N244);
or OR4 (N1444, N1443, N814, N737, N283);
xor XOR2 (N1445, N1425, N1055);
or OR2 (N1446, N1438, N646);
not NOT1 (N1447, N1435);
and AND4 (N1448, N1441, N1282, N848, N1246);
buf BUF1 (N1449, N1446);
nor NOR2 (N1450, N1400, N705);
or OR2 (N1451, N1449, N946);
nor NOR2 (N1452, N1450, N886);
not NOT1 (N1453, N1439);
not NOT1 (N1454, N1445);
and AND3 (N1455, N1410, N1050, N874);
and AND4 (N1456, N1454, N581, N267, N8);
not NOT1 (N1457, N1447);
xor XOR2 (N1458, N1444, N1151);
and AND3 (N1459, N1448, N269, N74);
not NOT1 (N1460, N1456);
and AND4 (N1461, N1453, N644, N963, N313);
not NOT1 (N1462, N1458);
buf BUF1 (N1463, N1461);
nand NAND3 (N1464, N1457, N529, N1323);
buf BUF1 (N1465, N1463);
xor XOR2 (N1466, N1455, N1171);
nor NOR3 (N1467, N1465, N1376, N533);
not NOT1 (N1468, N1452);
not NOT1 (N1469, N1460);
not NOT1 (N1470, N1469);
buf BUF1 (N1471, N1464);
and AND4 (N1472, N1471, N658, N834, N387);
or OR3 (N1473, N1470, N1087, N469);
not NOT1 (N1474, N1451);
and AND2 (N1475, N1429, N138);
or OR4 (N1476, N1473, N410, N1013, N1040);
not NOT1 (N1477, N1459);
xor XOR2 (N1478, N1468, N1404);
xor XOR2 (N1479, N1466, N1445);
nand NAND2 (N1480, N1462, N1003);
xor XOR2 (N1481, N1476, N764);
nand NAND2 (N1482, N1478, N159);
nand NAND4 (N1483, N1475, N1041, N1253, N1256);
nor NOR2 (N1484, N1480, N670);
buf BUF1 (N1485, N1474);
not NOT1 (N1486, N1483);
nand NAND4 (N1487, N1482, N994, N769, N939);
buf BUF1 (N1488, N1484);
and AND3 (N1489, N1477, N245, N1304);
or OR2 (N1490, N1472, N237);
nand NAND4 (N1491, N1442, N908, N279, N517);
and AND4 (N1492, N1485, N973, N231, N179);
and AND3 (N1493, N1488, N534, N374);
nor NOR2 (N1494, N1492, N831);
not NOT1 (N1495, N1486);
nand NAND3 (N1496, N1493, N219, N693);
xor XOR2 (N1497, N1481, N189);
xor XOR2 (N1498, N1490, N765);
buf BUF1 (N1499, N1467);
xor XOR2 (N1500, N1497, N52);
nor NOR3 (N1501, N1500, N1369, N48);
not NOT1 (N1502, N1487);
not NOT1 (N1503, N1496);
not NOT1 (N1504, N1479);
nor NOR3 (N1505, N1501, N264, N1307);
or OR3 (N1506, N1489, N596, N1106);
not NOT1 (N1507, N1502);
nor NOR3 (N1508, N1504, N222, N1274);
and AND3 (N1509, N1505, N462, N90);
xor XOR2 (N1510, N1508, N163);
or OR4 (N1511, N1503, N949, N136, N208);
or OR2 (N1512, N1506, N1489);
nor NOR3 (N1513, N1491, N343, N522);
not NOT1 (N1514, N1498);
nand NAND4 (N1515, N1509, N520, N101, N650);
and AND2 (N1516, N1494, N727);
or OR4 (N1517, N1514, N1098, N874, N1296);
xor XOR2 (N1518, N1507, N1501);
buf BUF1 (N1519, N1511);
buf BUF1 (N1520, N1510);
nand NAND2 (N1521, N1518, N1194);
xor XOR2 (N1522, N1521, N906);
not NOT1 (N1523, N1516);
buf BUF1 (N1524, N1512);
or OR3 (N1525, N1495, N1033, N612);
and AND4 (N1526, N1515, N659, N360, N1424);
nor NOR4 (N1527, N1524, N347, N1433, N312);
not NOT1 (N1528, N1519);
or OR2 (N1529, N1523, N1484);
xor XOR2 (N1530, N1513, N227);
nand NAND3 (N1531, N1527, N37, N928);
not NOT1 (N1532, N1530);
buf BUF1 (N1533, N1525);
and AND2 (N1534, N1531, N1159);
nand NAND2 (N1535, N1520, N510);
nor NOR3 (N1536, N1526, N541, N827);
or OR3 (N1537, N1532, N108, N1384);
not NOT1 (N1538, N1499);
nor NOR2 (N1539, N1537, N1043);
nand NAND4 (N1540, N1535, N449, N882, N233);
not NOT1 (N1541, N1533);
or OR3 (N1542, N1534, N1515, N1232);
and AND4 (N1543, N1536, N1426, N59, N1369);
and AND4 (N1544, N1540, N489, N1166, N491);
or OR2 (N1545, N1542, N1041);
nand NAND3 (N1546, N1544, N1478, N1181);
and AND3 (N1547, N1522, N239, N85);
xor XOR2 (N1548, N1539, N774);
or OR4 (N1549, N1547, N945, N669, N736);
and AND3 (N1550, N1538, N1113, N1440);
not NOT1 (N1551, N1545);
nand NAND3 (N1552, N1548, N64, N810);
xor XOR2 (N1553, N1550, N408);
not NOT1 (N1554, N1529);
buf BUF1 (N1555, N1541);
xor XOR2 (N1556, N1517, N1144);
and AND2 (N1557, N1552, N410);
and AND2 (N1558, N1551, N331);
nand NAND4 (N1559, N1557, N1115, N1232, N1254);
nand NAND4 (N1560, N1555, N491, N1514, N529);
nor NOR3 (N1561, N1558, N444, N410);
nand NAND2 (N1562, N1559, N698);
not NOT1 (N1563, N1549);
and AND3 (N1564, N1561, N1046, N1448);
and AND2 (N1565, N1560, N415);
not NOT1 (N1566, N1562);
not NOT1 (N1567, N1554);
and AND4 (N1568, N1553, N131, N807, N40);
buf BUF1 (N1569, N1528);
or OR4 (N1570, N1565, N813, N46, N91);
and AND3 (N1571, N1563, N580, N736);
nand NAND3 (N1572, N1567, N1252, N432);
or OR3 (N1573, N1556, N1282, N111);
buf BUF1 (N1574, N1571);
nand NAND2 (N1575, N1573, N914);
xor XOR2 (N1576, N1569, N783);
and AND4 (N1577, N1570, N5, N1281, N461);
xor XOR2 (N1578, N1577, N239);
or OR3 (N1579, N1576, N592, N1349);
or OR3 (N1580, N1572, N1353, N600);
or OR2 (N1581, N1574, N1505);
nor NOR2 (N1582, N1575, N1148);
buf BUF1 (N1583, N1566);
and AND4 (N1584, N1546, N1365, N932, N37);
buf BUF1 (N1585, N1579);
buf BUF1 (N1586, N1564);
nor NOR2 (N1587, N1586, N1075);
xor XOR2 (N1588, N1581, N847);
not NOT1 (N1589, N1587);
xor XOR2 (N1590, N1583, N1377);
nand NAND3 (N1591, N1568, N679, N543);
and AND2 (N1592, N1585, N917);
and AND2 (N1593, N1589, N1254);
xor XOR2 (N1594, N1593, N1505);
not NOT1 (N1595, N1580);
nor NOR4 (N1596, N1591, N1224, N1567, N872);
nand NAND4 (N1597, N1596, N1551, N241, N811);
nor NOR2 (N1598, N1582, N365);
xor XOR2 (N1599, N1595, N916);
nor NOR4 (N1600, N1588, N147, N547, N81);
nand NAND4 (N1601, N1594, N430, N315, N1266);
not NOT1 (N1602, N1597);
not NOT1 (N1603, N1601);
nor NOR3 (N1604, N1598, N843, N1477);
nor NOR3 (N1605, N1604, N1465, N549);
nor NOR4 (N1606, N1543, N1531, N1590, N1589);
not NOT1 (N1607, N775);
buf BUF1 (N1608, N1592);
nand NAND4 (N1609, N1600, N344, N21, N418);
nor NOR2 (N1610, N1605, N1492);
nand NAND2 (N1611, N1610, N354);
not NOT1 (N1612, N1578);
xor XOR2 (N1613, N1599, N306);
and AND4 (N1614, N1606, N398, N1260, N297);
and AND3 (N1615, N1614, N405, N1370);
not NOT1 (N1616, N1613);
or OR3 (N1617, N1608, N121, N1115);
buf BUF1 (N1618, N1616);
nand NAND4 (N1619, N1611, N312, N444, N794);
endmodule