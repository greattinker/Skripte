// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N16013,N15996,N16011,N16009,N16012,N16016,N16015,N15963,N16007,N16018;

nand NAND4 (N19, N12, N7, N3, N2);
and AND3 (N20, N13, N15, N7);
and AND3 (N21, N17, N8, N9);
nand NAND2 (N22, N10, N18);
or OR2 (N23, N13, N10);
xor XOR2 (N24, N6, N12);
or OR3 (N25, N23, N15, N11);
nor NOR2 (N26, N19, N15);
or OR3 (N27, N18, N3, N8);
nand NAND3 (N28, N20, N27, N6);
or OR2 (N29, N9, N24);
nand NAND2 (N30, N25, N23);
buf BUF1 (N31, N7);
or OR2 (N32, N15, N11);
not NOT1 (N33, N21);
nor NOR4 (N34, N10, N7, N5, N24);
and AND2 (N35, N34, N10);
nor NOR3 (N36, N11, N33, N7);
xor XOR2 (N37, N13, N8);
xor XOR2 (N38, N26, N3);
and AND3 (N39, N22, N32, N11);
or OR4 (N40, N27, N27, N38, N3);
nand NAND3 (N41, N25, N25, N16);
or OR4 (N42, N41, N35, N36, N41);
xor XOR2 (N43, N9, N40);
and AND4 (N44, N14, N41, N22, N2);
nand NAND2 (N45, N43, N33);
buf BUF1 (N46, N22);
or OR2 (N47, N37, N4);
nor NOR4 (N48, N42, N36, N16, N15);
nor NOR3 (N49, N30, N9, N3);
buf BUF1 (N50, N45);
xor XOR2 (N51, N28, N4);
and AND4 (N52, N48, N19, N42, N33);
xor XOR2 (N53, N46, N32);
buf BUF1 (N54, N49);
buf BUF1 (N55, N51);
not NOT1 (N56, N53);
buf BUF1 (N57, N39);
xor XOR2 (N58, N52, N28);
and AND2 (N59, N29, N48);
and AND3 (N60, N54, N31, N7);
nor NOR3 (N61, N57, N20, N50);
xor XOR2 (N62, N30, N12);
xor XOR2 (N63, N54, N45);
or OR3 (N64, N58, N32, N29);
nand NAND3 (N65, N47, N5, N64);
nand NAND4 (N66, N58, N8, N30, N50);
xor XOR2 (N67, N61, N43);
not NOT1 (N68, N56);
not NOT1 (N69, N59);
and AND4 (N70, N63, N21, N54, N62);
nand NAND3 (N71, N65, N61, N62);
and AND2 (N72, N42, N56);
xor XOR2 (N73, N66, N3);
not NOT1 (N74, N67);
not NOT1 (N75, N68);
and AND4 (N76, N73, N29, N11, N25);
not NOT1 (N77, N70);
nand NAND4 (N78, N76, N77, N11, N51);
not NOT1 (N79, N46);
xor XOR2 (N80, N75, N55);
and AND4 (N81, N10, N59, N14, N10);
nor NOR2 (N82, N80, N60);
buf BUF1 (N83, N23);
and AND2 (N84, N81, N17);
not NOT1 (N85, N74);
nor NOR3 (N86, N71, N22, N70);
buf BUF1 (N87, N79);
buf BUF1 (N88, N87);
buf BUF1 (N89, N84);
and AND2 (N90, N44, N15);
xor XOR2 (N91, N88, N2);
nor NOR2 (N92, N91, N7);
xor XOR2 (N93, N82, N21);
xor XOR2 (N94, N69, N62);
xor XOR2 (N95, N72, N42);
not NOT1 (N96, N78);
and AND3 (N97, N83, N44, N36);
and AND3 (N98, N92, N59, N70);
not NOT1 (N99, N94);
nor NOR4 (N100, N96, N65, N63, N9);
buf BUF1 (N101, N99);
xor XOR2 (N102, N93, N43);
not NOT1 (N103, N89);
nand NAND3 (N104, N100, N61, N50);
not NOT1 (N105, N95);
not NOT1 (N106, N86);
or OR2 (N107, N104, N100);
xor XOR2 (N108, N102, N46);
nor NOR2 (N109, N103, N28);
not NOT1 (N110, N108);
or OR3 (N111, N97, N87, N2);
nand NAND4 (N112, N85, N7, N73, N78);
nor NOR4 (N113, N111, N16, N10, N89);
not NOT1 (N114, N113);
buf BUF1 (N115, N106);
xor XOR2 (N116, N98, N115);
xor XOR2 (N117, N24, N58);
xor XOR2 (N118, N109, N50);
or OR2 (N119, N116, N34);
or OR4 (N120, N110, N8, N69, N47);
nor NOR4 (N121, N120, N116, N95, N53);
xor XOR2 (N122, N117, N76);
and AND3 (N123, N101, N50, N83);
nand NAND2 (N124, N122, N99);
not NOT1 (N125, N124);
and AND3 (N126, N118, N31, N120);
and AND4 (N127, N125, N25, N77, N107);
buf BUF1 (N128, N25);
xor XOR2 (N129, N128, N123);
buf BUF1 (N130, N105);
or OR4 (N131, N13, N74, N30, N83);
not NOT1 (N132, N130);
or OR4 (N133, N119, N85, N107, N107);
buf BUF1 (N134, N127);
xor XOR2 (N135, N131, N92);
and AND2 (N136, N135, N126);
and AND2 (N137, N16, N88);
not NOT1 (N138, N132);
and AND3 (N139, N137, N122, N86);
xor XOR2 (N140, N138, N116);
xor XOR2 (N141, N114, N96);
xor XOR2 (N142, N136, N124);
nor NOR2 (N143, N133, N26);
xor XOR2 (N144, N139, N77);
or OR2 (N145, N90, N140);
nor NOR2 (N146, N69, N85);
not NOT1 (N147, N145);
nand NAND2 (N148, N144, N81);
or OR2 (N149, N142, N33);
not NOT1 (N150, N134);
or OR3 (N151, N129, N143, N18);
buf BUF1 (N152, N74);
xor XOR2 (N153, N147, N131);
xor XOR2 (N154, N146, N29);
or OR4 (N155, N151, N73, N62, N57);
nor NOR3 (N156, N141, N116, N68);
nand NAND4 (N157, N155, N61, N40, N118);
buf BUF1 (N158, N156);
not NOT1 (N159, N152);
xor XOR2 (N160, N112, N57);
buf BUF1 (N161, N158);
buf BUF1 (N162, N148);
or OR2 (N163, N160, N18);
xor XOR2 (N164, N150, N149);
or OR4 (N165, N108, N145, N118, N73);
and AND4 (N166, N164, N155, N33, N73);
nand NAND3 (N167, N154, N71, N118);
and AND3 (N168, N163, N56, N85);
not NOT1 (N169, N166);
xor XOR2 (N170, N161, N53);
not NOT1 (N171, N169);
nor NOR3 (N172, N165, N53, N66);
and AND3 (N173, N171, N104, N164);
xor XOR2 (N174, N170, N64);
xor XOR2 (N175, N159, N52);
nor NOR2 (N176, N172, N70);
nor NOR3 (N177, N173, N126, N104);
buf BUF1 (N178, N175);
not NOT1 (N179, N177);
xor XOR2 (N180, N153, N131);
buf BUF1 (N181, N178);
xor XOR2 (N182, N167, N11);
xor XOR2 (N183, N181, N124);
xor XOR2 (N184, N179, N65);
xor XOR2 (N185, N182, N97);
not NOT1 (N186, N121);
xor XOR2 (N187, N183, N88);
or OR4 (N188, N174, N69, N34, N174);
and AND4 (N189, N162, N135, N158, N103);
or OR2 (N190, N168, N27);
nand NAND4 (N191, N187, N160, N61, N12);
nor NOR3 (N192, N188, N167, N98);
or OR4 (N193, N185, N131, N155, N172);
xor XOR2 (N194, N157, N187);
buf BUF1 (N195, N194);
or OR2 (N196, N190, N4);
nand NAND2 (N197, N195, N149);
buf BUF1 (N198, N191);
nand NAND3 (N199, N176, N89, N83);
or OR3 (N200, N196, N82, N115);
buf BUF1 (N201, N186);
not NOT1 (N202, N193);
and AND4 (N203, N180, N178, N166, N97);
xor XOR2 (N204, N199, N15);
nor NOR3 (N205, N203, N50, N138);
buf BUF1 (N206, N204);
nor NOR2 (N207, N206, N50);
and AND4 (N208, N207, N38, N147, N90);
xor XOR2 (N209, N201, N30);
or OR4 (N210, N208, N150, N140, N77);
and AND3 (N211, N198, N75, N120);
and AND3 (N212, N209, N47, N111);
not NOT1 (N213, N200);
nand NAND4 (N214, N192, N197, N19, N27);
and AND3 (N215, N168, N177, N122);
or OR4 (N216, N213, N147, N124, N96);
and AND4 (N217, N211, N29, N165, N160);
nand NAND2 (N218, N205, N17);
or OR2 (N219, N217, N131);
or OR2 (N220, N184, N22);
and AND4 (N221, N219, N118, N28, N127);
and AND2 (N222, N220, N157);
xor XOR2 (N223, N214, N165);
and AND3 (N224, N218, N21, N8);
and AND4 (N225, N189, N79, N152, N191);
xor XOR2 (N226, N224, N1);
xor XOR2 (N227, N225, N191);
nor NOR2 (N228, N210, N189);
xor XOR2 (N229, N222, N99);
not NOT1 (N230, N229);
xor XOR2 (N231, N227, N1);
not NOT1 (N232, N221);
or OR4 (N233, N230, N135, N200, N174);
nand NAND4 (N234, N223, N44, N212, N126);
or OR3 (N235, N45, N104, N128);
and AND4 (N236, N216, N106, N93, N19);
not NOT1 (N237, N236);
buf BUF1 (N238, N232);
not NOT1 (N239, N237);
not NOT1 (N240, N239);
not NOT1 (N241, N235);
buf BUF1 (N242, N234);
xor XOR2 (N243, N202, N82);
not NOT1 (N244, N238);
and AND2 (N245, N242, N9);
xor XOR2 (N246, N233, N124);
xor XOR2 (N247, N240, N29);
nand NAND3 (N248, N243, N154, N150);
buf BUF1 (N249, N244);
or OR3 (N250, N215, N231, N147);
nand NAND4 (N251, N104, N98, N90, N27);
nand NAND3 (N252, N247, N111, N135);
nand NAND4 (N253, N249, N218, N24, N159);
not NOT1 (N254, N248);
nor NOR4 (N255, N251, N135, N219, N48);
not NOT1 (N256, N241);
nor NOR2 (N257, N245, N20);
nand NAND2 (N258, N256, N209);
xor XOR2 (N259, N257, N198);
buf BUF1 (N260, N226);
nor NOR3 (N261, N246, N180, N204);
and AND2 (N262, N253, N10);
and AND4 (N263, N250, N90, N71, N154);
not NOT1 (N264, N260);
nor NOR3 (N265, N261, N158, N6);
buf BUF1 (N266, N228);
nor NOR2 (N267, N266, N158);
and AND3 (N268, N258, N231, N49);
not NOT1 (N269, N263);
buf BUF1 (N270, N265);
buf BUF1 (N271, N269);
xor XOR2 (N272, N264, N92);
xor XOR2 (N273, N255, N60);
not NOT1 (N274, N273);
nor NOR3 (N275, N259, N115, N191);
nand NAND4 (N276, N268, N176, N228, N84);
or OR2 (N277, N271, N141);
nand NAND4 (N278, N272, N45, N127, N192);
and AND4 (N279, N252, N168, N50, N36);
buf BUF1 (N280, N278);
nor NOR3 (N281, N254, N61, N232);
not NOT1 (N282, N267);
or OR4 (N283, N270, N184, N137, N34);
nand NAND4 (N284, N280, N95, N160, N169);
not NOT1 (N285, N284);
and AND3 (N286, N277, N2, N117);
buf BUF1 (N287, N285);
nand NAND3 (N288, N287, N266, N58);
buf BUF1 (N289, N276);
not NOT1 (N290, N283);
not NOT1 (N291, N288);
not NOT1 (N292, N289);
or OR2 (N293, N275, N174);
nor NOR2 (N294, N291, N27);
not NOT1 (N295, N274);
or OR4 (N296, N295, N256, N85, N14);
xor XOR2 (N297, N294, N28);
xor XOR2 (N298, N279, N14);
and AND4 (N299, N297, N28, N88, N199);
xor XOR2 (N300, N296, N101);
and AND4 (N301, N262, N174, N191, N140);
or OR4 (N302, N282, N76, N209, N201);
and AND4 (N303, N302, N39, N85, N290);
nor NOR4 (N304, N136, N22, N112, N113);
buf BUF1 (N305, N298);
nand NAND3 (N306, N305, N285, N43);
and AND4 (N307, N306, N257, N87, N278);
and AND3 (N308, N292, N296, N190);
buf BUF1 (N309, N286);
buf BUF1 (N310, N300);
nor NOR4 (N311, N299, N7, N183, N2);
nand NAND2 (N312, N301, N9);
buf BUF1 (N313, N312);
and AND3 (N314, N304, N32, N231);
buf BUF1 (N315, N303);
nand NAND3 (N316, N293, N8, N275);
not NOT1 (N317, N281);
nand NAND3 (N318, N317, N310, N110);
nand NAND2 (N319, N291, N105);
and AND2 (N320, N315, N138);
nor NOR2 (N321, N307, N282);
xor XOR2 (N322, N308, N19);
nor NOR3 (N323, N313, N83, N72);
nand NAND4 (N324, N321, N277, N201, N201);
nor NOR3 (N325, N309, N277, N165);
buf BUF1 (N326, N324);
buf BUF1 (N327, N318);
not NOT1 (N328, N320);
or OR4 (N329, N323, N13, N291, N85);
nor NOR4 (N330, N311, N222, N251, N122);
or OR4 (N331, N328, N206, N117, N10);
and AND2 (N332, N331, N206);
and AND3 (N333, N325, N15, N319);
nand NAND3 (N334, N272, N31, N40);
or OR4 (N335, N314, N94, N155, N239);
nand NAND4 (N336, N327, N58, N330, N67);
xor XOR2 (N337, N234, N168);
not NOT1 (N338, N322);
xor XOR2 (N339, N332, N182);
or OR4 (N340, N333, N195, N61, N249);
or OR2 (N341, N334, N165);
buf BUF1 (N342, N326);
nand NAND2 (N343, N316, N102);
buf BUF1 (N344, N336);
nand NAND4 (N345, N341, N33, N210, N254);
nor NOR3 (N346, N339, N280, N115);
buf BUF1 (N347, N344);
nand NAND4 (N348, N338, N140, N140, N40);
nor NOR4 (N349, N348, N212, N122, N334);
nand NAND4 (N350, N337, N60, N249, N4);
nand NAND4 (N351, N342, N308, N228, N7);
nor NOR4 (N352, N343, N44, N312, N331);
nand NAND4 (N353, N352, N334, N342, N15);
xor XOR2 (N354, N329, N130);
xor XOR2 (N355, N335, N345);
not NOT1 (N356, N165);
nor NOR4 (N357, N350, N313, N130, N225);
nor NOR4 (N358, N347, N185, N265, N39);
nor NOR3 (N359, N357, N312, N181);
not NOT1 (N360, N349);
and AND3 (N361, N355, N58, N20);
nand NAND3 (N362, N360, N294, N224);
and AND2 (N363, N354, N135);
or OR4 (N364, N358, N82, N98, N51);
nand NAND2 (N365, N351, N139);
and AND2 (N366, N340, N292);
nand NAND3 (N367, N366, N90, N252);
nor NOR3 (N368, N365, N318, N284);
nor NOR3 (N369, N356, N161, N301);
nand NAND2 (N370, N367, N34);
buf BUF1 (N371, N369);
buf BUF1 (N372, N371);
buf BUF1 (N373, N346);
not NOT1 (N374, N364);
nor NOR2 (N375, N368, N200);
xor XOR2 (N376, N374, N171);
nor NOR3 (N377, N375, N195, N172);
nor NOR4 (N378, N362, N61, N116, N153);
and AND2 (N379, N378, N16);
and AND4 (N380, N379, N129, N169, N8);
xor XOR2 (N381, N372, N353);
nand NAND4 (N382, N302, N337, N28, N28);
or OR2 (N383, N382, N87);
and AND2 (N384, N381, N138);
and AND2 (N385, N380, N305);
xor XOR2 (N386, N383, N169);
xor XOR2 (N387, N370, N321);
not NOT1 (N388, N386);
xor XOR2 (N389, N377, N358);
nor NOR2 (N390, N359, N308);
not NOT1 (N391, N363);
buf BUF1 (N392, N385);
and AND3 (N393, N388, N260, N307);
nand NAND2 (N394, N373, N145);
nand NAND2 (N395, N393, N377);
xor XOR2 (N396, N361, N152);
nand NAND2 (N397, N387, N312);
xor XOR2 (N398, N376, N244);
nand NAND2 (N399, N398, N343);
and AND2 (N400, N394, N241);
buf BUF1 (N401, N395);
nand NAND3 (N402, N384, N209, N205);
buf BUF1 (N403, N390);
and AND3 (N404, N391, N171, N45);
nor NOR4 (N405, N392, N137, N186, N204);
nor NOR3 (N406, N403, N142, N300);
and AND3 (N407, N405, N28, N84);
and AND2 (N408, N406, N135);
buf BUF1 (N409, N408);
nand NAND2 (N410, N397, N93);
nand NAND2 (N411, N401, N322);
nor NOR4 (N412, N402, N98, N196, N379);
not NOT1 (N413, N400);
and AND4 (N414, N412, N80, N209, N326);
buf BUF1 (N415, N389);
not NOT1 (N416, N404);
nor NOR3 (N417, N410, N304, N378);
and AND2 (N418, N399, N386);
not NOT1 (N419, N409);
or OR2 (N420, N415, N219);
nand NAND4 (N421, N411, N417, N352, N38);
or OR3 (N422, N5, N335, N271);
not NOT1 (N423, N421);
not NOT1 (N424, N407);
xor XOR2 (N425, N418, N37);
xor XOR2 (N426, N424, N251);
or OR2 (N427, N416, N41);
nand NAND3 (N428, N423, N257, N294);
buf BUF1 (N429, N427);
and AND4 (N430, N414, N40, N381, N189);
not NOT1 (N431, N413);
buf BUF1 (N432, N419);
not NOT1 (N433, N428);
xor XOR2 (N434, N433, N104);
or OR4 (N435, N429, N294, N201, N264);
nand NAND2 (N436, N422, N72);
xor XOR2 (N437, N425, N19);
nand NAND3 (N438, N434, N332, N322);
nand NAND3 (N439, N438, N210, N218);
and AND2 (N440, N432, N147);
nand NAND4 (N441, N436, N245, N422, N207);
xor XOR2 (N442, N435, N388);
not NOT1 (N443, N441);
or OR2 (N444, N420, N410);
or OR4 (N445, N431, N120, N425, N439);
not NOT1 (N446, N56);
buf BUF1 (N447, N445);
and AND2 (N448, N437, N193);
xor XOR2 (N449, N442, N272);
xor XOR2 (N450, N447, N284);
or OR3 (N451, N450, N183, N346);
nand NAND2 (N452, N443, N41);
and AND2 (N453, N440, N111);
nor NOR4 (N454, N452, N145, N332, N405);
nand NAND4 (N455, N448, N82, N53, N81);
buf BUF1 (N456, N396);
nand NAND4 (N457, N449, N225, N448, N16);
and AND2 (N458, N446, N331);
buf BUF1 (N459, N430);
not NOT1 (N460, N444);
not NOT1 (N461, N456);
xor XOR2 (N462, N458, N5);
and AND2 (N463, N453, N191);
nand NAND2 (N464, N460, N176);
not NOT1 (N465, N463);
and AND3 (N466, N464, N260, N185);
buf BUF1 (N467, N459);
nand NAND2 (N468, N467, N238);
nor NOR2 (N469, N468, N443);
xor XOR2 (N470, N451, N158);
xor XOR2 (N471, N457, N312);
buf BUF1 (N472, N469);
buf BUF1 (N473, N472);
nand NAND2 (N474, N473, N111);
xor XOR2 (N475, N454, N153);
xor XOR2 (N476, N462, N91);
xor XOR2 (N477, N474, N459);
not NOT1 (N478, N471);
xor XOR2 (N479, N470, N70);
nand NAND2 (N480, N465, N34);
xor XOR2 (N481, N480, N226);
and AND4 (N482, N466, N353, N93, N463);
nor NOR2 (N483, N461, N116);
buf BUF1 (N484, N426);
nor NOR2 (N485, N484, N307);
buf BUF1 (N486, N477);
xor XOR2 (N487, N475, N262);
xor XOR2 (N488, N455, N285);
xor XOR2 (N489, N486, N113);
not NOT1 (N490, N488);
nor NOR4 (N491, N479, N431, N447, N154);
buf BUF1 (N492, N482);
or OR3 (N493, N491, N23, N305);
or OR3 (N494, N483, N183, N462);
buf BUF1 (N495, N478);
nand NAND4 (N496, N481, N469, N219, N15);
nand NAND2 (N497, N489, N41);
and AND3 (N498, N487, N343, N288);
nor NOR3 (N499, N498, N339, N128);
or OR2 (N500, N496, N421);
not NOT1 (N501, N493);
nand NAND4 (N502, N495, N499, N71, N479);
xor XOR2 (N503, N118, N256);
not NOT1 (N504, N494);
nand NAND2 (N505, N490, N49);
and AND2 (N506, N476, N362);
and AND4 (N507, N503, N314, N21, N355);
xor XOR2 (N508, N506, N7);
nand NAND2 (N509, N508, N65);
xor XOR2 (N510, N502, N271);
nor NOR2 (N511, N501, N259);
buf BUF1 (N512, N509);
and AND3 (N513, N510, N387, N19);
and AND2 (N514, N504, N193);
xor XOR2 (N515, N511, N505);
not NOT1 (N516, N437);
xor XOR2 (N517, N513, N447);
xor XOR2 (N518, N515, N341);
not NOT1 (N519, N507);
or OR2 (N520, N518, N457);
or OR3 (N521, N517, N11, N103);
or OR3 (N522, N485, N154, N200);
xor XOR2 (N523, N492, N175);
nand NAND3 (N524, N512, N155, N364);
nand NAND2 (N525, N523, N233);
xor XOR2 (N526, N525, N318);
buf BUF1 (N527, N524);
nand NAND4 (N528, N500, N2, N453, N520);
or OR4 (N529, N122, N103, N454, N507);
not NOT1 (N530, N526);
xor XOR2 (N531, N529, N322);
buf BUF1 (N532, N530);
and AND4 (N533, N528, N287, N217, N33);
and AND4 (N534, N516, N90, N397, N526);
not NOT1 (N535, N531);
nand NAND2 (N536, N535, N158);
buf BUF1 (N537, N521);
buf BUF1 (N538, N527);
nand NAND2 (N539, N536, N127);
xor XOR2 (N540, N497, N120);
or OR4 (N541, N532, N346, N33, N178);
or OR4 (N542, N519, N206, N365, N495);
not NOT1 (N543, N534);
nor NOR2 (N544, N533, N441);
buf BUF1 (N545, N540);
nor NOR2 (N546, N542, N2);
and AND3 (N547, N546, N147, N426);
xor XOR2 (N548, N543, N7);
nor NOR2 (N549, N545, N119);
not NOT1 (N550, N538);
and AND2 (N551, N522, N58);
nor NOR4 (N552, N544, N79, N155, N266);
xor XOR2 (N553, N551, N454);
nand NAND2 (N554, N552, N277);
and AND2 (N555, N553, N237);
xor XOR2 (N556, N548, N392);
nor NOR2 (N557, N554, N515);
nor NOR4 (N558, N547, N239, N360, N383);
nand NAND2 (N559, N558, N330);
xor XOR2 (N560, N550, N190);
not NOT1 (N561, N557);
nand NAND2 (N562, N560, N555);
nor NOR3 (N563, N514, N481, N471);
or OR3 (N564, N68, N406, N512);
not NOT1 (N565, N556);
nand NAND3 (N566, N541, N391, N87);
nand NAND2 (N567, N565, N165);
and AND2 (N568, N564, N535);
nand NAND3 (N569, N562, N290, N62);
not NOT1 (N570, N549);
not NOT1 (N571, N568);
nand NAND3 (N572, N537, N227, N24);
nand NAND3 (N573, N566, N547, N47);
and AND3 (N574, N573, N296, N526);
nor NOR4 (N575, N572, N520, N285, N481);
and AND4 (N576, N571, N492, N501, N354);
xor XOR2 (N577, N539, N480);
not NOT1 (N578, N575);
buf BUF1 (N579, N563);
and AND4 (N580, N576, N62, N469, N273);
buf BUF1 (N581, N577);
and AND2 (N582, N569, N491);
nand NAND4 (N583, N559, N493, N47, N277);
xor XOR2 (N584, N578, N112);
xor XOR2 (N585, N567, N156);
nand NAND3 (N586, N580, N483, N374);
or OR2 (N587, N579, N344);
not NOT1 (N588, N585);
buf BUF1 (N589, N581);
or OR3 (N590, N584, N400, N311);
not NOT1 (N591, N589);
xor XOR2 (N592, N587, N241);
xor XOR2 (N593, N591, N572);
nand NAND3 (N594, N570, N159, N328);
nor NOR4 (N595, N590, N90, N236, N143);
not NOT1 (N596, N588);
xor XOR2 (N597, N595, N517);
nor NOR3 (N598, N593, N52, N86);
or OR2 (N599, N596, N3);
buf BUF1 (N600, N598);
and AND2 (N601, N599, N80);
buf BUF1 (N602, N586);
not NOT1 (N603, N597);
xor XOR2 (N604, N592, N562);
nand NAND2 (N605, N600, N87);
nand NAND2 (N606, N605, N421);
and AND3 (N607, N606, N66, N567);
or OR4 (N608, N607, N303, N42, N359);
nor NOR2 (N609, N602, N204);
and AND3 (N610, N601, N327, N603);
and AND2 (N611, N545, N455);
buf BUF1 (N612, N604);
or OR3 (N613, N582, N43, N237);
nor NOR4 (N614, N574, N475, N19, N136);
or OR2 (N615, N594, N239);
and AND4 (N616, N613, N615, N599, N229);
buf BUF1 (N617, N492);
not NOT1 (N618, N617);
xor XOR2 (N619, N618, N565);
xor XOR2 (N620, N619, N612);
and AND4 (N621, N74, N346, N569, N334);
buf BUF1 (N622, N620);
nand NAND3 (N623, N611, N494, N299);
not NOT1 (N624, N609);
and AND2 (N625, N608, N266);
or OR3 (N626, N610, N386, N393);
nor NOR2 (N627, N623, N120);
or OR3 (N628, N625, N291, N444);
xor XOR2 (N629, N622, N277);
nand NAND4 (N630, N614, N26, N117, N466);
and AND4 (N631, N628, N592, N534, N234);
and AND3 (N632, N631, N42, N631);
or OR2 (N633, N621, N22);
nand NAND4 (N634, N626, N20, N232, N49);
and AND4 (N635, N616, N381, N74, N569);
nor NOR3 (N636, N624, N370, N250);
xor XOR2 (N637, N632, N512);
xor XOR2 (N638, N636, N206);
xor XOR2 (N639, N638, N517);
or OR2 (N640, N627, N415);
nor NOR4 (N641, N583, N36, N294, N117);
buf BUF1 (N642, N634);
not NOT1 (N643, N629);
buf BUF1 (N644, N641);
nand NAND3 (N645, N637, N230, N386);
buf BUF1 (N646, N643);
xor XOR2 (N647, N633, N121);
nor NOR2 (N648, N640, N394);
or OR3 (N649, N639, N178, N419);
and AND2 (N650, N644, N594);
and AND4 (N651, N646, N350, N491, N197);
and AND4 (N652, N561, N161, N237, N453);
not NOT1 (N653, N648);
or OR3 (N654, N649, N285, N140);
nand NAND3 (N655, N650, N526, N284);
nand NAND2 (N656, N655, N297);
or OR3 (N657, N651, N214, N114);
or OR2 (N658, N635, N541);
nor NOR3 (N659, N658, N606, N110);
xor XOR2 (N660, N656, N638);
nand NAND3 (N661, N630, N420, N462);
or OR4 (N662, N642, N378, N41, N65);
nand NAND4 (N663, N657, N441, N354, N199);
or OR4 (N664, N645, N549, N472, N27);
nor NOR2 (N665, N654, N612);
and AND4 (N666, N660, N590, N80, N534);
and AND2 (N667, N659, N259);
or OR2 (N668, N664, N479);
not NOT1 (N669, N652);
or OR3 (N670, N647, N295, N363);
not NOT1 (N671, N667);
and AND4 (N672, N665, N406, N16, N34);
nand NAND3 (N673, N671, N41, N578);
not NOT1 (N674, N673);
nand NAND3 (N675, N661, N535, N99);
not NOT1 (N676, N672);
or OR3 (N677, N674, N291, N216);
not NOT1 (N678, N676);
nand NAND4 (N679, N663, N538, N24, N578);
nor NOR4 (N680, N669, N237, N171, N43);
xor XOR2 (N681, N662, N156);
buf BUF1 (N682, N668);
nor NOR2 (N683, N675, N589);
xor XOR2 (N684, N680, N19);
nor NOR3 (N685, N679, N338, N120);
not NOT1 (N686, N678);
nor NOR4 (N687, N686, N328, N679, N142);
nand NAND4 (N688, N666, N405, N179, N626);
or OR4 (N689, N683, N475, N100, N185);
or OR3 (N690, N684, N421, N83);
nor NOR2 (N691, N681, N213);
nand NAND4 (N692, N691, N576, N185, N89);
and AND4 (N693, N688, N33, N514, N448);
xor XOR2 (N694, N687, N331);
nand NAND2 (N695, N653, N671);
nand NAND4 (N696, N670, N180, N563, N190);
nand NAND4 (N697, N690, N354, N581, N9);
and AND2 (N698, N694, N90);
xor XOR2 (N699, N677, N427);
nand NAND2 (N700, N699, N669);
nor NOR3 (N701, N700, N146, N551);
or OR4 (N702, N693, N254, N635, N567);
nor NOR3 (N703, N698, N457, N131);
nand NAND3 (N704, N702, N543, N56);
buf BUF1 (N705, N697);
nand NAND3 (N706, N705, N601, N254);
or OR3 (N707, N704, N30, N133);
and AND3 (N708, N696, N544, N244);
nor NOR3 (N709, N689, N338, N575);
not NOT1 (N710, N685);
xor XOR2 (N711, N709, N491);
xor XOR2 (N712, N711, N592);
buf BUF1 (N713, N706);
nor NOR4 (N714, N710, N528, N440, N430);
buf BUF1 (N715, N695);
nor NOR3 (N716, N703, N555, N577);
or OR4 (N717, N701, N452, N547, N54);
nand NAND3 (N718, N717, N668, N516);
buf BUF1 (N719, N718);
and AND3 (N720, N708, N585, N283);
nor NOR2 (N721, N713, N77);
xor XOR2 (N722, N715, N12);
or OR4 (N723, N722, N6, N517, N334);
and AND4 (N724, N721, N203, N629, N686);
nand NAND3 (N725, N723, N651, N451);
and AND4 (N726, N707, N170, N120, N4);
nand NAND2 (N727, N692, N331);
not NOT1 (N728, N682);
and AND2 (N729, N724, N202);
and AND2 (N730, N714, N188);
not NOT1 (N731, N712);
nand NAND4 (N732, N726, N704, N99, N453);
nand NAND2 (N733, N720, N284);
not NOT1 (N734, N731);
nor NOR3 (N735, N725, N506, N371);
and AND2 (N736, N734, N489);
not NOT1 (N737, N730);
nand NAND3 (N738, N716, N459, N257);
not NOT1 (N739, N719);
or OR2 (N740, N736, N286);
not NOT1 (N741, N738);
nor NOR2 (N742, N728, N428);
xor XOR2 (N743, N742, N678);
nor NOR2 (N744, N729, N413);
nand NAND4 (N745, N740, N156, N29, N579);
nand NAND4 (N746, N739, N165, N381, N318);
or OR4 (N747, N727, N258, N584, N279);
or OR4 (N748, N743, N218, N405, N439);
nand NAND4 (N749, N733, N693, N60, N530);
not NOT1 (N750, N745);
xor XOR2 (N751, N735, N40);
and AND4 (N752, N744, N474, N326, N363);
nor NOR4 (N753, N748, N680, N380, N516);
xor XOR2 (N754, N751, N467);
and AND4 (N755, N747, N129, N699, N654);
nor NOR3 (N756, N750, N437, N593);
and AND3 (N757, N737, N366, N517);
and AND4 (N758, N753, N716, N594, N308);
xor XOR2 (N759, N741, N349);
nand NAND3 (N760, N752, N261, N491);
nor NOR2 (N761, N758, N708);
not NOT1 (N762, N754);
nand NAND3 (N763, N732, N285, N434);
xor XOR2 (N764, N762, N698);
buf BUF1 (N765, N763);
buf BUF1 (N766, N764);
not NOT1 (N767, N761);
nor NOR4 (N768, N759, N227, N265, N245);
or OR3 (N769, N746, N223, N320);
buf BUF1 (N770, N767);
nor NOR3 (N771, N770, N543, N264);
buf BUF1 (N772, N755);
and AND2 (N773, N768, N284);
or OR4 (N774, N756, N281, N26, N381);
and AND4 (N775, N757, N279, N591, N223);
nand NAND2 (N776, N773, N736);
nor NOR2 (N777, N769, N259);
nand NAND3 (N778, N760, N102, N599);
and AND3 (N779, N766, N82, N288);
buf BUF1 (N780, N779);
or OR4 (N781, N777, N276, N373, N767);
xor XOR2 (N782, N775, N764);
and AND4 (N783, N776, N349, N547, N518);
and AND2 (N784, N765, N537);
nor NOR2 (N785, N778, N50);
or OR4 (N786, N749, N22, N221, N636);
or OR2 (N787, N772, N42);
or OR3 (N788, N786, N451, N494);
nor NOR3 (N789, N781, N548, N179);
nor NOR4 (N790, N785, N138, N251, N747);
xor XOR2 (N791, N774, N458);
or OR3 (N792, N787, N234, N491);
not NOT1 (N793, N771);
nand NAND4 (N794, N792, N300, N314, N493);
xor XOR2 (N795, N789, N594);
buf BUF1 (N796, N794);
nand NAND3 (N797, N790, N223, N782);
or OR4 (N798, N194, N295, N683, N44);
buf BUF1 (N799, N795);
nor NOR2 (N800, N793, N28);
not NOT1 (N801, N788);
and AND4 (N802, N784, N721, N119, N419);
xor XOR2 (N803, N798, N363);
xor XOR2 (N804, N791, N717);
buf BUF1 (N805, N796);
buf BUF1 (N806, N802);
and AND2 (N807, N804, N218);
not NOT1 (N808, N807);
nand NAND2 (N809, N800, N368);
and AND2 (N810, N808, N420);
nand NAND4 (N811, N780, N479, N195, N710);
xor XOR2 (N812, N783, N394);
or OR2 (N813, N805, N614);
xor XOR2 (N814, N810, N313);
not NOT1 (N815, N797);
not NOT1 (N816, N814);
buf BUF1 (N817, N813);
not NOT1 (N818, N806);
and AND3 (N819, N799, N426, N410);
not NOT1 (N820, N818);
xor XOR2 (N821, N809, N70);
or OR2 (N822, N820, N349);
buf BUF1 (N823, N821);
xor XOR2 (N824, N817, N325);
buf BUF1 (N825, N824);
not NOT1 (N826, N816);
or OR4 (N827, N811, N319, N71, N358);
not NOT1 (N828, N823);
buf BUF1 (N829, N828);
nand NAND4 (N830, N827, N724, N53, N224);
nand NAND4 (N831, N825, N784, N344, N28);
not NOT1 (N832, N812);
nor NOR4 (N833, N801, N619, N442, N706);
nor NOR2 (N834, N822, N695);
not NOT1 (N835, N829);
or OR2 (N836, N830, N210);
nor NOR4 (N837, N834, N218, N616, N343);
buf BUF1 (N838, N819);
not NOT1 (N839, N826);
nand NAND2 (N840, N837, N668);
not NOT1 (N841, N836);
nor NOR2 (N842, N832, N307);
not NOT1 (N843, N840);
nand NAND3 (N844, N803, N446, N189);
and AND3 (N845, N835, N585, N527);
buf BUF1 (N846, N839);
nor NOR4 (N847, N838, N715, N831, N717);
or OR4 (N848, N456, N385, N606, N321);
nor NOR2 (N849, N845, N16);
xor XOR2 (N850, N847, N85);
not NOT1 (N851, N850);
buf BUF1 (N852, N815);
nand NAND4 (N853, N844, N591, N752, N91);
not NOT1 (N854, N848);
and AND4 (N855, N849, N39, N505, N260);
buf BUF1 (N856, N852);
xor XOR2 (N857, N853, N658);
nor NOR3 (N858, N843, N321, N451);
or OR4 (N859, N851, N611, N568, N664);
nand NAND2 (N860, N856, N88);
not NOT1 (N861, N833);
nor NOR2 (N862, N859, N201);
xor XOR2 (N863, N846, N118);
nor NOR4 (N864, N842, N153, N618, N349);
nand NAND3 (N865, N864, N630, N538);
or OR4 (N866, N858, N417, N355, N714);
not NOT1 (N867, N855);
nand NAND3 (N868, N857, N100, N406);
nor NOR2 (N869, N868, N260);
not NOT1 (N870, N861);
nand NAND4 (N871, N870, N828, N777, N359);
nand NAND4 (N872, N869, N501, N620, N511);
or OR2 (N873, N863, N177);
not NOT1 (N874, N862);
buf BUF1 (N875, N872);
and AND4 (N876, N871, N426, N662, N451);
or OR2 (N877, N873, N196);
buf BUF1 (N878, N865);
not NOT1 (N879, N878);
nor NOR4 (N880, N875, N133, N6, N428);
and AND2 (N881, N866, N425);
and AND2 (N882, N867, N473);
xor XOR2 (N883, N876, N401);
not NOT1 (N884, N854);
nand NAND2 (N885, N874, N462);
not NOT1 (N886, N885);
or OR3 (N887, N860, N400, N805);
or OR3 (N888, N877, N748, N527);
xor XOR2 (N889, N881, N427);
or OR4 (N890, N883, N678, N165, N801);
or OR4 (N891, N884, N887, N411, N633);
not NOT1 (N892, N664);
not NOT1 (N893, N841);
buf BUF1 (N894, N892);
xor XOR2 (N895, N879, N86);
not NOT1 (N896, N888);
nor NOR4 (N897, N882, N24, N113, N729);
nand NAND3 (N898, N895, N729, N342);
not NOT1 (N899, N894);
xor XOR2 (N900, N898, N274);
and AND2 (N901, N896, N495);
xor XOR2 (N902, N890, N244);
not NOT1 (N903, N889);
xor XOR2 (N904, N901, N737);
nand NAND4 (N905, N886, N595, N141, N501);
nor NOR2 (N906, N902, N304);
not NOT1 (N907, N880);
xor XOR2 (N908, N906, N375);
or OR3 (N909, N900, N845, N44);
buf BUF1 (N910, N905);
not NOT1 (N911, N904);
not NOT1 (N912, N909);
xor XOR2 (N913, N908, N342);
and AND3 (N914, N907, N335, N861);
not NOT1 (N915, N910);
and AND2 (N916, N903, N491);
nand NAND2 (N917, N899, N315);
xor XOR2 (N918, N893, N376);
nand NAND2 (N919, N911, N124);
xor XOR2 (N920, N919, N78);
nand NAND2 (N921, N897, N346);
and AND3 (N922, N918, N544, N611);
or OR2 (N923, N922, N615);
nor NOR3 (N924, N923, N135, N761);
nor NOR2 (N925, N924, N188);
and AND3 (N926, N921, N350, N212);
not NOT1 (N927, N916);
xor XOR2 (N928, N925, N743);
or OR4 (N929, N927, N277, N457, N354);
buf BUF1 (N930, N920);
xor XOR2 (N931, N913, N551);
and AND4 (N932, N912, N454, N733, N695);
nor NOR4 (N933, N928, N500, N894, N921);
not NOT1 (N934, N932);
xor XOR2 (N935, N931, N306);
xor XOR2 (N936, N933, N169);
nor NOR2 (N937, N936, N396);
xor XOR2 (N938, N937, N731);
nand NAND3 (N939, N929, N193, N235);
not NOT1 (N940, N914);
buf BUF1 (N941, N940);
nor NOR3 (N942, N917, N880, N854);
not NOT1 (N943, N941);
and AND4 (N944, N935, N504, N672, N363);
xor XOR2 (N945, N939, N166);
nand NAND4 (N946, N926, N308, N107, N332);
buf BUF1 (N947, N930);
buf BUF1 (N948, N891);
not NOT1 (N949, N915);
or OR2 (N950, N938, N921);
buf BUF1 (N951, N950);
not NOT1 (N952, N949);
buf BUF1 (N953, N948);
nor NOR4 (N954, N947, N196, N894, N384);
not NOT1 (N955, N945);
and AND4 (N956, N955, N575, N415, N646);
nor NOR2 (N957, N952, N51);
buf BUF1 (N958, N957);
xor XOR2 (N959, N954, N157);
buf BUF1 (N960, N934);
and AND4 (N961, N944, N491, N394, N951);
and AND4 (N962, N146, N808, N664, N523);
nor NOR3 (N963, N943, N504, N232);
or OR3 (N964, N946, N444, N282);
not NOT1 (N965, N953);
nand NAND2 (N966, N959, N236);
and AND3 (N967, N942, N132, N395);
not NOT1 (N968, N963);
nor NOR4 (N969, N961, N837, N811, N499);
not NOT1 (N970, N965);
nand NAND3 (N971, N958, N14, N272);
or OR4 (N972, N962, N599, N646, N615);
buf BUF1 (N973, N967);
nand NAND4 (N974, N966, N764, N154, N290);
xor XOR2 (N975, N970, N496);
nor NOR3 (N976, N971, N643, N768);
or OR2 (N977, N964, N971);
nand NAND4 (N978, N976, N686, N619, N380);
or OR4 (N979, N978, N323, N719, N421);
and AND2 (N980, N972, N381);
buf BUF1 (N981, N968);
buf BUF1 (N982, N975);
xor XOR2 (N983, N960, N664);
nor NOR3 (N984, N979, N83, N781);
buf BUF1 (N985, N969);
and AND2 (N986, N981, N967);
nor NOR2 (N987, N974, N486);
not NOT1 (N988, N987);
buf BUF1 (N989, N956);
nand NAND4 (N990, N983, N5, N929, N625);
or OR2 (N991, N973, N695);
and AND4 (N992, N982, N367, N105, N429);
nor NOR2 (N993, N980, N522);
buf BUF1 (N994, N993);
xor XOR2 (N995, N988, N146);
nand NAND4 (N996, N990, N287, N574, N125);
or OR3 (N997, N992, N302, N845);
not NOT1 (N998, N977);
xor XOR2 (N999, N996, N6);
or OR2 (N1000, N994, N685);
not NOT1 (N1001, N991);
and AND4 (N1002, N985, N213, N521, N216);
nand NAND2 (N1003, N1000, N797);
nand NAND3 (N1004, N1002, N649, N483);
nand NAND2 (N1005, N1004, N42);
nand NAND3 (N1006, N986, N14, N181);
nand NAND4 (N1007, N998, N256, N6, N944);
not NOT1 (N1008, N999);
buf BUF1 (N1009, N1008);
buf BUF1 (N1010, N989);
xor XOR2 (N1011, N1006, N306);
or OR2 (N1012, N1005, N956);
or OR3 (N1013, N1007, N436, N92);
not NOT1 (N1014, N1001);
xor XOR2 (N1015, N1009, N907);
buf BUF1 (N1016, N1015);
xor XOR2 (N1017, N997, N539);
not NOT1 (N1018, N995);
and AND4 (N1019, N1003, N205, N364, N978);
and AND4 (N1020, N1017, N948, N327, N916);
xor XOR2 (N1021, N1013, N513);
or OR3 (N1022, N984, N654, N408);
buf BUF1 (N1023, N1022);
and AND3 (N1024, N1012, N491, N366);
and AND3 (N1025, N1010, N471, N810);
buf BUF1 (N1026, N1019);
buf BUF1 (N1027, N1024);
buf BUF1 (N1028, N1011);
nor NOR4 (N1029, N1025, N614, N882, N833);
buf BUF1 (N1030, N1027);
nand NAND4 (N1031, N1030, N335, N651, N465);
nor NOR3 (N1032, N1014, N810, N228);
xor XOR2 (N1033, N1018, N396);
nand NAND4 (N1034, N1016, N681, N280, N576);
not NOT1 (N1035, N1034);
not NOT1 (N1036, N1023);
and AND4 (N1037, N1029, N943, N195, N785);
xor XOR2 (N1038, N1037, N537);
and AND3 (N1039, N1031, N681, N289);
and AND4 (N1040, N1026, N821, N692, N573);
not NOT1 (N1041, N1040);
not NOT1 (N1042, N1035);
buf BUF1 (N1043, N1036);
buf BUF1 (N1044, N1041);
not NOT1 (N1045, N1043);
buf BUF1 (N1046, N1020);
and AND2 (N1047, N1042, N438);
not NOT1 (N1048, N1039);
and AND3 (N1049, N1021, N119, N483);
or OR4 (N1050, N1046, N869, N673, N447);
nor NOR2 (N1051, N1045, N59);
not NOT1 (N1052, N1051);
or OR2 (N1053, N1047, N406);
nand NAND4 (N1054, N1033, N426, N789, N72);
or OR2 (N1055, N1054, N578);
nor NOR3 (N1056, N1055, N271, N952);
and AND3 (N1057, N1038, N111, N243);
buf BUF1 (N1058, N1049);
and AND2 (N1059, N1053, N612);
xor XOR2 (N1060, N1050, N105);
nor NOR4 (N1061, N1056, N890, N206, N327);
and AND2 (N1062, N1058, N448);
or OR4 (N1063, N1057, N964, N1018, N778);
and AND2 (N1064, N1044, N391);
nor NOR2 (N1065, N1063, N971);
buf BUF1 (N1066, N1048);
or OR2 (N1067, N1059, N615);
not NOT1 (N1068, N1065);
nor NOR2 (N1069, N1028, N558);
nand NAND3 (N1070, N1068, N758, N227);
xor XOR2 (N1071, N1062, N11);
nor NOR2 (N1072, N1060, N1007);
nand NAND4 (N1073, N1032, N120, N651, N950);
and AND2 (N1074, N1052, N566);
or OR4 (N1075, N1069, N490, N317, N894);
not NOT1 (N1076, N1075);
and AND4 (N1077, N1072, N104, N433, N93);
not NOT1 (N1078, N1071);
nor NOR3 (N1079, N1077, N185, N77);
nor NOR2 (N1080, N1070, N24);
xor XOR2 (N1081, N1064, N14);
and AND3 (N1082, N1074, N586, N682);
not NOT1 (N1083, N1079);
nand NAND2 (N1084, N1073, N925);
nor NOR4 (N1085, N1067, N744, N798, N156);
nand NAND3 (N1086, N1076, N399, N419);
nor NOR3 (N1087, N1066, N402, N404);
buf BUF1 (N1088, N1085);
buf BUF1 (N1089, N1088);
not NOT1 (N1090, N1081);
nor NOR3 (N1091, N1090, N61, N1033);
not NOT1 (N1092, N1078);
nor NOR2 (N1093, N1091, N443);
xor XOR2 (N1094, N1086, N230);
buf BUF1 (N1095, N1093);
not NOT1 (N1096, N1080);
and AND2 (N1097, N1082, N119);
not NOT1 (N1098, N1083);
and AND3 (N1099, N1097, N979, N994);
or OR2 (N1100, N1099, N1044);
xor XOR2 (N1101, N1087, N167);
nand NAND3 (N1102, N1095, N93, N245);
or OR2 (N1103, N1096, N711);
not NOT1 (N1104, N1103);
nor NOR2 (N1105, N1101, N433);
and AND4 (N1106, N1092, N794, N660, N35);
or OR4 (N1107, N1100, N1010, N802, N358);
buf BUF1 (N1108, N1098);
and AND4 (N1109, N1105, N814, N687, N622);
nor NOR3 (N1110, N1106, N499, N504);
not NOT1 (N1111, N1109);
or OR4 (N1112, N1108, N849, N387, N879);
buf BUF1 (N1113, N1089);
not NOT1 (N1114, N1094);
nor NOR4 (N1115, N1061, N789, N1080, N202);
nand NAND3 (N1116, N1115, N490, N576);
nor NOR4 (N1117, N1084, N1016, N464, N277);
nand NAND2 (N1118, N1116, N233);
or OR2 (N1119, N1102, N785);
not NOT1 (N1120, N1112);
buf BUF1 (N1121, N1104);
or OR3 (N1122, N1121, N581, N907);
buf BUF1 (N1123, N1111);
not NOT1 (N1124, N1113);
nor NOR2 (N1125, N1119, N1112);
nand NAND4 (N1126, N1125, N87, N111, N457);
nor NOR4 (N1127, N1107, N427, N854, N594);
xor XOR2 (N1128, N1120, N935);
not NOT1 (N1129, N1118);
and AND3 (N1130, N1129, N422, N222);
not NOT1 (N1131, N1117);
nor NOR4 (N1132, N1122, N150, N342, N782);
nand NAND2 (N1133, N1126, N871);
not NOT1 (N1134, N1114);
and AND3 (N1135, N1110, N978, N1072);
buf BUF1 (N1136, N1127);
and AND3 (N1137, N1132, N843, N181);
or OR2 (N1138, N1134, N1105);
nor NOR2 (N1139, N1130, N783);
or OR2 (N1140, N1138, N399);
nor NOR2 (N1141, N1128, N308);
not NOT1 (N1142, N1137);
not NOT1 (N1143, N1141);
xor XOR2 (N1144, N1143, N417);
nand NAND3 (N1145, N1123, N956, N373);
buf BUF1 (N1146, N1131);
nor NOR2 (N1147, N1124, N848);
or OR3 (N1148, N1135, N18, N642);
buf BUF1 (N1149, N1144);
and AND4 (N1150, N1133, N478, N720, N77);
buf BUF1 (N1151, N1148);
or OR2 (N1152, N1145, N594);
nor NOR2 (N1153, N1147, N819);
not NOT1 (N1154, N1142);
nand NAND3 (N1155, N1136, N238, N846);
nand NAND3 (N1156, N1155, N870, N534);
xor XOR2 (N1157, N1152, N268);
buf BUF1 (N1158, N1146);
and AND3 (N1159, N1150, N129, N442);
buf BUF1 (N1160, N1153);
nor NOR2 (N1161, N1151, N976);
and AND3 (N1162, N1158, N1009, N1147);
nor NOR3 (N1163, N1140, N494, N565);
and AND3 (N1164, N1156, N401, N1054);
nor NOR4 (N1165, N1164, N968, N6, N1022);
nor NOR4 (N1166, N1157, N754, N230, N73);
not NOT1 (N1167, N1139);
or OR4 (N1168, N1162, N912, N326, N658);
or OR4 (N1169, N1167, N174, N889, N515);
not NOT1 (N1170, N1154);
not NOT1 (N1171, N1169);
xor XOR2 (N1172, N1160, N1131);
xor XOR2 (N1173, N1163, N1123);
or OR2 (N1174, N1149, N1083);
nand NAND2 (N1175, N1159, N36);
xor XOR2 (N1176, N1172, N520);
xor XOR2 (N1177, N1173, N739);
xor XOR2 (N1178, N1165, N681);
or OR2 (N1179, N1177, N180);
xor XOR2 (N1180, N1176, N920);
buf BUF1 (N1181, N1170);
buf BUF1 (N1182, N1175);
nand NAND2 (N1183, N1181, N299);
nor NOR2 (N1184, N1182, N385);
buf BUF1 (N1185, N1166);
or OR3 (N1186, N1171, N81, N1126);
and AND4 (N1187, N1161, N100, N930, N294);
and AND2 (N1188, N1168, N74);
not NOT1 (N1189, N1178);
or OR2 (N1190, N1189, N1161);
xor XOR2 (N1191, N1183, N768);
and AND2 (N1192, N1184, N1036);
xor XOR2 (N1193, N1188, N971);
nand NAND2 (N1194, N1193, N540);
and AND2 (N1195, N1179, N544);
buf BUF1 (N1196, N1186);
xor XOR2 (N1197, N1187, N8);
xor XOR2 (N1198, N1180, N583);
nor NOR4 (N1199, N1174, N757, N377, N1033);
and AND4 (N1200, N1190, N104, N852, N159);
nand NAND4 (N1201, N1191, N910, N1003, N253);
or OR4 (N1202, N1197, N46, N723, N981);
buf BUF1 (N1203, N1200);
and AND3 (N1204, N1198, N465, N738);
or OR3 (N1205, N1203, N671, N363);
buf BUF1 (N1206, N1194);
or OR4 (N1207, N1199, N381, N928, N1141);
nor NOR4 (N1208, N1207, N128, N1135, N412);
or OR2 (N1209, N1202, N114);
not NOT1 (N1210, N1195);
or OR2 (N1211, N1210, N778);
or OR2 (N1212, N1196, N369);
or OR4 (N1213, N1206, N528, N994, N257);
nand NAND2 (N1214, N1185, N579);
and AND3 (N1215, N1212, N285, N1159);
or OR3 (N1216, N1208, N169, N72);
xor XOR2 (N1217, N1214, N369);
buf BUF1 (N1218, N1215);
xor XOR2 (N1219, N1217, N643);
or OR2 (N1220, N1213, N1054);
xor XOR2 (N1221, N1205, N1121);
nor NOR4 (N1222, N1204, N827, N637, N870);
buf BUF1 (N1223, N1221);
and AND4 (N1224, N1201, N734, N560, N138);
xor XOR2 (N1225, N1218, N197);
buf BUF1 (N1226, N1192);
buf BUF1 (N1227, N1223);
nand NAND4 (N1228, N1216, N1226, N922, N205);
xor XOR2 (N1229, N387, N9);
and AND3 (N1230, N1222, N914, N771);
or OR3 (N1231, N1227, N825, N722);
or OR3 (N1232, N1229, N531, N582);
or OR2 (N1233, N1209, N1164);
nor NOR2 (N1234, N1225, N1092);
and AND2 (N1235, N1219, N831);
not NOT1 (N1236, N1230);
buf BUF1 (N1237, N1224);
nor NOR2 (N1238, N1231, N873);
and AND3 (N1239, N1238, N1176, N1128);
nor NOR2 (N1240, N1234, N608);
nor NOR3 (N1241, N1239, N290, N316);
nor NOR2 (N1242, N1235, N537);
not NOT1 (N1243, N1236);
or OR3 (N1244, N1241, N511, N1148);
and AND2 (N1245, N1228, N192);
or OR3 (N1246, N1232, N569, N736);
or OR4 (N1247, N1220, N136, N947, N234);
and AND3 (N1248, N1211, N552, N590);
nor NOR4 (N1249, N1243, N502, N652, N953);
nand NAND4 (N1250, N1248, N1220, N797, N672);
buf BUF1 (N1251, N1244);
and AND2 (N1252, N1251, N759);
and AND4 (N1253, N1247, N381, N403, N31);
nor NOR2 (N1254, N1237, N1252);
xor XOR2 (N1255, N682, N1140);
or OR4 (N1256, N1253, N330, N622, N202);
nor NOR3 (N1257, N1254, N1235, N574);
or OR2 (N1258, N1233, N452);
nand NAND3 (N1259, N1258, N498, N853);
or OR4 (N1260, N1246, N658, N313, N545);
nand NAND2 (N1261, N1257, N773);
nand NAND4 (N1262, N1259, N203, N194, N556);
or OR4 (N1263, N1250, N817, N289, N583);
or OR4 (N1264, N1249, N271, N434, N187);
not NOT1 (N1265, N1260);
or OR2 (N1266, N1255, N345);
nor NOR4 (N1267, N1242, N89, N649, N86);
not NOT1 (N1268, N1265);
nor NOR2 (N1269, N1240, N1089);
xor XOR2 (N1270, N1263, N285);
xor XOR2 (N1271, N1261, N799);
or OR4 (N1272, N1264, N202, N279, N656);
nand NAND2 (N1273, N1272, N1144);
not NOT1 (N1274, N1256);
not NOT1 (N1275, N1262);
nand NAND3 (N1276, N1271, N10, N1173);
not NOT1 (N1277, N1269);
or OR4 (N1278, N1275, N740, N907, N934);
buf BUF1 (N1279, N1267);
nor NOR4 (N1280, N1278, N306, N893, N499);
xor XOR2 (N1281, N1270, N947);
xor XOR2 (N1282, N1276, N1256);
not NOT1 (N1283, N1245);
buf BUF1 (N1284, N1281);
nand NAND2 (N1285, N1277, N1212);
or OR2 (N1286, N1273, N482);
xor XOR2 (N1287, N1268, N1144);
and AND4 (N1288, N1287, N1074, N154, N759);
xor XOR2 (N1289, N1288, N828);
nand NAND4 (N1290, N1284, N2, N78, N1088);
nor NOR2 (N1291, N1266, N170);
nor NOR4 (N1292, N1280, N43, N989, N805);
xor XOR2 (N1293, N1289, N879);
and AND4 (N1294, N1279, N388, N1061, N979);
buf BUF1 (N1295, N1282);
buf BUF1 (N1296, N1293);
nand NAND3 (N1297, N1283, N1198, N80);
buf BUF1 (N1298, N1296);
and AND3 (N1299, N1298, N1186, N493);
and AND2 (N1300, N1286, N767);
nand NAND4 (N1301, N1274, N711, N405, N784);
not NOT1 (N1302, N1300);
nor NOR3 (N1303, N1290, N177, N954);
buf BUF1 (N1304, N1294);
buf BUF1 (N1305, N1304);
xor XOR2 (N1306, N1303, N722);
and AND4 (N1307, N1291, N221, N129, N893);
nand NAND4 (N1308, N1306, N1189, N1303, N570);
buf BUF1 (N1309, N1292);
nand NAND4 (N1310, N1302, N114, N622, N98);
and AND4 (N1311, N1295, N34, N25, N526);
nor NOR2 (N1312, N1309, N969);
xor XOR2 (N1313, N1310, N277);
xor XOR2 (N1314, N1307, N61);
nor NOR2 (N1315, N1311, N489);
or OR3 (N1316, N1312, N931, N763);
not NOT1 (N1317, N1316);
or OR2 (N1318, N1299, N170);
or OR4 (N1319, N1315, N293, N575, N708);
nand NAND3 (N1320, N1314, N113, N901);
or OR2 (N1321, N1318, N108);
nor NOR3 (N1322, N1285, N611, N414);
xor XOR2 (N1323, N1301, N335);
nand NAND4 (N1324, N1313, N1128, N454, N1204);
nand NAND2 (N1325, N1320, N205);
nor NOR2 (N1326, N1325, N47);
or OR4 (N1327, N1305, N1297, N885, N53);
not NOT1 (N1328, N1122);
or OR3 (N1329, N1317, N689, N545);
xor XOR2 (N1330, N1326, N321);
xor XOR2 (N1331, N1308, N1181);
buf BUF1 (N1332, N1331);
buf BUF1 (N1333, N1327);
and AND4 (N1334, N1329, N990, N1043, N588);
or OR2 (N1335, N1319, N805);
xor XOR2 (N1336, N1321, N1181);
or OR3 (N1337, N1336, N922, N61);
or OR2 (N1338, N1323, N210);
buf BUF1 (N1339, N1328);
nand NAND4 (N1340, N1322, N1112, N172, N261);
nor NOR4 (N1341, N1332, N239, N104, N1048);
not NOT1 (N1342, N1330);
and AND4 (N1343, N1324, N845, N122, N1290);
or OR4 (N1344, N1341, N460, N958, N61);
nand NAND3 (N1345, N1338, N1230, N1032);
xor XOR2 (N1346, N1337, N1262);
and AND2 (N1347, N1334, N710);
buf BUF1 (N1348, N1333);
or OR3 (N1349, N1348, N759, N709);
xor XOR2 (N1350, N1339, N394);
nor NOR4 (N1351, N1347, N395, N615, N864);
or OR3 (N1352, N1343, N177, N222);
xor XOR2 (N1353, N1350, N951);
xor XOR2 (N1354, N1344, N60);
xor XOR2 (N1355, N1351, N211);
and AND4 (N1356, N1346, N1188, N3, N789);
and AND4 (N1357, N1354, N715, N28, N1125);
or OR4 (N1358, N1345, N914, N709, N321);
buf BUF1 (N1359, N1355);
nor NOR3 (N1360, N1356, N352, N1113);
not NOT1 (N1361, N1352);
buf BUF1 (N1362, N1340);
buf BUF1 (N1363, N1358);
nor NOR2 (N1364, N1363, N177);
or OR3 (N1365, N1361, N1342, N604);
nor NOR4 (N1366, N245, N950, N1266, N207);
nand NAND4 (N1367, N1357, N1279, N68, N913);
xor XOR2 (N1368, N1367, N627);
buf BUF1 (N1369, N1335);
nor NOR3 (N1370, N1360, N586, N532);
and AND3 (N1371, N1349, N1078, N125);
buf BUF1 (N1372, N1371);
xor XOR2 (N1373, N1364, N926);
nor NOR4 (N1374, N1359, N867, N1165, N798);
xor XOR2 (N1375, N1362, N218);
xor XOR2 (N1376, N1368, N147);
xor XOR2 (N1377, N1373, N872);
not NOT1 (N1378, N1365);
xor XOR2 (N1379, N1353, N48);
or OR3 (N1380, N1366, N1334, N210);
buf BUF1 (N1381, N1375);
not NOT1 (N1382, N1377);
not NOT1 (N1383, N1381);
nand NAND3 (N1384, N1372, N1093, N435);
and AND3 (N1385, N1382, N650, N1217);
nor NOR2 (N1386, N1383, N1262);
buf BUF1 (N1387, N1376);
nand NAND4 (N1388, N1370, N958, N153, N970);
nand NAND3 (N1389, N1379, N1282, N524);
buf BUF1 (N1390, N1385);
nand NAND3 (N1391, N1388, N1284, N1066);
not NOT1 (N1392, N1391);
not NOT1 (N1393, N1384);
or OR4 (N1394, N1393, N916, N217, N978);
buf BUF1 (N1395, N1374);
buf BUF1 (N1396, N1387);
or OR4 (N1397, N1380, N302, N969, N541);
nor NOR2 (N1398, N1395, N1189);
or OR4 (N1399, N1390, N1328, N887, N441);
or OR3 (N1400, N1397, N378, N338);
xor XOR2 (N1401, N1386, N404);
buf BUF1 (N1402, N1389);
nor NOR3 (N1403, N1394, N1097, N1195);
and AND2 (N1404, N1396, N1238);
not NOT1 (N1405, N1369);
and AND3 (N1406, N1403, N1296, N1096);
xor XOR2 (N1407, N1398, N1309);
buf BUF1 (N1408, N1402);
xor XOR2 (N1409, N1400, N1028);
nand NAND4 (N1410, N1404, N1045, N689, N1274);
and AND3 (N1411, N1405, N861, N1157);
or OR3 (N1412, N1409, N1237, N1228);
and AND4 (N1413, N1378, N394, N647, N135);
buf BUF1 (N1414, N1407);
xor XOR2 (N1415, N1412, N701);
buf BUF1 (N1416, N1413);
nand NAND4 (N1417, N1401, N687, N246, N158);
xor XOR2 (N1418, N1406, N455);
or OR3 (N1419, N1417, N955, N453);
and AND2 (N1420, N1392, N84);
nand NAND4 (N1421, N1410, N1195, N1086, N1383);
not NOT1 (N1422, N1408);
nor NOR4 (N1423, N1422, N19, N394, N612);
nand NAND2 (N1424, N1416, N252);
xor XOR2 (N1425, N1414, N188);
buf BUF1 (N1426, N1418);
not NOT1 (N1427, N1419);
nand NAND3 (N1428, N1427, N81, N471);
not NOT1 (N1429, N1420);
or OR4 (N1430, N1428, N169, N1083, N567);
or OR3 (N1431, N1426, N843, N491);
nand NAND3 (N1432, N1425, N949, N763);
and AND2 (N1433, N1421, N1051);
nand NAND3 (N1434, N1432, N431, N488);
and AND3 (N1435, N1430, N887, N109);
xor XOR2 (N1436, N1415, N612);
nand NAND4 (N1437, N1423, N755, N1338, N920);
xor XOR2 (N1438, N1434, N480);
not NOT1 (N1439, N1424);
and AND2 (N1440, N1433, N334);
buf BUF1 (N1441, N1435);
and AND4 (N1442, N1431, N80, N397, N677);
xor XOR2 (N1443, N1441, N992);
nand NAND2 (N1444, N1436, N875);
or OR2 (N1445, N1440, N889);
and AND2 (N1446, N1429, N78);
nand NAND3 (N1447, N1399, N609, N1316);
nand NAND4 (N1448, N1438, N211, N570, N101);
or OR3 (N1449, N1411, N171, N609);
nand NAND2 (N1450, N1442, N254);
buf BUF1 (N1451, N1444);
nand NAND3 (N1452, N1445, N434, N548);
nand NAND3 (N1453, N1452, N455, N1386);
and AND2 (N1454, N1439, N1313);
buf BUF1 (N1455, N1451);
not NOT1 (N1456, N1446);
and AND4 (N1457, N1455, N162, N2, N825);
not NOT1 (N1458, N1437);
and AND3 (N1459, N1454, N1109, N637);
buf BUF1 (N1460, N1449);
nand NAND4 (N1461, N1460, N473, N1124, N978);
nand NAND3 (N1462, N1458, N1146, N693);
and AND2 (N1463, N1459, N495);
buf BUF1 (N1464, N1462);
not NOT1 (N1465, N1463);
not NOT1 (N1466, N1465);
buf BUF1 (N1467, N1457);
buf BUF1 (N1468, N1461);
nor NOR2 (N1469, N1443, N621);
buf BUF1 (N1470, N1468);
or OR2 (N1471, N1448, N607);
and AND3 (N1472, N1447, N226, N1338);
xor XOR2 (N1473, N1472, N867);
and AND2 (N1474, N1453, N138);
xor XOR2 (N1475, N1473, N1247);
nand NAND3 (N1476, N1466, N403, N997);
not NOT1 (N1477, N1471);
buf BUF1 (N1478, N1450);
and AND3 (N1479, N1467, N1355, N905);
xor XOR2 (N1480, N1469, N486);
nor NOR3 (N1481, N1478, N1133, N647);
nor NOR4 (N1482, N1479, N478, N716, N354);
xor XOR2 (N1483, N1475, N1174);
and AND4 (N1484, N1476, N818, N960, N32);
nor NOR2 (N1485, N1470, N631);
or OR2 (N1486, N1464, N1288);
nand NAND2 (N1487, N1477, N688);
buf BUF1 (N1488, N1483);
buf BUF1 (N1489, N1456);
xor XOR2 (N1490, N1487, N1428);
nor NOR3 (N1491, N1485, N1465, N846);
nand NAND2 (N1492, N1480, N237);
or OR3 (N1493, N1482, N676, N762);
or OR4 (N1494, N1488, N1138, N767, N1037);
nand NAND2 (N1495, N1474, N712);
nand NAND3 (N1496, N1492, N357, N1191);
and AND4 (N1497, N1494, N77, N1360, N683);
not NOT1 (N1498, N1491);
not NOT1 (N1499, N1484);
buf BUF1 (N1500, N1481);
nand NAND3 (N1501, N1497, N341, N825);
nor NOR2 (N1502, N1489, N113);
and AND2 (N1503, N1495, N527);
buf BUF1 (N1504, N1498);
nor NOR3 (N1505, N1501, N1431, N600);
nand NAND2 (N1506, N1500, N841);
not NOT1 (N1507, N1506);
nand NAND4 (N1508, N1504, N162, N395, N1068);
nor NOR3 (N1509, N1508, N576, N765);
buf BUF1 (N1510, N1503);
and AND3 (N1511, N1502, N1284, N1473);
xor XOR2 (N1512, N1509, N1276);
buf BUF1 (N1513, N1505);
or OR3 (N1514, N1511, N698, N1109);
buf BUF1 (N1515, N1510);
not NOT1 (N1516, N1490);
not NOT1 (N1517, N1499);
xor XOR2 (N1518, N1496, N1400);
buf BUF1 (N1519, N1513);
buf BUF1 (N1520, N1514);
nor NOR2 (N1521, N1512, N1168);
nand NAND4 (N1522, N1507, N342, N1027, N1510);
buf BUF1 (N1523, N1520);
not NOT1 (N1524, N1518);
and AND4 (N1525, N1516, N893, N1276, N1372);
buf BUF1 (N1526, N1525);
or OR3 (N1527, N1519, N191, N1354);
and AND2 (N1528, N1515, N1449);
and AND4 (N1529, N1523, N190, N125, N737);
nand NAND4 (N1530, N1486, N791, N728, N1361);
nand NAND3 (N1531, N1517, N1138, N67);
nor NOR4 (N1532, N1521, N981, N677, N113);
nor NOR3 (N1533, N1522, N334, N1329);
buf BUF1 (N1534, N1530);
buf BUF1 (N1535, N1527);
nor NOR3 (N1536, N1526, N66, N720);
xor XOR2 (N1537, N1533, N108);
nor NOR4 (N1538, N1535, N654, N315, N889);
and AND2 (N1539, N1536, N15);
or OR2 (N1540, N1532, N1196);
not NOT1 (N1541, N1524);
not NOT1 (N1542, N1538);
nor NOR2 (N1543, N1531, N1361);
and AND3 (N1544, N1493, N1275, N44);
nor NOR4 (N1545, N1534, N496, N798, N1043);
and AND2 (N1546, N1542, N1244);
and AND3 (N1547, N1546, N1213, N1170);
nor NOR4 (N1548, N1541, N781, N216, N1452);
buf BUF1 (N1549, N1545);
and AND3 (N1550, N1547, N1379, N907);
and AND4 (N1551, N1537, N184, N458, N218);
xor XOR2 (N1552, N1543, N1504);
nand NAND4 (N1553, N1540, N881, N859, N1105);
or OR3 (N1554, N1552, N1272, N688);
nor NOR4 (N1555, N1548, N1000, N1238, N638);
buf BUF1 (N1556, N1550);
buf BUF1 (N1557, N1544);
buf BUF1 (N1558, N1556);
buf BUF1 (N1559, N1551);
buf BUF1 (N1560, N1529);
not NOT1 (N1561, N1555);
and AND4 (N1562, N1560, N997, N1207, N1449);
xor XOR2 (N1563, N1561, N1110);
nand NAND3 (N1564, N1528, N1193, N1464);
not NOT1 (N1565, N1554);
nor NOR3 (N1566, N1558, N67, N1222);
not NOT1 (N1567, N1557);
and AND3 (N1568, N1553, N342, N493);
nand NAND3 (N1569, N1559, N1025, N793);
and AND4 (N1570, N1568, N1416, N459, N1298);
or OR3 (N1571, N1562, N1481, N67);
nand NAND2 (N1572, N1569, N136);
xor XOR2 (N1573, N1549, N1284);
xor XOR2 (N1574, N1572, N101);
not NOT1 (N1575, N1539);
or OR2 (N1576, N1566, N304);
xor XOR2 (N1577, N1575, N1146);
or OR2 (N1578, N1567, N492);
not NOT1 (N1579, N1574);
nand NAND2 (N1580, N1564, N1192);
nor NOR2 (N1581, N1578, N494);
nor NOR3 (N1582, N1573, N709, N501);
not NOT1 (N1583, N1580);
nor NOR2 (N1584, N1565, N875);
xor XOR2 (N1585, N1563, N289);
xor XOR2 (N1586, N1576, N1315);
and AND2 (N1587, N1570, N245);
or OR3 (N1588, N1585, N1350, N1579);
buf BUF1 (N1589, N615);
nand NAND3 (N1590, N1587, N1161, N393);
buf BUF1 (N1591, N1581);
or OR3 (N1592, N1590, N967, N980);
and AND3 (N1593, N1592, N413, N584);
nor NOR2 (N1594, N1588, N844);
and AND2 (N1595, N1584, N1313);
xor XOR2 (N1596, N1591, N262);
nor NOR4 (N1597, N1593, N255, N1193, N1274);
nor NOR4 (N1598, N1582, N294, N182, N1502);
xor XOR2 (N1599, N1596, N510);
not NOT1 (N1600, N1599);
nor NOR4 (N1601, N1571, N1224, N1551, N259);
nor NOR2 (N1602, N1595, N485);
nand NAND4 (N1603, N1594, N379, N1072, N334);
xor XOR2 (N1604, N1602, N381);
xor XOR2 (N1605, N1597, N535);
not NOT1 (N1606, N1603);
not NOT1 (N1607, N1589);
buf BUF1 (N1608, N1604);
or OR3 (N1609, N1598, N813, N894);
buf BUF1 (N1610, N1607);
nor NOR3 (N1611, N1610, N1306, N994);
nand NAND3 (N1612, N1586, N608, N20);
xor XOR2 (N1613, N1583, N510);
nor NOR4 (N1614, N1612, N1372, N1212, N1485);
buf BUF1 (N1615, N1608);
nand NAND4 (N1616, N1605, N205, N914, N253);
not NOT1 (N1617, N1613);
or OR4 (N1618, N1577, N1150, N1209, N1284);
not NOT1 (N1619, N1618);
and AND3 (N1620, N1616, N1292, N286);
nor NOR2 (N1621, N1606, N566);
buf BUF1 (N1622, N1615);
or OR4 (N1623, N1609, N1189, N649, N472);
nor NOR4 (N1624, N1600, N1149, N534, N1372);
or OR4 (N1625, N1617, N254, N962, N834);
and AND4 (N1626, N1619, N161, N89, N661);
not NOT1 (N1627, N1624);
nand NAND4 (N1628, N1622, N1511, N451, N933);
buf BUF1 (N1629, N1614);
not NOT1 (N1630, N1628);
nor NOR4 (N1631, N1623, N482, N436, N1231);
not NOT1 (N1632, N1631);
not NOT1 (N1633, N1625);
not NOT1 (N1634, N1627);
and AND4 (N1635, N1621, N537, N1588, N1121);
or OR4 (N1636, N1626, N1176, N932, N1449);
buf BUF1 (N1637, N1633);
and AND3 (N1638, N1620, N1153, N766);
not NOT1 (N1639, N1635);
or OR4 (N1640, N1632, N734, N640, N773);
nand NAND2 (N1641, N1630, N45);
nand NAND2 (N1642, N1636, N533);
nor NOR4 (N1643, N1640, N182, N113, N578);
buf BUF1 (N1644, N1639);
xor XOR2 (N1645, N1642, N424);
not NOT1 (N1646, N1645);
buf BUF1 (N1647, N1641);
not NOT1 (N1648, N1643);
or OR3 (N1649, N1648, N1049, N1588);
nor NOR3 (N1650, N1649, N9, N1054);
buf BUF1 (N1651, N1611);
nand NAND3 (N1652, N1637, N231, N1162);
nand NAND4 (N1653, N1647, N771, N749, N753);
nand NAND4 (N1654, N1651, N1052, N104, N473);
nor NOR2 (N1655, N1653, N789);
not NOT1 (N1656, N1655);
nand NAND4 (N1657, N1638, N633, N817, N168);
nor NOR3 (N1658, N1629, N1196, N155);
or OR3 (N1659, N1601, N611, N909);
or OR3 (N1660, N1656, N1321, N990);
xor XOR2 (N1661, N1659, N345);
nand NAND4 (N1662, N1650, N1614, N1415, N189);
not NOT1 (N1663, N1634);
or OR4 (N1664, N1652, N1441, N435, N1550);
or OR2 (N1665, N1661, N1481);
and AND4 (N1666, N1660, N54, N822, N393);
buf BUF1 (N1667, N1658);
nand NAND2 (N1668, N1667, N303);
nor NOR3 (N1669, N1644, N312, N1018);
xor XOR2 (N1670, N1646, N267);
nor NOR3 (N1671, N1657, N85, N1652);
nand NAND4 (N1672, N1666, N957, N1586, N1447);
not NOT1 (N1673, N1672);
nor NOR2 (N1674, N1664, N1078);
or OR2 (N1675, N1674, N1602);
buf BUF1 (N1676, N1668);
nor NOR2 (N1677, N1675, N1496);
nand NAND4 (N1678, N1677, N1197, N644, N709);
nor NOR3 (N1679, N1670, N204, N1413);
and AND3 (N1680, N1654, N1468, N1340);
or OR3 (N1681, N1665, N118, N387);
nor NOR3 (N1682, N1676, N464, N834);
nor NOR4 (N1683, N1671, N1288, N1519, N1241);
nand NAND3 (N1684, N1669, N146, N691);
buf BUF1 (N1685, N1662);
and AND3 (N1686, N1683, N798, N1103);
and AND3 (N1687, N1684, N1137, N246);
nor NOR3 (N1688, N1687, N646, N828);
not NOT1 (N1689, N1681);
nand NAND2 (N1690, N1682, N1647);
and AND2 (N1691, N1689, N198);
xor XOR2 (N1692, N1691, N1085);
not NOT1 (N1693, N1663);
and AND2 (N1694, N1690, N494);
nor NOR4 (N1695, N1673, N1339, N850, N1062);
and AND3 (N1696, N1693, N662, N482);
or OR2 (N1697, N1692, N397);
and AND2 (N1698, N1680, N1028);
or OR2 (N1699, N1698, N475);
not NOT1 (N1700, N1686);
or OR3 (N1701, N1688, N972, N1005);
nor NOR4 (N1702, N1700, N1551, N653, N1562);
and AND3 (N1703, N1697, N711, N612);
buf BUF1 (N1704, N1679);
nor NOR4 (N1705, N1696, N1370, N452, N1122);
buf BUF1 (N1706, N1703);
not NOT1 (N1707, N1705);
nand NAND3 (N1708, N1685, N1245, N422);
buf BUF1 (N1709, N1699);
nor NOR3 (N1710, N1709, N330, N30);
nor NOR3 (N1711, N1706, N1542, N593);
and AND3 (N1712, N1695, N823, N1566);
xor XOR2 (N1713, N1707, N946);
buf BUF1 (N1714, N1694);
nor NOR2 (N1715, N1702, N991);
or OR2 (N1716, N1710, N588);
buf BUF1 (N1717, N1716);
xor XOR2 (N1718, N1712, N1138);
buf BUF1 (N1719, N1715);
buf BUF1 (N1720, N1708);
xor XOR2 (N1721, N1719, N1480);
buf BUF1 (N1722, N1717);
and AND2 (N1723, N1678, N205);
not NOT1 (N1724, N1718);
buf BUF1 (N1725, N1722);
xor XOR2 (N1726, N1724, N950);
xor XOR2 (N1727, N1701, N1720);
xor XOR2 (N1728, N178, N182);
nand NAND4 (N1729, N1728, N926, N1057, N1386);
xor XOR2 (N1730, N1721, N284);
and AND2 (N1731, N1725, N852);
nand NAND3 (N1732, N1704, N1284, N533);
buf BUF1 (N1733, N1729);
xor XOR2 (N1734, N1726, N1712);
and AND4 (N1735, N1730, N1320, N472, N224);
or OR2 (N1736, N1711, N767);
not NOT1 (N1737, N1713);
xor XOR2 (N1738, N1732, N1597);
not NOT1 (N1739, N1731);
buf BUF1 (N1740, N1735);
buf BUF1 (N1741, N1723);
nand NAND3 (N1742, N1733, N149, N505);
buf BUF1 (N1743, N1741);
nand NAND3 (N1744, N1740, N181, N769);
buf BUF1 (N1745, N1734);
nand NAND3 (N1746, N1738, N472, N1319);
xor XOR2 (N1747, N1737, N1663);
not NOT1 (N1748, N1743);
nor NOR3 (N1749, N1739, N955, N947);
nand NAND2 (N1750, N1727, N1277);
nand NAND2 (N1751, N1736, N424);
buf BUF1 (N1752, N1748);
nor NOR3 (N1753, N1749, N1368, N1318);
and AND4 (N1754, N1752, N956, N1237, N62);
not NOT1 (N1755, N1745);
xor XOR2 (N1756, N1754, N273);
nand NAND2 (N1757, N1742, N1525);
nor NOR4 (N1758, N1757, N1058, N1166, N1179);
or OR4 (N1759, N1746, N384, N530, N308);
not NOT1 (N1760, N1750);
not NOT1 (N1761, N1755);
not NOT1 (N1762, N1714);
nand NAND4 (N1763, N1760, N122, N354, N597);
buf BUF1 (N1764, N1762);
and AND3 (N1765, N1761, N403, N315);
nor NOR4 (N1766, N1744, N1126, N1618, N628);
nand NAND4 (N1767, N1758, N506, N377, N619);
nand NAND2 (N1768, N1759, N1621);
nand NAND4 (N1769, N1751, N1400, N1443, N222);
not NOT1 (N1770, N1765);
or OR4 (N1771, N1766, N991, N658, N513);
buf BUF1 (N1772, N1769);
and AND2 (N1773, N1768, N257);
xor XOR2 (N1774, N1773, N1655);
not NOT1 (N1775, N1770);
or OR4 (N1776, N1767, N387, N586, N768);
buf BUF1 (N1777, N1753);
xor XOR2 (N1778, N1756, N1645);
xor XOR2 (N1779, N1776, N715);
not NOT1 (N1780, N1777);
buf BUF1 (N1781, N1764);
or OR3 (N1782, N1781, N825, N1735);
not NOT1 (N1783, N1774);
nor NOR3 (N1784, N1783, N708, N952);
or OR4 (N1785, N1778, N1444, N169, N1470);
buf BUF1 (N1786, N1785);
nand NAND4 (N1787, N1782, N1470, N104, N554);
xor XOR2 (N1788, N1786, N1210);
not NOT1 (N1789, N1780);
or OR3 (N1790, N1788, N660, N1274);
or OR4 (N1791, N1787, N471, N1255, N38);
nor NOR4 (N1792, N1747, N562, N718, N641);
not NOT1 (N1793, N1763);
and AND4 (N1794, N1790, N1168, N1085, N1283);
or OR4 (N1795, N1772, N736, N596, N1334);
or OR4 (N1796, N1784, N265, N998, N1723);
xor XOR2 (N1797, N1779, N1695);
or OR4 (N1798, N1795, N1462, N23, N1208);
nand NAND2 (N1799, N1789, N556);
and AND2 (N1800, N1775, N1259);
and AND2 (N1801, N1796, N805);
not NOT1 (N1802, N1797);
nor NOR2 (N1803, N1801, N1172);
and AND3 (N1804, N1803, N991, N1582);
not NOT1 (N1805, N1791);
xor XOR2 (N1806, N1794, N267);
buf BUF1 (N1807, N1804);
buf BUF1 (N1808, N1792);
nand NAND3 (N1809, N1805, N1459, N1401);
or OR3 (N1810, N1808, N1539, N403);
buf BUF1 (N1811, N1806);
nand NAND3 (N1812, N1800, N500, N735);
not NOT1 (N1813, N1809);
and AND2 (N1814, N1811, N1738);
nand NAND2 (N1815, N1807, N110);
nor NOR4 (N1816, N1813, N1045, N1025, N380);
nor NOR4 (N1817, N1814, N1695, N1076, N1155);
xor XOR2 (N1818, N1802, N272);
nor NOR4 (N1819, N1815, N252, N909, N1430);
nand NAND4 (N1820, N1810, N1605, N504, N1467);
not NOT1 (N1821, N1798);
not NOT1 (N1822, N1799);
nand NAND4 (N1823, N1822, N1212, N584, N218);
buf BUF1 (N1824, N1820);
nor NOR3 (N1825, N1817, N1666, N1023);
not NOT1 (N1826, N1824);
xor XOR2 (N1827, N1823, N1425);
not NOT1 (N1828, N1821);
or OR3 (N1829, N1812, N1626, N545);
or OR4 (N1830, N1771, N627, N1200, N1449);
nand NAND4 (N1831, N1829, N536, N214, N1649);
or OR2 (N1832, N1828, N1325);
nand NAND2 (N1833, N1832, N641);
nor NOR4 (N1834, N1831, N1183, N69, N53);
and AND2 (N1835, N1819, N915);
buf BUF1 (N1836, N1830);
xor XOR2 (N1837, N1833, N465);
nor NOR4 (N1838, N1793, N1618, N1651, N389);
xor XOR2 (N1839, N1826, N220);
buf BUF1 (N1840, N1816);
nor NOR4 (N1841, N1835, N125, N1545, N1658);
nand NAND2 (N1842, N1836, N1392);
not NOT1 (N1843, N1840);
and AND3 (N1844, N1825, N282, N48);
nor NOR4 (N1845, N1827, N1109, N1725, N737);
buf BUF1 (N1846, N1837);
not NOT1 (N1847, N1842);
nor NOR3 (N1848, N1847, N636, N684);
nand NAND4 (N1849, N1834, N598, N835, N1420);
not NOT1 (N1850, N1841);
nor NOR4 (N1851, N1846, N1705, N991, N498);
nor NOR3 (N1852, N1849, N1579, N764);
nand NAND2 (N1853, N1850, N701);
buf BUF1 (N1854, N1843);
nand NAND2 (N1855, N1854, N1506);
nand NAND4 (N1856, N1852, N1449, N1327, N63);
not NOT1 (N1857, N1853);
xor XOR2 (N1858, N1818, N396);
buf BUF1 (N1859, N1845);
xor XOR2 (N1860, N1838, N1789);
and AND4 (N1861, N1839, N1413, N330, N1498);
not NOT1 (N1862, N1859);
nor NOR3 (N1863, N1856, N846, N1363);
buf BUF1 (N1864, N1858);
or OR3 (N1865, N1848, N1473, N224);
and AND2 (N1866, N1844, N1572);
or OR4 (N1867, N1860, N1525, N238, N558);
buf BUF1 (N1868, N1863);
buf BUF1 (N1869, N1862);
not NOT1 (N1870, N1864);
nor NOR3 (N1871, N1869, N477, N1622);
and AND2 (N1872, N1855, N925);
buf BUF1 (N1873, N1865);
buf BUF1 (N1874, N1870);
xor XOR2 (N1875, N1857, N944);
buf BUF1 (N1876, N1866);
nand NAND4 (N1877, N1876, N210, N509, N481);
and AND2 (N1878, N1875, N383);
xor XOR2 (N1879, N1878, N1091);
or OR3 (N1880, N1871, N1048, N482);
nand NAND4 (N1881, N1867, N1550, N1091, N153);
not NOT1 (N1882, N1868);
or OR4 (N1883, N1882, N416, N341, N77);
and AND2 (N1884, N1883, N1034);
or OR4 (N1885, N1879, N697, N292, N1209);
nand NAND4 (N1886, N1881, N1801, N142, N815);
and AND2 (N1887, N1873, N816);
not NOT1 (N1888, N1872);
or OR3 (N1889, N1851, N1176, N366);
buf BUF1 (N1890, N1886);
xor XOR2 (N1891, N1885, N1628);
buf BUF1 (N1892, N1877);
nor NOR4 (N1893, N1861, N1874, N1726, N235);
or OR2 (N1894, N1249, N386);
buf BUF1 (N1895, N1893);
or OR3 (N1896, N1892, N952, N1653);
and AND4 (N1897, N1887, N1007, N1469, N193);
xor XOR2 (N1898, N1894, N1742);
and AND3 (N1899, N1888, N1252, N1770);
buf BUF1 (N1900, N1895);
nor NOR3 (N1901, N1900, N391, N1086);
not NOT1 (N1902, N1890);
nor NOR2 (N1903, N1901, N233);
nand NAND3 (N1904, N1891, N336, N1526);
nor NOR4 (N1905, N1903, N1371, N131, N480);
buf BUF1 (N1906, N1889);
xor XOR2 (N1907, N1896, N1857);
or OR2 (N1908, N1898, N1428);
buf BUF1 (N1909, N1907);
xor XOR2 (N1910, N1909, N1520);
nor NOR2 (N1911, N1902, N1574);
buf BUF1 (N1912, N1905);
xor XOR2 (N1913, N1908, N512);
and AND3 (N1914, N1904, N176, N1648);
buf BUF1 (N1915, N1880);
nand NAND2 (N1916, N1884, N920);
not NOT1 (N1917, N1897);
xor XOR2 (N1918, N1906, N1386);
buf BUF1 (N1919, N1912);
nor NOR2 (N1920, N1917, N1416);
and AND2 (N1921, N1914, N21);
and AND3 (N1922, N1913, N400, N1511);
not NOT1 (N1923, N1921);
and AND2 (N1924, N1915, N1698);
xor XOR2 (N1925, N1918, N809);
or OR3 (N1926, N1923, N347, N1323);
nand NAND2 (N1927, N1926, N315);
or OR3 (N1928, N1922, N1906, N1230);
nor NOR2 (N1929, N1920, N827);
nand NAND4 (N1930, N1911, N1344, N1689, N1268);
or OR2 (N1931, N1925, N252);
nor NOR3 (N1932, N1916, N1540, N804);
nor NOR4 (N1933, N1928, N1499, N1092, N1898);
nor NOR3 (N1934, N1930, N454, N523);
or OR4 (N1935, N1927, N1420, N168, N92);
or OR2 (N1936, N1910, N1792);
buf BUF1 (N1937, N1936);
nor NOR2 (N1938, N1919, N531);
not NOT1 (N1939, N1899);
nand NAND3 (N1940, N1931, N641, N947);
or OR4 (N1941, N1938, N1422, N590, N210);
not NOT1 (N1942, N1933);
nor NOR2 (N1943, N1937, N1821);
or OR2 (N1944, N1940, N1318);
xor XOR2 (N1945, N1934, N69);
or OR2 (N1946, N1932, N852);
or OR4 (N1947, N1944, N601, N532, N950);
and AND3 (N1948, N1929, N1821, N1480);
buf BUF1 (N1949, N1948);
and AND3 (N1950, N1947, N1830, N489);
nand NAND4 (N1951, N1941, N1628, N1583, N1920);
not NOT1 (N1952, N1945);
nand NAND4 (N1953, N1943, N1081, N1081, N248);
xor XOR2 (N1954, N1946, N1180);
not NOT1 (N1955, N1951);
xor XOR2 (N1956, N1924, N834);
xor XOR2 (N1957, N1935, N1173);
and AND2 (N1958, N1942, N256);
and AND4 (N1959, N1953, N578, N1624, N1155);
nor NOR4 (N1960, N1954, N970, N1365, N1704);
not NOT1 (N1961, N1957);
not NOT1 (N1962, N1960);
xor XOR2 (N1963, N1956, N1639);
nor NOR3 (N1964, N1949, N1766, N1213);
nor NOR4 (N1965, N1950, N60, N1672, N1097);
nor NOR2 (N1966, N1963, N1885);
not NOT1 (N1967, N1966);
buf BUF1 (N1968, N1939);
not NOT1 (N1969, N1965);
or OR2 (N1970, N1962, N1697);
xor XOR2 (N1971, N1955, N1585);
or OR2 (N1972, N1958, N1466);
nor NOR4 (N1973, N1969, N1711, N1264, N734);
nand NAND4 (N1974, N1972, N1750, N1646, N326);
xor XOR2 (N1975, N1961, N1620);
or OR2 (N1976, N1970, N1577);
xor XOR2 (N1977, N1967, N1147);
not NOT1 (N1978, N1968);
xor XOR2 (N1979, N1977, N1691);
nor NOR3 (N1980, N1975, N1803, N518);
xor XOR2 (N1981, N1978, N1968);
xor XOR2 (N1982, N1952, N822);
and AND2 (N1983, N1964, N323);
nand NAND3 (N1984, N1973, N966, N1333);
or OR3 (N1985, N1974, N1390, N951);
or OR2 (N1986, N1979, N1302);
nor NOR2 (N1987, N1980, N166);
buf BUF1 (N1988, N1983);
xor XOR2 (N1989, N1971, N479);
or OR2 (N1990, N1989, N162);
not NOT1 (N1991, N1986);
or OR2 (N1992, N1976, N1416);
nand NAND3 (N1993, N1959, N421, N627);
nor NOR4 (N1994, N1988, N1158, N1291, N436);
and AND2 (N1995, N1981, N598);
not NOT1 (N1996, N1987);
nand NAND3 (N1997, N1994, N1033, N123);
nor NOR2 (N1998, N1995, N901);
nand NAND4 (N1999, N1982, N447, N337, N1277);
xor XOR2 (N2000, N1990, N54);
nor NOR3 (N2001, N1997, N1258, N280);
xor XOR2 (N2002, N1993, N340);
or OR3 (N2003, N1992, N714, N83);
nand NAND3 (N2004, N1985, N1842, N1051);
buf BUF1 (N2005, N2001);
and AND3 (N2006, N2002, N149, N955);
nor NOR3 (N2007, N2006, N469, N663);
and AND2 (N2008, N1998, N744);
or OR3 (N2009, N2005, N1955, N19);
nand NAND4 (N2010, N2009, N1231, N384, N1940);
xor XOR2 (N2011, N1984, N666);
not NOT1 (N2012, N2000);
not NOT1 (N2013, N2003);
buf BUF1 (N2014, N2012);
not NOT1 (N2015, N1996);
buf BUF1 (N2016, N2013);
or OR2 (N2017, N2010, N792);
not NOT1 (N2018, N2017);
xor XOR2 (N2019, N2014, N1028);
xor XOR2 (N2020, N1991, N200);
buf BUF1 (N2021, N2018);
not NOT1 (N2022, N2008);
not NOT1 (N2023, N1999);
xor XOR2 (N2024, N2004, N556);
xor XOR2 (N2025, N2024, N759);
not NOT1 (N2026, N2021);
or OR3 (N2027, N2025, N1185, N1360);
and AND2 (N2028, N2023, N529);
and AND4 (N2029, N2020, N597, N1624, N159);
xor XOR2 (N2030, N2028, N1976);
nand NAND2 (N2031, N2007, N1444);
and AND4 (N2032, N2029, N848, N1334, N538);
nand NAND4 (N2033, N2027, N801, N611, N1799);
nand NAND3 (N2034, N2030, N462, N1294);
and AND3 (N2035, N2016, N51, N1819);
nor NOR4 (N2036, N2033, N69, N1884, N853);
xor XOR2 (N2037, N2034, N471);
not NOT1 (N2038, N2036);
not NOT1 (N2039, N2038);
xor XOR2 (N2040, N2022, N1124);
xor XOR2 (N2041, N2037, N1027);
and AND3 (N2042, N2019, N740, N380);
not NOT1 (N2043, N2026);
xor XOR2 (N2044, N2015, N684);
nand NAND4 (N2045, N2041, N1356, N563, N329);
nor NOR3 (N2046, N2011, N448, N1193);
xor XOR2 (N2047, N2035, N311);
and AND3 (N2048, N2039, N691, N1130);
not NOT1 (N2049, N2040);
xor XOR2 (N2050, N2043, N1332);
xor XOR2 (N2051, N2046, N153);
nor NOR3 (N2052, N2049, N808, N449);
and AND4 (N2053, N2048, N1406, N811, N613);
nor NOR2 (N2054, N2042, N565);
and AND4 (N2055, N2054, N1711, N1848, N301);
and AND3 (N2056, N2047, N469, N1083);
nand NAND3 (N2057, N2050, N406, N626);
and AND3 (N2058, N2044, N1356, N1185);
not NOT1 (N2059, N2057);
nand NAND4 (N2060, N2045, N1039, N1618, N1927);
nor NOR3 (N2061, N2058, N2034, N514);
not NOT1 (N2062, N2061);
buf BUF1 (N2063, N2056);
not NOT1 (N2064, N2032);
nand NAND2 (N2065, N2052, N1607);
and AND4 (N2066, N2051, N1726, N508, N1036);
buf BUF1 (N2067, N2066);
buf BUF1 (N2068, N2065);
xor XOR2 (N2069, N2068, N454);
buf BUF1 (N2070, N2060);
and AND3 (N2071, N2059, N1376, N1341);
nand NAND3 (N2072, N2053, N669, N1515);
or OR2 (N2073, N2071, N1964);
buf BUF1 (N2074, N2069);
not NOT1 (N2075, N2074);
xor XOR2 (N2076, N2063, N1793);
or OR3 (N2077, N2073, N809, N1545);
or OR3 (N2078, N2055, N1411, N612);
nand NAND3 (N2079, N2070, N1812, N1695);
xor XOR2 (N2080, N2031, N625);
xor XOR2 (N2081, N2076, N1662);
not NOT1 (N2082, N2077);
xor XOR2 (N2083, N2064, N1100);
nor NOR3 (N2084, N2082, N1337, N1522);
nor NOR4 (N2085, N2079, N1531, N822, N811);
xor XOR2 (N2086, N2080, N553);
nand NAND3 (N2087, N2078, N1019, N651);
buf BUF1 (N2088, N2084);
or OR3 (N2089, N2083, N713, N802);
not NOT1 (N2090, N2085);
not NOT1 (N2091, N2072);
xor XOR2 (N2092, N2088, N1815);
xor XOR2 (N2093, N2090, N1052);
not NOT1 (N2094, N2089);
and AND3 (N2095, N2087, N1884, N367);
and AND2 (N2096, N2093, N257);
nor NOR3 (N2097, N2081, N1822, N1006);
nor NOR3 (N2098, N2092, N1789, N1888);
nor NOR2 (N2099, N2067, N332);
xor XOR2 (N2100, N2099, N690);
not NOT1 (N2101, N2094);
or OR3 (N2102, N2062, N488, N961);
nand NAND3 (N2103, N2075, N2026, N14);
xor XOR2 (N2104, N2102, N444);
or OR3 (N2105, N2104, N1433, N1224);
nor NOR4 (N2106, N2105, N1825, N609, N770);
xor XOR2 (N2107, N2095, N942);
not NOT1 (N2108, N2091);
nand NAND4 (N2109, N2103, N1591, N1575, N1335);
xor XOR2 (N2110, N2109, N1502);
nand NAND3 (N2111, N2110, N459, N1830);
nor NOR2 (N2112, N2086, N814);
and AND3 (N2113, N2106, N1923, N281);
not NOT1 (N2114, N2100);
not NOT1 (N2115, N2108);
not NOT1 (N2116, N2114);
nor NOR4 (N2117, N2116, N1268, N1649, N926);
xor XOR2 (N2118, N2115, N301);
buf BUF1 (N2119, N2098);
or OR2 (N2120, N2096, N1411);
or OR4 (N2121, N2097, N1970, N1013, N102);
not NOT1 (N2122, N2111);
xor XOR2 (N2123, N2121, N1021);
and AND2 (N2124, N2112, N2051);
nor NOR4 (N2125, N2120, N2000, N1934, N740);
or OR4 (N2126, N2113, N334, N579, N2031);
buf BUF1 (N2127, N2124);
or OR4 (N2128, N2123, N1935, N232, N773);
or OR3 (N2129, N2125, N550, N1810);
and AND2 (N2130, N2122, N31);
or OR4 (N2131, N2119, N517, N2039, N1947);
xor XOR2 (N2132, N2130, N1298);
and AND2 (N2133, N2132, N1866);
nor NOR2 (N2134, N2131, N487);
or OR3 (N2135, N2126, N1350, N788);
or OR3 (N2136, N2107, N764, N1251);
nand NAND2 (N2137, N2118, N1176);
not NOT1 (N2138, N2127);
nor NOR3 (N2139, N2135, N2060, N2105);
not NOT1 (N2140, N2133);
buf BUF1 (N2141, N2137);
nor NOR4 (N2142, N2134, N1682, N1507, N475);
or OR2 (N2143, N2142, N1393);
buf BUF1 (N2144, N2138);
nand NAND3 (N2145, N2101, N1192, N226);
or OR3 (N2146, N2144, N1578, N469);
nand NAND2 (N2147, N2140, N284);
and AND2 (N2148, N2143, N1758);
not NOT1 (N2149, N2117);
or OR2 (N2150, N2148, N2087);
buf BUF1 (N2151, N2129);
xor XOR2 (N2152, N2141, N1185);
nor NOR3 (N2153, N2146, N118, N206);
or OR3 (N2154, N2150, N2119, N941);
and AND4 (N2155, N2147, N1051, N1116, N2139);
nor NOR3 (N2156, N1730, N1728, N265);
not NOT1 (N2157, N2155);
xor XOR2 (N2158, N2152, N958);
nor NOR3 (N2159, N2145, N731, N1468);
xor XOR2 (N2160, N2128, N789);
nor NOR4 (N2161, N2149, N1706, N1124, N1021);
nand NAND2 (N2162, N2158, N74);
xor XOR2 (N2163, N2136, N1941);
or OR2 (N2164, N2154, N179);
or OR2 (N2165, N2164, N1877);
not NOT1 (N2166, N2159);
and AND4 (N2167, N2156, N810, N1887, N1963);
or OR4 (N2168, N2151, N1489, N97, N1110);
xor XOR2 (N2169, N2153, N1747);
buf BUF1 (N2170, N2165);
xor XOR2 (N2171, N2160, N1886);
and AND2 (N2172, N2170, N1469);
xor XOR2 (N2173, N2163, N1555);
nor NOR2 (N2174, N2171, N1242);
and AND3 (N2175, N2167, N363, N346);
xor XOR2 (N2176, N2161, N463);
buf BUF1 (N2177, N2175);
not NOT1 (N2178, N2176);
and AND3 (N2179, N2169, N1536, N377);
nand NAND3 (N2180, N2162, N418, N829);
xor XOR2 (N2181, N2172, N1487);
or OR4 (N2182, N2178, N1366, N407, N883);
not NOT1 (N2183, N2168);
not NOT1 (N2184, N2179);
or OR2 (N2185, N2180, N1823);
and AND3 (N2186, N2166, N1518, N1259);
xor XOR2 (N2187, N2157, N2106);
and AND2 (N2188, N2182, N1442);
xor XOR2 (N2189, N2187, N1927);
nor NOR2 (N2190, N2186, N1268);
nand NAND4 (N2191, N2174, N1245, N682, N390);
not NOT1 (N2192, N2173);
not NOT1 (N2193, N2184);
xor XOR2 (N2194, N2191, N65);
buf BUF1 (N2195, N2189);
nand NAND3 (N2196, N2192, N101, N81);
not NOT1 (N2197, N2190);
xor XOR2 (N2198, N2177, N112);
and AND3 (N2199, N2198, N1454, N110);
not NOT1 (N2200, N2188);
xor XOR2 (N2201, N2183, N1427);
or OR4 (N2202, N2197, N1533, N199, N1917);
nor NOR3 (N2203, N2202, N72, N2001);
nor NOR2 (N2204, N2193, N596);
buf BUF1 (N2205, N2181);
buf BUF1 (N2206, N2185);
buf BUF1 (N2207, N2194);
and AND3 (N2208, N2203, N785, N798);
or OR3 (N2209, N2206, N2077, N1763);
or OR4 (N2210, N2205, N1136, N1196, N22);
nand NAND3 (N2211, N2204, N1327, N1865);
or OR4 (N2212, N2208, N1251, N940, N613);
not NOT1 (N2213, N2212);
or OR2 (N2214, N2200, N1681);
and AND3 (N2215, N2201, N675, N2117);
nor NOR2 (N2216, N2215, N1383);
buf BUF1 (N2217, N2214);
buf BUF1 (N2218, N2210);
xor XOR2 (N2219, N2213, N1504);
nand NAND4 (N2220, N2199, N2116, N1658, N46);
nand NAND3 (N2221, N2195, N1986, N2097);
nor NOR2 (N2222, N2221, N2056);
nor NOR4 (N2223, N2217, N1398, N1004, N171);
nor NOR4 (N2224, N2216, N2083, N64, N887);
or OR2 (N2225, N2220, N845);
buf BUF1 (N2226, N2209);
nor NOR2 (N2227, N2196, N370);
or OR3 (N2228, N2222, N1167, N1893);
buf BUF1 (N2229, N2228);
or OR4 (N2230, N2219, N1968, N1413, N290);
nor NOR4 (N2231, N2225, N2048, N843, N1848);
and AND4 (N2232, N2227, N1355, N1748, N811);
buf BUF1 (N2233, N2232);
not NOT1 (N2234, N2207);
or OR3 (N2235, N2230, N885, N389);
or OR3 (N2236, N2224, N1210, N1244);
not NOT1 (N2237, N2229);
and AND3 (N2238, N2218, N2110, N155);
or OR2 (N2239, N2235, N737);
not NOT1 (N2240, N2211);
xor XOR2 (N2241, N2236, N1350);
and AND4 (N2242, N2231, N830, N1766, N1000);
buf BUF1 (N2243, N2234);
not NOT1 (N2244, N2237);
nand NAND4 (N2245, N2242, N2031, N975, N1740);
xor XOR2 (N2246, N2243, N643);
xor XOR2 (N2247, N2223, N1367);
or OR4 (N2248, N2241, N2103, N707, N2215);
buf BUF1 (N2249, N2246);
not NOT1 (N2250, N2247);
and AND2 (N2251, N2244, N599);
and AND3 (N2252, N2250, N610, N1251);
and AND3 (N2253, N2240, N1070, N245);
not NOT1 (N2254, N2249);
not NOT1 (N2255, N2226);
and AND3 (N2256, N2252, N2173, N1772);
xor XOR2 (N2257, N2255, N767);
and AND3 (N2258, N2238, N388, N1492);
and AND3 (N2259, N2248, N376, N1502);
xor XOR2 (N2260, N2245, N1231);
nor NOR3 (N2261, N2233, N419, N2194);
nand NAND3 (N2262, N2258, N164, N154);
and AND3 (N2263, N2254, N1025, N1351);
buf BUF1 (N2264, N2259);
or OR4 (N2265, N2253, N1793, N761, N573);
nand NAND4 (N2266, N2263, N1203, N1274, N508);
and AND4 (N2267, N2257, N235, N1086, N1731);
not NOT1 (N2268, N2239);
not NOT1 (N2269, N2265);
buf BUF1 (N2270, N2261);
nor NOR2 (N2271, N2268, N355);
nand NAND4 (N2272, N2264, N9, N501, N81);
or OR4 (N2273, N2260, N855, N2053, N1975);
or OR2 (N2274, N2271, N162);
and AND4 (N2275, N2256, N262, N550, N1045);
nor NOR2 (N2276, N2270, N1447);
not NOT1 (N2277, N2251);
nand NAND3 (N2278, N2266, N1391, N1368);
or OR2 (N2279, N2274, N1210);
xor XOR2 (N2280, N2269, N1142);
nand NAND3 (N2281, N2279, N970, N1124);
and AND2 (N2282, N2278, N667);
buf BUF1 (N2283, N2276);
buf BUF1 (N2284, N2283);
buf BUF1 (N2285, N2275);
not NOT1 (N2286, N2262);
buf BUF1 (N2287, N2282);
not NOT1 (N2288, N2277);
nand NAND2 (N2289, N2273, N829);
xor XOR2 (N2290, N2289, N209);
buf BUF1 (N2291, N2290);
nand NAND4 (N2292, N2287, N567, N1938, N995);
or OR3 (N2293, N2280, N1877, N640);
not NOT1 (N2294, N2293);
not NOT1 (N2295, N2292);
nor NOR4 (N2296, N2285, N560, N2212, N886);
not NOT1 (N2297, N2294);
and AND2 (N2298, N2288, N1737);
or OR4 (N2299, N2295, N769, N1095, N1556);
nor NOR2 (N2300, N2267, N327);
buf BUF1 (N2301, N2284);
nand NAND3 (N2302, N2291, N1226, N1737);
xor XOR2 (N2303, N2281, N952);
and AND3 (N2304, N2298, N1676, N1337);
nor NOR3 (N2305, N2272, N2091, N518);
xor XOR2 (N2306, N2296, N1449);
buf BUF1 (N2307, N2286);
nand NAND3 (N2308, N2302, N1809, N2036);
nand NAND4 (N2309, N2307, N2297, N614, N2068);
not NOT1 (N2310, N1129);
or OR3 (N2311, N2305, N1422, N1810);
xor XOR2 (N2312, N2308, N861);
not NOT1 (N2313, N2303);
not NOT1 (N2314, N2306);
and AND4 (N2315, N2311, N1896, N2041, N257);
nor NOR3 (N2316, N2312, N704, N586);
and AND3 (N2317, N2301, N130, N38);
nand NAND2 (N2318, N2304, N2007);
not NOT1 (N2319, N2310);
or OR2 (N2320, N2314, N677);
buf BUF1 (N2321, N2319);
or OR4 (N2322, N2309, N2224, N1851, N1679);
buf BUF1 (N2323, N2320);
nor NOR4 (N2324, N2317, N1859, N2111, N574);
xor XOR2 (N2325, N2299, N570);
or OR2 (N2326, N2324, N1186);
or OR2 (N2327, N2321, N1686);
nand NAND2 (N2328, N2313, N128);
xor XOR2 (N2329, N2300, N282);
not NOT1 (N2330, N2322);
nand NAND3 (N2331, N2325, N668, N1967);
xor XOR2 (N2332, N2327, N1339);
buf BUF1 (N2333, N2326);
and AND2 (N2334, N2333, N2268);
nor NOR2 (N2335, N2331, N282);
and AND2 (N2336, N2329, N1999);
nor NOR4 (N2337, N2335, N1261, N850, N86);
buf BUF1 (N2338, N2323);
nor NOR3 (N2339, N2328, N1522, N1233);
not NOT1 (N2340, N2315);
xor XOR2 (N2341, N2332, N1660);
and AND2 (N2342, N2318, N1685);
and AND4 (N2343, N2316, N110, N830, N1161);
not NOT1 (N2344, N2340);
nor NOR2 (N2345, N2342, N561);
buf BUF1 (N2346, N2344);
nand NAND4 (N2347, N2336, N1557, N2098, N1277);
xor XOR2 (N2348, N2334, N908);
xor XOR2 (N2349, N2341, N1708);
and AND2 (N2350, N2349, N2193);
nand NAND4 (N2351, N2339, N1363, N632, N1746);
or OR3 (N2352, N2338, N1452, N769);
not NOT1 (N2353, N2351);
xor XOR2 (N2354, N2343, N643);
buf BUF1 (N2355, N2337);
xor XOR2 (N2356, N2354, N602);
buf BUF1 (N2357, N2345);
buf BUF1 (N2358, N2330);
or OR2 (N2359, N2353, N1341);
buf BUF1 (N2360, N2347);
nand NAND4 (N2361, N2355, N25, N1213, N19);
nand NAND3 (N2362, N2357, N646, N1055);
or OR3 (N2363, N2360, N1541, N710);
xor XOR2 (N2364, N2362, N1898);
or OR4 (N2365, N2352, N1183, N202, N1023);
xor XOR2 (N2366, N2346, N1118);
or OR2 (N2367, N2348, N182);
or OR3 (N2368, N2356, N1603, N1616);
nand NAND3 (N2369, N2361, N575, N1946);
nor NOR4 (N2370, N2368, N1777, N308, N704);
nor NOR3 (N2371, N2370, N1899, N1613);
nor NOR2 (N2372, N2350, N1621);
and AND4 (N2373, N2369, N1992, N584, N2132);
nand NAND2 (N2374, N2364, N153);
nand NAND4 (N2375, N2371, N111, N1744, N1894);
not NOT1 (N2376, N2373);
buf BUF1 (N2377, N2376);
buf BUF1 (N2378, N2377);
xor XOR2 (N2379, N2358, N1318);
xor XOR2 (N2380, N2367, N1693);
and AND2 (N2381, N2365, N799);
not NOT1 (N2382, N2363);
or OR2 (N2383, N2374, N1595);
not NOT1 (N2384, N2381);
not NOT1 (N2385, N2378);
nand NAND2 (N2386, N2383, N812);
buf BUF1 (N2387, N2379);
buf BUF1 (N2388, N2385);
not NOT1 (N2389, N2382);
or OR3 (N2390, N2380, N1938, N1947);
xor XOR2 (N2391, N2375, N416);
not NOT1 (N2392, N2359);
xor XOR2 (N2393, N2389, N2141);
nor NOR2 (N2394, N2392, N2179);
and AND2 (N2395, N2390, N1768);
nand NAND2 (N2396, N2395, N882);
xor XOR2 (N2397, N2384, N820);
xor XOR2 (N2398, N2372, N363);
nand NAND3 (N2399, N2386, N388, N2185);
xor XOR2 (N2400, N2396, N927);
nand NAND4 (N2401, N2397, N770, N2394, N2046);
and AND4 (N2402, N1776, N993, N1917, N90);
xor XOR2 (N2403, N2366, N610);
buf BUF1 (N2404, N2401);
buf BUF1 (N2405, N2393);
and AND4 (N2406, N2387, N2388, N2283, N278);
nand NAND4 (N2407, N628, N1159, N614, N1969);
buf BUF1 (N2408, N2402);
nor NOR3 (N2409, N2399, N481, N354);
nor NOR2 (N2410, N2405, N611);
xor XOR2 (N2411, N2403, N813);
buf BUF1 (N2412, N2391);
nor NOR2 (N2413, N2409, N1843);
not NOT1 (N2414, N2411);
nand NAND2 (N2415, N2404, N1318);
and AND4 (N2416, N2412, N1598, N545, N1704);
xor XOR2 (N2417, N2415, N1175);
not NOT1 (N2418, N2414);
or OR4 (N2419, N2418, N1265, N1881, N1152);
buf BUF1 (N2420, N2398);
buf BUF1 (N2421, N2419);
not NOT1 (N2422, N2407);
or OR2 (N2423, N2413, N2164);
or OR3 (N2424, N2422, N1379, N2124);
buf BUF1 (N2425, N2406);
not NOT1 (N2426, N2424);
buf BUF1 (N2427, N2420);
not NOT1 (N2428, N2425);
or OR3 (N2429, N2423, N176, N1346);
buf BUF1 (N2430, N2429);
xor XOR2 (N2431, N2417, N307);
buf BUF1 (N2432, N2426);
xor XOR2 (N2433, N2432, N817);
nand NAND4 (N2434, N2400, N142, N101, N116);
xor XOR2 (N2435, N2431, N624);
xor XOR2 (N2436, N2434, N2280);
xor XOR2 (N2437, N2416, N328);
not NOT1 (N2438, N2427);
buf BUF1 (N2439, N2438);
nand NAND3 (N2440, N2435, N2116, N450);
nor NOR4 (N2441, N2433, N290, N274, N1201);
nand NAND3 (N2442, N2440, N4, N1975);
not NOT1 (N2443, N2408);
xor XOR2 (N2444, N2439, N2190);
and AND3 (N2445, N2428, N1150, N2197);
nor NOR4 (N2446, N2444, N68, N1199, N169);
or OR3 (N2447, N2445, N2281, N443);
buf BUF1 (N2448, N2430);
or OR2 (N2449, N2421, N677);
buf BUF1 (N2450, N2443);
or OR2 (N2451, N2442, N1940);
nor NOR4 (N2452, N2436, N607, N2349, N1595);
and AND3 (N2453, N2448, N1911, N744);
or OR2 (N2454, N2452, N2385);
not NOT1 (N2455, N2447);
buf BUF1 (N2456, N2437);
buf BUF1 (N2457, N2453);
nor NOR2 (N2458, N2450, N1215);
buf BUF1 (N2459, N2456);
nand NAND2 (N2460, N2446, N1928);
not NOT1 (N2461, N2449);
xor XOR2 (N2462, N2451, N1329);
or OR3 (N2463, N2457, N2099, N257);
nor NOR3 (N2464, N2463, N884, N2);
buf BUF1 (N2465, N2441);
nand NAND2 (N2466, N2464, N256);
or OR4 (N2467, N2459, N135, N51, N361);
nor NOR2 (N2468, N2466, N2372);
nand NAND3 (N2469, N2462, N2009, N1785);
and AND3 (N2470, N2468, N150, N1847);
nand NAND3 (N2471, N2455, N1800, N1377);
xor XOR2 (N2472, N2465, N1251);
nand NAND3 (N2473, N2454, N245, N1050);
or OR4 (N2474, N2471, N1581, N532, N1577);
not NOT1 (N2475, N2469);
nor NOR2 (N2476, N2474, N1653);
or OR3 (N2477, N2470, N353, N856);
nand NAND2 (N2478, N2472, N517);
nand NAND2 (N2479, N2461, N722);
nand NAND3 (N2480, N2475, N1463, N1558);
xor XOR2 (N2481, N2467, N1305);
nand NAND4 (N2482, N2458, N139, N111, N1389);
xor XOR2 (N2483, N2460, N1911);
and AND2 (N2484, N2473, N1475);
and AND3 (N2485, N2484, N2120, N2118);
buf BUF1 (N2486, N2483);
not NOT1 (N2487, N2477);
nor NOR3 (N2488, N2481, N2068, N1715);
nor NOR3 (N2489, N2485, N2300, N896);
and AND2 (N2490, N2479, N1549);
nor NOR4 (N2491, N2480, N1185, N1356, N940);
or OR3 (N2492, N2482, N361, N1352);
buf BUF1 (N2493, N2486);
xor XOR2 (N2494, N2488, N1710);
buf BUF1 (N2495, N2478);
nand NAND4 (N2496, N2476, N347, N2487, N548);
not NOT1 (N2497, N1210);
buf BUF1 (N2498, N2494);
xor XOR2 (N2499, N2491, N1661);
not NOT1 (N2500, N2489);
nand NAND3 (N2501, N2497, N640, N785);
and AND2 (N2502, N2500, N1173);
xor XOR2 (N2503, N2498, N1212);
xor XOR2 (N2504, N2490, N1371);
buf BUF1 (N2505, N2504);
nor NOR4 (N2506, N2502, N413, N724, N586);
and AND4 (N2507, N2503, N2195, N1680, N1832);
nor NOR3 (N2508, N2493, N2447, N72);
not NOT1 (N2509, N2505);
nor NOR2 (N2510, N2507, N1616);
xor XOR2 (N2511, N2506, N1185);
xor XOR2 (N2512, N2509, N2166);
or OR3 (N2513, N2492, N1651, N353);
xor XOR2 (N2514, N2495, N2313);
not NOT1 (N2515, N2513);
not NOT1 (N2516, N2499);
xor XOR2 (N2517, N2511, N2242);
not NOT1 (N2518, N2501);
buf BUF1 (N2519, N2515);
and AND2 (N2520, N2519, N247);
not NOT1 (N2521, N2508);
buf BUF1 (N2522, N2520);
xor XOR2 (N2523, N2522, N2009);
not NOT1 (N2524, N2516);
nand NAND3 (N2525, N2521, N1545, N1070);
nor NOR2 (N2526, N2510, N1026);
xor XOR2 (N2527, N2518, N137);
nor NOR4 (N2528, N2410, N613, N759, N935);
nor NOR4 (N2529, N2514, N708, N1922, N710);
not NOT1 (N2530, N2528);
nand NAND3 (N2531, N2496, N1727, N1551);
or OR4 (N2532, N2517, N394, N1337, N53);
not NOT1 (N2533, N2526);
not NOT1 (N2534, N2533);
xor XOR2 (N2535, N2532, N978);
buf BUF1 (N2536, N2529);
nor NOR2 (N2537, N2534, N1953);
nand NAND2 (N2538, N2524, N1149);
xor XOR2 (N2539, N2538, N2232);
not NOT1 (N2540, N2535);
nand NAND3 (N2541, N2530, N7, N129);
nor NOR3 (N2542, N2539, N1561, N2350);
not NOT1 (N2543, N2542);
nor NOR4 (N2544, N2523, N876, N1592, N810);
buf BUF1 (N2545, N2540);
xor XOR2 (N2546, N2541, N2406);
buf BUF1 (N2547, N2544);
nor NOR2 (N2548, N2545, N2135);
nand NAND4 (N2549, N2548, N1374, N2391, N924);
nand NAND4 (N2550, N2537, N1096, N1902, N2436);
xor XOR2 (N2551, N2512, N698);
not NOT1 (N2552, N2551);
or OR2 (N2553, N2550, N1732);
and AND3 (N2554, N2531, N618, N296);
nand NAND4 (N2555, N2554, N1974, N2006, N1458);
and AND4 (N2556, N2555, N525, N1296, N1665);
nand NAND4 (N2557, N2543, N1726, N2071, N890);
nand NAND2 (N2558, N2536, N1043);
nor NOR4 (N2559, N2557, N2368, N2276, N504);
xor XOR2 (N2560, N2559, N954);
nand NAND2 (N2561, N2525, N2152);
xor XOR2 (N2562, N2553, N1635);
xor XOR2 (N2563, N2560, N1084);
and AND2 (N2564, N2527, N681);
xor XOR2 (N2565, N2549, N1359);
and AND2 (N2566, N2558, N1599);
xor XOR2 (N2567, N2561, N2356);
xor XOR2 (N2568, N2546, N905);
nand NAND4 (N2569, N2562, N1197, N1920, N2014);
nor NOR4 (N2570, N2569, N310, N52, N211);
not NOT1 (N2571, N2564);
buf BUF1 (N2572, N2547);
not NOT1 (N2573, N2568);
xor XOR2 (N2574, N2567, N2126);
nor NOR3 (N2575, N2570, N1314, N1157);
nand NAND4 (N2576, N2565, N1572, N1561, N2171);
buf BUF1 (N2577, N2563);
or OR4 (N2578, N2572, N1899, N1102, N437);
xor XOR2 (N2579, N2571, N172);
and AND3 (N2580, N2579, N1054, N871);
and AND3 (N2581, N2556, N1851, N1287);
not NOT1 (N2582, N2573);
nand NAND2 (N2583, N2577, N2007);
and AND3 (N2584, N2552, N1433, N1521);
not NOT1 (N2585, N2574);
buf BUF1 (N2586, N2566);
nand NAND3 (N2587, N2582, N1498, N1080);
nand NAND2 (N2588, N2586, N1961);
buf BUF1 (N2589, N2580);
xor XOR2 (N2590, N2584, N46);
or OR4 (N2591, N2578, N114, N1911, N529);
nor NOR4 (N2592, N2587, N596, N726, N663);
buf BUF1 (N2593, N2575);
xor XOR2 (N2594, N2576, N1524);
and AND3 (N2595, N2589, N2197, N1240);
and AND2 (N2596, N2590, N1587);
or OR4 (N2597, N2583, N1762, N1213, N132);
or OR3 (N2598, N2594, N1577, N1633);
or OR2 (N2599, N2598, N1253);
nor NOR2 (N2600, N2593, N2176);
buf BUF1 (N2601, N2595);
nand NAND3 (N2602, N2599, N1766, N2452);
buf BUF1 (N2603, N2585);
and AND3 (N2604, N2591, N1643, N2538);
not NOT1 (N2605, N2588);
nand NAND3 (N2606, N2592, N704, N964);
not NOT1 (N2607, N2605);
and AND2 (N2608, N2600, N1586);
xor XOR2 (N2609, N2602, N1178);
buf BUF1 (N2610, N2597);
buf BUF1 (N2611, N2610);
nand NAND2 (N2612, N2596, N2190);
nand NAND4 (N2613, N2604, N797, N438, N1881);
xor XOR2 (N2614, N2613, N1282);
buf BUF1 (N2615, N2614);
or OR2 (N2616, N2606, N2292);
or OR3 (N2617, N2609, N823, N311);
and AND3 (N2618, N2615, N1400, N1220);
not NOT1 (N2619, N2601);
nor NOR3 (N2620, N2608, N2021, N1741);
or OR4 (N2621, N2607, N2537, N245, N389);
nor NOR3 (N2622, N2619, N2090, N2287);
nor NOR2 (N2623, N2616, N321);
or OR4 (N2624, N2618, N2065, N2037, N1980);
xor XOR2 (N2625, N2612, N129);
buf BUF1 (N2626, N2617);
buf BUF1 (N2627, N2622);
nor NOR3 (N2628, N2625, N2276, N1476);
buf BUF1 (N2629, N2611);
xor XOR2 (N2630, N2626, N577);
buf BUF1 (N2631, N2623);
and AND4 (N2632, N2631, N1575, N1837, N2427);
or OR3 (N2633, N2632, N698, N1347);
and AND4 (N2634, N2629, N881, N1643, N1219);
and AND2 (N2635, N2627, N1089);
and AND4 (N2636, N2581, N364, N370, N1460);
xor XOR2 (N2637, N2628, N643);
nand NAND3 (N2638, N2634, N528, N2384);
not NOT1 (N2639, N2603);
or OR4 (N2640, N2624, N1126, N2104, N2580);
xor XOR2 (N2641, N2621, N1925);
or OR3 (N2642, N2640, N2320, N2248);
not NOT1 (N2643, N2636);
buf BUF1 (N2644, N2641);
buf BUF1 (N2645, N2635);
xor XOR2 (N2646, N2644, N742);
nand NAND3 (N2647, N2646, N1598, N558);
nor NOR3 (N2648, N2639, N1171, N1734);
or OR3 (N2649, N2620, N1859, N927);
and AND3 (N2650, N2642, N2368, N1506);
nand NAND3 (N2651, N2645, N1592, N428);
or OR4 (N2652, N2651, N13, N199, N1181);
not NOT1 (N2653, N2649);
nand NAND2 (N2654, N2643, N31);
buf BUF1 (N2655, N2654);
nor NOR3 (N2656, N2630, N1921, N2544);
buf BUF1 (N2657, N2648);
and AND3 (N2658, N2650, N2365, N417);
nand NAND3 (N2659, N2655, N621, N2293);
xor XOR2 (N2660, N2653, N887);
and AND3 (N2661, N2658, N1137, N2582);
buf BUF1 (N2662, N2638);
not NOT1 (N2663, N2637);
xor XOR2 (N2664, N2652, N2066);
nor NOR2 (N2665, N2656, N2160);
or OR3 (N2666, N2660, N2427, N2047);
and AND4 (N2667, N2659, N2168, N931, N2484);
or OR3 (N2668, N2657, N669, N2136);
buf BUF1 (N2669, N2647);
or OR2 (N2670, N2664, N802);
and AND2 (N2671, N2665, N1203);
and AND2 (N2672, N2669, N559);
buf BUF1 (N2673, N2661);
buf BUF1 (N2674, N2662);
buf BUF1 (N2675, N2670);
and AND3 (N2676, N2666, N588, N1786);
or OR4 (N2677, N2675, N1046, N698, N939);
nand NAND3 (N2678, N2668, N708, N10);
and AND4 (N2679, N2667, N1325, N2596, N291);
or OR3 (N2680, N2678, N789, N2030);
nor NOR2 (N2681, N2680, N179);
not NOT1 (N2682, N2671);
buf BUF1 (N2683, N2673);
buf BUF1 (N2684, N2681);
nand NAND3 (N2685, N2682, N2000, N903);
or OR2 (N2686, N2672, N361);
nor NOR4 (N2687, N2674, N2648, N1358, N1506);
not NOT1 (N2688, N2633);
not NOT1 (N2689, N2688);
nor NOR2 (N2690, N2676, N415);
xor XOR2 (N2691, N2677, N1462);
or OR3 (N2692, N2683, N2086, N1523);
buf BUF1 (N2693, N2684);
xor XOR2 (N2694, N2685, N1789);
nor NOR3 (N2695, N2691, N553, N1972);
xor XOR2 (N2696, N2695, N618);
nand NAND3 (N2697, N2689, N318, N2508);
or OR4 (N2698, N2693, N732, N890, N589);
nor NOR4 (N2699, N2687, N1108, N838, N508);
xor XOR2 (N2700, N2696, N700);
nor NOR2 (N2701, N2700, N2474);
nor NOR2 (N2702, N2692, N1719);
or OR3 (N2703, N2698, N2389, N1302);
nand NAND4 (N2704, N2699, N1903, N1760, N1136);
nand NAND4 (N2705, N2663, N1272, N1116, N1145);
or OR2 (N2706, N2701, N2465);
nor NOR2 (N2707, N2704, N2337);
or OR4 (N2708, N2707, N2006, N28, N634);
xor XOR2 (N2709, N2708, N777);
or OR2 (N2710, N2703, N1949);
and AND3 (N2711, N2706, N710, N932);
xor XOR2 (N2712, N2711, N1278);
nand NAND3 (N2713, N2705, N1394, N1362);
not NOT1 (N2714, N2713);
and AND3 (N2715, N2697, N580, N1439);
nor NOR3 (N2716, N2690, N2407, N1733);
or OR4 (N2717, N2694, N1540, N2069, N1904);
not NOT1 (N2718, N2709);
buf BUF1 (N2719, N2679);
and AND3 (N2720, N2702, N1390, N1944);
xor XOR2 (N2721, N2714, N1722);
buf BUF1 (N2722, N2719);
buf BUF1 (N2723, N2720);
xor XOR2 (N2724, N2722, N863);
xor XOR2 (N2725, N2715, N1766);
nand NAND4 (N2726, N2712, N2428, N976, N913);
and AND3 (N2727, N2723, N666, N2388);
and AND4 (N2728, N2725, N880, N679, N1360);
and AND2 (N2729, N2727, N2186);
nor NOR4 (N2730, N2717, N1044, N2652, N492);
or OR2 (N2731, N2726, N1807);
nand NAND2 (N2732, N2718, N2344);
nor NOR4 (N2733, N2729, N1365, N1824, N886);
nand NAND3 (N2734, N2733, N2488, N110);
nand NAND4 (N2735, N2730, N2003, N1981, N696);
nor NOR3 (N2736, N2716, N632, N288);
or OR2 (N2737, N2736, N2290);
nand NAND2 (N2738, N2731, N1793);
nor NOR3 (N2739, N2710, N182, N770);
xor XOR2 (N2740, N2737, N164);
nor NOR2 (N2741, N2739, N62);
not NOT1 (N2742, N2735);
not NOT1 (N2743, N2721);
nor NOR2 (N2744, N2740, N2378);
xor XOR2 (N2745, N2724, N1405);
nor NOR3 (N2746, N2742, N371, N1090);
xor XOR2 (N2747, N2728, N1868);
or OR2 (N2748, N2738, N150);
not NOT1 (N2749, N2686);
buf BUF1 (N2750, N2743);
and AND2 (N2751, N2750, N1752);
xor XOR2 (N2752, N2741, N1496);
not NOT1 (N2753, N2747);
or OR2 (N2754, N2745, N2);
nand NAND2 (N2755, N2746, N265);
xor XOR2 (N2756, N2753, N1068);
not NOT1 (N2757, N2732);
nor NOR3 (N2758, N2756, N1320, N1559);
nor NOR3 (N2759, N2752, N1500, N2742);
nand NAND4 (N2760, N2744, N2479, N2670, N2151);
buf BUF1 (N2761, N2758);
or OR3 (N2762, N2751, N2118, N1779);
xor XOR2 (N2763, N2748, N701);
and AND4 (N2764, N2754, N1235, N1923, N362);
and AND2 (N2765, N2749, N1294);
xor XOR2 (N2766, N2734, N1661);
or OR4 (N2767, N2761, N113, N1979, N1014);
buf BUF1 (N2768, N2762);
xor XOR2 (N2769, N2759, N791);
xor XOR2 (N2770, N2767, N1908);
or OR4 (N2771, N2763, N1429, N1962, N2468);
not NOT1 (N2772, N2769);
nand NAND3 (N2773, N2766, N472, N791);
not NOT1 (N2774, N2757);
and AND2 (N2775, N2760, N1577);
nor NOR3 (N2776, N2770, N668, N1554);
or OR4 (N2777, N2776, N1019, N1184, N1575);
nor NOR2 (N2778, N2755, N2094);
and AND3 (N2779, N2771, N2114, N2146);
xor XOR2 (N2780, N2773, N1470);
nand NAND3 (N2781, N2778, N2280, N1913);
and AND2 (N2782, N2768, N1561);
or OR3 (N2783, N2781, N384, N1229);
buf BUF1 (N2784, N2777);
not NOT1 (N2785, N2772);
and AND3 (N2786, N2782, N209, N935);
and AND2 (N2787, N2780, N221);
nor NOR3 (N2788, N2786, N933, N2446);
buf BUF1 (N2789, N2783);
nand NAND4 (N2790, N2774, N713, N2567, N843);
buf BUF1 (N2791, N2779);
buf BUF1 (N2792, N2789);
xor XOR2 (N2793, N2790, N902);
not NOT1 (N2794, N2792);
buf BUF1 (N2795, N2784);
xor XOR2 (N2796, N2795, N1830);
buf BUF1 (N2797, N2796);
nor NOR3 (N2798, N2788, N642, N1684);
or OR3 (N2799, N2793, N333, N486);
buf BUF1 (N2800, N2798);
buf BUF1 (N2801, N2799);
nand NAND2 (N2802, N2797, N1689);
buf BUF1 (N2803, N2775);
or OR2 (N2804, N2785, N748);
buf BUF1 (N2805, N2804);
buf BUF1 (N2806, N2765);
buf BUF1 (N2807, N2800);
nand NAND2 (N2808, N2787, N311);
not NOT1 (N2809, N2794);
nor NOR4 (N2810, N2801, N310, N554, N1018);
and AND4 (N2811, N2808, N41, N1582, N952);
xor XOR2 (N2812, N2802, N539);
nand NAND4 (N2813, N2810, N1142, N2153, N2280);
nor NOR3 (N2814, N2764, N781, N1628);
nor NOR2 (N2815, N2791, N1640);
xor XOR2 (N2816, N2815, N371);
nand NAND3 (N2817, N2806, N1839, N1420);
buf BUF1 (N2818, N2814);
not NOT1 (N2819, N2813);
buf BUF1 (N2820, N2809);
xor XOR2 (N2821, N2812, N2029);
and AND3 (N2822, N2819, N1373, N574);
not NOT1 (N2823, N2817);
or OR3 (N2824, N2805, N2531, N119);
nor NOR2 (N2825, N2824, N1341);
nor NOR2 (N2826, N2820, N853);
nand NAND4 (N2827, N2823, N132, N467, N2617);
not NOT1 (N2828, N2816);
nand NAND3 (N2829, N2807, N254, N1640);
or OR3 (N2830, N2818, N1047, N1336);
and AND2 (N2831, N2803, N1417);
and AND4 (N2832, N2831, N535, N1267, N2119);
or OR2 (N2833, N2828, N2309);
or OR4 (N2834, N2830, N2592, N2495, N339);
buf BUF1 (N2835, N2829);
buf BUF1 (N2836, N2825);
nor NOR4 (N2837, N2822, N966, N48, N1027);
and AND4 (N2838, N2833, N1154, N1177, N456);
xor XOR2 (N2839, N2827, N1301);
not NOT1 (N2840, N2839);
xor XOR2 (N2841, N2834, N98);
and AND4 (N2842, N2835, N2717, N282, N2549);
or OR2 (N2843, N2821, N1863);
xor XOR2 (N2844, N2843, N857);
xor XOR2 (N2845, N2838, N1613);
nor NOR2 (N2846, N2837, N665);
nand NAND4 (N2847, N2846, N1836, N1188, N2255);
xor XOR2 (N2848, N2841, N345);
not NOT1 (N2849, N2832);
and AND4 (N2850, N2845, N287, N1541, N259);
and AND2 (N2851, N2811, N1678);
and AND4 (N2852, N2842, N1446, N2025, N2725);
not NOT1 (N2853, N2848);
nor NOR4 (N2854, N2840, N608, N339, N2705);
buf BUF1 (N2855, N2854);
or OR3 (N2856, N2826, N1031, N1186);
buf BUF1 (N2857, N2847);
nand NAND3 (N2858, N2852, N2573, N2525);
nor NOR3 (N2859, N2851, N623, N651);
or OR3 (N2860, N2836, N895, N1440);
nor NOR3 (N2861, N2853, N988, N1994);
nor NOR4 (N2862, N2857, N2432, N1621, N2664);
or OR2 (N2863, N2859, N761);
nand NAND3 (N2864, N2861, N835, N959);
and AND3 (N2865, N2860, N1977, N281);
or OR3 (N2866, N2850, N821, N107);
nand NAND4 (N2867, N2849, N686, N186, N355);
buf BUF1 (N2868, N2856);
nor NOR2 (N2869, N2866, N1995);
buf BUF1 (N2870, N2867);
nor NOR3 (N2871, N2844, N2382, N2675);
xor XOR2 (N2872, N2870, N2810);
nor NOR2 (N2873, N2872, N2724);
nand NAND2 (N2874, N2862, N1772);
not NOT1 (N2875, N2871);
nand NAND3 (N2876, N2875, N1771, N915);
xor XOR2 (N2877, N2855, N786);
not NOT1 (N2878, N2858);
not NOT1 (N2879, N2874);
and AND3 (N2880, N2878, N2542, N247);
and AND3 (N2881, N2873, N2390, N2420);
and AND4 (N2882, N2881, N45, N188, N1756);
nor NOR3 (N2883, N2869, N2240, N756);
or OR2 (N2884, N2880, N1493);
buf BUF1 (N2885, N2877);
or OR2 (N2886, N2865, N1372);
not NOT1 (N2887, N2864);
nor NOR2 (N2888, N2882, N2476);
and AND3 (N2889, N2888, N2073, N1624);
nor NOR2 (N2890, N2883, N813);
nor NOR3 (N2891, N2884, N993, N1448);
buf BUF1 (N2892, N2887);
or OR4 (N2893, N2889, N2317, N1676, N417);
not NOT1 (N2894, N2868);
xor XOR2 (N2895, N2892, N2803);
or OR2 (N2896, N2886, N1667);
xor XOR2 (N2897, N2885, N485);
nor NOR3 (N2898, N2897, N402, N2545);
nand NAND4 (N2899, N2896, N1351, N1777, N1329);
nand NAND4 (N2900, N2876, N363, N2097, N727);
buf BUF1 (N2901, N2898);
not NOT1 (N2902, N2900);
nor NOR3 (N2903, N2863, N772, N1887);
or OR2 (N2904, N2902, N1363);
or OR2 (N2905, N2901, N1715);
or OR4 (N2906, N2893, N2117, N2007, N1492);
xor XOR2 (N2907, N2895, N1812);
nor NOR2 (N2908, N2903, N2319);
or OR4 (N2909, N2894, N424, N210, N1406);
xor XOR2 (N2910, N2890, N276);
or OR4 (N2911, N2906, N2328, N1240, N1134);
buf BUF1 (N2912, N2910);
nand NAND2 (N2913, N2879, N2189);
and AND4 (N2914, N2909, N2470, N2501, N1519);
not NOT1 (N2915, N2912);
not NOT1 (N2916, N2904);
nor NOR2 (N2917, N2907, N2131);
nor NOR4 (N2918, N2914, N2441, N543, N1484);
buf BUF1 (N2919, N2913);
nand NAND4 (N2920, N2905, N2436, N1777, N2591);
nor NOR4 (N2921, N2908, N1094, N710, N1197);
not NOT1 (N2922, N2921);
nor NOR2 (N2923, N2918, N1960);
buf BUF1 (N2924, N2911);
buf BUF1 (N2925, N2891);
nand NAND2 (N2926, N2916, N487);
and AND3 (N2927, N2925, N530, N1909);
buf BUF1 (N2928, N2899);
buf BUF1 (N2929, N2915);
not NOT1 (N2930, N2927);
or OR4 (N2931, N2930, N1103, N308, N1680);
nor NOR2 (N2932, N2928, N2053);
or OR3 (N2933, N2923, N2625, N464);
xor XOR2 (N2934, N2922, N2480);
nor NOR2 (N2935, N2919, N1682);
or OR4 (N2936, N2932, N2528, N2832, N776);
buf BUF1 (N2937, N2931);
nor NOR3 (N2938, N2936, N2839, N2197);
nand NAND3 (N2939, N2937, N1090, N2621);
or OR4 (N2940, N2939, N1316, N1544, N562);
buf BUF1 (N2941, N2917);
or OR2 (N2942, N2941, N1430);
nand NAND3 (N2943, N2942, N2813, N319);
nor NOR2 (N2944, N2929, N1638);
or OR4 (N2945, N2920, N995, N765, N1066);
xor XOR2 (N2946, N2944, N1692);
not NOT1 (N2947, N2934);
nand NAND2 (N2948, N2935, N2583);
nor NOR4 (N2949, N2938, N425, N761, N1809);
not NOT1 (N2950, N2933);
not NOT1 (N2951, N2945);
buf BUF1 (N2952, N2924);
nor NOR2 (N2953, N2952, N1962);
buf BUF1 (N2954, N2946);
not NOT1 (N2955, N2943);
and AND3 (N2956, N2926, N431, N2765);
xor XOR2 (N2957, N2954, N2477);
xor XOR2 (N2958, N2951, N814);
not NOT1 (N2959, N2956);
or OR2 (N2960, N2955, N2636);
nand NAND3 (N2961, N2947, N133, N2872);
nand NAND3 (N2962, N2958, N2820, N1690);
and AND2 (N2963, N2949, N2936);
buf BUF1 (N2964, N2948);
and AND2 (N2965, N2953, N1867);
not NOT1 (N2966, N2940);
and AND2 (N2967, N2959, N1608);
nor NOR3 (N2968, N2961, N169, N2321);
and AND3 (N2969, N2964, N129, N262);
xor XOR2 (N2970, N2963, N2467);
nor NOR2 (N2971, N2967, N2211);
nor NOR2 (N2972, N2969, N725);
nand NAND3 (N2973, N2971, N790, N1760);
and AND3 (N2974, N2957, N857, N71);
and AND3 (N2975, N2966, N1271, N306);
not NOT1 (N2976, N2950);
nand NAND2 (N2977, N2965, N1855);
nor NOR4 (N2978, N2970, N979, N2145, N756);
nor NOR2 (N2979, N2960, N2213);
buf BUF1 (N2980, N2972);
or OR4 (N2981, N2977, N2266, N2750, N2165);
xor XOR2 (N2982, N2981, N284);
nor NOR3 (N2983, N2962, N657, N2341);
or OR3 (N2984, N2978, N545, N1097);
nand NAND3 (N2985, N2982, N1327, N2648);
or OR4 (N2986, N2979, N1433, N845, N596);
nand NAND4 (N2987, N2974, N1047, N1491, N573);
and AND4 (N2988, N2973, N2833, N260, N1017);
not NOT1 (N2989, N2976);
and AND3 (N2990, N2985, N925, N2819);
not NOT1 (N2991, N2986);
xor XOR2 (N2992, N2991, N2747);
xor XOR2 (N2993, N2987, N1155);
and AND3 (N2994, N2983, N470, N677);
nand NAND4 (N2995, N2990, N1278, N2372, N2191);
xor XOR2 (N2996, N2980, N2555);
or OR4 (N2997, N2975, N1022, N2868, N335);
not NOT1 (N2998, N2989);
or OR4 (N2999, N2998, N1660, N2484, N781);
and AND2 (N3000, N2994, N2148);
not NOT1 (N3001, N2999);
nand NAND2 (N3002, N3001, N126);
xor XOR2 (N3003, N3000, N285);
buf BUF1 (N3004, N2993);
not NOT1 (N3005, N2996);
and AND3 (N3006, N2984, N1254, N802);
xor XOR2 (N3007, N2992, N962);
nand NAND3 (N3008, N3002, N591, N2144);
nand NAND3 (N3009, N2968, N2998, N384);
xor XOR2 (N3010, N2997, N601);
and AND2 (N3011, N2988, N661);
xor XOR2 (N3012, N3005, N1293);
or OR2 (N3013, N3003, N396);
buf BUF1 (N3014, N3009);
nor NOR4 (N3015, N3004, N1040, N2220, N952);
xor XOR2 (N3016, N3012, N15);
nand NAND4 (N3017, N3015, N2365, N1786, N640);
nand NAND3 (N3018, N3016, N1196, N1708);
not NOT1 (N3019, N3008);
nand NAND3 (N3020, N3007, N1183, N670);
nor NOR3 (N3021, N3020, N1745, N1150);
nand NAND4 (N3022, N3019, N2443, N520, N2032);
xor XOR2 (N3023, N3006, N2771);
xor XOR2 (N3024, N3023, N415);
buf BUF1 (N3025, N3014);
buf BUF1 (N3026, N3010);
buf BUF1 (N3027, N3024);
xor XOR2 (N3028, N3022, N1500);
xor XOR2 (N3029, N3018, N2796);
or OR4 (N3030, N3027, N1352, N573, N1291);
buf BUF1 (N3031, N3017);
nand NAND3 (N3032, N2995, N2560, N1662);
and AND3 (N3033, N3031, N1738, N2293);
not NOT1 (N3034, N3028);
buf BUF1 (N3035, N3032);
buf BUF1 (N3036, N3026);
nor NOR2 (N3037, N3025, N1997);
nand NAND2 (N3038, N3029, N2998);
not NOT1 (N3039, N3030);
xor XOR2 (N3040, N3034, N2666);
nand NAND4 (N3041, N3037, N1225, N144, N2529);
not NOT1 (N3042, N3013);
buf BUF1 (N3043, N3033);
buf BUF1 (N3044, N3035);
not NOT1 (N3045, N3011);
not NOT1 (N3046, N3044);
and AND3 (N3047, N3036, N1602, N2670);
xor XOR2 (N3048, N3043, N2765);
or OR3 (N3049, N3040, N560, N1588);
and AND4 (N3050, N3038, N621, N1145, N2831);
not NOT1 (N3051, N3045);
nand NAND4 (N3052, N3048, N1077, N613, N1390);
and AND4 (N3053, N3046, N1266, N977, N316);
xor XOR2 (N3054, N3047, N1855);
xor XOR2 (N3055, N3052, N1466);
and AND3 (N3056, N3041, N1102, N2936);
or OR4 (N3057, N3021, N2935, N2285, N841);
buf BUF1 (N3058, N3042);
or OR4 (N3059, N3058, N1801, N941, N2133);
nand NAND2 (N3060, N3053, N365);
xor XOR2 (N3061, N3049, N3024);
and AND2 (N3062, N3061, N1710);
or OR4 (N3063, N3050, N2334, N2997, N2456);
nor NOR2 (N3064, N3055, N383);
and AND2 (N3065, N3056, N2929);
and AND2 (N3066, N3039, N2806);
not NOT1 (N3067, N3063);
nor NOR3 (N3068, N3054, N1329, N1059);
nor NOR3 (N3069, N3059, N158, N2908);
nand NAND3 (N3070, N3068, N2511, N1620);
nor NOR3 (N3071, N3069, N866, N384);
buf BUF1 (N3072, N3060);
xor XOR2 (N3073, N3065, N1888);
nand NAND2 (N3074, N3070, N1408);
or OR4 (N3075, N3064, N303, N2658, N2048);
not NOT1 (N3076, N3073);
nand NAND4 (N3077, N3062, N376, N2124, N1195);
not NOT1 (N3078, N3072);
not NOT1 (N3079, N3077);
and AND4 (N3080, N3076, N1702, N1782, N2283);
nand NAND2 (N3081, N3080, N513);
buf BUF1 (N3082, N3067);
or OR4 (N3083, N3051, N1264, N1390, N189);
or OR2 (N3084, N3074, N1673);
nand NAND3 (N3085, N3057, N758, N1103);
nor NOR2 (N3086, N3079, N2350);
xor XOR2 (N3087, N3075, N1344);
and AND4 (N3088, N3087, N2908, N1036, N2252);
xor XOR2 (N3089, N3083, N468);
and AND4 (N3090, N3078, N1708, N362, N1664);
and AND3 (N3091, N3084, N1412, N3047);
and AND4 (N3092, N3085, N761, N1799, N2551);
or OR2 (N3093, N3092, N321);
and AND3 (N3094, N3082, N1540, N2321);
and AND3 (N3095, N3071, N894, N2175);
or OR2 (N3096, N3093, N1386);
buf BUF1 (N3097, N3091);
not NOT1 (N3098, N3096);
nand NAND2 (N3099, N3066, N857);
nand NAND4 (N3100, N3088, N1224, N978, N2635);
or OR4 (N3101, N3086, N2875, N1338, N2979);
nor NOR3 (N3102, N3081, N1362, N249);
or OR2 (N3103, N3095, N1848);
buf BUF1 (N3104, N3089);
nand NAND3 (N3105, N3101, N1792, N1645);
not NOT1 (N3106, N3102);
not NOT1 (N3107, N3103);
nand NAND3 (N3108, N3097, N1434, N635);
and AND4 (N3109, N3105, N588, N1861, N2777);
or OR2 (N3110, N3098, N1480);
not NOT1 (N3111, N3104);
xor XOR2 (N3112, N3111, N530);
nor NOR4 (N3113, N3100, N639, N141, N394);
not NOT1 (N3114, N3109);
or OR4 (N3115, N3113, N1631, N1145, N1671);
xor XOR2 (N3116, N3090, N1684);
and AND2 (N3117, N3115, N2402);
not NOT1 (N3118, N3094);
and AND2 (N3119, N3117, N1747);
nor NOR4 (N3120, N3108, N2113, N2886, N3037);
buf BUF1 (N3121, N3107);
xor XOR2 (N3122, N3118, N246);
or OR4 (N3123, N3112, N2218, N1177, N2101);
not NOT1 (N3124, N3122);
xor XOR2 (N3125, N3116, N458);
buf BUF1 (N3126, N3123);
xor XOR2 (N3127, N3099, N1373);
not NOT1 (N3128, N3124);
nand NAND2 (N3129, N3127, N2000);
nand NAND4 (N3130, N3129, N1771, N2118, N78);
or OR3 (N3131, N3126, N1833, N523);
buf BUF1 (N3132, N3121);
nand NAND3 (N3133, N3110, N2979, N1580);
xor XOR2 (N3134, N3132, N3131);
not NOT1 (N3135, N2272);
and AND4 (N3136, N3133, N1699, N99, N529);
not NOT1 (N3137, N3134);
and AND3 (N3138, N3119, N1270, N1623);
not NOT1 (N3139, N3114);
or OR4 (N3140, N3106, N1383, N2136, N1097);
and AND4 (N3141, N3140, N2812, N1051, N324);
or OR4 (N3142, N3128, N1183, N2258, N297);
nand NAND3 (N3143, N3141, N2888, N2234);
nand NAND3 (N3144, N3137, N1149, N2308);
not NOT1 (N3145, N3125);
or OR2 (N3146, N3120, N3038);
and AND4 (N3147, N3138, N1738, N2979, N866);
nor NOR2 (N3148, N3130, N136);
nand NAND2 (N3149, N3143, N2053);
or OR3 (N3150, N3142, N2376, N1063);
and AND3 (N3151, N3139, N2776, N954);
and AND2 (N3152, N3150, N2029);
not NOT1 (N3153, N3149);
xor XOR2 (N3154, N3153, N1141);
buf BUF1 (N3155, N3136);
and AND2 (N3156, N3155, N558);
and AND3 (N3157, N3156, N2512, N1002);
nand NAND4 (N3158, N3157, N2940, N2473, N154);
and AND3 (N3159, N3152, N979, N1249);
buf BUF1 (N3160, N3146);
and AND3 (N3161, N3151, N2774, N1216);
not NOT1 (N3162, N3154);
nor NOR2 (N3163, N3144, N1236);
buf BUF1 (N3164, N3161);
and AND3 (N3165, N3135, N2606, N886);
buf BUF1 (N3166, N3159);
xor XOR2 (N3167, N3166, N1398);
and AND2 (N3168, N3165, N2159);
nand NAND2 (N3169, N3160, N2999);
not NOT1 (N3170, N3158);
not NOT1 (N3171, N3164);
or OR4 (N3172, N3148, N1694, N2562, N2307);
buf BUF1 (N3173, N3145);
nand NAND3 (N3174, N3172, N2422, N2576);
or OR3 (N3175, N3162, N3051, N1896);
nor NOR4 (N3176, N3168, N1621, N3064, N999);
not NOT1 (N3177, N3170);
xor XOR2 (N3178, N3147, N2229);
xor XOR2 (N3179, N3174, N2493);
nand NAND3 (N3180, N3178, N1051, N360);
not NOT1 (N3181, N3176);
or OR3 (N3182, N3169, N2009, N746);
or OR3 (N3183, N3177, N1043, N368);
nand NAND3 (N3184, N3181, N657, N1497);
nand NAND2 (N3185, N3167, N2173);
nor NOR4 (N3186, N3185, N1054, N120, N1684);
and AND4 (N3187, N3186, N1958, N2369, N1453);
buf BUF1 (N3188, N3171);
and AND2 (N3189, N3184, N2255);
nand NAND4 (N3190, N3179, N3158, N2977, N589);
nor NOR3 (N3191, N3183, N48, N965);
nor NOR2 (N3192, N3163, N2235);
nor NOR4 (N3193, N3173, N517, N2435, N2589);
and AND3 (N3194, N3190, N63, N432);
xor XOR2 (N3195, N3194, N478);
buf BUF1 (N3196, N3195);
and AND4 (N3197, N3188, N1271, N881, N1809);
nor NOR2 (N3198, N3175, N2984);
nand NAND2 (N3199, N3198, N1387);
nand NAND4 (N3200, N3192, N1123, N1275, N2563);
xor XOR2 (N3201, N3200, N1119);
nand NAND4 (N3202, N3197, N126, N1944, N477);
xor XOR2 (N3203, N3202, N1989);
xor XOR2 (N3204, N3203, N676);
nor NOR2 (N3205, N3189, N2123);
xor XOR2 (N3206, N3205, N1543);
or OR2 (N3207, N3206, N722);
nand NAND2 (N3208, N3187, N2979);
not NOT1 (N3209, N3193);
and AND2 (N3210, N3180, N1156);
xor XOR2 (N3211, N3191, N2154);
or OR3 (N3212, N3182, N1119, N2298);
not NOT1 (N3213, N3207);
and AND3 (N3214, N3196, N630, N1453);
nand NAND2 (N3215, N3204, N2031);
and AND3 (N3216, N3209, N2751, N2435);
nor NOR4 (N3217, N3210, N1575, N304, N2606);
not NOT1 (N3218, N3201);
buf BUF1 (N3219, N3213);
not NOT1 (N3220, N3217);
xor XOR2 (N3221, N3219, N2896);
nand NAND2 (N3222, N3212, N3155);
nor NOR4 (N3223, N3214, N2147, N738, N3147);
xor XOR2 (N3224, N3222, N2726);
not NOT1 (N3225, N3220);
and AND2 (N3226, N3225, N2532);
and AND4 (N3227, N3226, N223, N3157, N2128);
buf BUF1 (N3228, N3224);
nand NAND2 (N3229, N3227, N1518);
or OR4 (N3230, N3216, N2199, N1198, N25);
and AND4 (N3231, N3211, N2581, N345, N644);
buf BUF1 (N3232, N3208);
or OR4 (N3233, N3229, N2017, N781, N578);
and AND4 (N3234, N3223, N2246, N1217, N595);
or OR2 (N3235, N3233, N2427);
and AND3 (N3236, N3221, N2412, N2555);
nand NAND2 (N3237, N3215, N124);
or OR4 (N3238, N3228, N2447, N1435, N839);
xor XOR2 (N3239, N3230, N532);
xor XOR2 (N3240, N3238, N2446);
or OR4 (N3241, N3239, N1903, N1493, N2293);
not NOT1 (N3242, N3218);
or OR4 (N3243, N3241, N2658, N1626, N1101);
not NOT1 (N3244, N3243);
buf BUF1 (N3245, N3242);
not NOT1 (N3246, N3231);
and AND2 (N3247, N3237, N2569);
or OR3 (N3248, N3234, N3093, N2483);
or OR2 (N3249, N3236, N2495);
not NOT1 (N3250, N3240);
not NOT1 (N3251, N3247);
and AND2 (N3252, N3232, N1786);
xor XOR2 (N3253, N3250, N1824);
xor XOR2 (N3254, N3244, N1837);
not NOT1 (N3255, N3199);
nand NAND4 (N3256, N3252, N1704, N2901, N2105);
not NOT1 (N3257, N3246);
nand NAND3 (N3258, N3254, N2300, N2616);
nand NAND3 (N3259, N3249, N302, N817);
xor XOR2 (N3260, N3235, N2208);
and AND2 (N3261, N3251, N3243);
nand NAND3 (N3262, N3258, N1371, N2967);
or OR2 (N3263, N3253, N1609);
xor XOR2 (N3264, N3257, N1314);
not NOT1 (N3265, N3263);
buf BUF1 (N3266, N3256);
or OR3 (N3267, N3265, N948, N1539);
xor XOR2 (N3268, N3266, N113);
buf BUF1 (N3269, N3245);
nand NAND3 (N3270, N3261, N2768, N3260);
or OR4 (N3271, N380, N581, N775, N1570);
and AND3 (N3272, N3270, N215, N1134);
nor NOR3 (N3273, N3267, N2773, N1858);
nand NAND3 (N3274, N3268, N803, N39);
buf BUF1 (N3275, N3274);
not NOT1 (N3276, N3275);
and AND4 (N3277, N3271, N369, N1428, N602);
or OR4 (N3278, N3255, N70, N2002, N3274);
nor NOR2 (N3279, N3272, N3156);
xor XOR2 (N3280, N3279, N1866);
xor XOR2 (N3281, N3264, N204);
not NOT1 (N3282, N3281);
not NOT1 (N3283, N3262);
nand NAND2 (N3284, N3280, N354);
nor NOR3 (N3285, N3273, N3034, N2582);
xor XOR2 (N3286, N3283, N304);
and AND2 (N3287, N3286, N548);
not NOT1 (N3288, N3287);
nand NAND3 (N3289, N3269, N2889, N1349);
nand NAND4 (N3290, N3284, N2232, N1532, N1891);
nor NOR2 (N3291, N3277, N1142);
xor XOR2 (N3292, N3248, N1516);
nor NOR4 (N3293, N3278, N881, N1704, N2624);
nand NAND4 (N3294, N3289, N659, N1439, N2183);
buf BUF1 (N3295, N3285);
xor XOR2 (N3296, N3276, N2975);
not NOT1 (N3297, N3291);
nor NOR4 (N3298, N3288, N1206, N2516, N976);
buf BUF1 (N3299, N3297);
buf BUF1 (N3300, N3296);
or OR2 (N3301, N3298, N755);
and AND4 (N3302, N3293, N1795, N2287, N1369);
and AND4 (N3303, N3259, N1602, N1320, N1606);
xor XOR2 (N3304, N3282, N1210);
not NOT1 (N3305, N3295);
or OR2 (N3306, N3305, N1645);
nor NOR4 (N3307, N3301, N1393, N1442, N1786);
and AND3 (N3308, N3300, N790, N1484);
or OR3 (N3309, N3303, N2923, N2721);
nand NAND2 (N3310, N3294, N413);
nand NAND4 (N3311, N3292, N1194, N1370, N1710);
and AND2 (N3312, N3299, N610);
not NOT1 (N3313, N3310);
or OR4 (N3314, N3306, N2548, N2607, N642);
xor XOR2 (N3315, N3290, N1893);
buf BUF1 (N3316, N3315);
not NOT1 (N3317, N3313);
not NOT1 (N3318, N3317);
xor XOR2 (N3319, N3311, N1705);
nor NOR4 (N3320, N3316, N1862, N582, N812);
not NOT1 (N3321, N3312);
buf BUF1 (N3322, N3302);
and AND2 (N3323, N3319, N400);
xor XOR2 (N3324, N3322, N1443);
or OR4 (N3325, N3321, N770, N1092, N1991);
nand NAND2 (N3326, N3323, N342);
not NOT1 (N3327, N3308);
not NOT1 (N3328, N3325);
or OR2 (N3329, N3307, N2342);
nand NAND4 (N3330, N3326, N557, N3101, N1185);
not NOT1 (N3331, N3304);
xor XOR2 (N3332, N3314, N433);
nand NAND3 (N3333, N3328, N1493, N269);
xor XOR2 (N3334, N3331, N2038);
buf BUF1 (N3335, N3309);
xor XOR2 (N3336, N3330, N1747);
buf BUF1 (N3337, N3332);
or OR3 (N3338, N3324, N280, N2918);
nand NAND3 (N3339, N3320, N2160, N2294);
or OR4 (N3340, N3329, N1935, N1242, N1670);
nor NOR3 (N3341, N3318, N2639, N2214);
nand NAND2 (N3342, N3340, N1222);
nor NOR4 (N3343, N3334, N893, N1737, N1065);
and AND4 (N3344, N3336, N123, N112, N1157);
or OR3 (N3345, N3339, N1948, N1779);
buf BUF1 (N3346, N3345);
and AND4 (N3347, N3342, N788, N784, N1769);
or OR3 (N3348, N3327, N1606, N213);
and AND3 (N3349, N3348, N2455, N2833);
buf BUF1 (N3350, N3341);
xor XOR2 (N3351, N3337, N2934);
and AND4 (N3352, N3346, N1457, N3290, N1938);
nor NOR3 (N3353, N3350, N1385, N3242);
xor XOR2 (N3354, N3349, N970);
not NOT1 (N3355, N3347);
and AND3 (N3356, N3351, N519, N610);
not NOT1 (N3357, N3352);
or OR4 (N3358, N3344, N3229, N1684, N2557);
not NOT1 (N3359, N3355);
xor XOR2 (N3360, N3357, N3051);
nand NAND2 (N3361, N3333, N3327);
nor NOR4 (N3362, N3356, N2726, N142, N2572);
buf BUF1 (N3363, N3358);
and AND2 (N3364, N3362, N2285);
buf BUF1 (N3365, N3343);
not NOT1 (N3366, N3365);
nor NOR2 (N3367, N3366, N522);
xor XOR2 (N3368, N3363, N1192);
nand NAND3 (N3369, N3368, N2512, N2049);
nor NOR2 (N3370, N3364, N1279);
nor NOR4 (N3371, N3338, N936, N3191, N3339);
and AND2 (N3372, N3359, N2266);
xor XOR2 (N3373, N3354, N2543);
buf BUF1 (N3374, N3367);
not NOT1 (N3375, N3335);
xor XOR2 (N3376, N3375, N368);
xor XOR2 (N3377, N3370, N2198);
and AND3 (N3378, N3376, N1832, N2432);
not NOT1 (N3379, N3378);
not NOT1 (N3380, N3379);
and AND4 (N3381, N3377, N3345, N1671, N2312);
nand NAND3 (N3382, N3374, N264, N652);
nor NOR2 (N3383, N3371, N1261);
xor XOR2 (N3384, N3381, N312);
buf BUF1 (N3385, N3384);
or OR3 (N3386, N3373, N1881, N2563);
or OR4 (N3387, N3382, N3250, N604, N2531);
buf BUF1 (N3388, N3380);
not NOT1 (N3389, N3369);
nand NAND3 (N3390, N3353, N1433, N2398);
nand NAND4 (N3391, N3386, N2880, N1033, N89);
and AND3 (N3392, N3387, N3329, N2327);
nand NAND2 (N3393, N3361, N3326);
nand NAND4 (N3394, N3393, N915, N428, N1638);
nor NOR3 (N3395, N3388, N1038, N1546);
nor NOR3 (N3396, N3360, N2290, N302);
nor NOR4 (N3397, N3392, N1960, N989, N1856);
not NOT1 (N3398, N3396);
or OR2 (N3399, N3383, N2850);
xor XOR2 (N3400, N3372, N760);
nand NAND3 (N3401, N3385, N2664, N193);
buf BUF1 (N3402, N3390);
or OR4 (N3403, N3395, N2970, N849, N3012);
nor NOR4 (N3404, N3391, N1643, N2299, N1045);
or OR4 (N3405, N3397, N1951, N2019, N1573);
xor XOR2 (N3406, N3402, N416);
or OR3 (N3407, N3405, N3324, N2622);
and AND3 (N3408, N3404, N416, N2595);
or OR2 (N3409, N3401, N3303);
and AND4 (N3410, N3389, N1672, N2506, N3016);
and AND2 (N3411, N3398, N453);
buf BUF1 (N3412, N3400);
nand NAND4 (N3413, N3399, N3364, N1526, N623);
not NOT1 (N3414, N3406);
or OR3 (N3415, N3411, N1445, N2152);
not NOT1 (N3416, N3414);
and AND4 (N3417, N3410, N755, N2391, N776);
nand NAND2 (N3418, N3413, N753);
nand NAND2 (N3419, N3408, N3319);
nor NOR2 (N3420, N3415, N212);
or OR3 (N3421, N3412, N1492, N371);
nand NAND4 (N3422, N3418, N2920, N1905, N1490);
buf BUF1 (N3423, N3416);
nor NOR4 (N3424, N3421, N3004, N848, N1020);
nand NAND4 (N3425, N3422, N2772, N2507, N1391);
not NOT1 (N3426, N3417);
xor XOR2 (N3427, N3420, N2749);
nor NOR4 (N3428, N3423, N3032, N2471, N82);
not NOT1 (N3429, N3427);
xor XOR2 (N3430, N3429, N1757);
nor NOR3 (N3431, N3409, N2405, N1469);
nor NOR2 (N3432, N3428, N221);
or OR2 (N3433, N3419, N1764);
nor NOR3 (N3434, N3433, N893, N68);
buf BUF1 (N3435, N3394);
buf BUF1 (N3436, N3407);
nor NOR4 (N3437, N3432, N480, N2615, N2906);
nand NAND2 (N3438, N3437, N956);
nand NAND3 (N3439, N3438, N1694, N1706);
or OR4 (N3440, N3425, N871, N2815, N1449);
nor NOR3 (N3441, N3434, N2233, N1514);
nor NOR3 (N3442, N3424, N1226, N1473);
nor NOR4 (N3443, N3431, N944, N1448, N609);
and AND4 (N3444, N3440, N1780, N3064, N2657);
nand NAND3 (N3445, N3430, N1879, N2706);
not NOT1 (N3446, N3445);
or OR4 (N3447, N3435, N2803, N3415, N853);
and AND2 (N3448, N3447, N2389);
or OR3 (N3449, N3426, N1018, N730);
or OR3 (N3450, N3443, N1252, N1311);
nor NOR4 (N3451, N3444, N2348, N2342, N608);
or OR2 (N3452, N3436, N2864);
nor NOR2 (N3453, N3452, N2200);
nor NOR4 (N3454, N3448, N631, N1607, N3241);
and AND4 (N3455, N3453, N489, N3134, N439);
nor NOR3 (N3456, N3446, N113, N423);
buf BUF1 (N3457, N3441);
and AND4 (N3458, N3403, N2462, N1345, N2263);
xor XOR2 (N3459, N3442, N2597);
and AND3 (N3460, N3455, N2018, N2638);
nand NAND4 (N3461, N3454, N2509, N2379, N1692);
not NOT1 (N3462, N3439);
buf BUF1 (N3463, N3456);
not NOT1 (N3464, N3463);
and AND2 (N3465, N3459, N2764);
buf BUF1 (N3466, N3458);
nand NAND3 (N3467, N3464, N225, N2114);
xor XOR2 (N3468, N3451, N3025);
or OR2 (N3469, N3465, N2654);
and AND2 (N3470, N3457, N1945);
buf BUF1 (N3471, N3461);
and AND4 (N3472, N3450, N884, N1199, N890);
buf BUF1 (N3473, N3471);
xor XOR2 (N3474, N3462, N1048);
not NOT1 (N3475, N3472);
xor XOR2 (N3476, N3466, N2591);
not NOT1 (N3477, N3474);
not NOT1 (N3478, N3460);
xor XOR2 (N3479, N3473, N3159);
buf BUF1 (N3480, N3470);
not NOT1 (N3481, N3469);
nor NOR2 (N3482, N3449, N2592);
xor XOR2 (N3483, N3468, N2579);
or OR3 (N3484, N3479, N2028, N2262);
buf BUF1 (N3485, N3482);
nand NAND3 (N3486, N3475, N1185, N2253);
buf BUF1 (N3487, N3478);
xor XOR2 (N3488, N3476, N2001);
nor NOR3 (N3489, N3480, N2386, N502);
xor XOR2 (N3490, N3477, N3399);
not NOT1 (N3491, N3490);
xor XOR2 (N3492, N3486, N2718);
and AND4 (N3493, N3491, N2193, N2151, N2384);
buf BUF1 (N3494, N3485);
not NOT1 (N3495, N3488);
nand NAND3 (N3496, N3494, N2383, N3381);
and AND3 (N3497, N3492, N963, N2058);
xor XOR2 (N3498, N3495, N1116);
nand NAND2 (N3499, N3484, N3464);
or OR3 (N3500, N3497, N1687, N3282);
or OR3 (N3501, N3496, N2899, N1811);
not NOT1 (N3502, N3500);
xor XOR2 (N3503, N3489, N3479);
buf BUF1 (N3504, N3498);
nand NAND2 (N3505, N3467, N551);
and AND4 (N3506, N3499, N1076, N634, N2234);
xor XOR2 (N3507, N3481, N2523);
nand NAND3 (N3508, N3506, N3487, N3444);
and AND4 (N3509, N1010, N1107, N2317, N1586);
and AND2 (N3510, N3508, N1457);
nand NAND4 (N3511, N3507, N3435, N517, N145);
nor NOR3 (N3512, N3501, N2408, N826);
xor XOR2 (N3513, N3493, N580);
nand NAND4 (N3514, N3504, N1021, N1302, N372);
nor NOR4 (N3515, N3503, N500, N76, N1374);
xor XOR2 (N3516, N3515, N202);
xor XOR2 (N3517, N3510, N367);
or OR2 (N3518, N3514, N2945);
nor NOR3 (N3519, N3509, N1949, N2639);
not NOT1 (N3520, N3512);
xor XOR2 (N3521, N3502, N2131);
buf BUF1 (N3522, N3519);
or OR2 (N3523, N3483, N782);
and AND4 (N3524, N3517, N819, N2114, N1961);
and AND2 (N3525, N3521, N3132);
not NOT1 (N3526, N3520);
nor NOR3 (N3527, N3505, N3122, N112);
and AND4 (N3528, N3523, N2470, N1353, N3002);
not NOT1 (N3529, N3511);
or OR2 (N3530, N3524, N1568);
nor NOR4 (N3531, N3516, N2477, N356, N2144);
nand NAND4 (N3532, N3526, N1098, N3027, N2923);
or OR2 (N3533, N3522, N3388);
xor XOR2 (N3534, N3532, N3290);
nand NAND3 (N3535, N3530, N1503, N291);
not NOT1 (N3536, N3531);
nand NAND3 (N3537, N3528, N1758, N672);
not NOT1 (N3538, N3529);
buf BUF1 (N3539, N3535);
or OR4 (N3540, N3513, N2345, N2066, N863);
or OR2 (N3541, N3527, N2547);
nor NOR2 (N3542, N3539, N241);
nor NOR3 (N3543, N3542, N1244, N1447);
nand NAND3 (N3544, N3525, N3508, N1242);
nor NOR4 (N3545, N3534, N1492, N1429, N768);
or OR2 (N3546, N3543, N3326);
nor NOR3 (N3547, N3545, N1559, N857);
not NOT1 (N3548, N3547);
not NOT1 (N3549, N3541);
not NOT1 (N3550, N3540);
buf BUF1 (N3551, N3549);
nor NOR3 (N3552, N3548, N2379, N33);
xor XOR2 (N3553, N3544, N1784);
or OR3 (N3554, N3518, N2213, N1534);
or OR2 (N3555, N3553, N684);
xor XOR2 (N3556, N3550, N770);
xor XOR2 (N3557, N3546, N1596);
or OR2 (N3558, N3557, N2681);
buf BUF1 (N3559, N3558);
buf BUF1 (N3560, N3536);
and AND3 (N3561, N3533, N2206, N3239);
nand NAND4 (N3562, N3537, N2129, N433, N2202);
or OR4 (N3563, N3552, N146, N1113, N772);
nor NOR3 (N3564, N3554, N538, N700);
or OR4 (N3565, N3559, N1216, N1601, N323);
xor XOR2 (N3566, N3562, N2880);
not NOT1 (N3567, N3561);
buf BUF1 (N3568, N3555);
and AND4 (N3569, N3567, N2625, N833, N1335);
and AND2 (N3570, N3556, N470);
buf BUF1 (N3571, N3538);
or OR3 (N3572, N3551, N2425, N1642);
buf BUF1 (N3573, N3564);
buf BUF1 (N3574, N3560);
nor NOR4 (N3575, N3568, N103, N3397, N1558);
or OR3 (N3576, N3571, N1220, N1355);
nand NAND4 (N3577, N3570, N2204, N2290, N3200);
nand NAND4 (N3578, N3575, N479, N373, N540);
buf BUF1 (N3579, N3569);
not NOT1 (N3580, N3574);
not NOT1 (N3581, N3576);
or OR2 (N3582, N3572, N1398);
nor NOR3 (N3583, N3565, N2797, N2462);
nand NAND4 (N3584, N3579, N3148, N2505, N965);
nand NAND2 (N3585, N3584, N3133);
or OR3 (N3586, N3585, N1277, N1012);
buf BUF1 (N3587, N3580);
not NOT1 (N3588, N3587);
buf BUF1 (N3589, N3563);
not NOT1 (N3590, N3578);
not NOT1 (N3591, N3586);
not NOT1 (N3592, N3591);
or OR4 (N3593, N3583, N942, N454, N2172);
or OR4 (N3594, N3592, N919, N402, N2556);
nor NOR4 (N3595, N3577, N2266, N1749, N2966);
not NOT1 (N3596, N3594);
nand NAND4 (N3597, N3588, N2860, N2022, N6);
or OR3 (N3598, N3589, N929, N1903);
and AND3 (N3599, N3598, N2363, N1158);
nor NOR2 (N3600, N3596, N3226);
buf BUF1 (N3601, N3590);
nand NAND3 (N3602, N3593, N3352, N2470);
and AND2 (N3603, N3602, N342);
nor NOR3 (N3604, N3566, N2952, N89);
not NOT1 (N3605, N3595);
nand NAND2 (N3606, N3599, N816);
and AND3 (N3607, N3603, N2157, N3092);
or OR2 (N3608, N3607, N58);
not NOT1 (N3609, N3601);
xor XOR2 (N3610, N3605, N3552);
and AND2 (N3611, N3604, N3341);
nor NOR4 (N3612, N3609, N238, N2864, N2771);
and AND4 (N3613, N3573, N1127, N2783, N900);
nor NOR2 (N3614, N3613, N1495);
xor XOR2 (N3615, N3606, N2939);
not NOT1 (N3616, N3610);
xor XOR2 (N3617, N3611, N1840);
buf BUF1 (N3618, N3615);
xor XOR2 (N3619, N3614, N992);
nor NOR3 (N3620, N3616, N1242, N3505);
xor XOR2 (N3621, N3620, N1145);
buf BUF1 (N3622, N3582);
nor NOR4 (N3623, N3621, N1099, N3601, N2975);
xor XOR2 (N3624, N3619, N1116);
nand NAND3 (N3625, N3617, N3004, N606);
xor XOR2 (N3626, N3597, N293);
and AND4 (N3627, N3612, N2043, N2623, N327);
xor XOR2 (N3628, N3623, N574);
and AND2 (N3629, N3626, N1521);
xor XOR2 (N3630, N3628, N778);
nor NOR4 (N3631, N3581, N2693, N2302, N1994);
or OR2 (N3632, N3608, N2751);
buf BUF1 (N3633, N3600);
buf BUF1 (N3634, N3622);
and AND2 (N3635, N3624, N2958);
xor XOR2 (N3636, N3629, N401);
nor NOR2 (N3637, N3618, N3215);
nand NAND3 (N3638, N3635, N2755, N2159);
buf BUF1 (N3639, N3638);
xor XOR2 (N3640, N3625, N232);
and AND3 (N3641, N3631, N1084, N542);
or OR4 (N3642, N3627, N3628, N1687, N2600);
xor XOR2 (N3643, N3630, N835);
nor NOR4 (N3644, N3639, N512, N2358, N1613);
buf BUF1 (N3645, N3643);
or OR3 (N3646, N3640, N2767, N1865);
nor NOR4 (N3647, N3632, N2126, N2459, N3306);
not NOT1 (N3648, N3637);
and AND2 (N3649, N3636, N815);
and AND4 (N3650, N3641, N3226, N3487, N3356);
or OR4 (N3651, N3650, N852, N3368, N785);
nor NOR4 (N3652, N3634, N233, N465, N3549);
and AND2 (N3653, N3647, N2471);
xor XOR2 (N3654, N3644, N2724);
or OR2 (N3655, N3648, N3232);
nor NOR2 (N3656, N3645, N1187);
buf BUF1 (N3657, N3652);
not NOT1 (N3658, N3642);
buf BUF1 (N3659, N3649);
buf BUF1 (N3660, N3654);
not NOT1 (N3661, N3659);
nor NOR2 (N3662, N3633, N3508);
nor NOR3 (N3663, N3660, N233, N2757);
buf BUF1 (N3664, N3653);
and AND3 (N3665, N3664, N1911, N3534);
not NOT1 (N3666, N3658);
xor XOR2 (N3667, N3661, N142);
and AND3 (N3668, N3651, N3272, N3658);
xor XOR2 (N3669, N3655, N1048);
not NOT1 (N3670, N3657);
nor NOR4 (N3671, N3668, N2246, N425, N1803);
nand NAND2 (N3672, N3671, N538);
xor XOR2 (N3673, N3665, N3464);
buf BUF1 (N3674, N3662);
xor XOR2 (N3675, N3666, N1501);
or OR4 (N3676, N3669, N1749, N381, N545);
not NOT1 (N3677, N3675);
buf BUF1 (N3678, N3646);
and AND2 (N3679, N3672, N3000);
nor NOR4 (N3680, N3676, N957, N1876, N3346);
nor NOR2 (N3681, N3673, N2536);
nand NAND4 (N3682, N3678, N979, N3188, N288);
not NOT1 (N3683, N3667);
not NOT1 (N3684, N3674);
buf BUF1 (N3685, N3682);
buf BUF1 (N3686, N3683);
or OR4 (N3687, N3681, N2327, N1867, N3101);
and AND4 (N3688, N3680, N2297, N2077, N1325);
and AND2 (N3689, N3685, N1794);
nand NAND3 (N3690, N3686, N1543, N2701);
nor NOR3 (N3691, N3677, N2113, N1123);
buf BUF1 (N3692, N3656);
and AND4 (N3693, N3688, N3107, N3183, N3093);
xor XOR2 (N3694, N3690, N963);
nand NAND2 (N3695, N3693, N3426);
not NOT1 (N3696, N3684);
nor NOR4 (N3697, N3663, N2140, N2453, N357);
nand NAND4 (N3698, N3689, N1689, N424, N1947);
or OR2 (N3699, N3679, N2652);
buf BUF1 (N3700, N3694);
not NOT1 (N3701, N3670);
not NOT1 (N3702, N3687);
xor XOR2 (N3703, N3695, N2916);
nor NOR4 (N3704, N3696, N2859, N1561, N1960);
nand NAND2 (N3705, N3700, N266);
nor NOR2 (N3706, N3704, N2340);
xor XOR2 (N3707, N3703, N3482);
nand NAND2 (N3708, N3706, N3372);
nor NOR4 (N3709, N3697, N2292, N437, N1236);
not NOT1 (N3710, N3701);
nor NOR3 (N3711, N3692, N29, N2761);
and AND3 (N3712, N3705, N2770, N1786);
not NOT1 (N3713, N3710);
nand NAND4 (N3714, N3712, N1266, N1355, N3083);
and AND4 (N3715, N3707, N3039, N2499, N2626);
or OR4 (N3716, N3709, N1021, N1565, N3001);
not NOT1 (N3717, N3698);
nand NAND2 (N3718, N3708, N2478);
nor NOR4 (N3719, N3699, N1333, N1571, N2331);
buf BUF1 (N3720, N3716);
or OR3 (N3721, N3720, N3610, N1351);
nor NOR3 (N3722, N3711, N2565, N1140);
nor NOR2 (N3723, N3719, N64);
buf BUF1 (N3724, N3723);
not NOT1 (N3725, N3718);
nand NAND3 (N3726, N3691, N3109, N3166);
and AND2 (N3727, N3702, N3289);
nand NAND4 (N3728, N3722, N2336, N1548, N1351);
nand NAND3 (N3729, N3727, N1421, N1170);
or OR2 (N3730, N3715, N2855);
xor XOR2 (N3731, N3717, N1990);
nand NAND2 (N3732, N3721, N2276);
nor NOR3 (N3733, N3725, N951, N1955);
or OR2 (N3734, N3733, N3002);
buf BUF1 (N3735, N3726);
buf BUF1 (N3736, N3732);
and AND3 (N3737, N3729, N669, N1863);
buf BUF1 (N3738, N3730);
buf BUF1 (N3739, N3738);
not NOT1 (N3740, N3713);
and AND4 (N3741, N3728, N20, N751, N2143);
xor XOR2 (N3742, N3734, N2953);
nand NAND4 (N3743, N3742, N536, N1587, N2524);
buf BUF1 (N3744, N3731);
xor XOR2 (N3745, N3714, N1998);
and AND2 (N3746, N3741, N774);
buf BUF1 (N3747, N3746);
or OR2 (N3748, N3743, N2983);
not NOT1 (N3749, N3737);
and AND4 (N3750, N3748, N3421, N1480, N143);
nand NAND2 (N3751, N3739, N1021);
or OR2 (N3752, N3735, N2018);
xor XOR2 (N3753, N3744, N3572);
not NOT1 (N3754, N3749);
xor XOR2 (N3755, N3724, N1777);
nand NAND4 (N3756, N3754, N1562, N1455, N2482);
or OR2 (N3757, N3750, N736);
or OR4 (N3758, N3752, N434, N567, N2707);
or OR3 (N3759, N3740, N769, N3042);
not NOT1 (N3760, N3757);
not NOT1 (N3761, N3753);
nand NAND3 (N3762, N3736, N832, N973);
buf BUF1 (N3763, N3760);
not NOT1 (N3764, N3756);
not NOT1 (N3765, N3764);
nor NOR4 (N3766, N3751, N1839, N2088, N510);
not NOT1 (N3767, N3766);
buf BUF1 (N3768, N3758);
nand NAND3 (N3769, N3745, N2684, N2679);
buf BUF1 (N3770, N3762);
or OR2 (N3771, N3763, N1115);
nor NOR4 (N3772, N3767, N2329, N112, N266);
xor XOR2 (N3773, N3761, N1795);
not NOT1 (N3774, N3769);
nor NOR2 (N3775, N3765, N415);
buf BUF1 (N3776, N3772);
or OR3 (N3777, N3775, N3307, N3150);
nand NAND4 (N3778, N3774, N2523, N256, N991);
xor XOR2 (N3779, N3773, N1528);
nor NOR4 (N3780, N3755, N2930, N2808, N1954);
or OR2 (N3781, N3768, N104);
nand NAND3 (N3782, N3770, N1752, N98);
nand NAND4 (N3783, N3776, N3052, N546, N1633);
nand NAND4 (N3784, N3777, N1059, N1363, N1030);
and AND4 (N3785, N3780, N2281, N3490, N3399);
xor XOR2 (N3786, N3779, N3315);
xor XOR2 (N3787, N3786, N56);
nor NOR4 (N3788, N3785, N2283, N2070, N462);
nand NAND2 (N3789, N3771, N3581);
nand NAND4 (N3790, N3759, N1244, N1817, N2887);
nor NOR3 (N3791, N3787, N588, N1863);
xor XOR2 (N3792, N3789, N963);
nand NAND2 (N3793, N3791, N596);
not NOT1 (N3794, N3783);
nor NOR2 (N3795, N3781, N1459);
not NOT1 (N3796, N3793);
nor NOR4 (N3797, N3747, N165, N2655, N271);
nand NAND3 (N3798, N3788, N1826, N3479);
nor NOR2 (N3799, N3795, N119);
buf BUF1 (N3800, N3796);
or OR4 (N3801, N3790, N1600, N2735, N3155);
nor NOR3 (N3802, N3784, N719, N1499);
buf BUF1 (N3803, N3800);
not NOT1 (N3804, N3792);
nor NOR2 (N3805, N3782, N168);
not NOT1 (N3806, N3799);
not NOT1 (N3807, N3803);
nor NOR3 (N3808, N3807, N3326, N2582);
or OR4 (N3809, N3794, N2429, N1941, N97);
nand NAND2 (N3810, N3797, N2680);
not NOT1 (N3811, N3809);
xor XOR2 (N3812, N3798, N3754);
nor NOR2 (N3813, N3801, N2269);
buf BUF1 (N3814, N3804);
xor XOR2 (N3815, N3811, N3669);
buf BUF1 (N3816, N3812);
nand NAND2 (N3817, N3806, N1257);
or OR3 (N3818, N3808, N2186, N448);
and AND2 (N3819, N3805, N3787);
nand NAND2 (N3820, N3815, N2081);
nor NOR2 (N3821, N3810, N117);
nand NAND2 (N3822, N3816, N3424);
buf BUF1 (N3823, N3814);
nand NAND4 (N3824, N3822, N916, N64, N1618);
xor XOR2 (N3825, N3821, N1151);
nand NAND3 (N3826, N3813, N3177, N541);
nor NOR2 (N3827, N3820, N213);
and AND3 (N3828, N3823, N44, N3450);
not NOT1 (N3829, N3824);
nor NOR4 (N3830, N3802, N71, N2477, N3087);
nand NAND3 (N3831, N3778, N2700, N1222);
not NOT1 (N3832, N3830);
and AND3 (N3833, N3817, N2725, N3008);
or OR4 (N3834, N3832, N2706, N1736, N3622);
buf BUF1 (N3835, N3825);
nand NAND4 (N3836, N3834, N530, N3095, N2785);
buf BUF1 (N3837, N3826);
buf BUF1 (N3838, N3827);
not NOT1 (N3839, N3837);
nor NOR2 (N3840, N3838, N1553);
or OR4 (N3841, N3840, N229, N575, N555);
and AND2 (N3842, N3829, N2262);
nand NAND3 (N3843, N3831, N26, N3264);
xor XOR2 (N3844, N3842, N2681);
and AND4 (N3845, N3819, N2528, N3414, N1985);
nor NOR3 (N3846, N3818, N2079, N1810);
not NOT1 (N3847, N3843);
buf BUF1 (N3848, N3835);
nor NOR2 (N3849, N3844, N2561);
buf BUF1 (N3850, N3845);
nand NAND2 (N3851, N3828, N3106);
and AND2 (N3852, N3836, N2080);
nor NOR2 (N3853, N3839, N834);
xor XOR2 (N3854, N3851, N3051);
and AND4 (N3855, N3833, N3707, N3519, N1066);
buf BUF1 (N3856, N3854);
buf BUF1 (N3857, N3841);
buf BUF1 (N3858, N3846);
or OR4 (N3859, N3847, N244, N2676, N706);
or OR4 (N3860, N3849, N1521, N2009, N2537);
not NOT1 (N3861, N3850);
buf BUF1 (N3862, N3852);
and AND4 (N3863, N3859, N3604, N3702, N345);
nand NAND4 (N3864, N3862, N1736, N324, N3256);
not NOT1 (N3865, N3861);
nor NOR3 (N3866, N3865, N3029, N2683);
nand NAND3 (N3867, N3856, N20, N1592);
and AND4 (N3868, N3864, N1715, N219, N2442);
xor XOR2 (N3869, N3848, N2324);
xor XOR2 (N3870, N3855, N1506);
not NOT1 (N3871, N3860);
xor XOR2 (N3872, N3853, N1903);
nand NAND3 (N3873, N3857, N2978, N3855);
buf BUF1 (N3874, N3873);
nor NOR4 (N3875, N3869, N1325, N1360, N1420);
or OR2 (N3876, N3875, N3356);
buf BUF1 (N3877, N3876);
or OR2 (N3878, N3866, N3021);
not NOT1 (N3879, N3872);
and AND2 (N3880, N3870, N3717);
nor NOR3 (N3881, N3858, N3016, N975);
nor NOR3 (N3882, N3880, N2756, N3210);
or OR2 (N3883, N3868, N3154);
or OR4 (N3884, N3883, N3413, N2346, N3655);
buf BUF1 (N3885, N3863);
buf BUF1 (N3886, N3885);
buf BUF1 (N3887, N3871);
xor XOR2 (N3888, N3887, N2830);
and AND4 (N3889, N3867, N2638, N1269, N3139);
or OR4 (N3890, N3874, N2730, N678, N610);
not NOT1 (N3891, N3878);
xor XOR2 (N3892, N3881, N3607);
nor NOR3 (N3893, N3891, N9, N2020);
xor XOR2 (N3894, N3884, N1744);
nand NAND3 (N3895, N3889, N1716, N2813);
and AND3 (N3896, N3888, N3087, N3550);
nand NAND3 (N3897, N3894, N764, N3237);
nor NOR4 (N3898, N3882, N2052, N3010, N1101);
xor XOR2 (N3899, N3896, N376);
not NOT1 (N3900, N3892);
not NOT1 (N3901, N3897);
nand NAND4 (N3902, N3890, N876, N49, N3231);
buf BUF1 (N3903, N3895);
buf BUF1 (N3904, N3877);
nand NAND3 (N3905, N3899, N3224, N3579);
xor XOR2 (N3906, N3903, N2955);
buf BUF1 (N3907, N3898);
and AND2 (N3908, N3886, N584);
not NOT1 (N3909, N3907);
and AND2 (N3910, N3902, N3741);
nand NAND3 (N3911, N3904, N3887, N16);
xor XOR2 (N3912, N3909, N2986);
and AND2 (N3913, N3908, N653);
xor XOR2 (N3914, N3910, N2952);
nand NAND2 (N3915, N3900, N126);
xor XOR2 (N3916, N3905, N973);
or OR2 (N3917, N3893, N1179);
xor XOR2 (N3918, N3913, N1095);
or OR3 (N3919, N3912, N440, N3372);
or OR3 (N3920, N3914, N2984, N2099);
and AND4 (N3921, N3879, N3506, N3840, N3048);
and AND3 (N3922, N3915, N471, N2905);
nor NOR2 (N3923, N3921, N912);
nand NAND4 (N3924, N3918, N837, N3261, N2749);
and AND2 (N3925, N3916, N1034);
or OR4 (N3926, N3924, N136, N1023, N448);
not NOT1 (N3927, N3923);
nand NAND2 (N3928, N3920, N3781);
nand NAND3 (N3929, N3926, N2015, N3702);
not NOT1 (N3930, N3925);
or OR4 (N3931, N3901, N281, N3091, N1232);
xor XOR2 (N3932, N3917, N321);
xor XOR2 (N3933, N3928, N3069);
xor XOR2 (N3934, N3927, N3741);
nor NOR4 (N3935, N3929, N767, N2489, N902);
xor XOR2 (N3936, N3922, N1757);
xor XOR2 (N3937, N3936, N953);
buf BUF1 (N3938, N3911);
nand NAND2 (N3939, N3919, N2204);
buf BUF1 (N3940, N3930);
xor XOR2 (N3941, N3938, N3779);
or OR2 (N3942, N3941, N891);
xor XOR2 (N3943, N3906, N1572);
nand NAND4 (N3944, N3935, N2996, N369, N2135);
not NOT1 (N3945, N3937);
nor NOR4 (N3946, N3944, N2952, N3285, N3695);
nor NOR3 (N3947, N3942, N2410, N1599);
xor XOR2 (N3948, N3933, N2104);
or OR4 (N3949, N3934, N3341, N3683, N3555);
not NOT1 (N3950, N3931);
buf BUF1 (N3951, N3940);
nor NOR4 (N3952, N3945, N42, N22, N2217);
nand NAND2 (N3953, N3948, N1539);
xor XOR2 (N3954, N3953, N3616);
xor XOR2 (N3955, N3947, N1316);
nor NOR4 (N3956, N3955, N2437, N3534, N1360);
nand NAND3 (N3957, N3939, N1548, N3852);
buf BUF1 (N3958, N3932);
xor XOR2 (N3959, N3949, N278);
xor XOR2 (N3960, N3959, N2892);
xor XOR2 (N3961, N3954, N1574);
buf BUF1 (N3962, N3957);
and AND4 (N3963, N3951, N1415, N2004, N3876);
buf BUF1 (N3964, N3962);
buf BUF1 (N3965, N3943);
buf BUF1 (N3966, N3956);
and AND3 (N3967, N3946, N1766, N2050);
xor XOR2 (N3968, N3967, N542);
or OR4 (N3969, N3950, N2247, N1643, N3017);
xor XOR2 (N3970, N3963, N1939);
not NOT1 (N3971, N3969);
buf BUF1 (N3972, N3961);
or OR3 (N3973, N3958, N120, N2404);
or OR2 (N3974, N3970, N8);
and AND3 (N3975, N3968, N1953, N3242);
nand NAND3 (N3976, N3960, N1897, N3066);
and AND3 (N3977, N3964, N3897, N209);
and AND3 (N3978, N3977, N426, N486);
and AND3 (N3979, N3971, N2045, N2514);
buf BUF1 (N3980, N3965);
buf BUF1 (N3981, N3952);
buf BUF1 (N3982, N3966);
nor NOR4 (N3983, N3978, N1074, N2703, N1562);
buf BUF1 (N3984, N3973);
nand NAND4 (N3985, N3984, N3408, N2053, N1688);
nand NAND4 (N3986, N3979, N2172, N992, N3714);
xor XOR2 (N3987, N3986, N536);
or OR4 (N3988, N3983, N3446, N1110, N3166);
nand NAND3 (N3989, N3985, N3499, N1388);
not NOT1 (N3990, N3976);
or OR3 (N3991, N3987, N3959, N997);
and AND4 (N3992, N3991, N1863, N831, N220);
buf BUF1 (N3993, N3990);
buf BUF1 (N3994, N3982);
or OR3 (N3995, N3981, N642, N1451);
nand NAND4 (N3996, N3980, N2451, N2326, N1516);
not NOT1 (N3997, N3994);
xor XOR2 (N3998, N3972, N1834);
xor XOR2 (N3999, N3989, N1056);
nand NAND2 (N4000, N3993, N3131);
and AND3 (N4001, N3974, N1775, N338);
or OR2 (N4002, N4000, N3096);
nand NAND4 (N4003, N3998, N3747, N1310, N2360);
nand NAND2 (N4004, N4001, N2848);
or OR3 (N4005, N3996, N957, N3181);
not NOT1 (N4006, N3999);
buf BUF1 (N4007, N4003);
or OR4 (N4008, N3992, N983, N1604, N3177);
nand NAND4 (N4009, N4002, N3936, N846, N3082);
xor XOR2 (N4010, N3975, N1016);
or OR4 (N4011, N4005, N1285, N92, N2143);
and AND2 (N4012, N4007, N2899);
nor NOR4 (N4013, N4012, N3238, N1924, N1353);
or OR2 (N4014, N4009, N1596);
xor XOR2 (N4015, N4013, N3023);
nor NOR3 (N4016, N3995, N3362, N2126);
xor XOR2 (N4017, N3997, N3782);
xor XOR2 (N4018, N4004, N44);
nor NOR2 (N4019, N3988, N2342);
or OR4 (N4020, N4018, N1238, N52, N2185);
and AND3 (N4021, N4020, N1522, N149);
and AND3 (N4022, N4010, N1808, N3517);
or OR4 (N4023, N4017, N251, N3382, N3973);
xor XOR2 (N4024, N4006, N2538);
buf BUF1 (N4025, N4024);
nand NAND2 (N4026, N4014, N1403);
nand NAND2 (N4027, N4021, N3660);
and AND4 (N4028, N4027, N1301, N460, N2856);
nor NOR3 (N4029, N4015, N1990, N887);
nand NAND4 (N4030, N4023, N275, N3168, N3586);
or OR2 (N4031, N4019, N1905);
buf BUF1 (N4032, N4008);
buf BUF1 (N4033, N4011);
or OR4 (N4034, N4025, N1671, N2757, N1527);
not NOT1 (N4035, N4032);
nor NOR2 (N4036, N4029, N1370);
or OR2 (N4037, N4036, N128);
buf BUF1 (N4038, N4016);
nor NOR3 (N4039, N4030, N1182, N2292);
nand NAND2 (N4040, N4035, N241);
buf BUF1 (N4041, N4040);
and AND2 (N4042, N4041, N3211);
or OR3 (N4043, N4042, N1620, N2491);
buf BUF1 (N4044, N4034);
nor NOR2 (N4045, N4039, N1969);
nand NAND2 (N4046, N4043, N3686);
nor NOR4 (N4047, N4022, N1752, N3342, N60);
nor NOR3 (N4048, N4046, N2747, N3460);
not NOT1 (N4049, N4031);
and AND4 (N4050, N4048, N3149, N3024, N789);
and AND3 (N4051, N4028, N1238, N2481);
xor XOR2 (N4052, N4026, N1491);
and AND2 (N4053, N4051, N362);
nand NAND3 (N4054, N4053, N3784, N3593);
nor NOR2 (N4055, N4044, N993);
nand NAND3 (N4056, N4038, N1269, N1949);
not NOT1 (N4057, N4045);
or OR4 (N4058, N4055, N636, N1176, N3039);
or OR4 (N4059, N4057, N4039, N2835, N1042);
or OR2 (N4060, N4058, N780);
nor NOR4 (N4061, N4049, N1849, N3719, N865);
not NOT1 (N4062, N4054);
and AND3 (N4063, N4060, N2348, N3152);
xor XOR2 (N4064, N4059, N3112);
not NOT1 (N4065, N4052);
not NOT1 (N4066, N4064);
nor NOR3 (N4067, N4065, N3080, N23);
or OR2 (N4068, N4066, N1155);
buf BUF1 (N4069, N4033);
nand NAND3 (N4070, N4063, N2063, N3506);
buf BUF1 (N4071, N4061);
nand NAND2 (N4072, N4037, N1226);
nor NOR3 (N4073, N4068, N1019, N3218);
and AND2 (N4074, N4072, N2476);
or OR4 (N4075, N4069, N3121, N2967, N1614);
and AND3 (N4076, N4062, N1347, N270);
and AND4 (N4077, N4050, N2445, N3298, N125);
buf BUF1 (N4078, N4071);
xor XOR2 (N4079, N4056, N2253);
or OR4 (N4080, N4067, N567, N3550, N4062);
or OR3 (N4081, N4079, N387, N704);
nand NAND4 (N4082, N4078, N4040, N2058, N2848);
not NOT1 (N4083, N4073);
xor XOR2 (N4084, N4082, N229);
or OR4 (N4085, N4081, N1714, N2191, N4082);
nor NOR4 (N4086, N4047, N2973, N3295, N1581);
and AND3 (N4087, N4080, N4037, N2011);
not NOT1 (N4088, N4077);
xor XOR2 (N4089, N4074, N2009);
not NOT1 (N4090, N4089);
buf BUF1 (N4091, N4086);
and AND2 (N4092, N4083, N2030);
and AND3 (N4093, N4084, N3845, N1550);
or OR4 (N4094, N4088, N2697, N574, N4006);
xor XOR2 (N4095, N4087, N3445);
nand NAND2 (N4096, N4075, N2832);
or OR4 (N4097, N4095, N965, N305, N1289);
buf BUF1 (N4098, N4090);
nand NAND3 (N4099, N4094, N2299, N2007);
not NOT1 (N4100, N4097);
xor XOR2 (N4101, N4091, N2980);
and AND2 (N4102, N4096, N2716);
and AND2 (N4103, N4085, N1617);
or OR3 (N4104, N4102, N1317, N1997);
buf BUF1 (N4105, N4092);
buf BUF1 (N4106, N4098);
or OR2 (N4107, N4093, N3669);
or OR2 (N4108, N4103, N2259);
and AND2 (N4109, N4105, N2895);
nand NAND3 (N4110, N4076, N2353, N3530);
buf BUF1 (N4111, N4104);
nor NOR3 (N4112, N4109, N2067, N2496);
xor XOR2 (N4113, N4110, N2762);
xor XOR2 (N4114, N4108, N866);
nor NOR2 (N4115, N4099, N3940);
not NOT1 (N4116, N4106);
xor XOR2 (N4117, N4115, N4011);
buf BUF1 (N4118, N4114);
not NOT1 (N4119, N4107);
or OR3 (N4120, N4111, N786, N2173);
xor XOR2 (N4121, N4120, N3648);
buf BUF1 (N4122, N4117);
nand NAND3 (N4123, N4100, N1652, N1753);
buf BUF1 (N4124, N4070);
or OR3 (N4125, N4123, N1120, N2573);
or OR4 (N4126, N4116, N2317, N2992, N3391);
xor XOR2 (N4127, N4126, N2847);
xor XOR2 (N4128, N4122, N2708);
and AND4 (N4129, N4121, N1893, N2339, N134);
buf BUF1 (N4130, N4118);
or OR4 (N4131, N4101, N589, N572, N10);
and AND4 (N4132, N4131, N2855, N466, N3012);
xor XOR2 (N4133, N4112, N1939);
and AND4 (N4134, N4119, N3004, N1359, N891);
xor XOR2 (N4135, N4127, N2155);
nor NOR3 (N4136, N4130, N2300, N1188);
not NOT1 (N4137, N4133);
nand NAND2 (N4138, N4113, N896);
xor XOR2 (N4139, N4125, N1352);
not NOT1 (N4140, N4136);
nand NAND4 (N4141, N4137, N2613, N1309, N3469);
xor XOR2 (N4142, N4138, N865);
nor NOR4 (N4143, N4129, N1068, N1379, N610);
and AND4 (N4144, N4140, N2503, N2773, N194);
nand NAND4 (N4145, N4124, N299, N1930, N578);
nand NAND2 (N4146, N4139, N2873);
nand NAND4 (N4147, N4143, N2660, N125, N493);
xor XOR2 (N4148, N4134, N3043);
nand NAND3 (N4149, N4148, N3759, N345);
and AND4 (N4150, N4128, N1630, N255, N4024);
buf BUF1 (N4151, N4135);
xor XOR2 (N4152, N4146, N1121);
nand NAND3 (N4153, N4145, N1910, N2751);
and AND4 (N4154, N4153, N3632, N1814, N565);
not NOT1 (N4155, N4150);
nand NAND2 (N4156, N4151, N669);
or OR4 (N4157, N4141, N215, N3406, N1905);
xor XOR2 (N4158, N4149, N3095);
not NOT1 (N4159, N4157);
buf BUF1 (N4160, N4147);
nor NOR4 (N4161, N4160, N2730, N2557, N3525);
or OR2 (N4162, N4132, N138);
buf BUF1 (N4163, N4162);
xor XOR2 (N4164, N4155, N2289);
or OR3 (N4165, N4156, N1541, N451);
nand NAND2 (N4166, N4165, N1497);
nand NAND2 (N4167, N4154, N3547);
and AND2 (N4168, N4144, N1741);
xor XOR2 (N4169, N4158, N55);
or OR2 (N4170, N4164, N194);
and AND3 (N4171, N4159, N2261, N2480);
and AND3 (N4172, N4170, N3120, N2238);
and AND3 (N4173, N4166, N845, N2129);
or OR3 (N4174, N4168, N2556, N1913);
nand NAND3 (N4175, N4172, N4161, N3187);
and AND4 (N4176, N1206, N1402, N3457, N2687);
nand NAND3 (N4177, N4176, N533, N3195);
and AND2 (N4178, N4163, N679);
nand NAND4 (N4179, N4152, N2531, N1569, N3769);
buf BUF1 (N4180, N4177);
nand NAND2 (N4181, N4169, N2804);
nand NAND4 (N4182, N4171, N507, N3661, N1136);
and AND2 (N4183, N4180, N2846);
and AND3 (N4184, N4183, N4121, N882);
and AND2 (N4185, N4175, N3402);
or OR4 (N4186, N4167, N2511, N1599, N2631);
and AND2 (N4187, N4178, N2898);
xor XOR2 (N4188, N4173, N1050);
nand NAND2 (N4189, N4184, N3834);
buf BUF1 (N4190, N4185);
or OR4 (N4191, N4179, N3607, N2521, N3684);
not NOT1 (N4192, N4191);
buf BUF1 (N4193, N4188);
and AND2 (N4194, N4190, N389);
nand NAND2 (N4195, N4193, N1042);
xor XOR2 (N4196, N4186, N18);
and AND4 (N4197, N4189, N3023, N1243, N1432);
nand NAND3 (N4198, N4182, N1553, N3754);
nand NAND4 (N4199, N4174, N2258, N3960, N486);
buf BUF1 (N4200, N4181);
or OR2 (N4201, N4142, N3052);
buf BUF1 (N4202, N4196);
or OR2 (N4203, N4187, N3183);
not NOT1 (N4204, N4203);
nand NAND3 (N4205, N4200, N440, N1968);
buf BUF1 (N4206, N4205);
nand NAND2 (N4207, N4201, N282);
not NOT1 (N4208, N4202);
not NOT1 (N4209, N4195);
buf BUF1 (N4210, N4207);
not NOT1 (N4211, N4204);
and AND4 (N4212, N4199, N1643, N1240, N3360);
not NOT1 (N4213, N4194);
or OR3 (N4214, N4211, N2719, N96);
or OR3 (N4215, N4198, N2423, N877);
not NOT1 (N4216, N4209);
nor NOR2 (N4217, N4192, N4030);
nand NAND4 (N4218, N4197, N2749, N1249, N1655);
not NOT1 (N4219, N4218);
xor XOR2 (N4220, N4212, N4180);
and AND4 (N4221, N4208, N3681, N3540, N3394);
and AND3 (N4222, N4206, N754, N3776);
buf BUF1 (N4223, N4217);
or OR3 (N4224, N4210, N629, N1632);
not NOT1 (N4225, N4213);
nor NOR3 (N4226, N4221, N524, N1401);
not NOT1 (N4227, N4225);
xor XOR2 (N4228, N4223, N936);
nor NOR2 (N4229, N4215, N3733);
or OR4 (N4230, N4214, N643, N3846, N1434);
not NOT1 (N4231, N4222);
not NOT1 (N4232, N4216);
and AND2 (N4233, N4232, N3824);
buf BUF1 (N4234, N4226);
or OR4 (N4235, N4227, N2516, N97, N3539);
and AND4 (N4236, N4234, N3447, N2067, N3902);
xor XOR2 (N4237, N4233, N860);
nand NAND4 (N4238, N4224, N1687, N4219, N3619);
nor NOR2 (N4239, N1968, N3771);
xor XOR2 (N4240, N4237, N2481);
nand NAND4 (N4241, N4220, N1472, N2852, N4114);
xor XOR2 (N4242, N4241, N3650);
and AND2 (N4243, N4229, N1258);
nor NOR3 (N4244, N4228, N2190, N3885);
xor XOR2 (N4245, N4243, N3025);
xor XOR2 (N4246, N4245, N3450);
nand NAND2 (N4247, N4244, N4179);
not NOT1 (N4248, N4246);
and AND3 (N4249, N4239, N2310, N950);
or OR4 (N4250, N4236, N1841, N624, N765);
not NOT1 (N4251, N4242);
or OR3 (N4252, N4251, N3344, N1013);
and AND4 (N4253, N4231, N1946, N1151, N3000);
nor NOR3 (N4254, N4235, N521, N4222);
or OR4 (N4255, N4240, N3975, N3986, N3444);
buf BUF1 (N4256, N4252);
xor XOR2 (N4257, N4253, N3519);
not NOT1 (N4258, N4250);
nor NOR4 (N4259, N4249, N2745, N937, N1531);
buf BUF1 (N4260, N4255);
or OR2 (N4261, N4247, N2174);
xor XOR2 (N4262, N4259, N3102);
or OR2 (N4263, N4254, N2178);
xor XOR2 (N4264, N4258, N3950);
buf BUF1 (N4265, N4256);
buf BUF1 (N4266, N4264);
and AND2 (N4267, N4257, N2955);
nand NAND2 (N4268, N4248, N923);
buf BUF1 (N4269, N4268);
nor NOR2 (N4270, N4260, N4058);
buf BUF1 (N4271, N4261);
and AND2 (N4272, N4269, N195);
and AND3 (N4273, N4272, N2595, N23);
and AND4 (N4274, N4267, N3520, N2868, N1139);
not NOT1 (N4275, N4274);
nor NOR2 (N4276, N4270, N2926);
or OR4 (N4277, N4276, N2708, N76, N1284);
nand NAND4 (N4278, N4265, N1061, N544, N4232);
nor NOR4 (N4279, N4273, N603, N2559, N3226);
buf BUF1 (N4280, N4266);
buf BUF1 (N4281, N4262);
nand NAND3 (N4282, N4230, N1335, N747);
buf BUF1 (N4283, N4275);
and AND4 (N4284, N4281, N3358, N3323, N2003);
xor XOR2 (N4285, N4284, N1602);
xor XOR2 (N4286, N4280, N879);
xor XOR2 (N4287, N4277, N3739);
xor XOR2 (N4288, N4278, N4167);
xor XOR2 (N4289, N4286, N2143);
and AND2 (N4290, N4283, N531);
not NOT1 (N4291, N4271);
and AND4 (N4292, N4287, N2315, N974, N3021);
and AND4 (N4293, N4285, N2414, N517, N2319);
not NOT1 (N4294, N4282);
or OR2 (N4295, N4238, N1905);
or OR2 (N4296, N4291, N1838);
nand NAND4 (N4297, N4288, N3895, N1968, N3731);
buf BUF1 (N4298, N4279);
nor NOR3 (N4299, N4293, N1340, N3864);
and AND3 (N4300, N4289, N703, N3392);
xor XOR2 (N4301, N4290, N4032);
not NOT1 (N4302, N4299);
buf BUF1 (N4303, N4263);
nor NOR3 (N4304, N4294, N705, N2490);
xor XOR2 (N4305, N4300, N1435);
nand NAND4 (N4306, N4302, N2008, N2224, N1548);
or OR4 (N4307, N4301, N3398, N505, N3104);
buf BUF1 (N4308, N4298);
xor XOR2 (N4309, N4303, N368);
nand NAND4 (N4310, N4307, N720, N1610, N647);
nor NOR2 (N4311, N4296, N1123);
xor XOR2 (N4312, N4305, N1008);
nand NAND4 (N4313, N4312, N1814, N868, N3196);
not NOT1 (N4314, N4310);
nand NAND2 (N4315, N4306, N2216);
xor XOR2 (N4316, N4313, N2468);
nand NAND2 (N4317, N4297, N2447);
buf BUF1 (N4318, N4314);
buf BUF1 (N4319, N4304);
nand NAND3 (N4320, N4308, N1281, N1718);
or OR2 (N4321, N4320, N790);
nand NAND2 (N4322, N4295, N240);
nor NOR4 (N4323, N4318, N4120, N3589, N3075);
xor XOR2 (N4324, N4315, N1758);
not NOT1 (N4325, N4321);
or OR4 (N4326, N4316, N306, N107, N1698);
or OR3 (N4327, N4326, N1463, N2613);
not NOT1 (N4328, N4309);
or OR4 (N4329, N4328, N884, N1987, N2670);
nor NOR4 (N4330, N4324, N1360, N3530, N2004);
nor NOR3 (N4331, N4292, N3882, N4325);
or OR2 (N4332, N3434, N2298);
nand NAND2 (N4333, N4311, N3142);
or OR2 (N4334, N4333, N104);
and AND4 (N4335, N4334, N3689, N3155, N1599);
buf BUF1 (N4336, N4335);
nand NAND3 (N4337, N4331, N1444, N1758);
nor NOR3 (N4338, N4336, N176, N404);
or OR3 (N4339, N4330, N4006, N3424);
or OR3 (N4340, N4339, N630, N2704);
or OR4 (N4341, N4340, N2754, N378, N3838);
buf BUF1 (N4342, N4319);
or OR3 (N4343, N4338, N2286, N3309);
or OR2 (N4344, N4332, N1668);
nand NAND2 (N4345, N4317, N866);
and AND2 (N4346, N4343, N508);
or OR2 (N4347, N4341, N52);
xor XOR2 (N4348, N4323, N2654);
xor XOR2 (N4349, N4329, N449);
nor NOR2 (N4350, N4345, N2407);
buf BUF1 (N4351, N4344);
buf BUF1 (N4352, N4342);
not NOT1 (N4353, N4349);
not NOT1 (N4354, N4346);
or OR4 (N4355, N4347, N1772, N27, N3393);
nand NAND4 (N4356, N4322, N908, N1027, N480);
and AND2 (N4357, N4352, N813);
not NOT1 (N4358, N4327);
nand NAND2 (N4359, N4351, N2715);
or OR4 (N4360, N4350, N1700, N2307, N3933);
and AND2 (N4361, N4356, N3069);
xor XOR2 (N4362, N4337, N4336);
xor XOR2 (N4363, N4358, N4290);
and AND2 (N4364, N4353, N134);
nand NAND4 (N4365, N4348, N2970, N2053, N196);
or OR4 (N4366, N4361, N406, N1079, N4266);
and AND2 (N4367, N4359, N2049);
xor XOR2 (N4368, N4367, N155);
buf BUF1 (N4369, N4366);
not NOT1 (N4370, N4364);
buf BUF1 (N4371, N4355);
and AND4 (N4372, N4371, N1073, N1782, N3963);
nand NAND2 (N4373, N4368, N1583);
xor XOR2 (N4374, N4365, N3268);
and AND4 (N4375, N4363, N1474, N2901, N4349);
xor XOR2 (N4376, N4360, N2867);
and AND2 (N4377, N4375, N4146);
buf BUF1 (N4378, N4362);
or OR2 (N4379, N4373, N2895);
nand NAND4 (N4380, N4374, N1961, N936, N1851);
not NOT1 (N4381, N4372);
or OR3 (N4382, N4379, N2973, N262);
nand NAND3 (N4383, N4380, N2608, N1139);
or OR3 (N4384, N4357, N1951, N3816);
nand NAND4 (N4385, N4381, N3745, N962, N1802);
and AND4 (N4386, N4370, N871, N2668, N75);
xor XOR2 (N4387, N4384, N2582);
or OR2 (N4388, N4377, N4255);
buf BUF1 (N4389, N4376);
and AND3 (N4390, N4387, N443, N3215);
buf BUF1 (N4391, N4389);
and AND2 (N4392, N4388, N3816);
xor XOR2 (N4393, N4382, N2984);
buf BUF1 (N4394, N4385);
buf BUF1 (N4395, N4390);
not NOT1 (N4396, N4354);
and AND4 (N4397, N4396, N3033, N3565, N3333);
or OR2 (N4398, N4369, N2560);
nor NOR2 (N4399, N4391, N2450);
xor XOR2 (N4400, N4386, N609);
nor NOR2 (N4401, N4399, N665);
or OR3 (N4402, N4378, N691, N8);
or OR2 (N4403, N4393, N1071);
and AND4 (N4404, N4394, N2176, N1519, N858);
and AND2 (N4405, N4402, N4233);
not NOT1 (N4406, N4401);
not NOT1 (N4407, N4397);
or OR3 (N4408, N4403, N4077, N3422);
and AND2 (N4409, N4404, N874);
xor XOR2 (N4410, N4407, N2552);
xor XOR2 (N4411, N4405, N3084);
nor NOR2 (N4412, N4400, N2179);
xor XOR2 (N4413, N4398, N2450);
buf BUF1 (N4414, N4406);
nor NOR4 (N4415, N4414, N66, N3325, N3586);
nand NAND3 (N4416, N4383, N2124, N3504);
nand NAND3 (N4417, N4409, N1355, N3332);
nand NAND3 (N4418, N4417, N2603, N2317);
not NOT1 (N4419, N4392);
nand NAND2 (N4420, N4415, N924);
xor XOR2 (N4421, N4408, N2123);
xor XOR2 (N4422, N4420, N2367);
buf BUF1 (N4423, N4413);
xor XOR2 (N4424, N4410, N1466);
and AND4 (N4425, N4416, N3682, N2003, N3692);
and AND3 (N4426, N4425, N507, N3330);
nand NAND2 (N4427, N4421, N570);
xor XOR2 (N4428, N4412, N4052);
buf BUF1 (N4429, N4418);
or OR4 (N4430, N4423, N2649, N1698, N4286);
xor XOR2 (N4431, N4411, N2049);
or OR2 (N4432, N4428, N2574);
buf BUF1 (N4433, N4427);
buf BUF1 (N4434, N4429);
and AND3 (N4435, N4431, N528, N2298);
buf BUF1 (N4436, N4430);
nand NAND3 (N4437, N4426, N1526, N1299);
and AND2 (N4438, N4395, N2358);
nand NAND3 (N4439, N4422, N577, N2186);
nor NOR3 (N4440, N4437, N442, N1742);
buf BUF1 (N4441, N4439);
or OR2 (N4442, N4432, N1381);
and AND4 (N4443, N4419, N458, N657, N1296);
xor XOR2 (N4444, N4424, N921);
or OR2 (N4445, N4436, N4026);
xor XOR2 (N4446, N4442, N844);
or OR4 (N4447, N4443, N3849, N2515, N2070);
xor XOR2 (N4448, N4441, N3904);
or OR2 (N4449, N4438, N3665);
nand NAND3 (N4450, N4440, N1845, N1060);
buf BUF1 (N4451, N4446);
nor NOR4 (N4452, N4434, N642, N1530, N3735);
or OR3 (N4453, N4447, N3006, N2316);
not NOT1 (N4454, N4448);
nor NOR2 (N4455, N4451, N2216);
xor XOR2 (N4456, N4445, N3341);
buf BUF1 (N4457, N4444);
not NOT1 (N4458, N4455);
buf BUF1 (N4459, N4433);
nor NOR2 (N4460, N4450, N3659);
nor NOR2 (N4461, N4454, N353);
xor XOR2 (N4462, N4456, N549);
buf BUF1 (N4463, N4459);
and AND4 (N4464, N4460, N2087, N3589, N2682);
or OR3 (N4465, N4461, N1812, N2083);
and AND4 (N4466, N4457, N3819, N3191, N1650);
and AND4 (N4467, N4453, N2476, N1749, N2159);
buf BUF1 (N4468, N4449);
or OR2 (N4469, N4467, N1240);
nor NOR4 (N4470, N4452, N2126, N331, N2836);
xor XOR2 (N4471, N4458, N3287);
and AND2 (N4472, N4470, N3826);
buf BUF1 (N4473, N4465);
or OR3 (N4474, N4469, N4204, N3152);
nor NOR3 (N4475, N4463, N970, N4357);
xor XOR2 (N4476, N4462, N4121);
and AND4 (N4477, N4471, N3973, N3367, N1064);
nor NOR4 (N4478, N4468, N1134, N3250, N495);
and AND2 (N4479, N4435, N1324);
or OR4 (N4480, N4475, N839, N867, N2465);
or OR2 (N4481, N4464, N182);
buf BUF1 (N4482, N4466);
and AND4 (N4483, N4482, N4393, N3897, N1747);
nor NOR2 (N4484, N4476, N4254);
xor XOR2 (N4485, N4479, N1354);
not NOT1 (N4486, N4474);
and AND3 (N4487, N4483, N3820, N1614);
xor XOR2 (N4488, N4472, N1908);
not NOT1 (N4489, N4481);
nand NAND3 (N4490, N4480, N249, N3788);
buf BUF1 (N4491, N4477);
buf BUF1 (N4492, N4491);
buf BUF1 (N4493, N4485);
nand NAND3 (N4494, N4484, N2058, N855);
buf BUF1 (N4495, N4494);
buf BUF1 (N4496, N4493);
buf BUF1 (N4497, N4490);
buf BUF1 (N4498, N4495);
xor XOR2 (N4499, N4487, N407);
buf BUF1 (N4500, N4499);
or OR3 (N4501, N4489, N2667, N1114);
or OR2 (N4502, N4501, N530);
buf BUF1 (N4503, N4486);
buf BUF1 (N4504, N4497);
or OR4 (N4505, N4502, N1427, N490, N3805);
and AND2 (N4506, N4503, N4041);
or OR4 (N4507, N4504, N2365, N2951, N248);
xor XOR2 (N4508, N4488, N1980);
xor XOR2 (N4509, N4507, N2989);
or OR3 (N4510, N4496, N1382, N2309);
nor NOR2 (N4511, N4505, N2611);
buf BUF1 (N4512, N4473);
xor XOR2 (N4513, N4498, N4101);
nand NAND3 (N4514, N4478, N538, N3064);
nand NAND2 (N4515, N4500, N3489);
buf BUF1 (N4516, N4492);
nand NAND3 (N4517, N4506, N418, N1656);
buf BUF1 (N4518, N4509);
or OR3 (N4519, N4511, N1861, N2064);
or OR4 (N4520, N4508, N3330, N121, N1801);
nor NOR4 (N4521, N4512, N1967, N3404, N3403);
nand NAND2 (N4522, N4513, N3958);
and AND2 (N4523, N4510, N4516);
buf BUF1 (N4524, N2881);
nand NAND4 (N4525, N4523, N3096, N836, N2155);
and AND4 (N4526, N4520, N2309, N3587, N430);
nand NAND2 (N4527, N4514, N1458);
xor XOR2 (N4528, N4519, N2476);
xor XOR2 (N4529, N4528, N2649);
and AND3 (N4530, N4518, N2102, N763);
or OR3 (N4531, N4527, N1629, N2552);
buf BUF1 (N4532, N4517);
not NOT1 (N4533, N4524);
xor XOR2 (N4534, N4529, N1516);
and AND2 (N4535, N4532, N2833);
xor XOR2 (N4536, N4534, N1553);
buf BUF1 (N4537, N4522);
not NOT1 (N4538, N4533);
not NOT1 (N4539, N4535);
nor NOR2 (N4540, N4537, N4405);
buf BUF1 (N4541, N4540);
xor XOR2 (N4542, N4525, N409);
buf BUF1 (N4543, N4526);
or OR4 (N4544, N4536, N2768, N1507, N2375);
or OR4 (N4545, N4543, N3259, N661, N764);
nand NAND2 (N4546, N4521, N3274);
xor XOR2 (N4547, N4545, N217);
buf BUF1 (N4548, N4538);
buf BUF1 (N4549, N4515);
and AND3 (N4550, N4531, N1636, N3650);
and AND2 (N4551, N4542, N1418);
and AND2 (N4552, N4547, N4502);
nand NAND2 (N4553, N4541, N4282);
nor NOR2 (N4554, N4539, N3122);
and AND3 (N4555, N4549, N3209, N2484);
or OR2 (N4556, N4544, N1357);
xor XOR2 (N4557, N4551, N3306);
nor NOR2 (N4558, N4550, N1991);
nor NOR2 (N4559, N4530, N3088);
not NOT1 (N4560, N4553);
or OR2 (N4561, N4555, N1470);
nand NAND4 (N4562, N4552, N2967, N3876, N2404);
nor NOR3 (N4563, N4556, N120, N3287);
or OR3 (N4564, N4554, N2829, N629);
nor NOR3 (N4565, N4548, N852, N128);
or OR4 (N4566, N4562, N615, N2333, N2905);
nor NOR4 (N4567, N4557, N3099, N1134, N2914);
buf BUF1 (N4568, N4559);
and AND4 (N4569, N4565, N400, N1582, N3138);
or OR2 (N4570, N4568, N951);
or OR4 (N4571, N4546, N2795, N1289, N426);
and AND4 (N4572, N4560, N4134, N2073, N2232);
xor XOR2 (N4573, N4561, N742);
and AND4 (N4574, N4567, N3605, N1516, N327);
not NOT1 (N4575, N4564);
xor XOR2 (N4576, N4574, N1816);
nor NOR2 (N4577, N4576, N3622);
and AND4 (N4578, N4570, N2470, N4096, N3510);
and AND3 (N4579, N4569, N3990, N386);
buf BUF1 (N4580, N4572);
xor XOR2 (N4581, N4573, N4316);
xor XOR2 (N4582, N4580, N2137);
not NOT1 (N4583, N4579);
nand NAND2 (N4584, N4558, N3158);
nand NAND4 (N4585, N4577, N3610, N703, N489);
nor NOR4 (N4586, N4575, N454, N3517, N2749);
nand NAND2 (N4587, N4563, N3524);
not NOT1 (N4588, N4586);
nand NAND4 (N4589, N4587, N1801, N2688, N252);
or OR2 (N4590, N4571, N3274);
or OR4 (N4591, N4584, N2036, N3280, N1214);
and AND3 (N4592, N4585, N4310, N465);
and AND2 (N4593, N4590, N1161);
not NOT1 (N4594, N4581);
buf BUF1 (N4595, N4582);
nand NAND2 (N4596, N4566, N3012);
xor XOR2 (N4597, N4593, N2298);
nand NAND2 (N4598, N4591, N932);
buf BUF1 (N4599, N4595);
not NOT1 (N4600, N4578);
xor XOR2 (N4601, N4589, N1067);
not NOT1 (N4602, N4601);
and AND2 (N4603, N4596, N2986);
or OR2 (N4604, N4588, N2338);
and AND2 (N4605, N4597, N4195);
buf BUF1 (N4606, N4592);
nor NOR4 (N4607, N4600, N659, N3256, N3537);
buf BUF1 (N4608, N4604);
nor NOR3 (N4609, N4602, N4266, N2927);
not NOT1 (N4610, N4605);
nor NOR2 (N4611, N4608, N2812);
nand NAND4 (N4612, N4603, N4206, N2919, N2794);
and AND4 (N4613, N4609, N394, N4218, N3505);
and AND2 (N4614, N4607, N636);
nand NAND4 (N4615, N4594, N1992, N2189, N424);
buf BUF1 (N4616, N4615);
xor XOR2 (N4617, N4616, N3648);
or OR2 (N4618, N4610, N4241);
and AND3 (N4619, N4618, N837, N566);
xor XOR2 (N4620, N4617, N2803);
or OR2 (N4621, N4598, N1599);
or OR3 (N4622, N4606, N3351, N4394);
not NOT1 (N4623, N4599);
nor NOR4 (N4624, N4613, N3666, N1026, N273);
or OR2 (N4625, N4622, N4399);
nand NAND2 (N4626, N4612, N2913);
nor NOR4 (N4627, N4625, N2072, N543, N4105);
not NOT1 (N4628, N4627);
buf BUF1 (N4629, N4614);
xor XOR2 (N4630, N4629, N1706);
or OR3 (N4631, N4624, N3763, N4047);
buf BUF1 (N4632, N4583);
or OR4 (N4633, N4630, N865, N2405, N3993);
not NOT1 (N4634, N4626);
and AND2 (N4635, N4633, N3748);
buf BUF1 (N4636, N4634);
not NOT1 (N4637, N4611);
not NOT1 (N4638, N4635);
or OR4 (N4639, N4623, N1702, N2534, N38);
nor NOR2 (N4640, N4637, N3379);
not NOT1 (N4641, N4638);
nand NAND4 (N4642, N4628, N2993, N688, N4092);
buf BUF1 (N4643, N4641);
buf BUF1 (N4644, N4620);
buf BUF1 (N4645, N4642);
or OR4 (N4646, N4621, N426, N3993, N169);
not NOT1 (N4647, N4645);
nor NOR2 (N4648, N4644, N3852);
xor XOR2 (N4649, N4643, N516);
not NOT1 (N4650, N4619);
or OR3 (N4651, N4650, N2920, N699);
buf BUF1 (N4652, N4647);
xor XOR2 (N4653, N4646, N2764);
and AND3 (N4654, N4648, N524, N1424);
and AND4 (N4655, N4639, N2160, N3890, N3909);
and AND4 (N4656, N4649, N666, N355, N761);
buf BUF1 (N4657, N4651);
and AND3 (N4658, N4654, N1581, N830);
nor NOR4 (N4659, N4657, N1294, N436, N865);
nor NOR3 (N4660, N4631, N867, N4424);
and AND3 (N4661, N4652, N4541, N4305);
not NOT1 (N4662, N4636);
nor NOR2 (N4663, N4658, N2287);
buf BUF1 (N4664, N4659);
or OR4 (N4665, N4656, N4390, N241, N2686);
xor XOR2 (N4666, N4661, N4030);
buf BUF1 (N4667, N4662);
nand NAND3 (N4668, N4666, N2377, N1639);
not NOT1 (N4669, N4655);
or OR4 (N4670, N4664, N2187, N1593, N3351);
nand NAND4 (N4671, N4663, N1611, N4195, N3136);
not NOT1 (N4672, N4670);
buf BUF1 (N4673, N4672);
or OR3 (N4674, N4660, N453, N2114);
not NOT1 (N4675, N4632);
buf BUF1 (N4676, N4653);
buf BUF1 (N4677, N4674);
not NOT1 (N4678, N4667);
xor XOR2 (N4679, N4676, N714);
buf BUF1 (N4680, N4673);
xor XOR2 (N4681, N4669, N2027);
and AND2 (N4682, N4668, N1042);
buf BUF1 (N4683, N4665);
and AND4 (N4684, N4679, N3611, N3593, N660);
and AND2 (N4685, N4684, N908);
not NOT1 (N4686, N4683);
buf BUF1 (N4687, N4682);
not NOT1 (N4688, N4681);
nand NAND4 (N4689, N4640, N1364, N1830, N2408);
nor NOR4 (N4690, N4671, N1649, N767, N1041);
and AND2 (N4691, N4690, N3236);
buf BUF1 (N4692, N4675);
xor XOR2 (N4693, N4688, N1640);
not NOT1 (N4694, N4685);
or OR4 (N4695, N4693, N2428, N1389, N3149);
or OR3 (N4696, N4694, N3222, N4122);
buf BUF1 (N4697, N4692);
or OR4 (N4698, N4697, N1581, N2895, N696);
and AND2 (N4699, N4689, N897);
nand NAND3 (N4700, N4696, N2724, N1767);
and AND3 (N4701, N4680, N4636, N3868);
nor NOR4 (N4702, N4700, N300, N2561, N415);
nand NAND4 (N4703, N4691, N197, N547, N2278);
or OR2 (N4704, N4677, N1027);
xor XOR2 (N4705, N4678, N2540);
nor NOR3 (N4706, N4695, N2261, N3482);
not NOT1 (N4707, N4702);
or OR2 (N4708, N4704, N1828);
or OR4 (N4709, N4708, N691, N4609, N424);
xor XOR2 (N4710, N4699, N584);
nor NOR4 (N4711, N4686, N2993, N3034, N17);
xor XOR2 (N4712, N4687, N280);
xor XOR2 (N4713, N4710, N3201);
nand NAND3 (N4714, N4701, N1924, N4641);
buf BUF1 (N4715, N4706);
and AND2 (N4716, N4709, N421);
and AND2 (N4717, N4711, N3913);
buf BUF1 (N4718, N4703);
not NOT1 (N4719, N4713);
buf BUF1 (N4720, N4715);
not NOT1 (N4721, N4720);
xor XOR2 (N4722, N4717, N3619);
and AND4 (N4723, N4721, N1744, N2264, N2490);
buf BUF1 (N4724, N4712);
not NOT1 (N4725, N4707);
and AND2 (N4726, N4722, N1537);
buf BUF1 (N4727, N4705);
or OR2 (N4728, N4714, N2338);
buf BUF1 (N4729, N4725);
buf BUF1 (N4730, N4718);
nor NOR3 (N4731, N4730, N481, N901);
or OR3 (N4732, N4698, N1734, N3216);
not NOT1 (N4733, N4716);
and AND3 (N4734, N4719, N646, N1541);
or OR3 (N4735, N4729, N1436, N3133);
not NOT1 (N4736, N4731);
nor NOR4 (N4737, N4727, N2983, N3740, N2730);
nor NOR4 (N4738, N4736, N1553, N4566, N2857);
nor NOR3 (N4739, N4732, N158, N3716);
not NOT1 (N4740, N4739);
or OR4 (N4741, N4728, N1921, N4436, N821);
nand NAND2 (N4742, N4738, N985);
and AND3 (N4743, N4724, N692, N1060);
nor NOR2 (N4744, N4734, N3135);
nor NOR2 (N4745, N4723, N2456);
nor NOR3 (N4746, N4737, N1722, N2439);
nor NOR4 (N4747, N4743, N2746, N333, N2198);
nor NOR2 (N4748, N4742, N3226);
nor NOR2 (N4749, N4747, N1652);
or OR2 (N4750, N4748, N1480);
nand NAND3 (N4751, N4746, N1912, N3641);
not NOT1 (N4752, N4745);
nor NOR4 (N4753, N4751, N1023, N2930, N4728);
xor XOR2 (N4754, N4740, N2561);
and AND3 (N4755, N4735, N443, N1082);
buf BUF1 (N4756, N4754);
or OR3 (N4757, N4750, N3125, N4046);
xor XOR2 (N4758, N4757, N4342);
nand NAND3 (N4759, N4753, N1244, N438);
xor XOR2 (N4760, N4756, N2078);
and AND2 (N4761, N4749, N1017);
nand NAND2 (N4762, N4726, N1359);
xor XOR2 (N4763, N4761, N1162);
nand NAND2 (N4764, N4762, N3449);
and AND3 (N4765, N4760, N2389, N1681);
not NOT1 (N4766, N4764);
xor XOR2 (N4767, N4759, N3294);
xor XOR2 (N4768, N4752, N4643);
nor NOR2 (N4769, N4755, N3532);
not NOT1 (N4770, N4768);
or OR2 (N4771, N4763, N1382);
and AND4 (N4772, N4766, N1102, N1439, N3080);
nor NOR4 (N4773, N4772, N54, N2340, N4382);
nand NAND2 (N4774, N4765, N1041);
xor XOR2 (N4775, N4769, N1797);
and AND2 (N4776, N4770, N1132);
and AND3 (N4777, N4744, N2192, N3964);
nor NOR2 (N4778, N4767, N1153);
xor XOR2 (N4779, N4776, N1713);
xor XOR2 (N4780, N4773, N1019);
buf BUF1 (N4781, N4771);
nand NAND4 (N4782, N4781, N4698, N180, N2255);
and AND4 (N4783, N4780, N3658, N3004, N1544);
not NOT1 (N4784, N4777);
nand NAND4 (N4785, N4782, N12, N3904, N4051);
xor XOR2 (N4786, N4778, N3131);
xor XOR2 (N4787, N4741, N2324);
buf BUF1 (N4788, N4779);
or OR2 (N4789, N4784, N1941);
not NOT1 (N4790, N4785);
xor XOR2 (N4791, N4790, N3606);
xor XOR2 (N4792, N4758, N2196);
buf BUF1 (N4793, N4774);
buf BUF1 (N4794, N4787);
buf BUF1 (N4795, N4788);
and AND4 (N4796, N4789, N681, N1659, N1142);
buf BUF1 (N4797, N4775);
buf BUF1 (N4798, N4795);
xor XOR2 (N4799, N4783, N2213);
buf BUF1 (N4800, N4799);
buf BUF1 (N4801, N4798);
xor XOR2 (N4802, N4794, N1283);
and AND2 (N4803, N4800, N3353);
or OR3 (N4804, N4791, N4728, N423);
xor XOR2 (N4805, N4786, N3183);
not NOT1 (N4806, N4796);
nand NAND4 (N4807, N4802, N3354, N2706, N1481);
not NOT1 (N4808, N4803);
nand NAND3 (N4809, N4797, N3081, N4283);
buf BUF1 (N4810, N4806);
not NOT1 (N4811, N4809);
not NOT1 (N4812, N4793);
buf BUF1 (N4813, N4811);
nor NOR2 (N4814, N4792, N4558);
and AND3 (N4815, N4801, N1785, N24);
nand NAND4 (N4816, N4815, N4628, N821, N2882);
nor NOR2 (N4817, N4814, N3508);
nor NOR3 (N4818, N4816, N4608, N3827);
buf BUF1 (N4819, N4808);
not NOT1 (N4820, N4807);
or OR3 (N4821, N4813, N4462, N1089);
xor XOR2 (N4822, N4817, N4249);
and AND2 (N4823, N4733, N847);
and AND4 (N4824, N4821, N663, N2557, N4808);
nand NAND3 (N4825, N4820, N18, N707);
nand NAND2 (N4826, N4819, N703);
nand NAND4 (N4827, N4804, N4343, N1594, N1377);
or OR3 (N4828, N4826, N1242, N2768);
and AND3 (N4829, N4812, N4405, N1460);
or OR3 (N4830, N4810, N3247, N964);
xor XOR2 (N4831, N4829, N2507);
nand NAND2 (N4832, N4831, N3598);
or OR3 (N4833, N4827, N555, N3777);
not NOT1 (N4834, N4818);
buf BUF1 (N4835, N4805);
and AND3 (N4836, N4832, N2223, N2811);
nor NOR3 (N4837, N4834, N1693, N2720);
xor XOR2 (N4838, N4830, N2090);
nand NAND3 (N4839, N4824, N1508, N2391);
nand NAND4 (N4840, N4833, N3451, N1953, N2341);
xor XOR2 (N4841, N4828, N19);
buf BUF1 (N4842, N4839);
xor XOR2 (N4843, N4835, N2903);
not NOT1 (N4844, N4823);
not NOT1 (N4845, N4825);
xor XOR2 (N4846, N4837, N2462);
xor XOR2 (N4847, N4842, N4262);
xor XOR2 (N4848, N4838, N421);
xor XOR2 (N4849, N4841, N1266);
nand NAND4 (N4850, N4845, N1906, N3510, N4399);
and AND2 (N4851, N4844, N1417);
xor XOR2 (N4852, N4847, N2788);
or OR4 (N4853, N4822, N863, N1772, N975);
not NOT1 (N4854, N4836);
buf BUF1 (N4855, N4846);
buf BUF1 (N4856, N4852);
not NOT1 (N4857, N4853);
nand NAND2 (N4858, N4857, N2903);
buf BUF1 (N4859, N4850);
nor NOR3 (N4860, N4840, N191, N3299);
nand NAND2 (N4861, N4858, N4409);
nand NAND3 (N4862, N4860, N3079, N1642);
or OR2 (N4863, N4859, N2277);
or OR3 (N4864, N4854, N1410, N879);
nand NAND3 (N4865, N4856, N2921, N1388);
xor XOR2 (N4866, N4851, N1281);
xor XOR2 (N4867, N4855, N4029);
nor NOR4 (N4868, N4863, N1584, N1002, N265);
buf BUF1 (N4869, N4866);
and AND3 (N4870, N4848, N4464, N2356);
nor NOR2 (N4871, N4865, N3308);
not NOT1 (N4872, N4869);
buf BUF1 (N4873, N4872);
or OR2 (N4874, N4849, N3617);
nor NOR2 (N4875, N4864, N2932);
xor XOR2 (N4876, N4871, N2689);
buf BUF1 (N4877, N4843);
or OR3 (N4878, N4870, N1474, N100);
nor NOR2 (N4879, N4874, N3615);
not NOT1 (N4880, N4877);
xor XOR2 (N4881, N4878, N2465);
nand NAND3 (N4882, N4868, N4375, N2964);
not NOT1 (N4883, N4867);
nor NOR4 (N4884, N4861, N1261, N3213, N217);
not NOT1 (N4885, N4881);
nor NOR3 (N4886, N4862, N2247, N2153);
not NOT1 (N4887, N4876);
nand NAND4 (N4888, N4882, N3929, N4155, N2762);
and AND4 (N4889, N4875, N1186, N553, N1137);
and AND3 (N4890, N4883, N184, N485);
and AND3 (N4891, N4888, N1370, N1694);
and AND4 (N4892, N4873, N268, N1040, N4219);
and AND4 (N4893, N4884, N1304, N3051, N3575);
xor XOR2 (N4894, N4890, N674);
xor XOR2 (N4895, N4894, N2916);
and AND3 (N4896, N4891, N2348, N1426);
nor NOR2 (N4897, N4885, N4659);
buf BUF1 (N4898, N4886);
nand NAND4 (N4899, N4896, N3463, N4634, N2853);
xor XOR2 (N4900, N4892, N3856);
nor NOR3 (N4901, N4897, N4289, N1798);
not NOT1 (N4902, N4900);
or OR2 (N4903, N4901, N3565);
nor NOR4 (N4904, N4893, N210, N3467, N855);
or OR4 (N4905, N4880, N3882, N1065, N2696);
and AND4 (N4906, N4904, N4392, N1894, N2390);
or OR4 (N4907, N4906, N1494, N4126, N3616);
nor NOR2 (N4908, N4898, N285);
not NOT1 (N4909, N4908);
not NOT1 (N4910, N4899);
or OR3 (N4911, N4909, N947, N446);
xor XOR2 (N4912, N4907, N3965);
and AND2 (N4913, N4889, N1455);
nor NOR4 (N4914, N4879, N1825, N87, N1229);
not NOT1 (N4915, N4905);
and AND4 (N4916, N4915, N51, N4377, N697);
nand NAND2 (N4917, N4913, N2785);
nor NOR2 (N4918, N4902, N3911);
or OR3 (N4919, N4910, N4747, N1177);
nor NOR3 (N4920, N4918, N1686, N1472);
and AND3 (N4921, N4919, N2526, N3154);
not NOT1 (N4922, N4914);
buf BUF1 (N4923, N4917);
not NOT1 (N4924, N4923);
and AND4 (N4925, N4916, N1952, N807, N429);
or OR3 (N4926, N4922, N4245, N1340);
not NOT1 (N4927, N4920);
xor XOR2 (N4928, N4895, N2902);
nor NOR2 (N4929, N4887, N2631);
nand NAND3 (N4930, N4927, N3954, N514);
xor XOR2 (N4931, N4928, N2047);
and AND2 (N4932, N4931, N1836);
or OR2 (N4933, N4924, N4795);
xor XOR2 (N4934, N4912, N2134);
xor XOR2 (N4935, N4934, N3347);
nor NOR2 (N4936, N4929, N3053);
xor XOR2 (N4937, N4933, N973);
xor XOR2 (N4938, N4925, N3276);
and AND3 (N4939, N4938, N2890, N2257);
nor NOR4 (N4940, N4937, N1798, N1240, N4882);
buf BUF1 (N4941, N4921);
buf BUF1 (N4942, N4930);
or OR3 (N4943, N4940, N725, N1703);
or OR4 (N4944, N4943, N3753, N2945, N94);
and AND4 (N4945, N4932, N3461, N3100, N4004);
nand NAND4 (N4946, N4911, N4584, N3736, N4177);
or OR2 (N4947, N4926, N2312);
and AND4 (N4948, N4944, N432, N2516, N4168);
or OR4 (N4949, N4948, N4845, N4618, N3201);
buf BUF1 (N4950, N4946);
not NOT1 (N4951, N4941);
nor NOR3 (N4952, N4951, N3366, N4900);
and AND2 (N4953, N4936, N3293);
nand NAND4 (N4954, N4950, N500, N4614, N2361);
nand NAND4 (N4955, N4945, N87, N1650, N3427);
nand NAND4 (N4956, N4942, N1956, N2397, N3058);
not NOT1 (N4957, N4947);
xor XOR2 (N4958, N4949, N2315);
nor NOR3 (N4959, N4955, N3922, N4615);
xor XOR2 (N4960, N4953, N2710);
or OR2 (N4961, N4958, N1438);
nand NAND2 (N4962, N4956, N145);
not NOT1 (N4963, N4939);
nand NAND4 (N4964, N4957, N2694, N2925, N790);
or OR3 (N4965, N4962, N256, N328);
nor NOR4 (N4966, N4960, N2821, N155, N1497);
nand NAND4 (N4967, N4903, N1451, N834, N2110);
and AND3 (N4968, N4966, N4346, N1458);
xor XOR2 (N4969, N4959, N4381);
nand NAND4 (N4970, N4965, N3933, N4148, N1274);
xor XOR2 (N4971, N4970, N4229);
xor XOR2 (N4972, N4969, N1180);
xor XOR2 (N4973, N4952, N126);
and AND4 (N4974, N4971, N453, N4933, N2334);
nor NOR3 (N4975, N4972, N4342, N3484);
and AND4 (N4976, N4968, N1120, N300, N2837);
or OR4 (N4977, N4963, N915, N1523, N4783);
nor NOR3 (N4978, N4977, N2332, N4709);
buf BUF1 (N4979, N4935);
or OR3 (N4980, N4973, N763, N2872);
nand NAND4 (N4981, N4967, N4330, N1840, N2589);
nand NAND2 (N4982, N4964, N3294);
buf BUF1 (N4983, N4981);
xor XOR2 (N4984, N4954, N1194);
nand NAND2 (N4985, N4980, N3005);
nor NOR4 (N4986, N4978, N138, N596, N4213);
nor NOR3 (N4987, N4979, N3978, N2117);
not NOT1 (N4988, N4983);
buf BUF1 (N4989, N4982);
xor XOR2 (N4990, N4974, N1195);
nor NOR4 (N4991, N4985, N673, N2542, N51);
xor XOR2 (N4992, N4976, N1);
nand NAND4 (N4993, N4984, N1137, N444, N235);
buf BUF1 (N4994, N4975);
not NOT1 (N4995, N4989);
nor NOR3 (N4996, N4994, N3865, N3686);
not NOT1 (N4997, N4990);
xor XOR2 (N4998, N4996, N471);
or OR3 (N4999, N4998, N2104, N1868);
nand NAND4 (N5000, N4961, N4909, N4731, N1711);
or OR4 (N5001, N4997, N1135, N1024, N1955);
and AND4 (N5002, N4999, N981, N4626, N4940);
xor XOR2 (N5003, N4987, N1250);
nand NAND2 (N5004, N5000, N3938);
nand NAND3 (N5005, N4993, N1469, N2342);
or OR2 (N5006, N5001, N3358);
nor NOR4 (N5007, N5006, N999, N3493, N549);
nand NAND2 (N5008, N5005, N4281);
or OR4 (N5009, N4986, N247, N2241, N4001);
and AND2 (N5010, N5009, N4558);
nand NAND4 (N5011, N5003, N4631, N2208, N3247);
and AND2 (N5012, N4991, N3731);
nand NAND4 (N5013, N5004, N4394, N1663, N3887);
or OR2 (N5014, N4988, N4404);
buf BUF1 (N5015, N5012);
and AND2 (N5016, N5014, N922);
buf BUF1 (N5017, N4992);
and AND2 (N5018, N5011, N4365);
not NOT1 (N5019, N5010);
buf BUF1 (N5020, N5013);
not NOT1 (N5021, N5019);
nand NAND2 (N5022, N5016, N1916);
nor NOR4 (N5023, N5020, N2989, N542, N915);
xor XOR2 (N5024, N4995, N1175);
or OR2 (N5025, N5002, N3646);
buf BUF1 (N5026, N5023);
buf BUF1 (N5027, N5026);
or OR3 (N5028, N5017, N498, N4718);
xor XOR2 (N5029, N5022, N1025);
buf BUF1 (N5030, N5015);
nand NAND2 (N5031, N5021, N941);
or OR4 (N5032, N5028, N2937, N419, N2687);
xor XOR2 (N5033, N5007, N2546);
buf BUF1 (N5034, N5029);
or OR3 (N5035, N5025, N3233, N3803);
and AND3 (N5036, N5033, N2990, N4150);
buf BUF1 (N5037, N5024);
nor NOR2 (N5038, N5018, N1525);
nand NAND3 (N5039, N5037, N291, N1652);
nand NAND4 (N5040, N5034, N2933, N1525, N4269);
buf BUF1 (N5041, N5036);
xor XOR2 (N5042, N5031, N4568);
not NOT1 (N5043, N5027);
nor NOR2 (N5044, N5038, N825);
and AND4 (N5045, N5039, N779, N4329, N3258);
nor NOR2 (N5046, N5032, N4569);
not NOT1 (N5047, N5030);
nor NOR4 (N5048, N5044, N2648, N4169, N4435);
xor XOR2 (N5049, N5047, N4791);
and AND3 (N5050, N5042, N151, N4445);
nand NAND4 (N5051, N5040, N4359, N925, N2678);
or OR4 (N5052, N5008, N2646, N1758, N1913);
nand NAND2 (N5053, N5050, N3050);
xor XOR2 (N5054, N5053, N2928);
buf BUF1 (N5055, N5048);
nand NAND3 (N5056, N5055, N2032, N1993);
or OR2 (N5057, N5046, N1417);
nor NOR3 (N5058, N5056, N3096, N387);
nand NAND4 (N5059, N5043, N1086, N1966, N4042);
nor NOR3 (N5060, N5041, N3510, N3682);
nor NOR4 (N5061, N5045, N3386, N4205, N4670);
nor NOR2 (N5062, N5059, N3547);
xor XOR2 (N5063, N5058, N742);
nand NAND4 (N5064, N5063, N3796, N3884, N1511);
buf BUF1 (N5065, N5060);
and AND3 (N5066, N5065, N4211, N3378);
buf BUF1 (N5067, N5054);
nor NOR3 (N5068, N5049, N4392, N4605);
or OR2 (N5069, N5052, N1971);
or OR2 (N5070, N5061, N415);
not NOT1 (N5071, N5066);
and AND2 (N5072, N5071, N3137);
buf BUF1 (N5073, N5068);
and AND3 (N5074, N5057, N863, N529);
xor XOR2 (N5075, N5069, N455);
xor XOR2 (N5076, N5075, N1210);
not NOT1 (N5077, N5051);
nand NAND3 (N5078, N5072, N3729, N1327);
nand NAND4 (N5079, N5078, N3984, N3304, N4483);
and AND4 (N5080, N5067, N334, N1418, N574);
nor NOR4 (N5081, N5076, N2289, N1657, N3067);
nor NOR3 (N5082, N5062, N2865, N1293);
buf BUF1 (N5083, N5081);
not NOT1 (N5084, N5077);
not NOT1 (N5085, N5070);
nand NAND4 (N5086, N5084, N171, N3746, N3053);
and AND4 (N5087, N5073, N1647, N970, N191);
not NOT1 (N5088, N5074);
or OR2 (N5089, N5086, N4551);
not NOT1 (N5090, N5064);
xor XOR2 (N5091, N5083, N3330);
nor NOR3 (N5092, N5085, N3307, N3934);
or OR4 (N5093, N5088, N576, N578, N4047);
and AND3 (N5094, N5090, N3575, N2419);
not NOT1 (N5095, N5035);
not NOT1 (N5096, N5093);
nor NOR3 (N5097, N5092, N637, N2025);
not NOT1 (N5098, N5082);
xor XOR2 (N5099, N5079, N126);
not NOT1 (N5100, N5094);
not NOT1 (N5101, N5089);
and AND4 (N5102, N5080, N2745, N4775, N59);
and AND4 (N5103, N5097, N712, N4874, N1753);
not NOT1 (N5104, N5100);
or OR2 (N5105, N5102, N1055);
buf BUF1 (N5106, N5101);
and AND2 (N5107, N5103, N4615);
xor XOR2 (N5108, N5099, N277);
buf BUF1 (N5109, N5105);
and AND3 (N5110, N5091, N915, N282);
buf BUF1 (N5111, N5098);
nand NAND2 (N5112, N5106, N1928);
not NOT1 (N5113, N5104);
not NOT1 (N5114, N5096);
or OR4 (N5115, N5087, N4665, N2074, N1);
not NOT1 (N5116, N5109);
and AND3 (N5117, N5114, N1314, N498);
nor NOR2 (N5118, N5111, N464);
buf BUF1 (N5119, N5118);
buf BUF1 (N5120, N5119);
xor XOR2 (N5121, N5120, N3534);
buf BUF1 (N5122, N5121);
and AND2 (N5123, N5113, N770);
xor XOR2 (N5124, N5108, N2898);
xor XOR2 (N5125, N5112, N3552);
buf BUF1 (N5126, N5117);
and AND4 (N5127, N5115, N3821, N4861, N880);
and AND3 (N5128, N5107, N316, N513);
not NOT1 (N5129, N5123);
not NOT1 (N5130, N5122);
or OR3 (N5131, N5127, N2385, N875);
nand NAND3 (N5132, N5128, N470, N1646);
and AND4 (N5133, N5124, N5027, N3528, N1323);
buf BUF1 (N5134, N5132);
nand NAND4 (N5135, N5110, N3697, N4619, N2563);
or OR2 (N5136, N5126, N3184);
not NOT1 (N5137, N5116);
or OR2 (N5138, N5129, N3951);
nand NAND2 (N5139, N5130, N1038);
and AND4 (N5140, N5131, N4500, N4925, N237);
and AND4 (N5141, N5138, N5051, N604, N4715);
xor XOR2 (N5142, N5125, N4111);
not NOT1 (N5143, N5137);
nor NOR4 (N5144, N5133, N4789, N2181, N2912);
and AND2 (N5145, N5141, N509);
buf BUF1 (N5146, N5142);
buf BUF1 (N5147, N5135);
not NOT1 (N5148, N5145);
buf BUF1 (N5149, N5134);
or OR2 (N5150, N5095, N593);
or OR4 (N5151, N5144, N2963, N2757, N4336);
buf BUF1 (N5152, N5140);
buf BUF1 (N5153, N5136);
nand NAND2 (N5154, N5139, N1138);
and AND4 (N5155, N5151, N5152, N4741, N3287);
nor NOR4 (N5156, N757, N4693, N53, N4173);
xor XOR2 (N5157, N5150, N3776);
or OR3 (N5158, N5148, N2817, N836);
xor XOR2 (N5159, N5143, N4243);
buf BUF1 (N5160, N5149);
nor NOR2 (N5161, N5147, N1233);
nor NOR4 (N5162, N5157, N1410, N4599, N1352);
not NOT1 (N5163, N5160);
or OR4 (N5164, N5146, N2543, N398, N3250);
xor XOR2 (N5165, N5161, N131);
xor XOR2 (N5166, N5162, N4722);
not NOT1 (N5167, N5156);
xor XOR2 (N5168, N5167, N1712);
nor NOR3 (N5169, N5154, N784, N4601);
buf BUF1 (N5170, N5163);
or OR3 (N5171, N5153, N1860, N3079);
and AND4 (N5172, N5165, N5067, N2921, N3930);
or OR2 (N5173, N5170, N3158);
nor NOR2 (N5174, N5159, N373);
nand NAND4 (N5175, N5168, N2470, N2828, N771);
not NOT1 (N5176, N5174);
and AND4 (N5177, N5171, N1921, N1371, N2926);
buf BUF1 (N5178, N5177);
buf BUF1 (N5179, N5175);
not NOT1 (N5180, N5172);
or OR2 (N5181, N5158, N4189);
nand NAND4 (N5182, N5166, N1098, N2067, N2675);
and AND4 (N5183, N5176, N430, N2939, N217);
xor XOR2 (N5184, N5183, N4695);
xor XOR2 (N5185, N5180, N751);
nand NAND2 (N5186, N5155, N3999);
xor XOR2 (N5187, N5184, N3504);
nor NOR3 (N5188, N5187, N554, N887);
xor XOR2 (N5189, N5173, N4234);
xor XOR2 (N5190, N5164, N1036);
nand NAND4 (N5191, N5169, N2040, N2543, N2373);
nand NAND4 (N5192, N5181, N4256, N3148, N4151);
xor XOR2 (N5193, N5186, N1857);
buf BUF1 (N5194, N5191);
buf BUF1 (N5195, N5194);
nor NOR2 (N5196, N5189, N4632);
and AND2 (N5197, N5192, N5180);
nand NAND4 (N5198, N5190, N1069, N3631, N144);
buf BUF1 (N5199, N5196);
nand NAND4 (N5200, N5182, N2882, N4397, N1032);
xor XOR2 (N5201, N5185, N1490);
buf BUF1 (N5202, N5188);
nor NOR2 (N5203, N5198, N5084);
nor NOR3 (N5204, N5199, N2671, N2531);
xor XOR2 (N5205, N5200, N2479);
xor XOR2 (N5206, N5205, N2412);
not NOT1 (N5207, N5204);
nand NAND3 (N5208, N5178, N780, N3020);
nand NAND2 (N5209, N5195, N4796);
nand NAND3 (N5210, N5203, N3361, N4423);
or OR4 (N5211, N5210, N1378, N1510, N3963);
nand NAND4 (N5212, N5179, N3922, N4071, N2568);
and AND3 (N5213, N5206, N1036, N4691);
nor NOR2 (N5214, N5208, N3032);
nor NOR2 (N5215, N5193, N210);
and AND3 (N5216, N5202, N3506, N2825);
nor NOR3 (N5217, N5209, N137, N3207);
nor NOR3 (N5218, N5201, N1125, N110);
xor XOR2 (N5219, N5213, N2523);
and AND3 (N5220, N5216, N5114, N3772);
buf BUF1 (N5221, N5217);
nor NOR3 (N5222, N5220, N230, N1204);
not NOT1 (N5223, N5212);
and AND2 (N5224, N5197, N3751);
nand NAND2 (N5225, N5222, N4842);
nor NOR4 (N5226, N5219, N4689, N1686, N1477);
or OR3 (N5227, N5211, N2812, N2220);
nand NAND2 (N5228, N5224, N5184);
or OR4 (N5229, N5225, N1899, N478, N4632);
nor NOR3 (N5230, N5228, N2282, N3172);
xor XOR2 (N5231, N5227, N483);
nor NOR4 (N5232, N5218, N1732, N4802, N2612);
xor XOR2 (N5233, N5229, N96);
buf BUF1 (N5234, N5207);
nor NOR2 (N5235, N5233, N5010);
xor XOR2 (N5236, N5232, N749);
nor NOR3 (N5237, N5231, N2141, N318);
nor NOR3 (N5238, N5223, N2417, N340);
xor XOR2 (N5239, N5236, N1944);
and AND3 (N5240, N5238, N4212, N3898);
not NOT1 (N5241, N5221);
or OR2 (N5242, N5237, N242);
buf BUF1 (N5243, N5235);
xor XOR2 (N5244, N5226, N554);
nor NOR3 (N5245, N5214, N2394, N2597);
nand NAND4 (N5246, N5240, N992, N1718, N1190);
nor NOR4 (N5247, N5246, N4298, N182, N4614);
buf BUF1 (N5248, N5215);
nor NOR3 (N5249, N5239, N4247, N853);
nor NOR3 (N5250, N5245, N402, N415);
buf BUF1 (N5251, N5234);
nand NAND2 (N5252, N5248, N1695);
and AND3 (N5253, N5241, N5095, N1715);
not NOT1 (N5254, N5253);
and AND3 (N5255, N5251, N359, N2831);
and AND2 (N5256, N5255, N4203);
nand NAND2 (N5257, N5242, N3716);
xor XOR2 (N5258, N5247, N4284);
and AND4 (N5259, N5243, N9, N576, N1349);
nand NAND2 (N5260, N5252, N895);
and AND4 (N5261, N5230, N3955, N5247, N1948);
and AND4 (N5262, N5259, N3562, N2703, N3208);
nand NAND3 (N5263, N5254, N604, N4964);
xor XOR2 (N5264, N5244, N742);
and AND2 (N5265, N5264, N1859);
nor NOR3 (N5266, N5256, N3967, N2087);
nor NOR3 (N5267, N5265, N1470, N504);
nor NOR4 (N5268, N5263, N3327, N1739, N2606);
not NOT1 (N5269, N5258);
xor XOR2 (N5270, N5262, N1311);
or OR2 (N5271, N5249, N2555);
nand NAND3 (N5272, N5268, N4097, N1314);
buf BUF1 (N5273, N5272);
buf BUF1 (N5274, N5260);
nand NAND3 (N5275, N5271, N157, N1673);
not NOT1 (N5276, N5270);
not NOT1 (N5277, N5275);
nor NOR2 (N5278, N5250, N4320);
and AND4 (N5279, N5278, N111, N2045, N1461);
and AND4 (N5280, N5257, N1914, N290, N4162);
or OR2 (N5281, N5279, N4789);
and AND2 (N5282, N5281, N4110);
nand NAND2 (N5283, N5266, N1261);
nor NOR2 (N5284, N5274, N2314);
nand NAND3 (N5285, N5282, N1961, N1413);
and AND4 (N5286, N5273, N2790, N5175, N1203);
xor XOR2 (N5287, N5286, N3662);
and AND4 (N5288, N5284, N887, N2463, N4760);
buf BUF1 (N5289, N5269);
nand NAND4 (N5290, N5285, N3269, N4434, N2584);
and AND3 (N5291, N5287, N4990, N2294);
or OR4 (N5292, N5291, N2528, N5132, N2363);
buf BUF1 (N5293, N5280);
or OR3 (N5294, N5293, N4671, N4729);
nand NAND2 (N5295, N5276, N2129);
nand NAND2 (N5296, N5294, N2734);
and AND4 (N5297, N5283, N1191, N984, N1164);
not NOT1 (N5298, N5296);
buf BUF1 (N5299, N5295);
not NOT1 (N5300, N5288);
nor NOR3 (N5301, N5277, N4600, N4193);
nor NOR3 (N5302, N5299, N991, N3360);
xor XOR2 (N5303, N5289, N4167);
nand NAND3 (N5304, N5297, N3511, N2691);
nand NAND4 (N5305, N5292, N3986, N1996, N941);
and AND4 (N5306, N5301, N3806, N3968, N2715);
nand NAND3 (N5307, N5302, N2973, N3917);
and AND4 (N5308, N5305, N4313, N3534, N2242);
buf BUF1 (N5309, N5267);
and AND2 (N5310, N5309, N945);
nand NAND2 (N5311, N5304, N3221);
nor NOR4 (N5312, N5303, N3460, N1929, N3163);
or OR3 (N5313, N5290, N2619, N2496);
nand NAND3 (N5314, N5306, N2399, N2746);
and AND2 (N5315, N5312, N1461);
buf BUF1 (N5316, N5313);
xor XOR2 (N5317, N5261, N2839);
xor XOR2 (N5318, N5314, N2259);
xor XOR2 (N5319, N5300, N1351);
buf BUF1 (N5320, N5319);
buf BUF1 (N5321, N5316);
nand NAND2 (N5322, N5320, N5274);
or OR4 (N5323, N5321, N469, N1786, N2627);
and AND3 (N5324, N5323, N3102, N5234);
buf BUF1 (N5325, N5322);
nand NAND2 (N5326, N5317, N1087);
buf BUF1 (N5327, N5326);
not NOT1 (N5328, N5307);
xor XOR2 (N5329, N5325, N5192);
not NOT1 (N5330, N5311);
xor XOR2 (N5331, N5324, N949);
nor NOR2 (N5332, N5330, N1923);
not NOT1 (N5333, N5308);
or OR4 (N5334, N5298, N3980, N2475, N4402);
xor XOR2 (N5335, N5315, N2846);
nor NOR3 (N5336, N5331, N1381, N2404);
or OR3 (N5337, N5333, N4325, N1016);
nand NAND3 (N5338, N5329, N1794, N1722);
xor XOR2 (N5339, N5337, N4355);
or OR3 (N5340, N5332, N5135, N1167);
nor NOR2 (N5341, N5327, N1446);
nand NAND3 (N5342, N5335, N2263, N4972);
not NOT1 (N5343, N5310);
not NOT1 (N5344, N5318);
xor XOR2 (N5345, N5328, N5067);
or OR4 (N5346, N5343, N3754, N3943, N3888);
xor XOR2 (N5347, N5339, N3450);
or OR3 (N5348, N5347, N2011, N1562);
buf BUF1 (N5349, N5346);
and AND4 (N5350, N5341, N4166, N4456, N309);
buf BUF1 (N5351, N5338);
xor XOR2 (N5352, N5345, N1510);
not NOT1 (N5353, N5340);
nor NOR2 (N5354, N5342, N1274);
nand NAND3 (N5355, N5336, N3449, N3817);
not NOT1 (N5356, N5351);
or OR3 (N5357, N5354, N2644, N4836);
nor NOR3 (N5358, N5350, N1244, N54);
or OR3 (N5359, N5357, N2654, N82);
buf BUF1 (N5360, N5352);
xor XOR2 (N5361, N5355, N2354);
buf BUF1 (N5362, N5358);
xor XOR2 (N5363, N5353, N1659);
nand NAND2 (N5364, N5356, N4686);
nand NAND4 (N5365, N5344, N3857, N281, N3989);
nand NAND4 (N5366, N5349, N253, N3548, N4384);
nand NAND4 (N5367, N5360, N5123, N1786, N2951);
buf BUF1 (N5368, N5367);
buf BUF1 (N5369, N5368);
buf BUF1 (N5370, N5369);
buf BUF1 (N5371, N5362);
or OR2 (N5372, N5370, N4578);
nor NOR4 (N5373, N5366, N4808, N2255, N3794);
not NOT1 (N5374, N5371);
buf BUF1 (N5375, N5361);
not NOT1 (N5376, N5372);
and AND2 (N5377, N5365, N3354);
not NOT1 (N5378, N5364);
xor XOR2 (N5379, N5378, N4295);
xor XOR2 (N5380, N5374, N3497);
nor NOR4 (N5381, N5348, N3202, N2688, N4851);
nor NOR3 (N5382, N5380, N3273, N3676);
or OR2 (N5383, N5375, N1445);
buf BUF1 (N5384, N5377);
buf BUF1 (N5385, N5383);
xor XOR2 (N5386, N5382, N5251);
not NOT1 (N5387, N5381);
and AND4 (N5388, N5379, N1655, N1926, N173);
and AND2 (N5389, N5384, N577);
buf BUF1 (N5390, N5389);
nor NOR3 (N5391, N5359, N3356, N3910);
or OR4 (N5392, N5385, N3588, N402, N3950);
not NOT1 (N5393, N5386);
or OR3 (N5394, N5388, N5327, N4468);
not NOT1 (N5395, N5391);
xor XOR2 (N5396, N5390, N5152);
not NOT1 (N5397, N5376);
not NOT1 (N5398, N5395);
buf BUF1 (N5399, N5393);
nand NAND2 (N5400, N5398, N4439);
or OR3 (N5401, N5387, N2227, N351);
buf BUF1 (N5402, N5392);
nand NAND3 (N5403, N5394, N3081, N225);
or OR4 (N5404, N5399, N2298, N2491, N3911);
xor XOR2 (N5405, N5397, N2944);
not NOT1 (N5406, N5403);
nor NOR3 (N5407, N5401, N514, N4632);
or OR3 (N5408, N5400, N4866, N16);
buf BUF1 (N5409, N5405);
or OR2 (N5410, N5409, N4986);
nand NAND3 (N5411, N5404, N4260, N3840);
and AND4 (N5412, N5411, N1964, N3282, N2386);
and AND4 (N5413, N5406, N1443, N1565, N1463);
nand NAND2 (N5414, N5408, N4764);
or OR2 (N5415, N5402, N4730);
xor XOR2 (N5416, N5363, N2387);
nor NOR4 (N5417, N5415, N1540, N1758, N1670);
nand NAND3 (N5418, N5412, N3638, N5246);
buf BUF1 (N5419, N5414);
nand NAND3 (N5420, N5410, N5327, N1984);
nand NAND3 (N5421, N5417, N5154, N1196);
not NOT1 (N5422, N5416);
nand NAND2 (N5423, N5407, N4361);
not NOT1 (N5424, N5419);
or OR2 (N5425, N5396, N328);
buf BUF1 (N5426, N5373);
and AND3 (N5427, N5425, N2474, N3619);
buf BUF1 (N5428, N5424);
not NOT1 (N5429, N5334);
and AND4 (N5430, N5423, N2255, N1000, N3082);
not NOT1 (N5431, N5428);
nor NOR3 (N5432, N5422, N1051, N2275);
not NOT1 (N5433, N5432);
nor NOR2 (N5434, N5429, N3525);
nand NAND3 (N5435, N5418, N2366, N542);
xor XOR2 (N5436, N5426, N3636);
nor NOR2 (N5437, N5434, N5420);
or OR2 (N5438, N4115, N3685);
or OR2 (N5439, N5433, N1551);
and AND2 (N5440, N5413, N4053);
or OR2 (N5441, N5438, N1259);
not NOT1 (N5442, N5441);
buf BUF1 (N5443, N5440);
xor XOR2 (N5444, N5431, N3022);
nor NOR2 (N5445, N5439, N4116);
nor NOR4 (N5446, N5436, N5322, N5427, N2158);
nand NAND4 (N5447, N213, N5147, N4240, N1273);
not NOT1 (N5448, N5437);
not NOT1 (N5449, N5442);
xor XOR2 (N5450, N5449, N3715);
or OR3 (N5451, N5430, N2107, N1746);
buf BUF1 (N5452, N5446);
buf BUF1 (N5453, N5448);
or OR4 (N5454, N5453, N2626, N3826, N3223);
buf BUF1 (N5455, N5444);
nor NOR2 (N5456, N5435, N3369);
xor XOR2 (N5457, N5454, N1001);
nand NAND2 (N5458, N5451, N1467);
nor NOR2 (N5459, N5421, N4850);
xor XOR2 (N5460, N5450, N2932);
xor XOR2 (N5461, N5457, N3190);
xor XOR2 (N5462, N5455, N4169);
nand NAND4 (N5463, N5456, N2902, N3967, N515);
buf BUF1 (N5464, N5452);
nor NOR4 (N5465, N5459, N2306, N4578, N3813);
nand NAND4 (N5466, N5460, N4942, N4710, N1858);
xor XOR2 (N5467, N5462, N1065);
or OR3 (N5468, N5465, N3221, N599);
or OR2 (N5469, N5443, N1209);
nand NAND4 (N5470, N5467, N966, N3335, N745);
xor XOR2 (N5471, N5469, N1251);
or OR4 (N5472, N5447, N2520, N802, N2376);
not NOT1 (N5473, N5470);
and AND4 (N5474, N5445, N1282, N4128, N3237);
or OR2 (N5475, N5474, N2492);
xor XOR2 (N5476, N5471, N3849);
and AND2 (N5477, N5472, N5047);
not NOT1 (N5478, N5473);
xor XOR2 (N5479, N5468, N2799);
xor XOR2 (N5480, N5464, N4030);
or OR2 (N5481, N5480, N4769);
xor XOR2 (N5482, N5478, N2060);
nand NAND2 (N5483, N5476, N1207);
and AND3 (N5484, N5461, N882, N2797);
xor XOR2 (N5485, N5463, N3100);
buf BUF1 (N5486, N5475);
xor XOR2 (N5487, N5458, N4548);
buf BUF1 (N5488, N5484);
nand NAND2 (N5489, N5481, N2431);
and AND2 (N5490, N5489, N1515);
buf BUF1 (N5491, N5485);
nor NOR3 (N5492, N5487, N2373, N559);
nand NAND4 (N5493, N5477, N1991, N4671, N5392);
or OR4 (N5494, N5483, N3185, N2103, N147);
nand NAND4 (N5495, N5493, N403, N4167, N4231);
nor NOR3 (N5496, N5479, N1688, N5484);
buf BUF1 (N5497, N5496);
xor XOR2 (N5498, N5490, N1303);
nand NAND2 (N5499, N5482, N966);
nand NAND2 (N5500, N5495, N2988);
not NOT1 (N5501, N5500);
or OR3 (N5502, N5498, N3883, N2159);
buf BUF1 (N5503, N5502);
and AND2 (N5504, N5494, N1007);
nand NAND4 (N5505, N5466, N3801, N3865, N883);
not NOT1 (N5506, N5503);
or OR3 (N5507, N5486, N1988, N740);
xor XOR2 (N5508, N5499, N5019);
xor XOR2 (N5509, N5504, N4698);
not NOT1 (N5510, N5505);
not NOT1 (N5511, N5501);
xor XOR2 (N5512, N5509, N2913);
or OR2 (N5513, N5491, N5475);
or OR3 (N5514, N5512, N3467, N2624);
or OR3 (N5515, N5511, N2351, N1891);
buf BUF1 (N5516, N5488);
xor XOR2 (N5517, N5513, N1769);
xor XOR2 (N5518, N5492, N4549);
not NOT1 (N5519, N5497);
and AND3 (N5520, N5507, N1023, N2032);
buf BUF1 (N5521, N5515);
and AND3 (N5522, N5514, N1750, N4342);
nor NOR4 (N5523, N5516, N4318, N4298, N3999);
not NOT1 (N5524, N5519);
not NOT1 (N5525, N5510);
or OR4 (N5526, N5520, N2416, N4179, N1618);
not NOT1 (N5527, N5518);
or OR4 (N5528, N5525, N3892, N671, N4854);
xor XOR2 (N5529, N5528, N4086);
nand NAND2 (N5530, N5521, N4179);
nor NOR2 (N5531, N5517, N3825);
xor XOR2 (N5532, N5508, N2400);
xor XOR2 (N5533, N5529, N1608);
buf BUF1 (N5534, N5532);
or OR4 (N5535, N5506, N3452, N1103, N3219);
and AND4 (N5536, N5530, N3988, N1747, N255);
or OR4 (N5537, N5531, N976, N1185, N17);
nand NAND3 (N5538, N5524, N3945, N334);
or OR4 (N5539, N5534, N1223, N3293, N2857);
nor NOR2 (N5540, N5523, N1277);
buf BUF1 (N5541, N5538);
xor XOR2 (N5542, N5537, N2900);
and AND2 (N5543, N5539, N1446);
xor XOR2 (N5544, N5526, N5188);
or OR4 (N5545, N5542, N14, N3640, N4811);
nor NOR3 (N5546, N5535, N577, N5303);
nor NOR4 (N5547, N5544, N485, N3820, N2212);
nor NOR2 (N5548, N5533, N4942);
not NOT1 (N5549, N5522);
not NOT1 (N5550, N5543);
not NOT1 (N5551, N5549);
nor NOR4 (N5552, N5547, N3077, N439, N4133);
buf BUF1 (N5553, N5548);
nand NAND3 (N5554, N5540, N3382, N4561);
and AND3 (N5555, N5551, N2360, N3604);
or OR4 (N5556, N5545, N1417, N2321, N91);
buf BUF1 (N5557, N5555);
xor XOR2 (N5558, N5553, N4435);
and AND3 (N5559, N5546, N2434, N5009);
buf BUF1 (N5560, N5556);
and AND4 (N5561, N5550, N2257, N3999, N5544);
or OR3 (N5562, N5561, N3964, N4410);
not NOT1 (N5563, N5559);
xor XOR2 (N5564, N5557, N2608);
not NOT1 (N5565, N5563);
buf BUF1 (N5566, N5565);
not NOT1 (N5567, N5536);
nor NOR4 (N5568, N5554, N972, N2565, N3381);
nor NOR3 (N5569, N5558, N2766, N2265);
nand NAND2 (N5570, N5541, N587);
buf BUF1 (N5571, N5562);
nor NOR2 (N5572, N5571, N4277);
xor XOR2 (N5573, N5560, N402);
nand NAND4 (N5574, N5567, N3829, N2517, N1415);
buf BUF1 (N5575, N5572);
or OR3 (N5576, N5575, N3603, N104);
and AND4 (N5577, N5527, N1590, N1424, N4583);
or OR2 (N5578, N5574, N83);
nand NAND2 (N5579, N5570, N1820);
not NOT1 (N5580, N5573);
or OR4 (N5581, N5579, N4810, N668, N4415);
nand NAND4 (N5582, N5577, N4531, N114, N4400);
buf BUF1 (N5583, N5578);
nand NAND3 (N5584, N5566, N2494, N370);
nor NOR3 (N5585, N5582, N3597, N3693);
and AND2 (N5586, N5552, N4385);
not NOT1 (N5587, N5584);
nand NAND4 (N5588, N5568, N2437, N4224, N1482);
nor NOR4 (N5589, N5588, N4060, N1482, N2416);
or OR2 (N5590, N5576, N848);
and AND4 (N5591, N5564, N5040, N4867, N2166);
not NOT1 (N5592, N5591);
not NOT1 (N5593, N5569);
not NOT1 (N5594, N5592);
xor XOR2 (N5595, N5585, N2221);
nand NAND3 (N5596, N5589, N625, N2691);
nor NOR2 (N5597, N5580, N4893);
buf BUF1 (N5598, N5593);
nor NOR2 (N5599, N5583, N4840);
or OR3 (N5600, N5587, N2960, N3611);
and AND3 (N5601, N5581, N3265, N2376);
and AND4 (N5602, N5594, N58, N4055, N4734);
or OR2 (N5603, N5586, N2985);
or OR3 (N5604, N5597, N5555, N1008);
or OR4 (N5605, N5600, N1221, N2679, N1548);
and AND4 (N5606, N5596, N4552, N3801, N4575);
buf BUF1 (N5607, N5606);
nand NAND2 (N5608, N5601, N1681);
xor XOR2 (N5609, N5602, N4356);
xor XOR2 (N5610, N5599, N2101);
buf BUF1 (N5611, N5590);
not NOT1 (N5612, N5610);
buf BUF1 (N5613, N5607);
not NOT1 (N5614, N5609);
buf BUF1 (N5615, N5598);
buf BUF1 (N5616, N5614);
not NOT1 (N5617, N5612);
nand NAND3 (N5618, N5605, N251, N711);
buf BUF1 (N5619, N5595);
nor NOR3 (N5620, N5618, N3048, N3525);
and AND2 (N5621, N5620, N1707);
buf BUF1 (N5622, N5611);
nand NAND2 (N5623, N5616, N1153);
buf BUF1 (N5624, N5621);
buf BUF1 (N5625, N5622);
nor NOR2 (N5626, N5604, N5001);
nand NAND2 (N5627, N5603, N4157);
buf BUF1 (N5628, N5623);
xor XOR2 (N5629, N5608, N999);
and AND4 (N5630, N5627, N797, N1812, N2430);
or OR3 (N5631, N5613, N4962, N2427);
or OR2 (N5632, N5624, N935);
buf BUF1 (N5633, N5615);
nor NOR4 (N5634, N5630, N1101, N5081, N5195);
nor NOR2 (N5635, N5628, N566);
nor NOR4 (N5636, N5626, N2398, N670, N3681);
nor NOR3 (N5637, N5625, N4307, N5122);
nor NOR4 (N5638, N5619, N3643, N3120, N4045);
and AND4 (N5639, N5635, N975, N4507, N19);
xor XOR2 (N5640, N5617, N2654);
buf BUF1 (N5641, N5639);
xor XOR2 (N5642, N5636, N5014);
and AND4 (N5643, N5637, N2057, N1483, N2286);
buf BUF1 (N5644, N5634);
and AND2 (N5645, N5640, N5301);
xor XOR2 (N5646, N5632, N2195);
not NOT1 (N5647, N5644);
not NOT1 (N5648, N5633);
nand NAND3 (N5649, N5645, N3368, N3876);
and AND2 (N5650, N5638, N2812);
nor NOR2 (N5651, N5648, N5552);
xor XOR2 (N5652, N5629, N3343);
buf BUF1 (N5653, N5650);
and AND2 (N5654, N5642, N1944);
not NOT1 (N5655, N5649);
nand NAND3 (N5656, N5654, N4108, N5068);
buf BUF1 (N5657, N5655);
nor NOR3 (N5658, N5647, N5033, N4143);
nor NOR3 (N5659, N5653, N1472, N5575);
nor NOR4 (N5660, N5652, N489, N3848, N2555);
and AND4 (N5661, N5646, N4118, N2840, N4770);
nand NAND3 (N5662, N5641, N915, N5106);
nor NOR2 (N5663, N5662, N1708);
and AND4 (N5664, N5656, N2894, N4289, N103);
nor NOR4 (N5665, N5664, N4320, N1025, N2870);
nor NOR4 (N5666, N5658, N1200, N2879, N4990);
and AND4 (N5667, N5665, N4920, N2514, N4729);
buf BUF1 (N5668, N5631);
nor NOR4 (N5669, N5659, N3451, N444, N4488);
buf BUF1 (N5670, N5661);
buf BUF1 (N5671, N5663);
xor XOR2 (N5672, N5670, N2383);
or OR2 (N5673, N5667, N2211);
or OR2 (N5674, N5672, N1314);
or OR4 (N5675, N5674, N3959, N5674, N1355);
and AND2 (N5676, N5657, N812);
or OR4 (N5677, N5660, N857, N3144, N1135);
buf BUF1 (N5678, N5669);
and AND3 (N5679, N5673, N1648, N4675);
and AND3 (N5680, N5668, N2263, N3872);
nor NOR4 (N5681, N5666, N604, N3454, N5502);
nor NOR2 (N5682, N5679, N1302);
nor NOR2 (N5683, N5678, N5364);
nand NAND3 (N5684, N5677, N5365, N719);
xor XOR2 (N5685, N5682, N1232);
nor NOR2 (N5686, N5680, N4052);
xor XOR2 (N5687, N5684, N801);
and AND4 (N5688, N5675, N5523, N2645, N1123);
and AND2 (N5689, N5671, N728);
not NOT1 (N5690, N5689);
xor XOR2 (N5691, N5683, N505);
or OR3 (N5692, N5685, N4147, N5424);
buf BUF1 (N5693, N5692);
and AND4 (N5694, N5693, N4450, N3264, N2801);
nor NOR3 (N5695, N5676, N945, N1549);
nor NOR3 (N5696, N5690, N4393, N1839);
xor XOR2 (N5697, N5691, N4570);
buf BUF1 (N5698, N5694);
not NOT1 (N5699, N5697);
nor NOR2 (N5700, N5686, N768);
not NOT1 (N5701, N5696);
nor NOR3 (N5702, N5701, N2891, N2749);
buf BUF1 (N5703, N5681);
not NOT1 (N5704, N5700);
or OR3 (N5705, N5699, N3168, N5224);
not NOT1 (N5706, N5703);
nor NOR4 (N5707, N5695, N4224, N1150, N4888);
nand NAND4 (N5708, N5704, N2859, N1524, N4957);
nor NOR4 (N5709, N5651, N5063, N2378, N13);
buf BUF1 (N5710, N5708);
and AND2 (N5711, N5687, N870);
buf BUF1 (N5712, N5711);
not NOT1 (N5713, N5706);
nand NAND4 (N5714, N5688, N4159, N5015, N4155);
xor XOR2 (N5715, N5714, N2937);
nor NOR4 (N5716, N5710, N3042, N525, N18);
or OR3 (N5717, N5702, N4092, N113);
not NOT1 (N5718, N5707);
xor XOR2 (N5719, N5715, N1064);
nor NOR4 (N5720, N5718, N4436, N4617, N127);
xor XOR2 (N5721, N5720, N3230);
or OR4 (N5722, N5713, N2868, N785, N1543);
or OR4 (N5723, N5716, N1538, N819, N461);
xor XOR2 (N5724, N5698, N1881);
or OR3 (N5725, N5721, N4100, N3140);
buf BUF1 (N5726, N5719);
nor NOR3 (N5727, N5717, N3308, N2046);
nor NOR2 (N5728, N5726, N1191);
nor NOR4 (N5729, N5727, N5557, N1877, N357);
or OR4 (N5730, N5709, N2801, N252, N2786);
xor XOR2 (N5731, N5729, N4363);
not NOT1 (N5732, N5723);
and AND2 (N5733, N5724, N3378);
nand NAND4 (N5734, N5731, N4631, N788, N4983);
or OR4 (N5735, N5722, N3311, N137, N5226);
xor XOR2 (N5736, N5725, N5552);
or OR4 (N5737, N5712, N935, N202, N3627);
or OR3 (N5738, N5736, N1186, N3901);
buf BUF1 (N5739, N5728);
or OR4 (N5740, N5738, N4016, N3309, N1914);
xor XOR2 (N5741, N5735, N1909);
nor NOR2 (N5742, N5739, N1217);
xor XOR2 (N5743, N5732, N974);
not NOT1 (N5744, N5740);
not NOT1 (N5745, N5744);
xor XOR2 (N5746, N5734, N1137);
buf BUF1 (N5747, N5733);
not NOT1 (N5748, N5730);
or OR2 (N5749, N5748, N2864);
and AND3 (N5750, N5749, N1200, N2807);
or OR2 (N5751, N5746, N4389);
nand NAND3 (N5752, N5643, N5105, N5609);
xor XOR2 (N5753, N5745, N4736);
buf BUF1 (N5754, N5742);
not NOT1 (N5755, N5751);
xor XOR2 (N5756, N5755, N777);
or OR4 (N5757, N5737, N3928, N1789, N5328);
not NOT1 (N5758, N5705);
xor XOR2 (N5759, N5752, N1819);
nand NAND2 (N5760, N5743, N5045);
not NOT1 (N5761, N5754);
buf BUF1 (N5762, N5753);
and AND4 (N5763, N5750, N5065, N839, N3804);
and AND3 (N5764, N5759, N2596, N988);
not NOT1 (N5765, N5764);
or OR4 (N5766, N5756, N1496, N26, N1400);
not NOT1 (N5767, N5760);
xor XOR2 (N5768, N5741, N1340);
nand NAND3 (N5769, N5765, N1798, N4676);
xor XOR2 (N5770, N5763, N4571);
and AND3 (N5771, N5768, N783, N4114);
xor XOR2 (N5772, N5762, N4806);
xor XOR2 (N5773, N5770, N1859);
nor NOR2 (N5774, N5771, N1968);
and AND3 (N5775, N5766, N2193, N2049);
or OR2 (N5776, N5773, N3452);
xor XOR2 (N5777, N5772, N508);
and AND3 (N5778, N5769, N938, N3586);
or OR2 (N5779, N5776, N397);
buf BUF1 (N5780, N5758);
and AND3 (N5781, N5775, N3797, N4597);
buf BUF1 (N5782, N5779);
nor NOR2 (N5783, N5777, N3434);
and AND2 (N5784, N5747, N4075);
buf BUF1 (N5785, N5761);
nand NAND3 (N5786, N5757, N1500, N3718);
not NOT1 (N5787, N5782);
buf BUF1 (N5788, N5767);
and AND3 (N5789, N5774, N2156, N2730);
buf BUF1 (N5790, N5789);
buf BUF1 (N5791, N5781);
nand NAND2 (N5792, N5787, N3928);
not NOT1 (N5793, N5788);
or OR3 (N5794, N5786, N102, N357);
nand NAND2 (N5795, N5793, N2491);
nor NOR3 (N5796, N5784, N3768, N4267);
buf BUF1 (N5797, N5795);
buf BUF1 (N5798, N5791);
nand NAND2 (N5799, N5797, N2821);
xor XOR2 (N5800, N5785, N78);
not NOT1 (N5801, N5780);
nor NOR3 (N5802, N5801, N4564, N4111);
xor XOR2 (N5803, N5783, N807);
and AND2 (N5804, N5790, N2724);
buf BUF1 (N5805, N5799);
nand NAND4 (N5806, N5800, N3855, N4380, N1324);
nor NOR2 (N5807, N5778, N5189);
or OR3 (N5808, N5806, N1114, N5482);
nand NAND4 (N5809, N5803, N2801, N3617, N2263);
not NOT1 (N5810, N5805);
buf BUF1 (N5811, N5804);
and AND3 (N5812, N5807, N5214, N3564);
nand NAND3 (N5813, N5811, N5119, N19);
nand NAND4 (N5814, N5798, N3299, N5017, N342);
nand NAND3 (N5815, N5792, N1412, N5079);
buf BUF1 (N5816, N5796);
buf BUF1 (N5817, N5808);
buf BUF1 (N5818, N5814);
nor NOR4 (N5819, N5794, N3766, N3709, N4661);
and AND2 (N5820, N5809, N78);
not NOT1 (N5821, N5812);
buf BUF1 (N5822, N5819);
xor XOR2 (N5823, N5822, N5739);
nand NAND3 (N5824, N5816, N1424, N895);
nor NOR3 (N5825, N5813, N5795, N374);
nor NOR3 (N5826, N5823, N2764, N5316);
buf BUF1 (N5827, N5820);
nor NOR4 (N5828, N5817, N3861, N1451, N1144);
nand NAND3 (N5829, N5818, N3718, N4697);
nand NAND3 (N5830, N5828, N2568, N2548);
buf BUF1 (N5831, N5830);
nand NAND3 (N5832, N5815, N2126, N5764);
or OR3 (N5833, N5810, N4073, N4979);
xor XOR2 (N5834, N5825, N2230);
not NOT1 (N5835, N5831);
not NOT1 (N5836, N5835);
or OR2 (N5837, N5824, N501);
nand NAND2 (N5838, N5832, N3313);
nor NOR4 (N5839, N5836, N825, N5039, N5022);
nand NAND2 (N5840, N5802, N3971);
buf BUF1 (N5841, N5826);
nand NAND4 (N5842, N5837, N3474, N1523, N5338);
or OR3 (N5843, N5838, N276, N1986);
nand NAND2 (N5844, N5834, N3585);
not NOT1 (N5845, N5841);
buf BUF1 (N5846, N5821);
buf BUF1 (N5847, N5827);
nand NAND2 (N5848, N5845, N1040);
not NOT1 (N5849, N5847);
not NOT1 (N5850, N5829);
buf BUF1 (N5851, N5839);
and AND2 (N5852, N5846, N5516);
buf BUF1 (N5853, N5842);
nor NOR4 (N5854, N5843, N5056, N100, N4045);
buf BUF1 (N5855, N5844);
nand NAND2 (N5856, N5855, N2715);
xor XOR2 (N5857, N5840, N4908);
or OR2 (N5858, N5853, N1293);
not NOT1 (N5859, N5850);
xor XOR2 (N5860, N5857, N587);
or OR2 (N5861, N5859, N3027);
nand NAND2 (N5862, N5860, N5595);
not NOT1 (N5863, N5858);
or OR3 (N5864, N5856, N5578, N1450);
nor NOR4 (N5865, N5854, N3898, N5365, N2420);
not NOT1 (N5866, N5833);
not NOT1 (N5867, N5861);
not NOT1 (N5868, N5867);
not NOT1 (N5869, N5849);
nand NAND4 (N5870, N5865, N3527, N5335, N3851);
not NOT1 (N5871, N5870);
xor XOR2 (N5872, N5848, N912);
or OR3 (N5873, N5851, N1557, N3489);
not NOT1 (N5874, N5866);
nand NAND4 (N5875, N5874, N777, N2916, N4289);
or OR3 (N5876, N5864, N4791, N3267);
or OR4 (N5877, N5876, N1206, N2618, N3748);
buf BUF1 (N5878, N5868);
xor XOR2 (N5879, N5878, N1030);
not NOT1 (N5880, N5877);
nor NOR4 (N5881, N5869, N5757, N3176, N5493);
not NOT1 (N5882, N5863);
not NOT1 (N5883, N5872);
xor XOR2 (N5884, N5879, N115);
xor XOR2 (N5885, N5881, N3616);
nor NOR2 (N5886, N5875, N2560);
not NOT1 (N5887, N5886);
buf BUF1 (N5888, N5887);
or OR2 (N5889, N5880, N468);
not NOT1 (N5890, N5882);
nor NOR3 (N5891, N5888, N3638, N3950);
and AND2 (N5892, N5862, N2320);
not NOT1 (N5893, N5885);
nand NAND2 (N5894, N5891, N3687);
nand NAND2 (N5895, N5893, N3828);
buf BUF1 (N5896, N5890);
buf BUF1 (N5897, N5889);
and AND3 (N5898, N5873, N5883, N60);
nand NAND2 (N5899, N2120, N5069);
nor NOR3 (N5900, N5884, N2949, N858);
nand NAND2 (N5901, N5899, N2202);
and AND4 (N5902, N5896, N4353, N2075, N990);
buf BUF1 (N5903, N5901);
not NOT1 (N5904, N5895);
not NOT1 (N5905, N5897);
and AND3 (N5906, N5852, N2293, N5427);
xor XOR2 (N5907, N5894, N1520);
or OR3 (N5908, N5904, N927, N1447);
nand NAND4 (N5909, N5908, N3151, N3294, N3550);
and AND2 (N5910, N5900, N621);
nor NOR2 (N5911, N5907, N2202);
or OR2 (N5912, N5871, N3286);
xor XOR2 (N5913, N5910, N718);
not NOT1 (N5914, N5909);
buf BUF1 (N5915, N5903);
nand NAND4 (N5916, N5912, N556, N5601, N645);
buf BUF1 (N5917, N5916);
nand NAND2 (N5918, N5905, N3960);
nor NOR4 (N5919, N5898, N1247, N5711, N3964);
xor XOR2 (N5920, N5915, N2875);
nor NOR4 (N5921, N5906, N3275, N4672, N5326);
xor XOR2 (N5922, N5919, N2595);
or OR2 (N5923, N5922, N1924);
buf BUF1 (N5924, N5913);
buf BUF1 (N5925, N5911);
not NOT1 (N5926, N5892);
nor NOR2 (N5927, N5926, N4052);
nand NAND4 (N5928, N5921, N194, N3486, N2050);
buf BUF1 (N5929, N5914);
nor NOR4 (N5930, N5918, N1322, N1292, N2615);
nand NAND3 (N5931, N5924, N2210, N4385);
not NOT1 (N5932, N5927);
buf BUF1 (N5933, N5928);
not NOT1 (N5934, N5932);
not NOT1 (N5935, N5934);
buf BUF1 (N5936, N5902);
nand NAND2 (N5937, N5923, N4247);
and AND3 (N5938, N5936, N3313, N5841);
and AND3 (N5939, N5931, N5791, N4543);
xor XOR2 (N5940, N5935, N1285);
xor XOR2 (N5941, N5939, N2483);
not NOT1 (N5942, N5933);
and AND3 (N5943, N5929, N2584, N4991);
or OR4 (N5944, N5937, N246, N4725, N3440);
or OR4 (N5945, N5942, N1340, N2224, N3307);
nor NOR4 (N5946, N5938, N5913, N1856, N4443);
nand NAND4 (N5947, N5941, N3305, N1440, N3503);
not NOT1 (N5948, N5945);
or OR4 (N5949, N5940, N4067, N4001, N92);
nand NAND4 (N5950, N5947, N4869, N2058, N1503);
buf BUF1 (N5951, N5925);
nand NAND2 (N5952, N5946, N1997);
buf BUF1 (N5953, N5949);
xor XOR2 (N5954, N5948, N3989);
buf BUF1 (N5955, N5953);
nand NAND3 (N5956, N5950, N2565, N1473);
nand NAND2 (N5957, N5952, N3850);
or OR3 (N5958, N5957, N3987, N5687);
and AND4 (N5959, N5958, N795, N2808, N4698);
and AND2 (N5960, N5920, N2984);
and AND3 (N5961, N5930, N973, N4985);
or OR3 (N5962, N5951, N2754, N5646);
nand NAND4 (N5963, N5959, N4052, N2116, N5382);
not NOT1 (N5964, N5962);
buf BUF1 (N5965, N5954);
or OR3 (N5966, N5964, N4994, N2325);
buf BUF1 (N5967, N5943);
and AND4 (N5968, N5966, N582, N1719, N3042);
or OR3 (N5969, N5956, N2459, N3964);
or OR3 (N5970, N5963, N1649, N65);
nor NOR2 (N5971, N5967, N4452);
nand NAND2 (N5972, N5969, N4501);
or OR4 (N5973, N5971, N2756, N4856, N1715);
not NOT1 (N5974, N5917);
not NOT1 (N5975, N5974);
not NOT1 (N5976, N5973);
and AND3 (N5977, N5955, N2364, N2107);
not NOT1 (N5978, N5976);
not NOT1 (N5979, N5977);
xor XOR2 (N5980, N5972, N5347);
or OR2 (N5981, N5978, N1683);
nor NOR2 (N5982, N5960, N4300);
nand NAND3 (N5983, N5970, N296, N1212);
xor XOR2 (N5984, N5983, N3677);
xor XOR2 (N5985, N5944, N5912);
not NOT1 (N5986, N5968);
nand NAND2 (N5987, N5985, N5558);
nand NAND2 (N5988, N5981, N831);
and AND4 (N5989, N5987, N1329, N3420, N4407);
nand NAND3 (N5990, N5982, N5939, N3762);
nand NAND2 (N5991, N5980, N3539);
nand NAND2 (N5992, N5965, N2637);
nor NOR4 (N5993, N5992, N2350, N4481, N2378);
xor XOR2 (N5994, N5991, N4533);
or OR2 (N5995, N5984, N2281);
nand NAND4 (N5996, N5994, N1892, N5412, N1435);
and AND3 (N5997, N5996, N5489, N5468);
not NOT1 (N5998, N5995);
and AND4 (N5999, N5961, N5262, N2684, N5455);
xor XOR2 (N6000, N5998, N2446);
and AND2 (N6001, N6000, N3026);
buf BUF1 (N6002, N5990);
nand NAND4 (N6003, N5988, N4222, N5986, N2668);
and AND2 (N6004, N944, N890);
nor NOR3 (N6005, N6003, N2575, N5611);
or OR2 (N6006, N5979, N2840);
not NOT1 (N6007, N6005);
buf BUF1 (N6008, N6004);
nand NAND4 (N6009, N6002, N2747, N2869, N1977);
and AND4 (N6010, N5975, N5165, N1440, N5344);
buf BUF1 (N6011, N5999);
nor NOR4 (N6012, N6006, N179, N266, N5126);
buf BUF1 (N6013, N6007);
not NOT1 (N6014, N6012);
nor NOR2 (N6015, N5997, N1551);
buf BUF1 (N6016, N6014);
buf BUF1 (N6017, N6008);
and AND3 (N6018, N6010, N1281, N3015);
and AND4 (N6019, N6017, N815, N5340, N4980);
xor XOR2 (N6020, N6016, N1805);
nor NOR3 (N6021, N6009, N45, N3230);
nand NAND4 (N6022, N6015, N4985, N3186, N1955);
buf BUF1 (N6023, N6011);
buf BUF1 (N6024, N6022);
nand NAND2 (N6025, N5989, N372);
not NOT1 (N6026, N6020);
xor XOR2 (N6027, N6021, N2224);
xor XOR2 (N6028, N6001, N1003);
not NOT1 (N6029, N6013);
not NOT1 (N6030, N6027);
or OR4 (N6031, N6025, N5009, N145, N3770);
or OR3 (N6032, N6018, N2490, N3896);
buf BUF1 (N6033, N6030);
or OR4 (N6034, N6023, N5889, N4371, N2102);
nor NOR3 (N6035, N6024, N5078, N5275);
nor NOR2 (N6036, N6019, N3611);
and AND2 (N6037, N6031, N5556);
buf BUF1 (N6038, N6035);
or OR2 (N6039, N6038, N1748);
and AND3 (N6040, N6037, N2194, N4067);
and AND2 (N6041, N6040, N2231);
buf BUF1 (N6042, N6028);
nand NAND3 (N6043, N6036, N1791, N2949);
buf BUF1 (N6044, N6041);
nor NOR4 (N6045, N6029, N5592, N4561, N2920);
buf BUF1 (N6046, N6032);
nand NAND4 (N6047, N6039, N4741, N6, N84);
buf BUF1 (N6048, N6026);
xor XOR2 (N6049, N6046, N3561);
xor XOR2 (N6050, N6034, N3432);
not NOT1 (N6051, N6042);
nand NAND3 (N6052, N6044, N1205, N591);
nand NAND3 (N6053, N6052, N3295, N4700);
and AND4 (N6054, N6048, N902, N2132, N1494);
and AND3 (N6055, N6045, N5779, N3385);
buf BUF1 (N6056, N5993);
not NOT1 (N6057, N6050);
xor XOR2 (N6058, N6055, N3462);
buf BUF1 (N6059, N6054);
nor NOR4 (N6060, N6053, N3659, N5896, N5726);
or OR2 (N6061, N6059, N5634);
xor XOR2 (N6062, N6057, N4921);
nand NAND2 (N6063, N6056, N2789);
and AND4 (N6064, N6063, N101, N4192, N3889);
or OR3 (N6065, N6047, N3892, N791);
nor NOR4 (N6066, N6058, N1806, N2353, N1896);
nand NAND4 (N6067, N6033, N3015, N3044, N1665);
xor XOR2 (N6068, N6064, N5065);
nor NOR3 (N6069, N6060, N2804, N4460);
xor XOR2 (N6070, N6067, N4952);
xor XOR2 (N6071, N6049, N2071);
nand NAND4 (N6072, N6062, N1417, N2956, N3287);
and AND3 (N6073, N6066, N617, N5019);
nand NAND2 (N6074, N6069, N5865);
buf BUF1 (N6075, N6068);
not NOT1 (N6076, N6065);
buf BUF1 (N6077, N6061);
nor NOR2 (N6078, N6075, N2947);
or OR3 (N6079, N6076, N351, N2424);
nand NAND2 (N6080, N6077, N4831);
nand NAND3 (N6081, N6074, N5061, N2276);
xor XOR2 (N6082, N6078, N2806);
nor NOR4 (N6083, N6072, N864, N1465, N2087);
not NOT1 (N6084, N6083);
or OR2 (N6085, N6043, N1831);
xor XOR2 (N6086, N6070, N5803);
or OR4 (N6087, N6086, N268, N2817, N2693);
buf BUF1 (N6088, N6079);
and AND4 (N6089, N6082, N4783, N250, N2992);
or OR2 (N6090, N6051, N399);
nor NOR3 (N6091, N6085, N2421, N4398);
nand NAND2 (N6092, N6090, N1940);
or OR3 (N6093, N6091, N437, N5438);
not NOT1 (N6094, N6089);
not NOT1 (N6095, N6080);
xor XOR2 (N6096, N6092, N5439);
xor XOR2 (N6097, N6087, N4985);
and AND2 (N6098, N6084, N1170);
xor XOR2 (N6099, N6073, N4488);
xor XOR2 (N6100, N6093, N1672);
nand NAND4 (N6101, N6096, N5484, N502, N4176);
and AND4 (N6102, N6094, N1429, N3950, N4130);
xor XOR2 (N6103, N6099, N1979);
not NOT1 (N6104, N6103);
nor NOR4 (N6105, N6100, N4435, N735, N5060);
nor NOR2 (N6106, N6105, N1318);
nor NOR4 (N6107, N6104, N4055, N6013, N930);
not NOT1 (N6108, N6095);
nand NAND3 (N6109, N6098, N4518, N5030);
nand NAND3 (N6110, N6071, N1380, N714);
and AND3 (N6111, N6110, N3562, N5302);
xor XOR2 (N6112, N6102, N1);
xor XOR2 (N6113, N6106, N560);
or OR2 (N6114, N6088, N1014);
or OR2 (N6115, N6109, N2862);
nor NOR4 (N6116, N6101, N3797, N5089, N4080);
or OR2 (N6117, N6116, N1420);
xor XOR2 (N6118, N6107, N371);
buf BUF1 (N6119, N6117);
buf BUF1 (N6120, N6114);
or OR4 (N6121, N6108, N3027, N3551, N3200);
nor NOR4 (N6122, N6118, N1143, N2500, N1640);
nor NOR2 (N6123, N6113, N1743);
nor NOR4 (N6124, N6123, N1106, N863, N4815);
xor XOR2 (N6125, N6115, N346);
buf BUF1 (N6126, N6120);
nand NAND3 (N6127, N6119, N5498, N5996);
or OR4 (N6128, N6081, N5997, N3730, N5864);
buf BUF1 (N6129, N6121);
not NOT1 (N6130, N6122);
not NOT1 (N6131, N6112);
or OR2 (N6132, N6127, N1523);
and AND4 (N6133, N6097, N3765, N5894, N5894);
and AND2 (N6134, N6129, N627);
not NOT1 (N6135, N6125);
or OR2 (N6136, N6128, N3508);
nand NAND2 (N6137, N6135, N283);
buf BUF1 (N6138, N6134);
or OR4 (N6139, N6138, N3203, N3768, N5338);
nand NAND3 (N6140, N6111, N2162, N915);
nand NAND3 (N6141, N6132, N1974, N118);
or OR4 (N6142, N6137, N5193, N2499, N159);
or OR3 (N6143, N6124, N4816, N2557);
and AND2 (N6144, N6143, N2112);
xor XOR2 (N6145, N6142, N2361);
buf BUF1 (N6146, N6130);
buf BUF1 (N6147, N6126);
or OR4 (N6148, N6133, N1732, N1965, N2056);
nor NOR3 (N6149, N6131, N4144, N2654);
and AND2 (N6150, N6139, N843);
or OR2 (N6151, N6145, N73);
buf BUF1 (N6152, N6150);
nand NAND3 (N6153, N6148, N292, N4092);
not NOT1 (N6154, N6144);
nand NAND3 (N6155, N6146, N5909, N1829);
buf BUF1 (N6156, N6151);
or OR3 (N6157, N6147, N11, N3385);
nor NOR2 (N6158, N6136, N5632);
nor NOR2 (N6159, N6156, N281);
xor XOR2 (N6160, N6157, N1720);
and AND2 (N6161, N6140, N992);
nor NOR3 (N6162, N6155, N2391, N441);
and AND3 (N6163, N6154, N148, N5153);
nand NAND2 (N6164, N6160, N1013);
not NOT1 (N6165, N6163);
nor NOR3 (N6166, N6164, N5764, N5651);
nor NOR3 (N6167, N6162, N3539, N5097);
nand NAND3 (N6168, N6166, N1542, N197);
nand NAND4 (N6169, N6149, N6046, N2197, N2839);
or OR4 (N6170, N6153, N3706, N5041, N4103);
and AND3 (N6171, N6167, N405, N3330);
and AND2 (N6172, N6171, N106);
not NOT1 (N6173, N6168);
buf BUF1 (N6174, N6172);
buf BUF1 (N6175, N6158);
buf BUF1 (N6176, N6175);
and AND4 (N6177, N6152, N833, N4474, N4637);
not NOT1 (N6178, N6170);
nor NOR3 (N6179, N6176, N4373, N1338);
or OR2 (N6180, N6177, N5654);
or OR3 (N6181, N6173, N529, N3670);
buf BUF1 (N6182, N6169);
or OR3 (N6183, N6141, N2216, N1534);
and AND4 (N6184, N6183, N5070, N6013, N2514);
nand NAND2 (N6185, N6161, N5605);
not NOT1 (N6186, N6165);
nand NAND4 (N6187, N6181, N1402, N5074, N1504);
or OR4 (N6188, N6186, N6070, N3391, N1245);
and AND4 (N6189, N6188, N4908, N2293, N5599);
buf BUF1 (N6190, N6179);
buf BUF1 (N6191, N6182);
nand NAND4 (N6192, N6191, N3741, N4209, N6034);
and AND4 (N6193, N6180, N3662, N345, N3780);
nand NAND3 (N6194, N6178, N3081, N5330);
buf BUF1 (N6195, N6174);
and AND3 (N6196, N6189, N4160, N751);
and AND3 (N6197, N6185, N4786, N5997);
and AND3 (N6198, N6190, N1776, N2011);
nor NOR2 (N6199, N6184, N2793);
not NOT1 (N6200, N6159);
nor NOR3 (N6201, N6196, N5916, N5605);
nor NOR3 (N6202, N6187, N1543, N3400);
not NOT1 (N6203, N6202);
and AND2 (N6204, N6192, N5985);
not NOT1 (N6205, N6204);
or OR4 (N6206, N6203, N1271, N3418, N2876);
or OR3 (N6207, N6197, N4298, N3522);
or OR4 (N6208, N6206, N1799, N38, N1221);
or OR4 (N6209, N6198, N4845, N3014, N340);
or OR3 (N6210, N6193, N1929, N3070);
or OR4 (N6211, N6209, N2480, N6057, N5391);
nor NOR4 (N6212, N6205, N389, N6045, N700);
buf BUF1 (N6213, N6211);
and AND4 (N6214, N6199, N3012, N3618, N4469);
buf BUF1 (N6215, N6210);
and AND4 (N6216, N6195, N4146, N1744, N4592);
or OR2 (N6217, N6212, N4894);
nor NOR2 (N6218, N6201, N1245);
and AND3 (N6219, N6194, N4009, N4681);
or OR2 (N6220, N6214, N3027);
not NOT1 (N6221, N6219);
nor NOR4 (N6222, N6217, N262, N2006, N5467);
buf BUF1 (N6223, N6213);
or OR3 (N6224, N6221, N234, N3112);
nand NAND3 (N6225, N6207, N5881, N695);
nand NAND2 (N6226, N6223, N1380);
and AND3 (N6227, N6225, N2315, N1802);
and AND2 (N6228, N6200, N4877);
or OR3 (N6229, N6215, N310, N5151);
and AND3 (N6230, N6227, N4106, N795);
or OR4 (N6231, N6228, N5469, N4858, N3217);
nor NOR3 (N6232, N6231, N164, N1302);
and AND4 (N6233, N6230, N5909, N3148, N2525);
nor NOR3 (N6234, N6226, N3767, N2049);
nand NAND2 (N6235, N6218, N960);
or OR4 (N6236, N6208, N528, N3513, N4544);
not NOT1 (N6237, N6233);
or OR2 (N6238, N6220, N4406);
nor NOR3 (N6239, N6238, N46, N5024);
nor NOR4 (N6240, N6216, N898, N29, N265);
and AND4 (N6241, N6239, N4407, N5025, N3209);
nand NAND2 (N6242, N6235, N1379);
xor XOR2 (N6243, N6232, N4877);
or OR3 (N6244, N6240, N1559, N4941);
or OR4 (N6245, N6241, N2562, N2176, N2023);
buf BUF1 (N6246, N6242);
or OR2 (N6247, N6246, N4284);
not NOT1 (N6248, N6224);
nand NAND4 (N6249, N6248, N4638, N5292, N3756);
xor XOR2 (N6250, N6229, N4424);
or OR3 (N6251, N6245, N1546, N2547);
buf BUF1 (N6252, N6249);
or OR3 (N6253, N6251, N3819, N794);
and AND2 (N6254, N6250, N5023);
or OR3 (N6255, N6253, N2562, N1868);
or OR3 (N6256, N6236, N4162, N3972);
and AND3 (N6257, N6255, N3065, N2669);
and AND2 (N6258, N6254, N356);
or OR4 (N6259, N6234, N2484, N4380, N2528);
and AND3 (N6260, N6252, N1168, N2602);
buf BUF1 (N6261, N6257);
xor XOR2 (N6262, N6243, N1087);
buf BUF1 (N6263, N6258);
nor NOR4 (N6264, N6237, N184, N1974, N1110);
or OR3 (N6265, N6222, N1013, N1407);
or OR4 (N6266, N6256, N3163, N5526, N790);
and AND3 (N6267, N6265, N1960, N2430);
and AND2 (N6268, N6259, N53);
or OR2 (N6269, N6264, N2014);
nand NAND2 (N6270, N6266, N5888);
and AND2 (N6271, N6269, N2227);
not NOT1 (N6272, N6268);
and AND4 (N6273, N6244, N6168, N853, N5254);
or OR3 (N6274, N6247, N2276, N5481);
not NOT1 (N6275, N6271);
nor NOR3 (N6276, N6275, N4223, N2590);
nor NOR2 (N6277, N6261, N2295);
not NOT1 (N6278, N6272);
nor NOR3 (N6279, N6263, N2579, N4310);
nor NOR3 (N6280, N6262, N4865, N3911);
nand NAND2 (N6281, N6276, N2778);
xor XOR2 (N6282, N6274, N3918);
xor XOR2 (N6283, N6278, N5599);
nand NAND3 (N6284, N6283, N1011, N429);
xor XOR2 (N6285, N6281, N1493);
nor NOR2 (N6286, N6277, N736);
buf BUF1 (N6287, N6260);
buf BUF1 (N6288, N6284);
and AND3 (N6289, N6287, N2056, N5566);
or OR3 (N6290, N6289, N3724, N771);
xor XOR2 (N6291, N6290, N3238);
and AND4 (N6292, N6270, N3358, N4760, N5683);
not NOT1 (N6293, N6282);
buf BUF1 (N6294, N6267);
or OR2 (N6295, N6292, N5365);
nand NAND4 (N6296, N6288, N2046, N6023, N2179);
or OR2 (N6297, N6296, N5661);
or OR4 (N6298, N6297, N3502, N540, N4278);
or OR2 (N6299, N6279, N2278);
xor XOR2 (N6300, N6286, N585);
xor XOR2 (N6301, N6298, N953);
not NOT1 (N6302, N6300);
or OR2 (N6303, N6302, N6261);
and AND2 (N6304, N6291, N1005);
not NOT1 (N6305, N6273);
xor XOR2 (N6306, N6305, N5813);
nand NAND3 (N6307, N6304, N3377, N5082);
nor NOR4 (N6308, N6294, N2368, N2202, N4889);
nor NOR4 (N6309, N6293, N1102, N1718, N1310);
nor NOR3 (N6310, N6299, N2555, N4073);
buf BUF1 (N6311, N6285);
not NOT1 (N6312, N6280);
or OR2 (N6313, N6307, N3482);
or OR2 (N6314, N6312, N4436);
and AND2 (N6315, N6311, N4134);
or OR3 (N6316, N6301, N18, N6002);
nand NAND3 (N6317, N6315, N3297, N5859);
xor XOR2 (N6318, N6303, N2576);
nand NAND3 (N6319, N6313, N3445, N4514);
nor NOR2 (N6320, N6295, N808);
xor XOR2 (N6321, N6309, N6166);
nor NOR4 (N6322, N6321, N3042, N5610, N1408);
nand NAND4 (N6323, N6318, N1294, N4601, N3232);
and AND3 (N6324, N6306, N1465, N1230);
buf BUF1 (N6325, N6308);
nand NAND4 (N6326, N6319, N6316, N215, N4588);
and AND4 (N6327, N6231, N5684, N1301, N4470);
and AND2 (N6328, N6317, N2274);
or OR2 (N6329, N6325, N1135);
not NOT1 (N6330, N6314);
nand NAND4 (N6331, N6328, N3272, N4764, N2146);
nor NOR4 (N6332, N6324, N5858, N4916, N627);
and AND3 (N6333, N6320, N3931, N3499);
buf BUF1 (N6334, N6329);
and AND2 (N6335, N6327, N4044);
or OR2 (N6336, N6322, N3094);
not NOT1 (N6337, N6333);
nand NAND3 (N6338, N6331, N6081, N5321);
not NOT1 (N6339, N6330);
xor XOR2 (N6340, N6334, N3239);
or OR4 (N6341, N6338, N4267, N5698, N4969);
buf BUF1 (N6342, N6341);
and AND2 (N6343, N6332, N3485);
xor XOR2 (N6344, N6326, N4830);
nand NAND4 (N6345, N6336, N4387, N239, N3334);
or OR2 (N6346, N6343, N719);
nor NOR4 (N6347, N6346, N5201, N151, N4275);
nor NOR2 (N6348, N6340, N1501);
buf BUF1 (N6349, N6323);
nand NAND4 (N6350, N6337, N5535, N5578, N714);
or OR2 (N6351, N6342, N5155);
not NOT1 (N6352, N6335);
not NOT1 (N6353, N6350);
buf BUF1 (N6354, N6349);
nor NOR3 (N6355, N6310, N97, N5064);
nand NAND3 (N6356, N6354, N3411, N400);
or OR2 (N6357, N6352, N3000);
nand NAND2 (N6358, N6353, N5902);
not NOT1 (N6359, N6355);
and AND2 (N6360, N6348, N1179);
xor XOR2 (N6361, N6345, N5403);
nor NOR3 (N6362, N6344, N518, N3268);
nand NAND4 (N6363, N6358, N2898, N1529, N3592);
buf BUF1 (N6364, N6339);
nand NAND4 (N6365, N6357, N261, N977, N1767);
nand NAND3 (N6366, N6351, N4351, N4756);
nand NAND2 (N6367, N6366, N2760);
nand NAND2 (N6368, N6363, N3156);
buf BUF1 (N6369, N6362);
nor NOR2 (N6370, N6360, N886);
not NOT1 (N6371, N6367);
nor NOR2 (N6372, N6369, N374);
or OR3 (N6373, N6371, N3609, N2372);
or OR4 (N6374, N6370, N4914, N906, N2201);
nor NOR4 (N6375, N6368, N2523, N2378, N2462);
nor NOR4 (N6376, N6375, N1163, N5233, N5388);
nand NAND4 (N6377, N6376, N5469, N774, N26);
and AND3 (N6378, N6347, N115, N859);
and AND2 (N6379, N6365, N4541);
nand NAND3 (N6380, N6378, N1484, N1446);
or OR4 (N6381, N6359, N4599, N4403, N3545);
not NOT1 (N6382, N6377);
xor XOR2 (N6383, N6381, N230);
or OR4 (N6384, N6356, N819, N4976, N3751);
buf BUF1 (N6385, N6373);
not NOT1 (N6386, N6374);
and AND4 (N6387, N6382, N5504, N1187, N2036);
or OR4 (N6388, N6386, N1424, N4075, N1530);
and AND2 (N6389, N6364, N6325);
and AND3 (N6390, N6380, N173, N3784);
nor NOR3 (N6391, N6384, N524, N3216);
not NOT1 (N6392, N6383);
or OR3 (N6393, N6361, N2679, N1368);
and AND4 (N6394, N6392, N404, N5404, N2258);
nand NAND2 (N6395, N6379, N4176);
and AND2 (N6396, N6393, N4992);
or OR2 (N6397, N6391, N1196);
nand NAND4 (N6398, N6389, N1564, N2362, N4430);
nand NAND2 (N6399, N6395, N2086);
nand NAND3 (N6400, N6387, N1547, N758);
or OR4 (N6401, N6388, N3166, N3597, N6113);
xor XOR2 (N6402, N6385, N237);
buf BUF1 (N6403, N6402);
nor NOR4 (N6404, N6372, N4012, N1016, N1382);
nand NAND2 (N6405, N6394, N2257);
nor NOR3 (N6406, N6403, N3643, N5228);
not NOT1 (N6407, N6405);
and AND2 (N6408, N6399, N2803);
buf BUF1 (N6409, N6404);
xor XOR2 (N6410, N6401, N3237);
nor NOR2 (N6411, N6408, N3746);
not NOT1 (N6412, N6410);
buf BUF1 (N6413, N6397);
xor XOR2 (N6414, N6413, N4250);
buf BUF1 (N6415, N6407);
nor NOR3 (N6416, N6409, N1605, N1535);
nand NAND2 (N6417, N6396, N5400);
buf BUF1 (N6418, N6411);
buf BUF1 (N6419, N6398);
or OR2 (N6420, N6412, N3);
xor XOR2 (N6421, N6414, N4552);
nand NAND2 (N6422, N6416, N5092);
nand NAND3 (N6423, N6418, N5684, N1395);
not NOT1 (N6424, N6390);
xor XOR2 (N6425, N6420, N5962);
not NOT1 (N6426, N6423);
nand NAND2 (N6427, N6426, N5504);
buf BUF1 (N6428, N6421);
buf BUF1 (N6429, N6415);
xor XOR2 (N6430, N6422, N1982);
or OR2 (N6431, N6430, N2733);
or OR2 (N6432, N6417, N4964);
nand NAND2 (N6433, N6429, N1111);
nand NAND2 (N6434, N6432, N1788);
and AND4 (N6435, N6431, N2959, N4973, N3877);
not NOT1 (N6436, N6435);
and AND3 (N6437, N6424, N2013, N3022);
or OR2 (N6438, N6400, N5747);
and AND4 (N6439, N6438, N4481, N5786, N434);
xor XOR2 (N6440, N6419, N3596);
not NOT1 (N6441, N6425);
and AND4 (N6442, N6406, N3804, N1232, N624);
not NOT1 (N6443, N6437);
buf BUF1 (N6444, N6428);
nand NAND2 (N6445, N6434, N5735);
and AND2 (N6446, N6443, N1575);
buf BUF1 (N6447, N6427);
and AND2 (N6448, N6445, N1011);
not NOT1 (N6449, N6447);
buf BUF1 (N6450, N6441);
nand NAND2 (N6451, N6448, N4405);
or OR2 (N6452, N6436, N4419);
nor NOR3 (N6453, N6433, N2570, N665);
not NOT1 (N6454, N6451);
nand NAND4 (N6455, N6454, N3613, N832, N6280);
nor NOR3 (N6456, N6452, N2800, N4709);
buf BUF1 (N6457, N6444);
nand NAND2 (N6458, N6449, N604);
nand NAND4 (N6459, N6453, N4459, N6071, N2389);
xor XOR2 (N6460, N6446, N437);
and AND2 (N6461, N6442, N6164);
or OR3 (N6462, N6440, N4555, N5937);
buf BUF1 (N6463, N6459);
or OR3 (N6464, N6455, N1392, N5727);
nand NAND3 (N6465, N6439, N2319, N188);
nor NOR4 (N6466, N6458, N6211, N660, N2178);
xor XOR2 (N6467, N6460, N5606);
nand NAND4 (N6468, N6465, N544, N4202, N6353);
buf BUF1 (N6469, N6466);
xor XOR2 (N6470, N6461, N388);
nor NOR3 (N6471, N6469, N32, N1323);
or OR4 (N6472, N6470, N4879, N1518, N4824);
or OR4 (N6473, N6463, N2307, N1587, N6403);
xor XOR2 (N6474, N6457, N2571);
nor NOR3 (N6475, N6450, N5457, N5167);
nor NOR2 (N6476, N6472, N2662);
and AND2 (N6477, N6475, N3172);
not NOT1 (N6478, N6471);
nand NAND3 (N6479, N6476, N2137, N5608);
nor NOR2 (N6480, N6467, N4382);
nand NAND3 (N6481, N6478, N4327, N3234);
nand NAND3 (N6482, N6462, N61, N5823);
and AND3 (N6483, N6482, N5759, N4123);
nor NOR4 (N6484, N6477, N978, N4223, N3153);
and AND4 (N6485, N6464, N5960, N159, N5129);
nor NOR3 (N6486, N6485, N443, N2361);
and AND4 (N6487, N6456, N1998, N4905, N5498);
xor XOR2 (N6488, N6481, N6446);
xor XOR2 (N6489, N6468, N3825);
buf BUF1 (N6490, N6474);
nand NAND2 (N6491, N6490, N5691);
nand NAND3 (N6492, N6479, N1632, N2186);
buf BUF1 (N6493, N6492);
nor NOR4 (N6494, N6483, N3927, N5549, N2422);
xor XOR2 (N6495, N6489, N5429);
and AND3 (N6496, N6491, N2809, N98);
not NOT1 (N6497, N6488);
xor XOR2 (N6498, N6497, N2969);
not NOT1 (N6499, N6494);
not NOT1 (N6500, N6498);
not NOT1 (N6501, N6473);
not NOT1 (N6502, N6499);
buf BUF1 (N6503, N6496);
or OR2 (N6504, N6495, N5096);
buf BUF1 (N6505, N6487);
or OR3 (N6506, N6504, N6450, N62);
nand NAND4 (N6507, N6505, N1928, N5238, N761);
or OR2 (N6508, N6500, N4459);
and AND3 (N6509, N6503, N4829, N4126);
nor NOR4 (N6510, N6484, N1972, N6295, N287);
and AND2 (N6511, N6510, N95);
xor XOR2 (N6512, N6502, N4600);
and AND2 (N6513, N6486, N3826);
xor XOR2 (N6514, N6509, N157);
or OR3 (N6515, N6507, N2213, N5024);
xor XOR2 (N6516, N6511, N1977);
nand NAND4 (N6517, N6480, N3224, N4918, N531);
not NOT1 (N6518, N6493);
buf BUF1 (N6519, N6501);
or OR3 (N6520, N6513, N4565, N3691);
nand NAND4 (N6521, N6516, N5460, N4885, N3269);
buf BUF1 (N6522, N6508);
or OR4 (N6523, N6506, N1457, N5447, N2022);
not NOT1 (N6524, N6520);
not NOT1 (N6525, N6521);
not NOT1 (N6526, N6515);
nor NOR4 (N6527, N6519, N1090, N1171, N4740);
nor NOR2 (N6528, N6524, N3427);
buf BUF1 (N6529, N6518);
xor XOR2 (N6530, N6526, N3791);
nor NOR4 (N6531, N6522, N3388, N2303, N3556);
xor XOR2 (N6532, N6512, N3723);
not NOT1 (N6533, N6527);
not NOT1 (N6534, N6531);
nand NAND3 (N6535, N6534, N5283, N5774);
nor NOR4 (N6536, N6528, N6501, N2553, N4469);
and AND3 (N6537, N6530, N5070, N5125);
not NOT1 (N6538, N6535);
or OR3 (N6539, N6532, N4882, N3270);
nor NOR3 (N6540, N6529, N1129, N4311);
or OR4 (N6541, N6537, N158, N2759, N5541);
xor XOR2 (N6542, N6517, N73);
nor NOR2 (N6543, N6525, N2164);
nand NAND2 (N6544, N6542, N1958);
and AND4 (N6545, N6543, N2603, N231, N2705);
not NOT1 (N6546, N6541);
xor XOR2 (N6547, N6533, N1641);
or OR2 (N6548, N6546, N6105);
nor NOR4 (N6549, N6536, N3582, N1934, N6004);
nand NAND3 (N6550, N6539, N3438, N2598);
nand NAND4 (N6551, N6548, N1952, N4421, N5216);
nand NAND2 (N6552, N6549, N2565);
not NOT1 (N6553, N6545);
nor NOR4 (N6554, N6553, N2597, N3786, N5946);
buf BUF1 (N6555, N6547);
or OR3 (N6556, N6550, N2934, N4045);
not NOT1 (N6557, N6540);
or OR4 (N6558, N6523, N3232, N6005, N4801);
not NOT1 (N6559, N6552);
nand NAND4 (N6560, N6544, N5901, N544, N4589);
or OR3 (N6561, N6560, N507, N4074);
nand NAND2 (N6562, N6514, N2938);
buf BUF1 (N6563, N6561);
nor NOR2 (N6564, N6551, N1523);
buf BUF1 (N6565, N6557);
not NOT1 (N6566, N6564);
nand NAND3 (N6567, N6563, N4138, N3554);
nor NOR3 (N6568, N6559, N747, N5067);
or OR3 (N6569, N6555, N20, N3431);
nand NAND2 (N6570, N6568, N1963);
and AND4 (N6571, N6562, N2520, N2110, N916);
nand NAND4 (N6572, N6565, N810, N3299, N2953);
and AND3 (N6573, N6554, N6033, N2013);
xor XOR2 (N6574, N6567, N4807);
not NOT1 (N6575, N6566);
or OR3 (N6576, N6570, N3924, N6235);
nor NOR3 (N6577, N6575, N682, N1985);
xor XOR2 (N6578, N6576, N3851);
and AND2 (N6579, N6556, N2563);
and AND3 (N6580, N6538, N467, N3551);
xor XOR2 (N6581, N6579, N642);
not NOT1 (N6582, N6571);
and AND2 (N6583, N6573, N5714);
not NOT1 (N6584, N6577);
not NOT1 (N6585, N6582);
nand NAND3 (N6586, N6585, N2204, N1420);
nand NAND3 (N6587, N6583, N1369, N1723);
nand NAND4 (N6588, N6587, N5315, N1503, N1411);
not NOT1 (N6589, N6558);
or OR2 (N6590, N6589, N1899);
and AND2 (N6591, N6569, N5907);
nand NAND2 (N6592, N6580, N2614);
nor NOR3 (N6593, N6578, N628, N5750);
xor XOR2 (N6594, N6590, N838);
nand NAND3 (N6595, N6588, N6476, N2825);
nand NAND3 (N6596, N6584, N3416, N3831);
nor NOR3 (N6597, N6574, N1240, N946);
nor NOR3 (N6598, N6592, N2605, N3261);
nor NOR3 (N6599, N6593, N1015, N1314);
or OR4 (N6600, N6595, N2976, N853, N83);
or OR2 (N6601, N6591, N3490);
xor XOR2 (N6602, N6596, N670);
nand NAND4 (N6603, N6598, N6583, N5536, N4372);
not NOT1 (N6604, N6603);
not NOT1 (N6605, N6594);
and AND4 (N6606, N6581, N5318, N2889, N2536);
and AND2 (N6607, N6597, N1912);
or OR2 (N6608, N6604, N171);
and AND4 (N6609, N6601, N2250, N6003, N2501);
nand NAND3 (N6610, N6606, N3543, N5600);
or OR2 (N6611, N6572, N5172);
nand NAND3 (N6612, N6586, N2348, N1445);
nor NOR4 (N6613, N6607, N4247, N1840, N1635);
and AND4 (N6614, N6599, N4756, N2274, N253);
nand NAND3 (N6615, N6613, N6552, N664);
buf BUF1 (N6616, N6609);
and AND3 (N6617, N6612, N2722, N467);
not NOT1 (N6618, N6602);
xor XOR2 (N6619, N6610, N1989);
and AND3 (N6620, N6611, N1664, N2877);
nand NAND4 (N6621, N6600, N3963, N3875, N852);
xor XOR2 (N6622, N6616, N5252);
not NOT1 (N6623, N6618);
nand NAND3 (N6624, N6617, N2601, N1915);
not NOT1 (N6625, N6619);
nand NAND3 (N6626, N6622, N5423, N3958);
not NOT1 (N6627, N6621);
nor NOR4 (N6628, N6626, N3651, N5504, N1454);
nor NOR4 (N6629, N6624, N5694, N5960, N5926);
buf BUF1 (N6630, N6620);
nand NAND2 (N6631, N6608, N6422);
nand NAND4 (N6632, N6628, N4541, N5533, N2403);
buf BUF1 (N6633, N6614);
or OR4 (N6634, N6615, N3103, N6539, N479);
buf BUF1 (N6635, N6627);
nor NOR2 (N6636, N6635, N2391);
or OR3 (N6637, N6630, N3491, N4293);
not NOT1 (N6638, N6629);
and AND4 (N6639, N6636, N2568, N3447, N5079);
and AND2 (N6640, N6637, N6636);
or OR2 (N6641, N6625, N2175);
not NOT1 (N6642, N6633);
or OR3 (N6643, N6642, N3850, N1091);
not NOT1 (N6644, N6641);
or OR3 (N6645, N6640, N2193, N60);
nand NAND4 (N6646, N6644, N6186, N5312, N748);
xor XOR2 (N6647, N6643, N3829);
nor NOR2 (N6648, N6605, N126);
nand NAND4 (N6649, N6623, N2840, N3125, N3430);
nand NAND4 (N6650, N6646, N829, N4921, N5101);
xor XOR2 (N6651, N6650, N5858);
or OR3 (N6652, N6648, N3259, N5495);
nor NOR4 (N6653, N6652, N1968, N1360, N5682);
and AND4 (N6654, N6632, N5374, N5791, N5601);
and AND4 (N6655, N6639, N1772, N316, N3034);
or OR2 (N6656, N6638, N2423);
buf BUF1 (N6657, N6647);
not NOT1 (N6658, N6653);
nand NAND2 (N6659, N6634, N1879);
buf BUF1 (N6660, N6656);
buf BUF1 (N6661, N6655);
xor XOR2 (N6662, N6631, N6225);
xor XOR2 (N6663, N6660, N2642);
buf BUF1 (N6664, N6663);
nor NOR2 (N6665, N6664, N4237);
buf BUF1 (N6666, N6665);
nor NOR4 (N6667, N6661, N1048, N3123, N3932);
buf BUF1 (N6668, N6658);
nor NOR2 (N6669, N6666, N1229);
not NOT1 (N6670, N6668);
nand NAND4 (N6671, N6654, N6088, N6043, N756);
buf BUF1 (N6672, N6651);
xor XOR2 (N6673, N6645, N5117);
buf BUF1 (N6674, N6662);
not NOT1 (N6675, N6669);
buf BUF1 (N6676, N6674);
xor XOR2 (N6677, N6670, N3936);
or OR2 (N6678, N6671, N1935);
xor XOR2 (N6679, N6657, N4560);
and AND2 (N6680, N6678, N5554);
not NOT1 (N6681, N6676);
or OR2 (N6682, N6649, N626);
and AND2 (N6683, N6659, N4060);
xor XOR2 (N6684, N6677, N921);
buf BUF1 (N6685, N6684);
nor NOR4 (N6686, N6673, N1746, N2555, N3607);
or OR3 (N6687, N6682, N1176, N5648);
nand NAND3 (N6688, N6680, N3255, N2646);
buf BUF1 (N6689, N6672);
or OR2 (N6690, N6686, N2177);
buf BUF1 (N6691, N6667);
and AND3 (N6692, N6685, N4394, N3883);
and AND4 (N6693, N6688, N4494, N3621, N2432);
nor NOR4 (N6694, N6679, N594, N1076, N3879);
or OR2 (N6695, N6687, N2756);
not NOT1 (N6696, N6681);
nand NAND2 (N6697, N6689, N4626);
buf BUF1 (N6698, N6696);
buf BUF1 (N6699, N6693);
not NOT1 (N6700, N6699);
or OR3 (N6701, N6690, N5183, N2635);
nand NAND3 (N6702, N6692, N2089, N5187);
or OR3 (N6703, N6697, N3166, N2232);
not NOT1 (N6704, N6683);
nand NAND2 (N6705, N6702, N3231);
and AND2 (N6706, N6704, N2030);
nand NAND4 (N6707, N6706, N2854, N5454, N4889);
xor XOR2 (N6708, N6698, N6301);
nor NOR2 (N6709, N6705, N4331);
and AND3 (N6710, N6701, N6149, N6537);
buf BUF1 (N6711, N6695);
and AND3 (N6712, N6710, N24, N3945);
nor NOR3 (N6713, N6703, N1206, N3250);
or OR4 (N6714, N6709, N3745, N642, N5175);
nand NAND3 (N6715, N6707, N3119, N5412);
nand NAND4 (N6716, N6712, N4955, N5445, N1008);
nand NAND2 (N6717, N6711, N4920);
nor NOR3 (N6718, N6691, N313, N2066);
nor NOR3 (N6719, N6713, N3212, N3743);
not NOT1 (N6720, N6719);
nor NOR4 (N6721, N6714, N5125, N2216, N4122);
or OR3 (N6722, N6715, N4914, N4301);
or OR3 (N6723, N6716, N3553, N5935);
or OR4 (N6724, N6722, N5903, N2315, N6461);
nor NOR2 (N6725, N6724, N993);
nor NOR2 (N6726, N6720, N174);
and AND2 (N6727, N6717, N4999);
not NOT1 (N6728, N6708);
buf BUF1 (N6729, N6727);
nand NAND2 (N6730, N6675, N5824);
buf BUF1 (N6731, N6694);
nand NAND3 (N6732, N6700, N3595, N2692);
xor XOR2 (N6733, N6726, N4522);
xor XOR2 (N6734, N6723, N2715);
or OR2 (N6735, N6732, N5715);
nor NOR3 (N6736, N6734, N3366, N1275);
xor XOR2 (N6737, N6736, N1328);
or OR2 (N6738, N6729, N1910);
or OR2 (N6739, N6737, N4623);
nand NAND4 (N6740, N6728, N3513, N6484, N244);
not NOT1 (N6741, N6718);
not NOT1 (N6742, N6735);
or OR3 (N6743, N6738, N1328, N579);
xor XOR2 (N6744, N6741, N4387);
nor NOR2 (N6745, N6742, N897);
and AND4 (N6746, N6740, N2798, N583, N5933);
and AND3 (N6747, N6745, N2634, N179);
and AND3 (N6748, N6739, N5002, N1136);
not NOT1 (N6749, N6747);
nor NOR2 (N6750, N6743, N4770);
xor XOR2 (N6751, N6750, N2709);
xor XOR2 (N6752, N6748, N5040);
and AND2 (N6753, N6721, N6214);
nor NOR4 (N6754, N6731, N271, N572, N334);
or OR3 (N6755, N6733, N6490, N339);
nor NOR2 (N6756, N6730, N5809);
not NOT1 (N6757, N6744);
not NOT1 (N6758, N6752);
nor NOR3 (N6759, N6755, N5645, N6);
or OR4 (N6760, N6749, N5566, N4993, N2753);
and AND2 (N6761, N6757, N6352);
nor NOR4 (N6762, N6758, N2440, N1226, N908);
buf BUF1 (N6763, N6754);
xor XOR2 (N6764, N6746, N4678);
not NOT1 (N6765, N6761);
not NOT1 (N6766, N6753);
not NOT1 (N6767, N6766);
nor NOR4 (N6768, N6725, N509, N3084, N2853);
nor NOR4 (N6769, N6763, N5335, N6348, N6708);
and AND3 (N6770, N6764, N6601, N4085);
xor XOR2 (N6771, N6760, N278);
buf BUF1 (N6772, N6762);
nand NAND4 (N6773, N6756, N654, N2896, N6056);
or OR3 (N6774, N6772, N3508, N4770);
or OR4 (N6775, N6770, N5786, N5950, N4466);
and AND3 (N6776, N6769, N2728, N4522);
nor NOR3 (N6777, N6775, N3656, N5795);
nand NAND2 (N6778, N6765, N1180);
and AND4 (N6779, N6777, N3295, N4628, N3205);
buf BUF1 (N6780, N6768);
nand NAND2 (N6781, N6778, N5180);
buf BUF1 (N6782, N6776);
nor NOR3 (N6783, N6782, N6148, N2830);
not NOT1 (N6784, N6783);
nand NAND2 (N6785, N6774, N5024);
not NOT1 (N6786, N6784);
and AND4 (N6787, N6759, N4539, N1583, N2977);
or OR4 (N6788, N6767, N2231, N1931, N609);
nand NAND3 (N6789, N6788, N1235, N6786);
not NOT1 (N6790, N4038);
and AND2 (N6791, N6780, N2009);
or OR3 (N6792, N6771, N3689, N884);
and AND4 (N6793, N6785, N3253, N5745, N4967);
nor NOR4 (N6794, N6793, N3920, N2735, N5649);
and AND4 (N6795, N6792, N2131, N67, N4437);
nor NOR4 (N6796, N6794, N2782, N476, N2015);
not NOT1 (N6797, N6781);
or OR4 (N6798, N6797, N5835, N19, N6195);
not NOT1 (N6799, N6796);
xor XOR2 (N6800, N6787, N6627);
and AND2 (N6801, N6773, N2255);
nand NAND3 (N6802, N6795, N1676, N6033);
xor XOR2 (N6803, N6802, N4546);
or OR2 (N6804, N6789, N4692);
nor NOR2 (N6805, N6791, N1678);
nand NAND4 (N6806, N6790, N4137, N5354, N1748);
nor NOR3 (N6807, N6798, N5144, N6152);
buf BUF1 (N6808, N6803);
and AND2 (N6809, N6805, N4605);
xor XOR2 (N6810, N6806, N5095);
xor XOR2 (N6811, N6800, N4034);
buf BUF1 (N6812, N6801);
not NOT1 (N6813, N6807);
nand NAND4 (N6814, N6779, N3212, N5522, N66);
and AND4 (N6815, N6809, N2698, N3933, N76);
and AND2 (N6816, N6812, N335);
nand NAND3 (N6817, N6813, N3712, N3778);
or OR4 (N6818, N6804, N1889, N2968, N3356);
buf BUF1 (N6819, N6814);
not NOT1 (N6820, N6818);
buf BUF1 (N6821, N6816);
buf BUF1 (N6822, N6817);
and AND4 (N6823, N6815, N6680, N3425, N1088);
and AND3 (N6824, N6811, N4133, N5033);
not NOT1 (N6825, N6821);
buf BUF1 (N6826, N6824);
and AND2 (N6827, N6822, N6771);
buf BUF1 (N6828, N6820);
buf BUF1 (N6829, N6808);
xor XOR2 (N6830, N6799, N6433);
or OR4 (N6831, N6810, N2781, N2323, N1568);
xor XOR2 (N6832, N6825, N1023);
xor XOR2 (N6833, N6829, N3627);
buf BUF1 (N6834, N6828);
xor XOR2 (N6835, N6834, N596);
and AND3 (N6836, N6833, N538, N4325);
nand NAND3 (N6837, N6826, N2674, N5414);
nor NOR4 (N6838, N6835, N2735, N6798, N5145);
and AND3 (N6839, N6823, N2351, N4383);
buf BUF1 (N6840, N6819);
buf BUF1 (N6841, N6838);
buf BUF1 (N6842, N6827);
not NOT1 (N6843, N6832);
buf BUF1 (N6844, N6843);
nand NAND3 (N6845, N6842, N1870, N2926);
xor XOR2 (N6846, N6839, N2152);
and AND2 (N6847, N6841, N3710);
nor NOR2 (N6848, N6845, N2774);
not NOT1 (N6849, N6831);
and AND2 (N6850, N6848, N258);
nand NAND4 (N6851, N6836, N6438, N4516, N2993);
xor XOR2 (N6852, N6850, N1253);
nand NAND2 (N6853, N6851, N655);
nand NAND3 (N6854, N6840, N3040, N3873);
and AND4 (N6855, N6849, N2814, N585, N1951);
xor XOR2 (N6856, N6844, N2880);
nand NAND4 (N6857, N6852, N2693, N5302, N2878);
nand NAND4 (N6858, N6837, N5230, N691, N840);
buf BUF1 (N6859, N6854);
buf BUF1 (N6860, N6858);
nor NOR2 (N6861, N6830, N1990);
or OR4 (N6862, N6847, N5885, N1036, N5302);
xor XOR2 (N6863, N6860, N3717);
xor XOR2 (N6864, N6855, N4005);
not NOT1 (N6865, N6853);
or OR2 (N6866, N6862, N6796);
not NOT1 (N6867, N6846);
buf BUF1 (N6868, N6867);
or OR2 (N6869, N6859, N5869);
not NOT1 (N6870, N6869);
nand NAND3 (N6871, N6751, N2708, N4144);
or OR2 (N6872, N6863, N3752);
nor NOR3 (N6873, N6870, N2164, N302);
buf BUF1 (N6874, N6856);
not NOT1 (N6875, N6868);
nand NAND2 (N6876, N6873, N4497);
and AND2 (N6877, N6865, N2272);
or OR4 (N6878, N6864, N3814, N6466, N1486);
xor XOR2 (N6879, N6877, N3140);
or OR4 (N6880, N6874, N2670, N279, N3354);
nand NAND2 (N6881, N6857, N3990);
xor XOR2 (N6882, N6881, N4113);
nor NOR2 (N6883, N6882, N4689);
nand NAND3 (N6884, N6872, N2280, N4812);
nor NOR3 (N6885, N6871, N962, N1354);
xor XOR2 (N6886, N6875, N1692);
xor XOR2 (N6887, N6879, N893);
nor NOR4 (N6888, N6885, N1880, N5809, N970);
nand NAND3 (N6889, N6887, N262, N144);
not NOT1 (N6890, N6878);
nand NAND4 (N6891, N6880, N3700, N179, N1974);
nor NOR4 (N6892, N6866, N4923, N685, N4359);
and AND3 (N6893, N6892, N4428, N879);
or OR4 (N6894, N6891, N2253, N5493, N5108);
nand NAND3 (N6895, N6884, N575, N4165);
and AND3 (N6896, N6893, N1081, N5773);
buf BUF1 (N6897, N6896);
not NOT1 (N6898, N6894);
or OR2 (N6899, N6883, N5444);
xor XOR2 (N6900, N6861, N2444);
and AND4 (N6901, N6890, N5488, N3394, N1408);
not NOT1 (N6902, N6899);
xor XOR2 (N6903, N6901, N4954);
or OR3 (N6904, N6903, N5661, N4847);
and AND3 (N6905, N6897, N2266, N5090);
xor XOR2 (N6906, N6876, N1034);
nor NOR3 (N6907, N6902, N1890, N2165);
xor XOR2 (N6908, N6906, N1238);
or OR2 (N6909, N6908, N6231);
nor NOR2 (N6910, N6889, N106);
or OR4 (N6911, N6898, N3530, N3069, N1415);
nand NAND4 (N6912, N6900, N2588, N1015, N765);
xor XOR2 (N6913, N6886, N435);
or OR4 (N6914, N6909, N2266, N1024, N3356);
or OR3 (N6915, N6907, N535, N4627);
nand NAND4 (N6916, N6911, N6400, N457, N2368);
nand NAND4 (N6917, N6913, N6718, N196, N2123);
buf BUF1 (N6918, N6915);
not NOT1 (N6919, N6888);
nand NAND3 (N6920, N6919, N1495, N3650);
nor NOR2 (N6921, N6920, N6796);
buf BUF1 (N6922, N6905);
nor NOR4 (N6923, N6914, N809, N1974, N4370);
nor NOR3 (N6924, N6910, N2790, N355);
not NOT1 (N6925, N6921);
and AND3 (N6926, N6904, N3509, N4825);
nor NOR2 (N6927, N6925, N5837);
buf BUF1 (N6928, N6923);
or OR3 (N6929, N6895, N3137, N2804);
nand NAND2 (N6930, N6918, N3827);
and AND2 (N6931, N6922, N1315);
nand NAND2 (N6932, N6917, N3829);
buf BUF1 (N6933, N6928);
or OR2 (N6934, N6930, N3945);
not NOT1 (N6935, N6912);
or OR4 (N6936, N6933, N3393, N3393, N3273);
buf BUF1 (N6937, N6916);
nor NOR3 (N6938, N6931, N5708, N3089);
buf BUF1 (N6939, N6936);
nor NOR2 (N6940, N6938, N5110);
buf BUF1 (N6941, N6926);
nand NAND3 (N6942, N6927, N6391, N3739);
not NOT1 (N6943, N6941);
or OR4 (N6944, N6929, N6302, N3064, N1430);
xor XOR2 (N6945, N6940, N3400);
and AND4 (N6946, N6924, N6352, N1602, N5969);
and AND2 (N6947, N6935, N1856);
xor XOR2 (N6948, N6939, N4687);
or OR4 (N6949, N6937, N5566, N3045, N2939);
or OR3 (N6950, N6948, N3689, N4732);
not NOT1 (N6951, N6934);
buf BUF1 (N6952, N6945);
xor XOR2 (N6953, N6947, N2436);
not NOT1 (N6954, N6953);
and AND2 (N6955, N6952, N2474);
buf BUF1 (N6956, N6949);
nand NAND3 (N6957, N6932, N2074, N987);
not NOT1 (N6958, N6955);
buf BUF1 (N6959, N6956);
and AND4 (N6960, N6943, N4387, N2439, N4352);
nor NOR4 (N6961, N6958, N6629, N597, N6932);
not NOT1 (N6962, N6946);
buf BUF1 (N6963, N6944);
buf BUF1 (N6964, N6959);
buf BUF1 (N6965, N6951);
buf BUF1 (N6966, N6960);
buf BUF1 (N6967, N6962);
nor NOR3 (N6968, N6957, N4220, N6545);
xor XOR2 (N6969, N6968, N1332);
xor XOR2 (N6970, N6950, N2578);
or OR3 (N6971, N6963, N1744, N775);
or OR4 (N6972, N6965, N5280, N38, N1315);
xor XOR2 (N6973, N6967, N4400);
nor NOR4 (N6974, N6973, N6292, N2090, N6235);
not NOT1 (N6975, N6961);
and AND3 (N6976, N6970, N5236, N1054);
nor NOR2 (N6977, N6969, N5092);
nor NOR3 (N6978, N6964, N6439, N1691);
or OR2 (N6979, N6978, N5520);
nand NAND4 (N6980, N6976, N6447, N6140, N3737);
not NOT1 (N6981, N6971);
or OR3 (N6982, N6980, N314, N650);
not NOT1 (N6983, N6966);
nor NOR3 (N6984, N6942, N2543, N6558);
buf BUF1 (N6985, N6972);
and AND2 (N6986, N6982, N5258);
nand NAND4 (N6987, N6983, N2657, N3524, N4216);
not NOT1 (N6988, N6954);
and AND2 (N6989, N6975, N3700);
and AND4 (N6990, N6977, N2020, N6350, N3995);
or OR2 (N6991, N6984, N5995);
nand NAND4 (N6992, N6979, N2743, N4730, N2940);
nor NOR2 (N6993, N6989, N5144);
nor NOR4 (N6994, N6988, N1447, N4888, N554);
or OR3 (N6995, N6985, N5285, N1977);
nand NAND3 (N6996, N6995, N468, N2999);
or OR3 (N6997, N6987, N1534, N4933);
nor NOR4 (N6998, N6994, N489, N3999, N1309);
xor XOR2 (N6999, N6974, N3395);
or OR2 (N7000, N6999, N5420);
xor XOR2 (N7001, N7000, N1435);
nand NAND4 (N7002, N6993, N265, N2885, N385);
or OR2 (N7003, N6992, N2544);
not NOT1 (N7004, N6986);
nand NAND3 (N7005, N6981, N6350, N1748);
xor XOR2 (N7006, N6998, N5830);
buf BUF1 (N7007, N6990);
not NOT1 (N7008, N7007);
nor NOR4 (N7009, N7001, N3965, N975, N345);
and AND3 (N7010, N7002, N4945, N1232);
xor XOR2 (N7011, N7005, N3261);
not NOT1 (N7012, N6997);
buf BUF1 (N7013, N7006);
nor NOR4 (N7014, N7012, N1435, N122, N2660);
and AND4 (N7015, N6996, N2641, N2291, N614);
nand NAND4 (N7016, N7010, N3740, N1017, N2164);
buf BUF1 (N7017, N7016);
not NOT1 (N7018, N7013);
xor XOR2 (N7019, N7008, N5078);
xor XOR2 (N7020, N7017, N6092);
or OR4 (N7021, N7003, N4456, N380, N2935);
or OR4 (N7022, N7021, N1885, N5336, N4505);
or OR2 (N7023, N6991, N2739);
and AND3 (N7024, N7004, N236, N5595);
not NOT1 (N7025, N7019);
xor XOR2 (N7026, N7011, N5347);
not NOT1 (N7027, N7024);
buf BUF1 (N7028, N7014);
nor NOR4 (N7029, N7023, N2396, N187, N5511);
not NOT1 (N7030, N7029);
and AND3 (N7031, N7022, N1847, N1109);
xor XOR2 (N7032, N7030, N6186);
xor XOR2 (N7033, N7026, N1418);
nor NOR2 (N7034, N7031, N6846);
or OR2 (N7035, N7020, N4740);
not NOT1 (N7036, N7028);
or OR3 (N7037, N7034, N3509, N5650);
xor XOR2 (N7038, N7035, N2412);
or OR4 (N7039, N7037, N5947, N4584, N3497);
nand NAND3 (N7040, N7009, N3768, N4395);
nor NOR2 (N7041, N7038, N5809);
or OR3 (N7042, N7032, N795, N5075);
nand NAND2 (N7043, N7039, N30);
or OR2 (N7044, N7040, N6002);
xor XOR2 (N7045, N7027, N3843);
nor NOR2 (N7046, N7041, N4121);
xor XOR2 (N7047, N7036, N6389);
xor XOR2 (N7048, N7045, N4066);
nor NOR3 (N7049, N7025, N3930, N6941);
or OR3 (N7050, N7046, N480, N7027);
buf BUF1 (N7051, N7018);
or OR4 (N7052, N7042, N3719, N6696, N6065);
xor XOR2 (N7053, N7033, N3409);
not NOT1 (N7054, N7050);
xor XOR2 (N7055, N7047, N6461);
not NOT1 (N7056, N7055);
nand NAND3 (N7057, N7048, N6641, N153);
or OR4 (N7058, N7052, N4227, N4427, N2222);
not NOT1 (N7059, N7053);
nand NAND4 (N7060, N7015, N1574, N6106, N3444);
nor NOR3 (N7061, N7057, N3128, N6172);
nor NOR3 (N7062, N7051, N2126, N6398);
nor NOR4 (N7063, N7049, N1888, N6254, N634);
not NOT1 (N7064, N7056);
or OR3 (N7065, N7061, N1803, N5901);
nor NOR2 (N7066, N7063, N442);
nor NOR4 (N7067, N7066, N3091, N5602, N275);
or OR2 (N7068, N7064, N4008);
nor NOR2 (N7069, N7058, N6196);
nor NOR4 (N7070, N7043, N1248, N351, N1854);
xor XOR2 (N7071, N7067, N852);
or OR4 (N7072, N7068, N5928, N1909, N4808);
xor XOR2 (N7073, N7072, N2631);
nand NAND2 (N7074, N7060, N2467);
nor NOR2 (N7075, N7062, N1615);
xor XOR2 (N7076, N7074, N6244);
xor XOR2 (N7077, N7065, N4824);
and AND4 (N7078, N7054, N1344, N6007, N2563);
buf BUF1 (N7079, N7044);
nand NAND4 (N7080, N7078, N3719, N4210, N4248);
and AND4 (N7081, N7069, N6739, N4357, N2093);
xor XOR2 (N7082, N7059, N5856);
buf BUF1 (N7083, N7070);
not NOT1 (N7084, N7075);
and AND2 (N7085, N7084, N5631);
not NOT1 (N7086, N7082);
and AND2 (N7087, N7079, N58);
buf BUF1 (N7088, N7076);
nand NAND3 (N7089, N7071, N4590, N4828);
nand NAND4 (N7090, N7080, N6455, N5405, N1525);
xor XOR2 (N7091, N7073, N1725);
nand NAND2 (N7092, N7088, N1553);
or OR4 (N7093, N7092, N1333, N6151, N5016);
or OR4 (N7094, N7085, N5904, N3337, N3335);
and AND2 (N7095, N7083, N1274);
nor NOR3 (N7096, N7081, N1915, N2826);
or OR2 (N7097, N7090, N4383);
not NOT1 (N7098, N7086);
buf BUF1 (N7099, N7093);
or OR4 (N7100, N7098, N3620, N3848, N4014);
xor XOR2 (N7101, N7091, N1021);
nor NOR3 (N7102, N7101, N4434, N2825);
and AND3 (N7103, N7095, N5943, N5434);
xor XOR2 (N7104, N7100, N153);
and AND3 (N7105, N7104, N1851, N97);
or OR4 (N7106, N7103, N519, N1682, N6631);
not NOT1 (N7107, N7105);
xor XOR2 (N7108, N7099, N931);
nand NAND4 (N7109, N7106, N3534, N549, N6713);
buf BUF1 (N7110, N7109);
or OR2 (N7111, N7096, N4146);
not NOT1 (N7112, N7077);
xor XOR2 (N7113, N7110, N6187);
nor NOR4 (N7114, N7094, N5738, N6366, N3629);
and AND4 (N7115, N7111, N1094, N1258, N2793);
nor NOR3 (N7116, N7107, N4585, N1637);
buf BUF1 (N7117, N7087);
nand NAND2 (N7118, N7108, N2861);
or OR4 (N7119, N7114, N252, N6601, N4682);
nor NOR2 (N7120, N7097, N3796);
or OR4 (N7121, N7117, N58, N5733, N2290);
nor NOR2 (N7122, N7112, N1690);
nor NOR3 (N7123, N7122, N3334, N5779);
and AND3 (N7124, N7113, N5926, N760);
or OR4 (N7125, N7123, N3828, N1977, N4035);
or OR3 (N7126, N7116, N5766, N5049);
not NOT1 (N7127, N7089);
nand NAND4 (N7128, N7119, N3121, N5041, N1460);
and AND4 (N7129, N7121, N2496, N1654, N902);
nor NOR4 (N7130, N7128, N1338, N4096, N4659);
nand NAND3 (N7131, N7127, N4576, N2990);
buf BUF1 (N7132, N7129);
xor XOR2 (N7133, N7132, N5217);
xor XOR2 (N7134, N7115, N5348);
buf BUF1 (N7135, N7124);
buf BUF1 (N7136, N7102);
and AND3 (N7137, N7133, N381, N5741);
and AND3 (N7138, N7118, N6696, N5842);
nor NOR3 (N7139, N7131, N6891, N2751);
and AND3 (N7140, N7136, N5168, N1429);
and AND2 (N7141, N7140, N578);
and AND2 (N7142, N7125, N2049);
not NOT1 (N7143, N7135);
nand NAND4 (N7144, N7134, N3935, N1125, N3962);
nor NOR2 (N7145, N7126, N5581);
buf BUF1 (N7146, N7145);
or OR4 (N7147, N7146, N2543, N44, N5157);
nand NAND4 (N7148, N7144, N2235, N4443, N2165);
or OR3 (N7149, N7143, N3275, N2887);
not NOT1 (N7150, N7147);
xor XOR2 (N7151, N7141, N3910);
nor NOR4 (N7152, N7130, N608, N5334, N4770);
and AND2 (N7153, N7138, N3231);
not NOT1 (N7154, N7153);
nand NAND2 (N7155, N7149, N461);
buf BUF1 (N7156, N7151);
not NOT1 (N7157, N7154);
xor XOR2 (N7158, N7150, N1572);
not NOT1 (N7159, N7158);
not NOT1 (N7160, N7148);
nand NAND4 (N7161, N7157, N4154, N1804, N5922);
not NOT1 (N7162, N7142);
and AND4 (N7163, N7139, N2765, N5187, N313);
xor XOR2 (N7164, N7137, N3473);
nand NAND3 (N7165, N7162, N3452, N592);
nand NAND3 (N7166, N7164, N2627, N1953);
xor XOR2 (N7167, N7160, N6679);
nand NAND3 (N7168, N7166, N6740, N2358);
nor NOR4 (N7169, N7165, N6432, N6938, N1744);
buf BUF1 (N7170, N7152);
buf BUF1 (N7171, N7169);
not NOT1 (N7172, N7163);
and AND3 (N7173, N7159, N4981, N3920);
nor NOR2 (N7174, N7168, N7121);
not NOT1 (N7175, N7173);
buf BUF1 (N7176, N7156);
not NOT1 (N7177, N7155);
xor XOR2 (N7178, N7172, N4093);
nand NAND2 (N7179, N7167, N5931);
or OR2 (N7180, N7120, N3324);
nand NAND2 (N7181, N7177, N6815);
not NOT1 (N7182, N7170);
nor NOR3 (N7183, N7161, N322, N5160);
and AND2 (N7184, N7183, N4694);
nand NAND3 (N7185, N7174, N5546, N2734);
not NOT1 (N7186, N7175);
nand NAND4 (N7187, N7178, N4487, N1162, N3407);
or OR4 (N7188, N7179, N3152, N5448, N5514);
or OR4 (N7189, N7188, N5437, N5655, N121);
xor XOR2 (N7190, N7180, N2113);
not NOT1 (N7191, N7176);
xor XOR2 (N7192, N7171, N6989);
nor NOR2 (N7193, N7185, N2337);
or OR4 (N7194, N7184, N3779, N5884, N3969);
not NOT1 (N7195, N7191);
or OR4 (N7196, N7190, N4159, N249, N6078);
nand NAND3 (N7197, N7196, N6066, N311);
nand NAND4 (N7198, N7194, N40, N1072, N2000);
and AND4 (N7199, N7195, N2313, N6531, N6266);
or OR2 (N7200, N7186, N4700);
buf BUF1 (N7201, N7200);
buf BUF1 (N7202, N7187);
not NOT1 (N7203, N7198);
not NOT1 (N7204, N7199);
and AND4 (N7205, N7193, N1135, N2864, N6104);
nand NAND4 (N7206, N7192, N1578, N6804, N5629);
buf BUF1 (N7207, N7206);
buf BUF1 (N7208, N7205);
xor XOR2 (N7209, N7201, N3477);
nand NAND4 (N7210, N7189, N1057, N2244, N904);
or OR4 (N7211, N7202, N5513, N3202, N1223);
buf BUF1 (N7212, N7182);
nand NAND3 (N7213, N7212, N682, N2513);
nand NAND4 (N7214, N7204, N2633, N5982, N4703);
not NOT1 (N7215, N7210);
nand NAND4 (N7216, N7215, N5720, N5541, N2469);
or OR2 (N7217, N7214, N6896);
or OR3 (N7218, N7209, N2215, N3950);
xor XOR2 (N7219, N7207, N1236);
buf BUF1 (N7220, N7219);
nor NOR2 (N7221, N7220, N5963);
not NOT1 (N7222, N7197);
nor NOR4 (N7223, N7221, N5739, N6627, N1688);
nand NAND2 (N7224, N7216, N6779);
or OR4 (N7225, N7208, N3509, N4287, N6141);
and AND4 (N7226, N7222, N4591, N417, N3484);
buf BUF1 (N7227, N7213);
nand NAND2 (N7228, N7224, N5233);
not NOT1 (N7229, N7217);
and AND3 (N7230, N7203, N5531, N5953);
buf BUF1 (N7231, N7211);
not NOT1 (N7232, N7223);
xor XOR2 (N7233, N7231, N1077);
not NOT1 (N7234, N7230);
and AND4 (N7235, N7232, N3978, N2398, N5245);
and AND3 (N7236, N7226, N6672, N4726);
not NOT1 (N7237, N7235);
or OR2 (N7238, N7218, N693);
xor XOR2 (N7239, N7228, N5050);
not NOT1 (N7240, N7233);
and AND4 (N7241, N7234, N6394, N2174, N6486);
buf BUF1 (N7242, N7225);
buf BUF1 (N7243, N7242);
not NOT1 (N7244, N7239);
and AND2 (N7245, N7238, N1846);
nand NAND4 (N7246, N7244, N5403, N2667, N5583);
buf BUF1 (N7247, N7241);
xor XOR2 (N7248, N7243, N6425);
nand NAND3 (N7249, N7181, N6916, N4683);
not NOT1 (N7250, N7237);
nor NOR3 (N7251, N7246, N6749, N4169);
xor XOR2 (N7252, N7236, N6001);
and AND4 (N7253, N7249, N6256, N4550, N2261);
nor NOR4 (N7254, N7253, N6604, N2745, N2115);
or OR3 (N7255, N7254, N1058, N2940);
or OR4 (N7256, N7227, N1369, N4598, N2720);
and AND2 (N7257, N7245, N5427);
nand NAND3 (N7258, N7229, N3196, N5890);
buf BUF1 (N7259, N7255);
or OR4 (N7260, N7252, N3239, N4277, N416);
nor NOR2 (N7261, N7248, N5228);
buf BUF1 (N7262, N7258);
nor NOR3 (N7263, N7250, N1917, N1501);
nor NOR4 (N7264, N7257, N2445, N3889, N801);
or OR3 (N7265, N7259, N1334, N3984);
nor NOR2 (N7266, N7240, N36);
and AND3 (N7267, N7262, N4210, N4845);
buf BUF1 (N7268, N7256);
xor XOR2 (N7269, N7267, N405);
and AND2 (N7270, N7265, N5164);
and AND3 (N7271, N7251, N7138, N4363);
nor NOR2 (N7272, N7261, N6498);
or OR4 (N7273, N7269, N6959, N305, N156);
buf BUF1 (N7274, N7273);
xor XOR2 (N7275, N7264, N1778);
or OR3 (N7276, N7271, N5127, N6462);
xor XOR2 (N7277, N7274, N2057);
or OR3 (N7278, N7270, N4518, N3940);
nand NAND3 (N7279, N7268, N6594, N2233);
and AND4 (N7280, N7247, N2114, N820, N4689);
or OR2 (N7281, N7280, N2533);
buf BUF1 (N7282, N7279);
buf BUF1 (N7283, N7277);
xor XOR2 (N7284, N7282, N3656);
nor NOR3 (N7285, N7283, N1902, N7163);
not NOT1 (N7286, N7263);
xor XOR2 (N7287, N7284, N1956);
xor XOR2 (N7288, N7272, N4736);
and AND2 (N7289, N7281, N1079);
nor NOR4 (N7290, N7260, N5205, N6833, N5795);
or OR2 (N7291, N7285, N2813);
nor NOR2 (N7292, N7278, N3391);
nand NAND3 (N7293, N7288, N3598, N6439);
not NOT1 (N7294, N7293);
nor NOR3 (N7295, N7266, N5288, N2710);
buf BUF1 (N7296, N7295);
or OR4 (N7297, N7290, N4866, N3759, N918);
xor XOR2 (N7298, N7296, N6950);
buf BUF1 (N7299, N7298);
buf BUF1 (N7300, N7292);
not NOT1 (N7301, N7287);
buf BUF1 (N7302, N7275);
xor XOR2 (N7303, N7291, N2164);
nand NAND3 (N7304, N7276, N6424, N2441);
or OR3 (N7305, N7294, N6737, N5037);
not NOT1 (N7306, N7297);
not NOT1 (N7307, N7299);
nor NOR3 (N7308, N7305, N913, N5676);
xor XOR2 (N7309, N7303, N2109);
not NOT1 (N7310, N7304);
or OR2 (N7311, N7310, N529);
buf BUF1 (N7312, N7308);
xor XOR2 (N7313, N7289, N4609);
not NOT1 (N7314, N7300);
nor NOR2 (N7315, N7312, N1479);
xor XOR2 (N7316, N7307, N449);
not NOT1 (N7317, N7316);
nor NOR4 (N7318, N7314, N2659, N664, N2266);
or OR2 (N7319, N7313, N1879);
xor XOR2 (N7320, N7306, N6215);
buf BUF1 (N7321, N7301);
buf BUF1 (N7322, N7311);
nand NAND2 (N7323, N7286, N6776);
nor NOR3 (N7324, N7321, N1739, N1992);
and AND2 (N7325, N7319, N6122);
and AND3 (N7326, N7320, N1768, N4337);
xor XOR2 (N7327, N7322, N601);
and AND4 (N7328, N7317, N6241, N2369, N2063);
or OR2 (N7329, N7327, N2554);
nor NOR3 (N7330, N7315, N6201, N1778);
nor NOR4 (N7331, N7328, N2559, N1390, N3493);
and AND4 (N7332, N7331, N3097, N2941, N5723);
and AND2 (N7333, N7323, N5753);
xor XOR2 (N7334, N7332, N4051);
xor XOR2 (N7335, N7333, N2988);
buf BUF1 (N7336, N7329);
xor XOR2 (N7337, N7309, N80);
nor NOR2 (N7338, N7326, N6501);
buf BUF1 (N7339, N7335);
not NOT1 (N7340, N7324);
and AND2 (N7341, N7330, N5003);
xor XOR2 (N7342, N7339, N1706);
or OR4 (N7343, N7341, N3645, N3901, N5704);
not NOT1 (N7344, N7338);
buf BUF1 (N7345, N7336);
and AND4 (N7346, N7345, N4219, N1989, N2998);
or OR4 (N7347, N7344, N2629, N5113, N6908);
xor XOR2 (N7348, N7347, N3495);
nor NOR2 (N7349, N7325, N3225);
nand NAND4 (N7350, N7346, N2673, N7275, N2705);
buf BUF1 (N7351, N7348);
nand NAND2 (N7352, N7342, N1157);
and AND4 (N7353, N7340, N4854, N2714, N6810);
nand NAND4 (N7354, N7352, N2029, N6128, N1200);
and AND4 (N7355, N7337, N3541, N6002, N1584);
or OR4 (N7356, N7350, N110, N329, N883);
not NOT1 (N7357, N7351);
nor NOR4 (N7358, N7334, N1278, N3568, N34);
xor XOR2 (N7359, N7349, N3194);
not NOT1 (N7360, N7357);
buf BUF1 (N7361, N7354);
buf BUF1 (N7362, N7302);
nor NOR2 (N7363, N7353, N6250);
nor NOR4 (N7364, N7343, N4031, N201, N716);
nand NAND4 (N7365, N7355, N3594, N7251, N5110);
and AND2 (N7366, N7358, N4790);
not NOT1 (N7367, N7363);
xor XOR2 (N7368, N7365, N6477);
and AND3 (N7369, N7360, N3611, N2430);
or OR2 (N7370, N7369, N6341);
nand NAND2 (N7371, N7362, N3014);
buf BUF1 (N7372, N7318);
nand NAND4 (N7373, N7359, N1613, N6803, N6269);
xor XOR2 (N7374, N7356, N2480);
and AND4 (N7375, N7374, N1402, N5317, N4054);
not NOT1 (N7376, N7370);
xor XOR2 (N7377, N7372, N1826);
not NOT1 (N7378, N7373);
xor XOR2 (N7379, N7361, N2007);
not NOT1 (N7380, N7368);
nand NAND2 (N7381, N7376, N7258);
not NOT1 (N7382, N7380);
or OR2 (N7383, N7378, N547);
nor NOR2 (N7384, N7371, N2778);
nand NAND2 (N7385, N7366, N5931);
nor NOR4 (N7386, N7375, N7245, N1383, N6258);
or OR4 (N7387, N7385, N5881, N6173, N7372);
nand NAND3 (N7388, N7381, N3274, N4559);
not NOT1 (N7389, N7377);
not NOT1 (N7390, N7386);
not NOT1 (N7391, N7382);
or OR2 (N7392, N7379, N1833);
and AND3 (N7393, N7384, N4990, N5225);
and AND3 (N7394, N7389, N2854, N2758);
nor NOR2 (N7395, N7392, N7249);
nor NOR3 (N7396, N7395, N3615, N848);
buf BUF1 (N7397, N7394);
not NOT1 (N7398, N7390);
xor XOR2 (N7399, N7388, N6216);
not NOT1 (N7400, N7396);
buf BUF1 (N7401, N7383);
nor NOR4 (N7402, N7401, N3811, N1843, N4564);
not NOT1 (N7403, N7398);
nand NAND2 (N7404, N7364, N28);
and AND4 (N7405, N7403, N2317, N3201, N6029);
or OR4 (N7406, N7404, N2076, N1168, N6158);
nor NOR2 (N7407, N7402, N809);
or OR4 (N7408, N7399, N5023, N288, N6226);
and AND3 (N7409, N7407, N2493, N3677);
not NOT1 (N7410, N7400);
nand NAND4 (N7411, N7387, N2398, N4569, N1946);
not NOT1 (N7412, N7411);
or OR2 (N7413, N7410, N3567);
buf BUF1 (N7414, N7391);
or OR2 (N7415, N7406, N4036);
nor NOR3 (N7416, N7393, N7087, N4481);
nand NAND4 (N7417, N7413, N56, N6688, N7415);
xor XOR2 (N7418, N5747, N6992);
buf BUF1 (N7419, N7405);
xor XOR2 (N7420, N7409, N3422);
nand NAND3 (N7421, N7417, N1904, N6414);
nor NOR3 (N7422, N7419, N3785, N5271);
nand NAND2 (N7423, N7408, N3163);
not NOT1 (N7424, N7423);
nor NOR4 (N7425, N7414, N4768, N5857, N1621);
or OR3 (N7426, N7420, N2883, N1274);
or OR3 (N7427, N7418, N2689, N1224);
nor NOR3 (N7428, N7421, N6539, N2008);
xor XOR2 (N7429, N7412, N4022);
not NOT1 (N7430, N7397);
buf BUF1 (N7431, N7367);
not NOT1 (N7432, N7426);
buf BUF1 (N7433, N7422);
nor NOR4 (N7434, N7416, N2860, N382, N3662);
and AND3 (N7435, N7424, N1650, N5215);
buf BUF1 (N7436, N7431);
or OR3 (N7437, N7428, N4153, N5926);
not NOT1 (N7438, N7435);
nor NOR3 (N7439, N7437, N7199, N1630);
buf BUF1 (N7440, N7430);
or OR3 (N7441, N7433, N6553, N3407);
and AND3 (N7442, N7432, N3289, N108);
nor NOR3 (N7443, N7436, N775, N5022);
xor XOR2 (N7444, N7425, N1394);
not NOT1 (N7445, N7438);
not NOT1 (N7446, N7429);
not NOT1 (N7447, N7434);
xor XOR2 (N7448, N7439, N5177);
nor NOR4 (N7449, N7427, N2743, N4033, N2354);
buf BUF1 (N7450, N7449);
nand NAND4 (N7451, N7442, N3393, N1882, N1474);
not NOT1 (N7452, N7441);
nor NOR4 (N7453, N7451, N6201, N886, N3636);
not NOT1 (N7454, N7443);
not NOT1 (N7455, N7440);
and AND2 (N7456, N7444, N6327);
or OR4 (N7457, N7456, N5106, N6982, N6486);
nor NOR2 (N7458, N7452, N7363);
or OR4 (N7459, N7457, N6712, N1131, N6526);
nand NAND4 (N7460, N7446, N6007, N6333, N21);
nand NAND2 (N7461, N7450, N6007);
and AND3 (N7462, N7455, N662, N4963);
nand NAND4 (N7463, N7460, N795, N1033, N3575);
buf BUF1 (N7464, N7462);
and AND4 (N7465, N7453, N1513, N654, N2441);
buf BUF1 (N7466, N7461);
and AND2 (N7467, N7445, N6530);
and AND4 (N7468, N7447, N391, N5148, N4656);
nor NOR4 (N7469, N7464, N6736, N5705, N16);
not NOT1 (N7470, N7459);
nand NAND3 (N7471, N7470, N3698, N6505);
or OR2 (N7472, N7471, N6429);
not NOT1 (N7473, N7465);
not NOT1 (N7474, N7458);
not NOT1 (N7475, N7469);
not NOT1 (N7476, N7466);
nor NOR3 (N7477, N7473, N5692, N4685);
not NOT1 (N7478, N7474);
xor XOR2 (N7479, N7463, N4276);
nand NAND3 (N7480, N7467, N7274, N4407);
nor NOR4 (N7481, N7480, N1485, N609, N1819);
not NOT1 (N7482, N7448);
nor NOR2 (N7483, N7482, N6257);
nand NAND4 (N7484, N7481, N5419, N4735, N5704);
and AND2 (N7485, N7472, N6155);
buf BUF1 (N7486, N7479);
xor XOR2 (N7487, N7475, N2865);
nand NAND3 (N7488, N7485, N4816, N3805);
not NOT1 (N7489, N7486);
and AND4 (N7490, N7488, N2967, N4627, N3317);
nor NOR2 (N7491, N7454, N6075);
nand NAND4 (N7492, N7483, N5884, N3997, N4640);
and AND3 (N7493, N7487, N2619, N3697);
buf BUF1 (N7494, N7478);
xor XOR2 (N7495, N7493, N6778);
and AND2 (N7496, N7477, N3216);
xor XOR2 (N7497, N7494, N4836);
not NOT1 (N7498, N7492);
or OR2 (N7499, N7490, N929);
nor NOR4 (N7500, N7489, N1724, N5619, N5772);
xor XOR2 (N7501, N7476, N2026);
nand NAND3 (N7502, N7499, N2186, N2514);
nor NOR4 (N7503, N7498, N5470, N1212, N5548);
and AND3 (N7504, N7501, N4535, N3299);
or OR4 (N7505, N7495, N4889, N2306, N4584);
not NOT1 (N7506, N7468);
buf BUF1 (N7507, N7504);
or OR4 (N7508, N7506, N6366, N3668, N3391);
not NOT1 (N7509, N7496);
and AND4 (N7510, N7491, N2300, N7060, N243);
and AND3 (N7511, N7484, N4641, N4270);
nor NOR4 (N7512, N7500, N1711, N3229, N4295);
xor XOR2 (N7513, N7505, N5722);
xor XOR2 (N7514, N7502, N6978);
nand NAND3 (N7515, N7511, N4227, N3041);
nor NOR2 (N7516, N7508, N1358);
nand NAND2 (N7517, N7507, N2329);
nor NOR4 (N7518, N7503, N1110, N5355, N4506);
nor NOR3 (N7519, N7516, N240, N2495);
nand NAND4 (N7520, N7509, N100, N5946, N5149);
buf BUF1 (N7521, N7519);
xor XOR2 (N7522, N7510, N3273);
nor NOR3 (N7523, N7522, N5769, N2462);
xor XOR2 (N7524, N7514, N4044);
nand NAND3 (N7525, N7515, N1609, N1377);
or OR3 (N7526, N7524, N3292, N3781);
and AND4 (N7527, N7520, N993, N566, N3795);
nor NOR3 (N7528, N7518, N4004, N2906);
nand NAND3 (N7529, N7525, N2312, N1231);
buf BUF1 (N7530, N7512);
xor XOR2 (N7531, N7528, N6576);
not NOT1 (N7532, N7527);
nand NAND3 (N7533, N7532, N4831, N2145);
nand NAND2 (N7534, N7533, N3523);
nor NOR3 (N7535, N7534, N3176, N2701);
not NOT1 (N7536, N7517);
nand NAND3 (N7537, N7535, N2558, N7438);
xor XOR2 (N7538, N7513, N4079);
buf BUF1 (N7539, N7497);
xor XOR2 (N7540, N7521, N5156);
and AND3 (N7541, N7530, N224, N5326);
nand NAND4 (N7542, N7537, N6407, N386, N5196);
nor NOR2 (N7543, N7542, N6440);
nand NAND2 (N7544, N7539, N5772);
nand NAND2 (N7545, N7536, N2950);
nand NAND4 (N7546, N7540, N3621, N1626, N7018);
nand NAND4 (N7547, N7546, N1340, N1459, N6115);
xor XOR2 (N7548, N7531, N5014);
buf BUF1 (N7549, N7523);
xor XOR2 (N7550, N7549, N1742);
and AND3 (N7551, N7550, N5840, N5139);
nand NAND3 (N7552, N7526, N7127, N4569);
or OR4 (N7553, N7551, N4328, N1710, N5950);
and AND3 (N7554, N7529, N1100, N852);
nor NOR4 (N7555, N7541, N2023, N388, N4930);
not NOT1 (N7556, N7548);
nand NAND2 (N7557, N7556, N992);
nand NAND2 (N7558, N7555, N6475);
not NOT1 (N7559, N7553);
buf BUF1 (N7560, N7558);
and AND4 (N7561, N7559, N4111, N5002, N909);
buf BUF1 (N7562, N7544);
not NOT1 (N7563, N7547);
xor XOR2 (N7564, N7560, N1573);
buf BUF1 (N7565, N7564);
buf BUF1 (N7566, N7563);
and AND2 (N7567, N7554, N4134);
xor XOR2 (N7568, N7561, N4031);
not NOT1 (N7569, N7557);
nand NAND2 (N7570, N7545, N2187);
nand NAND4 (N7571, N7543, N629, N7280, N6412);
or OR3 (N7572, N7562, N1723, N4119);
and AND4 (N7573, N7567, N2384, N2571, N3956);
nor NOR3 (N7574, N7573, N5379, N2065);
not NOT1 (N7575, N7538);
and AND2 (N7576, N7574, N670);
nor NOR4 (N7577, N7576, N6256, N6238, N2590);
buf BUF1 (N7578, N7569);
nor NOR3 (N7579, N7570, N902, N4687);
xor XOR2 (N7580, N7566, N5981);
or OR3 (N7581, N7571, N1098, N4821);
not NOT1 (N7582, N7565);
or OR2 (N7583, N7552, N5332);
nand NAND2 (N7584, N7581, N7300);
not NOT1 (N7585, N7579);
not NOT1 (N7586, N7578);
not NOT1 (N7587, N7586);
nand NAND4 (N7588, N7572, N1587, N5366, N3488);
nand NAND4 (N7589, N7575, N3909, N260, N1423);
xor XOR2 (N7590, N7583, N6685);
nor NOR4 (N7591, N7582, N1053, N3292, N7316);
nor NOR2 (N7592, N7584, N4462);
not NOT1 (N7593, N7591);
xor XOR2 (N7594, N7592, N2248);
and AND3 (N7595, N7589, N6477, N4884);
or OR2 (N7596, N7595, N4348);
nand NAND4 (N7597, N7580, N5124, N133, N1307);
and AND3 (N7598, N7597, N3419, N100);
buf BUF1 (N7599, N7587);
and AND4 (N7600, N7598, N4596, N3019, N160);
or OR3 (N7601, N7593, N2711, N7575);
buf BUF1 (N7602, N7585);
and AND3 (N7603, N7596, N2069, N7324);
and AND2 (N7604, N7599, N6313);
nand NAND2 (N7605, N7600, N6078);
nor NOR2 (N7606, N7568, N5578);
xor XOR2 (N7607, N7577, N1754);
and AND2 (N7608, N7590, N2730);
xor XOR2 (N7609, N7606, N3505);
buf BUF1 (N7610, N7608);
buf BUF1 (N7611, N7610);
not NOT1 (N7612, N7611);
not NOT1 (N7613, N7588);
and AND2 (N7614, N7612, N5943);
and AND2 (N7615, N7605, N245);
xor XOR2 (N7616, N7607, N3497);
nor NOR3 (N7617, N7603, N37, N1773);
buf BUF1 (N7618, N7614);
or OR2 (N7619, N7604, N6346);
and AND4 (N7620, N7615, N4647, N4902, N7543);
not NOT1 (N7621, N7602);
nor NOR3 (N7622, N7617, N5687, N4008);
not NOT1 (N7623, N7601);
nand NAND4 (N7624, N7621, N3381, N6898, N3159);
xor XOR2 (N7625, N7624, N436);
buf BUF1 (N7626, N7620);
nand NAND2 (N7627, N7622, N5129);
nand NAND3 (N7628, N7626, N6988, N6807);
or OR3 (N7629, N7619, N827, N4207);
not NOT1 (N7630, N7594);
and AND3 (N7631, N7609, N3248, N4235);
nand NAND3 (N7632, N7618, N3470, N7102);
nor NOR3 (N7633, N7623, N1477, N5812);
and AND2 (N7634, N7625, N519);
nand NAND3 (N7635, N7630, N6411, N1598);
not NOT1 (N7636, N7616);
or OR4 (N7637, N7631, N5194, N2432, N5648);
nor NOR2 (N7638, N7635, N3828);
nor NOR4 (N7639, N7613, N1649, N1257, N4970);
nand NAND3 (N7640, N7628, N2972, N1818);
xor XOR2 (N7641, N7633, N1674);
buf BUF1 (N7642, N7636);
or OR4 (N7643, N7629, N3452, N7620, N6395);
buf BUF1 (N7644, N7643);
or OR3 (N7645, N7638, N2592, N3156);
xor XOR2 (N7646, N7639, N4747);
buf BUF1 (N7647, N7645);
xor XOR2 (N7648, N7627, N3604);
nor NOR4 (N7649, N7637, N131, N4395, N6856);
and AND4 (N7650, N7634, N7256, N3016, N2588);
nor NOR2 (N7651, N7644, N7271);
and AND3 (N7652, N7642, N5123, N3882);
nor NOR3 (N7653, N7648, N6734, N1672);
not NOT1 (N7654, N7650);
buf BUF1 (N7655, N7651);
or OR3 (N7656, N7632, N4342, N3214);
nor NOR4 (N7657, N7653, N5830, N4373, N7474);
buf BUF1 (N7658, N7656);
buf BUF1 (N7659, N7640);
not NOT1 (N7660, N7641);
xor XOR2 (N7661, N7654, N7034);
nor NOR3 (N7662, N7659, N6593, N6985);
and AND4 (N7663, N7652, N2517, N6872, N1088);
nor NOR2 (N7664, N7660, N3131);
xor XOR2 (N7665, N7655, N4087);
nor NOR3 (N7666, N7661, N956, N6763);
nor NOR2 (N7667, N7666, N6433);
nand NAND2 (N7668, N7647, N3577);
or OR3 (N7669, N7663, N3210, N4553);
nor NOR2 (N7670, N7667, N2048);
or OR4 (N7671, N7657, N3470, N2716, N3688);
not NOT1 (N7672, N7668);
not NOT1 (N7673, N7669);
xor XOR2 (N7674, N7658, N7021);
buf BUF1 (N7675, N7646);
nand NAND2 (N7676, N7665, N3194);
nand NAND4 (N7677, N7672, N4709, N2656, N1591);
xor XOR2 (N7678, N7673, N6426);
or OR3 (N7679, N7677, N3565, N2645);
nor NOR2 (N7680, N7662, N4436);
nor NOR3 (N7681, N7649, N2623, N3998);
and AND4 (N7682, N7678, N874, N408, N7096);
buf BUF1 (N7683, N7680);
and AND3 (N7684, N7675, N7149, N208);
and AND4 (N7685, N7670, N6258, N3792, N7232);
xor XOR2 (N7686, N7681, N3635);
or OR3 (N7687, N7679, N3187, N6398);
or OR2 (N7688, N7676, N799);
nor NOR4 (N7689, N7687, N7275, N4095, N2031);
xor XOR2 (N7690, N7686, N3778);
xor XOR2 (N7691, N7674, N2516);
and AND2 (N7692, N7684, N847);
xor XOR2 (N7693, N7690, N4158);
and AND4 (N7694, N7691, N5421, N6327, N3421);
xor XOR2 (N7695, N7692, N5694);
buf BUF1 (N7696, N7693);
and AND3 (N7697, N7682, N1972, N543);
and AND2 (N7698, N7685, N725);
not NOT1 (N7699, N7671);
nor NOR2 (N7700, N7696, N3507);
buf BUF1 (N7701, N7700);
or OR4 (N7702, N7664, N6426, N937, N4539);
and AND3 (N7703, N7688, N7333, N5291);
nand NAND3 (N7704, N7689, N7067, N748);
nor NOR4 (N7705, N7701, N2145, N6868, N291);
nand NAND4 (N7706, N7695, N2231, N284, N7648);
and AND4 (N7707, N7704, N3368, N2413, N6980);
or OR2 (N7708, N7707, N6494);
and AND2 (N7709, N7703, N2606);
xor XOR2 (N7710, N7683, N1113);
nor NOR2 (N7711, N7709, N1815);
buf BUF1 (N7712, N7699);
or OR4 (N7713, N7698, N2156, N7629, N3908);
buf BUF1 (N7714, N7697);
and AND3 (N7715, N7708, N1867, N4828);
or OR2 (N7716, N7711, N1154);
nor NOR2 (N7717, N7716, N772);
and AND3 (N7718, N7710, N3251, N1311);
xor XOR2 (N7719, N7712, N2034);
or OR2 (N7720, N7705, N5638);
and AND4 (N7721, N7694, N3342, N1947, N6551);
or OR2 (N7722, N7713, N4982);
nor NOR4 (N7723, N7706, N984, N4401, N2576);
xor XOR2 (N7724, N7715, N6319);
xor XOR2 (N7725, N7719, N5221);
or OR4 (N7726, N7723, N348, N5196, N824);
nand NAND2 (N7727, N7722, N1207);
buf BUF1 (N7728, N7717);
nor NOR3 (N7729, N7724, N6593, N4740);
buf BUF1 (N7730, N7725);
or OR3 (N7731, N7714, N350, N2615);
nor NOR3 (N7732, N7730, N5773, N7709);
nand NAND4 (N7733, N7720, N5125, N4899, N2042);
not NOT1 (N7734, N7702);
not NOT1 (N7735, N7726);
or OR2 (N7736, N7734, N4325);
or OR4 (N7737, N7733, N7052, N2246, N1517);
buf BUF1 (N7738, N7731);
or OR4 (N7739, N7729, N2980, N3935, N4027);
nand NAND3 (N7740, N7735, N4173, N3116);
or OR2 (N7741, N7738, N3286);
or OR4 (N7742, N7741, N2830, N2970, N2049);
not NOT1 (N7743, N7736);
xor XOR2 (N7744, N7737, N2826);
nor NOR4 (N7745, N7743, N3553, N3427, N4293);
buf BUF1 (N7746, N7732);
or OR2 (N7747, N7727, N3652);
nand NAND3 (N7748, N7718, N5766, N5042);
nor NOR4 (N7749, N7746, N1525, N1709, N6632);
or OR3 (N7750, N7744, N5870, N440);
buf BUF1 (N7751, N7747);
nand NAND2 (N7752, N7751, N6830);
and AND3 (N7753, N7740, N3313, N6824);
xor XOR2 (N7754, N7748, N6965);
xor XOR2 (N7755, N7721, N6477);
or OR2 (N7756, N7742, N1113);
or OR2 (N7757, N7728, N6508);
xor XOR2 (N7758, N7757, N2147);
and AND3 (N7759, N7745, N3358, N6564);
not NOT1 (N7760, N7758);
nor NOR4 (N7761, N7754, N2083, N5677, N229);
not NOT1 (N7762, N7753);
xor XOR2 (N7763, N7759, N2647);
or OR4 (N7764, N7763, N1554, N2552, N1770);
and AND2 (N7765, N7756, N6177);
nor NOR2 (N7766, N7755, N2118);
or OR2 (N7767, N7749, N2399);
nand NAND3 (N7768, N7765, N610, N5132);
not NOT1 (N7769, N7766);
and AND2 (N7770, N7739, N3692);
xor XOR2 (N7771, N7764, N5608);
buf BUF1 (N7772, N7762);
nand NAND3 (N7773, N7760, N4138, N3551);
nor NOR3 (N7774, N7769, N4437, N2822);
not NOT1 (N7775, N7772);
nor NOR3 (N7776, N7761, N4337, N6774);
or OR4 (N7777, N7774, N6372, N2694, N6768);
or OR4 (N7778, N7775, N2448, N815, N6780);
and AND2 (N7779, N7777, N3376);
and AND2 (N7780, N7752, N5072);
and AND2 (N7781, N7771, N3384);
and AND3 (N7782, N7750, N7329, N7071);
buf BUF1 (N7783, N7778);
or OR4 (N7784, N7780, N802, N6991, N6161);
and AND3 (N7785, N7783, N7275, N5367);
nor NOR3 (N7786, N7782, N3858, N797);
not NOT1 (N7787, N7785);
xor XOR2 (N7788, N7786, N5697);
buf BUF1 (N7789, N7779);
nor NOR3 (N7790, N7781, N2877, N671);
nor NOR4 (N7791, N7789, N5523, N3750, N4371);
not NOT1 (N7792, N7770);
or OR2 (N7793, N7767, N1273);
not NOT1 (N7794, N7776);
buf BUF1 (N7795, N7788);
or OR4 (N7796, N7787, N5550, N1224, N3991);
or OR4 (N7797, N7794, N7108, N5174, N5205);
xor XOR2 (N7798, N7792, N4990);
nor NOR3 (N7799, N7791, N4957, N5875);
nand NAND2 (N7800, N7773, N7728);
or OR4 (N7801, N7796, N5324, N6445, N690);
or OR3 (N7802, N7801, N1996, N6628);
nand NAND4 (N7803, N7784, N5396, N4891, N6872);
buf BUF1 (N7804, N7795);
not NOT1 (N7805, N7802);
and AND3 (N7806, N7804, N1588, N7253);
xor XOR2 (N7807, N7793, N1180);
or OR3 (N7808, N7768, N4531, N5479);
and AND2 (N7809, N7807, N3204);
nor NOR2 (N7810, N7798, N25);
nand NAND3 (N7811, N7810, N517, N76);
buf BUF1 (N7812, N7811);
buf BUF1 (N7813, N7803);
or OR3 (N7814, N7790, N3220, N1321);
xor XOR2 (N7815, N7808, N2681);
not NOT1 (N7816, N7812);
xor XOR2 (N7817, N7806, N2908);
nand NAND4 (N7818, N7809, N5124, N3148, N5759);
or OR3 (N7819, N7815, N7394, N5834);
nor NOR4 (N7820, N7816, N3774, N2507, N3481);
xor XOR2 (N7821, N7814, N1046);
not NOT1 (N7822, N7797);
nand NAND4 (N7823, N7821, N1601, N3975, N1545);
nor NOR4 (N7824, N7818, N5714, N686, N2304);
or OR2 (N7825, N7800, N3374);
nor NOR4 (N7826, N7823, N247, N591, N2802);
not NOT1 (N7827, N7820);
buf BUF1 (N7828, N7805);
nand NAND2 (N7829, N7824, N2107);
and AND4 (N7830, N7813, N3736, N6791, N4349);
or OR4 (N7831, N7799, N3201, N373, N7775);
and AND3 (N7832, N7829, N665, N4319);
xor XOR2 (N7833, N7832, N2521);
buf BUF1 (N7834, N7825);
nor NOR4 (N7835, N7833, N4770, N2955, N5691);
not NOT1 (N7836, N7827);
buf BUF1 (N7837, N7830);
or OR4 (N7838, N7836, N3639, N5989, N5475);
not NOT1 (N7839, N7817);
buf BUF1 (N7840, N7831);
buf BUF1 (N7841, N7826);
xor XOR2 (N7842, N7837, N1892);
buf BUF1 (N7843, N7839);
or OR4 (N7844, N7828, N4960, N3949, N5176);
and AND2 (N7845, N7842, N5889);
nand NAND2 (N7846, N7834, N2263);
nand NAND3 (N7847, N7838, N3514, N2369);
xor XOR2 (N7848, N7845, N2070);
or OR3 (N7849, N7822, N1622, N7695);
nor NOR3 (N7850, N7848, N6175, N2659);
xor XOR2 (N7851, N7847, N6153);
or OR4 (N7852, N7844, N770, N3217, N3632);
nor NOR4 (N7853, N7849, N3107, N1921, N7599);
nand NAND3 (N7854, N7841, N1685, N5835);
nand NAND2 (N7855, N7843, N2855);
buf BUF1 (N7856, N7846);
nand NAND2 (N7857, N7819, N7400);
not NOT1 (N7858, N7850);
buf BUF1 (N7859, N7840);
nor NOR2 (N7860, N7853, N2690);
not NOT1 (N7861, N7859);
and AND3 (N7862, N7856, N7693, N6078);
nor NOR4 (N7863, N7861, N34, N1324, N6294);
not NOT1 (N7864, N7862);
and AND3 (N7865, N7851, N2040, N6491);
nor NOR3 (N7866, N7865, N2092, N3645);
not NOT1 (N7867, N7860);
nand NAND2 (N7868, N7835, N5216);
not NOT1 (N7869, N7867);
or OR2 (N7870, N7854, N2466);
and AND2 (N7871, N7870, N4856);
and AND4 (N7872, N7858, N6479, N7501, N7078);
or OR4 (N7873, N7869, N3274, N7811, N7780);
xor XOR2 (N7874, N7855, N7257);
nor NOR2 (N7875, N7871, N1932);
or OR4 (N7876, N7873, N2367, N5904, N5627);
and AND4 (N7877, N7874, N7362, N4186, N2594);
nand NAND3 (N7878, N7875, N3816, N6699);
nor NOR3 (N7879, N7857, N5228, N2022);
nand NAND3 (N7880, N7852, N4987, N4898);
and AND2 (N7881, N7866, N3010);
and AND4 (N7882, N7880, N3211, N7603, N1354);
or OR4 (N7883, N7878, N30, N7240, N3105);
buf BUF1 (N7884, N7868);
xor XOR2 (N7885, N7881, N7241);
nand NAND2 (N7886, N7863, N5540);
nor NOR3 (N7887, N7864, N3933, N6116);
buf BUF1 (N7888, N7886);
xor XOR2 (N7889, N7876, N1434);
and AND2 (N7890, N7877, N1083);
and AND4 (N7891, N7890, N5381, N7608, N6679);
buf BUF1 (N7892, N7891);
and AND3 (N7893, N7888, N6363, N4906);
or OR3 (N7894, N7879, N7347, N5945);
nand NAND3 (N7895, N7872, N5091, N7578);
nand NAND2 (N7896, N7885, N5008);
buf BUF1 (N7897, N7893);
nand NAND4 (N7898, N7882, N6766, N1035, N1478);
xor XOR2 (N7899, N7884, N5842);
buf BUF1 (N7900, N7899);
not NOT1 (N7901, N7900);
and AND2 (N7902, N7895, N3924);
buf BUF1 (N7903, N7902);
and AND2 (N7904, N7897, N1072);
not NOT1 (N7905, N7894);
not NOT1 (N7906, N7883);
not NOT1 (N7907, N7896);
not NOT1 (N7908, N7907);
xor XOR2 (N7909, N7887, N6684);
xor XOR2 (N7910, N7906, N96);
buf BUF1 (N7911, N7905);
not NOT1 (N7912, N7898);
not NOT1 (N7913, N7889);
nand NAND2 (N7914, N7901, N709);
nor NOR3 (N7915, N7910, N6600, N5726);
buf BUF1 (N7916, N7914);
or OR3 (N7917, N7913, N4622, N2803);
not NOT1 (N7918, N7911);
xor XOR2 (N7919, N7904, N3495);
or OR2 (N7920, N7919, N2238);
xor XOR2 (N7921, N7916, N1106);
nor NOR3 (N7922, N7915, N270, N2797);
and AND3 (N7923, N7912, N1500, N415);
and AND3 (N7924, N7917, N5490, N5490);
xor XOR2 (N7925, N7923, N2891);
not NOT1 (N7926, N7909);
nand NAND4 (N7927, N7918, N7347, N5638, N6278);
or OR3 (N7928, N7922, N4432, N4489);
xor XOR2 (N7929, N7892, N2185);
and AND4 (N7930, N7908, N6797, N3216, N3638);
or OR3 (N7931, N7920, N4458, N5895);
nor NOR2 (N7932, N7929, N821);
not NOT1 (N7933, N7921);
nand NAND3 (N7934, N7924, N2600, N6);
and AND4 (N7935, N7926, N2356, N5227, N5285);
buf BUF1 (N7936, N7927);
xor XOR2 (N7937, N7925, N2433);
buf BUF1 (N7938, N7930);
and AND2 (N7939, N7938, N5750);
and AND4 (N7940, N7937, N1500, N4117, N3766);
and AND4 (N7941, N7936, N4642, N4848, N447);
xor XOR2 (N7942, N7935, N5817);
buf BUF1 (N7943, N7939);
or OR2 (N7944, N7934, N6269);
nor NOR2 (N7945, N7903, N4466);
nor NOR3 (N7946, N7941, N5752, N3867);
not NOT1 (N7947, N7933);
and AND2 (N7948, N7931, N4472);
nand NAND3 (N7949, N7932, N3418, N4636);
not NOT1 (N7950, N7945);
not NOT1 (N7951, N7942);
xor XOR2 (N7952, N7950, N6702);
and AND4 (N7953, N7949, N474, N5509, N4331);
not NOT1 (N7954, N7940);
nand NAND4 (N7955, N7928, N4062, N1262, N7050);
or OR2 (N7956, N7946, N603);
or OR4 (N7957, N7951, N5908, N1647, N2491);
or OR2 (N7958, N7943, N6760);
nor NOR2 (N7959, N7953, N1447);
nor NOR2 (N7960, N7954, N1523);
not NOT1 (N7961, N7960);
and AND2 (N7962, N7957, N6617);
or OR3 (N7963, N7948, N6709, N4144);
buf BUF1 (N7964, N7962);
or OR4 (N7965, N7944, N500, N1273, N7662);
buf BUF1 (N7966, N7958);
nand NAND4 (N7967, N7952, N3231, N1878, N3142);
nor NOR4 (N7968, N7955, N1622, N3661, N6303);
and AND3 (N7969, N7964, N4761, N6530);
not NOT1 (N7970, N7956);
or OR2 (N7971, N7970, N6306);
and AND4 (N7972, N7961, N1145, N5910, N211);
nand NAND2 (N7973, N7959, N1965);
not NOT1 (N7974, N7968);
or OR3 (N7975, N7947, N108, N4802);
nor NOR3 (N7976, N7963, N2558, N7719);
nand NAND3 (N7977, N7974, N1669, N84);
xor XOR2 (N7978, N7975, N4590);
or OR3 (N7979, N7978, N1893, N3730);
buf BUF1 (N7980, N7979);
or OR3 (N7981, N7972, N2813, N2874);
buf BUF1 (N7982, N7965);
and AND4 (N7983, N7976, N7308, N3627, N3021);
nor NOR3 (N7984, N7983, N66, N6990);
not NOT1 (N7985, N7982);
or OR3 (N7986, N7973, N2015, N2195);
not NOT1 (N7987, N7981);
nand NAND2 (N7988, N7969, N7160);
nor NOR3 (N7989, N7985, N7323, N160);
or OR2 (N7990, N7967, N843);
not NOT1 (N7991, N7986);
nor NOR3 (N7992, N7977, N1650, N4791);
nor NOR4 (N7993, N7992, N5257, N7969, N5750);
or OR3 (N7994, N7984, N5967, N3597);
nand NAND4 (N7995, N7980, N7157, N1075, N863);
not NOT1 (N7996, N7971);
nand NAND3 (N7997, N7993, N7911, N386);
nand NAND4 (N7998, N7988, N2981, N6272, N1555);
not NOT1 (N7999, N7991);
xor XOR2 (N8000, N7987, N1281);
nand NAND2 (N8001, N7990, N7526);
nor NOR4 (N8002, N7999, N920, N415, N7626);
and AND3 (N8003, N8002, N3820, N5728);
nand NAND3 (N8004, N8003, N1598, N3406);
nor NOR4 (N8005, N7989, N1763, N989, N6106);
xor XOR2 (N8006, N8001, N2979);
xor XOR2 (N8007, N8000, N4040);
nand NAND2 (N8008, N7966, N5758);
nand NAND2 (N8009, N7996, N2903);
and AND4 (N8010, N8004, N7432, N5844, N6269);
not NOT1 (N8011, N8006);
not NOT1 (N8012, N8005);
not NOT1 (N8013, N8011);
and AND3 (N8014, N8013, N6756, N4671);
nor NOR2 (N8015, N8007, N2550);
and AND3 (N8016, N8015, N7641, N586);
buf BUF1 (N8017, N8014);
and AND3 (N8018, N8016, N6323, N4180);
and AND4 (N8019, N7995, N573, N2954, N3590);
or OR3 (N8020, N8017, N4429, N3100);
buf BUF1 (N8021, N8018);
not NOT1 (N8022, N8021);
or OR3 (N8023, N8022, N3575, N4881);
and AND3 (N8024, N8008, N2016, N7184);
or OR2 (N8025, N8020, N4764);
not NOT1 (N8026, N8012);
buf BUF1 (N8027, N8024);
not NOT1 (N8028, N7997);
nor NOR3 (N8029, N8023, N3661, N1487);
buf BUF1 (N8030, N8010);
buf BUF1 (N8031, N7994);
nand NAND4 (N8032, N8019, N4984, N6879, N2991);
nand NAND3 (N8033, N8029, N6635, N1570);
buf BUF1 (N8034, N8025);
xor XOR2 (N8035, N8032, N3859);
buf BUF1 (N8036, N8030);
xor XOR2 (N8037, N8026, N4425);
not NOT1 (N8038, N8037);
buf BUF1 (N8039, N8034);
and AND2 (N8040, N7998, N3108);
not NOT1 (N8041, N8038);
nor NOR4 (N8042, N8039, N4725, N5039, N5516);
or OR4 (N8043, N8027, N4299, N5612, N4071);
xor XOR2 (N8044, N8009, N3166);
xor XOR2 (N8045, N8044, N3943);
buf BUF1 (N8046, N8028);
not NOT1 (N8047, N8042);
buf BUF1 (N8048, N8035);
and AND4 (N8049, N8047, N4457, N789, N517);
or OR4 (N8050, N8040, N224, N5133, N2353);
and AND2 (N8051, N8041, N880);
nor NOR3 (N8052, N8048, N7066, N4258);
xor XOR2 (N8053, N8036, N3083);
nor NOR4 (N8054, N8053, N7377, N5359, N5169);
or OR2 (N8055, N8049, N3278);
or OR2 (N8056, N8054, N4423);
buf BUF1 (N8057, N8050);
nor NOR2 (N8058, N8056, N3720);
or OR2 (N8059, N8033, N5671);
and AND3 (N8060, N8045, N593, N6856);
nor NOR3 (N8061, N8057, N5081, N220);
buf BUF1 (N8062, N8060);
nor NOR2 (N8063, N8051, N4197);
xor XOR2 (N8064, N8031, N7999);
not NOT1 (N8065, N8064);
xor XOR2 (N8066, N8055, N7292);
nor NOR4 (N8067, N8062, N5914, N6665, N7732);
buf BUF1 (N8068, N8058);
buf BUF1 (N8069, N8046);
buf BUF1 (N8070, N8063);
and AND4 (N8071, N8043, N3251, N466, N2187);
and AND2 (N8072, N8061, N6703);
nor NOR4 (N8073, N8070, N3757, N6927, N5620);
or OR4 (N8074, N8068, N7109, N2506, N7632);
nand NAND3 (N8075, N8065, N1800, N3345);
nand NAND3 (N8076, N8072, N7402, N7491);
or OR2 (N8077, N8074, N5563);
or OR2 (N8078, N8077, N5518);
nand NAND4 (N8079, N8052, N5100, N6646, N5907);
and AND4 (N8080, N8066, N7136, N7588, N7260);
and AND3 (N8081, N8075, N4154, N7092);
not NOT1 (N8082, N8073);
and AND4 (N8083, N8059, N4728, N1525, N6740);
nand NAND2 (N8084, N8069, N178);
and AND3 (N8085, N8079, N2438, N6810);
buf BUF1 (N8086, N8084);
or OR3 (N8087, N8080, N3346, N4726);
nor NOR3 (N8088, N8086, N5086, N4027);
buf BUF1 (N8089, N8088);
xor XOR2 (N8090, N8067, N4694);
xor XOR2 (N8091, N8089, N4051);
or OR3 (N8092, N8076, N4408, N1734);
xor XOR2 (N8093, N8087, N7061);
nor NOR3 (N8094, N8078, N375, N5701);
not NOT1 (N8095, N8090);
xor XOR2 (N8096, N8091, N639);
nand NAND4 (N8097, N8071, N2487, N2331, N550);
or OR4 (N8098, N8081, N6901, N5347, N6045);
or OR4 (N8099, N8085, N2558, N6855, N7627);
nand NAND4 (N8100, N8082, N2229, N6964, N7125);
not NOT1 (N8101, N8097);
not NOT1 (N8102, N8101);
and AND4 (N8103, N8100, N2260, N3611, N2929);
nand NAND4 (N8104, N8096, N2577, N4211, N2058);
nor NOR4 (N8105, N8092, N4548, N5280, N586);
and AND4 (N8106, N8093, N7498, N5044, N6518);
buf BUF1 (N8107, N8103);
and AND4 (N8108, N8104, N631, N5125, N7368);
nor NOR3 (N8109, N8094, N3384, N7768);
buf BUF1 (N8110, N8102);
nand NAND3 (N8111, N8095, N8071, N4776);
and AND2 (N8112, N8106, N5306);
buf BUF1 (N8113, N8111);
not NOT1 (N8114, N8113);
and AND3 (N8115, N8107, N3964, N7476);
nor NOR2 (N8116, N8099, N7793);
nand NAND4 (N8117, N8116, N4502, N245, N3168);
or OR2 (N8118, N8105, N3587);
buf BUF1 (N8119, N8117);
xor XOR2 (N8120, N8118, N4940);
xor XOR2 (N8121, N8083, N3482);
not NOT1 (N8122, N8119);
or OR3 (N8123, N8108, N1948, N5299);
not NOT1 (N8124, N8121);
or OR3 (N8125, N8109, N1082, N2002);
or OR2 (N8126, N8110, N5991);
nand NAND3 (N8127, N8125, N7580, N5781);
or OR3 (N8128, N8115, N7752, N7926);
xor XOR2 (N8129, N8128, N2497);
or OR4 (N8130, N8126, N3236, N4990, N2823);
xor XOR2 (N8131, N8124, N2536);
or OR3 (N8132, N8122, N5358, N6302);
buf BUF1 (N8133, N8112);
and AND3 (N8134, N8132, N7767, N3943);
nand NAND4 (N8135, N8129, N407, N2322, N8100);
buf BUF1 (N8136, N8114);
xor XOR2 (N8137, N8131, N799);
not NOT1 (N8138, N8120);
xor XOR2 (N8139, N8130, N3134);
nor NOR2 (N8140, N8138, N828);
buf BUF1 (N8141, N8140);
and AND2 (N8142, N8123, N4178);
xor XOR2 (N8143, N8135, N4485);
nand NAND3 (N8144, N8127, N2561, N836);
nor NOR2 (N8145, N8143, N6803);
buf BUF1 (N8146, N8136);
xor XOR2 (N8147, N8146, N7379);
buf BUF1 (N8148, N8145);
nand NAND3 (N8149, N8098, N5374, N3251);
xor XOR2 (N8150, N8134, N2306);
nor NOR4 (N8151, N8133, N5337, N8134, N6209);
xor XOR2 (N8152, N8149, N6945);
or OR3 (N8153, N8139, N6668, N2204);
nand NAND3 (N8154, N8147, N1990, N8049);
xor XOR2 (N8155, N8150, N2467);
or OR4 (N8156, N8152, N2114, N5305, N746);
nand NAND3 (N8157, N8148, N4036, N7797);
nor NOR3 (N8158, N8155, N4177, N3661);
nor NOR4 (N8159, N8137, N553, N5708, N7026);
nor NOR3 (N8160, N8159, N5746, N3150);
not NOT1 (N8161, N8144);
nand NAND3 (N8162, N8161, N2742, N6588);
xor XOR2 (N8163, N8157, N7089);
not NOT1 (N8164, N8142);
and AND3 (N8165, N8151, N3677, N6230);
xor XOR2 (N8166, N8141, N6604);
not NOT1 (N8167, N8164);
buf BUF1 (N8168, N8154);
nand NAND3 (N8169, N8163, N1462, N4654);
buf BUF1 (N8170, N8167);
and AND2 (N8171, N8170, N1768);
not NOT1 (N8172, N8165);
buf BUF1 (N8173, N8158);
buf BUF1 (N8174, N8171);
xor XOR2 (N8175, N8168, N7751);
nand NAND2 (N8176, N8160, N1299);
nand NAND2 (N8177, N8153, N7769);
and AND4 (N8178, N8175, N5100, N7276, N1038);
or OR3 (N8179, N8178, N6579, N8110);
buf BUF1 (N8180, N8172);
nand NAND3 (N8181, N8166, N7654, N3018);
and AND3 (N8182, N8174, N1591, N7496);
nor NOR3 (N8183, N8169, N1914, N5615);
or OR3 (N8184, N8156, N2732, N4155);
and AND4 (N8185, N8183, N5177, N7421, N6627);
nand NAND4 (N8186, N8182, N1894, N3950, N1101);
not NOT1 (N8187, N8179);
buf BUF1 (N8188, N8184);
and AND2 (N8189, N8180, N736);
buf BUF1 (N8190, N8189);
and AND3 (N8191, N8177, N7324, N2949);
and AND3 (N8192, N8176, N2438, N2073);
nand NAND4 (N8193, N8187, N29, N4915, N3831);
buf BUF1 (N8194, N8193);
not NOT1 (N8195, N8186);
nor NOR2 (N8196, N8195, N7406);
xor XOR2 (N8197, N8190, N5808);
or OR2 (N8198, N8194, N2991);
nand NAND3 (N8199, N8181, N6247, N6549);
and AND3 (N8200, N8197, N1270, N6823);
nor NOR4 (N8201, N8185, N4477, N7909, N4382);
and AND3 (N8202, N8192, N1094, N1303);
buf BUF1 (N8203, N8173);
or OR4 (N8204, N8203, N1952, N2113, N6327);
or OR2 (N8205, N8199, N6874);
nor NOR4 (N8206, N8191, N6073, N258, N8005);
or OR4 (N8207, N8204, N3608, N4295, N8192);
xor XOR2 (N8208, N8205, N8021);
nand NAND4 (N8209, N8207, N2859, N5252, N6541);
and AND4 (N8210, N8196, N6628, N3443, N2276);
and AND2 (N8211, N8162, N3996);
nor NOR4 (N8212, N8209, N7961, N1036, N3588);
buf BUF1 (N8213, N8188);
buf BUF1 (N8214, N8211);
nand NAND4 (N8215, N8200, N5042, N5645, N2200);
nand NAND3 (N8216, N8214, N3911, N2135);
and AND4 (N8217, N8198, N3751, N4115, N937);
nor NOR2 (N8218, N8201, N3137);
and AND4 (N8219, N8208, N5766, N3821, N7513);
not NOT1 (N8220, N8218);
or OR2 (N8221, N8213, N6139);
buf BUF1 (N8222, N8206);
xor XOR2 (N8223, N8222, N2907);
nor NOR2 (N8224, N8217, N5575);
nor NOR2 (N8225, N8223, N2655);
buf BUF1 (N8226, N8216);
buf BUF1 (N8227, N8215);
nor NOR3 (N8228, N8227, N4713, N5270);
nor NOR4 (N8229, N8220, N1711, N2075, N4734);
nand NAND3 (N8230, N8229, N5254, N4446);
nand NAND3 (N8231, N8226, N854, N5896);
nor NOR3 (N8232, N8221, N1040, N6721);
buf BUF1 (N8233, N8202);
buf BUF1 (N8234, N8228);
or OR4 (N8235, N8225, N1288, N4466, N5800);
and AND4 (N8236, N8231, N134, N3217, N2916);
nor NOR3 (N8237, N8235, N1151, N7696);
nand NAND4 (N8238, N8224, N8077, N6971, N1521);
nor NOR3 (N8239, N8238, N4801, N5496);
xor XOR2 (N8240, N8210, N7392);
and AND4 (N8241, N8212, N4609, N593, N7514);
nor NOR2 (N8242, N8233, N2078);
buf BUF1 (N8243, N8234);
and AND4 (N8244, N8240, N4010, N4936, N4637);
not NOT1 (N8245, N8239);
xor XOR2 (N8246, N8230, N28);
nor NOR4 (N8247, N8245, N7729, N2567, N3123);
nor NOR3 (N8248, N8237, N4934, N1823);
nand NAND3 (N8249, N8243, N1675, N6305);
nand NAND3 (N8250, N8242, N2737, N5610);
nor NOR4 (N8251, N8248, N1936, N7533, N2922);
nand NAND3 (N8252, N8249, N6212, N8207);
or OR2 (N8253, N8251, N542);
not NOT1 (N8254, N8253);
nor NOR4 (N8255, N8219, N2579, N5938, N2611);
buf BUF1 (N8256, N8244);
and AND3 (N8257, N8241, N1580, N5967);
nor NOR2 (N8258, N8247, N7567);
nand NAND3 (N8259, N8257, N3193, N4699);
nand NAND2 (N8260, N8255, N5570);
nand NAND2 (N8261, N8236, N6224);
buf BUF1 (N8262, N8252);
not NOT1 (N8263, N8260);
nor NOR4 (N8264, N8262, N479, N5602, N3518);
or OR4 (N8265, N8232, N2846, N5751, N2751);
and AND3 (N8266, N8250, N8228, N5376);
not NOT1 (N8267, N8258);
and AND4 (N8268, N8266, N2156, N2535, N265);
and AND4 (N8269, N8254, N6860, N2057, N3371);
nand NAND3 (N8270, N8264, N6315, N8244);
nand NAND2 (N8271, N8256, N5182);
xor XOR2 (N8272, N8246, N6966);
buf BUF1 (N8273, N8263);
and AND2 (N8274, N8269, N1384);
buf BUF1 (N8275, N8261);
nor NOR3 (N8276, N8267, N8134, N7703);
xor XOR2 (N8277, N8274, N6681);
nand NAND3 (N8278, N8273, N6072, N3522);
nor NOR3 (N8279, N8270, N359, N2655);
buf BUF1 (N8280, N8276);
not NOT1 (N8281, N8280);
and AND3 (N8282, N8265, N1213, N5251);
nand NAND2 (N8283, N8272, N3269);
not NOT1 (N8284, N8268);
nor NOR3 (N8285, N8259, N1793, N302);
xor XOR2 (N8286, N8285, N2607);
xor XOR2 (N8287, N8286, N7838);
nor NOR3 (N8288, N8277, N1200, N7857);
xor XOR2 (N8289, N8275, N6189);
or OR4 (N8290, N8284, N3952, N514, N3539);
not NOT1 (N8291, N8279);
xor XOR2 (N8292, N8287, N4587);
nand NAND2 (N8293, N8282, N7197);
nor NOR4 (N8294, N8278, N696, N1752, N4796);
nand NAND3 (N8295, N8289, N2295, N6500);
xor XOR2 (N8296, N8281, N7698);
buf BUF1 (N8297, N8295);
buf BUF1 (N8298, N8296);
buf BUF1 (N8299, N8288);
xor XOR2 (N8300, N8293, N6653);
buf BUF1 (N8301, N8299);
and AND4 (N8302, N8294, N7905, N3645, N1687);
nor NOR4 (N8303, N8271, N4732, N2994, N5516);
buf BUF1 (N8304, N8300);
and AND3 (N8305, N8292, N6884, N8249);
nand NAND3 (N8306, N8304, N3300, N3573);
not NOT1 (N8307, N8305);
xor XOR2 (N8308, N8307, N7674);
nor NOR4 (N8309, N8303, N6180, N1981, N4172);
not NOT1 (N8310, N8302);
nand NAND4 (N8311, N8301, N6787, N4009, N256);
nor NOR4 (N8312, N8308, N6316, N8111, N4583);
nor NOR2 (N8313, N8297, N7331);
not NOT1 (N8314, N8283);
and AND3 (N8315, N8314, N756, N4489);
xor XOR2 (N8316, N8298, N5840);
nand NAND4 (N8317, N8313, N5118, N1915, N6656);
xor XOR2 (N8318, N8291, N1073);
and AND2 (N8319, N8306, N4060);
or OR3 (N8320, N8290, N6818, N7683);
xor XOR2 (N8321, N8320, N7490);
buf BUF1 (N8322, N8315);
buf BUF1 (N8323, N8312);
and AND3 (N8324, N8310, N5166, N4851);
not NOT1 (N8325, N8323);
buf BUF1 (N8326, N8316);
not NOT1 (N8327, N8325);
buf BUF1 (N8328, N8321);
or OR3 (N8329, N8311, N417, N7337);
xor XOR2 (N8330, N8319, N74);
not NOT1 (N8331, N8309);
or OR4 (N8332, N8328, N3120, N6474, N2208);
not NOT1 (N8333, N8322);
not NOT1 (N8334, N8327);
xor XOR2 (N8335, N8332, N1866);
buf BUF1 (N8336, N8331);
not NOT1 (N8337, N8324);
buf BUF1 (N8338, N8317);
nand NAND3 (N8339, N8337, N4899, N3234);
and AND2 (N8340, N8329, N187);
buf BUF1 (N8341, N8330);
not NOT1 (N8342, N8333);
buf BUF1 (N8343, N8339);
and AND3 (N8344, N8318, N1521, N7980);
buf BUF1 (N8345, N8340);
not NOT1 (N8346, N8335);
or OR3 (N8347, N8346, N6917, N1506);
not NOT1 (N8348, N8345);
and AND3 (N8349, N8336, N6670, N6019);
xor XOR2 (N8350, N8326, N1066);
xor XOR2 (N8351, N8342, N7776);
not NOT1 (N8352, N8338);
or OR4 (N8353, N8352, N5953, N3596, N7145);
or OR3 (N8354, N8353, N976, N410);
or OR3 (N8355, N8343, N7694, N7013);
xor XOR2 (N8356, N8354, N2242);
nand NAND2 (N8357, N8355, N2031);
not NOT1 (N8358, N8349);
and AND2 (N8359, N8350, N5837);
xor XOR2 (N8360, N8347, N7084);
or OR4 (N8361, N8334, N3235, N5857, N8176);
or OR3 (N8362, N8356, N2699, N1063);
not NOT1 (N8363, N8341);
xor XOR2 (N8364, N8361, N2499);
not NOT1 (N8365, N8359);
or OR2 (N8366, N8344, N6439);
or OR4 (N8367, N8365, N5132, N535, N1475);
or OR4 (N8368, N8358, N4877, N2732, N1220);
nand NAND3 (N8369, N8363, N5117, N1675);
or OR3 (N8370, N8351, N1641, N3899);
nor NOR2 (N8371, N8368, N8186);
and AND2 (N8372, N8367, N6295);
not NOT1 (N8373, N8371);
xor XOR2 (N8374, N8357, N922);
nand NAND2 (N8375, N8369, N977);
xor XOR2 (N8376, N8348, N6819);
nand NAND4 (N8377, N8376, N740, N8054, N6132);
or OR2 (N8378, N8375, N2497);
not NOT1 (N8379, N8364);
nor NOR3 (N8380, N8366, N1357, N95);
not NOT1 (N8381, N8380);
xor XOR2 (N8382, N8379, N2620);
nor NOR2 (N8383, N8378, N6989);
not NOT1 (N8384, N8382);
and AND2 (N8385, N8360, N1371);
nor NOR2 (N8386, N8362, N3075);
not NOT1 (N8387, N8383);
nor NOR3 (N8388, N8374, N1561, N3927);
not NOT1 (N8389, N8385);
nand NAND2 (N8390, N8388, N1954);
xor XOR2 (N8391, N8390, N2931);
buf BUF1 (N8392, N8373);
and AND2 (N8393, N8392, N1201);
xor XOR2 (N8394, N8391, N7470);
not NOT1 (N8395, N8389);
nor NOR2 (N8396, N8372, N5244);
not NOT1 (N8397, N8384);
and AND4 (N8398, N8394, N8058, N6060, N4708);
buf BUF1 (N8399, N8381);
not NOT1 (N8400, N8393);
nand NAND2 (N8401, N8387, N6774);
buf BUF1 (N8402, N8399);
nand NAND4 (N8403, N8398, N4388, N5970, N1602);
or OR4 (N8404, N8400, N3100, N2394, N6156);
nor NOR4 (N8405, N8386, N4856, N5726, N677);
buf BUF1 (N8406, N8397);
buf BUF1 (N8407, N8395);
xor XOR2 (N8408, N8406, N2191);
or OR4 (N8409, N8407, N272, N5593, N7697);
nand NAND3 (N8410, N8377, N3786, N4216);
and AND3 (N8411, N8370, N3440, N1746);
buf BUF1 (N8412, N8401);
nand NAND4 (N8413, N8411, N5487, N2210, N6565);
xor XOR2 (N8414, N8408, N7196);
or OR3 (N8415, N8414, N8368, N8109);
and AND2 (N8416, N8409, N5908);
and AND3 (N8417, N8396, N5550, N8039);
nor NOR4 (N8418, N8413, N6674, N3997, N2286);
buf BUF1 (N8419, N8410);
nand NAND3 (N8420, N8403, N3163, N6432);
nor NOR3 (N8421, N8416, N2696, N4284);
xor XOR2 (N8422, N8418, N120);
not NOT1 (N8423, N8422);
nor NOR4 (N8424, N8423, N5832, N4183, N8042);
nand NAND2 (N8425, N8419, N310);
xor XOR2 (N8426, N8425, N150);
buf BUF1 (N8427, N8412);
not NOT1 (N8428, N8405);
not NOT1 (N8429, N8427);
or OR3 (N8430, N8424, N4883, N2800);
xor XOR2 (N8431, N8402, N2494);
not NOT1 (N8432, N8415);
xor XOR2 (N8433, N8428, N6392);
or OR3 (N8434, N8429, N7487, N6309);
and AND4 (N8435, N8421, N1242, N4248, N740);
and AND4 (N8436, N8430, N1741, N415, N2543);
and AND2 (N8437, N8426, N6359);
and AND2 (N8438, N8435, N7970);
xor XOR2 (N8439, N8433, N8187);
not NOT1 (N8440, N8404);
buf BUF1 (N8441, N8420);
not NOT1 (N8442, N8436);
not NOT1 (N8443, N8439);
buf BUF1 (N8444, N8438);
nand NAND2 (N8445, N8442, N5707);
nor NOR2 (N8446, N8444, N6304);
nor NOR3 (N8447, N8445, N929, N5892);
nor NOR3 (N8448, N8432, N306, N7309);
or OR4 (N8449, N8448, N3486, N4385, N2185);
xor XOR2 (N8450, N8443, N3397);
and AND3 (N8451, N8450, N1191, N3634);
and AND3 (N8452, N8441, N8079, N254);
nor NOR4 (N8453, N8451, N4344, N6565, N7285);
nand NAND2 (N8454, N8447, N5303);
nor NOR4 (N8455, N8452, N5173, N4513, N3765);
buf BUF1 (N8456, N8431);
or OR3 (N8457, N8417, N8313, N671);
buf BUF1 (N8458, N8440);
nor NOR3 (N8459, N8457, N2169, N1298);
buf BUF1 (N8460, N8437);
not NOT1 (N8461, N8453);
buf BUF1 (N8462, N8446);
or OR3 (N8463, N8459, N8149, N5707);
buf BUF1 (N8464, N8461);
and AND3 (N8465, N8434, N6771, N2118);
nand NAND4 (N8466, N8454, N15, N5195, N4608);
not NOT1 (N8467, N8465);
not NOT1 (N8468, N8467);
or OR3 (N8469, N8449, N6401, N5321);
not NOT1 (N8470, N8468);
xor XOR2 (N8471, N8455, N3117);
and AND3 (N8472, N8462, N1687, N4397);
not NOT1 (N8473, N8458);
nand NAND4 (N8474, N8456, N2652, N400, N3123);
nor NOR4 (N8475, N8470, N6113, N692, N4121);
nor NOR2 (N8476, N8460, N3026);
buf BUF1 (N8477, N8464);
and AND2 (N8478, N8475, N4657);
xor XOR2 (N8479, N8474, N6924);
nand NAND2 (N8480, N8473, N5526);
nand NAND2 (N8481, N8469, N3);
nor NOR2 (N8482, N8478, N5310);
and AND4 (N8483, N8476, N5152, N2382, N4382);
and AND2 (N8484, N8466, N6210);
nor NOR2 (N8485, N8484, N5445);
buf BUF1 (N8486, N8485);
xor XOR2 (N8487, N8463, N1840);
buf BUF1 (N8488, N8481);
or OR2 (N8489, N8483, N3342);
not NOT1 (N8490, N8486);
nand NAND3 (N8491, N8482, N7992, N4680);
or OR3 (N8492, N8488, N7330, N1611);
not NOT1 (N8493, N8487);
buf BUF1 (N8494, N8471);
or OR2 (N8495, N8477, N6971);
or OR4 (N8496, N8491, N7439, N4564, N4677);
and AND4 (N8497, N8490, N4796, N1222, N4444);
buf BUF1 (N8498, N8479);
buf BUF1 (N8499, N8480);
xor XOR2 (N8500, N8494, N1073);
nand NAND3 (N8501, N8499, N7234, N8378);
and AND2 (N8502, N8497, N8456);
nor NOR4 (N8503, N8496, N2446, N5046, N7486);
xor XOR2 (N8504, N8503, N8462);
and AND3 (N8505, N8489, N7487, N2080);
not NOT1 (N8506, N8493);
or OR3 (N8507, N8498, N5206, N1394);
or OR3 (N8508, N8492, N209, N4841);
nand NAND4 (N8509, N8472, N6468, N7225, N5816);
nand NAND3 (N8510, N8495, N7772, N1681);
nor NOR4 (N8511, N8502, N1208, N1545, N1401);
or OR2 (N8512, N8504, N4968);
nand NAND3 (N8513, N8506, N3132, N6614);
nand NAND3 (N8514, N8510, N2022, N8505);
not NOT1 (N8515, N2188);
nor NOR4 (N8516, N8514, N4463, N1657, N6540);
nand NAND2 (N8517, N8516, N2283);
nand NAND4 (N8518, N8500, N6848, N6395, N2910);
nand NAND4 (N8519, N8517, N4016, N5448, N5424);
and AND2 (N8520, N8512, N451);
nor NOR3 (N8521, N8511, N5247, N7281);
nor NOR3 (N8522, N8521, N5763, N3597);
and AND3 (N8523, N8501, N6114, N3994);
nor NOR3 (N8524, N8508, N5093, N725);
not NOT1 (N8525, N8513);
xor XOR2 (N8526, N8507, N4939);
buf BUF1 (N8527, N8523);
buf BUF1 (N8528, N8515);
buf BUF1 (N8529, N8520);
nand NAND2 (N8530, N8524, N5354);
not NOT1 (N8531, N8529);
buf BUF1 (N8532, N8519);
or OR4 (N8533, N8522, N3411, N1391, N2664);
nor NOR4 (N8534, N8530, N3150, N2786, N5949);
and AND3 (N8535, N8533, N1437, N3137);
nand NAND3 (N8536, N8528, N1697, N6925);
nand NAND4 (N8537, N8532, N438, N4637, N7975);
xor XOR2 (N8538, N8527, N4562);
and AND4 (N8539, N8534, N3685, N7352, N6151);
nand NAND2 (N8540, N8538, N471);
nand NAND2 (N8541, N8526, N6577);
buf BUF1 (N8542, N8525);
nor NOR3 (N8543, N8541, N5488, N2000);
or OR2 (N8544, N8509, N3007);
and AND2 (N8545, N8544, N414);
nand NAND2 (N8546, N8539, N2606);
not NOT1 (N8547, N8545);
nand NAND4 (N8548, N8547, N5062, N3573, N2561);
and AND3 (N8549, N8536, N4927, N4509);
xor XOR2 (N8550, N8543, N4406);
not NOT1 (N8551, N8531);
nor NOR3 (N8552, N8540, N2831, N1799);
and AND3 (N8553, N8518, N5198, N1918);
nand NAND3 (N8554, N8537, N2196, N3600);
xor XOR2 (N8555, N8535, N6192);
and AND4 (N8556, N8553, N5392, N4137, N926);
or OR3 (N8557, N8548, N535, N7420);
buf BUF1 (N8558, N8542);
not NOT1 (N8559, N8550);
not NOT1 (N8560, N8554);
or OR3 (N8561, N8546, N5792, N83);
buf BUF1 (N8562, N8558);
xor XOR2 (N8563, N8551, N3656);
xor XOR2 (N8564, N8560, N1818);
nor NOR3 (N8565, N8559, N4468, N8422);
and AND2 (N8566, N8552, N1891);
nand NAND4 (N8567, N8557, N6212, N7422, N5512);
nand NAND2 (N8568, N8549, N5847);
nand NAND2 (N8569, N8564, N4194);
or OR2 (N8570, N8562, N8404);
or OR3 (N8571, N8556, N895, N2417);
nand NAND3 (N8572, N8570, N4969, N1555);
not NOT1 (N8573, N8572);
not NOT1 (N8574, N8563);
or OR4 (N8575, N8574, N4531, N8545, N7523);
xor XOR2 (N8576, N8575, N166);
xor XOR2 (N8577, N8567, N1182);
buf BUF1 (N8578, N8568);
xor XOR2 (N8579, N8573, N3952);
xor XOR2 (N8580, N8569, N3709);
buf BUF1 (N8581, N8566);
nor NOR3 (N8582, N8576, N3657, N3150);
nand NAND2 (N8583, N8555, N4229);
not NOT1 (N8584, N8580);
nor NOR3 (N8585, N8578, N4760, N6422);
xor XOR2 (N8586, N8584, N8427);
nor NOR2 (N8587, N8586, N6445);
xor XOR2 (N8588, N8577, N4095);
nor NOR2 (N8589, N8561, N3692);
xor XOR2 (N8590, N8585, N4254);
xor XOR2 (N8591, N8587, N4996);
nand NAND3 (N8592, N8565, N3734, N5698);
and AND2 (N8593, N8590, N8385);
and AND3 (N8594, N8579, N4730, N8126);
nand NAND3 (N8595, N8594, N2902, N7771);
xor XOR2 (N8596, N8571, N147);
or OR3 (N8597, N8588, N3054, N3102);
nand NAND3 (N8598, N8597, N7914, N4627);
not NOT1 (N8599, N8583);
buf BUF1 (N8600, N8593);
xor XOR2 (N8601, N8592, N2206);
and AND3 (N8602, N8596, N5667, N3121);
not NOT1 (N8603, N8581);
xor XOR2 (N8604, N8598, N1818);
xor XOR2 (N8605, N8602, N338);
xor XOR2 (N8606, N8604, N6742);
or OR4 (N8607, N8605, N7338, N610, N7979);
not NOT1 (N8608, N8591);
not NOT1 (N8609, N8600);
xor XOR2 (N8610, N8601, N7349);
nand NAND3 (N8611, N8610, N2824, N7371);
nand NAND3 (N8612, N8599, N5204, N6793);
not NOT1 (N8613, N8607);
xor XOR2 (N8614, N8589, N559);
xor XOR2 (N8615, N8609, N4017);
and AND3 (N8616, N8606, N5958, N6272);
and AND3 (N8617, N8613, N1041, N1430);
not NOT1 (N8618, N8617);
nor NOR4 (N8619, N8612, N4067, N1164, N6024);
nand NAND3 (N8620, N8614, N8129, N2083);
buf BUF1 (N8621, N8582);
nor NOR4 (N8622, N8620, N8163, N3619, N1930);
and AND2 (N8623, N8618, N3229);
nor NOR4 (N8624, N8608, N3473, N2172, N5930);
nor NOR4 (N8625, N8595, N6220, N5559, N6293);
nand NAND4 (N8626, N8611, N8438, N5955, N2020);
not NOT1 (N8627, N8621);
and AND4 (N8628, N8616, N8021, N981, N3161);
buf BUF1 (N8629, N8622);
nand NAND4 (N8630, N8627, N4982, N1427, N8462);
nand NAND4 (N8631, N8624, N1655, N2833, N7850);
nand NAND2 (N8632, N8628, N3201);
nand NAND2 (N8633, N8625, N3036);
xor XOR2 (N8634, N8630, N5692);
nand NAND2 (N8635, N8623, N6507);
nor NOR2 (N8636, N8634, N6149);
nand NAND3 (N8637, N8603, N5734, N4531);
and AND3 (N8638, N8631, N3046, N2821);
nand NAND3 (N8639, N8638, N1648, N434);
xor XOR2 (N8640, N8629, N1529);
xor XOR2 (N8641, N8635, N2914);
buf BUF1 (N8642, N8633);
nand NAND2 (N8643, N8641, N5528);
or OR3 (N8644, N8639, N406, N8364);
nand NAND3 (N8645, N8642, N8404, N5988);
buf BUF1 (N8646, N8615);
nand NAND2 (N8647, N8646, N4646);
not NOT1 (N8648, N8626);
nor NOR3 (N8649, N8644, N4550, N2307);
xor XOR2 (N8650, N8645, N3063);
or OR2 (N8651, N8636, N2825);
buf BUF1 (N8652, N8650);
nor NOR4 (N8653, N8643, N5319, N2171, N1850);
nand NAND2 (N8654, N8640, N6680);
nand NAND4 (N8655, N8652, N581, N2842, N949);
nand NAND2 (N8656, N8648, N7981);
not NOT1 (N8657, N8619);
or OR2 (N8658, N8647, N1805);
buf BUF1 (N8659, N8656);
and AND3 (N8660, N8651, N2364, N2196);
or OR4 (N8661, N8654, N5894, N3944, N6364);
nand NAND3 (N8662, N8637, N3904, N6489);
nand NAND3 (N8663, N8632, N800, N2855);
and AND3 (N8664, N8662, N2551, N1349);
xor XOR2 (N8665, N8658, N2300);
and AND4 (N8666, N8663, N2267, N6405, N587);
not NOT1 (N8667, N8666);
not NOT1 (N8668, N8661);
nor NOR3 (N8669, N8668, N4033, N560);
nand NAND4 (N8670, N8655, N2888, N3960, N455);
nor NOR3 (N8671, N8653, N2348, N1412);
xor XOR2 (N8672, N8670, N593);
nor NOR3 (N8673, N8665, N271, N4240);
or OR3 (N8674, N8669, N200, N6975);
nor NOR4 (N8675, N8674, N268, N5195, N1033);
nor NOR2 (N8676, N8664, N4144);
not NOT1 (N8677, N8675);
buf BUF1 (N8678, N8677);
not NOT1 (N8679, N8649);
xor XOR2 (N8680, N8660, N1021);
nand NAND4 (N8681, N8678, N6729, N6551, N8147);
buf BUF1 (N8682, N8680);
nand NAND3 (N8683, N8673, N5772, N2747);
not NOT1 (N8684, N8679);
or OR3 (N8685, N8676, N2538, N6436);
buf BUF1 (N8686, N8659);
and AND3 (N8687, N8683, N16, N7244);
not NOT1 (N8688, N8681);
or OR4 (N8689, N8685, N7998, N950, N2676);
xor XOR2 (N8690, N8671, N8246);
not NOT1 (N8691, N8689);
xor XOR2 (N8692, N8682, N3596);
nand NAND3 (N8693, N8686, N6593, N6194);
buf BUF1 (N8694, N8691);
and AND4 (N8695, N8694, N5362, N4171, N2229);
nand NAND3 (N8696, N8688, N8601, N3983);
or OR2 (N8697, N8695, N2853);
xor XOR2 (N8698, N8667, N930);
nand NAND2 (N8699, N8684, N1443);
buf BUF1 (N8700, N8696);
nor NOR3 (N8701, N8700, N7022, N2296);
xor XOR2 (N8702, N8701, N6115);
or OR3 (N8703, N8702, N3725, N8079);
and AND2 (N8704, N8693, N7270);
buf BUF1 (N8705, N8704);
xor XOR2 (N8706, N8692, N1757);
xor XOR2 (N8707, N8672, N7974);
nor NOR2 (N8708, N8657, N4677);
and AND2 (N8709, N8703, N5335);
not NOT1 (N8710, N8708);
not NOT1 (N8711, N8709);
nor NOR3 (N8712, N8687, N1612, N6647);
nand NAND2 (N8713, N8698, N6891);
and AND4 (N8714, N8697, N2503, N3443, N7517);
and AND2 (N8715, N8714, N1634);
buf BUF1 (N8716, N8705);
xor XOR2 (N8717, N8712, N28);
not NOT1 (N8718, N8710);
or OR3 (N8719, N8713, N6158, N4487);
buf BUF1 (N8720, N8715);
or OR3 (N8721, N8699, N8647, N5975);
or OR3 (N8722, N8706, N3177, N2947);
not NOT1 (N8723, N8722);
not NOT1 (N8724, N8718);
nor NOR3 (N8725, N8690, N3381, N8111);
not NOT1 (N8726, N8720);
buf BUF1 (N8727, N8725);
buf BUF1 (N8728, N8716);
nand NAND4 (N8729, N8711, N2820, N2016, N6854);
not NOT1 (N8730, N8721);
buf BUF1 (N8731, N8707);
xor XOR2 (N8732, N8731, N2052);
not NOT1 (N8733, N8723);
nand NAND3 (N8734, N8719, N1872, N5540);
or OR4 (N8735, N8727, N6506, N2993, N4441);
not NOT1 (N8736, N8726);
and AND4 (N8737, N8730, N4334, N3636, N2479);
nor NOR4 (N8738, N8735, N5900, N6285, N212);
nor NOR3 (N8739, N8729, N2227, N7653);
and AND4 (N8740, N8739, N711, N4, N6985);
buf BUF1 (N8741, N8738);
nand NAND3 (N8742, N8732, N1104, N8174);
not NOT1 (N8743, N8736);
and AND3 (N8744, N8740, N8313, N6547);
not NOT1 (N8745, N8733);
not NOT1 (N8746, N8744);
or OR2 (N8747, N8742, N5278);
nor NOR4 (N8748, N8747, N4615, N6727, N413);
and AND3 (N8749, N8728, N1785, N3437);
xor XOR2 (N8750, N8743, N2944);
buf BUF1 (N8751, N8741);
and AND3 (N8752, N8717, N5420, N6567);
buf BUF1 (N8753, N8752);
nand NAND2 (N8754, N8746, N2390);
nor NOR2 (N8755, N8734, N1391);
xor XOR2 (N8756, N8724, N2604);
and AND3 (N8757, N8754, N4023, N6119);
not NOT1 (N8758, N8756);
nor NOR2 (N8759, N8737, N4485);
not NOT1 (N8760, N8748);
or OR3 (N8761, N8760, N8634, N6643);
nand NAND4 (N8762, N8759, N1243, N496, N8426);
nor NOR4 (N8763, N8750, N4774, N1949, N3839);
or OR3 (N8764, N8762, N918, N7007);
nor NOR2 (N8765, N8757, N4322);
or OR2 (N8766, N8758, N1939);
xor XOR2 (N8767, N8764, N6881);
or OR4 (N8768, N8763, N3963, N4639, N2229);
nand NAND3 (N8769, N8768, N3260, N8056);
nand NAND2 (N8770, N8753, N7091);
xor XOR2 (N8771, N8770, N4996);
xor XOR2 (N8772, N8766, N1551);
and AND3 (N8773, N8749, N8236, N5297);
nor NOR3 (N8774, N8773, N1110, N7456);
nand NAND4 (N8775, N8767, N2618, N5647, N7198);
nand NAND4 (N8776, N8755, N390, N8492, N8017);
nor NOR2 (N8777, N8761, N6696);
xor XOR2 (N8778, N8771, N6269);
xor XOR2 (N8779, N8769, N2354);
not NOT1 (N8780, N8777);
not NOT1 (N8781, N8775);
or OR3 (N8782, N8781, N5786, N7458);
nor NOR2 (N8783, N8774, N7884);
not NOT1 (N8784, N8779);
nand NAND2 (N8785, N8745, N2186);
xor XOR2 (N8786, N8784, N2293);
or OR2 (N8787, N8786, N4042);
or OR2 (N8788, N8772, N5409);
xor XOR2 (N8789, N8782, N7057);
nor NOR3 (N8790, N8751, N5493, N5288);
and AND3 (N8791, N8778, N1374, N1517);
not NOT1 (N8792, N8791);
or OR3 (N8793, N8792, N6914, N3487);
nor NOR4 (N8794, N8765, N7123, N4803, N3710);
nand NAND4 (N8795, N8785, N2905, N7532, N5130);
buf BUF1 (N8796, N8794);
or OR2 (N8797, N8776, N6217);
xor XOR2 (N8798, N8793, N485);
not NOT1 (N8799, N8780);
and AND4 (N8800, N8788, N1256, N8337, N8699);
buf BUF1 (N8801, N8789);
not NOT1 (N8802, N8799);
not NOT1 (N8803, N8783);
and AND4 (N8804, N8801, N240, N3522, N5262);
and AND3 (N8805, N8804, N5939, N188);
or OR4 (N8806, N8803, N8776, N2463, N7338);
xor XOR2 (N8807, N8797, N1039);
and AND3 (N8808, N8807, N4180, N7464);
nand NAND4 (N8809, N8802, N1815, N7631, N3017);
buf BUF1 (N8810, N8796);
nor NOR4 (N8811, N8798, N659, N5934, N2544);
or OR4 (N8812, N8790, N2331, N374, N1010);
and AND3 (N8813, N8810, N4717, N7321);
or OR3 (N8814, N8787, N7210, N2363);
nand NAND3 (N8815, N8806, N1218, N5247);
and AND4 (N8816, N8805, N3348, N4551, N3231);
or OR2 (N8817, N8800, N4095);
buf BUF1 (N8818, N8795);
xor XOR2 (N8819, N8818, N7690);
not NOT1 (N8820, N8812);
and AND3 (N8821, N8813, N356, N4468);
nor NOR2 (N8822, N8816, N7517);
nor NOR3 (N8823, N8820, N5059, N7635);
nor NOR2 (N8824, N8811, N5887);
and AND3 (N8825, N8823, N1839, N8679);
nand NAND4 (N8826, N8819, N7556, N457, N2139);
xor XOR2 (N8827, N8809, N4434);
and AND3 (N8828, N8824, N5832, N3322);
nor NOR3 (N8829, N8827, N7511, N3701);
buf BUF1 (N8830, N8817);
and AND4 (N8831, N8825, N5025, N7676, N6392);
or OR4 (N8832, N8821, N2648, N4498, N871);
nand NAND3 (N8833, N8832, N5020, N6405);
not NOT1 (N8834, N8808);
not NOT1 (N8835, N8814);
or OR4 (N8836, N8829, N3926, N1907, N3834);
not NOT1 (N8837, N8815);
and AND4 (N8838, N8831, N3461, N2640, N3763);
nand NAND2 (N8839, N8826, N5993);
buf BUF1 (N8840, N8833);
nor NOR2 (N8841, N8838, N8566);
and AND2 (N8842, N8836, N213);
buf BUF1 (N8843, N8839);
buf BUF1 (N8844, N8842);
or OR4 (N8845, N8844, N8050, N3621, N2188);
buf BUF1 (N8846, N8837);
nor NOR2 (N8847, N8846, N504);
not NOT1 (N8848, N8822);
and AND4 (N8849, N8847, N8297, N4296, N7160);
nor NOR2 (N8850, N8841, N7718);
nand NAND4 (N8851, N8849, N2234, N6647, N1479);
and AND3 (N8852, N8843, N634, N5451);
and AND3 (N8853, N8851, N6375, N7133);
xor XOR2 (N8854, N8845, N5755);
and AND3 (N8855, N8853, N2911, N7321);
buf BUF1 (N8856, N8855);
or OR2 (N8857, N8840, N6494);
nor NOR3 (N8858, N8856, N187, N2180);
and AND2 (N8859, N8854, N5779);
buf BUF1 (N8860, N8828);
or OR2 (N8861, N8835, N21);
buf BUF1 (N8862, N8852);
nand NAND3 (N8863, N8862, N1539, N3022);
or OR4 (N8864, N8830, N4739, N6135, N5293);
and AND4 (N8865, N8864, N3374, N309, N5809);
or OR4 (N8866, N8865, N5352, N3227, N7282);
or OR3 (N8867, N8850, N7659, N152);
xor XOR2 (N8868, N8860, N3215);
not NOT1 (N8869, N8848);
not NOT1 (N8870, N8869);
nand NAND2 (N8871, N8834, N7715);
and AND4 (N8872, N8871, N3220, N8643, N1476);
nand NAND3 (N8873, N8861, N2236, N7872);
nand NAND2 (N8874, N8870, N7276);
nor NOR3 (N8875, N8859, N6408, N5697);
not NOT1 (N8876, N8868);
or OR4 (N8877, N8867, N7193, N913, N5738);
not NOT1 (N8878, N8875);
nor NOR4 (N8879, N8863, N2351, N7131, N1380);
nand NAND3 (N8880, N8866, N3324, N3868);
nor NOR3 (N8881, N8872, N608, N4);
xor XOR2 (N8882, N8874, N7569);
and AND4 (N8883, N8873, N171, N7402, N5415);
and AND3 (N8884, N8857, N8529, N5432);
not NOT1 (N8885, N8880);
and AND2 (N8886, N8883, N2231);
xor XOR2 (N8887, N8879, N5726);
buf BUF1 (N8888, N8886);
nand NAND2 (N8889, N8881, N2135);
buf BUF1 (N8890, N8878);
nor NOR2 (N8891, N8885, N7326);
xor XOR2 (N8892, N8858, N1231);
nor NOR4 (N8893, N8889, N3659, N6071, N763);
nor NOR2 (N8894, N8891, N2603);
or OR3 (N8895, N8894, N4053, N1625);
not NOT1 (N8896, N8890);
not NOT1 (N8897, N8884);
and AND4 (N8898, N8896, N4837, N1138, N7610);
buf BUF1 (N8899, N8897);
or OR2 (N8900, N8882, N7264);
or OR2 (N8901, N8898, N2385);
not NOT1 (N8902, N8888);
not NOT1 (N8903, N8900);
buf BUF1 (N8904, N8899);
xor XOR2 (N8905, N8877, N7784);
and AND4 (N8906, N8895, N7540, N7569, N4891);
not NOT1 (N8907, N8876);
nand NAND4 (N8908, N8904, N8883, N2298, N3396);
or OR4 (N8909, N8893, N1388, N667, N2893);
nand NAND2 (N8910, N8906, N1026);
xor XOR2 (N8911, N8903, N3186);
xor XOR2 (N8912, N8909, N3070);
or OR2 (N8913, N8902, N3546);
and AND3 (N8914, N8913, N5445, N3933);
not NOT1 (N8915, N8892);
buf BUF1 (N8916, N8915);
xor XOR2 (N8917, N8910, N8261);
nand NAND4 (N8918, N8917, N7966, N6990, N3501);
nor NOR3 (N8919, N8907, N5290, N8511);
and AND3 (N8920, N8911, N3274, N7233);
and AND4 (N8921, N8920, N1056, N5477, N3319);
buf BUF1 (N8922, N8919);
not NOT1 (N8923, N8887);
nand NAND2 (N8924, N8916, N606);
not NOT1 (N8925, N8905);
and AND4 (N8926, N8921, N3837, N4775, N8209);
nor NOR4 (N8927, N8908, N1408, N5609, N7875);
or OR4 (N8928, N8924, N8549, N5806, N1890);
nand NAND2 (N8929, N8928, N1747);
nand NAND4 (N8930, N8922, N6376, N3952, N7052);
or OR2 (N8931, N8929, N7934);
not NOT1 (N8932, N8925);
nor NOR3 (N8933, N8923, N6465, N7765);
or OR3 (N8934, N8926, N4663, N4322);
buf BUF1 (N8935, N8914);
and AND2 (N8936, N8934, N755);
and AND4 (N8937, N8927, N1268, N7807, N5461);
or OR4 (N8938, N8935, N7456, N7855, N4850);
nor NOR2 (N8939, N8931, N2969);
not NOT1 (N8940, N8936);
xor XOR2 (N8941, N8940, N3607);
not NOT1 (N8942, N8941);
nor NOR3 (N8943, N8918, N136, N695);
or OR3 (N8944, N8942, N6127, N6215);
xor XOR2 (N8945, N8938, N6810);
and AND3 (N8946, N8901, N7777, N4807);
not NOT1 (N8947, N8932);
or OR3 (N8948, N8945, N950, N3032);
xor XOR2 (N8949, N8948, N8283);
buf BUF1 (N8950, N8943);
buf BUF1 (N8951, N8912);
nor NOR4 (N8952, N8933, N8910, N5258, N629);
not NOT1 (N8953, N8946);
nand NAND2 (N8954, N8953, N6758);
and AND3 (N8955, N8939, N4804, N6914);
xor XOR2 (N8956, N8930, N6720);
and AND4 (N8957, N8949, N6238, N5624, N4045);
nand NAND3 (N8958, N8950, N4993, N48);
nor NOR2 (N8959, N8958, N7703);
buf BUF1 (N8960, N8944);
and AND3 (N8961, N8954, N2649, N1646);
nand NAND3 (N8962, N8960, N6154, N1166);
xor XOR2 (N8963, N8955, N2749);
xor XOR2 (N8964, N8957, N6223);
or OR3 (N8965, N8952, N5043, N7618);
not NOT1 (N8966, N8959);
not NOT1 (N8967, N8951);
nand NAND4 (N8968, N8947, N291, N4556, N6710);
or OR2 (N8969, N8937, N4758);
or OR2 (N8970, N8969, N3977);
and AND3 (N8971, N8964, N3436, N5494);
nand NAND4 (N8972, N8963, N1387, N2123, N3957);
and AND4 (N8973, N8965, N537, N8940, N3065);
or OR3 (N8974, N8956, N4760, N60);
buf BUF1 (N8975, N8974);
nor NOR2 (N8976, N8966, N6321);
and AND2 (N8977, N8972, N140);
and AND4 (N8978, N8962, N8061, N2302, N1047);
xor XOR2 (N8979, N8978, N840);
not NOT1 (N8980, N8973);
xor XOR2 (N8981, N8971, N8701);
nor NOR2 (N8982, N8981, N3452);
xor XOR2 (N8983, N8961, N3252);
and AND3 (N8984, N8977, N2032, N239);
buf BUF1 (N8985, N8979);
nand NAND4 (N8986, N8982, N3122, N8034, N6413);
not NOT1 (N8987, N8984);
or OR2 (N8988, N8980, N6567);
nor NOR2 (N8989, N8970, N4823);
xor XOR2 (N8990, N8983, N453);
nor NOR4 (N8991, N8985, N2742, N5049, N7640);
and AND4 (N8992, N8968, N7567, N5772, N8356);
not NOT1 (N8993, N8967);
or OR2 (N8994, N8986, N6688);
nor NOR2 (N8995, N8975, N1887);
not NOT1 (N8996, N8993);
nor NOR4 (N8997, N8994, N8677, N7763, N6223);
and AND4 (N8998, N8995, N8932, N5397, N3437);
nor NOR3 (N8999, N8992, N6634, N8841);
nor NOR2 (N9000, N8991, N2142);
not NOT1 (N9001, N8989);
or OR2 (N9002, N9000, N5317);
and AND3 (N9003, N8990, N4526, N4948);
and AND3 (N9004, N8996, N7473, N5954);
xor XOR2 (N9005, N9003, N5629);
nand NAND2 (N9006, N8999, N3221);
or OR2 (N9007, N8976, N6028);
and AND4 (N9008, N8997, N8761, N2596, N3211);
nand NAND2 (N9009, N9001, N3878);
not NOT1 (N9010, N9008);
or OR4 (N9011, N9007, N6441, N1864, N8214);
or OR2 (N9012, N9002, N6188);
buf BUF1 (N9013, N8998);
or OR4 (N9014, N9005, N2212, N7428, N5649);
nand NAND4 (N9015, N8988, N8426, N1626, N6455);
or OR4 (N9016, N9011, N2569, N8662, N256);
or OR4 (N9017, N9014, N1480, N2891, N6482);
xor XOR2 (N9018, N9009, N7784);
or OR4 (N9019, N9004, N7452, N5859, N5805);
or OR2 (N9020, N9019, N3144);
or OR2 (N9021, N9013, N2014);
buf BUF1 (N9022, N9015);
and AND3 (N9023, N9012, N5347, N3146);
or OR4 (N9024, N9017, N3003, N2757, N7932);
buf BUF1 (N9025, N9021);
or OR3 (N9026, N9010, N4883, N2388);
nand NAND2 (N9027, N9016, N7306);
nand NAND2 (N9028, N9027, N173);
nor NOR2 (N9029, N9023, N3548);
nor NOR3 (N9030, N9026, N2308, N4308);
nand NAND3 (N9031, N9024, N3207, N6253);
nand NAND3 (N9032, N9028, N5004, N6946);
not NOT1 (N9033, N9020);
or OR2 (N9034, N9032, N4018);
not NOT1 (N9035, N9033);
or OR4 (N9036, N9022, N5685, N2550, N6166);
nand NAND3 (N9037, N9006, N4103, N1340);
nand NAND2 (N9038, N9036, N578);
xor XOR2 (N9039, N9030, N8710);
xor XOR2 (N9040, N9031, N5346);
and AND4 (N9041, N9035, N4900, N7760, N6984);
nor NOR3 (N9042, N9025, N4973, N2850);
or OR4 (N9043, N9018, N8417, N6877, N5227);
buf BUF1 (N9044, N9041);
nand NAND3 (N9045, N9043, N1061, N8457);
nor NOR2 (N9046, N9037, N1653);
buf BUF1 (N9047, N9029);
or OR4 (N9048, N9045, N3158, N2267, N9015);
nand NAND2 (N9049, N9044, N7515);
xor XOR2 (N9050, N9039, N776);
and AND4 (N9051, N9049, N1953, N3403, N4302);
not NOT1 (N9052, N9046);
nor NOR2 (N9053, N9050, N4358);
or OR3 (N9054, N9040, N3608, N3204);
xor XOR2 (N9055, N9038, N4623);
buf BUF1 (N9056, N9054);
and AND2 (N9057, N8987, N5724);
xor XOR2 (N9058, N9055, N1276);
nand NAND4 (N9059, N9047, N7377, N8775, N3337);
not NOT1 (N9060, N9056);
nand NAND2 (N9061, N9048, N4974);
xor XOR2 (N9062, N9042, N625);
nor NOR3 (N9063, N9034, N5857, N3430);
nand NAND2 (N9064, N9051, N8268);
nor NOR3 (N9065, N9059, N1986, N6939);
not NOT1 (N9066, N9058);
xor XOR2 (N9067, N9063, N8592);
buf BUF1 (N9068, N9052);
xor XOR2 (N9069, N9062, N4071);
buf BUF1 (N9070, N9065);
and AND2 (N9071, N9057, N8837);
nor NOR3 (N9072, N9068, N2849, N8963);
not NOT1 (N9073, N9064);
nand NAND3 (N9074, N9060, N2537, N2440);
xor XOR2 (N9075, N9074, N5693);
and AND4 (N9076, N9073, N1277, N1956, N7725);
and AND3 (N9077, N9069, N8812, N998);
nor NOR3 (N9078, N9053, N7776, N5260);
xor XOR2 (N9079, N9066, N7716);
and AND2 (N9080, N9079, N7084);
buf BUF1 (N9081, N9076);
or OR3 (N9082, N9075, N6521, N9035);
nand NAND4 (N9083, N9078, N7681, N7614, N7698);
or OR2 (N9084, N9067, N5305);
or OR3 (N9085, N9081, N648, N6643);
buf BUF1 (N9086, N9083);
nor NOR4 (N9087, N9061, N7416, N1052, N6082);
buf BUF1 (N9088, N9080);
and AND4 (N9089, N9072, N2308, N1526, N6119);
or OR4 (N9090, N9082, N7464, N8657, N7777);
xor XOR2 (N9091, N9071, N5004);
xor XOR2 (N9092, N9090, N1754);
not NOT1 (N9093, N9086);
not NOT1 (N9094, N9070);
nand NAND2 (N9095, N9087, N3229);
and AND4 (N9096, N9089, N3551, N8389, N3766);
nor NOR4 (N9097, N9093, N5238, N8980, N1359);
not NOT1 (N9098, N9077);
buf BUF1 (N9099, N9088);
or OR4 (N9100, N9095, N5869, N2645, N8507);
nor NOR4 (N9101, N9100, N29, N5975, N4479);
xor XOR2 (N9102, N9092, N8886);
or OR4 (N9103, N9097, N8676, N92, N6706);
not NOT1 (N9104, N9098);
not NOT1 (N9105, N9096);
and AND4 (N9106, N9085, N8374, N5136, N3226);
or OR4 (N9107, N9084, N7301, N650, N5596);
or OR2 (N9108, N9101, N5031);
or OR2 (N9109, N9102, N2753);
not NOT1 (N9110, N9109);
or OR3 (N9111, N9105, N2994, N5883);
nor NOR2 (N9112, N9091, N7535);
xor XOR2 (N9113, N9106, N1574);
or OR2 (N9114, N9113, N975);
xor XOR2 (N9115, N9099, N2045);
buf BUF1 (N9116, N9115);
buf BUF1 (N9117, N9110);
nand NAND2 (N9118, N9107, N4181);
nor NOR2 (N9119, N9118, N7828);
xor XOR2 (N9120, N9104, N2441);
or OR3 (N9121, N9117, N5861, N4636);
and AND3 (N9122, N9103, N2219, N3615);
or OR3 (N9123, N9121, N7608, N1312);
xor XOR2 (N9124, N9111, N6851);
or OR3 (N9125, N9114, N4658, N4978);
and AND2 (N9126, N9120, N2691);
nor NOR4 (N9127, N9124, N382, N3778, N5226);
xor XOR2 (N9128, N9125, N2640);
nor NOR3 (N9129, N9094, N1789, N6503);
buf BUF1 (N9130, N9116);
not NOT1 (N9131, N9119);
and AND4 (N9132, N9130, N1110, N8757, N3078);
or OR2 (N9133, N9123, N5346);
xor XOR2 (N9134, N9108, N3896);
or OR3 (N9135, N9122, N7939, N4505);
or OR2 (N9136, N9112, N3155);
and AND2 (N9137, N9126, N5146);
xor XOR2 (N9138, N9131, N6399);
not NOT1 (N9139, N9134);
buf BUF1 (N9140, N9127);
xor XOR2 (N9141, N9132, N6495);
nand NAND4 (N9142, N9137, N1165, N4164, N6044);
nor NOR2 (N9143, N9140, N4358);
nor NOR3 (N9144, N9128, N4678, N6480);
not NOT1 (N9145, N9144);
not NOT1 (N9146, N9139);
or OR4 (N9147, N9133, N4340, N1202, N1989);
buf BUF1 (N9148, N9142);
xor XOR2 (N9149, N9129, N2903);
or OR2 (N9150, N9138, N2685);
xor XOR2 (N9151, N9141, N6049);
buf BUF1 (N9152, N9145);
nand NAND4 (N9153, N9135, N6744, N1900, N8039);
not NOT1 (N9154, N9136);
buf BUF1 (N9155, N9149);
buf BUF1 (N9156, N9155);
nand NAND4 (N9157, N9146, N2652, N5553, N2246);
and AND4 (N9158, N9152, N1274, N5202, N5388);
and AND4 (N9159, N9150, N2212, N6155, N2637);
nand NAND4 (N9160, N9147, N3486, N7124, N2059);
buf BUF1 (N9161, N9148);
nand NAND2 (N9162, N9143, N4154);
or OR3 (N9163, N9158, N1967, N7401);
or OR2 (N9164, N9163, N679);
not NOT1 (N9165, N9160);
nor NOR4 (N9166, N9156, N1526, N1135, N4154);
nand NAND2 (N9167, N9151, N1353);
nand NAND2 (N9168, N9164, N520);
buf BUF1 (N9169, N9165);
buf BUF1 (N9170, N9162);
or OR4 (N9171, N9154, N5114, N1784, N8993);
nor NOR4 (N9172, N9170, N7086, N7914, N252);
and AND2 (N9173, N9169, N3493);
xor XOR2 (N9174, N9173, N794);
nand NAND3 (N9175, N9157, N2118, N3807);
xor XOR2 (N9176, N9172, N4565);
nor NOR4 (N9177, N9166, N6418, N5687, N5686);
xor XOR2 (N9178, N9175, N6204);
xor XOR2 (N9179, N9168, N8112);
nor NOR2 (N9180, N9179, N8034);
not NOT1 (N9181, N9177);
and AND3 (N9182, N9153, N7890, N2287);
nor NOR2 (N9183, N9181, N4965);
xor XOR2 (N9184, N9159, N3146);
buf BUF1 (N9185, N9176);
nand NAND2 (N9186, N9161, N6934);
and AND3 (N9187, N9167, N3906, N8464);
not NOT1 (N9188, N9178);
xor XOR2 (N9189, N9182, N7848);
buf BUF1 (N9190, N9185);
buf BUF1 (N9191, N9188);
buf BUF1 (N9192, N9184);
not NOT1 (N9193, N9187);
not NOT1 (N9194, N9192);
or OR4 (N9195, N9180, N3108, N3677, N3559);
not NOT1 (N9196, N9191);
or OR2 (N9197, N9193, N230);
nand NAND4 (N9198, N9194, N3295, N3679, N8138);
buf BUF1 (N9199, N9190);
and AND3 (N9200, N9197, N604, N5202);
and AND3 (N9201, N9198, N339, N2833);
buf BUF1 (N9202, N9183);
not NOT1 (N9203, N9186);
nor NOR4 (N9204, N9189, N3854, N6958, N2538);
or OR2 (N9205, N9204, N2794);
not NOT1 (N9206, N9195);
nand NAND2 (N9207, N9205, N4130);
nor NOR4 (N9208, N9174, N4730, N4674, N3016);
buf BUF1 (N9209, N9202);
nor NOR4 (N9210, N9203, N3615, N750, N9099);
buf BUF1 (N9211, N9208);
nor NOR3 (N9212, N9200, N4445, N1431);
and AND3 (N9213, N9171, N6241, N4842);
not NOT1 (N9214, N9210);
xor XOR2 (N9215, N9201, N3651);
and AND3 (N9216, N9215, N5000, N4744);
buf BUF1 (N9217, N9211);
or OR4 (N9218, N9214, N1698, N7338, N6986);
nand NAND2 (N9219, N9196, N7166);
not NOT1 (N9220, N9216);
nand NAND2 (N9221, N9220, N5251);
buf BUF1 (N9222, N9221);
not NOT1 (N9223, N9207);
nand NAND4 (N9224, N9212, N4790, N2910, N5589);
or OR3 (N9225, N9224, N4954, N4526);
nand NAND3 (N9226, N9218, N353, N2167);
nand NAND2 (N9227, N9225, N6313);
nor NOR2 (N9228, N9219, N1042);
buf BUF1 (N9229, N9213);
nor NOR4 (N9230, N9226, N8977, N2699, N2729);
nand NAND4 (N9231, N9199, N8590, N7149, N1641);
nor NOR3 (N9232, N9217, N4310, N6031);
and AND4 (N9233, N9228, N1666, N4922, N5348);
nor NOR3 (N9234, N9223, N3551, N1403);
and AND3 (N9235, N9229, N15, N988);
buf BUF1 (N9236, N9231);
nand NAND2 (N9237, N9233, N9019);
nand NAND3 (N9238, N9232, N6058, N1234);
buf BUF1 (N9239, N9209);
or OR4 (N9240, N9237, N1417, N1820, N1523);
nor NOR2 (N9241, N9240, N3676);
not NOT1 (N9242, N9227);
or OR2 (N9243, N9230, N3392);
or OR2 (N9244, N9206, N9167);
xor XOR2 (N9245, N9238, N3414);
nor NOR2 (N9246, N9245, N2848);
nor NOR3 (N9247, N9243, N9164, N8955);
xor XOR2 (N9248, N9242, N1208);
buf BUF1 (N9249, N9234);
not NOT1 (N9250, N9248);
or OR4 (N9251, N9241, N8460, N607, N8953);
nor NOR2 (N9252, N9244, N6667);
or OR4 (N9253, N9249, N5704, N2730, N6607);
buf BUF1 (N9254, N9253);
nand NAND3 (N9255, N9254, N5098, N7574);
nand NAND2 (N9256, N9235, N918);
buf BUF1 (N9257, N9236);
nor NOR2 (N9258, N9222, N5837);
not NOT1 (N9259, N9256);
not NOT1 (N9260, N9250);
xor XOR2 (N9261, N9252, N1693);
nor NOR3 (N9262, N9239, N4308, N2848);
xor XOR2 (N9263, N9255, N8176);
buf BUF1 (N9264, N9260);
or OR2 (N9265, N9262, N4874);
or OR2 (N9266, N9257, N3129);
not NOT1 (N9267, N9246);
or OR4 (N9268, N9267, N4769, N880, N975);
xor XOR2 (N9269, N9261, N7968);
nor NOR4 (N9270, N9264, N7223, N5609, N1889);
or OR3 (N9271, N9259, N2194, N6920);
xor XOR2 (N9272, N9266, N7241);
and AND2 (N9273, N9258, N4708);
nor NOR4 (N9274, N9265, N229, N4936, N8547);
nand NAND3 (N9275, N9271, N8997, N4562);
buf BUF1 (N9276, N9270);
or OR3 (N9277, N9247, N294, N1840);
xor XOR2 (N9278, N9274, N6621);
nand NAND4 (N9279, N9278, N5234, N3455, N2170);
buf BUF1 (N9280, N9277);
nand NAND2 (N9281, N9273, N32);
nand NAND4 (N9282, N9275, N2542, N1654, N1979);
nor NOR2 (N9283, N9276, N3696);
nand NAND4 (N9284, N9251, N8634, N5822, N2123);
and AND3 (N9285, N9284, N7459, N4491);
or OR4 (N9286, N9280, N5522, N2988, N4643);
not NOT1 (N9287, N9285);
buf BUF1 (N9288, N9281);
or OR3 (N9289, N9282, N5472, N3923);
or OR3 (N9290, N9289, N3644, N7301);
buf BUF1 (N9291, N9283);
or OR3 (N9292, N9268, N6709, N5066);
nor NOR2 (N9293, N9279, N6291);
buf BUF1 (N9294, N9272);
buf BUF1 (N9295, N9290);
nand NAND3 (N9296, N9293, N7927, N6234);
not NOT1 (N9297, N9294);
not NOT1 (N9298, N9288);
not NOT1 (N9299, N9295);
nor NOR3 (N9300, N9297, N7651, N8028);
nand NAND4 (N9301, N9292, N75, N1370, N5227);
not NOT1 (N9302, N9296);
xor XOR2 (N9303, N9300, N8602);
buf BUF1 (N9304, N9298);
or OR4 (N9305, N9303, N1594, N8958, N7942);
xor XOR2 (N9306, N9301, N5817);
nor NOR2 (N9307, N9299, N8459);
not NOT1 (N9308, N9307);
and AND2 (N9309, N9306, N2533);
not NOT1 (N9310, N9302);
not NOT1 (N9311, N9269);
not NOT1 (N9312, N9311);
not NOT1 (N9313, N9287);
xor XOR2 (N9314, N9313, N6318);
and AND4 (N9315, N9310, N1669, N8512, N5080);
and AND2 (N9316, N9305, N802);
nand NAND3 (N9317, N9286, N2487, N3541);
buf BUF1 (N9318, N9309);
buf BUF1 (N9319, N9316);
buf BUF1 (N9320, N9315);
xor XOR2 (N9321, N9263, N205);
and AND4 (N9322, N9314, N7566, N1168, N6622);
nor NOR4 (N9323, N9322, N3437, N6237, N6119);
not NOT1 (N9324, N9321);
xor XOR2 (N9325, N9304, N6948);
not NOT1 (N9326, N9308);
xor XOR2 (N9327, N9325, N2645);
nor NOR3 (N9328, N9319, N860, N8522);
and AND3 (N9329, N9327, N2326, N6809);
xor XOR2 (N9330, N9323, N7454);
or OR2 (N9331, N9320, N979);
xor XOR2 (N9332, N9317, N8737);
buf BUF1 (N9333, N9330);
nor NOR4 (N9334, N9328, N7297, N8830, N2485);
nand NAND2 (N9335, N9329, N8680);
not NOT1 (N9336, N9318);
or OR4 (N9337, N9331, N1903, N1627, N6833);
or OR3 (N9338, N9334, N3419, N5742);
buf BUF1 (N9339, N9312);
nor NOR2 (N9340, N9339, N6756);
not NOT1 (N9341, N9340);
nand NAND3 (N9342, N9341, N1293, N429);
and AND2 (N9343, N9333, N4232);
buf BUF1 (N9344, N9342);
nor NOR3 (N9345, N9326, N1906, N7338);
nor NOR3 (N9346, N9324, N4500, N6823);
and AND3 (N9347, N9335, N222, N7178);
nor NOR3 (N9348, N9291, N6691, N931);
nor NOR4 (N9349, N9348, N1619, N1349, N5856);
nor NOR3 (N9350, N9345, N6352, N192);
or OR3 (N9351, N9344, N3307, N8719);
or OR3 (N9352, N9351, N7619, N1226);
and AND3 (N9353, N9338, N6268, N9177);
not NOT1 (N9354, N9347);
buf BUF1 (N9355, N9352);
nor NOR4 (N9356, N9350, N2384, N1396, N6370);
nor NOR2 (N9357, N9332, N8607);
nor NOR3 (N9358, N9337, N909, N4287);
buf BUF1 (N9359, N9354);
not NOT1 (N9360, N9357);
buf BUF1 (N9361, N9359);
nor NOR3 (N9362, N9336, N3436, N8448);
nor NOR2 (N9363, N9360, N2987);
nand NAND3 (N9364, N9363, N3719, N1759);
or OR3 (N9365, N9358, N7396, N8371);
and AND3 (N9366, N9364, N2998, N5653);
not NOT1 (N9367, N9343);
buf BUF1 (N9368, N9355);
buf BUF1 (N9369, N9368);
buf BUF1 (N9370, N9369);
and AND3 (N9371, N9361, N6203, N2336);
nand NAND4 (N9372, N9371, N4606, N2375, N2696);
xor XOR2 (N9373, N9367, N4339);
xor XOR2 (N9374, N9356, N5658);
buf BUF1 (N9375, N9366);
or OR4 (N9376, N9372, N2615, N7916, N7610);
nor NOR4 (N9377, N9375, N898, N3710, N6088);
nand NAND3 (N9378, N9346, N7823, N5741);
or OR4 (N9379, N9373, N3448, N2090, N40);
xor XOR2 (N9380, N9379, N9220);
xor XOR2 (N9381, N9349, N1090);
not NOT1 (N9382, N9365);
or OR3 (N9383, N9380, N4792, N7674);
nand NAND2 (N9384, N9382, N7914);
or OR4 (N9385, N9377, N6022, N4580, N6626);
nor NOR3 (N9386, N9376, N5028, N3027);
nand NAND3 (N9387, N9383, N1555, N9332);
nor NOR3 (N9388, N9353, N2955, N48);
or OR4 (N9389, N9381, N6914, N3536, N6648);
nor NOR2 (N9390, N9378, N953);
nor NOR3 (N9391, N9374, N3321, N4988);
xor XOR2 (N9392, N9386, N8928);
or OR2 (N9393, N9391, N3770);
or OR3 (N9394, N9384, N3183, N294);
or OR2 (N9395, N9385, N975);
buf BUF1 (N9396, N9390);
nor NOR4 (N9397, N9387, N7813, N4217, N2171);
or OR3 (N9398, N9370, N37, N7237);
and AND3 (N9399, N9392, N676, N2422);
nor NOR3 (N9400, N9397, N1855, N2440);
and AND4 (N9401, N9362, N3950, N6071, N9222);
buf BUF1 (N9402, N9401);
or OR2 (N9403, N9402, N7271);
xor XOR2 (N9404, N9396, N467);
or OR3 (N9405, N9388, N4581, N7315);
xor XOR2 (N9406, N9393, N6088);
not NOT1 (N9407, N9389);
buf BUF1 (N9408, N9400);
and AND3 (N9409, N9398, N3679, N4587);
or OR3 (N9410, N9409, N6230, N1844);
and AND2 (N9411, N9403, N1949);
xor XOR2 (N9412, N9406, N2944);
not NOT1 (N9413, N9410);
nand NAND3 (N9414, N9407, N3441, N8932);
buf BUF1 (N9415, N9405);
nor NOR4 (N9416, N9394, N343, N1705, N1451);
or OR2 (N9417, N9413, N5429);
buf BUF1 (N9418, N9411);
not NOT1 (N9419, N9408);
or OR2 (N9420, N9416, N1790);
or OR3 (N9421, N9414, N7798, N898);
and AND2 (N9422, N9419, N2325);
nor NOR3 (N9423, N9395, N7089, N2776);
not NOT1 (N9424, N9420);
buf BUF1 (N9425, N9418);
xor XOR2 (N9426, N9425, N4287);
buf BUF1 (N9427, N9415);
not NOT1 (N9428, N9424);
and AND3 (N9429, N9399, N3578, N2591);
nand NAND2 (N9430, N9426, N5348);
nor NOR2 (N9431, N9412, N5276);
xor XOR2 (N9432, N9417, N853);
xor XOR2 (N9433, N9422, N7590);
not NOT1 (N9434, N9421);
not NOT1 (N9435, N9404);
nor NOR4 (N9436, N9423, N3467, N7089, N3085);
or OR4 (N9437, N9433, N8022, N1293, N8467);
nor NOR4 (N9438, N9427, N4263, N3094, N2907);
xor XOR2 (N9439, N9436, N3634);
buf BUF1 (N9440, N9428);
or OR2 (N9441, N9440, N3569);
or OR2 (N9442, N9431, N7350);
xor XOR2 (N9443, N9437, N6905);
xor XOR2 (N9444, N9441, N6591);
nand NAND4 (N9445, N9443, N789, N7326, N8919);
or OR4 (N9446, N9445, N5447, N382, N5448);
or OR3 (N9447, N9430, N7003, N5345);
not NOT1 (N9448, N9439);
and AND3 (N9449, N9429, N9170, N1451);
buf BUF1 (N9450, N9432);
xor XOR2 (N9451, N9442, N8405);
buf BUF1 (N9452, N9446);
not NOT1 (N9453, N9434);
or OR2 (N9454, N9438, N3573);
not NOT1 (N9455, N9435);
and AND4 (N9456, N9455, N1160, N994, N3528);
xor XOR2 (N9457, N9449, N8769);
not NOT1 (N9458, N9451);
nor NOR4 (N9459, N9448, N9001, N2013, N7597);
xor XOR2 (N9460, N9453, N198);
nand NAND2 (N9461, N9450, N8143);
buf BUF1 (N9462, N9461);
nor NOR4 (N9463, N9462, N8960, N1071, N5756);
or OR3 (N9464, N9444, N9328, N7260);
and AND2 (N9465, N9458, N6747);
xor XOR2 (N9466, N9456, N5396);
nand NAND4 (N9467, N9465, N9450, N7003, N8039);
not NOT1 (N9468, N9452);
buf BUF1 (N9469, N9468);
nand NAND2 (N9470, N9447, N4902);
and AND4 (N9471, N9463, N686, N817, N269);
and AND4 (N9472, N9467, N6349, N7764, N726);
buf BUF1 (N9473, N9457);
and AND4 (N9474, N9466, N7950, N6590, N2074);
and AND2 (N9475, N9473, N9258);
nor NOR2 (N9476, N9459, N5745);
nand NAND4 (N9477, N9475, N6448, N3703, N582);
buf BUF1 (N9478, N9469);
nand NAND2 (N9479, N9460, N638);
buf BUF1 (N9480, N9464);
xor XOR2 (N9481, N9470, N6387);
nand NAND2 (N9482, N9474, N8356);
nor NOR4 (N9483, N9454, N4807, N4608, N989);
xor XOR2 (N9484, N9478, N7828);
or OR3 (N9485, N9481, N6859, N5932);
nor NOR2 (N9486, N9480, N2425);
not NOT1 (N9487, N9484);
nor NOR2 (N9488, N9487, N2645);
nand NAND4 (N9489, N9483, N3506, N6135, N4913);
nand NAND4 (N9490, N9477, N8948, N1582, N8038);
xor XOR2 (N9491, N9486, N5893);
nand NAND2 (N9492, N9482, N2313);
xor XOR2 (N9493, N9472, N3660);
and AND2 (N9494, N9493, N1366);
not NOT1 (N9495, N9471);
or OR2 (N9496, N9489, N812);
and AND3 (N9497, N9495, N310, N2537);
nand NAND2 (N9498, N9479, N5391);
not NOT1 (N9499, N9496);
nand NAND4 (N9500, N9497, N4202, N113, N9005);
xor XOR2 (N9501, N9499, N5456);
nand NAND3 (N9502, N9488, N9296, N8661);
nor NOR2 (N9503, N9494, N3146);
buf BUF1 (N9504, N9501);
buf BUF1 (N9505, N9500);
and AND4 (N9506, N9492, N3670, N6561, N1711);
buf BUF1 (N9507, N9476);
not NOT1 (N9508, N9506);
buf BUF1 (N9509, N9503);
or OR2 (N9510, N9490, N7915);
xor XOR2 (N9511, N9504, N7564);
nor NOR2 (N9512, N9505, N2492);
not NOT1 (N9513, N9508);
and AND3 (N9514, N9507, N6967, N821);
or OR4 (N9515, N9491, N5069, N3828, N6742);
nor NOR4 (N9516, N9485, N7615, N2903, N7543);
xor XOR2 (N9517, N9511, N5288);
and AND3 (N9518, N9509, N486, N6365);
nand NAND3 (N9519, N9515, N611, N8183);
nor NOR2 (N9520, N9519, N8872);
xor XOR2 (N9521, N9520, N3838);
and AND2 (N9522, N9518, N9240);
and AND3 (N9523, N9516, N3807, N2158);
and AND3 (N9524, N9521, N5173, N8866);
nand NAND4 (N9525, N9498, N3348, N3489, N9264);
not NOT1 (N9526, N9524);
nor NOR2 (N9527, N9522, N7529);
and AND2 (N9528, N9526, N292);
or OR4 (N9529, N9513, N8656, N7981, N413);
or OR3 (N9530, N9523, N5948, N2937);
buf BUF1 (N9531, N9529);
buf BUF1 (N9532, N9512);
nor NOR2 (N9533, N9528, N6228);
xor XOR2 (N9534, N9527, N7441);
nand NAND3 (N9535, N9510, N1960, N8376);
or OR2 (N9536, N9532, N1113);
and AND2 (N9537, N9502, N5513);
nor NOR4 (N9538, N9534, N65, N378, N8798);
not NOT1 (N9539, N9538);
not NOT1 (N9540, N9517);
buf BUF1 (N9541, N9514);
buf BUF1 (N9542, N9530);
and AND3 (N9543, N9533, N1150, N4888);
not NOT1 (N9544, N9543);
xor XOR2 (N9545, N9535, N1945);
buf BUF1 (N9546, N9539);
or OR4 (N9547, N9531, N1740, N5678, N8328);
nor NOR3 (N9548, N9537, N6864, N8464);
nor NOR4 (N9549, N9548, N2024, N6366, N6675);
or OR4 (N9550, N9547, N3505, N599, N6088);
not NOT1 (N9551, N9540);
or OR2 (N9552, N9550, N3711);
or OR2 (N9553, N9551, N4694);
buf BUF1 (N9554, N9544);
nor NOR3 (N9555, N9546, N7980, N2533);
nand NAND4 (N9556, N9541, N4043, N7822, N7862);
or OR2 (N9557, N9542, N5586);
nor NOR2 (N9558, N9545, N4682);
or OR4 (N9559, N9556, N6510, N5223, N8082);
or OR4 (N9560, N9559, N3319, N4039, N5809);
xor XOR2 (N9561, N9560, N3433);
or OR4 (N9562, N9536, N8234, N1314, N4748);
xor XOR2 (N9563, N9549, N4830);
not NOT1 (N9564, N9552);
not NOT1 (N9565, N9561);
or OR4 (N9566, N9565, N3940, N6180, N1961);
nor NOR3 (N9567, N9554, N3285, N8985);
nor NOR4 (N9568, N9525, N5895, N1370, N3378);
or OR4 (N9569, N9555, N2374, N4864, N6423);
buf BUF1 (N9570, N9566);
or OR4 (N9571, N9567, N1448, N6285, N6173);
xor XOR2 (N9572, N9558, N7548);
or OR2 (N9573, N9570, N5744);
nand NAND3 (N9574, N9568, N6766, N9107);
xor XOR2 (N9575, N9571, N7121);
not NOT1 (N9576, N9569);
nand NAND2 (N9577, N9562, N3108);
xor XOR2 (N9578, N9563, N7736);
nand NAND3 (N9579, N9573, N8097, N2356);
and AND4 (N9580, N9577, N1392, N8674, N7348);
not NOT1 (N9581, N9578);
and AND2 (N9582, N9575, N9157);
xor XOR2 (N9583, N9564, N1170);
xor XOR2 (N9584, N9581, N4491);
and AND2 (N9585, N9574, N4209);
xor XOR2 (N9586, N9557, N1473);
or OR2 (N9587, N9585, N4899);
not NOT1 (N9588, N9553);
xor XOR2 (N9589, N9582, N8982);
and AND4 (N9590, N9584, N103, N1114, N8858);
not NOT1 (N9591, N9590);
and AND3 (N9592, N9591, N6534, N5256);
not NOT1 (N9593, N9588);
nand NAND2 (N9594, N9586, N74);
or OR3 (N9595, N9593, N5850, N5984);
nand NAND4 (N9596, N9579, N1587, N1258, N4706);
or OR2 (N9597, N9592, N7388);
not NOT1 (N9598, N9576);
and AND2 (N9599, N9596, N3438);
nand NAND3 (N9600, N9594, N6155, N2996);
or OR4 (N9601, N9600, N7814, N3984, N1111);
not NOT1 (N9602, N9601);
or OR4 (N9603, N9587, N4154, N4648, N2583);
nand NAND2 (N9604, N9572, N916);
not NOT1 (N9605, N9604);
and AND3 (N9606, N9580, N8533, N9301);
nor NOR3 (N9607, N9605, N8877, N783);
not NOT1 (N9608, N9595);
xor XOR2 (N9609, N9599, N3573);
or OR4 (N9610, N9598, N9459, N4351, N1712);
nand NAND4 (N9611, N9608, N1183, N5470, N9457);
xor XOR2 (N9612, N9589, N5875);
not NOT1 (N9613, N9597);
not NOT1 (N9614, N9603);
or OR2 (N9615, N9614, N7765);
nor NOR3 (N9616, N9602, N7041, N873);
and AND4 (N9617, N9611, N5053, N3113, N3268);
and AND2 (N9618, N9613, N3643);
nor NOR3 (N9619, N9615, N4506, N3075);
nor NOR2 (N9620, N9612, N1353);
nor NOR3 (N9621, N9618, N4400, N2786);
not NOT1 (N9622, N9607);
nor NOR3 (N9623, N9610, N8511, N9354);
nand NAND4 (N9624, N9609, N8720, N4084, N6854);
buf BUF1 (N9625, N9617);
nand NAND2 (N9626, N9623, N4056);
nand NAND3 (N9627, N9622, N1297, N4917);
or OR3 (N9628, N9621, N5219, N3131);
nor NOR4 (N9629, N9583, N6026, N1393, N496);
nand NAND2 (N9630, N9629, N662);
xor XOR2 (N9631, N9628, N6823);
buf BUF1 (N9632, N9620);
or OR2 (N9633, N9616, N9349);
nand NAND2 (N9634, N9606, N851);
nand NAND2 (N9635, N9627, N5992);
nand NAND4 (N9636, N9626, N5469, N4445, N833);
buf BUF1 (N9637, N9635);
buf BUF1 (N9638, N9634);
nor NOR4 (N9639, N9632, N4147, N9465, N9227);
xor XOR2 (N9640, N9630, N5315);
or OR4 (N9641, N9631, N6972, N7446, N6277);
or OR4 (N9642, N9625, N6840, N2736, N2334);
buf BUF1 (N9643, N9633);
nor NOR3 (N9644, N9637, N8243, N6115);
nor NOR3 (N9645, N9639, N5202, N1767);
nor NOR4 (N9646, N9643, N6074, N8379, N4845);
not NOT1 (N9647, N9624);
buf BUF1 (N9648, N9640);
nor NOR4 (N9649, N9641, N8611, N9531, N2527);
or OR3 (N9650, N9636, N2030, N5410);
and AND2 (N9651, N9646, N5457);
nand NAND4 (N9652, N9648, N9547, N5506, N8443);
nor NOR4 (N9653, N9645, N9625, N8938, N4471);
nand NAND3 (N9654, N9653, N2668, N7968);
buf BUF1 (N9655, N9619);
nand NAND3 (N9656, N9651, N1401, N7599);
and AND3 (N9657, N9644, N1381, N357);
and AND3 (N9658, N9650, N1839, N672);
xor XOR2 (N9659, N9638, N8506);
nor NOR4 (N9660, N9652, N6172, N5849, N5165);
and AND4 (N9661, N9659, N6462, N2514, N8956);
nor NOR4 (N9662, N9642, N6491, N3808, N2935);
not NOT1 (N9663, N9647);
nor NOR2 (N9664, N9654, N4491);
buf BUF1 (N9665, N9657);
buf BUF1 (N9666, N9663);
buf BUF1 (N9667, N9665);
xor XOR2 (N9668, N9656, N5035);
or OR2 (N9669, N9664, N8826);
not NOT1 (N9670, N9649);
nand NAND2 (N9671, N9660, N5282);
not NOT1 (N9672, N9667);
and AND3 (N9673, N9669, N7449, N7282);
nand NAND3 (N9674, N9672, N2246, N2516);
xor XOR2 (N9675, N9662, N7078);
not NOT1 (N9676, N9658);
and AND3 (N9677, N9673, N7490, N7175);
and AND4 (N9678, N9675, N9109, N375, N2413);
or OR4 (N9679, N9670, N6587, N7724, N5338);
nand NAND4 (N9680, N9676, N7168, N2908, N1134);
nand NAND4 (N9681, N9674, N4784, N7060, N827);
or OR3 (N9682, N9671, N8611, N253);
nor NOR3 (N9683, N9682, N4107, N5027);
nand NAND3 (N9684, N9681, N5502, N755);
buf BUF1 (N9685, N9661);
buf BUF1 (N9686, N9678);
buf BUF1 (N9687, N9686);
xor XOR2 (N9688, N9668, N8543);
or OR2 (N9689, N9680, N4793);
not NOT1 (N9690, N9687);
buf BUF1 (N9691, N9684);
nor NOR2 (N9692, N9655, N7519);
buf BUF1 (N9693, N9679);
not NOT1 (N9694, N9693);
not NOT1 (N9695, N9692);
xor XOR2 (N9696, N9666, N729);
xor XOR2 (N9697, N9689, N1240);
not NOT1 (N9698, N9690);
xor XOR2 (N9699, N9677, N9003);
nor NOR2 (N9700, N9696, N6898);
buf BUF1 (N9701, N9695);
not NOT1 (N9702, N9701);
not NOT1 (N9703, N9691);
nor NOR3 (N9704, N9700, N871, N1652);
xor XOR2 (N9705, N9683, N2535);
nor NOR2 (N9706, N9704, N1519);
and AND3 (N9707, N9699, N3277, N2000);
buf BUF1 (N9708, N9694);
buf BUF1 (N9709, N9688);
xor XOR2 (N9710, N9698, N6194);
nand NAND2 (N9711, N9702, N894);
nor NOR2 (N9712, N9707, N5844);
or OR2 (N9713, N9697, N7738);
and AND3 (N9714, N9706, N1615, N602);
not NOT1 (N9715, N9711);
buf BUF1 (N9716, N9708);
nor NOR3 (N9717, N9712, N2151, N4696);
buf BUF1 (N9718, N9705);
not NOT1 (N9719, N9710);
and AND3 (N9720, N9703, N6740, N8183);
and AND2 (N9721, N9715, N78);
nor NOR4 (N9722, N9716, N5063, N2802, N4974);
xor XOR2 (N9723, N9714, N2497);
nor NOR2 (N9724, N9717, N5988);
xor XOR2 (N9725, N9713, N3779);
and AND3 (N9726, N9722, N4609, N5955);
xor XOR2 (N9727, N9724, N3411);
nand NAND2 (N9728, N9723, N4449);
nand NAND4 (N9729, N9719, N3551, N1343, N940);
nand NAND2 (N9730, N9718, N1139);
not NOT1 (N9731, N9729);
xor XOR2 (N9732, N9685, N2042);
and AND4 (N9733, N9731, N7951, N5313, N3889);
nor NOR4 (N9734, N9730, N881, N9578, N1652);
xor XOR2 (N9735, N9709, N7223);
xor XOR2 (N9736, N9725, N8646);
buf BUF1 (N9737, N9734);
nand NAND3 (N9738, N9720, N2400, N1135);
xor XOR2 (N9739, N9728, N5060);
xor XOR2 (N9740, N9737, N6342);
and AND2 (N9741, N9740, N7737);
nor NOR4 (N9742, N9741, N353, N9356, N3791);
nor NOR3 (N9743, N9739, N2157, N2613);
nand NAND3 (N9744, N9735, N2857, N566);
not NOT1 (N9745, N9736);
xor XOR2 (N9746, N9727, N6170);
or OR3 (N9747, N9726, N7334, N2243);
nand NAND4 (N9748, N9743, N8989, N3681, N7622);
buf BUF1 (N9749, N9748);
xor XOR2 (N9750, N9721, N6911);
and AND3 (N9751, N9733, N7234, N2236);
nor NOR3 (N9752, N9751, N274, N8238);
and AND4 (N9753, N9732, N7057, N1608, N1077);
buf BUF1 (N9754, N9738);
buf BUF1 (N9755, N9745);
or OR3 (N9756, N9746, N569, N4071);
nand NAND2 (N9757, N9756, N9446);
not NOT1 (N9758, N9753);
or OR3 (N9759, N9744, N7321, N8721);
and AND3 (N9760, N9755, N4015, N2104);
nor NOR3 (N9761, N9754, N9613, N2686);
buf BUF1 (N9762, N9760);
xor XOR2 (N9763, N9747, N8951);
buf BUF1 (N9764, N9742);
nor NOR2 (N9765, N9758, N6406);
buf BUF1 (N9766, N9759);
not NOT1 (N9767, N9763);
xor XOR2 (N9768, N9766, N9616);
nand NAND2 (N9769, N9749, N3350);
xor XOR2 (N9770, N9769, N6103);
not NOT1 (N9771, N9768);
buf BUF1 (N9772, N9765);
buf BUF1 (N9773, N9761);
or OR2 (N9774, N9770, N3586);
buf BUF1 (N9775, N9762);
nand NAND4 (N9776, N9757, N1471, N148, N2131);
buf BUF1 (N9777, N9772);
nand NAND3 (N9778, N9752, N1193, N7660);
and AND4 (N9779, N9775, N5654, N22, N8047);
nand NAND3 (N9780, N9773, N4376, N3017);
nand NAND4 (N9781, N9767, N2516, N1740, N8697);
xor XOR2 (N9782, N9779, N9715);
nand NAND3 (N9783, N9771, N1723, N2151);
buf BUF1 (N9784, N9778);
or OR2 (N9785, N9777, N1311);
nand NAND3 (N9786, N9781, N5659, N9155);
xor XOR2 (N9787, N9780, N1615);
buf BUF1 (N9788, N9774);
nand NAND4 (N9789, N9787, N5642, N8665, N9655);
and AND2 (N9790, N9750, N6675);
buf BUF1 (N9791, N9786);
or OR3 (N9792, N9788, N698, N2631);
nand NAND3 (N9793, N9785, N3200, N6263);
and AND4 (N9794, N9776, N2716, N5346, N8877);
nand NAND4 (N9795, N9790, N4182, N45, N6595);
and AND4 (N9796, N9784, N6799, N8788, N6561);
not NOT1 (N9797, N9782);
nand NAND2 (N9798, N9791, N5049);
or OR3 (N9799, N9764, N8733, N1850);
nor NOR3 (N9800, N9796, N5820, N7898);
nand NAND2 (N9801, N9800, N763);
not NOT1 (N9802, N9792);
nor NOR4 (N9803, N9789, N6713, N3325, N9324);
and AND2 (N9804, N9799, N6460);
nor NOR2 (N9805, N9801, N2415);
nor NOR4 (N9806, N9783, N4379, N3849, N1032);
nor NOR4 (N9807, N9797, N7892, N8539, N9765);
and AND3 (N9808, N9793, N6089, N4241);
or OR4 (N9809, N9804, N5188, N6075, N8423);
nand NAND3 (N9810, N9802, N4588, N9422);
nor NOR2 (N9811, N9808, N4355);
xor XOR2 (N9812, N9803, N4927);
nor NOR2 (N9813, N9794, N2061);
or OR4 (N9814, N9807, N113, N3070, N9174);
buf BUF1 (N9815, N9810);
or OR4 (N9816, N9805, N549, N9138, N3154);
buf BUF1 (N9817, N9816);
buf BUF1 (N9818, N9814);
xor XOR2 (N9819, N9818, N1689);
xor XOR2 (N9820, N9812, N5359);
not NOT1 (N9821, N9819);
nand NAND2 (N9822, N9821, N4336);
and AND3 (N9823, N9798, N5408, N4358);
or OR2 (N9824, N9823, N889);
xor XOR2 (N9825, N9809, N9076);
buf BUF1 (N9826, N9817);
nor NOR4 (N9827, N9815, N8084, N2106, N2977);
xor XOR2 (N9828, N9827, N8999);
nor NOR4 (N9829, N9826, N1012, N8491, N9228);
not NOT1 (N9830, N9829);
buf BUF1 (N9831, N9830);
nor NOR3 (N9832, N9825, N4171, N8179);
xor XOR2 (N9833, N9811, N6518);
nand NAND3 (N9834, N9824, N4007, N4826);
xor XOR2 (N9835, N9828, N3594);
not NOT1 (N9836, N9834);
not NOT1 (N9837, N9835);
and AND2 (N9838, N9806, N4806);
buf BUF1 (N9839, N9838);
xor XOR2 (N9840, N9822, N2769);
buf BUF1 (N9841, N9831);
xor XOR2 (N9842, N9837, N3364);
nand NAND2 (N9843, N9841, N797);
buf BUF1 (N9844, N9820);
xor XOR2 (N9845, N9813, N7960);
xor XOR2 (N9846, N9845, N8431);
buf BUF1 (N9847, N9844);
or OR3 (N9848, N9839, N6696, N4399);
and AND3 (N9849, N9832, N4963, N3028);
and AND3 (N9850, N9848, N6369, N3640);
not NOT1 (N9851, N9843);
nor NOR3 (N9852, N9846, N3993, N3199);
nand NAND3 (N9853, N9840, N8760, N163);
not NOT1 (N9854, N9853);
xor XOR2 (N9855, N9854, N3053);
nand NAND4 (N9856, N9836, N4068, N2999, N6034);
or OR4 (N9857, N9855, N8613, N6942, N4091);
or OR4 (N9858, N9847, N6932, N9266, N7771);
nand NAND2 (N9859, N9851, N7321);
or OR4 (N9860, N9842, N6789, N7626, N8273);
nor NOR2 (N9861, N9849, N3509);
nand NAND2 (N9862, N9857, N1421);
and AND3 (N9863, N9795, N4238, N9084);
not NOT1 (N9864, N9833);
not NOT1 (N9865, N9852);
buf BUF1 (N9866, N9861);
nor NOR3 (N9867, N9866, N1887, N6655);
nand NAND2 (N9868, N9867, N1062);
buf BUF1 (N9869, N9850);
and AND2 (N9870, N9868, N4840);
not NOT1 (N9871, N9858);
nor NOR4 (N9872, N9870, N3118, N9571, N8389);
not NOT1 (N9873, N9859);
nand NAND2 (N9874, N9856, N1453);
not NOT1 (N9875, N9864);
buf BUF1 (N9876, N9875);
nand NAND4 (N9877, N9873, N126, N1847, N5979);
and AND3 (N9878, N9862, N2016, N1399);
and AND4 (N9879, N9876, N6279, N1097, N3773);
or OR3 (N9880, N9863, N3664, N3575);
nor NOR3 (N9881, N9865, N697, N5339);
nand NAND2 (N9882, N9872, N6741);
buf BUF1 (N9883, N9869);
xor XOR2 (N9884, N9860, N2526);
not NOT1 (N9885, N9883);
not NOT1 (N9886, N9879);
nand NAND3 (N9887, N9881, N5845, N7382);
xor XOR2 (N9888, N9885, N969);
nor NOR2 (N9889, N9880, N1428);
not NOT1 (N9890, N9888);
nand NAND2 (N9891, N9886, N2509);
buf BUF1 (N9892, N9877);
nor NOR3 (N9893, N9878, N6622, N6664);
buf BUF1 (N9894, N9884);
and AND2 (N9895, N9882, N1723);
and AND3 (N9896, N9871, N273, N8706);
not NOT1 (N9897, N9874);
nand NAND3 (N9898, N9891, N228, N1839);
buf BUF1 (N9899, N9896);
buf BUF1 (N9900, N9892);
and AND3 (N9901, N9890, N5965, N1533);
or OR2 (N9902, N9889, N3007);
nor NOR2 (N9903, N9899, N9128);
and AND3 (N9904, N9898, N5961, N5264);
or OR4 (N9905, N9887, N7635, N9603, N6603);
not NOT1 (N9906, N9904);
xor XOR2 (N9907, N9906, N7479);
xor XOR2 (N9908, N9900, N46);
nand NAND2 (N9909, N9897, N8846);
nor NOR2 (N9910, N9905, N3396);
nor NOR2 (N9911, N9909, N3650);
and AND4 (N9912, N9902, N6495, N8728, N9861);
or OR4 (N9913, N9908, N4719, N9667, N6505);
or OR4 (N9914, N9895, N3437, N7918, N6754);
xor XOR2 (N9915, N9913, N1723);
xor XOR2 (N9916, N9911, N3405);
or OR4 (N9917, N9915, N3908, N3111, N2797);
not NOT1 (N9918, N9903);
or OR4 (N9919, N9894, N6407, N7380, N3398);
or OR4 (N9920, N9907, N732, N331, N6916);
or OR4 (N9921, N9901, N9903, N5881, N8912);
buf BUF1 (N9922, N9919);
xor XOR2 (N9923, N9912, N9388);
not NOT1 (N9924, N9914);
nor NOR3 (N9925, N9921, N8013, N5864);
or OR3 (N9926, N9925, N9032, N1424);
or OR4 (N9927, N9910, N737, N1346, N4594);
not NOT1 (N9928, N9926);
or OR3 (N9929, N9923, N2352, N9718);
buf BUF1 (N9930, N9918);
buf BUF1 (N9931, N9929);
nand NAND4 (N9932, N9931, N5071, N5647, N2451);
not NOT1 (N9933, N9922);
buf BUF1 (N9934, N9920);
and AND2 (N9935, N9933, N5190);
nand NAND4 (N9936, N9928, N264, N1468, N3786);
not NOT1 (N9937, N9917);
and AND2 (N9938, N9930, N9044);
nor NOR2 (N9939, N9893, N6760);
xor XOR2 (N9940, N9934, N9046);
nand NAND2 (N9941, N9937, N5791);
nand NAND3 (N9942, N9941, N9927, N2991);
xor XOR2 (N9943, N7642, N2874);
nand NAND3 (N9944, N9940, N9221, N7129);
nand NAND3 (N9945, N9935, N1237, N1624);
nor NOR4 (N9946, N9916, N5317, N4870, N4603);
xor XOR2 (N9947, N9945, N570);
nor NOR3 (N9948, N9943, N620, N2336);
buf BUF1 (N9949, N9924);
not NOT1 (N9950, N9936);
not NOT1 (N9951, N9949);
xor XOR2 (N9952, N9948, N5670);
or OR4 (N9953, N9939, N884, N5976, N694);
and AND4 (N9954, N9932, N6279, N5018, N8384);
not NOT1 (N9955, N9951);
buf BUF1 (N9956, N9950);
xor XOR2 (N9957, N9952, N9252);
xor XOR2 (N9958, N9956, N2178);
not NOT1 (N9959, N9954);
nor NOR4 (N9960, N9944, N954, N4884, N9874);
or OR3 (N9961, N9960, N4937, N8542);
or OR2 (N9962, N9953, N457);
xor XOR2 (N9963, N9938, N2528);
nand NAND4 (N9964, N9955, N7478, N3211, N5945);
buf BUF1 (N9965, N9964);
nor NOR2 (N9966, N9958, N6807);
or OR3 (N9967, N9942, N1209, N6593);
buf BUF1 (N9968, N9966);
nor NOR3 (N9969, N9967, N5358, N2457);
xor XOR2 (N9970, N9965, N5794);
and AND2 (N9971, N9959, N5379);
or OR3 (N9972, N9947, N3378, N448);
xor XOR2 (N9973, N9972, N200);
xor XOR2 (N9974, N9973, N6745);
or OR3 (N9975, N9969, N6032, N2120);
and AND2 (N9976, N9971, N9289);
and AND2 (N9977, N9961, N3980);
and AND3 (N9978, N9976, N1755, N6717);
nor NOR3 (N9979, N9963, N1015, N1143);
nand NAND3 (N9980, N9978, N6635, N8734);
and AND4 (N9981, N9977, N2309, N328, N6083);
nand NAND3 (N9982, N9957, N634, N8625);
xor XOR2 (N9983, N9981, N5156);
or OR2 (N9984, N9983, N5411);
and AND2 (N9985, N9968, N1874);
xor XOR2 (N9986, N9984, N2606);
not NOT1 (N9987, N9946);
or OR4 (N9988, N9979, N7049, N5355, N3034);
or OR4 (N9989, N9980, N6906, N8987, N449);
nor NOR3 (N9990, N9988, N6161, N2058);
and AND3 (N9991, N9982, N5501, N4457);
nand NAND3 (N9992, N9991, N6927, N5965);
or OR4 (N9993, N9992, N1234, N8466, N2604);
not NOT1 (N9994, N9990);
nand NAND3 (N9995, N9987, N8308, N9375);
xor XOR2 (N9996, N9993, N1789);
not NOT1 (N9997, N9995);
or OR4 (N9998, N9996, N2619, N6889, N5431);
nand NAND3 (N9999, N9970, N7943, N5411);
buf BUF1 (N10000, N9962);
nand NAND4 (N10001, N9975, N2233, N5807, N3918);
not NOT1 (N10002, N9986);
not NOT1 (N10003, N10000);
buf BUF1 (N10004, N9994);
buf BUF1 (N10005, N9998);
nor NOR4 (N10006, N9999, N2329, N9757, N1067);
and AND2 (N10007, N10005, N2242);
xor XOR2 (N10008, N9974, N206);
and AND2 (N10009, N10007, N7351);
nor NOR3 (N10010, N10001, N5922, N2423);
nand NAND4 (N10011, N10009, N3495, N7971, N2390);
xor XOR2 (N10012, N10010, N7761);
buf BUF1 (N10013, N10008);
nor NOR2 (N10014, N9997, N5219);
xor XOR2 (N10015, N10006, N8803);
nand NAND3 (N10016, N10004, N1052, N5214);
buf BUF1 (N10017, N10002);
xor XOR2 (N10018, N10017, N4800);
xor XOR2 (N10019, N10013, N4780);
and AND2 (N10020, N9985, N9905);
not NOT1 (N10021, N10003);
not NOT1 (N10022, N10011);
and AND2 (N10023, N10021, N2236);
nor NOR3 (N10024, N10022, N8575, N7280);
nand NAND2 (N10025, N10014, N5979);
buf BUF1 (N10026, N10025);
nand NAND4 (N10027, N10026, N2474, N3320, N5152);
nand NAND4 (N10028, N10012, N2307, N4258, N2760);
nand NAND4 (N10029, N10019, N8535, N2565, N8644);
nand NAND2 (N10030, N10024, N1825);
xor XOR2 (N10031, N10023, N2776);
xor XOR2 (N10032, N10031, N5628);
buf BUF1 (N10033, N10030);
nand NAND4 (N10034, N10033, N1961, N4328, N1731);
and AND2 (N10035, N10016, N656);
xor XOR2 (N10036, N10035, N5006);
or OR3 (N10037, N10036, N3168, N593);
buf BUF1 (N10038, N9989);
or OR3 (N10039, N10027, N3618, N31);
and AND2 (N10040, N10029, N6418);
xor XOR2 (N10041, N10034, N6618);
nor NOR3 (N10042, N10037, N47, N2669);
nand NAND3 (N10043, N10041, N4407, N9736);
nor NOR4 (N10044, N10028, N9639, N9734, N4674);
buf BUF1 (N10045, N10042);
not NOT1 (N10046, N10015);
xor XOR2 (N10047, N10046, N4314);
buf BUF1 (N10048, N10039);
xor XOR2 (N10049, N10038, N830);
xor XOR2 (N10050, N10020, N416);
xor XOR2 (N10051, N10040, N7369);
xor XOR2 (N10052, N10048, N1550);
nor NOR4 (N10053, N10043, N1861, N2287, N8542);
not NOT1 (N10054, N10053);
not NOT1 (N10055, N10032);
buf BUF1 (N10056, N10050);
buf BUF1 (N10057, N10051);
nor NOR4 (N10058, N10044, N8478, N8320, N2249);
xor XOR2 (N10059, N10058, N7611);
or OR4 (N10060, N10059, N8269, N9867, N6677);
xor XOR2 (N10061, N10056, N9977);
nand NAND2 (N10062, N10061, N1006);
not NOT1 (N10063, N10054);
not NOT1 (N10064, N10062);
not NOT1 (N10065, N10063);
and AND4 (N10066, N10018, N2806, N7308, N2886);
xor XOR2 (N10067, N10055, N7752);
buf BUF1 (N10068, N10057);
nand NAND3 (N10069, N10060, N1559, N8604);
nor NOR3 (N10070, N10052, N2150, N9468);
not NOT1 (N10071, N10066);
nor NOR4 (N10072, N10070, N6010, N5271, N8244);
nor NOR3 (N10073, N10045, N8926, N29);
and AND4 (N10074, N10072, N6292, N9151, N4765);
nor NOR3 (N10075, N10065, N2352, N4017);
nand NAND2 (N10076, N10068, N310);
nand NAND3 (N10077, N10064, N7902, N9513);
not NOT1 (N10078, N10047);
or OR4 (N10079, N10069, N5086, N9923, N4583);
and AND3 (N10080, N10073, N3250, N4169);
or OR3 (N10081, N10079, N3124, N9494);
xor XOR2 (N10082, N10077, N5590);
nor NOR3 (N10083, N10078, N2917, N7453);
nor NOR4 (N10084, N10081, N2972, N4136, N3254);
and AND3 (N10085, N10049, N5759, N6703);
not NOT1 (N10086, N10076);
xor XOR2 (N10087, N10067, N504);
buf BUF1 (N10088, N10082);
or OR2 (N10089, N10071, N3793);
xor XOR2 (N10090, N10080, N9559);
nor NOR3 (N10091, N10089, N3132, N3928);
and AND3 (N10092, N10090, N1766, N8021);
nand NAND3 (N10093, N10085, N796, N1879);
or OR3 (N10094, N10075, N6918, N6796);
buf BUF1 (N10095, N10093);
and AND2 (N10096, N10074, N3045);
buf BUF1 (N10097, N10088);
not NOT1 (N10098, N10087);
and AND3 (N10099, N10084, N2860, N8569);
nand NAND2 (N10100, N10098, N5813);
buf BUF1 (N10101, N10099);
xor XOR2 (N10102, N10083, N6220);
and AND2 (N10103, N10094, N3050);
xor XOR2 (N10104, N10097, N2635);
and AND4 (N10105, N10086, N79, N9457, N355);
or OR4 (N10106, N10101, N4673, N2865, N661);
nand NAND2 (N10107, N10106, N1630);
nor NOR3 (N10108, N10103, N7021, N2107);
or OR3 (N10109, N10105, N2328, N6330);
xor XOR2 (N10110, N10108, N6123);
xor XOR2 (N10111, N10095, N3619);
nor NOR4 (N10112, N10110, N7590, N4415, N8785);
nand NAND4 (N10113, N10100, N4389, N2648, N6084);
or OR4 (N10114, N10113, N8481, N1008, N1077);
xor XOR2 (N10115, N10107, N4109);
not NOT1 (N10116, N10104);
not NOT1 (N10117, N10091);
nor NOR2 (N10118, N10117, N886);
nand NAND4 (N10119, N10114, N2444, N3754, N3476);
nor NOR2 (N10120, N10102, N5967);
nor NOR2 (N10121, N10109, N1507);
nor NOR3 (N10122, N10119, N8500, N3937);
nand NAND4 (N10123, N10118, N483, N1977, N3739);
not NOT1 (N10124, N10123);
not NOT1 (N10125, N10112);
buf BUF1 (N10126, N10092);
and AND3 (N10127, N10125, N6293, N1187);
and AND4 (N10128, N10115, N2495, N6992, N3262);
or OR2 (N10129, N10126, N6510);
xor XOR2 (N10130, N10120, N9727);
xor XOR2 (N10131, N10129, N4483);
or OR4 (N10132, N10131, N3925, N7838, N8239);
not NOT1 (N10133, N10111);
and AND4 (N10134, N10130, N5776, N8274, N4908);
nand NAND3 (N10135, N10134, N1175, N796);
nor NOR3 (N10136, N10116, N6269, N6767);
nand NAND2 (N10137, N10133, N2968);
or OR4 (N10138, N10136, N9172, N8997, N7731);
and AND2 (N10139, N10132, N10074);
nand NAND2 (N10140, N10137, N989);
buf BUF1 (N10141, N10128);
or OR4 (N10142, N10139, N10061, N6474, N9782);
or OR4 (N10143, N10135, N7864, N845, N1859);
nand NAND4 (N10144, N10096, N5118, N1698, N1033);
buf BUF1 (N10145, N10127);
not NOT1 (N10146, N10144);
buf BUF1 (N10147, N10145);
or OR3 (N10148, N10147, N5091, N7348);
nand NAND2 (N10149, N10143, N2239);
or OR4 (N10150, N10141, N5545, N3546, N7723);
xor XOR2 (N10151, N10150, N2224);
and AND2 (N10152, N10138, N5310);
buf BUF1 (N10153, N10148);
or OR3 (N10154, N10140, N239, N7439);
nand NAND4 (N10155, N10142, N8727, N2277, N389);
nand NAND3 (N10156, N10152, N4751, N2119);
buf BUF1 (N10157, N10155);
buf BUF1 (N10158, N10124);
nor NOR3 (N10159, N10154, N1504, N8753);
nor NOR3 (N10160, N10149, N3007, N5458);
xor XOR2 (N10161, N10158, N7141);
not NOT1 (N10162, N10156);
nand NAND4 (N10163, N10161, N3250, N9116, N3953);
nor NOR2 (N10164, N10163, N4324);
buf BUF1 (N10165, N10159);
buf BUF1 (N10166, N10157);
nand NAND3 (N10167, N10153, N5982, N6786);
nor NOR2 (N10168, N10164, N963);
nand NAND2 (N10169, N10122, N6091);
not NOT1 (N10170, N10151);
not NOT1 (N10171, N10146);
buf BUF1 (N10172, N10168);
xor XOR2 (N10173, N10162, N4372);
or OR4 (N10174, N10167, N5983, N8355, N1111);
xor XOR2 (N10175, N10165, N3058);
nand NAND2 (N10176, N10169, N7441);
buf BUF1 (N10177, N10174);
nor NOR3 (N10178, N10173, N5816, N6255);
not NOT1 (N10179, N10166);
and AND3 (N10180, N10170, N8109, N9350);
or OR3 (N10181, N10160, N2505, N697);
nor NOR4 (N10182, N10172, N1745, N4193, N4597);
buf BUF1 (N10183, N10121);
buf BUF1 (N10184, N10178);
buf BUF1 (N10185, N10177);
or OR4 (N10186, N10183, N6758, N6366, N821);
and AND2 (N10187, N10185, N9332);
not NOT1 (N10188, N10182);
nand NAND2 (N10189, N10171, N8974);
nor NOR2 (N10190, N10175, N1347);
buf BUF1 (N10191, N10189);
not NOT1 (N10192, N10190);
buf BUF1 (N10193, N10184);
or OR2 (N10194, N10193, N984);
or OR3 (N10195, N10186, N9882, N8375);
and AND2 (N10196, N10187, N8492);
xor XOR2 (N10197, N10179, N7623);
and AND4 (N10198, N10192, N4069, N1627, N1348);
or OR4 (N10199, N10194, N4235, N3329, N6382);
nand NAND4 (N10200, N10180, N2791, N6124, N8137);
nand NAND4 (N10201, N10200, N7671, N2866, N6551);
and AND4 (N10202, N10198, N1191, N7980, N3886);
nand NAND3 (N10203, N10188, N4740, N2337);
xor XOR2 (N10204, N10181, N5368);
and AND2 (N10205, N10203, N4229);
and AND3 (N10206, N10201, N1383, N6398);
nor NOR4 (N10207, N10196, N3712, N6085, N509);
and AND4 (N10208, N10205, N7987, N8053, N691);
or OR3 (N10209, N10202, N5086, N6407);
buf BUF1 (N10210, N10197);
or OR2 (N10211, N10207, N7303);
or OR4 (N10212, N10176, N9425, N3376, N4753);
buf BUF1 (N10213, N10204);
or OR2 (N10214, N10211, N10191);
not NOT1 (N10215, N9521);
nor NOR4 (N10216, N10208, N4682, N6623, N2059);
and AND4 (N10217, N10216, N7438, N5062, N2367);
buf BUF1 (N10218, N10217);
xor XOR2 (N10219, N10215, N684);
or OR3 (N10220, N10219, N3111, N6385);
nand NAND3 (N10221, N10210, N8332, N7310);
nor NOR2 (N10222, N10218, N7942);
and AND4 (N10223, N10222, N8803, N9399, N5025);
xor XOR2 (N10224, N10213, N2909);
buf BUF1 (N10225, N10195);
nor NOR4 (N10226, N10199, N1487, N3540, N9618);
nand NAND3 (N10227, N10223, N1310, N4870);
xor XOR2 (N10228, N10227, N6249);
and AND3 (N10229, N10221, N5686, N7289);
xor XOR2 (N10230, N10224, N7244);
nand NAND2 (N10231, N10225, N3658);
buf BUF1 (N10232, N10229);
nor NOR2 (N10233, N10212, N849);
nand NAND2 (N10234, N10220, N6857);
xor XOR2 (N10235, N10230, N5925);
not NOT1 (N10236, N10226);
xor XOR2 (N10237, N10228, N3149);
nand NAND2 (N10238, N10236, N4870);
nand NAND3 (N10239, N10235, N308, N5371);
xor XOR2 (N10240, N10231, N9464);
xor XOR2 (N10241, N10206, N1751);
xor XOR2 (N10242, N10237, N3554);
or OR4 (N10243, N10233, N6833, N4439, N5692);
or OR3 (N10244, N10214, N3045, N3483);
nor NOR4 (N10245, N10232, N5857, N7182, N8468);
not NOT1 (N10246, N10240);
nor NOR3 (N10247, N10246, N3190, N5223);
nand NAND4 (N10248, N10241, N5728, N8700, N3410);
nor NOR4 (N10249, N10248, N3359, N3476, N6731);
nand NAND4 (N10250, N10238, N1037, N1190, N5722);
or OR4 (N10251, N10250, N7352, N6734, N1617);
or OR3 (N10252, N10247, N3091, N3320);
nand NAND3 (N10253, N10243, N5944, N1940);
nor NOR2 (N10254, N10251, N5688);
buf BUF1 (N10255, N10234);
nand NAND2 (N10256, N10245, N4304);
and AND3 (N10257, N10255, N4306, N6029);
and AND4 (N10258, N10242, N8723, N2203, N4338);
nor NOR2 (N10259, N10256, N4313);
buf BUF1 (N10260, N10244);
buf BUF1 (N10261, N10253);
nand NAND3 (N10262, N10259, N10035, N3636);
xor XOR2 (N10263, N10254, N5189);
and AND2 (N10264, N10262, N4203);
nand NAND2 (N10265, N10264, N8069);
nand NAND2 (N10266, N10260, N5532);
xor XOR2 (N10267, N10258, N2782);
not NOT1 (N10268, N10249);
nor NOR2 (N10269, N10267, N9946);
xor XOR2 (N10270, N10266, N2667);
buf BUF1 (N10271, N10252);
xor XOR2 (N10272, N10268, N9232);
and AND3 (N10273, N10263, N9643, N4206);
xor XOR2 (N10274, N10272, N1632);
nand NAND2 (N10275, N10265, N7899);
buf BUF1 (N10276, N10275);
and AND4 (N10277, N10276, N4197, N4419, N2731);
not NOT1 (N10278, N10239);
buf BUF1 (N10279, N10271);
and AND2 (N10280, N10261, N9923);
and AND3 (N10281, N10279, N10203, N9365);
nand NAND4 (N10282, N10278, N9339, N7392, N2664);
nor NOR2 (N10283, N10257, N8881);
and AND2 (N10284, N10281, N3302);
buf BUF1 (N10285, N10280);
and AND3 (N10286, N10277, N1896, N3462);
nand NAND2 (N10287, N10283, N8307);
xor XOR2 (N10288, N10270, N9221);
nor NOR3 (N10289, N10284, N3420, N2082);
buf BUF1 (N10290, N10273);
xor XOR2 (N10291, N10286, N329);
nand NAND2 (N10292, N10288, N1004);
nand NAND2 (N10293, N10274, N2523);
not NOT1 (N10294, N10291);
nand NAND4 (N10295, N10293, N3964, N2152, N2864);
buf BUF1 (N10296, N10292);
xor XOR2 (N10297, N10290, N1732);
nor NOR4 (N10298, N10209, N2222, N8973, N4468);
nand NAND3 (N10299, N10285, N3688, N5009);
nor NOR2 (N10300, N10298, N1793);
xor XOR2 (N10301, N10282, N7900);
buf BUF1 (N10302, N10299);
nand NAND2 (N10303, N10297, N6728);
xor XOR2 (N10304, N10300, N1106);
or OR4 (N10305, N10296, N9843, N9669, N7488);
xor XOR2 (N10306, N10295, N7116);
nor NOR4 (N10307, N10287, N6377, N6190, N8159);
nand NAND2 (N10308, N10305, N347);
or OR4 (N10309, N10304, N3164, N5483, N6);
buf BUF1 (N10310, N10309);
or OR2 (N10311, N10303, N4785);
or OR3 (N10312, N10289, N7061, N8991);
and AND2 (N10313, N10308, N2790);
xor XOR2 (N10314, N10302, N4920);
and AND2 (N10315, N10301, N1891);
nand NAND4 (N10316, N10311, N8566, N6345, N3790);
xor XOR2 (N10317, N10316, N799);
nor NOR4 (N10318, N10310, N8561, N2344, N4559);
nand NAND3 (N10319, N10269, N7792, N8136);
xor XOR2 (N10320, N10306, N6130);
or OR4 (N10321, N10312, N9007, N5112, N1799);
xor XOR2 (N10322, N10315, N8915);
not NOT1 (N10323, N10319);
or OR3 (N10324, N10321, N2537, N4079);
buf BUF1 (N10325, N10314);
nand NAND2 (N10326, N10317, N9036);
or OR2 (N10327, N10318, N5460);
nor NOR3 (N10328, N10320, N1672, N9991);
nand NAND3 (N10329, N10325, N577, N5690);
nor NOR2 (N10330, N10327, N6830);
nor NOR3 (N10331, N10322, N3223, N5033);
xor XOR2 (N10332, N10294, N572);
buf BUF1 (N10333, N10326);
buf BUF1 (N10334, N10307);
buf BUF1 (N10335, N10323);
and AND3 (N10336, N10332, N3472, N3713);
or OR2 (N10337, N10328, N3421);
and AND2 (N10338, N10337, N6143);
xor XOR2 (N10339, N10313, N5977);
xor XOR2 (N10340, N10338, N7720);
xor XOR2 (N10341, N10340, N1918);
and AND3 (N10342, N10330, N7808, N3976);
xor XOR2 (N10343, N10324, N3935);
xor XOR2 (N10344, N10334, N8225);
buf BUF1 (N10345, N10344);
nand NAND2 (N10346, N10331, N5225);
nand NAND4 (N10347, N10345, N3281, N8940, N478);
xor XOR2 (N10348, N10335, N4060);
or OR2 (N10349, N10339, N2513);
xor XOR2 (N10350, N10336, N2053);
buf BUF1 (N10351, N10341);
and AND4 (N10352, N10351, N10189, N8517, N1201);
nor NOR4 (N10353, N10349, N2471, N1076, N7897);
nand NAND2 (N10354, N10352, N8451);
nor NOR2 (N10355, N10348, N9845);
buf BUF1 (N10356, N10329);
nand NAND3 (N10357, N10347, N10230, N1590);
and AND3 (N10358, N10355, N4967, N1383);
buf BUF1 (N10359, N10346);
nor NOR3 (N10360, N10359, N2537, N981);
nor NOR4 (N10361, N10342, N7091, N2453, N5897);
buf BUF1 (N10362, N10357);
and AND2 (N10363, N10358, N864);
or OR4 (N10364, N10354, N6620, N5086, N7980);
and AND3 (N10365, N10362, N5958, N274);
or OR4 (N10366, N10361, N2840, N5719, N8356);
and AND2 (N10367, N10333, N3451);
buf BUF1 (N10368, N10353);
nand NAND4 (N10369, N10363, N7920, N8314, N3450);
not NOT1 (N10370, N10368);
buf BUF1 (N10371, N10369);
nor NOR2 (N10372, N10370, N7156);
or OR4 (N10373, N10343, N9134, N1413, N8282);
buf BUF1 (N10374, N10364);
buf BUF1 (N10375, N10366);
nor NOR2 (N10376, N10356, N4888);
nand NAND4 (N10377, N10365, N1235, N8073, N7263);
nor NOR4 (N10378, N10350, N426, N673, N4393);
nor NOR2 (N10379, N10377, N8353);
buf BUF1 (N10380, N10376);
and AND3 (N10381, N10375, N8499, N7605);
and AND4 (N10382, N10380, N7196, N9864, N451);
buf BUF1 (N10383, N10374);
or OR2 (N10384, N10360, N4236);
or OR2 (N10385, N10382, N3584);
xor XOR2 (N10386, N10383, N10209);
xor XOR2 (N10387, N10371, N1223);
or OR3 (N10388, N10372, N8886, N1594);
nor NOR3 (N10389, N10379, N7334, N9505);
not NOT1 (N10390, N10381);
buf BUF1 (N10391, N10390);
or OR4 (N10392, N10388, N3028, N128, N1542);
not NOT1 (N10393, N10387);
or OR4 (N10394, N10393, N7984, N319, N20);
not NOT1 (N10395, N10367);
not NOT1 (N10396, N10384);
and AND3 (N10397, N10396, N9032, N1048);
buf BUF1 (N10398, N10391);
buf BUF1 (N10399, N10398);
and AND3 (N10400, N10394, N722, N7865);
nand NAND2 (N10401, N10386, N1534);
buf BUF1 (N10402, N10385);
buf BUF1 (N10403, N10395);
or OR4 (N10404, N10392, N2840, N4331, N1868);
not NOT1 (N10405, N10400);
not NOT1 (N10406, N10401);
or OR3 (N10407, N10373, N7339, N9967);
not NOT1 (N10408, N10399);
or OR2 (N10409, N10406, N8703);
xor XOR2 (N10410, N10378, N1311);
buf BUF1 (N10411, N10405);
or OR2 (N10412, N10407, N6413);
buf BUF1 (N10413, N10412);
buf BUF1 (N10414, N10402);
nor NOR4 (N10415, N10404, N5196, N991, N3040);
nor NOR2 (N10416, N10397, N6601);
or OR3 (N10417, N10411, N7341, N8856);
not NOT1 (N10418, N10415);
nor NOR4 (N10419, N10417, N917, N8835, N6918);
or OR3 (N10420, N10419, N4747, N4087);
xor XOR2 (N10421, N10410, N9167);
xor XOR2 (N10422, N10408, N6474);
nand NAND4 (N10423, N10422, N9342, N5543, N1581);
nand NAND2 (N10424, N10420, N2917);
buf BUF1 (N10425, N10416);
nand NAND4 (N10426, N10413, N8658, N4310, N1858);
or OR2 (N10427, N10424, N3907);
nor NOR3 (N10428, N10425, N7405, N8727);
buf BUF1 (N10429, N10409);
not NOT1 (N10430, N10418);
and AND2 (N10431, N10427, N6306);
xor XOR2 (N10432, N10421, N2655);
buf BUF1 (N10433, N10414);
not NOT1 (N10434, N10431);
not NOT1 (N10435, N10428);
not NOT1 (N10436, N10430);
nor NOR3 (N10437, N10403, N1957, N7899);
nand NAND4 (N10438, N10435, N7987, N1193, N8933);
nand NAND3 (N10439, N10426, N9034, N2813);
or OR4 (N10440, N10423, N5799, N7866, N7334);
nor NOR2 (N10441, N10436, N1556);
xor XOR2 (N10442, N10437, N8421);
nand NAND4 (N10443, N10442, N9558, N8228, N8563);
nor NOR2 (N10444, N10439, N3962);
or OR4 (N10445, N10443, N1184, N5739, N2392);
nor NOR3 (N10446, N10441, N9191, N1669);
nand NAND2 (N10447, N10429, N9713);
not NOT1 (N10448, N10440);
not NOT1 (N10449, N10445);
or OR4 (N10450, N10449, N10331, N5393, N8740);
nand NAND3 (N10451, N10447, N10004, N5334);
buf BUF1 (N10452, N10446);
and AND2 (N10453, N10438, N1394);
nor NOR2 (N10454, N10433, N7656);
xor XOR2 (N10455, N10454, N5449);
and AND2 (N10456, N10448, N1827);
buf BUF1 (N10457, N10450);
and AND4 (N10458, N10453, N7980, N4330, N7866);
or OR2 (N10459, N10451, N6957);
xor XOR2 (N10460, N10459, N7797);
buf BUF1 (N10461, N10434);
nor NOR4 (N10462, N10460, N5270, N10069, N4614);
buf BUF1 (N10463, N10432);
xor XOR2 (N10464, N10463, N373);
or OR2 (N10465, N10389, N4497);
not NOT1 (N10466, N10452);
nor NOR2 (N10467, N10457, N5416);
xor XOR2 (N10468, N10444, N7418);
and AND2 (N10469, N10465, N8008);
buf BUF1 (N10470, N10466);
buf BUF1 (N10471, N10456);
buf BUF1 (N10472, N10455);
not NOT1 (N10473, N10472);
or OR3 (N10474, N10461, N7861, N10412);
xor XOR2 (N10475, N10467, N7472);
or OR2 (N10476, N10462, N8811);
buf BUF1 (N10477, N10473);
buf BUF1 (N10478, N10477);
or OR2 (N10479, N10464, N4283);
nand NAND2 (N10480, N10470, N7854);
nor NOR3 (N10481, N10468, N7963, N8756);
nor NOR3 (N10482, N10479, N4677, N1167);
or OR2 (N10483, N10458, N7089);
or OR2 (N10484, N10483, N820);
buf BUF1 (N10485, N10484);
xor XOR2 (N10486, N10478, N7523);
not NOT1 (N10487, N10485);
and AND4 (N10488, N10482, N1621, N10184, N5406);
nor NOR4 (N10489, N10471, N9802, N8548, N6034);
or OR2 (N10490, N10487, N8994);
or OR4 (N10491, N10480, N9327, N4986, N8168);
nand NAND2 (N10492, N10488, N8623);
nor NOR2 (N10493, N10481, N9348);
buf BUF1 (N10494, N10475);
nor NOR2 (N10495, N10490, N4113);
nand NAND4 (N10496, N10469, N8774, N4506, N2372);
not NOT1 (N10497, N10489);
xor XOR2 (N10498, N10495, N143);
or OR3 (N10499, N10496, N5105, N9232);
nand NAND3 (N10500, N10476, N2902, N7457);
or OR3 (N10501, N10500, N3443, N2069);
not NOT1 (N10502, N10501);
or OR4 (N10503, N10498, N7239, N125, N4117);
not NOT1 (N10504, N10492);
buf BUF1 (N10505, N10503);
nand NAND4 (N10506, N10474, N5073, N6404, N7577);
nor NOR4 (N10507, N10499, N96, N2456, N8535);
and AND4 (N10508, N10491, N4027, N31, N7997);
xor XOR2 (N10509, N10505, N9546);
xor XOR2 (N10510, N10507, N1848);
not NOT1 (N10511, N10502);
nor NOR4 (N10512, N10504, N3211, N7201, N8880);
and AND3 (N10513, N10510, N7459, N7237);
xor XOR2 (N10514, N10506, N4093);
and AND4 (N10515, N10511, N6631, N380, N8281);
not NOT1 (N10516, N10513);
nand NAND2 (N10517, N10493, N7267);
xor XOR2 (N10518, N10509, N4492);
or OR4 (N10519, N10494, N8611, N9754, N7957);
and AND4 (N10520, N10486, N10176, N9232, N8424);
and AND3 (N10521, N10516, N1934, N8927);
and AND4 (N10522, N10497, N8248, N9772, N8598);
or OR3 (N10523, N10512, N2356, N2736);
buf BUF1 (N10524, N10518);
nand NAND3 (N10525, N10508, N3332, N9197);
nor NOR4 (N10526, N10519, N2031, N6791, N10051);
nand NAND3 (N10527, N10521, N1837, N9249);
not NOT1 (N10528, N10525);
and AND2 (N10529, N10526, N2917);
nor NOR4 (N10530, N10520, N8928, N6972, N4292);
nand NAND3 (N10531, N10527, N8851, N6200);
not NOT1 (N10532, N10515);
nand NAND4 (N10533, N10529, N8947, N4163, N4307);
or OR2 (N10534, N10532, N5931);
nor NOR2 (N10535, N10528, N3810);
nand NAND3 (N10536, N10517, N2640, N5677);
and AND2 (N10537, N10534, N3264);
nand NAND2 (N10538, N10533, N8743);
nor NOR3 (N10539, N10523, N1623, N2372);
not NOT1 (N10540, N10530);
not NOT1 (N10541, N10540);
and AND2 (N10542, N10541, N8397);
and AND3 (N10543, N10531, N3139, N6077);
and AND2 (N10544, N10524, N5650);
nor NOR4 (N10545, N10542, N3894, N3918, N8855);
and AND3 (N10546, N10545, N4583, N3604);
buf BUF1 (N10547, N10514);
or OR2 (N10548, N10538, N634);
not NOT1 (N10549, N10535);
nand NAND2 (N10550, N10544, N156);
nor NOR3 (N10551, N10539, N4016, N3023);
xor XOR2 (N10552, N10546, N7733);
xor XOR2 (N10553, N10547, N8563);
and AND3 (N10554, N10522, N6488, N7167);
buf BUF1 (N10555, N10536);
xor XOR2 (N10556, N10543, N10402);
or OR2 (N10557, N10551, N3447);
or OR3 (N10558, N10553, N4678, N9168);
not NOT1 (N10559, N10549);
and AND2 (N10560, N10559, N7022);
nand NAND3 (N10561, N10548, N9969, N6214);
nand NAND4 (N10562, N10560, N1715, N439, N8898);
xor XOR2 (N10563, N10537, N2776);
nand NAND4 (N10564, N10555, N9487, N252, N1439);
xor XOR2 (N10565, N10562, N10055);
not NOT1 (N10566, N10557);
not NOT1 (N10567, N10552);
and AND3 (N10568, N10567, N7393, N1974);
or OR4 (N10569, N10550, N385, N7454, N8918);
nand NAND2 (N10570, N10563, N883);
not NOT1 (N10571, N10556);
not NOT1 (N10572, N10565);
nand NAND2 (N10573, N10570, N5849);
nor NOR4 (N10574, N10569, N4335, N9272, N4025);
xor XOR2 (N10575, N10574, N1959);
buf BUF1 (N10576, N10566);
buf BUF1 (N10577, N10561);
buf BUF1 (N10578, N10577);
or OR4 (N10579, N10575, N8707, N2808, N7879);
buf BUF1 (N10580, N10578);
not NOT1 (N10581, N10579);
buf BUF1 (N10582, N10558);
and AND2 (N10583, N10581, N9348);
nand NAND3 (N10584, N10573, N5905, N6846);
and AND4 (N10585, N10572, N2574, N8656, N10131);
xor XOR2 (N10586, N10564, N9779);
buf BUF1 (N10587, N10582);
xor XOR2 (N10588, N10586, N7207);
and AND4 (N10589, N10585, N3881, N9683, N1760);
xor XOR2 (N10590, N10584, N4185);
xor XOR2 (N10591, N10588, N6820);
or OR4 (N10592, N10587, N9189, N3588, N7939);
or OR2 (N10593, N10571, N8635);
or OR3 (N10594, N10554, N6409, N7308);
xor XOR2 (N10595, N10593, N1088);
nor NOR2 (N10596, N10594, N2066);
nor NOR4 (N10597, N10590, N8398, N3570, N1278);
nor NOR4 (N10598, N10595, N7377, N4885, N3344);
xor XOR2 (N10599, N10596, N10369);
not NOT1 (N10600, N10583);
buf BUF1 (N10601, N10591);
and AND3 (N10602, N10592, N9337, N5703);
not NOT1 (N10603, N10601);
not NOT1 (N10604, N10599);
not NOT1 (N10605, N10598);
not NOT1 (N10606, N10568);
and AND4 (N10607, N10606, N8307, N3762, N1288);
and AND3 (N10608, N10597, N10031, N9050);
xor XOR2 (N10609, N10608, N1214);
xor XOR2 (N10610, N10609, N5328);
and AND4 (N10611, N10580, N7270, N5922, N2797);
xor XOR2 (N10612, N10610, N8557);
nor NOR2 (N10613, N10602, N5318);
nor NOR4 (N10614, N10613, N10583, N3644, N4115);
or OR2 (N10615, N10600, N857);
nor NOR2 (N10616, N10589, N8507);
xor XOR2 (N10617, N10605, N6605);
or OR3 (N10618, N10615, N5190, N7957);
xor XOR2 (N10619, N10604, N1712);
nand NAND2 (N10620, N10607, N1147);
nand NAND4 (N10621, N10618, N2503, N10549, N10105);
xor XOR2 (N10622, N10614, N8549);
and AND2 (N10623, N10603, N7565);
and AND3 (N10624, N10620, N4361, N2668);
nor NOR3 (N10625, N10611, N91, N10235);
xor XOR2 (N10626, N10612, N6543);
not NOT1 (N10627, N10617);
not NOT1 (N10628, N10626);
not NOT1 (N10629, N10621);
and AND4 (N10630, N10623, N5012, N8474, N1037);
nor NOR2 (N10631, N10622, N1913);
and AND4 (N10632, N10576, N8169, N2487, N8935);
and AND2 (N10633, N10629, N9651);
nor NOR3 (N10634, N10625, N689, N10031);
nand NAND4 (N10635, N10634, N6231, N7600, N5348);
or OR4 (N10636, N10630, N6791, N5481, N9207);
xor XOR2 (N10637, N10624, N6722);
and AND3 (N10638, N10632, N1656, N439);
nor NOR4 (N10639, N10636, N328, N8056, N10298);
not NOT1 (N10640, N10637);
and AND4 (N10641, N10628, N505, N7063, N3245);
and AND2 (N10642, N10640, N9620);
xor XOR2 (N10643, N10639, N1220);
and AND2 (N10644, N10643, N7622);
buf BUF1 (N10645, N10635);
not NOT1 (N10646, N10627);
nand NAND4 (N10647, N10616, N8770, N7577, N4854);
xor XOR2 (N10648, N10631, N2941);
xor XOR2 (N10649, N10646, N577);
xor XOR2 (N10650, N10619, N3144);
buf BUF1 (N10651, N10645);
xor XOR2 (N10652, N10641, N2149);
buf BUF1 (N10653, N10651);
nor NOR2 (N10654, N10633, N375);
nor NOR2 (N10655, N10653, N9115);
or OR2 (N10656, N10655, N1302);
or OR4 (N10657, N10650, N5073, N7111, N42);
nor NOR2 (N10658, N10652, N6107);
or OR2 (N10659, N10656, N121);
and AND3 (N10660, N10638, N3383, N392);
not NOT1 (N10661, N10642);
or OR4 (N10662, N10654, N5878, N605, N8427);
and AND2 (N10663, N10657, N9798);
and AND3 (N10664, N10660, N8913, N6662);
and AND2 (N10665, N10644, N9542);
buf BUF1 (N10666, N10661);
or OR4 (N10667, N10648, N10069, N1569, N2214);
nand NAND3 (N10668, N10647, N9368, N8102);
xor XOR2 (N10669, N10658, N6254);
nand NAND3 (N10670, N10664, N1422, N988);
or OR2 (N10671, N10659, N2277);
xor XOR2 (N10672, N10665, N1327);
or OR4 (N10673, N10669, N2933, N9871, N2016);
nand NAND2 (N10674, N10649, N6665);
nor NOR2 (N10675, N10673, N6011);
or OR3 (N10676, N10666, N7107, N9581);
xor XOR2 (N10677, N10667, N2904);
and AND3 (N10678, N10668, N7069, N7290);
xor XOR2 (N10679, N10663, N124);
and AND2 (N10680, N10670, N6664);
nand NAND2 (N10681, N10674, N4967);
xor XOR2 (N10682, N10672, N7659);
nor NOR3 (N10683, N10682, N4828, N8674);
and AND2 (N10684, N10680, N9901);
xor XOR2 (N10685, N10675, N4173);
and AND4 (N10686, N10683, N5004, N834, N7683);
not NOT1 (N10687, N10662);
buf BUF1 (N10688, N10684);
and AND4 (N10689, N10681, N185, N4064, N9917);
or OR4 (N10690, N10685, N7915, N4895, N8319);
or OR2 (N10691, N10676, N2331);
not NOT1 (N10692, N10689);
not NOT1 (N10693, N10678);
and AND4 (N10694, N10690, N141, N2301, N4752);
not NOT1 (N10695, N10687);
and AND4 (N10696, N10677, N1655, N7589, N6051);
nand NAND2 (N10697, N10686, N6779);
or OR4 (N10698, N10679, N3202, N5307, N8191);
nor NOR2 (N10699, N10695, N9946);
nand NAND3 (N10700, N10671, N10145, N4593);
nor NOR3 (N10701, N10698, N3794, N7807);
xor XOR2 (N10702, N10691, N2417);
nand NAND4 (N10703, N10699, N376, N3293, N650);
not NOT1 (N10704, N10702);
and AND2 (N10705, N10696, N2893);
and AND4 (N10706, N10688, N10625, N8964, N10496);
buf BUF1 (N10707, N10697);
and AND4 (N10708, N10707, N96, N4174, N6356);
buf BUF1 (N10709, N10700);
xor XOR2 (N10710, N10694, N7675);
or OR2 (N10711, N10706, N3931);
or OR3 (N10712, N10703, N1762, N4083);
and AND4 (N10713, N10708, N8182, N6189, N9860);
buf BUF1 (N10714, N10710);
nor NOR3 (N10715, N10711, N9368, N6790);
and AND4 (N10716, N10701, N9895, N3907, N8673);
nand NAND4 (N10717, N10705, N4268, N3102, N4839);
or OR3 (N10718, N10714, N304, N2493);
nor NOR4 (N10719, N10704, N3468, N2548, N7586);
and AND4 (N10720, N10717, N1700, N2155, N1516);
nand NAND3 (N10721, N10716, N832, N1882);
not NOT1 (N10722, N10713);
buf BUF1 (N10723, N10719);
or OR4 (N10724, N10693, N3175, N8768, N2627);
xor XOR2 (N10725, N10718, N10038);
or OR2 (N10726, N10720, N7657);
buf BUF1 (N10727, N10722);
and AND2 (N10728, N10725, N2368);
nor NOR3 (N10729, N10727, N2323, N9943);
or OR4 (N10730, N10728, N7600, N9430, N5364);
xor XOR2 (N10731, N10721, N9200);
nand NAND4 (N10732, N10709, N2633, N4181, N3046);
or OR2 (N10733, N10715, N822);
buf BUF1 (N10734, N10730);
not NOT1 (N10735, N10733);
nor NOR2 (N10736, N10731, N603);
not NOT1 (N10737, N10723);
xor XOR2 (N10738, N10712, N2817);
nor NOR2 (N10739, N10738, N7321);
buf BUF1 (N10740, N10737);
nor NOR3 (N10741, N10726, N6690, N4158);
buf BUF1 (N10742, N10732);
buf BUF1 (N10743, N10735);
nand NAND4 (N10744, N10739, N2774, N7156, N1799);
buf BUF1 (N10745, N10743);
not NOT1 (N10746, N10741);
not NOT1 (N10747, N10736);
xor XOR2 (N10748, N10747, N134);
xor XOR2 (N10749, N10745, N1206);
nor NOR3 (N10750, N10734, N1482, N5493);
buf BUF1 (N10751, N10724);
nand NAND2 (N10752, N10746, N3439);
buf BUF1 (N10753, N10692);
nor NOR2 (N10754, N10753, N5822);
nor NOR3 (N10755, N10742, N304, N4772);
nor NOR2 (N10756, N10749, N10395);
buf BUF1 (N10757, N10756);
nor NOR2 (N10758, N10744, N7652);
not NOT1 (N10759, N10751);
nor NOR4 (N10760, N10748, N7941, N5520, N2443);
and AND2 (N10761, N10752, N3165);
or OR2 (N10762, N10755, N5975);
and AND3 (N10763, N10758, N327, N1684);
or OR2 (N10764, N10750, N6832);
nor NOR4 (N10765, N10764, N5060, N2637, N5365);
or OR3 (N10766, N10763, N887, N6204);
and AND3 (N10767, N10761, N10561, N1149);
and AND3 (N10768, N10740, N8743, N9233);
buf BUF1 (N10769, N10759);
nor NOR3 (N10770, N10729, N3672, N9801);
or OR3 (N10771, N10765, N5166, N7311);
nor NOR3 (N10772, N10762, N5934, N4165);
nor NOR3 (N10773, N10771, N1033, N519);
not NOT1 (N10774, N10760);
buf BUF1 (N10775, N10768);
buf BUF1 (N10776, N10770);
not NOT1 (N10777, N10767);
and AND4 (N10778, N10766, N3592, N1954, N7085);
and AND4 (N10779, N10769, N4243, N2207, N4347);
xor XOR2 (N10780, N10754, N4711);
nor NOR2 (N10781, N10780, N4373);
nand NAND3 (N10782, N10757, N2637, N518);
buf BUF1 (N10783, N10782);
and AND4 (N10784, N10779, N327, N2599, N8600);
and AND3 (N10785, N10772, N10270, N3547);
nand NAND3 (N10786, N10775, N3806, N5999);
buf BUF1 (N10787, N10776);
buf BUF1 (N10788, N10774);
and AND4 (N10789, N10784, N2299, N7353, N2629);
nor NOR4 (N10790, N10783, N7727, N4690, N889);
buf BUF1 (N10791, N10788);
buf BUF1 (N10792, N10781);
and AND3 (N10793, N10773, N8766, N849);
or OR3 (N10794, N10789, N1812, N4966);
not NOT1 (N10795, N10785);
or OR4 (N10796, N10778, N3215, N5407, N9906);
buf BUF1 (N10797, N10791);
nand NAND2 (N10798, N10793, N6005);
or OR3 (N10799, N10796, N1229, N5737);
not NOT1 (N10800, N10787);
nor NOR3 (N10801, N10790, N9162, N9869);
or OR3 (N10802, N10786, N4168, N6460);
xor XOR2 (N10803, N10794, N5757);
or OR3 (N10804, N10777, N2099, N4139);
nand NAND4 (N10805, N10800, N8086, N6766, N9682);
nor NOR2 (N10806, N10798, N9490);
nor NOR2 (N10807, N10799, N7793);
xor XOR2 (N10808, N10807, N893);
or OR2 (N10809, N10803, N7750);
nand NAND4 (N10810, N10808, N4654, N168, N7803);
buf BUF1 (N10811, N10806);
nand NAND3 (N10812, N10809, N2617, N5724);
xor XOR2 (N10813, N10810, N1865);
nand NAND3 (N10814, N10812, N3139, N9390);
nand NAND3 (N10815, N10805, N5704, N8551);
or OR4 (N10816, N10815, N3171, N9013, N281);
nand NAND4 (N10817, N10804, N2804, N1643, N4842);
nand NAND4 (N10818, N10813, N7476, N10327, N4017);
and AND4 (N10819, N10797, N2822, N90, N1735);
not NOT1 (N10820, N10814);
buf BUF1 (N10821, N10818);
nor NOR3 (N10822, N10792, N10265, N8317);
nor NOR4 (N10823, N10816, N4818, N6479, N1315);
and AND3 (N10824, N10801, N1375, N3193);
nor NOR3 (N10825, N10795, N2379, N2634);
nand NAND4 (N10826, N10817, N2824, N6827, N1058);
nand NAND4 (N10827, N10825, N2711, N8610, N5058);
and AND4 (N10828, N10826, N650, N1753, N3001);
xor XOR2 (N10829, N10827, N8841);
not NOT1 (N10830, N10828);
buf BUF1 (N10831, N10824);
or OR3 (N10832, N10821, N10704, N104);
or OR2 (N10833, N10820, N4674);
nor NOR4 (N10834, N10829, N2017, N6321, N553);
nand NAND4 (N10835, N10830, N6955, N4667, N1288);
buf BUF1 (N10836, N10833);
and AND3 (N10837, N10832, N4785, N7409);
or OR3 (N10838, N10802, N8234, N10777);
nand NAND4 (N10839, N10823, N2572, N7411, N2687);
buf BUF1 (N10840, N10836);
nand NAND4 (N10841, N10831, N4842, N8343, N7640);
nand NAND3 (N10842, N10811, N7723, N3225);
not NOT1 (N10843, N10840);
or OR4 (N10844, N10839, N4939, N7911, N10188);
nor NOR4 (N10845, N10822, N9306, N9916, N9081);
not NOT1 (N10846, N10844);
not NOT1 (N10847, N10842);
and AND4 (N10848, N10838, N5011, N10373, N6414);
or OR2 (N10849, N10819, N5841);
nand NAND3 (N10850, N10834, N3450, N4695);
nor NOR3 (N10851, N10841, N1482, N10542);
or OR3 (N10852, N10851, N8094, N10222);
nand NAND4 (N10853, N10843, N10352, N10629, N5899);
nand NAND4 (N10854, N10847, N2589, N398, N1633);
nor NOR4 (N10855, N10849, N516, N10047, N3567);
buf BUF1 (N10856, N10835);
not NOT1 (N10857, N10852);
not NOT1 (N10858, N10853);
or OR2 (N10859, N10858, N5901);
buf BUF1 (N10860, N10845);
or OR4 (N10861, N10846, N4137, N5995, N7988);
not NOT1 (N10862, N10856);
buf BUF1 (N10863, N10855);
buf BUF1 (N10864, N10857);
not NOT1 (N10865, N10837);
buf BUF1 (N10866, N10860);
or OR3 (N10867, N10854, N5570, N3815);
and AND4 (N10868, N10848, N2308, N8783, N470);
not NOT1 (N10869, N10864);
not NOT1 (N10870, N10866);
and AND4 (N10871, N10861, N294, N2091, N1372);
or OR3 (N10872, N10871, N3688, N7696);
not NOT1 (N10873, N10867);
or OR4 (N10874, N10850, N1182, N3592, N4329);
xor XOR2 (N10875, N10862, N9749);
xor XOR2 (N10876, N10870, N8950);
nor NOR4 (N10877, N10863, N7950, N1439, N2486);
not NOT1 (N10878, N10869);
or OR3 (N10879, N10868, N5707, N519);
nand NAND4 (N10880, N10873, N8380, N3522, N2516);
or OR4 (N10881, N10876, N5509, N2609, N5155);
nor NOR4 (N10882, N10881, N8961, N7739, N10493);
nand NAND2 (N10883, N10879, N5409);
and AND2 (N10884, N10865, N6181);
nor NOR4 (N10885, N10878, N8754, N9221, N7950);
nor NOR3 (N10886, N10872, N5301, N10744);
nand NAND2 (N10887, N10874, N6121);
or OR3 (N10888, N10859, N9195, N4486);
xor XOR2 (N10889, N10888, N1174);
or OR3 (N10890, N10886, N4149, N6275);
nand NAND4 (N10891, N10882, N6980, N5611, N795);
nand NAND4 (N10892, N10875, N848, N5071, N9506);
nand NAND3 (N10893, N10891, N2135, N7731);
and AND4 (N10894, N10884, N3266, N6879, N251);
nor NOR3 (N10895, N10880, N1363, N601);
or OR4 (N10896, N10892, N4938, N1524, N9770);
or OR3 (N10897, N10895, N4547, N9284);
buf BUF1 (N10898, N10890);
and AND3 (N10899, N10885, N10499, N10882);
buf BUF1 (N10900, N10893);
or OR3 (N10901, N10900, N6682, N337);
or OR2 (N10902, N10889, N9443);
and AND2 (N10903, N10899, N7620);
nand NAND3 (N10904, N10897, N8285, N7203);
nand NAND4 (N10905, N10903, N9988, N4893, N4001);
xor XOR2 (N10906, N10898, N7226);
nand NAND2 (N10907, N10901, N9271);
buf BUF1 (N10908, N10906);
nand NAND4 (N10909, N10883, N4319, N6702, N7669);
not NOT1 (N10910, N10894);
nand NAND2 (N10911, N10907, N2979);
not NOT1 (N10912, N10909);
xor XOR2 (N10913, N10910, N6891);
nand NAND3 (N10914, N10913, N2186, N2235);
nand NAND4 (N10915, N10887, N4398, N4082, N794);
nand NAND2 (N10916, N10905, N5307);
nand NAND3 (N10917, N10916, N6274, N3046);
buf BUF1 (N10918, N10917);
nand NAND4 (N10919, N10904, N10185, N6199, N2615);
not NOT1 (N10920, N10908);
and AND4 (N10921, N10911, N1718, N10181, N9603);
nor NOR2 (N10922, N10915, N2124);
nor NOR4 (N10923, N10902, N1246, N7951, N5565);
not NOT1 (N10924, N10923);
nor NOR3 (N10925, N10877, N4816, N2720);
xor XOR2 (N10926, N10912, N5863);
or OR4 (N10927, N10925, N7661, N640, N3655);
or OR3 (N10928, N10921, N5803, N9477);
xor XOR2 (N10929, N10896, N10461);
buf BUF1 (N10930, N10922);
and AND4 (N10931, N10929, N3522, N4804, N6757);
and AND4 (N10932, N10927, N6205, N8104, N6555);
not NOT1 (N10933, N10926);
not NOT1 (N10934, N10924);
nor NOR4 (N10935, N10928, N3480, N1571, N7017);
or OR2 (N10936, N10933, N4474);
and AND3 (N10937, N10919, N8172, N8614);
or OR2 (N10938, N10931, N6708);
xor XOR2 (N10939, N10918, N6332);
xor XOR2 (N10940, N10935, N10834);
or OR4 (N10941, N10934, N1481, N1164, N5692);
xor XOR2 (N10942, N10937, N6158);
nand NAND4 (N10943, N10941, N8689, N4659, N1514);
buf BUF1 (N10944, N10943);
buf BUF1 (N10945, N10944);
or OR4 (N10946, N10942, N7555, N2445, N832);
xor XOR2 (N10947, N10939, N7690);
nor NOR3 (N10948, N10938, N4575, N1346);
xor XOR2 (N10949, N10914, N8741);
and AND3 (N10950, N10932, N3188, N2224);
buf BUF1 (N10951, N10930);
not NOT1 (N10952, N10951);
and AND3 (N10953, N10946, N8565, N4073);
nand NAND3 (N10954, N10948, N5645, N4733);
xor XOR2 (N10955, N10952, N3306);
not NOT1 (N10956, N10949);
buf BUF1 (N10957, N10956);
buf BUF1 (N10958, N10940);
or OR3 (N10959, N10957, N2184, N4080);
buf BUF1 (N10960, N10958);
and AND4 (N10961, N10950, N1648, N9585, N3827);
buf BUF1 (N10962, N10947);
nand NAND2 (N10963, N10920, N403);
and AND2 (N10964, N10955, N7985);
buf BUF1 (N10965, N10963);
nand NAND4 (N10966, N10960, N4326, N2899, N1212);
and AND4 (N10967, N10959, N7202, N5602, N832);
nand NAND2 (N10968, N10962, N7854);
or OR4 (N10969, N10954, N9360, N10685, N7206);
or OR3 (N10970, N10965, N5163, N246);
nand NAND3 (N10971, N10969, N10441, N2832);
nand NAND3 (N10972, N10936, N1619, N10086);
nand NAND3 (N10973, N10945, N5035, N5765);
nor NOR3 (N10974, N10970, N2600, N8661);
and AND2 (N10975, N10971, N7124);
or OR4 (N10976, N10966, N9702, N4024, N261);
or OR4 (N10977, N10973, N22, N4752, N237);
buf BUF1 (N10978, N10964);
nand NAND2 (N10979, N10961, N5343);
xor XOR2 (N10980, N10976, N5741);
not NOT1 (N10981, N10975);
and AND4 (N10982, N10980, N473, N337, N8362);
or OR2 (N10983, N10953, N5100);
and AND3 (N10984, N10968, N3582, N8126);
and AND4 (N10985, N10982, N8058, N585, N1617);
and AND2 (N10986, N10985, N9340);
not NOT1 (N10987, N10977);
not NOT1 (N10988, N10978);
xor XOR2 (N10989, N10988, N10410);
xor XOR2 (N10990, N10989, N9718);
xor XOR2 (N10991, N10974, N7788);
or OR2 (N10992, N10972, N1797);
nor NOR4 (N10993, N10984, N3675, N1093, N769);
xor XOR2 (N10994, N10990, N6812);
not NOT1 (N10995, N10994);
nand NAND2 (N10996, N10993, N10134);
nor NOR3 (N10997, N10986, N7498, N1386);
and AND4 (N10998, N10996, N3527, N7638, N1836);
nand NAND4 (N10999, N10983, N3744, N5870, N10379);
nand NAND4 (N11000, N10995, N5354, N9739, N5675);
xor XOR2 (N11001, N10987, N3447);
nor NOR4 (N11002, N11001, N8296, N2108, N4038);
buf BUF1 (N11003, N11002);
nand NAND2 (N11004, N10981, N8284);
not NOT1 (N11005, N11003);
and AND3 (N11006, N11004, N723, N8036);
buf BUF1 (N11007, N11000);
or OR2 (N11008, N11005, N9754);
xor XOR2 (N11009, N10992, N497);
xor XOR2 (N11010, N10991, N1132);
nor NOR4 (N11011, N11006, N10533, N6149, N5808);
or OR2 (N11012, N11010, N9365);
xor XOR2 (N11013, N11009, N6366);
and AND2 (N11014, N11013, N3992);
not NOT1 (N11015, N10998);
buf BUF1 (N11016, N10967);
buf BUF1 (N11017, N10979);
xor XOR2 (N11018, N11007, N5269);
not NOT1 (N11019, N11017);
or OR2 (N11020, N11012, N2173);
xor XOR2 (N11021, N11011, N1313);
nor NOR2 (N11022, N11021, N2959);
not NOT1 (N11023, N11019);
nor NOR4 (N11024, N11018, N2579, N10377, N855);
xor XOR2 (N11025, N11015, N199);
not NOT1 (N11026, N11023);
and AND4 (N11027, N10999, N2215, N6566, N9004);
and AND3 (N11028, N11008, N9036, N6677);
or OR3 (N11029, N11024, N9522, N2706);
and AND3 (N11030, N11026, N6641, N9006);
or OR3 (N11031, N11027, N5921, N5914);
nor NOR3 (N11032, N11022, N2209, N5464);
nor NOR2 (N11033, N11014, N8231);
nor NOR2 (N11034, N11032, N2762);
buf BUF1 (N11035, N11029);
or OR2 (N11036, N11030, N6569);
nor NOR2 (N11037, N11016, N5877);
not NOT1 (N11038, N11034);
and AND4 (N11039, N11031, N2146, N6490, N8367);
nand NAND2 (N11040, N11037, N10597);
xor XOR2 (N11041, N11020, N7009);
or OR4 (N11042, N11039, N1984, N9232, N566);
nor NOR4 (N11043, N11038, N543, N5306, N7615);
or OR2 (N11044, N11043, N968);
and AND2 (N11045, N11028, N3610);
xor XOR2 (N11046, N11045, N1635);
nand NAND4 (N11047, N11033, N2277, N2488, N9472);
nor NOR4 (N11048, N10997, N8823, N8838, N3866);
buf BUF1 (N11049, N11036);
and AND3 (N11050, N11041, N8051, N8849);
xor XOR2 (N11051, N11042, N9849);
not NOT1 (N11052, N11047);
nor NOR2 (N11053, N11035, N10072);
nand NAND4 (N11054, N11051, N10045, N5589, N8771);
or OR2 (N11055, N11044, N8768);
buf BUF1 (N11056, N11025);
and AND2 (N11057, N11048, N6897);
nand NAND3 (N11058, N11046, N7004, N8709);
or OR3 (N11059, N11056, N9899, N2972);
xor XOR2 (N11060, N11058, N7535);
nor NOR3 (N11061, N11057, N6233, N4960);
or OR4 (N11062, N11061, N4737, N5546, N2612);
buf BUF1 (N11063, N11055);
buf BUF1 (N11064, N11060);
nor NOR3 (N11065, N11050, N9384, N767);
not NOT1 (N11066, N11064);
not NOT1 (N11067, N11052);
and AND2 (N11068, N11059, N2716);
and AND4 (N11069, N11066, N8950, N3871, N9233);
nor NOR2 (N11070, N11063, N506);
nor NOR2 (N11071, N11062, N89);
not NOT1 (N11072, N11054);
or OR3 (N11073, N11049, N2328, N7278);
and AND4 (N11074, N11065, N5142, N6944, N5295);
and AND3 (N11075, N11068, N6434, N1719);
nor NOR2 (N11076, N11053, N826);
nor NOR4 (N11077, N11076, N2498, N6560, N9562);
xor XOR2 (N11078, N11074, N4257);
xor XOR2 (N11079, N11072, N2459);
not NOT1 (N11080, N11067);
buf BUF1 (N11081, N11070);
and AND2 (N11082, N11069, N7343);
not NOT1 (N11083, N11081);
and AND4 (N11084, N11075, N2356, N8981, N5658);
nand NAND3 (N11085, N11040, N549, N1900);
or OR2 (N11086, N11077, N95);
buf BUF1 (N11087, N11082);
or OR4 (N11088, N11083, N5911, N2421, N1456);
not NOT1 (N11089, N11071);
and AND4 (N11090, N11086, N4521, N5203, N4753);
not NOT1 (N11091, N11085);
buf BUF1 (N11092, N11080);
or OR2 (N11093, N11090, N2163);
or OR2 (N11094, N11087, N5263);
and AND2 (N11095, N11093, N7554);
buf BUF1 (N11096, N11095);
nor NOR3 (N11097, N11079, N7714, N5077);
nor NOR2 (N11098, N11091, N2469);
buf BUF1 (N11099, N11084);
nor NOR4 (N11100, N11089, N9428, N4894, N6461);
not NOT1 (N11101, N11096);
or OR2 (N11102, N11073, N9888);
nor NOR4 (N11103, N11100, N4485, N10057, N10694);
nor NOR2 (N11104, N11099, N6848);
nand NAND2 (N11105, N11098, N6993);
or OR4 (N11106, N11102, N5041, N1023, N1762);
nor NOR2 (N11107, N11103, N4178);
nor NOR4 (N11108, N11097, N671, N3294, N10571);
or OR4 (N11109, N11108, N9994, N8309, N10115);
buf BUF1 (N11110, N11104);
or OR2 (N11111, N11092, N8133);
or OR4 (N11112, N11101, N9914, N7650, N1643);
buf BUF1 (N11113, N11106);
buf BUF1 (N11114, N11107);
buf BUF1 (N11115, N11111);
or OR2 (N11116, N11113, N5194);
and AND4 (N11117, N11088, N8537, N7165, N3438);
nand NAND3 (N11118, N11094, N5761, N2177);
nand NAND3 (N11119, N11116, N6498, N766);
or OR4 (N11120, N11105, N4171, N442, N4803);
not NOT1 (N11121, N11112);
buf BUF1 (N11122, N11109);
xor XOR2 (N11123, N11115, N10734);
nor NOR3 (N11124, N11117, N4693, N3148);
or OR4 (N11125, N11114, N6449, N189, N4388);
and AND3 (N11126, N11125, N3330, N6849);
or OR2 (N11127, N11119, N2062);
nand NAND2 (N11128, N11122, N10521);
nand NAND2 (N11129, N11118, N9984);
nand NAND2 (N11130, N11078, N7140);
and AND4 (N11131, N11126, N4977, N8531, N1322);
nor NOR2 (N11132, N11131, N1148);
nand NAND2 (N11133, N11132, N6216);
or OR2 (N11134, N11120, N10499);
nand NAND2 (N11135, N11128, N9328);
nand NAND4 (N11136, N11134, N11094, N5222, N1673);
xor XOR2 (N11137, N11135, N2046);
nor NOR3 (N11138, N11137, N4642, N10496);
xor XOR2 (N11139, N11124, N9363);
nor NOR4 (N11140, N11129, N9368, N6358, N6443);
not NOT1 (N11141, N11138);
and AND4 (N11142, N11123, N7396, N5373, N703);
or OR4 (N11143, N11130, N7644, N8542, N2077);
and AND3 (N11144, N11133, N7503, N6860);
not NOT1 (N11145, N11121);
and AND3 (N11146, N11141, N9346, N8297);
nand NAND3 (N11147, N11146, N4835, N2607);
not NOT1 (N11148, N11147);
nor NOR4 (N11149, N11110, N574, N3404, N6295);
nand NAND2 (N11150, N11143, N8910);
buf BUF1 (N11151, N11142);
nor NOR3 (N11152, N11148, N9196, N8128);
and AND2 (N11153, N11145, N2863);
xor XOR2 (N11154, N11149, N3460);
or OR3 (N11155, N11150, N7986, N6445);
nor NOR2 (N11156, N11153, N2907);
or OR3 (N11157, N11156, N9059, N4551);
nand NAND3 (N11158, N11136, N3650, N6196);
or OR2 (N11159, N11154, N7563);
and AND3 (N11160, N11155, N9026, N5822);
or OR4 (N11161, N11152, N4941, N2561, N5081);
not NOT1 (N11162, N11127);
or OR3 (N11163, N11160, N9803, N7753);
and AND3 (N11164, N11139, N4657, N10662);
nor NOR4 (N11165, N11161, N3949, N4330, N6220);
not NOT1 (N11166, N11157);
nor NOR4 (N11167, N11158, N1314, N10332, N4789);
nor NOR2 (N11168, N11167, N7189);
and AND2 (N11169, N11165, N10056);
and AND3 (N11170, N11140, N1317, N4749);
not NOT1 (N11171, N11163);
nand NAND2 (N11172, N11171, N9173);
nor NOR4 (N11173, N11159, N11043, N1735, N8159);
and AND4 (N11174, N11162, N8920, N905, N8918);
and AND2 (N11175, N11144, N3818);
not NOT1 (N11176, N11175);
xor XOR2 (N11177, N11173, N1164);
nand NAND4 (N11178, N11168, N802, N8920, N5149);
not NOT1 (N11179, N11174);
nor NOR4 (N11180, N11178, N3945, N6573, N3227);
buf BUF1 (N11181, N11166);
and AND2 (N11182, N11169, N3985);
or OR2 (N11183, N11182, N8245);
or OR3 (N11184, N11170, N4873, N10396);
not NOT1 (N11185, N11151);
or OR2 (N11186, N11164, N9183);
xor XOR2 (N11187, N11176, N9400);
nor NOR4 (N11188, N11185, N2461, N5111, N4733);
not NOT1 (N11189, N11188);
and AND3 (N11190, N11183, N7890, N6492);
xor XOR2 (N11191, N11190, N5363);
not NOT1 (N11192, N11191);
buf BUF1 (N11193, N11186);
not NOT1 (N11194, N11192);
nor NOR3 (N11195, N11181, N9507, N1328);
and AND3 (N11196, N11172, N11072, N1312);
buf BUF1 (N11197, N11195);
or OR3 (N11198, N11180, N254, N9626);
buf BUF1 (N11199, N11193);
xor XOR2 (N11200, N11177, N8162);
or OR3 (N11201, N11189, N2723, N9446);
or OR4 (N11202, N11197, N10251, N6985, N3761);
and AND3 (N11203, N11199, N4265, N5379);
and AND4 (N11204, N11196, N9541, N470, N6481);
or OR3 (N11205, N11198, N6948, N8786);
xor XOR2 (N11206, N11202, N3295);
nor NOR4 (N11207, N11179, N6005, N2971, N6806);
not NOT1 (N11208, N11206);
xor XOR2 (N11209, N11200, N3484);
buf BUF1 (N11210, N11208);
or OR3 (N11211, N11209, N3441, N5661);
nor NOR3 (N11212, N11205, N1731, N4453);
nor NOR2 (N11213, N11204, N1423);
buf BUF1 (N11214, N11210);
and AND4 (N11215, N11194, N3285, N658, N6240);
nand NAND4 (N11216, N11187, N4262, N10760, N5390);
xor XOR2 (N11217, N11214, N3396);
nand NAND4 (N11218, N11211, N1201, N9450, N7296);
or OR3 (N11219, N11218, N8423, N9005);
nor NOR4 (N11220, N11201, N4919, N4376, N7521);
not NOT1 (N11221, N11219);
buf BUF1 (N11222, N11184);
buf BUF1 (N11223, N11221);
nor NOR3 (N11224, N11212, N6080, N7742);
and AND2 (N11225, N11213, N8473);
buf BUF1 (N11226, N11217);
and AND4 (N11227, N11226, N9037, N5733, N10333);
not NOT1 (N11228, N11224);
not NOT1 (N11229, N11216);
nand NAND4 (N11230, N11223, N2805, N2586, N10842);
nor NOR2 (N11231, N11227, N6602);
or OR3 (N11232, N11230, N7380, N1605);
nor NOR2 (N11233, N11228, N6796);
nand NAND3 (N11234, N11231, N1749, N5520);
xor XOR2 (N11235, N11215, N1466);
nand NAND2 (N11236, N11229, N8916);
and AND4 (N11237, N11222, N6161, N5087, N1869);
or OR4 (N11238, N11233, N9380, N8635, N3219);
not NOT1 (N11239, N11225);
xor XOR2 (N11240, N11232, N3880);
not NOT1 (N11241, N11240);
not NOT1 (N11242, N11235);
xor XOR2 (N11243, N11203, N7742);
buf BUF1 (N11244, N11220);
not NOT1 (N11245, N11244);
or OR4 (N11246, N11241, N5715, N6618, N1779);
xor XOR2 (N11247, N11234, N5129);
not NOT1 (N11248, N11245);
buf BUF1 (N11249, N11207);
or OR4 (N11250, N11237, N5500, N10361, N5498);
buf BUF1 (N11251, N11236);
xor XOR2 (N11252, N11248, N10738);
not NOT1 (N11253, N11238);
nand NAND3 (N11254, N11253, N2878, N6401);
xor XOR2 (N11255, N11250, N3957);
buf BUF1 (N11256, N11255);
or OR4 (N11257, N11256, N1752, N2598, N9741);
buf BUF1 (N11258, N11249);
xor XOR2 (N11259, N11252, N3758);
xor XOR2 (N11260, N11257, N5926);
nor NOR3 (N11261, N11243, N6955, N5745);
nor NOR3 (N11262, N11254, N1753, N5197);
or OR3 (N11263, N11251, N7629, N148);
buf BUF1 (N11264, N11259);
nor NOR2 (N11265, N11264, N5893);
or OR3 (N11266, N11263, N7118, N3607);
xor XOR2 (N11267, N11247, N7395);
nand NAND4 (N11268, N11246, N9957, N2915, N9802);
and AND2 (N11269, N11262, N2925);
and AND3 (N11270, N11267, N6622, N553);
buf BUF1 (N11271, N11270);
and AND2 (N11272, N11266, N95);
nor NOR4 (N11273, N11269, N9075, N2559, N4527);
or OR2 (N11274, N11273, N3284);
buf BUF1 (N11275, N11258);
and AND4 (N11276, N11261, N1120, N3801, N3976);
or OR4 (N11277, N11275, N5143, N3499, N10609);
and AND4 (N11278, N11239, N1456, N8246, N9380);
not NOT1 (N11279, N11265);
xor XOR2 (N11280, N11277, N10624);
not NOT1 (N11281, N11276);
xor XOR2 (N11282, N11271, N4072);
nor NOR4 (N11283, N11260, N5674, N9370, N3921);
or OR4 (N11284, N11279, N2189, N1370, N4184);
and AND2 (N11285, N11268, N499);
not NOT1 (N11286, N11272);
xor XOR2 (N11287, N11281, N1545);
nor NOR4 (N11288, N11285, N1415, N5421, N8398);
xor XOR2 (N11289, N11278, N8064);
buf BUF1 (N11290, N11287);
or OR2 (N11291, N11284, N3175);
xor XOR2 (N11292, N11280, N1400);
not NOT1 (N11293, N11274);
nor NOR3 (N11294, N11293, N900, N6613);
xor XOR2 (N11295, N11288, N3191);
or OR3 (N11296, N11294, N1359, N7312);
nor NOR3 (N11297, N11289, N5216, N11257);
nor NOR3 (N11298, N11297, N6188, N1961);
or OR2 (N11299, N11290, N6925);
not NOT1 (N11300, N11295);
xor XOR2 (N11301, N11300, N534);
buf BUF1 (N11302, N11282);
nor NOR4 (N11303, N11286, N6006, N10501, N8449);
or OR3 (N11304, N11292, N2709, N8114);
or OR3 (N11305, N11298, N2022, N3815);
xor XOR2 (N11306, N11242, N689);
xor XOR2 (N11307, N11306, N5355);
buf BUF1 (N11308, N11291);
not NOT1 (N11309, N11301);
and AND3 (N11310, N11308, N9572, N777);
nor NOR3 (N11311, N11303, N5682, N8485);
buf BUF1 (N11312, N11283);
and AND2 (N11313, N11299, N6962);
not NOT1 (N11314, N11302);
buf BUF1 (N11315, N11313);
xor XOR2 (N11316, N11314, N1997);
nand NAND4 (N11317, N11307, N1359, N3300, N10385);
nand NAND2 (N11318, N11312, N2580);
or OR3 (N11319, N11311, N9399, N9575);
or OR4 (N11320, N11316, N6560, N8790, N9858);
buf BUF1 (N11321, N11317);
buf BUF1 (N11322, N11315);
and AND3 (N11323, N11304, N9270, N7435);
and AND3 (N11324, N11320, N3875, N10649);
and AND3 (N11325, N11321, N11106, N123);
and AND3 (N11326, N11318, N5746, N8453);
buf BUF1 (N11327, N11319);
nand NAND3 (N11328, N11327, N2503, N8190);
buf BUF1 (N11329, N11323);
and AND4 (N11330, N11305, N5206, N3214, N7401);
nand NAND2 (N11331, N11326, N1062);
not NOT1 (N11332, N11324);
not NOT1 (N11333, N11309);
or OR4 (N11334, N11329, N6795, N9583, N6667);
xor XOR2 (N11335, N11331, N6151);
buf BUF1 (N11336, N11335);
nand NAND3 (N11337, N11322, N824, N6518);
nor NOR4 (N11338, N11333, N1616, N7243, N8211);
nor NOR4 (N11339, N11336, N8217, N7158, N5789);
xor XOR2 (N11340, N11338, N9959);
or OR4 (N11341, N11310, N8120, N1270, N1441);
nand NAND3 (N11342, N11334, N10316, N3255);
or OR4 (N11343, N11296, N1177, N11219, N7507);
nor NOR4 (N11344, N11332, N6694, N8577, N7542);
buf BUF1 (N11345, N11337);
xor XOR2 (N11346, N11330, N11043);
and AND3 (N11347, N11343, N7332, N2093);
nor NOR2 (N11348, N11325, N8902);
nand NAND3 (N11349, N11348, N11204, N3318);
nand NAND3 (N11350, N11340, N4779, N3905);
buf BUF1 (N11351, N11342);
nor NOR2 (N11352, N11349, N10395);
buf BUF1 (N11353, N11341);
buf BUF1 (N11354, N11352);
nor NOR4 (N11355, N11345, N11231, N5748, N7417);
or OR4 (N11356, N11328, N6465, N10401, N2685);
or OR3 (N11357, N11356, N9731, N2897);
or OR4 (N11358, N11344, N1920, N9315, N2442);
buf BUF1 (N11359, N11353);
buf BUF1 (N11360, N11339);
and AND2 (N11361, N11346, N7090);
nand NAND2 (N11362, N11347, N9684);
buf BUF1 (N11363, N11357);
not NOT1 (N11364, N11362);
nor NOR3 (N11365, N11358, N10635, N9621);
not NOT1 (N11366, N11360);
nand NAND4 (N11367, N11355, N4473, N2227, N7585);
and AND3 (N11368, N11359, N7472, N6631);
xor XOR2 (N11369, N11367, N2776);
buf BUF1 (N11370, N11351);
not NOT1 (N11371, N11368);
nand NAND2 (N11372, N11371, N8666);
not NOT1 (N11373, N11372);
not NOT1 (N11374, N11361);
not NOT1 (N11375, N11369);
or OR4 (N11376, N11364, N5958, N7972, N2136);
nand NAND4 (N11377, N11354, N6218, N2939, N6399);
not NOT1 (N11378, N11350);
not NOT1 (N11379, N11363);
or OR4 (N11380, N11376, N7352, N1723, N7280);
not NOT1 (N11381, N11379);
and AND2 (N11382, N11377, N7744);
nor NOR4 (N11383, N11374, N8170, N10330, N10928);
or OR2 (N11384, N11370, N6849);
nand NAND3 (N11385, N11381, N7485, N2566);
nor NOR2 (N11386, N11382, N11331);
or OR4 (N11387, N11386, N5139, N845, N5410);
not NOT1 (N11388, N11373);
buf BUF1 (N11389, N11366);
buf BUF1 (N11390, N11385);
xor XOR2 (N11391, N11378, N3914);
nor NOR3 (N11392, N11384, N8946, N3152);
nor NOR4 (N11393, N11390, N2778, N6158, N1250);
or OR3 (N11394, N11393, N11066, N8509);
not NOT1 (N11395, N11365);
not NOT1 (N11396, N11388);
buf BUF1 (N11397, N11394);
buf BUF1 (N11398, N11380);
or OR4 (N11399, N11395, N276, N83, N2463);
or OR3 (N11400, N11398, N256, N11219);
nand NAND3 (N11401, N11383, N8107, N7181);
nor NOR4 (N11402, N11391, N10540, N3195, N1159);
or OR4 (N11403, N11402, N10556, N2208, N9417);
xor XOR2 (N11404, N11403, N2375);
nor NOR4 (N11405, N11397, N6082, N11084, N5820);
xor XOR2 (N11406, N11396, N6668);
xor XOR2 (N11407, N11406, N3560);
buf BUF1 (N11408, N11389);
not NOT1 (N11409, N11405);
nand NAND3 (N11410, N11392, N7783, N4841);
nor NOR4 (N11411, N11375, N1738, N1482, N967);
buf BUF1 (N11412, N11409);
xor XOR2 (N11413, N11404, N11189);
not NOT1 (N11414, N11401);
and AND4 (N11415, N11407, N3284, N7787, N579);
nand NAND2 (N11416, N11415, N5869);
xor XOR2 (N11417, N11412, N1174);
xor XOR2 (N11418, N11410, N2816);
buf BUF1 (N11419, N11387);
or OR3 (N11420, N11399, N3074, N8680);
buf BUF1 (N11421, N11420);
not NOT1 (N11422, N11413);
not NOT1 (N11423, N11408);
not NOT1 (N11424, N11422);
not NOT1 (N11425, N11421);
or OR3 (N11426, N11416, N843, N933);
nor NOR3 (N11427, N11424, N7836, N1515);
not NOT1 (N11428, N11417);
or OR2 (N11429, N11425, N7068);
or OR4 (N11430, N11429, N782, N10024, N1021);
xor XOR2 (N11431, N11418, N10578);
not NOT1 (N11432, N11426);
xor XOR2 (N11433, N11411, N3692);
not NOT1 (N11434, N11400);
and AND2 (N11435, N11419, N1745);
xor XOR2 (N11436, N11431, N5626);
not NOT1 (N11437, N11433);
or OR2 (N11438, N11434, N4111);
nor NOR3 (N11439, N11435, N2955, N989);
nor NOR2 (N11440, N11439, N10581);
or OR3 (N11441, N11438, N3875, N5599);
not NOT1 (N11442, N11430);
and AND3 (N11443, N11428, N7775, N4296);
or OR3 (N11444, N11423, N6064, N1874);
and AND4 (N11445, N11441, N8992, N33, N1021);
xor XOR2 (N11446, N11440, N5103);
nand NAND2 (N11447, N11446, N887);
nor NOR4 (N11448, N11427, N5881, N5368, N4577);
or OR4 (N11449, N11414, N6298, N6091, N2257);
or OR3 (N11450, N11443, N9224, N4287);
buf BUF1 (N11451, N11436);
not NOT1 (N11452, N11445);
nor NOR3 (N11453, N11448, N8678, N3739);
nand NAND3 (N11454, N11447, N3127, N3598);
buf BUF1 (N11455, N11454);
xor XOR2 (N11456, N11444, N9822);
buf BUF1 (N11457, N11452);
nor NOR3 (N11458, N11455, N340, N4131);
nor NOR2 (N11459, N11458, N670);
xor XOR2 (N11460, N11456, N1690);
nor NOR3 (N11461, N11437, N3283, N5643);
nor NOR4 (N11462, N11449, N5845, N4901, N75);
and AND2 (N11463, N11450, N1450);
nor NOR4 (N11464, N11461, N9341, N2122, N9448);
or OR2 (N11465, N11432, N3123);
nand NAND2 (N11466, N11451, N11121);
and AND3 (N11467, N11464, N6398, N7297);
xor XOR2 (N11468, N11457, N11330);
not NOT1 (N11469, N11460);
buf BUF1 (N11470, N11463);
nor NOR2 (N11471, N11466, N3794);
nand NAND4 (N11472, N11469, N9568, N10147, N6145);
nand NAND3 (N11473, N11471, N10683, N1337);
nor NOR3 (N11474, N11473, N7481, N8999);
not NOT1 (N11475, N11459);
and AND3 (N11476, N11453, N8587, N1348);
nor NOR4 (N11477, N11465, N2549, N4814, N8266);
not NOT1 (N11478, N11468);
or OR3 (N11479, N11475, N9433, N8289);
nand NAND3 (N11480, N11472, N9335, N1700);
or OR3 (N11481, N11470, N2290, N4951);
buf BUF1 (N11482, N11467);
buf BUF1 (N11483, N11462);
xor XOR2 (N11484, N11482, N3144);
nand NAND4 (N11485, N11481, N9723, N6715, N1234);
buf BUF1 (N11486, N11485);
or OR4 (N11487, N11483, N8106, N8627, N9485);
nand NAND2 (N11488, N11487, N5647);
and AND2 (N11489, N11486, N9244);
and AND4 (N11490, N11477, N7148, N1586, N4022);
xor XOR2 (N11491, N11480, N9800);
or OR2 (N11492, N11479, N6966);
nand NAND4 (N11493, N11478, N5251, N1306, N11363);
not NOT1 (N11494, N11492);
nor NOR2 (N11495, N11493, N7320);
nor NOR2 (N11496, N11474, N3434);
nand NAND2 (N11497, N11496, N5974);
not NOT1 (N11498, N11497);
buf BUF1 (N11499, N11484);
not NOT1 (N11500, N11488);
xor XOR2 (N11501, N11499, N9093);
and AND3 (N11502, N11442, N5914, N9242);
not NOT1 (N11503, N11498);
not NOT1 (N11504, N11495);
and AND3 (N11505, N11476, N11090, N9489);
nor NOR4 (N11506, N11502, N2242, N5422, N255);
nand NAND2 (N11507, N11505, N1349);
xor XOR2 (N11508, N11506, N4517);
xor XOR2 (N11509, N11508, N6671);
buf BUF1 (N11510, N11503);
nand NAND3 (N11511, N11489, N1037, N6487);
xor XOR2 (N11512, N11501, N8918);
buf BUF1 (N11513, N11491);
or OR2 (N11514, N11513, N11361);
buf BUF1 (N11515, N11494);
nor NOR4 (N11516, N11514, N1474, N5056, N5933);
xor XOR2 (N11517, N11510, N7211);
nor NOR3 (N11518, N11504, N2308, N8948);
and AND2 (N11519, N11518, N8850);
or OR4 (N11520, N11490, N7179, N8198, N394);
nor NOR4 (N11521, N11516, N1184, N1115, N5760);
and AND2 (N11522, N11511, N11030);
nand NAND3 (N11523, N11517, N10437, N3194);
or OR3 (N11524, N11507, N7672, N8020);
nand NAND3 (N11525, N11500, N5305, N2394);
and AND4 (N11526, N11509, N2780, N1841, N6455);
nand NAND3 (N11527, N11522, N3498, N923);
and AND3 (N11528, N11512, N10447, N2902);
xor XOR2 (N11529, N11527, N7862);
xor XOR2 (N11530, N11524, N1144);
xor XOR2 (N11531, N11530, N1509);
and AND3 (N11532, N11519, N193, N3168);
not NOT1 (N11533, N11515);
not NOT1 (N11534, N11529);
nor NOR3 (N11535, N11523, N11068, N8782);
xor XOR2 (N11536, N11520, N10576);
nand NAND3 (N11537, N11536, N11183, N7035);
nor NOR2 (N11538, N11537, N11524);
nor NOR2 (N11539, N11535, N5611);
xor XOR2 (N11540, N11531, N9102);
buf BUF1 (N11541, N11521);
nor NOR2 (N11542, N11528, N10649);
nor NOR3 (N11543, N11534, N7209, N1351);
and AND2 (N11544, N11540, N7007);
buf BUF1 (N11545, N11526);
and AND3 (N11546, N11542, N9151, N3764);
and AND2 (N11547, N11539, N7095);
buf BUF1 (N11548, N11538);
xor XOR2 (N11549, N11525, N3584);
and AND3 (N11550, N11532, N4994, N5377);
xor XOR2 (N11551, N11548, N6564);
not NOT1 (N11552, N11547);
xor XOR2 (N11553, N11546, N5032);
and AND4 (N11554, N11551, N11182, N1592, N1924);
buf BUF1 (N11555, N11545);
xor XOR2 (N11556, N11533, N3529);
nand NAND4 (N11557, N11553, N2272, N8947, N10036);
buf BUF1 (N11558, N11544);
and AND2 (N11559, N11549, N10006);
nor NOR4 (N11560, N11552, N211, N10048, N10379);
xor XOR2 (N11561, N11559, N2661);
buf BUF1 (N11562, N11555);
not NOT1 (N11563, N11554);
nand NAND3 (N11564, N11556, N577, N2435);
and AND4 (N11565, N11557, N9256, N2816, N3499);
not NOT1 (N11566, N11561);
buf BUF1 (N11567, N11565);
nor NOR2 (N11568, N11543, N5600);
nor NOR4 (N11569, N11567, N10628, N6445, N5327);
nand NAND4 (N11570, N11563, N10293, N7749, N8250);
or OR3 (N11571, N11541, N11007, N4162);
xor XOR2 (N11572, N11564, N7367);
or OR2 (N11573, N11558, N9424);
and AND2 (N11574, N11560, N9532);
or OR4 (N11575, N11569, N10947, N4162, N10885);
or OR2 (N11576, N11568, N2152);
buf BUF1 (N11577, N11572);
or OR2 (N11578, N11562, N8449);
not NOT1 (N11579, N11576);
and AND4 (N11580, N11574, N923, N1740, N581);
nand NAND4 (N11581, N11578, N2883, N6370, N3244);
nor NOR4 (N11582, N11571, N4470, N5607, N1255);
or OR4 (N11583, N11566, N8493, N11273, N790);
nor NOR2 (N11584, N11575, N5400);
and AND2 (N11585, N11550, N6226);
nor NOR3 (N11586, N11585, N9462, N2246);
not NOT1 (N11587, N11584);
nand NAND4 (N11588, N11586, N6802, N4056, N7127);
or OR2 (N11589, N11570, N10932);
buf BUF1 (N11590, N11587);
and AND2 (N11591, N11580, N7284);
nand NAND3 (N11592, N11589, N1145, N5240);
xor XOR2 (N11593, N11590, N1010);
nor NOR2 (N11594, N11588, N10427);
not NOT1 (N11595, N11579);
not NOT1 (N11596, N11582);
nor NOR3 (N11597, N11577, N10399, N7425);
not NOT1 (N11598, N11591);
not NOT1 (N11599, N11595);
xor XOR2 (N11600, N11581, N3035);
nand NAND2 (N11601, N11598, N591);
and AND3 (N11602, N11573, N7693, N4969);
nand NAND2 (N11603, N11600, N10168);
not NOT1 (N11604, N11602);
not NOT1 (N11605, N11593);
buf BUF1 (N11606, N11597);
buf BUF1 (N11607, N11603);
nor NOR3 (N11608, N11604, N8141, N595);
buf BUF1 (N11609, N11592);
not NOT1 (N11610, N11609);
not NOT1 (N11611, N11605);
or OR3 (N11612, N11599, N10718, N4983);
buf BUF1 (N11613, N11596);
not NOT1 (N11614, N11610);
not NOT1 (N11615, N11601);
nor NOR2 (N11616, N11606, N1880);
and AND2 (N11617, N11616, N1677);
nand NAND4 (N11618, N11617, N4510, N719, N428);
nor NOR4 (N11619, N11618, N1728, N2856, N4208);
buf BUF1 (N11620, N11608);
or OR4 (N11621, N11619, N10700, N7998, N924);
nor NOR2 (N11622, N11615, N10357);
nor NOR4 (N11623, N11614, N2861, N9992, N476);
nand NAND3 (N11624, N11611, N985, N4825);
xor XOR2 (N11625, N11621, N934);
and AND4 (N11626, N11583, N3172, N2002, N862);
or OR3 (N11627, N11625, N8963, N4604);
nand NAND4 (N11628, N11607, N10753, N5134, N8653);
not NOT1 (N11629, N11620);
buf BUF1 (N11630, N11622);
buf BUF1 (N11631, N11594);
not NOT1 (N11632, N11631);
buf BUF1 (N11633, N11612);
buf BUF1 (N11634, N11629);
xor XOR2 (N11635, N11633, N7610);
nand NAND3 (N11636, N11635, N2051, N3950);
not NOT1 (N11637, N11626);
and AND4 (N11638, N11634, N8651, N974, N7678);
and AND2 (N11639, N11623, N4386);
nand NAND2 (N11640, N11637, N5902);
nor NOR4 (N11641, N11627, N11584, N10981, N7666);
not NOT1 (N11642, N11613);
nand NAND3 (N11643, N11639, N6512, N8014);
buf BUF1 (N11644, N11630);
or OR3 (N11645, N11624, N635, N1746);
nor NOR3 (N11646, N11640, N6420, N2135);
buf BUF1 (N11647, N11646);
and AND2 (N11648, N11642, N2650);
nor NOR4 (N11649, N11638, N10615, N6404, N3414);
nor NOR3 (N11650, N11628, N760, N8828);
nor NOR2 (N11651, N11641, N8648);
nor NOR4 (N11652, N11636, N7467, N4468, N10809);
xor XOR2 (N11653, N11645, N9624);
xor XOR2 (N11654, N11651, N178);
xor XOR2 (N11655, N11648, N9112);
nor NOR2 (N11656, N11650, N125);
buf BUF1 (N11657, N11647);
buf BUF1 (N11658, N11653);
buf BUF1 (N11659, N11649);
or OR2 (N11660, N11632, N4407);
buf BUF1 (N11661, N11656);
xor XOR2 (N11662, N11654, N9273);
and AND4 (N11663, N11659, N10612, N6464, N1529);
and AND2 (N11664, N11658, N867);
nor NOR4 (N11665, N11655, N5730, N4834, N4190);
and AND4 (N11666, N11644, N164, N11083, N7093);
not NOT1 (N11667, N11660);
buf BUF1 (N11668, N11661);
or OR2 (N11669, N11665, N1441);
nor NOR4 (N11670, N11657, N5479, N3674, N1135);
nand NAND4 (N11671, N11662, N4975, N1729, N3735);
or OR4 (N11672, N11643, N5516, N3339, N9742);
nor NOR2 (N11673, N11669, N3871);
nor NOR3 (N11674, N11664, N10882, N7008);
not NOT1 (N11675, N11671);
xor XOR2 (N11676, N11672, N9684);
buf BUF1 (N11677, N11668);
and AND4 (N11678, N11663, N10239, N5281, N1805);
nand NAND2 (N11679, N11675, N6316);
nand NAND3 (N11680, N11678, N4692, N2848);
and AND3 (N11681, N11680, N9731, N10240);
not NOT1 (N11682, N11681);
or OR3 (N11683, N11677, N1474, N464);
and AND4 (N11684, N11673, N9793, N9501, N2490);
or OR4 (N11685, N11670, N3189, N1437, N6736);
or OR3 (N11686, N11682, N49, N3606);
and AND2 (N11687, N11667, N1636);
xor XOR2 (N11688, N11666, N727);
and AND4 (N11689, N11685, N1347, N6823, N8804);
buf BUF1 (N11690, N11676);
not NOT1 (N11691, N11687);
xor XOR2 (N11692, N11683, N2654);
not NOT1 (N11693, N11689);
or OR2 (N11694, N11693, N10013);
or OR2 (N11695, N11694, N2647);
and AND3 (N11696, N11692, N9812, N6982);
xor XOR2 (N11697, N11679, N269);
nand NAND2 (N11698, N11686, N3687);
xor XOR2 (N11699, N11696, N2753);
nand NAND3 (N11700, N11690, N8030, N2152);
nand NAND2 (N11701, N11699, N10489);
and AND2 (N11702, N11695, N230);
buf BUF1 (N11703, N11698);
xor XOR2 (N11704, N11688, N8286);
and AND2 (N11705, N11700, N3781);
nor NOR2 (N11706, N11691, N676);
buf BUF1 (N11707, N11702);
nand NAND4 (N11708, N11703, N8218, N8316, N11362);
xor XOR2 (N11709, N11697, N10784);
nand NAND4 (N11710, N11705, N4770, N2523, N5139);
nor NOR2 (N11711, N11706, N11383);
and AND3 (N11712, N11711, N5731, N9469);
not NOT1 (N11713, N11674);
not NOT1 (N11714, N11704);
nor NOR2 (N11715, N11714, N8526);
not NOT1 (N11716, N11710);
not NOT1 (N11717, N11712);
nor NOR3 (N11718, N11717, N8140, N7635);
or OR3 (N11719, N11684, N3413, N967);
buf BUF1 (N11720, N11716);
and AND2 (N11721, N11708, N7454);
xor XOR2 (N11722, N11719, N839);
buf BUF1 (N11723, N11721);
nor NOR3 (N11724, N11718, N10110, N9321);
and AND3 (N11725, N11720, N10430, N4477);
and AND4 (N11726, N11652, N4714, N7833, N11710);
nor NOR2 (N11727, N11726, N8870);
and AND4 (N11728, N11707, N10809, N6155, N1419);
nor NOR2 (N11729, N11713, N5324);
buf BUF1 (N11730, N11724);
not NOT1 (N11731, N11723);
or OR3 (N11732, N11730, N5793, N488);
nand NAND3 (N11733, N11715, N9197, N8482);
or OR4 (N11734, N11733, N9640, N8383, N7043);
nand NAND4 (N11735, N11734, N2749, N881, N10047);
nor NOR2 (N11736, N11722, N6820);
or OR4 (N11737, N11736, N5218, N9805, N4278);
not NOT1 (N11738, N11735);
and AND3 (N11739, N11728, N10363, N45);
buf BUF1 (N11740, N11727);
buf BUF1 (N11741, N11732);
and AND4 (N11742, N11709, N8696, N11572, N3712);
buf BUF1 (N11743, N11742);
or OR2 (N11744, N11739, N8666);
nor NOR2 (N11745, N11731, N2589);
or OR3 (N11746, N11740, N6877, N5509);
nor NOR4 (N11747, N11743, N6465, N6764, N2210);
nor NOR3 (N11748, N11744, N1624, N6833);
or OR3 (N11749, N11746, N3422, N2924);
not NOT1 (N11750, N11747);
nand NAND4 (N11751, N11749, N11090, N6748, N10517);
or OR3 (N11752, N11745, N42, N4335);
nor NOR4 (N11753, N11701, N11400, N4060, N1303);
buf BUF1 (N11754, N11725);
xor XOR2 (N11755, N11729, N5250);
not NOT1 (N11756, N11737);
or OR3 (N11757, N11754, N5863, N3772);
and AND2 (N11758, N11748, N3493);
buf BUF1 (N11759, N11753);
nor NOR3 (N11760, N11758, N616, N2611);
or OR2 (N11761, N11751, N1565);
buf BUF1 (N11762, N11756);
nand NAND2 (N11763, N11760, N2793);
or OR2 (N11764, N11755, N4029);
nor NOR3 (N11765, N11764, N7391, N9377);
nand NAND4 (N11766, N11741, N3978, N6300, N2032);
xor XOR2 (N11767, N11763, N1335);
nand NAND2 (N11768, N11767, N1505);
xor XOR2 (N11769, N11761, N3688);
xor XOR2 (N11770, N11765, N3171);
and AND4 (N11771, N11762, N6914, N5348, N8706);
or OR3 (N11772, N11766, N9880, N6520);
or OR4 (N11773, N11738, N2504, N5462, N3515);
nand NAND3 (N11774, N11773, N11628, N9792);
xor XOR2 (N11775, N11750, N6257);
buf BUF1 (N11776, N11771);
not NOT1 (N11777, N11776);
or OR2 (N11778, N11757, N1790);
nand NAND3 (N11779, N11772, N8488, N2242);
not NOT1 (N11780, N11779);
xor XOR2 (N11781, N11759, N1860);
nor NOR4 (N11782, N11774, N7695, N6541, N712);
nor NOR3 (N11783, N11769, N4228, N10259);
nand NAND4 (N11784, N11783, N296, N2828, N4798);
or OR2 (N11785, N11784, N7823);
xor XOR2 (N11786, N11777, N782);
buf BUF1 (N11787, N11782);
nand NAND4 (N11788, N11778, N2541, N5326, N2361);
nor NOR3 (N11789, N11780, N7530, N6019);
nand NAND4 (N11790, N11785, N2654, N2044, N4105);
nand NAND3 (N11791, N11770, N8766, N10523);
nand NAND3 (N11792, N11775, N11035, N9064);
or OR3 (N11793, N11792, N10319, N7672);
nor NOR2 (N11794, N11786, N3362);
buf BUF1 (N11795, N11791);
nand NAND3 (N11796, N11795, N11086, N6619);
nand NAND4 (N11797, N11796, N4171, N6566, N8950);
xor XOR2 (N11798, N11797, N3885);
and AND2 (N11799, N11793, N8737);
and AND3 (N11800, N11798, N9701, N8361);
xor XOR2 (N11801, N11790, N8717);
not NOT1 (N11802, N11800);
and AND4 (N11803, N11768, N4465, N5155, N153);
and AND3 (N11804, N11803, N3875, N6761);
nand NAND4 (N11805, N11801, N7223, N567, N3227);
buf BUF1 (N11806, N11799);
not NOT1 (N11807, N11804);
and AND4 (N11808, N11806, N625, N11349, N10421);
nand NAND2 (N11809, N11794, N2069);
buf BUF1 (N11810, N11802);
xor XOR2 (N11811, N11808, N6384);
nor NOR4 (N11812, N11805, N6140, N6802, N11329);
nand NAND3 (N11813, N11807, N960, N516);
xor XOR2 (N11814, N11788, N1177);
or OR4 (N11815, N11781, N8109, N7654, N9844);
buf BUF1 (N11816, N11789);
nor NOR2 (N11817, N11815, N9618);
not NOT1 (N11818, N11752);
buf BUF1 (N11819, N11809);
or OR4 (N11820, N11814, N2610, N5808, N10825);
xor XOR2 (N11821, N11819, N9449);
buf BUF1 (N11822, N11810);
nand NAND2 (N11823, N11816, N1601);
nand NAND2 (N11824, N11822, N10678);
nor NOR3 (N11825, N11812, N1119, N9579);
buf BUF1 (N11826, N11820);
or OR4 (N11827, N11821, N728, N9136, N1558);
nand NAND3 (N11828, N11824, N8976, N2325);
nor NOR3 (N11829, N11825, N387, N285);
not NOT1 (N11830, N11813);
not NOT1 (N11831, N11787);
not NOT1 (N11832, N11831);
nand NAND3 (N11833, N11832, N7871, N9975);
and AND4 (N11834, N11830, N1672, N7860, N7316);
and AND4 (N11835, N11818, N3594, N6369, N2614);
xor XOR2 (N11836, N11834, N2263);
not NOT1 (N11837, N11836);
or OR2 (N11838, N11835, N6509);
xor XOR2 (N11839, N11823, N8863);
nor NOR2 (N11840, N11837, N5253);
nor NOR2 (N11841, N11817, N4402);
or OR3 (N11842, N11840, N7013, N3185);
not NOT1 (N11843, N11828);
nand NAND2 (N11844, N11827, N11490);
buf BUF1 (N11845, N11838);
buf BUF1 (N11846, N11811);
not NOT1 (N11847, N11843);
nand NAND4 (N11848, N11846, N7545, N4878, N10425);
nor NOR3 (N11849, N11842, N8834, N9308);
buf BUF1 (N11850, N11844);
nor NOR2 (N11851, N11849, N9371);
not NOT1 (N11852, N11847);
nand NAND4 (N11853, N11852, N2662, N2639, N9433);
or OR3 (N11854, N11845, N807, N8064);
and AND3 (N11855, N11850, N7972, N7336);
buf BUF1 (N11856, N11841);
and AND2 (N11857, N11829, N6654);
nor NOR3 (N11858, N11855, N3322, N7513);
and AND4 (N11859, N11833, N8932, N4858, N8938);
nand NAND2 (N11860, N11848, N1823);
nor NOR2 (N11861, N11839, N5746);
and AND3 (N11862, N11851, N10513, N10151);
not NOT1 (N11863, N11859);
not NOT1 (N11864, N11858);
not NOT1 (N11865, N11861);
buf BUF1 (N11866, N11862);
nor NOR3 (N11867, N11866, N6904, N8886);
nor NOR2 (N11868, N11854, N9203);
not NOT1 (N11869, N11853);
xor XOR2 (N11870, N11856, N9258);
or OR3 (N11871, N11863, N9732, N3472);
or OR3 (N11872, N11867, N8735, N1804);
nor NOR4 (N11873, N11860, N9622, N9088, N724);
xor XOR2 (N11874, N11826, N8707);
or OR2 (N11875, N11874, N6836);
nand NAND2 (N11876, N11875, N7323);
nand NAND2 (N11877, N11871, N9101);
and AND3 (N11878, N11869, N212, N2978);
nand NAND3 (N11879, N11877, N5028, N3952);
nor NOR2 (N11880, N11870, N2574);
and AND3 (N11881, N11876, N8184, N9567);
buf BUF1 (N11882, N11881);
not NOT1 (N11883, N11864);
xor XOR2 (N11884, N11880, N7391);
nand NAND3 (N11885, N11879, N6991, N11713);
nor NOR4 (N11886, N11872, N2111, N7930, N7801);
or OR4 (N11887, N11878, N8914, N5276, N11382);
buf BUF1 (N11888, N11865);
nand NAND4 (N11889, N11882, N6167, N9835, N5894);
or OR4 (N11890, N11873, N9955, N2752, N1081);
and AND3 (N11891, N11890, N5702, N4384);
nor NOR4 (N11892, N11868, N342, N7620, N10478);
nor NOR2 (N11893, N11888, N4772);
buf BUF1 (N11894, N11886);
not NOT1 (N11895, N11883);
not NOT1 (N11896, N11887);
buf BUF1 (N11897, N11896);
or OR4 (N11898, N11894, N7446, N659, N10470);
and AND4 (N11899, N11892, N5873, N9119, N10232);
nor NOR4 (N11900, N11898, N821, N4861, N6237);
nand NAND2 (N11901, N11857, N1371);
or OR3 (N11902, N11897, N11241, N2009);
or OR4 (N11903, N11895, N7219, N5810, N8005);
nand NAND3 (N11904, N11903, N10533, N4733);
nor NOR3 (N11905, N11889, N10458, N4313);
xor XOR2 (N11906, N11884, N8652);
buf BUF1 (N11907, N11905);
buf BUF1 (N11908, N11906);
and AND3 (N11909, N11900, N6158, N10517);
xor XOR2 (N11910, N11909, N11602);
buf BUF1 (N11911, N11901);
not NOT1 (N11912, N11893);
buf BUF1 (N11913, N11902);
buf BUF1 (N11914, N11910);
and AND3 (N11915, N11911, N532, N8463);
or OR2 (N11916, N11891, N644);
xor XOR2 (N11917, N11885, N1243);
and AND2 (N11918, N11904, N1077);
nor NOR2 (N11919, N11917, N11321);
nand NAND2 (N11920, N11899, N6378);
not NOT1 (N11921, N11915);
or OR3 (N11922, N11921, N6516, N10728);
not NOT1 (N11923, N11908);
xor XOR2 (N11924, N11907, N5933);
not NOT1 (N11925, N11913);
buf BUF1 (N11926, N11918);
or OR3 (N11927, N11922, N1256, N112);
xor XOR2 (N11928, N11919, N1148);
xor XOR2 (N11929, N11926, N7517);
not NOT1 (N11930, N11912);
nand NAND4 (N11931, N11923, N8478, N9782, N5657);
and AND3 (N11932, N11929, N5495, N850);
nand NAND4 (N11933, N11920, N3966, N11766, N4699);
nand NAND2 (N11934, N11932, N5823);
nor NOR2 (N11935, N11930, N11499);
xor XOR2 (N11936, N11928, N7428);
not NOT1 (N11937, N11931);
nor NOR4 (N11938, N11927, N2125, N6672, N5502);
and AND4 (N11939, N11934, N4210, N10518, N2310);
not NOT1 (N11940, N11939);
buf BUF1 (N11941, N11937);
buf BUF1 (N11942, N11933);
not NOT1 (N11943, N11935);
buf BUF1 (N11944, N11924);
or OR3 (N11945, N11944, N3374, N7330);
or OR3 (N11946, N11941, N8707, N8070);
nand NAND4 (N11947, N11946, N10557, N5658, N3024);
nor NOR3 (N11948, N11943, N6356, N10828);
or OR3 (N11949, N11948, N2794, N8258);
buf BUF1 (N11950, N11945);
nand NAND4 (N11951, N11914, N10242, N5895, N2762);
xor XOR2 (N11952, N11916, N11235);
nor NOR2 (N11953, N11952, N9010);
and AND3 (N11954, N11950, N425, N1556);
or OR2 (N11955, N11938, N7133);
xor XOR2 (N11956, N11942, N7504);
nand NAND2 (N11957, N11956, N4432);
nor NOR2 (N11958, N11947, N7039);
or OR4 (N11959, N11949, N10189, N4826, N2660);
nor NOR3 (N11960, N11955, N1020, N4968);
xor XOR2 (N11961, N11959, N2826);
nor NOR3 (N11962, N11936, N5670, N8392);
or OR3 (N11963, N11940, N2942, N8915);
buf BUF1 (N11964, N11951);
nor NOR3 (N11965, N11954, N11378, N7940);
or OR3 (N11966, N11964, N2083, N9516);
xor XOR2 (N11967, N11961, N4275);
and AND2 (N11968, N11962, N1725);
buf BUF1 (N11969, N11963);
xor XOR2 (N11970, N11925, N6095);
or OR2 (N11971, N11969, N617);
and AND4 (N11972, N11970, N2314, N9567, N9705);
buf BUF1 (N11973, N11953);
nand NAND2 (N11974, N11960, N315);
nor NOR2 (N11975, N11965, N7947);
buf BUF1 (N11976, N11973);
nand NAND3 (N11977, N11968, N3752, N3009);
xor XOR2 (N11978, N11966, N9984);
or OR3 (N11979, N11976, N3165, N4947);
not NOT1 (N11980, N11957);
or OR4 (N11981, N11972, N3614, N11680, N3761);
and AND4 (N11982, N11981, N775, N5782, N1074);
and AND4 (N11983, N11977, N4115, N5680, N10580);
buf BUF1 (N11984, N11983);
or OR2 (N11985, N11971, N4053);
xor XOR2 (N11986, N11980, N9792);
nor NOR3 (N11987, N11958, N2141, N918);
nor NOR2 (N11988, N11985, N10010);
xor XOR2 (N11989, N11982, N11945);
xor XOR2 (N11990, N11978, N6850);
buf BUF1 (N11991, N11979);
not NOT1 (N11992, N11987);
or OR3 (N11993, N11990, N2444, N1860);
not NOT1 (N11994, N11991);
xor XOR2 (N11995, N11967, N3168);
and AND2 (N11996, N11975, N7107);
and AND4 (N11997, N11974, N11429, N9233, N2650);
buf BUF1 (N11998, N11997);
nor NOR4 (N11999, N11988, N11088, N3166, N2642);
xor XOR2 (N12000, N11989, N7640);
xor XOR2 (N12001, N11984, N3532);
and AND3 (N12002, N11996, N2462, N1655);
and AND2 (N12003, N12001, N6277);
nand NAND2 (N12004, N11994, N3253);
xor XOR2 (N12005, N11993, N163);
buf BUF1 (N12006, N12003);
xor XOR2 (N12007, N12005, N6721);
nand NAND3 (N12008, N11986, N9110, N5037);
not NOT1 (N12009, N12002);
or OR4 (N12010, N11995, N3414, N6917, N9544);
nand NAND3 (N12011, N12000, N4933, N11777);
nand NAND4 (N12012, N11992, N6351, N4903, N11111);
xor XOR2 (N12013, N12012, N1311);
buf BUF1 (N12014, N12010);
nor NOR2 (N12015, N11999, N10731);
and AND4 (N12016, N11998, N6303, N7536, N1173);
nor NOR2 (N12017, N12014, N6410);
buf BUF1 (N12018, N12008);
xor XOR2 (N12019, N12009, N11562);
buf BUF1 (N12020, N12019);
nor NOR4 (N12021, N12007, N7210, N10486, N8627);
xor XOR2 (N12022, N12011, N8622);
xor XOR2 (N12023, N12022, N7708);
or OR4 (N12024, N12020, N11171, N7833, N4864);
nor NOR2 (N12025, N12017, N4727);
nand NAND2 (N12026, N12024, N10562);
not NOT1 (N12027, N12015);
buf BUF1 (N12028, N12027);
xor XOR2 (N12029, N12021, N3296);
nor NOR4 (N12030, N12025, N7522, N1240, N5085);
not NOT1 (N12031, N12018);
nor NOR3 (N12032, N12026, N7522, N1981);
or OR4 (N12033, N12029, N7933, N3761, N5215);
buf BUF1 (N12034, N12023);
xor XOR2 (N12035, N12032, N9544);
xor XOR2 (N12036, N12030, N6054);
not NOT1 (N12037, N12013);
not NOT1 (N12038, N12037);
nor NOR2 (N12039, N12038, N11575);
not NOT1 (N12040, N12004);
buf BUF1 (N12041, N12035);
not NOT1 (N12042, N12036);
xor XOR2 (N12043, N12016, N4325);
nor NOR2 (N12044, N12040, N8782);
nor NOR4 (N12045, N12034, N2591, N8956, N3505);
and AND3 (N12046, N12006, N6214, N384);
or OR4 (N12047, N12028, N10828, N8131, N11715);
xor XOR2 (N12048, N12041, N103);
not NOT1 (N12049, N12039);
not NOT1 (N12050, N12046);
nor NOR4 (N12051, N12044, N1130, N6774, N11801);
xor XOR2 (N12052, N12031, N739);
nand NAND4 (N12053, N12047, N5524, N5485, N4829);
not NOT1 (N12054, N12053);
xor XOR2 (N12055, N12042, N9183);
nand NAND2 (N12056, N12051, N11651);
nand NAND4 (N12057, N12056, N933, N2147, N10237);
and AND2 (N12058, N12049, N6796);
nor NOR3 (N12059, N12050, N4909, N5983);
not NOT1 (N12060, N12054);
xor XOR2 (N12061, N12060, N7642);
buf BUF1 (N12062, N12058);
and AND2 (N12063, N12033, N2930);
and AND3 (N12064, N12063, N12033, N1216);
nand NAND3 (N12065, N12064, N11639, N11060);
buf BUF1 (N12066, N12055);
nand NAND3 (N12067, N12043, N882, N4694);
nor NOR4 (N12068, N12065, N2127, N9271, N1201);
buf BUF1 (N12069, N12052);
buf BUF1 (N12070, N12059);
and AND3 (N12071, N12068, N5050, N5474);
xor XOR2 (N12072, N12062, N7587);
and AND4 (N12073, N12066, N7379, N6676, N10553);
nor NOR3 (N12074, N12072, N4186, N11158);
not NOT1 (N12075, N12074);
or OR4 (N12076, N12057, N1627, N9045, N9969);
or OR2 (N12077, N12073, N2284);
and AND2 (N12078, N12075, N9452);
xor XOR2 (N12079, N12076, N1214);
nor NOR4 (N12080, N12048, N4809, N6458, N4419);
and AND3 (N12081, N12071, N1628, N1491);
nand NAND3 (N12082, N12045, N7029, N3788);
xor XOR2 (N12083, N12067, N9703);
buf BUF1 (N12084, N12077);
buf BUF1 (N12085, N12078);
nor NOR3 (N12086, N12069, N9646, N1063);
not NOT1 (N12087, N12079);
xor XOR2 (N12088, N12070, N10688);
or OR4 (N12089, N12080, N726, N10246, N688);
buf BUF1 (N12090, N12083);
or OR3 (N12091, N12061, N11567, N9604);
or OR3 (N12092, N12086, N2572, N2944);
buf BUF1 (N12093, N12092);
nand NAND2 (N12094, N12082, N4558);
nand NAND3 (N12095, N12081, N10782, N10127);
nor NOR2 (N12096, N12094, N11716);
xor XOR2 (N12097, N12096, N7214);
buf BUF1 (N12098, N12089);
and AND2 (N12099, N12095, N7371);
not NOT1 (N12100, N12098);
buf BUF1 (N12101, N12090);
buf BUF1 (N12102, N12097);
not NOT1 (N12103, N12099);
nor NOR2 (N12104, N12093, N5776);
xor XOR2 (N12105, N12102, N11131);
not NOT1 (N12106, N12087);
nor NOR3 (N12107, N12100, N6839, N7605);
nand NAND2 (N12108, N12104, N11672);
xor XOR2 (N12109, N12088, N3166);
nor NOR2 (N12110, N12109, N1080);
buf BUF1 (N12111, N12110);
buf BUF1 (N12112, N12106);
nor NOR4 (N12113, N12108, N724, N5216, N922);
xor XOR2 (N12114, N12101, N9140);
nand NAND4 (N12115, N12103, N5406, N8787, N2181);
nor NOR4 (N12116, N12084, N10919, N9606, N1565);
buf BUF1 (N12117, N12116);
and AND2 (N12118, N12107, N7363);
nor NOR4 (N12119, N12105, N2797, N10383, N6933);
nor NOR2 (N12120, N12117, N4240);
nor NOR3 (N12121, N12091, N7933, N5146);
and AND2 (N12122, N12115, N9470);
nor NOR2 (N12123, N12121, N3875);
xor XOR2 (N12124, N12118, N10237);
buf BUF1 (N12125, N12119);
not NOT1 (N12126, N12123);
not NOT1 (N12127, N12122);
xor XOR2 (N12128, N12120, N5474);
and AND3 (N12129, N12111, N1761, N8045);
not NOT1 (N12130, N12085);
and AND2 (N12131, N12125, N1263);
and AND2 (N12132, N12128, N7315);
nand NAND3 (N12133, N12114, N4733, N11223);
xor XOR2 (N12134, N12126, N1723);
nand NAND4 (N12135, N12113, N2618, N9559, N9168);
nand NAND2 (N12136, N12130, N4510);
nor NOR2 (N12137, N12134, N7420);
or OR3 (N12138, N12127, N384, N4784);
buf BUF1 (N12139, N12133);
or OR3 (N12140, N12112, N5066, N768);
or OR4 (N12141, N12140, N8055, N1546, N10784);
buf BUF1 (N12142, N12131);
and AND4 (N12143, N12136, N6001, N1773, N2695);
not NOT1 (N12144, N12143);
and AND2 (N12145, N12124, N3845);
and AND2 (N12146, N12137, N9208);
nor NOR4 (N12147, N12145, N10537, N7693, N2776);
buf BUF1 (N12148, N12144);
xor XOR2 (N12149, N12138, N6512);
or OR2 (N12150, N12129, N6577);
nand NAND4 (N12151, N12150, N3600, N7497, N6525);
not NOT1 (N12152, N12132);
buf BUF1 (N12153, N12146);
buf BUF1 (N12154, N12139);
not NOT1 (N12155, N12135);
nand NAND4 (N12156, N12151, N2775, N3767, N7825);
not NOT1 (N12157, N12141);
and AND2 (N12158, N12149, N3988);
and AND4 (N12159, N12158, N11074, N3559, N3963);
buf BUF1 (N12160, N12156);
nor NOR2 (N12161, N12154, N2090);
nand NAND3 (N12162, N12147, N11204, N7194);
nand NAND2 (N12163, N12152, N4390);
and AND4 (N12164, N12159, N8909, N2622, N5586);
buf BUF1 (N12165, N12161);
not NOT1 (N12166, N12163);
nand NAND3 (N12167, N12164, N7191, N8222);
or OR2 (N12168, N12167, N1488);
xor XOR2 (N12169, N12165, N11426);
nor NOR3 (N12170, N12157, N5200, N3665);
or OR3 (N12171, N12166, N1441, N2538);
not NOT1 (N12172, N12142);
and AND3 (N12173, N12172, N2557, N1514);
or OR4 (N12174, N12148, N2590, N3525, N6391);
nor NOR4 (N12175, N12170, N11276, N9520, N8379);
or OR4 (N12176, N12173, N7157, N2909, N2500);
nor NOR3 (N12177, N12175, N10463, N287);
xor XOR2 (N12178, N12169, N84);
and AND4 (N12179, N12174, N7428, N337, N5186);
nor NOR3 (N12180, N12179, N6973, N225);
xor XOR2 (N12181, N12171, N7876);
nand NAND2 (N12182, N12178, N8887);
nand NAND2 (N12183, N12180, N82);
not NOT1 (N12184, N12177);
nand NAND3 (N12185, N12153, N6799, N3431);
xor XOR2 (N12186, N12168, N6183);
or OR4 (N12187, N12185, N12136, N6291, N10358);
and AND2 (N12188, N12176, N7919);
nand NAND2 (N12189, N12183, N6520);
not NOT1 (N12190, N12188);
nor NOR2 (N12191, N12155, N7029);
nor NOR4 (N12192, N12191, N1884, N4804, N1321);
and AND2 (N12193, N12162, N10354);
xor XOR2 (N12194, N12190, N9330);
not NOT1 (N12195, N12182);
nand NAND2 (N12196, N12193, N3778);
not NOT1 (N12197, N12189);
xor XOR2 (N12198, N12184, N6073);
and AND4 (N12199, N12197, N9047, N675, N7119);
not NOT1 (N12200, N12195);
or OR3 (N12201, N12181, N5785, N6760);
and AND2 (N12202, N12200, N388);
nor NOR4 (N12203, N12202, N10593, N4945, N9161);
xor XOR2 (N12204, N12160, N9780);
and AND2 (N12205, N12196, N8023);
and AND3 (N12206, N12186, N2139, N8811);
not NOT1 (N12207, N12204);
nor NOR3 (N12208, N12206, N1507, N7604);
and AND4 (N12209, N12205, N12001, N1770, N11498);
or OR3 (N12210, N12198, N9484, N7117);
nand NAND3 (N12211, N12209, N5969, N1210);
nor NOR3 (N12212, N12201, N6977, N4448);
or OR2 (N12213, N12187, N11509);
and AND3 (N12214, N12210, N1789, N8834);
xor XOR2 (N12215, N12203, N10108);
not NOT1 (N12216, N12215);
nor NOR3 (N12217, N12194, N7789, N6488);
xor XOR2 (N12218, N12212, N3090);
or OR3 (N12219, N12213, N4028, N7893);
or OR2 (N12220, N12217, N10451);
nor NOR3 (N12221, N12199, N320, N4174);
nand NAND3 (N12222, N12216, N1304, N6308);
not NOT1 (N12223, N12192);
xor XOR2 (N12224, N12223, N8889);
xor XOR2 (N12225, N12220, N6321);
or OR3 (N12226, N12207, N9149, N4539);
or OR4 (N12227, N12208, N9632, N1008, N9881);
not NOT1 (N12228, N12224);
buf BUF1 (N12229, N12222);
nor NOR2 (N12230, N12218, N1942);
nor NOR4 (N12231, N12228, N8812, N10250, N5960);
buf BUF1 (N12232, N12219);
or OR4 (N12233, N12231, N996, N11314, N4621);
or OR2 (N12234, N12214, N3092);
buf BUF1 (N12235, N12227);
xor XOR2 (N12236, N12226, N7505);
nand NAND3 (N12237, N12221, N12050, N11325);
not NOT1 (N12238, N12229);
or OR3 (N12239, N12225, N1603, N6741);
not NOT1 (N12240, N12239);
nand NAND2 (N12241, N12230, N1860);
buf BUF1 (N12242, N12211);
nor NOR2 (N12243, N12234, N6737);
xor XOR2 (N12244, N12233, N484);
and AND3 (N12245, N12236, N4121, N3315);
nand NAND4 (N12246, N12238, N9285, N303, N9005);
not NOT1 (N12247, N12240);
nor NOR4 (N12248, N12242, N7111, N7446, N8972);
and AND3 (N12249, N12247, N1654, N2807);
not NOT1 (N12250, N12232);
nand NAND4 (N12251, N12243, N2027, N2141, N5717);
nand NAND4 (N12252, N12250, N8590, N10281, N2454);
or OR2 (N12253, N12235, N8347);
buf BUF1 (N12254, N12237);
nand NAND3 (N12255, N12254, N5949, N10898);
xor XOR2 (N12256, N12245, N5426);
not NOT1 (N12257, N12249);
nor NOR2 (N12258, N12251, N6498);
and AND4 (N12259, N12258, N7949, N11239, N1090);
nand NAND2 (N12260, N12255, N6816);
or OR4 (N12261, N12257, N8005, N10293, N3314);
or OR4 (N12262, N12256, N3480, N6622, N528);
or OR3 (N12263, N12261, N8316, N8994);
not NOT1 (N12264, N12246);
and AND4 (N12265, N12248, N3608, N5567, N10272);
nor NOR3 (N12266, N12253, N8967, N11152);
not NOT1 (N12267, N12265);
buf BUF1 (N12268, N12263);
buf BUF1 (N12269, N12241);
or OR4 (N12270, N12260, N2075, N2301, N9279);
xor XOR2 (N12271, N12266, N8736);
or OR3 (N12272, N12252, N1573, N5027);
and AND2 (N12273, N12271, N6523);
not NOT1 (N12274, N12259);
not NOT1 (N12275, N12262);
nand NAND3 (N12276, N12273, N8925, N1829);
not NOT1 (N12277, N12268);
nor NOR2 (N12278, N12270, N2033);
buf BUF1 (N12279, N12277);
and AND2 (N12280, N12272, N821);
buf BUF1 (N12281, N12274);
buf BUF1 (N12282, N12279);
nand NAND3 (N12283, N12281, N7223, N5279);
and AND3 (N12284, N12278, N8654, N5419);
buf BUF1 (N12285, N12282);
xor XOR2 (N12286, N12264, N825);
nor NOR4 (N12287, N12267, N11401, N5133, N333);
xor XOR2 (N12288, N12286, N4893);
nand NAND2 (N12289, N12244, N6081);
nor NOR3 (N12290, N12269, N1132, N2556);
nand NAND3 (N12291, N12290, N8624, N4569);
and AND2 (N12292, N12280, N4280);
nor NOR4 (N12293, N12291, N4522, N1238, N3780);
and AND3 (N12294, N12275, N11269, N9802);
xor XOR2 (N12295, N12288, N2760);
nor NOR4 (N12296, N12284, N8329, N4207, N9751);
xor XOR2 (N12297, N12296, N12229);
and AND3 (N12298, N12292, N5791, N5573);
not NOT1 (N12299, N12276);
nand NAND3 (N12300, N12297, N466, N9911);
or OR3 (N12301, N12289, N4792, N10568);
or OR3 (N12302, N12300, N2194, N10091);
not NOT1 (N12303, N12287);
not NOT1 (N12304, N12303);
nand NAND2 (N12305, N12302, N12216);
or OR2 (N12306, N12304, N7460);
nor NOR4 (N12307, N12305, N1459, N11024, N4918);
and AND2 (N12308, N12285, N303);
and AND2 (N12309, N12308, N9504);
xor XOR2 (N12310, N12301, N8360);
or OR4 (N12311, N12299, N1079, N7427, N9686);
nand NAND3 (N12312, N12294, N6375, N5734);
buf BUF1 (N12313, N12309);
buf BUF1 (N12314, N12307);
nand NAND3 (N12315, N12306, N9047, N5394);
nor NOR4 (N12316, N12310, N6591, N4165, N6787);
xor XOR2 (N12317, N12283, N8750);
xor XOR2 (N12318, N12293, N11692);
and AND3 (N12319, N12316, N6155, N2951);
xor XOR2 (N12320, N12313, N8854);
nor NOR4 (N12321, N12298, N8250, N6569, N2845);
and AND2 (N12322, N12321, N11296);
and AND4 (N12323, N12317, N421, N6261, N7304);
nand NAND4 (N12324, N12318, N9450, N1421, N1592);
nand NAND4 (N12325, N12324, N9316, N10781, N82);
or OR2 (N12326, N12319, N2161);
not NOT1 (N12327, N12322);
or OR3 (N12328, N12315, N3494, N10791);
or OR4 (N12329, N12295, N10467, N7258, N9241);
xor XOR2 (N12330, N12320, N4968);
or OR4 (N12331, N12314, N8368, N7807, N12140);
nand NAND2 (N12332, N12312, N11019);
xor XOR2 (N12333, N12323, N415);
or OR3 (N12334, N12329, N7046, N4216);
buf BUF1 (N12335, N12334);
and AND3 (N12336, N12325, N3559, N433);
and AND2 (N12337, N12311, N6557);
and AND3 (N12338, N12326, N9231, N7536);
and AND3 (N12339, N12328, N4089, N7008);
nor NOR4 (N12340, N12337, N8689, N11150, N5261);
and AND2 (N12341, N12340, N1320);
nand NAND4 (N12342, N12332, N9051, N3469, N1746);
or OR2 (N12343, N12336, N1623);
nor NOR4 (N12344, N12339, N158, N12211, N4508);
nor NOR3 (N12345, N12343, N11603, N7892);
and AND2 (N12346, N12344, N3945);
nand NAND4 (N12347, N12345, N2974, N276, N350);
nand NAND2 (N12348, N12338, N11900);
buf BUF1 (N12349, N12348);
nor NOR3 (N12350, N12333, N3259, N7813);
buf BUF1 (N12351, N12342);
or OR4 (N12352, N12327, N8966, N6050, N6111);
buf BUF1 (N12353, N12352);
buf BUF1 (N12354, N12351);
nand NAND4 (N12355, N12341, N10565, N2030, N10392);
and AND4 (N12356, N12349, N6278, N10681, N5422);
nand NAND3 (N12357, N12330, N10553, N1760);
not NOT1 (N12358, N12350);
not NOT1 (N12359, N12347);
or OR2 (N12360, N12357, N3822);
nand NAND4 (N12361, N12331, N2290, N2808, N9103);
buf BUF1 (N12362, N12354);
nor NOR3 (N12363, N12335, N3561, N5111);
or OR4 (N12364, N12353, N7842, N8053, N10);
xor XOR2 (N12365, N12361, N1008);
xor XOR2 (N12366, N12355, N5513);
nor NOR4 (N12367, N12362, N12294, N1986, N9576);
xor XOR2 (N12368, N12358, N10400);
nand NAND4 (N12369, N12365, N3744, N625, N3771);
and AND2 (N12370, N12360, N1058);
nand NAND4 (N12371, N12364, N12028, N3245, N9083);
not NOT1 (N12372, N12363);
xor XOR2 (N12373, N12346, N807);
and AND4 (N12374, N12366, N11843, N12152, N6626);
buf BUF1 (N12375, N12372);
nand NAND4 (N12376, N12367, N1810, N8092, N9648);
xor XOR2 (N12377, N12359, N6098);
not NOT1 (N12378, N12370);
and AND2 (N12379, N12356, N10621);
buf BUF1 (N12380, N12375);
buf BUF1 (N12381, N12369);
or OR4 (N12382, N12377, N6684, N12295, N8176);
and AND2 (N12383, N12379, N1514);
buf BUF1 (N12384, N12373);
nand NAND4 (N12385, N12384, N7757, N2931, N1676);
xor XOR2 (N12386, N12380, N7970);
xor XOR2 (N12387, N12386, N8518);
buf BUF1 (N12388, N12381);
not NOT1 (N12389, N12368);
xor XOR2 (N12390, N12371, N1765);
buf BUF1 (N12391, N12378);
nand NAND3 (N12392, N12389, N11564, N284);
or OR4 (N12393, N12376, N9691, N11280, N4799);
buf BUF1 (N12394, N12393);
xor XOR2 (N12395, N12374, N320);
buf BUF1 (N12396, N12385);
or OR4 (N12397, N12396, N6003, N4993, N2250);
or OR2 (N12398, N12387, N10342);
and AND2 (N12399, N12392, N7431);
or OR3 (N12400, N12399, N3184, N3697);
nor NOR2 (N12401, N12390, N6095);
buf BUF1 (N12402, N12382);
xor XOR2 (N12403, N12397, N11664);
not NOT1 (N12404, N12394);
xor XOR2 (N12405, N12404, N2305);
buf BUF1 (N12406, N12383);
or OR4 (N12407, N12401, N5308, N10943, N5161);
xor XOR2 (N12408, N12402, N4921);
and AND2 (N12409, N12391, N6530);
buf BUF1 (N12410, N12405);
nand NAND3 (N12411, N12410, N8131, N4702);
or OR4 (N12412, N12398, N9406, N6523, N6257);
nor NOR3 (N12413, N12411, N984, N11532);
xor XOR2 (N12414, N12400, N10081);
xor XOR2 (N12415, N12413, N699);
or OR2 (N12416, N12395, N5475);
buf BUF1 (N12417, N12403);
or OR4 (N12418, N12408, N5537, N9461, N6979);
or OR4 (N12419, N12418, N9794, N666, N2996);
not NOT1 (N12420, N12414);
and AND4 (N12421, N12409, N4329, N2505, N11701);
xor XOR2 (N12422, N12415, N6001);
buf BUF1 (N12423, N12420);
not NOT1 (N12424, N12407);
and AND4 (N12425, N12419, N10822, N10678, N4366);
xor XOR2 (N12426, N12425, N9425);
xor XOR2 (N12427, N12412, N8963);
xor XOR2 (N12428, N12426, N5058);
nor NOR3 (N12429, N12428, N3010, N10275);
and AND2 (N12430, N12388, N7912);
not NOT1 (N12431, N12422);
nor NOR4 (N12432, N12416, N12262, N3925, N6682);
nor NOR2 (N12433, N12432, N4975);
nand NAND4 (N12434, N12433, N11847, N6910, N12097);
and AND3 (N12435, N12423, N14, N1952);
buf BUF1 (N12436, N12421);
and AND2 (N12437, N12424, N7919);
xor XOR2 (N12438, N12406, N1543);
xor XOR2 (N12439, N12435, N747);
nand NAND4 (N12440, N12438, N4244, N384, N1986);
and AND4 (N12441, N12430, N8034, N5165, N12139);
buf BUF1 (N12442, N12417);
and AND4 (N12443, N12434, N10121, N5633, N9898);
buf BUF1 (N12444, N12439);
and AND3 (N12445, N12427, N3521, N10565);
buf BUF1 (N12446, N12431);
not NOT1 (N12447, N12440);
not NOT1 (N12448, N12447);
not NOT1 (N12449, N12444);
not NOT1 (N12450, N12446);
not NOT1 (N12451, N12449);
xor XOR2 (N12452, N12448, N902);
nor NOR3 (N12453, N12452, N11188, N12139);
xor XOR2 (N12454, N12451, N1118);
nand NAND4 (N12455, N12442, N193, N7988, N7927);
nor NOR4 (N12456, N12455, N7382, N6503, N6272);
or OR2 (N12457, N12441, N8850);
or OR3 (N12458, N12457, N4546, N9124);
not NOT1 (N12459, N12445);
nor NOR3 (N12460, N12429, N10569, N4991);
buf BUF1 (N12461, N12459);
nand NAND4 (N12462, N12453, N5840, N5750, N3713);
nand NAND3 (N12463, N12436, N346, N7805);
or OR3 (N12464, N12437, N7679, N5273);
nand NAND3 (N12465, N12454, N1716, N2087);
or OR2 (N12466, N12462, N10643);
not NOT1 (N12467, N12460);
nor NOR4 (N12468, N12461, N837, N11523, N1153);
nor NOR3 (N12469, N12465, N3224, N12323);
xor XOR2 (N12470, N12463, N11708);
buf BUF1 (N12471, N12450);
xor XOR2 (N12472, N12467, N9796);
not NOT1 (N12473, N12458);
nor NOR4 (N12474, N12468, N4181, N2551, N841);
xor XOR2 (N12475, N12469, N693);
nor NOR2 (N12476, N12471, N8367);
buf BUF1 (N12477, N12464);
xor XOR2 (N12478, N12475, N5006);
or OR2 (N12479, N12472, N4107);
nor NOR3 (N12480, N12456, N1621, N2664);
and AND4 (N12481, N12477, N5894, N9576, N3984);
not NOT1 (N12482, N12480);
buf BUF1 (N12483, N12473);
or OR4 (N12484, N12481, N11601, N5306, N2694);
or OR3 (N12485, N12474, N7409, N6268);
buf BUF1 (N12486, N12478);
or OR2 (N12487, N12479, N2966);
or OR3 (N12488, N12470, N9857, N9361);
nor NOR4 (N12489, N12443, N2434, N4662, N6849);
buf BUF1 (N12490, N12486);
or OR3 (N12491, N12484, N9355, N9811);
not NOT1 (N12492, N12466);
and AND3 (N12493, N12485, N8156, N12140);
buf BUF1 (N12494, N12476);
and AND3 (N12495, N12489, N3251, N4398);
xor XOR2 (N12496, N12495, N9610);
and AND4 (N12497, N12487, N7078, N6159, N2109);
buf BUF1 (N12498, N12482);
or OR3 (N12499, N12491, N5084, N354);
nor NOR4 (N12500, N12497, N4012, N1226, N2834);
or OR4 (N12501, N12499, N249, N3574, N4568);
xor XOR2 (N12502, N12496, N2886);
nand NAND2 (N12503, N12488, N2101);
xor XOR2 (N12504, N12494, N9102);
or OR4 (N12505, N12483, N203, N11563, N7047);
nand NAND4 (N12506, N12492, N4156, N194, N11576);
not NOT1 (N12507, N12500);
buf BUF1 (N12508, N12504);
and AND4 (N12509, N12501, N5119, N1939, N3270);
nand NAND3 (N12510, N12507, N10243, N4078);
nor NOR3 (N12511, N12498, N2862, N5591);
xor XOR2 (N12512, N12509, N7841);
not NOT1 (N12513, N12502);
or OR2 (N12514, N12506, N11389);
nor NOR2 (N12515, N12510, N6563);
nand NAND2 (N12516, N12505, N11971);
or OR4 (N12517, N12511, N10818, N8420, N10380);
buf BUF1 (N12518, N12490);
buf BUF1 (N12519, N12513);
not NOT1 (N12520, N12518);
xor XOR2 (N12521, N12517, N9703);
and AND3 (N12522, N12515, N9326, N1101);
nand NAND2 (N12523, N12508, N3416);
nor NOR3 (N12524, N12521, N3581, N10851);
nand NAND2 (N12525, N12493, N9049);
buf BUF1 (N12526, N12525);
buf BUF1 (N12527, N12522);
not NOT1 (N12528, N12514);
nand NAND3 (N12529, N12524, N7606, N11260);
and AND3 (N12530, N12512, N2217, N38);
not NOT1 (N12531, N12516);
not NOT1 (N12532, N12520);
nand NAND3 (N12533, N12531, N9454, N4120);
xor XOR2 (N12534, N12527, N2365);
not NOT1 (N12535, N12523);
not NOT1 (N12536, N12526);
and AND3 (N12537, N12528, N691, N8216);
not NOT1 (N12538, N12530);
buf BUF1 (N12539, N12538);
nand NAND3 (N12540, N12519, N1881, N12274);
buf BUF1 (N12541, N12537);
xor XOR2 (N12542, N12536, N8132);
not NOT1 (N12543, N12540);
or OR4 (N12544, N12532, N10332, N3480, N4208);
and AND3 (N12545, N12535, N1326, N9059);
buf BUF1 (N12546, N12543);
xor XOR2 (N12547, N12542, N8301);
nand NAND4 (N12548, N12547, N3645, N7965, N3126);
not NOT1 (N12549, N12544);
nor NOR4 (N12550, N12529, N2507, N12250, N11127);
nand NAND2 (N12551, N12550, N36);
nand NAND2 (N12552, N12503, N12210);
and AND2 (N12553, N12552, N2727);
buf BUF1 (N12554, N12546);
buf BUF1 (N12555, N12545);
xor XOR2 (N12556, N12554, N12322);
nand NAND4 (N12557, N12553, N116, N2953, N2826);
not NOT1 (N12558, N12539);
or OR3 (N12559, N12557, N10173, N8548);
xor XOR2 (N12560, N12558, N809);
xor XOR2 (N12561, N12548, N2566);
xor XOR2 (N12562, N12561, N9566);
buf BUF1 (N12563, N12559);
or OR2 (N12564, N12556, N122);
nor NOR2 (N12565, N12560, N5131);
and AND2 (N12566, N12533, N10229);
not NOT1 (N12567, N12549);
nand NAND3 (N12568, N12563, N4532, N7669);
xor XOR2 (N12569, N12555, N11428);
or OR4 (N12570, N12562, N12306, N8985, N10040);
buf BUF1 (N12571, N12570);
xor XOR2 (N12572, N12541, N3905);
and AND4 (N12573, N12567, N11377, N1583, N12095);
and AND3 (N12574, N12534, N1417, N1295);
not NOT1 (N12575, N12566);
buf BUF1 (N12576, N12569);
not NOT1 (N12577, N12568);
not NOT1 (N12578, N12551);
nand NAND2 (N12579, N12575, N10205);
and AND4 (N12580, N12579, N6040, N11294, N3839);
or OR4 (N12581, N12572, N8648, N11817, N9841);
buf BUF1 (N12582, N12565);
and AND4 (N12583, N12574, N10641, N6668, N1117);
nand NAND4 (N12584, N12576, N500, N1291, N3196);
buf BUF1 (N12585, N12584);
buf BUF1 (N12586, N12581);
not NOT1 (N12587, N12582);
nor NOR3 (N12588, N12578, N6024, N5176);
nor NOR4 (N12589, N12588, N9028, N11687, N6750);
and AND2 (N12590, N12573, N8167);
and AND3 (N12591, N12587, N12117, N388);
xor XOR2 (N12592, N12591, N6641);
buf BUF1 (N12593, N12585);
nand NAND3 (N12594, N12571, N8990, N261);
buf BUF1 (N12595, N12589);
and AND4 (N12596, N12586, N5364, N274, N3727);
or OR3 (N12597, N12577, N7403, N3451);
or OR4 (N12598, N12594, N4127, N3376, N1321);
or OR2 (N12599, N12583, N1978);
and AND3 (N12600, N12590, N7736, N10516);
not NOT1 (N12601, N12580);
and AND2 (N12602, N12593, N1343);
not NOT1 (N12603, N12598);
buf BUF1 (N12604, N12592);
nand NAND2 (N12605, N12599, N7394);
and AND2 (N12606, N12564, N3635);
nor NOR4 (N12607, N12602, N9516, N12574, N7158);
xor XOR2 (N12608, N12606, N10446);
not NOT1 (N12609, N12603);
not NOT1 (N12610, N12605);
xor XOR2 (N12611, N12600, N5935);
xor XOR2 (N12612, N12597, N12353);
buf BUF1 (N12613, N12601);
nand NAND2 (N12614, N12596, N329);
or OR3 (N12615, N12610, N11282, N4412);
or OR3 (N12616, N12613, N2974, N4487);
or OR2 (N12617, N12616, N1546);
nor NOR4 (N12618, N12609, N5130, N997, N5568);
or OR2 (N12619, N12618, N7957);
nor NOR3 (N12620, N12615, N9922, N6209);
not NOT1 (N12621, N12619);
nor NOR4 (N12622, N12617, N10674, N7153, N12152);
not NOT1 (N12623, N12621);
nand NAND2 (N12624, N12612, N2818);
not NOT1 (N12625, N12622);
xor XOR2 (N12626, N12620, N9376);
buf BUF1 (N12627, N12625);
or OR4 (N12628, N12611, N1882, N4431, N7851);
or OR2 (N12629, N12608, N11148);
and AND2 (N12630, N12595, N12522);
nand NAND4 (N12631, N12628, N7978, N4800, N4694);
nor NOR3 (N12632, N12604, N2904, N5917);
nand NAND3 (N12633, N12614, N2548, N228);
and AND4 (N12634, N12630, N9410, N62, N12179);
nand NAND2 (N12635, N12631, N8852);
nor NOR4 (N12636, N12607, N5422, N10783, N3037);
nand NAND4 (N12637, N12629, N8497, N694, N4670);
buf BUF1 (N12638, N12634);
nor NOR3 (N12639, N12637, N5915, N10086);
and AND3 (N12640, N12638, N2571, N5899);
xor XOR2 (N12641, N12640, N10358);
not NOT1 (N12642, N12641);
nand NAND3 (N12643, N12639, N10228, N98);
and AND3 (N12644, N12635, N11373, N2372);
and AND2 (N12645, N12632, N3076);
buf BUF1 (N12646, N12643);
not NOT1 (N12647, N12626);
xor XOR2 (N12648, N12646, N1161);
or OR3 (N12649, N12636, N5753, N1540);
and AND3 (N12650, N12642, N11061, N2032);
and AND2 (N12651, N12645, N5915);
nor NOR3 (N12652, N12648, N5998, N7204);
nand NAND2 (N12653, N12633, N4630);
or OR3 (N12654, N12623, N9953, N3731);
or OR2 (N12655, N12644, N6301);
buf BUF1 (N12656, N12651);
not NOT1 (N12657, N12653);
and AND3 (N12658, N12655, N7708, N6101);
nor NOR4 (N12659, N12652, N4980, N10180, N3818);
xor XOR2 (N12660, N12650, N6803);
nand NAND4 (N12661, N12658, N2538, N10417, N2512);
nand NAND3 (N12662, N12649, N3831, N4382);
nand NAND2 (N12663, N12654, N9030);
and AND2 (N12664, N12647, N9970);
not NOT1 (N12665, N12656);
nor NOR2 (N12666, N12664, N1136);
nand NAND3 (N12667, N12657, N5063, N9798);
nor NOR2 (N12668, N12624, N12275);
xor XOR2 (N12669, N12667, N3028);
xor XOR2 (N12670, N12665, N1962);
nand NAND3 (N12671, N12627, N8152, N8909);
buf BUF1 (N12672, N12661);
xor XOR2 (N12673, N12668, N7334);
or OR3 (N12674, N12669, N10944, N5417);
buf BUF1 (N12675, N12673);
xor XOR2 (N12676, N12672, N10516);
nand NAND2 (N12677, N12675, N10449);
xor XOR2 (N12678, N12662, N12203);
not NOT1 (N12679, N12663);
or OR3 (N12680, N12666, N7316, N1484);
not NOT1 (N12681, N12677);
not NOT1 (N12682, N12660);
or OR3 (N12683, N12676, N10909, N10016);
not NOT1 (N12684, N12682);
and AND4 (N12685, N12681, N9085, N8052, N7987);
or OR4 (N12686, N12671, N8580, N11689, N7392);
or OR4 (N12687, N12679, N10080, N7636, N7619);
and AND3 (N12688, N12680, N4800, N2527);
nor NOR3 (N12689, N12685, N10165, N10824);
nor NOR4 (N12690, N12678, N8055, N3076, N11958);
or OR4 (N12691, N12670, N7460, N5507, N11531);
or OR4 (N12692, N12674, N8330, N528, N595);
or OR3 (N12693, N12683, N2444, N7674);
xor XOR2 (N12694, N12684, N10484);
xor XOR2 (N12695, N12693, N482);
buf BUF1 (N12696, N12659);
not NOT1 (N12697, N12687);
and AND4 (N12698, N12690, N10583, N10906, N6563);
nand NAND4 (N12699, N12696, N1880, N6300, N4003);
nand NAND4 (N12700, N12686, N5730, N4530, N5282);
not NOT1 (N12701, N12691);
or OR3 (N12702, N12689, N236, N7220);
or OR4 (N12703, N12702, N7673, N3806, N783);
nor NOR3 (N12704, N12700, N9703, N2015);
buf BUF1 (N12705, N12698);
buf BUF1 (N12706, N12688);
xor XOR2 (N12707, N12704, N7820);
buf BUF1 (N12708, N12705);
nand NAND2 (N12709, N12701, N12108);
buf BUF1 (N12710, N12697);
and AND4 (N12711, N12699, N11947, N1138, N7369);
xor XOR2 (N12712, N12708, N6806);
nor NOR2 (N12713, N12711, N2578);
nor NOR4 (N12714, N12706, N6492, N2384, N1442);
buf BUF1 (N12715, N12694);
and AND2 (N12716, N12713, N7108);
and AND4 (N12717, N12715, N9877, N6992, N3010);
nor NOR3 (N12718, N12703, N350, N8231);
nand NAND2 (N12719, N12710, N9409);
xor XOR2 (N12720, N12716, N2927);
and AND2 (N12721, N12714, N1304);
buf BUF1 (N12722, N12707);
nand NAND3 (N12723, N12718, N5652, N8020);
or OR4 (N12724, N12720, N9248, N3442, N3336);
and AND4 (N12725, N12717, N1673, N3194, N4141);
not NOT1 (N12726, N12724);
not NOT1 (N12727, N12712);
or OR4 (N12728, N12725, N1324, N11403, N12447);
or OR4 (N12729, N12728, N5560, N10354, N12209);
nor NOR4 (N12730, N12729, N2086, N11625, N1347);
and AND3 (N12731, N12723, N8864, N2409);
nand NAND2 (N12732, N12727, N3165);
and AND3 (N12733, N12730, N8253, N12442);
and AND3 (N12734, N12695, N11262, N10190);
buf BUF1 (N12735, N12726);
buf BUF1 (N12736, N12709);
nor NOR4 (N12737, N12733, N3590, N9132, N10895);
nor NOR4 (N12738, N12737, N3033, N12494, N10705);
buf BUF1 (N12739, N12735);
or OR3 (N12740, N12736, N2896, N6945);
and AND2 (N12741, N12739, N11553);
nor NOR3 (N12742, N12738, N8694, N918);
nor NOR2 (N12743, N12719, N3169);
xor XOR2 (N12744, N12731, N6547);
nor NOR2 (N12745, N12692, N6266);
xor XOR2 (N12746, N12744, N5434);
nor NOR4 (N12747, N12745, N8732, N6004, N2121);
not NOT1 (N12748, N12740);
or OR2 (N12749, N12721, N5985);
xor XOR2 (N12750, N12734, N10624);
or OR2 (N12751, N12747, N12405);
nor NOR4 (N12752, N12746, N940, N5828, N655);
buf BUF1 (N12753, N12749);
not NOT1 (N12754, N12750);
buf BUF1 (N12755, N12743);
nand NAND2 (N12756, N12751, N11546);
and AND2 (N12757, N12748, N23);
not NOT1 (N12758, N12732);
buf BUF1 (N12759, N12756);
or OR2 (N12760, N12752, N4223);
nand NAND4 (N12761, N12741, N6014, N9464, N5508);
or OR2 (N12762, N12761, N2449);
buf BUF1 (N12763, N12759);
buf BUF1 (N12764, N12754);
nor NOR3 (N12765, N12764, N975, N11225);
buf BUF1 (N12766, N12760);
buf BUF1 (N12767, N12762);
and AND3 (N12768, N12766, N9862, N2635);
nand NAND3 (N12769, N12765, N3392, N10388);
and AND2 (N12770, N12768, N8500);
nand NAND4 (N12771, N12769, N403, N9822, N11563);
nor NOR4 (N12772, N12753, N10193, N2096, N5036);
or OR2 (N12773, N12742, N9093);
or OR4 (N12774, N12722, N4504, N8305, N8240);
buf BUF1 (N12775, N12755);
or OR4 (N12776, N12771, N2269, N6575, N2200);
nor NOR4 (N12777, N12767, N2449, N11016, N9709);
buf BUF1 (N12778, N12770);
not NOT1 (N12779, N12776);
xor XOR2 (N12780, N12772, N7989);
and AND3 (N12781, N12778, N997, N8253);
nand NAND4 (N12782, N12773, N9302, N6098, N6530);
buf BUF1 (N12783, N12779);
buf BUF1 (N12784, N12783);
nor NOR2 (N12785, N12777, N1153);
buf BUF1 (N12786, N12763);
not NOT1 (N12787, N12758);
nor NOR2 (N12788, N12774, N11191);
buf BUF1 (N12789, N12787);
and AND4 (N12790, N12788, N2750, N7627, N2421);
nand NAND2 (N12791, N12790, N11909);
not NOT1 (N12792, N12789);
buf BUF1 (N12793, N12791);
buf BUF1 (N12794, N12775);
nor NOR4 (N12795, N12785, N1159, N438, N5625);
or OR2 (N12796, N12794, N3910);
buf BUF1 (N12797, N12781);
or OR4 (N12798, N12757, N5609, N3961, N11780);
nand NAND2 (N12799, N12780, N12087);
or OR3 (N12800, N12793, N8340, N5857);
nand NAND2 (N12801, N12797, N10177);
or OR2 (N12802, N12782, N6689);
buf BUF1 (N12803, N12796);
nor NOR2 (N12804, N12798, N11343);
buf BUF1 (N12805, N12792);
nand NAND3 (N12806, N12799, N4083, N101);
nor NOR2 (N12807, N12800, N11628);
xor XOR2 (N12808, N12801, N8093);
nor NOR3 (N12809, N12804, N11460, N1180);
or OR4 (N12810, N12802, N9764, N3096, N8402);
nand NAND3 (N12811, N12806, N3387, N11661);
and AND4 (N12812, N12811, N11813, N5434, N10799);
not NOT1 (N12813, N12807);
and AND2 (N12814, N12803, N2198);
not NOT1 (N12815, N12812);
not NOT1 (N12816, N12805);
and AND2 (N12817, N12808, N10886);
and AND2 (N12818, N12817, N8819);
not NOT1 (N12819, N12816);
nor NOR3 (N12820, N12810, N7722, N4030);
not NOT1 (N12821, N12809);
or OR4 (N12822, N12819, N7980, N1259, N10837);
or OR3 (N12823, N12820, N8965, N5046);
not NOT1 (N12824, N12814);
or OR4 (N12825, N12824, N801, N12505, N730);
nor NOR3 (N12826, N12821, N5819, N688);
nor NOR4 (N12827, N12786, N4488, N1833, N3692);
nand NAND4 (N12828, N12822, N10206, N9527, N8739);
nand NAND2 (N12829, N12825, N3002);
not NOT1 (N12830, N12795);
and AND3 (N12831, N12813, N6749, N464);
nor NOR2 (N12832, N12829, N1502);
buf BUF1 (N12833, N12818);
nor NOR2 (N12834, N12832, N1363);
or OR2 (N12835, N12815, N3924);
and AND3 (N12836, N12823, N2521, N5555);
nand NAND2 (N12837, N12826, N7613);
nor NOR2 (N12838, N12836, N2148);
buf BUF1 (N12839, N12828);
nor NOR2 (N12840, N12834, N8982);
buf BUF1 (N12841, N12840);
buf BUF1 (N12842, N12837);
buf BUF1 (N12843, N12827);
nor NOR4 (N12844, N12843, N4325, N7445, N4393);
buf BUF1 (N12845, N12841);
xor XOR2 (N12846, N12835, N10951);
or OR2 (N12847, N12844, N12291);
nand NAND2 (N12848, N12839, N6447);
not NOT1 (N12849, N12845);
xor XOR2 (N12850, N12849, N1860);
and AND4 (N12851, N12842, N9112, N5810, N10027);
not NOT1 (N12852, N12831);
not NOT1 (N12853, N12830);
not NOT1 (N12854, N12851);
or OR4 (N12855, N12852, N10117, N2277, N12621);
buf BUF1 (N12856, N12853);
and AND4 (N12857, N12847, N8367, N1121, N5810);
not NOT1 (N12858, N12856);
or OR3 (N12859, N12833, N4557, N7526);
nor NOR3 (N12860, N12857, N6465, N1642);
nand NAND3 (N12861, N12859, N12000, N4648);
nor NOR4 (N12862, N12858, N7239, N1767, N6056);
not NOT1 (N12863, N12860);
not NOT1 (N12864, N12855);
nor NOR4 (N12865, N12848, N4425, N9324, N5022);
not NOT1 (N12866, N12865);
not NOT1 (N12867, N12863);
nand NAND3 (N12868, N12838, N1419, N610);
not NOT1 (N12869, N12868);
nor NOR3 (N12870, N12862, N2641, N896);
nor NOR3 (N12871, N12864, N5650, N5108);
and AND3 (N12872, N12866, N8113, N554);
nor NOR4 (N12873, N12861, N5629, N3373, N11580);
or OR3 (N12874, N12873, N4204, N3577);
buf BUF1 (N12875, N12846);
or OR3 (N12876, N12784, N7251, N5956);
xor XOR2 (N12877, N12869, N7172);
not NOT1 (N12878, N12876);
buf BUF1 (N12879, N12874);
buf BUF1 (N12880, N12879);
nand NAND2 (N12881, N12880, N4494);
buf BUF1 (N12882, N12881);
or OR4 (N12883, N12882, N7960, N6379, N3542);
nor NOR3 (N12884, N12867, N8563, N4758);
xor XOR2 (N12885, N12872, N10804);
nand NAND2 (N12886, N12883, N1472);
xor XOR2 (N12887, N12870, N1692);
not NOT1 (N12888, N12875);
nor NOR4 (N12889, N12878, N11116, N11349, N11015);
and AND2 (N12890, N12854, N2153);
not NOT1 (N12891, N12890);
and AND4 (N12892, N12884, N11214, N8114, N759);
buf BUF1 (N12893, N12891);
not NOT1 (N12894, N12889);
buf BUF1 (N12895, N12893);
nor NOR3 (N12896, N12886, N6553, N10480);
xor XOR2 (N12897, N12850, N6382);
and AND2 (N12898, N12877, N12090);
not NOT1 (N12899, N12898);
xor XOR2 (N12900, N12887, N9987);
nor NOR4 (N12901, N12871, N10481, N7074, N4257);
or OR4 (N12902, N12901, N244, N10243, N10951);
and AND2 (N12903, N12892, N9677);
and AND3 (N12904, N12894, N7539, N10850);
buf BUF1 (N12905, N12895);
buf BUF1 (N12906, N12888);
and AND4 (N12907, N12885, N9438, N167, N1120);
buf BUF1 (N12908, N12900);
not NOT1 (N12909, N12899);
or OR2 (N12910, N12908, N4660);
xor XOR2 (N12911, N12909, N4823);
and AND2 (N12912, N12904, N9636);
xor XOR2 (N12913, N12910, N1478);
xor XOR2 (N12914, N12905, N873);
buf BUF1 (N12915, N12914);
not NOT1 (N12916, N12913);
xor XOR2 (N12917, N12916, N10310);
and AND2 (N12918, N12906, N10234);
buf BUF1 (N12919, N12918);
and AND2 (N12920, N12917, N4513);
and AND3 (N12921, N12907, N2638, N1658);
nand NAND4 (N12922, N12920, N9288, N4745, N10372);
and AND4 (N12923, N12912, N1153, N10443, N2276);
not NOT1 (N12924, N12921);
or OR2 (N12925, N12897, N7505);
nor NOR3 (N12926, N12896, N487, N7833);
nand NAND2 (N12927, N12926, N3510);
or OR4 (N12928, N12927, N103, N1958, N7887);
or OR3 (N12929, N12919, N10795, N5961);
buf BUF1 (N12930, N12925);
nor NOR2 (N12931, N12915, N10259);
nand NAND2 (N12932, N12902, N1449);
xor XOR2 (N12933, N12932, N5316);
xor XOR2 (N12934, N12931, N11574);
buf BUF1 (N12935, N12911);
or OR4 (N12936, N12930, N7009, N11764, N4352);
not NOT1 (N12937, N12933);
xor XOR2 (N12938, N12924, N2897);
or OR3 (N12939, N12929, N124, N7503);
not NOT1 (N12940, N12935);
or OR3 (N12941, N12936, N7851, N6409);
nand NAND3 (N12942, N12940, N5325, N1450);
not NOT1 (N12943, N12934);
buf BUF1 (N12944, N12923);
nor NOR3 (N12945, N12941, N6327, N10454);
buf BUF1 (N12946, N12928);
and AND3 (N12947, N12939, N6130, N8348);
nand NAND4 (N12948, N12938, N6016, N6080, N8569);
or OR4 (N12949, N12946, N6022, N4406, N2938);
and AND3 (N12950, N12945, N3257, N3512);
nand NAND4 (N12951, N12942, N2869, N12861, N11845);
and AND3 (N12952, N12943, N10536, N8342);
nor NOR2 (N12953, N12944, N10399);
nand NAND2 (N12954, N12953, N3484);
or OR3 (N12955, N12947, N1423, N11571);
nand NAND4 (N12956, N12937, N253, N5396, N1439);
buf BUF1 (N12957, N12955);
and AND3 (N12958, N12922, N12888, N5884);
buf BUF1 (N12959, N12958);
or OR3 (N12960, N12948, N12866, N4656);
not NOT1 (N12961, N12903);
nand NAND3 (N12962, N12961, N8403, N12911);
not NOT1 (N12963, N12957);
nor NOR4 (N12964, N12952, N1314, N10987, N3759);
or OR4 (N12965, N12960, N10489, N31, N3733);
or OR3 (N12966, N12951, N10363, N12064);
or OR2 (N12967, N12962, N4077);
nand NAND2 (N12968, N12949, N7201);
nand NAND3 (N12969, N12966, N2286, N7378);
buf BUF1 (N12970, N12963);
or OR2 (N12971, N12967, N8032);
and AND3 (N12972, N12964, N3754, N2074);
nand NAND4 (N12973, N12970, N6515, N2887, N10832);
and AND3 (N12974, N12950, N1939, N6497);
not NOT1 (N12975, N12971);
and AND4 (N12976, N12969, N4824, N1874, N1125);
not NOT1 (N12977, N12956);
or OR4 (N12978, N12974, N2407, N5235, N6532);
or OR2 (N12979, N12975, N7109);
not NOT1 (N12980, N12977);
nand NAND2 (N12981, N12968, N9857);
buf BUF1 (N12982, N12965);
or OR3 (N12983, N12979, N5818, N284);
not NOT1 (N12984, N12983);
nor NOR4 (N12985, N12978, N2921, N733, N840);
or OR3 (N12986, N12954, N11020, N6789);
xor XOR2 (N12987, N12982, N9234);
and AND3 (N12988, N12980, N6290, N11684);
or OR2 (N12989, N12959, N8716);
buf BUF1 (N12990, N12988);
and AND2 (N12991, N12985, N8991);
and AND3 (N12992, N12984, N4260, N6355);
nand NAND2 (N12993, N12973, N10209);
xor XOR2 (N12994, N12981, N1593);
nand NAND2 (N12995, N12972, N1973);
and AND3 (N12996, N12991, N3124, N352);
and AND4 (N12997, N12993, N4735, N4030, N5893);
xor XOR2 (N12998, N12995, N5760);
and AND2 (N12999, N12987, N5405);
nand NAND2 (N13000, N12989, N2332);
or OR3 (N13001, N13000, N10761, N3560);
buf BUF1 (N13002, N12996);
buf BUF1 (N13003, N12994);
not NOT1 (N13004, N13001);
buf BUF1 (N13005, N12986);
and AND3 (N13006, N13004, N9766, N8030);
and AND4 (N13007, N13006, N434, N8261, N10734);
nand NAND3 (N13008, N12998, N920, N9415);
not NOT1 (N13009, N13003);
nor NOR2 (N13010, N13005, N235);
nand NAND3 (N13011, N12976, N2454, N8180);
not NOT1 (N13012, N12999);
xor XOR2 (N13013, N13010, N10451);
buf BUF1 (N13014, N13008);
nand NAND2 (N13015, N13014, N1199);
xor XOR2 (N13016, N13011, N11396);
or OR2 (N13017, N12990, N2803);
xor XOR2 (N13018, N12997, N8849);
xor XOR2 (N13019, N13016, N11724);
buf BUF1 (N13020, N13015);
nor NOR2 (N13021, N13002, N7141);
buf BUF1 (N13022, N13021);
nand NAND4 (N13023, N13012, N11667, N2609, N11173);
buf BUF1 (N13024, N13019);
xor XOR2 (N13025, N13013, N3738);
xor XOR2 (N13026, N13017, N1156);
nand NAND3 (N13027, N13022, N5955, N978);
nor NOR3 (N13028, N12992, N7796, N6598);
nor NOR4 (N13029, N13024, N680, N6325, N5801);
and AND2 (N13030, N13009, N5662);
nand NAND3 (N13031, N13029, N9086, N8345);
and AND4 (N13032, N13007, N6070, N1628, N2165);
not NOT1 (N13033, N13020);
nor NOR3 (N13034, N13027, N4542, N9155);
not NOT1 (N13035, N13025);
xor XOR2 (N13036, N13023, N4146);
buf BUF1 (N13037, N13018);
buf BUF1 (N13038, N13036);
nand NAND4 (N13039, N13033, N11601, N6921, N2446);
or OR2 (N13040, N13039, N7454);
or OR2 (N13041, N13032, N3310);
nand NAND2 (N13042, N13035, N2276);
buf BUF1 (N13043, N13040);
not NOT1 (N13044, N13041);
nand NAND2 (N13045, N13034, N2415);
not NOT1 (N13046, N13028);
buf BUF1 (N13047, N13026);
and AND3 (N13048, N13038, N2546, N12230);
xor XOR2 (N13049, N13042, N564);
and AND4 (N13050, N13049, N6828, N11119, N1726);
buf BUF1 (N13051, N13047);
not NOT1 (N13052, N13048);
nor NOR3 (N13053, N13050, N7150, N2783);
buf BUF1 (N13054, N13044);
xor XOR2 (N13055, N13054, N9707);
xor XOR2 (N13056, N13053, N781);
nor NOR2 (N13057, N13031, N8125);
or OR3 (N13058, N13037, N10938, N3382);
not NOT1 (N13059, N13051);
buf BUF1 (N13060, N13056);
nand NAND3 (N13061, N13057, N10783, N8274);
nor NOR4 (N13062, N13060, N10038, N9808, N7783);
not NOT1 (N13063, N13055);
buf BUF1 (N13064, N13063);
nor NOR4 (N13065, N13046, N6015, N2474, N5137);
xor XOR2 (N13066, N13043, N3941);
or OR4 (N13067, N13030, N361, N9577, N10997);
or OR3 (N13068, N13058, N7198, N12152);
xor XOR2 (N13069, N13066, N7941);
nand NAND2 (N13070, N13067, N10649);
or OR3 (N13071, N13069, N5042, N6447);
and AND2 (N13072, N13065, N1777);
nor NOR2 (N13073, N13052, N9260);
xor XOR2 (N13074, N13064, N8502);
not NOT1 (N13075, N13070);
buf BUF1 (N13076, N13061);
or OR2 (N13077, N13045, N9409);
nor NOR4 (N13078, N13071, N6998, N171, N11772);
buf BUF1 (N13079, N13077);
not NOT1 (N13080, N13068);
and AND4 (N13081, N13080, N2813, N1061, N140);
and AND4 (N13082, N13072, N9603, N10997, N4962);
nor NOR3 (N13083, N13079, N7378, N6573);
not NOT1 (N13084, N13076);
nand NAND3 (N13085, N13081, N12778, N3535);
or OR4 (N13086, N13073, N2434, N8343, N10419);
not NOT1 (N13087, N13059);
nand NAND3 (N13088, N13086, N4417, N6845);
buf BUF1 (N13089, N13078);
or OR4 (N13090, N13084, N11785, N10704, N2693);
not NOT1 (N13091, N13074);
and AND3 (N13092, N13085, N12102, N7369);
nand NAND2 (N13093, N13089, N3265);
or OR2 (N13094, N13083, N4428);
and AND3 (N13095, N13088, N5015, N3973);
nor NOR2 (N13096, N13090, N6734);
buf BUF1 (N13097, N13087);
nor NOR3 (N13098, N13075, N466, N4987);
xor XOR2 (N13099, N13082, N6454);
not NOT1 (N13100, N13099);
not NOT1 (N13101, N13100);
or OR2 (N13102, N13098, N3304);
and AND4 (N13103, N13095, N12795, N5338, N3418);
not NOT1 (N13104, N13093);
nor NOR2 (N13105, N13097, N12538);
not NOT1 (N13106, N13091);
nor NOR4 (N13107, N13101, N7679, N862, N5585);
xor XOR2 (N13108, N13105, N5875);
nor NOR2 (N13109, N13094, N9213);
and AND2 (N13110, N13104, N1583);
or OR2 (N13111, N13109, N11437);
or OR2 (N13112, N13103, N432);
or OR4 (N13113, N13111, N4420, N9581, N5009);
nand NAND2 (N13114, N13102, N11290);
not NOT1 (N13115, N13096);
not NOT1 (N13116, N13106);
nor NOR2 (N13117, N13062, N8446);
and AND4 (N13118, N13107, N9386, N9753, N3833);
and AND3 (N13119, N13108, N11357, N5548);
nand NAND4 (N13120, N13110, N12235, N75, N6909);
nand NAND4 (N13121, N13115, N7935, N4274, N8435);
nor NOR4 (N13122, N13113, N5302, N6072, N83);
xor XOR2 (N13123, N13117, N3402);
xor XOR2 (N13124, N13122, N9426);
nor NOR2 (N13125, N13116, N11037);
buf BUF1 (N13126, N13092);
or OR4 (N13127, N13114, N1289, N522, N10608);
and AND4 (N13128, N13124, N262, N10750, N6234);
not NOT1 (N13129, N13123);
xor XOR2 (N13130, N13121, N12200);
buf BUF1 (N13131, N13118);
nor NOR3 (N13132, N13119, N8374, N11048);
or OR2 (N13133, N13131, N12273);
nand NAND4 (N13134, N13112, N10680, N4692, N12870);
nor NOR4 (N13135, N13125, N10862, N651, N4973);
nor NOR3 (N13136, N13133, N1801, N8361);
buf BUF1 (N13137, N13127);
or OR2 (N13138, N13130, N6346);
nand NAND2 (N13139, N13126, N12294);
xor XOR2 (N13140, N13139, N6547);
xor XOR2 (N13141, N13135, N8662);
or OR3 (N13142, N13141, N3793, N2384);
xor XOR2 (N13143, N13128, N7726);
xor XOR2 (N13144, N13120, N2768);
and AND4 (N13145, N13142, N11074, N5067, N2582);
xor XOR2 (N13146, N13138, N3926);
xor XOR2 (N13147, N13140, N11780);
xor XOR2 (N13148, N13144, N8048);
nor NOR3 (N13149, N13136, N6616, N12807);
or OR4 (N13150, N13148, N6187, N7557, N4796);
nand NAND3 (N13151, N13137, N2917, N1322);
and AND4 (N13152, N13149, N11234, N6571, N2248);
not NOT1 (N13153, N13134);
nor NOR2 (N13154, N13132, N9863);
xor XOR2 (N13155, N13151, N5738);
or OR2 (N13156, N13129, N1424);
not NOT1 (N13157, N13145);
nor NOR3 (N13158, N13150, N4897, N10596);
and AND3 (N13159, N13143, N8810, N2342);
nor NOR2 (N13160, N13153, N8623);
buf BUF1 (N13161, N13146);
and AND3 (N13162, N13161, N4398, N11336);
not NOT1 (N13163, N13158);
nand NAND2 (N13164, N13155, N8924);
nand NAND4 (N13165, N13156, N1666, N4307, N12883);
xor XOR2 (N13166, N13163, N6627);
buf BUF1 (N13167, N13164);
not NOT1 (N13168, N13162);
nand NAND3 (N13169, N13165, N10207, N6635);
or OR2 (N13170, N13169, N473);
or OR2 (N13171, N13152, N10714);
xor XOR2 (N13172, N13159, N12834);
not NOT1 (N13173, N13171);
nand NAND4 (N13174, N13157, N599, N896, N2339);
xor XOR2 (N13175, N13160, N10844);
not NOT1 (N13176, N13173);
not NOT1 (N13177, N13175);
nand NAND2 (N13178, N13177, N5398);
and AND2 (N13179, N13176, N8486);
and AND4 (N13180, N13168, N6756, N2868, N5786);
xor XOR2 (N13181, N13166, N8118);
and AND3 (N13182, N13178, N9441, N7962);
nor NOR3 (N13183, N13170, N355, N2313);
and AND3 (N13184, N13172, N9962, N10522);
xor XOR2 (N13185, N13179, N6788);
nor NOR4 (N13186, N13147, N12530, N7067, N2634);
buf BUF1 (N13187, N13183);
nor NOR2 (N13188, N13184, N2267);
xor XOR2 (N13189, N13154, N11657);
or OR3 (N13190, N13186, N12639, N8690);
not NOT1 (N13191, N13187);
not NOT1 (N13192, N13191);
not NOT1 (N13193, N13182);
or OR4 (N13194, N13180, N3743, N12895, N6263);
nand NAND2 (N13195, N13192, N6755);
and AND3 (N13196, N13188, N8472, N8887);
not NOT1 (N13197, N13185);
xor XOR2 (N13198, N13174, N3630);
nor NOR4 (N13199, N13193, N9126, N1792, N6235);
nand NAND2 (N13200, N13196, N10034);
buf BUF1 (N13201, N13190);
or OR2 (N13202, N13189, N9044);
or OR4 (N13203, N13194, N7246, N10995, N1650);
nor NOR3 (N13204, N13200, N2061, N8784);
or OR2 (N13205, N13198, N12976);
and AND2 (N13206, N13203, N3665);
xor XOR2 (N13207, N13195, N1859);
or OR4 (N13208, N13167, N245, N12394, N11491);
nand NAND4 (N13209, N13199, N7839, N8246, N9300);
nand NAND2 (N13210, N13207, N737);
nor NOR4 (N13211, N13181, N10649, N4724, N1959);
nor NOR2 (N13212, N13204, N1966);
buf BUF1 (N13213, N13205);
nor NOR3 (N13214, N13202, N3258, N8653);
nand NAND2 (N13215, N13213, N11535);
nand NAND2 (N13216, N13211, N2786);
or OR3 (N13217, N13208, N4798, N513);
not NOT1 (N13218, N13217);
buf BUF1 (N13219, N13197);
nor NOR3 (N13220, N13216, N3438, N908);
not NOT1 (N13221, N13206);
and AND2 (N13222, N13215, N5097);
buf BUF1 (N13223, N13222);
or OR4 (N13224, N13220, N3406, N1430, N11252);
not NOT1 (N13225, N13210);
xor XOR2 (N13226, N13214, N1152);
nand NAND3 (N13227, N13209, N6316, N9134);
nand NAND3 (N13228, N13224, N7511, N1689);
and AND3 (N13229, N13221, N5029, N12465);
buf BUF1 (N13230, N13201);
nor NOR4 (N13231, N13212, N12726, N2224, N12470);
buf BUF1 (N13232, N13219);
or OR2 (N13233, N13225, N10809);
xor XOR2 (N13234, N13233, N8482);
nand NAND4 (N13235, N13232, N11791, N3284, N6824);
buf BUF1 (N13236, N13230);
nor NOR4 (N13237, N13228, N1748, N4204, N7957);
or OR2 (N13238, N13226, N9158);
xor XOR2 (N13239, N13229, N5087);
not NOT1 (N13240, N13223);
buf BUF1 (N13241, N13237);
and AND2 (N13242, N13231, N5937);
xor XOR2 (N13243, N13240, N62);
not NOT1 (N13244, N13236);
not NOT1 (N13245, N13244);
and AND2 (N13246, N13245, N2470);
buf BUF1 (N13247, N13241);
nor NOR2 (N13248, N13243, N7808);
buf BUF1 (N13249, N13239);
and AND2 (N13250, N13248, N8554);
buf BUF1 (N13251, N13249);
xor XOR2 (N13252, N13227, N6517);
not NOT1 (N13253, N13246);
xor XOR2 (N13254, N13235, N2866);
and AND4 (N13255, N13242, N2847, N7433, N8163);
and AND4 (N13256, N13251, N1122, N9274, N8747);
not NOT1 (N13257, N13252);
xor XOR2 (N13258, N13250, N2741);
not NOT1 (N13259, N13238);
xor XOR2 (N13260, N13256, N11231);
and AND4 (N13261, N13247, N9127, N4244, N9694);
xor XOR2 (N13262, N13260, N6776);
and AND3 (N13263, N13259, N7764, N12613);
or OR2 (N13264, N13255, N5189);
xor XOR2 (N13265, N13218, N2043);
or OR2 (N13266, N13263, N9812);
or OR2 (N13267, N13261, N12122);
and AND3 (N13268, N13262, N1600, N5037);
and AND4 (N13269, N13266, N9847, N7868, N6671);
nand NAND3 (N13270, N13253, N3420, N11027);
buf BUF1 (N13271, N13258);
nand NAND2 (N13272, N13268, N7378);
buf BUF1 (N13273, N13270);
not NOT1 (N13274, N13265);
buf BUF1 (N13275, N13234);
buf BUF1 (N13276, N13275);
or OR2 (N13277, N13272, N9833);
nor NOR3 (N13278, N13276, N4961, N3621);
nor NOR2 (N13279, N13271, N12969);
xor XOR2 (N13280, N13277, N2134);
xor XOR2 (N13281, N13264, N12731);
xor XOR2 (N13282, N13278, N13227);
buf BUF1 (N13283, N13269);
not NOT1 (N13284, N13257);
buf BUF1 (N13285, N13282);
or OR4 (N13286, N13285, N5796, N11012, N10346);
xor XOR2 (N13287, N13274, N2662);
xor XOR2 (N13288, N13254, N108);
nor NOR2 (N13289, N13280, N502);
or OR3 (N13290, N13281, N8975, N11723);
xor XOR2 (N13291, N13273, N2489);
and AND3 (N13292, N13286, N9536, N7284);
nor NOR3 (N13293, N13279, N3428, N3176);
and AND4 (N13294, N13289, N2466, N10188, N2011);
buf BUF1 (N13295, N13294);
buf BUF1 (N13296, N13288);
nand NAND3 (N13297, N13287, N3941, N10455);
nor NOR4 (N13298, N13295, N1419, N4553, N1271);
buf BUF1 (N13299, N13298);
or OR3 (N13300, N13293, N5738, N7014);
not NOT1 (N13301, N13267);
xor XOR2 (N13302, N13296, N2167);
and AND4 (N13303, N13300, N7865, N8667, N11234);
or OR2 (N13304, N13303, N3970);
not NOT1 (N13305, N13290);
or OR2 (N13306, N13305, N3457);
buf BUF1 (N13307, N13284);
nor NOR2 (N13308, N13292, N4352);
not NOT1 (N13309, N13297);
or OR4 (N13310, N13291, N2829, N11390, N6868);
nor NOR3 (N13311, N13309, N11980, N728);
and AND3 (N13312, N13301, N11746, N392);
or OR3 (N13313, N13312, N8370, N2208);
nor NOR2 (N13314, N13283, N10616);
xor XOR2 (N13315, N13304, N9049);
and AND4 (N13316, N13299, N8658, N8096, N7313);
nor NOR4 (N13317, N13307, N7235, N9313, N4687);
and AND2 (N13318, N13310, N12169);
nand NAND4 (N13319, N13314, N11404, N10448, N1615);
or OR4 (N13320, N13302, N664, N1258, N3293);
nand NAND4 (N13321, N13315, N6075, N11468, N3506);
and AND4 (N13322, N13320, N9468, N4667, N8896);
or OR2 (N13323, N13311, N2825);
nor NOR3 (N13324, N13317, N3395, N520);
buf BUF1 (N13325, N13316);
not NOT1 (N13326, N13321);
nor NOR2 (N13327, N13313, N4284);
and AND3 (N13328, N13326, N2086, N4486);
xor XOR2 (N13329, N13327, N5729);
nor NOR3 (N13330, N13306, N5843, N8215);
nor NOR4 (N13331, N13329, N9319, N11711, N6818);
not NOT1 (N13332, N13331);
nor NOR4 (N13333, N13318, N6379, N10697, N2084);
buf BUF1 (N13334, N13328);
nand NAND3 (N13335, N13334, N6538, N8856);
nor NOR4 (N13336, N13324, N9516, N13118, N279);
not NOT1 (N13337, N13325);
and AND4 (N13338, N13332, N6954, N5691, N12059);
or OR2 (N13339, N13323, N2474);
or OR2 (N13340, N13308, N4281);
or OR2 (N13341, N13338, N7546);
and AND3 (N13342, N13337, N10809, N10833);
not NOT1 (N13343, N13335);
not NOT1 (N13344, N13333);
buf BUF1 (N13345, N13340);
or OR3 (N13346, N13344, N8833, N5166);
and AND3 (N13347, N13343, N2512, N4227);
and AND3 (N13348, N13347, N5780, N169);
or OR2 (N13349, N13346, N541);
nand NAND3 (N13350, N13345, N4607, N11644);
nor NOR4 (N13351, N13322, N480, N3364, N9607);
xor XOR2 (N13352, N13350, N2324);
xor XOR2 (N13353, N13351, N7529);
or OR2 (N13354, N13330, N9067);
nor NOR4 (N13355, N13354, N13329, N5428, N2438);
nor NOR2 (N13356, N13352, N6729);
nor NOR4 (N13357, N13353, N11418, N10778, N6121);
buf BUF1 (N13358, N13341);
nor NOR3 (N13359, N13348, N12447, N10732);
and AND3 (N13360, N13342, N1594, N9789);
and AND3 (N13361, N13339, N5144, N536);
and AND2 (N13362, N13359, N4418);
and AND4 (N13363, N13349, N1253, N11770, N8579);
xor XOR2 (N13364, N13336, N4505);
nand NAND2 (N13365, N13358, N2656);
xor XOR2 (N13366, N13355, N3232);
buf BUF1 (N13367, N13366);
and AND3 (N13368, N13365, N7190, N9743);
and AND3 (N13369, N13357, N12701, N11440);
or OR3 (N13370, N13369, N6730, N1368);
or OR3 (N13371, N13356, N13110, N2558);
xor XOR2 (N13372, N13361, N5885);
xor XOR2 (N13373, N13363, N3232);
or OR3 (N13374, N13370, N8601, N9709);
nor NOR2 (N13375, N13373, N10521);
not NOT1 (N13376, N13374);
nor NOR3 (N13377, N13375, N950, N2596);
or OR4 (N13378, N13377, N12381, N12592, N12585);
not NOT1 (N13379, N13372);
xor XOR2 (N13380, N13368, N12170);
xor XOR2 (N13381, N13362, N4141);
not NOT1 (N13382, N13319);
buf BUF1 (N13383, N13380);
nand NAND4 (N13384, N13381, N5647, N7364, N4659);
nand NAND2 (N13385, N13367, N3800);
buf BUF1 (N13386, N13364);
buf BUF1 (N13387, N13386);
and AND4 (N13388, N13371, N12974, N3403, N7737);
nand NAND3 (N13389, N13387, N12944, N8498);
and AND4 (N13390, N13388, N4300, N8369, N3743);
nand NAND3 (N13391, N13390, N2867, N1392);
nand NAND2 (N13392, N13382, N10691);
nand NAND4 (N13393, N13383, N2726, N10821, N13);
buf BUF1 (N13394, N13384);
xor XOR2 (N13395, N13392, N6332);
nor NOR2 (N13396, N13360, N7233);
xor XOR2 (N13397, N13393, N2402);
or OR4 (N13398, N13385, N13044, N4577, N8905);
nand NAND4 (N13399, N13395, N13345, N7146, N8963);
and AND3 (N13400, N13391, N9750, N13145);
not NOT1 (N13401, N13396);
not NOT1 (N13402, N13378);
nand NAND2 (N13403, N13394, N6246);
buf BUF1 (N13404, N13401);
and AND4 (N13405, N13404, N5091, N8528, N6659);
and AND4 (N13406, N13403, N9928, N10490, N2363);
nor NOR4 (N13407, N13398, N6600, N2928, N6392);
or OR4 (N13408, N13399, N12092, N1692, N12899);
nor NOR2 (N13409, N13376, N9828);
and AND2 (N13410, N13397, N890);
or OR4 (N13411, N13409, N3958, N2721, N8941);
not NOT1 (N13412, N13407);
or OR4 (N13413, N13412, N355, N5064, N2207);
nand NAND3 (N13414, N13406, N3578, N718);
nand NAND3 (N13415, N13405, N985, N10021);
or OR2 (N13416, N13389, N1780);
or OR3 (N13417, N13400, N1139, N8354);
nor NOR2 (N13418, N13417, N6650);
not NOT1 (N13419, N13416);
xor XOR2 (N13420, N13379, N7357);
buf BUF1 (N13421, N13411);
nand NAND4 (N13422, N13421, N6090, N4995, N13098);
nand NAND2 (N13423, N13420, N6138);
buf BUF1 (N13424, N13402);
not NOT1 (N13425, N13422);
nor NOR2 (N13426, N13414, N11357);
or OR4 (N13427, N13410, N8591, N9431, N4272);
xor XOR2 (N13428, N13413, N2645);
and AND4 (N13429, N13408, N3781, N5684, N7969);
nor NOR4 (N13430, N13415, N10278, N10045, N202);
nand NAND2 (N13431, N13428, N1555);
and AND4 (N13432, N13418, N5448, N4131, N1671);
and AND4 (N13433, N13432, N1669, N6188, N9994);
not NOT1 (N13434, N13423);
and AND2 (N13435, N13427, N2431);
buf BUF1 (N13436, N13424);
nand NAND3 (N13437, N13429, N3165, N7742);
or OR4 (N13438, N13431, N10324, N2888, N6409);
and AND4 (N13439, N13435, N5237, N5009, N9980);
xor XOR2 (N13440, N13426, N10271);
nor NOR4 (N13441, N13430, N11386, N1540, N3648);
or OR4 (N13442, N13419, N8556, N12559, N1391);
and AND4 (N13443, N13433, N2565, N2748, N1292);
buf BUF1 (N13444, N13436);
nor NOR3 (N13445, N13440, N5856, N6906);
and AND4 (N13446, N13439, N5800, N2272, N10711);
nor NOR3 (N13447, N13441, N495, N1684);
or OR4 (N13448, N13444, N3360, N2542, N2231);
or OR4 (N13449, N13425, N9786, N5103, N2677);
and AND3 (N13450, N13448, N7301, N9603);
and AND2 (N13451, N13434, N12763);
not NOT1 (N13452, N13451);
and AND4 (N13453, N13437, N3041, N2055, N3545);
or OR4 (N13454, N13445, N10727, N10772, N9038);
or OR2 (N13455, N13454, N10063);
xor XOR2 (N13456, N13443, N8934);
nand NAND2 (N13457, N13456, N364);
and AND4 (N13458, N13446, N12192, N3754, N12921);
nor NOR3 (N13459, N13442, N8250, N7961);
and AND2 (N13460, N13455, N1905);
and AND2 (N13461, N13458, N10245);
not NOT1 (N13462, N13459);
nor NOR3 (N13463, N13457, N1087, N1802);
buf BUF1 (N13464, N13460);
xor XOR2 (N13465, N13453, N9271);
xor XOR2 (N13466, N13452, N9664);
buf BUF1 (N13467, N13461);
and AND2 (N13468, N13447, N7382);
and AND4 (N13469, N13462, N974, N10825, N5522);
xor XOR2 (N13470, N13468, N11747);
xor XOR2 (N13471, N13450, N5027);
and AND3 (N13472, N13463, N4231, N11092);
or OR2 (N13473, N13466, N5261);
and AND3 (N13474, N13449, N11531, N492);
not NOT1 (N13475, N13470);
and AND3 (N13476, N13469, N8010, N5044);
xor XOR2 (N13477, N13475, N715);
xor XOR2 (N13478, N13438, N1043);
and AND2 (N13479, N13477, N12836);
nor NOR4 (N13480, N13467, N4178, N2398, N12979);
nand NAND2 (N13481, N13480, N3975);
and AND2 (N13482, N13478, N5326);
buf BUF1 (N13483, N13481);
and AND3 (N13484, N13476, N247, N10252);
buf BUF1 (N13485, N13465);
not NOT1 (N13486, N13484);
or OR4 (N13487, N13485, N7377, N8355, N6287);
buf BUF1 (N13488, N13479);
not NOT1 (N13489, N13483);
not NOT1 (N13490, N13489);
nand NAND2 (N13491, N13464, N2632);
and AND3 (N13492, N13490, N12852, N6173);
nand NAND2 (N13493, N13471, N8402);
xor XOR2 (N13494, N13492, N6942);
nor NOR2 (N13495, N13487, N10327);
nor NOR3 (N13496, N13473, N9431, N11171);
nand NAND4 (N13497, N13482, N7176, N9065, N4942);
xor XOR2 (N13498, N13472, N1223);
and AND3 (N13499, N13496, N7405, N11333);
xor XOR2 (N13500, N13498, N10890);
buf BUF1 (N13501, N13494);
and AND4 (N13502, N13491, N6632, N11, N199);
nand NAND4 (N13503, N13495, N13369, N12167, N9808);
nor NOR4 (N13504, N13493, N4279, N294, N13252);
nand NAND4 (N13505, N13497, N5304, N6491, N9467);
and AND2 (N13506, N13504, N5862);
and AND2 (N13507, N13488, N8390);
nand NAND2 (N13508, N13503, N12719);
nor NOR3 (N13509, N13502, N11006, N7701);
and AND3 (N13510, N13506, N12616, N3363);
nand NAND2 (N13511, N13474, N8005);
nor NOR3 (N13512, N13510, N12872, N11066);
not NOT1 (N13513, N13486);
nand NAND2 (N13514, N13500, N6965);
not NOT1 (N13515, N13508);
nand NAND3 (N13516, N13514, N46, N7890);
not NOT1 (N13517, N13507);
buf BUF1 (N13518, N13515);
xor XOR2 (N13519, N13518, N4963);
not NOT1 (N13520, N13517);
xor XOR2 (N13521, N13519, N3454);
not NOT1 (N13522, N13505);
buf BUF1 (N13523, N13521);
xor XOR2 (N13524, N13501, N1966);
buf BUF1 (N13525, N13524);
xor XOR2 (N13526, N13522, N1573);
nand NAND2 (N13527, N13509, N9321);
nor NOR4 (N13528, N13513, N10583, N12558, N10739);
nor NOR2 (N13529, N13511, N12664);
buf BUF1 (N13530, N13527);
or OR2 (N13531, N13512, N4120);
not NOT1 (N13532, N13528);
or OR2 (N13533, N13531, N6454);
or OR3 (N13534, N13523, N12486, N4406);
nor NOR4 (N13535, N13533, N2776, N7852, N2053);
and AND3 (N13536, N13534, N1947, N5542);
nand NAND4 (N13537, N13529, N7235, N1802, N6012);
buf BUF1 (N13538, N13537);
buf BUF1 (N13539, N13536);
nor NOR2 (N13540, N13525, N10481);
xor XOR2 (N13541, N13526, N11766);
and AND4 (N13542, N13516, N6705, N12177, N6041);
buf BUF1 (N13543, N13542);
nor NOR3 (N13544, N13530, N11300, N4304);
nor NOR2 (N13545, N13539, N7878);
xor XOR2 (N13546, N13532, N5118);
not NOT1 (N13547, N13545);
nand NAND4 (N13548, N13543, N10704, N4089, N5614);
and AND3 (N13549, N13535, N10325, N5911);
not NOT1 (N13550, N13546);
nand NAND4 (N13551, N13547, N10545, N3120, N2452);
or OR2 (N13552, N13551, N7368);
or OR4 (N13553, N13549, N12710, N2890, N7619);
nand NAND4 (N13554, N13538, N7734, N12556, N8001);
buf BUF1 (N13555, N13552);
buf BUF1 (N13556, N13544);
nand NAND4 (N13557, N13550, N8532, N805, N7699);
nor NOR4 (N13558, N13554, N3814, N1757, N11677);
and AND2 (N13559, N13557, N10155);
not NOT1 (N13560, N13556);
buf BUF1 (N13561, N13555);
xor XOR2 (N13562, N13561, N10634);
xor XOR2 (N13563, N13540, N351);
buf BUF1 (N13564, N13559);
buf BUF1 (N13565, N13564);
buf BUF1 (N13566, N13499);
nand NAND4 (N13567, N13562, N1858, N5673, N9991);
or OR3 (N13568, N13567, N10077, N9976);
or OR3 (N13569, N13553, N7922, N11522);
nor NOR4 (N13570, N13560, N12267, N2922, N1715);
and AND3 (N13571, N13520, N13488, N1495);
nand NAND4 (N13572, N13558, N6182, N7122, N3799);
nor NOR3 (N13573, N13571, N7835, N6885);
nand NAND3 (N13574, N13570, N12233, N6561);
buf BUF1 (N13575, N13569);
not NOT1 (N13576, N13572);
buf BUF1 (N13577, N13574);
nand NAND4 (N13578, N13568, N10930, N4882, N5579);
and AND4 (N13579, N13565, N11055, N7619, N12584);
not NOT1 (N13580, N13566);
xor XOR2 (N13581, N13577, N2919);
or OR3 (N13582, N13581, N1802, N2018);
nand NAND4 (N13583, N13582, N5560, N790, N6721);
nor NOR4 (N13584, N13580, N9751, N745, N7127);
not NOT1 (N13585, N13548);
and AND3 (N13586, N13576, N7235, N7262);
or OR2 (N13587, N13585, N12911);
nand NAND4 (N13588, N13586, N5057, N4094, N8659);
or OR3 (N13589, N13541, N3922, N4954);
nor NOR4 (N13590, N13583, N7165, N1788, N13019);
xor XOR2 (N13591, N13587, N11547);
not NOT1 (N13592, N13563);
xor XOR2 (N13593, N13579, N912);
nor NOR3 (N13594, N13591, N11210, N11155);
and AND2 (N13595, N13590, N9208);
xor XOR2 (N13596, N13594, N5788);
and AND4 (N13597, N13589, N12739, N5591, N4742);
buf BUF1 (N13598, N13588);
not NOT1 (N13599, N13595);
nand NAND2 (N13600, N13596, N13270);
nor NOR2 (N13601, N13598, N13169);
xor XOR2 (N13602, N13578, N440);
xor XOR2 (N13603, N13599, N11637);
xor XOR2 (N13604, N13597, N3398);
buf BUF1 (N13605, N13600);
or OR4 (N13606, N13592, N7974, N417, N6094);
and AND2 (N13607, N13606, N7250);
nor NOR2 (N13608, N13573, N3290);
or OR2 (N13609, N13608, N13021);
nand NAND4 (N13610, N13609, N6382, N2059, N12000);
or OR2 (N13611, N13584, N5888);
and AND2 (N13612, N13604, N8979);
buf BUF1 (N13613, N13607);
and AND3 (N13614, N13603, N11416, N12483);
nand NAND4 (N13615, N13611, N13462, N8999, N388);
buf BUF1 (N13616, N13610);
nand NAND2 (N13617, N13616, N3703);
buf BUF1 (N13618, N13601);
buf BUF1 (N13619, N13614);
nand NAND2 (N13620, N13602, N8158);
nor NOR4 (N13621, N13619, N13544, N5913, N9892);
nor NOR4 (N13622, N13613, N9549, N9592, N8902);
nor NOR3 (N13623, N13620, N12838, N13447);
and AND2 (N13624, N13618, N9144);
buf BUF1 (N13625, N13624);
or OR4 (N13626, N13617, N11948, N2135, N5028);
not NOT1 (N13627, N13575);
nand NAND2 (N13628, N13625, N2806);
not NOT1 (N13629, N13626);
or OR2 (N13630, N13615, N9833);
buf BUF1 (N13631, N13629);
or OR2 (N13632, N13623, N7944);
nand NAND4 (N13633, N13630, N9411, N2902, N9017);
xor XOR2 (N13634, N13622, N7375);
nor NOR3 (N13635, N13605, N6140, N10143);
or OR2 (N13636, N13633, N10816);
xor XOR2 (N13637, N13636, N3022);
xor XOR2 (N13638, N13621, N5012);
nor NOR3 (N13639, N13634, N3550, N4383);
and AND4 (N13640, N13637, N4633, N10849, N4520);
buf BUF1 (N13641, N13593);
xor XOR2 (N13642, N13638, N8734);
xor XOR2 (N13643, N13612, N6295);
xor XOR2 (N13644, N13642, N8851);
buf BUF1 (N13645, N13643);
and AND4 (N13646, N13627, N8810, N625, N2540);
not NOT1 (N13647, N13641);
xor XOR2 (N13648, N13645, N5600);
or OR3 (N13649, N13640, N10205, N8047);
and AND4 (N13650, N13644, N3563, N11997, N12277);
buf BUF1 (N13651, N13628);
or OR3 (N13652, N13651, N7107, N8787);
and AND2 (N13653, N13648, N4379);
and AND2 (N13654, N13631, N13328);
nor NOR4 (N13655, N13652, N612, N1983, N2367);
or OR2 (N13656, N13655, N940);
nor NOR3 (N13657, N13639, N7074, N13475);
nand NAND2 (N13658, N13646, N12464);
nand NAND2 (N13659, N13657, N7618);
not NOT1 (N13660, N13658);
or OR2 (N13661, N13650, N6135);
nand NAND3 (N13662, N13632, N8719, N3909);
buf BUF1 (N13663, N13660);
not NOT1 (N13664, N13659);
nand NAND4 (N13665, N13635, N3967, N12635, N339);
nand NAND3 (N13666, N13662, N12039, N382);
xor XOR2 (N13667, N13649, N11473);
and AND2 (N13668, N13666, N7072);
nor NOR4 (N13669, N13663, N4859, N11809, N7540);
buf BUF1 (N13670, N13647);
nand NAND3 (N13671, N13664, N4746, N2513);
xor XOR2 (N13672, N13670, N80);
or OR3 (N13673, N13654, N13480, N8517);
xor XOR2 (N13674, N13672, N2557);
not NOT1 (N13675, N13665);
not NOT1 (N13676, N13661);
and AND2 (N13677, N13673, N12078);
and AND3 (N13678, N13677, N6283, N9413);
and AND3 (N13679, N13675, N6040, N11499);
nand NAND2 (N13680, N13653, N11955);
nand NAND3 (N13681, N13679, N2080, N3263);
or OR4 (N13682, N13681, N5156, N12409, N5348);
nor NOR2 (N13683, N13668, N5454);
not NOT1 (N13684, N13682);
buf BUF1 (N13685, N13674);
nor NOR4 (N13686, N13685, N6392, N4358, N1051);
or OR3 (N13687, N13667, N10506, N3052);
and AND3 (N13688, N13680, N6584, N2819);
nor NOR3 (N13689, N13684, N2390, N8654);
not NOT1 (N13690, N13687);
not NOT1 (N13691, N13656);
not NOT1 (N13692, N13676);
and AND3 (N13693, N13689, N10912, N7520);
and AND4 (N13694, N13693, N7620, N212, N3509);
nand NAND4 (N13695, N13686, N3241, N3536, N5244);
or OR4 (N13696, N13694, N7225, N4479, N8093);
nand NAND4 (N13697, N13691, N256, N12367, N2625);
buf BUF1 (N13698, N13678);
xor XOR2 (N13699, N13698, N10966);
and AND2 (N13700, N13699, N1657);
and AND2 (N13701, N13700, N10389);
not NOT1 (N13702, N13671);
nor NOR4 (N13703, N13690, N9689, N10067, N11681);
or OR2 (N13704, N13702, N1977);
buf BUF1 (N13705, N13683);
xor XOR2 (N13706, N13669, N6705);
xor XOR2 (N13707, N13692, N6302);
buf BUF1 (N13708, N13704);
xor XOR2 (N13709, N13695, N2314);
xor XOR2 (N13710, N13703, N12813);
or OR2 (N13711, N13696, N5507);
and AND2 (N13712, N13711, N3292);
not NOT1 (N13713, N13710);
nor NOR4 (N13714, N13709, N10697, N1633, N7657);
or OR3 (N13715, N13714, N11755, N3927);
or OR2 (N13716, N13707, N5807);
xor XOR2 (N13717, N13706, N8836);
buf BUF1 (N13718, N13715);
buf BUF1 (N13719, N13718);
buf BUF1 (N13720, N13708);
buf BUF1 (N13721, N13716);
or OR3 (N13722, N13697, N9005, N7305);
nand NAND4 (N13723, N13722, N7034, N3952, N2667);
and AND4 (N13724, N13705, N1834, N3420, N5836);
and AND3 (N13725, N13720, N893, N7665);
and AND4 (N13726, N13721, N2636, N5018, N915);
or OR2 (N13727, N13701, N2338);
nand NAND3 (N13728, N13726, N13656, N2292);
and AND4 (N13729, N13728, N8477, N10726, N11065);
not NOT1 (N13730, N13713);
or OR2 (N13731, N13688, N4769);
or OR4 (N13732, N13731, N12074, N11358, N6000);
or OR3 (N13733, N13712, N11796, N1722);
xor XOR2 (N13734, N13719, N3617);
and AND4 (N13735, N13733, N11871, N2134, N2514);
nor NOR2 (N13736, N13729, N7098);
nand NAND4 (N13737, N13735, N3864, N10727, N10910);
and AND4 (N13738, N13737, N4315, N6190, N1429);
xor XOR2 (N13739, N13734, N3278);
nand NAND4 (N13740, N13732, N13091, N6930, N12703);
buf BUF1 (N13741, N13727);
buf BUF1 (N13742, N13736);
not NOT1 (N13743, N13730);
not NOT1 (N13744, N13717);
or OR2 (N13745, N13740, N7684);
and AND3 (N13746, N13741, N5047, N7683);
and AND4 (N13747, N13723, N13175, N9783, N2919);
buf BUF1 (N13748, N13744);
buf BUF1 (N13749, N13747);
nor NOR4 (N13750, N13745, N8442, N1268, N463);
or OR3 (N13751, N13746, N12224, N4267);
and AND3 (N13752, N13738, N5796, N11753);
buf BUF1 (N13753, N13743);
or OR4 (N13754, N13750, N2797, N10902, N1191);
and AND2 (N13755, N13739, N8084);
xor XOR2 (N13756, N13754, N3348);
or OR2 (N13757, N13748, N2690);
or OR2 (N13758, N13742, N11795);
and AND4 (N13759, N13753, N3996, N11558, N12561);
xor XOR2 (N13760, N13757, N5121);
not NOT1 (N13761, N13749);
or OR2 (N13762, N13752, N8265);
nand NAND4 (N13763, N13762, N13602, N378, N7204);
nand NAND2 (N13764, N13761, N5477);
or OR2 (N13765, N13759, N3798);
xor XOR2 (N13766, N13764, N5717);
or OR4 (N13767, N13756, N9009, N4748, N10352);
or OR3 (N13768, N13763, N5113, N3478);
not NOT1 (N13769, N13760);
buf BUF1 (N13770, N13755);
not NOT1 (N13771, N13765);
nor NOR3 (N13772, N13751, N5430, N10977);
nor NOR4 (N13773, N13725, N11370, N966, N2909);
nand NAND3 (N13774, N13770, N5389, N5211);
and AND4 (N13775, N13774, N12273, N10529, N6207);
buf BUF1 (N13776, N13771);
buf BUF1 (N13777, N13758);
buf BUF1 (N13778, N13767);
nand NAND4 (N13779, N13776, N11416, N3737, N5646);
nand NAND4 (N13780, N13777, N7251, N13050, N5297);
or OR2 (N13781, N13780, N12876);
nor NOR2 (N13782, N13766, N1811);
nor NOR3 (N13783, N13775, N8969, N1844);
xor XOR2 (N13784, N13772, N5971);
buf BUF1 (N13785, N13773);
or OR2 (N13786, N13724, N5652);
buf BUF1 (N13787, N13781);
nor NOR2 (N13788, N13782, N4516);
buf BUF1 (N13789, N13783);
and AND3 (N13790, N13778, N2088, N6165);
nand NAND2 (N13791, N13790, N791);
not NOT1 (N13792, N13784);
and AND2 (N13793, N13788, N5266);
nand NAND2 (N13794, N13768, N4500);
nand NAND2 (N13795, N13793, N6520);
nand NAND3 (N13796, N13787, N13249, N6049);
and AND2 (N13797, N13795, N9926);
xor XOR2 (N13798, N13785, N556);
or OR2 (N13799, N13769, N12904);
xor XOR2 (N13800, N13791, N4985);
or OR4 (N13801, N13797, N11241, N10786, N8907);
buf BUF1 (N13802, N13801);
buf BUF1 (N13803, N13798);
or OR3 (N13804, N13779, N13664, N1565);
nand NAND3 (N13805, N13789, N6837, N3831);
nand NAND4 (N13806, N13792, N10749, N5348, N739);
nand NAND4 (N13807, N13796, N1220, N8718, N13539);
nor NOR2 (N13808, N13806, N1881);
not NOT1 (N13809, N13807);
and AND4 (N13810, N13786, N9787, N3722, N7133);
and AND2 (N13811, N13810, N10049);
not NOT1 (N13812, N13800);
xor XOR2 (N13813, N13799, N624);
buf BUF1 (N13814, N13811);
xor XOR2 (N13815, N13814, N7);
xor XOR2 (N13816, N13812, N155);
or OR2 (N13817, N13808, N3688);
xor XOR2 (N13818, N13805, N7359);
buf BUF1 (N13819, N13816);
not NOT1 (N13820, N13818);
or OR2 (N13821, N13802, N12009);
nand NAND4 (N13822, N13817, N9086, N10776, N6222);
or OR3 (N13823, N13809, N4048, N4798);
or OR2 (N13824, N13823, N12669);
buf BUF1 (N13825, N13804);
or OR4 (N13826, N13825, N7572, N7225, N6240);
and AND2 (N13827, N13822, N10013);
xor XOR2 (N13828, N13821, N2681);
xor XOR2 (N13829, N13794, N7458);
and AND2 (N13830, N13819, N11029);
nand NAND4 (N13831, N13828, N6640, N204, N11038);
buf BUF1 (N13832, N13827);
not NOT1 (N13833, N13815);
not NOT1 (N13834, N13830);
nand NAND4 (N13835, N13826, N6123, N11292, N13303);
or OR2 (N13836, N13820, N9017);
or OR4 (N13837, N13803, N1604, N4852, N2823);
xor XOR2 (N13838, N13824, N12123);
or OR3 (N13839, N13829, N12591, N11842);
buf BUF1 (N13840, N13813);
not NOT1 (N13841, N13835);
or OR2 (N13842, N13833, N10190);
xor XOR2 (N13843, N13841, N1336);
and AND3 (N13844, N13839, N12162, N2743);
nor NOR3 (N13845, N13840, N596, N5811);
and AND2 (N13846, N13837, N12257);
nand NAND2 (N13847, N13834, N5957);
nor NOR2 (N13848, N13846, N4959);
not NOT1 (N13849, N13847);
nor NOR2 (N13850, N13832, N9645);
and AND3 (N13851, N13845, N3285, N9404);
nor NOR3 (N13852, N13844, N9889, N9914);
not NOT1 (N13853, N13851);
or OR4 (N13854, N13852, N6193, N7453, N3353);
buf BUF1 (N13855, N13831);
nor NOR4 (N13856, N13854, N1513, N6067, N12953);
nor NOR3 (N13857, N13855, N10212, N13027);
buf BUF1 (N13858, N13838);
and AND2 (N13859, N13848, N6641);
xor XOR2 (N13860, N13850, N11625);
or OR3 (N13861, N13860, N9594, N10531);
nor NOR2 (N13862, N13853, N2409);
not NOT1 (N13863, N13842);
nand NAND3 (N13864, N13856, N9044, N12981);
not NOT1 (N13865, N13843);
nor NOR2 (N13866, N13865, N5747);
and AND4 (N13867, N13862, N3706, N1531, N4330);
or OR3 (N13868, N13859, N10060, N1761);
nand NAND2 (N13869, N13866, N12921);
nand NAND2 (N13870, N13858, N5161);
xor XOR2 (N13871, N13861, N1449);
nor NOR2 (N13872, N13870, N12941);
buf BUF1 (N13873, N13849);
not NOT1 (N13874, N13868);
and AND2 (N13875, N13867, N9601);
nor NOR3 (N13876, N13872, N351, N9159);
or OR3 (N13877, N13873, N4762, N650);
buf BUF1 (N13878, N13877);
not NOT1 (N13879, N13836);
nand NAND2 (N13880, N13857, N3838);
nand NAND2 (N13881, N13879, N301);
and AND3 (N13882, N13864, N1593, N3115);
or OR4 (N13883, N13878, N9946, N10859, N11224);
or OR2 (N13884, N13881, N488);
and AND2 (N13885, N13880, N6587);
and AND4 (N13886, N13869, N11991, N1207, N7921);
not NOT1 (N13887, N13886);
nand NAND2 (N13888, N13883, N11959);
buf BUF1 (N13889, N13888);
and AND3 (N13890, N13889, N11469, N664);
and AND4 (N13891, N13884, N6216, N7097, N975);
nor NOR4 (N13892, N13863, N9008, N11739, N3390);
or OR4 (N13893, N13887, N7191, N3339, N6059);
xor XOR2 (N13894, N13890, N10924);
buf BUF1 (N13895, N13874);
and AND3 (N13896, N13882, N8772, N3063);
xor XOR2 (N13897, N13885, N2878);
nand NAND2 (N13898, N13894, N12418);
buf BUF1 (N13899, N13896);
and AND2 (N13900, N13871, N11495);
xor XOR2 (N13901, N13899, N6184);
buf BUF1 (N13902, N13876);
not NOT1 (N13903, N13900);
nand NAND3 (N13904, N13893, N2498, N7127);
nand NAND4 (N13905, N13892, N2543, N10455, N7518);
nand NAND4 (N13906, N13898, N9736, N8061, N11322);
nand NAND2 (N13907, N13897, N328);
or OR2 (N13908, N13895, N2061);
and AND3 (N13909, N13907, N2548, N6116);
xor XOR2 (N13910, N13901, N10315);
and AND3 (N13911, N13904, N765, N3985);
or OR4 (N13912, N13905, N2893, N11460, N6169);
nand NAND4 (N13913, N13875, N13624, N7969, N12261);
nand NAND3 (N13914, N13913, N3161, N6340);
buf BUF1 (N13915, N13911);
buf BUF1 (N13916, N13906);
and AND4 (N13917, N13915, N11793, N3835, N3206);
xor XOR2 (N13918, N13910, N13770);
nand NAND2 (N13919, N13908, N21);
buf BUF1 (N13920, N13891);
buf BUF1 (N13921, N13914);
or OR4 (N13922, N13917, N7102, N1824, N12488);
or OR3 (N13923, N13921, N9451, N7896);
not NOT1 (N13924, N13902);
and AND2 (N13925, N13923, N2272);
or OR2 (N13926, N13916, N10803);
and AND2 (N13927, N13918, N13476);
not NOT1 (N13928, N13924);
nand NAND4 (N13929, N13903, N7217, N2633, N4752);
nor NOR3 (N13930, N13929, N9404, N8099);
and AND2 (N13931, N13920, N3390);
nor NOR2 (N13932, N13928, N490);
nand NAND2 (N13933, N13930, N762);
nand NAND3 (N13934, N13932, N4487, N11673);
or OR2 (N13935, N13927, N4542);
xor XOR2 (N13936, N13931, N7690);
buf BUF1 (N13937, N13925);
buf BUF1 (N13938, N13935);
not NOT1 (N13939, N13909);
and AND3 (N13940, N13939, N5197, N1597);
not NOT1 (N13941, N13933);
not NOT1 (N13942, N13941);
or OR3 (N13943, N13919, N4383, N2348);
and AND2 (N13944, N13943, N7895);
or OR4 (N13945, N13940, N1024, N3727, N12647);
nand NAND3 (N13946, N13942, N11582, N4318);
nand NAND3 (N13947, N13912, N3294, N13557);
nand NAND3 (N13948, N13934, N7539, N6071);
nand NAND2 (N13949, N13948, N6332);
xor XOR2 (N13950, N13945, N13684);
nor NOR4 (N13951, N13950, N11813, N7849, N6905);
xor XOR2 (N13952, N13949, N4634);
and AND2 (N13953, N13938, N11427);
not NOT1 (N13954, N13952);
not NOT1 (N13955, N13951);
nor NOR4 (N13956, N13926, N11745, N2615, N10580);
and AND2 (N13957, N13936, N8415);
xor XOR2 (N13958, N13953, N5732);
not NOT1 (N13959, N13922);
nor NOR3 (N13960, N13954, N13102, N8546);
nor NOR4 (N13961, N13956, N4749, N7402, N2119);
nand NAND2 (N13962, N13946, N6916);
or OR3 (N13963, N13947, N1332, N6963);
or OR2 (N13964, N13963, N2160);
or OR2 (N13965, N13964, N12146);
or OR2 (N13966, N13961, N7594);
not NOT1 (N13967, N13960);
and AND4 (N13968, N13962, N12145, N12876, N4957);
buf BUF1 (N13969, N13955);
nor NOR4 (N13970, N13969, N3661, N6276, N856);
nand NAND2 (N13971, N13957, N9323);
nor NOR2 (N13972, N13968, N8861);
buf BUF1 (N13973, N13966);
nor NOR4 (N13974, N13937, N9516, N10175, N8829);
nand NAND2 (N13975, N13972, N8789);
not NOT1 (N13976, N13965);
and AND3 (N13977, N13970, N8229, N4747);
and AND4 (N13978, N13975, N12056, N9651, N13060);
buf BUF1 (N13979, N13976);
xor XOR2 (N13980, N13944, N5019);
or OR4 (N13981, N13967, N9377, N7802, N1143);
nand NAND2 (N13982, N13974, N3677);
and AND3 (N13983, N13973, N5816, N10048);
nor NOR4 (N13984, N13980, N288, N6250, N357);
buf BUF1 (N13985, N13978);
and AND4 (N13986, N13982, N12393, N861, N10758);
xor XOR2 (N13987, N13981, N1843);
buf BUF1 (N13988, N13959);
or OR2 (N13989, N13979, N8760);
xor XOR2 (N13990, N13983, N2860);
and AND4 (N13991, N13958, N10346, N10313, N13183);
not NOT1 (N13992, N13971);
nand NAND3 (N13993, N13990, N961, N9122);
xor XOR2 (N13994, N13985, N6529);
nand NAND2 (N13995, N13988, N7281);
or OR2 (N13996, N13994, N3296);
not NOT1 (N13997, N13977);
nand NAND3 (N13998, N13989, N12020, N8924);
or OR4 (N13999, N13984, N6226, N5542, N3723);
buf BUF1 (N14000, N13987);
or OR3 (N14001, N13999, N3031, N13326);
nand NAND4 (N14002, N13986, N5899, N8011, N13261);
nor NOR3 (N14003, N14002, N6767, N423);
xor XOR2 (N14004, N14000, N3422);
or OR3 (N14005, N13996, N13063, N1335);
not NOT1 (N14006, N13991);
nor NOR4 (N14007, N14003, N11046, N2301, N12011);
or OR4 (N14008, N14001, N2034, N11965, N4278);
or OR3 (N14009, N13995, N762, N12618);
or OR2 (N14010, N13993, N7949);
and AND3 (N14011, N13997, N13398, N2093);
nand NAND4 (N14012, N14008, N11701, N108, N13285);
nand NAND4 (N14013, N14010, N10938, N3938, N2617);
nand NAND2 (N14014, N14006, N12999);
not NOT1 (N14015, N14007);
and AND4 (N14016, N13998, N13309, N12062, N13006);
buf BUF1 (N14017, N14009);
nor NOR2 (N14018, N14004, N1716);
nand NAND2 (N14019, N14018, N9172);
and AND4 (N14020, N14015, N13873, N8032, N11717);
nand NAND3 (N14021, N14020, N9965, N10785);
or OR4 (N14022, N14016, N7083, N5391, N8352);
not NOT1 (N14023, N14021);
nor NOR3 (N14024, N14017, N744, N304);
xor XOR2 (N14025, N14011, N12388);
nand NAND4 (N14026, N13992, N2973, N8635, N11740);
xor XOR2 (N14027, N14012, N2777);
and AND2 (N14028, N14019, N12904);
buf BUF1 (N14029, N14013);
or OR2 (N14030, N14026, N11260);
and AND3 (N14031, N14005, N6343, N10034);
nand NAND2 (N14032, N14029, N12956);
not NOT1 (N14033, N14014);
nor NOR2 (N14034, N14022, N8776);
and AND3 (N14035, N14030, N13009, N5708);
xor XOR2 (N14036, N14025, N319);
nor NOR4 (N14037, N14035, N211, N4599, N8227);
or OR3 (N14038, N14031, N6518, N10763);
nor NOR2 (N14039, N14034, N12357);
buf BUF1 (N14040, N14027);
xor XOR2 (N14041, N14023, N13717);
nor NOR2 (N14042, N14039, N12968);
nand NAND3 (N14043, N14037, N1197, N4487);
xor XOR2 (N14044, N14024, N12807);
nand NAND3 (N14045, N14041, N8908, N2039);
xor XOR2 (N14046, N14032, N6988);
or OR4 (N14047, N14040, N4212, N12609, N2644);
xor XOR2 (N14048, N14042, N155);
not NOT1 (N14049, N14048);
nor NOR4 (N14050, N14043, N486, N11330, N5694);
buf BUF1 (N14051, N14047);
not NOT1 (N14052, N14051);
not NOT1 (N14053, N14033);
nand NAND2 (N14054, N14028, N7953);
and AND4 (N14055, N14038, N4734, N13478, N13370);
nand NAND4 (N14056, N14045, N13756, N2079, N11169);
not NOT1 (N14057, N14050);
nor NOR2 (N14058, N14057, N6163);
and AND4 (N14059, N14049, N8435, N6513, N13668);
nand NAND2 (N14060, N14055, N9913);
buf BUF1 (N14061, N14059);
nand NAND4 (N14062, N14058, N14024, N5409, N722);
not NOT1 (N14063, N14036);
nor NOR3 (N14064, N14052, N13740, N12357);
nand NAND3 (N14065, N14064, N5421, N1982);
and AND4 (N14066, N14060, N11329, N308, N886);
not NOT1 (N14067, N14056);
xor XOR2 (N14068, N14044, N9827);
nor NOR2 (N14069, N14065, N4622);
and AND2 (N14070, N14053, N12176);
and AND3 (N14071, N14070, N11082, N9176);
buf BUF1 (N14072, N14061);
buf BUF1 (N14073, N14067);
or OR2 (N14074, N14062, N9319);
or OR2 (N14075, N14074, N10162);
and AND4 (N14076, N14054, N12057, N6406, N4229);
or OR4 (N14077, N14066, N12098, N12038, N11509);
or OR2 (N14078, N14046, N4004);
and AND2 (N14079, N14078, N9688);
and AND4 (N14080, N14071, N7247, N511, N4419);
or OR4 (N14081, N14077, N6743, N5473, N5531);
buf BUF1 (N14082, N14069);
or OR2 (N14083, N14079, N13675);
nor NOR3 (N14084, N14081, N13681, N3546);
nand NAND4 (N14085, N14083, N9012, N5874, N3288);
not NOT1 (N14086, N14085);
not NOT1 (N14087, N14068);
nor NOR2 (N14088, N14087, N1838);
buf BUF1 (N14089, N14076);
or OR3 (N14090, N14072, N7125, N2727);
nand NAND2 (N14091, N14063, N12197);
and AND4 (N14092, N14082, N5006, N5256, N2729);
or OR3 (N14093, N14086, N11342, N10759);
nand NAND2 (N14094, N14073, N7234);
and AND2 (N14095, N14075, N5688);
and AND2 (N14096, N14093, N5384);
not NOT1 (N14097, N14089);
or OR4 (N14098, N14091, N4111, N837, N13224);
or OR4 (N14099, N14094, N7910, N1705, N6135);
nor NOR4 (N14100, N14099, N3389, N3157, N4455);
nand NAND4 (N14101, N14097, N13832, N4333, N13450);
buf BUF1 (N14102, N14084);
not NOT1 (N14103, N14096);
buf BUF1 (N14104, N14080);
nor NOR3 (N14105, N14092, N2716, N4120);
not NOT1 (N14106, N14101);
or OR3 (N14107, N14103, N7431, N11728);
nor NOR4 (N14108, N14088, N10420, N7766, N2199);
xor XOR2 (N14109, N14105, N3789);
nand NAND2 (N14110, N14095, N12318);
and AND3 (N14111, N14102, N12572, N11832);
not NOT1 (N14112, N14106);
buf BUF1 (N14113, N14109);
xor XOR2 (N14114, N14090, N8773);
nor NOR2 (N14115, N14110, N8410);
xor XOR2 (N14116, N14115, N6344);
buf BUF1 (N14117, N14104);
xor XOR2 (N14118, N14113, N3929);
nand NAND2 (N14119, N14114, N8505);
and AND4 (N14120, N14116, N12906, N5561, N781);
nand NAND3 (N14121, N14120, N6672, N7502);
buf BUF1 (N14122, N14100);
nor NOR4 (N14123, N14117, N6826, N4679, N8720);
nor NOR3 (N14124, N14098, N8107, N8141);
xor XOR2 (N14125, N14122, N5716);
nor NOR3 (N14126, N14118, N2161, N3754);
nor NOR4 (N14127, N14125, N4480, N1605, N4988);
xor XOR2 (N14128, N14126, N13164);
or OR3 (N14129, N14108, N8913, N9670);
nor NOR3 (N14130, N14107, N10076, N2363);
buf BUF1 (N14131, N14119);
or OR3 (N14132, N14130, N2274, N11697);
not NOT1 (N14133, N14128);
and AND3 (N14134, N14111, N839, N6758);
not NOT1 (N14135, N14134);
buf BUF1 (N14136, N14135);
xor XOR2 (N14137, N14121, N2035);
nor NOR4 (N14138, N14124, N3634, N13669, N12150);
not NOT1 (N14139, N14127);
buf BUF1 (N14140, N14129);
buf BUF1 (N14141, N14139);
nand NAND3 (N14142, N14141, N5602, N8095);
nor NOR2 (N14143, N14123, N2962);
or OR3 (N14144, N14132, N9282, N10193);
not NOT1 (N14145, N14131);
buf BUF1 (N14146, N14138);
not NOT1 (N14147, N14142);
and AND2 (N14148, N14140, N3109);
buf BUF1 (N14149, N14133);
nor NOR4 (N14150, N14145, N4074, N1547, N2179);
not NOT1 (N14151, N14147);
xor XOR2 (N14152, N14150, N7261);
not NOT1 (N14153, N14144);
nor NOR3 (N14154, N14148, N11257, N6910);
nand NAND3 (N14155, N14149, N238, N182);
buf BUF1 (N14156, N14146);
xor XOR2 (N14157, N14136, N12853);
nor NOR3 (N14158, N14112, N11801, N13141);
and AND3 (N14159, N14158, N7952, N13431);
and AND4 (N14160, N14154, N5674, N11295, N1703);
xor XOR2 (N14161, N14152, N13847);
nand NAND4 (N14162, N14155, N7171, N6216, N4939);
and AND3 (N14163, N14151, N3674, N9016);
not NOT1 (N14164, N14143);
not NOT1 (N14165, N14160);
or OR3 (N14166, N14153, N337, N3716);
nor NOR4 (N14167, N14156, N3463, N10171, N11106);
buf BUF1 (N14168, N14164);
buf BUF1 (N14169, N14157);
nand NAND4 (N14170, N14165, N2687, N4687, N6882);
buf BUF1 (N14171, N14137);
nor NOR2 (N14172, N14162, N10689);
or OR2 (N14173, N14171, N10118);
nor NOR3 (N14174, N14169, N2972, N8166);
not NOT1 (N14175, N14167);
xor XOR2 (N14176, N14161, N6089);
not NOT1 (N14177, N14175);
not NOT1 (N14178, N14176);
nor NOR3 (N14179, N14170, N2157, N11832);
xor XOR2 (N14180, N14173, N3665);
nand NAND2 (N14181, N14172, N7489);
nand NAND2 (N14182, N14168, N13188);
nand NAND3 (N14183, N14180, N12426, N11481);
not NOT1 (N14184, N14163);
and AND2 (N14185, N14179, N10868);
nor NOR2 (N14186, N14159, N6091);
buf BUF1 (N14187, N14178);
or OR3 (N14188, N14166, N9201, N7426);
nand NAND3 (N14189, N14184, N6017, N6006);
buf BUF1 (N14190, N14181);
nand NAND2 (N14191, N14174, N13511);
buf BUF1 (N14192, N14188);
or OR3 (N14193, N14191, N10872, N10180);
nand NAND4 (N14194, N14193, N6556, N11831, N13806);
or OR3 (N14195, N14182, N11667, N13370);
nand NAND4 (N14196, N14195, N14012, N11139, N5464);
and AND2 (N14197, N14192, N405);
buf BUF1 (N14198, N14196);
xor XOR2 (N14199, N14183, N10095);
or OR4 (N14200, N14177, N199, N8445, N4073);
nand NAND2 (N14201, N14200, N14038);
nor NOR2 (N14202, N14198, N8012);
buf BUF1 (N14203, N14185);
buf BUF1 (N14204, N14190);
or OR3 (N14205, N14203, N9519, N13346);
nor NOR4 (N14206, N14199, N4113, N6144, N3528);
or OR2 (N14207, N14194, N11131);
xor XOR2 (N14208, N14189, N10874);
nor NOR2 (N14209, N14201, N10);
not NOT1 (N14210, N14208);
nand NAND3 (N14211, N14186, N8424, N1638);
and AND2 (N14212, N14197, N2861);
and AND3 (N14213, N14187, N4906, N1446);
nand NAND3 (N14214, N14202, N8370, N6586);
and AND2 (N14215, N14205, N6809);
and AND2 (N14216, N14214, N11057);
buf BUF1 (N14217, N14213);
buf BUF1 (N14218, N14207);
and AND2 (N14219, N14216, N7292);
and AND2 (N14220, N14218, N12574);
nor NOR2 (N14221, N14211, N2142);
xor XOR2 (N14222, N14219, N2326);
or OR4 (N14223, N14221, N5315, N12906, N8154);
not NOT1 (N14224, N14220);
buf BUF1 (N14225, N14223);
not NOT1 (N14226, N14209);
or OR4 (N14227, N14226, N12637, N12215, N8206);
nand NAND3 (N14228, N14217, N1462, N12984);
nor NOR4 (N14229, N14222, N5791, N72, N448);
not NOT1 (N14230, N14206);
nand NAND2 (N14231, N14230, N7775);
not NOT1 (N14232, N14224);
buf BUF1 (N14233, N14225);
not NOT1 (N14234, N14227);
not NOT1 (N14235, N14229);
buf BUF1 (N14236, N14235);
nand NAND3 (N14237, N14234, N9232, N11357);
buf BUF1 (N14238, N14212);
xor XOR2 (N14239, N14215, N12764);
nor NOR3 (N14240, N14236, N4386, N5856);
or OR4 (N14241, N14237, N389, N5376, N2624);
not NOT1 (N14242, N14233);
or OR4 (N14243, N14238, N7422, N10408, N13551);
buf BUF1 (N14244, N14210);
not NOT1 (N14245, N14232);
and AND2 (N14246, N14204, N3248);
nor NOR4 (N14247, N14239, N10957, N7203, N10338);
xor XOR2 (N14248, N14245, N2400);
or OR3 (N14249, N14244, N3478, N10232);
or OR4 (N14250, N14242, N1144, N3610, N9982);
buf BUF1 (N14251, N14241);
or OR2 (N14252, N14249, N1187);
or OR3 (N14253, N14250, N8457, N706);
not NOT1 (N14254, N14248);
or OR3 (N14255, N14251, N14167, N4074);
nand NAND2 (N14256, N14243, N7022);
nand NAND3 (N14257, N14256, N6949, N14243);
buf BUF1 (N14258, N14252);
xor XOR2 (N14259, N14254, N10547);
and AND2 (N14260, N14258, N8904);
buf BUF1 (N14261, N14247);
and AND2 (N14262, N14255, N13429);
nand NAND2 (N14263, N14231, N11623);
nor NOR4 (N14264, N14253, N59, N1626, N11453);
buf BUF1 (N14265, N14261);
buf BUF1 (N14266, N14240);
buf BUF1 (N14267, N14246);
not NOT1 (N14268, N14264);
xor XOR2 (N14269, N14260, N14161);
nor NOR3 (N14270, N14269, N7331, N14160);
nor NOR2 (N14271, N14262, N9386);
or OR3 (N14272, N14268, N1364, N7733);
buf BUF1 (N14273, N14270);
buf BUF1 (N14274, N14271);
and AND2 (N14275, N14257, N13453);
buf BUF1 (N14276, N14273);
nor NOR4 (N14277, N14228, N7056, N3016, N6494);
buf BUF1 (N14278, N14259);
buf BUF1 (N14279, N14275);
buf BUF1 (N14280, N14266);
and AND4 (N14281, N14276, N8386, N4649, N7085);
or OR2 (N14282, N14274, N8980);
or OR2 (N14283, N14278, N9298);
buf BUF1 (N14284, N14272);
buf BUF1 (N14285, N14283);
not NOT1 (N14286, N14280);
not NOT1 (N14287, N14263);
xor XOR2 (N14288, N14281, N7728);
nand NAND2 (N14289, N14267, N2509);
or OR3 (N14290, N14287, N5262, N7986);
xor XOR2 (N14291, N14289, N1599);
nor NOR2 (N14292, N14284, N3836);
or OR4 (N14293, N14277, N13760, N4815, N10431);
nand NAND4 (N14294, N14292, N11135, N5948, N5938);
or OR2 (N14295, N14282, N12618);
and AND4 (N14296, N14288, N3755, N6636, N13580);
or OR4 (N14297, N14294, N3441, N13500, N2348);
and AND2 (N14298, N14291, N13434);
not NOT1 (N14299, N14279);
or OR3 (N14300, N14285, N10712, N12996);
xor XOR2 (N14301, N14286, N6911);
xor XOR2 (N14302, N14265, N2468);
or OR4 (N14303, N14300, N9486, N14169, N10987);
not NOT1 (N14304, N14303);
buf BUF1 (N14305, N14298);
nor NOR4 (N14306, N14304, N5147, N11219, N13754);
and AND3 (N14307, N14301, N4219, N13329);
and AND2 (N14308, N14305, N4701);
nor NOR4 (N14309, N14296, N11638, N12685, N4153);
xor XOR2 (N14310, N14306, N4567);
xor XOR2 (N14311, N14295, N9002);
not NOT1 (N14312, N14302);
nor NOR2 (N14313, N14290, N14174);
xor XOR2 (N14314, N14308, N732);
nand NAND3 (N14315, N14299, N13902, N12610);
and AND3 (N14316, N14315, N10451, N6363);
buf BUF1 (N14317, N14313);
not NOT1 (N14318, N14314);
nor NOR3 (N14319, N14311, N7312, N11254);
nor NOR3 (N14320, N14316, N5884, N4149);
xor XOR2 (N14321, N14307, N6725);
and AND3 (N14322, N14321, N4219, N7454);
or OR3 (N14323, N14319, N10359, N3488);
or OR3 (N14324, N14293, N9510, N8713);
not NOT1 (N14325, N14317);
not NOT1 (N14326, N14322);
xor XOR2 (N14327, N14297, N12837);
not NOT1 (N14328, N14310);
buf BUF1 (N14329, N14327);
xor XOR2 (N14330, N14309, N11721);
not NOT1 (N14331, N14330);
xor XOR2 (N14332, N14325, N7537);
and AND4 (N14333, N14332, N11813, N6507, N2333);
nor NOR2 (N14334, N14312, N9794);
and AND4 (N14335, N14320, N4458, N2148, N1509);
buf BUF1 (N14336, N14331);
xor XOR2 (N14337, N14318, N12693);
not NOT1 (N14338, N14329);
or OR4 (N14339, N14337, N6240, N639, N13496);
xor XOR2 (N14340, N14323, N893);
or OR3 (N14341, N14333, N4292, N1579);
buf BUF1 (N14342, N14328);
not NOT1 (N14343, N14342);
nor NOR4 (N14344, N14334, N8367, N3371, N11669);
not NOT1 (N14345, N14343);
xor XOR2 (N14346, N14341, N13768);
or OR3 (N14347, N14339, N13825, N1194);
buf BUF1 (N14348, N14347);
not NOT1 (N14349, N14344);
not NOT1 (N14350, N14324);
and AND4 (N14351, N14346, N6452, N2236, N6094);
buf BUF1 (N14352, N14335);
nand NAND2 (N14353, N14348, N1743);
nand NAND3 (N14354, N14338, N10397, N4373);
buf BUF1 (N14355, N14349);
xor XOR2 (N14356, N14354, N1982);
not NOT1 (N14357, N14356);
not NOT1 (N14358, N14355);
nand NAND3 (N14359, N14358, N14099, N9360);
xor XOR2 (N14360, N14336, N4767);
buf BUF1 (N14361, N14340);
nand NAND4 (N14362, N14353, N7291, N6736, N8312);
xor XOR2 (N14363, N14362, N5884);
nor NOR2 (N14364, N14351, N13844);
or OR2 (N14365, N14357, N13714);
and AND2 (N14366, N14352, N608);
nand NAND3 (N14367, N14366, N3731, N11961);
and AND2 (N14368, N14350, N13145);
nand NAND4 (N14369, N14345, N7759, N4521, N5364);
not NOT1 (N14370, N14365);
nor NOR2 (N14371, N14361, N7351);
not NOT1 (N14372, N14363);
xor XOR2 (N14373, N14369, N9277);
and AND2 (N14374, N14359, N11729);
xor XOR2 (N14375, N14326, N10166);
buf BUF1 (N14376, N14370);
nor NOR3 (N14377, N14373, N11542, N1350);
buf BUF1 (N14378, N14368);
and AND3 (N14379, N14377, N7119, N14192);
xor XOR2 (N14380, N14374, N148);
not NOT1 (N14381, N14360);
and AND2 (N14382, N14379, N7327);
nor NOR2 (N14383, N14371, N1100);
or OR4 (N14384, N14364, N13005, N12939, N4457);
buf BUF1 (N14385, N14384);
nor NOR4 (N14386, N14367, N9474, N7017, N1536);
buf BUF1 (N14387, N14376);
buf BUF1 (N14388, N14385);
not NOT1 (N14389, N14375);
not NOT1 (N14390, N14389);
and AND2 (N14391, N14381, N8664);
and AND2 (N14392, N14386, N11232);
xor XOR2 (N14393, N14382, N11893);
or OR3 (N14394, N14393, N10384, N6373);
buf BUF1 (N14395, N14394);
buf BUF1 (N14396, N14388);
and AND3 (N14397, N14396, N1335, N4638);
and AND3 (N14398, N14395, N6566, N1497);
or OR3 (N14399, N14398, N30, N9725);
nor NOR2 (N14400, N14390, N2025);
buf BUF1 (N14401, N14372);
or OR4 (N14402, N14401, N11561, N10366, N2011);
nor NOR3 (N14403, N14383, N13131, N8904);
buf BUF1 (N14404, N14378);
nand NAND3 (N14405, N14387, N7984, N13523);
and AND4 (N14406, N14399, N4950, N3425, N8811);
or OR4 (N14407, N14403, N4303, N3864, N6807);
and AND4 (N14408, N14380, N4857, N2612, N1922);
or OR4 (N14409, N14406, N12752, N10458, N9865);
and AND2 (N14410, N14397, N11360);
nor NOR4 (N14411, N14408, N7595, N6920, N875);
or OR3 (N14412, N14405, N1956, N1901);
nand NAND4 (N14413, N14402, N3885, N11383, N1053);
or OR3 (N14414, N14391, N8861, N10956);
xor XOR2 (N14415, N14412, N7570);
nor NOR4 (N14416, N14409, N9606, N13357, N11755);
buf BUF1 (N14417, N14400);
nand NAND3 (N14418, N14410, N12039, N2859);
not NOT1 (N14419, N14418);
or OR4 (N14420, N14404, N2784, N7823, N2160);
nand NAND4 (N14421, N14420, N2860, N8508, N4094);
xor XOR2 (N14422, N14411, N3690);
not NOT1 (N14423, N14407);
xor XOR2 (N14424, N14416, N7718);
buf BUF1 (N14425, N14392);
buf BUF1 (N14426, N14424);
nor NOR3 (N14427, N14425, N2011, N11872);
or OR4 (N14428, N14417, N6104, N8023, N12259);
nor NOR3 (N14429, N14419, N4868, N11120);
and AND3 (N14430, N14423, N7079, N3060);
or OR3 (N14431, N14421, N11591, N13681);
not NOT1 (N14432, N14429);
xor XOR2 (N14433, N14428, N8120);
buf BUF1 (N14434, N14431);
and AND3 (N14435, N14414, N5196, N12627);
or OR3 (N14436, N14430, N2852, N12221);
xor XOR2 (N14437, N14426, N13026);
nor NOR2 (N14438, N14434, N3302);
nor NOR3 (N14439, N14422, N3561, N11759);
xor XOR2 (N14440, N14415, N12723);
xor XOR2 (N14441, N14435, N11992);
not NOT1 (N14442, N14441);
nand NAND2 (N14443, N14433, N5425);
nor NOR4 (N14444, N14413, N9361, N6563, N7883);
nor NOR2 (N14445, N14436, N250);
xor XOR2 (N14446, N14438, N3879);
or OR3 (N14447, N14437, N690, N6438);
and AND2 (N14448, N14445, N6697);
and AND2 (N14449, N14439, N13175);
nand NAND4 (N14450, N14448, N477, N8922, N5518);
buf BUF1 (N14451, N14449);
buf BUF1 (N14452, N14447);
and AND2 (N14453, N14452, N2335);
nor NOR2 (N14454, N14432, N5681);
xor XOR2 (N14455, N14444, N3681);
or OR2 (N14456, N14440, N13715);
or OR3 (N14457, N14446, N470, N13993);
nand NAND3 (N14458, N14450, N4823, N3274);
nand NAND4 (N14459, N14443, N9149, N1832, N8860);
xor XOR2 (N14460, N14455, N2246);
nor NOR2 (N14461, N14454, N5999);
not NOT1 (N14462, N14442);
not NOT1 (N14463, N14451);
not NOT1 (N14464, N14463);
nand NAND3 (N14465, N14462, N172, N6861);
xor XOR2 (N14466, N14458, N4433);
not NOT1 (N14467, N14457);
not NOT1 (N14468, N14464);
nor NOR2 (N14469, N14456, N13912);
nand NAND3 (N14470, N14427, N8781, N4392);
or OR4 (N14471, N14459, N13342, N6640, N3663);
xor XOR2 (N14472, N14469, N10370);
xor XOR2 (N14473, N14461, N11606);
xor XOR2 (N14474, N14472, N839);
xor XOR2 (N14475, N14470, N1673);
xor XOR2 (N14476, N14466, N4668);
and AND3 (N14477, N14471, N9248, N3904);
not NOT1 (N14478, N14465);
and AND2 (N14479, N14475, N5468);
xor XOR2 (N14480, N14476, N374);
nand NAND2 (N14481, N14460, N13513);
nor NOR2 (N14482, N14481, N7910);
nor NOR3 (N14483, N14482, N8560, N6096);
nor NOR4 (N14484, N14453, N8553, N3850, N2179);
nand NAND3 (N14485, N14479, N4486, N7093);
or OR2 (N14486, N14468, N3341);
not NOT1 (N14487, N14483);
buf BUF1 (N14488, N14487);
not NOT1 (N14489, N14478);
nor NOR2 (N14490, N14477, N2358);
nand NAND4 (N14491, N14467, N5389, N14410, N6656);
and AND3 (N14492, N14491, N9424, N5136);
or OR4 (N14493, N14484, N14089, N8892, N9705);
buf BUF1 (N14494, N14485);
nor NOR4 (N14495, N14486, N10323, N561, N559);
not NOT1 (N14496, N14489);
buf BUF1 (N14497, N14490);
xor XOR2 (N14498, N14496, N14329);
and AND3 (N14499, N14480, N1191, N10514);
buf BUF1 (N14500, N14474);
nor NOR2 (N14501, N14493, N1892);
and AND4 (N14502, N14501, N3457, N9727, N1321);
nand NAND3 (N14503, N14500, N11618, N4734);
and AND4 (N14504, N14492, N2421, N14304, N7873);
xor XOR2 (N14505, N14504, N2113);
xor XOR2 (N14506, N14473, N14323);
nand NAND4 (N14507, N14505, N6412, N1128, N8414);
or OR4 (N14508, N14502, N9278, N2585, N7666);
not NOT1 (N14509, N14498);
nand NAND3 (N14510, N14499, N12706, N1690);
not NOT1 (N14511, N14506);
and AND3 (N14512, N14503, N7967, N13855);
or OR2 (N14513, N14494, N12466);
xor XOR2 (N14514, N14512, N5810);
nor NOR3 (N14515, N14513, N7097, N11465);
nor NOR2 (N14516, N14497, N12335);
and AND4 (N14517, N14516, N3354, N10905, N1306);
and AND3 (N14518, N14515, N7357, N8782);
xor XOR2 (N14519, N14510, N1267);
nor NOR4 (N14520, N14507, N14432, N821, N6024);
not NOT1 (N14521, N14488);
xor XOR2 (N14522, N14521, N9537);
and AND2 (N14523, N14520, N12497);
and AND4 (N14524, N14523, N13846, N3218, N14144);
and AND2 (N14525, N14495, N9643);
and AND2 (N14526, N14514, N1274);
not NOT1 (N14527, N14524);
nand NAND2 (N14528, N14509, N13784);
xor XOR2 (N14529, N14528, N1040);
buf BUF1 (N14530, N14519);
or OR2 (N14531, N14518, N280);
nand NAND3 (N14532, N14525, N5251, N3640);
and AND2 (N14533, N14527, N6753);
nor NOR4 (N14534, N14508, N9728, N4402, N12013);
nand NAND4 (N14535, N14526, N2672, N10762, N8801);
xor XOR2 (N14536, N14511, N7783);
xor XOR2 (N14537, N14530, N5816);
xor XOR2 (N14538, N14535, N2430);
nor NOR4 (N14539, N14517, N9620, N10809, N6533);
and AND3 (N14540, N14529, N12968, N9052);
or OR2 (N14541, N14522, N1197);
not NOT1 (N14542, N14536);
buf BUF1 (N14543, N14540);
nor NOR2 (N14544, N14532, N13657);
xor XOR2 (N14545, N14541, N4799);
nand NAND4 (N14546, N14538, N14162, N4898, N11109);
nand NAND3 (N14547, N14544, N6582, N2210);
and AND4 (N14548, N14537, N13795, N2529, N1958);
nand NAND4 (N14549, N14542, N11101, N3861, N10997);
nand NAND4 (N14550, N14548, N10821, N7961, N5530);
xor XOR2 (N14551, N14545, N8892);
or OR3 (N14552, N14533, N12087, N6912);
not NOT1 (N14553, N14531);
buf BUF1 (N14554, N14547);
and AND4 (N14555, N14543, N13118, N10691, N6667);
xor XOR2 (N14556, N14553, N7836);
not NOT1 (N14557, N14539);
nor NOR4 (N14558, N14552, N9010, N6029, N12454);
nor NOR4 (N14559, N14558, N8155, N7652, N11610);
nor NOR2 (N14560, N14534, N12006);
nor NOR4 (N14561, N14546, N8831, N4660, N14344);
or OR4 (N14562, N14561, N3499, N938, N2838);
xor XOR2 (N14563, N14555, N3176);
or OR2 (N14564, N14562, N5532);
and AND3 (N14565, N14549, N2304, N8055);
buf BUF1 (N14566, N14557);
xor XOR2 (N14567, N14554, N6005);
xor XOR2 (N14568, N14551, N11324);
or OR2 (N14569, N14568, N8877);
buf BUF1 (N14570, N14567);
buf BUF1 (N14571, N14563);
nand NAND2 (N14572, N14565, N4748);
nor NOR4 (N14573, N14569, N8919, N3371, N8658);
buf BUF1 (N14574, N14573);
buf BUF1 (N14575, N14564);
or OR2 (N14576, N14560, N12076);
not NOT1 (N14577, N14576);
and AND4 (N14578, N14570, N14154, N5161, N5586);
or OR3 (N14579, N14574, N13092, N4835);
xor XOR2 (N14580, N14566, N11553);
nand NAND4 (N14581, N14556, N267, N2453, N8330);
nand NAND4 (N14582, N14578, N4276, N5512, N6944);
nor NOR4 (N14583, N14571, N5718, N7707, N4529);
buf BUF1 (N14584, N14581);
and AND4 (N14585, N14584, N2370, N8210, N10829);
buf BUF1 (N14586, N14579);
or OR2 (N14587, N14559, N7870);
nor NOR4 (N14588, N14585, N2205, N11802, N12845);
xor XOR2 (N14589, N14572, N1371);
xor XOR2 (N14590, N14586, N970);
or OR4 (N14591, N14580, N10386, N7769, N3707);
and AND2 (N14592, N14583, N12595);
or OR2 (N14593, N14575, N10109);
and AND3 (N14594, N14550, N3527, N12578);
buf BUF1 (N14595, N14590);
or OR4 (N14596, N14591, N13733, N3374, N4671);
buf BUF1 (N14597, N14594);
or OR4 (N14598, N14589, N4916, N6068, N11231);
xor XOR2 (N14599, N14592, N1845);
and AND3 (N14600, N14587, N14073, N10365);
nor NOR4 (N14601, N14598, N11325, N7964, N3297);
nor NOR4 (N14602, N14599, N8620, N12048, N103);
or OR3 (N14603, N14577, N5544, N456);
not NOT1 (N14604, N14595);
xor XOR2 (N14605, N14603, N10062);
not NOT1 (N14606, N14604);
not NOT1 (N14607, N14593);
and AND3 (N14608, N14601, N2233, N6028);
buf BUF1 (N14609, N14596);
and AND3 (N14610, N14588, N853, N12020);
nor NOR3 (N14611, N14610, N8674, N1733);
nor NOR4 (N14612, N14600, N2439, N9186, N14606);
xor XOR2 (N14613, N6434, N3878);
nor NOR4 (N14614, N14612, N9178, N9354, N4429);
xor XOR2 (N14615, N14607, N11584);
not NOT1 (N14616, N14597);
xor XOR2 (N14617, N14616, N11845);
and AND2 (N14618, N14608, N10551);
or OR4 (N14619, N14582, N13630, N12202, N10461);
xor XOR2 (N14620, N14617, N2870);
and AND4 (N14621, N14620, N9044, N7815, N14605);
nand NAND4 (N14622, N11774, N6480, N3918, N8224);
and AND3 (N14623, N14621, N5821, N1352);
nor NOR2 (N14624, N14613, N8576);
and AND2 (N14625, N14614, N7682);
xor XOR2 (N14626, N14622, N11498);
or OR2 (N14627, N14625, N7496);
xor XOR2 (N14628, N14624, N102);
xor XOR2 (N14629, N14602, N14368);
or OR3 (N14630, N14626, N191, N6773);
buf BUF1 (N14631, N14619);
not NOT1 (N14632, N14609);
or OR4 (N14633, N14611, N9600, N4373, N9646);
buf BUF1 (N14634, N14627);
xor XOR2 (N14635, N14634, N6329);
nand NAND4 (N14636, N14618, N9142, N9981, N7000);
buf BUF1 (N14637, N14631);
buf BUF1 (N14638, N14628);
xor XOR2 (N14639, N14637, N2462);
and AND4 (N14640, N14633, N13889, N7922, N6506);
nand NAND2 (N14641, N14640, N3719);
nand NAND4 (N14642, N14635, N12185, N10358, N5720);
or OR2 (N14643, N14642, N2202);
or OR2 (N14644, N14641, N4330);
xor XOR2 (N14645, N14623, N1369);
nand NAND4 (N14646, N14643, N7975, N13828, N3663);
nand NAND2 (N14647, N14630, N8624);
and AND3 (N14648, N14647, N11557, N6878);
nor NOR4 (N14649, N14615, N1611, N11776, N983);
not NOT1 (N14650, N14644);
and AND3 (N14651, N14645, N5574, N10903);
and AND3 (N14652, N14646, N8298, N10096);
not NOT1 (N14653, N14651);
and AND4 (N14654, N14636, N13165, N2655, N10777);
or OR3 (N14655, N14650, N12017, N3549);
or OR4 (N14656, N14639, N11240, N5685, N3322);
buf BUF1 (N14657, N14656);
xor XOR2 (N14658, N14657, N9159);
nor NOR4 (N14659, N14648, N11859, N1018, N9534);
nand NAND4 (N14660, N14653, N4280, N7940, N9983);
nor NOR3 (N14661, N14658, N3663, N6729);
not NOT1 (N14662, N14649);
nor NOR3 (N14663, N14632, N13824, N10831);
xor XOR2 (N14664, N14654, N1882);
nand NAND3 (N14665, N14661, N5227, N407);
nand NAND2 (N14666, N14655, N11606);
or OR4 (N14667, N14660, N11126, N3847, N13014);
or OR4 (N14668, N14652, N6105, N2864, N12669);
nor NOR2 (N14669, N14664, N8236);
and AND4 (N14670, N14659, N466, N3289, N11500);
and AND2 (N14671, N14668, N13138);
or OR2 (N14672, N14669, N10331);
not NOT1 (N14673, N14670);
nand NAND4 (N14674, N14662, N3516, N12427, N2078);
xor XOR2 (N14675, N14667, N5395);
nand NAND3 (N14676, N14672, N5836, N12385);
buf BUF1 (N14677, N14666);
and AND3 (N14678, N14671, N7823, N1895);
buf BUF1 (N14679, N14665);
xor XOR2 (N14680, N14674, N11060);
nand NAND2 (N14681, N14678, N14365);
not NOT1 (N14682, N14673);
or OR2 (N14683, N14676, N6236);
and AND4 (N14684, N14675, N9764, N6443, N10718);
not NOT1 (N14685, N14682);
and AND2 (N14686, N14663, N14417);
or OR3 (N14687, N14680, N3717, N13071);
or OR2 (N14688, N14687, N14611);
xor XOR2 (N14689, N14688, N5746);
xor XOR2 (N14690, N14638, N5234);
not NOT1 (N14691, N14683);
or OR3 (N14692, N14689, N3409, N6114);
and AND4 (N14693, N14684, N5604, N6228, N9988);
and AND2 (N14694, N14691, N8829);
nor NOR2 (N14695, N14685, N3018);
or OR4 (N14696, N14690, N8174, N8241, N3866);
nand NAND4 (N14697, N14677, N12147, N4312, N6066);
nor NOR3 (N14698, N14681, N6199, N6000);
and AND2 (N14699, N14692, N2976);
buf BUF1 (N14700, N14679);
not NOT1 (N14701, N14695);
not NOT1 (N14702, N14686);
nand NAND2 (N14703, N14697, N8956);
nor NOR2 (N14704, N14693, N2570);
or OR4 (N14705, N14629, N7971, N5337, N10585);
not NOT1 (N14706, N14701);
xor XOR2 (N14707, N14696, N10623);
and AND2 (N14708, N14704, N5228);
nand NAND3 (N14709, N14694, N6486, N12541);
buf BUF1 (N14710, N14702);
xor XOR2 (N14711, N14707, N325);
xor XOR2 (N14712, N14698, N13841);
buf BUF1 (N14713, N14700);
nor NOR2 (N14714, N14711, N6409);
and AND4 (N14715, N14709, N649, N12843, N1779);
nand NAND3 (N14716, N14699, N2322, N12199);
xor XOR2 (N14717, N14706, N6847);
xor XOR2 (N14718, N14715, N8853);
xor XOR2 (N14719, N14705, N10216);
not NOT1 (N14720, N14708);
and AND3 (N14721, N14716, N8085, N12273);
nor NOR2 (N14722, N14710, N6700);
buf BUF1 (N14723, N14712);
buf BUF1 (N14724, N14714);
or OR4 (N14725, N14721, N7354, N2434, N1981);
buf BUF1 (N14726, N14725);
not NOT1 (N14727, N14723);
nor NOR2 (N14728, N14722, N2308);
not NOT1 (N14729, N14713);
nor NOR4 (N14730, N14719, N8503, N10247, N6017);
nor NOR4 (N14731, N14718, N2334, N5053, N686);
xor XOR2 (N14732, N14730, N11770);
nor NOR3 (N14733, N14717, N5697, N11633);
xor XOR2 (N14734, N14720, N4870);
nand NAND3 (N14735, N14734, N603, N10704);
buf BUF1 (N14736, N14728);
and AND4 (N14737, N14703, N5387, N6105, N11310);
nand NAND2 (N14738, N14737, N5626);
not NOT1 (N14739, N14726);
xor XOR2 (N14740, N14738, N8259);
nor NOR3 (N14741, N14733, N4853, N9749);
and AND3 (N14742, N14735, N4076, N1951);
nor NOR3 (N14743, N14724, N13388, N13027);
or OR3 (N14744, N14732, N13981, N1998);
nor NOR2 (N14745, N14744, N10492);
nand NAND3 (N14746, N14727, N981, N9856);
buf BUF1 (N14747, N14729);
not NOT1 (N14748, N14739);
buf BUF1 (N14749, N14741);
buf BUF1 (N14750, N14736);
not NOT1 (N14751, N14742);
nand NAND4 (N14752, N14747, N13127, N5239, N2427);
xor XOR2 (N14753, N14745, N5026);
nor NOR2 (N14754, N14743, N6800);
nor NOR3 (N14755, N14746, N4040, N868);
buf BUF1 (N14756, N14754);
xor XOR2 (N14757, N14740, N912);
nor NOR2 (N14758, N14748, N7914);
xor XOR2 (N14759, N14753, N14702);
nor NOR3 (N14760, N14757, N9725, N6813);
not NOT1 (N14761, N14750);
xor XOR2 (N14762, N14751, N13500);
and AND3 (N14763, N14756, N907, N6370);
xor XOR2 (N14764, N14759, N12842);
nand NAND2 (N14765, N14764, N5877);
and AND4 (N14766, N14760, N1343, N3813, N2893);
not NOT1 (N14767, N14731);
buf BUF1 (N14768, N14762);
not NOT1 (N14769, N14752);
or OR3 (N14770, N14767, N797, N9182);
and AND3 (N14771, N14755, N4135, N7303);
buf BUF1 (N14772, N14769);
not NOT1 (N14773, N14770);
buf BUF1 (N14774, N14761);
or OR4 (N14775, N14771, N14652, N788, N12146);
or OR2 (N14776, N14774, N184);
and AND3 (N14777, N14749, N10635, N8933);
nand NAND2 (N14778, N14772, N12486);
and AND2 (N14779, N14777, N12492);
nor NOR3 (N14780, N14779, N11111, N12971);
xor XOR2 (N14781, N14763, N9501);
nor NOR4 (N14782, N14768, N5300, N8398, N7773);
not NOT1 (N14783, N14781);
buf BUF1 (N14784, N14783);
or OR3 (N14785, N14758, N13278, N7713);
xor XOR2 (N14786, N14773, N9115);
xor XOR2 (N14787, N14782, N11657);
nand NAND4 (N14788, N14786, N10915, N4509, N7336);
or OR3 (N14789, N14788, N11211, N6540);
and AND3 (N14790, N14787, N6271, N13346);
nor NOR4 (N14791, N14790, N3741, N13902, N9589);
not NOT1 (N14792, N14775);
or OR4 (N14793, N14778, N679, N1226, N6928);
buf BUF1 (N14794, N14791);
not NOT1 (N14795, N14789);
not NOT1 (N14796, N14784);
buf BUF1 (N14797, N14796);
nor NOR3 (N14798, N14794, N12545, N10943);
nand NAND4 (N14799, N14797, N5761, N14274, N10708);
not NOT1 (N14800, N14798);
or OR3 (N14801, N14765, N3609, N8718);
nand NAND2 (N14802, N14795, N2297);
nor NOR2 (N14803, N14793, N8823);
buf BUF1 (N14804, N14801);
and AND2 (N14805, N14799, N4263);
nor NOR2 (N14806, N14802, N12458);
xor XOR2 (N14807, N14800, N915);
not NOT1 (N14808, N14792);
nor NOR3 (N14809, N14806, N3592, N4883);
nand NAND2 (N14810, N14809, N7315);
and AND2 (N14811, N14804, N3203);
buf BUF1 (N14812, N14766);
nand NAND4 (N14813, N14776, N5073, N3479, N1916);
and AND2 (N14814, N14810, N7500);
not NOT1 (N14815, N14785);
and AND3 (N14816, N14807, N14055, N13080);
or OR4 (N14817, N14814, N9945, N9468, N3259);
or OR2 (N14818, N14812, N298);
buf BUF1 (N14819, N14803);
buf BUF1 (N14820, N14818);
buf BUF1 (N14821, N14808);
and AND4 (N14822, N14811, N11168, N6508, N1843);
not NOT1 (N14823, N14822);
or OR4 (N14824, N14819, N9174, N9655, N7466);
or OR2 (N14825, N14780, N6054);
nor NOR3 (N14826, N14821, N11665, N11013);
nor NOR3 (N14827, N14825, N14264, N6253);
and AND4 (N14828, N14823, N13097, N6790, N10588);
not NOT1 (N14829, N14817);
buf BUF1 (N14830, N14805);
and AND3 (N14831, N14829, N11821, N2509);
or OR3 (N14832, N14827, N1929, N3935);
nor NOR3 (N14833, N14832, N3597, N1869);
nor NOR2 (N14834, N14826, N13316);
and AND2 (N14835, N14831, N13121);
nand NAND2 (N14836, N14828, N2630);
or OR4 (N14837, N14813, N5121, N4297, N3540);
or OR2 (N14838, N14820, N9241);
and AND2 (N14839, N14835, N13582);
nand NAND3 (N14840, N14836, N6394, N8647);
or OR4 (N14841, N14830, N9379, N8227, N4725);
or OR3 (N14842, N14837, N10998, N5131);
not NOT1 (N14843, N14842);
nor NOR4 (N14844, N14815, N13589, N11408, N277);
nor NOR2 (N14845, N14841, N3743);
or OR2 (N14846, N14834, N10200);
and AND4 (N14847, N14844, N769, N9974, N7823);
buf BUF1 (N14848, N14838);
not NOT1 (N14849, N14847);
and AND3 (N14850, N14839, N5951, N11545);
nand NAND3 (N14851, N14816, N7553, N13779);
nand NAND3 (N14852, N14849, N11174, N8990);
buf BUF1 (N14853, N14850);
buf BUF1 (N14854, N14852);
nand NAND3 (N14855, N14854, N9178, N4641);
xor XOR2 (N14856, N14855, N8809);
nor NOR2 (N14857, N14856, N5366);
nand NAND3 (N14858, N14824, N14421, N11418);
nand NAND2 (N14859, N14845, N14449);
buf BUF1 (N14860, N14848);
nand NAND2 (N14861, N14859, N13223);
xor XOR2 (N14862, N14857, N5095);
nor NOR2 (N14863, N14840, N3236);
nand NAND2 (N14864, N14860, N4299);
and AND2 (N14865, N14833, N11031);
nor NOR3 (N14866, N14862, N3898, N5206);
xor XOR2 (N14867, N14843, N7815);
buf BUF1 (N14868, N14861);
not NOT1 (N14869, N14866);
or OR2 (N14870, N14865, N7997);
xor XOR2 (N14871, N14867, N3840);
buf BUF1 (N14872, N14864);
nor NOR4 (N14873, N14868, N3150, N8254, N1120);
nand NAND3 (N14874, N14863, N36, N6295);
buf BUF1 (N14875, N14873);
or OR4 (N14876, N14875, N2031, N2455, N10953);
or OR3 (N14877, N14874, N14218, N3897);
nand NAND2 (N14878, N14853, N1526);
nor NOR4 (N14879, N14871, N9811, N12239, N10716);
nor NOR2 (N14880, N14879, N11841);
buf BUF1 (N14881, N14878);
nand NAND2 (N14882, N14869, N5313);
nor NOR2 (N14883, N14880, N1666);
xor XOR2 (N14884, N14877, N14731);
not NOT1 (N14885, N14876);
or OR3 (N14886, N14883, N6089, N3792);
buf BUF1 (N14887, N14846);
and AND4 (N14888, N14882, N2391, N7225, N2089);
nor NOR2 (N14889, N14887, N2962);
and AND4 (N14890, N14872, N12625, N3260, N9504);
nor NOR4 (N14891, N14884, N13901, N12408, N5797);
xor XOR2 (N14892, N14891, N4358);
not NOT1 (N14893, N14870);
nor NOR2 (N14894, N14892, N11611);
and AND2 (N14895, N14888, N14739);
nand NAND4 (N14896, N14889, N13928, N3093, N1485);
not NOT1 (N14897, N14893);
or OR2 (N14898, N14851, N6334);
xor XOR2 (N14899, N14897, N12686);
not NOT1 (N14900, N14894);
or OR4 (N14901, N14881, N11822, N5494, N3064);
and AND2 (N14902, N14886, N10266);
nor NOR2 (N14903, N14885, N4618);
nor NOR3 (N14904, N14890, N9864, N5472);
or OR2 (N14905, N14903, N7063);
xor XOR2 (N14906, N14904, N2712);
buf BUF1 (N14907, N14906);
and AND3 (N14908, N14898, N13389, N4273);
nand NAND4 (N14909, N14896, N3108, N14463, N9218);
nand NAND2 (N14910, N14900, N2245);
xor XOR2 (N14911, N14907, N5782);
buf BUF1 (N14912, N14909);
not NOT1 (N14913, N14908);
nor NOR2 (N14914, N14899, N5222);
not NOT1 (N14915, N14901);
and AND3 (N14916, N14911, N12009, N12047);
and AND2 (N14917, N14915, N8517);
nand NAND2 (N14918, N14905, N1529);
nand NAND4 (N14919, N14895, N2004, N13035, N8007);
xor XOR2 (N14920, N14917, N381);
and AND2 (N14921, N14910, N7842);
and AND3 (N14922, N14919, N11511, N3363);
and AND3 (N14923, N14920, N4380, N13874);
nand NAND3 (N14924, N14912, N5481, N4599);
buf BUF1 (N14925, N14921);
nor NOR4 (N14926, N14916, N13307, N2786, N12917);
xor XOR2 (N14927, N14926, N9557);
xor XOR2 (N14928, N14918, N5480);
nor NOR2 (N14929, N14913, N10129);
or OR3 (N14930, N14922, N11353, N4063);
nor NOR2 (N14931, N14914, N14635);
or OR2 (N14932, N14924, N5754);
buf BUF1 (N14933, N14930);
xor XOR2 (N14934, N14929, N8641);
and AND4 (N14935, N14923, N11928, N13610, N5101);
or OR4 (N14936, N14931, N9192, N5507, N6831);
nand NAND4 (N14937, N14902, N6224, N12142, N8184);
and AND4 (N14938, N14935, N8043, N4337, N4439);
xor XOR2 (N14939, N14933, N5972);
not NOT1 (N14940, N14932);
xor XOR2 (N14941, N14937, N11977);
not NOT1 (N14942, N14928);
xor XOR2 (N14943, N14927, N8132);
not NOT1 (N14944, N14940);
nor NOR3 (N14945, N14939, N5118, N11256);
nor NOR2 (N14946, N14945, N928);
buf BUF1 (N14947, N14938);
nand NAND2 (N14948, N14944, N13310);
xor XOR2 (N14949, N14941, N1879);
not NOT1 (N14950, N14858);
not NOT1 (N14951, N14950);
buf BUF1 (N14952, N14947);
nor NOR4 (N14953, N14936, N8054, N6436, N12893);
buf BUF1 (N14954, N14925);
nor NOR4 (N14955, N14946, N12931, N3662, N2350);
nor NOR2 (N14956, N14955, N6098);
nor NOR3 (N14957, N14948, N4685, N3937);
or OR2 (N14958, N14954, N6008);
xor XOR2 (N14959, N14934, N13143);
or OR4 (N14960, N14952, N14476, N10403, N6582);
or OR2 (N14961, N14953, N12655);
and AND4 (N14962, N14958, N11088, N6477, N12779);
or OR2 (N14963, N14961, N1385);
buf BUF1 (N14964, N14959);
nor NOR3 (N14965, N14951, N13369, N14606);
buf BUF1 (N14966, N14960);
nand NAND4 (N14967, N14962, N3076, N8531, N7389);
and AND4 (N14968, N14949, N11400, N5428, N1206);
or OR2 (N14969, N14968, N3288);
not NOT1 (N14970, N14969);
or OR2 (N14971, N14957, N9496);
xor XOR2 (N14972, N14956, N14767);
xor XOR2 (N14973, N14966, N5810);
nor NOR4 (N14974, N14963, N9840, N11432, N4787);
nor NOR3 (N14975, N14974, N7145, N3957);
nor NOR3 (N14976, N14943, N14082, N14037);
nor NOR4 (N14977, N14967, N10107, N12249, N4756);
nor NOR4 (N14978, N14973, N11346, N10929, N5424);
buf BUF1 (N14979, N14975);
buf BUF1 (N14980, N14942);
nor NOR3 (N14981, N14971, N1348, N13926);
nor NOR2 (N14982, N14972, N7505);
nand NAND4 (N14983, N14976, N4777, N9357, N8250);
and AND3 (N14984, N14964, N13114, N10435);
xor XOR2 (N14985, N14981, N7329);
xor XOR2 (N14986, N14984, N4397);
nor NOR3 (N14987, N14965, N11133, N10232);
nor NOR3 (N14988, N14979, N3981, N6734);
nand NAND3 (N14989, N14988, N3667, N9878);
not NOT1 (N14990, N14982);
xor XOR2 (N14991, N14980, N10151);
and AND4 (N14992, N14978, N7354, N12819, N1070);
or OR4 (N14993, N14977, N14021, N10371, N8845);
nand NAND2 (N14994, N14992, N3431);
or OR3 (N14995, N14970, N1458, N13542);
or OR4 (N14996, N14986, N13821, N11157, N1829);
nor NOR4 (N14997, N14994, N5721, N7818, N10131);
nand NAND2 (N14998, N14991, N10187);
nor NOR3 (N14999, N14987, N6103, N3392);
or OR4 (N15000, N14989, N9364, N3259, N9154);
xor XOR2 (N15001, N14993, N1535);
buf BUF1 (N15002, N14999);
buf BUF1 (N15003, N14990);
nor NOR2 (N15004, N14985, N5326);
buf BUF1 (N15005, N14998);
and AND3 (N15006, N14983, N8891, N5752);
xor XOR2 (N15007, N15002, N1543);
nand NAND3 (N15008, N14996, N8183, N5359);
buf BUF1 (N15009, N15007);
or OR2 (N15010, N15006, N5652);
nor NOR4 (N15011, N14995, N6890, N12163, N1834);
xor XOR2 (N15012, N15003, N1184);
and AND3 (N15013, N14997, N13369, N11518);
nand NAND4 (N15014, N15013, N15000, N7043, N9904);
or OR4 (N15015, N3321, N10983, N2407, N3052);
nand NAND3 (N15016, N15005, N338, N1837);
buf BUF1 (N15017, N15009);
not NOT1 (N15018, N15010);
or OR3 (N15019, N15012, N2701, N13447);
and AND2 (N15020, N15015, N2180);
nor NOR4 (N15021, N15020, N6006, N1159, N13065);
or OR3 (N15022, N15011, N1033, N2423);
xor XOR2 (N15023, N15017, N8984);
nand NAND3 (N15024, N15019, N2752, N10978);
xor XOR2 (N15025, N15021, N11175);
nand NAND4 (N15026, N15023, N8808, N5648, N6240);
and AND3 (N15027, N15026, N6445, N646);
or OR3 (N15028, N15014, N6878, N3381);
nand NAND4 (N15029, N15028, N13748, N9639, N11073);
xor XOR2 (N15030, N15001, N8756);
and AND4 (N15031, N15030, N6061, N6021, N10331);
nand NAND3 (N15032, N15024, N14592, N2941);
nor NOR3 (N15033, N15029, N7774, N13663);
and AND2 (N15034, N15022, N8209);
buf BUF1 (N15035, N15032);
nor NOR4 (N15036, N15008, N1785, N5425, N10009);
nand NAND3 (N15037, N15025, N8813, N4079);
xor XOR2 (N15038, N15031, N14637);
nor NOR4 (N15039, N15034, N3275, N826, N5327);
buf BUF1 (N15040, N15035);
nor NOR4 (N15041, N15040, N3423, N10891, N12053);
or OR2 (N15042, N15027, N5363);
nand NAND2 (N15043, N15037, N14218);
nand NAND3 (N15044, N15042, N6840, N1743);
not NOT1 (N15045, N15039);
not NOT1 (N15046, N15004);
buf BUF1 (N15047, N15036);
buf BUF1 (N15048, N15043);
not NOT1 (N15049, N15038);
buf BUF1 (N15050, N15048);
or OR4 (N15051, N15049, N9652, N135, N13740);
xor XOR2 (N15052, N15041, N14893);
buf BUF1 (N15053, N15047);
nor NOR3 (N15054, N15050, N10434, N1880);
or OR3 (N15055, N15054, N3076, N14414);
or OR2 (N15056, N15044, N1403);
not NOT1 (N15057, N15046);
or OR4 (N15058, N15016, N10541, N12177, N14391);
nand NAND2 (N15059, N15053, N9155);
or OR3 (N15060, N15052, N5224, N11606);
or OR4 (N15061, N15057, N2702, N9499, N3080);
buf BUF1 (N15062, N15045);
nor NOR2 (N15063, N15059, N14873);
nand NAND3 (N15064, N15063, N8108, N12514);
and AND2 (N15065, N15064, N3025);
and AND3 (N15066, N15018, N10924, N14593);
or OR3 (N15067, N15056, N5525, N4480);
nor NOR2 (N15068, N15066, N8394);
nor NOR2 (N15069, N15061, N427);
or OR4 (N15070, N15055, N4572, N13046, N12030);
not NOT1 (N15071, N15058);
xor XOR2 (N15072, N15068, N561);
buf BUF1 (N15073, N15065);
or OR3 (N15074, N15051, N7882, N4508);
and AND2 (N15075, N15069, N599);
not NOT1 (N15076, N15060);
xor XOR2 (N15077, N15076, N7869);
not NOT1 (N15078, N15073);
buf BUF1 (N15079, N15077);
xor XOR2 (N15080, N15070, N1626);
not NOT1 (N15081, N15071);
not NOT1 (N15082, N15079);
not NOT1 (N15083, N15075);
not NOT1 (N15084, N15072);
or OR4 (N15085, N15081, N977, N6882, N12465);
xor XOR2 (N15086, N15082, N13863);
and AND4 (N15087, N15083, N2327, N7527, N11729);
buf BUF1 (N15088, N15085);
not NOT1 (N15089, N15074);
and AND4 (N15090, N15062, N12939, N14724, N5069);
xor XOR2 (N15091, N15089, N14054);
xor XOR2 (N15092, N15088, N9858);
or OR3 (N15093, N15086, N12949, N3075);
xor XOR2 (N15094, N15093, N3846);
and AND2 (N15095, N15033, N10552);
and AND3 (N15096, N15087, N10386, N1903);
nor NOR2 (N15097, N15080, N10839);
and AND2 (N15098, N15094, N4482);
nand NAND4 (N15099, N15091, N4464, N10497, N11839);
not NOT1 (N15100, N15096);
nor NOR2 (N15101, N15067, N764);
and AND4 (N15102, N15095, N3166, N713, N11224);
not NOT1 (N15103, N15097);
not NOT1 (N15104, N15078);
not NOT1 (N15105, N15090);
nand NAND3 (N15106, N15101, N4140, N13493);
xor XOR2 (N15107, N15105, N9043);
nor NOR3 (N15108, N15098, N6178, N2501);
buf BUF1 (N15109, N15103);
xor XOR2 (N15110, N15106, N8734);
and AND2 (N15111, N15100, N3210);
nand NAND2 (N15112, N15111, N587);
or OR2 (N15113, N15102, N12081);
nor NOR2 (N15114, N15109, N3817);
nand NAND4 (N15115, N15104, N3144, N6531, N14053);
not NOT1 (N15116, N15099);
nand NAND4 (N15117, N15108, N10822, N14496, N14810);
or OR4 (N15118, N15110, N2792, N977, N3754);
nand NAND4 (N15119, N15115, N7379, N2293, N13530);
and AND4 (N15120, N15117, N1106, N13144, N15104);
nor NOR4 (N15121, N15118, N14786, N12521, N8680);
xor XOR2 (N15122, N15084, N4623);
nor NOR4 (N15123, N15119, N9264, N6833, N10120);
and AND2 (N15124, N15114, N1710);
or OR4 (N15125, N15120, N3109, N5875, N3014);
nor NOR2 (N15126, N15112, N9751);
and AND4 (N15127, N15122, N11141, N8002, N4603);
nor NOR2 (N15128, N15126, N5619);
and AND4 (N15129, N15124, N7747, N3635, N3635);
buf BUF1 (N15130, N15092);
or OR4 (N15131, N15107, N12415, N14149, N7379);
nand NAND4 (N15132, N15125, N12763, N514, N656);
buf BUF1 (N15133, N15113);
buf BUF1 (N15134, N15128);
or OR3 (N15135, N15132, N3004, N12707);
xor XOR2 (N15136, N15135, N7882);
or OR2 (N15137, N15116, N2945);
nor NOR3 (N15138, N15136, N7925, N4015);
xor XOR2 (N15139, N15129, N7947);
and AND3 (N15140, N15130, N11830, N9453);
nand NAND2 (N15141, N15121, N4858);
not NOT1 (N15142, N15127);
or OR3 (N15143, N15139, N2747, N3980);
nor NOR3 (N15144, N15141, N6392, N6026);
buf BUF1 (N15145, N15123);
nand NAND2 (N15146, N15140, N1563);
and AND4 (N15147, N15137, N11783, N3868, N602);
not NOT1 (N15148, N15144);
or OR3 (N15149, N15142, N13908, N3904);
not NOT1 (N15150, N15145);
nand NAND4 (N15151, N15148, N11817, N9718, N5697);
not NOT1 (N15152, N15146);
or OR4 (N15153, N15133, N7624, N8125, N2060);
xor XOR2 (N15154, N15151, N7608);
and AND3 (N15155, N15149, N8884, N7087);
nand NAND3 (N15156, N15153, N14247, N1266);
nand NAND3 (N15157, N15134, N12952, N1366);
xor XOR2 (N15158, N15143, N14341);
and AND2 (N15159, N15157, N1671);
nor NOR4 (N15160, N15156, N9566, N5978, N4547);
not NOT1 (N15161, N15159);
or OR4 (N15162, N15131, N6233, N10087, N7339);
nor NOR3 (N15163, N15138, N5698, N5026);
buf BUF1 (N15164, N15161);
nor NOR4 (N15165, N15164, N3283, N3105, N9673);
nand NAND3 (N15166, N15147, N9909, N13336);
nor NOR2 (N15167, N15162, N456);
buf BUF1 (N15168, N15167);
xor XOR2 (N15169, N15166, N3497);
or OR4 (N15170, N15158, N3774, N8823, N1576);
or OR3 (N15171, N15152, N2133, N2219);
nor NOR4 (N15172, N15165, N9096, N5050, N2083);
buf BUF1 (N15173, N15170);
or OR2 (N15174, N15154, N10845);
buf BUF1 (N15175, N15172);
or OR4 (N15176, N15171, N8304, N14416, N8270);
and AND2 (N15177, N15163, N8672);
nor NOR4 (N15178, N15155, N4390, N14438, N14093);
buf BUF1 (N15179, N15173);
nor NOR3 (N15180, N15179, N2504, N8481);
and AND2 (N15181, N15174, N214);
not NOT1 (N15182, N15181);
nand NAND4 (N15183, N15176, N14332, N8763, N9968);
or OR4 (N15184, N15178, N8468, N3561, N9641);
nand NAND2 (N15185, N15177, N5617);
buf BUF1 (N15186, N15169);
and AND4 (N15187, N15175, N7776, N3865, N2982);
xor XOR2 (N15188, N15182, N9095);
buf BUF1 (N15189, N15168);
buf BUF1 (N15190, N15183);
buf BUF1 (N15191, N15189);
xor XOR2 (N15192, N15185, N9244);
xor XOR2 (N15193, N15160, N5708);
not NOT1 (N15194, N15188);
or OR4 (N15195, N15194, N13463, N7279, N4488);
not NOT1 (N15196, N15193);
nor NOR4 (N15197, N15196, N4135, N4915, N11933);
and AND2 (N15198, N15180, N10585);
and AND4 (N15199, N15197, N409, N10721, N15102);
nor NOR3 (N15200, N15191, N7242, N3644);
and AND2 (N15201, N15187, N11024);
xor XOR2 (N15202, N15192, N11097);
xor XOR2 (N15203, N15198, N12699);
nor NOR4 (N15204, N15150, N11733, N1017, N6436);
nand NAND2 (N15205, N15199, N14956);
not NOT1 (N15206, N15202);
buf BUF1 (N15207, N15205);
xor XOR2 (N15208, N15184, N9772);
xor XOR2 (N15209, N15201, N5379);
nand NAND4 (N15210, N15186, N2215, N10259, N11509);
buf BUF1 (N15211, N15207);
buf BUF1 (N15212, N15209);
and AND4 (N15213, N15200, N10706, N2326, N4101);
nor NOR2 (N15214, N15195, N14888);
nor NOR4 (N15215, N15214, N11369, N3440, N12874);
nand NAND4 (N15216, N15190, N3507, N13738, N5279);
or OR4 (N15217, N15216, N3926, N4566, N4183);
nand NAND3 (N15218, N15203, N9172, N10499);
or OR2 (N15219, N15211, N6545);
or OR3 (N15220, N15219, N6249, N11456);
not NOT1 (N15221, N15208);
xor XOR2 (N15222, N15206, N3710);
and AND3 (N15223, N15210, N12606, N1668);
nor NOR2 (N15224, N15213, N14739);
nand NAND4 (N15225, N15218, N9324, N15181, N10805);
and AND4 (N15226, N15222, N11751, N7544, N2416);
not NOT1 (N15227, N15220);
xor XOR2 (N15228, N15215, N11465);
buf BUF1 (N15229, N15204);
nand NAND3 (N15230, N15224, N12937, N5628);
not NOT1 (N15231, N15227);
nor NOR2 (N15232, N15217, N6983);
buf BUF1 (N15233, N15228);
and AND3 (N15234, N15229, N3863, N9135);
nand NAND3 (N15235, N15231, N13665, N4476);
buf BUF1 (N15236, N15233);
or OR4 (N15237, N15226, N12521, N6031, N11002);
nor NOR4 (N15238, N15236, N6459, N14634, N14441);
not NOT1 (N15239, N15234);
buf BUF1 (N15240, N15237);
not NOT1 (N15241, N15223);
and AND4 (N15242, N15221, N9890, N14954, N2298);
not NOT1 (N15243, N15225);
buf BUF1 (N15244, N15239);
nand NAND2 (N15245, N15244, N12685);
buf BUF1 (N15246, N15230);
and AND3 (N15247, N15238, N9995, N8552);
or OR2 (N15248, N15242, N8041);
not NOT1 (N15249, N15246);
buf BUF1 (N15250, N15243);
and AND2 (N15251, N15247, N3612);
nand NAND3 (N15252, N15248, N15008, N5753);
nand NAND3 (N15253, N15252, N5632, N3110);
and AND3 (N15254, N15250, N2863, N11361);
or OR3 (N15255, N15241, N11167, N1333);
nand NAND3 (N15256, N15253, N7853, N9775);
not NOT1 (N15257, N15255);
and AND2 (N15258, N15232, N12226);
or OR2 (N15259, N15245, N6405);
buf BUF1 (N15260, N15258);
or OR4 (N15261, N15256, N10352, N508, N10576);
nand NAND4 (N15262, N15254, N10182, N3035, N3567);
xor XOR2 (N15263, N15261, N3500);
and AND2 (N15264, N15257, N5805);
nand NAND3 (N15265, N15251, N14087, N12496);
or OR4 (N15266, N15265, N11803, N11214, N1245);
nor NOR2 (N15267, N15263, N5153);
nand NAND3 (N15268, N15212, N13982, N11514);
and AND4 (N15269, N15262, N4241, N14869, N9067);
buf BUF1 (N15270, N15235);
and AND4 (N15271, N15266, N9461, N1682, N14768);
or OR2 (N15272, N15267, N6812);
nor NOR2 (N15273, N15240, N14666);
or OR2 (N15274, N15268, N11027);
nor NOR4 (N15275, N15249, N1546, N14881, N10014);
nand NAND3 (N15276, N15273, N14636, N13365);
xor XOR2 (N15277, N15269, N1014);
and AND2 (N15278, N15277, N286);
not NOT1 (N15279, N15274);
not NOT1 (N15280, N15272);
and AND3 (N15281, N15270, N9081, N13019);
not NOT1 (N15282, N15275);
xor XOR2 (N15283, N15278, N3724);
nor NOR4 (N15284, N15282, N38, N11763, N576);
not NOT1 (N15285, N15259);
nor NOR2 (N15286, N15279, N4591);
and AND4 (N15287, N15276, N9559, N2006, N5210);
xor XOR2 (N15288, N15287, N10723);
xor XOR2 (N15289, N15280, N11531);
nor NOR4 (N15290, N15264, N6549, N7500, N4418);
and AND4 (N15291, N15281, N15016, N5242, N7001);
not NOT1 (N15292, N15291);
and AND3 (N15293, N15284, N2076, N569);
not NOT1 (N15294, N15286);
xor XOR2 (N15295, N15290, N13362);
buf BUF1 (N15296, N15295);
xor XOR2 (N15297, N15288, N3273);
buf BUF1 (N15298, N15289);
or OR3 (N15299, N15260, N877, N7285);
and AND3 (N15300, N15283, N1709, N1612);
or OR2 (N15301, N15285, N10705);
or OR4 (N15302, N15292, N6878, N6722, N5080);
nor NOR3 (N15303, N15299, N13004, N11589);
nor NOR3 (N15304, N15303, N13784, N3822);
and AND4 (N15305, N15294, N6898, N3442, N2728);
nor NOR4 (N15306, N15301, N869, N6440, N2398);
and AND2 (N15307, N15300, N1847);
nor NOR4 (N15308, N15306, N11511, N3737, N1388);
not NOT1 (N15309, N15304);
xor XOR2 (N15310, N15309, N12790);
and AND4 (N15311, N15293, N14633, N1736, N1359);
nand NAND2 (N15312, N15311, N3343);
or OR2 (N15313, N15302, N5603);
and AND2 (N15314, N15307, N2634);
nor NOR3 (N15315, N15312, N4585, N3121);
and AND3 (N15316, N15313, N1793, N15263);
not NOT1 (N15317, N15316);
buf BUF1 (N15318, N15317);
nand NAND3 (N15319, N15271, N3480, N866);
not NOT1 (N15320, N15319);
and AND3 (N15321, N15310, N1612, N15053);
nand NAND3 (N15322, N15296, N12754, N5618);
and AND2 (N15323, N15321, N14746);
and AND3 (N15324, N15314, N13562, N9351);
nor NOR3 (N15325, N15320, N1893, N13797);
nand NAND3 (N15326, N15298, N11362, N9657);
not NOT1 (N15327, N15308);
or OR3 (N15328, N15318, N14201, N9734);
not NOT1 (N15329, N15305);
xor XOR2 (N15330, N15328, N3337);
nor NOR2 (N15331, N15329, N6010);
buf BUF1 (N15332, N15326);
or OR4 (N15333, N15323, N9760, N10109, N1090);
or OR2 (N15334, N15327, N10425);
buf BUF1 (N15335, N15322);
nor NOR2 (N15336, N15324, N4188);
nor NOR4 (N15337, N15331, N12371, N14771, N7553);
nor NOR2 (N15338, N15297, N4384);
and AND4 (N15339, N15315, N1666, N4671, N5929);
buf BUF1 (N15340, N15335);
not NOT1 (N15341, N15333);
xor XOR2 (N15342, N15339, N8418);
xor XOR2 (N15343, N15337, N2397);
and AND4 (N15344, N15342, N2072, N11646, N12370);
and AND4 (N15345, N15344, N14749, N3138, N4181);
and AND3 (N15346, N15332, N155, N12739);
nor NOR3 (N15347, N15343, N9582, N7874);
nor NOR4 (N15348, N15336, N2453, N6346, N2389);
nand NAND4 (N15349, N15338, N8599, N1527, N10626);
nand NAND3 (N15350, N15346, N3256, N7602);
nor NOR3 (N15351, N15334, N906, N709);
not NOT1 (N15352, N15345);
not NOT1 (N15353, N15350);
and AND3 (N15354, N15352, N12732, N714);
or OR2 (N15355, N15354, N14455);
not NOT1 (N15356, N15340);
nand NAND4 (N15357, N15325, N13965, N431, N5012);
xor XOR2 (N15358, N15355, N12846);
or OR4 (N15359, N15349, N2272, N11783, N9284);
nor NOR3 (N15360, N15359, N6393, N1309);
nor NOR3 (N15361, N15357, N15106, N9823);
nor NOR4 (N15362, N15347, N915, N2369, N13259);
xor XOR2 (N15363, N15358, N5098);
nand NAND2 (N15364, N15330, N13732);
buf BUF1 (N15365, N15362);
nor NOR4 (N15366, N15353, N13882, N10170, N510);
nand NAND3 (N15367, N15360, N3266, N13734);
xor XOR2 (N15368, N15341, N11603);
buf BUF1 (N15369, N15361);
not NOT1 (N15370, N15367);
and AND3 (N15371, N15364, N14069, N1947);
not NOT1 (N15372, N15371);
xor XOR2 (N15373, N15368, N2858);
nor NOR3 (N15374, N15372, N11723, N13803);
and AND2 (N15375, N15370, N7531);
nor NOR3 (N15376, N15375, N1840, N819);
and AND3 (N15377, N15376, N12966, N13437);
nor NOR3 (N15378, N15366, N8352, N11902);
not NOT1 (N15379, N15378);
or OR4 (N15380, N15369, N7983, N8119, N9465);
not NOT1 (N15381, N15379);
xor XOR2 (N15382, N15373, N4204);
and AND4 (N15383, N15351, N2987, N13485, N3947);
or OR3 (N15384, N15381, N888, N8763);
and AND3 (N15385, N15365, N8862, N3500);
xor XOR2 (N15386, N15363, N13392);
nor NOR4 (N15387, N15380, N1125, N7318, N9649);
not NOT1 (N15388, N15386);
xor XOR2 (N15389, N15383, N11258);
nand NAND4 (N15390, N15377, N8726, N14907, N10029);
or OR2 (N15391, N15389, N6693);
buf BUF1 (N15392, N15387);
buf BUF1 (N15393, N15384);
xor XOR2 (N15394, N15393, N15237);
buf BUF1 (N15395, N15391);
or OR4 (N15396, N15348, N5735, N11393, N2910);
not NOT1 (N15397, N15356);
not NOT1 (N15398, N15396);
or OR4 (N15399, N15394, N11997, N3362, N10424);
nor NOR2 (N15400, N15374, N8458);
nor NOR2 (N15401, N15382, N12857);
xor XOR2 (N15402, N15401, N2325);
or OR4 (N15403, N15385, N5565, N14240, N15380);
xor XOR2 (N15404, N15397, N13932);
or OR2 (N15405, N15399, N3092);
not NOT1 (N15406, N15404);
xor XOR2 (N15407, N15395, N13699);
not NOT1 (N15408, N15405);
buf BUF1 (N15409, N15392);
nand NAND2 (N15410, N15402, N10527);
nor NOR4 (N15411, N15407, N10995, N6492, N5512);
and AND3 (N15412, N15406, N10486, N13223);
nor NOR2 (N15413, N15409, N7463);
nand NAND3 (N15414, N15388, N7239, N13691);
nand NAND3 (N15415, N15411, N12119, N7787);
not NOT1 (N15416, N15415);
or OR3 (N15417, N15416, N14526, N5855);
xor XOR2 (N15418, N15414, N1408);
nand NAND2 (N15419, N15408, N9066);
buf BUF1 (N15420, N15390);
nand NAND2 (N15421, N15420, N9906);
buf BUF1 (N15422, N15410);
nor NOR4 (N15423, N15419, N4411, N10057, N14028);
or OR2 (N15424, N15413, N14590);
nand NAND2 (N15425, N15422, N6276);
or OR2 (N15426, N15423, N7158);
or OR3 (N15427, N15426, N14468, N5702);
nor NOR3 (N15428, N15424, N10205, N3494);
nand NAND2 (N15429, N15412, N12172);
buf BUF1 (N15430, N15400);
buf BUF1 (N15431, N15398);
not NOT1 (N15432, N15425);
and AND4 (N15433, N15431, N8356, N760, N2431);
xor XOR2 (N15434, N15418, N8660);
xor XOR2 (N15435, N15434, N2261);
nand NAND4 (N15436, N15428, N3018, N9709, N592);
nand NAND2 (N15437, N15433, N11162);
nand NAND4 (N15438, N15435, N7654, N11615, N6483);
xor XOR2 (N15439, N15417, N14283);
and AND4 (N15440, N15439, N6894, N3138, N10197);
buf BUF1 (N15441, N15421);
xor XOR2 (N15442, N15436, N2124);
or OR2 (N15443, N15432, N12794);
and AND2 (N15444, N15429, N27);
and AND4 (N15445, N15442, N717, N8757, N11966);
nor NOR4 (N15446, N15440, N14763, N11925, N11038);
nor NOR3 (N15447, N15403, N10254, N124);
nor NOR2 (N15448, N15427, N1258);
not NOT1 (N15449, N15444);
xor XOR2 (N15450, N15446, N15238);
xor XOR2 (N15451, N15438, N14518);
nor NOR4 (N15452, N15441, N9668, N2067, N3173);
not NOT1 (N15453, N15437);
not NOT1 (N15454, N15430);
buf BUF1 (N15455, N15453);
nand NAND4 (N15456, N15455, N8305, N6447, N11226);
and AND2 (N15457, N15447, N14822);
buf BUF1 (N15458, N15448);
xor XOR2 (N15459, N15458, N11281);
xor XOR2 (N15460, N15456, N1147);
buf BUF1 (N15461, N15454);
nor NOR2 (N15462, N15461, N929);
xor XOR2 (N15463, N15457, N9669);
nand NAND2 (N15464, N15452, N7111);
or OR3 (N15465, N15450, N7873, N9370);
xor XOR2 (N15466, N15465, N7895);
nand NAND4 (N15467, N15464, N14507, N9036, N190);
and AND4 (N15468, N15467, N9199, N2349, N2378);
not NOT1 (N15469, N15462);
buf BUF1 (N15470, N15466);
buf BUF1 (N15471, N15445);
and AND3 (N15472, N15471, N1795, N13490);
xor XOR2 (N15473, N15451, N13247);
or OR2 (N15474, N15470, N179);
or OR2 (N15475, N15473, N7068);
nand NAND4 (N15476, N15469, N6296, N8751, N7103);
nor NOR2 (N15477, N15474, N12311);
or OR4 (N15478, N15472, N9200, N3812, N11025);
buf BUF1 (N15479, N15475);
or OR3 (N15480, N15478, N11939, N398);
buf BUF1 (N15481, N15479);
nand NAND4 (N15482, N15476, N2730, N7299, N1002);
not NOT1 (N15483, N15459);
or OR3 (N15484, N15449, N10487, N7812);
not NOT1 (N15485, N15463);
nand NAND4 (N15486, N15468, N14322, N5863, N14231);
buf BUF1 (N15487, N15460);
xor XOR2 (N15488, N15480, N10790);
nand NAND2 (N15489, N15483, N5157);
not NOT1 (N15490, N15485);
xor XOR2 (N15491, N15477, N13483);
nand NAND3 (N15492, N15484, N14861, N5013);
not NOT1 (N15493, N15492);
nand NAND4 (N15494, N15489, N13984, N6138, N658);
or OR4 (N15495, N15443, N5465, N5818, N15178);
xor XOR2 (N15496, N15482, N5343);
buf BUF1 (N15497, N15491);
not NOT1 (N15498, N15481);
not NOT1 (N15499, N15496);
xor XOR2 (N15500, N15498, N14579);
not NOT1 (N15501, N15497);
xor XOR2 (N15502, N15495, N7448);
nand NAND3 (N15503, N15500, N9090, N5329);
or OR3 (N15504, N15487, N6494, N15190);
nor NOR2 (N15505, N15494, N4127);
buf BUF1 (N15506, N15490);
xor XOR2 (N15507, N15488, N4198);
xor XOR2 (N15508, N15502, N12234);
nor NOR2 (N15509, N15499, N10809);
xor XOR2 (N15510, N15505, N14161);
not NOT1 (N15511, N15504);
and AND4 (N15512, N15507, N8864, N1244, N12230);
buf BUF1 (N15513, N15501);
buf BUF1 (N15514, N15493);
nor NOR2 (N15515, N15506, N11906);
xor XOR2 (N15516, N15515, N7675);
not NOT1 (N15517, N15509);
or OR2 (N15518, N15513, N10034);
or OR3 (N15519, N15508, N6070, N14241);
or OR2 (N15520, N15503, N4831);
not NOT1 (N15521, N15514);
nor NOR3 (N15522, N15512, N14194, N1782);
nand NAND3 (N15523, N15518, N5638, N15015);
nor NOR4 (N15524, N15523, N835, N995, N7242);
nor NOR4 (N15525, N15517, N4437, N208, N12543);
or OR3 (N15526, N15524, N3547, N7718);
and AND3 (N15527, N15511, N8284, N5442);
or OR4 (N15528, N15522, N14613, N14937, N5804);
buf BUF1 (N15529, N15510);
nor NOR2 (N15530, N15520, N9184);
not NOT1 (N15531, N15526);
or OR2 (N15532, N15528, N5603);
not NOT1 (N15533, N15532);
xor XOR2 (N15534, N15525, N7333);
not NOT1 (N15535, N15531);
not NOT1 (N15536, N15486);
or OR4 (N15537, N15527, N8732, N6559, N718);
nand NAND4 (N15538, N15521, N15170, N13047, N10152);
or OR2 (N15539, N15534, N12861);
not NOT1 (N15540, N15536);
xor XOR2 (N15541, N15519, N11118);
nand NAND3 (N15542, N15537, N3133, N12529);
buf BUF1 (N15543, N15535);
xor XOR2 (N15544, N15540, N5873);
and AND4 (N15545, N15539, N6526, N231, N12160);
nor NOR4 (N15546, N15516, N10901, N15131, N14160);
nand NAND4 (N15547, N15530, N12810, N3787, N1489);
and AND2 (N15548, N15547, N10435);
buf BUF1 (N15549, N15543);
and AND2 (N15550, N15533, N1397);
xor XOR2 (N15551, N15549, N4433);
nand NAND3 (N15552, N15548, N10771, N37);
xor XOR2 (N15553, N15529, N12602);
nand NAND4 (N15554, N15545, N8131, N10932, N1939);
nand NAND3 (N15555, N15553, N7511, N10310);
xor XOR2 (N15556, N15552, N11346);
nor NOR3 (N15557, N15542, N12179, N8553);
and AND4 (N15558, N15551, N539, N15519, N8505);
or OR4 (N15559, N15544, N1180, N3406, N4986);
buf BUF1 (N15560, N15541);
not NOT1 (N15561, N15550);
not NOT1 (N15562, N15557);
nand NAND3 (N15563, N15546, N13695, N2084);
and AND4 (N15564, N15559, N5697, N1710, N8333);
not NOT1 (N15565, N15561);
buf BUF1 (N15566, N15564);
or OR3 (N15567, N15560, N5660, N11681);
nand NAND3 (N15568, N15565, N1639, N192);
buf BUF1 (N15569, N15566);
not NOT1 (N15570, N15562);
xor XOR2 (N15571, N15556, N14087);
buf BUF1 (N15572, N15568);
nor NOR2 (N15573, N15563, N9795);
or OR3 (N15574, N15570, N4467, N2618);
buf BUF1 (N15575, N15567);
and AND3 (N15576, N15558, N3337, N13940);
and AND3 (N15577, N15554, N537, N5376);
nor NOR4 (N15578, N15576, N13365, N15274, N2371);
nand NAND4 (N15579, N15577, N11410, N10227, N7030);
nor NOR2 (N15580, N15575, N4380);
not NOT1 (N15581, N15574);
or OR4 (N15582, N15538, N1425, N12097, N13221);
not NOT1 (N15583, N15572);
nor NOR4 (N15584, N15571, N8541, N1020, N8986);
buf BUF1 (N15585, N15584);
or OR3 (N15586, N15583, N4873, N3447);
and AND3 (N15587, N15585, N2725, N6350);
or OR2 (N15588, N15586, N8889);
or OR4 (N15589, N15581, N15198, N11455, N5603);
and AND2 (N15590, N15569, N10848);
or OR4 (N15591, N15555, N12157, N10806, N13118);
and AND3 (N15592, N15587, N1589, N1693);
or OR4 (N15593, N15590, N12237, N3549, N518);
buf BUF1 (N15594, N15578);
not NOT1 (N15595, N15579);
not NOT1 (N15596, N15573);
nand NAND2 (N15597, N15592, N2002);
xor XOR2 (N15598, N15594, N6331);
nor NOR4 (N15599, N15597, N5493, N10364, N13543);
nand NAND4 (N15600, N15589, N9509, N3447, N11677);
nand NAND2 (N15601, N15588, N4621);
or OR3 (N15602, N15598, N12661, N2497);
xor XOR2 (N15603, N15601, N763);
buf BUF1 (N15604, N15596);
nor NOR4 (N15605, N15593, N5039, N9452, N5883);
buf BUF1 (N15606, N15604);
xor XOR2 (N15607, N15600, N9529);
and AND2 (N15608, N15603, N3668);
or OR3 (N15609, N15595, N7965, N4384);
buf BUF1 (N15610, N15602);
and AND2 (N15611, N15608, N1565);
not NOT1 (N15612, N15606);
not NOT1 (N15613, N15610);
xor XOR2 (N15614, N15609, N13094);
and AND4 (N15615, N15613, N15079, N2951, N15392);
nand NAND4 (N15616, N15615, N11457, N1540, N2948);
buf BUF1 (N15617, N15616);
buf BUF1 (N15618, N15611);
and AND4 (N15619, N15612, N9523, N11520, N11507);
or OR3 (N15620, N15605, N4545, N3243);
not NOT1 (N15621, N15599);
not NOT1 (N15622, N15607);
xor XOR2 (N15623, N15619, N1298);
nor NOR2 (N15624, N15622, N2991);
and AND2 (N15625, N15618, N9968);
xor XOR2 (N15626, N15591, N7158);
nand NAND4 (N15627, N15582, N3253, N10007, N12807);
or OR3 (N15628, N15580, N7294, N11046);
not NOT1 (N15629, N15626);
nor NOR3 (N15630, N15625, N2466, N963);
or OR3 (N15631, N15614, N2071, N2349);
xor XOR2 (N15632, N15621, N8751);
not NOT1 (N15633, N15627);
or OR4 (N15634, N15624, N3898, N9651, N12377);
and AND2 (N15635, N15620, N5384);
nand NAND4 (N15636, N15631, N4198, N2514, N5797);
nor NOR3 (N15637, N15632, N8994, N14452);
or OR3 (N15638, N15636, N14374, N1516);
and AND4 (N15639, N15628, N3314, N2715, N8304);
or OR2 (N15640, N15637, N4697);
and AND2 (N15641, N15640, N6645);
not NOT1 (N15642, N15635);
nor NOR4 (N15643, N15634, N9885, N1834, N3608);
not NOT1 (N15644, N15630);
not NOT1 (N15645, N15644);
and AND2 (N15646, N15639, N2971);
not NOT1 (N15647, N15617);
nand NAND2 (N15648, N15638, N4370);
nor NOR3 (N15649, N15629, N13856, N5519);
and AND2 (N15650, N15645, N15476);
buf BUF1 (N15651, N15648);
nand NAND2 (N15652, N15651, N615);
not NOT1 (N15653, N15623);
xor XOR2 (N15654, N15646, N11133);
buf BUF1 (N15655, N15642);
and AND3 (N15656, N15650, N6937, N10572);
xor XOR2 (N15657, N15656, N11458);
and AND4 (N15658, N15657, N13280, N13149, N1743);
and AND4 (N15659, N15643, N2672, N8582, N3237);
xor XOR2 (N15660, N15633, N2888);
not NOT1 (N15661, N15659);
buf BUF1 (N15662, N15654);
nor NOR4 (N15663, N15647, N10850, N4861, N1746);
or OR3 (N15664, N15649, N9915, N15212);
nor NOR3 (N15665, N15641, N8072, N12566);
and AND4 (N15666, N15660, N2352, N12877, N6785);
not NOT1 (N15667, N15653);
xor XOR2 (N15668, N15664, N15138);
xor XOR2 (N15669, N15666, N10461);
or OR4 (N15670, N15655, N14005, N7737, N7053);
not NOT1 (N15671, N15665);
not NOT1 (N15672, N15670);
nor NOR4 (N15673, N15663, N8523, N14707, N12210);
not NOT1 (N15674, N15652);
not NOT1 (N15675, N15668);
or OR3 (N15676, N15675, N11468, N1234);
buf BUF1 (N15677, N15658);
nor NOR3 (N15678, N15667, N3154, N10739);
xor XOR2 (N15679, N15661, N11242);
buf BUF1 (N15680, N15669);
and AND4 (N15681, N15679, N7058, N13901, N8739);
and AND4 (N15682, N15673, N13122, N2566, N7752);
buf BUF1 (N15683, N15662);
nor NOR3 (N15684, N15680, N12395, N2113);
nand NAND2 (N15685, N15676, N11695);
nor NOR4 (N15686, N15672, N14291, N2899, N11350);
nor NOR4 (N15687, N15674, N10422, N6696, N800);
nand NAND4 (N15688, N15671, N5846, N3180, N2140);
and AND4 (N15689, N15682, N11696, N9008, N3631);
not NOT1 (N15690, N15689);
and AND3 (N15691, N15677, N13168, N12219);
nand NAND4 (N15692, N15686, N3135, N5044, N5416);
nand NAND4 (N15693, N15691, N11178, N14425, N686);
or OR4 (N15694, N15693, N2523, N10372, N15525);
and AND3 (N15695, N15685, N9132, N715);
and AND4 (N15696, N15694, N14927, N526, N5288);
not NOT1 (N15697, N15696);
nand NAND4 (N15698, N15687, N14297, N8924, N12730);
nand NAND2 (N15699, N15684, N13619);
buf BUF1 (N15700, N15683);
nand NAND4 (N15701, N15681, N1087, N8637, N7637);
not NOT1 (N15702, N15701);
nor NOR3 (N15703, N15700, N14766, N11341);
nand NAND2 (N15704, N15703, N2995);
not NOT1 (N15705, N15704);
xor XOR2 (N15706, N15692, N295);
buf BUF1 (N15707, N15698);
nand NAND4 (N15708, N15706, N9438, N6877, N11623);
or OR2 (N15709, N15707, N5730);
xor XOR2 (N15710, N15708, N7013);
nor NOR4 (N15711, N15678, N508, N1960, N1875);
buf BUF1 (N15712, N15709);
buf BUF1 (N15713, N15712);
and AND2 (N15714, N15688, N1459);
or OR4 (N15715, N15713, N12918, N8305, N8988);
and AND2 (N15716, N15702, N11548);
xor XOR2 (N15717, N15690, N13256);
xor XOR2 (N15718, N15710, N11397);
not NOT1 (N15719, N15705);
buf BUF1 (N15720, N15715);
xor XOR2 (N15721, N15717, N9782);
nor NOR2 (N15722, N15721, N5033);
nand NAND2 (N15723, N15722, N9632);
not NOT1 (N15724, N15699);
nor NOR3 (N15725, N15697, N253, N5937);
nor NOR2 (N15726, N15723, N7033);
nand NAND2 (N15727, N15695, N8968);
nand NAND4 (N15728, N15714, N11669, N13208, N507);
xor XOR2 (N15729, N15716, N3567);
nor NOR3 (N15730, N15725, N10598, N2956);
xor XOR2 (N15731, N15720, N812);
or OR3 (N15732, N15724, N11104, N11820);
buf BUF1 (N15733, N15726);
or OR4 (N15734, N15719, N4327, N2316, N5121);
not NOT1 (N15735, N15711);
buf BUF1 (N15736, N15727);
or OR2 (N15737, N15731, N10747);
not NOT1 (N15738, N15733);
xor XOR2 (N15739, N15718, N6416);
xor XOR2 (N15740, N15729, N9575);
and AND3 (N15741, N15736, N716, N7172);
nand NAND2 (N15742, N15732, N702);
not NOT1 (N15743, N15728);
and AND4 (N15744, N15738, N3891, N12080, N5589);
nand NAND2 (N15745, N15730, N2849);
or OR3 (N15746, N15742, N4463, N2266);
nand NAND3 (N15747, N15734, N3333, N8866);
xor XOR2 (N15748, N15743, N7843);
or OR3 (N15749, N15740, N9163, N4729);
nor NOR3 (N15750, N15748, N3401, N14946);
or OR2 (N15751, N15749, N7170);
or OR2 (N15752, N15741, N2461);
nand NAND2 (N15753, N15752, N12820);
buf BUF1 (N15754, N15744);
buf BUF1 (N15755, N15746);
nand NAND3 (N15756, N15750, N13332, N542);
nand NAND4 (N15757, N15753, N4566, N13913, N15551);
or OR3 (N15758, N15737, N1763, N5553);
and AND3 (N15759, N15747, N4630, N658);
or OR2 (N15760, N15757, N7246);
nand NAND3 (N15761, N15758, N1348, N156);
nand NAND2 (N15762, N15756, N3546);
nor NOR4 (N15763, N15754, N3447, N4725, N4283);
nor NOR2 (N15764, N15760, N1034);
buf BUF1 (N15765, N15759);
nand NAND4 (N15766, N15765, N3504, N7448, N4756);
nor NOR3 (N15767, N15755, N14838, N11100);
nor NOR3 (N15768, N15766, N9370, N7899);
buf BUF1 (N15769, N15768);
buf BUF1 (N15770, N15769);
and AND2 (N15771, N15770, N82);
xor XOR2 (N15772, N15764, N4816);
nor NOR2 (N15773, N15772, N10144);
and AND4 (N15774, N15735, N7589, N10381, N7660);
and AND3 (N15775, N15774, N13898, N6468);
and AND3 (N15776, N15751, N3579, N9495);
xor XOR2 (N15777, N15773, N8180);
or OR4 (N15778, N15776, N4065, N11368, N1934);
and AND2 (N15779, N15771, N5916);
nand NAND2 (N15780, N15767, N13781);
nor NOR2 (N15781, N15778, N15721);
buf BUF1 (N15782, N15781);
xor XOR2 (N15783, N15780, N61);
nand NAND3 (N15784, N15745, N11722, N10637);
or OR2 (N15785, N15762, N12802);
and AND4 (N15786, N15763, N3726, N5036, N819);
not NOT1 (N15787, N15777);
buf BUF1 (N15788, N15784);
not NOT1 (N15789, N15787);
nor NOR3 (N15790, N15775, N5535, N15738);
nor NOR3 (N15791, N15785, N4187, N11999);
nand NAND2 (N15792, N15791, N4467);
or OR3 (N15793, N15779, N14526, N259);
buf BUF1 (N15794, N15793);
xor XOR2 (N15795, N15786, N4529);
nand NAND3 (N15796, N15795, N15458, N12540);
nand NAND3 (N15797, N15789, N14236, N2187);
not NOT1 (N15798, N15782);
nand NAND3 (N15799, N15794, N2246, N8027);
nor NOR4 (N15800, N15799, N6684, N4504, N9407);
xor XOR2 (N15801, N15797, N14003);
nor NOR3 (N15802, N15796, N6199, N14821);
and AND3 (N15803, N15792, N8815, N8115);
buf BUF1 (N15804, N15790);
or OR4 (N15805, N15783, N15129, N6437, N1995);
and AND2 (N15806, N15798, N3661);
nand NAND2 (N15807, N15788, N6675);
xor XOR2 (N15808, N15803, N3965);
buf BUF1 (N15809, N15761);
buf BUF1 (N15810, N15739);
buf BUF1 (N15811, N15805);
xor XOR2 (N15812, N15809, N270);
nor NOR3 (N15813, N15808, N4849, N3528);
nand NAND3 (N15814, N15810, N8863, N8442);
not NOT1 (N15815, N15811);
not NOT1 (N15816, N15804);
nand NAND2 (N15817, N15801, N14555);
and AND3 (N15818, N15800, N2829, N9125);
or OR4 (N15819, N15807, N3748, N3943, N6315);
and AND4 (N15820, N15806, N11015, N13431, N12579);
buf BUF1 (N15821, N15816);
xor XOR2 (N15822, N15813, N13879);
nor NOR4 (N15823, N15802, N2580, N1646, N14551);
or OR3 (N15824, N15820, N7990, N7591);
or OR2 (N15825, N15823, N988);
or OR2 (N15826, N15825, N14542);
nand NAND2 (N15827, N15824, N1143);
or OR3 (N15828, N15827, N10174, N875);
nand NAND4 (N15829, N15817, N2447, N7404, N12625);
not NOT1 (N15830, N15815);
nor NOR4 (N15831, N15829, N122, N15468, N14416);
nor NOR3 (N15832, N15831, N8691, N11978);
nor NOR4 (N15833, N15814, N887, N8357, N11476);
nor NOR2 (N15834, N15818, N9242);
not NOT1 (N15835, N15819);
nor NOR4 (N15836, N15828, N4785, N6609, N10094);
nand NAND2 (N15837, N15822, N8116);
not NOT1 (N15838, N15812);
xor XOR2 (N15839, N15821, N12761);
buf BUF1 (N15840, N15837);
xor XOR2 (N15841, N15840, N8000);
buf BUF1 (N15842, N15838);
and AND4 (N15843, N15832, N15146, N2817, N12866);
or OR4 (N15844, N15833, N8308, N1943, N1424);
nor NOR2 (N15845, N15835, N1883);
nand NAND3 (N15846, N15844, N7428, N11308);
buf BUF1 (N15847, N15845);
and AND3 (N15848, N15847, N14919, N7721);
nor NOR4 (N15849, N15846, N11416, N3352, N1698);
buf BUF1 (N15850, N15842);
or OR4 (N15851, N15843, N12390, N6508, N5560);
not NOT1 (N15852, N15849);
nand NAND3 (N15853, N15848, N2023, N4969);
and AND2 (N15854, N15830, N7510);
not NOT1 (N15855, N15850);
nor NOR2 (N15856, N15853, N14444);
buf BUF1 (N15857, N15851);
buf BUF1 (N15858, N15839);
not NOT1 (N15859, N15858);
xor XOR2 (N15860, N15852, N2685);
and AND3 (N15861, N15841, N12687, N1813);
nor NOR2 (N15862, N15826, N13332);
nand NAND2 (N15863, N15857, N12361);
or OR4 (N15864, N15856, N10821, N634, N8141);
nor NOR2 (N15865, N15861, N713);
and AND2 (N15866, N15854, N7722);
and AND4 (N15867, N15864, N4726, N6657, N12556);
not NOT1 (N15868, N15859);
not NOT1 (N15869, N15862);
not NOT1 (N15870, N15865);
xor XOR2 (N15871, N15834, N6613);
nor NOR4 (N15872, N15870, N12410, N13409, N4202);
not NOT1 (N15873, N15836);
nor NOR2 (N15874, N15871, N141);
not NOT1 (N15875, N15867);
xor XOR2 (N15876, N15872, N7776);
xor XOR2 (N15877, N15866, N11214);
and AND4 (N15878, N15863, N5120, N15765, N5693);
nand NAND2 (N15879, N15875, N7852);
nor NOR3 (N15880, N15855, N14970, N14362);
and AND2 (N15881, N15868, N11456);
and AND4 (N15882, N15874, N4093, N7458, N9911);
buf BUF1 (N15883, N15860);
xor XOR2 (N15884, N15882, N10541);
nor NOR4 (N15885, N15876, N5696, N15318, N2487);
xor XOR2 (N15886, N15880, N1037);
and AND4 (N15887, N15879, N9058, N8951, N5298);
buf BUF1 (N15888, N15887);
and AND3 (N15889, N15886, N9559, N9200);
not NOT1 (N15890, N15877);
buf BUF1 (N15891, N15888);
nand NAND3 (N15892, N15869, N2591, N10162);
and AND4 (N15893, N15891, N6459, N2320, N2519);
not NOT1 (N15894, N15884);
nor NOR2 (N15895, N15893, N2400);
not NOT1 (N15896, N15889);
and AND2 (N15897, N15894, N2572);
nor NOR4 (N15898, N15892, N2371, N13440, N11423);
nor NOR4 (N15899, N15885, N8949, N13341, N13506);
not NOT1 (N15900, N15895);
xor XOR2 (N15901, N15890, N4078);
and AND4 (N15902, N15899, N6813, N13293, N10770);
nand NAND4 (N15903, N15873, N1400, N930, N5409);
nand NAND2 (N15904, N15896, N3610);
buf BUF1 (N15905, N15881);
nand NAND3 (N15906, N15883, N6884, N590);
buf BUF1 (N15907, N15898);
nor NOR4 (N15908, N15907, N7963, N2237, N13052);
nand NAND3 (N15909, N15900, N6741, N9298);
or OR4 (N15910, N15903, N9252, N12004, N9538);
not NOT1 (N15911, N15897);
xor XOR2 (N15912, N15911, N12884);
xor XOR2 (N15913, N15901, N983);
xor XOR2 (N15914, N15908, N12887);
and AND3 (N15915, N15902, N3105, N7990);
xor XOR2 (N15916, N15878, N7902);
xor XOR2 (N15917, N15912, N1250);
xor XOR2 (N15918, N15916, N7303);
xor XOR2 (N15919, N15906, N5789);
xor XOR2 (N15920, N15904, N3222);
and AND3 (N15921, N15905, N15602, N11558);
xor XOR2 (N15922, N15917, N6377);
not NOT1 (N15923, N15913);
nand NAND2 (N15924, N15921, N1821);
and AND2 (N15925, N15919, N1);
and AND2 (N15926, N15918, N11776);
xor XOR2 (N15927, N15915, N6859);
not NOT1 (N15928, N15927);
nor NOR3 (N15929, N15909, N277, N2367);
nor NOR3 (N15930, N15928, N14130, N191);
not NOT1 (N15931, N15923);
xor XOR2 (N15932, N15931, N4095);
or OR3 (N15933, N15920, N11491, N6057);
nand NAND4 (N15934, N15933, N8807, N6614, N10609);
or OR4 (N15935, N15925, N441, N3911, N8261);
and AND4 (N15936, N15924, N185, N10489, N5668);
xor XOR2 (N15937, N15910, N12460);
not NOT1 (N15938, N15930);
or OR3 (N15939, N15922, N6468, N15426);
xor XOR2 (N15940, N15938, N3835);
not NOT1 (N15941, N15940);
nand NAND3 (N15942, N15929, N12286, N8210);
nand NAND2 (N15943, N15937, N5055);
nand NAND3 (N15944, N15942, N1237, N2147);
or OR4 (N15945, N15914, N7349, N4829, N14319);
or OR3 (N15946, N15939, N6885, N11494);
nor NOR4 (N15947, N15934, N1099, N11505, N513);
and AND4 (N15948, N15932, N5343, N8096, N12262);
nor NOR4 (N15949, N15947, N14884, N13988, N7386);
or OR2 (N15950, N15936, N5913);
buf BUF1 (N15951, N15950);
buf BUF1 (N15952, N15948);
not NOT1 (N15953, N15944);
xor XOR2 (N15954, N15945, N13137);
xor XOR2 (N15955, N15952, N5258);
nand NAND4 (N15956, N15935, N7698, N5351, N940);
and AND4 (N15957, N15956, N5884, N12128, N7544);
not NOT1 (N15958, N15957);
nand NAND2 (N15959, N15926, N14728);
and AND2 (N15960, N15958, N6506);
and AND3 (N15961, N15949, N5954, N13503);
and AND3 (N15962, N15951, N15676, N4654);
nand NAND4 (N15963, N15954, N15625, N7466, N4218);
not NOT1 (N15964, N15955);
or OR4 (N15965, N15960, N9919, N14299, N6746);
xor XOR2 (N15966, N15962, N1516);
nand NAND4 (N15967, N15964, N428, N4684, N15909);
xor XOR2 (N15968, N15966, N5786);
not NOT1 (N15969, N15941);
nand NAND2 (N15970, N15953, N9779);
not NOT1 (N15971, N15969);
nor NOR2 (N15972, N15961, N1866);
or OR2 (N15973, N15971, N250);
xor XOR2 (N15974, N15959, N12795);
and AND2 (N15975, N15974, N473);
xor XOR2 (N15976, N15968, N10672);
and AND4 (N15977, N15972, N4047, N9284, N9438);
not NOT1 (N15978, N15976);
xor XOR2 (N15979, N15975, N2457);
and AND2 (N15980, N15970, N10572);
buf BUF1 (N15981, N15943);
and AND3 (N15982, N15980, N5120, N9572);
nor NOR3 (N15983, N15977, N15635, N9785);
and AND4 (N15984, N15965, N5281, N2601, N204);
or OR2 (N15985, N15967, N1706);
not NOT1 (N15986, N15984);
xor XOR2 (N15987, N15985, N12198);
buf BUF1 (N15988, N15982);
or OR3 (N15989, N15978, N12764, N6788);
nor NOR2 (N15990, N15989, N4401);
and AND4 (N15991, N15988, N2907, N1814, N7119);
nand NAND3 (N15992, N15979, N12523, N7854);
xor XOR2 (N15993, N15990, N11507);
buf BUF1 (N15994, N15987);
nor NOR3 (N15995, N15991, N6876, N5796);
nor NOR2 (N15996, N15992, N6823);
buf BUF1 (N15997, N15983);
xor XOR2 (N15998, N15973, N22);
buf BUF1 (N15999, N15995);
buf BUF1 (N16000, N15981);
or OR4 (N16001, N15946, N6397, N11243, N12435);
nand NAND2 (N16002, N15999, N13314);
nand NAND2 (N16003, N15994, N3002);
and AND2 (N16004, N15997, N14330);
not NOT1 (N16005, N16003);
not NOT1 (N16006, N16000);
xor XOR2 (N16007, N15986, N15502);
buf BUF1 (N16008, N16001);
buf BUF1 (N16009, N16004);
nor NOR3 (N16010, N16002, N3179, N13181);
nor NOR4 (N16011, N16005, N2734, N7430, N15910);
nor NOR3 (N16012, N16010, N11765, N7961);
and AND2 (N16013, N15998, N5630);
or OR3 (N16014, N16008, N7692, N13685);
nor NOR4 (N16015, N16006, N1250, N4625, N5998);
xor XOR2 (N16016, N16014, N4531);
xor XOR2 (N16017, N15993, N15433);
buf BUF1 (N16018, N16017);
endmodule