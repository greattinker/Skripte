// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N25605,N25609,N25586,N25610,N25608,N25616,N25615,N25611,N25614,N25617;

xor XOR2 (N18, N11, N11);
buf BUF1 (N19, N3);
xor XOR2 (N20, N4, N1);
not NOT1 (N21, N17);
nor NOR2 (N22, N16, N20);
nor NOR2 (N23, N1, N18);
buf BUF1 (N24, N5);
buf BUF1 (N25, N5);
and AND4 (N26, N20, N16, N9, N19);
xor XOR2 (N27, N23, N15);
nand NAND3 (N28, N25, N12, N18);
xor XOR2 (N29, N6, N12);
nand NAND4 (N30, N26, N2, N22, N9);
buf BUF1 (N31, N25);
xor XOR2 (N32, N18, N9);
nor NOR4 (N33, N26, N19, N26, N32);
buf BUF1 (N34, N26);
not NOT1 (N35, N28);
or OR4 (N36, N25, N25, N4, N10);
nand NAND3 (N37, N27, N11, N26);
nand NAND2 (N38, N24, N25);
buf BUF1 (N39, N35);
nor NOR4 (N40, N36, N18, N26, N16);
nand NAND3 (N41, N39, N39, N22);
not NOT1 (N42, N37);
not NOT1 (N43, N38);
buf BUF1 (N44, N33);
xor XOR2 (N45, N40, N34);
or OR4 (N46, N31, N45, N11, N19);
not NOT1 (N47, N33);
nor NOR3 (N48, N45, N16, N29);
buf BUF1 (N49, N17);
nor NOR2 (N50, N30, N7);
nor NOR4 (N51, N44, N40, N45, N15);
and AND2 (N52, N41, N28);
not NOT1 (N53, N49);
not NOT1 (N54, N46);
not NOT1 (N55, N48);
nand NAND2 (N56, N55, N44);
buf BUF1 (N57, N53);
xor XOR2 (N58, N50, N32);
or OR2 (N59, N43, N7);
xor XOR2 (N60, N59, N34);
nor NOR3 (N61, N51, N32, N43);
nor NOR4 (N62, N61, N29, N3, N18);
not NOT1 (N63, N62);
or OR4 (N64, N60, N52, N23, N24);
and AND4 (N65, N37, N33, N25, N20);
nand NAND2 (N66, N63, N8);
buf BUF1 (N67, N64);
and AND2 (N68, N66, N14);
nor NOR4 (N69, N21, N17, N24, N36);
nor NOR4 (N70, N68, N36, N41, N68);
nand NAND3 (N71, N57, N69, N65);
and AND4 (N72, N68, N64, N36, N47);
buf BUF1 (N73, N72);
not NOT1 (N74, N3);
or OR3 (N75, N73, N48, N4);
or OR2 (N76, N10, N56);
xor XOR2 (N77, N49, N13);
nor NOR4 (N78, N67, N10, N13, N6);
buf BUF1 (N79, N74);
nand NAND3 (N80, N77, N36, N45);
buf BUF1 (N81, N80);
not NOT1 (N82, N79);
not NOT1 (N83, N54);
not NOT1 (N84, N81);
not NOT1 (N85, N76);
nand NAND2 (N86, N70, N18);
not NOT1 (N87, N82);
or OR4 (N88, N71, N45, N60, N20);
xor XOR2 (N89, N88, N63);
nor NOR2 (N90, N78, N86);
nor NOR3 (N91, N63, N45, N8);
nand NAND2 (N92, N90, N42);
and AND4 (N93, N61, N15, N26, N76);
nand NAND2 (N94, N85, N24);
nor NOR4 (N95, N83, N17, N31, N35);
buf BUF1 (N96, N87);
buf BUF1 (N97, N75);
or OR2 (N98, N96, N43);
buf BUF1 (N99, N98);
xor XOR2 (N100, N99, N63);
or OR3 (N101, N58, N35, N84);
nor NOR2 (N102, N61, N12);
buf BUF1 (N103, N102);
buf BUF1 (N104, N95);
not NOT1 (N105, N89);
nor NOR4 (N106, N100, N100, N1, N97);
nand NAND3 (N107, N40, N33, N25);
nor NOR4 (N108, N104, N41, N16, N99);
not NOT1 (N109, N108);
xor XOR2 (N110, N92, N47);
or OR4 (N111, N94, N48, N99, N78);
and AND3 (N112, N101, N35, N57);
xor XOR2 (N113, N110, N74);
not NOT1 (N114, N91);
buf BUF1 (N115, N103);
nor NOR2 (N116, N114, N14);
nor NOR4 (N117, N109, N58, N49, N50);
nand NAND3 (N118, N117, N66, N117);
not NOT1 (N119, N118);
xor XOR2 (N120, N105, N104);
nor NOR4 (N121, N115, N57, N25, N18);
and AND2 (N122, N121, N50);
buf BUF1 (N123, N107);
not NOT1 (N124, N120);
nor NOR2 (N125, N124, N109);
nor NOR2 (N126, N116, N38);
nor NOR3 (N127, N123, N82, N20);
and AND3 (N128, N122, N118, N41);
and AND4 (N129, N113, N126, N69, N61);
xor XOR2 (N130, N50, N91);
nand NAND3 (N131, N125, N85, N16);
or OR2 (N132, N128, N109);
and AND2 (N133, N127, N35);
xor XOR2 (N134, N93, N128);
or OR4 (N135, N131, N2, N78, N86);
and AND4 (N136, N130, N13, N24, N80);
xor XOR2 (N137, N133, N99);
nand NAND3 (N138, N112, N82, N10);
and AND3 (N139, N137, N45, N23);
and AND3 (N140, N111, N70, N85);
not NOT1 (N141, N119);
xor XOR2 (N142, N132, N4);
buf BUF1 (N143, N140);
nand NAND3 (N144, N141, N63, N37);
and AND3 (N145, N135, N13, N26);
nand NAND4 (N146, N145, N16, N97, N134);
nand NAND4 (N147, N141, N51, N47, N48);
xor XOR2 (N148, N129, N76);
or OR4 (N149, N146, N40, N107, N64);
xor XOR2 (N150, N148, N85);
not NOT1 (N151, N139);
nor NOR3 (N152, N106, N99, N13);
buf BUF1 (N153, N144);
or OR4 (N154, N138, N140, N18, N58);
nor NOR2 (N155, N149, N130);
buf BUF1 (N156, N155);
and AND3 (N157, N153, N58, N76);
nor NOR2 (N158, N143, N11);
nand NAND2 (N159, N150, N22);
buf BUF1 (N160, N142);
buf BUF1 (N161, N147);
nor NOR4 (N162, N160, N18, N159, N74);
xor XOR2 (N163, N115, N49);
nor NOR2 (N164, N156, N139);
and AND2 (N165, N154, N33);
nand NAND4 (N166, N136, N87, N136, N46);
buf BUF1 (N167, N165);
or OR2 (N168, N162, N126);
and AND3 (N169, N158, N24, N19);
nand NAND3 (N170, N161, N17, N90);
not NOT1 (N171, N152);
xor XOR2 (N172, N171, N124);
or OR4 (N173, N172, N27, N65, N172);
nor NOR4 (N174, N163, N142, N117, N50);
xor XOR2 (N175, N173, N58);
xor XOR2 (N176, N168, N115);
buf BUF1 (N177, N164);
not NOT1 (N178, N177);
nand NAND2 (N179, N170, N153);
or OR2 (N180, N174, N14);
nor NOR3 (N181, N157, N62, N54);
nand NAND2 (N182, N178, N143);
and AND3 (N183, N166, N14, N100);
buf BUF1 (N184, N180);
or OR2 (N185, N175, N84);
or OR2 (N186, N176, N166);
and AND4 (N187, N167, N85, N49, N105);
buf BUF1 (N188, N181);
or OR2 (N189, N179, N154);
nor NOR3 (N190, N182, N187, N113);
buf BUF1 (N191, N165);
buf BUF1 (N192, N185);
buf BUF1 (N193, N151);
not NOT1 (N194, N193);
and AND2 (N195, N184, N61);
nand NAND3 (N196, N191, N145, N49);
nand NAND2 (N197, N195, N55);
and AND3 (N198, N183, N176, N152);
nor NOR4 (N199, N190, N42, N156, N33);
nor NOR3 (N200, N169, N1, N44);
or OR4 (N201, N188, N22, N91, N62);
or OR4 (N202, N196, N45, N119, N26);
and AND2 (N203, N199, N109);
or OR2 (N204, N198, N108);
nand NAND3 (N205, N192, N143, N51);
or OR3 (N206, N202, N18, N35);
buf BUF1 (N207, N189);
nor NOR4 (N208, N203, N157, N67, N172);
buf BUF1 (N209, N201);
nor NOR3 (N210, N186, N187, N128);
nor NOR4 (N211, N209, N115, N118, N41);
xor XOR2 (N212, N210, N84);
not NOT1 (N213, N197);
buf BUF1 (N214, N207);
buf BUF1 (N215, N200);
and AND2 (N216, N215, N202);
nand NAND3 (N217, N216, N143, N120);
nor NOR3 (N218, N205, N131, N87);
nand NAND3 (N219, N214, N189, N203);
xor XOR2 (N220, N204, N42);
nand NAND3 (N221, N206, N192, N23);
nand NAND2 (N222, N220, N113);
not NOT1 (N223, N218);
not NOT1 (N224, N211);
and AND4 (N225, N224, N43, N63, N36);
xor XOR2 (N226, N222, N106);
xor XOR2 (N227, N194, N14);
xor XOR2 (N228, N212, N168);
or OR4 (N229, N228, N5, N189, N147);
buf BUF1 (N230, N208);
nand NAND2 (N231, N227, N108);
and AND2 (N232, N223, N153);
xor XOR2 (N233, N217, N201);
nand NAND3 (N234, N213, N70, N4);
or OR4 (N235, N231, N134, N219, N172);
or OR3 (N236, N2, N12, N40);
or OR4 (N237, N226, N206, N20, N97);
buf BUF1 (N238, N235);
and AND3 (N239, N237, N238, N61);
nor NOR4 (N240, N121, N218, N189, N60);
not NOT1 (N241, N233);
xor XOR2 (N242, N240, N192);
not NOT1 (N243, N230);
buf BUF1 (N244, N225);
and AND4 (N245, N239, N218, N238, N172);
xor XOR2 (N246, N221, N126);
or OR4 (N247, N236, N98, N173, N113);
nand NAND2 (N248, N242, N11);
buf BUF1 (N249, N229);
xor XOR2 (N250, N244, N51);
nor NOR2 (N251, N248, N126);
xor XOR2 (N252, N247, N10);
xor XOR2 (N253, N252, N70);
xor XOR2 (N254, N250, N52);
or OR4 (N255, N243, N143, N6, N207);
not NOT1 (N256, N246);
nand NAND4 (N257, N232, N179, N148, N58);
nand NAND2 (N258, N251, N39);
xor XOR2 (N259, N253, N191);
and AND3 (N260, N249, N100, N253);
nor NOR2 (N261, N257, N231);
xor XOR2 (N262, N255, N138);
or OR2 (N263, N262, N239);
not NOT1 (N264, N258);
buf BUF1 (N265, N261);
buf BUF1 (N266, N256);
xor XOR2 (N267, N241, N177);
xor XOR2 (N268, N265, N2);
or OR3 (N269, N264, N64, N68);
and AND4 (N270, N268, N87, N187, N18);
xor XOR2 (N271, N269, N173);
nand NAND4 (N272, N254, N259, N206, N4);
not NOT1 (N273, N95);
buf BUF1 (N274, N245);
and AND4 (N275, N270, N156, N259, N129);
nand NAND4 (N276, N234, N266, N207, N246);
buf BUF1 (N277, N208);
xor XOR2 (N278, N271, N161);
or OR2 (N279, N277, N11);
nand NAND3 (N280, N274, N195, N262);
not NOT1 (N281, N263);
or OR3 (N282, N281, N157, N181);
or OR2 (N283, N276, N108);
nand NAND3 (N284, N267, N93, N274);
nand NAND3 (N285, N283, N241, N16);
or OR4 (N286, N272, N146, N130, N95);
nor NOR3 (N287, N284, N173, N219);
or OR4 (N288, N273, N5, N222, N100);
not NOT1 (N289, N275);
or OR4 (N290, N286, N193, N130, N154);
xor XOR2 (N291, N278, N229);
and AND2 (N292, N287, N128);
xor XOR2 (N293, N290, N289);
and AND3 (N294, N140, N5, N189);
nand NAND3 (N295, N260, N216, N120);
nand NAND3 (N296, N294, N89, N33);
and AND3 (N297, N282, N288, N48);
nor NOR4 (N298, N199, N201, N97, N242);
nor NOR2 (N299, N298, N173);
nor NOR4 (N300, N295, N198, N284, N211);
nor NOR3 (N301, N296, N141, N95);
nand NAND3 (N302, N280, N189, N22);
xor XOR2 (N303, N300, N45);
xor XOR2 (N304, N297, N277);
nor NOR3 (N305, N299, N199, N267);
xor XOR2 (N306, N291, N105);
nand NAND3 (N307, N302, N290, N242);
nand NAND3 (N308, N292, N288, N28);
nor NOR3 (N309, N279, N202, N61);
xor XOR2 (N310, N304, N100);
xor XOR2 (N311, N285, N109);
and AND2 (N312, N307, N45);
nand NAND3 (N313, N301, N172, N211);
and AND3 (N314, N308, N112, N39);
and AND4 (N315, N312, N234, N219, N222);
xor XOR2 (N316, N314, N196);
and AND2 (N317, N305, N133);
and AND3 (N318, N309, N135, N96);
buf BUF1 (N319, N311);
buf BUF1 (N320, N313);
nor NOR2 (N321, N293, N268);
or OR4 (N322, N315, N58, N45, N281);
and AND4 (N323, N316, N312, N65, N247);
nor NOR2 (N324, N318, N301);
nor NOR3 (N325, N317, N110, N141);
nand NAND3 (N326, N303, N268, N102);
or OR4 (N327, N321, N22, N44, N14);
buf BUF1 (N328, N326);
or OR3 (N329, N310, N96, N2);
xor XOR2 (N330, N322, N35);
xor XOR2 (N331, N306, N26);
not NOT1 (N332, N319);
and AND3 (N333, N323, N15, N256);
nand NAND3 (N334, N325, N111, N185);
xor XOR2 (N335, N333, N265);
or OR2 (N336, N332, N127);
buf BUF1 (N337, N328);
buf BUF1 (N338, N331);
buf BUF1 (N339, N335);
nand NAND4 (N340, N338, N156, N267, N203);
nand NAND3 (N341, N327, N263, N302);
xor XOR2 (N342, N337, N6);
buf BUF1 (N343, N324);
nor NOR2 (N344, N330, N212);
xor XOR2 (N345, N341, N26);
not NOT1 (N346, N334);
nor NOR3 (N347, N344, N183, N264);
or OR3 (N348, N340, N35, N177);
or OR2 (N349, N336, N285);
xor XOR2 (N350, N320, N297);
nor NOR4 (N351, N347, N280, N163, N26);
or OR2 (N352, N351, N44);
and AND2 (N353, N349, N62);
nor NOR2 (N354, N348, N137);
nand NAND2 (N355, N343, N307);
not NOT1 (N356, N329);
nor NOR4 (N357, N339, N155, N238, N99);
not NOT1 (N358, N346);
xor XOR2 (N359, N356, N316);
xor XOR2 (N360, N359, N281);
or OR2 (N361, N353, N255);
nor NOR3 (N362, N345, N342, N306);
or OR2 (N363, N334, N197);
and AND4 (N364, N358, N188, N34, N313);
nor NOR4 (N365, N352, N77, N135, N361);
buf BUF1 (N366, N277);
not NOT1 (N367, N350);
not NOT1 (N368, N355);
nor NOR4 (N369, N367, N367, N63, N145);
xor XOR2 (N370, N368, N163);
or OR2 (N371, N370, N140);
nand NAND4 (N372, N360, N187, N298, N137);
nand NAND4 (N373, N362, N226, N295, N184);
or OR4 (N374, N357, N12, N262, N196);
and AND2 (N375, N369, N43);
or OR2 (N376, N375, N340);
buf BUF1 (N377, N372);
nand NAND2 (N378, N374, N282);
and AND4 (N379, N378, N336, N135, N89);
xor XOR2 (N380, N363, N43);
buf BUF1 (N381, N366);
nor NOR4 (N382, N365, N264, N27, N158);
not NOT1 (N383, N371);
and AND2 (N384, N381, N119);
and AND2 (N385, N354, N175);
and AND2 (N386, N373, N284);
and AND2 (N387, N383, N338);
nand NAND2 (N388, N386, N202);
nor NOR3 (N389, N385, N123, N261);
buf BUF1 (N390, N380);
not NOT1 (N391, N364);
not NOT1 (N392, N379);
nor NOR4 (N393, N391, N360, N156, N352);
nand NAND3 (N394, N387, N254, N208);
nand NAND3 (N395, N390, N118, N74);
xor XOR2 (N396, N394, N206);
buf BUF1 (N397, N382);
or OR3 (N398, N377, N34, N137);
not NOT1 (N399, N396);
buf BUF1 (N400, N393);
nor NOR3 (N401, N392, N293, N236);
or OR2 (N402, N397, N286);
or OR4 (N403, N398, N127, N214, N121);
and AND3 (N404, N395, N56, N42);
xor XOR2 (N405, N388, N135);
buf BUF1 (N406, N389);
or OR4 (N407, N403, N129, N209, N340);
and AND2 (N408, N400, N249);
nor NOR2 (N409, N399, N18);
nor NOR3 (N410, N409, N248, N167);
and AND2 (N411, N376, N132);
nand NAND3 (N412, N406, N67, N139);
not NOT1 (N413, N411);
nand NAND3 (N414, N407, N110, N261);
and AND4 (N415, N414, N390, N209, N160);
nand NAND3 (N416, N408, N82, N208);
or OR4 (N417, N412, N46, N68, N263);
and AND2 (N418, N404, N357);
and AND2 (N419, N384, N306);
nor NOR2 (N420, N401, N307);
xor XOR2 (N421, N419, N248);
buf BUF1 (N422, N420);
nor NOR4 (N423, N410, N36, N40, N197);
buf BUF1 (N424, N421);
buf BUF1 (N425, N413);
not NOT1 (N426, N425);
xor XOR2 (N427, N405, N216);
nand NAND4 (N428, N417, N143, N63, N295);
xor XOR2 (N429, N415, N145);
or OR3 (N430, N428, N337, N36);
xor XOR2 (N431, N427, N79);
buf BUF1 (N432, N426);
and AND3 (N433, N432, N213, N369);
nand NAND4 (N434, N430, N394, N365, N159);
or OR3 (N435, N429, N135, N217);
and AND3 (N436, N423, N325, N389);
and AND2 (N437, N422, N396);
nor NOR2 (N438, N436, N262);
xor XOR2 (N439, N437, N102);
nand NAND2 (N440, N418, N258);
or OR4 (N441, N424, N193, N192, N92);
not NOT1 (N442, N434);
and AND4 (N443, N438, N393, N406, N312);
not NOT1 (N444, N416);
or OR4 (N445, N402, N152, N107, N359);
nand NAND4 (N446, N443, N206, N105, N278);
buf BUF1 (N447, N439);
or OR3 (N448, N446, N141, N11);
or OR3 (N449, N448, N90, N182);
and AND2 (N450, N433, N197);
or OR3 (N451, N431, N79, N80);
or OR2 (N452, N447, N358);
not NOT1 (N453, N449);
buf BUF1 (N454, N453);
xor XOR2 (N455, N441, N367);
or OR3 (N456, N440, N89, N59);
nor NOR3 (N457, N456, N435, N348);
buf BUF1 (N458, N433);
xor XOR2 (N459, N444, N413);
not NOT1 (N460, N451);
not NOT1 (N461, N454);
nand NAND2 (N462, N459, N80);
buf BUF1 (N463, N452);
nor NOR2 (N464, N457, N443);
buf BUF1 (N465, N445);
nor NOR4 (N466, N461, N34, N30, N369);
xor XOR2 (N467, N464, N339);
nand NAND3 (N468, N463, N138, N6);
or OR4 (N469, N460, N37, N389, N195);
xor XOR2 (N470, N442, N443);
nor NOR4 (N471, N455, N15, N184, N84);
nand NAND4 (N472, N450, N362, N70, N337);
nand NAND3 (N473, N467, N154, N249);
or OR4 (N474, N468, N45, N29, N384);
or OR2 (N475, N465, N90);
not NOT1 (N476, N469);
buf BUF1 (N477, N472);
and AND3 (N478, N476, N266, N189);
nand NAND4 (N479, N477, N425, N459, N269);
or OR4 (N480, N462, N470, N37, N214);
xor XOR2 (N481, N49, N423);
buf BUF1 (N482, N466);
not NOT1 (N483, N473);
not NOT1 (N484, N483);
nor NOR3 (N485, N481, N403, N346);
or OR2 (N486, N458, N153);
or OR4 (N487, N484, N300, N424, N169);
nor NOR3 (N488, N475, N47, N287);
buf BUF1 (N489, N478);
xor XOR2 (N490, N474, N375);
buf BUF1 (N491, N482);
and AND2 (N492, N485, N1);
buf BUF1 (N493, N471);
and AND3 (N494, N487, N79, N376);
and AND2 (N495, N479, N78);
buf BUF1 (N496, N480);
and AND2 (N497, N492, N40);
nor NOR2 (N498, N497, N143);
xor XOR2 (N499, N489, N43);
nand NAND4 (N500, N498, N116, N39, N370);
buf BUF1 (N501, N500);
xor XOR2 (N502, N499, N190);
nor NOR4 (N503, N495, N282, N166, N45);
not NOT1 (N504, N493);
nand NAND2 (N505, N501, N125);
buf BUF1 (N506, N504);
nor NOR2 (N507, N503, N365);
buf BUF1 (N508, N494);
and AND4 (N509, N490, N286, N13, N347);
buf BUF1 (N510, N496);
nor NOR4 (N511, N505, N275, N124, N382);
nand NAND2 (N512, N507, N187);
nand NAND3 (N513, N509, N296, N232);
buf BUF1 (N514, N486);
and AND4 (N515, N488, N334, N169, N322);
xor XOR2 (N516, N508, N409);
not NOT1 (N517, N511);
nor NOR3 (N518, N512, N402, N15);
xor XOR2 (N519, N517, N286);
nor NOR3 (N520, N491, N481, N376);
not NOT1 (N521, N515);
not NOT1 (N522, N519);
not NOT1 (N523, N518);
nand NAND3 (N524, N506, N165, N406);
nor NOR4 (N525, N523, N24, N106, N373);
buf BUF1 (N526, N513);
and AND4 (N527, N525, N37, N119, N58);
not NOT1 (N528, N521);
not NOT1 (N529, N522);
or OR4 (N530, N526, N67, N281, N515);
or OR3 (N531, N514, N299, N396);
not NOT1 (N532, N527);
nor NOR2 (N533, N502, N55);
buf BUF1 (N534, N532);
nor NOR2 (N535, N530, N441);
and AND2 (N536, N516, N281);
not NOT1 (N537, N533);
nand NAND2 (N538, N537, N534);
nand NAND3 (N539, N388, N469, N235);
buf BUF1 (N540, N529);
xor XOR2 (N541, N538, N313);
not NOT1 (N542, N540);
and AND4 (N543, N510, N409, N303, N295);
xor XOR2 (N544, N536, N121);
not NOT1 (N545, N542);
or OR3 (N546, N541, N268, N252);
not NOT1 (N547, N535);
nor NOR4 (N548, N531, N296, N198, N525);
nor NOR2 (N549, N520, N491);
not NOT1 (N550, N524);
and AND3 (N551, N550, N374, N10);
nand NAND3 (N552, N539, N183, N491);
and AND4 (N553, N551, N416, N445, N334);
xor XOR2 (N554, N549, N449);
nand NAND4 (N555, N528, N388, N198, N55);
not NOT1 (N556, N545);
nor NOR3 (N557, N548, N252, N297);
xor XOR2 (N558, N555, N51);
buf BUF1 (N559, N547);
nand NAND2 (N560, N546, N282);
and AND4 (N561, N552, N295, N366, N92);
nand NAND2 (N562, N544, N187);
not NOT1 (N563, N557);
buf BUF1 (N564, N563);
or OR3 (N565, N562, N292, N53);
xor XOR2 (N566, N554, N125);
or OR2 (N567, N543, N137);
or OR4 (N568, N558, N32, N546, N323);
buf BUF1 (N569, N556);
nand NAND3 (N570, N568, N521, N51);
not NOT1 (N571, N570);
not NOT1 (N572, N567);
not NOT1 (N573, N572);
nand NAND4 (N574, N559, N495, N449, N552);
nand NAND2 (N575, N561, N255);
not NOT1 (N576, N575);
nor NOR3 (N577, N560, N267, N48);
and AND2 (N578, N564, N124);
nand NAND4 (N579, N574, N261, N101, N498);
nor NOR3 (N580, N578, N440, N429);
nand NAND3 (N581, N571, N420, N570);
nor NOR2 (N582, N566, N190);
xor XOR2 (N583, N582, N443);
nor NOR2 (N584, N553, N153);
not NOT1 (N585, N577);
nor NOR4 (N586, N569, N538, N149, N437);
not NOT1 (N587, N580);
nor NOR4 (N588, N587, N558, N92, N118);
xor XOR2 (N589, N586, N220);
nor NOR2 (N590, N581, N380);
buf BUF1 (N591, N588);
xor XOR2 (N592, N584, N20);
nand NAND2 (N593, N591, N308);
and AND2 (N594, N573, N246);
nand NAND4 (N595, N565, N316, N119, N534);
or OR3 (N596, N583, N140, N396);
nand NAND3 (N597, N593, N393, N121);
buf BUF1 (N598, N597);
nor NOR3 (N599, N596, N26, N260);
buf BUF1 (N600, N595);
and AND4 (N601, N598, N271, N67, N314);
nor NOR2 (N602, N592, N252);
and AND4 (N603, N599, N397, N410, N45);
not NOT1 (N604, N576);
or OR4 (N605, N589, N391, N352, N477);
not NOT1 (N606, N605);
or OR4 (N607, N600, N162, N433, N512);
nor NOR3 (N608, N601, N433, N25);
buf BUF1 (N609, N585);
nor NOR2 (N610, N590, N482);
not NOT1 (N611, N594);
xor XOR2 (N612, N607, N280);
buf BUF1 (N613, N579);
or OR2 (N614, N613, N599);
and AND4 (N615, N604, N420, N533, N550);
buf BUF1 (N616, N614);
or OR4 (N617, N612, N478, N307, N266);
or OR3 (N618, N606, N617, N442);
buf BUF1 (N619, N376);
or OR4 (N620, N608, N475, N315, N619);
nand NAND4 (N621, N123, N84, N442, N6);
buf BUF1 (N622, N609);
nand NAND4 (N623, N615, N556, N151, N32);
or OR2 (N624, N620, N412);
buf BUF1 (N625, N621);
nor NOR2 (N626, N616, N46);
not NOT1 (N627, N618);
and AND4 (N628, N626, N47, N278, N93);
and AND3 (N629, N625, N378, N87);
and AND3 (N630, N629, N257, N298);
nand NAND4 (N631, N611, N284, N107, N480);
nand NAND4 (N632, N622, N559, N159, N202);
not NOT1 (N633, N610);
buf BUF1 (N634, N633);
and AND2 (N635, N632, N623);
or OR3 (N636, N529, N289, N42);
xor XOR2 (N637, N636, N525);
and AND4 (N638, N603, N509, N589, N204);
not NOT1 (N639, N627);
and AND2 (N640, N631, N413);
or OR3 (N641, N628, N119, N507);
not NOT1 (N642, N630);
not NOT1 (N643, N641);
not NOT1 (N644, N624);
buf BUF1 (N645, N643);
buf BUF1 (N646, N639);
or OR3 (N647, N637, N420, N576);
xor XOR2 (N648, N645, N541);
nor NOR3 (N649, N634, N67, N243);
buf BUF1 (N650, N649);
buf BUF1 (N651, N635);
or OR3 (N652, N650, N628, N269);
xor XOR2 (N653, N638, N306);
nor NOR3 (N654, N640, N576, N443);
xor XOR2 (N655, N651, N154);
xor XOR2 (N656, N648, N473);
not NOT1 (N657, N652);
buf BUF1 (N658, N655);
not NOT1 (N659, N654);
nor NOR3 (N660, N657, N325, N428);
nand NAND3 (N661, N660, N478, N458);
not NOT1 (N662, N602);
buf BUF1 (N663, N656);
buf BUF1 (N664, N653);
not NOT1 (N665, N662);
xor XOR2 (N666, N646, N428);
nor NOR4 (N667, N642, N10, N465, N60);
xor XOR2 (N668, N664, N30);
xor XOR2 (N669, N659, N270);
or OR2 (N670, N661, N586);
nand NAND2 (N671, N644, N219);
or OR3 (N672, N647, N479, N172);
not NOT1 (N673, N670);
not NOT1 (N674, N672);
and AND3 (N675, N667, N213, N68);
not NOT1 (N676, N666);
nand NAND4 (N677, N668, N669, N46, N501);
buf BUF1 (N678, N572);
buf BUF1 (N679, N673);
buf BUF1 (N680, N665);
or OR2 (N681, N675, N637);
xor XOR2 (N682, N658, N504);
or OR2 (N683, N678, N446);
xor XOR2 (N684, N681, N503);
nand NAND4 (N685, N676, N568, N233, N61);
and AND3 (N686, N679, N684, N493);
nor NOR4 (N687, N685, N356, N223, N464);
nand NAND2 (N688, N564, N501);
xor XOR2 (N689, N671, N121);
nor NOR2 (N690, N677, N383);
nor NOR4 (N691, N687, N146, N639, N70);
nand NAND2 (N692, N682, N142);
buf BUF1 (N693, N663);
nand NAND4 (N694, N689, N43, N8, N438);
nor NOR3 (N695, N674, N118, N295);
or OR2 (N696, N688, N454);
xor XOR2 (N697, N690, N496);
buf BUF1 (N698, N693);
xor XOR2 (N699, N691, N123);
or OR2 (N700, N696, N476);
not NOT1 (N701, N686);
nand NAND2 (N702, N700, N660);
and AND2 (N703, N683, N132);
nand NAND2 (N704, N694, N646);
or OR2 (N705, N703, N328);
not NOT1 (N706, N698);
not NOT1 (N707, N697);
or OR4 (N708, N699, N542, N324, N5);
or OR2 (N709, N708, N526);
not NOT1 (N710, N707);
nand NAND4 (N711, N709, N9, N493, N589);
or OR4 (N712, N706, N626, N312, N155);
and AND2 (N713, N695, N97);
nand NAND4 (N714, N702, N586, N135, N362);
nor NOR2 (N715, N692, N52);
xor XOR2 (N716, N705, N27);
nor NOR4 (N717, N704, N91, N106, N507);
and AND4 (N718, N717, N7, N70, N541);
not NOT1 (N719, N701);
and AND2 (N720, N716, N236);
nand NAND2 (N721, N710, N118);
or OR4 (N722, N718, N584, N497, N310);
buf BUF1 (N723, N714);
not NOT1 (N724, N713);
not NOT1 (N725, N711);
nand NAND4 (N726, N720, N518, N495, N357);
or OR4 (N727, N724, N121, N576, N291);
xor XOR2 (N728, N723, N4);
buf BUF1 (N729, N727);
nand NAND3 (N730, N725, N443, N578);
buf BUF1 (N731, N722);
buf BUF1 (N732, N730);
or OR2 (N733, N719, N152);
not NOT1 (N734, N712);
xor XOR2 (N735, N732, N562);
xor XOR2 (N736, N729, N608);
nand NAND4 (N737, N721, N475, N456, N637);
xor XOR2 (N738, N735, N201);
nand NAND2 (N739, N733, N181);
or OR3 (N740, N738, N572, N582);
not NOT1 (N741, N728);
xor XOR2 (N742, N737, N481);
nand NAND2 (N743, N740, N142);
nor NOR3 (N744, N742, N295, N67);
nor NOR3 (N745, N731, N136, N451);
nand NAND3 (N746, N734, N583, N442);
nor NOR3 (N747, N736, N687, N349);
xor XOR2 (N748, N746, N109);
nor NOR4 (N749, N726, N378, N312, N27);
xor XOR2 (N750, N744, N511);
xor XOR2 (N751, N715, N25);
and AND2 (N752, N748, N525);
xor XOR2 (N753, N750, N304);
nor NOR2 (N754, N753, N568);
nor NOR3 (N755, N680, N156, N470);
nor NOR3 (N756, N755, N288, N325);
not NOT1 (N757, N739);
nand NAND2 (N758, N743, N241);
nor NOR4 (N759, N747, N91, N315, N300);
and AND2 (N760, N741, N686);
nand NAND3 (N761, N754, N64, N33);
or OR3 (N762, N745, N631, N326);
nor NOR3 (N763, N762, N190, N704);
not NOT1 (N764, N752);
nor NOR4 (N765, N764, N394, N215, N587);
and AND3 (N766, N758, N260, N366);
xor XOR2 (N767, N756, N620);
not NOT1 (N768, N751);
or OR2 (N769, N749, N117);
nor NOR2 (N770, N761, N178);
not NOT1 (N771, N768);
xor XOR2 (N772, N760, N464);
buf BUF1 (N773, N763);
or OR3 (N774, N771, N716, N353);
xor XOR2 (N775, N774, N734);
buf BUF1 (N776, N775);
xor XOR2 (N777, N766, N420);
and AND3 (N778, N776, N450, N218);
nor NOR4 (N779, N778, N410, N76, N501);
and AND4 (N780, N769, N244, N339, N276);
not NOT1 (N781, N772);
nor NOR3 (N782, N757, N187, N8);
xor XOR2 (N783, N767, N355);
nor NOR2 (N784, N782, N653);
nor NOR3 (N785, N784, N784, N330);
xor XOR2 (N786, N770, N406);
not NOT1 (N787, N783);
buf BUF1 (N788, N786);
or OR4 (N789, N765, N507, N267, N719);
nor NOR4 (N790, N773, N251, N11, N150);
buf BUF1 (N791, N781);
or OR3 (N792, N777, N583, N196);
and AND3 (N793, N780, N686, N573);
nor NOR3 (N794, N792, N189, N102);
nand NAND4 (N795, N793, N527, N73, N259);
and AND2 (N796, N787, N48);
and AND3 (N797, N794, N516, N128);
or OR3 (N798, N796, N73, N255);
buf BUF1 (N799, N779);
nor NOR3 (N800, N759, N42, N279);
xor XOR2 (N801, N795, N525);
nor NOR2 (N802, N791, N372);
not NOT1 (N803, N788);
or OR4 (N804, N802, N749, N658, N258);
buf BUF1 (N805, N804);
nand NAND2 (N806, N799, N519);
nand NAND3 (N807, N798, N774, N111);
and AND2 (N808, N807, N156);
xor XOR2 (N809, N800, N738);
nor NOR4 (N810, N808, N703, N228, N734);
not NOT1 (N811, N785);
nor NOR3 (N812, N790, N732, N61);
nor NOR4 (N813, N805, N60, N699, N701);
and AND4 (N814, N801, N659, N446, N217);
nand NAND2 (N815, N806, N684);
nor NOR4 (N816, N814, N641, N245, N561);
xor XOR2 (N817, N797, N546);
nand NAND2 (N818, N813, N84);
nor NOR2 (N819, N812, N239);
not NOT1 (N820, N809);
nand NAND4 (N821, N816, N9, N406, N761);
not NOT1 (N822, N789);
nand NAND2 (N823, N818, N140);
nor NOR4 (N824, N815, N328, N14, N743);
xor XOR2 (N825, N817, N464);
and AND2 (N826, N810, N32);
nand NAND4 (N827, N826, N132, N293, N293);
and AND4 (N828, N827, N157, N27, N473);
and AND3 (N829, N822, N275, N600);
xor XOR2 (N830, N829, N245);
not NOT1 (N831, N830);
nor NOR3 (N832, N811, N148, N575);
nor NOR2 (N833, N828, N783);
nor NOR4 (N834, N819, N640, N365, N398);
nor NOR2 (N835, N821, N572);
or OR4 (N836, N823, N231, N175, N497);
nand NAND3 (N837, N824, N761, N73);
buf BUF1 (N838, N825);
and AND4 (N839, N837, N575, N602, N752);
nand NAND4 (N840, N832, N437, N709, N359);
buf BUF1 (N841, N820);
not NOT1 (N842, N836);
not NOT1 (N843, N838);
nand NAND4 (N844, N843, N436, N67, N590);
and AND3 (N845, N835, N625, N192);
xor XOR2 (N846, N840, N754);
and AND2 (N847, N803, N706);
not NOT1 (N848, N847);
xor XOR2 (N849, N848, N16);
xor XOR2 (N850, N831, N549);
xor XOR2 (N851, N849, N749);
not NOT1 (N852, N844);
nand NAND4 (N853, N846, N656, N684, N444);
nor NOR2 (N854, N851, N811);
buf BUF1 (N855, N845);
xor XOR2 (N856, N833, N516);
and AND4 (N857, N855, N16, N830, N117);
nor NOR4 (N858, N852, N225, N508, N394);
nor NOR4 (N859, N834, N410, N623, N231);
and AND4 (N860, N857, N248, N338, N116);
not NOT1 (N861, N842);
or OR3 (N862, N859, N70, N318);
buf BUF1 (N863, N861);
nor NOR2 (N864, N863, N92);
and AND3 (N865, N858, N299, N140);
nand NAND3 (N866, N850, N340, N736);
and AND2 (N867, N853, N497);
nor NOR2 (N868, N865, N85);
buf BUF1 (N869, N868);
xor XOR2 (N870, N839, N198);
nand NAND4 (N871, N864, N95, N130, N332);
buf BUF1 (N872, N854);
nor NOR4 (N873, N860, N304, N276, N659);
nor NOR3 (N874, N856, N293, N228);
and AND2 (N875, N872, N226);
buf BUF1 (N876, N867);
not NOT1 (N877, N841);
and AND2 (N878, N866, N112);
and AND3 (N879, N877, N859, N688);
or OR4 (N880, N869, N753, N770, N865);
buf BUF1 (N881, N876);
not NOT1 (N882, N871);
xor XOR2 (N883, N875, N37);
or OR4 (N884, N878, N318, N498, N548);
not NOT1 (N885, N882);
buf BUF1 (N886, N881);
buf BUF1 (N887, N862);
not NOT1 (N888, N874);
buf BUF1 (N889, N883);
nand NAND4 (N890, N879, N481, N133, N356);
buf BUF1 (N891, N884);
buf BUF1 (N892, N873);
nor NOR3 (N893, N892, N118, N160);
not NOT1 (N894, N890);
not NOT1 (N895, N894);
not NOT1 (N896, N870);
xor XOR2 (N897, N887, N624);
buf BUF1 (N898, N888);
nor NOR2 (N899, N898, N195);
nor NOR2 (N900, N896, N660);
and AND4 (N901, N891, N632, N540, N783);
not NOT1 (N902, N885);
nand NAND2 (N903, N900, N693);
or OR2 (N904, N893, N683);
nor NOR4 (N905, N903, N126, N220, N861);
xor XOR2 (N906, N902, N244);
and AND4 (N907, N880, N566, N703, N854);
nand NAND2 (N908, N897, N131);
buf BUF1 (N909, N901);
buf BUF1 (N910, N895);
or OR3 (N911, N886, N246, N271);
or OR4 (N912, N899, N315, N524, N409);
nand NAND2 (N913, N910, N631);
not NOT1 (N914, N912);
xor XOR2 (N915, N914, N646);
and AND3 (N916, N909, N152, N763);
or OR3 (N917, N911, N114, N178);
nor NOR4 (N918, N908, N536, N310, N913);
nor NOR3 (N919, N62, N383, N852);
not NOT1 (N920, N917);
not NOT1 (N921, N919);
nor NOR3 (N922, N920, N502, N195);
not NOT1 (N923, N916);
nor NOR4 (N924, N921, N688, N270, N92);
and AND2 (N925, N924, N267);
nor NOR4 (N926, N889, N918, N426, N315);
buf BUF1 (N927, N34);
and AND4 (N928, N922, N843, N267, N90);
nand NAND2 (N929, N915, N198);
xor XOR2 (N930, N905, N247);
and AND4 (N931, N927, N573, N642, N919);
nand NAND3 (N932, N926, N402, N45);
nand NAND2 (N933, N904, N543);
not NOT1 (N934, N906);
not NOT1 (N935, N907);
not NOT1 (N936, N929);
nand NAND3 (N937, N923, N193, N486);
nor NOR4 (N938, N937, N215, N282, N822);
nand NAND2 (N939, N931, N275);
not NOT1 (N940, N935);
nor NOR2 (N941, N940, N889);
or OR4 (N942, N936, N185, N611, N368);
nor NOR3 (N943, N930, N844, N328);
xor XOR2 (N944, N938, N511);
nor NOR3 (N945, N928, N265, N57);
or OR2 (N946, N943, N597);
or OR4 (N947, N941, N747, N536, N61);
or OR3 (N948, N932, N519, N686);
not NOT1 (N949, N948);
nand NAND3 (N950, N934, N178, N709);
nand NAND2 (N951, N925, N715);
nor NOR2 (N952, N950, N774);
or OR2 (N953, N944, N595);
buf BUF1 (N954, N953);
or OR3 (N955, N949, N3, N630);
nand NAND4 (N956, N933, N474, N596, N643);
and AND3 (N957, N954, N237, N111);
nand NAND3 (N958, N957, N181, N75);
nor NOR2 (N959, N947, N339);
nand NAND4 (N960, N959, N613, N522, N314);
nor NOR3 (N961, N960, N337, N608);
nor NOR4 (N962, N951, N115, N453, N932);
xor XOR2 (N963, N939, N674);
or OR2 (N964, N956, N192);
or OR4 (N965, N942, N873, N891, N640);
buf BUF1 (N966, N946);
or OR2 (N967, N965, N104);
xor XOR2 (N968, N962, N693);
not NOT1 (N969, N952);
or OR2 (N970, N966, N478);
not NOT1 (N971, N968);
and AND4 (N972, N963, N9, N163, N794);
nand NAND2 (N973, N964, N334);
xor XOR2 (N974, N972, N24);
buf BUF1 (N975, N945);
or OR4 (N976, N973, N120, N236, N258);
not NOT1 (N977, N974);
and AND3 (N978, N955, N885, N225);
nand NAND2 (N979, N976, N353);
not NOT1 (N980, N961);
nor NOR4 (N981, N980, N220, N562, N330);
buf BUF1 (N982, N967);
not NOT1 (N983, N969);
buf BUF1 (N984, N977);
buf BUF1 (N985, N958);
or OR2 (N986, N985, N243);
and AND4 (N987, N970, N135, N182, N807);
nand NAND3 (N988, N971, N347, N186);
buf BUF1 (N989, N986);
and AND2 (N990, N984, N522);
or OR2 (N991, N975, N958);
or OR3 (N992, N988, N986, N880);
nor NOR3 (N993, N989, N721, N767);
xor XOR2 (N994, N993, N220);
nor NOR3 (N995, N981, N600, N80);
or OR2 (N996, N994, N250);
not NOT1 (N997, N987);
buf BUF1 (N998, N997);
xor XOR2 (N999, N978, N976);
nor NOR4 (N1000, N979, N227, N941, N782);
and AND3 (N1001, N992, N316, N134);
buf BUF1 (N1002, N990);
or OR3 (N1003, N998, N992, N228);
xor XOR2 (N1004, N995, N273);
and AND4 (N1005, N983, N294, N489, N649);
nand NAND4 (N1006, N991, N26, N83, N336);
xor XOR2 (N1007, N1003, N927);
not NOT1 (N1008, N982);
not NOT1 (N1009, N1005);
not NOT1 (N1010, N1009);
nand NAND3 (N1011, N1000, N780, N136);
not NOT1 (N1012, N1001);
or OR2 (N1013, N1011, N576);
nand NAND2 (N1014, N1008, N784);
not NOT1 (N1015, N999);
not NOT1 (N1016, N1007);
or OR4 (N1017, N1012, N674, N908, N675);
nor NOR4 (N1018, N1013, N285, N366, N905);
nor NOR2 (N1019, N1016, N122);
xor XOR2 (N1020, N1004, N540);
nand NAND4 (N1021, N1014, N146, N300, N265);
not NOT1 (N1022, N1015);
nor NOR3 (N1023, N1020, N653, N648);
or OR2 (N1024, N1018, N547);
nor NOR2 (N1025, N1017, N788);
xor XOR2 (N1026, N1010, N299);
or OR4 (N1027, N1023, N437, N699, N876);
nand NAND2 (N1028, N1002, N610);
buf BUF1 (N1029, N1025);
xor XOR2 (N1030, N1028, N522);
buf BUF1 (N1031, N1019);
not NOT1 (N1032, N1027);
not NOT1 (N1033, N1024);
xor XOR2 (N1034, N1029, N529);
nor NOR4 (N1035, N1031, N123, N233, N147);
nor NOR3 (N1036, N1032, N5, N976);
buf BUF1 (N1037, N996);
not NOT1 (N1038, N1035);
and AND4 (N1039, N1037, N66, N180, N45);
nor NOR4 (N1040, N1039, N924, N977, N95);
or OR2 (N1041, N1021, N131);
buf BUF1 (N1042, N1033);
nor NOR4 (N1043, N1034, N665, N735, N876);
not NOT1 (N1044, N1006);
not NOT1 (N1045, N1040);
not NOT1 (N1046, N1043);
xor XOR2 (N1047, N1038, N50);
and AND2 (N1048, N1044, N314);
not NOT1 (N1049, N1041);
nor NOR2 (N1050, N1030, N216);
or OR3 (N1051, N1050, N331, N571);
or OR4 (N1052, N1026, N722, N988, N698);
buf BUF1 (N1053, N1048);
not NOT1 (N1054, N1022);
xor XOR2 (N1055, N1046, N782);
not NOT1 (N1056, N1049);
not NOT1 (N1057, N1054);
or OR2 (N1058, N1052, N594);
nor NOR4 (N1059, N1058, N274, N309, N962);
nor NOR3 (N1060, N1055, N295, N941);
buf BUF1 (N1061, N1057);
xor XOR2 (N1062, N1045, N1052);
nand NAND2 (N1063, N1061, N509);
not NOT1 (N1064, N1060);
xor XOR2 (N1065, N1063, N197);
not NOT1 (N1066, N1064);
nor NOR2 (N1067, N1051, N904);
nor NOR4 (N1068, N1047, N886, N804, N983);
and AND4 (N1069, N1067, N836, N947, N53);
and AND4 (N1070, N1042, N967, N377, N367);
nor NOR4 (N1071, N1036, N85, N942, N365);
not NOT1 (N1072, N1071);
nand NAND4 (N1073, N1056, N369, N9, N1065);
buf BUF1 (N1074, N362);
xor XOR2 (N1075, N1053, N108);
or OR2 (N1076, N1066, N712);
or OR2 (N1077, N1075, N267);
nand NAND3 (N1078, N1072, N965, N465);
and AND3 (N1079, N1059, N5, N951);
not NOT1 (N1080, N1078);
nand NAND4 (N1081, N1077, N1068, N1049, N129);
or OR2 (N1082, N727, N772);
or OR3 (N1083, N1062, N766, N674);
not NOT1 (N1084, N1074);
nor NOR4 (N1085, N1083, N1040, N872, N862);
buf BUF1 (N1086, N1085);
and AND2 (N1087, N1070, N111);
xor XOR2 (N1088, N1076, N244);
xor XOR2 (N1089, N1086, N438);
nand NAND4 (N1090, N1081, N894, N595, N97);
nor NOR4 (N1091, N1084, N796, N296, N760);
or OR2 (N1092, N1079, N407);
nand NAND4 (N1093, N1082, N79, N726, N721);
and AND2 (N1094, N1069, N726);
or OR4 (N1095, N1087, N468, N917, N27);
nor NOR3 (N1096, N1090, N437, N921);
or OR4 (N1097, N1089, N484, N948, N967);
nor NOR4 (N1098, N1093, N216, N37, N875);
xor XOR2 (N1099, N1088, N742);
xor XOR2 (N1100, N1095, N673);
xor XOR2 (N1101, N1100, N960);
or OR3 (N1102, N1094, N395, N662);
nand NAND2 (N1103, N1092, N173);
buf BUF1 (N1104, N1097);
nand NAND4 (N1105, N1102, N266, N983, N984);
nand NAND2 (N1106, N1103, N616);
and AND3 (N1107, N1099, N872, N58);
or OR3 (N1108, N1107, N461, N460);
nand NAND4 (N1109, N1101, N67, N967, N501);
nand NAND2 (N1110, N1096, N179);
nand NAND3 (N1111, N1108, N552, N426);
not NOT1 (N1112, N1110);
and AND4 (N1113, N1112, N251, N83, N713);
nand NAND2 (N1114, N1073, N882);
nor NOR3 (N1115, N1114, N565, N669);
nand NAND4 (N1116, N1111, N562, N454, N154);
xor XOR2 (N1117, N1113, N1003);
and AND3 (N1118, N1098, N712, N307);
buf BUF1 (N1119, N1118);
nor NOR3 (N1120, N1109, N624, N1113);
not NOT1 (N1121, N1115);
buf BUF1 (N1122, N1116);
buf BUF1 (N1123, N1105);
buf BUF1 (N1124, N1091);
nor NOR4 (N1125, N1120, N784, N523, N312);
xor XOR2 (N1126, N1121, N1003);
not NOT1 (N1127, N1104);
nor NOR3 (N1128, N1106, N318, N173);
nor NOR3 (N1129, N1125, N441, N589);
xor XOR2 (N1130, N1123, N529);
buf BUF1 (N1131, N1126);
nand NAND2 (N1132, N1080, N251);
xor XOR2 (N1133, N1119, N599);
not NOT1 (N1134, N1117);
nor NOR2 (N1135, N1133, N184);
nand NAND4 (N1136, N1132, N986, N161, N189);
xor XOR2 (N1137, N1128, N425);
nand NAND4 (N1138, N1134, N282, N788, N975);
or OR3 (N1139, N1137, N1000, N25);
not NOT1 (N1140, N1139);
or OR4 (N1141, N1130, N667, N444, N555);
nor NOR2 (N1142, N1140, N388);
nor NOR3 (N1143, N1131, N771, N570);
or OR2 (N1144, N1124, N101);
nor NOR4 (N1145, N1143, N349, N1097, N701);
xor XOR2 (N1146, N1122, N540);
and AND2 (N1147, N1135, N482);
nor NOR4 (N1148, N1129, N315, N855, N1021);
xor XOR2 (N1149, N1146, N166);
or OR3 (N1150, N1148, N357, N1041);
or OR4 (N1151, N1138, N206, N1115, N538);
xor XOR2 (N1152, N1142, N372);
or OR2 (N1153, N1147, N519);
nand NAND3 (N1154, N1150, N879, N882);
and AND3 (N1155, N1136, N106, N520);
nor NOR2 (N1156, N1141, N194);
nor NOR3 (N1157, N1156, N581, N655);
and AND2 (N1158, N1145, N1070);
buf BUF1 (N1159, N1153);
xor XOR2 (N1160, N1155, N812);
nand NAND4 (N1161, N1157, N755, N828, N167);
and AND4 (N1162, N1151, N589, N417, N1132);
not NOT1 (N1163, N1152);
and AND3 (N1164, N1158, N59, N255);
not NOT1 (N1165, N1154);
nand NAND4 (N1166, N1162, N138, N1130, N764);
and AND3 (N1167, N1127, N55, N124);
nor NOR3 (N1168, N1161, N151, N1010);
nand NAND2 (N1169, N1149, N772);
and AND2 (N1170, N1144, N578);
buf BUF1 (N1171, N1169);
or OR2 (N1172, N1170, N754);
and AND4 (N1173, N1159, N1035, N602, N854);
nand NAND2 (N1174, N1168, N692);
and AND4 (N1175, N1167, N217, N324, N669);
and AND3 (N1176, N1175, N579, N498);
buf BUF1 (N1177, N1160);
nor NOR2 (N1178, N1166, N998);
not NOT1 (N1179, N1164);
or OR3 (N1180, N1171, N50, N95);
or OR2 (N1181, N1176, N162);
nor NOR4 (N1182, N1178, N1153, N513, N56);
nor NOR2 (N1183, N1179, N341);
nand NAND2 (N1184, N1183, N101);
or OR2 (N1185, N1173, N103);
nor NOR2 (N1186, N1181, N866);
nand NAND3 (N1187, N1184, N503, N1014);
and AND2 (N1188, N1163, N148);
xor XOR2 (N1189, N1174, N498);
not NOT1 (N1190, N1185);
nand NAND3 (N1191, N1188, N660, N586);
or OR4 (N1192, N1190, N700, N436, N657);
buf BUF1 (N1193, N1187);
nand NAND3 (N1194, N1186, N277, N124);
buf BUF1 (N1195, N1182);
xor XOR2 (N1196, N1172, N144);
or OR3 (N1197, N1180, N310, N137);
nor NOR2 (N1198, N1193, N1174);
nor NOR3 (N1199, N1195, N89, N1156);
not NOT1 (N1200, N1198);
or OR4 (N1201, N1165, N1021, N216, N565);
buf BUF1 (N1202, N1189);
nand NAND2 (N1203, N1200, N150);
nand NAND2 (N1204, N1192, N904);
xor XOR2 (N1205, N1191, N638);
xor XOR2 (N1206, N1196, N1120);
nand NAND4 (N1207, N1199, N51, N959, N1067);
and AND2 (N1208, N1201, N1194);
nand NAND2 (N1209, N792, N427);
not NOT1 (N1210, N1208);
or OR3 (N1211, N1205, N998, N1129);
and AND3 (N1212, N1197, N717, N939);
xor XOR2 (N1213, N1211, N878);
not NOT1 (N1214, N1204);
xor XOR2 (N1215, N1209, N661);
xor XOR2 (N1216, N1207, N256);
or OR4 (N1217, N1206, N124, N1163, N78);
or OR3 (N1218, N1212, N386, N830);
buf BUF1 (N1219, N1217);
nand NAND3 (N1220, N1210, N408, N580);
xor XOR2 (N1221, N1220, N32);
buf BUF1 (N1222, N1203);
and AND3 (N1223, N1222, N1166, N267);
or OR4 (N1224, N1221, N162, N311, N224);
or OR3 (N1225, N1218, N519, N98);
nand NAND4 (N1226, N1223, N112, N808, N595);
not NOT1 (N1227, N1225);
nand NAND3 (N1228, N1224, N140, N1067);
buf BUF1 (N1229, N1177);
xor XOR2 (N1230, N1214, N1087);
nor NOR4 (N1231, N1216, N1016, N1023, N1203);
and AND4 (N1232, N1229, N433, N688, N188);
not NOT1 (N1233, N1228);
buf BUF1 (N1234, N1232);
nor NOR3 (N1235, N1234, N512, N796);
or OR3 (N1236, N1202, N767, N723);
or OR3 (N1237, N1233, N939, N100);
nand NAND2 (N1238, N1230, N1200);
nand NAND2 (N1239, N1215, N501);
buf BUF1 (N1240, N1235);
not NOT1 (N1241, N1219);
and AND4 (N1242, N1236, N83, N1166, N75);
nor NOR2 (N1243, N1226, N697);
and AND3 (N1244, N1241, N448, N1104);
buf BUF1 (N1245, N1227);
nor NOR2 (N1246, N1245, N435);
xor XOR2 (N1247, N1246, N593);
nand NAND2 (N1248, N1239, N1093);
xor XOR2 (N1249, N1247, N887);
nor NOR2 (N1250, N1240, N974);
nor NOR4 (N1251, N1250, N473, N1076, N237);
and AND2 (N1252, N1231, N1243);
xor XOR2 (N1253, N147, N817);
xor XOR2 (N1254, N1249, N217);
and AND4 (N1255, N1238, N1210, N1023, N408);
buf BUF1 (N1256, N1255);
or OR2 (N1257, N1213, N490);
buf BUF1 (N1258, N1253);
nand NAND4 (N1259, N1257, N383, N1168, N452);
nand NAND2 (N1260, N1259, N416);
xor XOR2 (N1261, N1237, N1134);
not NOT1 (N1262, N1244);
buf BUF1 (N1263, N1262);
xor XOR2 (N1264, N1254, N1020);
not NOT1 (N1265, N1264);
xor XOR2 (N1266, N1251, N630);
xor XOR2 (N1267, N1265, N241);
nor NOR3 (N1268, N1266, N1267, N1167);
nand NAND3 (N1269, N600, N633, N1149);
not NOT1 (N1270, N1252);
not NOT1 (N1271, N1268);
or OR2 (N1272, N1270, N1131);
buf BUF1 (N1273, N1256);
nor NOR3 (N1274, N1273, N969, N1094);
or OR2 (N1275, N1258, N1139);
nor NOR2 (N1276, N1272, N142);
xor XOR2 (N1277, N1269, N763);
xor XOR2 (N1278, N1248, N153);
and AND3 (N1279, N1261, N894, N1254);
nand NAND4 (N1280, N1260, N711, N374, N963);
and AND3 (N1281, N1275, N415, N106);
nand NAND2 (N1282, N1277, N572);
xor XOR2 (N1283, N1281, N327);
buf BUF1 (N1284, N1242);
nor NOR3 (N1285, N1274, N565, N506);
not NOT1 (N1286, N1284);
nor NOR3 (N1287, N1286, N686, N827);
and AND3 (N1288, N1278, N1125, N368);
nor NOR3 (N1289, N1263, N346, N1129);
not NOT1 (N1290, N1287);
buf BUF1 (N1291, N1285);
nand NAND3 (N1292, N1279, N896, N550);
nand NAND2 (N1293, N1292, N545);
and AND3 (N1294, N1271, N974, N604);
buf BUF1 (N1295, N1282);
nand NAND4 (N1296, N1293, N1232, N578, N716);
or OR2 (N1297, N1294, N345);
nor NOR2 (N1298, N1276, N668);
buf BUF1 (N1299, N1295);
not NOT1 (N1300, N1290);
xor XOR2 (N1301, N1298, N995);
nand NAND3 (N1302, N1299, N988, N445);
xor XOR2 (N1303, N1300, N217);
or OR2 (N1304, N1283, N609);
not NOT1 (N1305, N1301);
and AND3 (N1306, N1291, N338, N554);
and AND3 (N1307, N1289, N1023, N572);
or OR2 (N1308, N1296, N391);
nor NOR4 (N1309, N1297, N447, N10, N178);
or OR3 (N1310, N1302, N796, N723);
or OR3 (N1311, N1280, N1278, N864);
nor NOR4 (N1312, N1310, N803, N330, N306);
xor XOR2 (N1313, N1304, N274);
not NOT1 (N1314, N1311);
nor NOR4 (N1315, N1308, N951, N1049, N118);
nand NAND3 (N1316, N1313, N1260, N1143);
buf BUF1 (N1317, N1307);
and AND2 (N1318, N1288, N710);
and AND3 (N1319, N1305, N1176, N1142);
not NOT1 (N1320, N1318);
not NOT1 (N1321, N1312);
nor NOR3 (N1322, N1306, N489, N1272);
xor XOR2 (N1323, N1315, N1037);
and AND2 (N1324, N1317, N959);
and AND4 (N1325, N1320, N1112, N1031, N40);
or OR3 (N1326, N1303, N502, N110);
or OR3 (N1327, N1309, N757, N861);
nand NAND4 (N1328, N1314, N869, N314, N476);
xor XOR2 (N1329, N1324, N1319);
or OR3 (N1330, N630, N900, N1149);
nor NOR3 (N1331, N1330, N987, N420);
not NOT1 (N1332, N1325);
nand NAND4 (N1333, N1316, N1053, N788, N1101);
xor XOR2 (N1334, N1323, N243);
buf BUF1 (N1335, N1329);
and AND2 (N1336, N1327, N772);
and AND4 (N1337, N1333, N498, N1131, N969);
and AND3 (N1338, N1328, N566, N49);
and AND4 (N1339, N1336, N856, N612, N806);
xor XOR2 (N1340, N1334, N773);
and AND3 (N1341, N1337, N848, N453);
buf BUF1 (N1342, N1322);
nand NAND4 (N1343, N1332, N1251, N566, N95);
and AND3 (N1344, N1326, N527, N944);
or OR2 (N1345, N1335, N378);
or OR2 (N1346, N1321, N101);
and AND2 (N1347, N1342, N191);
xor XOR2 (N1348, N1341, N964);
not NOT1 (N1349, N1346);
nor NOR3 (N1350, N1344, N1237, N118);
or OR3 (N1351, N1347, N286, N843);
not NOT1 (N1352, N1340);
or OR4 (N1353, N1339, N787, N366, N784);
and AND4 (N1354, N1343, N583, N831, N1290);
buf BUF1 (N1355, N1345);
nand NAND3 (N1356, N1351, N122, N683);
or OR2 (N1357, N1350, N815);
buf BUF1 (N1358, N1355);
and AND4 (N1359, N1354, N1229, N17, N946);
nor NOR3 (N1360, N1348, N341, N726);
not NOT1 (N1361, N1349);
nand NAND2 (N1362, N1357, N500);
xor XOR2 (N1363, N1358, N1299);
xor XOR2 (N1364, N1331, N859);
or OR2 (N1365, N1359, N5);
nand NAND2 (N1366, N1364, N595);
nor NOR3 (N1367, N1366, N614, N740);
not NOT1 (N1368, N1352);
buf BUF1 (N1369, N1360);
xor XOR2 (N1370, N1363, N310);
nor NOR2 (N1371, N1367, N1240);
not NOT1 (N1372, N1361);
not NOT1 (N1373, N1369);
not NOT1 (N1374, N1373);
nor NOR2 (N1375, N1353, N856);
xor XOR2 (N1376, N1372, N67);
nand NAND2 (N1377, N1365, N14);
not NOT1 (N1378, N1370);
and AND2 (N1379, N1375, N181);
or OR3 (N1380, N1374, N816, N568);
not NOT1 (N1381, N1356);
buf BUF1 (N1382, N1379);
nand NAND2 (N1383, N1376, N1248);
not NOT1 (N1384, N1381);
and AND2 (N1385, N1371, N647);
nand NAND2 (N1386, N1377, N430);
not NOT1 (N1387, N1380);
buf BUF1 (N1388, N1378);
xor XOR2 (N1389, N1386, N933);
xor XOR2 (N1390, N1385, N563);
or OR2 (N1391, N1388, N426);
buf BUF1 (N1392, N1382);
and AND2 (N1393, N1368, N599);
buf BUF1 (N1394, N1383);
or OR2 (N1395, N1394, N778);
xor XOR2 (N1396, N1392, N914);
xor XOR2 (N1397, N1396, N635);
or OR2 (N1398, N1393, N1213);
xor XOR2 (N1399, N1397, N566);
and AND4 (N1400, N1398, N505, N872, N196);
nand NAND4 (N1401, N1400, N990, N82, N69);
nor NOR3 (N1402, N1391, N1273, N652);
buf BUF1 (N1403, N1389);
and AND2 (N1404, N1338, N252);
and AND2 (N1405, N1390, N170);
and AND3 (N1406, N1387, N553, N510);
xor XOR2 (N1407, N1362, N259);
xor XOR2 (N1408, N1402, N1263);
nand NAND2 (N1409, N1407, N1121);
and AND4 (N1410, N1384, N550, N888, N412);
nand NAND2 (N1411, N1408, N1333);
nor NOR3 (N1412, N1404, N932, N613);
xor XOR2 (N1413, N1411, N412);
nand NAND4 (N1414, N1399, N506, N143, N1145);
nand NAND3 (N1415, N1395, N594, N551);
nand NAND4 (N1416, N1413, N1248, N1168, N18);
and AND4 (N1417, N1405, N1304, N1309, N638);
nor NOR4 (N1418, N1412, N633, N1182, N1009);
not NOT1 (N1419, N1415);
xor XOR2 (N1420, N1409, N527);
and AND3 (N1421, N1417, N16, N899);
and AND3 (N1422, N1403, N491, N229);
nor NOR4 (N1423, N1420, N615, N937, N503);
buf BUF1 (N1424, N1406);
and AND4 (N1425, N1418, N1249, N417, N730);
or OR4 (N1426, N1421, N1361, N1034, N1133);
buf BUF1 (N1427, N1410);
or OR4 (N1428, N1424, N1353, N992, N662);
and AND2 (N1429, N1401, N1275);
and AND2 (N1430, N1429, N834);
and AND4 (N1431, N1428, N52, N938, N590);
xor XOR2 (N1432, N1423, N1405);
and AND3 (N1433, N1419, N619, N689);
xor XOR2 (N1434, N1427, N1102);
nor NOR3 (N1435, N1414, N862, N958);
nor NOR4 (N1436, N1430, N91, N9, N810);
nand NAND3 (N1437, N1435, N1238, N308);
not NOT1 (N1438, N1431);
and AND3 (N1439, N1437, N236, N492);
buf BUF1 (N1440, N1416);
buf BUF1 (N1441, N1434);
nand NAND4 (N1442, N1433, N1384, N1355, N1364);
and AND3 (N1443, N1440, N994, N62);
xor XOR2 (N1444, N1436, N41);
nand NAND2 (N1445, N1438, N550);
buf BUF1 (N1446, N1425);
buf BUF1 (N1447, N1426);
buf BUF1 (N1448, N1441);
nor NOR3 (N1449, N1442, N1221, N768);
nor NOR4 (N1450, N1432, N777, N670, N598);
nand NAND4 (N1451, N1447, N819, N1132, N878);
or OR2 (N1452, N1449, N683);
buf BUF1 (N1453, N1451);
buf BUF1 (N1454, N1452);
and AND2 (N1455, N1445, N615);
or OR4 (N1456, N1454, N1159, N150, N775);
nand NAND3 (N1457, N1448, N134, N1023);
buf BUF1 (N1458, N1457);
buf BUF1 (N1459, N1453);
or OR4 (N1460, N1456, N385, N124, N1152);
buf BUF1 (N1461, N1459);
or OR4 (N1462, N1461, N833, N667, N1355);
buf BUF1 (N1463, N1450);
xor XOR2 (N1464, N1443, N434);
and AND4 (N1465, N1422, N1283, N298, N801);
nor NOR2 (N1466, N1455, N1243);
nor NOR4 (N1467, N1444, N1332, N14, N1283);
nor NOR4 (N1468, N1439, N397, N209, N1072);
buf BUF1 (N1469, N1446);
buf BUF1 (N1470, N1464);
xor XOR2 (N1471, N1462, N57);
or OR3 (N1472, N1458, N843, N805);
nor NOR2 (N1473, N1460, N308);
or OR4 (N1474, N1469, N699, N982, N1425);
nand NAND4 (N1475, N1473, N690, N1107, N727);
nand NAND4 (N1476, N1470, N489, N1059, N1082);
not NOT1 (N1477, N1475);
xor XOR2 (N1478, N1471, N387);
xor XOR2 (N1479, N1468, N781);
buf BUF1 (N1480, N1476);
buf BUF1 (N1481, N1479);
or OR4 (N1482, N1474, N925, N1076, N43);
or OR2 (N1483, N1472, N1316);
xor XOR2 (N1484, N1482, N291);
or OR4 (N1485, N1466, N1102, N1060, N384);
nand NAND3 (N1486, N1463, N1237, N1335);
not NOT1 (N1487, N1465);
xor XOR2 (N1488, N1477, N351);
nand NAND2 (N1489, N1481, N36);
nand NAND4 (N1490, N1484, N1058, N827, N249);
nand NAND3 (N1491, N1489, N73, N1355);
buf BUF1 (N1492, N1467);
nor NOR3 (N1493, N1478, N1270, N802);
nand NAND4 (N1494, N1488, N1421, N1268, N636);
xor XOR2 (N1495, N1486, N838);
buf BUF1 (N1496, N1494);
or OR4 (N1497, N1495, N219, N1017, N1495);
not NOT1 (N1498, N1492);
nor NOR4 (N1499, N1497, N1073, N1139, N114);
and AND4 (N1500, N1493, N640, N20, N1180);
not NOT1 (N1501, N1487);
and AND2 (N1502, N1483, N302);
or OR2 (N1503, N1502, N714);
buf BUF1 (N1504, N1499);
buf BUF1 (N1505, N1485);
or OR2 (N1506, N1490, N1054);
and AND4 (N1507, N1498, N1095, N111, N447);
or OR3 (N1508, N1504, N985, N1025);
nor NOR2 (N1509, N1496, N316);
buf BUF1 (N1510, N1501);
buf BUF1 (N1511, N1510);
not NOT1 (N1512, N1505);
not NOT1 (N1513, N1500);
buf BUF1 (N1514, N1503);
or OR3 (N1515, N1480, N362, N870);
buf BUF1 (N1516, N1515);
and AND3 (N1517, N1507, N1509, N1462);
nand NAND2 (N1518, N1257, N610);
and AND3 (N1519, N1512, N626, N194);
xor XOR2 (N1520, N1514, N335);
xor XOR2 (N1521, N1516, N890);
nand NAND4 (N1522, N1491, N875, N958, N200);
or OR2 (N1523, N1511, N292);
nor NOR4 (N1524, N1513, N520, N722, N5);
and AND3 (N1525, N1522, N293, N18);
not NOT1 (N1526, N1519);
nor NOR2 (N1527, N1521, N504);
not NOT1 (N1528, N1527);
not NOT1 (N1529, N1525);
xor XOR2 (N1530, N1517, N1259);
and AND4 (N1531, N1526, N32, N833, N439);
not NOT1 (N1532, N1508);
or OR4 (N1533, N1520, N313, N6, N502);
buf BUF1 (N1534, N1529);
nand NAND3 (N1535, N1524, N534, N293);
nand NAND4 (N1536, N1531, N152, N129, N575);
not NOT1 (N1537, N1518);
xor XOR2 (N1538, N1532, N602);
xor XOR2 (N1539, N1536, N103);
buf BUF1 (N1540, N1533);
nor NOR2 (N1541, N1523, N721);
not NOT1 (N1542, N1540);
not NOT1 (N1543, N1530);
xor XOR2 (N1544, N1535, N332);
buf BUF1 (N1545, N1539);
and AND2 (N1546, N1541, N288);
buf BUF1 (N1547, N1544);
and AND2 (N1548, N1545, N1420);
or OR3 (N1549, N1506, N1495, N377);
nor NOR4 (N1550, N1546, N1354, N1307, N261);
xor XOR2 (N1551, N1534, N1248);
or OR2 (N1552, N1548, N472);
nor NOR2 (N1553, N1549, N220);
xor XOR2 (N1554, N1542, N619);
xor XOR2 (N1555, N1543, N887);
and AND4 (N1556, N1554, N750, N718, N439);
nand NAND3 (N1557, N1528, N629, N236);
xor XOR2 (N1558, N1552, N1219);
nand NAND2 (N1559, N1555, N1134);
buf BUF1 (N1560, N1553);
buf BUF1 (N1561, N1551);
or OR3 (N1562, N1561, N1427, N825);
not NOT1 (N1563, N1556);
buf BUF1 (N1564, N1547);
or OR2 (N1565, N1557, N1201);
nand NAND4 (N1566, N1550, N398, N1006, N702);
buf BUF1 (N1567, N1565);
xor XOR2 (N1568, N1562, N577);
buf BUF1 (N1569, N1568);
or OR3 (N1570, N1559, N1051, N929);
and AND2 (N1571, N1560, N873);
xor XOR2 (N1572, N1564, N1342);
or OR2 (N1573, N1566, N1472);
buf BUF1 (N1574, N1558);
not NOT1 (N1575, N1569);
or OR3 (N1576, N1563, N920, N398);
and AND3 (N1577, N1538, N1543, N397);
or OR4 (N1578, N1574, N518, N1550, N404);
not NOT1 (N1579, N1578);
or OR3 (N1580, N1577, N537, N976);
nand NAND2 (N1581, N1567, N852);
or OR2 (N1582, N1571, N1231);
or OR4 (N1583, N1579, N1341, N1486, N1115);
and AND4 (N1584, N1573, N921, N1567, N985);
not NOT1 (N1585, N1576);
buf BUF1 (N1586, N1580);
and AND4 (N1587, N1581, N1353, N107, N585);
xor XOR2 (N1588, N1586, N1140);
not NOT1 (N1589, N1575);
xor XOR2 (N1590, N1589, N765);
nor NOR3 (N1591, N1588, N476, N305);
buf BUF1 (N1592, N1591);
xor XOR2 (N1593, N1585, N1269);
nor NOR3 (N1594, N1582, N483, N72);
or OR4 (N1595, N1590, N426, N768, N211);
xor XOR2 (N1596, N1572, N1466);
nand NAND2 (N1597, N1592, N221);
xor XOR2 (N1598, N1597, N1015);
nor NOR2 (N1599, N1537, N439);
not NOT1 (N1600, N1596);
not NOT1 (N1601, N1594);
nand NAND4 (N1602, N1600, N932, N783, N754);
nor NOR3 (N1603, N1595, N1197, N1126);
not NOT1 (N1604, N1599);
nand NAND4 (N1605, N1604, N221, N1217, N402);
not NOT1 (N1606, N1603);
nor NOR3 (N1607, N1587, N694, N191);
or OR2 (N1608, N1602, N462);
buf BUF1 (N1609, N1606);
nor NOR2 (N1610, N1601, N271);
buf BUF1 (N1611, N1609);
nor NOR2 (N1612, N1611, N112);
nor NOR4 (N1613, N1583, N1269, N1189, N421);
xor XOR2 (N1614, N1598, N580);
nor NOR4 (N1615, N1584, N563, N883, N1565);
and AND2 (N1616, N1605, N980);
or OR4 (N1617, N1593, N1262, N1234, N787);
and AND3 (N1618, N1614, N986, N729);
buf BUF1 (N1619, N1613);
buf BUF1 (N1620, N1607);
xor XOR2 (N1621, N1619, N880);
nand NAND4 (N1622, N1617, N311, N154, N777);
not NOT1 (N1623, N1615);
and AND4 (N1624, N1608, N1293, N218, N1228);
buf BUF1 (N1625, N1610);
not NOT1 (N1626, N1621);
nand NAND2 (N1627, N1620, N1565);
xor XOR2 (N1628, N1612, N1396);
nor NOR3 (N1629, N1625, N1514, N169);
buf BUF1 (N1630, N1618);
not NOT1 (N1631, N1630);
xor XOR2 (N1632, N1624, N1115);
xor XOR2 (N1633, N1622, N821);
xor XOR2 (N1634, N1628, N386);
and AND3 (N1635, N1570, N1521, N360);
or OR3 (N1636, N1629, N153, N802);
not NOT1 (N1637, N1634);
buf BUF1 (N1638, N1627);
and AND3 (N1639, N1637, N1490, N640);
nand NAND3 (N1640, N1616, N1615, N409);
not NOT1 (N1641, N1631);
or OR4 (N1642, N1623, N761, N415, N1293);
nor NOR2 (N1643, N1633, N35);
nor NOR3 (N1644, N1643, N71, N314);
nand NAND2 (N1645, N1644, N66);
xor XOR2 (N1646, N1635, N347);
and AND4 (N1647, N1636, N457, N1497, N1374);
nand NAND3 (N1648, N1647, N246, N1251);
buf BUF1 (N1649, N1639);
buf BUF1 (N1650, N1642);
not NOT1 (N1651, N1632);
and AND4 (N1652, N1648, N975, N1077, N945);
or OR4 (N1653, N1638, N1191, N166, N540);
xor XOR2 (N1654, N1653, N1053);
or OR4 (N1655, N1645, N357, N166, N1056);
xor XOR2 (N1656, N1651, N1643);
nand NAND2 (N1657, N1656, N302);
xor XOR2 (N1658, N1626, N21);
nand NAND2 (N1659, N1657, N802);
nand NAND3 (N1660, N1650, N822, N1292);
and AND2 (N1661, N1640, N148);
and AND4 (N1662, N1646, N663, N131, N568);
xor XOR2 (N1663, N1649, N893);
nor NOR2 (N1664, N1662, N1301);
nand NAND2 (N1665, N1663, N307);
or OR3 (N1666, N1659, N1166, N1052);
nor NOR2 (N1667, N1666, N48);
or OR4 (N1668, N1664, N172, N227, N1379);
and AND4 (N1669, N1641, N478, N1445, N289);
xor XOR2 (N1670, N1654, N601);
nand NAND3 (N1671, N1652, N936, N614);
or OR2 (N1672, N1671, N335);
buf BUF1 (N1673, N1658);
or OR4 (N1674, N1655, N721, N822, N132);
not NOT1 (N1675, N1668);
or OR3 (N1676, N1670, N259, N765);
and AND4 (N1677, N1669, N1390, N648, N67);
not NOT1 (N1678, N1672);
not NOT1 (N1679, N1667);
xor XOR2 (N1680, N1678, N1409);
not NOT1 (N1681, N1660);
nor NOR3 (N1682, N1665, N95, N175);
nand NAND3 (N1683, N1676, N1420, N1638);
nand NAND2 (N1684, N1674, N364);
nor NOR3 (N1685, N1683, N1282, N183);
xor XOR2 (N1686, N1681, N1530);
or OR4 (N1687, N1675, N222, N650, N1241);
nand NAND3 (N1688, N1677, N1125, N23);
nand NAND2 (N1689, N1682, N441);
nor NOR4 (N1690, N1673, N15, N616, N791);
and AND4 (N1691, N1687, N685, N921, N1030);
or OR3 (N1692, N1679, N1087, N473);
not NOT1 (N1693, N1680);
not NOT1 (N1694, N1693);
buf BUF1 (N1695, N1692);
nor NOR3 (N1696, N1689, N1547, N871);
and AND4 (N1697, N1690, N649, N931, N345);
nand NAND4 (N1698, N1691, N615, N280, N1489);
not NOT1 (N1699, N1695);
or OR3 (N1700, N1686, N1596, N1351);
or OR2 (N1701, N1661, N1665);
buf BUF1 (N1702, N1685);
buf BUF1 (N1703, N1700);
nor NOR4 (N1704, N1697, N671, N689, N28);
buf BUF1 (N1705, N1696);
xor XOR2 (N1706, N1698, N136);
not NOT1 (N1707, N1705);
or OR3 (N1708, N1706, N640, N711);
nand NAND2 (N1709, N1708, N1116);
not NOT1 (N1710, N1703);
or OR2 (N1711, N1707, N1380);
nand NAND4 (N1712, N1694, N871, N175, N1268);
xor XOR2 (N1713, N1684, N499);
not NOT1 (N1714, N1699);
nand NAND3 (N1715, N1701, N77, N185);
nand NAND4 (N1716, N1711, N395, N1635, N652);
xor XOR2 (N1717, N1715, N145);
and AND3 (N1718, N1714, N391, N1338);
not NOT1 (N1719, N1716);
xor XOR2 (N1720, N1713, N1563);
not NOT1 (N1721, N1688);
xor XOR2 (N1722, N1717, N1463);
and AND3 (N1723, N1721, N394, N46);
not NOT1 (N1724, N1720);
or OR2 (N1725, N1704, N127);
or OR2 (N1726, N1723, N482);
not NOT1 (N1727, N1718);
nor NOR2 (N1728, N1722, N1541);
nor NOR3 (N1729, N1712, N1175, N256);
or OR3 (N1730, N1729, N1108, N1252);
not NOT1 (N1731, N1710);
and AND2 (N1732, N1728, N646);
nand NAND3 (N1733, N1719, N1513, N907);
not NOT1 (N1734, N1725);
and AND4 (N1735, N1730, N169, N524, N1248);
or OR3 (N1736, N1727, N1646, N62);
buf BUF1 (N1737, N1734);
nor NOR3 (N1738, N1702, N777, N747);
nor NOR3 (N1739, N1731, N1018, N1170);
nor NOR2 (N1740, N1724, N519);
or OR3 (N1741, N1736, N1427, N928);
nand NAND3 (N1742, N1733, N254, N1364);
xor XOR2 (N1743, N1732, N94);
or OR2 (N1744, N1726, N1634);
nor NOR4 (N1745, N1735, N138, N1419, N156);
buf BUF1 (N1746, N1741);
xor XOR2 (N1747, N1738, N703);
buf BUF1 (N1748, N1709);
xor XOR2 (N1749, N1742, N224);
nand NAND3 (N1750, N1745, N722, N821);
and AND3 (N1751, N1750, N325, N1237);
nand NAND2 (N1752, N1751, N476);
nand NAND3 (N1753, N1737, N1076, N722);
not NOT1 (N1754, N1749);
not NOT1 (N1755, N1748);
and AND4 (N1756, N1743, N1088, N828, N728);
buf BUF1 (N1757, N1754);
xor XOR2 (N1758, N1756, N518);
and AND4 (N1759, N1758, N1398, N37, N893);
nor NOR3 (N1760, N1752, N343, N1548);
or OR4 (N1761, N1760, N1144, N1367, N671);
and AND2 (N1762, N1739, N506);
and AND4 (N1763, N1762, N99, N1463, N1701);
nand NAND4 (N1764, N1747, N1265, N988, N1050);
xor XOR2 (N1765, N1744, N879);
buf BUF1 (N1766, N1763);
xor XOR2 (N1767, N1740, N1747);
or OR3 (N1768, N1765, N1700, N697);
buf BUF1 (N1769, N1764);
nand NAND3 (N1770, N1761, N1443, N1420);
or OR2 (N1771, N1746, N1326);
buf BUF1 (N1772, N1757);
and AND2 (N1773, N1770, N1332);
or OR4 (N1774, N1769, N1759, N705, N1410);
nand NAND2 (N1775, N766, N684);
or OR3 (N1776, N1766, N409, N1440);
nand NAND4 (N1777, N1771, N1461, N1644, N69);
nand NAND3 (N1778, N1777, N364, N1606);
xor XOR2 (N1779, N1772, N116);
nand NAND3 (N1780, N1778, N1025, N1650);
nand NAND2 (N1781, N1753, N1118);
nand NAND2 (N1782, N1775, N349);
and AND2 (N1783, N1774, N1179);
buf BUF1 (N1784, N1776);
and AND3 (N1785, N1767, N1687, N1073);
or OR4 (N1786, N1768, N56, N68, N1708);
buf BUF1 (N1787, N1779);
xor XOR2 (N1788, N1785, N670);
nand NAND4 (N1789, N1783, N225, N341, N689);
not NOT1 (N1790, N1789);
xor XOR2 (N1791, N1782, N1703);
and AND4 (N1792, N1788, N1223, N52, N811);
nand NAND3 (N1793, N1755, N1264, N1039);
nor NOR3 (N1794, N1787, N285, N1146);
nand NAND3 (N1795, N1781, N494, N1773);
not NOT1 (N1796, N1589);
or OR4 (N1797, N1790, N1174, N1550, N912);
or OR3 (N1798, N1786, N623, N811);
or OR2 (N1799, N1792, N453);
xor XOR2 (N1800, N1796, N39);
nand NAND3 (N1801, N1784, N1786, N420);
and AND3 (N1802, N1799, N417, N644);
nand NAND4 (N1803, N1802, N1487, N428, N215);
nand NAND2 (N1804, N1800, N597);
nor NOR2 (N1805, N1795, N705);
and AND4 (N1806, N1798, N698, N1603, N662);
nor NOR2 (N1807, N1804, N35);
buf BUF1 (N1808, N1803);
or OR3 (N1809, N1793, N1245, N768);
not NOT1 (N1810, N1797);
buf BUF1 (N1811, N1809);
xor XOR2 (N1812, N1801, N482);
not NOT1 (N1813, N1780);
or OR4 (N1814, N1794, N1106, N795, N1335);
nand NAND2 (N1815, N1812, N1275);
not NOT1 (N1816, N1805);
xor XOR2 (N1817, N1815, N1242);
xor XOR2 (N1818, N1807, N963);
or OR2 (N1819, N1808, N1140);
buf BUF1 (N1820, N1806);
xor XOR2 (N1821, N1810, N719);
and AND4 (N1822, N1819, N1314, N1550, N1167);
not NOT1 (N1823, N1814);
buf BUF1 (N1824, N1811);
or OR4 (N1825, N1791, N1524, N831, N1331);
nor NOR4 (N1826, N1816, N1700, N1207, N49);
and AND2 (N1827, N1818, N671);
nand NAND3 (N1828, N1817, N158, N990);
xor XOR2 (N1829, N1821, N756);
not NOT1 (N1830, N1826);
nand NAND2 (N1831, N1830, N690);
not NOT1 (N1832, N1828);
nor NOR4 (N1833, N1822, N90, N65, N785);
nand NAND3 (N1834, N1813, N731, N307);
not NOT1 (N1835, N1833);
xor XOR2 (N1836, N1835, N1776);
nand NAND2 (N1837, N1832, N456);
not NOT1 (N1838, N1824);
and AND3 (N1839, N1820, N864, N518);
buf BUF1 (N1840, N1827);
nor NOR3 (N1841, N1838, N438, N1613);
nor NOR2 (N1842, N1834, N193);
and AND3 (N1843, N1831, N310, N988);
not NOT1 (N1844, N1825);
nor NOR4 (N1845, N1843, N79, N1329, N857);
nor NOR3 (N1846, N1844, N868, N1775);
and AND4 (N1847, N1837, N997, N1217, N1392);
nand NAND3 (N1848, N1823, N1644, N1737);
buf BUF1 (N1849, N1848);
buf BUF1 (N1850, N1840);
nand NAND2 (N1851, N1839, N244);
nor NOR2 (N1852, N1851, N316);
buf BUF1 (N1853, N1845);
nor NOR2 (N1854, N1836, N529);
nand NAND2 (N1855, N1847, N1613);
nor NOR2 (N1856, N1853, N27);
and AND2 (N1857, N1841, N347);
or OR4 (N1858, N1854, N746, N900, N764);
nor NOR3 (N1859, N1850, N1732, N435);
nand NAND3 (N1860, N1842, N574, N334);
not NOT1 (N1861, N1829);
or OR4 (N1862, N1860, N1124, N1216, N1722);
nor NOR2 (N1863, N1862, N1457);
buf BUF1 (N1864, N1846);
or OR3 (N1865, N1855, N1095, N1016);
nand NAND2 (N1866, N1856, N287);
and AND2 (N1867, N1866, N991);
not NOT1 (N1868, N1861);
and AND2 (N1869, N1852, N1650);
or OR4 (N1870, N1857, N1735, N1148, N1421);
buf BUF1 (N1871, N1869);
not NOT1 (N1872, N1858);
not NOT1 (N1873, N1868);
not NOT1 (N1874, N1870);
xor XOR2 (N1875, N1864, N1749);
and AND2 (N1876, N1873, N223);
nor NOR2 (N1877, N1871, N131);
or OR2 (N1878, N1867, N1876);
nand NAND2 (N1879, N939, N210);
nand NAND4 (N1880, N1879, N594, N1082, N1876);
nor NOR4 (N1881, N1849, N250, N1215, N70);
or OR4 (N1882, N1881, N1576, N1167, N840);
or OR2 (N1883, N1877, N66);
buf BUF1 (N1884, N1874);
buf BUF1 (N1885, N1880);
buf BUF1 (N1886, N1878);
or OR4 (N1887, N1884, N784, N703, N161);
xor XOR2 (N1888, N1887, N52);
buf BUF1 (N1889, N1859);
nor NOR3 (N1890, N1886, N909, N1505);
or OR4 (N1891, N1882, N85, N301, N1110);
xor XOR2 (N1892, N1891, N270);
xor XOR2 (N1893, N1875, N418);
xor XOR2 (N1894, N1890, N665);
xor XOR2 (N1895, N1883, N389);
nor NOR4 (N1896, N1865, N211, N348, N899);
not NOT1 (N1897, N1895);
buf BUF1 (N1898, N1889);
not NOT1 (N1899, N1896);
and AND2 (N1900, N1893, N1192);
or OR3 (N1901, N1872, N92, N456);
xor XOR2 (N1902, N1897, N209);
buf BUF1 (N1903, N1902);
buf BUF1 (N1904, N1885);
xor XOR2 (N1905, N1888, N451);
or OR3 (N1906, N1892, N636, N1056);
nor NOR3 (N1907, N1905, N1651, N79);
not NOT1 (N1908, N1899);
and AND4 (N1909, N1901, N385, N117, N1681);
and AND4 (N1910, N1907, N1008, N487, N206);
not NOT1 (N1911, N1900);
or OR3 (N1912, N1906, N1283, N1649);
nand NAND3 (N1913, N1903, N702, N1176);
buf BUF1 (N1914, N1911);
nand NAND3 (N1915, N1908, N1748, N1025);
and AND4 (N1916, N1894, N1907, N496, N1618);
or OR3 (N1917, N1898, N799, N615);
buf BUF1 (N1918, N1913);
buf BUF1 (N1919, N1916);
and AND4 (N1920, N1917, N1197, N1897, N46);
nand NAND4 (N1921, N1910, N1902, N763, N288);
nand NAND4 (N1922, N1909, N14, N66, N734);
and AND3 (N1923, N1922, N1211, N742);
nand NAND2 (N1924, N1919, N13);
nand NAND2 (N1925, N1904, N92);
buf BUF1 (N1926, N1914);
nand NAND4 (N1927, N1921, N531, N333, N793);
and AND2 (N1928, N1923, N940);
nor NOR4 (N1929, N1863, N1184, N1193, N908);
nor NOR4 (N1930, N1926, N680, N1915, N1454);
or OR2 (N1931, N1556, N21);
and AND2 (N1932, N1912, N1448);
buf BUF1 (N1933, N1920);
nand NAND2 (N1934, N1929, N760);
buf BUF1 (N1935, N1925);
and AND3 (N1936, N1918, N840, N816);
nor NOR3 (N1937, N1934, N266, N1367);
or OR2 (N1938, N1935, N884);
buf BUF1 (N1939, N1931);
buf BUF1 (N1940, N1924);
and AND4 (N1941, N1936, N1369, N1660, N631);
xor XOR2 (N1942, N1932, N759);
or OR2 (N1943, N1938, N602);
nor NOR3 (N1944, N1940, N516, N1613);
nor NOR3 (N1945, N1943, N1700, N573);
not NOT1 (N1946, N1939);
nand NAND3 (N1947, N1930, N1710, N1849);
buf BUF1 (N1948, N1933);
nand NAND3 (N1949, N1927, N1926, N1235);
nand NAND2 (N1950, N1941, N1568);
nor NOR3 (N1951, N1947, N371, N1419);
or OR3 (N1952, N1950, N1147, N624);
nor NOR2 (N1953, N1951, N497);
xor XOR2 (N1954, N1942, N1073);
nor NOR3 (N1955, N1948, N149, N482);
nand NAND3 (N1956, N1946, N1424, N1845);
buf BUF1 (N1957, N1955);
nor NOR3 (N1958, N1957, N1431, N619);
or OR3 (N1959, N1944, N1923, N1744);
nor NOR2 (N1960, N1959, N1239);
xor XOR2 (N1961, N1956, N1704);
or OR2 (N1962, N1954, N457);
nand NAND2 (N1963, N1953, N1592);
nor NOR3 (N1964, N1949, N1741, N178);
xor XOR2 (N1965, N1945, N750);
xor XOR2 (N1966, N1964, N607);
and AND4 (N1967, N1961, N1959, N1021, N1148);
xor XOR2 (N1968, N1960, N1546);
nor NOR2 (N1969, N1967, N462);
not NOT1 (N1970, N1969);
nor NOR3 (N1971, N1965, N248, N1416);
buf BUF1 (N1972, N1970);
and AND3 (N1973, N1962, N316, N1720);
xor XOR2 (N1974, N1958, N909);
xor XOR2 (N1975, N1972, N682);
and AND4 (N1976, N1974, N1623, N846, N1290);
nor NOR4 (N1977, N1968, N1860, N932, N1001);
nand NAND3 (N1978, N1971, N123, N49);
and AND2 (N1979, N1976, N506);
nand NAND2 (N1980, N1977, N1234);
and AND4 (N1981, N1980, N959, N26, N772);
not NOT1 (N1982, N1928);
not NOT1 (N1983, N1952);
buf BUF1 (N1984, N1975);
not NOT1 (N1985, N1984);
nand NAND2 (N1986, N1966, N89);
buf BUF1 (N1987, N1983);
not NOT1 (N1988, N1985);
nand NAND3 (N1989, N1979, N1522, N1314);
and AND4 (N1990, N1982, N1283, N460, N786);
nor NOR2 (N1991, N1937, N1827);
and AND2 (N1992, N1973, N947);
nand NAND2 (N1993, N1978, N1304);
buf BUF1 (N1994, N1989);
nand NAND3 (N1995, N1992, N411, N1052);
not NOT1 (N1996, N1963);
nand NAND4 (N1997, N1988, N60, N96, N1044);
buf BUF1 (N1998, N1993);
nor NOR3 (N1999, N1981, N1052, N1690);
xor XOR2 (N2000, N1995, N560);
not NOT1 (N2001, N1998);
buf BUF1 (N2002, N1990);
nor NOR3 (N2003, N1986, N262, N1985);
buf BUF1 (N2004, N1996);
and AND4 (N2005, N1991, N1870, N598, N275);
buf BUF1 (N2006, N1999);
nand NAND4 (N2007, N2005, N20, N1865, N488);
not NOT1 (N2008, N2004);
and AND2 (N2009, N2002, N1185);
nor NOR4 (N2010, N2008, N1798, N1102, N1312);
or OR4 (N2011, N2010, N1344, N872, N1331);
buf BUF1 (N2012, N2003);
buf BUF1 (N2013, N2007);
or OR3 (N2014, N2009, N1278, N1789);
xor XOR2 (N2015, N2014, N1928);
buf BUF1 (N2016, N1987);
not NOT1 (N2017, N2012);
and AND2 (N2018, N1997, N595);
buf BUF1 (N2019, N2006);
xor XOR2 (N2020, N1994, N1551);
nor NOR4 (N2021, N2000, N800, N527, N557);
xor XOR2 (N2022, N2018, N392);
xor XOR2 (N2023, N2022, N2021);
xor XOR2 (N2024, N1889, N910);
buf BUF1 (N2025, N2011);
or OR4 (N2026, N2019, N1137, N1496, N1067);
xor XOR2 (N2027, N2025, N1724);
not NOT1 (N2028, N2013);
not NOT1 (N2029, N2026);
and AND2 (N2030, N2028, N867);
buf BUF1 (N2031, N2027);
nor NOR3 (N2032, N2023, N1707, N361);
or OR4 (N2033, N2032, N145, N1565, N207);
nand NAND2 (N2034, N2017, N853);
not NOT1 (N2035, N2034);
buf BUF1 (N2036, N2030);
or OR3 (N2037, N2031, N1180, N1229);
nand NAND4 (N2038, N2029, N646, N944, N1479);
nand NAND4 (N2039, N2016, N632, N407, N1582);
nand NAND2 (N2040, N2037, N1818);
or OR2 (N2041, N2015, N1030);
nor NOR3 (N2042, N2038, N353, N816);
nand NAND3 (N2043, N2039, N220, N1507);
nand NAND2 (N2044, N2020, N882);
xor XOR2 (N2045, N2044, N107);
nor NOR2 (N2046, N2043, N1208);
and AND4 (N2047, N2036, N518, N1063, N799);
buf BUF1 (N2048, N2046);
nor NOR4 (N2049, N2048, N742, N1483, N1545);
xor XOR2 (N2050, N2045, N1867);
nand NAND2 (N2051, N2035, N269);
or OR4 (N2052, N2042, N134, N934, N1025);
xor XOR2 (N2053, N2001, N120);
and AND4 (N2054, N2053, N1181, N1278, N1904);
buf BUF1 (N2055, N2054);
xor XOR2 (N2056, N2047, N118);
nand NAND3 (N2057, N2055, N951, N666);
xor XOR2 (N2058, N2049, N1562);
not NOT1 (N2059, N2056);
nor NOR4 (N2060, N2057, N1457, N549, N687);
nor NOR2 (N2061, N2060, N1037);
xor XOR2 (N2062, N2059, N78);
nor NOR2 (N2063, N2050, N1112);
not NOT1 (N2064, N2041);
not NOT1 (N2065, N2033);
and AND3 (N2066, N2040, N112, N1946);
or OR3 (N2067, N2066, N1772, N330);
buf BUF1 (N2068, N2058);
or OR2 (N2069, N2067, N1899);
nand NAND3 (N2070, N2063, N86, N457);
not NOT1 (N2071, N2070);
nor NOR2 (N2072, N2062, N546);
not NOT1 (N2073, N2069);
nor NOR4 (N2074, N2065, N1944, N927, N248);
xor XOR2 (N2075, N2073, N1351);
and AND2 (N2076, N2024, N975);
or OR4 (N2077, N2068, N1283, N233, N954);
and AND3 (N2078, N2061, N679, N2029);
or OR4 (N2079, N2075, N873, N1564, N1437);
or OR4 (N2080, N2077, N1469, N289, N1086);
nor NOR3 (N2081, N2072, N809, N753);
buf BUF1 (N2082, N2052);
buf BUF1 (N2083, N2082);
and AND2 (N2084, N2080, N679);
buf BUF1 (N2085, N2051);
nor NOR3 (N2086, N2085, N805, N722);
not NOT1 (N2087, N2074);
and AND3 (N2088, N2084, N267, N65);
xor XOR2 (N2089, N2086, N1526);
and AND4 (N2090, N2089, N438, N881, N1502);
nand NAND4 (N2091, N2087, N1398, N1881, N487);
or OR3 (N2092, N2076, N1270, N746);
or OR3 (N2093, N2078, N781, N1115);
nand NAND4 (N2094, N2064, N374, N1568, N968);
nor NOR4 (N2095, N2090, N1861, N1566, N327);
or OR2 (N2096, N2083, N1652);
not NOT1 (N2097, N2088);
xor XOR2 (N2098, N2097, N788);
xor XOR2 (N2099, N2079, N365);
nand NAND2 (N2100, N2091, N1301);
and AND2 (N2101, N2071, N1456);
buf BUF1 (N2102, N2093);
buf BUF1 (N2103, N2095);
or OR4 (N2104, N2092, N197, N1845, N842);
nor NOR4 (N2105, N2094, N1345, N1208, N1662);
or OR4 (N2106, N2100, N1369, N1672, N1399);
buf BUF1 (N2107, N2081);
buf BUF1 (N2108, N2105);
buf BUF1 (N2109, N2106);
nand NAND3 (N2110, N2099, N1637, N1728);
nand NAND2 (N2111, N2109, N1658);
not NOT1 (N2112, N2096);
nor NOR2 (N2113, N2110, N1370);
xor XOR2 (N2114, N2108, N1177);
nor NOR2 (N2115, N2098, N1712);
not NOT1 (N2116, N2111);
or OR3 (N2117, N2102, N1135, N1219);
nor NOR3 (N2118, N2101, N1592, N628);
or OR2 (N2119, N2118, N1845);
not NOT1 (N2120, N2117);
nor NOR4 (N2121, N2120, N696, N928, N1005);
and AND4 (N2122, N2104, N1992, N734, N1979);
xor XOR2 (N2123, N2115, N1671);
not NOT1 (N2124, N2103);
nor NOR4 (N2125, N2113, N1553, N559, N933);
nor NOR2 (N2126, N2122, N1902);
xor XOR2 (N2127, N2124, N1197);
or OR3 (N2128, N2112, N1890, N563);
buf BUF1 (N2129, N2114);
nor NOR4 (N2130, N2116, N1162, N1575, N883);
and AND2 (N2131, N2107, N836);
xor XOR2 (N2132, N2121, N300);
nand NAND3 (N2133, N2125, N1045, N343);
nand NAND3 (N2134, N2130, N609, N2129);
buf BUF1 (N2135, N1369);
buf BUF1 (N2136, N2127);
not NOT1 (N2137, N2135);
nand NAND3 (N2138, N2134, N864, N1787);
or OR4 (N2139, N2132, N236, N502, N916);
nand NAND2 (N2140, N2133, N854);
not NOT1 (N2141, N2138);
nand NAND2 (N2142, N2119, N1511);
and AND4 (N2143, N2141, N1475, N707, N519);
or OR2 (N2144, N2136, N361);
and AND4 (N2145, N2142, N7, N2087, N153);
nand NAND3 (N2146, N2137, N1795, N744);
or OR4 (N2147, N2145, N261, N1793, N866);
or OR4 (N2148, N2139, N646, N1250, N1200);
and AND2 (N2149, N2123, N881);
or OR3 (N2150, N2128, N1542, N684);
buf BUF1 (N2151, N2148);
not NOT1 (N2152, N2147);
or OR4 (N2153, N2152, N1829, N875, N68);
nor NOR4 (N2154, N2149, N2112, N1332, N1150);
nor NOR3 (N2155, N2151, N2130, N1976);
nand NAND3 (N2156, N2143, N378, N751);
or OR4 (N2157, N2140, N151, N222, N1225);
not NOT1 (N2158, N2157);
buf BUF1 (N2159, N2150);
nand NAND2 (N2160, N2154, N1122);
not NOT1 (N2161, N2158);
nand NAND4 (N2162, N2161, N1667, N1978, N1905);
buf BUF1 (N2163, N2153);
and AND2 (N2164, N2126, N319);
xor XOR2 (N2165, N2144, N477);
nand NAND3 (N2166, N2159, N1266, N1673);
and AND2 (N2167, N2163, N900);
buf BUF1 (N2168, N2162);
not NOT1 (N2169, N2168);
and AND3 (N2170, N2155, N1362, N1931);
buf BUF1 (N2171, N2169);
and AND2 (N2172, N2165, N148);
nand NAND3 (N2173, N2171, N626, N1064);
nor NOR2 (N2174, N2166, N569);
xor XOR2 (N2175, N2174, N834);
not NOT1 (N2176, N2131);
nor NOR2 (N2177, N2156, N353);
and AND2 (N2178, N2160, N666);
nand NAND4 (N2179, N2172, N1073, N485, N808);
buf BUF1 (N2180, N2175);
and AND4 (N2181, N2177, N1149, N1426, N734);
and AND2 (N2182, N2146, N65);
buf BUF1 (N2183, N2182);
nor NOR2 (N2184, N2181, N914);
xor XOR2 (N2185, N2173, N1872);
or OR3 (N2186, N2179, N800, N1214);
buf BUF1 (N2187, N2186);
nand NAND2 (N2188, N2185, N1308);
not NOT1 (N2189, N2178);
and AND2 (N2190, N2176, N1515);
buf BUF1 (N2191, N2190);
nand NAND2 (N2192, N2180, N1617);
or OR3 (N2193, N2183, N722, N5);
not NOT1 (N2194, N2189);
buf BUF1 (N2195, N2167);
buf BUF1 (N2196, N2193);
nand NAND3 (N2197, N2170, N1716, N564);
nor NOR4 (N2198, N2188, N1207, N1321, N2152);
xor XOR2 (N2199, N2198, N1194);
buf BUF1 (N2200, N2187);
and AND4 (N2201, N2197, N1341, N224, N1366);
buf BUF1 (N2202, N2184);
xor XOR2 (N2203, N2195, N1461);
and AND3 (N2204, N2196, N568, N1391);
xor XOR2 (N2205, N2194, N2034);
or OR2 (N2206, N2203, N777);
xor XOR2 (N2207, N2202, N1087);
nand NAND2 (N2208, N2191, N821);
not NOT1 (N2209, N2199);
and AND4 (N2210, N2192, N1426, N1010, N1174);
or OR2 (N2211, N2204, N880);
not NOT1 (N2212, N2164);
buf BUF1 (N2213, N2209);
nand NAND4 (N2214, N2211, N1553, N1092, N1320);
not NOT1 (N2215, N2206);
not NOT1 (N2216, N2212);
nand NAND3 (N2217, N2216, N839, N2011);
nand NAND4 (N2218, N2208, N636, N429, N2207);
buf BUF1 (N2219, N2117);
nand NAND4 (N2220, N2210, N1478, N672, N361);
or OR3 (N2221, N2213, N1534, N1192);
buf BUF1 (N2222, N2215);
or OR4 (N2223, N2221, N1672, N118, N740);
buf BUF1 (N2224, N2201);
and AND3 (N2225, N2224, N566, N641);
nand NAND2 (N2226, N2223, N1304);
or OR2 (N2227, N2220, N982);
not NOT1 (N2228, N2218);
not NOT1 (N2229, N2200);
not NOT1 (N2230, N2219);
and AND3 (N2231, N2226, N588, N1012);
not NOT1 (N2232, N2214);
nand NAND3 (N2233, N2225, N1241, N583);
or OR2 (N2234, N2228, N1827);
not NOT1 (N2235, N2231);
nand NAND4 (N2236, N2234, N2071, N2204, N1762);
or OR2 (N2237, N2205, N1577);
not NOT1 (N2238, N2235);
or OR4 (N2239, N2232, N1570, N679, N705);
not NOT1 (N2240, N2217);
buf BUF1 (N2241, N2237);
or OR4 (N2242, N2227, N1189, N1369, N906);
and AND2 (N2243, N2229, N421);
or OR3 (N2244, N2230, N498, N681);
or OR4 (N2245, N2238, N334, N144, N145);
xor XOR2 (N2246, N2241, N1757);
or OR3 (N2247, N2246, N1802, N1656);
nor NOR4 (N2248, N2244, N1311, N713, N1474);
xor XOR2 (N2249, N2239, N1172);
not NOT1 (N2250, N2248);
and AND3 (N2251, N2233, N1954, N1657);
and AND4 (N2252, N2247, N1990, N663, N438);
xor XOR2 (N2253, N2249, N1687);
xor XOR2 (N2254, N2245, N1051);
nand NAND4 (N2255, N2240, N1647, N522, N1553);
or OR4 (N2256, N2253, N1918, N438, N711);
or OR3 (N2257, N2252, N833, N1);
xor XOR2 (N2258, N2222, N1292);
buf BUF1 (N2259, N2242);
nand NAND4 (N2260, N2256, N1985, N44, N1739);
or OR4 (N2261, N2236, N1123, N1422, N1185);
or OR4 (N2262, N2243, N996, N2072, N2169);
not NOT1 (N2263, N2255);
nand NAND2 (N2264, N2250, N2132);
or OR2 (N2265, N2257, N1730);
buf BUF1 (N2266, N2263);
not NOT1 (N2267, N2258);
buf BUF1 (N2268, N2264);
xor XOR2 (N2269, N2260, N736);
or OR2 (N2270, N2261, N1502);
or OR4 (N2271, N2266, N1557, N2201, N39);
nand NAND2 (N2272, N2259, N1280);
or OR2 (N2273, N2268, N2055);
buf BUF1 (N2274, N2271);
xor XOR2 (N2275, N2274, N520);
nor NOR2 (N2276, N2273, N1977);
nor NOR4 (N2277, N2251, N1587, N1728, N2045);
nor NOR4 (N2278, N2270, N1799, N15, N1390);
buf BUF1 (N2279, N2262);
not NOT1 (N2280, N2272);
and AND2 (N2281, N2265, N2040);
nand NAND3 (N2282, N2277, N1752, N2132);
not NOT1 (N2283, N2267);
or OR4 (N2284, N2282, N2068, N1544, N880);
or OR4 (N2285, N2279, N30, N930, N2190);
xor XOR2 (N2286, N2280, N1934);
not NOT1 (N2287, N2283);
nor NOR2 (N2288, N2284, N148);
buf BUF1 (N2289, N2288);
buf BUF1 (N2290, N2269);
or OR3 (N2291, N2276, N1433, N2070);
buf BUF1 (N2292, N2285);
nor NOR3 (N2293, N2287, N2242, N1405);
nor NOR2 (N2294, N2289, N2092);
not NOT1 (N2295, N2281);
and AND2 (N2296, N2254, N28);
and AND3 (N2297, N2278, N460, N2107);
and AND3 (N2298, N2290, N1759, N2024);
buf BUF1 (N2299, N2293);
not NOT1 (N2300, N2286);
buf BUF1 (N2301, N2294);
nand NAND2 (N2302, N2298, N2163);
buf BUF1 (N2303, N2275);
nand NAND2 (N2304, N2303, N485);
not NOT1 (N2305, N2291);
and AND3 (N2306, N2297, N846, N1048);
and AND2 (N2307, N2296, N87);
nor NOR4 (N2308, N2301, N1310, N2140, N956);
nand NAND3 (N2309, N2292, N1530, N2257);
nand NAND3 (N2310, N2304, N364, N2041);
nor NOR4 (N2311, N2306, N54, N460, N2101);
buf BUF1 (N2312, N2310);
xor XOR2 (N2313, N2312, N1153);
not NOT1 (N2314, N2309);
nor NOR4 (N2315, N2313, N1208, N238, N287);
not NOT1 (N2316, N2299);
buf BUF1 (N2317, N2316);
not NOT1 (N2318, N2305);
nand NAND2 (N2319, N2302, N2299);
not NOT1 (N2320, N2307);
not NOT1 (N2321, N2315);
nand NAND4 (N2322, N2318, N966, N2181, N408);
buf BUF1 (N2323, N2321);
xor XOR2 (N2324, N2323, N1294);
xor XOR2 (N2325, N2314, N1897);
nand NAND4 (N2326, N2325, N395, N384, N1139);
xor XOR2 (N2327, N2311, N929);
xor XOR2 (N2328, N2295, N596);
and AND2 (N2329, N2326, N195);
xor XOR2 (N2330, N2300, N1602);
nand NAND3 (N2331, N2308, N1872, N474);
buf BUF1 (N2332, N2319);
xor XOR2 (N2333, N2331, N1349);
buf BUF1 (N2334, N2330);
xor XOR2 (N2335, N2329, N1707);
buf BUF1 (N2336, N2327);
buf BUF1 (N2337, N2333);
and AND3 (N2338, N2322, N2267, N915);
nor NOR2 (N2339, N2335, N2109);
and AND2 (N2340, N2334, N1120);
xor XOR2 (N2341, N2336, N476);
not NOT1 (N2342, N2324);
nand NAND2 (N2343, N2339, N516);
buf BUF1 (N2344, N2317);
or OR3 (N2345, N2338, N2313, N690);
or OR4 (N2346, N2332, N792, N1401, N419);
not NOT1 (N2347, N2340);
xor XOR2 (N2348, N2337, N400);
xor XOR2 (N2349, N2346, N2341);
or OR4 (N2350, N535, N1930, N2245, N634);
and AND4 (N2351, N2348, N743, N225, N2085);
buf BUF1 (N2352, N2343);
xor XOR2 (N2353, N2345, N229);
nand NAND2 (N2354, N2349, N1874);
xor XOR2 (N2355, N2344, N934);
or OR4 (N2356, N2347, N1199, N856, N1874);
nand NAND2 (N2357, N2320, N137);
buf BUF1 (N2358, N2357);
nor NOR2 (N2359, N2358, N1751);
xor XOR2 (N2360, N2353, N1042);
or OR3 (N2361, N2351, N1812, N2112);
not NOT1 (N2362, N2356);
buf BUF1 (N2363, N2355);
not NOT1 (N2364, N2360);
buf BUF1 (N2365, N2362);
buf BUF1 (N2366, N2364);
nand NAND4 (N2367, N2350, N1518, N2208, N1272);
or OR3 (N2368, N2342, N2076, N49);
nand NAND2 (N2369, N2363, N3);
and AND2 (N2370, N2366, N235);
xor XOR2 (N2371, N2368, N2327);
nand NAND2 (N2372, N2365, N1972);
buf BUF1 (N2373, N2354);
buf BUF1 (N2374, N2373);
and AND4 (N2375, N2372, N650, N1560, N2109);
and AND4 (N2376, N2374, N365, N1981, N927);
or OR2 (N2377, N2370, N279);
xor XOR2 (N2378, N2371, N808);
nor NOR4 (N2379, N2369, N308, N1160, N436);
or OR3 (N2380, N2328, N17, N376);
nand NAND3 (N2381, N2378, N1417, N2180);
and AND2 (N2382, N2377, N2213);
or OR2 (N2383, N2361, N2131);
nor NOR2 (N2384, N2352, N90);
or OR4 (N2385, N2379, N1776, N2164, N1291);
nand NAND2 (N2386, N2367, N1998);
nand NAND2 (N2387, N2359, N1214);
or OR3 (N2388, N2383, N387, N2072);
buf BUF1 (N2389, N2375);
nor NOR4 (N2390, N2385, N1579, N2025, N2011);
xor XOR2 (N2391, N2386, N2278);
buf BUF1 (N2392, N2387);
or OR3 (N2393, N2381, N165, N1813);
buf BUF1 (N2394, N2390);
nand NAND4 (N2395, N2392, N1141, N1555, N818);
nand NAND4 (N2396, N2382, N117, N1677, N1206);
xor XOR2 (N2397, N2395, N2113);
nand NAND4 (N2398, N2397, N672, N248, N1776);
xor XOR2 (N2399, N2396, N2278);
nand NAND3 (N2400, N2391, N39, N1343);
nand NAND4 (N2401, N2393, N2196, N2044, N566);
buf BUF1 (N2402, N2389);
nand NAND4 (N2403, N2380, N593, N1104, N1723);
nand NAND3 (N2404, N2399, N2302, N1103);
or OR4 (N2405, N2404, N2254, N1882, N251);
nor NOR3 (N2406, N2401, N199, N1136);
or OR3 (N2407, N2400, N1468, N2394);
or OR2 (N2408, N589, N457);
nand NAND3 (N2409, N2407, N1008, N1173);
and AND3 (N2410, N2376, N287, N585);
buf BUF1 (N2411, N2410);
nor NOR2 (N2412, N2406, N385);
or OR2 (N2413, N2403, N2269);
nand NAND4 (N2414, N2409, N392, N733, N1767);
and AND4 (N2415, N2411, N252, N893, N1528);
or OR2 (N2416, N2413, N647);
nor NOR2 (N2417, N2412, N2188);
or OR2 (N2418, N2398, N1229);
and AND3 (N2419, N2384, N292, N1674);
or OR3 (N2420, N2405, N1745, N1198);
not NOT1 (N2421, N2415);
nor NOR3 (N2422, N2421, N1272, N1733);
xor XOR2 (N2423, N2402, N1295);
nand NAND4 (N2424, N2414, N110, N1011, N1874);
not NOT1 (N2425, N2418);
nor NOR3 (N2426, N2419, N863, N1945);
xor XOR2 (N2427, N2426, N1665);
xor XOR2 (N2428, N2420, N445);
or OR2 (N2429, N2417, N1524);
xor XOR2 (N2430, N2427, N699);
xor XOR2 (N2431, N2416, N17);
nor NOR2 (N2432, N2424, N552);
and AND2 (N2433, N2429, N2049);
xor XOR2 (N2434, N2432, N1378);
not NOT1 (N2435, N2434);
nor NOR3 (N2436, N2433, N1321, N1180);
buf BUF1 (N2437, N2422);
or OR2 (N2438, N2425, N1231);
and AND4 (N2439, N2436, N761, N99, N211);
buf BUF1 (N2440, N2423);
nor NOR4 (N2441, N2439, N389, N2363, N1595);
and AND3 (N2442, N2440, N1000, N1805);
nor NOR2 (N2443, N2435, N864);
not NOT1 (N2444, N2408);
or OR4 (N2445, N2428, N1010, N1393, N747);
and AND2 (N2446, N2388, N2075);
buf BUF1 (N2447, N2430);
or OR4 (N2448, N2446, N347, N1359, N896);
not NOT1 (N2449, N2447);
xor XOR2 (N2450, N2441, N1108);
or OR2 (N2451, N2449, N2253);
not NOT1 (N2452, N2431);
buf BUF1 (N2453, N2450);
and AND3 (N2454, N2438, N1420, N20);
and AND2 (N2455, N2452, N1219);
or OR3 (N2456, N2443, N843, N1753);
buf BUF1 (N2457, N2437);
buf BUF1 (N2458, N2442);
nor NOR4 (N2459, N2457, N269, N2168, N876);
nor NOR3 (N2460, N2455, N138, N610);
xor XOR2 (N2461, N2445, N578);
not NOT1 (N2462, N2460);
buf BUF1 (N2463, N2458);
not NOT1 (N2464, N2451);
xor XOR2 (N2465, N2459, N1258);
nand NAND3 (N2466, N2454, N2017, N1090);
or OR3 (N2467, N2463, N2212, N1789);
not NOT1 (N2468, N2465);
and AND3 (N2469, N2448, N1324, N334);
nand NAND2 (N2470, N2466, N885);
and AND4 (N2471, N2464, N79, N621, N1100);
and AND3 (N2472, N2471, N134, N633);
buf BUF1 (N2473, N2456);
not NOT1 (N2474, N2461);
nand NAND2 (N2475, N2453, N1107);
xor XOR2 (N2476, N2472, N1899);
nor NOR3 (N2477, N2462, N9, N1984);
not NOT1 (N2478, N2477);
and AND3 (N2479, N2476, N2392, N158);
xor XOR2 (N2480, N2475, N1334);
nor NOR2 (N2481, N2469, N614);
not NOT1 (N2482, N2467);
xor XOR2 (N2483, N2473, N861);
not NOT1 (N2484, N2481);
buf BUF1 (N2485, N2470);
and AND2 (N2486, N2483, N1249);
buf BUF1 (N2487, N2478);
nor NOR2 (N2488, N2484, N207);
xor XOR2 (N2489, N2474, N222);
buf BUF1 (N2490, N2485);
or OR4 (N2491, N2486, N790, N343, N423);
nand NAND3 (N2492, N2480, N722, N1404);
or OR4 (N2493, N2482, N1082, N1716, N2017);
nor NOR4 (N2494, N2468, N2274, N1723, N884);
nand NAND3 (N2495, N2493, N756, N983);
nand NAND3 (N2496, N2479, N2071, N535);
or OR2 (N2497, N2492, N499);
xor XOR2 (N2498, N2490, N1385);
buf BUF1 (N2499, N2444);
nor NOR4 (N2500, N2487, N110, N957, N838);
xor XOR2 (N2501, N2489, N1638);
or OR4 (N2502, N2499, N112, N2248, N1402);
nor NOR2 (N2503, N2502, N1662);
or OR3 (N2504, N2491, N860, N1817);
and AND4 (N2505, N2504, N2132, N832, N1726);
nor NOR4 (N2506, N2497, N1117, N1041, N2292);
or OR2 (N2507, N2500, N628);
not NOT1 (N2508, N2507);
buf BUF1 (N2509, N2496);
xor XOR2 (N2510, N2495, N2038);
and AND4 (N2511, N2505, N112, N967, N1106);
nand NAND4 (N2512, N2509, N1873, N715, N361);
not NOT1 (N2513, N2501);
not NOT1 (N2514, N2513);
and AND3 (N2515, N2506, N450, N1811);
or OR3 (N2516, N2511, N954, N1905);
not NOT1 (N2517, N2514);
nor NOR3 (N2518, N2494, N1676, N1064);
xor XOR2 (N2519, N2516, N1493);
and AND2 (N2520, N2517, N1850);
nand NAND4 (N2521, N2512, N1702, N414, N1861);
xor XOR2 (N2522, N2488, N2478);
and AND4 (N2523, N2519, N1539, N1220, N92);
xor XOR2 (N2524, N2521, N1769);
nand NAND3 (N2525, N2508, N897, N1125);
nor NOR4 (N2526, N2520, N450, N946, N2344);
buf BUF1 (N2527, N2518);
buf BUF1 (N2528, N2527);
nor NOR4 (N2529, N2515, N1487, N2170, N1728);
and AND4 (N2530, N2528, N265, N721, N842);
not NOT1 (N2531, N2526);
not NOT1 (N2532, N2523);
xor XOR2 (N2533, N2531, N2187);
nor NOR2 (N2534, N2503, N1391);
and AND3 (N2535, N2525, N824, N987);
or OR4 (N2536, N2535, N1475, N1298, N147);
and AND3 (N2537, N2534, N948, N252);
buf BUF1 (N2538, N2533);
not NOT1 (N2539, N2530);
not NOT1 (N2540, N2538);
nand NAND2 (N2541, N2529, N1409);
buf BUF1 (N2542, N2510);
xor XOR2 (N2543, N2539, N2275);
not NOT1 (N2544, N2536);
or OR4 (N2545, N2542, N1664, N384, N2125);
and AND4 (N2546, N2545, N526, N2313, N1441);
nor NOR3 (N2547, N2522, N814, N2241);
xor XOR2 (N2548, N2544, N2230);
and AND2 (N2549, N2543, N1400);
buf BUF1 (N2550, N2540);
and AND3 (N2551, N2498, N2146, N2206);
and AND4 (N2552, N2546, N1731, N2253, N1351);
or OR2 (N2553, N2551, N104);
buf BUF1 (N2554, N2547);
and AND2 (N2555, N2532, N582);
nor NOR2 (N2556, N2524, N1898);
and AND3 (N2557, N2537, N1749, N1835);
nor NOR3 (N2558, N2553, N232, N1971);
nor NOR2 (N2559, N2550, N2177);
nand NAND3 (N2560, N2549, N844, N1962);
nand NAND3 (N2561, N2548, N2429, N39);
or OR3 (N2562, N2557, N2007, N1959);
and AND4 (N2563, N2541, N2013, N2239, N1699);
xor XOR2 (N2564, N2563, N57);
nand NAND4 (N2565, N2559, N2388, N1570, N291);
not NOT1 (N2566, N2555);
not NOT1 (N2567, N2558);
nor NOR4 (N2568, N2567, N728, N1697, N924);
nand NAND4 (N2569, N2552, N764, N1070, N994);
and AND2 (N2570, N2561, N1332);
not NOT1 (N2571, N2570);
xor XOR2 (N2572, N2556, N1945);
nor NOR3 (N2573, N2560, N1666, N2421);
or OR4 (N2574, N2566, N589, N1987, N196);
nor NOR3 (N2575, N2574, N1427, N1556);
nor NOR3 (N2576, N2564, N133, N2029);
not NOT1 (N2577, N2576);
buf BUF1 (N2578, N2569);
nor NOR4 (N2579, N2572, N114, N921, N234);
nor NOR3 (N2580, N2577, N1978, N2076);
and AND4 (N2581, N2571, N2477, N634, N687);
or OR2 (N2582, N2565, N1084);
not NOT1 (N2583, N2582);
buf BUF1 (N2584, N2579);
nor NOR4 (N2585, N2578, N1365, N350, N1113);
xor XOR2 (N2586, N2585, N1650);
nor NOR2 (N2587, N2581, N1912);
not NOT1 (N2588, N2573);
nand NAND3 (N2589, N2554, N1639, N1203);
xor XOR2 (N2590, N2580, N525);
and AND3 (N2591, N2583, N2039, N2372);
xor XOR2 (N2592, N2587, N1518);
buf BUF1 (N2593, N2562);
buf BUF1 (N2594, N2589);
buf BUF1 (N2595, N2594);
and AND4 (N2596, N2590, N2388, N1580, N1001);
and AND2 (N2597, N2588, N1606);
buf BUF1 (N2598, N2597);
nor NOR4 (N2599, N2595, N249, N2534, N891);
buf BUF1 (N2600, N2575);
or OR3 (N2601, N2591, N93, N1769);
or OR4 (N2602, N2599, N429, N792, N1673);
and AND4 (N2603, N2592, N656, N368, N1422);
buf BUF1 (N2604, N2601);
nor NOR3 (N2605, N2593, N1607, N1654);
buf BUF1 (N2606, N2584);
nor NOR4 (N2607, N2603, N757, N2272, N640);
and AND4 (N2608, N2596, N2290, N654, N1356);
and AND2 (N2609, N2598, N1572);
or OR4 (N2610, N2607, N1303, N1318, N2220);
nand NAND3 (N2611, N2568, N695, N1703);
xor XOR2 (N2612, N2609, N1702);
nand NAND2 (N2613, N2608, N2367);
and AND2 (N2614, N2600, N1865);
or OR4 (N2615, N2605, N2534, N1260, N2367);
nor NOR2 (N2616, N2602, N1124);
xor XOR2 (N2617, N2616, N874);
nor NOR2 (N2618, N2615, N950);
and AND4 (N2619, N2618, N2321, N2345, N612);
xor XOR2 (N2620, N2604, N1355);
nand NAND2 (N2621, N2613, N2323);
nand NAND4 (N2622, N2610, N2153, N2057, N640);
and AND4 (N2623, N2619, N1532, N1537, N1047);
buf BUF1 (N2624, N2586);
and AND3 (N2625, N2623, N1061, N194);
not NOT1 (N2626, N2624);
nor NOR2 (N2627, N2626, N1707);
nor NOR2 (N2628, N2617, N1660);
nand NAND4 (N2629, N2606, N1668, N2159, N1756);
nand NAND4 (N2630, N2621, N1242, N1540, N1233);
xor XOR2 (N2631, N2627, N1031);
nand NAND2 (N2632, N2625, N872);
and AND4 (N2633, N2612, N676, N689, N2390);
nor NOR4 (N2634, N2611, N751, N1970, N2002);
nor NOR3 (N2635, N2630, N1039, N2342);
not NOT1 (N2636, N2631);
buf BUF1 (N2637, N2629);
not NOT1 (N2638, N2634);
or OR3 (N2639, N2622, N317, N2219);
or OR3 (N2640, N2636, N683, N1932);
or OR3 (N2641, N2628, N671, N1858);
nor NOR3 (N2642, N2635, N1140, N209);
and AND3 (N2643, N2639, N1804, N675);
not NOT1 (N2644, N2642);
nand NAND3 (N2645, N2632, N2405, N1750);
and AND3 (N2646, N2640, N121, N45);
not NOT1 (N2647, N2633);
xor XOR2 (N2648, N2638, N1954);
nand NAND4 (N2649, N2646, N941, N505, N120);
buf BUF1 (N2650, N2649);
xor XOR2 (N2651, N2644, N781);
xor XOR2 (N2652, N2650, N1874);
buf BUF1 (N2653, N2648);
and AND3 (N2654, N2653, N2301, N2201);
and AND4 (N2655, N2645, N2236, N1779, N715);
not NOT1 (N2656, N2620);
xor XOR2 (N2657, N2614, N582);
xor XOR2 (N2658, N2657, N2469);
buf BUF1 (N2659, N2655);
nand NAND3 (N2660, N2652, N1332, N887);
buf BUF1 (N2661, N2654);
and AND2 (N2662, N2656, N1812);
xor XOR2 (N2663, N2643, N2262);
or OR4 (N2664, N2651, N1562, N959, N980);
nor NOR4 (N2665, N2658, N396, N2593, N256);
nor NOR4 (N2666, N2659, N1568, N2201, N1224);
or OR2 (N2667, N2665, N2317);
nand NAND3 (N2668, N2661, N1563, N2140);
nand NAND4 (N2669, N2660, N1422, N1895, N753);
or OR2 (N2670, N2663, N2436);
nand NAND2 (N2671, N2670, N2032);
nand NAND2 (N2672, N2668, N2534);
xor XOR2 (N2673, N2672, N855);
and AND2 (N2674, N2664, N2186);
or OR4 (N2675, N2641, N1487, N1638, N2472);
or OR4 (N2676, N2674, N2123, N1955, N2029);
and AND2 (N2677, N2662, N1926);
and AND4 (N2678, N2673, N1341, N2346, N1462);
not NOT1 (N2679, N2677);
xor XOR2 (N2680, N2679, N1673);
buf BUF1 (N2681, N2680);
buf BUF1 (N2682, N2666);
nor NOR2 (N2683, N2682, N404);
and AND2 (N2684, N2681, N1621);
nor NOR3 (N2685, N2676, N29, N747);
xor XOR2 (N2686, N2678, N1485);
or OR2 (N2687, N2683, N173);
or OR2 (N2688, N2684, N2418);
xor XOR2 (N2689, N2669, N2499);
nand NAND2 (N2690, N2685, N1830);
not NOT1 (N2691, N2687);
buf BUF1 (N2692, N2691);
and AND3 (N2693, N2689, N593, N2263);
nand NAND2 (N2694, N2667, N1399);
or OR3 (N2695, N2694, N1843, N1186);
nand NAND4 (N2696, N2686, N1496, N1791, N1836);
not NOT1 (N2697, N2671);
nand NAND3 (N2698, N2693, N1646, N106);
nand NAND2 (N2699, N2697, N1111);
and AND3 (N2700, N2699, N2451, N2330);
buf BUF1 (N2701, N2637);
buf BUF1 (N2702, N2701);
buf BUF1 (N2703, N2675);
buf BUF1 (N2704, N2703);
xor XOR2 (N2705, N2692, N984);
and AND4 (N2706, N2698, N1223, N905, N1349);
nor NOR3 (N2707, N2688, N496, N157);
nand NAND2 (N2708, N2696, N2226);
xor XOR2 (N2709, N2695, N1925);
buf BUF1 (N2710, N2706);
and AND3 (N2711, N2705, N2055, N2531);
buf BUF1 (N2712, N2647);
xor XOR2 (N2713, N2707, N207);
nor NOR2 (N2714, N2713, N1626);
or OR4 (N2715, N2710, N1859, N2168, N1728);
nor NOR2 (N2716, N2702, N2598);
xor XOR2 (N2717, N2700, N1504);
xor XOR2 (N2718, N2704, N1661);
buf BUF1 (N2719, N2709);
buf BUF1 (N2720, N2708);
nand NAND2 (N2721, N2718, N1585);
nor NOR2 (N2722, N2721, N2150);
or OR3 (N2723, N2711, N1586, N1266);
xor XOR2 (N2724, N2714, N1933);
xor XOR2 (N2725, N2690, N604);
not NOT1 (N2726, N2724);
nand NAND4 (N2727, N2723, N991, N667, N1727);
and AND4 (N2728, N2720, N1895, N637, N2105);
xor XOR2 (N2729, N2722, N2468);
nor NOR2 (N2730, N2717, N1549);
or OR2 (N2731, N2729, N1956);
nor NOR4 (N2732, N2726, N198, N1424, N1893);
or OR3 (N2733, N2719, N919, N1447);
xor XOR2 (N2734, N2712, N881);
nand NAND2 (N2735, N2732, N2043);
not NOT1 (N2736, N2725);
nand NAND2 (N2737, N2716, N2048);
xor XOR2 (N2738, N2730, N517);
not NOT1 (N2739, N2738);
nand NAND4 (N2740, N2734, N51, N2330, N604);
or OR2 (N2741, N2731, N37);
not NOT1 (N2742, N2735);
not NOT1 (N2743, N2742);
buf BUF1 (N2744, N2739);
nand NAND3 (N2745, N2727, N2248, N1130);
not NOT1 (N2746, N2715);
nand NAND4 (N2747, N2745, N2104, N1257, N2556);
nor NOR4 (N2748, N2744, N832, N1641, N2517);
buf BUF1 (N2749, N2733);
xor XOR2 (N2750, N2743, N1549);
or OR4 (N2751, N2748, N2637, N2289, N2610);
nor NOR3 (N2752, N2750, N2561, N785);
or OR4 (N2753, N2751, N1523, N1849, N1543);
or OR4 (N2754, N2736, N1525, N2717, N775);
buf BUF1 (N2755, N2737);
nor NOR4 (N2756, N2749, N1711, N2732, N901);
not NOT1 (N2757, N2740);
xor XOR2 (N2758, N2746, N1548);
not NOT1 (N2759, N2747);
or OR2 (N2760, N2728, N185);
nor NOR2 (N2761, N2755, N2580);
or OR3 (N2762, N2758, N110, N1200);
or OR4 (N2763, N2760, N676, N1596, N1159);
or OR4 (N2764, N2759, N1640, N1670, N2254);
or OR4 (N2765, N2754, N214, N808, N1687);
buf BUF1 (N2766, N2762);
not NOT1 (N2767, N2763);
nor NOR4 (N2768, N2767, N2381, N739, N2431);
not NOT1 (N2769, N2761);
and AND2 (N2770, N2766, N1526);
nand NAND3 (N2771, N2756, N1868, N2231);
not NOT1 (N2772, N2753);
nor NOR3 (N2773, N2769, N2277, N2233);
xor XOR2 (N2774, N2773, N1073);
xor XOR2 (N2775, N2752, N2149);
buf BUF1 (N2776, N2771);
nand NAND4 (N2777, N2774, N739, N938, N490);
and AND3 (N2778, N2757, N88, N454);
and AND4 (N2779, N2776, N2671, N332, N161);
nand NAND2 (N2780, N2741, N1218);
buf BUF1 (N2781, N2764);
nor NOR2 (N2782, N2775, N165);
and AND3 (N2783, N2778, N2571, N890);
not NOT1 (N2784, N2782);
nand NAND3 (N2785, N2783, N179, N1790);
or OR4 (N2786, N2772, N2715, N834, N1710);
or OR4 (N2787, N2785, N1675, N2781, N2003);
nand NAND2 (N2788, N797, N2305);
or OR3 (N2789, N2765, N1723, N352);
nor NOR4 (N2790, N2784, N1771, N76, N1424);
xor XOR2 (N2791, N2786, N728);
and AND4 (N2792, N2791, N849, N1966, N199);
or OR2 (N2793, N2789, N2347);
buf BUF1 (N2794, N2779);
and AND3 (N2795, N2793, N1940, N863);
nor NOR4 (N2796, N2787, N841, N81, N2379);
or OR3 (N2797, N2792, N1567, N1692);
xor XOR2 (N2798, N2796, N574);
nand NAND4 (N2799, N2790, N2437, N80, N2701);
not NOT1 (N2800, N2795);
buf BUF1 (N2801, N2768);
or OR4 (N2802, N2797, N35, N2351, N1797);
nor NOR4 (N2803, N2801, N978, N2714, N88);
or OR2 (N2804, N2780, N1830);
buf BUF1 (N2805, N2788);
or OR2 (N2806, N2803, N2161);
xor XOR2 (N2807, N2800, N2026);
nand NAND2 (N2808, N2802, N128);
not NOT1 (N2809, N2794);
and AND2 (N2810, N2804, N1738);
or OR3 (N2811, N2805, N89, N2309);
not NOT1 (N2812, N2770);
or OR3 (N2813, N2812, N2384, N772);
or OR4 (N2814, N2808, N2559, N1124, N148);
not NOT1 (N2815, N2807);
and AND2 (N2816, N2809, N844);
or OR2 (N2817, N2813, N1766);
nand NAND4 (N2818, N2777, N2760, N288, N495);
nand NAND4 (N2819, N2814, N2221, N1649, N2428);
xor XOR2 (N2820, N2811, N1433);
or OR2 (N2821, N2818, N513);
or OR2 (N2822, N2806, N1562);
nand NAND3 (N2823, N2816, N2372, N2781);
nand NAND4 (N2824, N2810, N2614, N1778, N2806);
not NOT1 (N2825, N2821);
not NOT1 (N2826, N2824);
nor NOR3 (N2827, N2799, N2129, N665);
nor NOR3 (N2828, N2817, N2239, N1092);
nand NAND4 (N2829, N2828, N2495, N2244, N2551);
and AND4 (N2830, N2822, N2028, N2139, N1705);
nand NAND3 (N2831, N2815, N2212, N1781);
buf BUF1 (N2832, N2820);
or OR4 (N2833, N2832, N1907, N612, N125);
nand NAND3 (N2834, N2831, N1417, N1058);
and AND4 (N2835, N2825, N286, N1836, N1132);
and AND4 (N2836, N2829, N440, N653, N2661);
not NOT1 (N2837, N2833);
nor NOR3 (N2838, N2798, N1424, N535);
nand NAND3 (N2839, N2837, N2013, N541);
nand NAND2 (N2840, N2823, N1547);
buf BUF1 (N2841, N2819);
buf BUF1 (N2842, N2836);
nor NOR2 (N2843, N2841, N2517);
nor NOR3 (N2844, N2834, N1429, N335);
not NOT1 (N2845, N2839);
nor NOR3 (N2846, N2843, N361, N1946);
nand NAND3 (N2847, N2840, N471, N1441);
and AND2 (N2848, N2826, N2567);
buf BUF1 (N2849, N2848);
and AND4 (N2850, N2835, N264, N434, N468);
and AND4 (N2851, N2842, N1366, N272, N2069);
buf BUF1 (N2852, N2845);
nand NAND4 (N2853, N2827, N1257, N1274, N1246);
xor XOR2 (N2854, N2849, N1754);
and AND4 (N2855, N2846, N2196, N702, N419);
nor NOR3 (N2856, N2853, N2110, N1161);
or OR3 (N2857, N2847, N201, N1562);
or OR2 (N2858, N2851, N939);
buf BUF1 (N2859, N2855);
buf BUF1 (N2860, N2856);
xor XOR2 (N2861, N2844, N2756);
and AND2 (N2862, N2861, N1178);
buf BUF1 (N2863, N2862);
nand NAND4 (N2864, N2858, N1826, N2136, N439);
xor XOR2 (N2865, N2854, N832);
or OR3 (N2866, N2863, N2371, N2535);
and AND2 (N2867, N2866, N376);
and AND4 (N2868, N2859, N591, N1126, N2250);
nor NOR2 (N2869, N2864, N1705);
and AND4 (N2870, N2865, N1396, N1429, N1163);
and AND3 (N2871, N2838, N1414, N975);
xor XOR2 (N2872, N2868, N2666);
xor XOR2 (N2873, N2869, N846);
and AND4 (N2874, N2872, N2474, N540, N1939);
buf BUF1 (N2875, N2870);
or OR4 (N2876, N2850, N1479, N327, N1355);
buf BUF1 (N2877, N2830);
nor NOR3 (N2878, N2860, N1635, N2204);
nor NOR3 (N2879, N2874, N1896, N1847);
xor XOR2 (N2880, N2876, N767);
not NOT1 (N2881, N2871);
xor XOR2 (N2882, N2881, N2825);
nand NAND3 (N2883, N2867, N21, N622);
nor NOR4 (N2884, N2879, N1784, N1372, N946);
and AND4 (N2885, N2857, N2821, N1805, N43);
nor NOR2 (N2886, N2883, N530);
or OR4 (N2887, N2884, N522, N393, N1641);
nand NAND4 (N2888, N2886, N362, N401, N1925);
nand NAND4 (N2889, N2873, N439, N235, N497);
nand NAND4 (N2890, N2875, N391, N1701, N2164);
nand NAND2 (N2891, N2890, N1946);
nand NAND3 (N2892, N2852, N1974, N1092);
nand NAND3 (N2893, N2888, N2706, N2324);
not NOT1 (N2894, N2887);
nor NOR3 (N2895, N2885, N1237, N2079);
nand NAND3 (N2896, N2889, N2469, N1626);
and AND2 (N2897, N2892, N2686);
buf BUF1 (N2898, N2877);
nand NAND2 (N2899, N2898, N378);
or OR3 (N2900, N2895, N2623, N2876);
and AND4 (N2901, N2899, N374, N2263, N2787);
buf BUF1 (N2902, N2880);
not NOT1 (N2903, N2894);
and AND4 (N2904, N2901, N2747, N337, N2043);
not NOT1 (N2905, N2893);
xor XOR2 (N2906, N2903, N2531);
or OR3 (N2907, N2896, N2458, N2311);
not NOT1 (N2908, N2900);
and AND4 (N2909, N2907, N217, N1592, N2335);
and AND3 (N2910, N2904, N1078, N1943);
xor XOR2 (N2911, N2908, N1860);
xor XOR2 (N2912, N2878, N2889);
xor XOR2 (N2913, N2910, N21);
and AND2 (N2914, N2902, N1868);
buf BUF1 (N2915, N2909);
not NOT1 (N2916, N2914);
nand NAND3 (N2917, N2891, N2297, N1864);
or OR2 (N2918, N2882, N1007);
not NOT1 (N2919, N2916);
xor XOR2 (N2920, N2905, N1295);
nor NOR4 (N2921, N2917, N2501, N2377, N447);
buf BUF1 (N2922, N2906);
nor NOR3 (N2923, N2921, N362, N649);
or OR3 (N2924, N2915, N2428, N454);
nor NOR4 (N2925, N2912, N296, N2506, N1837);
and AND3 (N2926, N2911, N2179, N1090);
and AND3 (N2927, N2924, N2371, N813);
and AND2 (N2928, N2927, N1135);
nand NAND4 (N2929, N2926, N1323, N1786, N1990);
nor NOR3 (N2930, N2897, N1003, N2644);
or OR3 (N2931, N2928, N487, N2515);
or OR3 (N2932, N2931, N1168, N1644);
nor NOR4 (N2933, N2932, N437, N2363, N1208);
xor XOR2 (N2934, N2925, N2758);
buf BUF1 (N2935, N2920);
not NOT1 (N2936, N2929);
and AND3 (N2937, N2933, N2881, N1169);
or OR4 (N2938, N2937, N293, N803, N1860);
not NOT1 (N2939, N2923);
and AND4 (N2940, N2936, N1204, N127, N1509);
nor NOR4 (N2941, N2930, N502, N2283, N2343);
buf BUF1 (N2942, N2919);
nand NAND3 (N2943, N2941, N2874, N1983);
nor NOR2 (N2944, N2940, N526);
xor XOR2 (N2945, N2913, N1476);
xor XOR2 (N2946, N2939, N2043);
and AND2 (N2947, N2945, N1593);
nor NOR4 (N2948, N2942, N2003, N2733, N569);
or OR4 (N2949, N2935, N1099, N2947, N628);
buf BUF1 (N2950, N1147);
xor XOR2 (N2951, N2944, N2025);
buf BUF1 (N2952, N2922);
nor NOR2 (N2953, N2943, N2702);
or OR3 (N2954, N2946, N1624, N2633);
nor NOR3 (N2955, N2938, N393, N1772);
not NOT1 (N2956, N2934);
nor NOR4 (N2957, N2955, N818, N459, N2181);
and AND3 (N2958, N2951, N1288, N2481);
buf BUF1 (N2959, N2953);
nor NOR2 (N2960, N2948, N2166);
buf BUF1 (N2961, N2952);
nand NAND3 (N2962, N2959, N1177, N1710);
not NOT1 (N2963, N2956);
nand NAND3 (N2964, N2963, N224, N1140);
and AND2 (N2965, N2962, N368);
nor NOR2 (N2966, N2950, N2505);
not NOT1 (N2967, N2949);
nand NAND2 (N2968, N2965, N1736);
and AND3 (N2969, N2918, N1985, N2200);
buf BUF1 (N2970, N2967);
xor XOR2 (N2971, N2969, N2750);
and AND3 (N2972, N2957, N2602, N108);
or OR4 (N2973, N2961, N2426, N1618, N882);
buf BUF1 (N2974, N2968);
nand NAND3 (N2975, N2966, N906, N1963);
nor NOR3 (N2976, N2974, N1016, N1469);
xor XOR2 (N2977, N2958, N2366);
nor NOR2 (N2978, N2964, N2909);
nor NOR4 (N2979, N2954, N750, N2274, N2165);
buf BUF1 (N2980, N2960);
or OR3 (N2981, N2978, N486, N963);
not NOT1 (N2982, N2981);
buf BUF1 (N2983, N2971);
nand NAND2 (N2984, N2972, N1572);
and AND4 (N2985, N2982, N2762, N2477, N403);
and AND2 (N2986, N2983, N2900);
buf BUF1 (N2987, N2980);
and AND4 (N2988, N2975, N1486, N1609, N1753);
not NOT1 (N2989, N2985);
xor XOR2 (N2990, N2988, N1882);
buf BUF1 (N2991, N2979);
xor XOR2 (N2992, N2986, N2921);
and AND2 (N2993, N2970, N1031);
nor NOR3 (N2994, N2987, N1246, N2136);
xor XOR2 (N2995, N2984, N130);
nor NOR3 (N2996, N2990, N2322, N1007);
nand NAND2 (N2997, N2977, N1001);
buf BUF1 (N2998, N2989);
nand NAND2 (N2999, N2991, N483);
nand NAND3 (N3000, N2994, N2904, N1026);
nor NOR3 (N3001, N2997, N1833, N2771);
xor XOR2 (N3002, N2976, N513);
xor XOR2 (N3003, N2996, N656);
not NOT1 (N3004, N3000);
or OR3 (N3005, N3001, N918, N1187);
and AND2 (N3006, N3002, N664);
nor NOR4 (N3007, N2995, N2754, N631, N2899);
and AND3 (N3008, N2973, N1548, N2542);
nand NAND4 (N3009, N3005, N1169, N1502, N803);
and AND4 (N3010, N3006, N66, N539, N124);
buf BUF1 (N3011, N3003);
and AND2 (N3012, N3008, N2546);
or OR3 (N3013, N2992, N790, N76);
nor NOR4 (N3014, N2999, N143, N1210, N2181);
and AND2 (N3015, N3011, N1289);
not NOT1 (N3016, N3014);
xor XOR2 (N3017, N3016, N747);
and AND4 (N3018, N3009, N770, N452, N282);
nor NOR4 (N3019, N3015, N1672, N254, N1380);
nor NOR4 (N3020, N2998, N2204, N2069, N843);
xor XOR2 (N3021, N2993, N2905);
and AND4 (N3022, N3020, N2871, N2686, N399);
and AND2 (N3023, N3004, N760);
buf BUF1 (N3024, N3022);
buf BUF1 (N3025, N3021);
nor NOR2 (N3026, N3024, N1563);
nor NOR3 (N3027, N3018, N813, N891);
or OR2 (N3028, N3017, N1494);
xor XOR2 (N3029, N3007, N203);
not NOT1 (N3030, N3029);
nor NOR3 (N3031, N3030, N1238, N1805);
and AND2 (N3032, N3023, N1235);
nand NAND2 (N3033, N3013, N904);
xor XOR2 (N3034, N3025, N131);
buf BUF1 (N3035, N3027);
nor NOR4 (N3036, N3032, N1725, N2599, N1209);
buf BUF1 (N3037, N3012);
not NOT1 (N3038, N3031);
or OR4 (N3039, N3033, N1860, N1551, N393);
or OR3 (N3040, N3028, N672, N922);
and AND3 (N3041, N3010, N2723, N2856);
xor XOR2 (N3042, N3036, N480);
and AND2 (N3043, N3042, N2821);
buf BUF1 (N3044, N3019);
and AND2 (N3045, N3026, N2933);
nor NOR3 (N3046, N3045, N3015, N2604);
buf BUF1 (N3047, N3039);
nor NOR4 (N3048, N3035, N2132, N577, N61);
nand NAND4 (N3049, N3038, N2889, N106, N2949);
buf BUF1 (N3050, N3048);
nor NOR4 (N3051, N3044, N170, N1295, N1897);
nand NAND3 (N3052, N3034, N3027, N1082);
or OR4 (N3053, N3051, N943, N2323, N2056);
nand NAND2 (N3054, N3043, N2275);
xor XOR2 (N3055, N3046, N1954);
buf BUF1 (N3056, N3047);
nor NOR2 (N3057, N3052, N2243);
buf BUF1 (N3058, N3050);
or OR3 (N3059, N3041, N1452, N1052);
nand NAND2 (N3060, N3040, N38);
xor XOR2 (N3061, N3058, N466);
and AND3 (N3062, N3054, N27, N2271);
and AND3 (N3063, N3056, N2801, N1851);
not NOT1 (N3064, N3060);
xor XOR2 (N3065, N3053, N2527);
nor NOR4 (N3066, N3049, N13, N367, N1094);
nand NAND2 (N3067, N3055, N1943);
nand NAND4 (N3068, N3062, N4, N219, N3010);
and AND3 (N3069, N3057, N997, N1236);
not NOT1 (N3070, N3037);
buf BUF1 (N3071, N3066);
xor XOR2 (N3072, N3063, N2303);
nor NOR2 (N3073, N3068, N528);
or OR3 (N3074, N3071, N2437, N564);
nor NOR2 (N3075, N3069, N502);
nand NAND4 (N3076, N3059, N532, N2727, N1177);
buf BUF1 (N3077, N3073);
or OR2 (N3078, N3067, N1328);
nor NOR2 (N3079, N3078, N491);
buf BUF1 (N3080, N3079);
nor NOR2 (N3081, N3075, N1789);
buf BUF1 (N3082, N3077);
or OR4 (N3083, N3076, N2201, N1783, N2437);
or OR2 (N3084, N3072, N140);
not NOT1 (N3085, N3083);
nor NOR2 (N3086, N3065, N2658);
nor NOR4 (N3087, N3074, N2687, N1885, N2841);
not NOT1 (N3088, N3084);
or OR2 (N3089, N3086, N870);
xor XOR2 (N3090, N3080, N1630);
or OR4 (N3091, N3085, N2811, N1354, N979);
or OR3 (N3092, N3061, N801, N334);
xor XOR2 (N3093, N3089, N509);
xor XOR2 (N3094, N3092, N2548);
and AND4 (N3095, N3082, N1495, N675, N985);
not NOT1 (N3096, N3064);
nor NOR4 (N3097, N3093, N146, N870, N1701);
xor XOR2 (N3098, N3091, N622);
nand NAND2 (N3099, N3081, N2366);
nand NAND2 (N3100, N3098, N1228);
and AND2 (N3101, N3096, N786);
not NOT1 (N3102, N3099);
buf BUF1 (N3103, N3087);
not NOT1 (N3104, N3088);
xor XOR2 (N3105, N3104, N2464);
xor XOR2 (N3106, N3090, N1469);
buf BUF1 (N3107, N3101);
nand NAND2 (N3108, N3094, N810);
nor NOR4 (N3109, N3095, N1398, N2323, N2611);
xor XOR2 (N3110, N3105, N1733);
not NOT1 (N3111, N3106);
buf BUF1 (N3112, N3070);
nand NAND3 (N3113, N3111, N1394, N907);
nor NOR4 (N3114, N3097, N778, N601, N2005);
nor NOR4 (N3115, N3102, N1146, N562, N1486);
not NOT1 (N3116, N3103);
and AND4 (N3117, N3108, N2864, N2703, N678);
not NOT1 (N3118, N3117);
not NOT1 (N3119, N3100);
buf BUF1 (N3120, N3112);
nand NAND3 (N3121, N3110, N1155, N2907);
buf BUF1 (N3122, N3115);
nor NOR2 (N3123, N3120, N870);
not NOT1 (N3124, N3118);
not NOT1 (N3125, N3116);
not NOT1 (N3126, N3114);
or OR2 (N3127, N3124, N1846);
buf BUF1 (N3128, N3122);
buf BUF1 (N3129, N3127);
not NOT1 (N3130, N3123);
or OR2 (N3131, N3125, N1652);
xor XOR2 (N3132, N3131, N506);
or OR3 (N3133, N3109, N129, N889);
nor NOR4 (N3134, N3133, N422, N705, N2039);
xor XOR2 (N3135, N3126, N1460);
xor XOR2 (N3136, N3113, N1921);
buf BUF1 (N3137, N3119);
not NOT1 (N3138, N3107);
or OR4 (N3139, N3137, N1102, N2131, N113);
and AND3 (N3140, N3121, N1738, N1073);
nand NAND2 (N3141, N3129, N1528);
buf BUF1 (N3142, N3135);
buf BUF1 (N3143, N3128);
not NOT1 (N3144, N3143);
nand NAND3 (N3145, N3136, N553, N1468);
and AND4 (N3146, N3138, N3138, N3014, N870);
nor NOR3 (N3147, N3141, N2905, N2208);
xor XOR2 (N3148, N3140, N989);
not NOT1 (N3149, N3130);
and AND4 (N3150, N3144, N2856, N2553, N206);
not NOT1 (N3151, N3147);
and AND4 (N3152, N3146, N2549, N1861, N2906);
not NOT1 (N3153, N3152);
xor XOR2 (N3154, N3145, N2187);
and AND3 (N3155, N3132, N734, N3120);
and AND2 (N3156, N3148, N1150);
nand NAND3 (N3157, N3156, N1994, N2624);
nor NOR3 (N3158, N3151, N2827, N997);
or OR2 (N3159, N3153, N1835);
or OR2 (N3160, N3154, N703);
and AND2 (N3161, N3157, N2400);
not NOT1 (N3162, N3155);
xor XOR2 (N3163, N3159, N50);
nor NOR2 (N3164, N3162, N340);
xor XOR2 (N3165, N3164, N1168);
not NOT1 (N3166, N3150);
nand NAND3 (N3167, N3139, N2961, N133);
or OR3 (N3168, N3167, N2412, N284);
and AND2 (N3169, N3166, N1622);
not NOT1 (N3170, N3161);
nor NOR2 (N3171, N3165, N835);
buf BUF1 (N3172, N3168);
not NOT1 (N3173, N3134);
nand NAND2 (N3174, N3171, N2055);
and AND2 (N3175, N3163, N1524);
buf BUF1 (N3176, N3170);
buf BUF1 (N3177, N3175);
or OR2 (N3178, N3172, N2911);
not NOT1 (N3179, N3158);
nand NAND4 (N3180, N3177, N1156, N1017, N1686);
xor XOR2 (N3181, N3180, N2104);
nand NAND2 (N3182, N3176, N1569);
nand NAND3 (N3183, N3169, N890, N2800);
xor XOR2 (N3184, N3183, N1518);
nor NOR4 (N3185, N3182, N2405, N1530, N1049);
not NOT1 (N3186, N3179);
and AND3 (N3187, N3142, N1968, N1191);
or OR4 (N3188, N3174, N2474, N2588, N2022);
xor XOR2 (N3189, N3187, N1802);
and AND4 (N3190, N3184, N380, N1882, N1561);
or OR3 (N3191, N3178, N2381, N2297);
nor NOR3 (N3192, N3181, N2583, N3034);
not NOT1 (N3193, N3190);
nand NAND3 (N3194, N3189, N2634, N875);
nand NAND2 (N3195, N3193, N434);
nand NAND3 (N3196, N3191, N1488, N466);
or OR3 (N3197, N3195, N7, N2082);
xor XOR2 (N3198, N3192, N2901);
buf BUF1 (N3199, N3173);
not NOT1 (N3200, N3199);
and AND3 (N3201, N3197, N2265, N2707);
or OR3 (N3202, N3196, N147, N2912);
not NOT1 (N3203, N3194);
and AND3 (N3204, N3200, N551, N104);
nor NOR4 (N3205, N3186, N3016, N663, N742);
xor XOR2 (N3206, N3149, N1822);
nand NAND4 (N3207, N3160, N676, N287, N1955);
or OR2 (N3208, N3185, N162);
not NOT1 (N3209, N3198);
xor XOR2 (N3210, N3205, N1984);
and AND4 (N3211, N3204, N1950, N1342, N3035);
not NOT1 (N3212, N3208);
buf BUF1 (N3213, N3210);
xor XOR2 (N3214, N3202, N2590);
not NOT1 (N3215, N3203);
xor XOR2 (N3216, N3215, N556);
nand NAND2 (N3217, N3201, N2197);
nand NAND2 (N3218, N3217, N1462);
buf BUF1 (N3219, N3213);
xor XOR2 (N3220, N3214, N1736);
and AND2 (N3221, N3206, N2270);
nor NOR3 (N3222, N3211, N2083, N2019);
nor NOR3 (N3223, N3209, N1954, N2029);
buf BUF1 (N3224, N3219);
buf BUF1 (N3225, N3223);
and AND4 (N3226, N3221, N1166, N2770, N2325);
nand NAND3 (N3227, N3224, N2149, N1954);
nor NOR4 (N3228, N3220, N878, N2559, N257);
not NOT1 (N3229, N3222);
nor NOR2 (N3230, N3229, N1202);
or OR4 (N3231, N3207, N2703, N3052, N2375);
buf BUF1 (N3232, N3218);
and AND2 (N3233, N3232, N282);
buf BUF1 (N3234, N3188);
nand NAND4 (N3235, N3230, N3095, N637, N2661);
nand NAND4 (N3236, N3231, N2883, N1303, N686);
xor XOR2 (N3237, N3233, N3078);
buf BUF1 (N3238, N3237);
nand NAND2 (N3239, N3227, N260);
buf BUF1 (N3240, N3235);
xor XOR2 (N3241, N3240, N639);
nand NAND3 (N3242, N3225, N1835, N2212);
xor XOR2 (N3243, N3238, N2757);
buf BUF1 (N3244, N3212);
nor NOR4 (N3245, N3226, N2680, N1170, N2181);
buf BUF1 (N3246, N3243);
nand NAND4 (N3247, N3246, N2291, N1106, N1637);
nor NOR4 (N3248, N3236, N1353, N3106, N1562);
or OR2 (N3249, N3247, N2416);
or OR3 (N3250, N3244, N1238, N1357);
or OR3 (N3251, N3228, N2670, N699);
xor XOR2 (N3252, N3239, N2706);
nand NAND4 (N3253, N3248, N954, N2198, N2341);
nand NAND2 (N3254, N3216, N1607);
or OR3 (N3255, N3242, N828, N2053);
nor NOR4 (N3256, N3249, N39, N2702, N2785);
nor NOR2 (N3257, N3253, N2018);
xor XOR2 (N3258, N3256, N2256);
xor XOR2 (N3259, N3254, N288);
nand NAND4 (N3260, N3251, N2228, N2376, N1992);
xor XOR2 (N3261, N3234, N838);
buf BUF1 (N3262, N3255);
not NOT1 (N3263, N3258);
buf BUF1 (N3264, N3252);
nand NAND2 (N3265, N3263, N3142);
and AND3 (N3266, N3250, N1255, N2638);
or OR2 (N3267, N3261, N1611);
and AND3 (N3268, N3259, N1441, N3025);
buf BUF1 (N3269, N3241);
nor NOR4 (N3270, N3260, N349, N794, N1877);
nand NAND2 (N3271, N3267, N3032);
not NOT1 (N3272, N3264);
buf BUF1 (N3273, N3245);
nand NAND4 (N3274, N3268, N2534, N1439, N3077);
nor NOR2 (N3275, N3269, N1988);
xor XOR2 (N3276, N3273, N103);
xor XOR2 (N3277, N3265, N1618);
buf BUF1 (N3278, N3271);
buf BUF1 (N3279, N3270);
and AND2 (N3280, N3279, N1661);
xor XOR2 (N3281, N3262, N3142);
nor NOR3 (N3282, N3275, N3002, N387);
nand NAND4 (N3283, N3278, N2725, N2520, N2093);
nand NAND2 (N3284, N3276, N2360);
nor NOR4 (N3285, N3272, N1467, N1609, N1788);
nand NAND4 (N3286, N3280, N2774, N321, N1968);
nor NOR4 (N3287, N3283, N1390, N1760, N2621);
buf BUF1 (N3288, N3281);
buf BUF1 (N3289, N3257);
xor XOR2 (N3290, N3287, N697);
or OR2 (N3291, N3289, N3193);
not NOT1 (N3292, N3274);
nand NAND3 (N3293, N3277, N1867, N48);
nor NOR4 (N3294, N3290, N2593, N2727, N2012);
xor XOR2 (N3295, N3294, N47);
nor NOR2 (N3296, N3266, N480);
or OR4 (N3297, N3288, N3198, N1965, N2799);
not NOT1 (N3298, N3292);
buf BUF1 (N3299, N3298);
buf BUF1 (N3300, N3297);
or OR3 (N3301, N3284, N1064, N710);
xor XOR2 (N3302, N3299, N589);
nor NOR2 (N3303, N3286, N823);
nand NAND2 (N3304, N3300, N521);
nand NAND4 (N3305, N3291, N2857, N1059, N3052);
nor NOR3 (N3306, N3301, N319, N3028);
nor NOR2 (N3307, N3296, N1508);
and AND3 (N3308, N3305, N1571, N2461);
and AND2 (N3309, N3308, N2778);
nand NAND2 (N3310, N3307, N545);
not NOT1 (N3311, N3303);
xor XOR2 (N3312, N3285, N2083);
and AND4 (N3313, N3311, N533, N2849, N1827);
or OR2 (N3314, N3306, N198);
nand NAND4 (N3315, N3304, N2342, N2046, N1473);
and AND4 (N3316, N3282, N3056, N1032, N2347);
or OR4 (N3317, N3312, N902, N179, N2438);
and AND3 (N3318, N3315, N1215, N415);
nand NAND4 (N3319, N3293, N1500, N1395, N1878);
nor NOR3 (N3320, N3319, N439, N3289);
xor XOR2 (N3321, N3302, N2668);
buf BUF1 (N3322, N3318);
buf BUF1 (N3323, N3320);
nand NAND2 (N3324, N3309, N2981);
xor XOR2 (N3325, N3317, N809);
xor XOR2 (N3326, N3314, N853);
or OR4 (N3327, N3313, N1420, N2636, N396);
or OR2 (N3328, N3323, N1353);
not NOT1 (N3329, N3324);
not NOT1 (N3330, N3325);
nand NAND2 (N3331, N3328, N2234);
nor NOR4 (N3332, N3295, N367, N1941, N61);
buf BUF1 (N3333, N3322);
and AND3 (N3334, N3310, N2454, N1753);
xor XOR2 (N3335, N3329, N3243);
not NOT1 (N3336, N3316);
or OR2 (N3337, N3326, N3151);
xor XOR2 (N3338, N3332, N1539);
or OR2 (N3339, N3333, N1731);
nor NOR2 (N3340, N3334, N3317);
not NOT1 (N3341, N3340);
nand NAND3 (N3342, N3331, N1329, N961);
xor XOR2 (N3343, N3341, N2211);
buf BUF1 (N3344, N3338);
xor XOR2 (N3345, N3327, N1082);
not NOT1 (N3346, N3343);
or OR2 (N3347, N3344, N958);
buf BUF1 (N3348, N3321);
and AND3 (N3349, N3347, N1295, N2244);
nor NOR2 (N3350, N3349, N1877);
not NOT1 (N3351, N3339);
and AND3 (N3352, N3348, N974, N2808);
buf BUF1 (N3353, N3351);
and AND3 (N3354, N3353, N1852, N1545);
buf BUF1 (N3355, N3346);
and AND2 (N3356, N3350, N1427);
xor XOR2 (N3357, N3354, N1261);
or OR2 (N3358, N3357, N499);
nor NOR2 (N3359, N3345, N3116);
xor XOR2 (N3360, N3355, N1327);
buf BUF1 (N3361, N3359);
nor NOR4 (N3362, N3360, N289, N167, N546);
nor NOR3 (N3363, N3330, N3125, N3181);
nand NAND3 (N3364, N3358, N1454, N3231);
and AND2 (N3365, N3362, N3009);
xor XOR2 (N3366, N3356, N1541);
not NOT1 (N3367, N3342);
buf BUF1 (N3368, N3366);
not NOT1 (N3369, N3335);
buf BUF1 (N3370, N3363);
xor XOR2 (N3371, N3367, N1428);
buf BUF1 (N3372, N3361);
xor XOR2 (N3373, N3370, N2906);
xor XOR2 (N3374, N3372, N2384);
nor NOR4 (N3375, N3365, N1647, N1091, N1580);
not NOT1 (N3376, N3371);
not NOT1 (N3377, N3352);
nand NAND2 (N3378, N3364, N2300);
xor XOR2 (N3379, N3337, N1841);
xor XOR2 (N3380, N3376, N2446);
or OR3 (N3381, N3378, N3316, N3108);
xor XOR2 (N3382, N3375, N2445);
xor XOR2 (N3383, N3382, N2750);
nand NAND2 (N3384, N3379, N1229);
or OR2 (N3385, N3383, N3365);
and AND2 (N3386, N3380, N2797);
and AND3 (N3387, N3374, N512, N2775);
buf BUF1 (N3388, N3381);
xor XOR2 (N3389, N3336, N756);
xor XOR2 (N3390, N3388, N2592);
buf BUF1 (N3391, N3386);
buf BUF1 (N3392, N3373);
and AND2 (N3393, N3385, N429);
nand NAND3 (N3394, N3390, N1172, N557);
xor XOR2 (N3395, N3387, N3244);
nor NOR4 (N3396, N3395, N558, N1727, N2945);
not NOT1 (N3397, N3389);
xor XOR2 (N3398, N3394, N2442);
or OR2 (N3399, N3384, N102);
xor XOR2 (N3400, N3393, N2911);
xor XOR2 (N3401, N3368, N173);
nor NOR2 (N3402, N3397, N305);
and AND2 (N3403, N3396, N1932);
nor NOR4 (N3404, N3402, N1432, N3369, N2541);
buf BUF1 (N3405, N2202);
buf BUF1 (N3406, N3377);
or OR4 (N3407, N3398, N1667, N2287, N1618);
nor NOR4 (N3408, N3391, N2556, N1866, N2636);
nand NAND2 (N3409, N3406, N2784);
nand NAND2 (N3410, N3399, N812);
and AND2 (N3411, N3410, N1322);
xor XOR2 (N3412, N3408, N1684);
or OR3 (N3413, N3411, N239, N782);
nor NOR2 (N3414, N3407, N299);
and AND4 (N3415, N3401, N97, N707, N2408);
and AND4 (N3416, N3405, N3264, N239, N770);
buf BUF1 (N3417, N3416);
nor NOR2 (N3418, N3413, N864);
and AND2 (N3419, N3404, N3404);
and AND3 (N3420, N3417, N645, N192);
buf BUF1 (N3421, N3418);
nor NOR3 (N3422, N3419, N1011, N1393);
and AND3 (N3423, N3421, N3213, N1199);
and AND4 (N3424, N3422, N906, N636, N1373);
not NOT1 (N3425, N3412);
or OR4 (N3426, N3400, N1758, N2377, N2289);
and AND4 (N3427, N3424, N2511, N783, N2256);
buf BUF1 (N3428, N3409);
buf BUF1 (N3429, N3415);
or OR2 (N3430, N3427, N280);
or OR2 (N3431, N3403, N2445);
not NOT1 (N3432, N3392);
xor XOR2 (N3433, N3414, N1170);
nor NOR3 (N3434, N3431, N1059, N2462);
buf BUF1 (N3435, N3429);
nor NOR3 (N3436, N3435, N2710, N3199);
nor NOR3 (N3437, N3433, N3311, N1389);
nand NAND3 (N3438, N3432, N3219, N47);
nand NAND4 (N3439, N3423, N3179, N126, N2367);
not NOT1 (N3440, N3434);
xor XOR2 (N3441, N3420, N679);
or OR4 (N3442, N3437, N1549, N1136, N2271);
buf BUF1 (N3443, N3438);
not NOT1 (N3444, N3441);
buf BUF1 (N3445, N3430);
xor XOR2 (N3446, N3425, N2163);
buf BUF1 (N3447, N3428);
nand NAND4 (N3448, N3439, N1292, N3086, N2828);
nand NAND2 (N3449, N3447, N633);
or OR3 (N3450, N3444, N3221, N1821);
buf BUF1 (N3451, N3442);
or OR4 (N3452, N3446, N2257, N2414, N2535);
or OR4 (N3453, N3451, N1803, N62, N226);
or OR2 (N3454, N3449, N450);
xor XOR2 (N3455, N3454, N2336);
nor NOR4 (N3456, N3455, N3049, N557, N693);
buf BUF1 (N3457, N3450);
nand NAND4 (N3458, N3448, N2672, N1598, N3190);
or OR4 (N3459, N3457, N3173, N1270, N2974);
nand NAND2 (N3460, N3445, N2413);
nand NAND4 (N3461, N3436, N2268, N3055, N2696);
nand NAND2 (N3462, N3456, N1062);
xor XOR2 (N3463, N3462, N2130);
nor NOR4 (N3464, N3440, N1160, N1574, N483);
or OR4 (N3465, N3453, N334, N3055, N1340);
and AND2 (N3466, N3464, N2454);
nand NAND3 (N3467, N3461, N514, N3070);
not NOT1 (N3468, N3465);
xor XOR2 (N3469, N3466, N622);
nand NAND4 (N3470, N3443, N1695, N114, N2696);
and AND3 (N3471, N3467, N179, N3043);
nand NAND3 (N3472, N3452, N986, N2953);
xor XOR2 (N3473, N3458, N1736);
not NOT1 (N3474, N3463);
or OR4 (N3475, N3460, N2446, N2101, N3085);
or OR4 (N3476, N3474, N1968, N58, N1774);
xor XOR2 (N3477, N3459, N2308);
or OR2 (N3478, N3473, N298);
xor XOR2 (N3479, N3475, N1872);
not NOT1 (N3480, N3472);
nor NOR3 (N3481, N3480, N2599, N3307);
nand NAND4 (N3482, N3476, N3368, N1388, N253);
nor NOR2 (N3483, N3477, N1775);
buf BUF1 (N3484, N3478);
not NOT1 (N3485, N3426);
xor XOR2 (N3486, N3485, N2675);
nand NAND3 (N3487, N3483, N1704, N1772);
and AND4 (N3488, N3479, N103, N1230, N1593);
and AND3 (N3489, N3486, N1280, N541);
buf BUF1 (N3490, N3470);
and AND4 (N3491, N3488, N463, N312, N2503);
nor NOR4 (N3492, N3468, N1282, N372, N2591);
nor NOR3 (N3493, N3490, N1901, N3395);
not NOT1 (N3494, N3493);
xor XOR2 (N3495, N3471, N3354);
nand NAND2 (N3496, N3482, N445);
nor NOR3 (N3497, N3484, N1015, N1883);
not NOT1 (N3498, N3469);
not NOT1 (N3499, N3498);
nor NOR2 (N3500, N3489, N471);
not NOT1 (N3501, N3500);
or OR2 (N3502, N3481, N845);
buf BUF1 (N3503, N3492);
and AND4 (N3504, N3503, N1076, N2828, N2872);
and AND2 (N3505, N3504, N2455);
xor XOR2 (N3506, N3501, N2410);
nor NOR3 (N3507, N3487, N3231, N3338);
not NOT1 (N3508, N3495);
nor NOR4 (N3509, N3496, N2172, N586, N3505);
xor XOR2 (N3510, N235, N301);
or OR2 (N3511, N3510, N1271);
or OR4 (N3512, N3507, N2379, N2366, N2046);
nand NAND2 (N3513, N3509, N3363);
or OR2 (N3514, N3506, N3331);
nor NOR4 (N3515, N3499, N145, N3404, N53);
nand NAND3 (N3516, N3494, N1796, N2166);
buf BUF1 (N3517, N3491);
xor XOR2 (N3518, N3517, N1374);
not NOT1 (N3519, N3513);
and AND4 (N3520, N3519, N522, N2599, N3341);
not NOT1 (N3521, N3520);
and AND3 (N3522, N3512, N2595, N1890);
nand NAND4 (N3523, N3518, N99, N480, N1656);
and AND4 (N3524, N3515, N2369, N297, N2595);
nor NOR3 (N3525, N3508, N2840, N2011);
not NOT1 (N3526, N3514);
and AND4 (N3527, N3524, N1127, N2984, N3156);
not NOT1 (N3528, N3511);
nand NAND3 (N3529, N3497, N1084, N2003);
xor XOR2 (N3530, N3525, N481);
not NOT1 (N3531, N3516);
buf BUF1 (N3532, N3530);
xor XOR2 (N3533, N3523, N2938);
and AND3 (N3534, N3527, N1092, N1406);
buf BUF1 (N3535, N3531);
xor XOR2 (N3536, N3534, N1425);
or OR2 (N3537, N3536, N2816);
buf BUF1 (N3538, N3526);
nor NOR4 (N3539, N3502, N2009, N2975, N47);
buf BUF1 (N3540, N3522);
not NOT1 (N3541, N3533);
or OR2 (N3542, N3532, N2052);
xor XOR2 (N3543, N3521, N1076);
buf BUF1 (N3544, N3535);
nand NAND4 (N3545, N3542, N2108, N3410, N149);
xor XOR2 (N3546, N3537, N2064);
buf BUF1 (N3547, N3546);
nor NOR4 (N3548, N3547, N671, N2931, N3405);
and AND4 (N3549, N3539, N927, N1996, N1791);
and AND3 (N3550, N3548, N2466, N1852);
not NOT1 (N3551, N3543);
or OR4 (N3552, N3545, N3109, N2455, N340);
not NOT1 (N3553, N3541);
xor XOR2 (N3554, N3529, N1849);
nand NAND3 (N3555, N3528, N2540, N3528);
buf BUF1 (N3556, N3555);
not NOT1 (N3557, N3549);
and AND4 (N3558, N3554, N1000, N1656, N1097);
nand NAND3 (N3559, N3540, N656, N2113);
buf BUF1 (N3560, N3551);
xor XOR2 (N3561, N3557, N2932);
or OR2 (N3562, N3559, N1645);
not NOT1 (N3563, N3562);
nand NAND3 (N3564, N3556, N2762, N69);
buf BUF1 (N3565, N3558);
nand NAND2 (N3566, N3560, N2495);
nor NOR4 (N3567, N3550, N2110, N1553, N3556);
buf BUF1 (N3568, N3563);
or OR2 (N3569, N3552, N1418);
or OR3 (N3570, N3553, N3361, N1753);
nor NOR3 (N3571, N3538, N710, N2446);
buf BUF1 (N3572, N3561);
nor NOR2 (N3573, N3567, N2639);
buf BUF1 (N3574, N3573);
xor XOR2 (N3575, N3565, N2952);
nand NAND2 (N3576, N3544, N3105);
buf BUF1 (N3577, N3575);
buf BUF1 (N3578, N3569);
nand NAND2 (N3579, N3570, N2011);
buf BUF1 (N3580, N3574);
xor XOR2 (N3581, N3564, N1561);
or OR4 (N3582, N3579, N2826, N2463, N531);
nor NOR2 (N3583, N3566, N2284);
or OR2 (N3584, N3580, N2283);
not NOT1 (N3585, N3582);
xor XOR2 (N3586, N3584, N368);
and AND3 (N3587, N3578, N3323, N2301);
not NOT1 (N3588, N3587);
buf BUF1 (N3589, N3576);
buf BUF1 (N3590, N3586);
and AND2 (N3591, N3590, N363);
xor XOR2 (N3592, N3589, N2257);
nand NAND2 (N3593, N3591, N1703);
not NOT1 (N3594, N3583);
buf BUF1 (N3595, N3581);
nor NOR2 (N3596, N3571, N222);
or OR2 (N3597, N3588, N1284);
not NOT1 (N3598, N3596);
and AND2 (N3599, N3594, N2517);
buf BUF1 (N3600, N3585);
and AND4 (N3601, N3597, N589, N2587, N1666);
not NOT1 (N3602, N3577);
nor NOR3 (N3603, N3598, N187, N1793);
xor XOR2 (N3604, N3602, N4);
not NOT1 (N3605, N3600);
not NOT1 (N3606, N3603);
nand NAND4 (N3607, N3592, N168, N2904, N1276);
buf BUF1 (N3608, N3605);
buf BUF1 (N3609, N3607);
xor XOR2 (N3610, N3601, N893);
and AND4 (N3611, N3595, N1115, N2305, N1913);
xor XOR2 (N3612, N3599, N2914);
or OR4 (N3613, N3609, N3578, N3140, N630);
nand NAND2 (N3614, N3608, N2708);
nor NOR2 (N3615, N3612, N1696);
buf BUF1 (N3616, N3568);
xor XOR2 (N3617, N3611, N1671);
buf BUF1 (N3618, N3572);
nand NAND4 (N3619, N3610, N2931, N1495, N3491);
and AND3 (N3620, N3617, N2449, N2116);
not NOT1 (N3621, N3593);
nor NOR4 (N3622, N3614, N1436, N3079, N601);
buf BUF1 (N3623, N3618);
and AND4 (N3624, N3616, N550, N2375, N1682);
nand NAND2 (N3625, N3623, N1272);
and AND4 (N3626, N3621, N818, N1212, N3100);
not NOT1 (N3627, N3622);
nor NOR3 (N3628, N3615, N815, N429);
xor XOR2 (N3629, N3627, N1678);
buf BUF1 (N3630, N3619);
not NOT1 (N3631, N3630);
and AND2 (N3632, N3628, N1570);
xor XOR2 (N3633, N3625, N3028);
and AND2 (N3634, N3620, N3284);
not NOT1 (N3635, N3613);
or OR3 (N3636, N3633, N236, N1614);
xor XOR2 (N3637, N3632, N321);
nor NOR3 (N3638, N3635, N2081, N3278);
nor NOR3 (N3639, N3634, N1058, N3395);
not NOT1 (N3640, N3637);
not NOT1 (N3641, N3636);
xor XOR2 (N3642, N3638, N994);
not NOT1 (N3643, N3642);
xor XOR2 (N3644, N3639, N3279);
or OR3 (N3645, N3624, N2155, N259);
not NOT1 (N3646, N3645);
and AND2 (N3647, N3641, N3272);
and AND4 (N3648, N3629, N1472, N272, N3485);
buf BUF1 (N3649, N3643);
or OR2 (N3650, N3626, N968);
or OR3 (N3651, N3631, N931, N687);
buf BUF1 (N3652, N3604);
xor XOR2 (N3653, N3640, N435);
and AND2 (N3654, N3650, N1085);
nor NOR3 (N3655, N3653, N1661, N2243);
nand NAND4 (N3656, N3655, N3462, N3365, N3030);
or OR4 (N3657, N3647, N356, N1819, N3566);
not NOT1 (N3658, N3654);
nor NOR2 (N3659, N3648, N492);
buf BUF1 (N3660, N3606);
and AND2 (N3661, N3649, N3202);
or OR4 (N3662, N3652, N42, N1094, N473);
buf BUF1 (N3663, N3662);
buf BUF1 (N3664, N3644);
xor XOR2 (N3665, N3651, N27);
buf BUF1 (N3666, N3658);
buf BUF1 (N3667, N3657);
or OR2 (N3668, N3663, N1916);
xor XOR2 (N3669, N3656, N1116);
not NOT1 (N3670, N3660);
nand NAND3 (N3671, N3666, N1517, N348);
buf BUF1 (N3672, N3668);
nor NOR4 (N3673, N3646, N728, N671, N629);
nand NAND3 (N3674, N3667, N3327, N146);
not NOT1 (N3675, N3672);
or OR2 (N3676, N3670, N1924);
not NOT1 (N3677, N3665);
nor NOR3 (N3678, N3669, N2208, N1449);
nor NOR3 (N3679, N3675, N1483, N3581);
or OR2 (N3680, N3661, N932);
and AND2 (N3681, N3680, N3584);
nand NAND4 (N3682, N3677, N734, N1429, N85);
buf BUF1 (N3683, N3676);
buf BUF1 (N3684, N3683);
and AND2 (N3685, N3681, N3336);
not NOT1 (N3686, N3679);
nor NOR4 (N3687, N3684, N1694, N1031, N2500);
xor XOR2 (N3688, N3678, N2283);
xor XOR2 (N3689, N3673, N425);
or OR4 (N3690, N3682, N3459, N3314, N316);
and AND3 (N3691, N3687, N390, N2646);
not NOT1 (N3692, N3689);
xor XOR2 (N3693, N3690, N1080);
xor XOR2 (N3694, N3674, N2848);
buf BUF1 (N3695, N3691);
xor XOR2 (N3696, N3671, N3536);
xor XOR2 (N3697, N3693, N3374);
and AND2 (N3698, N3685, N2856);
nand NAND2 (N3699, N3659, N264);
xor XOR2 (N3700, N3697, N3353);
nor NOR3 (N3701, N3698, N292, N1068);
or OR2 (N3702, N3688, N2921);
not NOT1 (N3703, N3664);
buf BUF1 (N3704, N3692);
and AND2 (N3705, N3696, N1217);
nor NOR4 (N3706, N3695, N3136, N2833, N776);
not NOT1 (N3707, N3699);
not NOT1 (N3708, N3701);
nor NOR4 (N3709, N3707, N3189, N415, N1174);
not NOT1 (N3710, N3686);
xor XOR2 (N3711, N3704, N3196);
and AND2 (N3712, N3706, N3684);
not NOT1 (N3713, N3700);
nand NAND2 (N3714, N3709, N1844);
or OR3 (N3715, N3705, N2203, N2413);
nand NAND2 (N3716, N3702, N736);
nand NAND2 (N3717, N3716, N3038);
and AND3 (N3718, N3703, N449, N438);
not NOT1 (N3719, N3708);
and AND2 (N3720, N3719, N3291);
nor NOR4 (N3721, N3711, N592, N3239, N3685);
buf BUF1 (N3722, N3718);
nor NOR4 (N3723, N3713, N2867, N3009, N77);
xor XOR2 (N3724, N3720, N2456);
nor NOR4 (N3725, N3722, N1418, N1853, N3050);
xor XOR2 (N3726, N3712, N580);
or OR4 (N3727, N3721, N2545, N2491, N1507);
or OR2 (N3728, N3725, N2554);
not NOT1 (N3729, N3710);
or OR3 (N3730, N3724, N2435, N2698);
xor XOR2 (N3731, N3730, N3226);
nand NAND3 (N3732, N3727, N2038, N2150);
and AND4 (N3733, N3715, N1230, N1187, N2721);
buf BUF1 (N3734, N3726);
and AND2 (N3735, N3728, N3545);
buf BUF1 (N3736, N3729);
nand NAND2 (N3737, N3736, N1926);
not NOT1 (N3738, N3714);
xor XOR2 (N3739, N3723, N2036);
or OR4 (N3740, N3732, N1619, N696, N1107);
not NOT1 (N3741, N3735);
and AND2 (N3742, N3740, N3251);
buf BUF1 (N3743, N3717);
and AND2 (N3744, N3743, N3438);
and AND3 (N3745, N3744, N1719, N2023);
nand NAND2 (N3746, N3738, N3601);
and AND4 (N3747, N3742, N3302, N1476, N3677);
buf BUF1 (N3748, N3745);
buf BUF1 (N3749, N3747);
and AND4 (N3750, N3731, N3636, N1624, N1913);
nand NAND4 (N3751, N3741, N562, N1556, N1902);
or OR3 (N3752, N3746, N2742, N1822);
buf BUF1 (N3753, N3734);
nor NOR4 (N3754, N3733, N941, N606, N2328);
buf BUF1 (N3755, N3737);
and AND4 (N3756, N3694, N1760, N2193, N3637);
not NOT1 (N3757, N3755);
xor XOR2 (N3758, N3749, N1384);
xor XOR2 (N3759, N3753, N3541);
xor XOR2 (N3760, N3754, N2588);
or OR2 (N3761, N3758, N223);
nor NOR2 (N3762, N3756, N1924);
and AND4 (N3763, N3751, N2631, N400, N1771);
and AND2 (N3764, N3757, N3695);
nand NAND3 (N3765, N3764, N3098, N321);
not NOT1 (N3766, N3750);
not NOT1 (N3767, N3765);
nor NOR4 (N3768, N3759, N2236, N537, N2745);
nand NAND4 (N3769, N3739, N549, N778, N1785);
buf BUF1 (N3770, N3760);
nor NOR3 (N3771, N3762, N407, N1140);
nand NAND2 (N3772, N3748, N738);
not NOT1 (N3773, N3768);
and AND3 (N3774, N3773, N1050, N2803);
not NOT1 (N3775, N3769);
not NOT1 (N3776, N3771);
nor NOR2 (N3777, N3752, N843);
nor NOR4 (N3778, N3777, N2048, N1124, N3092);
xor XOR2 (N3779, N3767, N1379);
or OR3 (N3780, N3770, N977, N2583);
or OR4 (N3781, N3779, N3296, N1848, N2358);
not NOT1 (N3782, N3766);
nand NAND4 (N3783, N3781, N749, N1576, N2404);
buf BUF1 (N3784, N3782);
nor NOR4 (N3785, N3783, N2658, N1014, N878);
and AND3 (N3786, N3774, N1888, N2596);
not NOT1 (N3787, N3763);
and AND3 (N3788, N3776, N2195, N1287);
nand NAND4 (N3789, N3788, N3015, N2914, N885);
or OR3 (N3790, N3789, N2361, N3530);
xor XOR2 (N3791, N3775, N1992);
nor NOR4 (N3792, N3780, N2000, N77, N665);
and AND2 (N3793, N3784, N1631);
not NOT1 (N3794, N3792);
buf BUF1 (N3795, N3787);
xor XOR2 (N3796, N3794, N3414);
or OR3 (N3797, N3793, N357, N2327);
not NOT1 (N3798, N3795);
nand NAND2 (N3799, N3798, N2963);
or OR4 (N3800, N3772, N187, N1383, N113);
nand NAND3 (N3801, N3761, N2909, N3233);
or OR3 (N3802, N3786, N1402, N709);
xor XOR2 (N3803, N3790, N3228);
xor XOR2 (N3804, N3802, N1182);
nand NAND2 (N3805, N3801, N1258);
or OR3 (N3806, N3778, N8, N2943);
nor NOR3 (N3807, N3791, N729, N1855);
nand NAND2 (N3808, N3785, N3437);
nor NOR2 (N3809, N3803, N473);
and AND4 (N3810, N3805, N2924, N2613, N2058);
and AND3 (N3811, N3809, N1910, N579);
not NOT1 (N3812, N3800);
and AND4 (N3813, N3812, N3730, N843, N2978);
nand NAND4 (N3814, N3811, N3179, N1017, N3357);
xor XOR2 (N3815, N3804, N3265);
or OR3 (N3816, N3815, N1997, N3233);
nor NOR4 (N3817, N3796, N1888, N2366, N3095);
nand NAND2 (N3818, N3808, N2870);
nor NOR2 (N3819, N3814, N2301);
xor XOR2 (N3820, N3806, N2699);
not NOT1 (N3821, N3819);
xor XOR2 (N3822, N3820, N2759);
or OR4 (N3823, N3799, N2433, N2036, N628);
nor NOR4 (N3824, N3807, N3656, N2839, N548);
xor XOR2 (N3825, N3824, N1979);
nor NOR3 (N3826, N3822, N2748, N2240);
nand NAND2 (N3827, N3825, N3417);
nor NOR3 (N3828, N3817, N38, N3163);
not NOT1 (N3829, N3823);
or OR4 (N3830, N3827, N1235, N2987, N3262);
nor NOR4 (N3831, N3813, N1981, N16, N115);
and AND2 (N3832, N3821, N1362);
or OR4 (N3833, N3818, N3109, N2224, N2921);
xor XOR2 (N3834, N3816, N1989);
and AND4 (N3835, N3830, N1893, N1211, N3460);
and AND4 (N3836, N3826, N2231, N1271, N2918);
or OR4 (N3837, N3835, N1912, N208, N271);
and AND3 (N3838, N3836, N1306, N2539);
xor XOR2 (N3839, N3837, N2441);
nand NAND3 (N3840, N3828, N1134, N324);
nor NOR2 (N3841, N3839, N1590);
nand NAND2 (N3842, N3841, N733);
and AND2 (N3843, N3842, N547);
nor NOR4 (N3844, N3833, N1379, N2193, N3690);
xor XOR2 (N3845, N3840, N2543);
buf BUF1 (N3846, N3829);
xor XOR2 (N3847, N3846, N1618);
xor XOR2 (N3848, N3844, N748);
xor XOR2 (N3849, N3832, N413);
or OR3 (N3850, N3810, N1947, N3148);
or OR2 (N3851, N3831, N2865);
not NOT1 (N3852, N3834);
not NOT1 (N3853, N3851);
nand NAND2 (N3854, N3843, N2748);
buf BUF1 (N3855, N3848);
or OR2 (N3856, N3850, N3615);
nor NOR4 (N3857, N3854, N1072, N1931, N110);
buf BUF1 (N3858, N3857);
not NOT1 (N3859, N3853);
not NOT1 (N3860, N3856);
nand NAND2 (N3861, N3852, N3519);
and AND4 (N3862, N3855, N1499, N3555, N196);
or OR2 (N3863, N3859, N69);
not NOT1 (N3864, N3858);
or OR4 (N3865, N3797, N3029, N2891, N2749);
not NOT1 (N3866, N3864);
nand NAND2 (N3867, N3860, N243);
xor XOR2 (N3868, N3849, N2992);
nor NOR3 (N3869, N3866, N3418, N2853);
and AND3 (N3870, N3865, N832, N545);
or OR3 (N3871, N3869, N3248, N275);
xor XOR2 (N3872, N3862, N333);
or OR4 (N3873, N3872, N2417, N3465, N1785);
xor XOR2 (N3874, N3861, N2676);
or OR2 (N3875, N3873, N554);
or OR3 (N3876, N3870, N3850, N3642);
or OR3 (N3877, N3845, N1118, N582);
or OR4 (N3878, N3863, N3024, N3501, N795);
nand NAND2 (N3879, N3875, N128);
or OR2 (N3880, N3838, N2017);
xor XOR2 (N3881, N3871, N3258);
nand NAND2 (N3882, N3877, N2606);
xor XOR2 (N3883, N3868, N116);
buf BUF1 (N3884, N3867);
buf BUF1 (N3885, N3883);
nand NAND2 (N3886, N3878, N695);
not NOT1 (N3887, N3876);
and AND3 (N3888, N3882, N140, N1554);
buf BUF1 (N3889, N3847);
xor XOR2 (N3890, N3886, N497);
nand NAND2 (N3891, N3889, N2148);
nand NAND3 (N3892, N3891, N112, N2041);
nand NAND3 (N3893, N3888, N1470, N2346);
xor XOR2 (N3894, N3880, N183);
not NOT1 (N3895, N3884);
nand NAND3 (N3896, N3885, N1237, N2877);
or OR2 (N3897, N3879, N1120);
not NOT1 (N3898, N3892);
not NOT1 (N3899, N3898);
nor NOR3 (N3900, N3874, N724, N510);
nand NAND2 (N3901, N3890, N3319);
xor XOR2 (N3902, N3895, N939);
or OR4 (N3903, N3896, N2166, N2714, N141);
xor XOR2 (N3904, N3897, N1694);
buf BUF1 (N3905, N3887);
not NOT1 (N3906, N3881);
nand NAND3 (N3907, N3903, N644, N1170);
or OR2 (N3908, N3907, N3028);
not NOT1 (N3909, N3908);
and AND2 (N3910, N3904, N2404);
nor NOR4 (N3911, N3909, N3369, N3856, N257);
or OR2 (N3912, N3901, N2584);
nor NOR4 (N3913, N3912, N3617, N3163, N1755);
buf BUF1 (N3914, N3906);
or OR3 (N3915, N3913, N1895, N2795);
nand NAND3 (N3916, N3894, N2370, N2364);
buf BUF1 (N3917, N3900);
or OR2 (N3918, N3916, N2907);
or OR3 (N3919, N3902, N595, N2905);
and AND4 (N3920, N3918, N2661, N29, N2214);
nor NOR4 (N3921, N3920, N2117, N3131, N3468);
nand NAND4 (N3922, N3915, N1648, N3915, N1805);
buf BUF1 (N3923, N3911);
buf BUF1 (N3924, N3905);
nand NAND3 (N3925, N3914, N2278, N3401);
nor NOR4 (N3926, N3925, N2125, N54, N388);
or OR2 (N3927, N3923, N2663);
and AND2 (N3928, N3926, N919);
nand NAND2 (N3929, N3924, N2927);
and AND2 (N3930, N3922, N964);
not NOT1 (N3931, N3919);
buf BUF1 (N3932, N3910);
nand NAND4 (N3933, N3929, N580, N3500, N1768);
nor NOR2 (N3934, N3921, N1703);
not NOT1 (N3935, N3934);
xor XOR2 (N3936, N3935, N285);
buf BUF1 (N3937, N3893);
and AND3 (N3938, N3937, N2667, N3653);
nor NOR4 (N3939, N3936, N3069, N553, N1635);
nor NOR3 (N3940, N3928, N2752, N1304);
nand NAND2 (N3941, N3931, N1509);
not NOT1 (N3942, N3899);
and AND2 (N3943, N3917, N2203);
xor XOR2 (N3944, N3939, N587);
xor XOR2 (N3945, N3927, N3789);
xor XOR2 (N3946, N3945, N811);
and AND3 (N3947, N3940, N3488, N1154);
nor NOR2 (N3948, N3932, N2391);
and AND2 (N3949, N3933, N1860);
not NOT1 (N3950, N3942);
buf BUF1 (N3951, N3949);
nand NAND3 (N3952, N3948, N2845, N147);
or OR2 (N3953, N3947, N3468);
buf BUF1 (N3954, N3953);
buf BUF1 (N3955, N3954);
or OR2 (N3956, N3943, N1924);
or OR4 (N3957, N3955, N1737, N1592, N580);
and AND2 (N3958, N3946, N2747);
or OR2 (N3959, N3956, N1401);
and AND3 (N3960, N3944, N2113, N3949);
not NOT1 (N3961, N3958);
not NOT1 (N3962, N3930);
nand NAND4 (N3963, N3957, N2445, N1535, N591);
nor NOR3 (N3964, N3962, N725, N3676);
nand NAND3 (N3965, N3950, N764, N2609);
and AND3 (N3966, N3960, N3667, N1971);
not NOT1 (N3967, N3951);
not NOT1 (N3968, N3941);
or OR3 (N3969, N3965, N3243, N2905);
xor XOR2 (N3970, N3968, N3944);
not NOT1 (N3971, N3969);
not NOT1 (N3972, N3961);
xor XOR2 (N3973, N3970, N1526);
buf BUF1 (N3974, N3959);
nand NAND2 (N3975, N3964, N1246);
or OR2 (N3976, N3972, N1244);
buf BUF1 (N3977, N3971);
nor NOR4 (N3978, N3976, N924, N3442, N229);
and AND3 (N3979, N3963, N2515, N3893);
buf BUF1 (N3980, N3966);
xor XOR2 (N3981, N3977, N2401);
buf BUF1 (N3982, N3974);
and AND2 (N3983, N3978, N1886);
nor NOR2 (N3984, N3973, N3548);
xor XOR2 (N3985, N3952, N2071);
nand NAND2 (N3986, N3981, N603);
or OR4 (N3987, N3982, N681, N1955, N1426);
nand NAND3 (N3988, N3985, N1949, N54);
xor XOR2 (N3989, N3967, N1142);
not NOT1 (N3990, N3983);
xor XOR2 (N3991, N3988, N307);
xor XOR2 (N3992, N3987, N1857);
xor XOR2 (N3993, N3991, N3604);
not NOT1 (N3994, N3938);
and AND4 (N3995, N3979, N1879, N164, N3920);
and AND2 (N3996, N3989, N1831);
nand NAND2 (N3997, N3975, N292);
nor NOR3 (N3998, N3997, N2395, N3019);
nand NAND2 (N3999, N3998, N1226);
and AND4 (N4000, N3996, N1307, N3001, N301);
nor NOR2 (N4001, N3980, N2984);
buf BUF1 (N4002, N3993);
or OR3 (N4003, N3990, N636, N2975);
xor XOR2 (N4004, N3984, N1358);
buf BUF1 (N4005, N4001);
and AND4 (N4006, N3992, N3265, N1542, N754);
not NOT1 (N4007, N3999);
and AND4 (N4008, N4000, N171, N1253, N974);
not NOT1 (N4009, N4008);
nor NOR4 (N4010, N4006, N1220, N365, N771);
and AND4 (N4011, N4002, N3202, N3136, N883);
not NOT1 (N4012, N4007);
xor XOR2 (N4013, N4011, N176);
or OR4 (N4014, N3986, N2948, N2314, N4010);
xor XOR2 (N4015, N2447, N477);
nand NAND3 (N4016, N4013, N3629, N3134);
and AND2 (N4017, N4004, N3108);
buf BUF1 (N4018, N4014);
buf BUF1 (N4019, N4018);
xor XOR2 (N4020, N4003, N3419);
nor NOR2 (N4021, N4015, N1922);
xor XOR2 (N4022, N4005, N1941);
not NOT1 (N4023, N4009);
nand NAND4 (N4024, N4023, N3874, N604, N2143);
nor NOR2 (N4025, N3995, N1762);
buf BUF1 (N4026, N4022);
or OR4 (N4027, N4025, N2531, N2442, N3495);
buf BUF1 (N4028, N4012);
buf BUF1 (N4029, N4027);
nand NAND4 (N4030, N4019, N2047, N1983, N3618);
nand NAND4 (N4031, N4026, N1451, N1630, N1998);
xor XOR2 (N4032, N4024, N3774);
nand NAND3 (N4033, N4021, N3537, N3217);
xor XOR2 (N4034, N4030, N374);
or OR2 (N4035, N4029, N862);
buf BUF1 (N4036, N4020);
and AND2 (N4037, N3994, N1536);
nor NOR3 (N4038, N4034, N2383, N1681);
buf BUF1 (N4039, N4028);
or OR3 (N4040, N4017, N2915, N636);
buf BUF1 (N4041, N4031);
xor XOR2 (N4042, N4038, N3304);
xor XOR2 (N4043, N4016, N738);
nand NAND4 (N4044, N4043, N3680, N1489, N3169);
nor NOR4 (N4045, N4041, N357, N2447, N2947);
nor NOR2 (N4046, N4033, N2046);
nor NOR2 (N4047, N4046, N2545);
and AND3 (N4048, N4032, N3706, N1843);
and AND3 (N4049, N4044, N3567, N2738);
nor NOR3 (N4050, N4036, N3392, N3175);
xor XOR2 (N4051, N4049, N2932);
nor NOR3 (N4052, N4045, N3291, N3664);
nand NAND3 (N4053, N4051, N2403, N1912);
xor XOR2 (N4054, N4047, N1434);
or OR2 (N4055, N4037, N1253);
nand NAND2 (N4056, N4040, N17);
and AND2 (N4057, N4056, N3153);
nand NAND4 (N4058, N4050, N2383, N3244, N1235);
nor NOR4 (N4059, N4042, N1788, N301, N222);
nand NAND4 (N4060, N4048, N2487, N2463, N330);
xor XOR2 (N4061, N4057, N2396);
not NOT1 (N4062, N4059);
and AND4 (N4063, N4054, N3188, N1206, N1476);
or OR2 (N4064, N4039, N1015);
nand NAND3 (N4065, N4052, N1352, N1171);
xor XOR2 (N4066, N4061, N1740);
not NOT1 (N4067, N4053);
and AND2 (N4068, N4064, N2388);
nor NOR4 (N4069, N4035, N588, N1570, N155);
and AND4 (N4070, N4065, N3779, N2213, N2950);
and AND4 (N4071, N4060, N3659, N1237, N903);
xor XOR2 (N4072, N4071, N1669);
not NOT1 (N4073, N4063);
nand NAND4 (N4074, N4055, N2619, N1950, N2638);
or OR3 (N4075, N4073, N4001, N228);
nand NAND4 (N4076, N4067, N3446, N1524, N1028);
buf BUF1 (N4077, N4072);
buf BUF1 (N4078, N4068);
nand NAND4 (N4079, N4069, N38, N3045, N1199);
nand NAND3 (N4080, N4076, N1679, N820);
and AND2 (N4081, N4074, N2674);
or OR3 (N4082, N4058, N3142, N3483);
nand NAND3 (N4083, N4078, N2011, N1168);
xor XOR2 (N4084, N4062, N602);
and AND3 (N4085, N4079, N4046, N408);
or OR3 (N4086, N4077, N230, N2675);
nand NAND3 (N4087, N4085, N1945, N4047);
buf BUF1 (N4088, N4081);
or OR4 (N4089, N4086, N1499, N2559, N4019);
xor XOR2 (N4090, N4082, N2806);
buf BUF1 (N4091, N4066);
buf BUF1 (N4092, N4083);
nor NOR4 (N4093, N4089, N603, N3990, N3013);
nor NOR3 (N4094, N4080, N2326, N1602);
xor XOR2 (N4095, N4094, N3708);
nand NAND4 (N4096, N4092, N2230, N607, N1352);
xor XOR2 (N4097, N4090, N1255);
buf BUF1 (N4098, N4095);
xor XOR2 (N4099, N4087, N2942);
or OR3 (N4100, N4093, N4052, N2630);
nor NOR4 (N4101, N4096, N2006, N1302, N3225);
xor XOR2 (N4102, N4100, N1005);
xor XOR2 (N4103, N4098, N2680);
xor XOR2 (N4104, N4091, N1199);
not NOT1 (N4105, N4099);
nor NOR2 (N4106, N4097, N1034);
or OR4 (N4107, N4088, N934, N3187, N3984);
buf BUF1 (N4108, N4070);
xor XOR2 (N4109, N4102, N1397);
not NOT1 (N4110, N4106);
nor NOR2 (N4111, N4104, N1088);
xor XOR2 (N4112, N4084, N1932);
and AND4 (N4113, N4110, N3498, N1513, N2342);
nor NOR3 (N4114, N4101, N1762, N3480);
nor NOR4 (N4115, N4109, N3255, N3428, N1317);
and AND3 (N4116, N4115, N3952, N228);
and AND2 (N4117, N4108, N2138);
nor NOR3 (N4118, N4103, N3890, N3495);
nor NOR3 (N4119, N4107, N3857, N1246);
and AND4 (N4120, N4118, N3350, N2211, N3410);
not NOT1 (N4121, N4117);
nor NOR4 (N4122, N4120, N3346, N692, N2226);
or OR2 (N4123, N4121, N2860);
not NOT1 (N4124, N4113);
nor NOR3 (N4125, N4075, N4119, N4115);
buf BUF1 (N4126, N1292);
xor XOR2 (N4127, N4123, N2259);
nand NAND4 (N4128, N4112, N1279, N3690, N3109);
xor XOR2 (N4129, N4111, N2253);
not NOT1 (N4130, N4125);
not NOT1 (N4131, N4105);
or OR2 (N4132, N4124, N2727);
buf BUF1 (N4133, N4122);
nand NAND3 (N4134, N4131, N464, N1137);
xor XOR2 (N4135, N4130, N1514);
buf BUF1 (N4136, N4128);
buf BUF1 (N4137, N4136);
nor NOR3 (N4138, N4116, N298, N912);
or OR3 (N4139, N4114, N94, N1480);
or OR3 (N4140, N4139, N2216, N940);
or OR2 (N4141, N4140, N2070);
or OR4 (N4142, N4137, N1883, N3679, N3348);
xor XOR2 (N4143, N4133, N3204);
nor NOR4 (N4144, N4132, N1418, N3252, N3135);
or OR3 (N4145, N4126, N3380, N2785);
nor NOR2 (N4146, N4141, N3789);
xor XOR2 (N4147, N4146, N3523);
nor NOR2 (N4148, N4147, N486);
xor XOR2 (N4149, N4134, N2736);
and AND4 (N4150, N4143, N1905, N1133, N1515);
nand NAND4 (N4151, N4150, N1974, N748, N1357);
nand NAND4 (N4152, N4135, N3839, N2595, N1521);
xor XOR2 (N4153, N4149, N2389);
buf BUF1 (N4154, N4127);
not NOT1 (N4155, N4153);
and AND4 (N4156, N4152, N2380, N2857, N605);
nand NAND4 (N4157, N4142, N1858, N3331, N2928);
nand NAND4 (N4158, N4156, N2869, N710, N2136);
nor NOR4 (N4159, N4145, N981, N1528, N566);
nor NOR4 (N4160, N4159, N2790, N1950, N1863);
nand NAND4 (N4161, N4154, N3145, N2580, N1738);
not NOT1 (N4162, N4138);
or OR4 (N4163, N4144, N492, N1894, N162);
nand NAND3 (N4164, N4148, N3990, N2085);
buf BUF1 (N4165, N4155);
xor XOR2 (N4166, N4160, N951);
and AND2 (N4167, N4129, N2645);
buf BUF1 (N4168, N4162);
buf BUF1 (N4169, N4158);
and AND4 (N4170, N4166, N1872, N2671, N3197);
buf BUF1 (N4171, N4170);
xor XOR2 (N4172, N4161, N20);
buf BUF1 (N4173, N4168);
xor XOR2 (N4174, N4165, N4101);
nand NAND3 (N4175, N4169, N285, N2002);
or OR3 (N4176, N4157, N3898, N1009);
nor NOR3 (N4177, N4167, N2764, N1284);
buf BUF1 (N4178, N4176);
xor XOR2 (N4179, N4151, N3207);
nand NAND4 (N4180, N4178, N3121, N2318, N1474);
and AND3 (N4181, N4180, N1139, N2066);
and AND3 (N4182, N4179, N1865, N534);
buf BUF1 (N4183, N4171);
buf BUF1 (N4184, N4181);
buf BUF1 (N4185, N4175);
buf BUF1 (N4186, N4163);
not NOT1 (N4187, N4177);
nor NOR3 (N4188, N4164, N3974, N2884);
or OR3 (N4189, N4184, N3547, N1247);
xor XOR2 (N4190, N4186, N1196);
and AND3 (N4191, N4182, N3515, N358);
nor NOR2 (N4192, N4188, N3164);
nor NOR4 (N4193, N4189, N1196, N4084, N3953);
or OR4 (N4194, N4183, N1095, N2268, N2595);
xor XOR2 (N4195, N4187, N3938);
nand NAND3 (N4196, N4192, N2048, N1218);
and AND2 (N4197, N4185, N2650);
xor XOR2 (N4198, N4172, N1891);
nand NAND2 (N4199, N4173, N4174);
nor NOR3 (N4200, N423, N1317, N2627);
nor NOR4 (N4201, N4193, N261, N3818, N270);
xor XOR2 (N4202, N4199, N697);
nor NOR3 (N4203, N4190, N2110, N2633);
or OR2 (N4204, N4191, N3564);
and AND4 (N4205, N4196, N2169, N63, N1521);
buf BUF1 (N4206, N4203);
nor NOR4 (N4207, N4202, N2966, N1706, N1880);
nand NAND3 (N4208, N4207, N20, N1521);
xor XOR2 (N4209, N4194, N1506);
and AND2 (N4210, N4198, N2783);
nor NOR4 (N4211, N4205, N3318, N485, N3141);
not NOT1 (N4212, N4210);
or OR2 (N4213, N4204, N3570);
nand NAND2 (N4214, N4201, N112);
not NOT1 (N4215, N4209);
and AND2 (N4216, N4214, N1545);
not NOT1 (N4217, N4208);
nand NAND3 (N4218, N4215, N3666, N3683);
buf BUF1 (N4219, N4212);
and AND3 (N4220, N4218, N1551, N2146);
nand NAND3 (N4221, N4216, N1014, N2722);
or OR4 (N4222, N4211, N1926, N1447, N483);
nand NAND3 (N4223, N4197, N1791, N2465);
and AND3 (N4224, N4220, N1517, N2642);
and AND3 (N4225, N4219, N3715, N1450);
and AND4 (N4226, N4223, N1216, N4025, N458);
and AND2 (N4227, N4222, N246);
and AND3 (N4228, N4224, N3644, N177);
or OR3 (N4229, N4200, N1941, N1335);
nand NAND4 (N4230, N4225, N2882, N423, N2048);
xor XOR2 (N4231, N4229, N453);
xor XOR2 (N4232, N4206, N2470);
buf BUF1 (N4233, N4228);
and AND2 (N4234, N4233, N801);
or OR3 (N4235, N4213, N2023, N3887);
nor NOR4 (N4236, N4217, N3619, N3531, N25);
nor NOR2 (N4237, N4234, N3338);
nand NAND2 (N4238, N4226, N3508);
buf BUF1 (N4239, N4232);
buf BUF1 (N4240, N4231);
and AND4 (N4241, N4240, N767, N1283, N1110);
xor XOR2 (N4242, N4195, N1744);
or OR2 (N4243, N4239, N2090);
nand NAND2 (N4244, N4238, N117);
nor NOR2 (N4245, N4242, N2650);
or OR4 (N4246, N4230, N1995, N1060, N1212);
not NOT1 (N4247, N4236);
buf BUF1 (N4248, N4237);
or OR4 (N4249, N4246, N3231, N801, N160);
not NOT1 (N4250, N4235);
not NOT1 (N4251, N4248);
buf BUF1 (N4252, N4251);
nand NAND4 (N4253, N4221, N3413, N3048, N2599);
and AND4 (N4254, N4227, N3599, N2488, N900);
not NOT1 (N4255, N4253);
nor NOR4 (N4256, N4247, N4008, N4129, N2773);
or OR4 (N4257, N4244, N3028, N710, N907);
xor XOR2 (N4258, N4252, N4139);
buf BUF1 (N4259, N4257);
not NOT1 (N4260, N4245);
not NOT1 (N4261, N4250);
not NOT1 (N4262, N4241);
or OR3 (N4263, N4254, N2321, N3235);
or OR2 (N4264, N4262, N2435);
nand NAND3 (N4265, N4260, N2784, N2205);
nand NAND2 (N4266, N4264, N3848);
buf BUF1 (N4267, N4243);
nor NOR4 (N4268, N4267, N889, N3862, N1210);
and AND2 (N4269, N4263, N756);
and AND2 (N4270, N4265, N353);
nand NAND4 (N4271, N4258, N1992, N961, N1830);
xor XOR2 (N4272, N4256, N1718);
not NOT1 (N4273, N4261);
or OR3 (N4274, N4249, N1952, N1355);
or OR2 (N4275, N4274, N150);
and AND3 (N4276, N4269, N290, N1761);
or OR2 (N4277, N4276, N1668);
not NOT1 (N4278, N4270);
nor NOR4 (N4279, N4272, N3798, N2416, N3401);
or OR3 (N4280, N4271, N2671, N973);
or OR2 (N4281, N4273, N330);
nor NOR3 (N4282, N4266, N3008, N3029);
and AND4 (N4283, N4275, N98, N1048, N513);
nor NOR2 (N4284, N4279, N4);
xor XOR2 (N4285, N4278, N2798);
not NOT1 (N4286, N4280);
or OR3 (N4287, N4283, N1506, N2559);
xor XOR2 (N4288, N4286, N3522);
or OR2 (N4289, N4277, N2134);
and AND4 (N4290, N4255, N1221, N1518, N1470);
and AND4 (N4291, N4259, N3107, N3964, N3112);
not NOT1 (N4292, N4288);
or OR2 (N4293, N4268, N524);
not NOT1 (N4294, N4291);
buf BUF1 (N4295, N4284);
or OR2 (N4296, N4287, N138);
buf BUF1 (N4297, N4281);
nor NOR4 (N4298, N4289, N2621, N2908, N2755);
and AND4 (N4299, N4292, N3638, N2925, N3078);
nor NOR2 (N4300, N4282, N1954);
nor NOR4 (N4301, N4299, N1956, N1806, N3751);
buf BUF1 (N4302, N4301);
and AND4 (N4303, N4302, N2009, N717, N1627);
nand NAND2 (N4304, N4303, N1264);
or OR3 (N4305, N4300, N3349, N4057);
and AND4 (N4306, N4304, N51, N392, N1015);
and AND3 (N4307, N4297, N2003, N1708);
nand NAND3 (N4308, N4305, N959, N901);
nor NOR2 (N4309, N4296, N3473);
nor NOR3 (N4310, N4295, N1539, N2400);
not NOT1 (N4311, N4307);
nor NOR4 (N4312, N4290, N2039, N1054, N339);
xor XOR2 (N4313, N4298, N2381);
nor NOR4 (N4314, N4312, N1674, N1713, N1199);
xor XOR2 (N4315, N4293, N2601);
and AND3 (N4316, N4311, N1071, N172);
and AND4 (N4317, N4285, N2326, N2621, N571);
xor XOR2 (N4318, N4310, N817);
and AND2 (N4319, N4314, N1111);
or OR2 (N4320, N4313, N1064);
buf BUF1 (N4321, N4294);
xor XOR2 (N4322, N4309, N3006);
buf BUF1 (N4323, N4306);
and AND3 (N4324, N4315, N2549, N15);
or OR4 (N4325, N4317, N29, N2463, N3515);
or OR2 (N4326, N4321, N2722);
and AND2 (N4327, N4319, N4050);
and AND3 (N4328, N4325, N1588, N4172);
not NOT1 (N4329, N4323);
buf BUF1 (N4330, N4329);
not NOT1 (N4331, N4328);
buf BUF1 (N4332, N4318);
not NOT1 (N4333, N4331);
xor XOR2 (N4334, N4308, N1922);
not NOT1 (N4335, N4327);
and AND2 (N4336, N4320, N2420);
xor XOR2 (N4337, N4332, N1780);
buf BUF1 (N4338, N4334);
not NOT1 (N4339, N4338);
nor NOR3 (N4340, N4337, N2343, N3646);
xor XOR2 (N4341, N4326, N1904);
buf BUF1 (N4342, N4316);
nand NAND2 (N4343, N4341, N3532);
and AND4 (N4344, N4343, N2062, N1527, N4070);
buf BUF1 (N4345, N4336);
xor XOR2 (N4346, N4330, N2909);
buf BUF1 (N4347, N4342);
buf BUF1 (N4348, N4322);
and AND4 (N4349, N4347, N450, N3365, N2157);
xor XOR2 (N4350, N4339, N193);
buf BUF1 (N4351, N4350);
not NOT1 (N4352, N4351);
or OR4 (N4353, N4349, N2447, N1184, N2659);
nand NAND2 (N4354, N4335, N3138);
not NOT1 (N4355, N4344);
or OR4 (N4356, N4348, N2226, N1024, N3635);
and AND3 (N4357, N4333, N290, N2985);
not NOT1 (N4358, N4355);
buf BUF1 (N4359, N4340);
buf BUF1 (N4360, N4359);
and AND3 (N4361, N4346, N2509, N1758);
not NOT1 (N4362, N4352);
not NOT1 (N4363, N4353);
or OR3 (N4364, N4362, N4130, N2157);
xor XOR2 (N4365, N4345, N3911);
and AND4 (N4366, N4356, N639, N3656, N1761);
and AND3 (N4367, N4366, N3981, N1314);
buf BUF1 (N4368, N4367);
buf BUF1 (N4369, N4365);
buf BUF1 (N4370, N4354);
buf BUF1 (N4371, N4363);
or OR4 (N4372, N4371, N4105, N208, N3353);
buf BUF1 (N4373, N4372);
nand NAND3 (N4374, N4364, N130, N632);
not NOT1 (N4375, N4360);
and AND2 (N4376, N4324, N1524);
xor XOR2 (N4377, N4357, N2484);
buf BUF1 (N4378, N4368);
nor NOR2 (N4379, N4376, N2591);
buf BUF1 (N4380, N4379);
nor NOR2 (N4381, N4373, N4343);
or OR2 (N4382, N4358, N4215);
buf BUF1 (N4383, N4377);
nor NOR4 (N4384, N4374, N3152, N615, N4195);
not NOT1 (N4385, N4381);
or OR4 (N4386, N4380, N1401, N366, N1120);
xor XOR2 (N4387, N4375, N939);
buf BUF1 (N4388, N4361);
or OR4 (N4389, N4385, N959, N742, N3995);
nor NOR2 (N4390, N4378, N244);
not NOT1 (N4391, N4370);
not NOT1 (N4392, N4387);
not NOT1 (N4393, N4392);
nor NOR3 (N4394, N4391, N2459, N1384);
and AND2 (N4395, N4369, N4273);
not NOT1 (N4396, N4386);
and AND2 (N4397, N4388, N3958);
or OR3 (N4398, N4395, N3529, N1180);
not NOT1 (N4399, N4383);
and AND2 (N4400, N4384, N1723);
and AND3 (N4401, N4390, N401, N4158);
buf BUF1 (N4402, N4397);
buf BUF1 (N4403, N4394);
not NOT1 (N4404, N4399);
nand NAND3 (N4405, N4396, N4335, N2384);
and AND4 (N4406, N4405, N2242, N43, N800);
xor XOR2 (N4407, N4382, N2849);
not NOT1 (N4408, N4398);
and AND4 (N4409, N4408, N657, N3837, N4044);
and AND2 (N4410, N4404, N482);
nor NOR3 (N4411, N4410, N4075, N382);
xor XOR2 (N4412, N4407, N3152);
or OR2 (N4413, N4393, N1148);
or OR3 (N4414, N4413, N3218, N744);
not NOT1 (N4415, N4400);
nor NOR2 (N4416, N4402, N3419);
buf BUF1 (N4417, N4406);
xor XOR2 (N4418, N4417, N4301);
not NOT1 (N4419, N4389);
not NOT1 (N4420, N4419);
nand NAND3 (N4421, N4411, N876, N3764);
or OR3 (N4422, N4414, N782, N1128);
not NOT1 (N4423, N4418);
and AND2 (N4424, N4412, N2114);
not NOT1 (N4425, N4424);
nand NAND3 (N4426, N4425, N2858, N1262);
and AND2 (N4427, N4401, N1171);
not NOT1 (N4428, N4409);
buf BUF1 (N4429, N4427);
xor XOR2 (N4430, N4428, N1982);
and AND3 (N4431, N4416, N390, N1353);
not NOT1 (N4432, N4429);
or OR4 (N4433, N4426, N1336, N1315, N1354);
nand NAND4 (N4434, N4422, N2438, N943, N3555);
nand NAND3 (N4435, N4434, N3322, N1834);
xor XOR2 (N4436, N4423, N4328);
not NOT1 (N4437, N4433);
not NOT1 (N4438, N4430);
or OR2 (N4439, N4431, N3717);
or OR4 (N4440, N4439, N602, N1477, N502);
nor NOR3 (N4441, N4403, N71, N3722);
xor XOR2 (N4442, N4421, N2823);
and AND4 (N4443, N4442, N2506, N1148, N99);
nor NOR2 (N4444, N4437, N511);
xor XOR2 (N4445, N4432, N215);
not NOT1 (N4446, N4444);
nor NOR3 (N4447, N4445, N3353, N3510);
or OR4 (N4448, N4415, N4053, N2704, N1956);
nor NOR3 (N4449, N4440, N3737, N3351);
nand NAND2 (N4450, N4443, N663);
or OR2 (N4451, N4420, N4372);
or OR2 (N4452, N4441, N1275);
or OR2 (N4453, N4449, N736);
and AND4 (N4454, N4451, N2088, N1946, N2854);
and AND3 (N4455, N4453, N4225, N757);
or OR3 (N4456, N4446, N2615, N4298);
nor NOR4 (N4457, N4438, N1743, N1755, N1927);
nand NAND3 (N4458, N4448, N607, N167);
buf BUF1 (N4459, N4447);
and AND3 (N4460, N4436, N350, N249);
buf BUF1 (N4461, N4459);
xor XOR2 (N4462, N4461, N3851);
buf BUF1 (N4463, N4455);
xor XOR2 (N4464, N4458, N3928);
not NOT1 (N4465, N4450);
and AND4 (N4466, N4464, N2822, N97, N3207);
and AND3 (N4467, N4460, N1118, N808);
nand NAND3 (N4468, N4467, N1475, N3466);
xor XOR2 (N4469, N4466, N1917);
or OR4 (N4470, N4469, N2424, N3722, N2100);
and AND2 (N4471, N4465, N1283);
or OR3 (N4472, N4454, N2833, N924);
not NOT1 (N4473, N4435);
not NOT1 (N4474, N4463);
not NOT1 (N4475, N4471);
nand NAND4 (N4476, N4468, N2629, N949, N1555);
not NOT1 (N4477, N4472);
and AND4 (N4478, N4452, N3005, N2931, N4438);
or OR3 (N4479, N4457, N878, N2467);
nand NAND4 (N4480, N4475, N3012, N3112, N131);
and AND2 (N4481, N4476, N776);
or OR3 (N4482, N4474, N3761, N2734);
xor XOR2 (N4483, N4478, N2520);
not NOT1 (N4484, N4480);
buf BUF1 (N4485, N4484);
xor XOR2 (N4486, N4456, N1914);
nand NAND3 (N4487, N4482, N1370, N1352);
xor XOR2 (N4488, N4477, N2444);
nor NOR3 (N4489, N4473, N1369, N1260);
or OR4 (N4490, N4487, N729, N4131, N1955);
buf BUF1 (N4491, N4485);
nor NOR4 (N4492, N4486, N3214, N2018, N2243);
buf BUF1 (N4493, N4491);
not NOT1 (N4494, N4481);
buf BUF1 (N4495, N4479);
or OR3 (N4496, N4492, N1949, N3992);
nand NAND2 (N4497, N4462, N1296);
nand NAND2 (N4498, N4497, N725);
not NOT1 (N4499, N4483);
xor XOR2 (N4500, N4495, N4477);
not NOT1 (N4501, N4496);
buf BUF1 (N4502, N4500);
buf BUF1 (N4503, N4493);
and AND4 (N4504, N4488, N3406, N1474, N1307);
or OR4 (N4505, N4501, N2438, N2738, N2927);
nand NAND4 (N4506, N4498, N4148, N2792, N977);
nor NOR3 (N4507, N4504, N1565, N2700);
and AND3 (N4508, N4507, N1438, N1981);
xor XOR2 (N4509, N4494, N3625);
xor XOR2 (N4510, N4489, N2387);
and AND4 (N4511, N4502, N96, N825, N1143);
not NOT1 (N4512, N4499);
and AND2 (N4513, N4508, N979);
nand NAND3 (N4514, N4506, N1372, N884);
or OR3 (N4515, N4510, N3745, N1138);
buf BUF1 (N4516, N4509);
or OR4 (N4517, N4514, N330, N1420, N2866);
not NOT1 (N4518, N4505);
nand NAND2 (N4519, N4518, N4161);
nor NOR2 (N4520, N4511, N1402);
and AND3 (N4521, N4470, N3754, N1299);
nor NOR2 (N4522, N4515, N1892);
or OR2 (N4523, N4503, N1517);
nor NOR2 (N4524, N4523, N3107);
nor NOR3 (N4525, N4520, N3991, N566);
nand NAND2 (N4526, N4522, N1340);
nand NAND3 (N4527, N4517, N1450, N4044);
xor XOR2 (N4528, N4519, N3456);
nand NAND4 (N4529, N4527, N1878, N1613, N1189);
or OR2 (N4530, N4525, N2368);
buf BUF1 (N4531, N4529);
nor NOR2 (N4532, N4526, N4224);
or OR2 (N4533, N4531, N2385);
and AND2 (N4534, N4512, N2669);
xor XOR2 (N4535, N4530, N3245);
nor NOR2 (N4536, N4534, N2255);
nand NAND3 (N4537, N4532, N333, N4379);
nand NAND2 (N4538, N4521, N2455);
or OR3 (N4539, N4516, N3784, N1380);
nor NOR2 (N4540, N4533, N1801);
xor XOR2 (N4541, N4538, N2508);
not NOT1 (N4542, N4540);
xor XOR2 (N4543, N4542, N2600);
buf BUF1 (N4544, N4539);
buf BUF1 (N4545, N4541);
xor XOR2 (N4546, N4537, N68);
nor NOR2 (N4547, N4546, N224);
xor XOR2 (N4548, N4528, N483);
or OR2 (N4549, N4547, N4517);
and AND4 (N4550, N4536, N3751, N4050, N3594);
nor NOR3 (N4551, N4490, N5, N3679);
nor NOR2 (N4552, N4524, N3061);
xor XOR2 (N4553, N4513, N864);
not NOT1 (N4554, N4543);
nor NOR2 (N4555, N4549, N4168);
not NOT1 (N4556, N4555);
nor NOR4 (N4557, N4548, N3238, N60, N1494);
not NOT1 (N4558, N4545);
nand NAND4 (N4559, N4550, N2694, N3317, N3307);
nand NAND2 (N4560, N4551, N3176);
not NOT1 (N4561, N4558);
buf BUF1 (N4562, N4554);
and AND3 (N4563, N4561, N2505, N3646);
and AND3 (N4564, N4535, N2582, N1009);
nand NAND3 (N4565, N4556, N789, N3191);
xor XOR2 (N4566, N4564, N2994);
nor NOR3 (N4567, N4563, N2000, N2874);
and AND2 (N4568, N4566, N3620);
buf BUF1 (N4569, N4562);
xor XOR2 (N4570, N4569, N2584);
or OR3 (N4571, N4565, N144, N559);
xor XOR2 (N4572, N4570, N3605);
or OR3 (N4573, N4544, N1280, N4566);
and AND2 (N4574, N4553, N3530);
xor XOR2 (N4575, N4552, N881);
xor XOR2 (N4576, N4560, N3458);
or OR2 (N4577, N4576, N2276);
nand NAND4 (N4578, N4574, N463, N2123, N1676);
or OR2 (N4579, N4557, N2004);
and AND4 (N4580, N4571, N2589, N933, N2015);
and AND3 (N4581, N4573, N1060, N1603);
and AND4 (N4582, N4567, N1264, N2946, N4485);
nor NOR2 (N4583, N4559, N1513);
xor XOR2 (N4584, N4580, N3639);
xor XOR2 (N4585, N4568, N3564);
or OR4 (N4586, N4584, N2031, N3209, N2052);
buf BUF1 (N4587, N4581);
nand NAND4 (N4588, N4583, N340, N2391, N1130);
nor NOR4 (N4589, N4586, N3545, N1988, N2913);
buf BUF1 (N4590, N4578);
nand NAND4 (N4591, N4577, N3362, N2491, N829);
xor XOR2 (N4592, N4587, N2231);
nand NAND3 (N4593, N4589, N782, N3092);
or OR2 (N4594, N4572, N3696);
xor XOR2 (N4595, N4575, N816);
nand NAND3 (N4596, N4591, N4337, N2262);
nor NOR3 (N4597, N4588, N1622, N2957);
and AND3 (N4598, N4592, N3416, N3325);
nand NAND3 (N4599, N4596, N3558, N3302);
nor NOR3 (N4600, N4579, N1429, N3427);
or OR3 (N4601, N4597, N3981, N3844);
and AND2 (N4602, N4600, N3858);
buf BUF1 (N4603, N4590);
nor NOR4 (N4604, N4595, N3454, N1726, N4071);
and AND4 (N4605, N4602, N3857, N2314, N4023);
buf BUF1 (N4606, N4599);
nand NAND4 (N4607, N4594, N3508, N321, N1287);
xor XOR2 (N4608, N4598, N3809);
nand NAND2 (N4609, N4603, N4091);
or OR4 (N4610, N4604, N2988, N2208, N3651);
not NOT1 (N4611, N4585);
nand NAND3 (N4612, N4610, N1948, N1155);
and AND3 (N4613, N4606, N2805, N2445);
xor XOR2 (N4614, N4611, N3015);
or OR4 (N4615, N4612, N306, N2457, N4551);
and AND2 (N4616, N4582, N3716);
nand NAND2 (N4617, N4613, N4334);
nor NOR4 (N4618, N4617, N30, N4007, N2757);
nand NAND2 (N4619, N4616, N41);
or OR4 (N4620, N4618, N1619, N1282, N730);
xor XOR2 (N4621, N4607, N1634);
or OR2 (N4622, N4601, N2641);
buf BUF1 (N4623, N4615);
buf BUF1 (N4624, N4620);
or OR2 (N4625, N4621, N1554);
xor XOR2 (N4626, N4608, N1470);
or OR3 (N4627, N4626, N3969, N1518);
or OR4 (N4628, N4622, N3895, N4530, N813);
not NOT1 (N4629, N4605);
or OR3 (N4630, N4627, N3989, N3641);
nor NOR2 (N4631, N4593, N2096);
not NOT1 (N4632, N4623);
not NOT1 (N4633, N4632);
nor NOR3 (N4634, N4614, N1829, N764);
or OR2 (N4635, N4628, N638);
or OR2 (N4636, N4633, N1648);
xor XOR2 (N4637, N4625, N1398);
and AND2 (N4638, N4634, N349);
nand NAND3 (N4639, N4624, N3823, N2538);
or OR2 (N4640, N4630, N1339);
nand NAND3 (N4641, N4629, N3604, N54);
and AND3 (N4642, N4639, N2343, N3535);
buf BUF1 (N4643, N4631);
or OR2 (N4644, N4637, N4552);
xor XOR2 (N4645, N4636, N747);
and AND4 (N4646, N4645, N599, N2844, N3247);
buf BUF1 (N4647, N4642);
or OR3 (N4648, N4641, N1013, N835);
xor XOR2 (N4649, N4609, N3835);
and AND2 (N4650, N4644, N4033);
buf BUF1 (N4651, N4647);
buf BUF1 (N4652, N4643);
nand NAND4 (N4653, N4638, N2844, N2296, N1658);
buf BUF1 (N4654, N4648);
nand NAND4 (N4655, N4635, N4267, N2232, N3441);
nand NAND2 (N4656, N4652, N2195);
nand NAND4 (N4657, N4653, N3196, N23, N4502);
nor NOR2 (N4658, N4656, N2000);
nor NOR2 (N4659, N4640, N3826);
xor XOR2 (N4660, N4651, N3588);
not NOT1 (N4661, N4659);
or OR3 (N4662, N4619, N1729, N339);
nor NOR4 (N4663, N4660, N795, N4569, N3126);
and AND2 (N4664, N4662, N4643);
buf BUF1 (N4665, N4663);
nor NOR3 (N4666, N4658, N4517, N355);
nor NOR2 (N4667, N4654, N4071);
nand NAND3 (N4668, N4650, N1740, N1252);
buf BUF1 (N4669, N4665);
nor NOR3 (N4670, N4668, N1371, N3140);
not NOT1 (N4671, N4664);
xor XOR2 (N4672, N4657, N3843);
nor NOR4 (N4673, N4649, N3884, N4375, N4030);
buf BUF1 (N4674, N4666);
not NOT1 (N4675, N4646);
nor NOR3 (N4676, N4661, N1392, N1658);
and AND3 (N4677, N4673, N2588, N4191);
not NOT1 (N4678, N4669);
or OR2 (N4679, N4672, N3236);
and AND4 (N4680, N4667, N139, N941, N245);
and AND2 (N4681, N4680, N4614);
or OR4 (N4682, N4670, N1710, N2140, N1059);
buf BUF1 (N4683, N4655);
nand NAND3 (N4684, N4682, N3538, N627);
nor NOR3 (N4685, N4677, N4337, N80);
and AND3 (N4686, N4675, N141, N4511);
buf BUF1 (N4687, N4683);
not NOT1 (N4688, N4679);
xor XOR2 (N4689, N4671, N3809);
not NOT1 (N4690, N4674);
not NOT1 (N4691, N4690);
nand NAND2 (N4692, N4678, N892);
xor XOR2 (N4693, N4686, N2785);
xor XOR2 (N4694, N4693, N2566);
not NOT1 (N4695, N4688);
nor NOR2 (N4696, N4676, N2376);
or OR2 (N4697, N4694, N1696);
nor NOR4 (N4698, N4687, N3801, N4544, N3733);
buf BUF1 (N4699, N4681);
xor XOR2 (N4700, N4685, N4347);
not NOT1 (N4701, N4697);
not NOT1 (N4702, N4691);
or OR4 (N4703, N4692, N1648, N4352, N3048);
not NOT1 (N4704, N4696);
xor XOR2 (N4705, N4684, N2791);
not NOT1 (N4706, N4698);
nand NAND3 (N4707, N4700, N1297, N3547);
and AND4 (N4708, N4689, N476, N3422, N4430);
or OR3 (N4709, N4701, N3179, N95);
buf BUF1 (N4710, N4699);
or OR3 (N4711, N4704, N4698, N486);
and AND4 (N4712, N4706, N2942, N2877, N1130);
buf BUF1 (N4713, N4707);
nor NOR3 (N4714, N4710, N3832, N1384);
buf BUF1 (N4715, N4705);
xor XOR2 (N4716, N4702, N2575);
xor XOR2 (N4717, N4695, N3541);
buf BUF1 (N4718, N4711);
not NOT1 (N4719, N4703);
nor NOR3 (N4720, N4714, N1161, N1872);
not NOT1 (N4721, N4708);
xor XOR2 (N4722, N4709, N3335);
buf BUF1 (N4723, N4712);
xor XOR2 (N4724, N4716, N143);
not NOT1 (N4725, N4715);
and AND4 (N4726, N4719, N2598, N1662, N4371);
buf BUF1 (N4727, N4725);
not NOT1 (N4728, N4718);
not NOT1 (N4729, N4726);
or OR3 (N4730, N4723, N843, N3216);
and AND4 (N4731, N4730, N3390, N3264, N1391);
nor NOR2 (N4732, N4731, N780);
xor XOR2 (N4733, N4717, N980);
nand NAND2 (N4734, N4732, N2120);
not NOT1 (N4735, N4733);
nor NOR2 (N4736, N4734, N3630);
and AND2 (N4737, N4713, N273);
nand NAND2 (N4738, N4729, N2064);
xor XOR2 (N4739, N4722, N2329);
buf BUF1 (N4740, N4739);
or OR4 (N4741, N4736, N2786, N247, N233);
or OR4 (N4742, N4728, N945, N4693, N2548);
or OR4 (N4743, N4724, N2443, N3584, N3211);
buf BUF1 (N4744, N4727);
nand NAND3 (N4745, N4741, N4220, N1341);
xor XOR2 (N4746, N4735, N1080);
and AND2 (N4747, N4745, N2939);
and AND4 (N4748, N4721, N3456, N938, N2632);
buf BUF1 (N4749, N4737);
and AND4 (N4750, N4746, N258, N2435, N1611);
not NOT1 (N4751, N4748);
nand NAND3 (N4752, N4744, N4192, N910);
nand NAND2 (N4753, N4747, N2976);
not NOT1 (N4754, N4738);
or OR3 (N4755, N4742, N2058, N3032);
buf BUF1 (N4756, N4755);
not NOT1 (N4757, N4751);
and AND4 (N4758, N4743, N2422, N3042, N4010);
not NOT1 (N4759, N4749);
nor NOR3 (N4760, N4757, N3608, N3764);
buf BUF1 (N4761, N4759);
xor XOR2 (N4762, N4758, N1004);
not NOT1 (N4763, N4754);
and AND3 (N4764, N4762, N1981, N4763);
buf BUF1 (N4765, N2881);
not NOT1 (N4766, N4761);
or OR3 (N4767, N4756, N648, N3586);
and AND2 (N4768, N4766, N842);
nor NOR2 (N4769, N4768, N1646);
nand NAND3 (N4770, N4720, N4275, N98);
not NOT1 (N4771, N4767);
nor NOR3 (N4772, N4770, N1780, N2798);
not NOT1 (N4773, N4740);
not NOT1 (N4774, N4753);
buf BUF1 (N4775, N4752);
nor NOR2 (N4776, N4773, N2578);
nand NAND3 (N4777, N4771, N2554, N4397);
buf BUF1 (N4778, N4764);
and AND2 (N4779, N4769, N3405);
not NOT1 (N4780, N4772);
nand NAND4 (N4781, N4775, N1286, N3297, N2445);
or OR2 (N4782, N4781, N1887);
or OR3 (N4783, N4760, N2482, N1341);
not NOT1 (N4784, N4779);
and AND2 (N4785, N4780, N435);
and AND3 (N4786, N4750, N2767, N3306);
and AND3 (N4787, N4782, N2863, N909);
or OR4 (N4788, N4778, N307, N137, N1060);
xor XOR2 (N4789, N4774, N367);
not NOT1 (N4790, N4765);
xor XOR2 (N4791, N4776, N4749);
xor XOR2 (N4792, N4790, N3066);
not NOT1 (N4793, N4789);
nand NAND3 (N4794, N4793, N651, N2963);
nor NOR2 (N4795, N4794, N2680);
buf BUF1 (N4796, N4795);
nor NOR3 (N4797, N4784, N1840, N4290);
and AND4 (N4798, N4796, N1180, N1362, N1670);
and AND2 (N4799, N4786, N519);
and AND3 (N4800, N4785, N1076, N4438);
not NOT1 (N4801, N4787);
nor NOR4 (N4802, N4799, N3105, N542, N3308);
xor XOR2 (N4803, N4797, N1701);
nand NAND4 (N4804, N4800, N2232, N2606, N4774);
nor NOR4 (N4805, N4788, N4779, N3360, N3015);
or OR4 (N4806, N4801, N1993, N3227, N467);
not NOT1 (N4807, N4792);
xor XOR2 (N4808, N4802, N2152);
or OR2 (N4809, N4805, N2801);
and AND4 (N4810, N4791, N2583, N3073, N624);
or OR2 (N4811, N4798, N3555);
not NOT1 (N4812, N4810);
xor XOR2 (N4813, N4804, N3520);
buf BUF1 (N4814, N4808);
nand NAND2 (N4815, N4812, N693);
not NOT1 (N4816, N4783);
nand NAND4 (N4817, N4814, N1125, N253, N2670);
and AND4 (N4818, N4777, N2912, N1102, N4585);
or OR4 (N4819, N4809, N1938, N4208, N4273);
buf BUF1 (N4820, N4811);
or OR3 (N4821, N4817, N791, N3410);
nor NOR2 (N4822, N4816, N1526);
not NOT1 (N4823, N4807);
nand NAND3 (N4824, N4818, N2586, N2351);
or OR4 (N4825, N4803, N4488, N452, N2576);
nor NOR3 (N4826, N4821, N602, N4006);
or OR2 (N4827, N4822, N699);
buf BUF1 (N4828, N4826);
not NOT1 (N4829, N4827);
buf BUF1 (N4830, N4828);
or OR3 (N4831, N4820, N4245, N4475);
buf BUF1 (N4832, N4825);
or OR4 (N4833, N4813, N1751, N4282, N315);
not NOT1 (N4834, N4831);
nor NOR4 (N4835, N4824, N1490, N4054, N4068);
nor NOR3 (N4836, N4819, N2897, N1774);
nor NOR4 (N4837, N4835, N547, N3139, N434);
buf BUF1 (N4838, N4836);
nand NAND4 (N4839, N4829, N4158, N3123, N2878);
or OR3 (N4840, N4830, N1986, N2087);
buf BUF1 (N4841, N4833);
nor NOR2 (N4842, N4834, N542);
buf BUF1 (N4843, N4840);
nor NOR3 (N4844, N4832, N2127, N2476);
not NOT1 (N4845, N4844);
buf BUF1 (N4846, N4842);
nor NOR3 (N4847, N4838, N3651, N1319);
or OR2 (N4848, N4815, N828);
xor XOR2 (N4849, N4839, N2769);
and AND4 (N4850, N4847, N4374, N4271, N1382);
buf BUF1 (N4851, N4848);
xor XOR2 (N4852, N4851, N3115);
nand NAND4 (N4853, N4806, N140, N2082, N2252);
or OR4 (N4854, N4850, N1267, N2311, N2846);
and AND2 (N4855, N4837, N318);
and AND3 (N4856, N4843, N1000, N2004);
or OR3 (N4857, N4845, N3639, N422);
nand NAND3 (N4858, N4852, N2436, N3597);
nor NOR2 (N4859, N4856, N2189);
and AND4 (N4860, N4855, N4602, N2109, N815);
xor XOR2 (N4861, N4857, N4049);
or OR4 (N4862, N4854, N1596, N2222, N435);
nor NOR4 (N4863, N4860, N954, N3382, N20);
buf BUF1 (N4864, N4862);
and AND2 (N4865, N4849, N1536);
not NOT1 (N4866, N4865);
nand NAND4 (N4867, N4823, N3334, N2734, N1655);
not NOT1 (N4868, N4864);
not NOT1 (N4869, N4868);
buf BUF1 (N4870, N4861);
nand NAND2 (N4871, N4867, N420);
and AND4 (N4872, N4859, N834, N2418, N2099);
buf BUF1 (N4873, N4863);
and AND2 (N4874, N4870, N136);
nor NOR4 (N4875, N4869, N4089, N1908, N4104);
nor NOR4 (N4876, N4874, N654, N1933, N1898);
buf BUF1 (N4877, N4841);
not NOT1 (N4878, N4876);
or OR2 (N4879, N4846, N1477);
xor XOR2 (N4880, N4878, N1664);
and AND4 (N4881, N4877, N4299, N2267, N2150);
nor NOR3 (N4882, N4866, N4795, N3622);
xor XOR2 (N4883, N4858, N3960);
buf BUF1 (N4884, N4871);
or OR3 (N4885, N4882, N3580, N3201);
nor NOR4 (N4886, N4883, N2641, N484, N1919);
nor NOR4 (N4887, N4885, N1689, N2804, N3989);
not NOT1 (N4888, N4853);
buf BUF1 (N4889, N4886);
xor XOR2 (N4890, N4879, N2307);
xor XOR2 (N4891, N4887, N4695);
nand NAND3 (N4892, N4884, N826, N3141);
xor XOR2 (N4893, N4891, N3484);
not NOT1 (N4894, N4888);
not NOT1 (N4895, N4890);
nand NAND3 (N4896, N4875, N553, N2129);
buf BUF1 (N4897, N4873);
not NOT1 (N4898, N4897);
nor NOR4 (N4899, N4894, N1967, N2449, N322);
not NOT1 (N4900, N4898);
buf BUF1 (N4901, N4881);
buf BUF1 (N4902, N4889);
or OR2 (N4903, N4900, N4506);
nor NOR4 (N4904, N4896, N3568, N1627, N3042);
nor NOR4 (N4905, N4892, N2362, N813, N4892);
buf BUF1 (N4906, N4899);
xor XOR2 (N4907, N4904, N1191);
and AND2 (N4908, N4872, N2076);
nor NOR2 (N4909, N4893, N390);
buf BUF1 (N4910, N4909);
nand NAND3 (N4911, N4906, N4819, N1444);
nand NAND4 (N4912, N4910, N3573, N3812, N1027);
not NOT1 (N4913, N4880);
nor NOR2 (N4914, N4912, N3033);
not NOT1 (N4915, N4902);
or OR3 (N4916, N4895, N3782, N381);
nand NAND2 (N4917, N4908, N506);
or OR2 (N4918, N4903, N2498);
nand NAND4 (N4919, N4907, N823, N2364, N1071);
and AND2 (N4920, N4916, N2186);
or OR3 (N4921, N4915, N455, N4231);
and AND4 (N4922, N4921, N69, N2293, N4089);
xor XOR2 (N4923, N4913, N3901);
not NOT1 (N4924, N4920);
or OR3 (N4925, N4911, N4584, N623);
and AND4 (N4926, N4919, N1802, N3491, N3528);
nand NAND2 (N4927, N4918, N1812);
nand NAND4 (N4928, N4926, N829, N1960, N47);
and AND4 (N4929, N4928, N140, N3849, N4436);
xor XOR2 (N4930, N4924, N2511);
xor XOR2 (N4931, N4914, N1998);
buf BUF1 (N4932, N4905);
nor NOR2 (N4933, N4932, N4075);
and AND3 (N4934, N4901, N1518, N2679);
buf BUF1 (N4935, N4922);
or OR2 (N4936, N4934, N3134);
xor XOR2 (N4937, N4923, N1567);
or OR2 (N4938, N4935, N2987);
and AND2 (N4939, N4930, N2425);
not NOT1 (N4940, N4917);
buf BUF1 (N4941, N4933);
nor NOR2 (N4942, N4931, N451);
nand NAND2 (N4943, N4925, N3699);
not NOT1 (N4944, N4927);
xor XOR2 (N4945, N4939, N3787);
nor NOR4 (N4946, N4936, N1033, N2502, N3176);
buf BUF1 (N4947, N4945);
buf BUF1 (N4948, N4944);
or OR2 (N4949, N4946, N3583);
xor XOR2 (N4950, N4949, N999);
nand NAND3 (N4951, N4929, N4209, N3503);
and AND4 (N4952, N4938, N3064, N2820, N378);
nor NOR2 (N4953, N4947, N3796);
nor NOR2 (N4954, N4952, N4123);
nand NAND3 (N4955, N4943, N3387, N4173);
buf BUF1 (N4956, N4948);
or OR3 (N4957, N4954, N883, N3459);
nor NOR3 (N4958, N4955, N1232, N2319);
or OR4 (N4959, N4950, N3514, N1593, N1915);
or OR4 (N4960, N4937, N1911, N4516, N1933);
nor NOR3 (N4961, N4957, N1127, N655);
or OR2 (N4962, N4941, N1806);
nor NOR2 (N4963, N4940, N3400);
not NOT1 (N4964, N4956);
or OR4 (N4965, N4963, N4862, N3289, N1976);
nand NAND2 (N4966, N4958, N840);
or OR2 (N4967, N4961, N3806);
or OR4 (N4968, N4965, N3030, N4628, N1166);
and AND2 (N4969, N4959, N2433);
or OR3 (N4970, N4953, N498, N4223);
nor NOR4 (N4971, N4962, N88, N237, N4308);
and AND4 (N4972, N4971, N4915, N3576, N2411);
nand NAND2 (N4973, N4970, N2253);
xor XOR2 (N4974, N4969, N2798);
nor NOR2 (N4975, N4942, N1544);
buf BUF1 (N4976, N4966);
and AND2 (N4977, N4960, N1081);
or OR3 (N4978, N4964, N3508, N85);
xor XOR2 (N4979, N4968, N2965);
nor NOR2 (N4980, N4976, N4387);
and AND2 (N4981, N4951, N3431);
not NOT1 (N4982, N4973);
xor XOR2 (N4983, N4981, N2368);
not NOT1 (N4984, N4974);
buf BUF1 (N4985, N4975);
buf BUF1 (N4986, N4977);
buf BUF1 (N4987, N4979);
not NOT1 (N4988, N4987);
not NOT1 (N4989, N4985);
and AND2 (N4990, N4978, N2939);
nor NOR2 (N4991, N4984, N3997);
and AND2 (N4992, N4982, N3721);
buf BUF1 (N4993, N4967);
buf BUF1 (N4994, N4989);
and AND3 (N4995, N4972, N1869, N1258);
buf BUF1 (N4996, N4986);
and AND2 (N4997, N4988, N10);
nand NAND3 (N4998, N4983, N1238, N3993);
buf BUF1 (N4999, N4997);
and AND2 (N5000, N4998, N1839);
nor NOR2 (N5001, N4996, N1781);
nor NOR4 (N5002, N4990, N1693, N810, N1063);
nand NAND2 (N5003, N5001, N3568);
not NOT1 (N5004, N4992);
or OR3 (N5005, N4999, N1146, N56);
nand NAND4 (N5006, N5000, N2759, N4729, N174);
or OR2 (N5007, N5005, N1829);
nor NOR2 (N5008, N5003, N4692);
buf BUF1 (N5009, N4993);
or OR2 (N5010, N5004, N3523);
buf BUF1 (N5011, N4980);
not NOT1 (N5012, N4991);
and AND3 (N5013, N5011, N3843, N3345);
and AND2 (N5014, N5012, N1604);
and AND3 (N5015, N5013, N858, N2630);
nand NAND4 (N5016, N4995, N1825, N4579, N4200);
nor NOR4 (N5017, N5009, N2543, N2571, N3809);
not NOT1 (N5018, N5008);
xor XOR2 (N5019, N5015, N4568);
not NOT1 (N5020, N5018);
xor XOR2 (N5021, N5016, N1631);
xor XOR2 (N5022, N5002, N2770);
not NOT1 (N5023, N5010);
not NOT1 (N5024, N5007);
not NOT1 (N5025, N5021);
or OR3 (N5026, N5014, N740, N2094);
nor NOR4 (N5027, N5025, N2615, N2364, N1107);
xor XOR2 (N5028, N5026, N4617);
xor XOR2 (N5029, N5028, N2696);
nor NOR2 (N5030, N5023, N4492);
nor NOR2 (N5031, N4994, N129);
nand NAND2 (N5032, N5027, N1439);
buf BUF1 (N5033, N5032);
buf BUF1 (N5034, N5031);
xor XOR2 (N5035, N5029, N2335);
nand NAND2 (N5036, N5020, N4117);
not NOT1 (N5037, N5006);
buf BUF1 (N5038, N5034);
buf BUF1 (N5039, N5036);
nand NAND3 (N5040, N5033, N2543, N2299);
nor NOR3 (N5041, N5038, N506, N1049);
or OR3 (N5042, N5024, N4164, N4391);
not NOT1 (N5043, N5035);
or OR2 (N5044, N5039, N718);
nor NOR2 (N5045, N5017, N2574);
nand NAND3 (N5046, N5022, N643, N2548);
nor NOR3 (N5047, N5045, N1877, N4361);
and AND3 (N5048, N5044, N354, N3358);
or OR2 (N5049, N5048, N4362);
nor NOR2 (N5050, N5047, N2468);
not NOT1 (N5051, N5030);
nand NAND4 (N5052, N5049, N4789, N942, N2892);
or OR4 (N5053, N5051, N4257, N198, N2162);
and AND4 (N5054, N5052, N3162, N1974, N2935);
and AND2 (N5055, N5019, N2168);
nor NOR3 (N5056, N5054, N4047, N3782);
or OR4 (N5057, N5055, N2723, N1103, N4239);
nand NAND4 (N5058, N5046, N2810, N400, N1801);
and AND3 (N5059, N5057, N3128, N4821);
and AND3 (N5060, N5043, N3528, N4685);
nor NOR4 (N5061, N5041, N2777, N1970, N1998);
nor NOR3 (N5062, N5061, N2658, N2189);
nand NAND2 (N5063, N5062, N4026);
or OR3 (N5064, N5040, N3610, N2656);
xor XOR2 (N5065, N5037, N2242);
not NOT1 (N5066, N5064);
nand NAND3 (N5067, N5056, N715, N248);
or OR2 (N5068, N5067, N4385);
and AND3 (N5069, N5066, N4983, N2012);
buf BUF1 (N5070, N5068);
buf BUF1 (N5071, N5065);
xor XOR2 (N5072, N5060, N1410);
nor NOR4 (N5073, N5053, N4604, N3180, N1800);
nand NAND3 (N5074, N5059, N3037, N1097);
buf BUF1 (N5075, N5074);
nand NAND2 (N5076, N5050, N3710);
nor NOR2 (N5077, N5063, N2265);
nand NAND4 (N5078, N5071, N1705, N1872, N2559);
and AND2 (N5079, N5058, N3571);
nor NOR3 (N5080, N5070, N3471, N2861);
and AND4 (N5081, N5079, N2943, N3513, N2764);
not NOT1 (N5082, N5076);
and AND3 (N5083, N5072, N2131, N3636);
nand NAND4 (N5084, N5077, N3606, N4460, N4205);
nor NOR3 (N5085, N5083, N1982, N3596);
or OR3 (N5086, N5082, N1075, N719);
nand NAND2 (N5087, N5042, N1333);
buf BUF1 (N5088, N5086);
or OR4 (N5089, N5073, N2534, N972, N4340);
buf BUF1 (N5090, N5087);
or OR4 (N5091, N5084, N3851, N3524, N3634);
xor XOR2 (N5092, N5080, N2566);
not NOT1 (N5093, N5069);
nor NOR2 (N5094, N5075, N1550);
xor XOR2 (N5095, N5094, N3845);
not NOT1 (N5096, N5091);
and AND2 (N5097, N5078, N755);
buf BUF1 (N5098, N5088);
nand NAND3 (N5099, N5085, N3211, N4755);
xor XOR2 (N5100, N5090, N2524);
not NOT1 (N5101, N5096);
xor XOR2 (N5102, N5098, N2752);
or OR3 (N5103, N5099, N3745, N1534);
not NOT1 (N5104, N5103);
nor NOR3 (N5105, N5097, N131, N932);
not NOT1 (N5106, N5081);
nor NOR4 (N5107, N5101, N2254, N3683, N1344);
buf BUF1 (N5108, N5089);
nor NOR3 (N5109, N5107, N2413, N1130);
nand NAND3 (N5110, N5109, N3774, N3221);
nor NOR4 (N5111, N5092, N1418, N1753, N2487);
buf BUF1 (N5112, N5111);
buf BUF1 (N5113, N5110);
xor XOR2 (N5114, N5113, N994);
buf BUF1 (N5115, N5100);
nor NOR2 (N5116, N5115, N1074);
buf BUF1 (N5117, N5112);
nand NAND3 (N5118, N5095, N1022, N3848);
and AND4 (N5119, N5106, N815, N2549, N2928);
nand NAND4 (N5120, N5108, N3781, N2960, N4375);
xor XOR2 (N5121, N5104, N3375);
or OR4 (N5122, N5120, N3052, N2213, N4521);
or OR2 (N5123, N5093, N4628);
not NOT1 (N5124, N5122);
and AND4 (N5125, N5114, N1839, N1968, N951);
not NOT1 (N5126, N5118);
nor NOR4 (N5127, N5124, N3501, N4560, N409);
xor XOR2 (N5128, N5126, N2868);
or OR4 (N5129, N5105, N2941, N3012, N339);
xor XOR2 (N5130, N5117, N1682);
not NOT1 (N5131, N5123);
nand NAND3 (N5132, N5128, N4683, N886);
buf BUF1 (N5133, N5129);
xor XOR2 (N5134, N5131, N143);
nand NAND2 (N5135, N5116, N907);
not NOT1 (N5136, N5121);
buf BUF1 (N5137, N5125);
or OR2 (N5138, N5127, N4916);
not NOT1 (N5139, N5102);
nor NOR3 (N5140, N5132, N2168, N4632);
xor XOR2 (N5141, N5137, N3378);
or OR2 (N5142, N5134, N1189);
or OR4 (N5143, N5138, N1092, N3033, N473);
not NOT1 (N5144, N5140);
not NOT1 (N5145, N5136);
nor NOR2 (N5146, N5139, N2936);
or OR4 (N5147, N5133, N1067, N4770, N2903);
and AND3 (N5148, N5144, N2276, N985);
nand NAND2 (N5149, N5146, N2227);
not NOT1 (N5150, N5149);
nor NOR3 (N5151, N5145, N2194, N4673);
nand NAND2 (N5152, N5135, N1386);
nand NAND4 (N5153, N5147, N4449, N1378, N5061);
and AND4 (N5154, N5142, N5110, N624, N2464);
not NOT1 (N5155, N5153);
and AND2 (N5156, N5151, N279);
nand NAND4 (N5157, N5148, N4, N4791, N1435);
nand NAND4 (N5158, N5157, N290, N195, N3856);
nor NOR2 (N5159, N5156, N119);
and AND3 (N5160, N5141, N2078, N3532);
and AND4 (N5161, N5159, N538, N227, N1507);
nand NAND2 (N5162, N5152, N2058);
nand NAND2 (N5163, N5154, N1777);
or OR4 (N5164, N5130, N26, N1782, N4304);
buf BUF1 (N5165, N5161);
and AND4 (N5166, N5150, N2751, N2564, N2533);
not NOT1 (N5167, N5163);
nor NOR3 (N5168, N5119, N3047, N4092);
not NOT1 (N5169, N5165);
buf BUF1 (N5170, N5162);
and AND4 (N5171, N5158, N2025, N4762, N3026);
nand NAND3 (N5172, N5171, N117, N2329);
and AND4 (N5173, N5143, N2362, N1404, N2140);
and AND2 (N5174, N5164, N1827);
not NOT1 (N5175, N5170);
and AND2 (N5176, N5155, N3557);
or OR3 (N5177, N5173, N1389, N3972);
buf BUF1 (N5178, N5168);
not NOT1 (N5179, N5178);
xor XOR2 (N5180, N5167, N4763);
not NOT1 (N5181, N5177);
nand NAND2 (N5182, N5180, N4382);
and AND4 (N5183, N5176, N3707, N2065, N1856);
buf BUF1 (N5184, N5182);
and AND3 (N5185, N5169, N966, N229);
nor NOR3 (N5186, N5181, N4276, N4371);
and AND3 (N5187, N5179, N4327, N1626);
and AND4 (N5188, N5183, N2720, N4732, N504);
or OR3 (N5189, N5184, N5102, N209);
nor NOR4 (N5190, N5174, N4426, N3745, N2794);
buf BUF1 (N5191, N5187);
nor NOR2 (N5192, N5189, N3050);
or OR2 (N5193, N5188, N277);
or OR4 (N5194, N5172, N1934, N3469, N2407);
buf BUF1 (N5195, N5192);
or OR2 (N5196, N5166, N1378);
buf BUF1 (N5197, N5191);
buf BUF1 (N5198, N5175);
buf BUF1 (N5199, N5186);
nand NAND4 (N5200, N5198, N3674, N188, N4907);
or OR4 (N5201, N5194, N4580, N1910, N4040);
or OR3 (N5202, N5185, N304, N770);
nor NOR3 (N5203, N5193, N3511, N5019);
not NOT1 (N5204, N5202);
not NOT1 (N5205, N5190);
not NOT1 (N5206, N5203);
xor XOR2 (N5207, N5206, N2814);
buf BUF1 (N5208, N5201);
and AND2 (N5209, N5204, N3471);
nor NOR3 (N5210, N5199, N5092, N3389);
nand NAND4 (N5211, N5200, N2735, N4263, N5006);
and AND4 (N5212, N5208, N632, N2525, N2535);
not NOT1 (N5213, N5209);
nand NAND4 (N5214, N5210, N3597, N1841, N2538);
nand NAND4 (N5215, N5214, N3403, N346, N4883);
nand NAND4 (N5216, N5205, N817, N4485, N210);
xor XOR2 (N5217, N5160, N2622);
and AND3 (N5218, N5215, N276, N1831);
not NOT1 (N5219, N5195);
nor NOR4 (N5220, N5218, N4953, N326, N942);
nand NAND3 (N5221, N5207, N4948, N3370);
nand NAND3 (N5222, N5213, N4220, N222);
nor NOR2 (N5223, N5212, N3286);
xor XOR2 (N5224, N5211, N1429);
xor XOR2 (N5225, N5224, N835);
nor NOR4 (N5226, N5220, N953, N201, N2232);
or OR2 (N5227, N5221, N1304);
nand NAND3 (N5228, N5217, N159, N2237);
or OR4 (N5229, N5225, N2300, N3811, N1010);
not NOT1 (N5230, N5226);
not NOT1 (N5231, N5197);
xor XOR2 (N5232, N5227, N4805);
or OR3 (N5233, N5216, N2614, N2161);
buf BUF1 (N5234, N5219);
buf BUF1 (N5235, N5234);
nor NOR2 (N5236, N5228, N3249);
nor NOR2 (N5237, N5229, N4648);
not NOT1 (N5238, N5231);
and AND3 (N5239, N5237, N2266, N4889);
or OR3 (N5240, N5238, N4987, N4837);
or OR4 (N5241, N5222, N3499, N3270, N1069);
or OR4 (N5242, N5239, N3773, N3291, N4124);
not NOT1 (N5243, N5230);
buf BUF1 (N5244, N5236);
xor XOR2 (N5245, N5196, N4113);
xor XOR2 (N5246, N5245, N1916);
not NOT1 (N5247, N5243);
not NOT1 (N5248, N5232);
not NOT1 (N5249, N5223);
buf BUF1 (N5250, N5248);
buf BUF1 (N5251, N5250);
not NOT1 (N5252, N5251);
nand NAND4 (N5253, N5241, N1838, N3543, N2204);
buf BUF1 (N5254, N5240);
or OR2 (N5255, N5249, N4705);
or OR2 (N5256, N5235, N1686);
and AND3 (N5257, N5246, N96, N4408);
and AND4 (N5258, N5244, N689, N2066, N756);
or OR3 (N5259, N5254, N4349, N3593);
nand NAND2 (N5260, N5252, N4115);
and AND2 (N5261, N5247, N3834);
not NOT1 (N5262, N5233);
nand NAND3 (N5263, N5257, N2141, N1927);
not NOT1 (N5264, N5261);
and AND2 (N5265, N5262, N1640);
or OR3 (N5266, N5263, N4832, N2050);
not NOT1 (N5267, N5264);
and AND4 (N5268, N5265, N1725, N2412, N4720);
buf BUF1 (N5269, N5260);
or OR2 (N5270, N5256, N4704);
and AND3 (N5271, N5270, N2141, N4052);
xor XOR2 (N5272, N5266, N4958);
nand NAND4 (N5273, N5269, N2731, N4646, N2297);
and AND4 (N5274, N5271, N919, N1160, N3538);
xor XOR2 (N5275, N5242, N235);
nand NAND2 (N5276, N5253, N4999);
nand NAND2 (N5277, N5276, N454);
and AND3 (N5278, N5272, N3717, N359);
or OR3 (N5279, N5278, N3960, N826);
xor XOR2 (N5280, N5273, N580);
buf BUF1 (N5281, N5259);
and AND2 (N5282, N5280, N2313);
and AND4 (N5283, N5281, N5220, N4792, N1581);
buf BUF1 (N5284, N5283);
buf BUF1 (N5285, N5282);
and AND2 (N5286, N5277, N3056);
nor NOR2 (N5287, N5275, N1197);
nor NOR4 (N5288, N5284, N5002, N1801, N4175);
not NOT1 (N5289, N5286);
and AND4 (N5290, N5258, N2689, N2365, N4729);
nand NAND3 (N5291, N5267, N3722, N4688);
nand NAND2 (N5292, N5279, N891);
xor XOR2 (N5293, N5285, N4174);
nand NAND2 (N5294, N5292, N2778);
buf BUF1 (N5295, N5294);
not NOT1 (N5296, N5290);
or OR2 (N5297, N5288, N661);
nor NOR3 (N5298, N5296, N4127, N1637);
or OR3 (N5299, N5255, N1985, N792);
nand NAND3 (N5300, N5299, N1376, N3160);
nand NAND4 (N5301, N5297, N3189, N3360, N3705);
nand NAND3 (N5302, N5301, N253, N1517);
nor NOR2 (N5303, N5298, N2874);
nor NOR3 (N5304, N5274, N4931, N350);
nor NOR3 (N5305, N5287, N2064, N2618);
and AND2 (N5306, N5295, N1818);
not NOT1 (N5307, N5305);
buf BUF1 (N5308, N5306);
nor NOR2 (N5309, N5307, N4942);
buf BUF1 (N5310, N5304);
xor XOR2 (N5311, N5308, N2994);
buf BUF1 (N5312, N5303);
buf BUF1 (N5313, N5311);
or OR3 (N5314, N5302, N3930, N559);
nor NOR3 (N5315, N5309, N4986, N2491);
buf BUF1 (N5316, N5268);
buf BUF1 (N5317, N5289);
and AND3 (N5318, N5313, N1002, N3427);
nand NAND2 (N5319, N5310, N1504);
and AND2 (N5320, N5293, N4660);
or OR2 (N5321, N5300, N447);
buf BUF1 (N5322, N5314);
nor NOR4 (N5323, N5318, N5117, N4958, N4184);
and AND4 (N5324, N5322, N5025, N1828, N2373);
or OR2 (N5325, N5321, N2908);
and AND2 (N5326, N5312, N4583);
nand NAND2 (N5327, N5315, N4984);
and AND2 (N5328, N5326, N1555);
not NOT1 (N5329, N5324);
buf BUF1 (N5330, N5291);
buf BUF1 (N5331, N5325);
buf BUF1 (N5332, N5316);
nor NOR3 (N5333, N5317, N3896, N3551);
not NOT1 (N5334, N5331);
xor XOR2 (N5335, N5320, N1131);
not NOT1 (N5336, N5319);
nand NAND4 (N5337, N5328, N4519, N5194, N1441);
nor NOR4 (N5338, N5334, N3846, N1352, N1898);
xor XOR2 (N5339, N5333, N1152);
nor NOR3 (N5340, N5329, N3513, N1661);
not NOT1 (N5341, N5335);
nor NOR3 (N5342, N5323, N4659, N5214);
not NOT1 (N5343, N5340);
nor NOR4 (N5344, N5343, N1298, N2805, N709);
xor XOR2 (N5345, N5339, N1838);
nand NAND2 (N5346, N5337, N2377);
not NOT1 (N5347, N5332);
or OR3 (N5348, N5327, N5293, N5182);
buf BUF1 (N5349, N5342);
or OR2 (N5350, N5349, N3308);
or OR3 (N5351, N5336, N3160, N4486);
buf BUF1 (N5352, N5347);
nand NAND2 (N5353, N5338, N35);
buf BUF1 (N5354, N5350);
nand NAND3 (N5355, N5344, N1049, N1826);
or OR3 (N5356, N5353, N4156, N2602);
nand NAND3 (N5357, N5355, N2968, N2933);
or OR2 (N5358, N5351, N4570);
nor NOR3 (N5359, N5348, N835, N2516);
buf BUF1 (N5360, N5358);
nand NAND3 (N5361, N5352, N2463, N3728);
not NOT1 (N5362, N5360);
and AND4 (N5363, N5357, N5184, N4163, N1648);
xor XOR2 (N5364, N5354, N5120);
buf BUF1 (N5365, N5330);
buf BUF1 (N5366, N5359);
not NOT1 (N5367, N5365);
nor NOR3 (N5368, N5366, N1936, N3233);
not NOT1 (N5369, N5364);
buf BUF1 (N5370, N5345);
buf BUF1 (N5371, N5370);
and AND2 (N5372, N5368, N5065);
or OR2 (N5373, N5356, N2691);
or OR4 (N5374, N5363, N394, N188, N4688);
nand NAND2 (N5375, N5371, N2062);
or OR3 (N5376, N5362, N2567, N779);
or OR2 (N5377, N5369, N1745);
and AND4 (N5378, N5361, N3808, N708, N2546);
nand NAND2 (N5379, N5378, N3204);
nor NOR3 (N5380, N5367, N4915, N1494);
or OR4 (N5381, N5374, N3779, N3363, N2208);
not NOT1 (N5382, N5375);
and AND3 (N5383, N5376, N2008, N1928);
nor NOR3 (N5384, N5382, N2238, N4824);
nor NOR3 (N5385, N5346, N4360, N123);
nor NOR4 (N5386, N5341, N5108, N3437, N1836);
or OR3 (N5387, N5372, N551, N4578);
xor XOR2 (N5388, N5387, N301);
nor NOR2 (N5389, N5384, N4871);
not NOT1 (N5390, N5373);
nor NOR2 (N5391, N5383, N1638);
or OR2 (N5392, N5390, N941);
nand NAND3 (N5393, N5386, N2908, N4154);
buf BUF1 (N5394, N5388);
and AND4 (N5395, N5381, N5227, N175, N928);
or OR3 (N5396, N5385, N4052, N4486);
buf BUF1 (N5397, N5392);
xor XOR2 (N5398, N5397, N1118);
buf BUF1 (N5399, N5380);
not NOT1 (N5400, N5395);
nor NOR3 (N5401, N5400, N1036, N1958);
not NOT1 (N5402, N5399);
and AND3 (N5403, N5401, N529, N175);
or OR2 (N5404, N5403, N4704);
xor XOR2 (N5405, N5404, N321);
nor NOR4 (N5406, N5391, N3892, N3232, N3802);
and AND2 (N5407, N5396, N344);
buf BUF1 (N5408, N5377);
nor NOR2 (N5409, N5393, N2734);
xor XOR2 (N5410, N5406, N3425);
xor XOR2 (N5411, N5409, N3347);
nor NOR4 (N5412, N5408, N4316, N3772, N5036);
and AND3 (N5413, N5405, N3484, N119);
xor XOR2 (N5414, N5379, N2727);
xor XOR2 (N5415, N5402, N1824);
nand NAND4 (N5416, N5415, N3808, N4856, N5172);
or OR4 (N5417, N5407, N5029, N2229, N2746);
and AND4 (N5418, N5389, N4513, N1678, N1416);
buf BUF1 (N5419, N5413);
not NOT1 (N5420, N5418);
and AND4 (N5421, N5410, N2603, N831, N2959);
xor XOR2 (N5422, N5414, N704);
and AND3 (N5423, N5419, N3764, N2566);
not NOT1 (N5424, N5422);
not NOT1 (N5425, N5411);
nand NAND2 (N5426, N5416, N5416);
buf BUF1 (N5427, N5412);
not NOT1 (N5428, N5423);
xor XOR2 (N5429, N5421, N2422);
nor NOR4 (N5430, N5428, N1164, N565, N4919);
or OR4 (N5431, N5417, N1451, N3133, N514);
nor NOR4 (N5432, N5425, N2934, N1141, N1599);
and AND4 (N5433, N5429, N4762, N2409, N2327);
not NOT1 (N5434, N5432);
buf BUF1 (N5435, N5398);
buf BUF1 (N5436, N5431);
nor NOR3 (N5437, N5433, N3389, N1555);
nand NAND3 (N5438, N5424, N3309, N944);
or OR4 (N5439, N5430, N1726, N3792, N4652);
and AND4 (N5440, N5420, N5144, N3699, N5134);
buf BUF1 (N5441, N5434);
or OR4 (N5442, N5426, N1003, N5359, N1862);
nor NOR3 (N5443, N5442, N4529, N1316);
xor XOR2 (N5444, N5427, N4514);
nor NOR4 (N5445, N5437, N3295, N3491, N2270);
and AND4 (N5446, N5440, N39, N5350, N4972);
xor XOR2 (N5447, N5394, N2807);
or OR3 (N5448, N5435, N4562, N892);
xor XOR2 (N5449, N5439, N2728);
or OR3 (N5450, N5444, N1862, N5056);
not NOT1 (N5451, N5436);
buf BUF1 (N5452, N5443);
or OR3 (N5453, N5446, N942, N4799);
or OR4 (N5454, N5450, N3412, N5360, N4439);
nand NAND2 (N5455, N5451, N1917);
buf BUF1 (N5456, N5453);
buf BUF1 (N5457, N5452);
xor XOR2 (N5458, N5448, N5044);
xor XOR2 (N5459, N5447, N2577);
or OR3 (N5460, N5458, N2076, N2845);
nor NOR3 (N5461, N5460, N3222, N5278);
nor NOR3 (N5462, N5461, N985, N1144);
nand NAND3 (N5463, N5457, N3293, N5086);
not NOT1 (N5464, N5438);
nor NOR2 (N5465, N5459, N4608);
buf BUF1 (N5466, N5449);
buf BUF1 (N5467, N5454);
nand NAND4 (N5468, N5441, N1200, N3351, N5191);
or OR4 (N5469, N5455, N2305, N5158, N3406);
xor XOR2 (N5470, N5467, N4216);
buf BUF1 (N5471, N5466);
not NOT1 (N5472, N5468);
and AND4 (N5473, N5456, N977, N148, N2695);
nor NOR3 (N5474, N5473, N2458, N2804);
buf BUF1 (N5475, N5470);
nand NAND2 (N5476, N5463, N3474);
xor XOR2 (N5477, N5469, N552);
nor NOR2 (N5478, N5471, N4927);
buf BUF1 (N5479, N5445);
and AND2 (N5480, N5472, N3469);
not NOT1 (N5481, N5475);
xor XOR2 (N5482, N5478, N4136);
not NOT1 (N5483, N5479);
or OR3 (N5484, N5465, N2093, N2729);
nand NAND2 (N5485, N5482, N3942);
nor NOR4 (N5486, N5476, N5442, N1887, N3536);
not NOT1 (N5487, N5462);
buf BUF1 (N5488, N5487);
nand NAND3 (N5489, N5477, N52, N3185);
buf BUF1 (N5490, N5486);
buf BUF1 (N5491, N5490);
and AND3 (N5492, N5464, N452, N951);
nand NAND2 (N5493, N5489, N4457);
and AND4 (N5494, N5483, N380, N5346, N1494);
not NOT1 (N5495, N5488);
not NOT1 (N5496, N5485);
nor NOR2 (N5497, N5481, N2153);
buf BUF1 (N5498, N5474);
and AND4 (N5499, N5496, N2165, N460, N3620);
nor NOR2 (N5500, N5498, N4502);
buf BUF1 (N5501, N5497);
xor XOR2 (N5502, N5501, N4910);
or OR3 (N5503, N5502, N2962, N448);
xor XOR2 (N5504, N5503, N4957);
xor XOR2 (N5505, N5494, N1030);
and AND3 (N5506, N5493, N1682, N1518);
buf BUF1 (N5507, N5484);
or OR4 (N5508, N5480, N8, N1202, N4692);
or OR3 (N5509, N5505, N3796, N3597);
buf BUF1 (N5510, N5495);
xor XOR2 (N5511, N5504, N1541);
nand NAND2 (N5512, N5507, N2241);
not NOT1 (N5513, N5491);
nand NAND4 (N5514, N5506, N2145, N177, N1115);
xor XOR2 (N5515, N5500, N3561);
or OR4 (N5516, N5512, N31, N4537, N1048);
not NOT1 (N5517, N5509);
and AND4 (N5518, N5514, N1103, N5345, N2807);
or OR4 (N5519, N5517, N3493, N253, N2239);
not NOT1 (N5520, N5515);
not NOT1 (N5521, N5513);
nand NAND2 (N5522, N5518, N5256);
nand NAND3 (N5523, N5508, N585, N1346);
and AND2 (N5524, N5521, N1283);
nand NAND2 (N5525, N5516, N2077);
xor XOR2 (N5526, N5510, N4442);
nor NOR3 (N5527, N5525, N3737, N1968);
not NOT1 (N5528, N5522);
buf BUF1 (N5529, N5527);
xor XOR2 (N5530, N5528, N3515);
buf BUF1 (N5531, N5499);
nor NOR2 (N5532, N5529, N5035);
nor NOR3 (N5533, N5531, N3912, N1608);
nor NOR4 (N5534, N5492, N893, N1429, N284);
buf BUF1 (N5535, N5534);
and AND4 (N5536, N5520, N1444, N2050, N4289);
xor XOR2 (N5537, N5532, N537);
or OR4 (N5538, N5526, N4542, N2078, N4534);
xor XOR2 (N5539, N5523, N1374);
nor NOR4 (N5540, N5536, N5298, N1758, N3285);
nor NOR2 (N5541, N5519, N3968);
nor NOR3 (N5542, N5533, N3796, N299);
not NOT1 (N5543, N5542);
not NOT1 (N5544, N5535);
not NOT1 (N5545, N5530);
and AND4 (N5546, N5539, N928, N3811, N3897);
nor NOR2 (N5547, N5544, N872);
nand NAND2 (N5548, N5540, N3417);
and AND4 (N5549, N5547, N2711, N4913, N3972);
nand NAND4 (N5550, N5545, N3850, N91, N3425);
buf BUF1 (N5551, N5546);
buf BUF1 (N5552, N5538);
nor NOR2 (N5553, N5541, N3619);
buf BUF1 (N5554, N5551);
not NOT1 (N5555, N5537);
xor XOR2 (N5556, N5552, N5413);
not NOT1 (N5557, N5556);
and AND4 (N5558, N5549, N4073, N1243, N1181);
nand NAND3 (N5559, N5557, N5181, N1856);
not NOT1 (N5560, N5555);
nand NAND4 (N5561, N5511, N4513, N4536, N4392);
nor NOR3 (N5562, N5560, N3492, N2294);
nor NOR2 (N5563, N5553, N4596);
nand NAND4 (N5564, N5554, N2619, N1369, N1353);
not NOT1 (N5565, N5558);
or OR4 (N5566, N5559, N3269, N1852, N3816);
nand NAND4 (N5567, N5561, N997, N2820, N3094);
or OR4 (N5568, N5567, N1397, N895, N4981);
or OR2 (N5569, N5543, N2402);
xor XOR2 (N5570, N5568, N1771);
nor NOR4 (N5571, N5524, N3763, N4232, N3738);
not NOT1 (N5572, N5564);
buf BUF1 (N5573, N5569);
buf BUF1 (N5574, N5563);
xor XOR2 (N5575, N5574, N5390);
xor XOR2 (N5576, N5548, N4323);
or OR4 (N5577, N5575, N4435, N2492, N2659);
nand NAND4 (N5578, N5573, N4790, N2591, N4657);
and AND2 (N5579, N5572, N2822);
nand NAND2 (N5580, N5579, N3121);
and AND4 (N5581, N5570, N3667, N519, N5514);
not NOT1 (N5582, N5580);
and AND2 (N5583, N5566, N1);
not NOT1 (N5584, N5577);
not NOT1 (N5585, N5581);
buf BUF1 (N5586, N5578);
not NOT1 (N5587, N5550);
buf BUF1 (N5588, N5587);
and AND3 (N5589, N5588, N4296, N3714);
and AND4 (N5590, N5571, N4934, N1688, N4791);
nor NOR4 (N5591, N5590, N4173, N5355, N3787);
not NOT1 (N5592, N5584);
or OR3 (N5593, N5582, N4707, N926);
nor NOR2 (N5594, N5589, N3458);
or OR2 (N5595, N5592, N1406);
not NOT1 (N5596, N5595);
or OR3 (N5597, N5594, N3022, N2933);
nand NAND2 (N5598, N5585, N782);
or OR4 (N5599, N5562, N5348, N5111, N2339);
nor NOR2 (N5600, N5591, N403);
and AND2 (N5601, N5565, N3659);
buf BUF1 (N5602, N5593);
and AND4 (N5603, N5583, N4522, N4139, N3);
and AND4 (N5604, N5586, N1639, N4640, N2571);
or OR4 (N5605, N5597, N766, N1762, N835);
xor XOR2 (N5606, N5598, N5299);
or OR2 (N5607, N5600, N2342);
or OR4 (N5608, N5599, N3552, N4442, N247);
buf BUF1 (N5609, N5606);
or OR2 (N5610, N5576, N817);
xor XOR2 (N5611, N5596, N1829);
xor XOR2 (N5612, N5602, N3979);
nand NAND3 (N5613, N5608, N1767, N1155);
nand NAND4 (N5614, N5611, N5174, N4568, N178);
nand NAND3 (N5615, N5609, N4009, N1102);
or OR2 (N5616, N5605, N358);
nor NOR4 (N5617, N5603, N408, N3472, N3593);
or OR3 (N5618, N5604, N2077, N1995);
xor XOR2 (N5619, N5614, N398);
not NOT1 (N5620, N5613);
and AND4 (N5621, N5616, N4538, N1881, N4383);
buf BUF1 (N5622, N5621);
not NOT1 (N5623, N5610);
not NOT1 (N5624, N5619);
and AND2 (N5625, N5623, N3059);
nor NOR4 (N5626, N5607, N756, N4958, N944);
xor XOR2 (N5627, N5625, N5268);
buf BUF1 (N5628, N5618);
nand NAND3 (N5629, N5624, N1158, N4715);
and AND3 (N5630, N5629, N2202, N2708);
buf BUF1 (N5631, N5626);
buf BUF1 (N5632, N5622);
xor XOR2 (N5633, N5627, N1566);
nor NOR4 (N5634, N5615, N4427, N3680, N4875);
buf BUF1 (N5635, N5617);
not NOT1 (N5636, N5601);
nand NAND2 (N5637, N5634, N1702);
xor XOR2 (N5638, N5630, N2761);
nor NOR4 (N5639, N5633, N73, N745, N3178);
buf BUF1 (N5640, N5638);
or OR4 (N5641, N5635, N5602, N2829, N3716);
buf BUF1 (N5642, N5620);
or OR4 (N5643, N5631, N5056, N963, N2066);
and AND3 (N5644, N5640, N4454, N4963);
or OR3 (N5645, N5628, N3552, N2857);
and AND4 (N5646, N5636, N1469, N3410, N981);
nor NOR2 (N5647, N5632, N4587);
nand NAND3 (N5648, N5642, N3432, N434);
xor XOR2 (N5649, N5641, N3129);
buf BUF1 (N5650, N5648);
not NOT1 (N5651, N5649);
nor NOR2 (N5652, N5644, N3119);
and AND2 (N5653, N5647, N529);
nor NOR3 (N5654, N5639, N2433, N612);
or OR2 (N5655, N5650, N3418);
and AND2 (N5656, N5655, N4227);
not NOT1 (N5657, N5654);
xor XOR2 (N5658, N5657, N5246);
nor NOR4 (N5659, N5637, N1257, N3322, N3626);
and AND2 (N5660, N5656, N5216);
nor NOR3 (N5661, N5645, N2620, N1900);
nand NAND3 (N5662, N5661, N102, N248);
xor XOR2 (N5663, N5651, N4311);
buf BUF1 (N5664, N5612);
buf BUF1 (N5665, N5664);
buf BUF1 (N5666, N5663);
nand NAND2 (N5667, N5659, N2588);
and AND3 (N5668, N5667, N2507, N3575);
and AND2 (N5669, N5662, N2562);
nor NOR2 (N5670, N5660, N4034);
xor XOR2 (N5671, N5670, N1046);
nor NOR4 (N5672, N5669, N5484, N5290, N409);
buf BUF1 (N5673, N5646);
nand NAND2 (N5674, N5665, N1320);
or OR4 (N5675, N5668, N3163, N1135, N3042);
not NOT1 (N5676, N5643);
buf BUF1 (N5677, N5666);
not NOT1 (N5678, N5652);
and AND4 (N5679, N5672, N1348, N2055, N2827);
xor XOR2 (N5680, N5678, N400);
and AND2 (N5681, N5680, N1433);
nor NOR4 (N5682, N5675, N5314, N119, N4155);
or OR4 (N5683, N5658, N406, N3421, N1752);
or OR2 (N5684, N5681, N1542);
or OR3 (N5685, N5674, N5053, N3121);
buf BUF1 (N5686, N5676);
and AND4 (N5687, N5673, N2815, N560, N5376);
buf BUF1 (N5688, N5685);
not NOT1 (N5689, N5684);
or OR4 (N5690, N5689, N5667, N2039, N3726);
buf BUF1 (N5691, N5688);
nand NAND3 (N5692, N5679, N3152, N2775);
nor NOR3 (N5693, N5671, N524, N5298);
nor NOR2 (N5694, N5693, N3671);
and AND2 (N5695, N5690, N3969);
and AND2 (N5696, N5682, N1964);
not NOT1 (N5697, N5653);
and AND3 (N5698, N5696, N2488, N3977);
not NOT1 (N5699, N5686);
buf BUF1 (N5700, N5698);
and AND3 (N5701, N5697, N5330, N674);
not NOT1 (N5702, N5687);
nor NOR3 (N5703, N5677, N963, N3465);
nand NAND4 (N5704, N5695, N3839, N569, N4186);
and AND4 (N5705, N5699, N587, N5600, N2746);
nor NOR4 (N5706, N5692, N3118, N4849, N5324);
and AND4 (N5707, N5703, N1885, N4419, N1881);
nor NOR4 (N5708, N5702, N4936, N2895, N2445);
not NOT1 (N5709, N5706);
and AND4 (N5710, N5691, N2246, N1409, N705);
xor XOR2 (N5711, N5700, N4919);
and AND3 (N5712, N5694, N5103, N4631);
buf BUF1 (N5713, N5708);
nand NAND4 (N5714, N5711, N1904, N2882, N1530);
or OR2 (N5715, N5712, N341);
xor XOR2 (N5716, N5713, N3828);
nor NOR4 (N5717, N5701, N1511, N4189, N1875);
or OR2 (N5718, N5707, N1427);
buf BUF1 (N5719, N5710);
or OR3 (N5720, N5683, N4294, N185);
nand NAND4 (N5721, N5714, N3733, N1829, N1011);
buf BUF1 (N5722, N5720);
and AND2 (N5723, N5716, N1388);
xor XOR2 (N5724, N5718, N3034);
xor XOR2 (N5725, N5724, N1175);
nand NAND3 (N5726, N5709, N5375, N4603);
or OR4 (N5727, N5723, N2837, N4174, N3800);
nand NAND2 (N5728, N5705, N5654);
xor XOR2 (N5729, N5725, N3251);
not NOT1 (N5730, N5717);
or OR2 (N5731, N5726, N572);
nand NAND2 (N5732, N5727, N2812);
xor XOR2 (N5733, N5721, N4773);
or OR4 (N5734, N5729, N2831, N2548, N4967);
and AND2 (N5735, N5728, N1068);
and AND2 (N5736, N5732, N2095);
or OR3 (N5737, N5719, N2722, N346);
and AND3 (N5738, N5704, N4107, N3271);
not NOT1 (N5739, N5722);
nand NAND3 (N5740, N5735, N4155, N2187);
nor NOR3 (N5741, N5738, N313, N5338);
nor NOR4 (N5742, N5733, N1627, N4132, N4169);
not NOT1 (N5743, N5736);
not NOT1 (N5744, N5730);
not NOT1 (N5745, N5741);
not NOT1 (N5746, N5737);
or OR4 (N5747, N5744, N3534, N503, N2997);
nand NAND4 (N5748, N5731, N4056, N3603, N1745);
nand NAND3 (N5749, N5745, N2034, N253);
and AND2 (N5750, N5740, N5358);
or OR4 (N5751, N5743, N4726, N5411, N2786);
buf BUF1 (N5752, N5751);
or OR3 (N5753, N5752, N2872, N5748);
not NOT1 (N5754, N4301);
or OR4 (N5755, N5734, N4476, N4909, N4510);
buf BUF1 (N5756, N5715);
or OR3 (N5757, N5739, N4757, N4207);
or OR2 (N5758, N5742, N871);
buf BUF1 (N5759, N5750);
not NOT1 (N5760, N5758);
or OR2 (N5761, N5755, N738);
or OR4 (N5762, N5753, N2069, N5308, N173);
xor XOR2 (N5763, N5756, N2029);
and AND4 (N5764, N5762, N564, N923, N1548);
and AND2 (N5765, N5759, N1211);
buf BUF1 (N5766, N5765);
or OR4 (N5767, N5763, N111, N5471, N5673);
nand NAND4 (N5768, N5757, N3426, N4083, N2359);
buf BUF1 (N5769, N5760);
not NOT1 (N5770, N5761);
not NOT1 (N5771, N5754);
or OR2 (N5772, N5764, N973);
nor NOR2 (N5773, N5772, N3069);
nor NOR4 (N5774, N5749, N4991, N2667, N4406);
nor NOR3 (N5775, N5774, N317, N5207);
nor NOR4 (N5776, N5746, N2602, N5420, N1652);
and AND2 (N5777, N5771, N4007);
nand NAND2 (N5778, N5777, N2779);
nor NOR4 (N5779, N5767, N2767, N690, N2141);
buf BUF1 (N5780, N5779);
or OR4 (N5781, N5769, N5198, N3918, N2463);
and AND3 (N5782, N5768, N2852, N356);
xor XOR2 (N5783, N5766, N2828);
nand NAND4 (N5784, N5783, N3514, N21, N1165);
nor NOR3 (N5785, N5784, N3756, N3389);
buf BUF1 (N5786, N5776);
xor XOR2 (N5787, N5775, N153);
xor XOR2 (N5788, N5780, N1382);
nor NOR3 (N5789, N5787, N4622, N4407);
nand NAND2 (N5790, N5782, N605);
xor XOR2 (N5791, N5785, N2580);
not NOT1 (N5792, N5786);
buf BUF1 (N5793, N5789);
not NOT1 (N5794, N5791);
nand NAND4 (N5795, N5770, N875, N792, N1449);
nor NOR4 (N5796, N5747, N2116, N4097, N4860);
not NOT1 (N5797, N5773);
xor XOR2 (N5798, N5794, N2638);
nor NOR2 (N5799, N5788, N3030);
not NOT1 (N5800, N5793);
not NOT1 (N5801, N5797);
nand NAND2 (N5802, N5798, N449);
nor NOR3 (N5803, N5781, N3457, N407);
nand NAND2 (N5804, N5799, N2897);
nor NOR4 (N5805, N5795, N5029, N1503, N963);
or OR3 (N5806, N5800, N4948, N3405);
or OR3 (N5807, N5778, N5237, N1798);
buf BUF1 (N5808, N5805);
nor NOR3 (N5809, N5792, N3458, N147);
buf BUF1 (N5810, N5804);
buf BUF1 (N5811, N5801);
and AND3 (N5812, N5810, N758, N4061);
and AND4 (N5813, N5796, N4446, N111, N1643);
not NOT1 (N5814, N5812);
nor NOR3 (N5815, N5808, N2265, N2097);
buf BUF1 (N5816, N5803);
or OR3 (N5817, N5811, N732, N1079);
nor NOR4 (N5818, N5790, N5679, N5512, N2233);
not NOT1 (N5819, N5807);
nand NAND2 (N5820, N5816, N1639);
not NOT1 (N5821, N5817);
and AND2 (N5822, N5802, N5498);
nor NOR4 (N5823, N5809, N1084, N2010, N4424);
xor XOR2 (N5824, N5806, N3191);
not NOT1 (N5825, N5818);
nor NOR3 (N5826, N5822, N177, N3988);
xor XOR2 (N5827, N5825, N1695);
buf BUF1 (N5828, N5824);
buf BUF1 (N5829, N5828);
nor NOR4 (N5830, N5819, N2041, N275, N1049);
or OR3 (N5831, N5830, N806, N2141);
nand NAND4 (N5832, N5826, N2820, N2879, N5204);
not NOT1 (N5833, N5815);
buf BUF1 (N5834, N5833);
nand NAND4 (N5835, N5834, N2798, N422, N3290);
not NOT1 (N5836, N5827);
nor NOR3 (N5837, N5820, N775, N5261);
buf BUF1 (N5838, N5836);
buf BUF1 (N5839, N5838);
xor XOR2 (N5840, N5829, N5108);
and AND3 (N5841, N5821, N5708, N497);
buf BUF1 (N5842, N5814);
xor XOR2 (N5843, N5837, N1265);
nor NOR4 (N5844, N5832, N278, N5731, N4037);
or OR2 (N5845, N5831, N1277);
and AND2 (N5846, N5835, N691);
or OR2 (N5847, N5843, N4254);
and AND3 (N5848, N5840, N2022, N1349);
and AND3 (N5849, N5848, N1800, N460);
not NOT1 (N5850, N5842);
or OR4 (N5851, N5844, N252, N4490, N3610);
and AND2 (N5852, N5839, N5181);
xor XOR2 (N5853, N5813, N4134);
or OR3 (N5854, N5852, N158, N4521);
or OR4 (N5855, N5853, N1899, N1372, N2127);
xor XOR2 (N5856, N5847, N1545);
nand NAND3 (N5857, N5856, N387, N1442);
xor XOR2 (N5858, N5841, N3537);
or OR2 (N5859, N5854, N5348);
and AND2 (N5860, N5823, N3578);
buf BUF1 (N5861, N5858);
not NOT1 (N5862, N5845);
xor XOR2 (N5863, N5862, N5476);
or OR3 (N5864, N5850, N4295, N2101);
nor NOR4 (N5865, N5855, N1331, N5311, N5125);
or OR4 (N5866, N5857, N275, N2336, N1395);
nand NAND3 (N5867, N5863, N3986, N3234);
xor XOR2 (N5868, N5860, N5391);
buf BUF1 (N5869, N5868);
nor NOR2 (N5870, N5851, N1299);
or OR3 (N5871, N5864, N945, N536);
xor XOR2 (N5872, N5861, N2692);
nand NAND3 (N5873, N5849, N3681, N5494);
or OR3 (N5874, N5872, N2320, N2839);
and AND4 (N5875, N5871, N3011, N4889, N1821);
not NOT1 (N5876, N5875);
and AND4 (N5877, N5866, N4546, N2109, N1150);
not NOT1 (N5878, N5846);
not NOT1 (N5879, N5865);
not NOT1 (N5880, N5867);
or OR3 (N5881, N5870, N4156, N1557);
not NOT1 (N5882, N5873);
and AND4 (N5883, N5877, N2676, N5648, N4355);
and AND4 (N5884, N5879, N3905, N597, N2984);
not NOT1 (N5885, N5878);
nand NAND4 (N5886, N5874, N2201, N4829, N251);
not NOT1 (N5887, N5869);
buf BUF1 (N5888, N5883);
nor NOR2 (N5889, N5886, N5489);
xor XOR2 (N5890, N5882, N1001);
nor NOR3 (N5891, N5887, N3942, N595);
nor NOR2 (N5892, N5888, N3074);
nand NAND2 (N5893, N5859, N5273);
xor XOR2 (N5894, N5892, N4145);
nor NOR4 (N5895, N5880, N5834, N5727, N3029);
xor XOR2 (N5896, N5876, N5328);
nor NOR2 (N5897, N5894, N4926);
xor XOR2 (N5898, N5895, N221);
or OR3 (N5899, N5896, N4076, N5383);
xor XOR2 (N5900, N5897, N3936);
or OR2 (N5901, N5898, N5176);
nand NAND2 (N5902, N5891, N845);
buf BUF1 (N5903, N5881);
buf BUF1 (N5904, N5885);
nand NAND3 (N5905, N5904, N982, N1274);
nand NAND4 (N5906, N5890, N2373, N5822, N1328);
xor XOR2 (N5907, N5893, N3665);
xor XOR2 (N5908, N5901, N4808);
not NOT1 (N5909, N5908);
nor NOR4 (N5910, N5905, N2244, N639, N5153);
buf BUF1 (N5911, N5910);
nand NAND2 (N5912, N5906, N1402);
or OR3 (N5913, N5911, N1523, N5035);
or OR4 (N5914, N5884, N1743, N4073, N2804);
or OR3 (N5915, N5889, N877, N5709);
nor NOR2 (N5916, N5915, N319);
not NOT1 (N5917, N5909);
xor XOR2 (N5918, N5903, N5585);
xor XOR2 (N5919, N5914, N2809);
and AND3 (N5920, N5918, N5902, N2043);
buf BUF1 (N5921, N4306);
nand NAND2 (N5922, N5920, N3242);
buf BUF1 (N5923, N5921);
nor NOR3 (N5924, N5900, N3316, N5775);
or OR4 (N5925, N5919, N415, N3479, N3125);
nand NAND4 (N5926, N5923, N2924, N4689, N1595);
or OR3 (N5927, N5926, N109, N1200);
buf BUF1 (N5928, N5912);
and AND3 (N5929, N5927, N204, N2845);
or OR2 (N5930, N5922, N4004);
xor XOR2 (N5931, N5928, N2875);
not NOT1 (N5932, N5925);
nor NOR3 (N5933, N5916, N5811, N5326);
not NOT1 (N5934, N5907);
and AND3 (N5935, N5930, N2469, N522);
buf BUF1 (N5936, N5913);
not NOT1 (N5937, N5936);
or OR3 (N5938, N5932, N5799, N5718);
xor XOR2 (N5939, N5924, N5767);
nand NAND2 (N5940, N5933, N3757);
nand NAND4 (N5941, N5929, N1742, N3304, N5659);
or OR2 (N5942, N5940, N5414);
not NOT1 (N5943, N5937);
xor XOR2 (N5944, N5935, N2355);
and AND3 (N5945, N5941, N2951, N4651);
or OR2 (N5946, N5939, N5317);
not NOT1 (N5947, N5938);
and AND2 (N5948, N5917, N5838);
not NOT1 (N5949, N5944);
nand NAND4 (N5950, N5931, N2029, N3069, N2097);
nor NOR4 (N5951, N5945, N2321, N2600, N919);
nand NAND2 (N5952, N5951, N4653);
nor NOR4 (N5953, N5943, N190, N4909, N4975);
xor XOR2 (N5954, N5948, N5183);
nor NOR3 (N5955, N5899, N2188, N4292);
nor NOR4 (N5956, N5954, N3332, N74, N4260);
not NOT1 (N5957, N5955);
nor NOR2 (N5958, N5957, N2594);
and AND2 (N5959, N5934, N5384);
nor NOR4 (N5960, N5947, N1885, N3002, N3784);
buf BUF1 (N5961, N5942);
nand NAND2 (N5962, N5961, N3594);
and AND4 (N5963, N5952, N5842, N5065, N5757);
buf BUF1 (N5964, N5963);
nor NOR3 (N5965, N5946, N3612, N231);
or OR4 (N5966, N5960, N4795, N1533, N4896);
nor NOR2 (N5967, N5964, N4877);
xor XOR2 (N5968, N5949, N450);
nor NOR4 (N5969, N5962, N1431, N2790, N2932);
or OR4 (N5970, N5966, N1545, N2608, N5638);
buf BUF1 (N5971, N5967);
not NOT1 (N5972, N5970);
buf BUF1 (N5973, N5965);
nand NAND3 (N5974, N5959, N4273, N4799);
xor XOR2 (N5975, N5950, N3787);
xor XOR2 (N5976, N5968, N4753);
nand NAND4 (N5977, N5969, N1619, N2790, N5828);
xor XOR2 (N5978, N5977, N2567);
nand NAND3 (N5979, N5975, N4657, N4336);
buf BUF1 (N5980, N5958);
buf BUF1 (N5981, N5956);
nand NAND4 (N5982, N5953, N235, N1563, N2100);
not NOT1 (N5983, N5972);
nor NOR2 (N5984, N5982, N3004);
buf BUF1 (N5985, N5984);
xor XOR2 (N5986, N5979, N1638);
nand NAND4 (N5987, N5971, N3955, N4295, N4377);
nand NAND4 (N5988, N5978, N1530, N5440, N1144);
nand NAND3 (N5989, N5973, N933, N5301);
nand NAND3 (N5990, N5983, N5162, N4560);
not NOT1 (N5991, N5988);
nand NAND3 (N5992, N5985, N212, N1801);
xor XOR2 (N5993, N5976, N2472);
buf BUF1 (N5994, N5986);
not NOT1 (N5995, N5991);
nor NOR3 (N5996, N5994, N4966, N498);
buf BUF1 (N5997, N5996);
and AND4 (N5998, N5987, N5081, N3476, N4581);
not NOT1 (N5999, N5990);
nor NOR2 (N6000, N5989, N104);
and AND3 (N6001, N5974, N3404, N2021);
xor XOR2 (N6002, N5999, N3133);
buf BUF1 (N6003, N5995);
or OR4 (N6004, N6003, N2775, N2079, N4478);
nand NAND2 (N6005, N6004, N228);
and AND2 (N6006, N5992, N2360);
nand NAND4 (N6007, N6006, N1898, N3032, N5004);
nor NOR3 (N6008, N6002, N863, N1497);
nor NOR4 (N6009, N5981, N1651, N5464, N1417);
and AND4 (N6010, N5980, N3311, N4230, N5920);
xor XOR2 (N6011, N6008, N1943);
nand NAND4 (N6012, N6010, N3147, N748, N5282);
and AND2 (N6013, N5997, N5349);
nand NAND2 (N6014, N6001, N3634);
and AND2 (N6015, N6009, N440);
or OR4 (N6016, N6014, N2041, N816, N5326);
xor XOR2 (N6017, N6015, N4041);
and AND2 (N6018, N6000, N2209);
not NOT1 (N6019, N6005);
xor XOR2 (N6020, N5993, N3441);
nor NOR2 (N6021, N6018, N1828);
buf BUF1 (N6022, N6013);
or OR3 (N6023, N6007, N4842, N1674);
or OR3 (N6024, N6016, N1708, N164);
or OR2 (N6025, N6011, N927);
not NOT1 (N6026, N6021);
or OR4 (N6027, N6022, N4654, N3798, N5055);
nor NOR3 (N6028, N6017, N1948, N5162);
xor XOR2 (N6029, N5998, N3049);
buf BUF1 (N6030, N6027);
nand NAND3 (N6031, N6026, N5913, N870);
or OR3 (N6032, N6031, N767, N5269);
not NOT1 (N6033, N6012);
nand NAND2 (N6034, N6028, N624);
or OR4 (N6035, N6019, N35, N3551, N2420);
not NOT1 (N6036, N6020);
and AND4 (N6037, N6023, N2203, N1840, N2725);
not NOT1 (N6038, N6036);
or OR3 (N6039, N6033, N3095, N2721);
nand NAND4 (N6040, N6034, N3552, N3665, N1861);
not NOT1 (N6041, N6037);
or OR3 (N6042, N6035, N173, N766);
xor XOR2 (N6043, N6039, N3898);
nor NOR4 (N6044, N6024, N14, N3653, N535);
nor NOR4 (N6045, N6040, N2399, N2322, N5552);
buf BUF1 (N6046, N6045);
xor XOR2 (N6047, N6043, N5197);
nor NOR3 (N6048, N6046, N932, N3687);
nand NAND3 (N6049, N6048, N2232, N1227);
and AND2 (N6050, N6030, N930);
xor XOR2 (N6051, N6050, N880);
xor XOR2 (N6052, N6038, N1033);
not NOT1 (N6053, N6041);
buf BUF1 (N6054, N6052);
buf BUF1 (N6055, N6053);
or OR3 (N6056, N6051, N3705, N5707);
or OR4 (N6057, N6032, N1004, N1316, N1215);
nand NAND2 (N6058, N6042, N295);
nand NAND4 (N6059, N6054, N5474, N903, N324);
nand NAND3 (N6060, N6047, N4273, N3818);
not NOT1 (N6061, N6058);
nand NAND2 (N6062, N6055, N589);
and AND4 (N6063, N6049, N5243, N2387, N5876);
nor NOR3 (N6064, N6060, N5027, N759);
nand NAND2 (N6065, N6061, N5001);
xor XOR2 (N6066, N6062, N2582);
nor NOR4 (N6067, N6057, N5030, N1453, N1584);
xor XOR2 (N6068, N6065, N4426);
xor XOR2 (N6069, N6067, N1340);
nor NOR2 (N6070, N6029, N2397);
not NOT1 (N6071, N6069);
not NOT1 (N6072, N6064);
and AND3 (N6073, N6056, N2374, N3365);
not NOT1 (N6074, N6068);
nand NAND4 (N6075, N6025, N2633, N4961, N1948);
and AND4 (N6076, N6075, N5482, N5117, N3175);
or OR4 (N6077, N6076, N5468, N4079, N606);
or OR2 (N6078, N6063, N3252);
or OR3 (N6079, N6059, N720, N4460);
nand NAND3 (N6080, N6077, N854, N4032);
or OR4 (N6081, N6071, N3553, N2692, N878);
nand NAND3 (N6082, N6079, N4021, N2867);
not NOT1 (N6083, N6072);
nand NAND4 (N6084, N6073, N3210, N1235, N3654);
buf BUF1 (N6085, N6083);
and AND3 (N6086, N6074, N2808, N1289);
nor NOR2 (N6087, N6081, N5943);
nand NAND4 (N6088, N6080, N2720, N500, N5830);
buf BUF1 (N6089, N6078);
not NOT1 (N6090, N6066);
not NOT1 (N6091, N6082);
buf BUF1 (N6092, N6090);
nand NAND4 (N6093, N6086, N4815, N5500, N3418);
not NOT1 (N6094, N6088);
nor NOR3 (N6095, N6093, N3617, N2819);
xor XOR2 (N6096, N6091, N682);
and AND4 (N6097, N6085, N450, N2375, N4142);
nand NAND4 (N6098, N6096, N1018, N5373, N1383);
or OR2 (N6099, N6092, N1756);
and AND3 (N6100, N6070, N333, N5332);
or OR3 (N6101, N6097, N2682, N3666);
and AND2 (N6102, N6101, N1573);
or OR2 (N6103, N6102, N1160);
xor XOR2 (N6104, N6103, N2844);
and AND2 (N6105, N6098, N576);
buf BUF1 (N6106, N6105);
and AND2 (N6107, N6089, N2069);
and AND3 (N6108, N6084, N2084, N3545);
xor XOR2 (N6109, N6044, N1867);
xor XOR2 (N6110, N6107, N1643);
or OR3 (N6111, N6109, N4560, N1121);
xor XOR2 (N6112, N6094, N4566);
xor XOR2 (N6113, N6110, N3435);
nor NOR4 (N6114, N6099, N5454, N2674, N4358);
and AND3 (N6115, N6100, N3531, N1860);
nand NAND4 (N6116, N6087, N2596, N5669, N81);
nor NOR3 (N6117, N6113, N1340, N4594);
nand NAND3 (N6118, N6114, N5125, N1465);
xor XOR2 (N6119, N6095, N4061);
or OR2 (N6120, N6116, N1175);
not NOT1 (N6121, N6111);
buf BUF1 (N6122, N6104);
buf BUF1 (N6123, N6115);
xor XOR2 (N6124, N6117, N3596);
nor NOR2 (N6125, N6118, N6079);
xor XOR2 (N6126, N6121, N605);
nor NOR3 (N6127, N6123, N5978, N1716);
nand NAND2 (N6128, N6120, N4561);
nor NOR3 (N6129, N6124, N5415, N3908);
or OR2 (N6130, N6108, N822);
not NOT1 (N6131, N6128);
and AND2 (N6132, N6126, N1222);
nor NOR3 (N6133, N6131, N2005, N3703);
nor NOR2 (N6134, N6133, N4369);
and AND3 (N6135, N6127, N1287, N5165);
nor NOR2 (N6136, N6112, N1579);
or OR4 (N6137, N6122, N5584, N4769, N5958);
nand NAND3 (N6138, N6137, N2942, N4048);
and AND3 (N6139, N6134, N3757, N3052);
nand NAND3 (N6140, N6139, N5261, N3411);
or OR2 (N6141, N6130, N3213);
nand NAND4 (N6142, N6106, N2204, N1431, N3879);
not NOT1 (N6143, N6136);
nand NAND3 (N6144, N6132, N3368, N3919);
buf BUF1 (N6145, N6119);
buf BUF1 (N6146, N6143);
nand NAND4 (N6147, N6146, N1755, N4222, N3946);
nand NAND2 (N6148, N6145, N60);
nand NAND4 (N6149, N6125, N2730, N5550, N4859);
not NOT1 (N6150, N6135);
buf BUF1 (N6151, N6129);
and AND2 (N6152, N6151, N5524);
not NOT1 (N6153, N6152);
and AND4 (N6154, N6149, N5528, N5903, N3113);
or OR3 (N6155, N6142, N112, N967);
buf BUF1 (N6156, N6141);
or OR4 (N6157, N6140, N1672, N2849, N2096);
and AND2 (N6158, N6138, N5340);
not NOT1 (N6159, N6158);
and AND4 (N6160, N6148, N4474, N3478, N6057);
nor NOR4 (N6161, N6159, N3597, N5268, N2077);
xor XOR2 (N6162, N6157, N3136);
buf BUF1 (N6163, N6156);
or OR2 (N6164, N6160, N458);
or OR4 (N6165, N6154, N224, N2261, N192);
buf BUF1 (N6166, N6147);
nand NAND4 (N6167, N6144, N2637, N2532, N1552);
or OR2 (N6168, N6164, N3016);
buf BUF1 (N6169, N6166);
nor NOR4 (N6170, N6167, N5044, N5503, N3765);
xor XOR2 (N6171, N6169, N769);
or OR3 (N6172, N6163, N1304, N1335);
not NOT1 (N6173, N6155);
nor NOR4 (N6174, N6173, N6004, N1837, N1061);
or OR4 (N6175, N6165, N6125, N3617, N2171);
nand NAND2 (N6176, N6150, N3378);
and AND4 (N6177, N6174, N2825, N1165, N2726);
xor XOR2 (N6178, N6153, N2927);
nor NOR3 (N6179, N6178, N2612, N3872);
and AND4 (N6180, N6168, N4119, N1233, N4466);
and AND4 (N6181, N6172, N2828, N4417, N64);
and AND4 (N6182, N6175, N3727, N1770, N5092);
nor NOR3 (N6183, N6181, N1005, N442);
nand NAND2 (N6184, N6182, N1751);
and AND2 (N6185, N6180, N4568);
and AND3 (N6186, N6162, N4187, N197);
nand NAND4 (N6187, N6185, N5670, N6050, N2942);
nor NOR2 (N6188, N6170, N3284);
nand NAND2 (N6189, N6177, N531);
or OR4 (N6190, N6184, N1413, N470, N4686);
nand NAND3 (N6191, N6187, N1909, N3906);
not NOT1 (N6192, N6186);
not NOT1 (N6193, N6171);
nand NAND4 (N6194, N6191, N3145, N278, N3233);
and AND3 (N6195, N6183, N4828, N5587);
nor NOR4 (N6196, N6194, N4098, N2829, N3744);
not NOT1 (N6197, N6190);
buf BUF1 (N6198, N6189);
or OR4 (N6199, N6179, N5871, N955, N3567);
or OR3 (N6200, N6198, N5454, N3225);
and AND3 (N6201, N6192, N4716, N1242);
xor XOR2 (N6202, N6199, N4900);
and AND3 (N6203, N6197, N3644, N1317);
not NOT1 (N6204, N6195);
not NOT1 (N6205, N6202);
nor NOR4 (N6206, N6196, N1457, N153, N790);
nand NAND2 (N6207, N6204, N3686);
or OR2 (N6208, N6205, N569);
and AND4 (N6209, N6176, N1971, N5000, N505);
nand NAND2 (N6210, N6201, N3572);
nand NAND4 (N6211, N6203, N341, N2328, N1743);
not NOT1 (N6212, N6207);
nor NOR2 (N6213, N6209, N2646);
buf BUF1 (N6214, N6200);
xor XOR2 (N6215, N6206, N1679);
nand NAND3 (N6216, N6161, N5408, N5537);
buf BUF1 (N6217, N6216);
buf BUF1 (N6218, N6211);
buf BUF1 (N6219, N6210);
xor XOR2 (N6220, N6193, N2048);
xor XOR2 (N6221, N6212, N1873);
buf BUF1 (N6222, N6214);
nand NAND3 (N6223, N6220, N4262, N2663);
nor NOR3 (N6224, N6215, N3420, N4989);
xor XOR2 (N6225, N6188, N3904);
and AND2 (N6226, N6222, N5482);
and AND2 (N6227, N6223, N468);
nor NOR2 (N6228, N6213, N3873);
not NOT1 (N6229, N6224);
xor XOR2 (N6230, N6227, N4811);
and AND2 (N6231, N6230, N658);
xor XOR2 (N6232, N6228, N1100);
nand NAND3 (N6233, N6231, N1495, N5486);
nand NAND3 (N6234, N6219, N4310, N1258);
and AND3 (N6235, N6234, N2857, N3158);
buf BUF1 (N6236, N6225);
nor NOR3 (N6237, N6226, N5225, N5201);
buf BUF1 (N6238, N6232);
and AND2 (N6239, N6236, N2979);
nand NAND4 (N6240, N6218, N4129, N3302, N5192);
or OR3 (N6241, N6208, N537, N4763);
xor XOR2 (N6242, N6239, N77);
buf BUF1 (N6243, N6217);
and AND4 (N6244, N6238, N5533, N2966, N3908);
xor XOR2 (N6245, N6221, N5181);
xor XOR2 (N6246, N6242, N2382);
nand NAND4 (N6247, N6243, N4824, N424, N4388);
xor XOR2 (N6248, N6246, N5044);
not NOT1 (N6249, N6245);
nor NOR2 (N6250, N6241, N5607);
nand NAND3 (N6251, N6229, N5278, N1654);
not NOT1 (N6252, N6248);
xor XOR2 (N6253, N6249, N4180);
nor NOR3 (N6254, N6247, N2372, N3749);
nand NAND3 (N6255, N6237, N6066, N2579);
not NOT1 (N6256, N6254);
nand NAND2 (N6257, N6250, N5083);
buf BUF1 (N6258, N6240);
nor NOR3 (N6259, N6235, N5680, N3605);
buf BUF1 (N6260, N6255);
not NOT1 (N6261, N6253);
nand NAND4 (N6262, N6233, N4772, N5152, N2988);
nand NAND4 (N6263, N6259, N5418, N2392, N546);
nor NOR2 (N6264, N6251, N1744);
and AND3 (N6265, N6263, N1192, N2960);
nor NOR2 (N6266, N6258, N6065);
nand NAND2 (N6267, N6265, N5787);
buf BUF1 (N6268, N6244);
not NOT1 (N6269, N6256);
nand NAND4 (N6270, N6266, N3357, N4869, N52);
or OR3 (N6271, N6262, N1806, N593);
buf BUF1 (N6272, N6264);
not NOT1 (N6273, N6269);
or OR4 (N6274, N6260, N2150, N6247, N6140);
buf BUF1 (N6275, N6268);
nand NAND4 (N6276, N6252, N4796, N5627, N4781);
nor NOR2 (N6277, N6275, N2661);
buf BUF1 (N6278, N6257);
and AND4 (N6279, N6278, N2857, N1639, N4415);
and AND4 (N6280, N6273, N620, N4844, N2568);
and AND2 (N6281, N6279, N3926);
nand NAND4 (N6282, N6276, N499, N1762, N5653);
or OR2 (N6283, N6274, N2140);
buf BUF1 (N6284, N6282);
nor NOR2 (N6285, N6284, N4443);
buf BUF1 (N6286, N6272);
or OR2 (N6287, N6267, N1979);
nor NOR3 (N6288, N6286, N794, N2083);
nand NAND2 (N6289, N6287, N5144);
nor NOR3 (N6290, N6288, N3577, N3154);
not NOT1 (N6291, N6277);
nor NOR3 (N6292, N6281, N4826, N1018);
not NOT1 (N6293, N6261);
not NOT1 (N6294, N6291);
and AND3 (N6295, N6270, N5516, N4712);
not NOT1 (N6296, N6271);
xor XOR2 (N6297, N6294, N4450);
and AND4 (N6298, N6296, N6067, N2612, N4156);
and AND2 (N6299, N6297, N1025);
and AND4 (N6300, N6290, N1664, N4926, N4480);
nand NAND4 (N6301, N6298, N1702, N87, N2700);
nand NAND3 (N6302, N6285, N84, N625);
xor XOR2 (N6303, N6280, N855);
or OR4 (N6304, N6299, N5797, N222, N4691);
and AND3 (N6305, N6303, N5683, N3308);
or OR3 (N6306, N6300, N4054, N5572);
not NOT1 (N6307, N6301);
nand NAND3 (N6308, N6307, N439, N3757);
nand NAND2 (N6309, N6306, N2491);
or OR2 (N6310, N6289, N5415);
buf BUF1 (N6311, N6283);
nor NOR2 (N6312, N6295, N2095);
and AND4 (N6313, N6302, N2220, N4541, N5045);
buf BUF1 (N6314, N6313);
nand NAND4 (N6315, N6305, N5681, N3893, N5592);
and AND4 (N6316, N6314, N6224, N4976, N6259);
or OR4 (N6317, N6293, N1918, N4719, N922);
buf BUF1 (N6318, N6304);
buf BUF1 (N6319, N6315);
nor NOR4 (N6320, N6311, N1586, N2879, N262);
nor NOR2 (N6321, N6316, N5439);
nor NOR2 (N6322, N6319, N4491);
nand NAND4 (N6323, N6322, N4862, N3756, N2277);
nor NOR4 (N6324, N6320, N4486, N345, N423);
and AND2 (N6325, N6324, N5174);
or OR2 (N6326, N6317, N88);
not NOT1 (N6327, N6321);
nor NOR4 (N6328, N6327, N1022, N5266, N1499);
nand NAND4 (N6329, N6309, N6126, N3247, N354);
not NOT1 (N6330, N6326);
and AND4 (N6331, N6292, N1284, N3998, N3460);
buf BUF1 (N6332, N6312);
or OR2 (N6333, N6310, N5442);
nor NOR3 (N6334, N6329, N4241, N523);
or OR4 (N6335, N6323, N1022, N505, N2136);
nor NOR4 (N6336, N6330, N2494, N2889, N3802);
buf BUF1 (N6337, N6328);
and AND2 (N6338, N6331, N3479);
not NOT1 (N6339, N6308);
buf BUF1 (N6340, N6334);
buf BUF1 (N6341, N6339);
nand NAND4 (N6342, N6338, N3984, N4946, N17);
nand NAND2 (N6343, N6341, N5729);
xor XOR2 (N6344, N6335, N6319);
xor XOR2 (N6345, N6337, N6144);
xor XOR2 (N6346, N6342, N2449);
nand NAND2 (N6347, N6340, N1300);
nand NAND3 (N6348, N6325, N3781, N3168);
nor NOR2 (N6349, N6343, N5702);
or OR3 (N6350, N6333, N2623, N5525);
nor NOR4 (N6351, N6349, N445, N4500, N319);
buf BUF1 (N6352, N6332);
and AND4 (N6353, N6336, N5349, N91, N3440);
xor XOR2 (N6354, N6348, N71);
not NOT1 (N6355, N6318);
and AND4 (N6356, N6353, N510, N5233, N6031);
nand NAND2 (N6357, N6355, N1401);
buf BUF1 (N6358, N6346);
nor NOR3 (N6359, N6350, N5453, N2079);
and AND3 (N6360, N6344, N6244, N1123);
or OR3 (N6361, N6347, N1449, N2371);
nor NOR3 (N6362, N6361, N1427, N610);
not NOT1 (N6363, N6362);
buf BUF1 (N6364, N6359);
and AND2 (N6365, N6352, N4180);
xor XOR2 (N6366, N6363, N2149);
and AND3 (N6367, N6357, N4602, N2670);
nor NOR2 (N6368, N6354, N3621);
nor NOR3 (N6369, N6358, N185, N1473);
or OR4 (N6370, N6351, N5817, N4090, N4562);
not NOT1 (N6371, N6365);
buf BUF1 (N6372, N6370);
or OR2 (N6373, N6372, N3848);
xor XOR2 (N6374, N6366, N3900);
xor XOR2 (N6375, N6345, N6334);
and AND2 (N6376, N6374, N1641);
xor XOR2 (N6377, N6375, N702);
not NOT1 (N6378, N6360);
or OR3 (N6379, N6373, N3000, N2089);
not NOT1 (N6380, N6377);
or OR4 (N6381, N6378, N5517, N3841, N1298);
xor XOR2 (N6382, N6381, N6352);
nand NAND3 (N6383, N6371, N4533, N96);
buf BUF1 (N6384, N6379);
or OR2 (N6385, N6382, N1807);
buf BUF1 (N6386, N6380);
buf BUF1 (N6387, N6368);
and AND3 (N6388, N6386, N5203, N3325);
buf BUF1 (N6389, N6388);
nand NAND4 (N6390, N6389, N5388, N5506, N3084);
not NOT1 (N6391, N6367);
xor XOR2 (N6392, N6383, N3536);
and AND3 (N6393, N6384, N6094, N4723);
or OR2 (N6394, N6393, N1844);
not NOT1 (N6395, N6385);
or OR3 (N6396, N6395, N2047, N365);
buf BUF1 (N6397, N6356);
and AND4 (N6398, N6397, N3966, N5855, N4383);
or OR4 (N6399, N6392, N3590, N1210, N3455);
xor XOR2 (N6400, N6399, N3144);
or OR2 (N6401, N6369, N6043);
or OR2 (N6402, N6394, N2374);
buf BUF1 (N6403, N6400);
or OR2 (N6404, N6364, N5792);
xor XOR2 (N6405, N6401, N372);
xor XOR2 (N6406, N6376, N5097);
not NOT1 (N6407, N6398);
nor NOR2 (N6408, N6403, N3888);
buf BUF1 (N6409, N6404);
nand NAND3 (N6410, N6387, N646, N5242);
xor XOR2 (N6411, N6406, N3898);
or OR4 (N6412, N6411, N5442, N6406, N2731);
xor XOR2 (N6413, N6405, N517);
xor XOR2 (N6414, N6412, N5534);
or OR3 (N6415, N6391, N2565, N4914);
buf BUF1 (N6416, N6396);
nand NAND2 (N6417, N6408, N123);
or OR3 (N6418, N6414, N3978, N5412);
and AND4 (N6419, N6415, N5184, N1752, N3836);
or OR2 (N6420, N6407, N5722);
buf BUF1 (N6421, N6416);
nand NAND2 (N6422, N6410, N4995);
nor NOR2 (N6423, N6418, N87);
buf BUF1 (N6424, N6420);
and AND3 (N6425, N6409, N959, N3332);
nand NAND2 (N6426, N6402, N2194);
nand NAND4 (N6427, N6426, N4683, N3094, N4103);
buf BUF1 (N6428, N6423);
and AND2 (N6429, N6425, N5013);
and AND3 (N6430, N6429, N6287, N285);
not NOT1 (N6431, N6417);
nor NOR3 (N6432, N6427, N2134, N3664);
or OR3 (N6433, N6419, N69, N2443);
not NOT1 (N6434, N6424);
nor NOR4 (N6435, N6390, N1822, N1363, N3218);
xor XOR2 (N6436, N6434, N3953);
nand NAND2 (N6437, N6413, N2230);
not NOT1 (N6438, N6437);
not NOT1 (N6439, N6438);
buf BUF1 (N6440, N6421);
nand NAND4 (N6441, N6436, N2056, N817, N2587);
nand NAND4 (N6442, N6431, N4156, N1724, N3502);
buf BUF1 (N6443, N6435);
not NOT1 (N6444, N6422);
or OR4 (N6445, N6444, N6328, N6024, N886);
or OR2 (N6446, N6432, N4961);
not NOT1 (N6447, N6430);
not NOT1 (N6448, N6441);
xor XOR2 (N6449, N6447, N4311);
xor XOR2 (N6450, N6445, N2700);
nor NOR3 (N6451, N6433, N5619, N617);
nand NAND2 (N6452, N6428, N1885);
not NOT1 (N6453, N6440);
nand NAND4 (N6454, N6439, N1318, N4838, N228);
and AND4 (N6455, N6453, N5429, N148, N5174);
nand NAND3 (N6456, N6450, N4265, N3939);
nand NAND3 (N6457, N6442, N4499, N2395);
buf BUF1 (N6458, N6446);
nand NAND2 (N6459, N6443, N4600);
not NOT1 (N6460, N6451);
nor NOR3 (N6461, N6457, N3487, N5446);
or OR4 (N6462, N6458, N3581, N6394, N3322);
nor NOR4 (N6463, N6452, N804, N2012, N4203);
buf BUF1 (N6464, N6460);
nand NAND4 (N6465, N6448, N2072, N6031, N187);
xor XOR2 (N6466, N6465, N3804);
buf BUF1 (N6467, N6463);
or OR2 (N6468, N6464, N3828);
and AND3 (N6469, N6466, N1594, N3471);
or OR2 (N6470, N6467, N3726);
or OR2 (N6471, N6459, N5793);
xor XOR2 (N6472, N6461, N4809);
xor XOR2 (N6473, N6472, N2374);
and AND3 (N6474, N6449, N2777, N1972);
nor NOR2 (N6475, N6455, N6307);
nand NAND3 (N6476, N6471, N1660, N4884);
nor NOR4 (N6477, N6456, N585, N898, N646);
nor NOR4 (N6478, N6475, N2372, N2402, N2825);
not NOT1 (N6479, N6468);
or OR2 (N6480, N6474, N54);
xor XOR2 (N6481, N6469, N3143);
and AND3 (N6482, N6476, N1748, N5609);
buf BUF1 (N6483, N6478);
not NOT1 (N6484, N6481);
not NOT1 (N6485, N6473);
xor XOR2 (N6486, N6477, N4859);
or OR4 (N6487, N6462, N252, N2413, N4630);
xor XOR2 (N6488, N6480, N2461);
buf BUF1 (N6489, N6486);
xor XOR2 (N6490, N6483, N3994);
nand NAND3 (N6491, N6485, N3615, N2906);
not NOT1 (N6492, N6490);
or OR4 (N6493, N6492, N1892, N5860, N242);
and AND2 (N6494, N6493, N5860);
buf BUF1 (N6495, N6489);
nor NOR4 (N6496, N6488, N3271, N1715, N3295);
xor XOR2 (N6497, N6454, N2364);
nor NOR3 (N6498, N6491, N1508, N5973);
or OR3 (N6499, N6484, N4785, N3883);
or OR3 (N6500, N6479, N1958, N343);
nor NOR2 (N6501, N6494, N3308);
and AND2 (N6502, N6498, N4466);
buf BUF1 (N6503, N6500);
or OR4 (N6504, N6502, N5505, N6305, N1924);
xor XOR2 (N6505, N6482, N2502);
nor NOR2 (N6506, N6505, N3510);
nor NOR2 (N6507, N6497, N2711);
and AND2 (N6508, N6496, N6421);
and AND2 (N6509, N6506, N6303);
xor XOR2 (N6510, N6508, N1521);
nand NAND4 (N6511, N6470, N1764, N6125, N1834);
xor XOR2 (N6512, N6501, N4064);
xor XOR2 (N6513, N6510, N4776);
or OR4 (N6514, N6513, N1755, N74, N782);
and AND4 (N6515, N6504, N4267, N6414, N6016);
or OR2 (N6516, N6515, N2298);
and AND2 (N6517, N6511, N6135);
not NOT1 (N6518, N6514);
not NOT1 (N6519, N6487);
buf BUF1 (N6520, N6495);
nor NOR4 (N6521, N6517, N4169, N5232, N5324);
xor XOR2 (N6522, N6512, N573);
nor NOR2 (N6523, N6509, N110);
and AND3 (N6524, N6503, N4740, N399);
xor XOR2 (N6525, N6521, N1859);
not NOT1 (N6526, N6499);
nand NAND3 (N6527, N6507, N4286, N2043);
xor XOR2 (N6528, N6525, N5667);
nor NOR3 (N6529, N6520, N3744, N6406);
not NOT1 (N6530, N6518);
or OR3 (N6531, N6522, N1329, N4801);
xor XOR2 (N6532, N6527, N3298);
xor XOR2 (N6533, N6531, N5931);
xor XOR2 (N6534, N6524, N6532);
not NOT1 (N6535, N1256);
not NOT1 (N6536, N6519);
and AND2 (N6537, N6526, N4466);
or OR2 (N6538, N6529, N1626);
xor XOR2 (N6539, N6538, N5331);
nor NOR2 (N6540, N6539, N5613);
nor NOR4 (N6541, N6537, N5187, N1996, N2791);
buf BUF1 (N6542, N6516);
not NOT1 (N6543, N6523);
and AND4 (N6544, N6528, N6100, N1431, N6412);
or OR4 (N6545, N6541, N4901, N1382, N837);
and AND3 (N6546, N6536, N4789, N6417);
buf BUF1 (N6547, N6535);
not NOT1 (N6548, N6540);
nor NOR3 (N6549, N6547, N1733, N4154);
nor NOR3 (N6550, N6544, N3095, N655);
or OR3 (N6551, N6550, N5052, N5849);
xor XOR2 (N6552, N6548, N3916);
buf BUF1 (N6553, N6552);
and AND2 (N6554, N6549, N3716);
and AND2 (N6555, N6546, N924);
or OR3 (N6556, N6534, N2131, N189);
nand NAND2 (N6557, N6543, N5603);
nand NAND3 (N6558, N6542, N2888, N2725);
not NOT1 (N6559, N6553);
nand NAND3 (N6560, N6559, N125, N3366);
nor NOR2 (N6561, N6530, N1600);
nor NOR2 (N6562, N6556, N5236);
or OR2 (N6563, N6557, N3518);
xor XOR2 (N6564, N6563, N5658);
nor NOR2 (N6565, N6561, N898);
and AND4 (N6566, N6562, N4209, N4158, N2899);
and AND4 (N6567, N6558, N476, N2059, N4200);
or OR4 (N6568, N6545, N5925, N5066, N1488);
buf BUF1 (N6569, N6533);
xor XOR2 (N6570, N6555, N6564);
or OR3 (N6571, N4942, N2260, N1273);
buf BUF1 (N6572, N6569);
or OR3 (N6573, N6565, N3036, N5218);
or OR2 (N6574, N6560, N2975);
not NOT1 (N6575, N6572);
not NOT1 (N6576, N6568);
nand NAND2 (N6577, N6575, N5808);
nor NOR2 (N6578, N6554, N1816);
nor NOR2 (N6579, N6566, N964);
not NOT1 (N6580, N6570);
nand NAND2 (N6581, N6567, N5061);
nand NAND4 (N6582, N6581, N4126, N3881, N1340);
nor NOR2 (N6583, N6578, N2938);
nand NAND3 (N6584, N6583, N6055, N3518);
buf BUF1 (N6585, N6577);
nor NOR4 (N6586, N6573, N4943, N1076, N3939);
xor XOR2 (N6587, N6551, N483);
nor NOR3 (N6588, N6574, N5381, N4904);
nor NOR2 (N6589, N6582, N2709);
buf BUF1 (N6590, N6587);
not NOT1 (N6591, N6588);
not NOT1 (N6592, N6585);
or OR3 (N6593, N6592, N6446, N1694);
buf BUF1 (N6594, N6590);
nand NAND2 (N6595, N6576, N5217);
nand NAND3 (N6596, N6571, N5843, N1552);
buf BUF1 (N6597, N6589);
or OR2 (N6598, N6594, N3678);
not NOT1 (N6599, N6598);
xor XOR2 (N6600, N6591, N948);
xor XOR2 (N6601, N6596, N2983);
xor XOR2 (N6602, N6593, N2311);
and AND2 (N6603, N6599, N5367);
xor XOR2 (N6604, N6595, N2812);
or OR2 (N6605, N6603, N2933);
nor NOR4 (N6606, N6586, N5958, N1512, N2808);
nor NOR3 (N6607, N6604, N6156, N8);
nor NOR3 (N6608, N6580, N5137, N5591);
or OR4 (N6609, N6602, N1904, N4878, N4661);
and AND4 (N6610, N6608, N3304, N306, N1538);
nor NOR3 (N6611, N6605, N6412, N2965);
nor NOR2 (N6612, N6609, N2520);
or OR3 (N6613, N6606, N4441, N3268);
or OR3 (N6614, N6601, N4877, N1448);
nand NAND4 (N6615, N6579, N5305, N3710, N4037);
and AND3 (N6616, N6600, N6025, N6274);
xor XOR2 (N6617, N6612, N2737);
buf BUF1 (N6618, N6611);
or OR3 (N6619, N6616, N5476, N1811);
not NOT1 (N6620, N6615);
xor XOR2 (N6621, N6613, N4363);
or OR2 (N6622, N6597, N1482);
or OR3 (N6623, N6620, N2395, N3947);
not NOT1 (N6624, N6614);
not NOT1 (N6625, N6618);
nand NAND3 (N6626, N6607, N92, N3501);
buf BUF1 (N6627, N6619);
nor NOR2 (N6628, N6624, N3433);
not NOT1 (N6629, N6610);
xor XOR2 (N6630, N6626, N3942);
buf BUF1 (N6631, N6584);
xor XOR2 (N6632, N6625, N721);
not NOT1 (N6633, N6623);
and AND2 (N6634, N6630, N4903);
buf BUF1 (N6635, N6633);
and AND3 (N6636, N6622, N5752, N4707);
not NOT1 (N6637, N6631);
nand NAND3 (N6638, N6627, N3949, N3291);
nor NOR2 (N6639, N6636, N6541);
or OR4 (N6640, N6629, N6299, N4733, N4687);
nand NAND2 (N6641, N6634, N5336);
and AND2 (N6642, N6628, N6416);
xor XOR2 (N6643, N6639, N5163);
or OR4 (N6644, N6638, N2097, N3765, N1793);
buf BUF1 (N6645, N6632);
and AND4 (N6646, N6617, N5586, N841, N4342);
not NOT1 (N6647, N6641);
nor NOR4 (N6648, N6642, N295, N2029, N5749);
or OR2 (N6649, N6635, N1812);
buf BUF1 (N6650, N6646);
and AND2 (N6651, N6649, N5451);
not NOT1 (N6652, N6644);
nor NOR3 (N6653, N6637, N4562, N3355);
xor XOR2 (N6654, N6648, N2928);
nor NOR4 (N6655, N6640, N6003, N633, N3485);
and AND3 (N6656, N6645, N2676, N357);
nand NAND2 (N6657, N6654, N90);
xor XOR2 (N6658, N6621, N1016);
or OR4 (N6659, N6657, N5289, N4243, N6106);
or OR4 (N6660, N6643, N1371, N3823, N1976);
not NOT1 (N6661, N6660);
and AND3 (N6662, N6661, N2278, N3228);
or OR4 (N6663, N6658, N3249, N2604, N1624);
and AND2 (N6664, N6662, N5741);
nor NOR2 (N6665, N6651, N474);
buf BUF1 (N6666, N6664);
not NOT1 (N6667, N6663);
and AND4 (N6668, N6667, N5657, N2132, N5884);
buf BUF1 (N6669, N6656);
buf BUF1 (N6670, N6653);
or OR2 (N6671, N6652, N3499);
nand NAND2 (N6672, N6668, N3961);
and AND2 (N6673, N6650, N2229);
not NOT1 (N6674, N6647);
or OR2 (N6675, N6673, N6027);
not NOT1 (N6676, N6674);
not NOT1 (N6677, N6666);
and AND2 (N6678, N6675, N2063);
or OR4 (N6679, N6670, N3621, N311, N508);
nor NOR4 (N6680, N6677, N3415, N4612, N2258);
nor NOR3 (N6681, N6672, N3565, N2046);
nor NOR3 (N6682, N6676, N4048, N603);
nand NAND4 (N6683, N6678, N913, N3756, N275);
not NOT1 (N6684, N6683);
buf BUF1 (N6685, N6669);
nand NAND4 (N6686, N6665, N4479, N1985, N6631);
or OR2 (N6687, N6680, N4595);
or OR3 (N6688, N6671, N2290, N4931);
or OR2 (N6689, N6686, N2237);
nor NOR3 (N6690, N6682, N6425, N3447);
xor XOR2 (N6691, N6685, N3997);
xor XOR2 (N6692, N6688, N1284);
xor XOR2 (N6693, N6692, N137);
not NOT1 (N6694, N6691);
and AND4 (N6695, N6679, N1963, N5222, N4113);
xor XOR2 (N6696, N6693, N393);
nor NOR4 (N6697, N6690, N145, N6609, N4354);
and AND2 (N6698, N6689, N5582);
not NOT1 (N6699, N6696);
and AND2 (N6700, N6694, N349);
not NOT1 (N6701, N6695);
not NOT1 (N6702, N6701);
not NOT1 (N6703, N6698);
not NOT1 (N6704, N6703);
nor NOR2 (N6705, N6659, N6224);
nor NOR2 (N6706, N6681, N1767);
xor XOR2 (N6707, N6700, N1700);
xor XOR2 (N6708, N6655, N4186);
or OR4 (N6709, N6707, N2036, N3160, N4438);
nand NAND3 (N6710, N6704, N190, N3362);
buf BUF1 (N6711, N6709);
buf BUF1 (N6712, N6710);
xor XOR2 (N6713, N6711, N6236);
not NOT1 (N6714, N6712);
and AND3 (N6715, N6699, N5049, N1568);
nand NAND3 (N6716, N6697, N3405, N607);
nor NOR2 (N6717, N6706, N4275);
and AND3 (N6718, N6702, N1994, N360);
and AND3 (N6719, N6705, N3641, N2385);
or OR4 (N6720, N6715, N3603, N4955, N1229);
nor NOR2 (N6721, N6687, N5395);
nand NAND4 (N6722, N6717, N6260, N6547, N2884);
buf BUF1 (N6723, N6714);
xor XOR2 (N6724, N6723, N6625);
nor NOR4 (N6725, N6719, N482, N5950, N2768);
nor NOR4 (N6726, N6716, N1145, N3619, N4381);
not NOT1 (N6727, N6724);
buf BUF1 (N6728, N6726);
not NOT1 (N6729, N6718);
xor XOR2 (N6730, N6729, N6420);
nor NOR4 (N6731, N6725, N4131, N1784, N3720);
nand NAND2 (N6732, N6722, N3536);
buf BUF1 (N6733, N6721);
and AND3 (N6734, N6684, N5857, N4082);
nor NOR3 (N6735, N6734, N85, N6602);
not NOT1 (N6736, N6733);
not NOT1 (N6737, N6735);
nand NAND3 (N6738, N6720, N1953, N6372);
nand NAND3 (N6739, N6713, N3439, N4133);
buf BUF1 (N6740, N6736);
xor XOR2 (N6741, N6731, N2238);
or OR3 (N6742, N6732, N1954, N3157);
nand NAND4 (N6743, N6742, N3920, N3812, N2612);
nor NOR4 (N6744, N6739, N3980, N2620, N3102);
nor NOR3 (N6745, N6743, N3700, N968);
buf BUF1 (N6746, N6738);
nor NOR4 (N6747, N6730, N4990, N1139, N6144);
not NOT1 (N6748, N6745);
and AND4 (N6749, N6740, N4383, N5958, N6426);
buf BUF1 (N6750, N6744);
nand NAND4 (N6751, N6708, N2242, N4993, N482);
nand NAND4 (N6752, N6728, N1175, N1633, N6498);
and AND3 (N6753, N6748, N1744, N2613);
nand NAND2 (N6754, N6737, N2699);
buf BUF1 (N6755, N6746);
nand NAND4 (N6756, N6747, N4145, N3601, N639);
nor NOR2 (N6757, N6727, N1097);
or OR2 (N6758, N6757, N2304);
and AND2 (N6759, N6751, N4217);
buf BUF1 (N6760, N6755);
not NOT1 (N6761, N6759);
not NOT1 (N6762, N6758);
xor XOR2 (N6763, N6750, N5983);
nand NAND2 (N6764, N6760, N6613);
nand NAND4 (N6765, N6753, N3290, N2770, N1067);
and AND2 (N6766, N6764, N3196);
and AND3 (N6767, N6756, N2275, N3429);
nand NAND2 (N6768, N6766, N1836);
nand NAND3 (N6769, N6767, N541, N4302);
nor NOR2 (N6770, N6741, N3663);
not NOT1 (N6771, N6749);
nor NOR2 (N6772, N6754, N4712);
or OR4 (N6773, N6765, N2651, N3996, N4368);
nand NAND3 (N6774, N6769, N2792, N4160);
xor XOR2 (N6775, N6763, N2492);
buf BUF1 (N6776, N6768);
not NOT1 (N6777, N6775);
or OR2 (N6778, N6776, N3651);
nand NAND3 (N6779, N6761, N471, N141);
not NOT1 (N6780, N6770);
nor NOR4 (N6781, N6780, N1974, N2836, N6144);
buf BUF1 (N6782, N6778);
or OR2 (N6783, N6774, N2885);
nand NAND4 (N6784, N6783, N3237, N4618, N5606);
and AND4 (N6785, N6773, N3923, N5308, N3782);
nor NOR2 (N6786, N6784, N1802);
nor NOR2 (N6787, N6786, N5429);
nand NAND4 (N6788, N6752, N3933, N3000, N1020);
not NOT1 (N6789, N6787);
nand NAND2 (N6790, N6772, N495);
xor XOR2 (N6791, N6771, N701);
and AND4 (N6792, N6785, N4081, N2793, N6502);
buf BUF1 (N6793, N6779);
not NOT1 (N6794, N6762);
buf BUF1 (N6795, N6781);
and AND2 (N6796, N6792, N3352);
xor XOR2 (N6797, N6790, N2819);
nor NOR3 (N6798, N6797, N1449, N5214);
buf BUF1 (N6799, N6789);
and AND2 (N6800, N6791, N2844);
nand NAND3 (N6801, N6799, N5482, N3451);
not NOT1 (N6802, N6795);
not NOT1 (N6803, N6801);
not NOT1 (N6804, N6788);
not NOT1 (N6805, N6777);
nand NAND2 (N6806, N6803, N2562);
nand NAND4 (N6807, N6804, N4634, N3006, N1118);
or OR4 (N6808, N6805, N3207, N1573, N266);
buf BUF1 (N6809, N6802);
nor NOR4 (N6810, N6809, N3897, N1478, N3903);
xor XOR2 (N6811, N6800, N6476);
or OR3 (N6812, N6810, N2410, N4280);
nand NAND2 (N6813, N6782, N1315);
buf BUF1 (N6814, N6808);
and AND4 (N6815, N6812, N4221, N6020, N5969);
nor NOR2 (N6816, N6793, N2802);
or OR4 (N6817, N6807, N1974, N1518, N910);
nor NOR3 (N6818, N6811, N4626, N3253);
and AND3 (N6819, N6806, N2879, N2320);
nor NOR3 (N6820, N6818, N1194, N6508);
nand NAND4 (N6821, N6815, N5499, N6044, N298);
nand NAND4 (N6822, N6796, N4130, N2562, N5666);
and AND3 (N6823, N6822, N2820, N3195);
nand NAND3 (N6824, N6816, N6753, N623);
nand NAND3 (N6825, N6823, N5088, N1525);
not NOT1 (N6826, N6817);
nand NAND4 (N6827, N6820, N4398, N239, N6131);
buf BUF1 (N6828, N6794);
not NOT1 (N6829, N6824);
xor XOR2 (N6830, N6798, N3685);
nand NAND4 (N6831, N6821, N5709, N359, N4969);
nor NOR3 (N6832, N6830, N6052, N1211);
not NOT1 (N6833, N6826);
xor XOR2 (N6834, N6813, N4600);
nor NOR2 (N6835, N6819, N5439);
nor NOR2 (N6836, N6829, N1962);
and AND3 (N6837, N6827, N1414, N2912);
or OR4 (N6838, N6831, N6062, N1733, N4108);
xor XOR2 (N6839, N6836, N304);
buf BUF1 (N6840, N6825);
or OR2 (N6841, N6832, N973);
xor XOR2 (N6842, N6814, N5124);
not NOT1 (N6843, N6842);
not NOT1 (N6844, N6843);
nor NOR2 (N6845, N6837, N6508);
nand NAND4 (N6846, N6841, N2060, N6702, N201);
nand NAND2 (N6847, N6835, N1562);
not NOT1 (N6848, N6845);
not NOT1 (N6849, N6839);
nand NAND4 (N6850, N6834, N6803, N2722, N1936);
xor XOR2 (N6851, N6849, N3657);
or OR3 (N6852, N6847, N6789, N147);
nand NAND4 (N6853, N6844, N270, N6476, N3033);
xor XOR2 (N6854, N6840, N4673);
not NOT1 (N6855, N6854);
and AND4 (N6856, N6850, N878, N3439, N5294);
and AND3 (N6857, N6838, N999, N6718);
not NOT1 (N6858, N6857);
or OR4 (N6859, N6856, N5517, N5739, N5896);
nor NOR4 (N6860, N6852, N1848, N5642, N4950);
buf BUF1 (N6861, N6860);
and AND3 (N6862, N6855, N648, N6473);
nand NAND4 (N6863, N6846, N4482, N728, N2622);
not NOT1 (N6864, N6858);
nor NOR4 (N6865, N6828, N5000, N3894, N1939);
xor XOR2 (N6866, N6865, N2627);
and AND3 (N6867, N6851, N1657, N2157);
or OR3 (N6868, N6867, N5444, N1216);
or OR4 (N6869, N6863, N4916, N926, N5995);
nor NOR2 (N6870, N6833, N5333);
xor XOR2 (N6871, N6870, N2655);
nor NOR3 (N6872, N6859, N6802, N1957);
and AND3 (N6873, N6868, N6017, N6234);
xor XOR2 (N6874, N6872, N5453);
nor NOR3 (N6875, N6853, N3590, N336);
nor NOR3 (N6876, N6861, N6185, N192);
xor XOR2 (N6877, N6848, N5292);
nand NAND4 (N6878, N6874, N3194, N6042, N122);
and AND2 (N6879, N6877, N711);
or OR3 (N6880, N6875, N2321, N2935);
nand NAND2 (N6881, N6866, N4387);
nand NAND3 (N6882, N6879, N4260, N4962);
nor NOR4 (N6883, N6878, N3911, N3406, N6793);
and AND4 (N6884, N6876, N5213, N4788, N1613);
buf BUF1 (N6885, N6883);
nor NOR2 (N6886, N6880, N1948);
or OR3 (N6887, N6881, N2383, N610);
not NOT1 (N6888, N6884);
not NOT1 (N6889, N6864);
nor NOR2 (N6890, N6888, N1343);
or OR4 (N6891, N6885, N957, N812, N564);
xor XOR2 (N6892, N6886, N3248);
or OR3 (N6893, N6873, N2272, N3702);
nand NAND3 (N6894, N6871, N2601, N3678);
not NOT1 (N6895, N6892);
xor XOR2 (N6896, N6882, N4124);
and AND4 (N6897, N6890, N3063, N2987, N1922);
and AND4 (N6898, N6893, N881, N2285, N3643);
and AND4 (N6899, N6869, N4826, N2666, N6512);
nand NAND3 (N6900, N6862, N3166, N4608);
nor NOR3 (N6901, N6900, N3415, N5600);
nand NAND2 (N6902, N6896, N4874);
nand NAND2 (N6903, N6902, N5640);
not NOT1 (N6904, N6895);
buf BUF1 (N6905, N6898);
xor XOR2 (N6906, N6903, N1507);
not NOT1 (N6907, N6906);
or OR2 (N6908, N6904, N6111);
nor NOR3 (N6909, N6901, N6711, N4860);
nor NOR2 (N6910, N6909, N3179);
or OR3 (N6911, N6891, N3173, N2750);
nand NAND3 (N6912, N6887, N3591, N671);
buf BUF1 (N6913, N6894);
nand NAND4 (N6914, N6912, N1439, N6512, N4557);
xor XOR2 (N6915, N6914, N6844);
not NOT1 (N6916, N6910);
nor NOR2 (N6917, N6889, N2483);
not NOT1 (N6918, N6916);
or OR2 (N6919, N6908, N2456);
xor XOR2 (N6920, N6907, N5231);
or OR4 (N6921, N6905, N2950, N5075, N5423);
not NOT1 (N6922, N6921);
and AND2 (N6923, N6915, N6101);
nor NOR2 (N6924, N6920, N1283);
not NOT1 (N6925, N6899);
nand NAND4 (N6926, N6897, N1138, N4156, N2750);
buf BUF1 (N6927, N6923);
nor NOR2 (N6928, N6918, N1841);
or OR3 (N6929, N6926, N6166, N4843);
nor NOR4 (N6930, N6919, N2939, N3686, N3352);
nand NAND4 (N6931, N6930, N5109, N2977, N2740);
or OR3 (N6932, N6925, N5505, N847);
not NOT1 (N6933, N6932);
nor NOR2 (N6934, N6913, N4911);
buf BUF1 (N6935, N6929);
buf BUF1 (N6936, N6931);
xor XOR2 (N6937, N6933, N2312);
nand NAND3 (N6938, N6922, N3158, N1816);
not NOT1 (N6939, N6924);
not NOT1 (N6940, N6938);
nor NOR3 (N6941, N6936, N3917, N3196);
or OR2 (N6942, N6935, N6395);
buf BUF1 (N6943, N6941);
or OR2 (N6944, N6917, N2419);
or OR3 (N6945, N6943, N3706, N3120);
and AND4 (N6946, N6911, N6904, N6077, N551);
and AND4 (N6947, N6939, N231, N4630, N3542);
or OR3 (N6948, N6946, N5488, N334);
nand NAND3 (N6949, N6947, N3767, N3429);
nor NOR2 (N6950, N6928, N277);
not NOT1 (N6951, N6945);
and AND4 (N6952, N6927, N2606, N5987, N5819);
or OR4 (N6953, N6949, N4084, N1202, N3182);
nand NAND2 (N6954, N6953, N894);
xor XOR2 (N6955, N6952, N6379);
or OR2 (N6956, N6942, N3283);
or OR3 (N6957, N6955, N2224, N3190);
and AND2 (N6958, N6934, N3011);
nand NAND4 (N6959, N6957, N6065, N3477, N1257);
nand NAND4 (N6960, N6944, N1139, N3500, N1045);
nor NOR2 (N6961, N6948, N4759);
or OR4 (N6962, N6950, N362, N6621, N442);
not NOT1 (N6963, N6958);
and AND2 (N6964, N6959, N131);
buf BUF1 (N6965, N6951);
xor XOR2 (N6966, N6956, N1691);
and AND4 (N6967, N6960, N3384, N4442, N4976);
and AND4 (N6968, N6961, N5711, N941, N1820);
buf BUF1 (N6969, N6965);
nor NOR3 (N6970, N6937, N808, N2375);
and AND2 (N6971, N6963, N564);
nand NAND2 (N6972, N6970, N2517);
xor XOR2 (N6973, N6967, N5534);
nand NAND3 (N6974, N6973, N3911, N424);
or OR4 (N6975, N6966, N4768, N6612, N2260);
not NOT1 (N6976, N6962);
or OR4 (N6977, N6976, N4888, N754, N465);
or OR3 (N6978, N6974, N1488, N986);
not NOT1 (N6979, N6940);
not NOT1 (N6980, N6964);
or OR2 (N6981, N6969, N3802);
and AND4 (N6982, N6981, N5877, N4318, N6514);
xor XOR2 (N6983, N6977, N951);
nor NOR3 (N6984, N6980, N3919, N3803);
buf BUF1 (N6985, N6982);
not NOT1 (N6986, N6985);
xor XOR2 (N6987, N6978, N3244);
and AND4 (N6988, N6983, N3575, N1183, N6492);
xor XOR2 (N6989, N6971, N5575);
and AND2 (N6990, N6987, N246);
not NOT1 (N6991, N6986);
buf BUF1 (N6992, N6954);
not NOT1 (N6993, N6988);
nor NOR3 (N6994, N6990, N3150, N6861);
and AND4 (N6995, N6975, N962, N2223, N1171);
and AND3 (N6996, N6994, N979, N4502);
nor NOR3 (N6997, N6992, N6643, N2434);
or OR2 (N6998, N6993, N1368);
nor NOR4 (N6999, N6998, N4647, N4724, N3668);
nand NAND2 (N7000, N6972, N6981);
not NOT1 (N7001, N6999);
and AND4 (N7002, N6996, N6448, N1015, N5917);
xor XOR2 (N7003, N7002, N422);
nand NAND4 (N7004, N6997, N1526, N5248, N4261);
nor NOR4 (N7005, N6984, N5350, N5749, N3252);
nor NOR2 (N7006, N7005, N1957);
xor XOR2 (N7007, N6995, N3496);
and AND3 (N7008, N7000, N2423, N6274);
not NOT1 (N7009, N7004);
nor NOR4 (N7010, N6991, N189, N3938, N1639);
nor NOR4 (N7011, N7007, N5998, N3070, N4537);
buf BUF1 (N7012, N7009);
not NOT1 (N7013, N7003);
nor NOR4 (N7014, N7001, N3791, N3962, N3705);
not NOT1 (N7015, N7006);
not NOT1 (N7016, N7008);
or OR2 (N7017, N7012, N3107);
and AND4 (N7018, N7015, N1762, N2910, N958);
xor XOR2 (N7019, N7010, N5092);
nor NOR4 (N7020, N7019, N3956, N3479, N1913);
and AND3 (N7021, N7018, N4992, N2775);
not NOT1 (N7022, N7017);
xor XOR2 (N7023, N7022, N1485);
not NOT1 (N7024, N6979);
xor XOR2 (N7025, N7024, N3161);
xor XOR2 (N7026, N7014, N5408);
nor NOR2 (N7027, N7021, N1439);
not NOT1 (N7028, N7013);
nor NOR4 (N7029, N7011, N3063, N797, N4542);
nor NOR2 (N7030, N7020, N1313);
nand NAND2 (N7031, N7029, N3591);
not NOT1 (N7032, N7023);
buf BUF1 (N7033, N7027);
buf BUF1 (N7034, N7030);
buf BUF1 (N7035, N7016);
nand NAND2 (N7036, N6989, N4978);
xor XOR2 (N7037, N7032, N1787);
xor XOR2 (N7038, N7025, N3712);
nand NAND4 (N7039, N7031, N2840, N6154, N1227);
nand NAND4 (N7040, N7034, N2207, N6050, N3591);
or OR4 (N7041, N7040, N4715, N5888, N3384);
and AND4 (N7042, N7033, N4576, N3016, N2841);
not NOT1 (N7043, N7039);
buf BUF1 (N7044, N7026);
nand NAND4 (N7045, N7036, N2390, N4418, N5680);
buf BUF1 (N7046, N7043);
buf BUF1 (N7047, N6968);
nand NAND2 (N7048, N7041, N1116);
and AND2 (N7049, N7047, N4153);
buf BUF1 (N7050, N7035);
or OR4 (N7051, N7042, N4169, N1764, N5566);
nand NAND2 (N7052, N7044, N4695);
not NOT1 (N7053, N7028);
or OR2 (N7054, N7050, N6463);
buf BUF1 (N7055, N7046);
or OR4 (N7056, N7055, N1559, N5600, N256);
buf BUF1 (N7057, N7049);
not NOT1 (N7058, N7051);
nor NOR2 (N7059, N7057, N5372);
nor NOR3 (N7060, N7056, N5113, N1482);
buf BUF1 (N7061, N7060);
buf BUF1 (N7062, N7052);
nor NOR2 (N7063, N7037, N1152);
xor XOR2 (N7064, N7053, N6578);
and AND3 (N7065, N7045, N6334, N3888);
and AND4 (N7066, N7048, N4777, N6689, N2108);
or OR3 (N7067, N7061, N7058, N4954);
buf BUF1 (N7068, N5481);
buf BUF1 (N7069, N7067);
nor NOR3 (N7070, N7063, N6651, N4057);
xor XOR2 (N7071, N7065, N6385);
not NOT1 (N7072, N7066);
not NOT1 (N7073, N7062);
xor XOR2 (N7074, N7070, N4407);
or OR4 (N7075, N7059, N2375, N3237, N5032);
and AND4 (N7076, N7054, N4115, N358, N3976);
buf BUF1 (N7077, N7075);
nand NAND3 (N7078, N7076, N4304, N7012);
xor XOR2 (N7079, N7071, N5451);
or OR2 (N7080, N7072, N2640);
xor XOR2 (N7081, N7074, N7022);
and AND4 (N7082, N7077, N2834, N6575, N1657);
and AND4 (N7083, N7078, N6178, N2993, N4267);
buf BUF1 (N7084, N7073);
xor XOR2 (N7085, N7082, N925);
nand NAND2 (N7086, N7085, N212);
or OR4 (N7087, N7069, N2307, N3887, N5032);
nor NOR3 (N7088, N7038, N2838, N5224);
not NOT1 (N7089, N7080);
not NOT1 (N7090, N7064);
and AND3 (N7091, N7084, N5287, N6888);
xor XOR2 (N7092, N7081, N1499);
and AND2 (N7093, N7079, N4212);
nand NAND2 (N7094, N7086, N2885);
or OR3 (N7095, N7091, N3553, N5124);
and AND4 (N7096, N7083, N4650, N3846, N205);
not NOT1 (N7097, N7088);
nor NOR3 (N7098, N7094, N3466, N4105);
not NOT1 (N7099, N7087);
or OR4 (N7100, N7090, N3172, N1760, N4160);
xor XOR2 (N7101, N7068, N6937);
nand NAND4 (N7102, N7095, N528, N5770, N2785);
nand NAND2 (N7103, N7092, N842);
nand NAND4 (N7104, N7101, N917, N5138, N1734);
not NOT1 (N7105, N7104);
xor XOR2 (N7106, N7103, N5000);
xor XOR2 (N7107, N7100, N1184);
nor NOR4 (N7108, N7106, N1321, N3186, N1891);
and AND2 (N7109, N7093, N3161);
and AND2 (N7110, N7096, N1438);
not NOT1 (N7111, N7109);
and AND2 (N7112, N7110, N3906);
nor NOR3 (N7113, N7098, N1911, N1717);
and AND4 (N7114, N7102, N5023, N2757, N6405);
and AND2 (N7115, N7112, N3162);
buf BUF1 (N7116, N7089);
buf BUF1 (N7117, N7099);
nor NOR3 (N7118, N7116, N3365, N2090);
buf BUF1 (N7119, N7114);
nor NOR2 (N7120, N7108, N1285);
or OR4 (N7121, N7120, N1876, N6091, N1163);
nor NOR2 (N7122, N7115, N5432);
nor NOR2 (N7123, N7105, N2827);
or OR2 (N7124, N7118, N5266);
or OR4 (N7125, N7119, N3383, N6280, N3236);
nand NAND4 (N7126, N7121, N3260, N1594, N1911);
not NOT1 (N7127, N7097);
xor XOR2 (N7128, N7124, N801);
nor NOR4 (N7129, N7127, N971, N2516, N5032);
or OR4 (N7130, N7113, N5899, N1888, N3690);
buf BUF1 (N7131, N7126);
xor XOR2 (N7132, N7107, N5908);
and AND2 (N7133, N7125, N1740);
nand NAND2 (N7134, N7122, N5444);
xor XOR2 (N7135, N7123, N2398);
nor NOR3 (N7136, N7129, N5282, N3531);
or OR2 (N7137, N7136, N2247);
nor NOR2 (N7138, N7137, N4980);
and AND3 (N7139, N7133, N4027, N6205);
nand NAND3 (N7140, N7134, N2152, N6824);
nor NOR4 (N7141, N7140, N269, N1857, N3848);
not NOT1 (N7142, N7138);
nor NOR3 (N7143, N7111, N2982, N5149);
or OR4 (N7144, N7143, N3588, N5281, N6602);
or OR2 (N7145, N7142, N500);
nand NAND2 (N7146, N7144, N6676);
nand NAND4 (N7147, N7132, N4505, N6941, N994);
buf BUF1 (N7148, N7117);
not NOT1 (N7149, N7146);
xor XOR2 (N7150, N7130, N4107);
buf BUF1 (N7151, N7128);
xor XOR2 (N7152, N7131, N7055);
buf BUF1 (N7153, N7135);
or OR2 (N7154, N7145, N2636);
or OR4 (N7155, N7148, N1600, N6868, N3947);
xor XOR2 (N7156, N7154, N2432);
nor NOR2 (N7157, N7156, N2058);
nand NAND3 (N7158, N7157, N4127, N74);
or OR4 (N7159, N7147, N5068, N3531, N6373);
not NOT1 (N7160, N7139);
nand NAND4 (N7161, N7152, N4074, N6072, N351);
not NOT1 (N7162, N7141);
nand NAND4 (N7163, N7153, N4725, N3521, N32);
nand NAND3 (N7164, N7155, N1862, N1624);
nand NAND4 (N7165, N7160, N4348, N4322, N1833);
nor NOR3 (N7166, N7161, N6826, N5271);
and AND2 (N7167, N7159, N1817);
and AND4 (N7168, N7167, N4537, N256, N7164);
buf BUF1 (N7169, N5929);
not NOT1 (N7170, N7151);
nor NOR2 (N7171, N7166, N3731);
not NOT1 (N7172, N7171);
or OR4 (N7173, N7168, N3702, N5768, N5085);
and AND3 (N7174, N7158, N1772, N816);
nor NOR2 (N7175, N7162, N716);
not NOT1 (N7176, N7173);
or OR4 (N7177, N7149, N206, N1433, N2103);
buf BUF1 (N7178, N7175);
nand NAND2 (N7179, N7178, N5658);
not NOT1 (N7180, N7177);
not NOT1 (N7181, N7180);
nor NOR3 (N7182, N7174, N3747, N1234);
and AND4 (N7183, N7176, N1946, N3161, N2187);
and AND2 (N7184, N7172, N6765);
buf BUF1 (N7185, N7169);
and AND4 (N7186, N7163, N1112, N6374, N4638);
xor XOR2 (N7187, N7170, N1047);
nor NOR3 (N7188, N7182, N6828, N5409);
nor NOR4 (N7189, N7188, N276, N5914, N5428);
not NOT1 (N7190, N7165);
and AND3 (N7191, N7186, N2989, N4847);
and AND4 (N7192, N7184, N3737, N1036, N3106);
or OR4 (N7193, N7189, N7064, N2541, N2609);
nand NAND4 (N7194, N7191, N5001, N4541, N3370);
and AND3 (N7195, N7179, N4995, N3903);
nand NAND4 (N7196, N7195, N2586, N948, N5596);
nand NAND4 (N7197, N7192, N144, N811, N3391);
xor XOR2 (N7198, N7185, N4309);
and AND4 (N7199, N7194, N2934, N1777, N2440);
buf BUF1 (N7200, N7193);
xor XOR2 (N7201, N7181, N5090);
nand NAND3 (N7202, N7183, N2910, N6884);
buf BUF1 (N7203, N7190);
xor XOR2 (N7204, N7199, N4541);
buf BUF1 (N7205, N7187);
xor XOR2 (N7206, N7203, N2932);
not NOT1 (N7207, N7206);
nor NOR4 (N7208, N7207, N1400, N3492, N2059);
nand NAND4 (N7209, N7196, N4659, N80, N4694);
nor NOR2 (N7210, N7200, N669);
or OR2 (N7211, N7197, N5643);
buf BUF1 (N7212, N7202);
not NOT1 (N7213, N7205);
and AND4 (N7214, N7150, N4933, N5765, N1168);
nor NOR4 (N7215, N7198, N6433, N3912, N6309);
buf BUF1 (N7216, N7210);
buf BUF1 (N7217, N7215);
and AND3 (N7218, N7213, N7201, N1235);
or OR2 (N7219, N2301, N1504);
and AND2 (N7220, N7208, N3447);
and AND2 (N7221, N7209, N3767);
and AND4 (N7222, N7218, N5435, N1710, N3894);
nor NOR4 (N7223, N7221, N1237, N5535, N5250);
nand NAND3 (N7224, N7219, N2655, N7146);
nand NAND3 (N7225, N7212, N2612, N1691);
nand NAND3 (N7226, N7222, N325, N5539);
buf BUF1 (N7227, N7226);
and AND4 (N7228, N7211, N6222, N3622, N4942);
xor XOR2 (N7229, N7214, N3296);
not NOT1 (N7230, N7229);
nand NAND3 (N7231, N7228, N1400, N2596);
nor NOR3 (N7232, N7220, N580, N5475);
or OR2 (N7233, N7204, N3004);
nand NAND3 (N7234, N7224, N6941, N146);
not NOT1 (N7235, N7234);
and AND3 (N7236, N7233, N4968, N6651);
and AND4 (N7237, N7235, N2478, N5571, N5833);
or OR2 (N7238, N7223, N3036);
xor XOR2 (N7239, N7236, N2001);
not NOT1 (N7240, N7239);
nor NOR2 (N7241, N7231, N2864);
and AND2 (N7242, N7238, N6335);
or OR4 (N7243, N7242, N5833, N3174, N2557);
nand NAND3 (N7244, N7225, N6475, N974);
nor NOR4 (N7245, N7244, N1937, N1890, N6661);
xor XOR2 (N7246, N7216, N2496);
nand NAND4 (N7247, N7232, N3067, N5421, N4853);
or OR3 (N7248, N7243, N5013, N6460);
and AND4 (N7249, N7248, N2297, N6064, N7146);
not NOT1 (N7250, N7217);
nor NOR3 (N7251, N7249, N4453, N698);
xor XOR2 (N7252, N7250, N4029);
or OR3 (N7253, N7241, N1139, N3505);
buf BUF1 (N7254, N7247);
buf BUF1 (N7255, N7251);
or OR3 (N7256, N7237, N4356, N3547);
not NOT1 (N7257, N7240);
nand NAND3 (N7258, N7256, N2292, N1916);
buf BUF1 (N7259, N7230);
nor NOR2 (N7260, N7254, N3922);
buf BUF1 (N7261, N7259);
not NOT1 (N7262, N7252);
or OR3 (N7263, N7255, N2640, N955);
nor NOR3 (N7264, N7261, N6341, N3756);
and AND3 (N7265, N7227, N6590, N4979);
and AND2 (N7266, N7262, N383);
or OR3 (N7267, N7263, N3035, N6008);
nand NAND4 (N7268, N7267, N1319, N2005, N4638);
nand NAND3 (N7269, N7258, N2595, N6122);
xor XOR2 (N7270, N7266, N1344);
or OR2 (N7271, N7253, N828);
nand NAND2 (N7272, N7260, N6973);
nand NAND2 (N7273, N7264, N943);
buf BUF1 (N7274, N7265);
and AND4 (N7275, N7270, N4820, N1641, N4206);
and AND2 (N7276, N7275, N1945);
or OR4 (N7277, N7257, N4030, N6743, N5718);
nand NAND2 (N7278, N7273, N377);
nor NOR4 (N7279, N7246, N2112, N4128, N6363);
nand NAND4 (N7280, N7277, N5370, N7257, N4245);
nand NAND2 (N7281, N7276, N4669);
or OR3 (N7282, N7272, N5480, N831);
nor NOR3 (N7283, N7271, N2209, N2231);
or OR2 (N7284, N7274, N3260);
and AND4 (N7285, N7269, N2405, N906, N140);
not NOT1 (N7286, N7279);
xor XOR2 (N7287, N7268, N3113);
or OR2 (N7288, N7280, N869);
and AND4 (N7289, N7288, N5077, N6779, N6223);
buf BUF1 (N7290, N7289);
nand NAND3 (N7291, N7287, N793, N4589);
or OR3 (N7292, N7286, N5317, N847);
nand NAND3 (N7293, N7292, N7127, N4289);
xor XOR2 (N7294, N7278, N1773);
buf BUF1 (N7295, N7283);
buf BUF1 (N7296, N7295);
nand NAND4 (N7297, N7291, N2934, N5764, N3715);
and AND4 (N7298, N7293, N1945, N5703, N6437);
nor NOR4 (N7299, N7245, N3370, N6982, N5197);
or OR3 (N7300, N7299, N1409, N2343);
not NOT1 (N7301, N7282);
not NOT1 (N7302, N7300);
or OR3 (N7303, N7297, N3524, N1554);
nor NOR4 (N7304, N7301, N6065, N1769, N4549);
nand NAND4 (N7305, N7296, N1018, N621, N3477);
not NOT1 (N7306, N7298);
nor NOR2 (N7307, N7285, N1996);
buf BUF1 (N7308, N7303);
nor NOR3 (N7309, N7308, N2053, N1953);
buf BUF1 (N7310, N7294);
nand NAND4 (N7311, N7306, N4108, N3837, N7000);
nand NAND2 (N7312, N7284, N5265);
or OR4 (N7313, N7311, N2223, N698, N4690);
xor XOR2 (N7314, N7313, N4818);
nand NAND2 (N7315, N7307, N2783);
nand NAND4 (N7316, N7305, N3235, N4283, N2451);
and AND2 (N7317, N7314, N4103);
or OR4 (N7318, N7309, N1679, N4528, N3531);
not NOT1 (N7319, N7312);
xor XOR2 (N7320, N7304, N3764);
xor XOR2 (N7321, N7315, N5010);
xor XOR2 (N7322, N7320, N3396);
nor NOR4 (N7323, N7321, N1434, N4181, N4009);
buf BUF1 (N7324, N7322);
not NOT1 (N7325, N7319);
buf BUF1 (N7326, N7317);
not NOT1 (N7327, N7310);
nor NOR3 (N7328, N7290, N5674, N6218);
nor NOR3 (N7329, N7318, N7293, N1);
xor XOR2 (N7330, N7325, N1396);
or OR3 (N7331, N7281, N1205, N6796);
nor NOR4 (N7332, N7302, N2962, N5228, N4366);
or OR4 (N7333, N7324, N702, N1314, N984);
or OR2 (N7334, N7328, N6832);
buf BUF1 (N7335, N7330);
nor NOR4 (N7336, N7332, N2521, N2234, N3175);
buf BUF1 (N7337, N7336);
nor NOR3 (N7338, N7323, N4400, N4708);
buf BUF1 (N7339, N7327);
nor NOR2 (N7340, N7334, N6081);
and AND3 (N7341, N7326, N364, N7048);
not NOT1 (N7342, N7329);
or OR4 (N7343, N7339, N6086, N6246, N5614);
and AND4 (N7344, N7341, N6292, N3851, N4300);
nand NAND2 (N7345, N7343, N3162);
not NOT1 (N7346, N7344);
buf BUF1 (N7347, N7342);
nor NOR2 (N7348, N7347, N5163);
or OR2 (N7349, N7331, N4417);
nor NOR3 (N7350, N7345, N1288, N3269);
buf BUF1 (N7351, N7340);
xor XOR2 (N7352, N7348, N182);
or OR2 (N7353, N7346, N5537);
nor NOR2 (N7354, N7351, N4642);
nand NAND2 (N7355, N7335, N1062);
not NOT1 (N7356, N7349);
and AND2 (N7357, N7316, N5674);
xor XOR2 (N7358, N7354, N2030);
and AND3 (N7359, N7353, N1759, N1444);
nand NAND4 (N7360, N7357, N1019, N6057, N3685);
xor XOR2 (N7361, N7360, N6758);
nand NAND2 (N7362, N7361, N5055);
not NOT1 (N7363, N7358);
nand NAND2 (N7364, N7362, N4220);
nand NAND2 (N7365, N7333, N2985);
nor NOR3 (N7366, N7365, N1680, N4719);
and AND4 (N7367, N7366, N756, N7144, N848);
and AND3 (N7368, N7337, N4533, N794);
or OR4 (N7369, N7352, N1516, N6804, N5621);
or OR2 (N7370, N7359, N4780);
nand NAND3 (N7371, N7355, N3180, N7230);
buf BUF1 (N7372, N7371);
and AND4 (N7373, N7369, N1149, N4407, N3218);
and AND4 (N7374, N7350, N2264, N4063, N35);
buf BUF1 (N7375, N7368);
nor NOR4 (N7376, N7364, N5153, N5318, N7231);
nand NAND3 (N7377, N7356, N4502, N221);
buf BUF1 (N7378, N7374);
nor NOR4 (N7379, N7363, N345, N5118, N1688);
nand NAND4 (N7380, N7379, N2804, N1560, N4250);
xor XOR2 (N7381, N7372, N1806);
not NOT1 (N7382, N7376);
and AND4 (N7383, N7338, N6424, N719, N4175);
buf BUF1 (N7384, N7370);
not NOT1 (N7385, N7382);
and AND4 (N7386, N7385, N5965, N5000, N1953);
buf BUF1 (N7387, N7377);
and AND2 (N7388, N7381, N6549);
xor XOR2 (N7389, N7387, N5721);
or OR3 (N7390, N7367, N1268, N5092);
nor NOR4 (N7391, N7388, N5633, N2799, N2299);
or OR3 (N7392, N7378, N5191, N1855);
nand NAND4 (N7393, N7391, N2030, N4099, N5745);
or OR3 (N7394, N7389, N7200, N2683);
buf BUF1 (N7395, N7392);
buf BUF1 (N7396, N7383);
or OR3 (N7397, N7394, N120, N4589);
nor NOR3 (N7398, N7386, N1555, N1240);
nand NAND4 (N7399, N7393, N5679, N4694, N4250);
nor NOR4 (N7400, N7375, N1832, N5589, N3654);
and AND4 (N7401, N7384, N2847, N3787, N1162);
buf BUF1 (N7402, N7390);
buf BUF1 (N7403, N7399);
nor NOR2 (N7404, N7403, N3503);
buf BUF1 (N7405, N7404);
xor XOR2 (N7406, N7401, N3312);
and AND3 (N7407, N7397, N4038, N173);
xor XOR2 (N7408, N7380, N3419);
nor NOR4 (N7409, N7400, N4702, N6799, N6681);
nor NOR3 (N7410, N7407, N1960, N5341);
nand NAND2 (N7411, N7373, N1404);
buf BUF1 (N7412, N7410);
buf BUF1 (N7413, N7402);
and AND2 (N7414, N7398, N4082);
and AND2 (N7415, N7396, N5453);
and AND4 (N7416, N7408, N5128, N7098, N4079);
or OR3 (N7417, N7405, N4475, N4413);
buf BUF1 (N7418, N7411);
buf BUF1 (N7419, N7413);
buf BUF1 (N7420, N7414);
and AND4 (N7421, N7418, N4817, N51, N5491);
and AND2 (N7422, N7416, N4694);
nor NOR4 (N7423, N7409, N2548, N3201, N2859);
buf BUF1 (N7424, N7423);
xor XOR2 (N7425, N7419, N941);
buf BUF1 (N7426, N7424);
and AND2 (N7427, N7415, N576);
xor XOR2 (N7428, N7425, N962);
nand NAND3 (N7429, N7421, N6030, N5411);
nand NAND2 (N7430, N7406, N373);
or OR4 (N7431, N7395, N6799, N6634, N6757);
and AND2 (N7432, N7417, N4490);
xor XOR2 (N7433, N7426, N35);
and AND4 (N7434, N7412, N550, N3911, N3664);
and AND3 (N7435, N7428, N5436, N6383);
and AND3 (N7436, N7422, N3731, N6460);
or OR4 (N7437, N7432, N1603, N2560, N1447);
not NOT1 (N7438, N7436);
or OR2 (N7439, N7431, N3969);
nand NAND4 (N7440, N7420, N242, N6246, N1404);
not NOT1 (N7441, N7435);
or OR2 (N7442, N7433, N3253);
nor NOR3 (N7443, N7437, N6321, N5057);
nand NAND4 (N7444, N7443, N5606, N5528, N7296);
and AND4 (N7445, N7438, N6485, N2764, N2707);
nand NAND2 (N7446, N7430, N1747);
xor XOR2 (N7447, N7434, N107);
or OR3 (N7448, N7444, N1954, N124);
nand NAND2 (N7449, N7429, N2566);
xor XOR2 (N7450, N7442, N5269);
xor XOR2 (N7451, N7450, N2116);
buf BUF1 (N7452, N7447);
and AND3 (N7453, N7445, N368, N986);
not NOT1 (N7454, N7449);
and AND2 (N7455, N7453, N4802);
or OR4 (N7456, N7455, N4024, N4655, N3781);
or OR4 (N7457, N7446, N5497, N7005, N4900);
or OR4 (N7458, N7454, N3385, N2928, N5757);
not NOT1 (N7459, N7439);
xor XOR2 (N7460, N7456, N7118);
buf BUF1 (N7461, N7441);
not NOT1 (N7462, N7458);
xor XOR2 (N7463, N7460, N734);
nor NOR2 (N7464, N7448, N960);
and AND4 (N7465, N7440, N3224, N6824, N4100);
xor XOR2 (N7466, N7459, N804);
nand NAND2 (N7467, N7452, N6439);
or OR3 (N7468, N7465, N494, N5294);
buf BUF1 (N7469, N7462);
or OR4 (N7470, N7467, N6951, N2511, N2010);
and AND2 (N7471, N7464, N1706);
nor NOR3 (N7472, N7471, N2622, N6260);
nor NOR3 (N7473, N7472, N4738, N4402);
and AND4 (N7474, N7473, N837, N6628, N1804);
or OR4 (N7475, N7463, N4567, N95, N6823);
xor XOR2 (N7476, N7427, N1580);
or OR3 (N7477, N7461, N2796, N772);
xor XOR2 (N7478, N7475, N1163);
and AND4 (N7479, N7457, N5758, N7058, N6028);
xor XOR2 (N7480, N7470, N6116);
or OR2 (N7481, N7474, N5354);
and AND4 (N7482, N7477, N31, N1465, N954);
and AND4 (N7483, N7478, N493, N138, N1233);
nand NAND2 (N7484, N7483, N1891);
or OR2 (N7485, N7484, N5905);
and AND2 (N7486, N7479, N5350);
buf BUF1 (N7487, N7481);
or OR4 (N7488, N7485, N491, N290, N1418);
buf BUF1 (N7489, N7480);
nor NOR2 (N7490, N7488, N6177);
and AND4 (N7491, N7490, N253, N3350, N4222);
not NOT1 (N7492, N7451);
buf BUF1 (N7493, N7492);
buf BUF1 (N7494, N7482);
nor NOR4 (N7495, N7491, N732, N7326, N6325);
or OR2 (N7496, N7469, N3064);
xor XOR2 (N7497, N7468, N3624);
nor NOR2 (N7498, N7489, N1348);
nor NOR4 (N7499, N7476, N537, N4660, N4807);
not NOT1 (N7500, N7466);
nand NAND2 (N7501, N7486, N5161);
xor XOR2 (N7502, N7493, N4565);
not NOT1 (N7503, N7494);
xor XOR2 (N7504, N7503, N6881);
not NOT1 (N7505, N7498);
xor XOR2 (N7506, N7505, N1428);
nor NOR3 (N7507, N7504, N4719, N1662);
or OR3 (N7508, N7500, N1008, N6951);
xor XOR2 (N7509, N7506, N4136);
xor XOR2 (N7510, N7507, N7267);
not NOT1 (N7511, N7497);
nand NAND2 (N7512, N7499, N5300);
nand NAND4 (N7513, N7495, N1538, N5683, N3838);
xor XOR2 (N7514, N7502, N1838);
and AND3 (N7515, N7511, N3933, N6969);
or OR4 (N7516, N7501, N3769, N4726, N5351);
not NOT1 (N7517, N7487);
and AND2 (N7518, N7513, N3092);
and AND4 (N7519, N7515, N5098, N2374, N2708);
nor NOR2 (N7520, N7514, N6196);
or OR4 (N7521, N7517, N2682, N4241, N3708);
buf BUF1 (N7522, N7520);
nand NAND2 (N7523, N7521, N5688);
and AND2 (N7524, N7510, N1434);
not NOT1 (N7525, N7524);
not NOT1 (N7526, N7522);
xor XOR2 (N7527, N7509, N1702);
nor NOR4 (N7528, N7526, N4393, N456, N6145);
nand NAND4 (N7529, N7496, N3697, N5352, N1998);
nor NOR2 (N7530, N7512, N4905);
or OR3 (N7531, N7519, N1700, N1625);
nor NOR2 (N7532, N7523, N3009);
xor XOR2 (N7533, N7532, N1837);
and AND3 (N7534, N7528, N2857, N1071);
not NOT1 (N7535, N7533);
or OR2 (N7536, N7518, N2004);
and AND2 (N7537, N7531, N7084);
or OR3 (N7538, N7525, N6391, N144);
nor NOR4 (N7539, N7516, N2629, N4832, N2417);
buf BUF1 (N7540, N7527);
nor NOR2 (N7541, N7508, N1275);
buf BUF1 (N7542, N7539);
nor NOR3 (N7543, N7530, N6068, N1950);
nor NOR2 (N7544, N7541, N5617);
buf BUF1 (N7545, N7534);
nand NAND4 (N7546, N7540, N5710, N1795, N6014);
nand NAND3 (N7547, N7538, N2829, N922);
and AND4 (N7548, N7529, N2424, N6051, N1997);
or OR3 (N7549, N7547, N7472, N6767);
and AND2 (N7550, N7545, N6977);
and AND4 (N7551, N7543, N2836, N6410, N40);
xor XOR2 (N7552, N7546, N1789);
or OR4 (N7553, N7549, N2884, N85, N7243);
xor XOR2 (N7554, N7550, N1082);
and AND3 (N7555, N7553, N7295, N3671);
buf BUF1 (N7556, N7542);
nor NOR4 (N7557, N7544, N4330, N973, N5825);
xor XOR2 (N7558, N7535, N353);
and AND3 (N7559, N7558, N5210, N2505);
buf BUF1 (N7560, N7559);
not NOT1 (N7561, N7551);
and AND2 (N7562, N7556, N5495);
not NOT1 (N7563, N7548);
and AND3 (N7564, N7560, N3403, N831);
and AND2 (N7565, N7564, N4349);
nor NOR2 (N7566, N7563, N7065);
buf BUF1 (N7567, N7562);
and AND2 (N7568, N7566, N7328);
buf BUF1 (N7569, N7536);
xor XOR2 (N7570, N7557, N2566);
and AND2 (N7571, N7554, N1302);
xor XOR2 (N7572, N7565, N339);
and AND3 (N7573, N7555, N6796, N4996);
not NOT1 (N7574, N7567);
buf BUF1 (N7575, N7574);
and AND3 (N7576, N7571, N3795, N382);
xor XOR2 (N7577, N7552, N2750);
or OR3 (N7578, N7572, N2733, N2136);
nand NAND2 (N7579, N7578, N4979);
or OR3 (N7580, N7569, N1010, N6688);
nand NAND3 (N7581, N7575, N6131, N904);
xor XOR2 (N7582, N7573, N3715);
nor NOR4 (N7583, N7568, N7036, N1458, N6785);
buf BUF1 (N7584, N7581);
buf BUF1 (N7585, N7577);
xor XOR2 (N7586, N7583, N1626);
buf BUF1 (N7587, N7579);
not NOT1 (N7588, N7580);
or OR3 (N7589, N7584, N1638, N5095);
nand NAND3 (N7590, N7570, N4115, N4576);
nand NAND2 (N7591, N7587, N2925);
buf BUF1 (N7592, N7591);
nor NOR3 (N7593, N7585, N1720, N6015);
or OR2 (N7594, N7593, N5749);
nand NAND3 (N7595, N7594, N4732, N2718);
not NOT1 (N7596, N7537);
buf BUF1 (N7597, N7590);
and AND2 (N7598, N7576, N2213);
xor XOR2 (N7599, N7597, N7208);
buf BUF1 (N7600, N7561);
or OR3 (N7601, N7599, N2762, N2858);
buf BUF1 (N7602, N7601);
and AND3 (N7603, N7595, N1574, N6763);
not NOT1 (N7604, N7600);
or OR2 (N7605, N7603, N718);
nand NAND2 (N7606, N7582, N6513);
not NOT1 (N7607, N7592);
not NOT1 (N7608, N7586);
or OR2 (N7609, N7598, N3855);
nor NOR3 (N7610, N7589, N4915, N2611);
nand NAND4 (N7611, N7610, N4502, N7058, N1755);
or OR3 (N7612, N7606, N7387, N2159);
nor NOR2 (N7613, N7604, N3571);
xor XOR2 (N7614, N7607, N4640);
xor XOR2 (N7615, N7588, N3494);
nor NOR2 (N7616, N7605, N2700);
not NOT1 (N7617, N7615);
not NOT1 (N7618, N7616);
xor XOR2 (N7619, N7612, N5352);
nor NOR2 (N7620, N7602, N1601);
nor NOR2 (N7621, N7611, N872);
xor XOR2 (N7622, N7609, N4378);
buf BUF1 (N7623, N7608);
not NOT1 (N7624, N7623);
nor NOR4 (N7625, N7622, N775, N1357, N5726);
xor XOR2 (N7626, N7624, N2250);
or OR2 (N7627, N7618, N989);
buf BUF1 (N7628, N7596);
buf BUF1 (N7629, N7619);
nand NAND3 (N7630, N7614, N7184, N3875);
buf BUF1 (N7631, N7613);
nand NAND2 (N7632, N7625, N4175);
nand NAND3 (N7633, N7617, N5102, N6885);
buf BUF1 (N7634, N7632);
xor XOR2 (N7635, N7631, N2550);
and AND4 (N7636, N7621, N6178, N3472, N339);
and AND3 (N7637, N7634, N7384, N3851);
nor NOR2 (N7638, N7630, N4703);
nand NAND2 (N7639, N7636, N2968);
buf BUF1 (N7640, N7628);
and AND4 (N7641, N7633, N3511, N6864, N2056);
or OR4 (N7642, N7639, N1980, N2103, N4973);
nand NAND4 (N7643, N7637, N2527, N4934, N1188);
nor NOR2 (N7644, N7635, N6477);
nand NAND4 (N7645, N7627, N2320, N4756, N1628);
xor XOR2 (N7646, N7641, N7357);
buf BUF1 (N7647, N7626);
not NOT1 (N7648, N7629);
not NOT1 (N7649, N7642);
xor XOR2 (N7650, N7643, N992);
nor NOR4 (N7651, N7646, N4014, N775, N3142);
nand NAND2 (N7652, N7651, N6261);
not NOT1 (N7653, N7645);
nor NOR2 (N7654, N7650, N3968);
or OR4 (N7655, N7652, N2240, N4113, N4507);
xor XOR2 (N7656, N7648, N4372);
and AND4 (N7657, N7647, N3955, N7034, N633);
and AND3 (N7658, N7640, N2203, N4345);
xor XOR2 (N7659, N7658, N4920);
xor XOR2 (N7660, N7638, N3545);
xor XOR2 (N7661, N7644, N6796);
buf BUF1 (N7662, N7657);
not NOT1 (N7663, N7649);
not NOT1 (N7664, N7660);
nand NAND3 (N7665, N7662, N3089, N125);
nor NOR2 (N7666, N7653, N7290);
nor NOR3 (N7667, N7665, N4066, N6128);
xor XOR2 (N7668, N7620, N1731);
xor XOR2 (N7669, N7666, N1534);
nor NOR3 (N7670, N7661, N1989, N5337);
and AND3 (N7671, N7669, N6382, N1502);
buf BUF1 (N7672, N7664);
nor NOR4 (N7673, N7668, N548, N2964, N5058);
buf BUF1 (N7674, N7663);
and AND4 (N7675, N7671, N2138, N2048, N996);
nor NOR3 (N7676, N7674, N2711, N6779);
and AND4 (N7677, N7670, N3448, N85, N1431);
nand NAND4 (N7678, N7659, N7646, N455, N4863);
or OR3 (N7679, N7678, N7187, N5358);
nor NOR2 (N7680, N7675, N3986);
and AND3 (N7681, N7654, N6053, N3177);
buf BUF1 (N7682, N7655);
buf BUF1 (N7683, N7680);
and AND4 (N7684, N7673, N5326, N1110, N4589);
and AND4 (N7685, N7683, N1677, N2060, N311);
buf BUF1 (N7686, N7672);
and AND4 (N7687, N7684, N7274, N3369, N1505);
and AND3 (N7688, N7682, N2636, N6470);
nor NOR3 (N7689, N7667, N4327, N3078);
not NOT1 (N7690, N7679);
and AND4 (N7691, N7686, N1733, N1246, N3929);
or OR2 (N7692, N7685, N5546);
not NOT1 (N7693, N7691);
nand NAND2 (N7694, N7676, N1640);
buf BUF1 (N7695, N7687);
and AND4 (N7696, N7681, N2257, N2891, N4565);
nand NAND4 (N7697, N7694, N2832, N543, N1474);
xor XOR2 (N7698, N7689, N2342);
and AND2 (N7699, N7688, N6699);
buf BUF1 (N7700, N7693);
not NOT1 (N7701, N7695);
xor XOR2 (N7702, N7700, N1109);
not NOT1 (N7703, N7702);
nand NAND2 (N7704, N7699, N1817);
not NOT1 (N7705, N7690);
xor XOR2 (N7706, N7692, N4879);
not NOT1 (N7707, N7677);
nor NOR2 (N7708, N7698, N947);
not NOT1 (N7709, N7701);
not NOT1 (N7710, N7706);
nand NAND2 (N7711, N7696, N189);
xor XOR2 (N7712, N7708, N3389);
and AND2 (N7713, N7656, N737);
and AND4 (N7714, N7704, N2846, N6325, N1684);
and AND4 (N7715, N7705, N5238, N1067, N6094);
not NOT1 (N7716, N7715);
buf BUF1 (N7717, N7712);
not NOT1 (N7718, N7703);
and AND2 (N7719, N7697, N7147);
and AND4 (N7720, N7710, N3032, N7290, N4095);
or OR4 (N7721, N7711, N5772, N1464, N7654);
buf BUF1 (N7722, N7720);
nor NOR3 (N7723, N7707, N5309, N7366);
and AND2 (N7724, N7721, N5739);
or OR3 (N7725, N7718, N1133, N3396);
nor NOR3 (N7726, N7722, N5210, N262);
and AND3 (N7727, N7709, N4251, N412);
nor NOR2 (N7728, N7723, N322);
nand NAND3 (N7729, N7716, N4846, N4154);
nor NOR3 (N7730, N7714, N3194, N6379);
buf BUF1 (N7731, N7727);
not NOT1 (N7732, N7729);
buf BUF1 (N7733, N7724);
not NOT1 (N7734, N7728);
or OR3 (N7735, N7734, N4933, N4542);
nand NAND4 (N7736, N7713, N7611, N5398, N3757);
nor NOR2 (N7737, N7717, N3260);
buf BUF1 (N7738, N7730);
nand NAND3 (N7739, N7731, N1584, N5456);
nand NAND3 (N7740, N7733, N756, N1127);
nand NAND4 (N7741, N7740, N7514, N6013, N5078);
nor NOR3 (N7742, N7736, N6138, N4282);
nand NAND2 (N7743, N7739, N7716);
and AND2 (N7744, N7741, N7050);
not NOT1 (N7745, N7737);
xor XOR2 (N7746, N7743, N4507);
nor NOR3 (N7747, N7738, N4598, N5238);
and AND3 (N7748, N7719, N1716, N1399);
not NOT1 (N7749, N7742);
nor NOR4 (N7750, N7749, N2638, N5891, N6736);
xor XOR2 (N7751, N7744, N1610);
xor XOR2 (N7752, N7747, N3378);
nor NOR3 (N7753, N7750, N2383, N6077);
or OR2 (N7754, N7735, N4406);
nand NAND3 (N7755, N7746, N5889, N4908);
buf BUF1 (N7756, N7745);
or OR3 (N7757, N7725, N2015, N4218);
and AND2 (N7758, N7726, N3532);
and AND4 (N7759, N7748, N3028, N1368, N1190);
buf BUF1 (N7760, N7751);
or OR4 (N7761, N7756, N4288, N4640, N4827);
nand NAND4 (N7762, N7761, N5641, N182, N2477);
nor NOR4 (N7763, N7760, N3940, N7055, N1148);
xor XOR2 (N7764, N7762, N3364);
nor NOR2 (N7765, N7763, N6504);
and AND4 (N7766, N7764, N5533, N477, N6640);
nand NAND3 (N7767, N7754, N3365, N6168);
or OR4 (N7768, N7767, N4998, N224, N698);
xor XOR2 (N7769, N7766, N5150);
nor NOR2 (N7770, N7755, N4010);
not NOT1 (N7771, N7732);
or OR2 (N7772, N7771, N7057);
xor XOR2 (N7773, N7753, N4754);
nor NOR4 (N7774, N7759, N1854, N2321, N749);
not NOT1 (N7775, N7765);
nand NAND3 (N7776, N7752, N1986, N5928);
nor NOR2 (N7777, N7757, N5921);
not NOT1 (N7778, N7777);
nand NAND2 (N7779, N7778, N1902);
and AND4 (N7780, N7768, N6889, N2102, N3915);
buf BUF1 (N7781, N7779);
xor XOR2 (N7782, N7776, N3779);
buf BUF1 (N7783, N7769);
not NOT1 (N7784, N7770);
nand NAND2 (N7785, N7775, N6732);
not NOT1 (N7786, N7758);
or OR4 (N7787, N7786, N7581, N6559, N6530);
and AND3 (N7788, N7782, N7608, N3756);
nand NAND3 (N7789, N7788, N2051, N4510);
nand NAND2 (N7790, N7785, N5899);
nor NOR3 (N7791, N7783, N901, N4457);
not NOT1 (N7792, N7791);
not NOT1 (N7793, N7792);
nor NOR2 (N7794, N7790, N7762);
xor XOR2 (N7795, N7773, N849);
xor XOR2 (N7796, N7772, N5082);
and AND4 (N7797, N7780, N5273, N7668, N3954);
not NOT1 (N7798, N7787);
nor NOR2 (N7799, N7798, N5444);
or OR4 (N7800, N7796, N6405, N2685, N4844);
or OR2 (N7801, N7774, N5090);
not NOT1 (N7802, N7793);
xor XOR2 (N7803, N7784, N6976);
and AND4 (N7804, N7789, N2215, N5545, N5625);
not NOT1 (N7805, N7801);
nor NOR2 (N7806, N7805, N7726);
nor NOR3 (N7807, N7795, N1988, N5391);
nand NAND3 (N7808, N7802, N3096, N2557);
or OR4 (N7809, N7794, N882, N2260, N3333);
not NOT1 (N7810, N7809);
buf BUF1 (N7811, N7807);
xor XOR2 (N7812, N7800, N1367);
nor NOR3 (N7813, N7810, N109, N2258);
not NOT1 (N7814, N7806);
nand NAND3 (N7815, N7804, N69, N4389);
buf BUF1 (N7816, N7813);
xor XOR2 (N7817, N7797, N6114);
not NOT1 (N7818, N7814);
nor NOR4 (N7819, N7818, N2224, N3055, N5888);
and AND2 (N7820, N7781, N6191);
not NOT1 (N7821, N7819);
xor XOR2 (N7822, N7816, N2344);
nor NOR2 (N7823, N7817, N5640);
nor NOR4 (N7824, N7803, N400, N181, N2608);
buf BUF1 (N7825, N7824);
nand NAND3 (N7826, N7822, N2810, N5256);
or OR2 (N7827, N7823, N6424);
buf BUF1 (N7828, N7826);
xor XOR2 (N7829, N7799, N287);
nand NAND3 (N7830, N7829, N3647, N807);
nor NOR4 (N7831, N7828, N5014, N389, N737);
buf BUF1 (N7832, N7827);
xor XOR2 (N7833, N7812, N4540);
and AND4 (N7834, N7825, N5458, N7514, N1913);
nor NOR3 (N7835, N7831, N5201, N2215);
nor NOR4 (N7836, N7835, N2014, N4274, N3694);
or OR2 (N7837, N7834, N5235);
buf BUF1 (N7838, N7820);
nand NAND2 (N7839, N7821, N2612);
buf BUF1 (N7840, N7839);
nor NOR3 (N7841, N7832, N2099, N535);
or OR2 (N7842, N7811, N992);
buf BUF1 (N7843, N7837);
or OR3 (N7844, N7838, N6719, N2350);
and AND3 (N7845, N7843, N7283, N4822);
nand NAND3 (N7846, N7842, N3952, N5612);
xor XOR2 (N7847, N7846, N2502);
not NOT1 (N7848, N7836);
not NOT1 (N7849, N7847);
buf BUF1 (N7850, N7840);
xor XOR2 (N7851, N7808, N3184);
or OR3 (N7852, N7851, N6239, N992);
and AND2 (N7853, N7844, N137);
nand NAND3 (N7854, N7850, N5633, N4547);
and AND3 (N7855, N7853, N3345, N929);
or OR4 (N7856, N7848, N968, N3101, N6848);
buf BUF1 (N7857, N7854);
buf BUF1 (N7858, N7833);
or OR2 (N7859, N7855, N6596);
nand NAND4 (N7860, N7859, N4618, N7838, N7103);
buf BUF1 (N7861, N7815);
and AND3 (N7862, N7849, N4480, N4296);
not NOT1 (N7863, N7858);
nor NOR3 (N7864, N7845, N5702, N3537);
nor NOR4 (N7865, N7852, N2456, N288, N4239);
nand NAND4 (N7866, N7841, N5508, N6056, N5106);
xor XOR2 (N7867, N7860, N3354);
nand NAND4 (N7868, N7865, N2230, N4384, N7563);
and AND4 (N7869, N7867, N856, N5846, N6257);
and AND3 (N7870, N7830, N3756, N5233);
buf BUF1 (N7871, N7866);
nand NAND3 (N7872, N7871, N2865, N5271);
or OR2 (N7873, N7868, N3992);
or OR3 (N7874, N7872, N3392, N493);
buf BUF1 (N7875, N7856);
nor NOR3 (N7876, N7864, N4157, N1547);
and AND3 (N7877, N7870, N2459, N3676);
nor NOR4 (N7878, N7877, N4515, N2137, N1670);
or OR3 (N7879, N7857, N4678, N7405);
nor NOR4 (N7880, N7878, N2338, N4182, N1855);
and AND3 (N7881, N7873, N1782, N1948);
nand NAND4 (N7882, N7874, N379, N3352, N5707);
or OR3 (N7883, N7881, N2409, N496);
not NOT1 (N7884, N7861);
nand NAND4 (N7885, N7875, N6619, N5203, N108);
and AND2 (N7886, N7879, N6826);
not NOT1 (N7887, N7882);
nand NAND2 (N7888, N7884, N1171);
or OR4 (N7889, N7883, N5628, N2547, N6201);
not NOT1 (N7890, N7886);
or OR3 (N7891, N7888, N248, N2269);
nand NAND3 (N7892, N7862, N6012, N2925);
or OR3 (N7893, N7889, N3880, N162);
nand NAND2 (N7894, N7887, N7439);
not NOT1 (N7895, N7863);
or OR4 (N7896, N7893, N6648, N6824, N2202);
xor XOR2 (N7897, N7894, N2724);
buf BUF1 (N7898, N7897);
buf BUF1 (N7899, N7895);
not NOT1 (N7900, N7876);
and AND4 (N7901, N7890, N5933, N4908, N4690);
and AND2 (N7902, N7901, N6926);
and AND2 (N7903, N7880, N2291);
xor XOR2 (N7904, N7885, N7619);
and AND4 (N7905, N7903, N2723, N5664, N6005);
xor XOR2 (N7906, N7899, N5152);
xor XOR2 (N7907, N7869, N1175);
nor NOR3 (N7908, N7905, N7564, N6422);
or OR4 (N7909, N7908, N6012, N660, N1128);
buf BUF1 (N7910, N7898);
nor NOR3 (N7911, N7896, N182, N1521);
not NOT1 (N7912, N7911);
buf BUF1 (N7913, N7891);
nand NAND3 (N7914, N7906, N6972, N3303);
not NOT1 (N7915, N7900);
nor NOR4 (N7916, N7912, N6317, N6670, N3062);
xor XOR2 (N7917, N7902, N4411);
nor NOR2 (N7918, N7914, N127);
buf BUF1 (N7919, N7909);
and AND4 (N7920, N7913, N437, N558, N4763);
nand NAND3 (N7921, N7920, N170, N6342);
or OR4 (N7922, N7921, N110, N7869, N4254);
nand NAND2 (N7923, N7917, N6189);
not NOT1 (N7924, N7904);
nor NOR4 (N7925, N7907, N1508, N1685, N4970);
xor XOR2 (N7926, N7892, N7799);
not NOT1 (N7927, N7926);
and AND2 (N7928, N7925, N4177);
and AND4 (N7929, N7928, N7445, N3539, N3019);
xor XOR2 (N7930, N7929, N2849);
nor NOR4 (N7931, N7918, N520, N4645, N7597);
nand NAND4 (N7932, N7930, N6762, N7346, N2876);
nand NAND3 (N7933, N7915, N2897, N6203);
not NOT1 (N7934, N7932);
nor NOR3 (N7935, N7934, N556, N7649);
and AND2 (N7936, N7923, N3799);
not NOT1 (N7937, N7935);
nor NOR4 (N7938, N7919, N5321, N3192, N1080);
nor NOR4 (N7939, N7931, N2947, N1654, N1257);
buf BUF1 (N7940, N7927);
xor XOR2 (N7941, N7939, N1865);
nor NOR3 (N7942, N7916, N552, N7604);
or OR3 (N7943, N7938, N7149, N2659);
or OR2 (N7944, N7942, N4202);
or OR4 (N7945, N7933, N2082, N3954, N4938);
xor XOR2 (N7946, N7922, N3395);
not NOT1 (N7947, N7944);
not NOT1 (N7948, N7946);
nor NOR4 (N7949, N7948, N5027, N5143, N3599);
and AND3 (N7950, N7910, N1579, N1960);
xor XOR2 (N7951, N7945, N6731);
nor NOR4 (N7952, N7936, N6416, N2454, N181);
nor NOR2 (N7953, N7947, N3979);
buf BUF1 (N7954, N7952);
xor XOR2 (N7955, N7951, N635);
nand NAND2 (N7956, N7954, N2300);
not NOT1 (N7957, N7949);
and AND2 (N7958, N7940, N7000);
buf BUF1 (N7959, N7950);
nor NOR4 (N7960, N7957, N4337, N7398, N6803);
not NOT1 (N7961, N7955);
not NOT1 (N7962, N7960);
and AND3 (N7963, N7956, N4516, N7425);
nor NOR3 (N7964, N7953, N2397, N4260);
nand NAND3 (N7965, N7958, N2417, N4428);
not NOT1 (N7966, N7959);
and AND2 (N7967, N7966, N7422);
nor NOR2 (N7968, N7962, N6994);
buf BUF1 (N7969, N7968);
xor XOR2 (N7970, N7965, N651);
buf BUF1 (N7971, N7943);
nand NAND3 (N7972, N7963, N1272, N2318);
or OR4 (N7973, N7969, N1489, N4118, N94);
buf BUF1 (N7974, N7973);
nor NOR4 (N7975, N7967, N6734, N1272, N6054);
xor XOR2 (N7976, N7972, N4963);
not NOT1 (N7977, N7961);
nand NAND3 (N7978, N7975, N2417, N2037);
xor XOR2 (N7979, N7976, N719);
not NOT1 (N7980, N7974);
nand NAND2 (N7981, N7980, N5820);
xor XOR2 (N7982, N7964, N6879);
not NOT1 (N7983, N7978);
nor NOR3 (N7984, N7924, N1534, N3703);
not NOT1 (N7985, N7937);
not NOT1 (N7986, N7982);
or OR2 (N7987, N7977, N1632);
and AND3 (N7988, N7984, N6316, N874);
nand NAND3 (N7989, N7986, N5959, N1908);
nor NOR2 (N7990, N7971, N4780);
or OR3 (N7991, N7979, N7963, N2738);
not NOT1 (N7992, N7989);
not NOT1 (N7993, N7987);
nand NAND4 (N7994, N7991, N1031, N2086, N7877);
xor XOR2 (N7995, N7985, N6382);
and AND4 (N7996, N7994, N916, N6674, N2097);
or OR3 (N7997, N7941, N712, N7806);
buf BUF1 (N7998, N7990);
not NOT1 (N7999, N7997);
xor XOR2 (N8000, N7999, N5973);
xor XOR2 (N8001, N7981, N225);
or OR2 (N8002, N7970, N2943);
and AND4 (N8003, N7992, N4825, N2187, N806);
nor NOR4 (N8004, N7983, N5224, N3038, N1);
or OR2 (N8005, N8000, N4279);
xor XOR2 (N8006, N7988, N6169);
nor NOR4 (N8007, N8005, N3981, N7, N3917);
not NOT1 (N8008, N7998);
buf BUF1 (N8009, N8002);
buf BUF1 (N8010, N8001);
xor XOR2 (N8011, N8006, N1816);
buf BUF1 (N8012, N8009);
or OR4 (N8013, N8004, N2653, N5002, N2675);
nor NOR2 (N8014, N8003, N4406);
nor NOR2 (N8015, N7993, N5844);
nand NAND3 (N8016, N8011, N4224, N1611);
nor NOR3 (N8017, N8007, N7988, N6517);
buf BUF1 (N8018, N8010);
and AND4 (N8019, N7996, N1773, N703, N519);
buf BUF1 (N8020, N8015);
not NOT1 (N8021, N8013);
not NOT1 (N8022, N7995);
and AND3 (N8023, N8017, N54, N5976);
nor NOR3 (N8024, N8016, N4908, N1046);
nand NAND4 (N8025, N8019, N6228, N701, N4284);
not NOT1 (N8026, N8020);
xor XOR2 (N8027, N8018, N5844);
xor XOR2 (N8028, N8026, N3129);
or OR4 (N8029, N8022, N4272, N2418, N6024);
or OR2 (N8030, N8029, N7763);
or OR4 (N8031, N8024, N4098, N5567, N7883);
buf BUF1 (N8032, N8008);
and AND3 (N8033, N8030, N759, N1107);
not NOT1 (N8034, N8033);
not NOT1 (N8035, N8031);
nand NAND3 (N8036, N8032, N5613, N4259);
xor XOR2 (N8037, N8023, N2557);
buf BUF1 (N8038, N8035);
buf BUF1 (N8039, N8037);
and AND3 (N8040, N8025, N4481, N2836);
or OR3 (N8041, N8027, N4619, N2616);
nand NAND4 (N8042, N8041, N7537, N3880, N539);
nand NAND4 (N8043, N8040, N4480, N3660, N2106);
nor NOR2 (N8044, N8014, N5591);
and AND2 (N8045, N8012, N1572);
nand NAND2 (N8046, N8039, N1669);
not NOT1 (N8047, N8028);
not NOT1 (N8048, N8047);
nand NAND3 (N8049, N8043, N418, N3773);
nand NAND2 (N8050, N8044, N1213);
nand NAND2 (N8051, N8038, N6930);
nand NAND2 (N8052, N8042, N1921);
buf BUF1 (N8053, N8036);
not NOT1 (N8054, N8045);
or OR2 (N8055, N8050, N361);
nand NAND3 (N8056, N8034, N1307, N4803);
xor XOR2 (N8057, N8052, N1193);
and AND3 (N8058, N8056, N4807, N3240);
or OR3 (N8059, N8057, N2884, N8057);
xor XOR2 (N8060, N8053, N7941);
and AND4 (N8061, N8060, N3374, N7072, N5926);
or OR2 (N8062, N8059, N4412);
or OR2 (N8063, N8049, N2256);
nor NOR4 (N8064, N8046, N6272, N129, N7800);
and AND2 (N8065, N8062, N1905);
nand NAND2 (N8066, N8021, N2743);
and AND2 (N8067, N8061, N3250);
or OR3 (N8068, N8063, N4709, N1324);
xor XOR2 (N8069, N8055, N6388);
or OR4 (N8070, N8066, N6261, N3557, N787);
buf BUF1 (N8071, N8054);
buf BUF1 (N8072, N8065);
and AND2 (N8073, N8068, N3205);
nand NAND4 (N8074, N8070, N1839, N7987, N623);
not NOT1 (N8075, N8073);
buf BUF1 (N8076, N8058);
nor NOR4 (N8077, N8067, N1884, N7673, N5640);
xor XOR2 (N8078, N8071, N915);
and AND2 (N8079, N8069, N1963);
not NOT1 (N8080, N8051);
buf BUF1 (N8081, N8072);
nor NOR2 (N8082, N8074, N5160);
nor NOR2 (N8083, N8082, N3418);
and AND2 (N8084, N8064, N2128);
nand NAND2 (N8085, N8083, N1731);
xor XOR2 (N8086, N8076, N7738);
or OR4 (N8087, N8085, N4772, N7097, N7645);
not NOT1 (N8088, N8084);
buf BUF1 (N8089, N8086);
buf BUF1 (N8090, N8078);
not NOT1 (N8091, N8081);
or OR3 (N8092, N8090, N5952, N1467);
buf BUF1 (N8093, N8048);
nor NOR3 (N8094, N8075, N171, N2504);
and AND2 (N8095, N8087, N5369);
and AND3 (N8096, N8079, N3418, N2286);
xor XOR2 (N8097, N8094, N5662);
nand NAND3 (N8098, N8093, N215, N7480);
or OR3 (N8099, N8098, N1250, N6369);
or OR2 (N8100, N8080, N2953);
buf BUF1 (N8101, N8091);
or OR2 (N8102, N8100, N4596);
nand NAND2 (N8103, N8077, N2426);
nor NOR2 (N8104, N8102, N4506);
xor XOR2 (N8105, N8089, N29);
or OR2 (N8106, N8092, N3061);
nand NAND4 (N8107, N8106, N2579, N7146, N5861);
and AND4 (N8108, N8095, N2207, N3803, N7331);
xor XOR2 (N8109, N8104, N6523);
and AND2 (N8110, N8108, N4107);
not NOT1 (N8111, N8107);
not NOT1 (N8112, N8105);
or OR3 (N8113, N8101, N6390, N6323);
or OR4 (N8114, N8112, N7846, N2148, N2506);
xor XOR2 (N8115, N8097, N136);
or OR2 (N8116, N8110, N5355);
nor NOR2 (N8117, N8116, N119);
or OR4 (N8118, N8113, N3993, N3396, N2950);
and AND2 (N8119, N8111, N5785);
buf BUF1 (N8120, N8118);
nand NAND3 (N8121, N8109, N8061, N4814);
nor NOR3 (N8122, N8114, N4857, N6523);
and AND3 (N8123, N8088, N5784, N6863);
not NOT1 (N8124, N8123);
or OR2 (N8125, N8121, N2270);
buf BUF1 (N8126, N8099);
nor NOR4 (N8127, N8096, N1960, N3191, N4017);
buf BUF1 (N8128, N8124);
nand NAND4 (N8129, N8115, N5480, N4747, N7013);
nand NAND3 (N8130, N8128, N2041, N7537);
and AND2 (N8131, N8120, N2151);
xor XOR2 (N8132, N8131, N7696);
buf BUF1 (N8133, N8126);
or OR4 (N8134, N8130, N1146, N4348, N3307);
nor NOR4 (N8135, N8129, N4551, N5892, N4617);
and AND4 (N8136, N8103, N1278, N8118, N2490);
buf BUF1 (N8137, N8119);
and AND3 (N8138, N8117, N1908, N6409);
or OR2 (N8139, N8138, N1215);
buf BUF1 (N8140, N8133);
xor XOR2 (N8141, N8134, N1785);
xor XOR2 (N8142, N8139, N6637);
and AND2 (N8143, N8125, N7144);
nor NOR3 (N8144, N8135, N923, N6804);
nand NAND2 (N8145, N8132, N3264);
nand NAND3 (N8146, N8144, N7071, N1959);
and AND2 (N8147, N8141, N5676);
nand NAND3 (N8148, N8140, N6072, N607);
or OR3 (N8149, N8142, N1710, N3197);
xor XOR2 (N8150, N8127, N3716);
or OR3 (N8151, N8149, N1326, N438);
nand NAND3 (N8152, N8143, N8022, N4351);
xor XOR2 (N8153, N8151, N4551);
and AND4 (N8154, N8136, N8062, N4146, N5799);
buf BUF1 (N8155, N8153);
and AND3 (N8156, N8146, N2328, N2116);
buf BUF1 (N8157, N8148);
nand NAND3 (N8158, N8147, N5627, N4489);
nor NOR3 (N8159, N8137, N1058, N1551);
not NOT1 (N8160, N8157);
and AND2 (N8161, N8145, N2523);
not NOT1 (N8162, N8155);
nor NOR2 (N8163, N8162, N4005);
nor NOR4 (N8164, N8122, N5864, N1210, N405);
and AND3 (N8165, N8163, N4604, N1532);
nor NOR4 (N8166, N8161, N6956, N1456, N1773);
or OR2 (N8167, N8156, N3732);
buf BUF1 (N8168, N8154);
xor XOR2 (N8169, N8165, N7086);
or OR4 (N8170, N8169, N5436, N4473, N5084);
not NOT1 (N8171, N8152);
nor NOR3 (N8172, N8170, N1103, N7218);
xor XOR2 (N8173, N8172, N6294);
or OR4 (N8174, N8164, N6398, N5921, N7490);
buf BUF1 (N8175, N8166);
or OR3 (N8176, N8171, N7824, N6699);
nor NOR4 (N8177, N8167, N4665, N1733, N3108);
not NOT1 (N8178, N8174);
xor XOR2 (N8179, N8177, N1541);
and AND4 (N8180, N8178, N599, N1621, N3144);
or OR3 (N8181, N8180, N4369, N6469);
xor XOR2 (N8182, N8150, N4275);
and AND3 (N8183, N8158, N7292, N7341);
nor NOR4 (N8184, N8181, N6357, N1432, N5804);
or OR4 (N8185, N8182, N2441, N4253, N6732);
xor XOR2 (N8186, N8168, N3624);
nor NOR3 (N8187, N8183, N1838, N6019);
xor XOR2 (N8188, N8179, N1295);
nand NAND4 (N8189, N8188, N2176, N1015, N6700);
buf BUF1 (N8190, N8187);
buf BUF1 (N8191, N8189);
buf BUF1 (N8192, N8191);
nand NAND3 (N8193, N8159, N7772, N712);
buf BUF1 (N8194, N8184);
and AND2 (N8195, N8193, N983);
xor XOR2 (N8196, N8192, N7184);
nand NAND4 (N8197, N8173, N887, N5840, N3942);
buf BUF1 (N8198, N8195);
buf BUF1 (N8199, N8185);
xor XOR2 (N8200, N8199, N4673);
nor NOR2 (N8201, N8196, N5183);
buf BUF1 (N8202, N8194);
nor NOR2 (N8203, N8202, N6232);
nand NAND2 (N8204, N8175, N531);
and AND4 (N8205, N8160, N4592, N3320, N5332);
not NOT1 (N8206, N8186);
nor NOR3 (N8207, N8204, N6830, N3911);
xor XOR2 (N8208, N8200, N7559);
xor XOR2 (N8209, N8197, N1351);
or OR4 (N8210, N8198, N8122, N6109, N7730);
or OR3 (N8211, N8190, N2707, N5924);
buf BUF1 (N8212, N8211);
nand NAND2 (N8213, N8201, N7910);
xor XOR2 (N8214, N8206, N4135);
nand NAND2 (N8215, N8176, N3147);
or OR2 (N8216, N8207, N469);
xor XOR2 (N8217, N8208, N7778);
not NOT1 (N8218, N8203);
xor XOR2 (N8219, N8218, N5158);
nand NAND4 (N8220, N8205, N2004, N5677, N2298);
and AND2 (N8221, N8217, N5040);
and AND2 (N8222, N8210, N6915);
nand NAND3 (N8223, N8213, N717, N5590);
and AND3 (N8224, N8212, N2544, N7569);
buf BUF1 (N8225, N8223);
xor XOR2 (N8226, N8215, N7287);
nand NAND3 (N8227, N8226, N383, N6983);
or OR2 (N8228, N8214, N7027);
xor XOR2 (N8229, N8221, N7857);
not NOT1 (N8230, N8225);
xor XOR2 (N8231, N8224, N5100);
or OR3 (N8232, N8219, N7484, N7514);
buf BUF1 (N8233, N8220);
nor NOR3 (N8234, N8231, N2630, N783);
nand NAND2 (N8235, N8230, N2865);
xor XOR2 (N8236, N8228, N4773);
not NOT1 (N8237, N8229);
nor NOR3 (N8238, N8236, N4281, N1960);
nor NOR4 (N8239, N8235, N7654, N2684, N5052);
or OR4 (N8240, N8233, N5698, N5906, N382);
nor NOR2 (N8241, N8239, N1140);
and AND2 (N8242, N8232, N5387);
nand NAND4 (N8243, N8234, N1031, N845, N7909);
and AND2 (N8244, N8243, N6426);
nand NAND3 (N8245, N8240, N5372, N317);
and AND2 (N8246, N8237, N7881);
xor XOR2 (N8247, N8241, N3971);
or OR4 (N8248, N8216, N4462, N5514, N7904);
nor NOR2 (N8249, N8238, N3317);
and AND4 (N8250, N8244, N6486, N4530, N1777);
or OR3 (N8251, N8248, N5248, N899);
nand NAND2 (N8252, N8246, N3906);
xor XOR2 (N8253, N8242, N1895);
nor NOR4 (N8254, N8245, N3990, N819, N7212);
not NOT1 (N8255, N8227);
and AND2 (N8256, N8254, N248);
nand NAND3 (N8257, N8256, N4422, N3114);
or OR3 (N8258, N8250, N3507, N3653);
or OR4 (N8259, N8222, N7055, N7926, N1466);
buf BUF1 (N8260, N8258);
buf BUF1 (N8261, N8255);
and AND3 (N8262, N8247, N2966, N466);
nor NOR2 (N8263, N8257, N7322);
nand NAND4 (N8264, N8260, N2195, N6727, N4372);
xor XOR2 (N8265, N8263, N7494);
or OR4 (N8266, N8252, N4425, N1719, N760);
and AND3 (N8267, N8261, N3036, N176);
nand NAND2 (N8268, N8253, N3216);
or OR2 (N8269, N8251, N6503);
or OR2 (N8270, N8264, N2889);
or OR2 (N8271, N8265, N2416);
buf BUF1 (N8272, N8209);
nand NAND4 (N8273, N8269, N2149, N3925, N880);
buf BUF1 (N8274, N8262);
not NOT1 (N8275, N8259);
buf BUF1 (N8276, N8266);
nor NOR4 (N8277, N8268, N7774, N378, N431);
not NOT1 (N8278, N8277);
nor NOR3 (N8279, N8272, N7287, N4895);
buf BUF1 (N8280, N8275);
not NOT1 (N8281, N8276);
not NOT1 (N8282, N8270);
xor XOR2 (N8283, N8281, N4738);
not NOT1 (N8284, N8271);
and AND4 (N8285, N8274, N1809, N3837, N1107);
buf BUF1 (N8286, N8279);
xor XOR2 (N8287, N8285, N4136);
and AND2 (N8288, N8267, N3879);
buf BUF1 (N8289, N8282);
nand NAND3 (N8290, N8280, N6598, N5383);
buf BUF1 (N8291, N8283);
nor NOR2 (N8292, N8286, N2244);
and AND2 (N8293, N8289, N1561);
xor XOR2 (N8294, N8291, N6231);
nand NAND2 (N8295, N8278, N6682);
nor NOR4 (N8296, N8293, N3971, N5525, N3002);
buf BUF1 (N8297, N8249);
nor NOR4 (N8298, N8295, N6537, N6986, N2223);
not NOT1 (N8299, N8287);
xor XOR2 (N8300, N8297, N4203);
buf BUF1 (N8301, N8298);
buf BUF1 (N8302, N8290);
or OR3 (N8303, N8301, N3731, N4204);
nor NOR2 (N8304, N8288, N3241);
buf BUF1 (N8305, N8304);
and AND4 (N8306, N8300, N5809, N259, N3335);
buf BUF1 (N8307, N8305);
nor NOR3 (N8308, N8296, N5310, N6726);
nor NOR3 (N8309, N8292, N738, N8209);
and AND4 (N8310, N8308, N5975, N496, N5498);
nand NAND3 (N8311, N8307, N139, N1338);
nand NAND2 (N8312, N8309, N7061);
not NOT1 (N8313, N8311);
nor NOR4 (N8314, N8303, N3117, N992, N4893);
and AND3 (N8315, N8284, N2198, N3300);
buf BUF1 (N8316, N8313);
nand NAND2 (N8317, N8314, N433);
buf BUF1 (N8318, N8310);
nor NOR2 (N8319, N8299, N3353);
not NOT1 (N8320, N8312);
or OR4 (N8321, N8302, N7962, N1540, N2515);
nor NOR3 (N8322, N8320, N2090, N6314);
not NOT1 (N8323, N8294);
and AND2 (N8324, N8315, N4835);
or OR2 (N8325, N8319, N4295);
xor XOR2 (N8326, N8317, N5923);
and AND3 (N8327, N8321, N4945, N4303);
nand NAND3 (N8328, N8325, N2048, N6452);
xor XOR2 (N8329, N8323, N335);
xor XOR2 (N8330, N8273, N20);
xor XOR2 (N8331, N8322, N3942);
buf BUF1 (N8332, N8324);
xor XOR2 (N8333, N8329, N3813);
nor NOR3 (N8334, N8331, N4789, N957);
nand NAND3 (N8335, N8306, N420, N3838);
or OR4 (N8336, N8327, N1914, N6370, N6054);
buf BUF1 (N8337, N8330);
or OR3 (N8338, N8337, N1160, N4110);
and AND3 (N8339, N8316, N4142, N5673);
buf BUF1 (N8340, N8332);
not NOT1 (N8341, N8338);
nor NOR2 (N8342, N8318, N7004);
or OR2 (N8343, N8335, N714);
buf BUF1 (N8344, N8342);
buf BUF1 (N8345, N8336);
and AND4 (N8346, N8340, N7952, N7106, N4902);
nand NAND4 (N8347, N8339, N1735, N5308, N680);
or OR4 (N8348, N8328, N604, N3892, N7619);
buf BUF1 (N8349, N8344);
buf BUF1 (N8350, N8341);
and AND2 (N8351, N8343, N8258);
nand NAND4 (N8352, N8345, N2444, N1365, N5228);
nand NAND2 (N8353, N8351, N1026);
or OR3 (N8354, N8352, N1777, N2865);
nor NOR2 (N8355, N8353, N5377);
xor XOR2 (N8356, N8349, N4490);
nand NAND2 (N8357, N8334, N2013);
nand NAND4 (N8358, N8347, N1684, N3414, N4725);
or OR4 (N8359, N8346, N5432, N1368, N6569);
not NOT1 (N8360, N8350);
buf BUF1 (N8361, N8333);
nor NOR2 (N8362, N8348, N7037);
nand NAND3 (N8363, N8361, N2085, N978);
nor NOR2 (N8364, N8363, N5108);
not NOT1 (N8365, N8354);
or OR3 (N8366, N8355, N725, N4361);
nand NAND4 (N8367, N8365, N7953, N1159, N1740);
or OR4 (N8368, N8360, N5984, N1682, N3654);
nand NAND3 (N8369, N8368, N1998, N3491);
xor XOR2 (N8370, N8362, N5426);
nor NOR4 (N8371, N8367, N8128, N441, N6606);
nand NAND3 (N8372, N8358, N2658, N7615);
xor XOR2 (N8373, N8356, N7659);
or OR2 (N8374, N8371, N1191);
or OR2 (N8375, N8369, N5710);
or OR4 (N8376, N8366, N6529, N253, N5427);
nand NAND4 (N8377, N8374, N5112, N5571, N6436);
xor XOR2 (N8378, N8373, N5404);
nor NOR3 (N8379, N8357, N6141, N1331);
nand NAND3 (N8380, N8370, N889, N5664);
nor NOR3 (N8381, N8359, N6273, N1885);
or OR4 (N8382, N8375, N7608, N2897, N78);
not NOT1 (N8383, N8382);
xor XOR2 (N8384, N8326, N7162);
nand NAND2 (N8385, N8384, N7826);
buf BUF1 (N8386, N8372);
nand NAND3 (N8387, N8383, N1143, N1998);
not NOT1 (N8388, N8364);
nand NAND4 (N8389, N8387, N8021, N6757, N691);
or OR2 (N8390, N8389, N5962);
and AND4 (N8391, N8390, N4286, N7528, N1676);
or OR4 (N8392, N8388, N5859, N4876, N1093);
nand NAND3 (N8393, N8392, N1783, N684);
not NOT1 (N8394, N8379);
nand NAND4 (N8395, N8381, N6405, N7936, N4305);
or OR2 (N8396, N8391, N2593);
nor NOR4 (N8397, N8385, N3779, N3091, N6261);
xor XOR2 (N8398, N8393, N4522);
and AND4 (N8399, N8376, N2689, N6296, N1664);
buf BUF1 (N8400, N8398);
and AND2 (N8401, N8378, N5891);
buf BUF1 (N8402, N8396);
buf BUF1 (N8403, N8377);
xor XOR2 (N8404, N8402, N4724);
and AND3 (N8405, N8399, N3187, N2338);
xor XOR2 (N8406, N8405, N3812);
or OR3 (N8407, N8397, N1532, N7856);
nand NAND3 (N8408, N8403, N1165, N5707);
or OR2 (N8409, N8401, N6342);
not NOT1 (N8410, N8400);
buf BUF1 (N8411, N8380);
xor XOR2 (N8412, N8395, N2433);
xor XOR2 (N8413, N8386, N4966);
buf BUF1 (N8414, N8409);
buf BUF1 (N8415, N8412);
and AND2 (N8416, N8404, N6246);
nor NOR4 (N8417, N8394, N334, N2300, N2930);
nor NOR4 (N8418, N8413, N1926, N10, N5044);
nand NAND2 (N8419, N8410, N5101);
nor NOR4 (N8420, N8419, N720, N1896, N5238);
xor XOR2 (N8421, N8417, N6);
and AND4 (N8422, N8420, N3017, N5876, N4621);
nand NAND4 (N8423, N8415, N821, N1529, N5110);
xor XOR2 (N8424, N8411, N6019);
xor XOR2 (N8425, N8406, N5423);
nor NOR2 (N8426, N8423, N6137);
buf BUF1 (N8427, N8408);
or OR4 (N8428, N8427, N1955, N4448, N3920);
or OR2 (N8429, N8428, N7723);
and AND3 (N8430, N8421, N6945, N7496);
or OR3 (N8431, N8424, N6152, N1574);
xor XOR2 (N8432, N8407, N3204);
nand NAND4 (N8433, N8416, N187, N2913, N2276);
xor XOR2 (N8434, N8426, N4388);
nand NAND3 (N8435, N8434, N2707, N5626);
and AND4 (N8436, N8433, N7186, N1286, N1962);
buf BUF1 (N8437, N8431);
nor NOR3 (N8438, N8429, N6164, N7664);
not NOT1 (N8439, N8418);
nor NOR2 (N8440, N8438, N2179);
nor NOR4 (N8441, N8436, N4202, N2905, N1245);
or OR4 (N8442, N8422, N5313, N5779, N3030);
not NOT1 (N8443, N8414);
nor NOR2 (N8444, N8443, N3994);
nor NOR2 (N8445, N8432, N2318);
nor NOR2 (N8446, N8439, N726);
buf BUF1 (N8447, N8441);
buf BUF1 (N8448, N8445);
nor NOR4 (N8449, N8444, N5646, N5719, N5344);
nand NAND4 (N8450, N8437, N3969, N8271, N1593);
and AND2 (N8451, N8448, N477);
or OR4 (N8452, N8440, N4124, N4912, N762);
nor NOR3 (N8453, N8430, N1820, N4506);
nand NAND3 (N8454, N8453, N7414, N998);
nor NOR4 (N8455, N8446, N7231, N3668, N1620);
or OR2 (N8456, N8450, N258);
and AND3 (N8457, N8425, N6902, N153);
nand NAND3 (N8458, N8455, N2950, N30);
or OR4 (N8459, N8449, N7330, N7479, N8160);
or OR3 (N8460, N8442, N3285, N6337);
not NOT1 (N8461, N8459);
not NOT1 (N8462, N8460);
buf BUF1 (N8463, N8457);
not NOT1 (N8464, N8452);
nand NAND3 (N8465, N8454, N274, N2698);
buf BUF1 (N8466, N8451);
and AND3 (N8467, N8464, N1805, N3430);
nand NAND4 (N8468, N8467, N2244, N2813, N5853);
nand NAND3 (N8469, N8435, N2781, N6998);
and AND4 (N8470, N8461, N7889, N4702, N2899);
or OR3 (N8471, N8470, N6112, N2342);
not NOT1 (N8472, N8468);
buf BUF1 (N8473, N8471);
buf BUF1 (N8474, N8473);
and AND3 (N8475, N8466, N1723, N6696);
and AND3 (N8476, N8472, N5877, N6732);
nand NAND3 (N8477, N8474, N3386, N7859);
buf BUF1 (N8478, N8475);
nand NAND3 (N8479, N8447, N8209, N4707);
xor XOR2 (N8480, N8478, N427);
or OR2 (N8481, N8479, N424);
and AND2 (N8482, N8458, N6690);
nand NAND2 (N8483, N8477, N7965);
nand NAND2 (N8484, N8465, N6348);
buf BUF1 (N8485, N8482);
not NOT1 (N8486, N8485);
xor XOR2 (N8487, N8456, N7618);
nand NAND4 (N8488, N8462, N5606, N3768, N7252);
nor NOR2 (N8489, N8487, N6168);
xor XOR2 (N8490, N8476, N2694);
buf BUF1 (N8491, N8488);
xor XOR2 (N8492, N8469, N2094);
not NOT1 (N8493, N8486);
not NOT1 (N8494, N8493);
and AND3 (N8495, N8494, N3131, N2186);
nor NOR2 (N8496, N8489, N6946);
nand NAND2 (N8497, N8480, N6787);
nand NAND2 (N8498, N8490, N3874);
and AND2 (N8499, N8497, N6298);
xor XOR2 (N8500, N8483, N7974);
or OR3 (N8501, N8484, N4895, N2055);
not NOT1 (N8502, N8500);
and AND2 (N8503, N8481, N1443);
not NOT1 (N8504, N8503);
or OR2 (N8505, N8502, N7374);
or OR2 (N8506, N8498, N7172);
nand NAND2 (N8507, N8491, N1795);
not NOT1 (N8508, N8499);
xor XOR2 (N8509, N8504, N2086);
not NOT1 (N8510, N8495);
not NOT1 (N8511, N8463);
buf BUF1 (N8512, N8506);
not NOT1 (N8513, N8512);
nand NAND3 (N8514, N8511, N4468, N6955);
or OR4 (N8515, N8513, N7171, N5384, N911);
not NOT1 (N8516, N8508);
and AND3 (N8517, N8515, N3731, N8071);
or OR3 (N8518, N8514, N6548, N6328);
nor NOR2 (N8519, N8496, N5230);
not NOT1 (N8520, N8517);
not NOT1 (N8521, N8510);
nand NAND2 (N8522, N8507, N2215);
nor NOR3 (N8523, N8492, N1637, N5761);
buf BUF1 (N8524, N8501);
nand NAND2 (N8525, N8523, N2910);
or OR4 (N8526, N8519, N1128, N6276, N8412);
nand NAND4 (N8527, N8520, N4074, N7923, N1101);
buf BUF1 (N8528, N8518);
nand NAND4 (N8529, N8516, N5413, N7115, N1479);
nor NOR3 (N8530, N8525, N1882, N5534);
nand NAND4 (N8531, N8509, N7681, N1855, N4416);
nand NAND3 (N8532, N8530, N8412, N273);
nor NOR2 (N8533, N8528, N3517);
not NOT1 (N8534, N8521);
nor NOR4 (N8535, N8531, N449, N3277, N3796);
or OR2 (N8536, N8527, N2616);
and AND3 (N8537, N8505, N2462, N5879);
buf BUF1 (N8538, N8522);
buf BUF1 (N8539, N8529);
nor NOR4 (N8540, N8535, N8284, N3772, N675);
not NOT1 (N8541, N8532);
nor NOR3 (N8542, N8536, N4442, N7981);
nor NOR3 (N8543, N8524, N5759, N4016);
buf BUF1 (N8544, N8543);
buf BUF1 (N8545, N8538);
xor XOR2 (N8546, N8541, N2410);
nor NOR3 (N8547, N8542, N8336, N3073);
and AND4 (N8548, N8526, N2761, N3875, N1478);
xor XOR2 (N8549, N8534, N6638);
xor XOR2 (N8550, N8547, N4089);
xor XOR2 (N8551, N8537, N1691);
xor XOR2 (N8552, N8546, N3627);
or OR4 (N8553, N8539, N6470, N1896, N2117);
buf BUF1 (N8554, N8533);
not NOT1 (N8555, N8554);
nor NOR3 (N8556, N8544, N4144, N8436);
xor XOR2 (N8557, N8552, N4335);
or OR4 (N8558, N8550, N4978, N1480, N5565);
xor XOR2 (N8559, N8555, N2055);
xor XOR2 (N8560, N8559, N4624);
and AND3 (N8561, N8553, N1178, N1332);
not NOT1 (N8562, N8545);
nor NOR3 (N8563, N8556, N2381, N4694);
or OR2 (N8564, N8560, N186);
buf BUF1 (N8565, N8561);
or OR3 (N8566, N8558, N4877, N1147);
not NOT1 (N8567, N8566);
nand NAND4 (N8568, N8562, N811, N2645, N2214);
and AND4 (N8569, N8540, N7445, N6729, N8140);
nand NAND2 (N8570, N8568, N6369);
buf BUF1 (N8571, N8557);
xor XOR2 (N8572, N8551, N1399);
buf BUF1 (N8573, N8565);
not NOT1 (N8574, N8563);
not NOT1 (N8575, N8569);
buf BUF1 (N8576, N8548);
nand NAND2 (N8577, N8572, N903);
not NOT1 (N8578, N8567);
and AND4 (N8579, N8578, N5948, N3265, N3708);
buf BUF1 (N8580, N8576);
or OR2 (N8581, N8570, N1483);
buf BUF1 (N8582, N8577);
xor XOR2 (N8583, N8549, N2862);
buf BUF1 (N8584, N8583);
nor NOR2 (N8585, N8564, N6570);
xor XOR2 (N8586, N8580, N3358);
xor XOR2 (N8587, N8575, N195);
or OR3 (N8588, N8587, N6014, N5742);
nor NOR2 (N8589, N8585, N2498);
and AND3 (N8590, N8581, N3342, N3238);
and AND3 (N8591, N8586, N4881, N3570);
and AND4 (N8592, N8589, N5273, N4344, N7896);
buf BUF1 (N8593, N8574);
xor XOR2 (N8594, N8579, N8543);
nor NOR2 (N8595, N8588, N402);
nand NAND4 (N8596, N8592, N6842, N2964, N4678);
nand NAND4 (N8597, N8594, N3927, N8300, N2552);
not NOT1 (N8598, N8593);
and AND2 (N8599, N8584, N6235);
nor NOR4 (N8600, N8582, N3774, N2165, N3780);
xor XOR2 (N8601, N8591, N1431);
or OR3 (N8602, N8590, N7377, N4872);
not NOT1 (N8603, N8599);
nand NAND3 (N8604, N8603, N3116, N7751);
buf BUF1 (N8605, N8601);
and AND4 (N8606, N8598, N5008, N5853, N7020);
xor XOR2 (N8607, N8602, N1844);
nor NOR3 (N8608, N8606, N1404, N3655);
nand NAND4 (N8609, N8600, N3140, N1701, N2383);
or OR3 (N8610, N8573, N7477, N6861);
and AND3 (N8611, N8609, N8277, N4180);
and AND3 (N8612, N8610, N4624, N1582);
nor NOR4 (N8613, N8604, N7760, N1749, N2329);
nor NOR4 (N8614, N8571, N828, N7805, N5787);
not NOT1 (N8615, N8597);
nand NAND3 (N8616, N8607, N5930, N1346);
and AND4 (N8617, N8616, N6729, N3373, N4519);
and AND4 (N8618, N8608, N1068, N4462, N3192);
not NOT1 (N8619, N8613);
not NOT1 (N8620, N8618);
xor XOR2 (N8621, N8619, N1816);
nand NAND4 (N8622, N8617, N4784, N2836, N7139);
buf BUF1 (N8623, N8605);
not NOT1 (N8624, N8620);
buf BUF1 (N8625, N8623);
buf BUF1 (N8626, N8614);
and AND2 (N8627, N8625, N5368);
xor XOR2 (N8628, N8621, N680);
nor NOR2 (N8629, N8627, N151);
buf BUF1 (N8630, N8629);
nand NAND2 (N8631, N8612, N3570);
buf BUF1 (N8632, N8622);
not NOT1 (N8633, N8628);
or OR4 (N8634, N8632, N6068, N3276, N2350);
nor NOR4 (N8635, N8630, N8286, N4408, N5100);
nor NOR2 (N8636, N8633, N2511);
and AND2 (N8637, N8636, N6885);
or OR2 (N8638, N8634, N935);
xor XOR2 (N8639, N8626, N4761);
not NOT1 (N8640, N8631);
xor XOR2 (N8641, N8595, N6881);
xor XOR2 (N8642, N8596, N2338);
or OR3 (N8643, N8641, N4187, N2467);
and AND4 (N8644, N8639, N1822, N5254, N8233);
nor NOR4 (N8645, N8615, N1628, N4183, N2684);
buf BUF1 (N8646, N8638);
xor XOR2 (N8647, N8624, N5870);
buf BUF1 (N8648, N8647);
xor XOR2 (N8649, N8611, N864);
not NOT1 (N8650, N8646);
nor NOR4 (N8651, N8637, N7968, N3821, N7982);
or OR4 (N8652, N8644, N5327, N518, N805);
nor NOR3 (N8653, N8649, N1145, N6496);
not NOT1 (N8654, N8650);
nand NAND2 (N8655, N8651, N446);
xor XOR2 (N8656, N8635, N2362);
buf BUF1 (N8657, N8642);
buf BUF1 (N8658, N8656);
nand NAND2 (N8659, N8645, N7272);
buf BUF1 (N8660, N8640);
and AND3 (N8661, N8648, N66, N2882);
xor XOR2 (N8662, N8659, N332);
xor XOR2 (N8663, N8654, N555);
and AND3 (N8664, N8662, N1007, N6404);
and AND2 (N8665, N8663, N2466);
nand NAND4 (N8666, N8665, N2694, N2505, N6830);
and AND4 (N8667, N8652, N1509, N8520, N8485);
xor XOR2 (N8668, N8661, N4711);
nor NOR2 (N8669, N8668, N8100);
or OR2 (N8670, N8669, N2231);
nor NOR3 (N8671, N8667, N423, N4187);
or OR3 (N8672, N8653, N2806, N8558);
nand NAND2 (N8673, N8670, N5859);
not NOT1 (N8674, N8643);
nor NOR4 (N8675, N8658, N3143, N8603, N6090);
buf BUF1 (N8676, N8660);
not NOT1 (N8677, N8674);
buf BUF1 (N8678, N8655);
and AND3 (N8679, N8673, N2079, N375);
nor NOR4 (N8680, N8679, N6059, N2979, N7665);
nand NAND4 (N8681, N8664, N6181, N5326, N699);
nand NAND3 (N8682, N8666, N4472, N2004);
nand NAND2 (N8683, N8675, N6738);
or OR2 (N8684, N8672, N5755);
nor NOR4 (N8685, N8682, N345, N2766, N4932);
xor XOR2 (N8686, N8680, N6132);
and AND3 (N8687, N8657, N6292, N2937);
xor XOR2 (N8688, N8687, N5251);
nand NAND4 (N8689, N8678, N6572, N7962, N5222);
and AND4 (N8690, N8684, N6463, N113, N6769);
nand NAND4 (N8691, N8676, N1443, N4237, N7171);
xor XOR2 (N8692, N8688, N8180);
and AND2 (N8693, N8692, N754);
buf BUF1 (N8694, N8677);
and AND3 (N8695, N8691, N4381, N6913);
nor NOR4 (N8696, N8690, N390, N5729, N93);
and AND2 (N8697, N8695, N3203);
and AND4 (N8698, N8686, N5153, N7063, N3822);
nand NAND4 (N8699, N8693, N4680, N3686, N1840);
xor XOR2 (N8700, N8698, N5626);
and AND4 (N8701, N8696, N1344, N2543, N3381);
not NOT1 (N8702, N8699);
xor XOR2 (N8703, N8694, N4573);
or OR3 (N8704, N8697, N6400, N851);
not NOT1 (N8705, N8702);
or OR3 (N8706, N8704, N490, N6954);
nor NOR4 (N8707, N8701, N8360, N6582, N5108);
xor XOR2 (N8708, N8683, N2324);
nand NAND3 (N8709, N8703, N3055, N671);
or OR2 (N8710, N8671, N5691);
nand NAND4 (N8711, N8708, N4032, N4090, N116);
nand NAND2 (N8712, N8709, N7222);
nor NOR2 (N8713, N8681, N1000);
and AND4 (N8714, N8706, N8358, N1270, N6251);
buf BUF1 (N8715, N8714);
nand NAND3 (N8716, N8689, N6535, N1530);
nand NAND3 (N8717, N8710, N2183, N7692);
nor NOR3 (N8718, N8707, N6797, N4880);
nand NAND2 (N8719, N8718, N410);
and AND4 (N8720, N8715, N277, N8305, N6331);
or OR4 (N8721, N8713, N7144, N4437, N3972);
xor XOR2 (N8722, N8717, N8005);
buf BUF1 (N8723, N8685);
and AND3 (N8724, N8712, N2842, N8331);
or OR3 (N8725, N8719, N2284, N1022);
not NOT1 (N8726, N8725);
nand NAND2 (N8727, N8724, N3492);
not NOT1 (N8728, N8721);
and AND4 (N8729, N8711, N7805, N103, N8225);
xor XOR2 (N8730, N8729, N3422);
buf BUF1 (N8731, N8723);
nand NAND4 (N8732, N8716, N8576, N1054, N4198);
not NOT1 (N8733, N8731);
nand NAND3 (N8734, N8728, N8013, N7986);
xor XOR2 (N8735, N8727, N7726);
or OR4 (N8736, N8730, N2634, N3821, N7920);
or OR4 (N8737, N8732, N1392, N783, N7838);
nand NAND2 (N8738, N8733, N5964);
or OR4 (N8739, N8737, N1814, N7161, N4606);
or OR3 (N8740, N8720, N5480, N3322);
not NOT1 (N8741, N8735);
nand NAND2 (N8742, N8738, N5493);
xor XOR2 (N8743, N8705, N2780);
not NOT1 (N8744, N8740);
nand NAND4 (N8745, N8741, N6585, N3767, N8435);
or OR4 (N8746, N8734, N1268, N7163, N1645);
buf BUF1 (N8747, N8745);
buf BUF1 (N8748, N8736);
buf BUF1 (N8749, N8748);
and AND4 (N8750, N8749, N829, N3646, N3094);
nand NAND3 (N8751, N8742, N7842, N3462);
xor XOR2 (N8752, N8751, N3770);
not NOT1 (N8753, N8739);
buf BUF1 (N8754, N8722);
and AND2 (N8755, N8750, N3906);
buf BUF1 (N8756, N8746);
xor XOR2 (N8757, N8754, N3840);
nand NAND4 (N8758, N8744, N7310, N4712, N3583);
nor NOR2 (N8759, N8726, N1332);
or OR4 (N8760, N8747, N7856, N5017, N7368);
nand NAND4 (N8761, N8752, N6779, N330, N6075);
and AND4 (N8762, N8759, N5048, N6695, N2882);
not NOT1 (N8763, N8762);
buf BUF1 (N8764, N8753);
and AND4 (N8765, N8757, N37, N3553, N3766);
or OR3 (N8766, N8764, N4850, N355);
nand NAND4 (N8767, N8756, N2477, N1671, N1823);
xor XOR2 (N8768, N8763, N4291);
or OR4 (N8769, N8743, N8195, N6074, N4609);
nor NOR3 (N8770, N8767, N110, N5775);
nor NOR3 (N8771, N8761, N8667, N3298);
buf BUF1 (N8772, N8771);
xor XOR2 (N8773, N8755, N1878);
nand NAND3 (N8774, N8768, N3050, N6728);
buf BUF1 (N8775, N8769);
not NOT1 (N8776, N8773);
or OR2 (N8777, N8700, N5441);
xor XOR2 (N8778, N8776, N8706);
nand NAND2 (N8779, N8775, N3965);
buf BUF1 (N8780, N8778);
nand NAND2 (N8781, N8765, N4289);
and AND2 (N8782, N8780, N6325);
xor XOR2 (N8783, N8770, N8104);
nor NOR2 (N8784, N8781, N1664);
nand NAND2 (N8785, N8779, N3660);
buf BUF1 (N8786, N8782);
and AND3 (N8787, N8784, N3227, N5772);
buf BUF1 (N8788, N8777);
nand NAND2 (N8789, N8786, N966);
xor XOR2 (N8790, N8788, N5039);
nand NAND4 (N8791, N8772, N208, N5331, N8441);
not NOT1 (N8792, N8758);
not NOT1 (N8793, N8766);
nand NAND4 (N8794, N8787, N515, N3565, N8752);
and AND3 (N8795, N8783, N7628, N971);
not NOT1 (N8796, N8792);
not NOT1 (N8797, N8790);
not NOT1 (N8798, N8796);
nand NAND3 (N8799, N8774, N7238, N6287);
buf BUF1 (N8800, N8789);
buf BUF1 (N8801, N8798);
xor XOR2 (N8802, N8800, N5137);
buf BUF1 (N8803, N8793);
nand NAND3 (N8804, N8795, N7017, N7027);
and AND2 (N8805, N8760, N6563);
nand NAND2 (N8806, N8804, N2454);
xor XOR2 (N8807, N8806, N716);
or OR2 (N8808, N8805, N7302);
or OR2 (N8809, N8801, N568);
buf BUF1 (N8810, N8808);
nor NOR4 (N8811, N8799, N8372, N6901, N3628);
nand NAND3 (N8812, N8810, N2428, N1484);
xor XOR2 (N8813, N8791, N7165);
nand NAND3 (N8814, N8785, N1662, N5750);
buf BUF1 (N8815, N8794);
or OR4 (N8816, N8802, N8275, N7954, N6476);
nand NAND3 (N8817, N8811, N8751, N3979);
or OR3 (N8818, N8813, N1799, N2800);
not NOT1 (N8819, N8797);
buf BUF1 (N8820, N8812);
not NOT1 (N8821, N8807);
nor NOR4 (N8822, N8819, N115, N386, N5807);
and AND3 (N8823, N8809, N1865, N2768);
buf BUF1 (N8824, N8803);
and AND4 (N8825, N8816, N2123, N8452, N4754);
or OR2 (N8826, N8822, N651);
or OR3 (N8827, N8818, N7856, N1430);
not NOT1 (N8828, N8825);
nor NOR4 (N8829, N8826, N6380, N2761, N1701);
buf BUF1 (N8830, N8817);
or OR2 (N8831, N8830, N5793);
buf BUF1 (N8832, N8815);
nand NAND2 (N8833, N8820, N5808);
buf BUF1 (N8834, N8832);
nand NAND4 (N8835, N8828, N3058, N6825, N8098);
and AND3 (N8836, N8823, N4303, N2289);
nor NOR3 (N8837, N8836, N1392, N8033);
or OR2 (N8838, N8829, N8000);
not NOT1 (N8839, N8821);
not NOT1 (N8840, N8831);
not NOT1 (N8841, N8814);
xor XOR2 (N8842, N8837, N3548);
buf BUF1 (N8843, N8838);
and AND2 (N8844, N8840, N43);
xor XOR2 (N8845, N8835, N6058);
not NOT1 (N8846, N8843);
xor XOR2 (N8847, N8834, N8135);
and AND3 (N8848, N8845, N5347, N6438);
or OR2 (N8849, N8847, N1142);
not NOT1 (N8850, N8839);
buf BUF1 (N8851, N8844);
nand NAND2 (N8852, N8833, N8161);
not NOT1 (N8853, N8848);
buf BUF1 (N8854, N8852);
buf BUF1 (N8855, N8824);
and AND2 (N8856, N8853, N1444);
nand NAND3 (N8857, N8856, N4781, N186);
xor XOR2 (N8858, N8849, N5867);
and AND3 (N8859, N8851, N1780, N2857);
xor XOR2 (N8860, N8858, N5158);
xor XOR2 (N8861, N8850, N4618);
buf BUF1 (N8862, N8827);
xor XOR2 (N8863, N8860, N8431);
or OR4 (N8864, N8861, N8362, N1182, N7284);
buf BUF1 (N8865, N8863);
or OR4 (N8866, N8855, N3959, N6830, N2902);
buf BUF1 (N8867, N8842);
and AND3 (N8868, N8866, N7125, N8663);
or OR2 (N8869, N8854, N5485);
nand NAND2 (N8870, N8868, N54);
nand NAND3 (N8871, N8862, N2136, N3772);
buf BUF1 (N8872, N8841);
buf BUF1 (N8873, N8865);
or OR4 (N8874, N8859, N384, N2890, N3558);
nor NOR3 (N8875, N8846, N2143, N5199);
nor NOR4 (N8876, N8869, N2218, N4638, N1646);
not NOT1 (N8877, N8872);
and AND2 (N8878, N8876, N412);
nor NOR3 (N8879, N8870, N8133, N8631);
and AND2 (N8880, N8867, N4157);
and AND3 (N8881, N8857, N5337, N1894);
and AND3 (N8882, N8875, N6522, N5417);
buf BUF1 (N8883, N8878);
nand NAND4 (N8884, N8883, N5832, N4546, N4482);
nand NAND4 (N8885, N8882, N1889, N2295, N2391);
xor XOR2 (N8886, N8879, N8228);
nand NAND2 (N8887, N8881, N2544);
buf BUF1 (N8888, N8884);
nand NAND4 (N8889, N8886, N5224, N5850, N3214);
buf BUF1 (N8890, N8885);
xor XOR2 (N8891, N8890, N2387);
and AND2 (N8892, N8873, N8031);
and AND4 (N8893, N8891, N5964, N5961, N7530);
nor NOR3 (N8894, N8888, N1019, N3864);
and AND3 (N8895, N8892, N1952, N6240);
xor XOR2 (N8896, N8887, N3296);
nand NAND4 (N8897, N8864, N2442, N8847, N8565);
nand NAND3 (N8898, N8877, N2199, N7798);
nor NOR4 (N8899, N8898, N1259, N554, N1735);
not NOT1 (N8900, N8893);
or OR3 (N8901, N8894, N3180, N6315);
xor XOR2 (N8902, N8880, N7647);
or OR4 (N8903, N8871, N1743, N7564, N1346);
nor NOR4 (N8904, N8901, N7400, N4027, N1197);
not NOT1 (N8905, N8902);
buf BUF1 (N8906, N8896);
nand NAND2 (N8907, N8905, N3525);
nor NOR2 (N8908, N8889, N7639);
and AND4 (N8909, N8895, N6673, N6259, N8532);
and AND2 (N8910, N8897, N6467);
nor NOR4 (N8911, N8907, N7681, N7481, N3197);
nor NOR4 (N8912, N8911, N5990, N977, N5089);
not NOT1 (N8913, N8909);
xor XOR2 (N8914, N8906, N8403);
buf BUF1 (N8915, N8903);
and AND2 (N8916, N8904, N4090);
nor NOR2 (N8917, N8874, N6302);
xor XOR2 (N8918, N8912, N1236);
or OR2 (N8919, N8910, N4741);
not NOT1 (N8920, N8913);
and AND3 (N8921, N8917, N6938, N7925);
xor XOR2 (N8922, N8915, N3416);
and AND2 (N8923, N8919, N4819);
buf BUF1 (N8924, N8918);
xor XOR2 (N8925, N8920, N3814);
nor NOR2 (N8926, N8924, N2729);
and AND3 (N8927, N8921, N8437, N8615);
nor NOR4 (N8928, N8926, N7790, N7031, N2228);
and AND2 (N8929, N8927, N8804);
xor XOR2 (N8930, N8899, N2670);
buf BUF1 (N8931, N8925);
not NOT1 (N8932, N8923);
not NOT1 (N8933, N8916);
not NOT1 (N8934, N8933);
and AND4 (N8935, N8930, N4448, N1552, N4768);
nand NAND2 (N8936, N8929, N1953);
xor XOR2 (N8937, N8922, N710);
buf BUF1 (N8938, N8928);
nor NOR3 (N8939, N8908, N3047, N8724);
or OR4 (N8940, N8932, N8380, N1805, N5627);
xor XOR2 (N8941, N8939, N7670);
or OR3 (N8942, N8938, N1174, N2723);
buf BUF1 (N8943, N8900);
nor NOR4 (N8944, N8935, N4824, N6842, N2431);
or OR2 (N8945, N8934, N8456);
nor NOR2 (N8946, N8937, N6642);
xor XOR2 (N8947, N8942, N1011);
not NOT1 (N8948, N8940);
not NOT1 (N8949, N8947);
or OR3 (N8950, N8914, N7155, N2886);
xor XOR2 (N8951, N8941, N7125);
or OR2 (N8952, N8945, N5110);
nand NAND2 (N8953, N8949, N4040);
or OR2 (N8954, N8951, N1201);
or OR3 (N8955, N8953, N4887, N5210);
not NOT1 (N8956, N8946);
buf BUF1 (N8957, N8954);
buf BUF1 (N8958, N8931);
or OR4 (N8959, N8957, N6962, N6196, N2372);
or OR4 (N8960, N8948, N7537, N7378, N7974);
nor NOR4 (N8961, N8952, N3421, N4593, N5980);
buf BUF1 (N8962, N8955);
and AND2 (N8963, N8962, N987);
buf BUF1 (N8964, N8960);
nor NOR2 (N8965, N8950, N1816);
buf BUF1 (N8966, N8965);
buf BUF1 (N8967, N8943);
nand NAND4 (N8968, N8964, N6370, N3953, N8794);
nor NOR2 (N8969, N8963, N2033);
nand NAND4 (N8970, N8944, N6474, N4000, N3885);
buf BUF1 (N8971, N8936);
or OR2 (N8972, N8966, N7353);
nand NAND3 (N8973, N8961, N5361, N391);
nor NOR2 (N8974, N8972, N4901);
not NOT1 (N8975, N8959);
buf BUF1 (N8976, N8973);
not NOT1 (N8977, N8970);
nand NAND2 (N8978, N8969, N4107);
or OR3 (N8979, N8971, N4300, N59);
nand NAND2 (N8980, N8968, N3510);
nand NAND4 (N8981, N8977, N685, N1279, N1969);
and AND3 (N8982, N8956, N3369, N5627);
not NOT1 (N8983, N8979);
and AND3 (N8984, N8974, N8563, N1248);
buf BUF1 (N8985, N8978);
nand NAND4 (N8986, N8980, N8441, N3306, N106);
xor XOR2 (N8987, N8982, N6197);
and AND3 (N8988, N8984, N8686, N4556);
and AND4 (N8989, N8967, N6301, N2042, N462);
or OR3 (N8990, N8981, N4695, N4606);
not NOT1 (N8991, N8989);
not NOT1 (N8992, N8975);
not NOT1 (N8993, N8987);
nor NOR2 (N8994, N8988, N3603);
buf BUF1 (N8995, N8976);
buf BUF1 (N8996, N8958);
not NOT1 (N8997, N8994);
not NOT1 (N8998, N8995);
or OR2 (N8999, N8992, N6414);
and AND2 (N9000, N8983, N6740);
nor NOR2 (N9001, N8986, N5433);
xor XOR2 (N9002, N8991, N8676);
xor XOR2 (N9003, N9001, N5440);
xor XOR2 (N9004, N8993, N593);
nor NOR3 (N9005, N9002, N924, N881);
nand NAND3 (N9006, N8997, N575, N3486);
buf BUF1 (N9007, N8996);
xor XOR2 (N9008, N9007, N3037);
nand NAND2 (N9009, N9004, N6510);
nor NOR3 (N9010, N9008, N4935, N3851);
and AND2 (N9011, N9003, N4114);
not NOT1 (N9012, N9005);
nor NOR3 (N9013, N9012, N6162, N2723);
not NOT1 (N9014, N8990);
buf BUF1 (N9015, N9009);
and AND4 (N9016, N9015, N6326, N1263, N3233);
or OR2 (N9017, N9000, N8017);
or OR2 (N9018, N9013, N2043);
nand NAND4 (N9019, N9018, N6172, N6861, N3465);
nand NAND2 (N9020, N8985, N6187);
xor XOR2 (N9021, N8998, N718);
nor NOR2 (N9022, N9010, N2342);
xor XOR2 (N9023, N9020, N7911);
not NOT1 (N9024, N9014);
nand NAND2 (N9025, N9024, N1832);
and AND3 (N9026, N9016, N1444, N5026);
buf BUF1 (N9027, N9006);
not NOT1 (N9028, N9017);
nand NAND2 (N9029, N9027, N1570);
xor XOR2 (N9030, N9026, N4952);
buf BUF1 (N9031, N9025);
nor NOR2 (N9032, N9028, N1604);
or OR3 (N9033, N9011, N7714, N1362);
nor NOR3 (N9034, N9033, N1112, N4713);
and AND3 (N9035, N9030, N4358, N6411);
not NOT1 (N9036, N9019);
buf BUF1 (N9037, N9034);
nor NOR2 (N9038, N9035, N518);
not NOT1 (N9039, N9036);
and AND4 (N9040, N9037, N2341, N4998, N4020);
or OR3 (N9041, N9039, N4719, N1131);
nor NOR3 (N9042, N9038, N5154, N3202);
buf BUF1 (N9043, N9041);
nand NAND3 (N9044, N9031, N7782, N3323);
xor XOR2 (N9045, N9029, N7534);
buf BUF1 (N9046, N9021);
and AND4 (N9047, N9040, N7031, N4372, N4507);
and AND2 (N9048, N9046, N8107);
not NOT1 (N9049, N9022);
or OR4 (N9050, N9023, N2695, N5333, N2666);
or OR2 (N9051, N9049, N7916);
nand NAND4 (N9052, N8999, N7594, N3216, N7059);
xor XOR2 (N9053, N9052, N1539);
not NOT1 (N9054, N9048);
not NOT1 (N9055, N9045);
nor NOR3 (N9056, N9043, N7629, N2775);
or OR2 (N9057, N9054, N22);
nand NAND3 (N9058, N9057, N8384, N124);
nand NAND2 (N9059, N9053, N810);
nor NOR3 (N9060, N9047, N5440, N3931);
buf BUF1 (N9061, N9058);
or OR2 (N9062, N9059, N6923);
and AND3 (N9063, N9044, N572, N3732);
nor NOR2 (N9064, N9063, N4383);
nand NAND4 (N9065, N9060, N805, N6772, N3412);
not NOT1 (N9066, N9056);
xor XOR2 (N9067, N9050, N1734);
nor NOR2 (N9068, N9061, N4313);
or OR4 (N9069, N9064, N7992, N3497, N673);
nand NAND2 (N9070, N9055, N5129);
nand NAND2 (N9071, N9062, N7290);
nor NOR4 (N9072, N9042, N5379, N9025, N5191);
nand NAND4 (N9073, N9069, N4163, N4721, N8393);
xor XOR2 (N9074, N9067, N6623);
buf BUF1 (N9075, N9065);
nor NOR3 (N9076, N9066, N8330, N2963);
buf BUF1 (N9077, N9032);
nand NAND2 (N9078, N9076, N959);
nor NOR4 (N9079, N9070, N8771, N582, N7163);
or OR3 (N9080, N9078, N5169, N6389);
and AND2 (N9081, N9074, N2353);
and AND2 (N9082, N9081, N8402);
or OR3 (N9083, N9051, N1251, N2699);
not NOT1 (N9084, N9073);
nand NAND4 (N9085, N9079, N792, N2895, N3573);
not NOT1 (N9086, N9083);
and AND2 (N9087, N9082, N3812);
and AND2 (N9088, N9068, N5052);
nor NOR2 (N9089, N9072, N8858);
nand NAND3 (N9090, N9080, N3568, N3551);
buf BUF1 (N9091, N9071);
and AND3 (N9092, N9084, N1184, N3906);
or OR4 (N9093, N9092, N4792, N8639, N1746);
and AND4 (N9094, N9093, N5294, N6693, N8610);
or OR4 (N9095, N9089, N4687, N4615, N7546);
buf BUF1 (N9096, N9075);
and AND3 (N9097, N9094, N1948, N8617);
buf BUF1 (N9098, N9087);
nor NOR2 (N9099, N9086, N5706);
or OR3 (N9100, N9091, N4950, N2655);
and AND2 (N9101, N9095, N5059);
nand NAND2 (N9102, N9101, N2943);
not NOT1 (N9103, N9098);
not NOT1 (N9104, N9103);
not NOT1 (N9105, N9104);
buf BUF1 (N9106, N9099);
buf BUF1 (N9107, N9102);
nand NAND3 (N9108, N9105, N2975, N3325);
xor XOR2 (N9109, N9088, N4982);
nand NAND4 (N9110, N9085, N2927, N3863, N5726);
not NOT1 (N9111, N9107);
nand NAND3 (N9112, N9110, N8553, N7805);
or OR3 (N9113, N9108, N3243, N1665);
nand NAND4 (N9114, N9113, N8543, N6243, N1487);
and AND2 (N9115, N9106, N3473);
not NOT1 (N9116, N9100);
and AND3 (N9117, N9090, N984, N4223);
or OR3 (N9118, N9117, N3694, N6070);
nor NOR2 (N9119, N9097, N5842);
xor XOR2 (N9120, N9096, N1012);
or OR4 (N9121, N9111, N7825, N762, N3449);
and AND3 (N9122, N9120, N238, N842);
or OR3 (N9123, N9115, N2443, N5289);
or OR2 (N9124, N9109, N6508);
buf BUF1 (N9125, N9122);
nor NOR2 (N9126, N9121, N3444);
buf BUF1 (N9127, N9112);
nand NAND2 (N9128, N9119, N7629);
and AND3 (N9129, N9127, N6094, N2306);
or OR3 (N9130, N9126, N3009, N5976);
and AND2 (N9131, N9125, N5574);
nor NOR3 (N9132, N9129, N3526, N6350);
not NOT1 (N9133, N9123);
and AND4 (N9134, N9130, N4715, N4426, N267);
and AND3 (N9135, N9124, N3138, N1458);
xor XOR2 (N9136, N9118, N2028);
not NOT1 (N9137, N9135);
buf BUF1 (N9138, N9132);
xor XOR2 (N9139, N9133, N5051);
and AND3 (N9140, N9131, N914, N8670);
or OR4 (N9141, N9114, N8742, N2748, N6735);
nor NOR2 (N9142, N9128, N6145);
nand NAND3 (N9143, N9137, N6783, N1335);
or OR4 (N9144, N9139, N4881, N3048, N3386);
nor NOR3 (N9145, N9136, N3707, N4718);
nand NAND3 (N9146, N9077, N4756, N5848);
nor NOR3 (N9147, N9141, N3429, N3099);
nand NAND3 (N9148, N9138, N56, N691);
xor XOR2 (N9149, N9142, N8050);
buf BUF1 (N9150, N9134);
nand NAND3 (N9151, N9144, N4370, N5644);
nor NOR3 (N9152, N9116, N7622, N5140);
nor NOR3 (N9153, N9150, N6292, N6260);
or OR3 (N9154, N9143, N8748, N4151);
not NOT1 (N9155, N9147);
and AND2 (N9156, N9151, N5894);
nor NOR3 (N9157, N9152, N4894, N2459);
nand NAND2 (N9158, N9156, N1097);
nand NAND2 (N9159, N9157, N6172);
nand NAND4 (N9160, N9149, N4492, N5927, N4554);
or OR2 (N9161, N9148, N7317);
xor XOR2 (N9162, N9161, N6068);
or OR4 (N9163, N9158, N1321, N4501, N8088);
not NOT1 (N9164, N9155);
nor NOR3 (N9165, N9145, N1531, N5034);
nor NOR4 (N9166, N9165, N2380, N208, N2481);
not NOT1 (N9167, N9162);
not NOT1 (N9168, N9166);
buf BUF1 (N9169, N9163);
and AND3 (N9170, N9153, N4555, N2198);
nor NOR4 (N9171, N9168, N6431, N4664, N252);
nor NOR4 (N9172, N9140, N1947, N5642, N2586);
and AND2 (N9173, N9159, N8908);
or OR2 (N9174, N9154, N8206);
and AND4 (N9175, N9164, N1446, N7735, N5082);
or OR2 (N9176, N9173, N5048);
or OR2 (N9177, N9146, N8110);
nand NAND2 (N9178, N9169, N6503);
buf BUF1 (N9179, N9177);
and AND3 (N9180, N9176, N726, N8643);
nor NOR2 (N9181, N9167, N8318);
nor NOR2 (N9182, N9175, N8863);
or OR4 (N9183, N9174, N6584, N4601, N2700);
or OR4 (N9184, N9181, N2156, N1997, N1176);
xor XOR2 (N9185, N9183, N99);
nor NOR4 (N9186, N9184, N2342, N8315, N4387);
or OR3 (N9187, N9182, N4655, N8034);
and AND3 (N9188, N9180, N4117, N4569);
nor NOR4 (N9189, N9188, N6977, N8390, N5395);
or OR4 (N9190, N9178, N4082, N4281, N889);
nor NOR2 (N9191, N9189, N1784);
not NOT1 (N9192, N9170);
nand NAND4 (N9193, N9187, N1064, N6260, N7314);
nand NAND4 (N9194, N9191, N54, N496, N3189);
buf BUF1 (N9195, N9186);
not NOT1 (N9196, N9171);
and AND3 (N9197, N9196, N4035, N4409);
not NOT1 (N9198, N9179);
nand NAND2 (N9199, N9194, N4880);
nor NOR4 (N9200, N9192, N5886, N8644, N3446);
nand NAND4 (N9201, N9172, N3012, N8855, N7041);
not NOT1 (N9202, N9200);
xor XOR2 (N9203, N9201, N7999);
nand NAND2 (N9204, N9160, N779);
buf BUF1 (N9205, N9204);
buf BUF1 (N9206, N9205);
not NOT1 (N9207, N9197);
nor NOR3 (N9208, N9207, N5017, N2322);
and AND4 (N9209, N9185, N8206, N5979, N1069);
buf BUF1 (N9210, N9203);
buf BUF1 (N9211, N9208);
or OR2 (N9212, N9210, N565);
buf BUF1 (N9213, N9195);
and AND3 (N9214, N9212, N3769, N2802);
nor NOR4 (N9215, N9190, N7311, N8220, N7301);
xor XOR2 (N9216, N9202, N6868);
buf BUF1 (N9217, N9198);
or OR4 (N9218, N9215, N4447, N6514, N92);
nand NAND3 (N9219, N9206, N3237, N6728);
xor XOR2 (N9220, N9219, N1116);
not NOT1 (N9221, N9193);
buf BUF1 (N9222, N9216);
xor XOR2 (N9223, N9218, N2841);
buf BUF1 (N9224, N9221);
or OR4 (N9225, N9209, N8314, N5349, N2805);
not NOT1 (N9226, N9213);
nand NAND4 (N9227, N9211, N2862, N5628, N7957);
nand NAND4 (N9228, N9222, N8890, N3724, N7548);
buf BUF1 (N9229, N9199);
buf BUF1 (N9230, N9224);
not NOT1 (N9231, N9214);
xor XOR2 (N9232, N9227, N8340);
and AND3 (N9233, N9229, N6157, N9226);
or OR2 (N9234, N3506, N6088);
xor XOR2 (N9235, N9233, N2285);
and AND2 (N9236, N9217, N2979);
buf BUF1 (N9237, N9232);
xor XOR2 (N9238, N9228, N5242);
or OR3 (N9239, N9235, N1325, N4768);
nand NAND4 (N9240, N9234, N6465, N7270, N4224);
or OR3 (N9241, N9236, N3515, N8616);
not NOT1 (N9242, N9225);
not NOT1 (N9243, N9239);
not NOT1 (N9244, N9237);
buf BUF1 (N9245, N9240);
and AND2 (N9246, N9220, N6066);
not NOT1 (N9247, N9230);
buf BUF1 (N9248, N9241);
not NOT1 (N9249, N9247);
not NOT1 (N9250, N9242);
buf BUF1 (N9251, N9249);
nor NOR4 (N9252, N9238, N2743, N5605, N276);
or OR2 (N9253, N9223, N4729);
buf BUF1 (N9254, N9248);
and AND2 (N9255, N9246, N9154);
or OR4 (N9256, N9254, N4664, N6584, N6632);
nand NAND2 (N9257, N9244, N7260);
xor XOR2 (N9258, N9250, N2262);
xor XOR2 (N9259, N9231, N1391);
buf BUF1 (N9260, N9258);
nor NOR2 (N9261, N9256, N5454);
nand NAND2 (N9262, N9260, N3782);
nor NOR3 (N9263, N9261, N4247, N3993);
buf BUF1 (N9264, N9252);
or OR4 (N9265, N9262, N8285, N9185, N45);
nor NOR2 (N9266, N9255, N7381);
or OR2 (N9267, N9263, N5670);
buf BUF1 (N9268, N9257);
not NOT1 (N9269, N9243);
buf BUF1 (N9270, N9259);
and AND3 (N9271, N9267, N2487, N4587);
nand NAND2 (N9272, N9264, N738);
buf BUF1 (N9273, N9253);
not NOT1 (N9274, N9270);
and AND4 (N9275, N9273, N2198, N3911, N8120);
xor XOR2 (N9276, N9275, N4672);
not NOT1 (N9277, N9274);
nor NOR4 (N9278, N9272, N7019, N4633, N323);
and AND2 (N9279, N9271, N7958);
xor XOR2 (N9280, N9245, N1156);
nand NAND2 (N9281, N9277, N1250);
buf BUF1 (N9282, N9279);
nor NOR2 (N9283, N9278, N472);
buf BUF1 (N9284, N9276);
not NOT1 (N9285, N9269);
or OR4 (N9286, N9280, N8496, N7224, N8290);
nor NOR4 (N9287, N9285, N5676, N7947, N8349);
or OR4 (N9288, N9266, N8088, N3029, N2187);
not NOT1 (N9289, N9288);
buf BUF1 (N9290, N9283);
nor NOR4 (N9291, N9286, N2208, N4276, N7756);
and AND2 (N9292, N9289, N6864);
xor XOR2 (N9293, N9287, N4564);
xor XOR2 (N9294, N9293, N1370);
or OR2 (N9295, N9290, N7226);
or OR3 (N9296, N9292, N9214, N2691);
or OR3 (N9297, N9251, N7866, N4701);
nand NAND4 (N9298, N9297, N8436, N2329, N9214);
xor XOR2 (N9299, N9281, N7233);
nor NOR2 (N9300, N9268, N66);
not NOT1 (N9301, N9296);
not NOT1 (N9302, N9291);
xor XOR2 (N9303, N9301, N1757);
nand NAND4 (N9304, N9282, N2690, N2285, N9232);
and AND4 (N9305, N9302, N6284, N6455, N6693);
buf BUF1 (N9306, N9298);
buf BUF1 (N9307, N9295);
buf BUF1 (N9308, N9305);
nand NAND3 (N9309, N9300, N4859, N7449);
or OR4 (N9310, N9307, N2350, N6112, N1924);
nor NOR2 (N9311, N9308, N1281);
not NOT1 (N9312, N9310);
nand NAND2 (N9313, N9299, N4611);
and AND3 (N9314, N9311, N7983, N4120);
or OR2 (N9315, N9265, N6431);
and AND4 (N9316, N9309, N9192, N4441, N3795);
nand NAND2 (N9317, N9294, N47);
or OR4 (N9318, N9315, N2081, N4376, N4069);
xor XOR2 (N9319, N9304, N5286);
xor XOR2 (N9320, N9313, N4792);
xor XOR2 (N9321, N9319, N2016);
xor XOR2 (N9322, N9320, N7191);
and AND3 (N9323, N9306, N3694, N3079);
xor XOR2 (N9324, N9303, N6717);
nor NOR4 (N9325, N9321, N4554, N6448, N2699);
nand NAND2 (N9326, N9316, N1157);
or OR3 (N9327, N9312, N3286, N3144);
or OR3 (N9328, N9314, N3151, N2539);
or OR2 (N9329, N9318, N6623);
not NOT1 (N9330, N9329);
nand NAND4 (N9331, N9325, N6184, N2731, N8198);
and AND4 (N9332, N9322, N5447, N9277, N2446);
xor XOR2 (N9333, N9284, N1762);
xor XOR2 (N9334, N9332, N7140);
and AND3 (N9335, N9326, N3385, N7714);
buf BUF1 (N9336, N9334);
and AND2 (N9337, N9333, N800);
or OR2 (N9338, N9327, N8057);
buf BUF1 (N9339, N9328);
or OR4 (N9340, N9336, N1438, N2677, N4410);
nor NOR4 (N9341, N9331, N7869, N6101, N333);
not NOT1 (N9342, N9335);
nor NOR3 (N9343, N9330, N8690, N2587);
nor NOR2 (N9344, N9343, N4123);
and AND4 (N9345, N9323, N6875, N7405, N3731);
nand NAND4 (N9346, N9340, N515, N7961, N78);
or OR4 (N9347, N9317, N4269, N1778, N1771);
or OR2 (N9348, N9339, N531);
nor NOR2 (N9349, N9342, N5217);
and AND3 (N9350, N9348, N1930, N1426);
and AND2 (N9351, N9341, N8858);
buf BUF1 (N9352, N9344);
or OR3 (N9353, N9349, N529, N7178);
xor XOR2 (N9354, N9352, N377);
and AND3 (N9355, N9351, N6564, N5167);
and AND2 (N9356, N9350, N4733);
nand NAND3 (N9357, N9324, N6214, N1177);
nand NAND3 (N9358, N9346, N8520, N6202);
nand NAND2 (N9359, N9354, N1702);
xor XOR2 (N9360, N9357, N4426);
xor XOR2 (N9361, N9355, N8929);
buf BUF1 (N9362, N9360);
nor NOR4 (N9363, N9362, N3281, N156, N716);
nor NOR2 (N9364, N9347, N4701);
and AND4 (N9365, N9363, N4162, N7263, N7077);
and AND2 (N9366, N9358, N8754);
nor NOR4 (N9367, N9345, N3735, N6137, N9336);
nand NAND3 (N9368, N9365, N2875, N345);
nor NOR3 (N9369, N9368, N7063, N313);
nor NOR2 (N9370, N9364, N2779);
nor NOR4 (N9371, N9370, N2759, N3439, N831);
buf BUF1 (N9372, N9366);
or OR4 (N9373, N9356, N8685, N7184, N165);
not NOT1 (N9374, N9337);
and AND2 (N9375, N9369, N7349);
buf BUF1 (N9376, N9353);
nor NOR2 (N9377, N9361, N2933);
xor XOR2 (N9378, N9374, N1882);
buf BUF1 (N9379, N9376);
nand NAND2 (N9380, N9377, N7129);
xor XOR2 (N9381, N9378, N5386);
and AND4 (N9382, N9367, N7479, N9292, N6473);
or OR4 (N9383, N9372, N3752, N9226, N4462);
nand NAND3 (N9384, N9359, N3355, N516);
xor XOR2 (N9385, N9384, N232);
buf BUF1 (N9386, N9338);
nor NOR2 (N9387, N9385, N1931);
buf BUF1 (N9388, N9382);
nor NOR3 (N9389, N9388, N8252, N2798);
buf BUF1 (N9390, N9373);
and AND3 (N9391, N9383, N5724, N4184);
buf BUF1 (N9392, N9375);
or OR3 (N9393, N9387, N4141, N643);
nor NOR2 (N9394, N9386, N1977);
not NOT1 (N9395, N9394);
buf BUF1 (N9396, N9392);
not NOT1 (N9397, N9389);
or OR4 (N9398, N9380, N5570, N4617, N629);
nor NOR3 (N9399, N9379, N3384, N543);
not NOT1 (N9400, N9390);
not NOT1 (N9401, N9398);
xor XOR2 (N9402, N9399, N3475);
buf BUF1 (N9403, N9397);
or OR4 (N9404, N9396, N2715, N6407, N6428);
buf BUF1 (N9405, N9395);
or OR4 (N9406, N9404, N1222, N6534, N4510);
not NOT1 (N9407, N9400);
and AND4 (N9408, N9405, N7961, N4284, N3423);
not NOT1 (N9409, N9381);
nor NOR3 (N9410, N9403, N5771, N2285);
xor XOR2 (N9411, N9408, N2206);
or OR3 (N9412, N9371, N8480, N9196);
xor XOR2 (N9413, N9409, N4528);
nor NOR2 (N9414, N9406, N4818);
xor XOR2 (N9415, N9391, N4818);
and AND4 (N9416, N9411, N9121, N9183, N3643);
nor NOR3 (N9417, N9415, N7730, N2708);
or OR2 (N9418, N9413, N4415);
xor XOR2 (N9419, N9414, N1796);
xor XOR2 (N9420, N9417, N5876);
nor NOR3 (N9421, N9418, N7456, N7569);
and AND3 (N9422, N9402, N5664, N7223);
not NOT1 (N9423, N9412);
or OR2 (N9424, N9422, N4607);
buf BUF1 (N9425, N9407);
xor XOR2 (N9426, N9420, N4279);
or OR3 (N9427, N9421, N4393, N4443);
or OR3 (N9428, N9423, N3440, N3376);
nor NOR2 (N9429, N9416, N5660);
buf BUF1 (N9430, N9427);
nand NAND3 (N9431, N9430, N3427, N4700);
not NOT1 (N9432, N9425);
nor NOR2 (N9433, N9429, N7332);
or OR3 (N9434, N9432, N1758, N1775);
nor NOR4 (N9435, N9433, N6217, N4403, N8410);
buf BUF1 (N9436, N9410);
or OR4 (N9437, N9393, N6569, N9228, N6438);
buf BUF1 (N9438, N9431);
xor XOR2 (N9439, N9424, N2727);
not NOT1 (N9440, N9434);
or OR3 (N9441, N9440, N7337, N8431);
nand NAND4 (N9442, N9419, N6104, N5264, N4261);
nand NAND3 (N9443, N9442, N882, N1051);
xor XOR2 (N9444, N9401, N4828);
not NOT1 (N9445, N9438);
not NOT1 (N9446, N9426);
nor NOR4 (N9447, N9441, N3317, N2619, N1745);
nand NAND4 (N9448, N9439, N8654, N5947, N1126);
not NOT1 (N9449, N9436);
nor NOR4 (N9450, N9444, N4538, N8099, N7260);
buf BUF1 (N9451, N9428);
buf BUF1 (N9452, N9450);
nor NOR2 (N9453, N9445, N3083);
and AND2 (N9454, N9437, N2486);
and AND2 (N9455, N9447, N7956);
xor XOR2 (N9456, N9451, N8840);
xor XOR2 (N9457, N9435, N8548);
or OR3 (N9458, N9456, N9452, N6708);
or OR4 (N9459, N2936, N804, N2397, N6317);
and AND4 (N9460, N9455, N1851, N666, N2341);
xor XOR2 (N9461, N9458, N3020);
xor XOR2 (N9462, N9454, N7944);
and AND3 (N9463, N9460, N7857, N5179);
and AND3 (N9464, N9463, N5070, N60);
buf BUF1 (N9465, N9462);
buf BUF1 (N9466, N9448);
buf BUF1 (N9467, N9461);
not NOT1 (N9468, N9464);
or OR3 (N9469, N9466, N3571, N7346);
nand NAND4 (N9470, N9465, N7748, N193, N5609);
nor NOR4 (N9471, N9453, N4717, N1516, N8887);
and AND3 (N9472, N9470, N8851, N3681);
xor XOR2 (N9473, N9443, N8142);
xor XOR2 (N9474, N9457, N9209);
or OR3 (N9475, N9473, N4799, N5565);
and AND2 (N9476, N9474, N5247);
xor XOR2 (N9477, N9446, N6707);
nand NAND4 (N9478, N9468, N7206, N2131, N5633);
buf BUF1 (N9479, N9472);
and AND4 (N9480, N9467, N1292, N7915, N8218);
nand NAND2 (N9481, N9477, N2778);
and AND4 (N9482, N9476, N9431, N4872, N8848);
nor NOR2 (N9483, N9478, N7167);
and AND2 (N9484, N9481, N1013);
buf BUF1 (N9485, N9484);
or OR4 (N9486, N9459, N7150, N6851, N5108);
xor XOR2 (N9487, N9471, N3101);
xor XOR2 (N9488, N9482, N6710);
nor NOR2 (N9489, N9449, N6185);
nor NOR4 (N9490, N9469, N7131, N7751, N1499);
not NOT1 (N9491, N9490);
nand NAND3 (N9492, N9488, N116, N5420);
or OR4 (N9493, N9492, N185, N1907, N695);
nor NOR3 (N9494, N9491, N5554, N6262);
buf BUF1 (N9495, N9483);
or OR2 (N9496, N9487, N1072);
xor XOR2 (N9497, N9495, N2789);
buf BUF1 (N9498, N9496);
nor NOR4 (N9499, N9493, N2939, N1770, N3533);
and AND4 (N9500, N9485, N5364, N4970, N18);
buf BUF1 (N9501, N9494);
nand NAND2 (N9502, N9498, N5193);
nand NAND4 (N9503, N9500, N7153, N8494, N3227);
nor NOR2 (N9504, N9503, N2410);
buf BUF1 (N9505, N9499);
or OR4 (N9506, N9480, N1834, N1669, N2841);
not NOT1 (N9507, N9475);
not NOT1 (N9508, N9506);
nand NAND3 (N9509, N9489, N1607, N4980);
nand NAND2 (N9510, N9508, N1499);
or OR2 (N9511, N9510, N8088);
xor XOR2 (N9512, N9511, N433);
or OR4 (N9513, N9507, N6553, N3798, N5803);
not NOT1 (N9514, N9486);
not NOT1 (N9515, N9509);
buf BUF1 (N9516, N9505);
and AND2 (N9517, N9479, N4650);
nand NAND2 (N9518, N9501, N7117);
buf BUF1 (N9519, N9504);
not NOT1 (N9520, N9502);
xor XOR2 (N9521, N9519, N5763);
or OR2 (N9522, N9512, N3360);
nand NAND2 (N9523, N9497, N1609);
not NOT1 (N9524, N9515);
buf BUF1 (N9525, N9524);
nor NOR2 (N9526, N9521, N8780);
nor NOR4 (N9527, N9522, N8812, N9291, N444);
or OR2 (N9528, N9517, N995);
or OR2 (N9529, N9525, N5733);
nor NOR4 (N9530, N9526, N3973, N3949, N7706);
buf BUF1 (N9531, N9527);
nor NOR4 (N9532, N9520, N8494, N286, N5326);
not NOT1 (N9533, N9529);
and AND3 (N9534, N9528, N9110, N3815);
buf BUF1 (N9535, N9514);
not NOT1 (N9536, N9531);
nor NOR2 (N9537, N9532, N2194);
nand NAND2 (N9538, N9518, N8740);
and AND2 (N9539, N9538, N9154);
xor XOR2 (N9540, N9536, N2533);
nor NOR4 (N9541, N9533, N9285, N8236, N2004);
and AND3 (N9542, N9537, N9259, N7050);
or OR4 (N9543, N9540, N6062, N3270, N3550);
or OR2 (N9544, N9523, N87);
buf BUF1 (N9545, N9534);
nand NAND3 (N9546, N9530, N3300, N8075);
and AND3 (N9547, N9542, N7040, N1535);
or OR2 (N9548, N9516, N2296);
nand NAND2 (N9549, N9541, N9252);
or OR4 (N9550, N9513, N4387, N9289, N1315);
and AND2 (N9551, N9549, N3871);
nor NOR2 (N9552, N9539, N1895);
nand NAND3 (N9553, N9544, N7798, N9139);
or OR2 (N9554, N9546, N6872);
or OR4 (N9555, N9550, N1549, N7557, N7351);
xor XOR2 (N9556, N9552, N188);
buf BUF1 (N9557, N9556);
buf BUF1 (N9558, N9547);
not NOT1 (N9559, N9551);
xor XOR2 (N9560, N9555, N2575);
xor XOR2 (N9561, N9548, N4540);
nand NAND4 (N9562, N9545, N9354, N7611, N9370);
buf BUF1 (N9563, N9562);
nand NAND2 (N9564, N9554, N5934);
not NOT1 (N9565, N9543);
buf BUF1 (N9566, N9535);
buf BUF1 (N9567, N9558);
xor XOR2 (N9568, N9564, N2053);
xor XOR2 (N9569, N9561, N2117);
nor NOR3 (N9570, N9553, N9335, N4383);
nor NOR2 (N9571, N9568, N2523);
buf BUF1 (N9572, N9569);
and AND3 (N9573, N9565, N4566, N6647);
xor XOR2 (N9574, N9560, N9463);
and AND3 (N9575, N9557, N7050, N5307);
not NOT1 (N9576, N9570);
not NOT1 (N9577, N9573);
and AND3 (N9578, N9571, N4617, N8171);
buf BUF1 (N9579, N9559);
and AND3 (N9580, N9572, N4645, N6326);
xor XOR2 (N9581, N9578, N4965);
nor NOR4 (N9582, N9576, N8127, N210, N8996);
and AND3 (N9583, N9575, N5250, N4418);
xor XOR2 (N9584, N9583, N6103);
or OR3 (N9585, N9567, N6240, N4256);
xor XOR2 (N9586, N9577, N6656);
and AND4 (N9587, N9581, N988, N6972, N7610);
nand NAND4 (N9588, N9580, N2850, N5138, N1685);
or OR3 (N9589, N9588, N5811, N5888);
not NOT1 (N9590, N9579);
xor XOR2 (N9591, N9566, N5025);
xor XOR2 (N9592, N9585, N2588);
or OR3 (N9593, N9590, N8307, N2057);
buf BUF1 (N9594, N9591);
not NOT1 (N9595, N9587);
not NOT1 (N9596, N9586);
nand NAND2 (N9597, N9592, N5926);
xor XOR2 (N9598, N9582, N8896);
xor XOR2 (N9599, N9594, N330);
or OR4 (N9600, N9593, N4440, N9389, N5129);
or OR2 (N9601, N9599, N5445);
buf BUF1 (N9602, N9601);
xor XOR2 (N9603, N9589, N1681);
buf BUF1 (N9604, N9596);
xor XOR2 (N9605, N9604, N4167);
not NOT1 (N9606, N9602);
nand NAND2 (N9607, N9595, N2457);
buf BUF1 (N9608, N9563);
xor XOR2 (N9609, N9605, N7621);
buf BUF1 (N9610, N9609);
not NOT1 (N9611, N9610);
and AND4 (N9612, N9607, N7666, N6040, N8993);
nand NAND4 (N9613, N9612, N8684, N627, N3742);
not NOT1 (N9614, N9574);
and AND2 (N9615, N9597, N8428);
nor NOR4 (N9616, N9603, N2538, N2428, N3767);
not NOT1 (N9617, N9616);
or OR2 (N9618, N9614, N6949);
or OR4 (N9619, N9617, N2260, N6699, N4863);
nand NAND2 (N9620, N9600, N3687);
nand NAND2 (N9621, N9615, N1876);
or OR3 (N9622, N9598, N3507, N6745);
or OR3 (N9623, N9622, N4204, N5746);
or OR4 (N9624, N9623, N8951, N767, N4888);
xor XOR2 (N9625, N9606, N6359);
and AND3 (N9626, N9624, N4722, N321);
nand NAND4 (N9627, N9625, N7500, N583, N6052);
buf BUF1 (N9628, N9627);
buf BUF1 (N9629, N9626);
buf BUF1 (N9630, N9628);
or OR2 (N9631, N9629, N4832);
or OR3 (N9632, N9611, N1819, N1877);
not NOT1 (N9633, N9618);
or OR4 (N9634, N9620, N6524, N3959, N3172);
buf BUF1 (N9635, N9634);
not NOT1 (N9636, N9621);
buf BUF1 (N9637, N9631);
not NOT1 (N9638, N9637);
nand NAND3 (N9639, N9584, N4896, N6008);
xor XOR2 (N9640, N9635, N2435);
and AND3 (N9641, N9636, N4267, N864);
and AND3 (N9642, N9641, N9041, N7229);
xor XOR2 (N9643, N9608, N8772);
not NOT1 (N9644, N9619);
or OR4 (N9645, N9613, N8356, N261, N3994);
xor XOR2 (N9646, N9638, N1894);
or OR2 (N9647, N9642, N31);
or OR2 (N9648, N9647, N751);
xor XOR2 (N9649, N9645, N8974);
nand NAND3 (N9650, N9632, N6938, N3088);
not NOT1 (N9651, N9646);
xor XOR2 (N9652, N9648, N3250);
or OR2 (N9653, N9644, N4714);
nor NOR3 (N9654, N9651, N5030, N2697);
buf BUF1 (N9655, N9652);
or OR4 (N9656, N9640, N7018, N7176, N4951);
not NOT1 (N9657, N9643);
and AND4 (N9658, N9649, N2181, N3180, N9502);
not NOT1 (N9659, N9655);
buf BUF1 (N9660, N9659);
or OR4 (N9661, N9630, N8704, N3049, N5446);
buf BUF1 (N9662, N9654);
not NOT1 (N9663, N9658);
nand NAND2 (N9664, N9653, N5673);
or OR2 (N9665, N9656, N4140);
nor NOR3 (N9666, N9663, N1934, N4152);
nor NOR4 (N9667, N9666, N5674, N2856, N6770);
not NOT1 (N9668, N9664);
xor XOR2 (N9669, N9660, N1732);
buf BUF1 (N9670, N9650);
not NOT1 (N9671, N9633);
nand NAND2 (N9672, N9665, N6527);
nand NAND4 (N9673, N9657, N5525, N6054, N8287);
not NOT1 (N9674, N9667);
or OR3 (N9675, N9673, N4977, N5483);
nand NAND2 (N9676, N9670, N8670);
and AND2 (N9677, N9639, N6589);
and AND4 (N9678, N9677, N4924, N2738, N1334);
and AND3 (N9679, N9661, N8772, N9288);
xor XOR2 (N9680, N9671, N9234);
and AND3 (N9681, N9675, N614, N2790);
not NOT1 (N9682, N9680);
not NOT1 (N9683, N9669);
nand NAND3 (N9684, N9678, N5758, N1181);
nor NOR2 (N9685, N9679, N1705);
nand NAND2 (N9686, N9683, N1884);
not NOT1 (N9687, N9674);
or OR2 (N9688, N9676, N9270);
or OR2 (N9689, N9686, N5842);
not NOT1 (N9690, N9668);
not NOT1 (N9691, N9688);
buf BUF1 (N9692, N9687);
or OR2 (N9693, N9684, N3060);
xor XOR2 (N9694, N9672, N199);
and AND4 (N9695, N9691, N4109, N7346, N6762);
not NOT1 (N9696, N9694);
buf BUF1 (N9697, N9681);
not NOT1 (N9698, N9690);
and AND2 (N9699, N9662, N1111);
and AND4 (N9700, N9699, N6345, N8062, N6760);
and AND3 (N9701, N9692, N2544, N1114);
xor XOR2 (N9702, N9685, N6795);
not NOT1 (N9703, N9702);
buf BUF1 (N9704, N9682);
or OR2 (N9705, N9700, N725);
xor XOR2 (N9706, N9693, N4607);
xor XOR2 (N9707, N9697, N5047);
buf BUF1 (N9708, N9701);
not NOT1 (N9709, N9706);
or OR3 (N9710, N9696, N369, N5128);
or OR4 (N9711, N9710, N3602, N2055, N2033);
buf BUF1 (N9712, N9705);
and AND3 (N9713, N9708, N3278, N3298);
nand NAND2 (N9714, N9712, N1374);
nor NOR2 (N9715, N9695, N9218);
xor XOR2 (N9716, N9714, N7181);
nor NOR2 (N9717, N9703, N519);
or OR3 (N9718, N9717, N4080, N4473);
nor NOR2 (N9719, N9698, N5749);
nor NOR2 (N9720, N9719, N3279);
buf BUF1 (N9721, N9718);
and AND4 (N9722, N9711, N6016, N6304, N8710);
nor NOR3 (N9723, N9722, N7792, N605);
nand NAND3 (N9724, N9721, N8657, N3515);
or OR4 (N9725, N9716, N7424, N4528, N85);
nand NAND3 (N9726, N9689, N1199, N4254);
not NOT1 (N9727, N9724);
buf BUF1 (N9728, N9726);
nor NOR2 (N9729, N9725, N5017);
or OR2 (N9730, N9713, N3751);
not NOT1 (N9731, N9723);
or OR3 (N9732, N9729, N5033, N8171);
and AND2 (N9733, N9728, N9529);
xor XOR2 (N9734, N9730, N7273);
nand NAND3 (N9735, N9707, N9561, N4547);
nand NAND4 (N9736, N9735, N4886, N5056, N9480);
or OR3 (N9737, N9704, N253, N1794);
xor XOR2 (N9738, N9720, N3176);
or OR3 (N9739, N9731, N5233, N8182);
buf BUF1 (N9740, N9737);
or OR3 (N9741, N9715, N2667, N6098);
nand NAND2 (N9742, N9732, N13);
nand NAND3 (N9743, N9736, N469, N9243);
nand NAND3 (N9744, N9740, N4751, N2622);
not NOT1 (N9745, N9733);
buf BUF1 (N9746, N9741);
and AND3 (N9747, N9739, N6910, N1148);
xor XOR2 (N9748, N9742, N1);
nor NOR2 (N9749, N9746, N7982);
xor XOR2 (N9750, N9749, N1429);
or OR2 (N9751, N9727, N5089);
nand NAND3 (N9752, N9748, N599, N8298);
nand NAND4 (N9753, N9747, N407, N6246, N5697);
not NOT1 (N9754, N9752);
nor NOR4 (N9755, N9754, N4959, N8391, N3572);
nand NAND3 (N9756, N9744, N117, N229);
or OR4 (N9757, N9734, N8225, N958, N7683);
nand NAND3 (N9758, N9738, N1027, N9039);
xor XOR2 (N9759, N9755, N5322);
xor XOR2 (N9760, N9756, N280);
nand NAND3 (N9761, N9709, N6578, N1059);
and AND3 (N9762, N9743, N7678, N9595);
buf BUF1 (N9763, N9750);
xor XOR2 (N9764, N9751, N939);
or OR4 (N9765, N9761, N3268, N29, N5867);
or OR3 (N9766, N9765, N8474, N9317);
xor XOR2 (N9767, N9760, N2269);
or OR2 (N9768, N9745, N6001);
not NOT1 (N9769, N9768);
buf BUF1 (N9770, N9762);
not NOT1 (N9771, N9759);
buf BUF1 (N9772, N9766);
nand NAND3 (N9773, N9769, N9655, N2780);
xor XOR2 (N9774, N9753, N5723);
nor NOR4 (N9775, N9767, N8494, N7998, N6636);
nor NOR4 (N9776, N9757, N7818, N4874, N3336);
and AND2 (N9777, N9770, N6768);
nand NAND2 (N9778, N9763, N6065);
and AND3 (N9779, N9774, N7154, N1831);
nand NAND4 (N9780, N9764, N2732, N6841, N8828);
nor NOR4 (N9781, N9780, N3275, N7491, N3645);
and AND3 (N9782, N9771, N5120, N4370);
xor XOR2 (N9783, N9772, N6955);
buf BUF1 (N9784, N9776);
and AND3 (N9785, N9781, N4424, N5521);
nor NOR2 (N9786, N9779, N5186);
and AND3 (N9787, N9786, N4662, N7034);
nor NOR2 (N9788, N9773, N2726);
nor NOR2 (N9789, N9777, N6296);
buf BUF1 (N9790, N9785);
or OR3 (N9791, N9790, N2348, N5094);
xor XOR2 (N9792, N9775, N2945);
and AND4 (N9793, N9787, N1509, N4897, N5683);
not NOT1 (N9794, N9784);
buf BUF1 (N9795, N9789);
nor NOR3 (N9796, N9793, N6059, N2897);
or OR4 (N9797, N9796, N8042, N9229, N5299);
buf BUF1 (N9798, N9797);
buf BUF1 (N9799, N9778);
or OR4 (N9800, N9792, N2335, N1265, N4158);
nand NAND2 (N9801, N9795, N8439);
buf BUF1 (N9802, N9800);
xor XOR2 (N9803, N9794, N6766);
and AND4 (N9804, N9803, N2776, N2674, N686);
buf BUF1 (N9805, N9802);
not NOT1 (N9806, N9798);
not NOT1 (N9807, N9783);
not NOT1 (N9808, N9804);
and AND3 (N9809, N9758, N4422, N3348);
nor NOR3 (N9810, N9807, N2189, N3155);
nand NAND4 (N9811, N9801, N1386, N7233, N684);
nand NAND2 (N9812, N9782, N6805);
nand NAND4 (N9813, N9812, N5560, N3565, N6503);
nand NAND4 (N9814, N9791, N4978, N2122, N7644);
nand NAND2 (N9815, N9808, N3792);
or OR4 (N9816, N9811, N7440, N6348, N2176);
xor XOR2 (N9817, N9805, N2988);
or OR4 (N9818, N9788, N7141, N128, N640);
nand NAND4 (N9819, N9817, N2542, N6924, N1979);
or OR2 (N9820, N9809, N1704);
and AND2 (N9821, N9814, N6562);
nand NAND4 (N9822, N9815, N9040, N3096, N3499);
not NOT1 (N9823, N9806);
buf BUF1 (N9824, N9821);
nand NAND2 (N9825, N9816, N8074);
nand NAND3 (N9826, N9824, N3523, N9261);
nand NAND4 (N9827, N9823, N5423, N1976, N8838);
or OR4 (N9828, N9826, N5391, N2637, N1533);
xor XOR2 (N9829, N9827, N3490);
nand NAND4 (N9830, N9813, N1378, N9125, N8212);
nor NOR2 (N9831, N9822, N1229);
xor XOR2 (N9832, N9820, N464);
or OR2 (N9833, N9799, N3152);
not NOT1 (N9834, N9819);
or OR2 (N9835, N9818, N8850);
and AND4 (N9836, N9834, N4673, N604, N4967);
nand NAND4 (N9837, N9810, N3150, N8261, N910);
buf BUF1 (N9838, N9837);
and AND2 (N9839, N9828, N1128);
nor NOR2 (N9840, N9830, N7851);
and AND3 (N9841, N9835, N1702, N6231);
nand NAND3 (N9842, N9833, N824, N4293);
xor XOR2 (N9843, N9841, N1809);
nand NAND2 (N9844, N9843, N911);
not NOT1 (N9845, N9838);
nor NOR3 (N9846, N9836, N657, N2475);
buf BUF1 (N9847, N9844);
and AND2 (N9848, N9845, N867);
buf BUF1 (N9849, N9825);
nor NOR2 (N9850, N9847, N1399);
xor XOR2 (N9851, N9839, N3024);
xor XOR2 (N9852, N9850, N9543);
buf BUF1 (N9853, N9851);
not NOT1 (N9854, N9846);
and AND2 (N9855, N9831, N9781);
nor NOR2 (N9856, N9853, N448);
xor XOR2 (N9857, N9840, N3505);
xor XOR2 (N9858, N9842, N6532);
nor NOR2 (N9859, N9857, N1810);
or OR4 (N9860, N9855, N3189, N7157, N677);
nand NAND2 (N9861, N9848, N229);
not NOT1 (N9862, N9832);
nor NOR2 (N9863, N9852, N7665);
or OR4 (N9864, N9861, N5067, N3669, N270);
buf BUF1 (N9865, N9858);
not NOT1 (N9866, N9856);
nor NOR3 (N9867, N9860, N6968, N9643);
xor XOR2 (N9868, N9849, N2181);
or OR2 (N9869, N9862, N5666);
not NOT1 (N9870, N9866);
nand NAND3 (N9871, N9863, N81, N1325);
buf BUF1 (N9872, N9854);
nor NOR3 (N9873, N9859, N6652, N8782);
xor XOR2 (N9874, N9872, N4692);
xor XOR2 (N9875, N9871, N5420);
not NOT1 (N9876, N9869);
buf BUF1 (N9877, N9865);
and AND4 (N9878, N9875, N1073, N1996, N7987);
buf BUF1 (N9879, N9878);
xor XOR2 (N9880, N9877, N4220);
nand NAND2 (N9881, N9880, N3730);
or OR4 (N9882, N9870, N9805, N1166, N4143);
or OR2 (N9883, N9829, N4268);
xor XOR2 (N9884, N9883, N4266);
nor NOR4 (N9885, N9874, N5277, N1428, N9370);
buf BUF1 (N9886, N9867);
and AND4 (N9887, N9868, N1638, N689, N3928);
buf BUF1 (N9888, N9864);
buf BUF1 (N9889, N9888);
buf BUF1 (N9890, N9886);
nor NOR3 (N9891, N9882, N1628, N3230);
buf BUF1 (N9892, N9891);
xor XOR2 (N9893, N9889, N3826);
buf BUF1 (N9894, N9892);
buf BUF1 (N9895, N9873);
nand NAND2 (N9896, N9893, N9294);
not NOT1 (N9897, N9879);
nor NOR3 (N9898, N9876, N7254, N4215);
nor NOR2 (N9899, N9887, N2034);
nor NOR3 (N9900, N9899, N1663, N7972);
nand NAND4 (N9901, N9898, N387, N8393, N9715);
nor NOR2 (N9902, N9901, N6510);
and AND4 (N9903, N9885, N2334, N6758, N1433);
nand NAND4 (N9904, N9881, N6879, N5125, N7032);
and AND2 (N9905, N9890, N2051);
xor XOR2 (N9906, N9903, N2316);
nor NOR3 (N9907, N9897, N7736, N7261);
and AND3 (N9908, N9900, N8608, N917);
nor NOR3 (N9909, N9904, N6371, N830);
xor XOR2 (N9910, N9894, N1332);
not NOT1 (N9911, N9907);
and AND3 (N9912, N9905, N1920, N2583);
nor NOR4 (N9913, N9911, N4412, N1216, N6043);
and AND2 (N9914, N9910, N9436);
and AND2 (N9915, N9914, N1619);
not NOT1 (N9916, N9902);
or OR3 (N9917, N9896, N2687, N992);
nand NAND2 (N9918, N9908, N6398);
or OR3 (N9919, N9909, N7963, N7613);
nand NAND2 (N9920, N9918, N9491);
xor XOR2 (N9921, N9895, N9342);
nand NAND3 (N9922, N9906, N6916, N8387);
xor XOR2 (N9923, N9884, N4923);
and AND4 (N9924, N9919, N8067, N8491, N7998);
nand NAND2 (N9925, N9912, N5706);
nor NOR3 (N9926, N9915, N1416, N1030);
and AND2 (N9927, N9921, N195);
not NOT1 (N9928, N9924);
not NOT1 (N9929, N9913);
or OR3 (N9930, N9927, N5311, N6);
and AND4 (N9931, N9929, N1588, N2499, N757);
or OR4 (N9932, N9931, N3701, N929, N9323);
buf BUF1 (N9933, N9926);
and AND3 (N9934, N9928, N4558, N251);
nand NAND3 (N9935, N9923, N2687, N2053);
and AND2 (N9936, N9922, N4061);
buf BUF1 (N9937, N9933);
or OR3 (N9938, N9925, N7399, N6530);
or OR3 (N9939, N9935, N9276, N4477);
not NOT1 (N9940, N9916);
xor XOR2 (N9941, N9940, N661);
nor NOR2 (N9942, N9937, N2812);
nor NOR2 (N9943, N9930, N4318);
xor XOR2 (N9944, N9936, N6190);
not NOT1 (N9945, N9942);
or OR3 (N9946, N9941, N1272, N9185);
buf BUF1 (N9947, N9938);
xor XOR2 (N9948, N9944, N1648);
nor NOR4 (N9949, N9932, N653, N3203, N1372);
nand NAND4 (N9950, N9934, N4528, N7651, N1088);
and AND2 (N9951, N9943, N1210);
xor XOR2 (N9952, N9951, N812);
nand NAND3 (N9953, N9917, N2151, N3300);
not NOT1 (N9954, N9949);
nor NOR4 (N9955, N9954, N1309, N1483, N7770);
and AND2 (N9956, N9950, N2650);
nor NOR2 (N9957, N9945, N8346);
xor XOR2 (N9958, N9957, N2118);
nand NAND4 (N9959, N9956, N6827, N7041, N4622);
or OR2 (N9960, N9952, N4920);
nor NOR3 (N9961, N9947, N6103, N5249);
not NOT1 (N9962, N9955);
xor XOR2 (N9963, N9939, N7610);
nand NAND2 (N9964, N9960, N9667);
xor XOR2 (N9965, N9958, N4824);
buf BUF1 (N9966, N9964);
buf BUF1 (N9967, N9920);
not NOT1 (N9968, N9962);
buf BUF1 (N9969, N9968);
and AND4 (N9970, N9967, N6642, N1845, N6949);
nor NOR2 (N9971, N9959, N3512);
buf BUF1 (N9972, N9966);
buf BUF1 (N9973, N9963);
not NOT1 (N9974, N9971);
not NOT1 (N9975, N9970);
not NOT1 (N9976, N9969);
or OR2 (N9977, N9953, N3108);
nand NAND2 (N9978, N9948, N4304);
and AND2 (N9979, N9965, N5310);
and AND3 (N9980, N9972, N5121, N808);
nor NOR4 (N9981, N9980, N435, N7833, N6629);
nand NAND4 (N9982, N9978, N1117, N1832, N8983);
nand NAND2 (N9983, N9981, N6674);
nor NOR4 (N9984, N9982, N7203, N1614, N3791);
nor NOR3 (N9985, N9976, N3374, N6012);
buf BUF1 (N9986, N9975);
and AND4 (N9987, N9985, N626, N5708, N9194);
not NOT1 (N9988, N9977);
xor XOR2 (N9989, N9983, N6815);
xor XOR2 (N9990, N9987, N3953);
nor NOR4 (N9991, N9979, N3623, N1388, N8367);
buf BUF1 (N9992, N9986);
buf BUF1 (N9993, N9946);
and AND3 (N9994, N9974, N3513, N471);
and AND4 (N9995, N9961, N7046, N8670, N9126);
nand NAND4 (N9996, N9990, N8110, N7805, N7833);
buf BUF1 (N9997, N9995);
buf BUF1 (N9998, N9988);
not NOT1 (N9999, N9984);
and AND4 (N10000, N9993, N5612, N2946, N1239);
xor XOR2 (N10001, N9989, N1948);
nand NAND3 (N10002, N9997, N3236, N5003);
nor NOR3 (N10003, N9998, N4687, N5260);
nand NAND4 (N10004, N10003, N5138, N367, N1223);
or OR2 (N10005, N10000, N5405);
xor XOR2 (N10006, N9992, N2013);
nor NOR3 (N10007, N10005, N7490, N8303);
or OR4 (N10008, N9991, N6833, N6918, N1067);
nand NAND3 (N10009, N9996, N5311, N8694);
buf BUF1 (N10010, N9994);
xor XOR2 (N10011, N9973, N7237);
not NOT1 (N10012, N10009);
buf BUF1 (N10013, N10010);
or OR3 (N10014, N10004, N4193, N1356);
buf BUF1 (N10015, N10006);
not NOT1 (N10016, N9999);
not NOT1 (N10017, N10012);
not NOT1 (N10018, N10015);
nor NOR4 (N10019, N10008, N6107, N2481, N2690);
nand NAND3 (N10020, N10007, N600, N52);
buf BUF1 (N10021, N10011);
nor NOR2 (N10022, N10014, N247);
and AND2 (N10023, N10016, N4090);
nor NOR4 (N10024, N10001, N2455, N4014, N3158);
and AND3 (N10025, N10021, N231, N3813);
not NOT1 (N10026, N10013);
nand NAND3 (N10027, N10017, N4611, N5048);
nand NAND2 (N10028, N10022, N6840);
nor NOR3 (N10029, N10023, N3851, N8642);
buf BUF1 (N10030, N10024);
xor XOR2 (N10031, N10025, N2082);
or OR3 (N10032, N10029, N5289, N3289);
buf BUF1 (N10033, N10030);
xor XOR2 (N10034, N10028, N4964);
or OR2 (N10035, N10027, N8892);
xor XOR2 (N10036, N10020, N8786);
buf BUF1 (N10037, N10002);
or OR2 (N10038, N10032, N5386);
and AND3 (N10039, N10036, N2421, N5046);
or OR3 (N10040, N10031, N3724, N3344);
buf BUF1 (N10041, N10026);
nor NOR3 (N10042, N10040, N5266, N2226);
or OR2 (N10043, N10019, N3996);
not NOT1 (N10044, N10035);
nor NOR4 (N10045, N10039, N6365, N2064, N6065);
not NOT1 (N10046, N10038);
buf BUF1 (N10047, N10018);
nor NOR2 (N10048, N10042, N8464);
nand NAND4 (N10049, N10034, N3555, N6452, N6995);
and AND2 (N10050, N10033, N3767);
or OR3 (N10051, N10045, N183, N2511);
buf BUF1 (N10052, N10050);
nand NAND4 (N10053, N10052, N3586, N4110, N6616);
buf BUF1 (N10054, N10046);
and AND4 (N10055, N10043, N8217, N8658, N6827);
nand NAND3 (N10056, N10055, N10, N7238);
nand NAND3 (N10057, N10041, N7641, N4651);
or OR4 (N10058, N10047, N5443, N6472, N2190);
buf BUF1 (N10059, N10058);
and AND2 (N10060, N10056, N4658);
not NOT1 (N10061, N10048);
nor NOR4 (N10062, N10051, N6882, N6790, N3864);
buf BUF1 (N10063, N10059);
buf BUF1 (N10064, N10063);
nor NOR2 (N10065, N10053, N6878);
or OR3 (N10066, N10057, N7190, N2999);
nor NOR3 (N10067, N10061, N2171, N7496);
buf BUF1 (N10068, N10054);
xor XOR2 (N10069, N10065, N695);
nor NOR4 (N10070, N10049, N4762, N2897, N9920);
not NOT1 (N10071, N10064);
nand NAND4 (N10072, N10066, N1432, N6605, N7786);
xor XOR2 (N10073, N10037, N2259);
buf BUF1 (N10074, N10073);
nor NOR2 (N10075, N10069, N3998);
buf BUF1 (N10076, N10060);
and AND3 (N10077, N10074, N1684, N9588);
nor NOR4 (N10078, N10068, N8583, N2676, N8870);
and AND4 (N10079, N10076, N3150, N9991, N6176);
nand NAND2 (N10080, N10078, N622);
not NOT1 (N10081, N10044);
or OR4 (N10082, N10077, N7141, N7968, N462);
and AND3 (N10083, N10081, N7637, N6904);
or OR3 (N10084, N10071, N4386, N2512);
nor NOR3 (N10085, N10062, N29, N7169);
not NOT1 (N10086, N10085);
nand NAND4 (N10087, N10075, N4530, N1170, N6655);
buf BUF1 (N10088, N10082);
buf BUF1 (N10089, N10072);
nor NOR2 (N10090, N10089, N2368);
or OR4 (N10091, N10083, N6629, N6718, N1755);
nor NOR4 (N10092, N10079, N9400, N3949, N1709);
nand NAND4 (N10093, N10090, N2221, N8013, N709);
nand NAND4 (N10094, N10084, N1992, N5972, N8404);
and AND2 (N10095, N10070, N5144);
nor NOR4 (N10096, N10094, N9210, N5890, N2345);
not NOT1 (N10097, N10080);
nand NAND3 (N10098, N10092, N2797, N8241);
nand NAND2 (N10099, N10091, N3548);
xor XOR2 (N10100, N10099, N7397);
nor NOR4 (N10101, N10086, N240, N7025, N7952);
nand NAND2 (N10102, N10088, N1837);
and AND3 (N10103, N10098, N5068, N9327);
nor NOR4 (N10104, N10095, N2318, N1613, N2580);
and AND2 (N10105, N10096, N112);
nor NOR3 (N10106, N10093, N5571, N6629);
nor NOR4 (N10107, N10100, N8841, N1631, N7008);
nand NAND4 (N10108, N10106, N281, N975, N1652);
buf BUF1 (N10109, N10108);
nor NOR3 (N10110, N10104, N691, N2897);
and AND4 (N10111, N10097, N4900, N4141, N6243);
buf BUF1 (N10112, N10101);
and AND3 (N10113, N10102, N3774, N1599);
and AND2 (N10114, N10113, N7911);
or OR2 (N10115, N10087, N4899);
buf BUF1 (N10116, N10115);
xor XOR2 (N10117, N10116, N9570);
xor XOR2 (N10118, N10067, N3454);
or OR4 (N10119, N10110, N8834, N5511, N2033);
xor XOR2 (N10120, N10109, N8360);
xor XOR2 (N10121, N10120, N8392);
nor NOR2 (N10122, N10114, N8510);
not NOT1 (N10123, N10119);
not NOT1 (N10124, N10107);
and AND4 (N10125, N10121, N672, N3788, N8564);
nor NOR3 (N10126, N10111, N259, N2936);
buf BUF1 (N10127, N10125);
not NOT1 (N10128, N10122);
and AND2 (N10129, N10103, N6774);
nor NOR3 (N10130, N10105, N2817, N6501);
xor XOR2 (N10131, N10124, N6543);
buf BUF1 (N10132, N10112);
nor NOR3 (N10133, N10131, N1858, N196);
not NOT1 (N10134, N10129);
xor XOR2 (N10135, N10127, N9058);
not NOT1 (N10136, N10132);
nor NOR3 (N10137, N10126, N299, N6342);
buf BUF1 (N10138, N10137);
not NOT1 (N10139, N10128);
xor XOR2 (N10140, N10135, N8047);
buf BUF1 (N10141, N10134);
xor XOR2 (N10142, N10118, N4646);
not NOT1 (N10143, N10117);
not NOT1 (N10144, N10136);
and AND3 (N10145, N10140, N3549, N9383);
nor NOR4 (N10146, N10145, N9409, N6052, N9889);
and AND3 (N10147, N10143, N4579, N9338);
or OR2 (N10148, N10139, N2109);
xor XOR2 (N10149, N10146, N1167);
not NOT1 (N10150, N10123);
nand NAND2 (N10151, N10147, N905);
nand NAND2 (N10152, N10150, N3874);
buf BUF1 (N10153, N10142);
and AND2 (N10154, N10133, N5077);
nand NAND3 (N10155, N10152, N2846, N5443);
xor XOR2 (N10156, N10148, N9756);
or OR2 (N10157, N10153, N4219);
nand NAND2 (N10158, N10157, N4682);
not NOT1 (N10159, N10141);
buf BUF1 (N10160, N10151);
or OR4 (N10161, N10138, N9484, N8143, N2935);
xor XOR2 (N10162, N10160, N1705);
xor XOR2 (N10163, N10154, N4048);
xor XOR2 (N10164, N10156, N8592);
nand NAND3 (N10165, N10161, N2049, N1339);
buf BUF1 (N10166, N10155);
and AND2 (N10167, N10164, N6820);
buf BUF1 (N10168, N10144);
buf BUF1 (N10169, N10158);
buf BUF1 (N10170, N10166);
xor XOR2 (N10171, N10162, N469);
buf BUF1 (N10172, N10163);
nand NAND4 (N10173, N10149, N6640, N6662, N5837);
nand NAND2 (N10174, N10171, N3036);
buf BUF1 (N10175, N10169);
and AND4 (N10176, N10170, N5297, N9667, N5864);
not NOT1 (N10177, N10172);
or OR3 (N10178, N10176, N1632, N9616);
buf BUF1 (N10179, N10168);
not NOT1 (N10180, N10173);
and AND4 (N10181, N10167, N136, N8150, N6297);
buf BUF1 (N10182, N10179);
or OR2 (N10183, N10165, N5105);
nand NAND4 (N10184, N10177, N7726, N1157, N6319);
buf BUF1 (N10185, N10181);
nor NOR2 (N10186, N10180, N5267);
xor XOR2 (N10187, N10183, N301);
nor NOR4 (N10188, N10178, N3886, N5132, N3189);
or OR2 (N10189, N10174, N4616);
not NOT1 (N10190, N10187);
and AND4 (N10191, N10182, N5606, N9527, N8688);
nor NOR2 (N10192, N10190, N246);
nand NAND2 (N10193, N10192, N4130);
nand NAND4 (N10194, N10130, N2492, N7207, N2166);
or OR4 (N10195, N10191, N1075, N5439, N3242);
not NOT1 (N10196, N10185);
or OR3 (N10197, N10184, N5944, N3346);
xor XOR2 (N10198, N10175, N3743);
nand NAND3 (N10199, N10194, N4106, N9334);
and AND3 (N10200, N10188, N5594, N9725);
nand NAND3 (N10201, N10196, N4700, N3680);
and AND4 (N10202, N10199, N8859, N3075, N6322);
nor NOR3 (N10203, N10197, N3961, N5191);
not NOT1 (N10204, N10201);
not NOT1 (N10205, N10202);
nand NAND2 (N10206, N10189, N4215);
nand NAND2 (N10207, N10186, N7276);
xor XOR2 (N10208, N10206, N1824);
xor XOR2 (N10209, N10198, N2239);
nor NOR2 (N10210, N10200, N870);
not NOT1 (N10211, N10204);
or OR3 (N10212, N10203, N6163, N4295);
not NOT1 (N10213, N10195);
buf BUF1 (N10214, N10159);
buf BUF1 (N10215, N10213);
and AND2 (N10216, N10205, N2375);
nor NOR4 (N10217, N10214, N2043, N5897, N2449);
nand NAND4 (N10218, N10193, N3052, N6166, N4719);
buf BUF1 (N10219, N10212);
or OR2 (N10220, N10218, N210);
xor XOR2 (N10221, N10210, N8415);
xor XOR2 (N10222, N10215, N4098);
xor XOR2 (N10223, N10209, N2106);
xor XOR2 (N10224, N10208, N9408);
or OR3 (N10225, N10220, N5771, N9127);
nand NAND2 (N10226, N10216, N5094);
xor XOR2 (N10227, N10211, N7878);
nand NAND4 (N10228, N10224, N1509, N9078, N10195);
not NOT1 (N10229, N10226);
or OR4 (N10230, N10229, N5996, N6295, N1881);
nand NAND3 (N10231, N10228, N7547, N7031);
not NOT1 (N10232, N10231);
xor XOR2 (N10233, N10217, N4361);
nor NOR3 (N10234, N10225, N2088, N4323);
buf BUF1 (N10235, N10207);
and AND4 (N10236, N10232, N183, N5101, N8557);
not NOT1 (N10237, N10222);
buf BUF1 (N10238, N10234);
buf BUF1 (N10239, N10221);
buf BUF1 (N10240, N10236);
nor NOR2 (N10241, N10219, N5114);
buf BUF1 (N10242, N10233);
and AND3 (N10243, N10238, N5714, N7463);
not NOT1 (N10244, N10240);
buf BUF1 (N10245, N10242);
or OR4 (N10246, N10245, N4467, N3120, N8794);
xor XOR2 (N10247, N10223, N9431);
buf BUF1 (N10248, N10241);
xor XOR2 (N10249, N10244, N2850);
or OR4 (N10250, N10235, N633, N6568, N7679);
and AND3 (N10251, N10239, N8145, N3759);
or OR3 (N10252, N10230, N7707, N1250);
buf BUF1 (N10253, N10251);
and AND4 (N10254, N10253, N7860, N3339, N7216);
or OR2 (N10255, N10248, N7708);
nand NAND4 (N10256, N10249, N171, N3258, N9355);
and AND4 (N10257, N10254, N9788, N9663, N9596);
not NOT1 (N10258, N10247);
nand NAND4 (N10259, N10246, N4513, N5011, N2911);
or OR2 (N10260, N10259, N471);
nand NAND3 (N10261, N10256, N9301, N4633);
or OR4 (N10262, N10243, N7690, N9448, N2929);
not NOT1 (N10263, N10227);
and AND2 (N10264, N10250, N2110);
nand NAND3 (N10265, N10255, N831, N9846);
buf BUF1 (N10266, N10252);
buf BUF1 (N10267, N10264);
xor XOR2 (N10268, N10265, N9417);
nand NAND2 (N10269, N10257, N8710);
xor XOR2 (N10270, N10237, N8828);
nor NOR4 (N10271, N10261, N4675, N9909, N3513);
xor XOR2 (N10272, N10270, N8325);
buf BUF1 (N10273, N10268);
and AND3 (N10274, N10262, N2022, N8183);
xor XOR2 (N10275, N10269, N7119);
xor XOR2 (N10276, N10266, N7415);
buf BUF1 (N10277, N10274);
and AND4 (N10278, N10273, N6487, N6496, N5866);
buf BUF1 (N10279, N10260);
nand NAND2 (N10280, N10267, N10172);
or OR3 (N10281, N10277, N9838, N4147);
xor XOR2 (N10282, N10281, N441);
not NOT1 (N10283, N10278);
and AND2 (N10284, N10258, N5161);
not NOT1 (N10285, N10271);
buf BUF1 (N10286, N10280);
buf BUF1 (N10287, N10263);
not NOT1 (N10288, N10283);
not NOT1 (N10289, N10282);
or OR3 (N10290, N10286, N1301, N8350);
xor XOR2 (N10291, N10287, N5844);
not NOT1 (N10292, N10284);
buf BUF1 (N10293, N10276);
buf BUF1 (N10294, N10289);
and AND4 (N10295, N10291, N3196, N9783, N253);
nand NAND3 (N10296, N10279, N3190, N3367);
or OR2 (N10297, N10293, N7868);
xor XOR2 (N10298, N10292, N1842);
xor XOR2 (N10299, N10295, N4357);
and AND3 (N10300, N10288, N3119, N3018);
not NOT1 (N10301, N10298);
buf BUF1 (N10302, N10275);
nand NAND2 (N10303, N10300, N10039);
nand NAND3 (N10304, N10296, N514, N1704);
nor NOR4 (N10305, N10297, N7012, N524, N2943);
not NOT1 (N10306, N10272);
not NOT1 (N10307, N10305);
xor XOR2 (N10308, N10285, N5931);
and AND4 (N10309, N10299, N8780, N9411, N8564);
nor NOR3 (N10310, N10304, N5822, N558);
not NOT1 (N10311, N10307);
and AND3 (N10312, N10303, N5351, N10257);
buf BUF1 (N10313, N10311);
buf BUF1 (N10314, N10313);
and AND4 (N10315, N10294, N4782, N4607, N4566);
and AND4 (N10316, N10301, N4079, N681, N4547);
nand NAND4 (N10317, N10314, N1748, N1504, N8632);
nand NAND2 (N10318, N10316, N1319);
or OR3 (N10319, N10312, N8819, N8525);
nand NAND2 (N10320, N10308, N4178);
or OR4 (N10321, N10306, N2947, N4821, N9845);
xor XOR2 (N10322, N10309, N3294);
nand NAND3 (N10323, N10315, N4128, N2839);
nand NAND4 (N10324, N10320, N70, N352, N3881);
xor XOR2 (N10325, N10324, N979);
nor NOR2 (N10326, N10310, N7597);
nor NOR2 (N10327, N10326, N3595);
buf BUF1 (N10328, N10317);
nand NAND4 (N10329, N10318, N3171, N8375, N9515);
nand NAND3 (N10330, N10319, N7000, N6500);
xor XOR2 (N10331, N10328, N3616);
nand NAND2 (N10332, N10321, N8247);
and AND3 (N10333, N10302, N5640, N5985);
or OR3 (N10334, N10331, N4645, N2466);
xor XOR2 (N10335, N10333, N1519);
not NOT1 (N10336, N10334);
nand NAND2 (N10337, N10329, N5164);
nand NAND3 (N10338, N10325, N10039, N8278);
xor XOR2 (N10339, N10290, N6340);
buf BUF1 (N10340, N10330);
or OR2 (N10341, N10335, N8998);
or OR2 (N10342, N10340, N1773);
or OR2 (N10343, N10323, N6900);
nand NAND4 (N10344, N10322, N4297, N7141, N9880);
nand NAND3 (N10345, N10344, N58, N8538);
nor NOR4 (N10346, N10336, N7938, N7910, N5689);
or OR2 (N10347, N10345, N3232);
nor NOR2 (N10348, N10342, N7907);
xor XOR2 (N10349, N10348, N4068);
and AND2 (N10350, N10338, N10142);
nand NAND2 (N10351, N10347, N5652);
nor NOR4 (N10352, N10349, N323, N1530, N3581);
not NOT1 (N10353, N10350);
not NOT1 (N10354, N10343);
xor XOR2 (N10355, N10339, N7710);
not NOT1 (N10356, N10337);
nand NAND2 (N10357, N10356, N2589);
not NOT1 (N10358, N10341);
xor XOR2 (N10359, N10351, N718);
buf BUF1 (N10360, N10359);
nor NOR3 (N10361, N10357, N694, N1808);
nand NAND2 (N10362, N10327, N7260);
or OR3 (N10363, N10346, N8189, N6872);
and AND2 (N10364, N10352, N732);
or OR4 (N10365, N10358, N2295, N3971, N7667);
buf BUF1 (N10366, N10355);
not NOT1 (N10367, N10332);
and AND2 (N10368, N10354, N1852);
or OR2 (N10369, N10368, N1055);
or OR3 (N10370, N10366, N7233, N3722);
xor XOR2 (N10371, N10353, N2174);
or OR2 (N10372, N10361, N6299);
not NOT1 (N10373, N10372);
nor NOR4 (N10374, N10369, N2781, N4940, N9341);
buf BUF1 (N10375, N10370);
nand NAND3 (N10376, N10373, N2705, N3986);
not NOT1 (N10377, N10365);
not NOT1 (N10378, N10374);
or OR2 (N10379, N10371, N3377);
nor NOR3 (N10380, N10377, N1312, N1753);
nor NOR3 (N10381, N10375, N984, N4845);
or OR3 (N10382, N10381, N9833, N3972);
nand NAND2 (N10383, N10364, N4212);
buf BUF1 (N10384, N10367);
nor NOR3 (N10385, N10363, N6727, N8329);
buf BUF1 (N10386, N10360);
and AND4 (N10387, N10378, N5064, N6228, N2928);
not NOT1 (N10388, N10382);
and AND4 (N10389, N10385, N7752, N6663, N2505);
and AND2 (N10390, N10387, N3846);
nand NAND3 (N10391, N10386, N3039, N7500);
and AND2 (N10392, N10379, N7708);
and AND4 (N10393, N10389, N5866, N4485, N2579);
nand NAND2 (N10394, N10383, N1055);
not NOT1 (N10395, N10384);
xor XOR2 (N10396, N10380, N4514);
buf BUF1 (N10397, N10362);
xor XOR2 (N10398, N10396, N2180);
or OR4 (N10399, N10395, N2018, N8694, N440);
buf BUF1 (N10400, N10392);
and AND4 (N10401, N10376, N9986, N6626, N1008);
nor NOR4 (N10402, N10388, N5721, N7476, N1659);
not NOT1 (N10403, N10400);
and AND3 (N10404, N10399, N2356, N6625);
or OR4 (N10405, N10401, N9612, N3606, N9656);
xor XOR2 (N10406, N10402, N3209);
not NOT1 (N10407, N10406);
buf BUF1 (N10408, N10394);
and AND4 (N10409, N10391, N9221, N745, N5935);
or OR2 (N10410, N10398, N2206);
or OR2 (N10411, N10407, N8115);
not NOT1 (N10412, N10404);
xor XOR2 (N10413, N10411, N5114);
or OR2 (N10414, N10412, N1842);
xor XOR2 (N10415, N10393, N1440);
nor NOR2 (N10416, N10408, N10228);
buf BUF1 (N10417, N10413);
and AND4 (N10418, N10415, N6775, N8203, N6053);
nor NOR2 (N10419, N10409, N1697);
xor XOR2 (N10420, N10397, N61);
xor XOR2 (N10421, N10414, N7671);
or OR2 (N10422, N10419, N157);
not NOT1 (N10423, N10405);
not NOT1 (N10424, N10423);
nor NOR4 (N10425, N10417, N8218, N7172, N3041);
nand NAND4 (N10426, N10421, N5001, N8299, N4167);
or OR3 (N10427, N10403, N5469, N5446);
nand NAND3 (N10428, N10422, N3295, N5544);
and AND3 (N10429, N10418, N6035, N6143);
and AND3 (N10430, N10429, N5525, N6460);
nand NAND3 (N10431, N10430, N3981, N3439);
or OR3 (N10432, N10427, N10180, N5311);
or OR4 (N10433, N10424, N1531, N7476, N237);
and AND3 (N10434, N10426, N6747, N7805);
or OR3 (N10435, N10428, N3750, N5467);
buf BUF1 (N10436, N10416);
nand NAND4 (N10437, N10433, N2214, N4918, N1149);
nand NAND4 (N10438, N10425, N3991, N9488, N2600);
xor XOR2 (N10439, N10435, N431);
or OR3 (N10440, N10410, N9996, N7872);
and AND3 (N10441, N10439, N8998, N707);
xor XOR2 (N10442, N10436, N2412);
and AND3 (N10443, N10390, N8282, N9887);
xor XOR2 (N10444, N10441, N853);
nand NAND2 (N10445, N10434, N7575);
or OR2 (N10446, N10444, N3884);
and AND4 (N10447, N10443, N1749, N10339, N10166);
not NOT1 (N10448, N10431);
nor NOR2 (N10449, N10445, N965);
nor NOR4 (N10450, N10438, N7042, N9470, N4241);
nand NAND2 (N10451, N10432, N5079);
and AND2 (N10452, N10440, N1178);
or OR3 (N10453, N10442, N8683, N2679);
xor XOR2 (N10454, N10449, N7656);
and AND3 (N10455, N10451, N7681, N3051);
buf BUF1 (N10456, N10450);
or OR2 (N10457, N10447, N4382);
and AND4 (N10458, N10456, N3405, N1633, N1366);
xor XOR2 (N10459, N10453, N4381);
xor XOR2 (N10460, N10455, N1625);
xor XOR2 (N10461, N10446, N10135);
and AND2 (N10462, N10420, N3022);
not NOT1 (N10463, N10459);
nor NOR2 (N10464, N10448, N8341);
nor NOR2 (N10465, N10457, N5138);
xor XOR2 (N10466, N10454, N6984);
buf BUF1 (N10467, N10458);
and AND2 (N10468, N10463, N9638);
buf BUF1 (N10469, N10468);
buf BUF1 (N10470, N10452);
buf BUF1 (N10471, N10465);
not NOT1 (N10472, N10461);
not NOT1 (N10473, N10437);
not NOT1 (N10474, N10462);
nor NOR3 (N10475, N10474, N426, N9196);
not NOT1 (N10476, N10466);
nor NOR4 (N10477, N10460, N5735, N9443, N4245);
buf BUF1 (N10478, N10475);
nand NAND3 (N10479, N10471, N6074, N3453);
xor XOR2 (N10480, N10476, N4471);
nor NOR4 (N10481, N10478, N6794, N9506, N8267);
or OR3 (N10482, N10480, N5752, N8786);
and AND4 (N10483, N10472, N10462, N8837, N1457);
and AND4 (N10484, N10482, N4185, N9100, N9144);
nand NAND2 (N10485, N10479, N1601);
xor XOR2 (N10486, N10464, N6606);
xor XOR2 (N10487, N10469, N3210);
or OR2 (N10488, N10481, N4876);
buf BUF1 (N10489, N10467);
buf BUF1 (N10490, N10483);
nand NAND3 (N10491, N10473, N446, N9564);
and AND3 (N10492, N10470, N7141, N4156);
nand NAND3 (N10493, N10487, N9516, N3890);
xor XOR2 (N10494, N10489, N119);
nor NOR4 (N10495, N10492, N936, N7703, N7216);
or OR3 (N10496, N10488, N2983, N3168);
nor NOR4 (N10497, N10486, N1307, N4070, N10232);
not NOT1 (N10498, N10494);
nor NOR3 (N10499, N10498, N1769, N6088);
and AND3 (N10500, N10491, N2299, N2688);
not NOT1 (N10501, N10499);
xor XOR2 (N10502, N10477, N8746);
and AND2 (N10503, N10484, N2823);
nor NOR3 (N10504, N10503, N3781, N6607);
xor XOR2 (N10505, N10497, N8810);
and AND3 (N10506, N10500, N3176, N9637);
or OR4 (N10507, N10485, N9843, N3730, N5050);
or OR4 (N10508, N10507, N5062, N9790, N6600);
xor XOR2 (N10509, N10506, N4465);
or OR2 (N10510, N10509, N8773);
and AND4 (N10511, N10493, N3587, N7107, N9005);
not NOT1 (N10512, N10496);
nor NOR3 (N10513, N10490, N6332, N6053);
not NOT1 (N10514, N10508);
buf BUF1 (N10515, N10510);
buf BUF1 (N10516, N10495);
or OR3 (N10517, N10511, N6456, N6143);
and AND2 (N10518, N10515, N1569);
buf BUF1 (N10519, N10505);
buf BUF1 (N10520, N10501);
buf BUF1 (N10521, N10519);
nand NAND4 (N10522, N10516, N9554, N5843, N2923);
nor NOR3 (N10523, N10520, N1855, N214);
or OR4 (N10524, N10512, N2004, N6818, N1418);
and AND4 (N10525, N10521, N7004, N4155, N1412);
or OR4 (N10526, N10524, N6699, N5453, N68);
and AND4 (N10527, N10514, N2256, N2230, N10375);
buf BUF1 (N10528, N10504);
nand NAND4 (N10529, N10517, N6357, N5965, N3920);
nand NAND4 (N10530, N10528, N4161, N1311, N149);
nand NAND4 (N10531, N10527, N2862, N7660, N6283);
nor NOR3 (N10532, N10513, N8342, N8889);
and AND2 (N10533, N10530, N7526);
nor NOR4 (N10534, N10522, N6454, N3471, N3550);
xor XOR2 (N10535, N10533, N5588);
nor NOR4 (N10536, N10535, N212, N5596, N2957);
xor XOR2 (N10537, N10518, N8784);
buf BUF1 (N10538, N10536);
not NOT1 (N10539, N10538);
buf BUF1 (N10540, N10523);
nand NAND4 (N10541, N10534, N2545, N1568, N5861);
nand NAND3 (N10542, N10537, N1543, N658);
nor NOR3 (N10543, N10539, N6156, N3241);
or OR2 (N10544, N10502, N41);
nor NOR2 (N10545, N10540, N1612);
xor XOR2 (N10546, N10542, N7973);
or OR2 (N10547, N10525, N7877);
nand NAND4 (N10548, N10529, N3453, N8546, N5019);
buf BUF1 (N10549, N10531);
or OR2 (N10550, N10548, N8715);
and AND4 (N10551, N10547, N7280, N3658, N9277);
and AND3 (N10552, N10526, N4747, N1584);
nor NOR3 (N10553, N10551, N3817, N1309);
nand NAND2 (N10554, N10545, N2654);
xor XOR2 (N10555, N10532, N7188);
and AND2 (N10556, N10543, N9830);
not NOT1 (N10557, N10554);
or OR4 (N10558, N10541, N3372, N5651, N1133);
and AND4 (N10559, N10553, N7705, N7354, N5381);
xor XOR2 (N10560, N10557, N2301);
or OR3 (N10561, N10558, N8138, N3302);
and AND4 (N10562, N10561, N8900, N5224, N1026);
not NOT1 (N10563, N10556);
nand NAND3 (N10564, N10562, N6695, N6405);
nand NAND3 (N10565, N10560, N5015, N1058);
or OR3 (N10566, N10550, N7414, N5988);
buf BUF1 (N10567, N10565);
or OR3 (N10568, N10544, N7386, N2049);
nand NAND2 (N10569, N10566, N8465);
nand NAND3 (N10570, N10568, N3375, N1352);
nand NAND3 (N10571, N10563, N322, N3090);
and AND3 (N10572, N10564, N6012, N5260);
not NOT1 (N10573, N10559);
xor XOR2 (N10574, N10572, N8623);
nand NAND2 (N10575, N10573, N9288);
xor XOR2 (N10576, N10567, N165);
nand NAND3 (N10577, N10570, N10359, N5461);
nand NAND3 (N10578, N10575, N1083, N5188);
xor XOR2 (N10579, N10549, N733);
or OR2 (N10580, N10571, N9977);
nor NOR2 (N10581, N10555, N9995);
nor NOR2 (N10582, N10569, N57);
or OR4 (N10583, N10576, N4630, N6492, N357);
not NOT1 (N10584, N10546);
or OR4 (N10585, N10583, N1799, N9803, N2008);
buf BUF1 (N10586, N10581);
xor XOR2 (N10587, N10578, N4911);
or OR2 (N10588, N10587, N1064);
and AND2 (N10589, N10584, N2157);
nand NAND4 (N10590, N10589, N6858, N1439, N691);
nor NOR3 (N10591, N10585, N9721, N9464);
nor NOR2 (N10592, N10574, N911);
buf BUF1 (N10593, N10591);
xor XOR2 (N10594, N10580, N2380);
nor NOR4 (N10595, N10579, N8639, N5282, N2555);
not NOT1 (N10596, N10552);
xor XOR2 (N10597, N10586, N2292);
and AND2 (N10598, N10593, N9748);
xor XOR2 (N10599, N10598, N9094);
nand NAND3 (N10600, N10582, N3001, N8121);
nor NOR2 (N10601, N10596, N4559);
not NOT1 (N10602, N10599);
and AND4 (N10603, N10602, N6798, N8287, N4666);
or OR2 (N10604, N10597, N212);
nor NOR3 (N10605, N10604, N7861, N1984);
or OR3 (N10606, N10595, N4083, N2075);
nand NAND4 (N10607, N10603, N10163, N8043, N6789);
xor XOR2 (N10608, N10594, N784);
nand NAND2 (N10609, N10590, N2207);
nand NAND2 (N10610, N10605, N2662);
or OR2 (N10611, N10607, N3462);
nand NAND2 (N10612, N10609, N8683);
nor NOR3 (N10613, N10592, N7771, N5096);
xor XOR2 (N10614, N10577, N10159);
or OR4 (N10615, N10610, N4148, N4082, N3587);
nand NAND4 (N10616, N10613, N9270, N2227, N10485);
and AND2 (N10617, N10601, N6053);
or OR2 (N10618, N10611, N5953);
not NOT1 (N10619, N10588);
nand NAND3 (N10620, N10612, N1568, N4672);
not NOT1 (N10621, N10600);
not NOT1 (N10622, N10617);
and AND4 (N10623, N10620, N6783, N6001, N3495);
or OR3 (N10624, N10622, N9251, N5925);
nand NAND2 (N10625, N10616, N2726);
buf BUF1 (N10626, N10621);
nand NAND4 (N10627, N10623, N1528, N163, N6690);
or OR4 (N10628, N10619, N6050, N7905, N6398);
or OR2 (N10629, N10618, N605);
buf BUF1 (N10630, N10625);
nand NAND2 (N10631, N10624, N6701);
nand NAND4 (N10632, N10627, N2701, N4091, N4118);
nand NAND2 (N10633, N10628, N9533);
buf BUF1 (N10634, N10629);
not NOT1 (N10635, N10606);
or OR2 (N10636, N10614, N8803);
nand NAND2 (N10637, N10626, N5662);
or OR3 (N10638, N10608, N6592, N6263);
buf BUF1 (N10639, N10633);
buf BUF1 (N10640, N10615);
xor XOR2 (N10641, N10638, N7939);
not NOT1 (N10642, N10641);
buf BUF1 (N10643, N10639);
buf BUF1 (N10644, N10637);
not NOT1 (N10645, N10632);
nand NAND3 (N10646, N10640, N7830, N3550);
and AND4 (N10647, N10646, N892, N7372, N3601);
nor NOR4 (N10648, N10644, N1632, N9987, N3993);
and AND2 (N10649, N10635, N9295);
and AND2 (N10650, N10647, N5167);
and AND3 (N10651, N10642, N10080, N4746);
nor NOR3 (N10652, N10650, N3969, N2620);
buf BUF1 (N10653, N10643);
nand NAND2 (N10654, N10649, N7993);
nand NAND2 (N10655, N10634, N5848);
and AND2 (N10656, N10648, N6075);
xor XOR2 (N10657, N10630, N7782);
not NOT1 (N10658, N10645);
or OR4 (N10659, N10658, N4766, N2136, N4605);
nand NAND4 (N10660, N10655, N9964, N1554, N9156);
buf BUF1 (N10661, N10659);
or OR3 (N10662, N10653, N7599, N4304);
xor XOR2 (N10663, N10654, N3058);
nand NAND2 (N10664, N10660, N9759);
nand NAND3 (N10665, N10661, N3141, N3943);
not NOT1 (N10666, N10664);
not NOT1 (N10667, N10651);
nor NOR4 (N10668, N10666, N7148, N9285, N455);
buf BUF1 (N10669, N10665);
nor NOR4 (N10670, N10656, N4072, N3727, N10667);
buf BUF1 (N10671, N4484);
xor XOR2 (N10672, N10670, N5975);
or OR3 (N10673, N10668, N5074, N8453);
nor NOR3 (N10674, N10673, N6940, N3804);
nor NOR3 (N10675, N10652, N7919, N16);
nor NOR4 (N10676, N10672, N4269, N4525, N9012);
buf BUF1 (N10677, N10631);
and AND3 (N10678, N10671, N3166, N9244);
nand NAND4 (N10679, N10657, N8072, N9406, N2508);
xor XOR2 (N10680, N10662, N6206);
buf BUF1 (N10681, N10678);
or OR4 (N10682, N10676, N8550, N9058, N8177);
nor NOR2 (N10683, N10674, N7719);
xor XOR2 (N10684, N10677, N3787);
not NOT1 (N10685, N10675);
not NOT1 (N10686, N10681);
xor XOR2 (N10687, N10686, N659);
xor XOR2 (N10688, N10684, N4125);
buf BUF1 (N10689, N10669);
or OR4 (N10690, N10689, N9017, N10025, N4171);
not NOT1 (N10691, N10663);
nor NOR3 (N10692, N10685, N7793, N8984);
buf BUF1 (N10693, N10636);
buf BUF1 (N10694, N10693);
not NOT1 (N10695, N10680);
buf BUF1 (N10696, N10690);
not NOT1 (N10697, N10688);
and AND2 (N10698, N10691, N2947);
xor XOR2 (N10699, N10683, N7907);
nand NAND3 (N10700, N10699, N75, N6298);
and AND3 (N10701, N10698, N3728, N10608);
nor NOR2 (N10702, N10679, N9569);
nand NAND4 (N10703, N10687, N4703, N2397, N2658);
buf BUF1 (N10704, N10692);
nor NOR4 (N10705, N10682, N1694, N8586, N3577);
or OR3 (N10706, N10702, N5846, N1641);
nand NAND4 (N10707, N10695, N7212, N503, N1633);
nor NOR3 (N10708, N10706, N2331, N10670);
or OR3 (N10709, N10697, N7648, N2004);
xor XOR2 (N10710, N10704, N8812);
nand NAND4 (N10711, N10710, N6254, N2421, N4258);
not NOT1 (N10712, N10701);
buf BUF1 (N10713, N10694);
xor XOR2 (N10714, N10709, N3086);
nand NAND3 (N10715, N10696, N7241, N10343);
and AND2 (N10716, N10714, N6303);
buf BUF1 (N10717, N10716);
buf BUF1 (N10718, N10713);
and AND2 (N10719, N10711, N5342);
xor XOR2 (N10720, N10708, N3478);
nor NOR2 (N10721, N10717, N1744);
and AND3 (N10722, N10703, N9556, N9208);
not NOT1 (N10723, N10722);
nand NAND3 (N10724, N10719, N895, N86);
and AND2 (N10725, N10718, N9359);
nor NOR2 (N10726, N10723, N4792);
or OR4 (N10727, N10720, N2947, N10660, N3369);
nand NAND4 (N10728, N10707, N592, N6547, N1768);
nor NOR2 (N10729, N10724, N9718);
nand NAND2 (N10730, N10725, N6053);
not NOT1 (N10731, N10728);
xor XOR2 (N10732, N10705, N2933);
buf BUF1 (N10733, N10729);
not NOT1 (N10734, N10733);
not NOT1 (N10735, N10727);
and AND2 (N10736, N10721, N190);
not NOT1 (N10737, N10700);
or OR3 (N10738, N10731, N3052, N8006);
xor XOR2 (N10739, N10734, N467);
buf BUF1 (N10740, N10730);
nand NAND4 (N10741, N10738, N10684, N450, N8211);
xor XOR2 (N10742, N10712, N117);
and AND4 (N10743, N10736, N9548, N10063, N4359);
not NOT1 (N10744, N10737);
or OR3 (N10745, N10740, N1507, N3870);
nor NOR4 (N10746, N10745, N10606, N9747, N9146);
nand NAND2 (N10747, N10726, N5927);
not NOT1 (N10748, N10747);
not NOT1 (N10749, N10741);
buf BUF1 (N10750, N10742);
buf BUF1 (N10751, N10743);
or OR3 (N10752, N10750, N7903, N5905);
nor NOR4 (N10753, N10739, N6261, N5354, N2113);
xor XOR2 (N10754, N10735, N7818);
not NOT1 (N10755, N10732);
and AND4 (N10756, N10752, N190, N5847, N8327);
nor NOR2 (N10757, N10753, N8098);
not NOT1 (N10758, N10748);
buf BUF1 (N10759, N10754);
or OR4 (N10760, N10751, N9082, N6164, N1958);
or OR3 (N10761, N10746, N2453, N10027);
or OR3 (N10762, N10749, N6968, N9096);
not NOT1 (N10763, N10758);
not NOT1 (N10764, N10761);
not NOT1 (N10765, N10760);
xor XOR2 (N10766, N10755, N177);
and AND4 (N10767, N10763, N7476, N7166, N1946);
or OR4 (N10768, N10744, N10742, N4793, N238);
buf BUF1 (N10769, N10757);
or OR3 (N10770, N10765, N9588, N3596);
not NOT1 (N10771, N10768);
nand NAND4 (N10772, N10769, N6386, N780, N9567);
nand NAND2 (N10773, N10766, N4897);
nor NOR3 (N10774, N10772, N9350, N9015);
and AND3 (N10775, N10770, N9480, N2440);
nor NOR2 (N10776, N10764, N2594);
buf BUF1 (N10777, N10756);
buf BUF1 (N10778, N10762);
nor NOR2 (N10779, N10715, N8459);
buf BUF1 (N10780, N10767);
xor XOR2 (N10781, N10773, N7297);
nand NAND4 (N10782, N10775, N1752, N1242, N308);
nand NAND3 (N10783, N10759, N9793, N9580);
xor XOR2 (N10784, N10778, N7730);
or OR4 (N10785, N10783, N452, N6711, N37);
xor XOR2 (N10786, N10774, N10412);
and AND3 (N10787, N10781, N5308, N126);
nor NOR2 (N10788, N10771, N10644);
and AND4 (N10789, N10784, N7765, N5206, N7406);
buf BUF1 (N10790, N10779);
and AND2 (N10791, N10777, N1770);
not NOT1 (N10792, N10787);
or OR4 (N10793, N10791, N9767, N1518, N9485);
buf BUF1 (N10794, N10786);
not NOT1 (N10795, N10785);
xor XOR2 (N10796, N10794, N6942);
nor NOR2 (N10797, N10776, N3666);
nor NOR4 (N10798, N10793, N5382, N3479, N5108);
xor XOR2 (N10799, N10798, N4575);
nor NOR2 (N10800, N10792, N2884);
or OR2 (N10801, N10799, N3455);
and AND3 (N10802, N10780, N7976, N8890);
xor XOR2 (N10803, N10801, N2856);
or OR2 (N10804, N10790, N7388);
buf BUF1 (N10805, N10795);
or OR3 (N10806, N10796, N5628, N5288);
buf BUF1 (N10807, N10800);
not NOT1 (N10808, N10797);
xor XOR2 (N10809, N10803, N1781);
xor XOR2 (N10810, N10806, N8899);
buf BUF1 (N10811, N10809);
buf BUF1 (N10812, N10789);
not NOT1 (N10813, N10807);
xor XOR2 (N10814, N10788, N592);
or OR4 (N10815, N10810, N10354, N4855, N1798);
buf BUF1 (N10816, N10802);
nor NOR2 (N10817, N10813, N3175);
nor NOR4 (N10818, N10805, N4585, N6750, N4489);
buf BUF1 (N10819, N10804);
xor XOR2 (N10820, N10812, N8402);
not NOT1 (N10821, N10782);
or OR2 (N10822, N10816, N706);
nor NOR3 (N10823, N10814, N5590, N9657);
nand NAND4 (N10824, N10819, N5521, N1782, N6843);
or OR2 (N10825, N10820, N4526);
or OR2 (N10826, N10818, N8407);
not NOT1 (N10827, N10815);
not NOT1 (N10828, N10808);
buf BUF1 (N10829, N10822);
not NOT1 (N10830, N10829);
buf BUF1 (N10831, N10817);
nand NAND4 (N10832, N10821, N2438, N4749, N9564);
buf BUF1 (N10833, N10830);
not NOT1 (N10834, N10827);
xor XOR2 (N10835, N10826, N3551);
xor XOR2 (N10836, N10824, N2408);
xor XOR2 (N10837, N10834, N4766);
buf BUF1 (N10838, N10823);
not NOT1 (N10839, N10828);
and AND3 (N10840, N10836, N4765, N4053);
buf BUF1 (N10841, N10831);
xor XOR2 (N10842, N10825, N10003);
nand NAND4 (N10843, N10840, N8864, N5521, N9039);
nand NAND3 (N10844, N10843, N2141, N9068);
xor XOR2 (N10845, N10842, N5332);
or OR3 (N10846, N10845, N2738, N9506);
xor XOR2 (N10847, N10837, N9327);
nor NOR3 (N10848, N10811, N10161, N72);
not NOT1 (N10849, N10839);
xor XOR2 (N10850, N10847, N2790);
or OR3 (N10851, N10844, N3298, N5506);
nand NAND3 (N10852, N10850, N4334, N2775);
and AND2 (N10853, N10838, N8539);
or OR2 (N10854, N10852, N10662);
and AND2 (N10855, N10846, N6142);
not NOT1 (N10856, N10833);
nand NAND2 (N10857, N10841, N9938);
and AND2 (N10858, N10854, N224);
buf BUF1 (N10859, N10835);
buf BUF1 (N10860, N10855);
not NOT1 (N10861, N10853);
or OR2 (N10862, N10856, N8939);
nor NOR4 (N10863, N10857, N2229, N4375, N4106);
and AND2 (N10864, N10849, N5807);
not NOT1 (N10865, N10861);
nand NAND4 (N10866, N10832, N8637, N7433, N2510);
not NOT1 (N10867, N10865);
xor XOR2 (N10868, N10866, N7573);
xor XOR2 (N10869, N10868, N10077);
buf BUF1 (N10870, N10848);
and AND2 (N10871, N10863, N4083);
or OR3 (N10872, N10851, N9297, N1468);
nand NAND4 (N10873, N10860, N1839, N6852, N6458);
and AND4 (N10874, N10873, N6460, N7780, N9676);
buf BUF1 (N10875, N10869);
not NOT1 (N10876, N10867);
nand NAND4 (N10877, N10859, N5617, N5952, N4441);
xor XOR2 (N10878, N10874, N8451);
nand NAND2 (N10879, N10876, N5282);
and AND3 (N10880, N10878, N1089, N9211);
xor XOR2 (N10881, N10879, N1766);
or OR2 (N10882, N10877, N4602);
xor XOR2 (N10883, N10881, N4870);
buf BUF1 (N10884, N10862);
or OR4 (N10885, N10880, N3373, N9419, N9175);
or OR2 (N10886, N10875, N3066);
nor NOR3 (N10887, N10870, N7854, N9777);
buf BUF1 (N10888, N10885);
nor NOR2 (N10889, N10871, N3856);
xor XOR2 (N10890, N10889, N9637);
nand NAND2 (N10891, N10864, N7409);
and AND4 (N10892, N10882, N368, N1567, N1904);
and AND2 (N10893, N10887, N486);
buf BUF1 (N10894, N10858);
not NOT1 (N10895, N10891);
or OR2 (N10896, N10893, N10879);
or OR3 (N10897, N10892, N5432, N5769);
nand NAND3 (N10898, N10895, N9728, N9225);
nor NOR3 (N10899, N10890, N10649, N2443);
or OR2 (N10900, N10883, N847);
nand NAND4 (N10901, N10897, N4869, N3798, N5022);
buf BUF1 (N10902, N10886);
and AND2 (N10903, N10901, N2912);
xor XOR2 (N10904, N10872, N2427);
buf BUF1 (N10905, N10894);
xor XOR2 (N10906, N10905, N5249);
and AND2 (N10907, N10904, N7354);
not NOT1 (N10908, N10896);
xor XOR2 (N10909, N10900, N5090);
nor NOR3 (N10910, N10888, N3867, N10020);
not NOT1 (N10911, N10902);
and AND4 (N10912, N10908, N6086, N4373, N1632);
or OR4 (N10913, N10903, N9060, N10525, N7625);
buf BUF1 (N10914, N10913);
nor NOR4 (N10915, N10910, N2935, N8400, N10305);
nor NOR3 (N10916, N10884, N3068, N2683);
xor XOR2 (N10917, N10915, N259);
buf BUF1 (N10918, N10912);
or OR2 (N10919, N10909, N5523);
and AND3 (N10920, N10899, N10366, N8444);
not NOT1 (N10921, N10919);
nand NAND2 (N10922, N10921, N8947);
buf BUF1 (N10923, N10911);
xor XOR2 (N10924, N10920, N7518);
nand NAND4 (N10925, N10907, N2109, N9696, N4633);
not NOT1 (N10926, N10923);
or OR4 (N10927, N10898, N4550, N9667, N4487);
or OR3 (N10928, N10925, N4946, N10886);
not NOT1 (N10929, N10918);
buf BUF1 (N10930, N10929);
nand NAND4 (N10931, N10906, N9001, N10879, N4075);
and AND3 (N10932, N10930, N3096, N7385);
buf BUF1 (N10933, N10917);
buf BUF1 (N10934, N10928);
and AND2 (N10935, N10926, N2958);
or OR3 (N10936, N10935, N297, N365);
xor XOR2 (N10937, N10934, N9942);
buf BUF1 (N10938, N10936);
xor XOR2 (N10939, N10922, N9394);
not NOT1 (N10940, N10938);
buf BUF1 (N10941, N10924);
and AND4 (N10942, N10932, N8502, N1485, N9520);
nand NAND3 (N10943, N10937, N3420, N6517);
xor XOR2 (N10944, N10940, N9686);
nand NAND4 (N10945, N10943, N6422, N10811, N1162);
not NOT1 (N10946, N10931);
buf BUF1 (N10947, N10942);
buf BUF1 (N10948, N10946);
buf BUF1 (N10949, N10914);
or OR3 (N10950, N10948, N2743, N8502);
not NOT1 (N10951, N10916);
buf BUF1 (N10952, N10939);
nor NOR2 (N10953, N10944, N1304);
buf BUF1 (N10954, N10933);
nor NOR2 (N10955, N10947, N1543);
nor NOR2 (N10956, N10927, N316);
buf BUF1 (N10957, N10956);
nand NAND4 (N10958, N10952, N5394, N4817, N10197);
not NOT1 (N10959, N10955);
nor NOR4 (N10960, N10959, N1202, N10054, N1436);
not NOT1 (N10961, N10953);
or OR2 (N10962, N10949, N1779);
nand NAND3 (N10963, N10945, N7164, N702);
and AND4 (N10964, N10954, N5059, N9845, N2129);
nor NOR3 (N10965, N10950, N4332, N6329);
xor XOR2 (N10966, N10964, N10432);
or OR2 (N10967, N10961, N2556);
not NOT1 (N10968, N10967);
not NOT1 (N10969, N10966);
nand NAND4 (N10970, N10951, N1252, N8148, N10451);
not NOT1 (N10971, N10941);
nor NOR2 (N10972, N10971, N3664);
buf BUF1 (N10973, N10960);
and AND3 (N10974, N10962, N8397, N8235);
nor NOR2 (N10975, N10973, N9547);
nand NAND4 (N10976, N10970, N6147, N632, N10227);
or OR4 (N10977, N10958, N2078, N8127, N514);
or OR3 (N10978, N10976, N9511, N5489);
nor NOR2 (N10979, N10957, N8855);
not NOT1 (N10980, N10972);
not NOT1 (N10981, N10968);
nor NOR2 (N10982, N10969, N1335);
nor NOR3 (N10983, N10978, N1822, N10695);
xor XOR2 (N10984, N10981, N10651);
xor XOR2 (N10985, N10975, N6434);
nor NOR3 (N10986, N10985, N7143, N7360);
or OR3 (N10987, N10986, N10523, N6494);
or OR3 (N10988, N10987, N1543, N3564);
nor NOR2 (N10989, N10979, N4372);
nand NAND3 (N10990, N10989, N288, N9053);
nand NAND2 (N10991, N10980, N3238);
xor XOR2 (N10992, N10965, N3643);
nand NAND3 (N10993, N10982, N2186, N5104);
xor XOR2 (N10994, N10992, N8298);
or OR2 (N10995, N10984, N159);
not NOT1 (N10996, N10988);
nand NAND4 (N10997, N10993, N10987, N2519, N9445);
or OR4 (N10998, N10977, N4043, N5717, N3039);
nor NOR2 (N10999, N10983, N6042);
xor XOR2 (N11000, N10999, N2812);
nor NOR3 (N11001, N10991, N7492, N3024);
not NOT1 (N11002, N10974);
xor XOR2 (N11003, N11000, N1900);
nand NAND4 (N11004, N10963, N1859, N8798, N7400);
or OR3 (N11005, N10994, N6556, N4309);
and AND2 (N11006, N10998, N9758);
and AND3 (N11007, N11006, N3120, N8921);
nor NOR3 (N11008, N11005, N8068, N1227);
nand NAND3 (N11009, N10995, N1053, N893);
or OR3 (N11010, N11002, N234, N10450);
buf BUF1 (N11011, N11004);
nor NOR3 (N11012, N11008, N5170, N9193);
or OR2 (N11013, N11007, N10513);
nand NAND2 (N11014, N11001, N5403);
or OR4 (N11015, N10997, N7058, N10090, N1925);
and AND3 (N11016, N11015, N5951, N4775);
nor NOR4 (N11017, N10996, N2418, N9928, N7914);
buf BUF1 (N11018, N11010);
nor NOR2 (N11019, N10990, N4951);
and AND2 (N11020, N11017, N6668);
nand NAND4 (N11021, N11014, N1680, N4147, N5179);
xor XOR2 (N11022, N11020, N2307);
buf BUF1 (N11023, N11013);
buf BUF1 (N11024, N11018);
not NOT1 (N11025, N11019);
or OR2 (N11026, N11021, N5799);
and AND4 (N11027, N11023, N700, N4074, N9967);
nor NOR4 (N11028, N11012, N2429, N5139, N2283);
and AND3 (N11029, N11009, N10353, N613);
or OR3 (N11030, N11011, N9862, N9314);
nor NOR3 (N11031, N11027, N6515, N6928);
not NOT1 (N11032, N11024);
xor XOR2 (N11033, N11003, N7595);
and AND3 (N11034, N11026, N2911, N39);
buf BUF1 (N11035, N11032);
not NOT1 (N11036, N11031);
and AND4 (N11037, N11022, N5215, N3802, N10244);
nand NAND3 (N11038, N11028, N10038, N10118);
buf BUF1 (N11039, N11030);
nand NAND2 (N11040, N11037, N9991);
not NOT1 (N11041, N11035);
nor NOR4 (N11042, N11040, N5423, N9183, N6235);
and AND4 (N11043, N11041, N2226, N7647, N9477);
nor NOR4 (N11044, N11034, N1922, N9289, N8273);
nand NAND3 (N11045, N11033, N652, N9320);
nor NOR2 (N11046, N11045, N8495);
nand NAND3 (N11047, N11025, N4850, N8137);
nor NOR2 (N11048, N11046, N8554);
and AND3 (N11049, N11042, N1449, N9969);
buf BUF1 (N11050, N11029);
nand NAND4 (N11051, N11050, N4063, N10209, N5579);
buf BUF1 (N11052, N11039);
buf BUF1 (N11053, N11043);
and AND2 (N11054, N11051, N2593);
or OR4 (N11055, N11038, N1583, N4560, N4686);
and AND4 (N11056, N11052, N7416, N8539, N3896);
not NOT1 (N11057, N11047);
xor XOR2 (N11058, N11048, N1400);
or OR3 (N11059, N11055, N8147, N1848);
or OR2 (N11060, N11036, N4100);
nand NAND4 (N11061, N11053, N3399, N4647, N8153);
buf BUF1 (N11062, N11054);
not NOT1 (N11063, N11057);
buf BUF1 (N11064, N11060);
and AND4 (N11065, N11059, N7143, N3346, N5493);
nor NOR2 (N11066, N11044, N10616);
or OR3 (N11067, N11062, N9648, N7015);
not NOT1 (N11068, N11067);
nand NAND4 (N11069, N11063, N10492, N943, N7241);
nor NOR3 (N11070, N11065, N1904, N1591);
and AND3 (N11071, N11069, N8176, N2011);
xor XOR2 (N11072, N11056, N1368);
nor NOR3 (N11073, N11068, N5023, N6589);
not NOT1 (N11074, N11066);
buf BUF1 (N11075, N11061);
nor NOR3 (N11076, N11049, N8389, N6192);
and AND3 (N11077, N11073, N6158, N9616);
xor XOR2 (N11078, N11072, N7643);
xor XOR2 (N11079, N11077, N7407);
and AND2 (N11080, N11075, N1642);
not NOT1 (N11081, N11076);
or OR4 (N11082, N11078, N7964, N2230, N11009);
nand NAND4 (N11083, N11074, N665, N10438, N3381);
nand NAND4 (N11084, N11080, N713, N6684, N7293);
buf BUF1 (N11085, N11070);
and AND4 (N11086, N11016, N8283, N5817, N1808);
nor NOR2 (N11087, N11083, N5776);
not NOT1 (N11088, N11058);
and AND2 (N11089, N11087, N8004);
and AND4 (N11090, N11082, N6596, N6169, N321);
nor NOR4 (N11091, N11081, N3329, N6920, N6831);
or OR3 (N11092, N11084, N6214, N5665);
or OR3 (N11093, N11092, N10762, N2006);
buf BUF1 (N11094, N11091);
nand NAND3 (N11095, N11071, N10200, N356);
nand NAND3 (N11096, N11094, N1433, N3603);
or OR4 (N11097, N11088, N5911, N10251, N10048);
not NOT1 (N11098, N11085);
nand NAND3 (N11099, N11095, N6682, N1666);
nor NOR3 (N11100, N11086, N10772, N105);
not NOT1 (N11101, N11089);
or OR2 (N11102, N11079, N430);
xor XOR2 (N11103, N11090, N4409);
and AND2 (N11104, N11102, N217);
xor XOR2 (N11105, N11093, N7304);
nor NOR2 (N11106, N11104, N7223);
nand NAND2 (N11107, N11098, N5619);
xor XOR2 (N11108, N11101, N5641);
buf BUF1 (N11109, N11107);
not NOT1 (N11110, N11106);
nand NAND3 (N11111, N11110, N3216, N8640);
not NOT1 (N11112, N11099);
xor XOR2 (N11113, N11100, N10193);
nand NAND4 (N11114, N11105, N5653, N6720, N9839);
not NOT1 (N11115, N11112);
not NOT1 (N11116, N11114);
xor XOR2 (N11117, N11116, N4887);
not NOT1 (N11118, N11096);
buf BUF1 (N11119, N11064);
not NOT1 (N11120, N11097);
and AND4 (N11121, N11113, N688, N1601, N3614);
not NOT1 (N11122, N11118);
nor NOR4 (N11123, N11122, N4303, N1869, N6762);
and AND2 (N11124, N11108, N6990);
not NOT1 (N11125, N11115);
xor XOR2 (N11126, N11124, N8354);
and AND4 (N11127, N11125, N4535, N2107, N7360);
not NOT1 (N11128, N11111);
and AND3 (N11129, N11128, N9188, N897);
or OR4 (N11130, N11109, N2592, N4662, N10503);
buf BUF1 (N11131, N11103);
buf BUF1 (N11132, N11126);
not NOT1 (N11133, N11129);
nand NAND3 (N11134, N11121, N10236, N7974);
nand NAND2 (N11135, N11119, N9153);
xor XOR2 (N11136, N11131, N7540);
nor NOR4 (N11137, N11135, N453, N678, N1580);
nand NAND3 (N11138, N11132, N4428, N3226);
nor NOR4 (N11139, N11138, N9258, N6149, N2480);
nor NOR2 (N11140, N11127, N10372);
buf BUF1 (N11141, N11133);
not NOT1 (N11142, N11117);
and AND4 (N11143, N11139, N890, N198, N8280);
not NOT1 (N11144, N11136);
and AND2 (N11145, N11123, N5846);
xor XOR2 (N11146, N11134, N10796);
buf BUF1 (N11147, N11142);
and AND2 (N11148, N11146, N299);
not NOT1 (N11149, N11137);
xor XOR2 (N11150, N11120, N1728);
nor NOR3 (N11151, N11147, N758, N9336);
not NOT1 (N11152, N11141);
buf BUF1 (N11153, N11130);
and AND4 (N11154, N11149, N6206, N1241, N4249);
and AND4 (N11155, N11144, N1157, N9138, N3283);
not NOT1 (N11156, N11154);
nor NOR4 (N11157, N11155, N1132, N6879, N9431);
not NOT1 (N11158, N11148);
nor NOR3 (N11159, N11153, N5920, N5369);
or OR2 (N11160, N11157, N8458);
and AND2 (N11161, N11145, N3984);
xor XOR2 (N11162, N11158, N6288);
and AND2 (N11163, N11140, N8372);
not NOT1 (N11164, N11159);
nor NOR4 (N11165, N11160, N289, N5155, N1976);
buf BUF1 (N11166, N11164);
buf BUF1 (N11167, N11156);
nor NOR2 (N11168, N11151, N2601);
nand NAND4 (N11169, N11166, N9680, N9208, N10056);
not NOT1 (N11170, N11162);
and AND2 (N11171, N11152, N1457);
or OR4 (N11172, N11161, N9111, N312, N5938);
and AND3 (N11173, N11169, N8975, N6244);
nor NOR2 (N11174, N11163, N6479);
nor NOR3 (N11175, N11173, N10031, N4950);
and AND4 (N11176, N11167, N640, N8260, N7997);
xor XOR2 (N11177, N11165, N5039);
and AND4 (N11178, N11170, N1235, N10056, N1998);
not NOT1 (N11179, N11177);
not NOT1 (N11180, N11172);
and AND4 (N11181, N11176, N7123, N6595, N6012);
nand NAND3 (N11182, N11181, N4855, N6225);
or OR2 (N11183, N11182, N7462);
nor NOR3 (N11184, N11175, N841, N7823);
xor XOR2 (N11185, N11178, N4916);
buf BUF1 (N11186, N11150);
and AND2 (N11187, N11186, N6239);
nor NOR4 (N11188, N11180, N9223, N3537, N6774);
nor NOR4 (N11189, N11183, N345, N7060, N8408);
or OR2 (N11190, N11189, N5724);
and AND4 (N11191, N11185, N4839, N2429, N4886);
not NOT1 (N11192, N11143);
or OR4 (N11193, N11184, N767, N9152, N2313);
buf BUF1 (N11194, N11190);
nor NOR3 (N11195, N11194, N6170, N10254);
nor NOR4 (N11196, N11192, N11067, N7508, N10116);
or OR4 (N11197, N11193, N4752, N4931, N55);
nand NAND3 (N11198, N11195, N6597, N3371);
or OR4 (N11199, N11171, N4521, N8496, N3422);
nor NOR2 (N11200, N11198, N10025);
nor NOR2 (N11201, N11187, N9119);
buf BUF1 (N11202, N11197);
xor XOR2 (N11203, N11200, N9587);
nor NOR3 (N11204, N11188, N1021, N9075);
or OR2 (N11205, N11174, N216);
nand NAND3 (N11206, N11202, N7850, N2058);
xor XOR2 (N11207, N11168, N5214);
or OR3 (N11208, N11196, N8571, N5294);
buf BUF1 (N11209, N11201);
and AND3 (N11210, N11208, N9534, N10020);
nor NOR4 (N11211, N11205, N5393, N1903, N4109);
buf BUF1 (N11212, N11207);
and AND4 (N11213, N11211, N3613, N2100, N4074);
and AND4 (N11214, N11212, N3697, N5947, N4129);
not NOT1 (N11215, N11210);
not NOT1 (N11216, N11203);
xor XOR2 (N11217, N11199, N11010);
xor XOR2 (N11218, N11206, N3544);
buf BUF1 (N11219, N11218);
not NOT1 (N11220, N11216);
or OR2 (N11221, N11179, N7142);
buf BUF1 (N11222, N11215);
nor NOR4 (N11223, N11220, N5145, N7666, N8028);
nor NOR4 (N11224, N11214, N6955, N9725, N10939);
or OR3 (N11225, N11224, N9127, N9689);
nor NOR3 (N11226, N11209, N10729, N5990);
buf BUF1 (N11227, N11217);
not NOT1 (N11228, N11191);
not NOT1 (N11229, N11219);
and AND3 (N11230, N11225, N2231, N9775);
nor NOR4 (N11231, N11229, N1732, N4128, N6473);
nand NAND4 (N11232, N11213, N2296, N723, N5001);
nor NOR2 (N11233, N11232, N7394);
not NOT1 (N11234, N11223);
or OR3 (N11235, N11221, N1998, N5519);
and AND2 (N11236, N11235, N6326);
xor XOR2 (N11237, N11236, N5816);
buf BUF1 (N11238, N11227);
xor XOR2 (N11239, N11228, N10958);
buf BUF1 (N11240, N11226);
xor XOR2 (N11241, N11230, N3621);
buf BUF1 (N11242, N11231);
nor NOR4 (N11243, N11238, N3408, N3661, N3834);
buf BUF1 (N11244, N11241);
and AND4 (N11245, N11222, N9101, N6956, N6);
nor NOR3 (N11246, N11240, N2185, N8484);
nand NAND4 (N11247, N11246, N260, N3195, N8336);
nor NOR2 (N11248, N11239, N8080);
nor NOR4 (N11249, N11244, N493, N9648, N41);
and AND3 (N11250, N11242, N10766, N7258);
not NOT1 (N11251, N11247);
buf BUF1 (N11252, N11243);
and AND4 (N11253, N11245, N1365, N2618, N592);
nor NOR3 (N11254, N11253, N2619, N8575);
buf BUF1 (N11255, N11204);
not NOT1 (N11256, N11237);
nand NAND4 (N11257, N11252, N8679, N10669, N3742);
nor NOR4 (N11258, N11254, N6157, N2758, N1835);
buf BUF1 (N11259, N11255);
not NOT1 (N11260, N11256);
xor XOR2 (N11261, N11250, N4101);
or OR3 (N11262, N11248, N1700, N11229);
buf BUF1 (N11263, N11261);
xor XOR2 (N11264, N11260, N8097);
buf BUF1 (N11265, N11259);
or OR3 (N11266, N11264, N9427, N8238);
xor XOR2 (N11267, N11265, N7782);
or OR2 (N11268, N11263, N204);
not NOT1 (N11269, N11262);
buf BUF1 (N11270, N11249);
not NOT1 (N11271, N11234);
nand NAND2 (N11272, N11233, N10549);
buf BUF1 (N11273, N11272);
and AND4 (N11274, N11271, N9011, N3247, N4821);
nand NAND4 (N11275, N11274, N4546, N196, N10922);
and AND3 (N11276, N11266, N3943, N6086);
buf BUF1 (N11277, N11257);
not NOT1 (N11278, N11276);
not NOT1 (N11279, N11267);
or OR3 (N11280, N11279, N9807, N3600);
or OR3 (N11281, N11273, N3779, N4530);
nor NOR2 (N11282, N11251, N6283);
or OR3 (N11283, N11270, N5451, N5180);
not NOT1 (N11284, N11277);
buf BUF1 (N11285, N11268);
and AND3 (N11286, N11285, N533, N390);
or OR2 (N11287, N11281, N4847);
or OR2 (N11288, N11284, N6195);
nor NOR4 (N11289, N11286, N8548, N4056, N9484);
or OR2 (N11290, N11280, N3511);
nand NAND3 (N11291, N11289, N7127, N5347);
nor NOR4 (N11292, N11288, N2197, N10231, N5053);
buf BUF1 (N11293, N11291);
and AND4 (N11294, N11275, N5368, N6364, N502);
nand NAND4 (N11295, N11294, N7022, N1924, N10450);
xor XOR2 (N11296, N11292, N10311);
xor XOR2 (N11297, N11287, N3077);
nand NAND2 (N11298, N11295, N787);
not NOT1 (N11299, N11278);
xor XOR2 (N11300, N11283, N653);
nand NAND3 (N11301, N11293, N9630, N10882);
nor NOR4 (N11302, N11301, N2238, N742, N647);
nand NAND3 (N11303, N11299, N10208, N891);
nand NAND3 (N11304, N11298, N6966, N2862);
buf BUF1 (N11305, N11304);
xor XOR2 (N11306, N11302, N222);
and AND4 (N11307, N11269, N11214, N1678, N9532);
and AND4 (N11308, N11307, N1473, N6433, N1076);
not NOT1 (N11309, N11303);
and AND3 (N11310, N11309, N6226, N8917);
xor XOR2 (N11311, N11282, N6237);
not NOT1 (N11312, N11297);
and AND3 (N11313, N11300, N9276, N2686);
nor NOR3 (N11314, N11306, N3871, N10113);
and AND2 (N11315, N11296, N7552);
not NOT1 (N11316, N11315);
nor NOR3 (N11317, N11316, N3735, N1772);
xor XOR2 (N11318, N11313, N7525);
and AND3 (N11319, N11305, N10555, N724);
buf BUF1 (N11320, N11310);
or OR2 (N11321, N11311, N3651);
not NOT1 (N11322, N11320);
buf BUF1 (N11323, N11312);
buf BUF1 (N11324, N11319);
buf BUF1 (N11325, N11317);
and AND4 (N11326, N11325, N2624, N5272, N2773);
buf BUF1 (N11327, N11322);
not NOT1 (N11328, N11324);
nor NOR3 (N11329, N11314, N6258, N8457);
nor NOR3 (N11330, N11321, N6131, N254);
not NOT1 (N11331, N11328);
or OR2 (N11332, N11327, N5397);
nor NOR2 (N11333, N11326, N6382);
nor NOR4 (N11334, N11308, N2732, N9117, N4374);
not NOT1 (N11335, N11323);
nor NOR3 (N11336, N11331, N4097, N2586);
buf BUF1 (N11337, N11290);
not NOT1 (N11338, N11337);
nor NOR4 (N11339, N11258, N3558, N2409, N7094);
nor NOR2 (N11340, N11329, N8793);
buf BUF1 (N11341, N11335);
xor XOR2 (N11342, N11333, N7530);
nor NOR2 (N11343, N11318, N7242);
not NOT1 (N11344, N11339);
nor NOR4 (N11345, N11338, N6935, N6689, N3308);
or OR4 (N11346, N11344, N434, N7249, N4043);
or OR3 (N11347, N11340, N7861, N7389);
xor XOR2 (N11348, N11330, N4009);
or OR4 (N11349, N11332, N4535, N2798, N10977);
nand NAND4 (N11350, N11341, N10796, N1614, N4155);
or OR4 (N11351, N11342, N6923, N2089, N135);
buf BUF1 (N11352, N11350);
nor NOR4 (N11353, N11346, N1798, N4674, N10161);
or OR4 (N11354, N11348, N4586, N10032, N2273);
and AND3 (N11355, N11334, N6961, N5128);
nor NOR2 (N11356, N11347, N485);
xor XOR2 (N11357, N11345, N5305);
and AND2 (N11358, N11349, N2030);
buf BUF1 (N11359, N11358);
xor XOR2 (N11360, N11359, N10407);
buf BUF1 (N11361, N11360);
xor XOR2 (N11362, N11351, N9138);
or OR4 (N11363, N11354, N8597, N7395, N11114);
nor NOR4 (N11364, N11352, N4951, N10608, N7332);
or OR4 (N11365, N11355, N2743, N5519, N8814);
or OR3 (N11366, N11336, N6595, N3590);
nand NAND3 (N11367, N11343, N8859, N3325);
not NOT1 (N11368, N11356);
nand NAND3 (N11369, N11361, N5010, N9076);
nor NOR4 (N11370, N11362, N1260, N8198, N895);
or OR4 (N11371, N11365, N385, N2799, N5121);
nor NOR3 (N11372, N11370, N4907, N2219);
not NOT1 (N11373, N11371);
nand NAND3 (N11374, N11372, N4144, N3738);
buf BUF1 (N11375, N11367);
and AND3 (N11376, N11369, N1110, N3742);
buf BUF1 (N11377, N11375);
nand NAND3 (N11378, N11366, N4678, N11124);
or OR2 (N11379, N11376, N6826);
nand NAND3 (N11380, N11377, N7825, N7622);
xor XOR2 (N11381, N11373, N4412);
xor XOR2 (N11382, N11380, N8459);
or OR4 (N11383, N11353, N1396, N7536, N4385);
nor NOR2 (N11384, N11381, N9486);
nand NAND3 (N11385, N11357, N10091, N9892);
not NOT1 (N11386, N11378);
or OR4 (N11387, N11364, N9756, N4725, N734);
buf BUF1 (N11388, N11384);
or OR3 (N11389, N11383, N3825, N5967);
nand NAND2 (N11390, N11363, N7282);
xor XOR2 (N11391, N11389, N2732);
nor NOR3 (N11392, N11387, N8885, N5265);
xor XOR2 (N11393, N11368, N2623);
and AND3 (N11394, N11390, N948, N842);
or OR4 (N11395, N11391, N10786, N1669, N5819);
buf BUF1 (N11396, N11394);
buf BUF1 (N11397, N11393);
and AND4 (N11398, N11379, N1645, N9999, N3208);
or OR4 (N11399, N11398, N3540, N7175, N8647);
nor NOR4 (N11400, N11397, N1846, N8090, N5165);
nor NOR4 (N11401, N11382, N3478, N6876, N3238);
nand NAND3 (N11402, N11401, N9846, N2474);
and AND3 (N11403, N11400, N7556, N60);
and AND2 (N11404, N11399, N2593);
buf BUF1 (N11405, N11396);
xor XOR2 (N11406, N11385, N6135);
or OR2 (N11407, N11405, N6112);
xor XOR2 (N11408, N11402, N8625);
nand NAND4 (N11409, N11374, N10228, N8127, N1038);
nor NOR4 (N11410, N11395, N5890, N7894, N9175);
nand NAND2 (N11411, N11407, N1061);
buf BUF1 (N11412, N11406);
and AND3 (N11413, N11410, N6928, N7664);
buf BUF1 (N11414, N11411);
nand NAND3 (N11415, N11413, N3787, N5184);
and AND4 (N11416, N11412, N8238, N5980, N2759);
and AND2 (N11417, N11386, N3311);
or OR3 (N11418, N11416, N7241, N10479);
xor XOR2 (N11419, N11408, N7222);
not NOT1 (N11420, N11403);
buf BUF1 (N11421, N11419);
not NOT1 (N11422, N11388);
buf BUF1 (N11423, N11417);
and AND2 (N11424, N11420, N394);
or OR4 (N11425, N11418, N2104, N5118, N5914);
buf BUF1 (N11426, N11423);
or OR4 (N11427, N11426, N5957, N555, N8151);
buf BUF1 (N11428, N11415);
buf BUF1 (N11429, N11414);
or OR2 (N11430, N11425, N1774);
xor XOR2 (N11431, N11428, N9540);
nand NAND4 (N11432, N11404, N6696, N1079, N516);
nor NOR3 (N11433, N11431, N8302, N4645);
or OR3 (N11434, N11409, N5038, N3273);
not NOT1 (N11435, N11392);
nand NAND2 (N11436, N11430, N2333);
not NOT1 (N11437, N11432);
and AND4 (N11438, N11434, N263, N9966, N7110);
xor XOR2 (N11439, N11421, N4877);
nor NOR3 (N11440, N11429, N2842, N6621);
nand NAND4 (N11441, N11422, N9037, N4337, N4884);
and AND4 (N11442, N11440, N1767, N2657, N8062);
nand NAND4 (N11443, N11427, N2124, N6581, N7636);
nand NAND3 (N11444, N11435, N9875, N7122);
nor NOR2 (N11445, N11444, N8319);
nand NAND3 (N11446, N11443, N8846, N1598);
or OR2 (N11447, N11436, N1816);
xor XOR2 (N11448, N11424, N6001);
nand NAND2 (N11449, N11441, N8880);
not NOT1 (N11450, N11446);
xor XOR2 (N11451, N11442, N9934);
or OR4 (N11452, N11439, N8223, N699, N7310);
and AND3 (N11453, N11451, N9308, N6143);
not NOT1 (N11454, N11433);
or OR3 (N11455, N11449, N6127, N4887);
buf BUF1 (N11456, N11454);
xor XOR2 (N11457, N11448, N330);
or OR2 (N11458, N11437, N2572);
buf BUF1 (N11459, N11452);
nor NOR3 (N11460, N11459, N6771, N4766);
or OR4 (N11461, N11456, N10549, N7396, N5373);
and AND2 (N11462, N11458, N2618);
nor NOR2 (N11463, N11450, N7448);
and AND2 (N11464, N11463, N4651);
not NOT1 (N11465, N11464);
not NOT1 (N11466, N11461);
buf BUF1 (N11467, N11466);
or OR3 (N11468, N11465, N209, N6075);
or OR3 (N11469, N11445, N8407, N6654);
nor NOR4 (N11470, N11453, N8422, N4730, N1234);
buf BUF1 (N11471, N11469);
or OR2 (N11472, N11467, N5865);
and AND3 (N11473, N11468, N5990, N2262);
nor NOR4 (N11474, N11455, N6534, N3073, N7414);
xor XOR2 (N11475, N11474, N7125);
nor NOR4 (N11476, N11462, N107, N9240, N1930);
buf BUF1 (N11477, N11447);
nor NOR4 (N11478, N11475, N7579, N1609, N3002);
buf BUF1 (N11479, N11476);
or OR4 (N11480, N11473, N1803, N11038, N2660);
buf BUF1 (N11481, N11438);
buf BUF1 (N11482, N11472);
or OR3 (N11483, N11460, N10618, N4713);
xor XOR2 (N11484, N11482, N8175);
or OR4 (N11485, N11481, N10929, N10739, N5849);
xor XOR2 (N11486, N11479, N1833);
buf BUF1 (N11487, N11470);
and AND2 (N11488, N11485, N8478);
xor XOR2 (N11489, N11478, N2391);
or OR3 (N11490, N11486, N10695, N6802);
or OR3 (N11491, N11490, N5230, N11063);
xor XOR2 (N11492, N11477, N30);
buf BUF1 (N11493, N11484);
nor NOR3 (N11494, N11483, N9784, N7737);
not NOT1 (N11495, N11494);
xor XOR2 (N11496, N11495, N1837);
not NOT1 (N11497, N11496);
not NOT1 (N11498, N11480);
or OR2 (N11499, N11493, N9646);
nor NOR2 (N11500, N11499, N7064);
buf BUF1 (N11501, N11457);
nor NOR3 (N11502, N11489, N3834, N9744);
or OR4 (N11503, N11491, N2703, N4743, N6755);
and AND2 (N11504, N11492, N4379);
or OR4 (N11505, N11497, N8653, N4002, N6895);
xor XOR2 (N11506, N11504, N3163);
and AND4 (N11507, N11502, N310, N9092, N1352);
not NOT1 (N11508, N11506);
nor NOR3 (N11509, N11500, N10805, N4943);
buf BUF1 (N11510, N11507);
and AND2 (N11511, N11505, N10493);
or OR2 (N11512, N11487, N1168);
buf BUF1 (N11513, N11511);
nand NAND2 (N11514, N11488, N1805);
or OR2 (N11515, N11509, N407);
nand NAND3 (N11516, N11501, N8724, N10298);
buf BUF1 (N11517, N11471);
xor XOR2 (N11518, N11516, N5598);
nor NOR2 (N11519, N11515, N8944);
not NOT1 (N11520, N11498);
and AND2 (N11521, N11514, N9991);
buf BUF1 (N11522, N11518);
not NOT1 (N11523, N11522);
nor NOR2 (N11524, N11521, N718);
not NOT1 (N11525, N11508);
xor XOR2 (N11526, N11523, N1710);
nand NAND3 (N11527, N11519, N542, N8156);
nor NOR2 (N11528, N11525, N6272);
buf BUF1 (N11529, N11512);
nand NAND3 (N11530, N11510, N5773, N11064);
buf BUF1 (N11531, N11529);
buf BUF1 (N11532, N11513);
or OR4 (N11533, N11520, N2363, N92, N9994);
nand NAND4 (N11534, N11524, N6733, N4656, N9728);
and AND4 (N11535, N11532, N1941, N4892, N1445);
and AND4 (N11536, N11526, N8452, N8008, N5350);
xor XOR2 (N11537, N11535, N1048);
or OR4 (N11538, N11527, N11136, N699, N4211);
not NOT1 (N11539, N11538);
nor NOR3 (N11540, N11536, N3042, N10757);
and AND4 (N11541, N11517, N3479, N10450, N6466);
xor XOR2 (N11542, N11540, N10563);
or OR3 (N11543, N11530, N229, N10665);
buf BUF1 (N11544, N11503);
or OR2 (N11545, N11543, N3395);
or OR3 (N11546, N11533, N7441, N4324);
buf BUF1 (N11547, N11534);
nand NAND3 (N11548, N11546, N9962, N105);
or OR2 (N11549, N11548, N7288);
and AND2 (N11550, N11528, N752);
nor NOR2 (N11551, N11544, N9016);
or OR3 (N11552, N11549, N3875, N9157);
nand NAND2 (N11553, N11545, N9057);
nor NOR2 (N11554, N11550, N9069);
or OR3 (N11555, N11541, N6715, N11102);
or OR4 (N11556, N11539, N4223, N8801, N5695);
nor NOR4 (N11557, N11552, N9580, N10607, N4940);
not NOT1 (N11558, N11542);
buf BUF1 (N11559, N11554);
not NOT1 (N11560, N11553);
nand NAND3 (N11561, N11558, N9653, N5193);
not NOT1 (N11562, N11537);
nor NOR2 (N11563, N11531, N4018);
buf BUF1 (N11564, N11547);
and AND3 (N11565, N11562, N3930, N3782);
and AND4 (N11566, N11555, N8705, N401, N6854);
buf BUF1 (N11567, N11556);
buf BUF1 (N11568, N11551);
buf BUF1 (N11569, N11563);
xor XOR2 (N11570, N11560, N5253);
xor XOR2 (N11571, N11566, N155);
buf BUF1 (N11572, N11570);
buf BUF1 (N11573, N11571);
not NOT1 (N11574, N11559);
not NOT1 (N11575, N11567);
and AND3 (N11576, N11569, N1421, N3792);
buf BUF1 (N11577, N11568);
xor XOR2 (N11578, N11561, N10026);
or OR2 (N11579, N11577, N5343);
xor XOR2 (N11580, N11564, N6729);
not NOT1 (N11581, N11565);
buf BUF1 (N11582, N11576);
or OR3 (N11583, N11580, N495, N1199);
not NOT1 (N11584, N11572);
xor XOR2 (N11585, N11557, N7584);
or OR4 (N11586, N11578, N4562, N348, N7508);
nor NOR2 (N11587, N11573, N10683);
not NOT1 (N11588, N11585);
nand NAND2 (N11589, N11574, N9445);
and AND2 (N11590, N11588, N6061);
nor NOR3 (N11591, N11579, N1662, N9912);
buf BUF1 (N11592, N11589);
buf BUF1 (N11593, N11586);
nand NAND3 (N11594, N11587, N6268, N11518);
nor NOR4 (N11595, N11583, N9414, N9281, N1487);
nand NAND3 (N11596, N11582, N3830, N8238);
and AND2 (N11597, N11595, N7111);
nand NAND3 (N11598, N11575, N2697, N6136);
not NOT1 (N11599, N11590);
buf BUF1 (N11600, N11581);
not NOT1 (N11601, N11596);
not NOT1 (N11602, N11592);
xor XOR2 (N11603, N11593, N10239);
nand NAND4 (N11604, N11584, N10807, N5835, N9154);
buf BUF1 (N11605, N11601);
nand NAND2 (N11606, N11598, N6327);
or OR4 (N11607, N11602, N2027, N5798, N8913);
and AND3 (N11608, N11605, N8556, N730);
nand NAND4 (N11609, N11600, N4545, N2281, N690);
or OR2 (N11610, N11608, N10284);
and AND4 (N11611, N11607, N4414, N9484, N9462);
nor NOR3 (N11612, N11603, N9377, N8835);
or OR2 (N11613, N11591, N5322);
or OR4 (N11614, N11610, N9740, N760, N8141);
xor XOR2 (N11615, N11609, N10043);
nand NAND3 (N11616, N11594, N9192, N11181);
and AND2 (N11617, N11604, N8178);
and AND4 (N11618, N11599, N2977, N2271, N4645);
xor XOR2 (N11619, N11613, N1577);
xor XOR2 (N11620, N11597, N4721);
or OR4 (N11621, N11614, N1460, N8453, N3844);
not NOT1 (N11622, N11615);
and AND3 (N11623, N11621, N9372, N9007);
and AND4 (N11624, N11622, N2750, N3807, N6365);
not NOT1 (N11625, N11618);
and AND3 (N11626, N11620, N4939, N731);
or OR3 (N11627, N11606, N1406, N4558);
buf BUF1 (N11628, N11619);
or OR4 (N11629, N11616, N1395, N5996, N312);
nor NOR3 (N11630, N11625, N9793, N11463);
xor XOR2 (N11631, N11626, N544);
and AND3 (N11632, N11611, N6900, N759);
or OR2 (N11633, N11629, N2350);
nand NAND2 (N11634, N11631, N1107);
not NOT1 (N11635, N11634);
buf BUF1 (N11636, N11628);
and AND3 (N11637, N11630, N1653, N5607);
nor NOR2 (N11638, N11623, N959);
and AND2 (N11639, N11635, N9468);
not NOT1 (N11640, N11624);
or OR2 (N11641, N11636, N7587);
buf BUF1 (N11642, N11633);
buf BUF1 (N11643, N11637);
xor XOR2 (N11644, N11632, N11112);
or OR2 (N11645, N11644, N6783);
xor XOR2 (N11646, N11627, N795);
buf BUF1 (N11647, N11638);
and AND3 (N11648, N11639, N11112, N247);
nand NAND3 (N11649, N11641, N7248, N2386);
or OR3 (N11650, N11643, N6393, N8258);
not NOT1 (N11651, N11612);
nand NAND4 (N11652, N11650, N2146, N6247, N8205);
xor XOR2 (N11653, N11642, N11331);
and AND4 (N11654, N11647, N4421, N7284, N7775);
not NOT1 (N11655, N11649);
xor XOR2 (N11656, N11648, N3398);
nor NOR4 (N11657, N11651, N11585, N4163, N5104);
not NOT1 (N11658, N11654);
nand NAND3 (N11659, N11655, N3089, N7635);
not NOT1 (N11660, N11653);
nor NOR2 (N11661, N11659, N8330);
nor NOR2 (N11662, N11658, N7913);
xor XOR2 (N11663, N11646, N1937);
not NOT1 (N11664, N11660);
nand NAND2 (N11665, N11640, N2857);
or OR3 (N11666, N11617, N11308, N2699);
nor NOR3 (N11667, N11656, N4398, N9893);
not NOT1 (N11668, N11666);
nor NOR2 (N11669, N11657, N8452);
nand NAND2 (N11670, N11667, N4581);
or OR4 (N11671, N11661, N9275, N6366, N10208);
and AND2 (N11672, N11669, N297);
not NOT1 (N11673, N11662);
or OR2 (N11674, N11663, N615);
nor NOR2 (N11675, N11665, N1);
not NOT1 (N11676, N11673);
nor NOR4 (N11677, N11664, N7413, N3468, N277);
or OR3 (N11678, N11676, N4449, N4680);
or OR2 (N11679, N11645, N10309);
and AND4 (N11680, N11679, N7323, N4222, N4217);
or OR3 (N11681, N11675, N7400, N11182);
and AND2 (N11682, N11671, N6209);
not NOT1 (N11683, N11668);
nor NOR3 (N11684, N11680, N8151, N200);
nand NAND3 (N11685, N11678, N6942, N5411);
nand NAND3 (N11686, N11672, N6536, N2800);
xor XOR2 (N11687, N11652, N4088);
xor XOR2 (N11688, N11687, N6385);
not NOT1 (N11689, N11686);
nand NAND3 (N11690, N11684, N4223, N7277);
and AND3 (N11691, N11670, N10765, N3435);
buf BUF1 (N11692, N11691);
or OR2 (N11693, N11692, N6010);
xor XOR2 (N11694, N11683, N6210);
xor XOR2 (N11695, N11682, N8205);
not NOT1 (N11696, N11690);
or OR4 (N11697, N11674, N5002, N10284, N11448);
xor XOR2 (N11698, N11688, N1419);
xor XOR2 (N11699, N11693, N7982);
xor XOR2 (N11700, N11695, N10055);
nor NOR3 (N11701, N11685, N10098, N11229);
or OR2 (N11702, N11700, N4093);
and AND2 (N11703, N11694, N3934);
buf BUF1 (N11704, N11703);
buf BUF1 (N11705, N11681);
nand NAND2 (N11706, N11704, N11162);
and AND3 (N11707, N11677, N1471, N8468);
nand NAND4 (N11708, N11698, N473, N10747, N6282);
xor XOR2 (N11709, N11705, N2519);
buf BUF1 (N11710, N11689);
xor XOR2 (N11711, N11709, N6806);
not NOT1 (N11712, N11699);
and AND3 (N11713, N11707, N5880, N3960);
not NOT1 (N11714, N11712);
xor XOR2 (N11715, N11708, N3686);
and AND4 (N11716, N11702, N8051, N11376, N9841);
buf BUF1 (N11717, N11716);
buf BUF1 (N11718, N11696);
xor XOR2 (N11719, N11715, N3717);
nand NAND4 (N11720, N11697, N9309, N3557, N4839);
xor XOR2 (N11721, N11717, N11252);
buf BUF1 (N11722, N11718);
and AND4 (N11723, N11710, N6984, N2405, N4050);
not NOT1 (N11724, N11706);
nor NOR4 (N11725, N11711, N4781, N3179, N8951);
and AND4 (N11726, N11723, N6538, N7289, N7116);
nand NAND2 (N11727, N11725, N1731);
nor NOR2 (N11728, N11713, N5597);
not NOT1 (N11729, N11719);
or OR2 (N11730, N11722, N11316);
buf BUF1 (N11731, N11720);
buf BUF1 (N11732, N11728);
and AND2 (N11733, N11727, N10299);
not NOT1 (N11734, N11714);
nor NOR2 (N11735, N11733, N9667);
xor XOR2 (N11736, N11735, N5178);
xor XOR2 (N11737, N11731, N5133);
buf BUF1 (N11738, N11729);
buf BUF1 (N11739, N11738);
or OR4 (N11740, N11721, N4428, N7808, N1532);
nor NOR2 (N11741, N11701, N7615);
and AND4 (N11742, N11730, N5655, N364, N8501);
xor XOR2 (N11743, N11726, N9913);
not NOT1 (N11744, N11734);
not NOT1 (N11745, N11744);
nand NAND2 (N11746, N11742, N10750);
buf BUF1 (N11747, N11746);
nor NOR4 (N11748, N11747, N3959, N4033, N5641);
nor NOR3 (N11749, N11724, N9408, N1518);
not NOT1 (N11750, N11736);
and AND4 (N11751, N11745, N6534, N5114, N6637);
nor NOR2 (N11752, N11743, N5156);
buf BUF1 (N11753, N11749);
and AND3 (N11754, N11750, N588, N11689);
buf BUF1 (N11755, N11753);
nor NOR4 (N11756, N11740, N9441, N10163, N6082);
buf BUF1 (N11757, N11737);
nand NAND3 (N11758, N11748, N3619, N11616);
xor XOR2 (N11759, N11751, N7169);
xor XOR2 (N11760, N11756, N7069);
buf BUF1 (N11761, N11759);
and AND2 (N11762, N11739, N7844);
or OR4 (N11763, N11754, N4553, N8460, N1974);
buf BUF1 (N11764, N11741);
nor NOR3 (N11765, N11764, N11340, N1075);
or OR4 (N11766, N11732, N8283, N5747, N2404);
nand NAND2 (N11767, N11757, N1015);
or OR3 (N11768, N11760, N940, N11630);
nand NAND4 (N11769, N11763, N1409, N916, N2779);
nor NOR2 (N11770, N11766, N3803);
nor NOR4 (N11771, N11752, N6741, N11097, N11515);
buf BUF1 (N11772, N11768);
nand NAND4 (N11773, N11761, N10518, N7076, N4933);
buf BUF1 (N11774, N11755);
nand NAND2 (N11775, N11769, N6665);
buf BUF1 (N11776, N11770);
xor XOR2 (N11777, N11772, N7060);
or OR2 (N11778, N11771, N5253);
buf BUF1 (N11779, N11765);
and AND4 (N11780, N11767, N10849, N7966, N11042);
not NOT1 (N11781, N11774);
not NOT1 (N11782, N11780);
not NOT1 (N11783, N11776);
nor NOR4 (N11784, N11762, N5766, N8643, N2740);
xor XOR2 (N11785, N11778, N7229);
nand NAND4 (N11786, N11785, N515, N7638, N5297);
nor NOR2 (N11787, N11784, N2474);
xor XOR2 (N11788, N11773, N3620);
and AND2 (N11789, N11779, N2299);
and AND4 (N11790, N11758, N9886, N3378, N746);
and AND4 (N11791, N11777, N10282, N2902, N2775);
buf BUF1 (N11792, N11775);
buf BUF1 (N11793, N11786);
and AND2 (N11794, N11791, N9272);
buf BUF1 (N11795, N11782);
buf BUF1 (N11796, N11788);
and AND4 (N11797, N11792, N204, N9134, N9893);
xor XOR2 (N11798, N11797, N9379);
or OR2 (N11799, N11794, N3819);
or OR2 (N11800, N11796, N5744);
and AND3 (N11801, N11793, N9071, N11633);
xor XOR2 (N11802, N11798, N5827);
and AND3 (N11803, N11790, N1506, N11528);
buf BUF1 (N11804, N11801);
xor XOR2 (N11805, N11783, N4091);
and AND2 (N11806, N11795, N6161);
nand NAND4 (N11807, N11804, N7753, N722, N10564);
buf BUF1 (N11808, N11806);
nor NOR4 (N11809, N11799, N1526, N10171, N11212);
not NOT1 (N11810, N11802);
not NOT1 (N11811, N11787);
nand NAND3 (N11812, N11809, N8466, N9544);
not NOT1 (N11813, N11807);
buf BUF1 (N11814, N11800);
not NOT1 (N11815, N11781);
and AND2 (N11816, N11808, N9552);
or OR2 (N11817, N11815, N6289);
and AND3 (N11818, N11817, N170, N9889);
xor XOR2 (N11819, N11814, N10773);
xor XOR2 (N11820, N11819, N7665);
not NOT1 (N11821, N11805);
or OR3 (N11822, N11816, N7132, N7994);
buf BUF1 (N11823, N11810);
and AND4 (N11824, N11813, N9638, N7452, N2624);
and AND3 (N11825, N11812, N2501, N3200);
or OR4 (N11826, N11824, N3575, N9871, N593);
nor NOR4 (N11827, N11803, N9011, N2156, N1528);
xor XOR2 (N11828, N11820, N1386);
nand NAND3 (N11829, N11818, N9064, N3509);
nor NOR3 (N11830, N11811, N8573, N9377);
xor XOR2 (N11831, N11821, N489);
xor XOR2 (N11832, N11789, N9406);
buf BUF1 (N11833, N11832);
or OR2 (N11834, N11822, N1619);
not NOT1 (N11835, N11829);
buf BUF1 (N11836, N11827);
nand NAND2 (N11837, N11825, N4442);
not NOT1 (N11838, N11833);
buf BUF1 (N11839, N11835);
not NOT1 (N11840, N11838);
not NOT1 (N11841, N11837);
nor NOR3 (N11842, N11831, N2334, N4790);
not NOT1 (N11843, N11823);
nor NOR4 (N11844, N11840, N4817, N9301, N7303);
nor NOR3 (N11845, N11844, N2208, N4943);
xor XOR2 (N11846, N11836, N3483);
and AND2 (N11847, N11839, N6543);
buf BUF1 (N11848, N11834);
not NOT1 (N11849, N11846);
not NOT1 (N11850, N11826);
not NOT1 (N11851, N11830);
nand NAND3 (N11852, N11842, N4976, N10151);
buf BUF1 (N11853, N11850);
nor NOR3 (N11854, N11852, N8183, N2535);
nor NOR3 (N11855, N11853, N3652, N4605);
or OR4 (N11856, N11848, N10089, N4855, N9782);
buf BUF1 (N11857, N11841);
or OR3 (N11858, N11845, N3366, N8934);
and AND3 (N11859, N11849, N3667, N10741);
and AND3 (N11860, N11828, N721, N438);
and AND3 (N11861, N11860, N2499, N8165);
buf BUF1 (N11862, N11854);
xor XOR2 (N11863, N11862, N2089);
xor XOR2 (N11864, N11858, N2504);
nand NAND2 (N11865, N11855, N3908);
nand NAND3 (N11866, N11859, N3245, N1754);
and AND2 (N11867, N11863, N11167);
or OR3 (N11868, N11857, N6972, N640);
or OR3 (N11869, N11861, N8164, N1242);
and AND3 (N11870, N11851, N3435, N8568);
or OR2 (N11871, N11843, N11305);
nand NAND4 (N11872, N11867, N2120, N451, N723);
nor NOR3 (N11873, N11856, N1658, N11834);
not NOT1 (N11874, N11872);
nor NOR3 (N11875, N11868, N3228, N10038);
buf BUF1 (N11876, N11875);
or OR2 (N11877, N11871, N3506);
nor NOR4 (N11878, N11865, N10067, N9684, N1435);
and AND3 (N11879, N11847, N1085, N3057);
xor XOR2 (N11880, N11874, N6109);
not NOT1 (N11881, N11873);
xor XOR2 (N11882, N11880, N10830);
buf BUF1 (N11883, N11876);
nor NOR3 (N11884, N11866, N5516, N5112);
buf BUF1 (N11885, N11864);
and AND4 (N11886, N11878, N4508, N3032, N9150);
xor XOR2 (N11887, N11870, N7881);
xor XOR2 (N11888, N11887, N9729);
nand NAND4 (N11889, N11883, N855, N4608, N7122);
xor XOR2 (N11890, N11869, N710);
not NOT1 (N11891, N11884);
nor NOR4 (N11892, N11891, N4586, N519, N11493);
and AND2 (N11893, N11892, N3077);
nand NAND4 (N11894, N11881, N10615, N9930, N4364);
nor NOR2 (N11895, N11886, N4851);
buf BUF1 (N11896, N11879);
not NOT1 (N11897, N11895);
or OR3 (N11898, N11890, N7697, N6470);
nor NOR3 (N11899, N11893, N11738, N1271);
not NOT1 (N11900, N11889);
xor XOR2 (N11901, N11897, N1752);
nor NOR3 (N11902, N11901, N3634, N8376);
not NOT1 (N11903, N11882);
xor XOR2 (N11904, N11902, N2338);
buf BUF1 (N11905, N11888);
and AND3 (N11906, N11896, N759, N8208);
not NOT1 (N11907, N11877);
nor NOR3 (N11908, N11903, N11775, N9408);
nand NAND3 (N11909, N11900, N2769, N7781);
buf BUF1 (N11910, N11898);
buf BUF1 (N11911, N11907);
nand NAND4 (N11912, N11906, N9734, N8002, N6647);
buf BUF1 (N11913, N11910);
nand NAND4 (N11914, N11885, N8302, N539, N971);
not NOT1 (N11915, N11905);
not NOT1 (N11916, N11894);
buf BUF1 (N11917, N11908);
and AND2 (N11918, N11909, N4557);
nor NOR4 (N11919, N11913, N9230, N4287, N658);
nand NAND4 (N11920, N11915, N3, N3378, N9472);
not NOT1 (N11921, N11920);
nor NOR4 (N11922, N11912, N4338, N5420, N11093);
or OR3 (N11923, N11899, N11858, N11281);
xor XOR2 (N11924, N11919, N754);
xor XOR2 (N11925, N11916, N4522);
buf BUF1 (N11926, N11917);
not NOT1 (N11927, N11923);
and AND2 (N11928, N11925, N4902);
xor XOR2 (N11929, N11911, N11229);
or OR2 (N11930, N11904, N11909);
nor NOR3 (N11931, N11930, N2989, N2233);
not NOT1 (N11932, N11921);
buf BUF1 (N11933, N11926);
not NOT1 (N11934, N11914);
nand NAND4 (N11935, N11932, N6584, N7707, N7851);
not NOT1 (N11936, N11933);
nand NAND2 (N11937, N11918, N8512);
and AND3 (N11938, N11929, N3700, N9445);
nor NOR2 (N11939, N11922, N7373);
nor NOR2 (N11940, N11927, N4773);
nand NAND2 (N11941, N11934, N4095);
or OR2 (N11942, N11937, N5305);
xor XOR2 (N11943, N11935, N7805);
xor XOR2 (N11944, N11924, N8289);
nand NAND3 (N11945, N11941, N2267, N10260);
or OR2 (N11946, N11931, N4272);
and AND3 (N11947, N11946, N10982, N6336);
and AND3 (N11948, N11939, N1950, N9641);
not NOT1 (N11949, N11936);
or OR2 (N11950, N11938, N6091);
buf BUF1 (N11951, N11948);
xor XOR2 (N11952, N11947, N6185);
and AND3 (N11953, N11944, N2262, N10411);
nor NOR4 (N11954, N11943, N4975, N11885, N5189);
nor NOR2 (N11955, N11928, N8559);
nor NOR3 (N11956, N11950, N7925, N9619);
not NOT1 (N11957, N11940);
buf BUF1 (N11958, N11942);
not NOT1 (N11959, N11953);
xor XOR2 (N11960, N11949, N1864);
buf BUF1 (N11961, N11952);
nor NOR3 (N11962, N11951, N7367, N3848);
and AND4 (N11963, N11962, N11796, N2797, N10169);
nand NAND2 (N11964, N11963, N3959);
or OR2 (N11965, N11960, N5076);
not NOT1 (N11966, N11965);
and AND2 (N11967, N11966, N7954);
nand NAND3 (N11968, N11967, N865, N2886);
nand NAND4 (N11969, N11956, N8670, N5090, N7219);
buf BUF1 (N11970, N11968);
xor XOR2 (N11971, N11970, N9331);
or OR3 (N11972, N11964, N7955, N168);
and AND3 (N11973, N11954, N2867, N8782);
buf BUF1 (N11974, N11961);
and AND4 (N11975, N11969, N6327, N6391, N4001);
nor NOR4 (N11976, N11973, N7734, N10895, N1634);
xor XOR2 (N11977, N11972, N7244);
nand NAND2 (N11978, N11958, N4);
or OR2 (N11979, N11959, N950);
xor XOR2 (N11980, N11977, N11621);
xor XOR2 (N11981, N11945, N803);
xor XOR2 (N11982, N11975, N8286);
and AND2 (N11983, N11979, N4337);
nand NAND2 (N11984, N11978, N862);
nor NOR2 (N11985, N11982, N228);
nor NOR4 (N11986, N11976, N1569, N2389, N1888);
not NOT1 (N11987, N11983);
xor XOR2 (N11988, N11981, N9390);
or OR2 (N11989, N11957, N5081);
nor NOR4 (N11990, N11986, N1047, N11547, N2052);
buf BUF1 (N11991, N11985);
buf BUF1 (N11992, N11989);
nand NAND2 (N11993, N11987, N11250);
or OR2 (N11994, N11988, N11602);
nand NAND2 (N11995, N11993, N9005);
not NOT1 (N11996, N11984);
and AND3 (N11997, N11992, N9058, N10410);
or OR3 (N11998, N11980, N10766, N4737);
and AND2 (N11999, N11974, N11392);
nand NAND2 (N12000, N11995, N3097);
not NOT1 (N12001, N11994);
xor XOR2 (N12002, N11997, N10212);
and AND3 (N12003, N11990, N8000, N6467);
buf BUF1 (N12004, N12003);
nor NOR3 (N12005, N11999, N2249, N4949);
nand NAND2 (N12006, N11991, N9927);
nand NAND4 (N12007, N12001, N3252, N8800, N4591);
xor XOR2 (N12008, N11998, N5589);
not NOT1 (N12009, N11971);
not NOT1 (N12010, N11955);
nor NOR2 (N12011, N12004, N9973);
buf BUF1 (N12012, N12007);
not NOT1 (N12013, N12005);
nand NAND2 (N12014, N12000, N8305);
xor XOR2 (N12015, N12012, N7215);
buf BUF1 (N12016, N12006);
not NOT1 (N12017, N12016);
or OR2 (N12018, N12014, N466);
nand NAND2 (N12019, N12018, N9087);
nor NOR3 (N12020, N12015, N3368, N8776);
nand NAND4 (N12021, N12013, N3646, N10089, N9040);
xor XOR2 (N12022, N12020, N1463);
or OR3 (N12023, N12002, N9565, N10017);
nor NOR3 (N12024, N12011, N9358, N4962);
xor XOR2 (N12025, N12010, N8407);
not NOT1 (N12026, N12019);
nand NAND4 (N12027, N12009, N799, N5358, N925);
nand NAND3 (N12028, N12025, N11898, N5808);
and AND4 (N12029, N12023, N9280, N2873, N7947);
xor XOR2 (N12030, N12017, N10236);
or OR2 (N12031, N12028, N4932);
nand NAND2 (N12032, N12030, N11817);
nand NAND2 (N12033, N12032, N5227);
not NOT1 (N12034, N12033);
buf BUF1 (N12035, N12024);
or OR4 (N12036, N12034, N2041, N232, N8626);
or OR2 (N12037, N12031, N9920);
nor NOR3 (N12038, N12029, N2180, N8551);
xor XOR2 (N12039, N12035, N6176);
nand NAND2 (N12040, N12027, N4672);
and AND3 (N12041, N11996, N2060, N9421);
not NOT1 (N12042, N12038);
nor NOR2 (N12043, N12037, N4937);
or OR2 (N12044, N12039, N9821);
or OR3 (N12045, N12042, N445, N5130);
not NOT1 (N12046, N12040);
nor NOR2 (N12047, N12022, N7474);
and AND4 (N12048, N12036, N10777, N3077, N9938);
nand NAND2 (N12049, N12043, N5247);
not NOT1 (N12050, N12008);
not NOT1 (N12051, N12046);
or OR2 (N12052, N12041, N4412);
or OR4 (N12053, N12049, N5394, N1149, N6951);
and AND4 (N12054, N12021, N1278, N1269, N354);
xor XOR2 (N12055, N12052, N5697);
nor NOR2 (N12056, N12048, N6805);
xor XOR2 (N12057, N12054, N1147);
buf BUF1 (N12058, N12053);
nand NAND3 (N12059, N12058, N3870, N4368);
not NOT1 (N12060, N12056);
and AND2 (N12061, N12060, N5558);
buf BUF1 (N12062, N12055);
not NOT1 (N12063, N12044);
nor NOR4 (N12064, N12045, N10988, N5369, N6027);
and AND2 (N12065, N12057, N6185);
or OR3 (N12066, N12065, N2352, N6241);
xor XOR2 (N12067, N12062, N2720);
or OR2 (N12068, N12059, N6205);
and AND4 (N12069, N12050, N8613, N6864, N1501);
and AND3 (N12070, N12068, N10115, N3597);
nand NAND4 (N12071, N12069, N5292, N7466, N9771);
nor NOR3 (N12072, N12067, N3039, N1726);
not NOT1 (N12073, N12026);
nand NAND4 (N12074, N12072, N5479, N4722, N5155);
xor XOR2 (N12075, N12074, N6249);
nand NAND4 (N12076, N12071, N2249, N457, N6326);
or OR4 (N12077, N12066, N217, N2261, N236);
and AND4 (N12078, N12075, N5548, N2621, N205);
nand NAND2 (N12079, N12047, N3035);
xor XOR2 (N12080, N12079, N9919);
and AND3 (N12081, N12080, N7081, N1775);
and AND3 (N12082, N12073, N437, N6893);
nand NAND3 (N12083, N12061, N3586, N6379);
not NOT1 (N12084, N12051);
buf BUF1 (N12085, N12063);
nand NAND2 (N12086, N12078, N10867);
xor XOR2 (N12087, N12082, N1215);
buf BUF1 (N12088, N12064);
nand NAND2 (N12089, N12077, N11820);
nor NOR4 (N12090, N12070, N8502, N8453, N11428);
buf BUF1 (N12091, N12086);
not NOT1 (N12092, N12089);
not NOT1 (N12093, N12084);
nor NOR3 (N12094, N12087, N5157, N1814);
or OR2 (N12095, N12094, N1708);
nor NOR4 (N12096, N12093, N3750, N1069, N11175);
or OR2 (N12097, N12088, N5395);
nor NOR4 (N12098, N12097, N3025, N6735, N7329);
nor NOR4 (N12099, N12096, N1140, N552, N9954);
nor NOR4 (N12100, N12081, N549, N10684, N5557);
and AND2 (N12101, N12091, N9150);
nand NAND3 (N12102, N12083, N7614, N2644);
or OR4 (N12103, N12099, N2168, N94, N8955);
not NOT1 (N12104, N12098);
nor NOR4 (N12105, N12095, N9324, N3623, N7185);
and AND3 (N12106, N12092, N6239, N2538);
or OR3 (N12107, N12102, N6832, N10910);
buf BUF1 (N12108, N12107);
not NOT1 (N12109, N12090);
and AND2 (N12110, N12108, N7596);
nand NAND3 (N12111, N12076, N1485, N1608);
and AND4 (N12112, N12085, N8830, N10353, N7368);
or OR2 (N12113, N12105, N9086);
or OR4 (N12114, N12100, N11373, N7587, N3260);
and AND2 (N12115, N12104, N9280);
not NOT1 (N12116, N12109);
and AND2 (N12117, N12112, N4411);
xor XOR2 (N12118, N12106, N3227);
nand NAND2 (N12119, N12116, N11354);
not NOT1 (N12120, N12114);
nor NOR3 (N12121, N12111, N2238, N6542);
or OR4 (N12122, N12121, N7127, N6246, N137);
xor XOR2 (N12123, N12122, N10855);
or OR4 (N12124, N12123, N9268, N1754, N9315);
nand NAND2 (N12125, N12110, N3968);
not NOT1 (N12126, N12117);
nor NOR2 (N12127, N12120, N3715);
xor XOR2 (N12128, N12103, N870);
xor XOR2 (N12129, N12126, N12100);
nor NOR4 (N12130, N12124, N8947, N10558, N5537);
buf BUF1 (N12131, N12115);
or OR2 (N12132, N12101, N6470);
nand NAND2 (N12133, N12119, N8593);
xor XOR2 (N12134, N12113, N4130);
xor XOR2 (N12135, N12128, N9083);
nor NOR2 (N12136, N12135, N5786);
xor XOR2 (N12137, N12134, N2629);
not NOT1 (N12138, N12118);
nand NAND3 (N12139, N12130, N10181, N3478);
and AND2 (N12140, N12139, N6241);
and AND3 (N12141, N12136, N4659, N11266);
buf BUF1 (N12142, N12129);
not NOT1 (N12143, N12127);
nand NAND3 (N12144, N12141, N10825, N3510);
not NOT1 (N12145, N12142);
nor NOR3 (N12146, N12132, N9245, N662);
and AND3 (N12147, N12133, N11110, N4468);
not NOT1 (N12148, N12140);
not NOT1 (N12149, N12137);
nand NAND2 (N12150, N12146, N9161);
nor NOR4 (N12151, N12145, N8308, N9963, N9157);
or OR4 (N12152, N12148, N10417, N789, N1174);
not NOT1 (N12153, N12147);
nor NOR2 (N12154, N12151, N11190);
nor NOR4 (N12155, N12131, N9742, N1365, N1101);
nand NAND4 (N12156, N12155, N1291, N2130, N5823);
or OR2 (N12157, N12152, N10901);
and AND2 (N12158, N12138, N10006);
not NOT1 (N12159, N12153);
nor NOR3 (N12160, N12159, N7964, N7627);
not NOT1 (N12161, N12157);
not NOT1 (N12162, N12161);
or OR3 (N12163, N12158, N10714, N114);
nor NOR2 (N12164, N12160, N6404);
and AND2 (N12165, N12154, N6747);
not NOT1 (N12166, N12163);
buf BUF1 (N12167, N12125);
nand NAND4 (N12168, N12156, N2404, N6329, N2059);
xor XOR2 (N12169, N12167, N9566);
nand NAND4 (N12170, N12162, N5891, N296, N10451);
or OR3 (N12171, N12149, N3386, N5640);
xor XOR2 (N12172, N12169, N11101);
not NOT1 (N12173, N12165);
xor XOR2 (N12174, N12144, N10679);
xor XOR2 (N12175, N12172, N7285);
xor XOR2 (N12176, N12150, N11827);
and AND3 (N12177, N12168, N805, N1138);
nand NAND2 (N12178, N12173, N756);
not NOT1 (N12179, N12143);
or OR2 (N12180, N12164, N7018);
xor XOR2 (N12181, N12166, N10119);
nor NOR3 (N12182, N12180, N1531, N7946);
nand NAND3 (N12183, N12174, N5872, N6260);
xor XOR2 (N12184, N12175, N4325);
buf BUF1 (N12185, N12183);
and AND4 (N12186, N12184, N7187, N4322, N10489);
or OR3 (N12187, N12171, N10760, N10846);
and AND4 (N12188, N12179, N10510, N8115, N6645);
buf BUF1 (N12189, N12170);
xor XOR2 (N12190, N12181, N7117);
xor XOR2 (N12191, N12190, N9962);
nor NOR3 (N12192, N12189, N1027, N3019);
xor XOR2 (N12193, N12187, N4966);
or OR3 (N12194, N12176, N9252, N1452);
nor NOR2 (N12195, N12193, N1618);
not NOT1 (N12196, N12185);
or OR2 (N12197, N12195, N9451);
xor XOR2 (N12198, N12197, N5996);
or OR3 (N12199, N12188, N5114, N8808);
buf BUF1 (N12200, N12194);
not NOT1 (N12201, N12182);
and AND2 (N12202, N12201, N2979);
nand NAND2 (N12203, N12200, N10245);
or OR2 (N12204, N12186, N8929);
xor XOR2 (N12205, N12177, N10176);
or OR3 (N12206, N12202, N4214, N11471);
nand NAND3 (N12207, N12196, N7230, N2416);
buf BUF1 (N12208, N12205);
xor XOR2 (N12209, N12208, N6877);
and AND3 (N12210, N12199, N4114, N11303);
xor XOR2 (N12211, N12206, N10570);
or OR4 (N12212, N12209, N10632, N8357, N3190);
nor NOR3 (N12213, N12198, N10198, N1168);
and AND4 (N12214, N12191, N7392, N2916, N1);
not NOT1 (N12215, N12178);
nor NOR3 (N12216, N12213, N7043, N4625);
and AND4 (N12217, N12211, N3980, N995, N8840);
xor XOR2 (N12218, N12204, N9173);
not NOT1 (N12219, N12214);
buf BUF1 (N12220, N12207);
xor XOR2 (N12221, N12218, N4402);
nor NOR2 (N12222, N12212, N11598);
and AND4 (N12223, N12210, N5167, N3063, N11119);
xor XOR2 (N12224, N12220, N11456);
or OR2 (N12225, N12221, N7705);
buf BUF1 (N12226, N12224);
or OR2 (N12227, N12216, N7056);
or OR2 (N12228, N12226, N5321);
buf BUF1 (N12229, N12228);
not NOT1 (N12230, N12227);
buf BUF1 (N12231, N12203);
xor XOR2 (N12232, N12192, N3701);
not NOT1 (N12233, N12230);
or OR4 (N12234, N12219, N3288, N5751, N4775);
or OR4 (N12235, N12231, N2326, N10693, N294);
and AND4 (N12236, N12233, N2336, N3592, N2231);
nor NOR3 (N12237, N12236, N3006, N5610);
nand NAND2 (N12238, N12234, N6155);
not NOT1 (N12239, N12229);
or OR4 (N12240, N12225, N2199, N10320, N5493);
and AND2 (N12241, N12223, N10616);
xor XOR2 (N12242, N12237, N11598);
not NOT1 (N12243, N12235);
nor NOR3 (N12244, N12241, N10972, N6839);
xor XOR2 (N12245, N12222, N11084);
buf BUF1 (N12246, N12245);
not NOT1 (N12247, N12242);
or OR4 (N12248, N12240, N8935, N10638, N4334);
or OR3 (N12249, N12243, N11892, N7408);
not NOT1 (N12250, N12232);
buf BUF1 (N12251, N12217);
nor NOR4 (N12252, N12249, N6818, N2026, N2542);
or OR3 (N12253, N12247, N1674, N3022);
nor NOR2 (N12254, N12251, N7798);
not NOT1 (N12255, N12248);
xor XOR2 (N12256, N12215, N4399);
xor XOR2 (N12257, N12246, N644);
buf BUF1 (N12258, N12256);
nor NOR2 (N12259, N12257, N11450);
and AND2 (N12260, N12252, N224);
and AND2 (N12261, N12239, N7057);
xor XOR2 (N12262, N12253, N6839);
and AND3 (N12263, N12258, N5938, N3016);
or OR4 (N12264, N12262, N10778, N1281, N10295);
or OR4 (N12265, N12250, N7436, N8376, N10744);
and AND2 (N12266, N12264, N6365);
or OR4 (N12267, N12265, N8074, N566, N1377);
and AND4 (N12268, N12263, N685, N11889, N4164);
or OR3 (N12269, N12244, N4978, N8125);
xor XOR2 (N12270, N12267, N1693);
and AND3 (N12271, N12255, N5722, N3015);
buf BUF1 (N12272, N12270);
xor XOR2 (N12273, N12259, N5561);
nor NOR2 (N12274, N12269, N3287);
nand NAND4 (N12275, N12268, N1788, N4853, N347);
and AND3 (N12276, N12266, N4354, N2829);
or OR4 (N12277, N12272, N8845, N2004, N10063);
and AND3 (N12278, N12238, N9546, N1452);
buf BUF1 (N12279, N12276);
buf BUF1 (N12280, N12254);
nand NAND4 (N12281, N12280, N8802, N956, N2231);
xor XOR2 (N12282, N12277, N8680);
or OR2 (N12283, N12281, N1308);
nor NOR3 (N12284, N12278, N9343, N6401);
or OR2 (N12285, N12271, N3858);
and AND3 (N12286, N12279, N4883, N11088);
not NOT1 (N12287, N12261);
nand NAND2 (N12288, N12275, N5291);
xor XOR2 (N12289, N12288, N297);
or OR4 (N12290, N12284, N2671, N4782, N1119);
or OR4 (N12291, N12290, N6251, N7879, N11314);
nor NOR2 (N12292, N12283, N8766);
not NOT1 (N12293, N12285);
not NOT1 (N12294, N12291);
nor NOR4 (N12295, N12286, N606, N6629, N5022);
xor XOR2 (N12296, N12294, N5256);
not NOT1 (N12297, N12260);
nor NOR2 (N12298, N12293, N5849);
or OR2 (N12299, N12287, N6601);
nand NAND4 (N12300, N12295, N9377, N11053, N1158);
nor NOR2 (N12301, N12297, N3179);
xor XOR2 (N12302, N12282, N10333);
and AND3 (N12303, N12302, N2335, N11636);
xor XOR2 (N12304, N12289, N427);
nor NOR3 (N12305, N12292, N9772, N8184);
nor NOR3 (N12306, N12299, N8974, N9866);
nor NOR3 (N12307, N12298, N3059, N3737);
and AND4 (N12308, N12301, N2929, N11241, N5207);
not NOT1 (N12309, N12305);
xor XOR2 (N12310, N12274, N11352);
nor NOR2 (N12311, N12304, N5854);
or OR2 (N12312, N12296, N11840);
buf BUF1 (N12313, N12306);
nor NOR3 (N12314, N12310, N7119, N2801);
and AND3 (N12315, N12300, N9305, N10632);
buf BUF1 (N12316, N12309);
nor NOR4 (N12317, N12315, N9936, N3162, N7581);
xor XOR2 (N12318, N12312, N11528);
buf BUF1 (N12319, N12313);
not NOT1 (N12320, N12316);
xor XOR2 (N12321, N12311, N10133);
xor XOR2 (N12322, N12317, N45);
or OR2 (N12323, N12322, N4156);
nor NOR2 (N12324, N12323, N7990);
and AND3 (N12325, N12308, N10081, N2897);
nand NAND3 (N12326, N12318, N8574, N2239);
buf BUF1 (N12327, N12307);
and AND2 (N12328, N12319, N7601);
nand NAND3 (N12329, N12324, N11156, N1681);
or OR4 (N12330, N12303, N5768, N4396, N11131);
and AND3 (N12331, N12330, N11349, N2315);
buf BUF1 (N12332, N12331);
nor NOR3 (N12333, N12329, N5352, N2733);
nand NAND2 (N12334, N12273, N2545);
nand NAND2 (N12335, N12332, N7908);
or OR2 (N12336, N12320, N4275);
or OR4 (N12337, N12314, N4570, N3587, N8266);
xor XOR2 (N12338, N12333, N232);
and AND2 (N12339, N12336, N11672);
not NOT1 (N12340, N12328);
buf BUF1 (N12341, N12335);
buf BUF1 (N12342, N12321);
not NOT1 (N12343, N12334);
nor NOR3 (N12344, N12325, N4198, N2327);
buf BUF1 (N12345, N12338);
buf BUF1 (N12346, N12344);
not NOT1 (N12347, N12346);
or OR2 (N12348, N12326, N6562);
buf BUF1 (N12349, N12348);
and AND3 (N12350, N12340, N11098, N9864);
buf BUF1 (N12351, N12339);
or OR2 (N12352, N12342, N495);
and AND2 (N12353, N12341, N3739);
not NOT1 (N12354, N12351);
and AND2 (N12355, N12353, N8939);
buf BUF1 (N12356, N12355);
not NOT1 (N12357, N12343);
and AND4 (N12358, N12354, N11087, N9871, N2299);
and AND3 (N12359, N12337, N11844, N1664);
or OR2 (N12360, N12327, N5101);
nor NOR2 (N12361, N12349, N2439);
nor NOR3 (N12362, N12357, N555, N10090);
not NOT1 (N12363, N12358);
and AND2 (N12364, N12356, N11834);
xor XOR2 (N12365, N12347, N7276);
nor NOR4 (N12366, N12352, N3343, N9807, N6812);
xor XOR2 (N12367, N12366, N2072);
xor XOR2 (N12368, N12350, N4303);
xor XOR2 (N12369, N12359, N9639);
or OR3 (N12370, N12368, N8901, N1786);
buf BUF1 (N12371, N12361);
nand NAND4 (N12372, N12370, N5776, N5608, N2031);
xor XOR2 (N12373, N12369, N3073);
not NOT1 (N12374, N12345);
buf BUF1 (N12375, N12363);
buf BUF1 (N12376, N12360);
buf BUF1 (N12377, N12372);
not NOT1 (N12378, N12362);
buf BUF1 (N12379, N12373);
not NOT1 (N12380, N12374);
nand NAND2 (N12381, N12364, N5495);
or OR2 (N12382, N12376, N11532);
nor NOR4 (N12383, N12365, N6981, N7168, N5704);
xor XOR2 (N12384, N12382, N11890);
xor XOR2 (N12385, N12371, N1705);
xor XOR2 (N12386, N12383, N2246);
and AND4 (N12387, N12385, N12374, N6655, N1478);
or OR4 (N12388, N12377, N4973, N6595, N11484);
or OR4 (N12389, N12380, N3727, N1952, N3473);
nand NAND2 (N12390, N12378, N9123);
or OR2 (N12391, N12386, N7402);
not NOT1 (N12392, N12381);
xor XOR2 (N12393, N12375, N12017);
nor NOR2 (N12394, N12390, N4956);
or OR2 (N12395, N12384, N5217);
nand NAND3 (N12396, N12393, N3421, N9700);
and AND2 (N12397, N12395, N2360);
xor XOR2 (N12398, N12389, N1690);
nand NAND3 (N12399, N12398, N8050, N3135);
nand NAND3 (N12400, N12379, N8263, N3425);
buf BUF1 (N12401, N12397);
not NOT1 (N12402, N12399);
nor NOR2 (N12403, N12367, N507);
nand NAND4 (N12404, N12394, N7809, N9740, N11766);
or OR2 (N12405, N12400, N7588);
and AND2 (N12406, N12405, N632);
not NOT1 (N12407, N12403);
buf BUF1 (N12408, N12392);
and AND2 (N12409, N12402, N5794);
or OR4 (N12410, N12391, N7937, N6799, N7311);
or OR3 (N12411, N12407, N10679, N5396);
or OR3 (N12412, N12408, N5814, N1011);
not NOT1 (N12413, N12411);
and AND3 (N12414, N12401, N7466, N11846);
nor NOR4 (N12415, N12414, N11392, N171, N9307);
buf BUF1 (N12416, N12406);
xor XOR2 (N12417, N12387, N3895);
not NOT1 (N12418, N12412);
xor XOR2 (N12419, N12417, N7926);
nor NOR3 (N12420, N12416, N11921, N4814);
or OR3 (N12421, N12413, N11552, N12331);
or OR3 (N12422, N12410, N2337, N11903);
xor XOR2 (N12423, N12409, N3612);
or OR4 (N12424, N12419, N1338, N6036, N7720);
nor NOR2 (N12425, N12420, N2283);
xor XOR2 (N12426, N12415, N1201);
xor XOR2 (N12427, N12423, N6422);
and AND3 (N12428, N12421, N5570, N5513);
buf BUF1 (N12429, N12422);
buf BUF1 (N12430, N12427);
or OR3 (N12431, N12430, N5899, N4953);
or OR3 (N12432, N12431, N9190, N916);
buf BUF1 (N12433, N12424);
buf BUF1 (N12434, N12426);
buf BUF1 (N12435, N12396);
nand NAND2 (N12436, N12433, N8735);
nand NAND4 (N12437, N12404, N1494, N5766, N4288);
not NOT1 (N12438, N12436);
xor XOR2 (N12439, N12432, N7057);
nand NAND4 (N12440, N12438, N7242, N7176, N4829);
not NOT1 (N12441, N12439);
and AND3 (N12442, N12428, N5475, N574);
or OR2 (N12443, N12418, N3777);
nor NOR3 (N12444, N12425, N8584, N9860);
nand NAND3 (N12445, N12434, N4809, N3721);
xor XOR2 (N12446, N12445, N330);
and AND3 (N12447, N12435, N9217, N3349);
and AND3 (N12448, N12443, N10637, N11617);
nor NOR3 (N12449, N12448, N5416, N8441);
and AND2 (N12450, N12449, N3555);
xor XOR2 (N12451, N12447, N10150);
nor NOR3 (N12452, N12444, N3351, N974);
nand NAND4 (N12453, N12451, N3280, N9825, N6857);
nand NAND3 (N12454, N12429, N4691, N4358);
buf BUF1 (N12455, N12450);
nand NAND4 (N12456, N12441, N698, N9682, N11273);
nor NOR4 (N12457, N12452, N8988, N3961, N7682);
and AND3 (N12458, N12388, N5703, N10453);
not NOT1 (N12459, N12456);
buf BUF1 (N12460, N12442);
nand NAND4 (N12461, N12457, N8602, N8998, N9066);
and AND4 (N12462, N12461, N2329, N3477, N10819);
xor XOR2 (N12463, N12446, N9966);
xor XOR2 (N12464, N12455, N11711);
nor NOR2 (N12465, N12462, N968);
not NOT1 (N12466, N12440);
not NOT1 (N12467, N12453);
buf BUF1 (N12468, N12467);
xor XOR2 (N12469, N12460, N10851);
or OR4 (N12470, N12454, N10241, N5424, N2781);
nand NAND3 (N12471, N12469, N2093, N11428);
nor NOR3 (N12472, N12465, N10454, N11469);
buf BUF1 (N12473, N12470);
and AND4 (N12474, N12464, N10284, N6227, N4124);
or OR3 (N12475, N12471, N8888, N1057);
not NOT1 (N12476, N12472);
and AND4 (N12477, N12459, N4429, N6117, N3805);
not NOT1 (N12478, N12477);
xor XOR2 (N12479, N12476, N8513);
nand NAND2 (N12480, N12473, N10232);
not NOT1 (N12481, N12480);
and AND4 (N12482, N12458, N7787, N7580, N10703);
nor NOR4 (N12483, N12481, N12033, N859, N5987);
or OR2 (N12484, N12437, N10504);
or OR3 (N12485, N12483, N12174, N10692);
not NOT1 (N12486, N12485);
nor NOR3 (N12487, N12479, N275, N10142);
and AND3 (N12488, N12468, N2374, N1105);
not NOT1 (N12489, N12475);
and AND2 (N12490, N12486, N12379);
or OR4 (N12491, N12490, N868, N2468, N3757);
nand NAND4 (N12492, N12491, N1112, N4608, N3004);
not NOT1 (N12493, N12489);
or OR3 (N12494, N12466, N12117, N1554);
or OR3 (N12495, N12493, N6644, N9429);
nand NAND3 (N12496, N12492, N7111, N10019);
or OR4 (N12497, N12487, N4400, N6655, N12165);
or OR2 (N12498, N12482, N4471);
xor XOR2 (N12499, N12488, N4157);
not NOT1 (N12500, N12474);
or OR4 (N12501, N12478, N3796, N2771, N10406);
nand NAND2 (N12502, N12499, N10059);
buf BUF1 (N12503, N12497);
and AND3 (N12504, N12498, N70, N9975);
or OR3 (N12505, N12503, N3305, N5166);
not NOT1 (N12506, N12496);
xor XOR2 (N12507, N12484, N331);
xor XOR2 (N12508, N12505, N2247);
xor XOR2 (N12509, N12507, N6112);
and AND4 (N12510, N12502, N9208, N2225, N1528);
buf BUF1 (N12511, N12510);
nor NOR2 (N12512, N12501, N11156);
buf BUF1 (N12513, N12494);
not NOT1 (N12514, N12495);
xor XOR2 (N12515, N12463, N1353);
or OR4 (N12516, N12500, N8933, N10223, N6722);
xor XOR2 (N12517, N12516, N1675);
nand NAND3 (N12518, N12512, N8658, N2812);
not NOT1 (N12519, N12513);
not NOT1 (N12520, N12518);
nor NOR3 (N12521, N12517, N9824, N5128);
buf BUF1 (N12522, N12515);
buf BUF1 (N12523, N12520);
and AND2 (N12524, N12506, N3374);
nand NAND2 (N12525, N12523, N10703);
or OR2 (N12526, N12514, N10300);
nand NAND3 (N12527, N12508, N3268, N9150);
not NOT1 (N12528, N12522);
or OR4 (N12529, N12526, N2687, N2990, N3018);
nand NAND4 (N12530, N12527, N2046, N7391, N7404);
nor NOR3 (N12531, N12504, N6333, N7271);
not NOT1 (N12532, N12525);
xor XOR2 (N12533, N12532, N9682);
nand NAND2 (N12534, N12524, N7145);
nand NAND3 (N12535, N12531, N4362, N7743);
not NOT1 (N12536, N12528);
nand NAND3 (N12537, N12535, N9931, N12459);
not NOT1 (N12538, N12536);
nor NOR2 (N12539, N12537, N4669);
or OR4 (N12540, N12521, N12280, N4171, N2641);
nand NAND4 (N12541, N12533, N12540, N2873, N11154);
nand NAND2 (N12542, N11405, N6619);
nor NOR3 (N12543, N12530, N11292, N8525);
and AND3 (N12544, N12511, N11636, N6613);
not NOT1 (N12545, N12534);
nor NOR4 (N12546, N12545, N5365, N7450, N7049);
not NOT1 (N12547, N12542);
or OR2 (N12548, N12539, N5889);
xor XOR2 (N12549, N12548, N3251);
not NOT1 (N12550, N12547);
not NOT1 (N12551, N12519);
buf BUF1 (N12552, N12551);
nand NAND4 (N12553, N12538, N2894, N7173, N3001);
not NOT1 (N12554, N12509);
nor NOR3 (N12555, N12544, N7113, N9980);
not NOT1 (N12556, N12549);
xor XOR2 (N12557, N12555, N12129);
and AND4 (N12558, N12554, N2770, N3496, N6494);
xor XOR2 (N12559, N12556, N11988);
nor NOR2 (N12560, N12541, N7690);
and AND2 (N12561, N12557, N1859);
nand NAND2 (N12562, N12553, N12401);
nand NAND4 (N12563, N12560, N2093, N5651, N12159);
nor NOR3 (N12564, N12562, N1400, N5689);
not NOT1 (N12565, N12564);
not NOT1 (N12566, N12529);
nand NAND4 (N12567, N12552, N9739, N583, N8456);
nand NAND4 (N12568, N12546, N8166, N6529, N9030);
and AND2 (N12569, N12568, N9506);
buf BUF1 (N12570, N12550);
or OR3 (N12571, N12561, N3955, N1390);
xor XOR2 (N12572, N12565, N5054);
nor NOR3 (N12573, N12572, N10258, N4638);
nor NOR2 (N12574, N12563, N5925);
or OR4 (N12575, N12569, N8656, N7648, N11058);
xor XOR2 (N12576, N12574, N3847);
buf BUF1 (N12577, N12558);
nor NOR4 (N12578, N12570, N4350, N2385, N8744);
nand NAND2 (N12579, N12559, N4015);
not NOT1 (N12580, N12573);
nand NAND3 (N12581, N12579, N1655, N4571);
xor XOR2 (N12582, N12567, N8095);
or OR4 (N12583, N12581, N4065, N743, N743);
not NOT1 (N12584, N12543);
buf BUF1 (N12585, N12577);
not NOT1 (N12586, N12585);
or OR3 (N12587, N12575, N819, N2088);
and AND3 (N12588, N12584, N8780, N3088);
buf BUF1 (N12589, N12576);
nand NAND2 (N12590, N12566, N8859);
buf BUF1 (N12591, N12588);
not NOT1 (N12592, N12578);
and AND2 (N12593, N12587, N9694);
nor NOR4 (N12594, N12593, N11157, N2197, N9834);
buf BUF1 (N12595, N12594);
or OR4 (N12596, N12580, N7103, N11471, N1814);
or OR3 (N12597, N12595, N2224, N3650);
and AND2 (N12598, N12582, N7846);
or OR4 (N12599, N12583, N11533, N8277, N10894);
nor NOR3 (N12600, N12599, N2400, N3228);
and AND4 (N12601, N12590, N12182, N10221, N1975);
xor XOR2 (N12602, N12571, N9785);
buf BUF1 (N12603, N12600);
nand NAND3 (N12604, N12597, N9959, N557);
and AND2 (N12605, N12603, N11128);
nand NAND3 (N12606, N12592, N9056, N473);
nor NOR3 (N12607, N12586, N10426, N7506);
nand NAND3 (N12608, N12598, N5660, N5882);
nand NAND4 (N12609, N12596, N6445, N5448, N12287);
nand NAND3 (N12610, N12607, N9140, N2972);
nand NAND2 (N12611, N12609, N9268);
not NOT1 (N12612, N12591);
nand NAND3 (N12613, N12601, N6597, N6397);
and AND3 (N12614, N12611, N2736, N773);
not NOT1 (N12615, N12614);
or OR4 (N12616, N12610, N5729, N2876, N6557);
and AND4 (N12617, N12613, N1948, N5354, N6070);
nor NOR2 (N12618, N12605, N9884);
nand NAND2 (N12619, N12604, N9956);
or OR2 (N12620, N12618, N1372);
or OR3 (N12621, N12608, N12441, N4699);
not NOT1 (N12622, N12606);
buf BUF1 (N12623, N12621);
or OR4 (N12624, N12622, N7114, N3683, N7223);
buf BUF1 (N12625, N12602);
buf BUF1 (N12626, N12620);
nor NOR2 (N12627, N12617, N6387);
not NOT1 (N12628, N12615);
not NOT1 (N12629, N12624);
xor XOR2 (N12630, N12625, N9747);
or OR4 (N12631, N12626, N12026, N1679, N1329);
not NOT1 (N12632, N12589);
not NOT1 (N12633, N12619);
nor NOR2 (N12634, N12629, N11968);
nor NOR2 (N12635, N12634, N4464);
xor XOR2 (N12636, N12612, N12344);
buf BUF1 (N12637, N12623);
nand NAND4 (N12638, N12628, N12023, N11076, N5017);
xor XOR2 (N12639, N12630, N9831);
buf BUF1 (N12640, N12616);
xor XOR2 (N12641, N12632, N2712);
and AND4 (N12642, N12635, N5935, N1772, N2925);
nand NAND4 (N12643, N12627, N4873, N8000, N1209);
not NOT1 (N12644, N12633);
or OR4 (N12645, N12640, N10239, N4334, N3636);
not NOT1 (N12646, N12643);
xor XOR2 (N12647, N12636, N10286);
xor XOR2 (N12648, N12639, N1681);
or OR4 (N12649, N12648, N7979, N8638, N1357);
or OR3 (N12650, N12647, N4353, N7436);
buf BUF1 (N12651, N12637);
xor XOR2 (N12652, N12631, N1528);
xor XOR2 (N12653, N12645, N11947);
and AND2 (N12654, N12638, N7804);
xor XOR2 (N12655, N12650, N7483);
nand NAND2 (N12656, N12654, N10702);
and AND2 (N12657, N12642, N3905);
and AND3 (N12658, N12655, N10951, N1642);
xor XOR2 (N12659, N12658, N5407);
or OR3 (N12660, N12649, N8854, N2001);
or OR2 (N12661, N12656, N8213);
xor XOR2 (N12662, N12644, N5053);
and AND2 (N12663, N12646, N11020);
nor NOR2 (N12664, N12641, N5606);
nor NOR4 (N12665, N12661, N1604, N11710, N5617);
or OR3 (N12666, N12652, N10154, N12309);
or OR3 (N12667, N12657, N4746, N9884);
or OR2 (N12668, N12659, N9613);
not NOT1 (N12669, N12653);
and AND2 (N12670, N12665, N1888);
or OR4 (N12671, N12666, N1837, N4737, N9600);
nor NOR4 (N12672, N12664, N7321, N5545, N11108);
nor NOR4 (N12673, N12670, N8676, N7767, N5177);
nand NAND4 (N12674, N12671, N10086, N2222, N8131);
xor XOR2 (N12675, N12663, N4253);
or OR3 (N12676, N12672, N5142, N885);
nand NAND3 (N12677, N12675, N496, N8241);
nand NAND2 (N12678, N12651, N3952);
buf BUF1 (N12679, N12676);
buf BUF1 (N12680, N12667);
nor NOR3 (N12681, N12668, N142, N4377);
buf BUF1 (N12682, N12680);
and AND2 (N12683, N12681, N9701);
not NOT1 (N12684, N12673);
xor XOR2 (N12685, N12683, N4402);
buf BUF1 (N12686, N12685);
xor XOR2 (N12687, N12678, N1480);
nor NOR3 (N12688, N12682, N5582, N3651);
nor NOR4 (N12689, N12687, N4525, N4697, N10932);
not NOT1 (N12690, N12679);
and AND4 (N12691, N12690, N1701, N8360, N6026);
or OR2 (N12692, N12688, N7961);
or OR4 (N12693, N12692, N11204, N1804, N10056);
xor XOR2 (N12694, N12669, N1904);
or OR2 (N12695, N12686, N10447);
nand NAND2 (N12696, N12677, N7211);
nor NOR2 (N12697, N12660, N6924);
and AND2 (N12698, N12693, N554);
xor XOR2 (N12699, N12691, N2938);
not NOT1 (N12700, N12695);
buf BUF1 (N12701, N12662);
and AND4 (N12702, N12694, N6674, N5498, N4094);
or OR4 (N12703, N12684, N11810, N2658, N821);
not NOT1 (N12704, N12699);
nand NAND4 (N12705, N12674, N629, N11704, N7222);
or OR3 (N12706, N12704, N7979, N2383);
not NOT1 (N12707, N12703);
buf BUF1 (N12708, N12696);
xor XOR2 (N12709, N12697, N9089);
nand NAND4 (N12710, N12698, N3183, N987, N6506);
and AND4 (N12711, N12708, N5295, N8594, N12023);
buf BUF1 (N12712, N12711);
nor NOR3 (N12713, N12689, N1488, N12355);
not NOT1 (N12714, N12713);
not NOT1 (N12715, N12710);
nor NOR4 (N12716, N12709, N66, N11061, N9937);
or OR2 (N12717, N12707, N8412);
or OR2 (N12718, N12702, N2857);
nand NAND4 (N12719, N12717, N10573, N813, N9508);
or OR3 (N12720, N12706, N3936, N8387);
nor NOR2 (N12721, N12705, N12245);
nand NAND3 (N12722, N12721, N8964, N758);
nor NOR2 (N12723, N12715, N3956);
or OR4 (N12724, N12700, N7284, N11875, N1438);
xor XOR2 (N12725, N12712, N11515);
not NOT1 (N12726, N12724);
nor NOR4 (N12727, N12726, N3506, N2620, N6391);
buf BUF1 (N12728, N12714);
or OR3 (N12729, N12716, N2879, N4827);
or OR4 (N12730, N12728, N4654, N10187, N608);
nor NOR4 (N12731, N12723, N10531, N8660, N6478);
and AND3 (N12732, N12719, N2773, N6878);
nand NAND4 (N12733, N12731, N5490, N6503, N1013);
xor XOR2 (N12734, N12720, N8754);
nand NAND2 (N12735, N12733, N4048);
or OR3 (N12736, N12725, N2830, N6309);
and AND2 (N12737, N12718, N85);
or OR2 (N12738, N12737, N2113);
nor NOR4 (N12739, N12735, N2182, N12681, N4000);
nor NOR4 (N12740, N12734, N622, N9789, N1565);
not NOT1 (N12741, N12738);
xor XOR2 (N12742, N12741, N6704);
or OR3 (N12743, N12740, N449, N7879);
nor NOR4 (N12744, N12730, N7788, N4945, N2229);
nand NAND3 (N12745, N12744, N3024, N369);
not NOT1 (N12746, N12729);
nor NOR4 (N12747, N12722, N6835, N10666, N1382);
and AND4 (N12748, N12743, N7578, N9526, N11663);
xor XOR2 (N12749, N12746, N576);
buf BUF1 (N12750, N12747);
nor NOR3 (N12751, N12742, N10443, N4348);
not NOT1 (N12752, N12739);
nor NOR3 (N12753, N12748, N8553, N6795);
buf BUF1 (N12754, N12732);
and AND3 (N12755, N12751, N1491, N8227);
and AND4 (N12756, N12736, N5215, N4455, N12147);
or OR3 (N12757, N12750, N9477, N10047);
nor NOR2 (N12758, N12749, N6066);
buf BUF1 (N12759, N12745);
buf BUF1 (N12760, N12727);
nand NAND2 (N12761, N12757, N11309);
and AND3 (N12762, N12755, N6949, N10075);
not NOT1 (N12763, N12760);
nor NOR2 (N12764, N12756, N9577);
or OR4 (N12765, N12752, N3666, N321, N9479);
nor NOR2 (N12766, N12701, N12273);
xor XOR2 (N12767, N12763, N5030);
xor XOR2 (N12768, N12758, N2866);
nor NOR2 (N12769, N12761, N5638);
and AND2 (N12770, N12754, N2251);
nand NAND4 (N12771, N12762, N1512, N1758, N3139);
nand NAND2 (N12772, N12766, N636);
and AND2 (N12773, N12771, N1627);
nand NAND4 (N12774, N12769, N11960, N4417, N7903);
buf BUF1 (N12775, N12764);
nor NOR2 (N12776, N12759, N3424);
nor NOR2 (N12777, N12772, N11453);
and AND3 (N12778, N12753, N9513, N10409);
and AND4 (N12779, N12777, N10709, N17, N7634);
xor XOR2 (N12780, N12765, N2278);
nand NAND4 (N12781, N12767, N7209, N666, N112);
nor NOR4 (N12782, N12773, N11597, N10584, N7340);
not NOT1 (N12783, N12782);
or OR3 (N12784, N12774, N6742, N618);
or OR4 (N12785, N12770, N7033, N6222, N9051);
nor NOR3 (N12786, N12776, N8012, N7152);
buf BUF1 (N12787, N12785);
or OR4 (N12788, N12783, N12028, N11899, N93);
and AND2 (N12789, N12780, N8255);
nand NAND3 (N12790, N12775, N2284, N5447);
not NOT1 (N12791, N12790);
xor XOR2 (N12792, N12768, N329);
xor XOR2 (N12793, N12788, N3669);
nor NOR3 (N12794, N12781, N11226, N10159);
buf BUF1 (N12795, N12784);
buf BUF1 (N12796, N12789);
or OR4 (N12797, N12794, N8547, N3881, N12365);
or OR2 (N12798, N12796, N4586);
not NOT1 (N12799, N12797);
xor XOR2 (N12800, N12793, N11457);
or OR3 (N12801, N12800, N5419, N4607);
xor XOR2 (N12802, N12779, N8297);
and AND4 (N12803, N12778, N5448, N9757, N3962);
buf BUF1 (N12804, N12787);
buf BUF1 (N12805, N12804);
or OR3 (N12806, N12805, N4278, N9921);
xor XOR2 (N12807, N12798, N11253);
not NOT1 (N12808, N12803);
nand NAND4 (N12809, N12795, N5667, N4003, N6559);
xor XOR2 (N12810, N12809, N11781);
buf BUF1 (N12811, N12799);
xor XOR2 (N12812, N12792, N4981);
or OR2 (N12813, N12812, N8360);
buf BUF1 (N12814, N12791);
not NOT1 (N12815, N12807);
not NOT1 (N12816, N12815);
or OR4 (N12817, N12814, N1516, N11640, N11473);
nor NOR3 (N12818, N12816, N10428, N1522);
or OR3 (N12819, N12806, N658, N5901);
nor NOR2 (N12820, N12813, N2941);
nor NOR2 (N12821, N12819, N9598);
not NOT1 (N12822, N12818);
nand NAND4 (N12823, N12822, N11140, N10003, N6038);
xor XOR2 (N12824, N12811, N8624);
or OR2 (N12825, N12823, N9044);
nor NOR4 (N12826, N12801, N8407, N5451, N2404);
not NOT1 (N12827, N12817);
and AND3 (N12828, N12808, N1578, N8531);
buf BUF1 (N12829, N12825);
and AND2 (N12830, N12827, N12201);
nand NAND2 (N12831, N12829, N10269);
and AND2 (N12832, N12830, N4807);
or OR3 (N12833, N12831, N5045, N1053);
buf BUF1 (N12834, N12826);
nor NOR2 (N12835, N12820, N7619);
xor XOR2 (N12836, N12821, N9150);
and AND2 (N12837, N12802, N5561);
buf BUF1 (N12838, N12832);
nor NOR2 (N12839, N12836, N4834);
or OR3 (N12840, N12834, N10078, N7558);
and AND4 (N12841, N12810, N5012, N7746, N506);
not NOT1 (N12842, N12828);
xor XOR2 (N12843, N12838, N390);
nand NAND2 (N12844, N12837, N5930);
buf BUF1 (N12845, N12824);
nor NOR2 (N12846, N12840, N7202);
not NOT1 (N12847, N12845);
nand NAND2 (N12848, N12786, N6556);
buf BUF1 (N12849, N12843);
or OR2 (N12850, N12847, N12582);
xor XOR2 (N12851, N12839, N1999);
xor XOR2 (N12852, N12846, N8826);
or OR2 (N12853, N12835, N5250);
or OR2 (N12854, N12848, N5645);
or OR2 (N12855, N12854, N2758);
or OR3 (N12856, N12844, N6744, N4498);
xor XOR2 (N12857, N12856, N8714);
and AND2 (N12858, N12850, N2418);
nor NOR2 (N12859, N12855, N10770);
xor XOR2 (N12860, N12857, N1474);
or OR2 (N12861, N12853, N613);
xor XOR2 (N12862, N12841, N9269);
nand NAND3 (N12863, N12851, N6169, N1322);
not NOT1 (N12864, N12849);
nand NAND3 (N12865, N12858, N2686, N1720);
nand NAND3 (N12866, N12860, N1126, N637);
buf BUF1 (N12867, N12862);
and AND2 (N12868, N12852, N6326);
nor NOR2 (N12869, N12833, N7081);
nor NOR2 (N12870, N12842, N246);
not NOT1 (N12871, N12863);
nand NAND4 (N12872, N12864, N7071, N5147, N10213);
buf BUF1 (N12873, N12872);
and AND4 (N12874, N12866, N6015, N5924, N187);
nor NOR4 (N12875, N12867, N4535, N8151, N156);
and AND4 (N12876, N12870, N4328, N11261, N7179);
or OR4 (N12877, N12865, N10870, N10004, N11376);
nor NOR2 (N12878, N12871, N8775);
nor NOR4 (N12879, N12859, N1806, N12507, N3300);
xor XOR2 (N12880, N12861, N5768);
xor XOR2 (N12881, N12868, N3924);
and AND3 (N12882, N12874, N2325, N9031);
nor NOR3 (N12883, N12869, N1806, N2674);
or OR2 (N12884, N12876, N11616);
xor XOR2 (N12885, N12877, N2188);
buf BUF1 (N12886, N12879);
not NOT1 (N12887, N12881);
buf BUF1 (N12888, N12880);
nand NAND4 (N12889, N12884, N2340, N6545, N12205);
buf BUF1 (N12890, N12878);
or OR4 (N12891, N12875, N2781, N4589, N12112);
buf BUF1 (N12892, N12886);
and AND2 (N12893, N12887, N5562);
nor NOR3 (N12894, N12890, N11890, N1087);
buf BUF1 (N12895, N12891);
not NOT1 (N12896, N12889);
xor XOR2 (N12897, N12895, N12126);
and AND3 (N12898, N12897, N9556, N3280);
nor NOR2 (N12899, N12882, N10300);
and AND2 (N12900, N12892, N4703);
nand NAND3 (N12901, N12885, N10184, N11753);
not NOT1 (N12902, N12893);
not NOT1 (N12903, N12898);
and AND2 (N12904, N12901, N12609);
and AND2 (N12905, N12894, N9458);
nand NAND4 (N12906, N12896, N7604, N4099, N6948);
xor XOR2 (N12907, N12888, N3779);
buf BUF1 (N12908, N12873);
nor NOR3 (N12909, N12899, N596, N468);
and AND3 (N12910, N12907, N7191, N4101);
not NOT1 (N12911, N12906);
or OR4 (N12912, N12908, N4374, N791, N9426);
or OR3 (N12913, N12909, N7182, N3770);
or OR4 (N12914, N12910, N3851, N7465, N6584);
not NOT1 (N12915, N12900);
not NOT1 (N12916, N12911);
or OR4 (N12917, N12905, N11585, N12539, N7894);
not NOT1 (N12918, N12915);
and AND2 (N12919, N12902, N11374);
and AND2 (N12920, N12914, N5194);
and AND2 (N12921, N12920, N534);
buf BUF1 (N12922, N12921);
xor XOR2 (N12923, N12916, N11088);
and AND3 (N12924, N12883, N274, N8827);
buf BUF1 (N12925, N12912);
and AND2 (N12926, N12913, N4155);
not NOT1 (N12927, N12923);
nand NAND3 (N12928, N12903, N826, N9405);
and AND2 (N12929, N12904, N1581);
xor XOR2 (N12930, N12928, N9872);
or OR4 (N12931, N12922, N11744, N10412, N2529);
and AND2 (N12932, N12931, N11153);
and AND3 (N12933, N12926, N4536, N9331);
or OR3 (N12934, N12929, N460, N5371);
or OR3 (N12935, N12919, N10450, N5676);
xor XOR2 (N12936, N12935, N1951);
buf BUF1 (N12937, N12927);
and AND4 (N12938, N12930, N11128, N2790, N2853);
buf BUF1 (N12939, N12936);
nor NOR3 (N12940, N12933, N9062, N2665);
buf BUF1 (N12941, N12918);
nor NOR4 (N12942, N12937, N6730, N4151, N6128);
or OR4 (N12943, N12934, N9607, N7364, N2955);
nor NOR4 (N12944, N12917, N6472, N10250, N4739);
nand NAND2 (N12945, N12932, N12262);
or OR3 (N12946, N12925, N8551, N5893);
and AND3 (N12947, N12942, N3168, N6456);
and AND2 (N12948, N12940, N8823);
not NOT1 (N12949, N12947);
not NOT1 (N12950, N12943);
nor NOR4 (N12951, N12938, N9401, N3129, N5090);
and AND2 (N12952, N12945, N10741);
and AND2 (N12953, N12944, N5885);
nand NAND3 (N12954, N12951, N7478, N10149);
buf BUF1 (N12955, N12939);
buf BUF1 (N12956, N12941);
nand NAND2 (N12957, N12955, N725);
nor NOR3 (N12958, N12950, N12435, N6383);
or OR4 (N12959, N12948, N7619, N5688, N8111);
nor NOR4 (N12960, N12958, N12635, N2040, N9618);
nand NAND2 (N12961, N12957, N1664);
buf BUF1 (N12962, N12956);
buf BUF1 (N12963, N12954);
xor XOR2 (N12964, N12963, N7680);
not NOT1 (N12965, N12959);
and AND3 (N12966, N12961, N7593, N7945);
or OR3 (N12967, N12966, N8455, N530);
nor NOR2 (N12968, N12949, N6060);
or OR3 (N12969, N12962, N9111, N7766);
nor NOR3 (N12970, N12967, N5164, N4724);
or OR4 (N12971, N12964, N12549, N10893, N2441);
or OR3 (N12972, N12971, N8263, N11771);
not NOT1 (N12973, N12953);
not NOT1 (N12974, N12970);
nor NOR2 (N12975, N12946, N5750);
nand NAND3 (N12976, N12974, N4298, N5062);
or OR2 (N12977, N12952, N11748);
not NOT1 (N12978, N12924);
or OR4 (N12979, N12965, N5797, N1535, N3916);
xor XOR2 (N12980, N12977, N10348);
xor XOR2 (N12981, N12976, N1523);
and AND2 (N12982, N12968, N2626);
nand NAND3 (N12983, N12973, N4008, N11369);
or OR3 (N12984, N12980, N607, N3728);
and AND3 (N12985, N12981, N10645, N11559);
or OR2 (N12986, N12960, N1027);
nor NOR4 (N12987, N12986, N5764, N4502, N9428);
nand NAND2 (N12988, N12979, N781);
nor NOR2 (N12989, N12984, N8353);
nand NAND4 (N12990, N12989, N2058, N11648, N12710);
and AND4 (N12991, N12990, N4202, N6413, N5045);
nand NAND3 (N12992, N12987, N12037, N5956);
not NOT1 (N12993, N12983);
xor XOR2 (N12994, N12992, N3519);
buf BUF1 (N12995, N12991);
buf BUF1 (N12996, N12994);
nor NOR4 (N12997, N12985, N6154, N11230, N5741);
nand NAND3 (N12998, N12969, N9548, N10109);
and AND4 (N12999, N12982, N12086, N563, N2372);
nand NAND2 (N13000, N12996, N6407);
and AND4 (N13001, N12993, N1270, N2893, N4133);
not NOT1 (N13002, N12995);
nand NAND4 (N13003, N12988, N5122, N1051, N6209);
xor XOR2 (N13004, N13002, N10950);
nor NOR4 (N13005, N12998, N3222, N12825, N6515);
and AND4 (N13006, N12997, N6293, N8306, N281);
not NOT1 (N13007, N13004);
xor XOR2 (N13008, N13006, N10478);
not NOT1 (N13009, N13001);
nor NOR2 (N13010, N12999, N4254);
xor XOR2 (N13011, N13000, N1513);
xor XOR2 (N13012, N13005, N10013);
or OR3 (N13013, N13009, N9493, N6254);
nand NAND4 (N13014, N13003, N4296, N7918, N1830);
or OR3 (N13015, N13013, N3367, N2255);
nor NOR4 (N13016, N13011, N4564, N7996, N12177);
buf BUF1 (N13017, N13008);
buf BUF1 (N13018, N12972);
or OR2 (N13019, N13007, N8487);
buf BUF1 (N13020, N13017);
buf BUF1 (N13021, N13010);
xor XOR2 (N13022, N12978, N11940);
not NOT1 (N13023, N13014);
not NOT1 (N13024, N13020);
buf BUF1 (N13025, N13016);
buf BUF1 (N13026, N13023);
buf BUF1 (N13027, N13025);
or OR3 (N13028, N13012, N6633, N1791);
not NOT1 (N13029, N13015);
and AND3 (N13030, N13021, N11654, N2407);
buf BUF1 (N13031, N13019);
nand NAND2 (N13032, N13024, N255);
not NOT1 (N13033, N13031);
nand NAND2 (N13034, N12975, N4902);
xor XOR2 (N13035, N13027, N7278);
buf BUF1 (N13036, N13022);
nor NOR4 (N13037, N13026, N4723, N9503, N6742);
xor XOR2 (N13038, N13018, N8800);
buf BUF1 (N13039, N13032);
buf BUF1 (N13040, N13033);
xor XOR2 (N13041, N13029, N12362);
not NOT1 (N13042, N13037);
not NOT1 (N13043, N13028);
and AND3 (N13044, N13035, N12423, N8719);
nand NAND3 (N13045, N13041, N12662, N178);
nand NAND3 (N13046, N13044, N11094, N429);
buf BUF1 (N13047, N13036);
xor XOR2 (N13048, N13045, N7505);
and AND2 (N13049, N13047, N2300);
not NOT1 (N13050, N13043);
nand NAND3 (N13051, N13046, N6433, N1276);
buf BUF1 (N13052, N13048);
not NOT1 (N13053, N13030);
nor NOR3 (N13054, N13038, N10775, N7236);
buf BUF1 (N13055, N13051);
not NOT1 (N13056, N13034);
nor NOR2 (N13057, N13054, N10);
nand NAND3 (N13058, N13050, N10447, N9665);
or OR4 (N13059, N13058, N9037, N8128, N2738);
xor XOR2 (N13060, N13042, N3651);
not NOT1 (N13061, N13052);
not NOT1 (N13062, N13053);
and AND4 (N13063, N13049, N10229, N4237, N6854);
and AND3 (N13064, N13063, N7265, N9388);
not NOT1 (N13065, N13060);
and AND2 (N13066, N13039, N3453);
not NOT1 (N13067, N13062);
xor XOR2 (N13068, N13065, N7812);
nor NOR3 (N13069, N13067, N10771, N4870);
xor XOR2 (N13070, N13066, N470);
or OR4 (N13071, N13057, N5110, N1020, N1741);
nand NAND3 (N13072, N13064, N3775, N1659);
not NOT1 (N13073, N13061);
nor NOR4 (N13074, N13073, N12805, N1717, N10248);
nand NAND4 (N13075, N13071, N6299, N3760, N6654);
and AND3 (N13076, N13069, N3220, N1193);
xor XOR2 (N13077, N13056, N4204);
or OR4 (N13078, N13059, N8859, N6801, N5408);
nand NAND4 (N13079, N13055, N6668, N7612, N10578);
buf BUF1 (N13080, N13074);
xor XOR2 (N13081, N13068, N8459);
buf BUF1 (N13082, N13077);
or OR2 (N13083, N13082, N5331);
xor XOR2 (N13084, N13083, N11146);
and AND2 (N13085, N13080, N11869);
nor NOR3 (N13086, N13078, N11045, N5300);
buf BUF1 (N13087, N13086);
xor XOR2 (N13088, N13072, N469);
or OR2 (N13089, N13088, N1933);
and AND4 (N13090, N13084, N7330, N9648, N12865);
nor NOR3 (N13091, N13075, N434, N3897);
buf BUF1 (N13092, N13081);
not NOT1 (N13093, N13070);
nand NAND2 (N13094, N13087, N868);
nor NOR3 (N13095, N13085, N10163, N939);
nor NOR4 (N13096, N13093, N5177, N2819, N3657);
nand NAND4 (N13097, N13095, N4813, N6990, N9000);
xor XOR2 (N13098, N13089, N2652);
or OR3 (N13099, N13096, N2290, N4664);
not NOT1 (N13100, N13099);
nor NOR4 (N13101, N13098, N5622, N8401, N2346);
or OR2 (N13102, N13079, N10040);
xor XOR2 (N13103, N13092, N5075);
and AND2 (N13104, N13102, N7960);
nor NOR2 (N13105, N13040, N6215);
not NOT1 (N13106, N13100);
nor NOR4 (N13107, N13097, N1656, N7486, N11730);
not NOT1 (N13108, N13091);
and AND4 (N13109, N13107, N5894, N11674, N9493);
nand NAND3 (N13110, N13105, N91, N207);
not NOT1 (N13111, N13106);
buf BUF1 (N13112, N13111);
not NOT1 (N13113, N13104);
and AND2 (N13114, N13094, N12483);
and AND4 (N13115, N13113, N1122, N10132, N8363);
nand NAND4 (N13116, N13076, N7994, N4989, N975);
nand NAND4 (N13117, N13108, N8090, N6810, N5342);
not NOT1 (N13118, N13116);
xor XOR2 (N13119, N13118, N7930);
or OR2 (N13120, N13112, N3958);
xor XOR2 (N13121, N13110, N1839);
buf BUF1 (N13122, N13090);
nand NAND4 (N13123, N13122, N425, N8512, N12775);
buf BUF1 (N13124, N13123);
nand NAND4 (N13125, N13101, N9417, N12698, N1307);
not NOT1 (N13126, N13124);
not NOT1 (N13127, N13125);
buf BUF1 (N13128, N13103);
nand NAND2 (N13129, N13115, N13045);
or OR2 (N13130, N13109, N5468);
or OR2 (N13131, N13117, N5790);
buf BUF1 (N13132, N13128);
and AND4 (N13133, N13119, N159, N12033, N12524);
nor NOR2 (N13134, N13121, N12712);
nand NAND2 (N13135, N13134, N8870);
not NOT1 (N13136, N13120);
and AND4 (N13137, N13130, N4849, N5852, N4906);
and AND3 (N13138, N13129, N1595, N1110);
not NOT1 (N13139, N13133);
or OR2 (N13140, N13132, N6343);
not NOT1 (N13141, N13114);
buf BUF1 (N13142, N13126);
and AND4 (N13143, N13140, N6929, N7471, N6209);
nand NAND2 (N13144, N13136, N13010);
or OR4 (N13145, N13143, N9416, N5711, N282);
nand NAND2 (N13146, N13141, N13109);
buf BUF1 (N13147, N13127);
or OR3 (N13148, N13147, N1554, N11775);
nand NAND3 (N13149, N13131, N8056, N4523);
or OR3 (N13150, N13142, N11720, N11507);
and AND2 (N13151, N13144, N5786);
buf BUF1 (N13152, N13137);
buf BUF1 (N13153, N13151);
buf BUF1 (N13154, N13138);
nor NOR4 (N13155, N13152, N4396, N12735, N11258);
or OR4 (N13156, N13135, N8419, N2713, N3527);
or OR2 (N13157, N13139, N5996);
and AND2 (N13158, N13155, N965);
nand NAND3 (N13159, N13148, N1519, N7566);
or OR2 (N13160, N13156, N6058);
or OR4 (N13161, N13153, N2370, N12521, N11888);
xor XOR2 (N13162, N13161, N6729);
xor XOR2 (N13163, N13160, N12767);
not NOT1 (N13164, N13158);
nand NAND3 (N13165, N13164, N2883, N9282);
not NOT1 (N13166, N13145);
nor NOR2 (N13167, N13149, N5504);
xor XOR2 (N13168, N13150, N6699);
nor NOR2 (N13169, N13167, N4255);
buf BUF1 (N13170, N13162);
nor NOR4 (N13171, N13146, N12818, N2211, N10477);
nor NOR3 (N13172, N13170, N3991, N4698);
nor NOR3 (N13173, N13159, N11848, N6831);
and AND4 (N13174, N13163, N8447, N5362, N5603);
not NOT1 (N13175, N13169);
nor NOR4 (N13176, N13175, N8905, N11727, N11807);
nand NAND3 (N13177, N13176, N12284, N5952);
and AND2 (N13178, N13174, N12426);
nand NAND4 (N13179, N13171, N8325, N5912, N3312);
or OR4 (N13180, N13154, N5877, N6355, N10123);
buf BUF1 (N13181, N13179);
buf BUF1 (N13182, N13157);
xor XOR2 (N13183, N13181, N7253);
buf BUF1 (N13184, N13166);
nor NOR3 (N13185, N13178, N9773, N12306);
not NOT1 (N13186, N13180);
nor NOR2 (N13187, N13185, N7438);
not NOT1 (N13188, N13165);
not NOT1 (N13189, N13188);
xor XOR2 (N13190, N13168, N5809);
nand NAND2 (N13191, N13186, N6688);
xor XOR2 (N13192, N13183, N7636);
xor XOR2 (N13193, N13191, N9763);
buf BUF1 (N13194, N13173);
nand NAND4 (N13195, N13189, N2141, N11356, N9291);
xor XOR2 (N13196, N13192, N3688);
buf BUF1 (N13197, N13193);
nand NAND3 (N13198, N13177, N2280, N7339);
or OR2 (N13199, N13198, N5642);
not NOT1 (N13200, N13187);
nor NOR3 (N13201, N13190, N9166, N4000);
buf BUF1 (N13202, N13197);
buf BUF1 (N13203, N13202);
nand NAND4 (N13204, N13203, N7637, N1450, N4490);
buf BUF1 (N13205, N13200);
nor NOR3 (N13206, N13196, N4836, N3174);
or OR4 (N13207, N13205, N8802, N12326, N2323);
buf BUF1 (N13208, N13206);
buf BUF1 (N13209, N13194);
nor NOR2 (N13210, N13207, N3494);
not NOT1 (N13211, N13172);
xor XOR2 (N13212, N13204, N8458);
buf BUF1 (N13213, N13211);
xor XOR2 (N13214, N13195, N12448);
nand NAND2 (N13215, N13184, N3482);
not NOT1 (N13216, N13213);
xor XOR2 (N13217, N13212, N5069);
nand NAND2 (N13218, N13210, N11781);
and AND2 (N13219, N13214, N9505);
not NOT1 (N13220, N13199);
nand NAND4 (N13221, N13201, N6000, N8880, N646);
or OR4 (N13222, N13217, N8595, N11468, N2811);
buf BUF1 (N13223, N13220);
not NOT1 (N13224, N13219);
nand NAND2 (N13225, N13209, N1819);
nor NOR2 (N13226, N13182, N5050);
xor XOR2 (N13227, N13216, N12634);
buf BUF1 (N13228, N13227);
buf BUF1 (N13229, N13218);
buf BUF1 (N13230, N13229);
nand NAND2 (N13231, N13215, N12436);
and AND2 (N13232, N13224, N7393);
not NOT1 (N13233, N13226);
nor NOR2 (N13234, N13223, N4254);
or OR4 (N13235, N13221, N2791, N4898, N2530);
buf BUF1 (N13236, N13231);
nor NOR4 (N13237, N13228, N998, N2890, N9535);
buf BUF1 (N13238, N13235);
nand NAND4 (N13239, N13234, N1437, N2986, N8218);
nand NAND4 (N13240, N13233, N1933, N11030, N4250);
buf BUF1 (N13241, N13232);
not NOT1 (N13242, N13222);
and AND3 (N13243, N13225, N10151, N6578);
nand NAND3 (N13244, N13230, N5999, N8352);
nand NAND4 (N13245, N13241, N6871, N12446, N12918);
nand NAND3 (N13246, N13237, N9645, N6827);
nand NAND3 (N13247, N13236, N4332, N2862);
or OR2 (N13248, N13247, N9715);
buf BUF1 (N13249, N13239);
buf BUF1 (N13250, N13240);
nor NOR4 (N13251, N13244, N11112, N6395, N8596);
not NOT1 (N13252, N13242);
nand NAND2 (N13253, N13246, N7067);
buf BUF1 (N13254, N13249);
not NOT1 (N13255, N13250);
xor XOR2 (N13256, N13251, N3267);
or OR3 (N13257, N13248, N10227, N6884);
and AND4 (N13258, N13256, N4554, N9123, N1792);
nand NAND4 (N13259, N13253, N193, N12016, N8815);
nor NOR4 (N13260, N13255, N6159, N11054, N1843);
nor NOR2 (N13261, N13245, N12037);
buf BUF1 (N13262, N13260);
nand NAND3 (N13263, N13262, N2565, N2729);
buf BUF1 (N13264, N13261);
not NOT1 (N13265, N13208);
or OR3 (N13266, N13258, N9446, N2426);
buf BUF1 (N13267, N13254);
or OR2 (N13268, N13267, N5209);
nand NAND2 (N13269, N13238, N5607);
or OR4 (N13270, N13264, N12589, N10838, N5595);
buf BUF1 (N13271, N13263);
not NOT1 (N13272, N13259);
nor NOR2 (N13273, N13272, N10709);
buf BUF1 (N13274, N13271);
not NOT1 (N13275, N13269);
not NOT1 (N13276, N13257);
nand NAND3 (N13277, N13273, N3622, N6875);
not NOT1 (N13278, N13275);
nand NAND4 (N13279, N13268, N5806, N12651, N2146);
not NOT1 (N13280, N13276);
and AND3 (N13281, N13266, N9734, N12592);
and AND2 (N13282, N13280, N2319);
and AND4 (N13283, N13279, N7923, N11443, N8321);
buf BUF1 (N13284, N13274);
nor NOR4 (N13285, N13281, N6993, N10034, N1848);
or OR2 (N13286, N13285, N1492);
or OR3 (N13287, N13282, N717, N2398);
not NOT1 (N13288, N13270);
or OR2 (N13289, N13278, N2417);
nand NAND2 (N13290, N13287, N3270);
xor XOR2 (N13291, N13286, N1741);
buf BUF1 (N13292, N13289);
xor XOR2 (N13293, N13252, N2439);
or OR3 (N13294, N13292, N11284, N7881);
buf BUF1 (N13295, N13290);
xor XOR2 (N13296, N13293, N508);
xor XOR2 (N13297, N13284, N616);
nor NOR4 (N13298, N13243, N8244, N4169, N6839);
and AND3 (N13299, N13295, N7874, N8089);
xor XOR2 (N13300, N13297, N12503);
nor NOR3 (N13301, N13299, N11473, N3519);
buf BUF1 (N13302, N13277);
nand NAND2 (N13303, N13265, N11221);
not NOT1 (N13304, N13302);
and AND4 (N13305, N13298, N11452, N10216, N111);
nand NAND3 (N13306, N13294, N400, N5960);
buf BUF1 (N13307, N13296);
buf BUF1 (N13308, N13300);
xor XOR2 (N13309, N13308, N1188);
or OR4 (N13310, N13305, N7249, N5541, N537);
or OR4 (N13311, N13291, N254, N12343, N10925);
not NOT1 (N13312, N13310);
xor XOR2 (N13313, N13309, N4928);
nor NOR2 (N13314, N13313, N10278);
or OR2 (N13315, N13306, N3384);
and AND3 (N13316, N13315, N6925, N692);
and AND2 (N13317, N13314, N9555);
nand NAND2 (N13318, N13317, N12183);
and AND4 (N13319, N13318, N2083, N4709, N3600);
nor NOR4 (N13320, N13303, N11265, N7121, N11321);
and AND4 (N13321, N13288, N3390, N5507, N6538);
and AND2 (N13322, N13319, N3591);
nor NOR3 (N13323, N13311, N13034, N10363);
or OR3 (N13324, N13307, N8021, N3310);
or OR3 (N13325, N13283, N6504, N11206);
or OR3 (N13326, N13320, N1668, N2250);
or OR2 (N13327, N13322, N8082);
nand NAND3 (N13328, N13325, N11038, N10683);
and AND4 (N13329, N13324, N9125, N8883, N5504);
and AND4 (N13330, N13327, N4618, N9500, N834);
buf BUF1 (N13331, N13312);
not NOT1 (N13332, N13326);
or OR4 (N13333, N13329, N13230, N2642, N11090);
not NOT1 (N13334, N13304);
or OR2 (N13335, N13333, N8966);
and AND3 (N13336, N13321, N4711, N6769);
nor NOR4 (N13337, N13330, N9015, N1228, N4820);
nor NOR2 (N13338, N13323, N7032);
xor XOR2 (N13339, N13335, N11902);
buf BUF1 (N13340, N13338);
and AND2 (N13341, N13316, N9356);
buf BUF1 (N13342, N13340);
and AND3 (N13343, N13301, N11401, N1076);
xor XOR2 (N13344, N13343, N5697);
nand NAND2 (N13345, N13334, N8633);
nor NOR2 (N13346, N13331, N10937);
xor XOR2 (N13347, N13328, N8906);
xor XOR2 (N13348, N13332, N8062);
or OR3 (N13349, N13345, N4890, N12473);
not NOT1 (N13350, N13344);
and AND3 (N13351, N13347, N10956, N6121);
nor NOR4 (N13352, N13350, N5706, N13188, N3225);
not NOT1 (N13353, N13342);
buf BUF1 (N13354, N13351);
nand NAND3 (N13355, N13346, N9896, N1045);
and AND3 (N13356, N13336, N9071, N2246);
and AND2 (N13357, N13355, N9212);
nand NAND4 (N13358, N13339, N10500, N6528, N225);
nand NAND2 (N13359, N13349, N9716);
not NOT1 (N13360, N13354);
nand NAND3 (N13361, N13337, N8719, N7015);
nand NAND4 (N13362, N13348, N3974, N7827, N310);
not NOT1 (N13363, N13352);
not NOT1 (N13364, N13362);
nand NAND3 (N13365, N13360, N1651, N3039);
buf BUF1 (N13366, N13358);
nor NOR2 (N13367, N13341, N4512);
or OR2 (N13368, N13364, N8970);
and AND3 (N13369, N13353, N1509, N5163);
not NOT1 (N13370, N13363);
and AND4 (N13371, N13366, N8564, N6707, N10146);
not NOT1 (N13372, N13365);
buf BUF1 (N13373, N13372);
nand NAND3 (N13374, N13359, N4356, N5775);
nand NAND3 (N13375, N13371, N9095, N8059);
or OR2 (N13376, N13368, N11193);
and AND3 (N13377, N13367, N7409, N311);
nand NAND2 (N13378, N13376, N6569);
and AND2 (N13379, N13356, N12858);
nor NOR3 (N13380, N13361, N11183, N1996);
buf BUF1 (N13381, N13357);
or OR2 (N13382, N13377, N7088);
buf BUF1 (N13383, N13378);
nor NOR3 (N13384, N13383, N5014, N8475);
not NOT1 (N13385, N13369);
xor XOR2 (N13386, N13375, N9492);
nor NOR2 (N13387, N13381, N3407);
nand NAND3 (N13388, N13384, N2787, N5153);
buf BUF1 (N13389, N13388);
or OR2 (N13390, N13370, N515);
nand NAND2 (N13391, N13382, N12610);
buf BUF1 (N13392, N13385);
buf BUF1 (N13393, N13380);
and AND2 (N13394, N13374, N2087);
or OR2 (N13395, N13390, N693);
nand NAND2 (N13396, N13379, N9750);
nand NAND2 (N13397, N13396, N8);
buf BUF1 (N13398, N13389);
and AND4 (N13399, N13397, N4749, N888, N3275);
buf BUF1 (N13400, N13393);
nor NOR4 (N13401, N13400, N12422, N8563, N6754);
nand NAND2 (N13402, N13386, N7955);
nand NAND4 (N13403, N13392, N172, N8659, N61);
nor NOR4 (N13404, N13399, N12304, N1607, N6885);
not NOT1 (N13405, N13373);
not NOT1 (N13406, N13404);
buf BUF1 (N13407, N13406);
buf BUF1 (N13408, N13387);
and AND3 (N13409, N13403, N13260, N7440);
and AND4 (N13410, N13394, N4648, N6691, N4173);
nand NAND2 (N13411, N13409, N12678);
xor XOR2 (N13412, N13402, N11955);
not NOT1 (N13413, N13395);
nand NAND3 (N13414, N13410, N7527, N1871);
or OR4 (N13415, N13391, N8074, N12, N8961);
nand NAND3 (N13416, N13408, N9306, N5920);
xor XOR2 (N13417, N13407, N7237);
and AND4 (N13418, N13412, N4159, N11381, N10377);
or OR4 (N13419, N13405, N5134, N10917, N2693);
nand NAND4 (N13420, N13417, N5845, N3692, N6767);
nand NAND3 (N13421, N13419, N3578, N806);
or OR4 (N13422, N13411, N12255, N10621, N10272);
buf BUF1 (N13423, N13414);
buf BUF1 (N13424, N13420);
nor NOR3 (N13425, N13415, N581, N13418);
nor NOR2 (N13426, N5748, N13131);
nand NAND2 (N13427, N13426, N11381);
buf BUF1 (N13428, N13421);
or OR4 (N13429, N13413, N6297, N6628, N10768);
nand NAND2 (N13430, N13425, N773);
nand NAND4 (N13431, N13429, N4324, N2336, N8452);
or OR3 (N13432, N13431, N7051, N2628);
and AND2 (N13433, N13401, N1695);
not NOT1 (N13434, N13423);
nand NAND4 (N13435, N13427, N8309, N6647, N3723);
xor XOR2 (N13436, N13422, N2087);
not NOT1 (N13437, N13398);
not NOT1 (N13438, N13424);
buf BUF1 (N13439, N13438);
or OR3 (N13440, N13432, N1868, N1206);
or OR2 (N13441, N13430, N10927);
buf BUF1 (N13442, N13440);
and AND4 (N13443, N13437, N7519, N7521, N510);
not NOT1 (N13444, N13436);
nand NAND3 (N13445, N13443, N5776, N338);
and AND4 (N13446, N13442, N9845, N8125, N6128);
not NOT1 (N13447, N13416);
nand NAND4 (N13448, N13447, N3828, N5591, N6612);
nor NOR4 (N13449, N13445, N3709, N4618, N3751);
and AND3 (N13450, N13433, N5723, N8190);
xor XOR2 (N13451, N13444, N3631);
buf BUF1 (N13452, N13435);
or OR4 (N13453, N13451, N1527, N2614, N7024);
nand NAND3 (N13454, N13441, N2966, N7166);
xor XOR2 (N13455, N13450, N9830);
or OR2 (N13456, N13446, N4404);
xor XOR2 (N13457, N13456, N6301);
not NOT1 (N13458, N13434);
and AND3 (N13459, N13454, N11631, N3328);
not NOT1 (N13460, N13457);
nor NOR2 (N13461, N13459, N11610);
or OR4 (N13462, N13448, N11399, N8534, N10271);
xor XOR2 (N13463, N13460, N9974);
not NOT1 (N13464, N13453);
and AND3 (N13465, N13455, N141, N4754);
xor XOR2 (N13466, N13452, N2834);
or OR3 (N13467, N13462, N4940, N3847);
and AND2 (N13468, N13439, N10980);
xor XOR2 (N13469, N13468, N8198);
and AND4 (N13470, N13469, N10576, N722, N12128);
or OR3 (N13471, N13449, N12809, N7665);
xor XOR2 (N13472, N13465, N1991);
buf BUF1 (N13473, N13470);
nand NAND2 (N13474, N13466, N5692);
nor NOR4 (N13475, N13467, N10840, N3746, N286);
and AND2 (N13476, N13458, N3233);
nand NAND3 (N13477, N13474, N6405, N8505);
and AND4 (N13478, N13464, N1451, N2050, N8883);
buf BUF1 (N13479, N13463);
buf BUF1 (N13480, N13471);
and AND3 (N13481, N13480, N3576, N564);
or OR3 (N13482, N13478, N8883, N4704);
not NOT1 (N13483, N13479);
not NOT1 (N13484, N13428);
nor NOR2 (N13485, N13475, N3162);
or OR4 (N13486, N13483, N5700, N11317, N5401);
and AND2 (N13487, N13477, N13306);
buf BUF1 (N13488, N13486);
nand NAND2 (N13489, N13481, N2960);
or OR3 (N13490, N13482, N11439, N10216);
and AND4 (N13491, N13476, N1585, N3721, N4185);
not NOT1 (N13492, N13488);
nor NOR2 (N13493, N13487, N1711);
buf BUF1 (N13494, N13492);
not NOT1 (N13495, N13472);
and AND4 (N13496, N13495, N614, N5228, N7003);
not NOT1 (N13497, N13494);
nand NAND4 (N13498, N13497, N10758, N11280, N4916);
nor NOR4 (N13499, N13491, N8817, N6103, N2165);
not NOT1 (N13500, N13489);
nor NOR2 (N13501, N13498, N1082);
nor NOR3 (N13502, N13500, N6844, N947);
or OR2 (N13503, N13461, N12454);
and AND3 (N13504, N13493, N8241, N4648);
and AND2 (N13505, N13490, N7717);
buf BUF1 (N13506, N13504);
nand NAND2 (N13507, N13503, N9505);
or OR3 (N13508, N13484, N2543, N12116);
nand NAND4 (N13509, N13506, N12282, N4360, N8195);
or OR3 (N13510, N13509, N4473, N4458);
and AND2 (N13511, N13510, N10422);
not NOT1 (N13512, N13496);
xor XOR2 (N13513, N13499, N5645);
xor XOR2 (N13514, N13513, N3150);
not NOT1 (N13515, N13502);
nor NOR3 (N13516, N13507, N13189, N2029);
buf BUF1 (N13517, N13511);
or OR2 (N13518, N13485, N8993);
nor NOR4 (N13519, N13516, N6306, N12298, N7247);
buf BUF1 (N13520, N13512);
buf BUF1 (N13521, N13473);
xor XOR2 (N13522, N13508, N11090);
or OR3 (N13523, N13514, N2077, N8868);
buf BUF1 (N13524, N13515);
or OR3 (N13525, N13522, N2988, N956);
not NOT1 (N13526, N13521);
and AND2 (N13527, N13519, N12656);
xor XOR2 (N13528, N13523, N8128);
nand NAND4 (N13529, N13518, N2133, N12881, N5383);
not NOT1 (N13530, N13529);
and AND3 (N13531, N13526, N11621, N3534);
nor NOR3 (N13532, N13525, N6175, N4668);
not NOT1 (N13533, N13520);
buf BUF1 (N13534, N13517);
nor NOR3 (N13535, N13505, N10036, N1257);
and AND2 (N13536, N13501, N2614);
or OR4 (N13537, N13527, N13227, N5760, N12890);
buf BUF1 (N13538, N13530);
nor NOR3 (N13539, N13535, N12725, N7300);
not NOT1 (N13540, N13539);
buf BUF1 (N13541, N13534);
nand NAND2 (N13542, N13533, N7998);
nand NAND2 (N13543, N13541, N13253);
buf BUF1 (N13544, N13540);
xor XOR2 (N13545, N13531, N7354);
not NOT1 (N13546, N13538);
nor NOR2 (N13547, N13524, N7572);
buf BUF1 (N13548, N13543);
nor NOR2 (N13549, N13532, N6722);
or OR2 (N13550, N13546, N914);
nor NOR4 (N13551, N13536, N3678, N3854, N1667);
and AND4 (N13552, N13544, N7226, N5835, N13232);
nor NOR4 (N13553, N13550, N11707, N3503, N2366);
xor XOR2 (N13554, N13542, N6125);
not NOT1 (N13555, N13547);
and AND2 (N13556, N13552, N5171);
buf BUF1 (N13557, N13549);
xor XOR2 (N13558, N13537, N3477);
xor XOR2 (N13559, N13557, N7490);
nor NOR3 (N13560, N13559, N3735, N1167);
buf BUF1 (N13561, N13554);
nor NOR3 (N13562, N13545, N1674, N7733);
nor NOR4 (N13563, N13553, N7790, N3796, N9406);
buf BUF1 (N13564, N13562);
nand NAND4 (N13565, N13555, N1007, N2900, N8551);
nand NAND2 (N13566, N13563, N2188);
nand NAND4 (N13567, N13551, N7677, N1984, N9349);
or OR3 (N13568, N13567, N1345, N11309);
nor NOR4 (N13569, N13560, N10548, N9334, N8198);
and AND2 (N13570, N13548, N12895);
nor NOR3 (N13571, N13561, N2119, N4631);
or OR4 (N13572, N13556, N2851, N12336, N7725);
nor NOR4 (N13573, N13568, N3148, N2914, N7680);
not NOT1 (N13574, N13573);
xor XOR2 (N13575, N13571, N2766);
xor XOR2 (N13576, N13572, N8757);
not NOT1 (N13577, N13574);
nor NOR2 (N13578, N13570, N3240);
xor XOR2 (N13579, N13565, N5254);
or OR3 (N13580, N13569, N102, N9947);
nand NAND2 (N13581, N13528, N12260);
or OR2 (N13582, N13581, N12780);
or OR4 (N13583, N13579, N1233, N9704, N322);
or OR2 (N13584, N13566, N13366);
buf BUF1 (N13585, N13578);
nor NOR3 (N13586, N13576, N8867, N7931);
nor NOR2 (N13587, N13580, N9741);
or OR3 (N13588, N13586, N12748, N13423);
and AND3 (N13589, N13583, N8468, N3988);
or OR4 (N13590, N13584, N3690, N8878, N6790);
and AND3 (N13591, N13577, N6426, N11244);
or OR4 (N13592, N13558, N2864, N1164, N3422);
or OR3 (N13593, N13590, N12271, N9958);
and AND4 (N13594, N13575, N3610, N3924, N801);
nand NAND3 (N13595, N13587, N4384, N9545);
and AND2 (N13596, N13592, N12075);
nor NOR2 (N13597, N13582, N8913);
or OR3 (N13598, N13593, N10132, N6335);
buf BUF1 (N13599, N13598);
and AND3 (N13600, N13591, N2253, N13455);
not NOT1 (N13601, N13599);
or OR2 (N13602, N13589, N6535);
nand NAND2 (N13603, N13597, N9297);
nand NAND3 (N13604, N13588, N2243, N11878);
nand NAND2 (N13605, N13603, N8616);
not NOT1 (N13606, N13594);
and AND2 (N13607, N13595, N6721);
nand NAND2 (N13608, N13605, N6637);
buf BUF1 (N13609, N13607);
or OR4 (N13610, N13600, N4134, N4489, N4915);
or OR3 (N13611, N13610, N8592, N6512);
nand NAND4 (N13612, N13585, N48, N11393, N4712);
and AND3 (N13613, N13564, N5672, N3428);
not NOT1 (N13614, N13596);
or OR4 (N13615, N13614, N2463, N9415, N5737);
buf BUF1 (N13616, N13609);
xor XOR2 (N13617, N13608, N11592);
or OR3 (N13618, N13613, N10506, N7556);
xor XOR2 (N13619, N13601, N7540);
or OR2 (N13620, N13606, N606);
nand NAND3 (N13621, N13618, N3205, N1741);
nand NAND4 (N13622, N13617, N4548, N13209, N7709);
and AND2 (N13623, N13616, N3756);
and AND3 (N13624, N13623, N4641, N5990);
or OR2 (N13625, N13620, N5317);
xor XOR2 (N13626, N13611, N13073);
nor NOR2 (N13627, N13624, N5915);
and AND3 (N13628, N13625, N9910, N11329);
or OR3 (N13629, N13615, N809, N4586);
xor XOR2 (N13630, N13612, N7613);
xor XOR2 (N13631, N13629, N12035);
or OR3 (N13632, N13602, N12142, N11882);
not NOT1 (N13633, N13630);
nand NAND3 (N13634, N13621, N13052, N356);
and AND3 (N13635, N13622, N2451, N7423);
not NOT1 (N13636, N13619);
and AND2 (N13637, N13626, N9343);
and AND2 (N13638, N13627, N2701);
not NOT1 (N13639, N13635);
nand NAND3 (N13640, N13632, N5056, N9068);
nand NAND3 (N13641, N13604, N9161, N9115);
or OR2 (N13642, N13641, N7842);
xor XOR2 (N13643, N13628, N6477);
nand NAND2 (N13644, N13638, N13626);
and AND4 (N13645, N13637, N2931, N9940, N7380);
not NOT1 (N13646, N13639);
xor XOR2 (N13647, N13631, N2914);
nor NOR2 (N13648, N13645, N2690);
nand NAND4 (N13649, N13643, N11101, N13174, N2969);
and AND3 (N13650, N13640, N10368, N983);
buf BUF1 (N13651, N13644);
nand NAND2 (N13652, N13636, N7250);
buf BUF1 (N13653, N13634);
not NOT1 (N13654, N13653);
or OR2 (N13655, N13651, N6726);
nor NOR4 (N13656, N13650, N8450, N8455, N3361);
and AND2 (N13657, N13642, N12215);
nand NAND3 (N13658, N13648, N4711, N6892);
nand NAND4 (N13659, N13655, N6248, N7114, N12616);
nand NAND2 (N13660, N13652, N6123);
nor NOR3 (N13661, N13649, N2089, N9646);
xor XOR2 (N13662, N13661, N1539);
buf BUF1 (N13663, N13633);
nand NAND3 (N13664, N13654, N13659, N12096);
xor XOR2 (N13665, N7481, N12659);
buf BUF1 (N13666, N13646);
not NOT1 (N13667, N13664);
and AND3 (N13668, N13656, N6404, N3664);
and AND2 (N13669, N13662, N4638);
xor XOR2 (N13670, N13668, N11486);
not NOT1 (N13671, N13669);
not NOT1 (N13672, N13657);
not NOT1 (N13673, N13667);
xor XOR2 (N13674, N13672, N12135);
or OR4 (N13675, N13663, N10936, N3331, N9910);
or OR4 (N13676, N13671, N10695, N11774, N342);
nand NAND4 (N13677, N13675, N7575, N2555, N7069);
not NOT1 (N13678, N13658);
xor XOR2 (N13679, N13677, N12729);
xor XOR2 (N13680, N13665, N7202);
not NOT1 (N13681, N13673);
nor NOR4 (N13682, N13660, N11539, N6278, N13019);
buf BUF1 (N13683, N13676);
not NOT1 (N13684, N13683);
nand NAND3 (N13685, N13680, N10079, N13179);
and AND3 (N13686, N13666, N5375, N12103);
not NOT1 (N13687, N13686);
nor NOR4 (N13688, N13678, N3479, N12907, N3777);
not NOT1 (N13689, N13688);
or OR2 (N13690, N13684, N1373);
or OR4 (N13691, N13647, N887, N11259, N2791);
and AND2 (N13692, N13679, N6468);
and AND4 (N13693, N13681, N83, N6270, N10847);
not NOT1 (N13694, N13691);
nor NOR3 (N13695, N13690, N11716, N10693);
not NOT1 (N13696, N13695);
and AND3 (N13697, N13692, N8575, N1448);
xor XOR2 (N13698, N13689, N1771);
not NOT1 (N13699, N13693);
buf BUF1 (N13700, N13682);
and AND3 (N13701, N13700, N4725, N10502);
and AND2 (N13702, N13687, N6194);
nor NOR4 (N13703, N13674, N5085, N7697, N3032);
buf BUF1 (N13704, N13702);
buf BUF1 (N13705, N13685);
nor NOR2 (N13706, N13703, N6527);
and AND4 (N13707, N13698, N10674, N1249, N954);
not NOT1 (N13708, N13670);
nand NAND2 (N13709, N13696, N730);
and AND3 (N13710, N13699, N164, N6439);
or OR2 (N13711, N13708, N736);
xor XOR2 (N13712, N13710, N7493);
nor NOR4 (N13713, N13707, N3339, N12964, N12459);
xor XOR2 (N13714, N13709, N13707);
or OR4 (N13715, N13712, N6049, N13123, N6907);
not NOT1 (N13716, N13714);
nand NAND4 (N13717, N13704, N12177, N3669, N12067);
and AND4 (N13718, N13717, N5300, N8763, N8827);
or OR4 (N13719, N13715, N4465, N301, N13583);
and AND4 (N13720, N13716, N4012, N2162, N515);
not NOT1 (N13721, N13713);
not NOT1 (N13722, N13718);
nor NOR3 (N13723, N13705, N7911, N1799);
nand NAND4 (N13724, N13722, N6705, N5996, N8649);
buf BUF1 (N13725, N13724);
not NOT1 (N13726, N13723);
nand NAND3 (N13727, N13701, N7634, N11837);
not NOT1 (N13728, N13726);
nand NAND4 (N13729, N13711, N3125, N7250, N11096);
buf BUF1 (N13730, N13719);
and AND2 (N13731, N13721, N3549);
or OR3 (N13732, N13694, N8693, N9276);
nand NAND2 (N13733, N13720, N5290);
or OR3 (N13734, N13697, N12855, N11445);
nor NOR4 (N13735, N13727, N1490, N11849, N5353);
nand NAND3 (N13736, N13730, N10888, N7004);
buf BUF1 (N13737, N13731);
and AND2 (N13738, N13737, N7590);
or OR4 (N13739, N13734, N9747, N7962, N3759);
or OR4 (N13740, N13736, N13152, N3887, N11773);
or OR2 (N13741, N13740, N11749);
nand NAND3 (N13742, N13728, N3035, N623);
nand NAND2 (N13743, N13738, N3181);
xor XOR2 (N13744, N13742, N8307);
nand NAND2 (N13745, N13725, N3179);
nor NOR2 (N13746, N13739, N12394);
not NOT1 (N13747, N13745);
buf BUF1 (N13748, N13747);
nor NOR4 (N13749, N13746, N2271, N6509, N11152);
and AND2 (N13750, N13732, N1226);
nand NAND2 (N13751, N13729, N11785);
or OR2 (N13752, N13748, N4464);
nand NAND4 (N13753, N13733, N11586, N10887, N9813);
nor NOR3 (N13754, N13735, N6049, N10589);
or OR2 (N13755, N13744, N9487);
xor XOR2 (N13756, N13706, N8511);
nand NAND3 (N13757, N13755, N13079, N6463);
and AND2 (N13758, N13754, N3402);
buf BUF1 (N13759, N13750);
or OR2 (N13760, N13749, N11538);
nor NOR3 (N13761, N13753, N4334, N9754);
buf BUF1 (N13762, N13759);
buf BUF1 (N13763, N13757);
nor NOR3 (N13764, N13751, N6825, N12401);
or OR2 (N13765, N13763, N13040);
or OR2 (N13766, N13756, N5262);
nand NAND4 (N13767, N13741, N2433, N11710, N4020);
xor XOR2 (N13768, N13743, N3328);
not NOT1 (N13769, N13761);
xor XOR2 (N13770, N13764, N667);
or OR2 (N13771, N13758, N11449);
and AND3 (N13772, N13770, N6234, N11756);
or OR2 (N13773, N13752, N13330);
xor XOR2 (N13774, N13762, N3486);
nand NAND3 (N13775, N13774, N5455, N4046);
buf BUF1 (N13776, N13767);
not NOT1 (N13777, N13769);
not NOT1 (N13778, N13766);
buf BUF1 (N13779, N13765);
nand NAND4 (N13780, N13778, N11583, N10352, N4722);
nor NOR3 (N13781, N13771, N450, N12068);
and AND4 (N13782, N13780, N9995, N8188, N10940);
buf BUF1 (N13783, N13775);
xor XOR2 (N13784, N13760, N4322);
buf BUF1 (N13785, N13784);
xor XOR2 (N13786, N13783, N4277);
xor XOR2 (N13787, N13777, N6567);
and AND4 (N13788, N13776, N8177, N5891, N4671);
not NOT1 (N13789, N13772);
nand NAND4 (N13790, N13773, N705, N1556, N12510);
xor XOR2 (N13791, N13789, N1888);
not NOT1 (N13792, N13790);
xor XOR2 (N13793, N13768, N11516);
nor NOR4 (N13794, N13787, N235, N1013, N269);
buf BUF1 (N13795, N13792);
nor NOR2 (N13796, N13794, N343);
xor XOR2 (N13797, N13785, N12580);
or OR2 (N13798, N13791, N7855);
nand NAND3 (N13799, N13793, N5570, N7029);
nor NOR2 (N13800, N13782, N2556);
and AND3 (N13801, N13799, N12745, N2194);
and AND3 (N13802, N13796, N9410, N1628);
not NOT1 (N13803, N13788);
not NOT1 (N13804, N13779);
buf BUF1 (N13805, N13800);
or OR2 (N13806, N13786, N2527);
and AND3 (N13807, N13802, N13439, N2376);
not NOT1 (N13808, N13806);
xor XOR2 (N13809, N13804, N9937);
nor NOR3 (N13810, N13797, N8758, N13612);
or OR3 (N13811, N13805, N88, N817);
or OR3 (N13812, N13811, N786, N8537);
nor NOR4 (N13813, N13801, N2879, N8958, N11450);
xor XOR2 (N13814, N13807, N2041);
nor NOR4 (N13815, N13798, N8232, N3484, N2879);
nor NOR3 (N13816, N13803, N10610, N570);
and AND3 (N13817, N13815, N2286, N2759);
buf BUF1 (N13818, N13809);
and AND4 (N13819, N13808, N8, N13649, N11899);
not NOT1 (N13820, N13795);
xor XOR2 (N13821, N13812, N8597);
xor XOR2 (N13822, N13821, N3634);
xor XOR2 (N13823, N13813, N8755);
and AND2 (N13824, N13810, N8539);
and AND2 (N13825, N13819, N2115);
nor NOR3 (N13826, N13824, N12846, N4292);
nand NAND2 (N13827, N13825, N8962);
buf BUF1 (N13828, N13822);
and AND4 (N13829, N13817, N10367, N9037, N6313);
or OR3 (N13830, N13814, N11179, N8703);
buf BUF1 (N13831, N13816);
or OR4 (N13832, N13828, N11541, N4922, N12226);
not NOT1 (N13833, N13832);
buf BUF1 (N13834, N13826);
or OR3 (N13835, N13827, N9034, N10940);
not NOT1 (N13836, N13831);
and AND4 (N13837, N13818, N12590, N13570, N3476);
buf BUF1 (N13838, N13820);
or OR4 (N13839, N13833, N1734, N4608, N268);
nor NOR3 (N13840, N13836, N4038, N5834);
buf BUF1 (N13841, N13829);
xor XOR2 (N13842, N13830, N4721);
xor XOR2 (N13843, N13839, N11112);
or OR3 (N13844, N13838, N1288, N10600);
buf BUF1 (N13845, N13835);
buf BUF1 (N13846, N13837);
nand NAND3 (N13847, N13842, N6473, N3308);
or OR4 (N13848, N13846, N3575, N8473, N2230);
or OR2 (N13849, N13843, N5241);
and AND4 (N13850, N13849, N8413, N8803, N1424);
nand NAND4 (N13851, N13844, N8257, N7855, N13133);
xor XOR2 (N13852, N13841, N13142);
xor XOR2 (N13853, N13850, N4311);
or OR2 (N13854, N13823, N4914);
nor NOR3 (N13855, N13834, N6058, N992);
not NOT1 (N13856, N13854);
xor XOR2 (N13857, N13781, N464);
buf BUF1 (N13858, N13857);
or OR4 (N13859, N13852, N6604, N2976, N6937);
not NOT1 (N13860, N13840);
not NOT1 (N13861, N13847);
xor XOR2 (N13862, N13860, N2268);
buf BUF1 (N13863, N13853);
or OR4 (N13864, N13863, N6902, N1925, N802);
nand NAND2 (N13865, N13864, N610);
not NOT1 (N13866, N13862);
not NOT1 (N13867, N13856);
nand NAND3 (N13868, N13858, N9042, N13099);
buf BUF1 (N13869, N13868);
xor XOR2 (N13870, N13861, N5497);
nor NOR3 (N13871, N13851, N2548, N10783);
nand NAND4 (N13872, N13867, N9049, N12371, N976);
xor XOR2 (N13873, N13866, N11784);
nor NOR4 (N13874, N13869, N10920, N10112, N5561);
nand NAND2 (N13875, N13872, N1469);
or OR4 (N13876, N13845, N13742, N12093, N9296);
or OR2 (N13877, N13848, N11863);
and AND2 (N13878, N13876, N11955);
buf BUF1 (N13879, N13855);
nand NAND4 (N13880, N13879, N6723, N12842, N8164);
and AND2 (N13881, N13880, N13457);
xor XOR2 (N13882, N13881, N10416);
not NOT1 (N13883, N13877);
nand NAND2 (N13884, N13871, N9151);
or OR2 (N13885, N13875, N1324);
xor XOR2 (N13886, N13865, N8591);
xor XOR2 (N13887, N13873, N12863);
not NOT1 (N13888, N13874);
or OR3 (N13889, N13888, N7803, N5302);
nor NOR3 (N13890, N13878, N9461, N7644);
not NOT1 (N13891, N13883);
nor NOR2 (N13892, N13889, N5217);
xor XOR2 (N13893, N13882, N6300);
xor XOR2 (N13894, N13891, N3075);
buf BUF1 (N13895, N13893);
not NOT1 (N13896, N13870);
not NOT1 (N13897, N13885);
or OR3 (N13898, N13890, N9727, N8236);
and AND3 (N13899, N13898, N12247, N12148);
nor NOR4 (N13900, N13899, N5186, N4879, N1971);
xor XOR2 (N13901, N13884, N230);
buf BUF1 (N13902, N13901);
buf BUF1 (N13903, N13900);
buf BUF1 (N13904, N13902);
not NOT1 (N13905, N13903);
buf BUF1 (N13906, N13905);
or OR2 (N13907, N13892, N3821);
and AND3 (N13908, N13886, N11877, N11990);
xor XOR2 (N13909, N13887, N7567);
nor NOR3 (N13910, N13894, N10446, N5425);
not NOT1 (N13911, N13910);
or OR2 (N13912, N13908, N2242);
xor XOR2 (N13913, N13897, N10492);
buf BUF1 (N13914, N13906);
nor NOR2 (N13915, N13909, N987);
nor NOR4 (N13916, N13896, N7755, N12583, N11904);
or OR2 (N13917, N13916, N12520);
xor XOR2 (N13918, N13904, N1047);
or OR3 (N13919, N13918, N8625, N7016);
nand NAND3 (N13920, N13912, N2617, N9089);
nand NAND3 (N13921, N13895, N11031, N13227);
or OR4 (N13922, N13917, N8276, N2978, N13806);
xor XOR2 (N13923, N13922, N13237);
or OR3 (N13924, N13914, N5276, N7958);
or OR3 (N13925, N13924, N9573, N4698);
and AND4 (N13926, N13919, N4211, N6961, N13659);
nor NOR4 (N13927, N13907, N1683, N2140, N8208);
buf BUF1 (N13928, N13859);
nand NAND3 (N13929, N13925, N12030, N5994);
not NOT1 (N13930, N13920);
and AND3 (N13931, N13915, N2147, N12573);
nor NOR2 (N13932, N13927, N5);
nand NAND4 (N13933, N13911, N1399, N9870, N2951);
and AND3 (N13934, N13913, N6953, N13709);
buf BUF1 (N13935, N13921);
nand NAND3 (N13936, N13934, N7657, N7305);
not NOT1 (N13937, N13931);
not NOT1 (N13938, N13936);
nor NOR3 (N13939, N13928, N11798, N118);
buf BUF1 (N13940, N13938);
xor XOR2 (N13941, N13926, N11163);
xor XOR2 (N13942, N13939, N2921);
buf BUF1 (N13943, N13932);
xor XOR2 (N13944, N13940, N6024);
buf BUF1 (N13945, N13929);
not NOT1 (N13946, N13933);
or OR3 (N13947, N13942, N8652, N3400);
xor XOR2 (N13948, N13935, N10411);
nand NAND4 (N13949, N13945, N264, N6153, N9369);
nand NAND3 (N13950, N13941, N6475, N1433);
nor NOR2 (N13951, N13943, N6898);
buf BUF1 (N13952, N13948);
buf BUF1 (N13953, N13944);
buf BUF1 (N13954, N13949);
nand NAND3 (N13955, N13950, N5342, N9788);
not NOT1 (N13956, N13937);
nor NOR2 (N13957, N13923, N1257);
or OR2 (N13958, N13956, N10978);
buf BUF1 (N13959, N13958);
xor XOR2 (N13960, N13957, N11858);
or OR3 (N13961, N13952, N2865, N13459);
and AND2 (N13962, N13954, N1776);
xor XOR2 (N13963, N13955, N8050);
nor NOR4 (N13964, N13961, N8781, N7838, N8135);
buf BUF1 (N13965, N13947);
buf BUF1 (N13966, N13965);
or OR2 (N13967, N13953, N7353);
and AND4 (N13968, N13946, N10077, N1222, N4300);
and AND2 (N13969, N13966, N3169);
or OR4 (N13970, N13964, N5520, N2239, N10192);
xor XOR2 (N13971, N13962, N3250);
and AND3 (N13972, N13960, N2352, N8825);
or OR4 (N13973, N13959, N2790, N7419, N8883);
or OR2 (N13974, N13970, N5903);
nand NAND4 (N13975, N13951, N10976, N1001, N3281);
nand NAND4 (N13976, N13972, N12744, N10586, N7600);
xor XOR2 (N13977, N13976, N3107);
not NOT1 (N13978, N13973);
buf BUF1 (N13979, N13967);
or OR2 (N13980, N13979, N9457);
and AND3 (N13981, N13974, N11774, N8434);
buf BUF1 (N13982, N13977);
and AND4 (N13983, N13963, N3231, N3627, N6815);
or OR4 (N13984, N13978, N13124, N7591, N13727);
not NOT1 (N13985, N13968);
buf BUF1 (N13986, N13985);
not NOT1 (N13987, N13982);
nand NAND2 (N13988, N13981, N3085);
and AND4 (N13989, N13930, N8171, N1188, N5076);
nor NOR2 (N13990, N13987, N8815);
buf BUF1 (N13991, N13983);
or OR3 (N13992, N13990, N10779, N2141);
nor NOR3 (N13993, N13980, N9368, N6387);
nor NOR4 (N13994, N13971, N12806, N11156, N9410);
xor XOR2 (N13995, N13986, N12126);
nand NAND4 (N13996, N13994, N6286, N2373, N9967);
xor XOR2 (N13997, N13996, N3896);
or OR4 (N13998, N13993, N10722, N3847, N3167);
not NOT1 (N13999, N13992);
not NOT1 (N14000, N13997);
nor NOR2 (N14001, N13969, N4943);
not NOT1 (N14002, N13984);
nand NAND3 (N14003, N13999, N6636, N1453);
and AND4 (N14004, N14000, N5999, N3892, N10786);
and AND4 (N14005, N13989, N6873, N10545, N1256);
and AND4 (N14006, N13988, N12360, N13319, N7678);
nor NOR4 (N14007, N14004, N1592, N7743, N2962);
nand NAND2 (N14008, N14005, N5030);
xor XOR2 (N14009, N14006, N1564);
and AND4 (N14010, N14008, N12221, N12750, N3035);
nand NAND3 (N14011, N14007, N7176, N2600);
not NOT1 (N14012, N14003);
nor NOR4 (N14013, N13991, N2293, N10728, N7118);
nor NOR3 (N14014, N14009, N7601, N1917);
nand NAND2 (N14015, N14013, N1661);
or OR2 (N14016, N14011, N7335);
nand NAND3 (N14017, N13998, N11488, N11297);
or OR3 (N14018, N14014, N1936, N13092);
or OR4 (N14019, N14001, N2016, N10516, N841);
or OR3 (N14020, N13975, N9394, N1508);
or OR4 (N14021, N13995, N5318, N3861, N654);
not NOT1 (N14022, N14002);
xor XOR2 (N14023, N14015, N12057);
nand NAND2 (N14024, N14010, N99);
buf BUF1 (N14025, N14024);
nor NOR4 (N14026, N14023, N8109, N11711, N13011);
and AND2 (N14027, N14018, N8911);
xor XOR2 (N14028, N14027, N13169);
or OR3 (N14029, N14016, N5937, N10381);
nor NOR2 (N14030, N14019, N14026);
buf BUF1 (N14031, N5007);
xor XOR2 (N14032, N14030, N14023);
nor NOR2 (N14033, N14021, N5701);
or OR4 (N14034, N14031, N8502, N9739, N4042);
and AND3 (N14035, N14022, N10400, N792);
or OR3 (N14036, N14034, N13953, N13197);
xor XOR2 (N14037, N14035, N11264);
and AND2 (N14038, N14025, N10966);
not NOT1 (N14039, N14029);
or OR4 (N14040, N14036, N13767, N12966, N4564);
nand NAND4 (N14041, N14012, N7572, N7150, N10420);
xor XOR2 (N14042, N14039, N2743);
buf BUF1 (N14043, N14017);
buf BUF1 (N14044, N14042);
or OR2 (N14045, N14032, N3018);
or OR3 (N14046, N14028, N10320, N13123);
or OR4 (N14047, N14043, N386, N2929, N7861);
buf BUF1 (N14048, N14045);
not NOT1 (N14049, N14048);
and AND2 (N14050, N14047, N9889);
nand NAND2 (N14051, N14046, N9125);
nand NAND4 (N14052, N14038, N11433, N6260, N2405);
or OR3 (N14053, N14050, N3364, N12970);
and AND3 (N14054, N14020, N5089, N8311);
and AND2 (N14055, N14037, N7935);
buf BUF1 (N14056, N14055);
nor NOR2 (N14057, N14049, N8075);
or OR2 (N14058, N14033, N8199);
or OR3 (N14059, N14058, N1715, N10881);
xor XOR2 (N14060, N14052, N12667);
nand NAND4 (N14061, N14059, N12029, N8783, N2789);
not NOT1 (N14062, N14061);
buf BUF1 (N14063, N14054);
xor XOR2 (N14064, N14057, N8350);
nor NOR2 (N14065, N14041, N2341);
and AND3 (N14066, N14063, N6486, N9867);
buf BUF1 (N14067, N14060);
nand NAND4 (N14068, N14066, N3487, N13724, N2645);
or OR4 (N14069, N14051, N13068, N13402, N2554);
or OR3 (N14070, N14064, N4890, N4457);
xor XOR2 (N14071, N14044, N8450);
not NOT1 (N14072, N14065);
nor NOR4 (N14073, N14062, N12525, N4744, N7567);
buf BUF1 (N14074, N14072);
xor XOR2 (N14075, N14053, N1893);
and AND3 (N14076, N14075, N4001, N9450);
and AND2 (N14077, N14074, N4879);
buf BUF1 (N14078, N14073);
or OR2 (N14079, N14070, N9677);
not NOT1 (N14080, N14056);
not NOT1 (N14081, N14067);
and AND3 (N14082, N14076, N6394, N677);
buf BUF1 (N14083, N14071);
buf BUF1 (N14084, N14069);
xor XOR2 (N14085, N14078, N4151);
buf BUF1 (N14086, N14083);
nand NAND2 (N14087, N14081, N12019);
nand NAND4 (N14088, N14087, N3929, N5826, N13403);
or OR2 (N14089, N14079, N12814);
or OR4 (N14090, N14077, N10626, N11495, N5311);
and AND4 (N14091, N14086, N4879, N1457, N8960);
or OR2 (N14092, N14088, N10281);
xor XOR2 (N14093, N14092, N4278);
nand NAND4 (N14094, N14040, N3097, N5576, N4869);
and AND2 (N14095, N14084, N11518);
and AND2 (N14096, N14095, N8162);
or OR4 (N14097, N14093, N1331, N11519, N6694);
nand NAND2 (N14098, N14089, N1393);
nand NAND3 (N14099, N14091, N2045, N1481);
nand NAND3 (N14100, N14097, N8244, N4757);
nor NOR2 (N14101, N14098, N6597);
not NOT1 (N14102, N14082);
and AND4 (N14103, N14080, N4249, N10928, N13074);
and AND3 (N14104, N14101, N12472, N6886);
or OR3 (N14105, N14096, N3232, N12998);
nor NOR3 (N14106, N14094, N245, N9691);
xor XOR2 (N14107, N14090, N12317);
buf BUF1 (N14108, N14104);
nor NOR3 (N14109, N14108, N13804, N11051);
and AND4 (N14110, N14109, N2628, N9856, N10524);
xor XOR2 (N14111, N14106, N6854);
and AND4 (N14112, N14102, N1666, N2840, N2463);
nor NOR2 (N14113, N14068, N4262);
xor XOR2 (N14114, N14105, N2639);
nor NOR3 (N14115, N14110, N1743, N3614);
nand NAND4 (N14116, N14100, N671, N2086, N12484);
nand NAND2 (N14117, N14113, N12675);
nand NAND2 (N14118, N14112, N3302);
xor XOR2 (N14119, N14107, N7802);
nor NOR2 (N14120, N14119, N3281);
or OR4 (N14121, N14118, N10447, N6319, N3828);
and AND3 (N14122, N14116, N11337, N12243);
nand NAND2 (N14123, N14122, N12007);
or OR4 (N14124, N14117, N11715, N2024, N3093);
nand NAND3 (N14125, N14085, N7964, N11896);
nor NOR2 (N14126, N14103, N6701);
and AND2 (N14127, N14121, N142);
nor NOR3 (N14128, N14123, N13219, N7066);
or OR4 (N14129, N14127, N5657, N7252, N10436);
xor XOR2 (N14130, N14129, N9239);
nor NOR2 (N14131, N14124, N9902);
buf BUF1 (N14132, N14126);
not NOT1 (N14133, N14125);
and AND3 (N14134, N14131, N8324, N12934);
and AND2 (N14135, N14134, N13211);
buf BUF1 (N14136, N14120);
and AND4 (N14137, N14130, N9799, N5401, N2809);
or OR2 (N14138, N14135, N4113);
xor XOR2 (N14139, N14137, N11900);
xor XOR2 (N14140, N14114, N10553);
and AND4 (N14141, N14133, N4059, N6385, N3000);
and AND2 (N14142, N14132, N10845);
nor NOR2 (N14143, N14139, N6003);
nor NOR4 (N14144, N14143, N2254, N7423, N13894);
nor NOR3 (N14145, N14136, N6250, N2458);
nand NAND3 (N14146, N14099, N11890, N11822);
not NOT1 (N14147, N14144);
nor NOR4 (N14148, N14138, N11387, N2546, N2);
or OR3 (N14149, N14111, N11239, N8011);
nor NOR2 (N14150, N14142, N6352);
nor NOR4 (N14151, N14146, N3351, N10744, N11760);
buf BUF1 (N14152, N14128);
buf BUF1 (N14153, N14151);
and AND2 (N14154, N14150, N9338);
not NOT1 (N14155, N14149);
buf BUF1 (N14156, N14152);
or OR3 (N14157, N14141, N6122, N9025);
nor NOR3 (N14158, N14156, N3416, N68);
buf BUF1 (N14159, N14147);
or OR4 (N14160, N14157, N7136, N12090, N12039);
not NOT1 (N14161, N14145);
xor XOR2 (N14162, N14161, N4896);
nor NOR3 (N14163, N14154, N9055, N3479);
or OR4 (N14164, N14159, N2035, N4201, N6284);
xor XOR2 (N14165, N14115, N11235);
buf BUF1 (N14166, N14160);
or OR3 (N14167, N14140, N4115, N9649);
nand NAND4 (N14168, N14158, N7299, N9370, N1002);
not NOT1 (N14169, N14164);
nand NAND3 (N14170, N14162, N7397, N12415);
not NOT1 (N14171, N14169);
nand NAND3 (N14172, N14163, N10368, N1866);
nor NOR3 (N14173, N14167, N12693, N285);
not NOT1 (N14174, N14148);
xor XOR2 (N14175, N14174, N13041);
buf BUF1 (N14176, N14173);
and AND3 (N14177, N14170, N10647, N13218);
and AND3 (N14178, N14155, N5574, N12855);
not NOT1 (N14179, N14171);
nand NAND4 (N14180, N14172, N6886, N11693, N5677);
nand NAND4 (N14181, N14175, N10813, N1747, N10739);
xor XOR2 (N14182, N14179, N4000);
buf BUF1 (N14183, N14153);
or OR3 (N14184, N14182, N1708, N14116);
nand NAND4 (N14185, N14165, N11207, N9212, N13457);
buf BUF1 (N14186, N14166);
not NOT1 (N14187, N14183);
buf BUF1 (N14188, N14178);
and AND2 (N14189, N14187, N12790);
not NOT1 (N14190, N14189);
nand NAND3 (N14191, N14180, N11309, N12844);
buf BUF1 (N14192, N14181);
buf BUF1 (N14193, N14176);
not NOT1 (N14194, N14185);
xor XOR2 (N14195, N14177, N6688);
not NOT1 (N14196, N14191);
buf BUF1 (N14197, N14192);
nand NAND3 (N14198, N14194, N704, N12390);
or OR2 (N14199, N14186, N8303);
xor XOR2 (N14200, N14197, N5976);
xor XOR2 (N14201, N14200, N11319);
buf BUF1 (N14202, N14184);
nor NOR3 (N14203, N14199, N5825, N10651);
nor NOR2 (N14204, N14196, N4298);
and AND2 (N14205, N14195, N3738);
or OR2 (N14206, N14190, N11717);
xor XOR2 (N14207, N14202, N5690);
nor NOR2 (N14208, N14188, N8107);
and AND3 (N14209, N14204, N4989, N2878);
nor NOR3 (N14210, N14201, N11311, N1437);
or OR3 (N14211, N14209, N9205, N2020);
not NOT1 (N14212, N14208);
or OR3 (N14213, N14203, N8285, N7826);
buf BUF1 (N14214, N14213);
not NOT1 (N14215, N14198);
not NOT1 (N14216, N14207);
xor XOR2 (N14217, N14216, N13135);
or OR4 (N14218, N14212, N4376, N5177, N9464);
xor XOR2 (N14219, N14210, N5798);
and AND4 (N14220, N14218, N4999, N13984, N10254);
xor XOR2 (N14221, N14219, N12262);
not NOT1 (N14222, N14211);
not NOT1 (N14223, N14214);
and AND2 (N14224, N14223, N2260);
or OR3 (N14225, N14168, N2546, N5199);
and AND2 (N14226, N14217, N7851);
and AND2 (N14227, N14226, N2101);
xor XOR2 (N14228, N14206, N2866);
not NOT1 (N14229, N14222);
xor XOR2 (N14230, N14215, N8304);
nor NOR2 (N14231, N14224, N8381);
or OR4 (N14232, N14229, N608, N5660, N3524);
nor NOR2 (N14233, N14221, N5189);
nor NOR4 (N14234, N14193, N9640, N2572, N13947);
buf BUF1 (N14235, N14220);
and AND2 (N14236, N14233, N3431);
not NOT1 (N14237, N14205);
xor XOR2 (N14238, N14228, N7363);
nand NAND2 (N14239, N14236, N10);
buf BUF1 (N14240, N14235);
buf BUF1 (N14241, N14239);
nor NOR4 (N14242, N14238, N8901, N5944, N6493);
xor XOR2 (N14243, N14241, N3104);
and AND3 (N14244, N14227, N14084, N7919);
or OR2 (N14245, N14240, N11025);
nor NOR3 (N14246, N14232, N6969, N2954);
not NOT1 (N14247, N14244);
xor XOR2 (N14248, N14245, N3499);
or OR4 (N14249, N14237, N11427, N10561, N6909);
or OR2 (N14250, N14249, N8463);
buf BUF1 (N14251, N14246);
not NOT1 (N14252, N14225);
nor NOR3 (N14253, N14230, N12491, N13967);
xor XOR2 (N14254, N14250, N2549);
nor NOR3 (N14255, N14243, N5830, N3805);
or OR3 (N14256, N14254, N7529, N10351);
xor XOR2 (N14257, N14253, N1208);
xor XOR2 (N14258, N14257, N11314);
and AND4 (N14259, N14255, N317, N6869, N9656);
nand NAND2 (N14260, N14248, N6415);
nand NAND2 (N14261, N14260, N814);
buf BUF1 (N14262, N14258);
and AND3 (N14263, N14242, N12082, N12695);
nor NOR3 (N14264, N14231, N7202, N4723);
nand NAND2 (N14265, N14234, N854);
buf BUF1 (N14266, N14256);
not NOT1 (N14267, N14251);
nand NAND4 (N14268, N14261, N9118, N1498, N7408);
nand NAND2 (N14269, N14267, N5416);
xor XOR2 (N14270, N14263, N1991);
and AND4 (N14271, N14264, N304, N7041, N6075);
not NOT1 (N14272, N14262);
buf BUF1 (N14273, N14259);
nand NAND4 (N14274, N14273, N13599, N13849, N12073);
or OR4 (N14275, N14268, N4596, N11827, N7670);
and AND3 (N14276, N14272, N12564, N11249);
nor NOR4 (N14277, N14270, N4098, N7785, N10126);
or OR2 (N14278, N14276, N10018);
buf BUF1 (N14279, N14274);
or OR4 (N14280, N14265, N12177, N6178, N14219);
and AND2 (N14281, N14275, N1046);
nor NOR2 (N14282, N14252, N5762);
or OR3 (N14283, N14266, N678, N3629);
nor NOR4 (N14284, N14278, N11414, N9159, N9096);
xor XOR2 (N14285, N14277, N47);
nand NAND4 (N14286, N14247, N1642, N7713, N12117);
and AND4 (N14287, N14285, N4006, N2007, N4610);
and AND4 (N14288, N14271, N7945, N4884, N9521);
and AND2 (N14289, N14269, N3226);
nor NOR4 (N14290, N14284, N9123, N844, N12796);
not NOT1 (N14291, N14283);
or OR3 (N14292, N14286, N13820, N6991);
xor XOR2 (N14293, N14279, N6298);
or OR4 (N14294, N14289, N795, N533, N13966);
buf BUF1 (N14295, N14280);
and AND2 (N14296, N14291, N4260);
buf BUF1 (N14297, N14292);
nor NOR4 (N14298, N14293, N2180, N7056, N5590);
nor NOR3 (N14299, N14281, N12924, N13478);
or OR2 (N14300, N14287, N314);
or OR4 (N14301, N14282, N12267, N6754, N9362);
buf BUF1 (N14302, N14295);
or OR3 (N14303, N14298, N8037, N1312);
buf BUF1 (N14304, N14288);
or OR2 (N14305, N14302, N3372);
not NOT1 (N14306, N14296);
xor XOR2 (N14307, N14290, N12289);
and AND4 (N14308, N14297, N3280, N7026, N8744);
nand NAND3 (N14309, N14307, N12973, N3928);
not NOT1 (N14310, N14294);
xor XOR2 (N14311, N14301, N4247);
and AND3 (N14312, N14299, N4315, N7521);
nand NAND4 (N14313, N14306, N3720, N9371, N11772);
and AND2 (N14314, N14311, N2696);
nor NOR2 (N14315, N14309, N9701);
not NOT1 (N14316, N14303);
nor NOR2 (N14317, N14308, N3217);
not NOT1 (N14318, N14300);
and AND3 (N14319, N14310, N5290, N6270);
and AND4 (N14320, N14319, N2703, N9555, N7481);
nand NAND2 (N14321, N14317, N6095);
nand NAND2 (N14322, N14315, N9697);
xor XOR2 (N14323, N14313, N1673);
nor NOR4 (N14324, N14312, N1278, N8441, N2904);
and AND2 (N14325, N14324, N3908);
nor NOR4 (N14326, N14321, N5085, N10390, N3641);
not NOT1 (N14327, N14325);
or OR3 (N14328, N14318, N8660, N4489);
or OR4 (N14329, N14316, N13566, N6180, N7721);
and AND2 (N14330, N14305, N4510);
or OR3 (N14331, N14320, N13461, N4249);
xor XOR2 (N14332, N14327, N9957);
and AND3 (N14333, N14326, N5305, N4473);
nor NOR3 (N14334, N14330, N1260, N10803);
nand NAND4 (N14335, N14314, N195, N1377, N7957);
or OR3 (N14336, N14329, N9026, N3386);
buf BUF1 (N14337, N14331);
or OR3 (N14338, N14336, N3883, N8605);
nand NAND2 (N14339, N14335, N2585);
or OR4 (N14340, N14328, N1090, N6635, N742);
and AND2 (N14341, N14323, N12534);
nand NAND3 (N14342, N14322, N970, N4126);
and AND2 (N14343, N14342, N8631);
not NOT1 (N14344, N14332);
buf BUF1 (N14345, N14334);
xor XOR2 (N14346, N14343, N2218);
nor NOR4 (N14347, N14304, N2375, N7386, N14177);
nand NAND4 (N14348, N14341, N11534, N8031, N6602);
and AND2 (N14349, N14338, N9619);
and AND3 (N14350, N14345, N7268, N1343);
nand NAND2 (N14351, N14346, N5415);
or OR3 (N14352, N14340, N11536, N14237);
xor XOR2 (N14353, N14352, N6688);
or OR4 (N14354, N14333, N3301, N12881, N8430);
nand NAND4 (N14355, N14344, N119, N12557, N10818);
not NOT1 (N14356, N14348);
or OR4 (N14357, N14347, N7189, N9586, N9402);
and AND4 (N14358, N14353, N2446, N12490, N3773);
xor XOR2 (N14359, N14337, N5921);
nand NAND2 (N14360, N14357, N12033);
nor NOR3 (N14361, N14358, N9265, N11822);
nor NOR3 (N14362, N14356, N7287, N8984);
and AND3 (N14363, N14354, N2671, N1496);
buf BUF1 (N14364, N14351);
nand NAND4 (N14365, N14355, N7617, N11396, N9937);
nor NOR3 (N14366, N14339, N9163, N4154);
xor XOR2 (N14367, N14365, N7862);
xor XOR2 (N14368, N14349, N13934);
or OR2 (N14369, N14367, N12129);
or OR3 (N14370, N14361, N8473, N10002);
not NOT1 (N14371, N14363);
xor XOR2 (N14372, N14360, N13576);
buf BUF1 (N14373, N14364);
buf BUF1 (N14374, N14368);
and AND2 (N14375, N14359, N4111);
xor XOR2 (N14376, N14370, N11736);
nor NOR2 (N14377, N14372, N5849);
nor NOR2 (N14378, N14374, N2470);
not NOT1 (N14379, N14373);
xor XOR2 (N14380, N14350, N1300);
xor XOR2 (N14381, N14362, N10163);
nand NAND3 (N14382, N14366, N10412, N1328);
and AND3 (N14383, N14378, N4458, N5983);
and AND4 (N14384, N14376, N1286, N8606, N7391);
buf BUF1 (N14385, N14379);
not NOT1 (N14386, N14385);
xor XOR2 (N14387, N14371, N11683);
xor XOR2 (N14388, N14377, N6980);
or OR4 (N14389, N14386, N2418, N8998, N3659);
nand NAND3 (N14390, N14383, N13490, N12961);
or OR2 (N14391, N14382, N12825);
not NOT1 (N14392, N14381);
xor XOR2 (N14393, N14380, N8056);
nor NOR4 (N14394, N14393, N13492, N7006, N187);
buf BUF1 (N14395, N14394);
nand NAND2 (N14396, N14384, N12831);
xor XOR2 (N14397, N14390, N10763);
nor NOR2 (N14398, N14395, N313);
xor XOR2 (N14399, N14398, N10212);
nor NOR3 (N14400, N14396, N4746, N9469);
or OR4 (N14401, N14388, N9313, N9501, N682);
nand NAND3 (N14402, N14375, N133, N7535);
and AND3 (N14403, N14391, N1328, N3599);
not NOT1 (N14404, N14401);
not NOT1 (N14405, N14400);
and AND2 (N14406, N14389, N12389);
nor NOR4 (N14407, N14397, N7960, N237, N3280);
and AND3 (N14408, N14369, N3198, N4693);
and AND4 (N14409, N14404, N13629, N7796, N2048);
nor NOR2 (N14410, N14403, N10161);
not NOT1 (N14411, N14410);
nor NOR4 (N14412, N14409, N12548, N595, N8387);
not NOT1 (N14413, N14408);
or OR4 (N14414, N14406, N13134, N11688, N14305);
xor XOR2 (N14415, N14387, N7414);
or OR4 (N14416, N14407, N5400, N14408, N2826);
and AND3 (N14417, N14415, N5690, N14024);
buf BUF1 (N14418, N14411);
not NOT1 (N14419, N14416);
nand NAND4 (N14420, N14405, N3933, N9218, N8336);
nor NOR2 (N14421, N14412, N2095);
and AND2 (N14422, N14414, N12955);
xor XOR2 (N14423, N14421, N7298);
nor NOR4 (N14424, N14392, N8864, N4781, N10543);
nand NAND2 (N14425, N14417, N7231);
or OR4 (N14426, N14399, N11714, N5968, N5945);
xor XOR2 (N14427, N14419, N329);
nor NOR3 (N14428, N14427, N12228, N8167);
buf BUF1 (N14429, N14426);
nand NAND4 (N14430, N14402, N7853, N3158, N7800);
nand NAND2 (N14431, N14420, N11579);
and AND3 (N14432, N14423, N5743, N7975);
nand NAND3 (N14433, N14418, N1849, N2399);
not NOT1 (N14434, N14433);
xor XOR2 (N14435, N14413, N7683);
nand NAND3 (N14436, N14428, N3641, N11995);
and AND2 (N14437, N14422, N6278);
or OR2 (N14438, N14434, N13010);
buf BUF1 (N14439, N14436);
and AND4 (N14440, N14429, N4481, N5249, N2201);
not NOT1 (N14441, N14437);
xor XOR2 (N14442, N14431, N4881);
nand NAND4 (N14443, N14442, N5818, N6749, N7033);
xor XOR2 (N14444, N14435, N4227);
or OR2 (N14445, N14430, N1872);
nand NAND3 (N14446, N14443, N3837, N6827);
and AND3 (N14447, N14444, N12305, N13268);
or OR3 (N14448, N14445, N6433, N7484);
buf BUF1 (N14449, N14439);
nor NOR3 (N14450, N14449, N5658, N11188);
or OR2 (N14451, N14424, N1809);
and AND3 (N14452, N14438, N9529, N10318);
or OR2 (N14453, N14446, N14326);
buf BUF1 (N14454, N14451);
nor NOR3 (N14455, N14454, N10078, N4474);
xor XOR2 (N14456, N14432, N4494);
nor NOR2 (N14457, N14455, N13971);
nand NAND2 (N14458, N14450, N7126);
nand NAND4 (N14459, N14453, N6034, N9810, N8583);
not NOT1 (N14460, N14447);
and AND2 (N14461, N14448, N9634);
buf BUF1 (N14462, N14440);
nand NAND4 (N14463, N14458, N1672, N9140, N3551);
nand NAND2 (N14464, N14425, N2490);
xor XOR2 (N14465, N14452, N1910);
and AND4 (N14466, N14441, N9631, N1230, N11043);
xor XOR2 (N14467, N14459, N4773);
or OR2 (N14468, N14466, N5677);
or OR4 (N14469, N14468, N8156, N2841, N10671);
buf BUF1 (N14470, N14463);
not NOT1 (N14471, N14469);
buf BUF1 (N14472, N14470);
buf BUF1 (N14473, N14464);
not NOT1 (N14474, N14462);
or OR2 (N14475, N14461, N11889);
and AND4 (N14476, N14471, N11738, N11278, N9072);
not NOT1 (N14477, N14456);
xor XOR2 (N14478, N14476, N10316);
xor XOR2 (N14479, N14457, N8152);
nor NOR3 (N14480, N14460, N13826, N12488);
nor NOR4 (N14481, N14474, N6275, N12454, N9888);
and AND4 (N14482, N14477, N10444, N6655, N5535);
buf BUF1 (N14483, N14472);
nand NAND2 (N14484, N14478, N902);
or OR3 (N14485, N14465, N9511, N3805);
or OR4 (N14486, N14473, N11918, N5620, N1727);
nand NAND4 (N14487, N14480, N2634, N9674, N11228);
xor XOR2 (N14488, N14484, N11342);
nand NAND4 (N14489, N14479, N5198, N8346, N757);
or OR4 (N14490, N14467, N125, N8654, N13883);
xor XOR2 (N14491, N14486, N1025);
xor XOR2 (N14492, N14475, N837);
nor NOR2 (N14493, N14490, N721);
xor XOR2 (N14494, N14483, N5059);
buf BUF1 (N14495, N14488);
or OR4 (N14496, N14491, N7095, N2188, N4384);
nor NOR3 (N14497, N14485, N11812, N9562);
or OR4 (N14498, N14497, N13895, N12268, N5587);
nor NOR3 (N14499, N14494, N10871, N2462);
nand NAND2 (N14500, N14496, N3184);
and AND4 (N14501, N14492, N10032, N6911, N1167);
or OR4 (N14502, N14500, N9379, N353, N9642);
or OR2 (N14503, N14498, N14198);
not NOT1 (N14504, N14482);
nor NOR3 (N14505, N14487, N12959, N2748);
xor XOR2 (N14506, N14502, N14127);
or OR2 (N14507, N14499, N1359);
and AND4 (N14508, N14504, N8173, N11490, N9063);
buf BUF1 (N14509, N14505);
nand NAND2 (N14510, N14509, N14157);
xor XOR2 (N14511, N14503, N4899);
and AND4 (N14512, N14506, N11773, N3284, N11560);
buf BUF1 (N14513, N14512);
nand NAND2 (N14514, N14507, N11172);
nor NOR4 (N14515, N14513, N10522, N12044, N12703);
nand NAND2 (N14516, N14501, N8937);
not NOT1 (N14517, N14489);
and AND4 (N14518, N14508, N5054, N8244, N440);
xor XOR2 (N14519, N14511, N3584);
nand NAND3 (N14520, N14514, N8457, N13618);
or OR2 (N14521, N14519, N13945);
or OR2 (N14522, N14481, N2214);
and AND2 (N14523, N14510, N8569);
and AND4 (N14524, N14515, N5391, N6424, N14365);
nor NOR4 (N14525, N14493, N10271, N9053, N6881);
or OR4 (N14526, N14520, N80, N5803, N8628);
nor NOR3 (N14527, N14516, N5122, N3917);
buf BUF1 (N14528, N14525);
not NOT1 (N14529, N14517);
and AND4 (N14530, N14518, N11802, N1831, N7936);
nand NAND2 (N14531, N14495, N2252);
and AND2 (N14532, N14528, N5743);
nor NOR3 (N14533, N14527, N11747, N2520);
nand NAND4 (N14534, N14526, N11826, N9877, N11965);
nand NAND3 (N14535, N14533, N14272, N10736);
nor NOR2 (N14536, N14529, N4737);
xor XOR2 (N14537, N14522, N218);
xor XOR2 (N14538, N14523, N3478);
not NOT1 (N14539, N14536);
not NOT1 (N14540, N14537);
xor XOR2 (N14541, N14534, N4058);
or OR4 (N14542, N14539, N1694, N13344, N12092);
xor XOR2 (N14543, N14521, N12113);
and AND3 (N14544, N14530, N2650, N650);
or OR3 (N14545, N14524, N9947, N138);
xor XOR2 (N14546, N14542, N12108);
nand NAND4 (N14547, N14535, N9135, N3255, N11279);
xor XOR2 (N14548, N14541, N12039);
or OR4 (N14549, N14545, N13429, N14500, N3265);
and AND2 (N14550, N14540, N7616);
or OR4 (N14551, N14531, N8538, N6472, N7492);
xor XOR2 (N14552, N14547, N14127);
or OR2 (N14553, N14551, N4884);
and AND2 (N14554, N14543, N6596);
nor NOR3 (N14555, N14549, N8198, N9738);
nor NOR2 (N14556, N14538, N11869);
nand NAND3 (N14557, N14546, N169, N2183);
nor NOR3 (N14558, N14553, N3415, N14315);
nor NOR4 (N14559, N14558, N14350, N3816, N3614);
and AND4 (N14560, N14550, N7873, N11870, N9109);
and AND2 (N14561, N14548, N4334);
nand NAND3 (N14562, N14561, N11892, N192);
nor NOR2 (N14563, N14555, N13383);
buf BUF1 (N14564, N14544);
nand NAND3 (N14565, N14564, N7488, N12217);
xor XOR2 (N14566, N14554, N2814);
or OR3 (N14567, N14565, N2354, N216);
or OR3 (N14568, N14560, N12617, N4424);
or OR3 (N14569, N14556, N6431, N11850);
not NOT1 (N14570, N14567);
buf BUF1 (N14571, N14569);
or OR4 (N14572, N14571, N6066, N8486, N1127);
and AND2 (N14573, N14532, N103);
nand NAND3 (N14574, N14562, N13505, N3081);
nand NAND4 (N14575, N14559, N11288, N4854, N7274);
nor NOR3 (N14576, N14573, N4351, N1904);
nor NOR2 (N14577, N14572, N13855);
nand NAND4 (N14578, N14577, N9580, N2412, N11150);
not NOT1 (N14579, N14576);
nand NAND3 (N14580, N14574, N9571, N11296);
xor XOR2 (N14581, N14579, N4540);
nand NAND3 (N14582, N14570, N10061, N14213);
xor XOR2 (N14583, N14581, N2141);
xor XOR2 (N14584, N14557, N11346);
and AND3 (N14585, N14568, N1209, N3422);
nor NOR4 (N14586, N14583, N10070, N2618, N1777);
buf BUF1 (N14587, N14578);
nor NOR3 (N14588, N14552, N3597, N5030);
or OR4 (N14589, N14587, N11107, N2589, N4893);
xor XOR2 (N14590, N14566, N12940);
not NOT1 (N14591, N14590);
buf BUF1 (N14592, N14591);
xor XOR2 (N14593, N14582, N5919);
and AND2 (N14594, N14575, N5350);
nor NOR4 (N14595, N14593, N3738, N9145, N8367);
nand NAND3 (N14596, N14588, N12425, N2300);
buf BUF1 (N14597, N14596);
or OR4 (N14598, N14580, N12857, N6797, N12821);
or OR3 (N14599, N14586, N13127, N14228);
nand NAND4 (N14600, N14598, N5217, N12057, N14580);
nor NOR4 (N14601, N14597, N10623, N2913, N5168);
not NOT1 (N14602, N14592);
buf BUF1 (N14603, N14563);
not NOT1 (N14604, N14585);
not NOT1 (N14605, N14600);
nand NAND2 (N14606, N14595, N7664);
xor XOR2 (N14607, N14601, N13572);
or OR4 (N14608, N14606, N5092, N12908, N3576);
nor NOR2 (N14609, N14604, N8463);
not NOT1 (N14610, N14608);
not NOT1 (N14611, N14584);
nor NOR4 (N14612, N14611, N5426, N13756, N1511);
buf BUF1 (N14613, N14612);
xor XOR2 (N14614, N14599, N3154);
buf BUF1 (N14615, N14602);
and AND4 (N14616, N14589, N5390, N5763, N14399);
buf BUF1 (N14617, N14616);
or OR2 (N14618, N14614, N313);
not NOT1 (N14619, N14618);
or OR4 (N14620, N14615, N12570, N12685, N3674);
xor XOR2 (N14621, N14603, N4706);
and AND4 (N14622, N14617, N5586, N1747, N1266);
xor XOR2 (N14623, N14609, N12650);
nor NOR4 (N14624, N14607, N8438, N2782, N5938);
and AND4 (N14625, N14605, N1777, N4501, N9421);
buf BUF1 (N14626, N14619);
nor NOR3 (N14627, N14625, N13692, N9762);
not NOT1 (N14628, N14624);
and AND4 (N14629, N14613, N78, N8279, N5639);
or OR3 (N14630, N14623, N10140, N13821);
not NOT1 (N14631, N14626);
nor NOR3 (N14632, N14629, N7606, N13457);
buf BUF1 (N14633, N14610);
nand NAND2 (N14634, N14594, N7478);
not NOT1 (N14635, N14627);
and AND3 (N14636, N14633, N11035, N13973);
nor NOR2 (N14637, N14631, N5780);
and AND2 (N14638, N14630, N8569);
nor NOR2 (N14639, N14635, N3603);
and AND2 (N14640, N14637, N13318);
nor NOR3 (N14641, N14639, N13474, N5087);
xor XOR2 (N14642, N14632, N12044);
buf BUF1 (N14643, N14638);
nor NOR3 (N14644, N14620, N6512, N3298);
not NOT1 (N14645, N14640);
not NOT1 (N14646, N14642);
or OR3 (N14647, N14628, N5759, N9478);
or OR4 (N14648, N14634, N8395, N1637, N7998);
not NOT1 (N14649, N14648);
nor NOR4 (N14650, N14645, N8576, N12113, N5417);
buf BUF1 (N14651, N14649);
buf BUF1 (N14652, N14646);
nand NAND4 (N14653, N14644, N5329, N10734, N7236);
and AND4 (N14654, N14622, N7965, N1808, N6922);
nor NOR2 (N14655, N14643, N6216);
nand NAND3 (N14656, N14636, N6231, N9112);
nor NOR3 (N14657, N14651, N181, N1787);
and AND3 (N14658, N14653, N4381, N4992);
buf BUF1 (N14659, N14654);
nand NAND4 (N14660, N14657, N11741, N11374, N8134);
or OR3 (N14661, N14650, N13477, N7629);
nor NOR4 (N14662, N14656, N10285, N11484, N1293);
xor XOR2 (N14663, N14658, N14400);
nor NOR4 (N14664, N14660, N11468, N8490, N12244);
xor XOR2 (N14665, N14662, N2253);
nand NAND2 (N14666, N14641, N11363);
buf BUF1 (N14667, N14665);
not NOT1 (N14668, N14647);
nor NOR4 (N14669, N14661, N5701, N3952, N1604);
nand NAND2 (N14670, N14621, N13187);
and AND4 (N14671, N14663, N12062, N7656, N6276);
and AND2 (N14672, N14667, N4143);
xor XOR2 (N14673, N14668, N8470);
or OR3 (N14674, N14671, N10353, N13452);
buf BUF1 (N14675, N14659);
or OR3 (N14676, N14652, N13875, N4713);
xor XOR2 (N14677, N14655, N4220);
nor NOR2 (N14678, N14666, N172);
and AND3 (N14679, N14676, N2226, N9882);
not NOT1 (N14680, N14678);
xor XOR2 (N14681, N14664, N5973);
xor XOR2 (N14682, N14680, N13797);
nand NAND2 (N14683, N14677, N1469);
nor NOR4 (N14684, N14669, N13599, N12609, N11875);
and AND4 (N14685, N14670, N691, N7908, N6008);
buf BUF1 (N14686, N14684);
buf BUF1 (N14687, N14681);
nor NOR4 (N14688, N14686, N2209, N5492, N5071);
nand NAND2 (N14689, N14673, N1610);
buf BUF1 (N14690, N14685);
nor NOR4 (N14691, N14679, N5304, N1079, N6810);
nor NOR4 (N14692, N14687, N14200, N11619, N4438);
nand NAND4 (N14693, N14692, N9654, N14638, N11519);
and AND3 (N14694, N14672, N4419, N5407);
or OR4 (N14695, N14674, N11275, N7663, N14434);
or OR3 (N14696, N14675, N541, N13014);
nand NAND4 (N14697, N14693, N8104, N8066, N4141);
not NOT1 (N14698, N14696);
buf BUF1 (N14699, N14682);
not NOT1 (N14700, N14694);
or OR2 (N14701, N14688, N2668);
not NOT1 (N14702, N14689);
nor NOR3 (N14703, N14702, N9902, N9119);
nand NAND4 (N14704, N14683, N7269, N3017, N12634);
nor NOR4 (N14705, N14690, N10355, N7252, N8318);
nand NAND3 (N14706, N14698, N14484, N5282);
and AND4 (N14707, N14701, N4186, N437, N6053);
or OR2 (N14708, N14691, N14568);
nand NAND2 (N14709, N14700, N12918);
nor NOR3 (N14710, N14705, N4886, N5307);
xor XOR2 (N14711, N14695, N11519);
xor XOR2 (N14712, N14703, N12822);
or OR3 (N14713, N14710, N10860, N14607);
and AND4 (N14714, N14713, N7172, N1598, N1523);
nor NOR2 (N14715, N14709, N688);
and AND4 (N14716, N14707, N4913, N7021, N6725);
not NOT1 (N14717, N14712);
xor XOR2 (N14718, N14704, N9938);
and AND3 (N14719, N14708, N8401, N1464);
or OR2 (N14720, N14719, N1738);
xor XOR2 (N14721, N14699, N10275);
not NOT1 (N14722, N14718);
xor XOR2 (N14723, N14697, N2490);
nor NOR4 (N14724, N14720, N4676, N3611, N14451);
or OR2 (N14725, N14716, N11131);
not NOT1 (N14726, N14725);
and AND3 (N14727, N14714, N9403, N4403);
or OR4 (N14728, N14715, N5557, N5192, N6211);
not NOT1 (N14729, N14722);
and AND2 (N14730, N14726, N8878);
xor XOR2 (N14731, N14728, N13351);
buf BUF1 (N14732, N14717);
nand NAND3 (N14733, N14711, N14226, N809);
or OR3 (N14734, N14721, N14150, N2903);
nand NAND4 (N14735, N14734, N5050, N3619, N13652);
not NOT1 (N14736, N14733);
xor XOR2 (N14737, N14706, N13411);
buf BUF1 (N14738, N14729);
nor NOR3 (N14739, N14738, N3120, N1265);
or OR2 (N14740, N14736, N11449);
or OR4 (N14741, N14732, N5040, N9519, N373);
and AND2 (N14742, N14727, N4438);
xor XOR2 (N14743, N14735, N1636);
nand NAND3 (N14744, N14742, N7543, N9694);
not NOT1 (N14745, N14724);
nor NOR2 (N14746, N14740, N1165);
buf BUF1 (N14747, N14730);
xor XOR2 (N14748, N14743, N3728);
nand NAND3 (N14749, N14739, N11359, N10057);
buf BUF1 (N14750, N14749);
and AND2 (N14751, N14723, N13420);
or OR4 (N14752, N14744, N5980, N1054, N3836);
not NOT1 (N14753, N14731);
not NOT1 (N14754, N14751);
buf BUF1 (N14755, N14748);
or OR3 (N14756, N14755, N2658, N8643);
nor NOR2 (N14757, N14747, N9420);
buf BUF1 (N14758, N14750);
xor XOR2 (N14759, N14752, N8650);
nand NAND3 (N14760, N14753, N737, N11626);
or OR4 (N14761, N14741, N4900, N9732, N14334);
buf BUF1 (N14762, N14757);
and AND4 (N14763, N14759, N5004, N7883, N12463);
nand NAND4 (N14764, N14760, N2939, N3397, N10297);
not NOT1 (N14765, N14745);
and AND3 (N14766, N14737, N1899, N13203);
and AND3 (N14767, N14758, N10040, N9061);
and AND4 (N14768, N14756, N3110, N9347, N3867);
nand NAND3 (N14769, N14767, N7456, N12443);
nor NOR2 (N14770, N14746, N14344);
or OR4 (N14771, N14763, N7888, N804, N12218);
and AND3 (N14772, N14768, N10121, N487);
or OR4 (N14773, N14754, N645, N5667, N1665);
and AND3 (N14774, N14772, N1118, N14519);
nand NAND3 (N14775, N14765, N5003, N7361);
or OR2 (N14776, N14766, N1769);
buf BUF1 (N14777, N14775);
nor NOR4 (N14778, N14762, N6769, N12692, N7443);
nand NAND3 (N14779, N14776, N9663, N9938);
not NOT1 (N14780, N14777);
nand NAND3 (N14781, N14780, N10665, N11885);
nor NOR4 (N14782, N14778, N11102, N10187, N2826);
nand NAND3 (N14783, N14769, N10523, N3766);
or OR2 (N14784, N14773, N8251);
nor NOR3 (N14785, N14784, N5994, N3075);
buf BUF1 (N14786, N14761);
and AND2 (N14787, N14786, N8041);
xor XOR2 (N14788, N14783, N1791);
and AND2 (N14789, N14779, N10449);
not NOT1 (N14790, N14782);
buf BUF1 (N14791, N14785);
not NOT1 (N14792, N14771);
or OR2 (N14793, N14770, N588);
and AND3 (N14794, N14790, N6112, N67);
or OR4 (N14795, N14764, N2357, N9427, N9110);
xor XOR2 (N14796, N14787, N11026);
buf BUF1 (N14797, N14794);
nand NAND2 (N14798, N14774, N7293);
and AND2 (N14799, N14781, N9639);
nor NOR4 (N14800, N14795, N6926, N11995, N4618);
nand NAND2 (N14801, N14791, N4269);
nor NOR2 (N14802, N14793, N13275);
nand NAND3 (N14803, N14789, N8919, N3656);
xor XOR2 (N14804, N14801, N3345);
buf BUF1 (N14805, N14799);
buf BUF1 (N14806, N14797);
and AND4 (N14807, N14798, N10505, N4615, N7633);
and AND3 (N14808, N14788, N9631, N1793);
nor NOR4 (N14809, N14796, N12336, N6036, N13004);
nor NOR2 (N14810, N14807, N13159);
nand NAND2 (N14811, N14792, N104);
buf BUF1 (N14812, N14802);
or OR4 (N14813, N14809, N14117, N5572, N13729);
or OR3 (N14814, N14812, N11554, N8233);
xor XOR2 (N14815, N14811, N8772);
buf BUF1 (N14816, N14810);
or OR2 (N14817, N14813, N9943);
or OR3 (N14818, N14814, N13323, N1061);
buf BUF1 (N14819, N14817);
buf BUF1 (N14820, N14808);
nand NAND3 (N14821, N14800, N13832, N9844);
nand NAND2 (N14822, N14819, N13213);
buf BUF1 (N14823, N14806);
nor NOR4 (N14824, N14815, N14402, N11721, N1788);
or OR2 (N14825, N14818, N12209);
nor NOR4 (N14826, N14805, N10526, N2089, N10222);
xor XOR2 (N14827, N14820, N2678);
xor XOR2 (N14828, N14824, N4696);
nand NAND4 (N14829, N14828, N6305, N6526, N8750);
or OR3 (N14830, N14816, N8226, N3437);
xor XOR2 (N14831, N14830, N14314);
or OR3 (N14832, N14825, N11669, N742);
xor XOR2 (N14833, N14822, N7357);
buf BUF1 (N14834, N14827);
or OR4 (N14835, N14803, N11654, N8507, N13245);
not NOT1 (N14836, N14826);
xor XOR2 (N14837, N14831, N11841);
buf BUF1 (N14838, N14829);
nand NAND4 (N14839, N14821, N11221, N2690, N9706);
nand NAND2 (N14840, N14823, N12048);
or OR4 (N14841, N14838, N2695, N6978, N3237);
not NOT1 (N14842, N14840);
xor XOR2 (N14843, N14836, N13053);
xor XOR2 (N14844, N14841, N2321);
not NOT1 (N14845, N14804);
not NOT1 (N14846, N14835);
buf BUF1 (N14847, N14842);
or OR2 (N14848, N14839, N1362);
buf BUF1 (N14849, N14847);
xor XOR2 (N14850, N14845, N11338);
buf BUF1 (N14851, N14834);
buf BUF1 (N14852, N14846);
or OR4 (N14853, N14848, N14135, N3053, N13551);
nor NOR2 (N14854, N14833, N9376);
or OR2 (N14855, N14854, N3475);
nor NOR3 (N14856, N14844, N9133, N10849);
and AND3 (N14857, N14832, N7879, N5861);
nand NAND2 (N14858, N14849, N4119);
xor XOR2 (N14859, N14855, N1475);
and AND3 (N14860, N14853, N10580, N3218);
buf BUF1 (N14861, N14837);
not NOT1 (N14862, N14851);
nand NAND2 (N14863, N14859, N13939);
not NOT1 (N14864, N14860);
not NOT1 (N14865, N14858);
xor XOR2 (N14866, N14856, N8933);
xor XOR2 (N14867, N14852, N9101);
and AND4 (N14868, N14843, N13383, N10259, N5250);
or OR3 (N14869, N14861, N698, N8580);
buf BUF1 (N14870, N14862);
or OR4 (N14871, N14870, N8824, N5097, N2846);
nand NAND2 (N14872, N14865, N439);
buf BUF1 (N14873, N14850);
xor XOR2 (N14874, N14868, N1532);
and AND3 (N14875, N14869, N8263, N9250);
buf BUF1 (N14876, N14866);
nand NAND3 (N14877, N14872, N4490, N5328);
not NOT1 (N14878, N14873);
not NOT1 (N14879, N14867);
nand NAND2 (N14880, N14879, N12011);
nor NOR4 (N14881, N14878, N9283, N1882, N708);
not NOT1 (N14882, N14881);
or OR3 (N14883, N14880, N12036, N3506);
not NOT1 (N14884, N14863);
or OR4 (N14885, N14882, N12270, N2581, N13183);
xor XOR2 (N14886, N14864, N5203);
nand NAND2 (N14887, N14886, N3737);
xor XOR2 (N14888, N14883, N11155);
or OR2 (N14889, N14887, N9257);
nand NAND2 (N14890, N14876, N12595);
or OR2 (N14891, N14888, N12659);
buf BUF1 (N14892, N14884);
buf BUF1 (N14893, N14891);
not NOT1 (N14894, N14875);
and AND3 (N14895, N14890, N892, N10150);
buf BUF1 (N14896, N14892);
xor XOR2 (N14897, N14885, N14717);
and AND2 (N14898, N14896, N3790);
buf BUF1 (N14899, N14898);
buf BUF1 (N14900, N14897);
not NOT1 (N14901, N14895);
not NOT1 (N14902, N14874);
or OR3 (N14903, N14894, N4382, N1338);
buf BUF1 (N14904, N14889);
or OR3 (N14905, N14893, N3377, N143);
nand NAND4 (N14906, N14871, N13566, N235, N10788);
and AND2 (N14907, N14877, N5732);
nor NOR3 (N14908, N14903, N5785, N10463);
xor XOR2 (N14909, N14907, N9488);
xor XOR2 (N14910, N14909, N6977);
and AND3 (N14911, N14857, N9400, N9328);
not NOT1 (N14912, N14905);
and AND3 (N14913, N14911, N8791, N7872);
xor XOR2 (N14914, N14900, N72);
buf BUF1 (N14915, N14914);
buf BUF1 (N14916, N14913);
nor NOR2 (N14917, N14912, N1964);
buf BUF1 (N14918, N14906);
nand NAND4 (N14919, N14915, N9678, N8851, N1661);
not NOT1 (N14920, N14918);
xor XOR2 (N14921, N14904, N9094);
or OR2 (N14922, N14899, N4782);
not NOT1 (N14923, N14910);
and AND3 (N14924, N14902, N2923, N1080);
or OR4 (N14925, N14923, N14351, N1165, N1981);
or OR3 (N14926, N14924, N5825, N9468);
nor NOR2 (N14927, N14921, N3594);
nand NAND2 (N14928, N14908, N5416);
buf BUF1 (N14929, N14919);
xor XOR2 (N14930, N14901, N9695);
not NOT1 (N14931, N14916);
nand NAND3 (N14932, N14920, N12661, N5888);
nor NOR3 (N14933, N14928, N3618, N642);
and AND2 (N14934, N14931, N6688);
or OR2 (N14935, N14930, N8803);
or OR2 (N14936, N14925, N4128);
not NOT1 (N14937, N14934);
and AND4 (N14938, N14935, N6473, N12822, N17);
xor XOR2 (N14939, N14922, N10813);
nor NOR2 (N14940, N14929, N8713);
or OR2 (N14941, N14927, N11399);
nand NAND2 (N14942, N14939, N12795);
xor XOR2 (N14943, N14936, N5709);
buf BUF1 (N14944, N14932);
or OR2 (N14945, N14943, N10057);
or OR2 (N14946, N14933, N2697);
and AND4 (N14947, N14941, N4262, N6049, N3360);
nand NAND2 (N14948, N14917, N5161);
buf BUF1 (N14949, N14938);
or OR2 (N14950, N14947, N7300);
or OR3 (N14951, N14948, N9286, N1336);
not NOT1 (N14952, N14937);
buf BUF1 (N14953, N14944);
xor XOR2 (N14954, N14951, N9757);
nor NOR3 (N14955, N14926, N7251, N8683);
buf BUF1 (N14956, N14940);
or OR4 (N14957, N14950, N10724, N7302, N8490);
buf BUF1 (N14958, N14956);
buf BUF1 (N14959, N14955);
or OR2 (N14960, N14945, N987);
and AND4 (N14961, N14958, N3082, N11276, N12487);
nor NOR3 (N14962, N14952, N6271, N4636);
nand NAND3 (N14963, N14953, N6588, N8159);
nand NAND3 (N14964, N14960, N6805, N3356);
buf BUF1 (N14965, N14959);
buf BUF1 (N14966, N14962);
xor XOR2 (N14967, N14949, N12253);
xor XOR2 (N14968, N14961, N390);
nor NOR2 (N14969, N14968, N8978);
nor NOR3 (N14970, N14967, N6815, N6738);
not NOT1 (N14971, N14970);
nor NOR4 (N14972, N14942, N2855, N6737, N5934);
not NOT1 (N14973, N14972);
nor NOR2 (N14974, N14973, N8497);
xor XOR2 (N14975, N14965, N13502);
buf BUF1 (N14976, N14946);
nor NOR4 (N14977, N14957, N1957, N7831, N14064);
xor XOR2 (N14978, N14969, N10514);
not NOT1 (N14979, N14974);
xor XOR2 (N14980, N14979, N7322);
not NOT1 (N14981, N14977);
nor NOR2 (N14982, N14971, N8258);
nand NAND3 (N14983, N14975, N14290, N6270);
or OR3 (N14984, N14964, N11694, N5557);
or OR3 (N14985, N14963, N2752, N10479);
not NOT1 (N14986, N14954);
nand NAND2 (N14987, N14983, N1265);
and AND4 (N14988, N14982, N12248, N14323, N5911);
and AND2 (N14989, N14986, N2895);
not NOT1 (N14990, N14976);
buf BUF1 (N14991, N14980);
and AND4 (N14992, N14978, N13191, N13699, N673);
buf BUF1 (N14993, N14984);
not NOT1 (N14994, N14988);
xor XOR2 (N14995, N14981, N12244);
nor NOR2 (N14996, N14987, N1476);
nor NOR4 (N14997, N14990, N6970, N13546, N559);
nor NOR3 (N14998, N14991, N7674, N5071);
and AND3 (N14999, N14966, N9022, N9892);
nand NAND2 (N15000, N14989, N12931);
nand NAND2 (N15001, N14995, N12086);
xor XOR2 (N15002, N14994, N14689);
and AND4 (N15003, N15001, N11155, N13537, N3808);
or OR3 (N15004, N14997, N10705, N5886);
and AND4 (N15005, N15002, N2622, N921, N1745);
buf BUF1 (N15006, N14996);
and AND2 (N15007, N14998, N12375);
and AND3 (N15008, N15006, N13463, N12829);
not NOT1 (N15009, N15000);
or OR4 (N15010, N14999, N14473, N11294, N12337);
nor NOR2 (N15011, N15004, N4191);
nand NAND4 (N15012, N15008, N2889, N7731, N2577);
nor NOR3 (N15013, N15010, N6933, N2645);
nand NAND3 (N15014, N15007, N6970, N5767);
nand NAND4 (N15015, N15005, N5497, N6032, N6743);
nor NOR3 (N15016, N15011, N640, N3083);
nor NOR3 (N15017, N15016, N14547, N10772);
nand NAND2 (N15018, N14993, N9802);
or OR4 (N15019, N15012, N2557, N11426, N9274);
nand NAND2 (N15020, N15019, N5383);
xor XOR2 (N15021, N15014, N11603);
xor XOR2 (N15022, N15017, N7131);
xor XOR2 (N15023, N15015, N7058);
xor XOR2 (N15024, N15013, N8476);
not NOT1 (N15025, N15024);
buf BUF1 (N15026, N15003);
or OR3 (N15027, N15009, N9295, N3033);
nor NOR3 (N15028, N15018, N10656, N1658);
nor NOR3 (N15029, N15025, N7232, N1167);
or OR3 (N15030, N15022, N4604, N2061);
not NOT1 (N15031, N15030);
and AND3 (N15032, N15021, N4321, N11272);
or OR3 (N15033, N15020, N5514, N14145);
buf BUF1 (N15034, N15031);
xor XOR2 (N15035, N14992, N13308);
and AND4 (N15036, N15035, N10480, N5697, N14304);
nand NAND2 (N15037, N15027, N665);
nand NAND2 (N15038, N15034, N7242);
nor NOR4 (N15039, N15038, N10674, N3165, N5597);
or OR3 (N15040, N15029, N4971, N3873);
nand NAND4 (N15041, N15040, N2281, N5147, N9032);
or OR2 (N15042, N15039, N7479);
xor XOR2 (N15043, N15026, N14215);
nand NAND3 (N15044, N15037, N12300, N7387);
buf BUF1 (N15045, N14985);
nand NAND2 (N15046, N15032, N1933);
buf BUF1 (N15047, N15033);
nor NOR4 (N15048, N15041, N10052, N9298, N3111);
or OR2 (N15049, N15044, N7294);
or OR3 (N15050, N15028, N3593, N14482);
nand NAND2 (N15051, N15023, N1445);
xor XOR2 (N15052, N15047, N9848);
buf BUF1 (N15053, N15048);
or OR4 (N15054, N15046, N8384, N7193, N6923);
buf BUF1 (N15055, N15049);
not NOT1 (N15056, N15043);
buf BUF1 (N15057, N15052);
nor NOR4 (N15058, N15053, N14861, N471, N2655);
or OR2 (N15059, N15042, N7646);
xor XOR2 (N15060, N15051, N3792);
and AND2 (N15061, N15036, N794);
or OR3 (N15062, N15060, N10295, N9967);
nor NOR4 (N15063, N15055, N9840, N6915, N6685);
and AND2 (N15064, N15050, N5704);
and AND4 (N15065, N15056, N11646, N6780, N7870);
buf BUF1 (N15066, N15045);
or OR4 (N15067, N15054, N9438, N7239, N4102);
not NOT1 (N15068, N15059);
or OR4 (N15069, N15067, N7500, N14925, N3447);
or OR4 (N15070, N15065, N8036, N257, N13186);
nand NAND3 (N15071, N15061, N2511, N13351);
and AND2 (N15072, N15071, N4127);
nand NAND2 (N15073, N15068, N8792);
nand NAND2 (N15074, N15073, N935);
or OR4 (N15075, N15066, N4994, N9386, N12276);
nor NOR2 (N15076, N15075, N2810);
nand NAND4 (N15077, N15069, N9761, N12261, N12361);
buf BUF1 (N15078, N15064);
or OR2 (N15079, N15063, N2914);
nand NAND2 (N15080, N15058, N10543);
nand NAND4 (N15081, N15079, N10306, N4051, N8914);
buf BUF1 (N15082, N15080);
xor XOR2 (N15083, N15057, N10160);
not NOT1 (N15084, N15077);
xor XOR2 (N15085, N15062, N4199);
not NOT1 (N15086, N15085);
buf BUF1 (N15087, N15076);
nand NAND4 (N15088, N15072, N10971, N8687, N11350);
nand NAND4 (N15089, N15086, N6977, N9924, N8514);
or OR2 (N15090, N15089, N8195);
or OR3 (N15091, N15070, N14412, N14296);
not NOT1 (N15092, N15083);
xor XOR2 (N15093, N15088, N6899);
xor XOR2 (N15094, N15092, N11069);
nand NAND3 (N15095, N15094, N13908, N12948);
nor NOR3 (N15096, N15091, N10356, N14299);
xor XOR2 (N15097, N15082, N6271);
nand NAND4 (N15098, N15084, N8778, N12326, N13283);
buf BUF1 (N15099, N15074);
and AND2 (N15100, N15095, N13894);
not NOT1 (N15101, N15100);
nand NAND4 (N15102, N15081, N14697, N1677, N7094);
xor XOR2 (N15103, N15102, N6953);
xor XOR2 (N15104, N15096, N8719);
or OR4 (N15105, N15101, N12990, N2596, N7547);
nand NAND2 (N15106, N15098, N10011);
nand NAND2 (N15107, N15103, N9004);
nand NAND4 (N15108, N15093, N1719, N6816, N6370);
nand NAND4 (N15109, N15090, N10945, N9504, N8695);
or OR3 (N15110, N15106, N8255, N1629);
and AND4 (N15111, N15108, N3875, N2515, N5643);
or OR4 (N15112, N15111, N14041, N11534, N9480);
xor XOR2 (N15113, N15097, N13696);
nor NOR2 (N15114, N15107, N9237);
or OR4 (N15115, N15109, N7233, N5754, N1584);
nor NOR4 (N15116, N15112, N8547, N2175, N10195);
xor XOR2 (N15117, N15113, N404);
buf BUF1 (N15118, N15104);
nand NAND2 (N15119, N15099, N5299);
buf BUF1 (N15120, N15105);
or OR4 (N15121, N15115, N9498, N2859, N3461);
nand NAND3 (N15122, N15119, N14470, N10358);
buf BUF1 (N15123, N15114);
buf BUF1 (N15124, N15118);
nand NAND4 (N15125, N15078, N10989, N11161, N8086);
not NOT1 (N15126, N15123);
nand NAND2 (N15127, N15124, N1817);
nor NOR3 (N15128, N15121, N529, N11380);
not NOT1 (N15129, N15117);
and AND4 (N15130, N15087, N7355, N9939, N6025);
or OR2 (N15131, N15116, N7154);
or OR4 (N15132, N15131, N2255, N13860, N4563);
not NOT1 (N15133, N15129);
or OR3 (N15134, N15110, N3409, N1133);
xor XOR2 (N15135, N15132, N1529);
nor NOR4 (N15136, N15133, N4060, N4083, N4126);
or OR3 (N15137, N15125, N1244, N1733);
xor XOR2 (N15138, N15120, N14785);
nor NOR2 (N15139, N15138, N14802);
or OR3 (N15140, N15126, N9875, N11683);
nor NOR3 (N15141, N15136, N2145, N7924);
not NOT1 (N15142, N15127);
or OR3 (N15143, N15140, N15088, N9117);
nand NAND4 (N15144, N15122, N9622, N12844, N10335);
and AND3 (N15145, N15139, N5319, N10960);
and AND3 (N15146, N15128, N7326, N5525);
and AND3 (N15147, N15141, N2736, N5222);
and AND3 (N15148, N15144, N8627, N12910);
or OR4 (N15149, N15145, N3695, N13270, N1498);
xor XOR2 (N15150, N15130, N12540);
nor NOR2 (N15151, N15137, N7609);
buf BUF1 (N15152, N15147);
or OR2 (N15153, N15151, N1705);
nand NAND4 (N15154, N15149, N11242, N7463, N5458);
or OR4 (N15155, N15142, N2375, N4399, N1735);
and AND3 (N15156, N15148, N8974, N5195);
xor XOR2 (N15157, N15156, N12085);
not NOT1 (N15158, N15154);
nand NAND2 (N15159, N15135, N5307);
buf BUF1 (N15160, N15143);
xor XOR2 (N15161, N15153, N13668);
xor XOR2 (N15162, N15158, N5001);
xor XOR2 (N15163, N15160, N12626);
not NOT1 (N15164, N15150);
and AND4 (N15165, N15163, N1351, N3191, N13598);
and AND2 (N15166, N15134, N13138);
nand NAND2 (N15167, N15161, N3001);
and AND2 (N15168, N15167, N2625);
not NOT1 (N15169, N15155);
not NOT1 (N15170, N15166);
nor NOR3 (N15171, N15152, N4561, N14197);
nand NAND4 (N15172, N15170, N3492, N3067, N4855);
xor XOR2 (N15173, N15169, N9670);
nand NAND2 (N15174, N15172, N6478);
xor XOR2 (N15175, N15162, N11737);
xor XOR2 (N15176, N15165, N11050);
nor NOR4 (N15177, N15174, N9334, N12877, N1834);
not NOT1 (N15178, N15171);
nand NAND2 (N15179, N15173, N12208);
not NOT1 (N15180, N15168);
nor NOR3 (N15181, N15164, N9181, N8850);
and AND3 (N15182, N15146, N14027, N6754);
buf BUF1 (N15183, N15159);
nor NOR3 (N15184, N15182, N14266, N9284);
or OR3 (N15185, N15179, N10842, N2839);
and AND2 (N15186, N15177, N10888);
or OR3 (N15187, N15178, N1291, N1734);
nor NOR4 (N15188, N15183, N3466, N14867, N4906);
not NOT1 (N15189, N15184);
buf BUF1 (N15190, N15181);
nand NAND4 (N15191, N15189, N2958, N716, N6195);
xor XOR2 (N15192, N15190, N13394);
nor NOR2 (N15193, N15157, N67);
not NOT1 (N15194, N15185);
nor NOR4 (N15195, N15191, N11929, N7314, N703);
not NOT1 (N15196, N15195);
buf BUF1 (N15197, N15186);
nor NOR4 (N15198, N15176, N6614, N10521, N12001);
nor NOR2 (N15199, N15193, N496);
or OR2 (N15200, N15199, N13010);
nand NAND2 (N15201, N15188, N13781);
or OR4 (N15202, N15175, N2939, N887, N4958);
not NOT1 (N15203, N15200);
not NOT1 (N15204, N15197);
not NOT1 (N15205, N15204);
nand NAND2 (N15206, N15201, N3406);
not NOT1 (N15207, N15202);
xor XOR2 (N15208, N15196, N1726);
and AND4 (N15209, N15192, N2479, N8490, N14446);
not NOT1 (N15210, N15207);
not NOT1 (N15211, N15209);
nor NOR4 (N15212, N15205, N9006, N13732, N315);
nand NAND2 (N15213, N15206, N4680);
not NOT1 (N15214, N15203);
nand NAND3 (N15215, N15187, N2716, N842);
or OR4 (N15216, N15214, N13055, N6431, N1872);
nand NAND3 (N15217, N15213, N3654, N3442);
nand NAND4 (N15218, N15198, N8040, N2133, N1130);
xor XOR2 (N15219, N15208, N11300);
nor NOR3 (N15220, N15211, N6114, N8602);
buf BUF1 (N15221, N15220);
not NOT1 (N15222, N15218);
or OR2 (N15223, N15180, N1947);
not NOT1 (N15224, N15216);
nand NAND3 (N15225, N15219, N6027, N13674);
not NOT1 (N15226, N15217);
nand NAND4 (N15227, N15221, N5021, N441, N12952);
or OR2 (N15228, N15222, N66);
not NOT1 (N15229, N15215);
nor NOR4 (N15230, N15225, N2909, N11038, N12534);
xor XOR2 (N15231, N15212, N3292);
nor NOR3 (N15232, N15194, N4507, N2684);
xor XOR2 (N15233, N15227, N3596);
not NOT1 (N15234, N15223);
nor NOR4 (N15235, N15234, N5860, N4091, N12269);
nand NAND4 (N15236, N15228, N10701, N9994, N1587);
buf BUF1 (N15237, N15230);
nand NAND3 (N15238, N15231, N8052, N11265);
nor NOR3 (N15239, N15224, N2895, N7315);
or OR2 (N15240, N15239, N10502);
xor XOR2 (N15241, N15235, N13659);
or OR3 (N15242, N15229, N5060, N854);
xor XOR2 (N15243, N15240, N13138);
not NOT1 (N15244, N15232);
buf BUF1 (N15245, N15210);
and AND4 (N15246, N15238, N780, N9498, N11875);
or OR4 (N15247, N15237, N10044, N8488, N14265);
and AND4 (N15248, N15244, N3248, N5974, N11823);
and AND2 (N15249, N15242, N15189);
not NOT1 (N15250, N15236);
nor NOR2 (N15251, N15226, N14774);
nand NAND2 (N15252, N15250, N5017);
or OR2 (N15253, N15243, N7666);
nor NOR4 (N15254, N15248, N3527, N3910, N7054);
and AND2 (N15255, N15254, N2489);
and AND2 (N15256, N15251, N7537);
xor XOR2 (N15257, N15247, N3326);
xor XOR2 (N15258, N15246, N2257);
nand NAND4 (N15259, N15253, N1645, N4759, N7641);
and AND2 (N15260, N15249, N8505);
nor NOR3 (N15261, N15258, N10419, N6793);
nand NAND3 (N15262, N15261, N652, N5455);
and AND4 (N15263, N15260, N10258, N1361, N10571);
xor XOR2 (N15264, N15256, N7346);
or OR4 (N15265, N15233, N7178, N234, N5349);
xor XOR2 (N15266, N15262, N6087);
nand NAND2 (N15267, N15257, N9121);
or OR2 (N15268, N15264, N7051);
nor NOR3 (N15269, N15267, N3354, N13483);
not NOT1 (N15270, N15269);
or OR2 (N15271, N15252, N8090);
and AND3 (N15272, N15241, N8328, N12268);
and AND4 (N15273, N15272, N13105, N9344, N7565);
nor NOR2 (N15274, N15265, N14120);
nand NAND2 (N15275, N15263, N5586);
and AND2 (N15276, N15274, N10307);
xor XOR2 (N15277, N15275, N10078);
buf BUF1 (N15278, N15268);
or OR4 (N15279, N15266, N6027, N862, N596);
buf BUF1 (N15280, N15259);
nor NOR3 (N15281, N15277, N6619, N13185);
buf BUF1 (N15282, N15255);
nand NAND2 (N15283, N15276, N4632);
xor XOR2 (N15284, N15278, N13541);
buf BUF1 (N15285, N15282);
xor XOR2 (N15286, N15245, N2336);
and AND4 (N15287, N15271, N11382, N4957, N10318);
nand NAND3 (N15288, N15287, N7879, N14189);
not NOT1 (N15289, N15281);
nor NOR4 (N15290, N15288, N4194, N2466, N13958);
nand NAND2 (N15291, N15279, N8580);
nand NAND4 (N15292, N15273, N159, N3714, N11046);
or OR3 (N15293, N15289, N5361, N4319);
nand NAND3 (N15294, N15285, N5819, N1384);
or OR3 (N15295, N15286, N2485, N3519);
and AND2 (N15296, N15292, N12001);
nand NAND4 (N15297, N15295, N3357, N5546, N9435);
not NOT1 (N15298, N15294);
nor NOR4 (N15299, N15291, N8328, N2048, N14859);
nand NAND3 (N15300, N15284, N5858, N14419);
nor NOR4 (N15301, N15299, N1956, N13919, N12605);
xor XOR2 (N15302, N15296, N1260);
and AND3 (N15303, N15290, N14116, N12960);
nor NOR3 (N15304, N15300, N2198, N5489);
not NOT1 (N15305, N15302);
nand NAND3 (N15306, N15293, N5349, N6668);
buf BUF1 (N15307, N15301);
xor XOR2 (N15308, N15283, N13484);
or OR2 (N15309, N15298, N14112);
or OR2 (N15310, N15307, N7611);
xor XOR2 (N15311, N15297, N5007);
or OR2 (N15312, N15310, N7592);
and AND4 (N15313, N15306, N9170, N12359, N9692);
nand NAND3 (N15314, N15305, N8768, N8126);
nor NOR2 (N15315, N15314, N1252);
xor XOR2 (N15316, N15309, N4996);
not NOT1 (N15317, N15308);
and AND4 (N15318, N15280, N11095, N11208, N12182);
or OR4 (N15319, N15315, N2408, N264, N10898);
and AND4 (N15320, N15312, N3926, N1793, N6616);
xor XOR2 (N15321, N15317, N7201);
not NOT1 (N15322, N15320);
buf BUF1 (N15323, N15311);
not NOT1 (N15324, N15323);
xor XOR2 (N15325, N15316, N10898);
or OR4 (N15326, N15324, N7735, N5212, N14258);
nand NAND3 (N15327, N15270, N57, N9543);
or OR3 (N15328, N15322, N5053, N1777);
nor NOR3 (N15329, N15303, N4645, N9369);
buf BUF1 (N15330, N15321);
and AND2 (N15331, N15313, N271);
and AND4 (N15332, N15327, N6551, N7486, N3434);
nand NAND4 (N15333, N15304, N13447, N9737, N8632);
not NOT1 (N15334, N15333);
xor XOR2 (N15335, N15332, N4492);
or OR3 (N15336, N15331, N7226, N13694);
and AND4 (N15337, N15318, N4653, N7772, N12653);
buf BUF1 (N15338, N15328);
and AND2 (N15339, N15319, N7190);
nand NAND3 (N15340, N15334, N5690, N12854);
nand NAND3 (N15341, N15338, N799, N6679);
nand NAND2 (N15342, N15340, N5810);
nor NOR3 (N15343, N15341, N10705, N14881);
xor XOR2 (N15344, N15342, N14234);
buf BUF1 (N15345, N15343);
nand NAND2 (N15346, N15337, N3101);
or OR4 (N15347, N15344, N9123, N14472, N8074);
not NOT1 (N15348, N15335);
nand NAND4 (N15349, N15330, N7166, N409, N11572);
not NOT1 (N15350, N15348);
not NOT1 (N15351, N15336);
buf BUF1 (N15352, N15339);
nor NOR4 (N15353, N15345, N15140, N11519, N11037);
nand NAND3 (N15354, N15349, N14092, N1912);
not NOT1 (N15355, N15346);
nor NOR2 (N15356, N15355, N13633);
and AND4 (N15357, N15352, N1639, N12538, N14074);
and AND2 (N15358, N15326, N6459);
nand NAND4 (N15359, N15329, N14719, N5534, N5421);
nand NAND2 (N15360, N15358, N11813);
nand NAND4 (N15361, N15351, N775, N3891, N12688);
nand NAND2 (N15362, N15360, N6258);
nor NOR2 (N15363, N15354, N13826);
nor NOR3 (N15364, N15325, N7739, N7564);
buf BUF1 (N15365, N15362);
and AND2 (N15366, N15353, N12347);
or OR4 (N15367, N15359, N1627, N15132, N2333);
and AND2 (N15368, N15350, N12113);
not NOT1 (N15369, N15363);
or OR2 (N15370, N15368, N5727);
and AND2 (N15371, N15357, N6048);
nand NAND4 (N15372, N15371, N11739, N2123, N5274);
nor NOR4 (N15373, N15365, N11607, N6312, N11133);
buf BUF1 (N15374, N15364);
not NOT1 (N15375, N15367);
or OR3 (N15376, N15366, N2905, N11619);
nor NOR3 (N15377, N15347, N5946, N4601);
nand NAND2 (N15378, N15370, N1162);
xor XOR2 (N15379, N15375, N7971);
nand NAND4 (N15380, N15374, N11348, N5624, N7742);
and AND2 (N15381, N15379, N982);
not NOT1 (N15382, N15369);
nor NOR4 (N15383, N15376, N626, N5281, N10154);
nand NAND2 (N15384, N15361, N7943);
buf BUF1 (N15385, N15373);
or OR2 (N15386, N15385, N11336);
nand NAND4 (N15387, N15378, N2809, N7286, N14141);
nor NOR2 (N15388, N15356, N14257);
nor NOR4 (N15389, N15381, N1122, N704, N3210);
nor NOR2 (N15390, N15384, N4327);
not NOT1 (N15391, N15390);
nand NAND3 (N15392, N15387, N1269, N6946);
nand NAND2 (N15393, N15392, N6540);
nor NOR2 (N15394, N15393, N139);
and AND3 (N15395, N15386, N13751, N12025);
not NOT1 (N15396, N15391);
or OR4 (N15397, N15395, N14568, N4502, N6680);
and AND2 (N15398, N15380, N235);
not NOT1 (N15399, N15398);
buf BUF1 (N15400, N15389);
and AND3 (N15401, N15383, N3287, N669);
xor XOR2 (N15402, N15399, N13872);
xor XOR2 (N15403, N15400, N11695);
nand NAND4 (N15404, N15394, N2011, N12839, N444);
xor XOR2 (N15405, N15401, N14647);
not NOT1 (N15406, N15403);
not NOT1 (N15407, N15404);
not NOT1 (N15408, N15377);
nor NOR2 (N15409, N15397, N7934);
nand NAND2 (N15410, N15372, N13048);
nand NAND2 (N15411, N15396, N6540);
nand NAND2 (N15412, N15388, N7387);
nor NOR3 (N15413, N15402, N8697, N6963);
nor NOR3 (N15414, N15411, N13887, N12534);
or OR2 (N15415, N15413, N12948);
or OR3 (N15416, N15382, N13326, N7308);
buf BUF1 (N15417, N15407);
buf BUF1 (N15418, N15414);
and AND3 (N15419, N15410, N6058, N14548);
nand NAND3 (N15420, N15415, N8067, N1217);
or OR3 (N15421, N15419, N8239, N10846);
and AND2 (N15422, N15409, N9291);
not NOT1 (N15423, N15406);
buf BUF1 (N15424, N15416);
not NOT1 (N15425, N15423);
nor NOR4 (N15426, N15412, N2390, N10421, N5610);
and AND3 (N15427, N15425, N745, N3177);
and AND3 (N15428, N15422, N5650, N15036);
xor XOR2 (N15429, N15427, N3792);
not NOT1 (N15430, N15426);
or OR4 (N15431, N15421, N8712, N6719, N14486);
xor XOR2 (N15432, N15420, N7391);
and AND3 (N15433, N15408, N1641, N3471);
and AND3 (N15434, N15431, N7, N4238);
buf BUF1 (N15435, N15424);
buf BUF1 (N15436, N15428);
or OR3 (N15437, N15432, N1796, N1852);
nand NAND4 (N15438, N15437, N9793, N3246, N3097);
or OR2 (N15439, N15418, N9318);
or OR4 (N15440, N15434, N12231, N8782, N13703);
nor NOR3 (N15441, N15439, N4997, N7170);
nand NAND3 (N15442, N15435, N3788, N12828);
xor XOR2 (N15443, N15405, N6568);
nor NOR3 (N15444, N15436, N13954, N1113);
and AND4 (N15445, N15433, N5244, N7670, N2366);
nand NAND3 (N15446, N15430, N2619, N9512);
or OR3 (N15447, N15445, N7271, N14699);
xor XOR2 (N15448, N15440, N10326);
nor NOR2 (N15449, N15429, N4471);
or OR3 (N15450, N15441, N7006, N4095);
nor NOR3 (N15451, N15446, N4040, N12500);
nand NAND3 (N15452, N15447, N13077, N14991);
nand NAND2 (N15453, N15451, N3908);
or OR2 (N15454, N15444, N5147);
nor NOR4 (N15455, N15452, N568, N1778, N13212);
or OR2 (N15456, N15442, N8268);
nor NOR2 (N15457, N15455, N7564);
nor NOR4 (N15458, N15457, N6024, N10809, N14141);
buf BUF1 (N15459, N15443);
not NOT1 (N15460, N15417);
xor XOR2 (N15461, N15454, N3915);
nor NOR3 (N15462, N15453, N13865, N859);
not NOT1 (N15463, N15450);
buf BUF1 (N15464, N15459);
xor XOR2 (N15465, N15458, N3519);
not NOT1 (N15466, N15449);
not NOT1 (N15467, N15462);
and AND4 (N15468, N15464, N12878, N15337, N8614);
or OR2 (N15469, N15448, N10190);
not NOT1 (N15470, N15456);
nor NOR3 (N15471, N15469, N10026, N13634);
or OR4 (N15472, N15438, N3965, N352, N3018);
nor NOR4 (N15473, N15465, N13006, N8492, N13798);
and AND4 (N15474, N15473, N1994, N2441, N6794);
and AND3 (N15475, N15460, N8302, N7816);
buf BUF1 (N15476, N15474);
nand NAND2 (N15477, N15468, N219);
and AND4 (N15478, N15471, N4368, N1122, N4813);
buf BUF1 (N15479, N15466);
not NOT1 (N15480, N15472);
or OR3 (N15481, N15477, N13516, N2874);
buf BUF1 (N15482, N15476);
nor NOR2 (N15483, N15481, N5404);
and AND3 (N15484, N15461, N4076, N1861);
nand NAND3 (N15485, N15480, N3567, N6247);
and AND3 (N15486, N15463, N14441, N14884);
buf BUF1 (N15487, N15482);
nand NAND4 (N15488, N15470, N5860, N9620, N11751);
not NOT1 (N15489, N15467);
xor XOR2 (N15490, N15484, N3893);
buf BUF1 (N15491, N15483);
not NOT1 (N15492, N15491);
buf BUF1 (N15493, N15479);
nor NOR3 (N15494, N15488, N4917, N10976);
or OR2 (N15495, N15486, N256);
nor NOR3 (N15496, N15494, N9677, N7216);
nand NAND3 (N15497, N15487, N12693, N9691);
or OR3 (N15498, N15490, N12014, N13883);
nand NAND2 (N15499, N15485, N12137);
or OR4 (N15500, N15496, N7923, N3732, N7087);
nand NAND3 (N15501, N15489, N6224, N7284);
xor XOR2 (N15502, N15501, N8014);
and AND3 (N15503, N15499, N4489, N9355);
xor XOR2 (N15504, N15497, N6795);
or OR4 (N15505, N15498, N2640, N12896, N8336);
xor XOR2 (N15506, N15478, N8512);
and AND2 (N15507, N15504, N9377);
xor XOR2 (N15508, N15503, N1273);
xor XOR2 (N15509, N15506, N14259);
xor XOR2 (N15510, N15507, N7148);
or OR3 (N15511, N15500, N12878, N5117);
not NOT1 (N15512, N15493);
nor NOR3 (N15513, N15510, N11048, N10096);
and AND2 (N15514, N15505, N9971);
not NOT1 (N15515, N15514);
xor XOR2 (N15516, N15509, N10269);
nor NOR4 (N15517, N15502, N8262, N15287, N12749);
nor NOR3 (N15518, N15495, N12311, N8322);
or OR4 (N15519, N15517, N7628, N14828, N3244);
not NOT1 (N15520, N15519);
or OR2 (N15521, N15508, N5825);
nor NOR3 (N15522, N15520, N2815, N12451);
buf BUF1 (N15523, N15522);
nand NAND3 (N15524, N15515, N15293, N5446);
not NOT1 (N15525, N15475);
not NOT1 (N15526, N15513);
nor NOR3 (N15527, N15523, N5737, N11185);
xor XOR2 (N15528, N15521, N4813);
not NOT1 (N15529, N15525);
or OR4 (N15530, N15526, N7550, N6585, N7788);
or OR3 (N15531, N15492, N6998, N8931);
xor XOR2 (N15532, N15512, N1368);
nor NOR2 (N15533, N15516, N7705);
not NOT1 (N15534, N15532);
buf BUF1 (N15535, N15534);
nor NOR4 (N15536, N15511, N435, N7516, N10875);
xor XOR2 (N15537, N15528, N4188);
not NOT1 (N15538, N15533);
nand NAND4 (N15539, N15529, N11768, N8553, N8949);
buf BUF1 (N15540, N15537);
nand NAND4 (N15541, N15535, N1791, N8048, N244);
nor NOR2 (N15542, N15538, N3971);
nor NOR2 (N15543, N15527, N7053);
nor NOR2 (N15544, N15518, N11532);
and AND3 (N15545, N15541, N12701, N14453);
or OR2 (N15546, N15524, N8848);
not NOT1 (N15547, N15530);
nor NOR2 (N15548, N15544, N9055);
not NOT1 (N15549, N15536);
nor NOR2 (N15550, N15540, N11007);
or OR4 (N15551, N15547, N2048, N13287, N5590);
nand NAND4 (N15552, N15545, N6845, N11665, N7163);
nand NAND2 (N15553, N15542, N523);
xor XOR2 (N15554, N15551, N9421);
not NOT1 (N15555, N15548);
xor XOR2 (N15556, N15553, N693);
and AND3 (N15557, N15539, N3831, N12158);
and AND4 (N15558, N15550, N8344, N10222, N7221);
nand NAND2 (N15559, N15543, N14507);
nand NAND2 (N15560, N15557, N1438);
and AND3 (N15561, N15531, N10712, N15281);
and AND2 (N15562, N15558, N1416);
and AND4 (N15563, N15561, N4041, N4443, N10869);
xor XOR2 (N15564, N15562, N5854);
or OR4 (N15565, N15559, N1890, N15412, N10150);
nor NOR2 (N15566, N15556, N7175);
nand NAND4 (N15567, N15546, N2789, N2074, N1249);
nand NAND4 (N15568, N15565, N14167, N7422, N7517);
nand NAND4 (N15569, N15566, N8008, N4568, N4638);
and AND2 (N15570, N15554, N4862);
and AND4 (N15571, N15560, N2799, N13373, N839);
buf BUF1 (N15572, N15567);
nor NOR4 (N15573, N15569, N6698, N1334, N90);
buf BUF1 (N15574, N15572);
xor XOR2 (N15575, N15555, N2255);
and AND2 (N15576, N15552, N11598);
buf BUF1 (N15577, N15574);
and AND4 (N15578, N15575, N5416, N4697, N1548);
nand NAND2 (N15579, N15577, N15071);
buf BUF1 (N15580, N15576);
and AND2 (N15581, N15580, N14685);
xor XOR2 (N15582, N15573, N15231);
buf BUF1 (N15583, N15571);
or OR3 (N15584, N15579, N13641, N2578);
xor XOR2 (N15585, N15584, N11388);
nor NOR4 (N15586, N15549, N14786, N173, N3901);
xor XOR2 (N15587, N15578, N14827);
nor NOR4 (N15588, N15585, N10087, N3850, N9488);
nand NAND3 (N15589, N15586, N3597, N3953);
not NOT1 (N15590, N15588);
or OR3 (N15591, N15583, N5674, N2156);
or OR3 (N15592, N15582, N10304, N7516);
not NOT1 (N15593, N15564);
nor NOR2 (N15594, N15589, N1810);
or OR2 (N15595, N15563, N11115);
nor NOR3 (N15596, N15587, N10312, N3498);
buf BUF1 (N15597, N15591);
xor XOR2 (N15598, N15592, N1609);
xor XOR2 (N15599, N15590, N3045);
or OR2 (N15600, N15568, N8259);
nor NOR2 (N15601, N15600, N4901);
or OR2 (N15602, N15593, N2528);
nand NAND3 (N15603, N15598, N6235, N695);
nor NOR2 (N15604, N15602, N9021);
nor NOR2 (N15605, N15599, N3837);
or OR4 (N15606, N15594, N10743, N2195, N10112);
nor NOR2 (N15607, N15603, N10681);
buf BUF1 (N15608, N15604);
buf BUF1 (N15609, N15581);
nand NAND2 (N15610, N15601, N12430);
nor NOR2 (N15611, N15605, N9404);
xor XOR2 (N15612, N15609, N5906);
xor XOR2 (N15613, N15610, N9413);
and AND2 (N15614, N15611, N545);
nand NAND3 (N15615, N15596, N12496, N2619);
or OR4 (N15616, N15612, N6305, N6455, N11746);
nand NAND4 (N15617, N15615, N11973, N12278, N2695);
nand NAND3 (N15618, N15608, N1934, N13678);
and AND3 (N15619, N15597, N284, N4507);
nor NOR2 (N15620, N15595, N5811);
and AND2 (N15621, N15570, N15001);
not NOT1 (N15622, N15617);
nand NAND3 (N15623, N15620, N8537, N11143);
not NOT1 (N15624, N15619);
xor XOR2 (N15625, N15616, N2341);
xor XOR2 (N15626, N15618, N8672);
and AND3 (N15627, N15624, N4760, N10107);
or OR2 (N15628, N15627, N3446);
and AND2 (N15629, N15607, N3255);
or OR3 (N15630, N15626, N4302, N4132);
not NOT1 (N15631, N15613);
or OR4 (N15632, N15625, N783, N7231, N13442);
nor NOR4 (N15633, N15631, N3971, N2660, N10375);
nand NAND3 (N15634, N15630, N5026, N115);
and AND3 (N15635, N15614, N5179, N10984);
or OR2 (N15636, N15628, N2696);
buf BUF1 (N15637, N15621);
nand NAND3 (N15638, N15635, N865, N11094);
and AND4 (N15639, N15622, N6359, N443, N8855);
nor NOR2 (N15640, N15639, N5008);
nor NOR3 (N15641, N15637, N10318, N8607);
xor XOR2 (N15642, N15640, N1584);
or OR4 (N15643, N15636, N12565, N13904, N9838);
and AND4 (N15644, N15643, N8832, N10870, N15413);
and AND2 (N15645, N15641, N9487);
buf BUF1 (N15646, N15632);
not NOT1 (N15647, N15629);
nor NOR2 (N15648, N15606, N2563);
nor NOR4 (N15649, N15644, N951, N8393, N4533);
not NOT1 (N15650, N15638);
xor XOR2 (N15651, N15633, N9744);
buf BUF1 (N15652, N15623);
or OR3 (N15653, N15648, N3549, N6928);
buf BUF1 (N15654, N15642);
xor XOR2 (N15655, N15652, N10811);
nand NAND3 (N15656, N15651, N2984, N11567);
nand NAND3 (N15657, N15646, N15261, N3810);
xor XOR2 (N15658, N15647, N13815);
xor XOR2 (N15659, N15653, N8442);
nand NAND4 (N15660, N15658, N6206, N5264, N3872);
xor XOR2 (N15661, N15649, N13984);
buf BUF1 (N15662, N15660);
xor XOR2 (N15663, N15659, N4061);
xor XOR2 (N15664, N15656, N9716);
buf BUF1 (N15665, N15645);
xor XOR2 (N15666, N15650, N8501);
nor NOR4 (N15667, N15662, N7020, N4908, N10525);
nor NOR3 (N15668, N15667, N15436, N5772);
nor NOR3 (N15669, N15668, N6163, N6748);
buf BUF1 (N15670, N15665);
or OR2 (N15671, N15664, N13848);
nor NOR3 (N15672, N15654, N612, N5508);
or OR3 (N15673, N15634, N11736, N4235);
or OR3 (N15674, N15671, N3980, N8898);
xor XOR2 (N15675, N15663, N9573);
and AND4 (N15676, N15655, N370, N2489, N15589);
buf BUF1 (N15677, N15670);
xor XOR2 (N15678, N15661, N7500);
xor XOR2 (N15679, N15657, N3622);
or OR3 (N15680, N15675, N13042, N8269);
and AND4 (N15681, N15672, N11715, N7297, N8393);
nor NOR3 (N15682, N15680, N14000, N14804);
nor NOR3 (N15683, N15676, N3450, N5970);
or OR3 (N15684, N15669, N9228, N2059);
xor XOR2 (N15685, N15679, N5286);
not NOT1 (N15686, N15684);
nand NAND3 (N15687, N15678, N11366, N6235);
xor XOR2 (N15688, N15687, N12410);
and AND2 (N15689, N15681, N11);
nor NOR2 (N15690, N15673, N3994);
nand NAND4 (N15691, N15682, N12450, N15427, N7991);
nand NAND2 (N15692, N15691, N12245);
nor NOR3 (N15693, N15685, N9528, N6468);
and AND3 (N15694, N15683, N12037, N5483);
nand NAND4 (N15695, N15689, N14981, N9628, N14254);
nand NAND2 (N15696, N15686, N9300);
nand NAND4 (N15697, N15695, N8883, N14264, N5725);
nand NAND3 (N15698, N15696, N2473, N12640);
xor XOR2 (N15699, N15688, N1611);
buf BUF1 (N15700, N15692);
xor XOR2 (N15701, N15694, N14500);
or OR2 (N15702, N15677, N295);
xor XOR2 (N15703, N15666, N14976);
nand NAND4 (N15704, N15703, N12534, N7946, N9108);
not NOT1 (N15705, N15704);
buf BUF1 (N15706, N15700);
xor XOR2 (N15707, N15698, N7082);
xor XOR2 (N15708, N15706, N5607);
nor NOR3 (N15709, N15705, N14953, N1585);
not NOT1 (N15710, N15709);
or OR3 (N15711, N15674, N3131, N2168);
xor XOR2 (N15712, N15707, N14182);
buf BUF1 (N15713, N15702);
nor NOR4 (N15714, N15713, N15364, N9276, N3874);
or OR4 (N15715, N15711, N5315, N9812, N8280);
buf BUF1 (N15716, N15699);
xor XOR2 (N15717, N15716, N4857);
buf BUF1 (N15718, N15712);
xor XOR2 (N15719, N15693, N6238);
and AND2 (N15720, N15690, N3417);
and AND3 (N15721, N15718, N4564, N14435);
not NOT1 (N15722, N15715);
or OR4 (N15723, N15714, N12825, N13149, N10772);
buf BUF1 (N15724, N15710);
nor NOR4 (N15725, N15701, N338, N15503, N15493);
nand NAND4 (N15726, N15723, N4153, N3635, N12918);
buf BUF1 (N15727, N15697);
not NOT1 (N15728, N15720);
not NOT1 (N15729, N15719);
nand NAND3 (N15730, N15727, N14788, N10942);
nor NOR2 (N15731, N15730, N13524);
xor XOR2 (N15732, N15721, N1910);
xor XOR2 (N15733, N15725, N8614);
buf BUF1 (N15734, N15717);
buf BUF1 (N15735, N15722);
nand NAND4 (N15736, N15729, N2102, N3791, N4539);
not NOT1 (N15737, N15734);
and AND3 (N15738, N15726, N668, N7605);
and AND4 (N15739, N15724, N6609, N10450, N319);
and AND4 (N15740, N15733, N967, N15454, N8650);
xor XOR2 (N15741, N15735, N8233);
or OR2 (N15742, N15731, N10109);
and AND3 (N15743, N15728, N13471, N8556);
and AND2 (N15744, N15737, N7378);
or OR3 (N15745, N15732, N5385, N12759);
nand NAND4 (N15746, N15744, N13976, N15573, N13161);
nand NAND3 (N15747, N15745, N7141, N6807);
not NOT1 (N15748, N15708);
nor NOR4 (N15749, N15738, N13867, N3610, N15229);
nand NAND3 (N15750, N15739, N12321, N13017);
xor XOR2 (N15751, N15749, N10490);
nand NAND2 (N15752, N15742, N3978);
buf BUF1 (N15753, N15750);
not NOT1 (N15754, N15748);
or OR4 (N15755, N15741, N7415, N10206, N4659);
xor XOR2 (N15756, N15755, N12314);
buf BUF1 (N15757, N15747);
and AND2 (N15758, N15757, N8648);
and AND4 (N15759, N15754, N11141, N6463, N5021);
and AND4 (N15760, N15759, N10311, N10481, N13208);
nor NOR2 (N15761, N15746, N7427);
or OR3 (N15762, N15743, N2823, N12973);
nand NAND2 (N15763, N15753, N9858);
xor XOR2 (N15764, N15752, N13703);
not NOT1 (N15765, N15760);
nor NOR4 (N15766, N15762, N12614, N8751, N7756);
xor XOR2 (N15767, N15758, N2655);
not NOT1 (N15768, N15767);
or OR3 (N15769, N15751, N4578, N14308);
nor NOR3 (N15770, N15769, N7163, N13309);
not NOT1 (N15771, N15736);
and AND3 (N15772, N15763, N1389, N3913);
nor NOR4 (N15773, N15765, N10585, N8692, N7507);
nor NOR4 (N15774, N15756, N6262, N1732, N572);
nand NAND2 (N15775, N15770, N12374);
nor NOR4 (N15776, N15772, N11288, N12886, N11064);
and AND3 (N15777, N15768, N7631, N7011);
xor XOR2 (N15778, N15761, N11972);
not NOT1 (N15779, N15740);
nor NOR2 (N15780, N15778, N4764);
nand NAND2 (N15781, N15777, N13917);
or OR2 (N15782, N15764, N10802);
buf BUF1 (N15783, N15771);
not NOT1 (N15784, N15775);
xor XOR2 (N15785, N15784, N658);
not NOT1 (N15786, N15776);
xor XOR2 (N15787, N15782, N6258);
or OR2 (N15788, N15783, N12268);
or OR2 (N15789, N15773, N14538);
xor XOR2 (N15790, N15780, N372);
buf BUF1 (N15791, N15789);
nand NAND3 (N15792, N15787, N6113, N6015);
or OR3 (N15793, N15792, N2704, N13724);
nand NAND2 (N15794, N15766, N6778);
nand NAND3 (N15795, N15788, N5456, N13781);
or OR2 (N15796, N15785, N9799);
buf BUF1 (N15797, N15781);
or OR2 (N15798, N15793, N4719);
or OR2 (N15799, N15796, N762);
and AND3 (N15800, N15786, N8285, N7572);
or OR3 (N15801, N15798, N11847, N15387);
xor XOR2 (N15802, N15790, N7506);
not NOT1 (N15803, N15802);
and AND3 (N15804, N15774, N11883, N6618);
not NOT1 (N15805, N15800);
not NOT1 (N15806, N15805);
or OR4 (N15807, N15791, N2627, N8674, N10262);
xor XOR2 (N15808, N15801, N7143);
not NOT1 (N15809, N15795);
not NOT1 (N15810, N15794);
xor XOR2 (N15811, N15804, N7560);
nand NAND4 (N15812, N15809, N4985, N2365, N14384);
xor XOR2 (N15813, N15810, N448);
xor XOR2 (N15814, N15803, N1822);
not NOT1 (N15815, N15808);
not NOT1 (N15816, N15814);
and AND2 (N15817, N15806, N769);
or OR4 (N15818, N15812, N12253, N9585, N2141);
and AND4 (N15819, N15817, N6585, N4939, N5695);
and AND3 (N15820, N15811, N15663, N8166);
nor NOR4 (N15821, N15813, N15007, N7097, N2001);
buf BUF1 (N15822, N15820);
nand NAND4 (N15823, N15815, N1660, N7611, N14923);
and AND4 (N15824, N15819, N12594, N15706, N3659);
not NOT1 (N15825, N15821);
buf BUF1 (N15826, N15816);
buf BUF1 (N15827, N15826);
nor NOR2 (N15828, N15823, N3);
nand NAND2 (N15829, N15818, N5148);
buf BUF1 (N15830, N15829);
nor NOR3 (N15831, N15828, N6937, N3458);
or OR4 (N15832, N15827, N669, N14066, N13242);
buf BUF1 (N15833, N15807);
xor XOR2 (N15834, N15779, N6328);
and AND3 (N15835, N15797, N2319, N4482);
not NOT1 (N15836, N15834);
not NOT1 (N15837, N15836);
buf BUF1 (N15838, N15837);
xor XOR2 (N15839, N15833, N1922);
not NOT1 (N15840, N15831);
nor NOR3 (N15841, N15830, N551, N5414);
nor NOR2 (N15842, N15824, N4017);
buf BUF1 (N15843, N15840);
and AND2 (N15844, N15839, N6813);
xor XOR2 (N15845, N15841, N10636);
nand NAND3 (N15846, N15845, N859, N12786);
xor XOR2 (N15847, N15835, N5064);
or OR2 (N15848, N15843, N15830);
nand NAND4 (N15849, N15822, N13983, N2137, N4194);
and AND4 (N15850, N15799, N201, N3260, N9312);
nor NOR2 (N15851, N15846, N461);
and AND3 (N15852, N15849, N12934, N9064);
nand NAND3 (N15853, N15852, N3555, N3610);
xor XOR2 (N15854, N15853, N8559);
or OR4 (N15855, N15832, N6422, N551, N5455);
buf BUF1 (N15856, N15850);
buf BUF1 (N15857, N15851);
buf BUF1 (N15858, N15857);
xor XOR2 (N15859, N15855, N6516);
and AND4 (N15860, N15844, N9497, N8102, N3121);
nand NAND4 (N15861, N15825, N11947, N15265, N1214);
or OR2 (N15862, N15847, N991);
and AND4 (N15863, N15861, N3301, N964, N10848);
buf BUF1 (N15864, N15842);
or OR2 (N15865, N15863, N13030);
nor NOR4 (N15866, N15865, N10123, N10191, N12396);
not NOT1 (N15867, N15848);
xor XOR2 (N15868, N15854, N7736);
and AND2 (N15869, N15864, N13504);
nand NAND3 (N15870, N15862, N10944, N7535);
not NOT1 (N15871, N15856);
or OR3 (N15872, N15867, N5793, N15454);
or OR2 (N15873, N15838, N13851);
xor XOR2 (N15874, N15868, N13282);
nor NOR3 (N15875, N15859, N3154, N11737);
nor NOR3 (N15876, N15866, N9576, N4220);
nand NAND3 (N15877, N15875, N6721, N3821);
and AND3 (N15878, N15871, N5996, N3529);
nand NAND3 (N15879, N15873, N10655, N2444);
nor NOR2 (N15880, N15869, N4121);
and AND4 (N15881, N15870, N549, N8991, N15226);
nor NOR3 (N15882, N15878, N3632, N15365);
xor XOR2 (N15883, N15877, N10762);
nand NAND4 (N15884, N15858, N10376, N5258, N964);
and AND4 (N15885, N15876, N14729, N4838, N10183);
and AND3 (N15886, N15860, N5801, N14419);
nand NAND4 (N15887, N15886, N15632, N4533, N1303);
not NOT1 (N15888, N15883);
not NOT1 (N15889, N15881);
not NOT1 (N15890, N15887);
not NOT1 (N15891, N15884);
and AND4 (N15892, N15879, N9424, N10866, N6838);
xor XOR2 (N15893, N15891, N4950);
or OR2 (N15894, N15874, N5661);
not NOT1 (N15895, N15872);
or OR2 (N15896, N15890, N3300);
nor NOR4 (N15897, N15894, N14420, N3203, N309);
and AND4 (N15898, N15885, N14319, N5360, N13533);
xor XOR2 (N15899, N15882, N8285);
nand NAND3 (N15900, N15896, N5966, N5184);
not NOT1 (N15901, N15893);
not NOT1 (N15902, N15901);
buf BUF1 (N15903, N15902);
or OR2 (N15904, N15900, N6703);
not NOT1 (N15905, N15895);
buf BUF1 (N15906, N15897);
and AND2 (N15907, N15889, N8883);
not NOT1 (N15908, N15904);
or OR2 (N15909, N15908, N10407);
and AND3 (N15910, N15909, N5164, N10546);
xor XOR2 (N15911, N15892, N13145);
nor NOR3 (N15912, N15907, N4223, N1745);
buf BUF1 (N15913, N15911);
xor XOR2 (N15914, N15888, N2835);
nand NAND2 (N15915, N15906, N1181);
nor NOR3 (N15916, N15903, N7839, N546);
or OR2 (N15917, N15910, N668);
xor XOR2 (N15918, N15912, N11136);
nand NAND2 (N15919, N15913, N9171);
buf BUF1 (N15920, N15918);
and AND4 (N15921, N15917, N1299, N6917, N2551);
not NOT1 (N15922, N15898);
nor NOR4 (N15923, N15915, N3246, N13727, N11627);
nor NOR3 (N15924, N15914, N410, N14159);
nand NAND2 (N15925, N15905, N10843);
not NOT1 (N15926, N15924);
not NOT1 (N15927, N15920);
buf BUF1 (N15928, N15925);
xor XOR2 (N15929, N15926, N3289);
or OR4 (N15930, N15929, N2712, N11073, N2190);
or OR2 (N15931, N15880, N3509);
and AND4 (N15932, N15916, N3588, N338, N13061);
nor NOR3 (N15933, N15899, N5393, N7165);
or OR2 (N15934, N15931, N13118);
not NOT1 (N15935, N15923);
buf BUF1 (N15936, N15935);
or OR3 (N15937, N15928, N2956, N95);
buf BUF1 (N15938, N15932);
and AND3 (N15939, N15919, N13792, N10700);
xor XOR2 (N15940, N15921, N3581);
xor XOR2 (N15941, N15927, N5138);
and AND4 (N15942, N15936, N11060, N2497, N5482);
buf BUF1 (N15943, N15937);
buf BUF1 (N15944, N15941);
or OR2 (N15945, N15930, N13845);
buf BUF1 (N15946, N15942);
not NOT1 (N15947, N15933);
or OR3 (N15948, N15939, N36, N9178);
nand NAND2 (N15949, N15934, N4255);
buf BUF1 (N15950, N15949);
xor XOR2 (N15951, N15948, N1960);
xor XOR2 (N15952, N15922, N6214);
not NOT1 (N15953, N15946);
or OR2 (N15954, N15951, N1772);
not NOT1 (N15955, N15940);
xor XOR2 (N15956, N15943, N736);
nor NOR3 (N15957, N15945, N7890, N12447);
nand NAND2 (N15958, N15950, N13442);
or OR3 (N15959, N15955, N5975, N15815);
or OR2 (N15960, N15959, N86);
buf BUF1 (N15961, N15938);
xor XOR2 (N15962, N15960, N8780);
not NOT1 (N15963, N15944);
xor XOR2 (N15964, N15956, N4675);
and AND2 (N15965, N15953, N8437);
nor NOR3 (N15966, N15962, N15203, N4746);
not NOT1 (N15967, N15957);
and AND4 (N15968, N15961, N5946, N10395, N4567);
nand NAND3 (N15969, N15947, N14442, N27);
buf BUF1 (N15970, N15963);
nor NOR2 (N15971, N15969, N11906);
or OR3 (N15972, N15964, N15311, N11038);
xor XOR2 (N15973, N15967, N11936);
nor NOR3 (N15974, N15972, N15849, N10814);
not NOT1 (N15975, N15954);
nor NOR3 (N15976, N15952, N14227, N13988);
nor NOR2 (N15977, N15973, N11473);
nand NAND4 (N15978, N15970, N13698, N11908, N7173);
or OR2 (N15979, N15958, N14893);
or OR2 (N15980, N15968, N8146);
or OR4 (N15981, N15974, N1052, N6605, N13693);
not NOT1 (N15982, N15976);
nand NAND4 (N15983, N15971, N9655, N7887, N6414);
nand NAND4 (N15984, N15980, N6668, N10243, N14920);
nor NOR3 (N15985, N15983, N3334, N15061);
nand NAND4 (N15986, N15978, N9866, N2121, N5075);
xor XOR2 (N15987, N15986, N8591);
nor NOR2 (N15988, N15984, N15351);
and AND3 (N15989, N15985, N12351, N206);
or OR2 (N15990, N15965, N4622);
xor XOR2 (N15991, N15977, N4924);
xor XOR2 (N15992, N15979, N8575);
not NOT1 (N15993, N15981);
xor XOR2 (N15994, N15975, N14145);
and AND3 (N15995, N15994, N15810, N4806);
or OR2 (N15996, N15966, N8254);
xor XOR2 (N15997, N15989, N13735);
and AND2 (N15998, N15991, N2181);
not NOT1 (N15999, N15987);
nor NOR2 (N16000, N15999, N11258);
or OR2 (N16001, N16000, N12778);
or OR2 (N16002, N15995, N1063);
or OR2 (N16003, N15993, N13910);
or OR3 (N16004, N15992, N13119, N7272);
not NOT1 (N16005, N15997);
and AND3 (N16006, N16004, N4871, N12276);
buf BUF1 (N16007, N16003);
or OR3 (N16008, N15996, N1822, N14791);
xor XOR2 (N16009, N15982, N15239);
xor XOR2 (N16010, N16005, N9189);
buf BUF1 (N16011, N15998);
not NOT1 (N16012, N16011);
nor NOR4 (N16013, N16009, N12979, N15443, N15125);
nor NOR2 (N16014, N16008, N12540);
xor XOR2 (N16015, N15990, N9662);
not NOT1 (N16016, N16013);
buf BUF1 (N16017, N15988);
nor NOR2 (N16018, N16006, N12778);
nor NOR3 (N16019, N16015, N2743, N10165);
not NOT1 (N16020, N16016);
not NOT1 (N16021, N16017);
nand NAND2 (N16022, N16019, N1779);
xor XOR2 (N16023, N16018, N8351);
xor XOR2 (N16024, N16007, N14235);
xor XOR2 (N16025, N16021, N8212);
nand NAND3 (N16026, N16024, N4190, N15715);
buf BUF1 (N16027, N16002);
xor XOR2 (N16028, N16010, N13800);
and AND3 (N16029, N16001, N7349, N4281);
nand NAND3 (N16030, N16029, N7181, N9709);
buf BUF1 (N16031, N16025);
nand NAND3 (N16032, N16028, N8057, N433);
or OR3 (N16033, N16012, N13999, N10934);
not NOT1 (N16034, N16014);
nand NAND4 (N16035, N16031, N895, N11966, N8932);
xor XOR2 (N16036, N16032, N4042);
not NOT1 (N16037, N16027);
nand NAND3 (N16038, N16035, N555, N3051);
or OR3 (N16039, N16034, N655, N8740);
nand NAND2 (N16040, N16036, N11988);
and AND2 (N16041, N16026, N12099);
nor NOR2 (N16042, N16022, N4632);
or OR3 (N16043, N16030, N1311, N956);
nor NOR4 (N16044, N16023, N9397, N1398, N8571);
nor NOR2 (N16045, N16038, N10369);
and AND4 (N16046, N16044, N12881, N14589, N12197);
xor XOR2 (N16047, N16043, N14658);
xor XOR2 (N16048, N16042, N15442);
not NOT1 (N16049, N16048);
nand NAND4 (N16050, N16020, N3752, N5471, N1828);
buf BUF1 (N16051, N16033);
buf BUF1 (N16052, N16049);
xor XOR2 (N16053, N16051, N2505);
and AND2 (N16054, N16053, N1879);
or OR3 (N16055, N16050, N10608, N8944);
buf BUF1 (N16056, N16045);
nand NAND4 (N16057, N16037, N4116, N5331, N3110);
or OR2 (N16058, N16056, N10524);
or OR3 (N16059, N16039, N11143, N473);
buf BUF1 (N16060, N16054);
not NOT1 (N16061, N16055);
nor NOR4 (N16062, N16052, N13154, N2433, N9792);
nand NAND2 (N16063, N16040, N679);
nor NOR4 (N16064, N16046, N11887, N5385, N6563);
or OR3 (N16065, N16064, N647, N12351);
nand NAND3 (N16066, N16063, N3787, N3302);
or OR3 (N16067, N16060, N5555, N9293);
and AND3 (N16068, N16062, N5991, N8457);
not NOT1 (N16069, N16058);
nand NAND3 (N16070, N16069, N12164, N14757);
nand NAND2 (N16071, N16047, N5701);
and AND2 (N16072, N16059, N2130);
and AND3 (N16073, N16041, N6227, N1035);
and AND3 (N16074, N16067, N9485, N15257);
nand NAND4 (N16075, N16074, N8391, N7129, N9550);
buf BUF1 (N16076, N16075);
nor NOR3 (N16077, N16057, N10286, N14526);
xor XOR2 (N16078, N16072, N719);
nor NOR4 (N16079, N16073, N15287, N14976, N2788);
nor NOR3 (N16080, N16077, N10322, N12879);
not NOT1 (N16081, N16070);
xor XOR2 (N16082, N16080, N3865);
buf BUF1 (N16083, N16071);
xor XOR2 (N16084, N16082, N8338);
or OR2 (N16085, N16079, N13064);
nor NOR2 (N16086, N16081, N12475);
and AND3 (N16087, N16076, N4012, N1181);
or OR2 (N16088, N16078, N2868);
nand NAND4 (N16089, N16085, N10461, N6042, N5348);
and AND2 (N16090, N16088, N6275);
and AND2 (N16091, N16090, N2675);
buf BUF1 (N16092, N16089);
nor NOR3 (N16093, N16068, N6422, N10553);
nand NAND2 (N16094, N16086, N12210);
nand NAND2 (N16095, N16092, N972);
xor XOR2 (N16096, N16095, N10429);
nor NOR3 (N16097, N16083, N10435, N13390);
not NOT1 (N16098, N16065);
or OR2 (N16099, N16087, N12107);
nor NOR3 (N16100, N16084, N5540, N12864);
buf BUF1 (N16101, N16099);
xor XOR2 (N16102, N16098, N391);
xor XOR2 (N16103, N16102, N12616);
and AND2 (N16104, N16100, N3395);
or OR4 (N16105, N16104, N2320, N10999, N15489);
not NOT1 (N16106, N16101);
nor NOR2 (N16107, N16105, N1604);
nand NAND4 (N16108, N16094, N1860, N15291, N15735);
nor NOR2 (N16109, N16066, N7590);
nand NAND2 (N16110, N16061, N5569);
or OR4 (N16111, N16108, N9320, N7730, N4034);
buf BUF1 (N16112, N16111);
buf BUF1 (N16113, N16091);
buf BUF1 (N16114, N16093);
xor XOR2 (N16115, N16097, N3539);
not NOT1 (N16116, N16109);
or OR3 (N16117, N16113, N5609, N10535);
xor XOR2 (N16118, N16110, N16019);
buf BUF1 (N16119, N16114);
buf BUF1 (N16120, N16115);
buf BUF1 (N16121, N16117);
xor XOR2 (N16122, N16120, N13612);
buf BUF1 (N16123, N16121);
nor NOR2 (N16124, N16123, N7150);
not NOT1 (N16125, N16112);
buf BUF1 (N16126, N16119);
buf BUF1 (N16127, N16122);
xor XOR2 (N16128, N16125, N12076);
not NOT1 (N16129, N16103);
or OR3 (N16130, N16128, N4993, N15555);
xor XOR2 (N16131, N16116, N3569);
xor XOR2 (N16132, N16126, N15708);
xor XOR2 (N16133, N16131, N14459);
xor XOR2 (N16134, N16107, N10545);
xor XOR2 (N16135, N16118, N13334);
nand NAND3 (N16136, N16132, N9324, N13670);
not NOT1 (N16137, N16130);
buf BUF1 (N16138, N16106);
or OR3 (N16139, N16135, N7267, N12389);
nor NOR2 (N16140, N16137, N14906);
nor NOR3 (N16141, N16140, N9895, N15075);
xor XOR2 (N16142, N16134, N2142);
buf BUF1 (N16143, N16139);
nand NAND2 (N16144, N16136, N10705);
nand NAND4 (N16145, N16143, N10866, N3137, N2838);
buf BUF1 (N16146, N16129);
or OR3 (N16147, N16146, N14575, N7040);
or OR2 (N16148, N16138, N739);
buf BUF1 (N16149, N16096);
nor NOR3 (N16150, N16145, N13064, N8795);
or OR2 (N16151, N16149, N3095);
or OR3 (N16152, N16144, N7728, N10933);
or OR3 (N16153, N16124, N13044, N14101);
or OR3 (N16154, N16147, N11478, N12927);
not NOT1 (N16155, N16152);
and AND2 (N16156, N16142, N6040);
nor NOR2 (N16157, N16150, N5527);
or OR3 (N16158, N16156, N977, N1809);
buf BUF1 (N16159, N16155);
not NOT1 (N16160, N16159);
buf BUF1 (N16161, N16133);
nor NOR3 (N16162, N16153, N140, N6032);
nand NAND4 (N16163, N16148, N6129, N14366, N1406);
or OR3 (N16164, N16157, N14537, N1642);
nand NAND4 (N16165, N16127, N316, N14120, N15987);
buf BUF1 (N16166, N16162);
and AND3 (N16167, N16158, N599, N7591);
or OR2 (N16168, N16163, N3668);
xor XOR2 (N16169, N16166, N287);
xor XOR2 (N16170, N16167, N6637);
not NOT1 (N16171, N16169);
and AND2 (N16172, N16141, N3397);
xor XOR2 (N16173, N16164, N8166);
nor NOR3 (N16174, N16170, N14300, N1491);
nand NAND3 (N16175, N16173, N13347, N6900);
xor XOR2 (N16176, N16165, N2826);
xor XOR2 (N16177, N16161, N2651);
xor XOR2 (N16178, N16154, N2560);
xor XOR2 (N16179, N16151, N5253);
or OR2 (N16180, N16177, N4766);
and AND3 (N16181, N16176, N4614, N7630);
buf BUF1 (N16182, N16181);
nor NOR4 (N16183, N16178, N8349, N10341, N13566);
buf BUF1 (N16184, N16175);
xor XOR2 (N16185, N16168, N814);
not NOT1 (N16186, N16182);
and AND4 (N16187, N16179, N8349, N8792, N4402);
nand NAND4 (N16188, N16174, N4020, N15878, N11936);
nor NOR3 (N16189, N16187, N2136, N6081);
or OR3 (N16190, N16180, N6854, N3743);
buf BUF1 (N16191, N16188);
nand NAND4 (N16192, N16172, N2707, N10560, N11142);
or OR3 (N16193, N16192, N2109, N14980);
nor NOR2 (N16194, N16191, N11818);
buf BUF1 (N16195, N16183);
nor NOR2 (N16196, N16185, N3454);
nor NOR4 (N16197, N16190, N11286, N16002, N5767);
and AND3 (N16198, N16171, N8503, N14398);
or OR2 (N16199, N16198, N16172);
and AND4 (N16200, N16196, N3509, N3814, N5830);
or OR4 (N16201, N16199, N4257, N5279, N4320);
or OR4 (N16202, N16193, N5484, N8735, N5528);
not NOT1 (N16203, N16186);
buf BUF1 (N16204, N16197);
nand NAND3 (N16205, N16200, N1672, N6949);
nor NOR2 (N16206, N16195, N2816);
nand NAND4 (N16207, N16201, N7542, N7810, N3804);
not NOT1 (N16208, N16205);
xor XOR2 (N16209, N16207, N11934);
buf BUF1 (N16210, N16203);
and AND2 (N16211, N16194, N11578);
or OR2 (N16212, N16211, N14264);
buf BUF1 (N16213, N16206);
or OR4 (N16214, N16209, N13752, N802, N7737);
xor XOR2 (N16215, N16160, N2177);
xor XOR2 (N16216, N16202, N5903);
not NOT1 (N16217, N16213);
nor NOR2 (N16218, N16215, N15833);
xor XOR2 (N16219, N16212, N14065);
or OR3 (N16220, N16208, N3362, N12149);
nor NOR3 (N16221, N16214, N9603, N8033);
nand NAND2 (N16222, N16220, N11029);
nor NOR4 (N16223, N16217, N15990, N12932, N2372);
and AND4 (N16224, N16216, N8240, N11238, N2186);
not NOT1 (N16225, N16189);
nand NAND3 (N16226, N16219, N4498, N8643);
nor NOR3 (N16227, N16224, N15048, N4012);
and AND3 (N16228, N16225, N11896, N11675);
xor XOR2 (N16229, N16222, N13215);
and AND2 (N16230, N16226, N12694);
nand NAND2 (N16231, N16223, N13614);
buf BUF1 (N16232, N16204);
and AND3 (N16233, N16221, N7926, N2222);
or OR4 (N16234, N16232, N5190, N14093, N6357);
not NOT1 (N16235, N16227);
or OR4 (N16236, N16233, N7084, N12118, N14131);
buf BUF1 (N16237, N16230);
xor XOR2 (N16238, N16229, N582);
nor NOR4 (N16239, N16236, N7207, N7574, N2954);
or OR2 (N16240, N16218, N7265);
xor XOR2 (N16241, N16235, N8773);
nand NAND2 (N16242, N16237, N2613);
or OR3 (N16243, N16240, N1957, N3025);
not NOT1 (N16244, N16242);
or OR2 (N16245, N16210, N1751);
not NOT1 (N16246, N16234);
xor XOR2 (N16247, N16228, N10606);
and AND2 (N16248, N16247, N9259);
xor XOR2 (N16249, N16239, N13673);
buf BUF1 (N16250, N16231);
buf BUF1 (N16251, N16243);
buf BUF1 (N16252, N16245);
buf BUF1 (N16253, N16252);
and AND2 (N16254, N16241, N10111);
or OR3 (N16255, N16248, N14521, N4334);
nand NAND3 (N16256, N16253, N4104, N13350);
or OR4 (N16257, N16251, N6008, N6432, N9461);
buf BUF1 (N16258, N16244);
or OR3 (N16259, N16249, N5277, N6382);
or OR3 (N16260, N16256, N3, N2516);
xor XOR2 (N16261, N16254, N13142);
or OR4 (N16262, N16257, N13247, N4753, N1718);
nor NOR3 (N16263, N16261, N2212, N5666);
and AND3 (N16264, N16250, N12849, N1901);
nand NAND4 (N16265, N16260, N3128, N6900, N15404);
buf BUF1 (N16266, N16258);
nor NOR2 (N16267, N16255, N15037);
nand NAND4 (N16268, N16265, N4246, N2523, N353);
nand NAND3 (N16269, N16267, N13820, N6523);
not NOT1 (N16270, N16184);
buf BUF1 (N16271, N16262);
and AND4 (N16272, N16268, N8387, N7763, N4528);
buf BUF1 (N16273, N16270);
xor XOR2 (N16274, N16269, N14232);
and AND2 (N16275, N16264, N15554);
xor XOR2 (N16276, N16238, N14179);
or OR4 (N16277, N16259, N3840, N5489, N12889);
nor NOR4 (N16278, N16276, N15732, N5906, N13791);
not NOT1 (N16279, N16274);
and AND2 (N16280, N16278, N8362);
or OR2 (N16281, N16272, N1760);
buf BUF1 (N16282, N16273);
xor XOR2 (N16283, N16280, N5215);
nor NOR4 (N16284, N16263, N15733, N6299, N7750);
xor XOR2 (N16285, N16284, N11216);
and AND3 (N16286, N16246, N2264, N15990);
nor NOR4 (N16287, N16283, N9114, N9482, N4792);
buf BUF1 (N16288, N16285);
xor XOR2 (N16289, N16275, N11732);
buf BUF1 (N16290, N16281);
or OR3 (N16291, N16277, N3394, N1302);
and AND3 (N16292, N16291, N5938, N10187);
nand NAND3 (N16293, N16286, N4998, N5284);
nand NAND4 (N16294, N16271, N16175, N69, N4678);
not NOT1 (N16295, N16290);
or OR2 (N16296, N16289, N14989);
nor NOR2 (N16297, N16293, N15472);
buf BUF1 (N16298, N16292);
buf BUF1 (N16299, N16296);
or OR4 (N16300, N16282, N15532, N5872, N5563);
nand NAND4 (N16301, N16279, N7621, N7787, N6662);
xor XOR2 (N16302, N16301, N9546);
buf BUF1 (N16303, N16302);
buf BUF1 (N16304, N16266);
not NOT1 (N16305, N16295);
and AND3 (N16306, N16298, N3243, N7495);
buf BUF1 (N16307, N16287);
buf BUF1 (N16308, N16306);
nor NOR2 (N16309, N16305, N9048);
nand NAND4 (N16310, N16304, N8138, N14766, N1755);
buf BUF1 (N16311, N16310);
nor NOR4 (N16312, N16300, N129, N6887, N15217);
nor NOR2 (N16313, N16288, N10826);
nand NAND4 (N16314, N16307, N9210, N6595, N14104);
or OR3 (N16315, N16309, N11327, N13008);
xor XOR2 (N16316, N16311, N3655);
nand NAND2 (N16317, N16316, N11276);
xor XOR2 (N16318, N16317, N2889);
nor NOR4 (N16319, N16299, N15521, N16203, N6242);
xor XOR2 (N16320, N16318, N7002);
nand NAND4 (N16321, N16314, N6654, N9782, N1992);
buf BUF1 (N16322, N16312);
or OR4 (N16323, N16319, N3341, N9495, N6227);
xor XOR2 (N16324, N16294, N9651);
nand NAND4 (N16325, N16315, N8780, N16093, N10485);
not NOT1 (N16326, N16313);
nor NOR4 (N16327, N16321, N7554, N8723, N10439);
and AND4 (N16328, N16297, N8207, N7627, N12194);
and AND3 (N16329, N16326, N11385, N2779);
xor XOR2 (N16330, N16322, N12646);
buf BUF1 (N16331, N16327);
not NOT1 (N16332, N16323);
xor XOR2 (N16333, N16320, N11707);
xor XOR2 (N16334, N16331, N13488);
or OR2 (N16335, N16303, N47);
buf BUF1 (N16336, N16332);
nor NOR3 (N16337, N16325, N8441, N15267);
or OR2 (N16338, N16335, N11221);
not NOT1 (N16339, N16333);
not NOT1 (N16340, N16336);
nor NOR2 (N16341, N16329, N8377);
buf BUF1 (N16342, N16308);
and AND2 (N16343, N16337, N443);
nand NAND2 (N16344, N16341, N4228);
nor NOR2 (N16345, N16338, N15004);
xor XOR2 (N16346, N16340, N12834);
and AND3 (N16347, N16346, N6798, N2746);
nand NAND2 (N16348, N16345, N10994);
xor XOR2 (N16349, N16328, N3673);
nor NOR3 (N16350, N16343, N10541, N3632);
or OR2 (N16351, N16350, N8722);
and AND2 (N16352, N16344, N2721);
nand NAND2 (N16353, N16349, N11527);
and AND4 (N16354, N16339, N2014, N7256, N1555);
nand NAND4 (N16355, N16353, N11827, N10852, N15310);
nor NOR2 (N16356, N16347, N6520);
not NOT1 (N16357, N16348);
nor NOR3 (N16358, N16356, N7122, N3824);
not NOT1 (N16359, N16334);
or OR3 (N16360, N16357, N9044, N10333);
or OR3 (N16361, N16355, N13500, N15381);
buf BUF1 (N16362, N16351);
not NOT1 (N16363, N16362);
nand NAND2 (N16364, N16324, N1376);
xor XOR2 (N16365, N16361, N5662);
and AND3 (N16366, N16359, N6713, N8944);
or OR2 (N16367, N16358, N10249);
buf BUF1 (N16368, N16364);
not NOT1 (N16369, N16354);
and AND4 (N16370, N16342, N10723, N8480, N12524);
and AND4 (N16371, N16366, N3815, N8653, N2684);
and AND2 (N16372, N16371, N6643);
and AND4 (N16373, N16360, N1307, N10595, N9057);
xor XOR2 (N16374, N16369, N889);
not NOT1 (N16375, N16367);
and AND2 (N16376, N16368, N10);
buf BUF1 (N16377, N16370);
not NOT1 (N16378, N16376);
or OR4 (N16379, N16363, N15452, N14389, N6556);
buf BUF1 (N16380, N16352);
not NOT1 (N16381, N16380);
nor NOR3 (N16382, N16379, N15469, N1753);
buf BUF1 (N16383, N16374);
and AND3 (N16384, N16330, N8136, N3781);
or OR2 (N16385, N16365, N1365);
not NOT1 (N16386, N16373);
xor XOR2 (N16387, N16384, N9269);
or OR2 (N16388, N16385, N140);
or OR2 (N16389, N16382, N15942);
not NOT1 (N16390, N16381);
nand NAND2 (N16391, N16389, N9844);
buf BUF1 (N16392, N16391);
and AND4 (N16393, N16375, N940, N3152, N15745);
or OR4 (N16394, N16378, N8868, N8369, N6212);
nor NOR3 (N16395, N16393, N7463, N15507);
or OR2 (N16396, N16387, N13958);
not NOT1 (N16397, N16383);
xor XOR2 (N16398, N16396, N2072);
xor XOR2 (N16399, N16372, N8823);
buf BUF1 (N16400, N16394);
nand NAND3 (N16401, N16395, N4088, N10492);
or OR2 (N16402, N16400, N12521);
or OR2 (N16403, N16398, N8586);
nand NAND4 (N16404, N16388, N5698, N9645, N11505);
buf BUF1 (N16405, N16392);
nand NAND2 (N16406, N16390, N2781);
buf BUF1 (N16407, N16405);
nand NAND4 (N16408, N16404, N11757, N11571, N11720);
not NOT1 (N16409, N16408);
xor XOR2 (N16410, N16406, N8242);
buf BUF1 (N16411, N16410);
nor NOR3 (N16412, N16402, N3835, N14822);
xor XOR2 (N16413, N16412, N3101);
nor NOR2 (N16414, N16413, N2297);
nand NAND2 (N16415, N16409, N7787);
buf BUF1 (N16416, N16386);
and AND3 (N16417, N16403, N11681, N15671);
or OR3 (N16418, N16417, N96, N12341);
not NOT1 (N16419, N16377);
or OR2 (N16420, N16415, N15860);
nor NOR3 (N16421, N16399, N5055, N357);
buf BUF1 (N16422, N16421);
not NOT1 (N16423, N16407);
nand NAND2 (N16424, N16420, N7531);
xor XOR2 (N16425, N16422, N2838);
xor XOR2 (N16426, N16423, N9434);
or OR4 (N16427, N16411, N3380, N5165, N7728);
nand NAND3 (N16428, N16419, N8250, N9582);
xor XOR2 (N16429, N16424, N12621);
nor NOR2 (N16430, N16418, N10372);
not NOT1 (N16431, N16430);
xor XOR2 (N16432, N16425, N10952);
xor XOR2 (N16433, N16426, N5933);
or OR4 (N16434, N16397, N5053, N2279, N14616);
not NOT1 (N16435, N16401);
xor XOR2 (N16436, N16431, N1703);
buf BUF1 (N16437, N16436);
buf BUF1 (N16438, N16429);
or OR2 (N16439, N16435, N3443);
or OR2 (N16440, N16438, N7922);
and AND3 (N16441, N16432, N4403, N3620);
nor NOR2 (N16442, N16428, N1044);
or OR2 (N16443, N16440, N3098);
xor XOR2 (N16444, N16434, N1348);
or OR3 (N16445, N16443, N9362, N1202);
not NOT1 (N16446, N16437);
xor XOR2 (N16447, N16414, N983);
nor NOR4 (N16448, N16444, N3261, N13204, N12477);
buf BUF1 (N16449, N16446);
not NOT1 (N16450, N16449);
buf BUF1 (N16451, N16450);
nand NAND4 (N16452, N16433, N7942, N839, N2871);
or OR4 (N16453, N16439, N5565, N1213, N9340);
and AND3 (N16454, N16451, N3050, N15265);
nand NAND3 (N16455, N16445, N13670, N4855);
nor NOR4 (N16456, N16447, N2854, N16002, N13012);
not NOT1 (N16457, N16455);
buf BUF1 (N16458, N16448);
nand NAND4 (N16459, N16453, N12462, N7332, N9690);
buf BUF1 (N16460, N16459);
nand NAND2 (N16461, N16456, N7764);
not NOT1 (N16462, N16460);
buf BUF1 (N16463, N16442);
nor NOR4 (N16464, N16427, N8500, N10364, N1745);
not NOT1 (N16465, N16463);
nand NAND3 (N16466, N16458, N8822, N11498);
or OR3 (N16467, N16441, N5086, N13690);
or OR4 (N16468, N16454, N11649, N13249, N5049);
or OR2 (N16469, N16466, N11789);
buf BUF1 (N16470, N16462);
nand NAND4 (N16471, N16416, N5259, N9609, N12502);
buf BUF1 (N16472, N16461);
buf BUF1 (N16473, N16470);
buf BUF1 (N16474, N16471);
buf BUF1 (N16475, N16464);
and AND2 (N16476, N16468, N12894);
not NOT1 (N16477, N16475);
buf BUF1 (N16478, N16472);
nand NAND4 (N16479, N16465, N13421, N1705, N9723);
xor XOR2 (N16480, N16452, N12128);
not NOT1 (N16481, N16476);
nand NAND3 (N16482, N16481, N4305, N7749);
nor NOR3 (N16483, N16478, N3092, N15512);
or OR2 (N16484, N16469, N4542);
not NOT1 (N16485, N16479);
xor XOR2 (N16486, N16473, N11824);
not NOT1 (N16487, N16482);
or OR4 (N16488, N16485, N7119, N14029, N5647);
not NOT1 (N16489, N16486);
or OR2 (N16490, N16480, N12769);
and AND4 (N16491, N16457, N7666, N11894, N6052);
xor XOR2 (N16492, N16491, N11975);
nand NAND2 (N16493, N16490, N14305);
not NOT1 (N16494, N16484);
xor XOR2 (N16495, N16493, N5656);
not NOT1 (N16496, N16495);
nand NAND3 (N16497, N16487, N15087, N13656);
buf BUF1 (N16498, N16477);
nand NAND3 (N16499, N16489, N15273, N16403);
not NOT1 (N16500, N16498);
nand NAND2 (N16501, N16497, N3085);
and AND3 (N16502, N16483, N6678, N9638);
xor XOR2 (N16503, N16492, N12221);
nand NAND3 (N16504, N16500, N7921, N10343);
buf BUF1 (N16505, N16504);
not NOT1 (N16506, N16474);
buf BUF1 (N16507, N16501);
nand NAND2 (N16508, N16499, N1915);
nand NAND2 (N16509, N16505, N713);
or OR4 (N16510, N16502, N12801, N3737, N16373);
xor XOR2 (N16511, N16508, N7933);
not NOT1 (N16512, N16506);
not NOT1 (N16513, N16507);
and AND4 (N16514, N16509, N673, N408, N3319);
xor XOR2 (N16515, N16488, N15708);
buf BUF1 (N16516, N16496);
xor XOR2 (N16517, N16467, N9652);
not NOT1 (N16518, N16494);
xor XOR2 (N16519, N16514, N8031);
nor NOR3 (N16520, N16519, N5183, N638);
and AND3 (N16521, N16510, N15856, N15020);
not NOT1 (N16522, N16503);
nand NAND3 (N16523, N16515, N4495, N8399);
or OR2 (N16524, N16520, N3560);
and AND2 (N16525, N16524, N10517);
buf BUF1 (N16526, N16523);
and AND2 (N16527, N16521, N16368);
not NOT1 (N16528, N16527);
buf BUF1 (N16529, N16528);
xor XOR2 (N16530, N16526, N11982);
nand NAND3 (N16531, N16517, N14607, N13800);
nor NOR2 (N16532, N16516, N1200);
and AND2 (N16533, N16532, N10769);
nor NOR2 (N16534, N16530, N13440);
and AND2 (N16535, N16525, N15157);
nor NOR4 (N16536, N16518, N4293, N5851, N10272);
and AND3 (N16537, N16512, N3263, N15025);
not NOT1 (N16538, N16534);
buf BUF1 (N16539, N16531);
not NOT1 (N16540, N16536);
not NOT1 (N16541, N16540);
and AND4 (N16542, N16539, N14318, N1937, N5661);
buf BUF1 (N16543, N16537);
buf BUF1 (N16544, N16533);
buf BUF1 (N16545, N16511);
or OR3 (N16546, N16545, N16359, N3305);
nand NAND4 (N16547, N16543, N5634, N5118, N11042);
or OR4 (N16548, N16544, N5067, N13769, N14723);
not NOT1 (N16549, N16548);
or OR2 (N16550, N16535, N16350);
and AND2 (N16551, N16513, N13816);
nor NOR2 (N16552, N16547, N8837);
not NOT1 (N16553, N16522);
buf BUF1 (N16554, N16552);
buf BUF1 (N16555, N16549);
xor XOR2 (N16556, N16550, N1213);
or OR2 (N16557, N16554, N14527);
nor NOR3 (N16558, N16538, N11151, N14673);
nor NOR3 (N16559, N16553, N15472, N2068);
or OR3 (N16560, N16546, N9929, N7902);
or OR4 (N16561, N16556, N13908, N8926, N12201);
xor XOR2 (N16562, N16542, N6082);
not NOT1 (N16563, N16555);
buf BUF1 (N16564, N16557);
xor XOR2 (N16565, N16541, N13810);
nand NAND4 (N16566, N16560, N2117, N8669, N12590);
and AND2 (N16567, N16558, N12718);
not NOT1 (N16568, N16529);
nand NAND4 (N16569, N16567, N7671, N1903, N810);
buf BUF1 (N16570, N16563);
nand NAND3 (N16571, N16568, N14031, N1600);
xor XOR2 (N16572, N16559, N16418);
not NOT1 (N16573, N16562);
xor XOR2 (N16574, N16551, N14090);
buf BUF1 (N16575, N16566);
buf BUF1 (N16576, N16569);
or OR2 (N16577, N16573, N3876);
nand NAND2 (N16578, N16561, N10139);
buf BUF1 (N16579, N16578);
xor XOR2 (N16580, N16571, N3577);
nand NAND2 (N16581, N16579, N515);
or OR4 (N16582, N16580, N837, N3507, N5313);
xor XOR2 (N16583, N16564, N457);
or OR2 (N16584, N16582, N11014);
xor XOR2 (N16585, N16570, N1725);
xor XOR2 (N16586, N16565, N13507);
nor NOR3 (N16587, N16581, N6583, N3427);
nand NAND4 (N16588, N16574, N10227, N2542, N9573);
and AND3 (N16589, N16572, N8657, N2176);
not NOT1 (N16590, N16586);
or OR2 (N16591, N16588, N13757);
nor NOR3 (N16592, N16583, N2638, N10125);
buf BUF1 (N16593, N16575);
and AND2 (N16594, N16585, N8284);
buf BUF1 (N16595, N16594);
not NOT1 (N16596, N16595);
not NOT1 (N16597, N16577);
nand NAND4 (N16598, N16589, N8167, N2688, N4565);
and AND2 (N16599, N16592, N5217);
and AND2 (N16600, N16599, N13466);
buf BUF1 (N16601, N16600);
nor NOR4 (N16602, N16593, N5176, N4171, N7618);
nor NOR4 (N16603, N16601, N12213, N13016, N6716);
or OR4 (N16604, N16587, N5697, N12081, N6742);
and AND3 (N16605, N16590, N11863, N6044);
xor XOR2 (N16606, N16604, N11513);
or OR2 (N16607, N16602, N2420);
buf BUF1 (N16608, N16607);
nor NOR2 (N16609, N16584, N14177);
not NOT1 (N16610, N16576);
or OR4 (N16611, N16606, N6727, N5254, N4442);
not NOT1 (N16612, N16591);
xor XOR2 (N16613, N16611, N3731);
xor XOR2 (N16614, N16608, N15027);
xor XOR2 (N16615, N16613, N11352);
and AND2 (N16616, N16612, N10160);
nand NAND3 (N16617, N16597, N5134, N7252);
nor NOR2 (N16618, N16616, N5990);
xor XOR2 (N16619, N16609, N14655);
not NOT1 (N16620, N16605);
nand NAND3 (N16621, N16618, N10508, N4422);
and AND2 (N16622, N16621, N12009);
xor XOR2 (N16623, N16615, N10935);
not NOT1 (N16624, N16603);
nor NOR3 (N16625, N16598, N14684, N7707);
nor NOR4 (N16626, N16623, N16246, N9370, N11529);
and AND2 (N16627, N16614, N11590);
nand NAND4 (N16628, N16617, N7770, N4804, N15908);
not NOT1 (N16629, N16619);
or OR2 (N16630, N16610, N13348);
nor NOR4 (N16631, N16626, N11320, N2744, N10519);
nor NOR4 (N16632, N16631, N10284, N15942, N5963);
nand NAND2 (N16633, N16622, N12058);
nor NOR4 (N16634, N16632, N10060, N2094, N15733);
buf BUF1 (N16635, N16625);
or OR4 (N16636, N16627, N6215, N10405, N5131);
not NOT1 (N16637, N16624);
or OR2 (N16638, N16620, N9900);
and AND4 (N16639, N16633, N4191, N464, N12060);
nand NAND3 (N16640, N16596, N594, N1794);
or OR2 (N16641, N16638, N7542);
xor XOR2 (N16642, N16628, N9471);
not NOT1 (N16643, N16642);
nor NOR4 (N16644, N16630, N5396, N2597, N13892);
not NOT1 (N16645, N16629);
buf BUF1 (N16646, N16640);
and AND2 (N16647, N16634, N7808);
nand NAND4 (N16648, N16647, N4588, N493, N3764);
nor NOR4 (N16649, N16641, N6307, N4400, N11606);
not NOT1 (N16650, N16637);
not NOT1 (N16651, N16644);
xor XOR2 (N16652, N16650, N4369);
xor XOR2 (N16653, N16646, N3736);
nor NOR2 (N16654, N16653, N392);
buf BUF1 (N16655, N16654);
or OR3 (N16656, N16645, N1377, N1833);
not NOT1 (N16657, N16649);
or OR3 (N16658, N16652, N2500, N12261);
or OR3 (N16659, N16648, N10623, N14395);
nor NOR2 (N16660, N16636, N12272);
nand NAND2 (N16661, N16635, N7701);
xor XOR2 (N16662, N16656, N13087);
or OR4 (N16663, N16651, N4989, N979, N13435);
xor XOR2 (N16664, N16643, N2153);
xor XOR2 (N16665, N16661, N5975);
buf BUF1 (N16666, N16660);
xor XOR2 (N16667, N16664, N10618);
and AND2 (N16668, N16665, N6891);
nand NAND3 (N16669, N16668, N14135, N13806);
xor XOR2 (N16670, N16662, N9523);
or OR4 (N16671, N16670, N6423, N16642, N12869);
or OR4 (N16672, N16655, N5175, N14082, N1350);
not NOT1 (N16673, N16659);
nand NAND3 (N16674, N16671, N11999, N580);
nor NOR4 (N16675, N16666, N1329, N12871, N4542);
and AND2 (N16676, N16639, N6203);
and AND4 (N16677, N16669, N8850, N14086, N1733);
and AND4 (N16678, N16673, N3363, N12283, N6645);
xor XOR2 (N16679, N16667, N7216);
or OR2 (N16680, N16663, N15058);
not NOT1 (N16681, N16674);
or OR4 (N16682, N16675, N8117, N853, N6573);
nor NOR2 (N16683, N16678, N5229);
or OR4 (N16684, N16680, N10778, N11039, N6087);
nor NOR4 (N16685, N16684, N7889, N11511, N2346);
nor NOR4 (N16686, N16681, N8123, N16236, N13151);
nand NAND4 (N16687, N16672, N16265, N3467, N3212);
and AND4 (N16688, N16677, N15949, N6856, N8504);
or OR4 (N16689, N16685, N6602, N279, N1176);
nand NAND3 (N16690, N16676, N2247, N6920);
xor XOR2 (N16691, N16686, N2054);
and AND4 (N16692, N16679, N9724, N11898, N8214);
nor NOR3 (N16693, N16683, N568, N3974);
buf BUF1 (N16694, N16658);
buf BUF1 (N16695, N16693);
nand NAND3 (N16696, N16694, N7996, N15822);
buf BUF1 (N16697, N16695);
not NOT1 (N16698, N16682);
and AND4 (N16699, N16691, N14396, N1133, N3005);
or OR3 (N16700, N16687, N7613, N10198);
xor XOR2 (N16701, N16697, N6245);
nand NAND2 (N16702, N16692, N9624);
and AND3 (N16703, N16657, N12152, N3097);
nand NAND4 (N16704, N16701, N6141, N11629, N468);
buf BUF1 (N16705, N16696);
and AND2 (N16706, N16704, N13580);
or OR4 (N16707, N16689, N2213, N11085, N6567);
not NOT1 (N16708, N16690);
or OR4 (N16709, N16688, N12151, N9795, N10268);
not NOT1 (N16710, N16707);
not NOT1 (N16711, N16699);
not NOT1 (N16712, N16698);
buf BUF1 (N16713, N16703);
xor XOR2 (N16714, N16702, N2597);
nor NOR3 (N16715, N16706, N8121, N8132);
not NOT1 (N16716, N16710);
or OR2 (N16717, N16712, N15038);
or OR2 (N16718, N16713, N7305);
or OR3 (N16719, N16705, N5614, N3092);
nor NOR3 (N16720, N16719, N2251, N13486);
nor NOR4 (N16721, N16700, N6874, N2097, N12889);
and AND2 (N16722, N16721, N15118);
or OR3 (N16723, N16711, N16218, N11921);
nand NAND2 (N16724, N16709, N3214);
nor NOR2 (N16725, N16723, N2877);
buf BUF1 (N16726, N16720);
or OR3 (N16727, N16725, N15070, N14645);
xor XOR2 (N16728, N16722, N8433);
nor NOR3 (N16729, N16728, N799, N872);
nand NAND3 (N16730, N16716, N7205, N11441);
or OR4 (N16731, N16715, N13720, N1049, N8280);
buf BUF1 (N16732, N16717);
xor XOR2 (N16733, N16729, N8636);
not NOT1 (N16734, N16708);
or OR4 (N16735, N16734, N14450, N2946, N7935);
not NOT1 (N16736, N16727);
buf BUF1 (N16737, N16726);
or OR4 (N16738, N16718, N16329, N5560, N11307);
nor NOR3 (N16739, N16724, N13215, N403);
nor NOR2 (N16740, N16733, N8795);
nand NAND3 (N16741, N16737, N11417, N5729);
not NOT1 (N16742, N16738);
nand NAND2 (N16743, N16732, N1759);
or OR2 (N16744, N16735, N4457);
buf BUF1 (N16745, N16743);
buf BUF1 (N16746, N16730);
not NOT1 (N16747, N16714);
and AND3 (N16748, N16747, N9605, N873);
and AND3 (N16749, N16740, N6429, N2689);
nand NAND3 (N16750, N16748, N15635, N5872);
or OR2 (N16751, N16746, N9134);
not NOT1 (N16752, N16736);
not NOT1 (N16753, N16752);
or OR2 (N16754, N16741, N1988);
nor NOR2 (N16755, N16753, N9102);
not NOT1 (N16756, N16744);
and AND4 (N16757, N16756, N596, N5597, N2793);
not NOT1 (N16758, N16749);
or OR4 (N16759, N16731, N11162, N7670, N4609);
and AND3 (N16760, N16759, N2229, N9551);
and AND3 (N16761, N16760, N4724, N1276);
buf BUF1 (N16762, N16739);
buf BUF1 (N16763, N16761);
nand NAND4 (N16764, N16755, N6952, N5783, N8583);
buf BUF1 (N16765, N16742);
xor XOR2 (N16766, N16765, N5902);
nor NOR4 (N16767, N16766, N5634, N4193, N15239);
nand NAND4 (N16768, N16745, N10370, N9356, N1606);
or OR3 (N16769, N16751, N8755, N13961);
xor XOR2 (N16770, N16768, N7394);
and AND4 (N16771, N16767, N2474, N6805, N4283);
not NOT1 (N16772, N16769);
nor NOR3 (N16773, N16762, N12872, N6474);
nand NAND2 (N16774, N16750, N2496);
or OR2 (N16775, N16758, N7369);
or OR3 (N16776, N16757, N5023, N3238);
buf BUF1 (N16777, N16770);
or OR4 (N16778, N16771, N1769, N3247, N6361);
nor NOR4 (N16779, N16776, N3261, N12001, N13086);
buf BUF1 (N16780, N16754);
nand NAND4 (N16781, N16779, N15508, N16057, N4028);
not NOT1 (N16782, N16773);
and AND2 (N16783, N16782, N6896);
buf BUF1 (N16784, N16781);
xor XOR2 (N16785, N16778, N9992);
nor NOR2 (N16786, N16775, N15933);
nor NOR2 (N16787, N16784, N13493);
buf BUF1 (N16788, N16786);
nand NAND4 (N16789, N16788, N5318, N5402, N14533);
not NOT1 (N16790, N16774);
xor XOR2 (N16791, N16764, N15901);
nor NOR2 (N16792, N16785, N1142);
buf BUF1 (N16793, N16789);
nand NAND2 (N16794, N16763, N13098);
xor XOR2 (N16795, N16783, N10837);
or OR2 (N16796, N16792, N5827);
buf BUF1 (N16797, N16777);
buf BUF1 (N16798, N16796);
xor XOR2 (N16799, N16798, N10391);
or OR2 (N16800, N16799, N15238);
xor XOR2 (N16801, N16787, N6954);
buf BUF1 (N16802, N16780);
nand NAND4 (N16803, N16801, N12587, N2118, N15933);
and AND3 (N16804, N16791, N1751, N14688);
or OR3 (N16805, N16797, N6754, N15340);
or OR4 (N16806, N16803, N253, N8187, N10456);
and AND2 (N16807, N16805, N11742);
xor XOR2 (N16808, N16807, N14939);
nor NOR4 (N16809, N16802, N9242, N1983, N15048);
buf BUF1 (N16810, N16795);
xor XOR2 (N16811, N16800, N13172);
not NOT1 (N16812, N16809);
buf BUF1 (N16813, N16808);
nor NOR4 (N16814, N16804, N15828, N11730, N8267);
or OR2 (N16815, N16814, N2629);
nand NAND3 (N16816, N16813, N11143, N6188);
buf BUF1 (N16817, N16816);
nor NOR4 (N16818, N16790, N12910, N12935, N2393);
xor XOR2 (N16819, N16811, N14231);
nand NAND3 (N16820, N16793, N14632, N4777);
nand NAND4 (N16821, N16818, N6589, N8088, N2844);
xor XOR2 (N16822, N16794, N15035);
not NOT1 (N16823, N16815);
and AND3 (N16824, N16823, N9305, N2223);
nand NAND4 (N16825, N16821, N15216, N15975, N9579);
buf BUF1 (N16826, N16810);
or OR3 (N16827, N16806, N968, N2519);
or OR2 (N16828, N16822, N4330);
nor NOR2 (N16829, N16828, N15462);
buf BUF1 (N16830, N16824);
and AND2 (N16831, N16830, N5055);
buf BUF1 (N16832, N16819);
nand NAND4 (N16833, N16772, N1830, N1010, N11581);
xor XOR2 (N16834, N16832, N12529);
nor NOR3 (N16835, N16829, N6721, N8888);
nand NAND3 (N16836, N16820, N8349, N9776);
buf BUF1 (N16837, N16833);
nand NAND2 (N16838, N16835, N15514);
or OR3 (N16839, N16831, N5009, N7237);
xor XOR2 (N16840, N16812, N8285);
xor XOR2 (N16841, N16827, N15206);
and AND3 (N16842, N16825, N14101, N14315);
and AND4 (N16843, N16826, N6151, N10193, N14294);
or OR3 (N16844, N16834, N12964, N15247);
or OR3 (N16845, N16844, N7616, N8893);
nor NOR2 (N16846, N16836, N12455);
xor XOR2 (N16847, N16817, N7220);
xor XOR2 (N16848, N16843, N6436);
or OR4 (N16849, N16846, N13744, N10143, N13277);
xor XOR2 (N16850, N16847, N5706);
buf BUF1 (N16851, N16849);
nand NAND3 (N16852, N16845, N3298, N16378);
nand NAND2 (N16853, N16840, N13137);
and AND4 (N16854, N16850, N3830, N6758, N7270);
nor NOR2 (N16855, N16848, N4211);
not NOT1 (N16856, N16855);
or OR4 (N16857, N16853, N15796, N5174, N16798);
or OR3 (N16858, N16854, N2036, N624);
nand NAND4 (N16859, N16852, N16806, N4495, N7832);
nor NOR4 (N16860, N16851, N16242, N11826, N962);
not NOT1 (N16861, N16858);
nand NAND3 (N16862, N16857, N11212, N13524);
xor XOR2 (N16863, N16837, N2190);
not NOT1 (N16864, N16841);
nand NAND3 (N16865, N16861, N14277, N6875);
buf BUF1 (N16866, N16838);
nor NOR3 (N16867, N16862, N16425, N1278);
buf BUF1 (N16868, N16864);
nand NAND2 (N16869, N16839, N2284);
not NOT1 (N16870, N16865);
nand NAND4 (N16871, N16863, N11731, N6646, N9212);
not NOT1 (N16872, N16868);
buf BUF1 (N16873, N16871);
or OR3 (N16874, N16860, N3234, N7443);
xor XOR2 (N16875, N16842, N15961);
nand NAND3 (N16876, N16872, N3053, N2240);
and AND3 (N16877, N16870, N13422, N349);
buf BUF1 (N16878, N16877);
not NOT1 (N16879, N16873);
buf BUF1 (N16880, N16875);
not NOT1 (N16881, N16876);
buf BUF1 (N16882, N16869);
nand NAND2 (N16883, N16856, N2934);
or OR4 (N16884, N16859, N7544, N16263, N16383);
or OR2 (N16885, N16882, N538);
not NOT1 (N16886, N16878);
not NOT1 (N16887, N16879);
nand NAND4 (N16888, N16887, N8457, N4219, N11206);
and AND2 (N16889, N16880, N584);
nand NAND4 (N16890, N16874, N4198, N13588, N3827);
xor XOR2 (N16891, N16881, N5909);
not NOT1 (N16892, N16888);
buf BUF1 (N16893, N16884);
nor NOR2 (N16894, N16891, N12422);
not NOT1 (N16895, N16886);
or OR3 (N16896, N16892, N3172, N9079);
and AND2 (N16897, N16867, N16159);
nand NAND2 (N16898, N16890, N9129);
or OR2 (N16899, N16898, N8980);
or OR2 (N16900, N16894, N14124);
nor NOR2 (N16901, N16896, N13739);
or OR2 (N16902, N16866, N2946);
nor NOR4 (N16903, N16893, N5868, N8424, N9714);
buf BUF1 (N16904, N16883);
not NOT1 (N16905, N16904);
not NOT1 (N16906, N16899);
xor XOR2 (N16907, N16905, N4895);
xor XOR2 (N16908, N16885, N6688);
and AND4 (N16909, N16889, N1787, N10691, N4860);
or OR4 (N16910, N16906, N10647, N4023, N13610);
or OR4 (N16911, N16903, N10287, N5573, N7705);
buf BUF1 (N16912, N16902);
nand NAND3 (N16913, N16908, N7193, N12395);
and AND3 (N16914, N16900, N800, N7234);
not NOT1 (N16915, N16895);
xor XOR2 (N16916, N16907, N11839);
nand NAND4 (N16917, N16901, N6294, N13169, N2781);
buf BUF1 (N16918, N16916);
buf BUF1 (N16919, N16912);
not NOT1 (N16920, N16913);
buf BUF1 (N16921, N16915);
nor NOR4 (N16922, N16911, N7527, N15998, N6755);
xor XOR2 (N16923, N16914, N10433);
and AND2 (N16924, N16920, N14315);
xor XOR2 (N16925, N16922, N587);
and AND2 (N16926, N16925, N11449);
nand NAND2 (N16927, N16921, N2736);
or OR4 (N16928, N16919, N8737, N15184, N1424);
xor XOR2 (N16929, N16897, N1793);
buf BUF1 (N16930, N16927);
buf BUF1 (N16931, N16930);
buf BUF1 (N16932, N16910);
or OR2 (N16933, N16931, N662);
nand NAND4 (N16934, N16932, N6451, N15060, N11422);
nor NOR2 (N16935, N16917, N2788);
xor XOR2 (N16936, N16935, N14996);
xor XOR2 (N16937, N16936, N12556);
buf BUF1 (N16938, N16928);
nand NAND4 (N16939, N16909, N11991, N15659, N2224);
or OR4 (N16940, N16933, N1011, N2708, N10716);
nor NOR2 (N16941, N16940, N9355);
buf BUF1 (N16942, N16918);
nor NOR4 (N16943, N16938, N12154, N15549, N4517);
buf BUF1 (N16944, N16923);
nor NOR4 (N16945, N16924, N14349, N1459, N5179);
or OR3 (N16946, N16926, N9896, N15425);
not NOT1 (N16947, N16929);
or OR2 (N16948, N16942, N4958);
nor NOR2 (N16949, N16945, N5193);
xor XOR2 (N16950, N16941, N1965);
nand NAND4 (N16951, N16937, N16081, N16734, N15815);
not NOT1 (N16952, N16946);
nor NOR3 (N16953, N16950, N7570, N14721);
xor XOR2 (N16954, N16952, N4454);
buf BUF1 (N16955, N16947);
and AND2 (N16956, N16934, N12613);
or OR3 (N16957, N16949, N8309, N14984);
buf BUF1 (N16958, N16951);
nor NOR3 (N16959, N16953, N2903, N4357);
and AND4 (N16960, N16954, N3551, N2972, N14023);
not NOT1 (N16961, N16957);
buf BUF1 (N16962, N16948);
nor NOR3 (N16963, N16961, N2715, N4031);
and AND3 (N16964, N16956, N2231, N2100);
nor NOR3 (N16965, N16962, N16962, N5414);
nand NAND2 (N16966, N16965, N1750);
nor NOR2 (N16967, N16955, N2599);
and AND3 (N16968, N16966, N2974, N13947);
xor XOR2 (N16969, N16959, N10593);
nand NAND2 (N16970, N16958, N15079);
or OR3 (N16971, N16967, N10411, N7503);
nor NOR4 (N16972, N16971, N14866, N5749, N16722);
nor NOR3 (N16973, N16963, N6479, N3753);
xor XOR2 (N16974, N16969, N6577);
not NOT1 (N16975, N16970);
or OR4 (N16976, N16974, N10096, N10683, N13125);
nor NOR4 (N16977, N16968, N10228, N15444, N12426);
nor NOR2 (N16978, N16977, N6108);
and AND2 (N16979, N16978, N7630);
or OR3 (N16980, N16939, N14346, N11335);
or OR4 (N16981, N16960, N7814, N11147, N3239);
nor NOR3 (N16982, N16980, N5250, N2795);
xor XOR2 (N16983, N16944, N15083);
nand NAND3 (N16984, N16982, N9345, N13035);
not NOT1 (N16985, N16973);
nor NOR2 (N16986, N16964, N5431);
or OR3 (N16987, N16985, N9707, N8294);
buf BUF1 (N16988, N16984);
buf BUF1 (N16989, N16983);
nand NAND2 (N16990, N16979, N7866);
or OR4 (N16991, N16989, N9388, N10360, N13741);
nor NOR4 (N16992, N16988, N14288, N10888, N2707);
and AND3 (N16993, N16987, N16752, N379);
nor NOR3 (N16994, N16943, N11040, N1621);
nand NAND4 (N16995, N16976, N4742, N8646, N6928);
nand NAND4 (N16996, N16991, N10245, N11331, N6356);
and AND3 (N16997, N16996, N15794, N14203);
not NOT1 (N16998, N16990);
nand NAND3 (N16999, N16998, N3790, N619);
buf BUF1 (N17000, N16986);
nand NAND3 (N17001, N17000, N11511, N16064);
or OR2 (N17002, N16972, N2467);
and AND4 (N17003, N17001, N15571, N502, N13656);
buf BUF1 (N17004, N16981);
and AND4 (N17005, N16975, N10090, N7612, N8366);
or OR3 (N17006, N17004, N12572, N10851);
buf BUF1 (N17007, N16994);
and AND2 (N17008, N16992, N7825);
not NOT1 (N17009, N17002);
xor XOR2 (N17010, N16995, N13665);
nor NOR2 (N17011, N16993, N12692);
nand NAND2 (N17012, N17005, N13015);
nand NAND2 (N17013, N17011, N9681);
or OR3 (N17014, N16997, N12039, N7687);
xor XOR2 (N17015, N17012, N7597);
and AND4 (N17016, N17003, N16234, N15591, N12237);
nand NAND3 (N17017, N17008, N9335, N4970);
nand NAND4 (N17018, N17010, N3713, N856, N8774);
xor XOR2 (N17019, N17016, N6494);
nor NOR4 (N17020, N17014, N1928, N14876, N15084);
xor XOR2 (N17021, N17018, N3485);
buf BUF1 (N17022, N17021);
nand NAND4 (N17023, N17013, N12345, N11881, N4196);
or OR2 (N17024, N17020, N13931);
buf BUF1 (N17025, N17023);
and AND2 (N17026, N17022, N9520);
or OR4 (N17027, N17017, N7121, N5688, N2428);
nand NAND3 (N17028, N17006, N7880, N5054);
nor NOR2 (N17029, N16999, N7434);
nand NAND2 (N17030, N17026, N10788);
nor NOR3 (N17031, N17015, N15512, N14344);
nor NOR4 (N17032, N17024, N16163, N15242, N14532);
nor NOR2 (N17033, N17019, N2276);
not NOT1 (N17034, N17032);
and AND2 (N17035, N17007, N13562);
buf BUF1 (N17036, N17033);
not NOT1 (N17037, N17027);
nor NOR4 (N17038, N17031, N5799, N6958, N985);
xor XOR2 (N17039, N17035, N13157);
or OR4 (N17040, N17037, N10835, N7314, N6846);
nand NAND3 (N17041, N17030, N13719, N5525);
nor NOR2 (N17042, N17009, N2462);
nor NOR4 (N17043, N17029, N4509, N7352, N15912);
nor NOR3 (N17044, N17042, N9213, N6487);
buf BUF1 (N17045, N17038);
or OR3 (N17046, N17044, N8413, N12065);
nor NOR3 (N17047, N17043, N8665, N11875);
xor XOR2 (N17048, N17034, N12153);
not NOT1 (N17049, N17047);
buf BUF1 (N17050, N17039);
xor XOR2 (N17051, N17036, N3346);
nor NOR2 (N17052, N17028, N15073);
not NOT1 (N17053, N17045);
nand NAND2 (N17054, N17040, N17003);
and AND2 (N17055, N17051, N6854);
or OR2 (N17056, N17041, N4147);
buf BUF1 (N17057, N17048);
not NOT1 (N17058, N17055);
nand NAND4 (N17059, N17056, N11352, N4428, N11890);
and AND3 (N17060, N17057, N6175, N14355);
or OR4 (N17061, N17050, N9048, N15168, N8383);
not NOT1 (N17062, N17060);
xor XOR2 (N17063, N17052, N13545);
not NOT1 (N17064, N17061);
buf BUF1 (N17065, N17062);
not NOT1 (N17066, N17058);
and AND3 (N17067, N17066, N15671, N16243);
buf BUF1 (N17068, N17064);
and AND3 (N17069, N17049, N7126, N8385);
nand NAND4 (N17070, N17053, N1193, N413, N11509);
buf BUF1 (N17071, N17068);
and AND4 (N17072, N17071, N16433, N12134, N15835);
and AND3 (N17073, N17046, N15594, N15602);
and AND3 (N17074, N17067, N4513, N15529);
not NOT1 (N17075, N17065);
nand NAND2 (N17076, N17074, N12443);
buf BUF1 (N17077, N17072);
nor NOR4 (N17078, N17059, N13410, N6878, N10862);
xor XOR2 (N17079, N17054, N11999);
xor XOR2 (N17080, N17075, N8943);
buf BUF1 (N17081, N17078);
or OR4 (N17082, N17081, N1943, N16187, N14244);
not NOT1 (N17083, N17069);
xor XOR2 (N17084, N17073, N6694);
nor NOR4 (N17085, N17082, N14407, N3534, N16917);
or OR3 (N17086, N17085, N15719, N9347);
nor NOR3 (N17087, N17086, N6295, N14403);
and AND4 (N17088, N17084, N2664, N8406, N15684);
not NOT1 (N17089, N17063);
and AND4 (N17090, N17087, N2625, N15351, N9863);
xor XOR2 (N17091, N17077, N16126);
not NOT1 (N17092, N17025);
not NOT1 (N17093, N17070);
and AND3 (N17094, N17080, N2862, N5455);
xor XOR2 (N17095, N17089, N10013);
not NOT1 (N17096, N17091);
or OR4 (N17097, N17092, N16108, N14307, N13800);
and AND3 (N17098, N17095, N1227, N525);
or OR4 (N17099, N17090, N1033, N13381, N5210);
nand NAND3 (N17100, N17088, N3958, N9703);
not NOT1 (N17101, N17097);
nand NAND4 (N17102, N17093, N10584, N5050, N1530);
buf BUF1 (N17103, N17100);
buf BUF1 (N17104, N17096);
or OR4 (N17105, N17104, N3928, N14455, N3123);
not NOT1 (N17106, N17103);
or OR2 (N17107, N17106, N130);
nor NOR2 (N17108, N17079, N880);
not NOT1 (N17109, N17083);
or OR2 (N17110, N17101, N11083);
and AND3 (N17111, N17105, N16337, N4767);
nand NAND2 (N17112, N17109, N1030);
or OR4 (N17113, N17107, N2091, N16926, N2734);
not NOT1 (N17114, N17076);
nor NOR3 (N17115, N17114, N16286, N9674);
or OR3 (N17116, N17102, N15187, N11329);
or OR4 (N17117, N17110, N4440, N12066, N13353);
not NOT1 (N17118, N17098);
nand NAND2 (N17119, N17115, N15986);
nor NOR2 (N17120, N17099, N2448);
nand NAND2 (N17121, N17119, N4830);
or OR3 (N17122, N17121, N5598, N12128);
nand NAND4 (N17123, N17112, N4224, N5123, N383);
not NOT1 (N17124, N17123);
xor XOR2 (N17125, N17120, N14989);
and AND2 (N17126, N17111, N8896);
buf BUF1 (N17127, N17116);
or OR3 (N17128, N17124, N13133, N11210);
buf BUF1 (N17129, N17117);
or OR3 (N17130, N17118, N3550, N16463);
xor XOR2 (N17131, N17129, N10654);
nand NAND2 (N17132, N17131, N11158);
or OR4 (N17133, N17113, N8446, N8918, N1475);
or OR2 (N17134, N17132, N7995);
nand NAND4 (N17135, N17130, N13293, N15900, N33);
or OR2 (N17136, N17133, N10375);
not NOT1 (N17137, N17136);
nand NAND3 (N17138, N17125, N6449, N6958);
or OR4 (N17139, N17126, N9720, N13715, N9241);
nand NAND4 (N17140, N17094, N10632, N3353, N1591);
or OR2 (N17141, N17135, N7535);
xor XOR2 (N17142, N17140, N12428);
and AND2 (N17143, N17139, N9328);
not NOT1 (N17144, N17137);
or OR2 (N17145, N17144, N17032);
and AND4 (N17146, N17143, N11135, N16133, N14573);
or OR4 (N17147, N17142, N2593, N2997, N13162);
and AND4 (N17148, N17108, N11707, N5596, N4107);
not NOT1 (N17149, N17145);
or OR3 (N17150, N17149, N3972, N12595);
xor XOR2 (N17151, N17122, N14556);
buf BUF1 (N17152, N17148);
nand NAND2 (N17153, N17138, N8637);
nand NAND2 (N17154, N17134, N14238);
nand NAND4 (N17155, N17153, N15845, N701, N4218);
xor XOR2 (N17156, N17147, N937);
nand NAND4 (N17157, N17156, N12436, N3810, N14289);
buf BUF1 (N17158, N17128);
buf BUF1 (N17159, N17157);
buf BUF1 (N17160, N17159);
or OR3 (N17161, N17155, N10213, N6447);
and AND2 (N17162, N17150, N5811);
or OR2 (N17163, N17152, N4909);
and AND4 (N17164, N17151, N3393, N7319, N449);
nand NAND3 (N17165, N17161, N13537, N8490);
and AND3 (N17166, N17164, N5039, N803);
buf BUF1 (N17167, N17165);
buf BUF1 (N17168, N17162);
or OR4 (N17169, N17154, N1236, N8315, N9710);
buf BUF1 (N17170, N17163);
nor NOR3 (N17171, N17167, N11748, N7902);
xor XOR2 (N17172, N17168, N6120);
not NOT1 (N17173, N17160);
nand NAND2 (N17174, N17173, N15626);
and AND2 (N17175, N17158, N16850);
and AND2 (N17176, N17146, N12229);
nor NOR4 (N17177, N17176, N14754, N12306, N9199);
xor XOR2 (N17178, N17166, N5076);
not NOT1 (N17179, N17175);
and AND2 (N17180, N17174, N8724);
not NOT1 (N17181, N17141);
xor XOR2 (N17182, N17172, N15887);
not NOT1 (N17183, N17169);
buf BUF1 (N17184, N17171);
or OR2 (N17185, N17179, N16433);
nand NAND2 (N17186, N17127, N4276);
nor NOR3 (N17187, N17186, N3914, N4205);
and AND4 (N17188, N17183, N6271, N7041, N1001);
nand NAND4 (N17189, N17188, N11492, N10960, N1689);
xor XOR2 (N17190, N17170, N16651);
nand NAND4 (N17191, N17178, N3619, N6872, N6330);
nand NAND3 (N17192, N17182, N13760, N10456);
not NOT1 (N17193, N17192);
nand NAND3 (N17194, N17190, N8899, N5786);
or OR4 (N17195, N17180, N5050, N1994, N8929);
buf BUF1 (N17196, N17193);
and AND2 (N17197, N17191, N4611);
and AND4 (N17198, N17181, N15812, N6782, N16057);
and AND3 (N17199, N17195, N14435, N112);
nand NAND3 (N17200, N17198, N16054, N14227);
nor NOR4 (N17201, N17200, N1187, N548, N9611);
xor XOR2 (N17202, N17201, N15248);
buf BUF1 (N17203, N17194);
nor NOR2 (N17204, N17189, N4464);
nor NOR2 (N17205, N17177, N14187);
buf BUF1 (N17206, N17185);
buf BUF1 (N17207, N17196);
not NOT1 (N17208, N17202);
and AND2 (N17209, N17199, N11385);
nand NAND4 (N17210, N17184, N12369, N17016, N1027);
nor NOR4 (N17211, N17203, N3128, N9463, N11372);
not NOT1 (N17212, N17208);
or OR4 (N17213, N17209, N8663, N2919, N13072);
nand NAND4 (N17214, N17197, N8110, N8686, N4725);
or OR2 (N17215, N17211, N17009);
not NOT1 (N17216, N17206);
or OR3 (N17217, N17210, N6430, N8274);
nand NAND4 (N17218, N17212, N743, N3250, N13932);
buf BUF1 (N17219, N17218);
xor XOR2 (N17220, N17217, N3550);
and AND4 (N17221, N17216, N3787, N4781, N5943);
xor XOR2 (N17222, N17221, N9891);
nand NAND3 (N17223, N17222, N1688, N8102);
nor NOR2 (N17224, N17187, N14369);
not NOT1 (N17225, N17223);
nand NAND2 (N17226, N17214, N8716);
not NOT1 (N17227, N17204);
buf BUF1 (N17228, N17227);
nor NOR3 (N17229, N17228, N28, N10315);
nor NOR4 (N17230, N17219, N14139, N4283, N6010);
xor XOR2 (N17231, N17205, N16222);
nor NOR2 (N17232, N17207, N4814);
not NOT1 (N17233, N17224);
xor XOR2 (N17234, N17233, N15019);
buf BUF1 (N17235, N17220);
and AND3 (N17236, N17229, N10992, N7321);
xor XOR2 (N17237, N17234, N1450);
xor XOR2 (N17238, N17225, N12731);
buf BUF1 (N17239, N17231);
nor NOR4 (N17240, N17239, N6247, N15981, N10351);
nand NAND3 (N17241, N17235, N2490, N3753);
xor XOR2 (N17242, N17241, N147);
nand NAND3 (N17243, N17237, N10774, N11337);
nand NAND3 (N17244, N17213, N2225, N9369);
or OR3 (N17245, N17242, N3414, N13081);
nor NOR4 (N17246, N17232, N359, N4418, N247);
xor XOR2 (N17247, N17243, N8978);
not NOT1 (N17248, N17230);
xor XOR2 (N17249, N17240, N14662);
not NOT1 (N17250, N17226);
not NOT1 (N17251, N17236);
nor NOR3 (N17252, N17215, N3334, N12179);
or OR2 (N17253, N17245, N271);
and AND3 (N17254, N17252, N10132, N14808);
xor XOR2 (N17255, N17238, N15014);
nor NOR3 (N17256, N17247, N2783, N2937);
nand NAND2 (N17257, N17254, N16681);
nand NAND3 (N17258, N17257, N16307, N6248);
nor NOR3 (N17259, N17251, N13681, N3857);
and AND2 (N17260, N17259, N591);
nand NAND4 (N17261, N17249, N12396, N7801, N9996);
or OR4 (N17262, N17258, N6317, N14288, N12531);
not NOT1 (N17263, N17248);
and AND3 (N17264, N17246, N1547, N10214);
not NOT1 (N17265, N17255);
not NOT1 (N17266, N17256);
xor XOR2 (N17267, N17263, N10208);
or OR4 (N17268, N17262, N1737, N8905, N14213);
nor NOR4 (N17269, N17250, N6178, N11099, N15361);
nor NOR3 (N17270, N17266, N2441, N9124);
nand NAND2 (N17271, N17260, N14469);
or OR3 (N17272, N17261, N572, N11765);
nand NAND2 (N17273, N17244, N10025);
xor XOR2 (N17274, N17269, N16545);
nand NAND4 (N17275, N17273, N7258, N1555, N1616);
or OR2 (N17276, N17268, N17127);
or OR4 (N17277, N17253, N412, N5524, N1713);
nand NAND4 (N17278, N17275, N16422, N17169, N423);
not NOT1 (N17279, N17272);
or OR3 (N17280, N17276, N10120, N9915);
buf BUF1 (N17281, N17264);
xor XOR2 (N17282, N17277, N7769);
nor NOR3 (N17283, N17270, N11666, N3109);
buf BUF1 (N17284, N17280);
or OR3 (N17285, N17284, N16348, N5645);
and AND4 (N17286, N17281, N8947, N10018, N5181);
nand NAND2 (N17287, N17279, N3990);
and AND4 (N17288, N17267, N6579, N1363, N17081);
not NOT1 (N17289, N17285);
and AND4 (N17290, N17283, N14578, N5554, N15699);
xor XOR2 (N17291, N17271, N13977);
buf BUF1 (N17292, N17265);
buf BUF1 (N17293, N17291);
nand NAND3 (N17294, N17274, N2574, N5738);
nor NOR3 (N17295, N17289, N3006, N15365);
buf BUF1 (N17296, N17292);
xor XOR2 (N17297, N17294, N3872);
buf BUF1 (N17298, N17278);
buf BUF1 (N17299, N17288);
xor XOR2 (N17300, N17287, N1636);
not NOT1 (N17301, N17290);
nand NAND2 (N17302, N17299, N3802);
xor XOR2 (N17303, N17282, N11240);
and AND2 (N17304, N17297, N6223);
nand NAND4 (N17305, N17300, N1463, N3489, N16884);
nand NAND2 (N17306, N17293, N15172);
xor XOR2 (N17307, N17304, N7260);
buf BUF1 (N17308, N17306);
or OR3 (N17309, N17301, N5287, N3015);
or OR4 (N17310, N17298, N6140, N16044, N11682);
nand NAND4 (N17311, N17308, N5890, N3733, N7860);
buf BUF1 (N17312, N17295);
nand NAND4 (N17313, N17303, N1553, N16344, N1880);
or OR2 (N17314, N17313, N13594);
nand NAND2 (N17315, N17312, N6719);
buf BUF1 (N17316, N17302);
nand NAND2 (N17317, N17315, N7859);
not NOT1 (N17318, N17305);
and AND3 (N17319, N17318, N3162, N1116);
and AND2 (N17320, N17296, N5715);
or OR3 (N17321, N17317, N15202, N8045);
and AND2 (N17322, N17310, N15747);
buf BUF1 (N17323, N17319);
buf BUF1 (N17324, N17307);
buf BUF1 (N17325, N17309);
buf BUF1 (N17326, N17311);
buf BUF1 (N17327, N17321);
buf BUF1 (N17328, N17286);
and AND3 (N17329, N17327, N8093, N8914);
nor NOR3 (N17330, N17320, N8297, N62);
nand NAND4 (N17331, N17322, N6018, N3135, N16844);
not NOT1 (N17332, N17328);
and AND4 (N17333, N17329, N1197, N12306, N16037);
xor XOR2 (N17334, N17316, N3312);
nor NOR2 (N17335, N17332, N13871);
nand NAND2 (N17336, N17335, N3527);
and AND4 (N17337, N17334, N13420, N13133, N5236);
or OR4 (N17338, N17324, N10351, N15328, N13774);
and AND4 (N17339, N17336, N12516, N734, N4771);
or OR2 (N17340, N17338, N664);
xor XOR2 (N17341, N17314, N14597);
xor XOR2 (N17342, N17337, N9767);
buf BUF1 (N17343, N17339);
not NOT1 (N17344, N17341);
or OR2 (N17345, N17323, N9066);
buf BUF1 (N17346, N17345);
or OR2 (N17347, N17340, N5045);
or OR2 (N17348, N17346, N5545);
or OR3 (N17349, N17326, N12608, N3417);
nand NAND4 (N17350, N17344, N13261, N4768, N7944);
and AND3 (N17351, N17333, N12385, N12648);
nor NOR3 (N17352, N17325, N7828, N3835);
and AND4 (N17353, N17343, N4453, N10840, N9793);
or OR2 (N17354, N17348, N1482);
or OR3 (N17355, N17351, N15901, N8046);
or OR2 (N17356, N17342, N10017);
not NOT1 (N17357, N17330);
and AND4 (N17358, N17355, N1357, N8674, N1917);
or OR4 (N17359, N17352, N11910, N9725, N5709);
not NOT1 (N17360, N17350);
and AND2 (N17361, N17357, N4397);
nand NAND4 (N17362, N17361, N6083, N8887, N4846);
xor XOR2 (N17363, N17354, N5402);
not NOT1 (N17364, N17347);
and AND3 (N17365, N17358, N5927, N15796);
or OR2 (N17366, N17356, N2116);
buf BUF1 (N17367, N17362);
not NOT1 (N17368, N17349);
xor XOR2 (N17369, N17363, N5526);
not NOT1 (N17370, N17366);
or OR4 (N17371, N17365, N12260, N2413, N8063);
or OR3 (N17372, N17360, N12856, N1107);
nor NOR3 (N17373, N17369, N1734, N17267);
or OR2 (N17374, N17367, N13403);
nand NAND4 (N17375, N17368, N16324, N11260, N3142);
not NOT1 (N17376, N17375);
not NOT1 (N17377, N17364);
or OR3 (N17378, N17374, N16177, N323);
buf BUF1 (N17379, N17371);
buf BUF1 (N17380, N17372);
nand NAND3 (N17381, N17353, N13621, N5234);
and AND2 (N17382, N17359, N6290);
not NOT1 (N17383, N17377);
not NOT1 (N17384, N17331);
buf BUF1 (N17385, N17378);
nand NAND2 (N17386, N17380, N1114);
not NOT1 (N17387, N17379);
xor XOR2 (N17388, N17376, N12255);
not NOT1 (N17389, N17383);
nand NAND3 (N17390, N17381, N6219, N14872);
and AND3 (N17391, N17387, N13591, N3410);
nand NAND2 (N17392, N17388, N838);
or OR4 (N17393, N17370, N8299, N17142, N1617);
or OR3 (N17394, N17389, N15939, N9327);
buf BUF1 (N17395, N17391);
and AND4 (N17396, N17373, N12695, N3372, N12963);
not NOT1 (N17397, N17393);
xor XOR2 (N17398, N17386, N3676);
not NOT1 (N17399, N17398);
nor NOR2 (N17400, N17399, N11927);
nor NOR3 (N17401, N17394, N12298, N5533);
xor XOR2 (N17402, N17384, N8952);
and AND4 (N17403, N17382, N2392, N7138, N10205);
nor NOR4 (N17404, N17403, N3154, N12193, N4166);
xor XOR2 (N17405, N17392, N14973);
and AND3 (N17406, N17395, N5410, N12513);
buf BUF1 (N17407, N17401);
nand NAND3 (N17408, N17400, N3089, N10832);
xor XOR2 (N17409, N17405, N13718);
nand NAND3 (N17410, N17407, N8951, N11155);
not NOT1 (N17411, N17397);
nand NAND2 (N17412, N17396, N16735);
nor NOR4 (N17413, N17412, N5265, N16419, N24);
nand NAND2 (N17414, N17409, N15831);
xor XOR2 (N17415, N17411, N15515);
not NOT1 (N17416, N17414);
buf BUF1 (N17417, N17410);
xor XOR2 (N17418, N17413, N16890);
and AND2 (N17419, N17417, N12766);
and AND3 (N17420, N17419, N300, N7673);
nor NOR4 (N17421, N17416, N1934, N17013, N2483);
and AND3 (N17422, N17421, N1448, N2337);
nand NAND4 (N17423, N17422, N4996, N4600, N3492);
not NOT1 (N17424, N17408);
or OR3 (N17425, N17415, N12983, N6715);
nand NAND3 (N17426, N17390, N9777, N3521);
nor NOR2 (N17427, N17425, N8549);
buf BUF1 (N17428, N17423);
nand NAND2 (N17429, N17385, N14505);
and AND4 (N17430, N17426, N3713, N13592, N4380);
nand NAND2 (N17431, N17429, N1007);
nor NOR3 (N17432, N17428, N10669, N8948);
xor XOR2 (N17433, N17430, N13426);
and AND2 (N17434, N17431, N14068);
buf BUF1 (N17435, N17433);
nand NAND4 (N17436, N17435, N6604, N8089, N2997);
not NOT1 (N17437, N17406);
not NOT1 (N17438, N17436);
and AND2 (N17439, N17437, N5121);
and AND3 (N17440, N17424, N11895, N5774);
buf BUF1 (N17441, N17438);
and AND2 (N17442, N17432, N11176);
not NOT1 (N17443, N17418);
xor XOR2 (N17444, N17443, N3539);
xor XOR2 (N17445, N17427, N4590);
or OR4 (N17446, N17434, N11918, N6882, N6209);
and AND4 (N17447, N17445, N5168, N12386, N14810);
and AND2 (N17448, N17441, N11898);
nand NAND4 (N17449, N17447, N16886, N15408, N16654);
xor XOR2 (N17450, N17420, N5043);
not NOT1 (N17451, N17448);
not NOT1 (N17452, N17451);
nor NOR2 (N17453, N17402, N2189);
or OR2 (N17454, N17453, N4266);
not NOT1 (N17455, N17446);
nand NAND4 (N17456, N17444, N2562, N5721, N2655);
not NOT1 (N17457, N17449);
and AND3 (N17458, N17455, N7584, N3324);
and AND4 (N17459, N17458, N2250, N12665, N16596);
nand NAND2 (N17460, N17452, N17140);
and AND3 (N17461, N17439, N15172, N6444);
buf BUF1 (N17462, N17450);
buf BUF1 (N17463, N17459);
nand NAND4 (N17464, N17461, N4361, N3207, N6379);
not NOT1 (N17465, N17457);
nand NAND3 (N17466, N17442, N3272, N5224);
xor XOR2 (N17467, N17462, N15932);
xor XOR2 (N17468, N17456, N13033);
or OR4 (N17469, N17404, N5408, N10985, N4148);
and AND3 (N17470, N17468, N12068, N5671);
not NOT1 (N17471, N17460);
and AND3 (N17472, N17440, N4819, N7432);
nor NOR4 (N17473, N17454, N17432, N11779, N16559);
nor NOR4 (N17474, N17472, N12108, N16974, N8228);
and AND2 (N17475, N17465, N11221);
nor NOR2 (N17476, N17464, N5485);
nand NAND4 (N17477, N17475, N16677, N5318, N2120);
buf BUF1 (N17478, N17471);
buf BUF1 (N17479, N17470);
xor XOR2 (N17480, N17476, N6444);
xor XOR2 (N17481, N17479, N10915);
buf BUF1 (N17482, N17474);
and AND4 (N17483, N17473, N17455, N1968, N1114);
nand NAND2 (N17484, N17477, N7009);
nor NOR3 (N17485, N17469, N14552, N305);
or OR4 (N17486, N17484, N204, N9791, N12921);
nor NOR3 (N17487, N17486, N14033, N11116);
or OR2 (N17488, N17481, N12181);
xor XOR2 (N17489, N17463, N13957);
or OR3 (N17490, N17467, N9659, N5282);
buf BUF1 (N17491, N17488);
xor XOR2 (N17492, N17466, N15467);
or OR3 (N17493, N17478, N10387, N16179);
xor XOR2 (N17494, N17489, N11309);
xor XOR2 (N17495, N17483, N4414);
buf BUF1 (N17496, N17487);
or OR2 (N17497, N17493, N7830);
buf BUF1 (N17498, N17480);
and AND2 (N17499, N17482, N2243);
and AND4 (N17500, N17498, N13411, N9748, N11076);
nor NOR3 (N17501, N17495, N16034, N13219);
not NOT1 (N17502, N17499);
not NOT1 (N17503, N17494);
nor NOR2 (N17504, N17491, N10774);
xor XOR2 (N17505, N17500, N11954);
buf BUF1 (N17506, N17496);
nand NAND3 (N17507, N17505, N16791, N1886);
nor NOR4 (N17508, N17485, N2459, N8524, N12113);
buf BUF1 (N17509, N17492);
and AND2 (N17510, N17490, N2530);
and AND2 (N17511, N17506, N13739);
xor XOR2 (N17512, N17507, N4044);
and AND4 (N17513, N17503, N2389, N4767, N7450);
buf BUF1 (N17514, N17497);
or OR2 (N17515, N17513, N8123);
or OR4 (N17516, N17504, N12590, N3808, N16338);
nand NAND3 (N17517, N17514, N9168, N9629);
nor NOR4 (N17518, N17516, N10109, N14938, N3220);
and AND4 (N17519, N17502, N16859, N1378, N3514);
xor XOR2 (N17520, N17508, N2902);
not NOT1 (N17521, N17512);
xor XOR2 (N17522, N17510, N17231);
not NOT1 (N17523, N17511);
nand NAND2 (N17524, N17509, N8869);
not NOT1 (N17525, N17515);
xor XOR2 (N17526, N17523, N1583);
nand NAND4 (N17527, N17518, N3684, N431, N14432);
and AND2 (N17528, N17501, N17134);
xor XOR2 (N17529, N17528, N1521);
buf BUF1 (N17530, N17517);
and AND3 (N17531, N17530, N4324, N11160);
or OR2 (N17532, N17522, N3407);
nand NAND2 (N17533, N17521, N6113);
or OR4 (N17534, N17525, N4698, N2994, N4027);
not NOT1 (N17535, N17526);
xor XOR2 (N17536, N17519, N10399);
xor XOR2 (N17537, N17532, N7740);
xor XOR2 (N17538, N17537, N16222);
buf BUF1 (N17539, N17524);
nor NOR2 (N17540, N17536, N6429);
nand NAND2 (N17541, N17538, N14965);
not NOT1 (N17542, N17541);
buf BUF1 (N17543, N17535);
xor XOR2 (N17544, N17531, N4084);
or OR2 (N17545, N17544, N4663);
xor XOR2 (N17546, N17533, N15921);
nor NOR4 (N17547, N17545, N160, N12502, N4584);
xor XOR2 (N17548, N17529, N1161);
not NOT1 (N17549, N17534);
nor NOR4 (N17550, N17539, N10943, N12988, N5033);
not NOT1 (N17551, N17542);
xor XOR2 (N17552, N17550, N11448);
not NOT1 (N17553, N17527);
and AND4 (N17554, N17547, N15821, N14371, N6202);
nor NOR2 (N17555, N17554, N5882);
nor NOR4 (N17556, N17540, N3272, N11758, N10345);
not NOT1 (N17557, N17553);
nand NAND2 (N17558, N17555, N8848);
xor XOR2 (N17559, N17546, N1573);
not NOT1 (N17560, N17558);
xor XOR2 (N17561, N17559, N15253);
buf BUF1 (N17562, N17552);
not NOT1 (N17563, N17520);
and AND4 (N17564, N17560, N16372, N9010, N17409);
and AND4 (N17565, N17556, N15184, N11795, N14832);
xor XOR2 (N17566, N17562, N8164);
not NOT1 (N17567, N17543);
buf BUF1 (N17568, N17565);
or OR3 (N17569, N17561, N13620, N5971);
nor NOR2 (N17570, N17569, N8839);
nor NOR3 (N17571, N17570, N9745, N4204);
or OR4 (N17572, N17557, N3088, N6812, N6992);
or OR3 (N17573, N17567, N1596, N14472);
and AND3 (N17574, N17571, N8035, N3404);
and AND3 (N17575, N17551, N15371, N17069);
or OR4 (N17576, N17575, N9583, N2410, N8131);
nand NAND4 (N17577, N17572, N11833, N1016, N2025);
buf BUF1 (N17578, N17548);
xor XOR2 (N17579, N17576, N15062);
not NOT1 (N17580, N17564);
buf BUF1 (N17581, N17566);
nor NOR2 (N17582, N17573, N11359);
nor NOR3 (N17583, N17568, N12186, N16236);
or OR4 (N17584, N17574, N1420, N359, N177);
buf BUF1 (N17585, N17563);
xor XOR2 (N17586, N17580, N6117);
buf BUF1 (N17587, N17586);
xor XOR2 (N17588, N17549, N7731);
not NOT1 (N17589, N17578);
nor NOR2 (N17590, N17589, N1910);
nor NOR2 (N17591, N17588, N347);
and AND4 (N17592, N17577, N12900, N96, N62);
and AND2 (N17593, N17585, N8869);
or OR2 (N17594, N17590, N13752);
buf BUF1 (N17595, N17594);
buf BUF1 (N17596, N17595);
or OR4 (N17597, N17581, N8431, N1994, N1622);
nor NOR2 (N17598, N17591, N10526);
or OR3 (N17599, N17584, N7099, N16718);
nor NOR4 (N17600, N17598, N9106, N8131, N9753);
nor NOR3 (N17601, N17593, N1708, N14315);
or OR4 (N17602, N17582, N15742, N3418, N6143);
or OR4 (N17603, N17592, N954, N9395, N5256);
nand NAND4 (N17604, N17603, N4926, N5466, N11560);
nand NAND4 (N17605, N17601, N5423, N4818, N4748);
xor XOR2 (N17606, N17599, N16129);
xor XOR2 (N17607, N17596, N16313);
not NOT1 (N17608, N17587);
nor NOR4 (N17609, N17583, N4138, N8973, N1499);
nand NAND3 (N17610, N17609, N6699, N789);
or OR3 (N17611, N17602, N1340, N16441);
xor XOR2 (N17612, N17605, N7543);
not NOT1 (N17613, N17607);
buf BUF1 (N17614, N17610);
nor NOR2 (N17615, N17606, N10217);
xor XOR2 (N17616, N17614, N15329);
nand NAND2 (N17617, N17604, N7639);
and AND4 (N17618, N17608, N6027, N7429, N11962);
nand NAND4 (N17619, N17617, N1566, N17147, N16435);
nor NOR4 (N17620, N17619, N5883, N12011, N12375);
xor XOR2 (N17621, N17579, N16320);
or OR2 (N17622, N17597, N14634);
nand NAND4 (N17623, N17615, N11580, N6917, N16965);
nor NOR2 (N17624, N17612, N6607);
nor NOR3 (N17625, N17616, N13145, N2850);
nand NAND2 (N17626, N17620, N12193);
buf BUF1 (N17627, N17622);
or OR2 (N17628, N17627, N359);
nand NAND2 (N17629, N17628, N17402);
xor XOR2 (N17630, N17600, N14917);
and AND2 (N17631, N17613, N16711);
xor XOR2 (N17632, N17629, N7728);
nor NOR2 (N17633, N17626, N9201);
and AND2 (N17634, N17631, N7792);
not NOT1 (N17635, N17634);
or OR3 (N17636, N17625, N6427, N11825);
or OR2 (N17637, N17633, N1934);
or OR2 (N17638, N17632, N12594);
nand NAND3 (N17639, N17621, N10929, N13496);
not NOT1 (N17640, N17635);
not NOT1 (N17641, N17611);
not NOT1 (N17642, N17640);
nor NOR3 (N17643, N17624, N2168, N11204);
xor XOR2 (N17644, N17637, N15872);
not NOT1 (N17645, N17639);
buf BUF1 (N17646, N17638);
buf BUF1 (N17647, N17618);
nor NOR4 (N17648, N17630, N6005, N1512, N731);
nor NOR3 (N17649, N17642, N9233, N1026);
or OR3 (N17650, N17645, N1930, N2577);
nor NOR2 (N17651, N17646, N8771);
not NOT1 (N17652, N17623);
nand NAND4 (N17653, N17650, N9660, N17216, N8254);
nor NOR3 (N17654, N17651, N14429, N11945);
nand NAND2 (N17655, N17648, N510);
nand NAND4 (N17656, N17649, N6133, N7386, N14885);
and AND4 (N17657, N17653, N499, N12100, N17411);
or OR3 (N17658, N17647, N16375, N6745);
buf BUF1 (N17659, N17636);
buf BUF1 (N17660, N17659);
xor XOR2 (N17661, N17655, N4048);
and AND3 (N17662, N17641, N6841, N4450);
nand NAND3 (N17663, N17660, N3829, N3089);
buf BUF1 (N17664, N17657);
nand NAND3 (N17665, N17663, N9670, N5136);
or OR4 (N17666, N17658, N1730, N14708, N5629);
nand NAND3 (N17667, N17661, N15238, N10040);
and AND4 (N17668, N17643, N4835, N2763, N12284);
nor NOR2 (N17669, N17665, N4994);
xor XOR2 (N17670, N17669, N7243);
not NOT1 (N17671, N17656);
nor NOR2 (N17672, N17671, N5684);
not NOT1 (N17673, N17654);
or OR3 (N17674, N17664, N10876, N17294);
or OR3 (N17675, N17670, N13094, N6439);
xor XOR2 (N17676, N17675, N9753);
not NOT1 (N17677, N17666);
xor XOR2 (N17678, N17644, N3434);
or OR3 (N17679, N17677, N14859, N16689);
and AND2 (N17680, N17662, N6940);
nor NOR3 (N17681, N17676, N1856, N8703);
nand NAND3 (N17682, N17672, N6882, N9887);
nand NAND3 (N17683, N17682, N5466, N12863);
and AND4 (N17684, N17652, N7309, N1150, N6451);
nand NAND3 (N17685, N17681, N16843, N8994);
xor XOR2 (N17686, N17668, N3335);
not NOT1 (N17687, N17680);
xor XOR2 (N17688, N17674, N4861);
and AND3 (N17689, N17673, N2510, N14511);
nand NAND2 (N17690, N17679, N17509);
or OR2 (N17691, N17684, N11537);
xor XOR2 (N17692, N17691, N5138);
not NOT1 (N17693, N17667);
nand NAND4 (N17694, N17688, N16703, N14553, N4597);
buf BUF1 (N17695, N17689);
nand NAND3 (N17696, N17687, N14909, N13845);
not NOT1 (N17697, N17694);
xor XOR2 (N17698, N17683, N17003);
xor XOR2 (N17699, N17678, N13331);
and AND4 (N17700, N17685, N8037, N13432, N6052);
buf BUF1 (N17701, N17695);
nand NAND4 (N17702, N17692, N738, N9984, N4187);
buf BUF1 (N17703, N17699);
nand NAND4 (N17704, N17702, N7874, N15421, N3847);
nor NOR3 (N17705, N17690, N4135, N351);
nor NOR4 (N17706, N17697, N11629, N10708, N7393);
not NOT1 (N17707, N17696);
buf BUF1 (N17708, N17700);
xor XOR2 (N17709, N17707, N12614);
or OR3 (N17710, N17709, N15154, N15508);
and AND2 (N17711, N17710, N5270);
not NOT1 (N17712, N17705);
xor XOR2 (N17713, N17712, N1585);
not NOT1 (N17714, N17698);
not NOT1 (N17715, N17704);
nand NAND4 (N17716, N17715, N2092, N14826, N4095);
buf BUF1 (N17717, N17701);
xor XOR2 (N17718, N17706, N7852);
xor XOR2 (N17719, N17693, N7446);
not NOT1 (N17720, N17714);
not NOT1 (N17721, N17718);
nor NOR4 (N17722, N17721, N3031, N4995, N7991);
buf BUF1 (N17723, N17711);
nand NAND3 (N17724, N17686, N8064, N8481);
buf BUF1 (N17725, N17716);
or OR2 (N17726, N17724, N10305);
nand NAND2 (N17727, N17703, N17075);
and AND4 (N17728, N17720, N1115, N17531, N17480);
and AND3 (N17729, N17708, N14046, N14235);
and AND4 (N17730, N17729, N6587, N5158, N9207);
or OR3 (N17731, N17717, N6939, N13844);
nor NOR4 (N17732, N17730, N3376, N10993, N3344);
xor XOR2 (N17733, N17732, N13246);
or OR4 (N17734, N17731, N7209, N9819, N4971);
nand NAND4 (N17735, N17734, N7992, N1407, N10525);
not NOT1 (N17736, N17722);
nand NAND4 (N17737, N17728, N7520, N12754, N4616);
buf BUF1 (N17738, N17719);
nand NAND3 (N17739, N17726, N7967, N2134);
xor XOR2 (N17740, N17736, N11869);
and AND3 (N17741, N17740, N6599, N8296);
and AND4 (N17742, N17738, N11772, N2068, N13464);
nor NOR3 (N17743, N17742, N14324, N3607);
or OR4 (N17744, N17723, N10925, N3233, N14455);
not NOT1 (N17745, N17737);
not NOT1 (N17746, N17741);
xor XOR2 (N17747, N17713, N7851);
or OR3 (N17748, N17739, N11768, N11385);
xor XOR2 (N17749, N17727, N13961);
nor NOR4 (N17750, N17725, N3717, N8343, N1999);
and AND4 (N17751, N17744, N13983, N13351, N6383);
nand NAND4 (N17752, N17749, N8595, N16926, N5023);
xor XOR2 (N17753, N17745, N16324);
nand NAND4 (N17754, N17743, N57, N8915, N7478);
and AND4 (N17755, N17735, N11714, N8019, N16271);
xor XOR2 (N17756, N17750, N8246);
nand NAND2 (N17757, N17751, N14573);
xor XOR2 (N17758, N17752, N11078);
xor XOR2 (N17759, N17746, N4868);
nand NAND4 (N17760, N17754, N7472, N7913, N6882);
xor XOR2 (N17761, N17747, N8400);
xor XOR2 (N17762, N17758, N7921);
nand NAND2 (N17763, N17733, N8693);
not NOT1 (N17764, N17763);
buf BUF1 (N17765, N17760);
buf BUF1 (N17766, N17757);
buf BUF1 (N17767, N17766);
nand NAND2 (N17768, N17756, N7322);
or OR3 (N17769, N17755, N15480, N12787);
xor XOR2 (N17770, N17767, N12816);
xor XOR2 (N17771, N17764, N7410);
buf BUF1 (N17772, N17769);
not NOT1 (N17773, N17772);
nor NOR2 (N17774, N17748, N3675);
not NOT1 (N17775, N17770);
nor NOR3 (N17776, N17774, N785, N7589);
nor NOR3 (N17777, N17773, N7023, N16982);
not NOT1 (N17778, N17775);
or OR2 (N17779, N17759, N12049);
and AND2 (N17780, N17762, N17750);
not NOT1 (N17781, N17779);
or OR4 (N17782, N17761, N6731, N16570, N1335);
buf BUF1 (N17783, N17782);
nand NAND3 (N17784, N17765, N3443, N15506);
or OR2 (N17785, N17777, N8175);
not NOT1 (N17786, N17783);
nor NOR2 (N17787, N17778, N16573);
xor XOR2 (N17788, N17787, N2135);
buf BUF1 (N17789, N17785);
nor NOR3 (N17790, N17780, N14123, N7854);
or OR2 (N17791, N17771, N8436);
and AND2 (N17792, N17791, N15406);
and AND4 (N17793, N17776, N7152, N9498, N3620);
nor NOR2 (N17794, N17753, N12915);
buf BUF1 (N17795, N17786);
or OR4 (N17796, N17768, N13864, N2788, N6673);
not NOT1 (N17797, N17794);
nand NAND2 (N17798, N17795, N4614);
and AND3 (N17799, N17798, N4389, N3365);
or OR4 (N17800, N17793, N7158, N2751, N5790);
xor XOR2 (N17801, N17784, N12668);
buf BUF1 (N17802, N17800);
not NOT1 (N17803, N17792);
nand NAND4 (N17804, N17781, N4471, N16027, N11045);
nand NAND2 (N17805, N17796, N15672);
and AND4 (N17806, N17797, N12158, N3664, N14970);
nor NOR3 (N17807, N17788, N3943, N3912);
nand NAND4 (N17808, N17801, N10891, N15927, N1816);
not NOT1 (N17809, N17808);
and AND2 (N17810, N17807, N7347);
and AND3 (N17811, N17790, N3614, N10527);
buf BUF1 (N17812, N17810);
buf BUF1 (N17813, N17811);
nor NOR2 (N17814, N17799, N5056);
nor NOR3 (N17815, N17802, N11638, N13163);
nor NOR2 (N17816, N17789, N13536);
and AND3 (N17817, N17813, N1716, N15239);
not NOT1 (N17818, N17804);
and AND2 (N17819, N17806, N1441);
buf BUF1 (N17820, N17817);
not NOT1 (N17821, N17812);
nor NOR3 (N17822, N17818, N12607, N12291);
buf BUF1 (N17823, N17803);
nand NAND2 (N17824, N17809, N5691);
or OR4 (N17825, N17814, N15854, N3942, N10437);
not NOT1 (N17826, N17819);
buf BUF1 (N17827, N17816);
not NOT1 (N17828, N17824);
nor NOR3 (N17829, N17823, N78, N7244);
not NOT1 (N17830, N17825);
nor NOR4 (N17831, N17826, N13485, N2997, N6484);
not NOT1 (N17832, N17828);
or OR3 (N17833, N17829, N14016, N13740);
buf BUF1 (N17834, N17821);
and AND4 (N17835, N17815, N17201, N3433, N2493);
xor XOR2 (N17836, N17827, N14030);
not NOT1 (N17837, N17834);
buf BUF1 (N17838, N17835);
nand NAND4 (N17839, N17833, N5267, N763, N16018);
and AND4 (N17840, N17822, N8170, N10195, N7056);
nor NOR2 (N17841, N17840, N33);
and AND4 (N17842, N17837, N2517, N335, N8214);
nand NAND4 (N17843, N17839, N7719, N9454, N14039);
buf BUF1 (N17844, N17836);
and AND3 (N17845, N17820, N7792, N16500);
not NOT1 (N17846, N17831);
or OR3 (N17847, N17842, N6543, N9554);
not NOT1 (N17848, N17844);
not NOT1 (N17849, N17846);
buf BUF1 (N17850, N17845);
xor XOR2 (N17851, N17838, N6230);
nand NAND2 (N17852, N17832, N13557);
and AND2 (N17853, N17849, N12736);
xor XOR2 (N17854, N17850, N4925);
xor XOR2 (N17855, N17848, N5424);
nand NAND4 (N17856, N17805, N16903, N6501, N7300);
nand NAND3 (N17857, N17853, N8460, N384);
and AND2 (N17858, N17851, N7783);
or OR3 (N17859, N17830, N6358, N1381);
or OR4 (N17860, N17856, N12724, N4434, N8417);
not NOT1 (N17861, N17841);
nor NOR3 (N17862, N17855, N8454, N11100);
nand NAND4 (N17863, N17861, N7758, N1336, N2059);
or OR2 (N17864, N17859, N3361);
nand NAND2 (N17865, N17858, N16648);
buf BUF1 (N17866, N17854);
xor XOR2 (N17867, N17866, N13731);
and AND3 (N17868, N17852, N9120, N7731);
xor XOR2 (N17869, N17868, N9711);
nand NAND4 (N17870, N17867, N4089, N11853, N9797);
buf BUF1 (N17871, N17865);
not NOT1 (N17872, N17847);
not NOT1 (N17873, N17864);
or OR2 (N17874, N17870, N13858);
nand NAND4 (N17875, N17871, N3792, N5973, N10738);
xor XOR2 (N17876, N17860, N5102);
not NOT1 (N17877, N17869);
or OR2 (N17878, N17863, N9625);
nor NOR2 (N17879, N17877, N1452);
xor XOR2 (N17880, N17874, N17266);
and AND2 (N17881, N17879, N6136);
not NOT1 (N17882, N17881);
not NOT1 (N17883, N17876);
not NOT1 (N17884, N17862);
nand NAND3 (N17885, N17843, N7832, N7237);
not NOT1 (N17886, N17878);
and AND4 (N17887, N17884, N11228, N10819, N6312);
nand NAND3 (N17888, N17886, N346, N7199);
buf BUF1 (N17889, N17880);
nand NAND4 (N17890, N17882, N10969, N9390, N16946);
buf BUF1 (N17891, N17883);
buf BUF1 (N17892, N17857);
or OR3 (N17893, N17890, N1417, N5443);
or OR3 (N17894, N17887, N17458, N5647);
buf BUF1 (N17895, N17888);
and AND3 (N17896, N17875, N9037, N17687);
buf BUF1 (N17897, N17894);
buf BUF1 (N17898, N17889);
nor NOR2 (N17899, N17892, N6156);
nand NAND4 (N17900, N17873, N687, N3171, N16764);
buf BUF1 (N17901, N17898);
xor XOR2 (N17902, N17897, N15753);
xor XOR2 (N17903, N17885, N14270);
and AND3 (N17904, N17901, N15408, N3845);
xor XOR2 (N17905, N17904, N4202);
not NOT1 (N17906, N17896);
not NOT1 (N17907, N17900);
or OR3 (N17908, N17907, N10015, N12775);
nor NOR2 (N17909, N17905, N16576);
and AND3 (N17910, N17872, N12034, N418);
not NOT1 (N17911, N17906);
and AND3 (N17912, N17902, N10944, N9138);
or OR4 (N17913, N17908, N13934, N3983, N10801);
or OR3 (N17914, N17913, N2596, N1218);
buf BUF1 (N17915, N17912);
and AND2 (N17916, N17914, N1772);
xor XOR2 (N17917, N17891, N8611);
not NOT1 (N17918, N17916);
buf BUF1 (N17919, N17909);
xor XOR2 (N17920, N17911, N11856);
not NOT1 (N17921, N17893);
buf BUF1 (N17922, N17895);
buf BUF1 (N17923, N17918);
nand NAND3 (N17924, N17917, N9247, N6805);
not NOT1 (N17925, N17922);
not NOT1 (N17926, N17915);
nor NOR3 (N17927, N17903, N14200, N9810);
nor NOR2 (N17928, N17921, N3325);
not NOT1 (N17929, N17925);
not NOT1 (N17930, N17929);
and AND3 (N17931, N17928, N14631, N12431);
not NOT1 (N17932, N17923);
nor NOR4 (N17933, N17920, N3571, N2784, N10997);
and AND3 (N17934, N17924, N16977, N7845);
and AND2 (N17935, N17910, N4459);
buf BUF1 (N17936, N17933);
buf BUF1 (N17937, N17927);
xor XOR2 (N17938, N17899, N5792);
and AND2 (N17939, N17934, N13115);
not NOT1 (N17940, N17939);
nor NOR4 (N17941, N17931, N10033, N16972, N12578);
not NOT1 (N17942, N17930);
or OR4 (N17943, N17940, N5814, N14701, N2544);
nand NAND3 (N17944, N17937, N10364, N13041);
nor NOR3 (N17945, N17935, N13804, N10453);
xor XOR2 (N17946, N17932, N16567);
xor XOR2 (N17947, N17946, N2531);
xor XOR2 (N17948, N17943, N16983);
buf BUF1 (N17949, N17948);
buf BUF1 (N17950, N17938);
and AND4 (N17951, N17950, N9826, N16777, N8033);
not NOT1 (N17952, N17941);
xor XOR2 (N17953, N17949, N2127);
nand NAND3 (N17954, N17953, N14939, N5213);
not NOT1 (N17955, N17919);
or OR4 (N17956, N17954, N1630, N5010, N4697);
buf BUF1 (N17957, N17926);
xor XOR2 (N17958, N17947, N2342);
buf BUF1 (N17959, N17955);
nor NOR4 (N17960, N17952, N9270, N7336, N9583);
or OR4 (N17961, N17942, N16948, N7797, N2370);
not NOT1 (N17962, N17961);
nor NOR4 (N17963, N17936, N10019, N16646, N16924);
buf BUF1 (N17964, N17944);
xor XOR2 (N17965, N17963, N14469);
nand NAND2 (N17966, N17965, N3825);
xor XOR2 (N17967, N17956, N10978);
nor NOR2 (N17968, N17962, N14491);
xor XOR2 (N17969, N17945, N37);
nor NOR4 (N17970, N17957, N12706, N2110, N8901);
xor XOR2 (N17971, N17959, N3245);
nor NOR3 (N17972, N17964, N1517, N4385);
nor NOR4 (N17973, N17967, N15955, N8095, N6417);
or OR3 (N17974, N17970, N9497, N10284);
not NOT1 (N17975, N17972);
and AND3 (N17976, N17974, N5787, N64);
nor NOR3 (N17977, N17951, N171, N9357);
nor NOR4 (N17978, N17968, N17687, N2595, N14458);
or OR2 (N17979, N17973, N961);
and AND3 (N17980, N17969, N12053, N5467);
nand NAND3 (N17981, N17975, N9835, N11433);
buf BUF1 (N17982, N17979);
nand NAND2 (N17983, N17971, N6609);
and AND2 (N17984, N17958, N6413);
and AND3 (N17985, N17976, N15014, N4356);
nor NOR2 (N17986, N17966, N10298);
not NOT1 (N17987, N17982);
nand NAND2 (N17988, N17977, N8410);
and AND4 (N17989, N17981, N12613, N2588, N3478);
nor NOR4 (N17990, N17986, N12983, N6939, N9599);
and AND4 (N17991, N17988, N4337, N7123, N12608);
nand NAND2 (N17992, N17978, N8230);
nor NOR2 (N17993, N17980, N15317);
not NOT1 (N17994, N17993);
nor NOR2 (N17995, N17990, N1558);
xor XOR2 (N17996, N17985, N17459);
and AND3 (N17997, N17960, N4084, N6254);
or OR4 (N17998, N17984, N14818, N12495, N11093);
or OR4 (N17999, N17996, N8567, N4600, N2151);
nand NAND3 (N18000, N17983, N2579, N7311);
and AND4 (N18001, N17998, N2546, N3111, N1869);
xor XOR2 (N18002, N17999, N7750);
or OR4 (N18003, N17994, N13924, N13698, N278);
not NOT1 (N18004, N18000);
not NOT1 (N18005, N17987);
or OR2 (N18006, N17992, N2456);
or OR2 (N18007, N17995, N6980);
xor XOR2 (N18008, N18003, N10821);
nor NOR3 (N18009, N17997, N7932, N343);
xor XOR2 (N18010, N18005, N16488);
nand NAND4 (N18011, N18006, N4710, N16438, N4267);
or OR2 (N18012, N17989, N15520);
buf BUF1 (N18013, N18011);
nor NOR4 (N18014, N18001, N17419, N12042, N8945);
and AND2 (N18015, N18008, N7860);
or OR3 (N18016, N18004, N11347, N16320);
not NOT1 (N18017, N18014);
buf BUF1 (N18018, N18013);
nor NOR2 (N18019, N18002, N2031);
and AND2 (N18020, N18012, N1302);
and AND3 (N18021, N18017, N468, N11880);
buf BUF1 (N18022, N18016);
or OR3 (N18023, N18010, N16582, N2695);
and AND4 (N18024, N17991, N12471, N11851, N1761);
xor XOR2 (N18025, N18018, N5280);
nand NAND2 (N18026, N18007, N8458);
and AND2 (N18027, N18025, N2322);
buf BUF1 (N18028, N18015);
nand NAND4 (N18029, N18028, N6295, N1695, N11366);
or OR2 (N18030, N18022, N11490);
nor NOR4 (N18031, N18021, N7288, N6088, N15340);
and AND4 (N18032, N18020, N9445, N10950, N5357);
or OR4 (N18033, N18027, N7849, N8438, N14856);
and AND2 (N18034, N18032, N13375);
or OR4 (N18035, N18033, N5905, N7158, N4660);
nand NAND2 (N18036, N18031, N6387);
nor NOR4 (N18037, N18030, N12611, N4547, N7348);
and AND2 (N18038, N18009, N15408);
nand NAND2 (N18039, N18034, N13554);
buf BUF1 (N18040, N18029);
and AND4 (N18041, N18040, N3559, N5173, N1931);
not NOT1 (N18042, N18019);
and AND4 (N18043, N18026, N5248, N4290, N11179);
or OR2 (N18044, N18043, N6374);
buf BUF1 (N18045, N18023);
or OR2 (N18046, N18042, N4794);
buf BUF1 (N18047, N18046);
nor NOR3 (N18048, N18037, N15920, N15168);
and AND4 (N18049, N18038, N714, N16068, N7979);
buf BUF1 (N18050, N18041);
or OR2 (N18051, N18024, N11696);
nand NAND4 (N18052, N18047, N12777, N1160, N4159);
nand NAND3 (N18053, N18039, N4614, N17197);
and AND4 (N18054, N18053, N13773, N14712, N1023);
and AND3 (N18055, N18052, N2852, N2543);
buf BUF1 (N18056, N18048);
buf BUF1 (N18057, N18049);
and AND2 (N18058, N18035, N16179);
or OR4 (N18059, N18058, N12201, N119, N5466);
not NOT1 (N18060, N18059);
not NOT1 (N18061, N18055);
and AND2 (N18062, N18050, N7664);
and AND2 (N18063, N18056, N11941);
xor XOR2 (N18064, N18045, N5946);
buf BUF1 (N18065, N18060);
nand NAND3 (N18066, N18054, N6480, N7944);
or OR4 (N18067, N18036, N16824, N7773, N11389);
xor XOR2 (N18068, N18064, N8634);
buf BUF1 (N18069, N18057);
and AND4 (N18070, N18044, N13492, N18042, N5562);
buf BUF1 (N18071, N18065);
nand NAND2 (N18072, N18068, N3717);
nand NAND4 (N18073, N18071, N12707, N3501, N7170);
xor XOR2 (N18074, N18072, N9722);
buf BUF1 (N18075, N18066);
nor NOR2 (N18076, N18067, N16891);
not NOT1 (N18077, N18062);
not NOT1 (N18078, N18074);
xor XOR2 (N18079, N18075, N7560);
nor NOR2 (N18080, N18069, N6062);
xor XOR2 (N18081, N18076, N10692);
nand NAND4 (N18082, N18077, N17272, N16966, N6524);
nand NAND4 (N18083, N18082, N4449, N7335, N14427);
and AND4 (N18084, N18073, N15559, N3944, N5935);
buf BUF1 (N18085, N18080);
xor XOR2 (N18086, N18083, N13703);
buf BUF1 (N18087, N18086);
or OR4 (N18088, N18070, N17310, N15266, N6524);
buf BUF1 (N18089, N18063);
nand NAND3 (N18090, N18079, N5959, N11276);
or OR2 (N18091, N18089, N1363);
nand NAND4 (N18092, N18078, N12826, N7401, N3352);
not NOT1 (N18093, N18090);
xor XOR2 (N18094, N18061, N17361);
nor NOR4 (N18095, N18091, N10969, N5848, N7881);
xor XOR2 (N18096, N18084, N12671);
and AND3 (N18097, N18087, N14566, N16396);
and AND4 (N18098, N18095, N14207, N14983, N6122);
buf BUF1 (N18099, N18093);
xor XOR2 (N18100, N18098, N9008);
and AND2 (N18101, N18097, N17716);
buf BUF1 (N18102, N18051);
nor NOR2 (N18103, N18081, N15916);
buf BUF1 (N18104, N18096);
and AND4 (N18105, N18101, N3352, N5173, N16336);
and AND2 (N18106, N18094, N13721);
or OR4 (N18107, N18085, N1921, N13892, N8216);
buf BUF1 (N18108, N18092);
or OR2 (N18109, N18099, N6214);
nand NAND2 (N18110, N18108, N3004);
nor NOR4 (N18111, N18100, N5435, N10959, N8614);
or OR4 (N18112, N18105, N15293, N11037, N1502);
nand NAND4 (N18113, N18088, N4801, N5737, N6783);
xor XOR2 (N18114, N18111, N16366);
nand NAND3 (N18115, N18114, N10581, N2313);
not NOT1 (N18116, N18113);
nor NOR2 (N18117, N18112, N7749);
nor NOR2 (N18118, N18109, N13593);
buf BUF1 (N18119, N18104);
not NOT1 (N18120, N18106);
and AND3 (N18121, N18116, N15360, N16485);
or OR4 (N18122, N18107, N14019, N14664, N7216);
and AND4 (N18123, N18121, N13925, N8040, N8734);
buf BUF1 (N18124, N18120);
buf BUF1 (N18125, N18119);
nand NAND4 (N18126, N18102, N2596, N6824, N854);
buf BUF1 (N18127, N18117);
buf BUF1 (N18128, N18103);
not NOT1 (N18129, N18118);
nand NAND4 (N18130, N18124, N2540, N5041, N6379);
nand NAND3 (N18131, N18129, N17011, N8748);
nor NOR2 (N18132, N18125, N8683);
nand NAND4 (N18133, N18122, N8760, N5285, N16383);
and AND4 (N18134, N18110, N7367, N3708, N16757);
not NOT1 (N18135, N18131);
xor XOR2 (N18136, N18132, N16902);
or OR2 (N18137, N18133, N169);
and AND3 (N18138, N18127, N4481, N2297);
or OR3 (N18139, N18134, N13234, N14829);
or OR4 (N18140, N18136, N1491, N7887, N8640);
nor NOR4 (N18141, N18130, N13812, N2290, N2635);
buf BUF1 (N18142, N18135);
and AND2 (N18143, N18115, N5837);
and AND4 (N18144, N18137, N11036, N1845, N2589);
buf BUF1 (N18145, N18126);
or OR2 (N18146, N18139, N9283);
buf BUF1 (N18147, N18123);
xor XOR2 (N18148, N18140, N3484);
nor NOR2 (N18149, N18138, N1855);
nand NAND3 (N18150, N18128, N4149, N13026);
and AND2 (N18151, N18149, N5131);
xor XOR2 (N18152, N18150, N14399);
or OR3 (N18153, N18145, N12781, N10010);
nor NOR2 (N18154, N18152, N5005);
xor XOR2 (N18155, N18142, N2940);
nand NAND2 (N18156, N18151, N1712);
xor XOR2 (N18157, N18147, N7712);
not NOT1 (N18158, N18144);
xor XOR2 (N18159, N18148, N5173);
buf BUF1 (N18160, N18143);
nor NOR2 (N18161, N18153, N11264);
and AND2 (N18162, N18146, N16953);
or OR3 (N18163, N18161, N977, N2604);
not NOT1 (N18164, N18163);
not NOT1 (N18165, N18159);
nand NAND2 (N18166, N18155, N9372);
buf BUF1 (N18167, N18141);
not NOT1 (N18168, N18157);
nor NOR2 (N18169, N18154, N10702);
and AND4 (N18170, N18158, N7779, N17442, N11323);
nor NOR4 (N18171, N18168, N12515, N2671, N14927);
xor XOR2 (N18172, N18165, N5681);
not NOT1 (N18173, N18162);
buf BUF1 (N18174, N18164);
or OR4 (N18175, N18172, N5768, N13728, N1495);
or OR4 (N18176, N18170, N8020, N16464, N16549);
xor XOR2 (N18177, N18175, N6947);
buf BUF1 (N18178, N18156);
and AND2 (N18179, N18177, N18131);
buf BUF1 (N18180, N18160);
and AND2 (N18181, N18166, N5738);
or OR3 (N18182, N18171, N11002, N8997);
or OR2 (N18183, N18169, N17073);
or OR4 (N18184, N18181, N3227, N18181, N2100);
and AND3 (N18185, N18167, N6831, N6601);
xor XOR2 (N18186, N18183, N1563);
nor NOR2 (N18187, N18184, N6289);
buf BUF1 (N18188, N18186);
nor NOR3 (N18189, N18176, N4199, N13420);
or OR4 (N18190, N18174, N598, N17254, N13948);
nand NAND3 (N18191, N18178, N14371, N5405);
not NOT1 (N18192, N18180);
not NOT1 (N18193, N18190);
nand NAND4 (N18194, N18189, N17947, N3842, N2384);
nand NAND4 (N18195, N18193, N16301, N14943, N16738);
xor XOR2 (N18196, N18195, N6203);
or OR2 (N18197, N18179, N1648);
buf BUF1 (N18198, N18187);
buf BUF1 (N18199, N18188);
not NOT1 (N18200, N18182);
or OR4 (N18201, N18192, N14576, N4982, N6756);
or OR4 (N18202, N18201, N17573, N6029, N9942);
or OR2 (N18203, N18199, N4130);
or OR3 (N18204, N18185, N14128, N6901);
nand NAND4 (N18205, N18196, N8403, N14054, N3709);
xor XOR2 (N18206, N18198, N2455);
buf BUF1 (N18207, N18205);
nand NAND2 (N18208, N18202, N8376);
xor XOR2 (N18209, N18208, N16346);
buf BUF1 (N18210, N18191);
nand NAND2 (N18211, N18200, N736);
buf BUF1 (N18212, N18210);
nor NOR4 (N18213, N18211, N8248, N11181, N9355);
xor XOR2 (N18214, N18206, N10532);
xor XOR2 (N18215, N18213, N6809);
nand NAND4 (N18216, N18203, N196, N13270, N7603);
or OR4 (N18217, N18197, N2474, N16054, N17796);
or OR3 (N18218, N18216, N18193, N9057);
and AND3 (N18219, N18209, N17495, N7147);
buf BUF1 (N18220, N18173);
nor NOR3 (N18221, N18212, N5675, N5390);
buf BUF1 (N18222, N18219);
xor XOR2 (N18223, N18218, N15692);
not NOT1 (N18224, N18217);
or OR3 (N18225, N18214, N14740, N10556);
nand NAND2 (N18226, N18221, N16506);
and AND3 (N18227, N18207, N12569, N618);
xor XOR2 (N18228, N18204, N3784);
or OR3 (N18229, N18225, N9317, N12927);
or OR4 (N18230, N18220, N5028, N627, N576);
xor XOR2 (N18231, N18224, N11374);
nor NOR2 (N18232, N18215, N6360);
buf BUF1 (N18233, N18194);
and AND3 (N18234, N18230, N5958, N1059);
and AND4 (N18235, N18228, N9563, N17899, N6908);
buf BUF1 (N18236, N18232);
buf BUF1 (N18237, N18231);
not NOT1 (N18238, N18223);
nor NOR2 (N18239, N18226, N13182);
nand NAND2 (N18240, N18222, N6107);
nor NOR2 (N18241, N18235, N17722);
xor XOR2 (N18242, N18234, N3002);
or OR2 (N18243, N18233, N5844);
buf BUF1 (N18244, N18240);
nor NOR3 (N18245, N18241, N5933, N2904);
or OR2 (N18246, N18237, N14054);
buf BUF1 (N18247, N18244);
nand NAND2 (N18248, N18239, N7302);
nand NAND4 (N18249, N18242, N2975, N8206, N4977);
or OR3 (N18250, N18227, N11572, N7223);
xor XOR2 (N18251, N18238, N11029);
nand NAND4 (N18252, N18245, N14180, N6765, N6452);
or OR2 (N18253, N18236, N2814);
nand NAND3 (N18254, N18243, N14756, N17222);
or OR3 (N18255, N18248, N14224, N11106);
not NOT1 (N18256, N18246);
nor NOR4 (N18257, N18255, N15510, N3204, N3643);
nor NOR3 (N18258, N18256, N11467, N15944);
nor NOR4 (N18259, N18229, N4850, N7796, N10229);
and AND3 (N18260, N18251, N9261, N11299);
not NOT1 (N18261, N18257);
not NOT1 (N18262, N18253);
or OR4 (N18263, N18262, N15586, N4317, N7301);
xor XOR2 (N18264, N18260, N11631);
not NOT1 (N18265, N18261);
buf BUF1 (N18266, N18254);
or OR2 (N18267, N18258, N9718);
not NOT1 (N18268, N18263);
nor NOR4 (N18269, N18266, N10541, N18148, N1303);
nand NAND3 (N18270, N18252, N3592, N16373);
nand NAND4 (N18271, N18247, N4331, N274, N5391);
buf BUF1 (N18272, N18265);
nor NOR2 (N18273, N18270, N3381);
xor XOR2 (N18274, N18271, N14365);
nor NOR2 (N18275, N18273, N12469);
or OR2 (N18276, N18249, N8656);
nand NAND2 (N18277, N18274, N15878);
xor XOR2 (N18278, N18267, N13878);
and AND2 (N18279, N18278, N6549);
or OR3 (N18280, N18268, N12079, N10619);
nor NOR3 (N18281, N18250, N17918, N4664);
and AND3 (N18282, N18269, N755, N11039);
xor XOR2 (N18283, N18264, N5214);
not NOT1 (N18284, N18277);
nand NAND2 (N18285, N18281, N15658);
and AND2 (N18286, N18284, N4834);
and AND3 (N18287, N18286, N2627, N10199);
not NOT1 (N18288, N18279);
nand NAND4 (N18289, N18272, N12996, N13998, N7356);
not NOT1 (N18290, N18283);
buf BUF1 (N18291, N18290);
nand NAND3 (N18292, N18275, N8975, N7301);
nor NOR2 (N18293, N18285, N9120);
not NOT1 (N18294, N18287);
or OR2 (N18295, N18288, N14401);
xor XOR2 (N18296, N18280, N695);
or OR3 (N18297, N18289, N15086, N12994);
or OR3 (N18298, N18293, N16284, N946);
not NOT1 (N18299, N18292);
xor XOR2 (N18300, N18296, N13893);
not NOT1 (N18301, N18300);
nor NOR4 (N18302, N18291, N8609, N13487, N15746);
not NOT1 (N18303, N18299);
nor NOR4 (N18304, N18303, N2498, N7762, N12271);
or OR3 (N18305, N18276, N17485, N6931);
or OR3 (N18306, N18282, N8784, N5645);
xor XOR2 (N18307, N18305, N2065);
nand NAND3 (N18308, N18306, N7999, N10288);
and AND3 (N18309, N18298, N15613, N3067);
nor NOR3 (N18310, N18307, N1899, N11706);
xor XOR2 (N18311, N18309, N15588);
buf BUF1 (N18312, N18294);
nand NAND3 (N18313, N18302, N16008, N14064);
not NOT1 (N18314, N18295);
and AND2 (N18315, N18297, N347);
nand NAND4 (N18316, N18308, N18246, N8527, N16374);
and AND2 (N18317, N18315, N17122);
and AND3 (N18318, N18259, N4304, N9595);
or OR3 (N18319, N18314, N11480, N1345);
nand NAND2 (N18320, N18316, N11259);
nand NAND2 (N18321, N18304, N4926);
nor NOR2 (N18322, N18318, N10812);
or OR3 (N18323, N18310, N3756, N14823);
buf BUF1 (N18324, N18323);
not NOT1 (N18325, N18312);
or OR3 (N18326, N18301, N16013, N3940);
buf BUF1 (N18327, N18325);
nor NOR3 (N18328, N18326, N11123, N13546);
and AND2 (N18329, N18322, N3622);
buf BUF1 (N18330, N18327);
nand NAND3 (N18331, N18329, N16682, N8154);
xor XOR2 (N18332, N18313, N16459);
not NOT1 (N18333, N18311);
buf BUF1 (N18334, N18333);
and AND2 (N18335, N18332, N14714);
not NOT1 (N18336, N18321);
buf BUF1 (N18337, N18324);
nand NAND4 (N18338, N18335, N7312, N4836, N3617);
nor NOR4 (N18339, N18337, N3521, N10791, N4718);
and AND2 (N18340, N18331, N3993);
xor XOR2 (N18341, N18317, N1896);
or OR4 (N18342, N18334, N4965, N9251, N3342);
and AND4 (N18343, N18340, N3266, N3781, N2588);
nand NAND4 (N18344, N18338, N3838, N17139, N15160);
and AND3 (N18345, N18343, N14841, N4920);
not NOT1 (N18346, N18320);
and AND2 (N18347, N18330, N15556);
xor XOR2 (N18348, N18328, N10781);
nor NOR2 (N18349, N18341, N13993);
buf BUF1 (N18350, N18344);
nor NOR3 (N18351, N18347, N5798, N11952);
and AND3 (N18352, N18348, N6963, N12937);
or OR3 (N18353, N18352, N10270, N5728);
nand NAND4 (N18354, N18351, N2513, N8187, N3220);
nor NOR4 (N18355, N18353, N13609, N2826, N15832);
nand NAND3 (N18356, N18350, N10710, N4210);
or OR3 (N18357, N18342, N15279, N3086);
nand NAND4 (N18358, N18349, N15281, N9194, N7234);
nand NAND2 (N18359, N18319, N18073);
or OR2 (N18360, N18345, N3139);
xor XOR2 (N18361, N18339, N6778);
buf BUF1 (N18362, N18336);
nor NOR3 (N18363, N18360, N13460, N11216);
buf BUF1 (N18364, N18354);
nor NOR4 (N18365, N18364, N11637, N12277, N15688);
nor NOR3 (N18366, N18361, N13633, N17397);
xor XOR2 (N18367, N18355, N7744);
buf BUF1 (N18368, N18358);
nor NOR2 (N18369, N18346, N3928);
nor NOR2 (N18370, N18356, N15997);
not NOT1 (N18371, N18359);
and AND4 (N18372, N18366, N13308, N6746, N12823);
nor NOR3 (N18373, N18370, N16885, N3779);
not NOT1 (N18374, N18365);
or OR3 (N18375, N18368, N16244, N8106);
or OR4 (N18376, N18362, N4989, N10836, N420);
and AND3 (N18377, N18375, N14280, N18285);
not NOT1 (N18378, N18367);
not NOT1 (N18379, N18378);
and AND4 (N18380, N18377, N18182, N8320, N5676);
nand NAND3 (N18381, N18376, N6255, N3559);
nor NOR2 (N18382, N18357, N9843);
buf BUF1 (N18383, N18382);
not NOT1 (N18384, N18381);
or OR3 (N18385, N18369, N17700, N6985);
not NOT1 (N18386, N18374);
not NOT1 (N18387, N18384);
buf BUF1 (N18388, N18363);
nand NAND4 (N18389, N18371, N3069, N10802, N17338);
or OR4 (N18390, N18385, N17705, N6297, N1174);
nor NOR2 (N18391, N18386, N1291);
nand NAND3 (N18392, N18391, N7321, N7868);
xor XOR2 (N18393, N18383, N5718);
nor NOR4 (N18394, N18392, N1325, N14417, N969);
not NOT1 (N18395, N18373);
buf BUF1 (N18396, N18387);
buf BUF1 (N18397, N18388);
xor XOR2 (N18398, N18390, N17569);
nor NOR4 (N18399, N18389, N12759, N12713, N1158);
buf BUF1 (N18400, N18394);
not NOT1 (N18401, N18380);
and AND3 (N18402, N18393, N2915, N7286);
xor XOR2 (N18403, N18400, N1699);
nand NAND4 (N18404, N18372, N11889, N8497, N13071);
not NOT1 (N18405, N18401);
not NOT1 (N18406, N18403);
not NOT1 (N18407, N18405);
nand NAND2 (N18408, N18404, N1520);
nand NAND2 (N18409, N18407, N7975);
nand NAND2 (N18410, N18397, N4336);
nand NAND2 (N18411, N18399, N14166);
buf BUF1 (N18412, N18396);
buf BUF1 (N18413, N18408);
nand NAND2 (N18414, N18402, N3370);
xor XOR2 (N18415, N18395, N13256);
and AND2 (N18416, N18413, N71);
buf BUF1 (N18417, N18409);
nand NAND2 (N18418, N18415, N6806);
and AND4 (N18419, N18410, N2150, N14183, N15133);
not NOT1 (N18420, N18398);
not NOT1 (N18421, N18411);
or OR3 (N18422, N18419, N6250, N4348);
or OR4 (N18423, N18420, N6695, N16278, N9138);
nand NAND4 (N18424, N18422, N5323, N2222, N11481);
xor XOR2 (N18425, N18418, N12820);
buf BUF1 (N18426, N18417);
nor NOR2 (N18427, N18425, N4597);
nor NOR2 (N18428, N18414, N10206);
nor NOR2 (N18429, N18426, N7685);
not NOT1 (N18430, N18429);
nand NAND3 (N18431, N18406, N11525, N17104);
nand NAND4 (N18432, N18430, N4112, N7852, N9456);
buf BUF1 (N18433, N18416);
or OR2 (N18434, N18428, N13990);
buf BUF1 (N18435, N18379);
and AND3 (N18436, N18423, N7908, N8962);
xor XOR2 (N18437, N18434, N12333);
buf BUF1 (N18438, N18431);
and AND4 (N18439, N18412, N8901, N7980, N2625);
nand NAND3 (N18440, N18421, N12588, N13779);
nand NAND2 (N18441, N18424, N12889);
buf BUF1 (N18442, N18436);
xor XOR2 (N18443, N18435, N12013);
xor XOR2 (N18444, N18439, N6887);
and AND3 (N18445, N18440, N12831, N4608);
nand NAND3 (N18446, N18445, N1476, N12896);
nor NOR4 (N18447, N18441, N1198, N17368, N4653);
nor NOR4 (N18448, N18444, N4507, N4484, N2883);
and AND3 (N18449, N18446, N554, N5632);
nand NAND2 (N18450, N18442, N6054);
or OR3 (N18451, N18438, N1893, N11593);
buf BUF1 (N18452, N18433);
nor NOR2 (N18453, N18427, N14758);
not NOT1 (N18454, N18450);
nor NOR4 (N18455, N18451, N14995, N13903, N1196);
and AND4 (N18456, N18447, N8555, N1424, N15840);
and AND4 (N18457, N18449, N10846, N10977, N8703);
xor XOR2 (N18458, N18456, N15441);
and AND3 (N18459, N18453, N13323, N5357);
nand NAND4 (N18460, N18454, N18242, N3325, N6329);
buf BUF1 (N18461, N18443);
not NOT1 (N18462, N18452);
and AND3 (N18463, N18461, N8946, N14785);
and AND2 (N18464, N18437, N12260);
not NOT1 (N18465, N18432);
nand NAND3 (N18466, N18462, N13537, N6019);
nor NOR2 (N18467, N18465, N3634);
buf BUF1 (N18468, N18457);
and AND4 (N18469, N18460, N16209, N13614, N8181);
or OR3 (N18470, N18466, N452, N4413);
and AND2 (N18471, N18468, N3197);
xor XOR2 (N18472, N18463, N191);
nor NOR3 (N18473, N18459, N2295, N8548);
nor NOR3 (N18474, N18464, N7398, N1219);
and AND2 (N18475, N18469, N13051);
buf BUF1 (N18476, N18475);
and AND2 (N18477, N18470, N15443);
nand NAND4 (N18478, N18476, N15199, N3348, N4752);
buf BUF1 (N18479, N18471);
nand NAND4 (N18480, N18473, N18184, N8293, N637);
not NOT1 (N18481, N18472);
xor XOR2 (N18482, N18480, N3295);
or OR3 (N18483, N18448, N8391, N12434);
or OR4 (N18484, N18482, N13560, N2638, N18363);
xor XOR2 (N18485, N18478, N5721);
nor NOR3 (N18486, N18455, N13922, N16738);
not NOT1 (N18487, N18484);
not NOT1 (N18488, N18479);
nand NAND4 (N18489, N18481, N1891, N16301, N9741);
or OR2 (N18490, N18489, N8893);
buf BUF1 (N18491, N18486);
xor XOR2 (N18492, N18477, N3178);
not NOT1 (N18493, N18490);
buf BUF1 (N18494, N18485);
xor XOR2 (N18495, N18467, N17080);
buf BUF1 (N18496, N18483);
nand NAND3 (N18497, N18496, N9442, N10404);
or OR2 (N18498, N18487, N1456);
not NOT1 (N18499, N18492);
nor NOR2 (N18500, N18499, N14613);
xor XOR2 (N18501, N18474, N14451);
and AND3 (N18502, N18494, N17279, N14598);
or OR4 (N18503, N18495, N12500, N18478, N14090);
xor XOR2 (N18504, N18491, N14969);
or OR3 (N18505, N18503, N14271, N12732);
xor XOR2 (N18506, N18497, N2740);
buf BUF1 (N18507, N18501);
not NOT1 (N18508, N18507);
not NOT1 (N18509, N18504);
xor XOR2 (N18510, N18509, N6068);
or OR4 (N18511, N18502, N3676, N5526, N1552);
not NOT1 (N18512, N18510);
xor XOR2 (N18513, N18458, N8468);
not NOT1 (N18514, N18506);
nor NOR3 (N18515, N18498, N2385, N18127);
and AND2 (N18516, N18500, N7493);
nand NAND4 (N18517, N18515, N17459, N12245, N13445);
nor NOR2 (N18518, N18511, N11495);
xor XOR2 (N18519, N18493, N310);
nor NOR2 (N18520, N18519, N1663);
not NOT1 (N18521, N18514);
and AND4 (N18522, N18520, N11045, N1681, N8991);
and AND4 (N18523, N18517, N8231, N6244, N5672);
xor XOR2 (N18524, N18488, N14437);
and AND2 (N18525, N18505, N1186);
and AND2 (N18526, N18521, N15911);
xor XOR2 (N18527, N18518, N17013);
and AND3 (N18528, N18508, N8178, N2765);
xor XOR2 (N18529, N18524, N6518);
not NOT1 (N18530, N18512);
nand NAND2 (N18531, N18523, N12457);
nand NAND4 (N18532, N18530, N6481, N7579, N14165);
nand NAND3 (N18533, N18513, N9796, N10163);
buf BUF1 (N18534, N18532);
and AND3 (N18535, N18529, N2674, N2159);
not NOT1 (N18536, N18527);
nor NOR2 (N18537, N18525, N17373);
nor NOR2 (N18538, N18536, N2783);
buf BUF1 (N18539, N18538);
buf BUF1 (N18540, N18531);
buf BUF1 (N18541, N18533);
nor NOR4 (N18542, N18526, N13558, N16016, N8076);
nor NOR4 (N18543, N18528, N5913, N927, N12274);
nor NOR4 (N18544, N18541, N4869, N10596, N6600);
xor XOR2 (N18545, N18522, N7961);
xor XOR2 (N18546, N18543, N2341);
nor NOR3 (N18547, N18544, N17615, N4005);
buf BUF1 (N18548, N18535);
buf BUF1 (N18549, N18547);
and AND3 (N18550, N18537, N14402, N4852);
nand NAND3 (N18551, N18550, N7215, N12843);
nor NOR3 (N18552, N18534, N10920, N7747);
nor NOR3 (N18553, N18549, N1411, N1494);
nor NOR3 (N18554, N18542, N14876, N14944);
nor NOR2 (N18555, N18539, N17017);
nor NOR4 (N18556, N18540, N16957, N14205, N7894);
nor NOR3 (N18557, N18553, N3257, N17486);
and AND3 (N18558, N18554, N16140, N16718);
and AND2 (N18559, N18558, N15378);
or OR2 (N18560, N18556, N10215);
nand NAND2 (N18561, N18555, N11927);
nand NAND2 (N18562, N18552, N2015);
or OR4 (N18563, N18561, N9613, N13627, N9097);
xor XOR2 (N18564, N18545, N1573);
xor XOR2 (N18565, N18551, N17659);
nor NOR3 (N18566, N18563, N7265, N16003);
nor NOR4 (N18567, N18557, N18309, N10571, N1417);
nand NAND2 (N18568, N18566, N7097);
buf BUF1 (N18569, N18559);
nand NAND2 (N18570, N18568, N14538);
nor NOR3 (N18571, N18516, N18301, N5037);
nand NAND2 (N18572, N18548, N12027);
xor XOR2 (N18573, N18571, N4566);
nand NAND3 (N18574, N18546, N583, N18002);
nor NOR2 (N18575, N18570, N9955);
not NOT1 (N18576, N18575);
not NOT1 (N18577, N18573);
buf BUF1 (N18578, N18562);
and AND2 (N18579, N18576, N5849);
not NOT1 (N18580, N18578);
and AND3 (N18581, N18564, N7130, N7293);
not NOT1 (N18582, N18565);
nor NOR2 (N18583, N18580, N18072);
buf BUF1 (N18584, N18560);
xor XOR2 (N18585, N18572, N15030);
xor XOR2 (N18586, N18581, N15254);
not NOT1 (N18587, N18586);
and AND4 (N18588, N18569, N10956, N5702, N9178);
and AND3 (N18589, N18577, N13555, N17158);
and AND3 (N18590, N18589, N7432, N7609);
not NOT1 (N18591, N18582);
xor XOR2 (N18592, N18574, N5003);
nand NAND3 (N18593, N18567, N3410, N16737);
not NOT1 (N18594, N18584);
or OR3 (N18595, N18587, N8495, N5238);
or OR3 (N18596, N18583, N1815, N1672);
nand NAND2 (N18597, N18595, N1866);
nor NOR4 (N18598, N18585, N1786, N462, N3582);
or OR4 (N18599, N18593, N1064, N3103, N693);
or OR4 (N18600, N18594, N16815, N9374, N5371);
or OR3 (N18601, N18590, N2849, N6333);
buf BUF1 (N18602, N18601);
or OR3 (N18603, N18600, N17347, N11379);
and AND3 (N18604, N18597, N9230, N5334);
not NOT1 (N18605, N18602);
or OR3 (N18606, N18579, N4303, N378);
and AND2 (N18607, N18598, N7981);
not NOT1 (N18608, N18591);
or OR3 (N18609, N18606, N2101, N1732);
buf BUF1 (N18610, N18596);
and AND2 (N18611, N18605, N14103);
or OR3 (N18612, N18603, N3338, N12025);
buf BUF1 (N18613, N18607);
xor XOR2 (N18614, N18609, N8275);
buf BUF1 (N18615, N18611);
buf BUF1 (N18616, N18599);
or OR3 (N18617, N18614, N17372, N11695);
nand NAND3 (N18618, N18608, N4894, N10670);
and AND2 (N18619, N18618, N3505);
xor XOR2 (N18620, N18617, N10469);
buf BUF1 (N18621, N18610);
nand NAND3 (N18622, N18613, N3664, N17407);
nor NOR3 (N18623, N18615, N7249, N3489);
xor XOR2 (N18624, N18592, N2298);
buf BUF1 (N18625, N18621);
and AND2 (N18626, N18588, N5467);
buf BUF1 (N18627, N18625);
nor NOR2 (N18628, N18622, N5041);
buf BUF1 (N18629, N18624);
not NOT1 (N18630, N18626);
nor NOR3 (N18631, N18628, N4675, N11070);
nand NAND2 (N18632, N18604, N17174);
buf BUF1 (N18633, N18631);
xor XOR2 (N18634, N18632, N5280);
nor NOR4 (N18635, N18629, N2287, N6224, N9811);
not NOT1 (N18636, N18627);
or OR4 (N18637, N18619, N12503, N14344, N11586);
and AND2 (N18638, N18630, N285);
or OR4 (N18639, N18620, N4308, N12734, N5760);
nor NOR2 (N18640, N18638, N9263);
nand NAND3 (N18641, N18635, N15886, N12407);
buf BUF1 (N18642, N18612);
and AND4 (N18643, N18642, N8956, N1864, N11749);
and AND4 (N18644, N18639, N4813, N7496, N13714);
nor NOR3 (N18645, N18644, N16894, N16091);
nor NOR2 (N18646, N18645, N6914);
and AND2 (N18647, N18641, N13788);
buf BUF1 (N18648, N18643);
nor NOR4 (N18649, N18634, N925, N10743, N6618);
and AND3 (N18650, N18636, N4771, N6219);
xor XOR2 (N18651, N18623, N18089);
or OR3 (N18652, N18637, N4260, N18391);
not NOT1 (N18653, N18652);
xor XOR2 (N18654, N18651, N16093);
or OR4 (N18655, N18649, N13619, N8059, N4586);
and AND3 (N18656, N18654, N16113, N3724);
nand NAND3 (N18657, N18653, N6913, N10706);
and AND4 (N18658, N18646, N13688, N14332, N12201);
xor XOR2 (N18659, N18657, N13294);
xor XOR2 (N18660, N18616, N3813);
not NOT1 (N18661, N18658);
or OR2 (N18662, N18661, N18539);
not NOT1 (N18663, N18648);
and AND2 (N18664, N18662, N18433);
nand NAND3 (N18665, N18660, N10906, N12642);
not NOT1 (N18666, N18664);
nor NOR2 (N18667, N18656, N6015);
buf BUF1 (N18668, N18663);
nand NAND2 (N18669, N18659, N11054);
nor NOR2 (N18670, N18669, N15613);
not NOT1 (N18671, N18668);
not NOT1 (N18672, N18665);
xor XOR2 (N18673, N18672, N2924);
or OR4 (N18674, N18647, N10004, N12065, N11792);
or OR4 (N18675, N18671, N1394, N7824, N16881);
or OR2 (N18676, N18655, N1357);
buf BUF1 (N18677, N18666);
buf BUF1 (N18678, N18650);
not NOT1 (N18679, N18633);
nand NAND2 (N18680, N18676, N12689);
or OR4 (N18681, N18667, N8246, N11652, N18654);
buf BUF1 (N18682, N18679);
nor NOR4 (N18683, N18674, N15680, N3278, N550);
or OR3 (N18684, N18675, N7543, N11678);
xor XOR2 (N18685, N18677, N9853);
not NOT1 (N18686, N18684);
and AND4 (N18687, N18686, N1345, N14368, N3400);
nand NAND3 (N18688, N18673, N12531, N11173);
and AND2 (N18689, N18670, N9329);
and AND3 (N18690, N18689, N18009, N12835);
or OR4 (N18691, N18685, N10928, N9726, N9099);
buf BUF1 (N18692, N18678);
nand NAND2 (N18693, N18688, N887);
nand NAND2 (N18694, N18682, N16008);
buf BUF1 (N18695, N18681);
buf BUF1 (N18696, N18690);
not NOT1 (N18697, N18696);
and AND2 (N18698, N18691, N18370);
not NOT1 (N18699, N18695);
nand NAND3 (N18700, N18687, N14839, N5300);
buf BUF1 (N18701, N18640);
xor XOR2 (N18702, N18701, N463);
nand NAND2 (N18703, N18698, N5471);
not NOT1 (N18704, N18694);
not NOT1 (N18705, N18693);
xor XOR2 (N18706, N18705, N5399);
buf BUF1 (N18707, N18699);
or OR3 (N18708, N18707, N13910, N946);
nand NAND2 (N18709, N18697, N16757);
and AND3 (N18710, N18704, N12238, N1406);
nand NAND4 (N18711, N18683, N12105, N8735, N15777);
nor NOR3 (N18712, N18709, N8283, N3546);
nor NOR3 (N18713, N18680, N1011, N12402);
and AND2 (N18714, N18706, N10734);
not NOT1 (N18715, N18712);
nand NAND4 (N18716, N18711, N8446, N2270, N3539);
buf BUF1 (N18717, N18702);
nand NAND3 (N18718, N18708, N6478, N11236);
and AND2 (N18719, N18692, N12525);
buf BUF1 (N18720, N18714);
or OR4 (N18721, N18718, N12824, N4422, N17570);
not NOT1 (N18722, N18717);
not NOT1 (N18723, N18715);
nor NOR3 (N18724, N18720, N1113, N16504);
not NOT1 (N18725, N18716);
not NOT1 (N18726, N18723);
xor XOR2 (N18727, N18722, N292);
not NOT1 (N18728, N18726);
and AND3 (N18729, N18703, N13964, N14696);
or OR3 (N18730, N18729, N15928, N4648);
or OR2 (N18731, N18730, N16779);
nor NOR2 (N18732, N18727, N8295);
nor NOR2 (N18733, N18728, N7381);
xor XOR2 (N18734, N18719, N6237);
and AND3 (N18735, N18710, N267, N14463);
and AND3 (N18736, N18735, N3214, N2272);
and AND2 (N18737, N18725, N3963);
and AND3 (N18738, N18737, N9411, N18310);
xor XOR2 (N18739, N18732, N16834);
and AND2 (N18740, N18736, N17325);
nand NAND2 (N18741, N18721, N14209);
and AND4 (N18742, N18713, N18497, N12969, N5491);
and AND2 (N18743, N18733, N9592);
or OR3 (N18744, N18700, N14577, N3544);
not NOT1 (N18745, N18740);
buf BUF1 (N18746, N18738);
nand NAND3 (N18747, N18742, N9594, N5703);
buf BUF1 (N18748, N18724);
or OR3 (N18749, N18731, N17444, N10483);
nand NAND4 (N18750, N18734, N6086, N2148, N12153);
or OR3 (N18751, N18743, N17968, N11745);
or OR4 (N18752, N18747, N14669, N9082, N3851);
or OR4 (N18753, N18739, N16760, N14313, N6514);
or OR3 (N18754, N18752, N3606, N8650);
and AND2 (N18755, N18745, N4290);
not NOT1 (N18756, N18744);
not NOT1 (N18757, N18748);
not NOT1 (N18758, N18754);
and AND2 (N18759, N18746, N13100);
buf BUF1 (N18760, N18753);
or OR3 (N18761, N18758, N9596, N4854);
xor XOR2 (N18762, N18761, N18652);
xor XOR2 (N18763, N18760, N444);
nand NAND2 (N18764, N18741, N11613);
buf BUF1 (N18765, N18763);
or OR3 (N18766, N18762, N1215, N376);
nand NAND3 (N18767, N18750, N10320, N13484);
or OR2 (N18768, N18749, N3607);
or OR2 (N18769, N18765, N15467);
nor NOR4 (N18770, N18751, N3019, N17873, N2653);
not NOT1 (N18771, N18768);
nor NOR2 (N18772, N18766, N15101);
nand NAND3 (N18773, N18755, N7267, N18635);
buf BUF1 (N18774, N18756);
nand NAND2 (N18775, N18769, N12468);
or OR4 (N18776, N18775, N1693, N14745, N10355);
nand NAND2 (N18777, N18774, N11589);
nand NAND4 (N18778, N18767, N3988, N17995, N4833);
nor NOR3 (N18779, N18776, N12618, N6542);
or OR3 (N18780, N18764, N573, N4440);
xor XOR2 (N18781, N18759, N13877);
nand NAND2 (N18782, N18773, N1086);
and AND2 (N18783, N18771, N155);
not NOT1 (N18784, N18782);
nand NAND2 (N18785, N18778, N17191);
xor XOR2 (N18786, N18779, N16844);
xor XOR2 (N18787, N18772, N6515);
not NOT1 (N18788, N18780);
and AND4 (N18789, N18781, N8947, N7120, N7922);
nand NAND3 (N18790, N18786, N6539, N11698);
not NOT1 (N18791, N18770);
and AND3 (N18792, N18789, N8095, N6853);
nor NOR3 (N18793, N18757, N11106, N6903);
not NOT1 (N18794, N18788);
buf BUF1 (N18795, N18785);
xor XOR2 (N18796, N18777, N4748);
nor NOR3 (N18797, N18792, N16443, N10993);
and AND2 (N18798, N18790, N11663);
and AND4 (N18799, N18791, N8094, N18268, N4829);
nand NAND2 (N18800, N18796, N9886);
xor XOR2 (N18801, N18787, N11100);
and AND3 (N18802, N18801, N14950, N12834);
not NOT1 (N18803, N18795);
not NOT1 (N18804, N18783);
and AND4 (N18805, N18784, N7652, N5959, N16285);
not NOT1 (N18806, N18799);
xor XOR2 (N18807, N18805, N16173);
nand NAND3 (N18808, N18806, N11158, N5311);
or OR3 (N18809, N18807, N740, N13019);
or OR4 (N18810, N18804, N16240, N745, N7390);
or OR3 (N18811, N18803, N4582, N311);
or OR3 (N18812, N18802, N14345, N3903);
not NOT1 (N18813, N18794);
or OR4 (N18814, N18810, N8354, N9834, N10552);
xor XOR2 (N18815, N18808, N1579);
xor XOR2 (N18816, N18797, N13424);
nor NOR4 (N18817, N18814, N12536, N1775, N1538);
nor NOR2 (N18818, N18812, N14582);
or OR2 (N18819, N18809, N6219);
nor NOR4 (N18820, N18800, N17290, N18029, N14843);
nor NOR4 (N18821, N18820, N10806, N5075, N17546);
and AND4 (N18822, N18816, N6872, N5021, N4753);
xor XOR2 (N18823, N18815, N9793);
buf BUF1 (N18824, N18813);
and AND4 (N18825, N18818, N14507, N13211, N13522);
and AND2 (N18826, N18819, N14103);
nand NAND2 (N18827, N18824, N7169);
xor XOR2 (N18828, N18823, N15622);
buf BUF1 (N18829, N18822);
and AND2 (N18830, N18829, N10593);
buf BUF1 (N18831, N18827);
buf BUF1 (N18832, N18811);
and AND2 (N18833, N18830, N7971);
not NOT1 (N18834, N18826);
or OR2 (N18835, N18825, N8360);
nor NOR2 (N18836, N18831, N8373);
and AND4 (N18837, N18832, N9745, N18589, N16248);
buf BUF1 (N18838, N18837);
nand NAND4 (N18839, N18838, N14571, N16219, N17541);
xor XOR2 (N18840, N18835, N12796);
not NOT1 (N18841, N18839);
or OR2 (N18842, N18798, N7796);
nor NOR4 (N18843, N18840, N14188, N15602, N17051);
nand NAND2 (N18844, N18842, N7503);
not NOT1 (N18845, N18843);
xor XOR2 (N18846, N18821, N1290);
not NOT1 (N18847, N18793);
or OR4 (N18848, N18841, N18763, N8564, N14426);
nand NAND3 (N18849, N18828, N15760, N5699);
nor NOR3 (N18850, N18834, N16011, N13117);
and AND4 (N18851, N18848, N1101, N7471, N17672);
nor NOR3 (N18852, N18833, N16260, N3614);
not NOT1 (N18853, N18836);
buf BUF1 (N18854, N18851);
nand NAND3 (N18855, N18817, N8414, N3213);
and AND3 (N18856, N18845, N3414, N10752);
not NOT1 (N18857, N18846);
and AND3 (N18858, N18855, N5640, N7542);
nor NOR3 (N18859, N18856, N12424, N16793);
xor XOR2 (N18860, N18852, N15033);
buf BUF1 (N18861, N18849);
nand NAND3 (N18862, N18854, N11139, N878);
nand NAND4 (N18863, N18860, N18147, N13773, N16522);
xor XOR2 (N18864, N18850, N5259);
not NOT1 (N18865, N18857);
and AND2 (N18866, N18861, N241);
nor NOR2 (N18867, N18863, N8);
or OR3 (N18868, N18867, N1259, N10342);
nand NAND3 (N18869, N18866, N10377, N4808);
buf BUF1 (N18870, N18853);
not NOT1 (N18871, N18865);
nand NAND3 (N18872, N18868, N3712, N9738);
not NOT1 (N18873, N18847);
nor NOR4 (N18874, N18871, N6668, N3618, N4008);
xor XOR2 (N18875, N18872, N18834);
xor XOR2 (N18876, N18858, N17128);
xor XOR2 (N18877, N18870, N1211);
and AND2 (N18878, N18876, N15109);
not NOT1 (N18879, N18862);
nand NAND4 (N18880, N18875, N7576, N9086, N7768);
or OR4 (N18881, N18869, N17156, N3989, N7331);
not NOT1 (N18882, N18880);
nand NAND3 (N18883, N18881, N9384, N12527);
xor XOR2 (N18884, N18859, N8252);
or OR2 (N18885, N18884, N8048);
xor XOR2 (N18886, N18864, N14937);
nand NAND3 (N18887, N18878, N5170, N15841);
xor XOR2 (N18888, N18879, N11010);
or OR3 (N18889, N18883, N11543, N6454);
nor NOR3 (N18890, N18887, N5055, N5157);
and AND3 (N18891, N18882, N16951, N12726);
not NOT1 (N18892, N18844);
nor NOR4 (N18893, N18885, N14850, N18510, N15658);
buf BUF1 (N18894, N18892);
nor NOR2 (N18895, N18886, N10188);
buf BUF1 (N18896, N18891);
buf BUF1 (N18897, N18890);
buf BUF1 (N18898, N18895);
nor NOR2 (N18899, N18894, N14488);
and AND2 (N18900, N18889, N18851);
and AND2 (N18901, N18896, N16324);
or OR2 (N18902, N18888, N7187);
buf BUF1 (N18903, N18901);
buf BUF1 (N18904, N18874);
buf BUF1 (N18905, N18873);
not NOT1 (N18906, N18899);
and AND2 (N18907, N18893, N17440);
xor XOR2 (N18908, N18906, N5417);
nor NOR2 (N18909, N18907, N10062);
and AND2 (N18910, N18897, N9640);
not NOT1 (N18911, N18904);
nor NOR2 (N18912, N18877, N3756);
and AND4 (N18913, N18912, N6691, N1777, N18411);
or OR2 (N18914, N18905, N10658);
buf BUF1 (N18915, N18898);
and AND2 (N18916, N18911, N15817);
nand NAND3 (N18917, N18902, N4812, N13978);
and AND4 (N18918, N18903, N4607, N7184, N15344);
buf BUF1 (N18919, N18916);
and AND2 (N18920, N18913, N7110);
and AND3 (N18921, N18908, N12569, N11942);
buf BUF1 (N18922, N18909);
buf BUF1 (N18923, N18914);
not NOT1 (N18924, N18920);
nor NOR2 (N18925, N18919, N16449);
buf BUF1 (N18926, N18923);
buf BUF1 (N18927, N18918);
buf BUF1 (N18928, N18917);
xor XOR2 (N18929, N18928, N18429);
nand NAND4 (N18930, N18900, N7203, N15389, N8628);
xor XOR2 (N18931, N18929, N16652);
nand NAND4 (N18932, N18926, N3631, N8575, N7376);
or OR4 (N18933, N18927, N6759, N4516, N11876);
not NOT1 (N18934, N18933);
nor NOR4 (N18935, N18934, N3211, N15348, N2226);
not NOT1 (N18936, N18924);
and AND2 (N18937, N18931, N10049);
and AND3 (N18938, N18930, N652, N15813);
nor NOR2 (N18939, N18915, N13337);
nor NOR4 (N18940, N18921, N17353, N850, N9856);
not NOT1 (N18941, N18925);
not NOT1 (N18942, N18910);
nand NAND4 (N18943, N18937, N6033, N11932, N1260);
nor NOR3 (N18944, N18922, N255, N3525);
buf BUF1 (N18945, N18940);
buf BUF1 (N18946, N18944);
buf BUF1 (N18947, N18942);
xor XOR2 (N18948, N18943, N6535);
nand NAND3 (N18949, N18948, N4512, N1894);
nor NOR4 (N18950, N18945, N16121, N15576, N12189);
xor XOR2 (N18951, N18947, N6134);
buf BUF1 (N18952, N18932);
and AND4 (N18953, N18950, N2555, N11681, N14578);
and AND2 (N18954, N18936, N14634);
xor XOR2 (N18955, N18946, N10486);
buf BUF1 (N18956, N18939);
buf BUF1 (N18957, N18935);
nor NOR3 (N18958, N18952, N4218, N14077);
or OR4 (N18959, N18957, N9815, N16780, N1973);
buf BUF1 (N18960, N18956);
buf BUF1 (N18961, N18941);
and AND2 (N18962, N18951, N9130);
or OR4 (N18963, N18958, N5466, N9075, N13960);
nor NOR4 (N18964, N18963, N6463, N5252, N17644);
buf BUF1 (N18965, N18938);
not NOT1 (N18966, N18965);
or OR3 (N18967, N18953, N6780, N10149);
xor XOR2 (N18968, N18949, N11759);
and AND3 (N18969, N18964, N9898, N15030);
nand NAND3 (N18970, N18954, N16210, N9808);
and AND4 (N18971, N18955, N3486, N9683, N18372);
nor NOR3 (N18972, N18961, N8349, N4249);
and AND3 (N18973, N18967, N7953, N10563);
nand NAND2 (N18974, N18962, N5807);
buf BUF1 (N18975, N18970);
buf BUF1 (N18976, N18975);
and AND2 (N18977, N18972, N8336);
or OR3 (N18978, N18966, N8908, N5877);
or OR4 (N18979, N18978, N8429, N2322, N8684);
and AND3 (N18980, N18979, N16820, N3910);
and AND2 (N18981, N18980, N9336);
nand NAND4 (N18982, N18971, N13913, N1099, N15257);
and AND4 (N18983, N18976, N5778, N13040, N14695);
not NOT1 (N18984, N18977);
xor XOR2 (N18985, N18973, N12049);
nor NOR2 (N18986, N18960, N12965);
not NOT1 (N18987, N18984);
buf BUF1 (N18988, N18959);
nor NOR4 (N18989, N18981, N6284, N6788, N7196);
buf BUF1 (N18990, N18974);
xor XOR2 (N18991, N18990, N13435);
buf BUF1 (N18992, N18991);
buf BUF1 (N18993, N18988);
not NOT1 (N18994, N18992);
and AND3 (N18995, N18982, N13835, N5823);
nor NOR2 (N18996, N18989, N9903);
and AND4 (N18997, N18969, N16038, N18556, N6901);
not NOT1 (N18998, N18997);
or OR2 (N18999, N18987, N14687);
buf BUF1 (N19000, N18968);
not NOT1 (N19001, N18995);
xor XOR2 (N19002, N18986, N12675);
not NOT1 (N19003, N18999);
nor NOR3 (N19004, N18983, N18091, N8297);
nand NAND2 (N19005, N18994, N9342);
xor XOR2 (N19006, N19001, N10425);
or OR3 (N19007, N19000, N7469, N5984);
or OR2 (N19008, N19005, N12905);
buf BUF1 (N19009, N19002);
nand NAND3 (N19010, N19008, N8744, N15784);
xor XOR2 (N19011, N18996, N5280);
nand NAND3 (N19012, N19009, N6180, N2524);
xor XOR2 (N19013, N18993, N12521);
nor NOR4 (N19014, N19003, N16316, N8857, N13195);
nand NAND4 (N19015, N19004, N1126, N10480, N18042);
xor XOR2 (N19016, N19010, N15229);
or OR4 (N19017, N19012, N17844, N14253, N18008);
and AND3 (N19018, N18985, N9011, N11940);
not NOT1 (N19019, N19007);
and AND2 (N19020, N19015, N14617);
not NOT1 (N19021, N19006);
xor XOR2 (N19022, N19016, N16489);
and AND2 (N19023, N19013, N1464);
not NOT1 (N19024, N19017);
and AND4 (N19025, N19014, N9231, N4334, N3899);
buf BUF1 (N19026, N19024);
or OR3 (N19027, N19018, N14030, N6725);
nor NOR4 (N19028, N19027, N17846, N6721, N9043);
or OR2 (N19029, N19021, N3503);
or OR4 (N19030, N19028, N2770, N15869, N11562);
and AND2 (N19031, N18998, N11515);
or OR4 (N19032, N19011, N15767, N13746, N615);
nor NOR2 (N19033, N19025, N3272);
xor XOR2 (N19034, N19031, N8469);
or OR4 (N19035, N19019, N1498, N18773, N17609);
buf BUF1 (N19036, N19034);
nor NOR3 (N19037, N19023, N17184, N2896);
buf BUF1 (N19038, N19036);
or OR4 (N19039, N19022, N9441, N9903, N8698);
buf BUF1 (N19040, N19037);
and AND2 (N19041, N19035, N8617);
not NOT1 (N19042, N19026);
xor XOR2 (N19043, N19029, N9396);
buf BUF1 (N19044, N19041);
buf BUF1 (N19045, N19032);
nor NOR2 (N19046, N19033, N14682);
buf BUF1 (N19047, N19042);
nor NOR4 (N19048, N19020, N8649, N15158, N1101);
nor NOR2 (N19049, N19030, N3107);
and AND3 (N19050, N19049, N5103, N3032);
xor XOR2 (N19051, N19048, N15592);
or OR2 (N19052, N19051, N18225);
and AND3 (N19053, N19050, N2689, N2045);
xor XOR2 (N19054, N19045, N15421);
xor XOR2 (N19055, N19047, N9196);
or OR4 (N19056, N19039, N16426, N17933, N16540);
and AND4 (N19057, N19056, N16880, N14206, N11000);
not NOT1 (N19058, N19053);
nand NAND2 (N19059, N19052, N12815);
or OR4 (N19060, N19057, N2838, N6230, N6148);
or OR2 (N19061, N19055, N4896);
and AND4 (N19062, N19038, N1674, N12100, N4835);
not NOT1 (N19063, N19059);
not NOT1 (N19064, N19054);
or OR2 (N19065, N19040, N16733);
xor XOR2 (N19066, N19046, N53);
or OR2 (N19067, N19065, N11947);
nand NAND4 (N19068, N19060, N11170, N13753, N18261);
and AND3 (N19069, N19064, N1628, N5650);
xor XOR2 (N19070, N19066, N15136);
and AND3 (N19071, N19070, N4041, N17770);
or OR4 (N19072, N19058, N9714, N17542, N3797);
or OR4 (N19073, N19072, N15578, N10841, N12505);
nand NAND4 (N19074, N19069, N7919, N5425, N11403);
nand NAND2 (N19075, N19073, N10665);
or OR2 (N19076, N19043, N9340);
nor NOR3 (N19077, N19062, N5960, N10395);
not NOT1 (N19078, N19068);
xor XOR2 (N19079, N19074, N1818);
not NOT1 (N19080, N19079);
not NOT1 (N19081, N19078);
buf BUF1 (N19082, N19080);
nor NOR4 (N19083, N19067, N7227, N1761, N11161);
xor XOR2 (N19084, N19082, N15401);
nand NAND2 (N19085, N19061, N16421);
buf BUF1 (N19086, N19071);
not NOT1 (N19087, N19076);
nand NAND2 (N19088, N19083, N10372);
and AND4 (N19089, N19077, N16453, N140, N15311);
and AND3 (N19090, N19081, N2288, N17348);
not NOT1 (N19091, N19090);
not NOT1 (N19092, N19089);
buf BUF1 (N19093, N19088);
and AND2 (N19094, N19075, N18184);
buf BUF1 (N19095, N19086);
not NOT1 (N19096, N19044);
and AND4 (N19097, N19093, N8738, N14100, N2572);
xor XOR2 (N19098, N19091, N7797);
and AND3 (N19099, N19098, N6578, N9871);
nor NOR3 (N19100, N19087, N19077, N11295);
and AND3 (N19101, N19096, N5197, N11019);
not NOT1 (N19102, N19085);
and AND4 (N19103, N19063, N1661, N11471, N14040);
buf BUF1 (N19104, N19101);
nand NAND2 (N19105, N19103, N6820);
not NOT1 (N19106, N19104);
nand NAND4 (N19107, N19099, N1352, N15064, N18034);
nor NOR3 (N19108, N19100, N1607, N17791);
xor XOR2 (N19109, N19105, N365);
nor NOR2 (N19110, N19107, N5388);
nand NAND2 (N19111, N19084, N525);
buf BUF1 (N19112, N19092);
and AND3 (N19113, N19111, N14637, N18429);
xor XOR2 (N19114, N19095, N9126);
buf BUF1 (N19115, N19110);
xor XOR2 (N19116, N19108, N14175);
not NOT1 (N19117, N19116);
xor XOR2 (N19118, N19097, N12649);
xor XOR2 (N19119, N19109, N11871);
nor NOR2 (N19120, N19119, N943);
and AND4 (N19121, N19114, N3330, N13381, N3435);
or OR3 (N19122, N19112, N1834, N3880);
nand NAND4 (N19123, N19122, N154, N17730, N2560);
buf BUF1 (N19124, N19106);
nand NAND3 (N19125, N19113, N11847, N13116);
nor NOR4 (N19126, N19118, N7363, N7079, N6049);
or OR3 (N19127, N19123, N2900, N2070);
nand NAND3 (N19128, N19117, N18054, N13568);
and AND3 (N19129, N19125, N7577, N17809);
xor XOR2 (N19130, N19094, N6711);
nand NAND3 (N19131, N19121, N666, N13268);
nor NOR4 (N19132, N19127, N12107, N12154, N17572);
and AND2 (N19133, N19129, N15520);
nor NOR4 (N19134, N19124, N14604, N18667, N12742);
buf BUF1 (N19135, N19126);
xor XOR2 (N19136, N19135, N6181);
not NOT1 (N19137, N19120);
xor XOR2 (N19138, N19136, N3927);
or OR2 (N19139, N19115, N3145);
nand NAND4 (N19140, N19132, N12214, N1053, N17803);
not NOT1 (N19141, N19131);
xor XOR2 (N19142, N19141, N99);
nand NAND4 (N19143, N19102, N7817, N1221, N9429);
buf BUF1 (N19144, N19139);
not NOT1 (N19145, N19128);
nand NAND3 (N19146, N19134, N8461, N15712);
nand NAND4 (N19147, N19137, N17857, N11493, N902);
not NOT1 (N19148, N19147);
and AND2 (N19149, N19145, N6021);
buf BUF1 (N19150, N19143);
buf BUF1 (N19151, N19148);
xor XOR2 (N19152, N19140, N7249);
xor XOR2 (N19153, N19152, N10672);
not NOT1 (N19154, N19146);
or OR3 (N19155, N19151, N12367, N5562);
buf BUF1 (N19156, N19138);
nor NOR4 (N19157, N19156, N7907, N11566, N17930);
and AND4 (N19158, N19144, N8176, N466, N12961);
buf BUF1 (N19159, N19157);
xor XOR2 (N19160, N19133, N15781);
nand NAND4 (N19161, N19158, N13784, N15941, N14575);
buf BUF1 (N19162, N19130);
and AND3 (N19163, N19161, N12185, N8512);
and AND2 (N19164, N19142, N572);
not NOT1 (N19165, N19154);
nand NAND4 (N19166, N19155, N6381, N3233, N312);
nor NOR3 (N19167, N19163, N11695, N13745);
and AND2 (N19168, N19166, N8105);
xor XOR2 (N19169, N19153, N2361);
or OR3 (N19170, N19168, N5248, N15399);
xor XOR2 (N19171, N19160, N15226);
nand NAND2 (N19172, N19165, N11180);
and AND3 (N19173, N19167, N5324, N15378);
nor NOR3 (N19174, N19171, N4694, N15832);
nor NOR3 (N19175, N19173, N15298, N17001);
xor XOR2 (N19176, N19150, N13040);
not NOT1 (N19177, N19162);
xor XOR2 (N19178, N19164, N11151);
nand NAND2 (N19179, N19174, N5194);
or OR4 (N19180, N19159, N5139, N8278, N11672);
buf BUF1 (N19181, N19175);
not NOT1 (N19182, N19181);
xor XOR2 (N19183, N19178, N1941);
nor NOR4 (N19184, N19170, N5079, N10313, N16728);
or OR2 (N19185, N19149, N13718);
and AND3 (N19186, N19177, N2591, N17004);
xor XOR2 (N19187, N19172, N14978);
or OR3 (N19188, N19179, N9328, N7632);
not NOT1 (N19189, N19183);
xor XOR2 (N19190, N19186, N1761);
not NOT1 (N19191, N19169);
nor NOR3 (N19192, N19190, N5267, N12826);
or OR3 (N19193, N19180, N10120, N1432);
buf BUF1 (N19194, N19185);
buf BUF1 (N19195, N19187);
nor NOR3 (N19196, N19176, N13297, N6706);
not NOT1 (N19197, N19192);
nor NOR4 (N19198, N19197, N7641, N231, N12572);
nand NAND2 (N19199, N19194, N14042);
or OR4 (N19200, N19193, N15725, N11843, N7433);
and AND3 (N19201, N19189, N7889, N1803);
nand NAND3 (N19202, N19198, N3396, N18824);
nand NAND4 (N19203, N19196, N7361, N7024, N2357);
nor NOR3 (N19204, N19188, N18880, N17962);
buf BUF1 (N19205, N19202);
nand NAND3 (N19206, N19205, N6931, N6001);
not NOT1 (N19207, N19184);
buf BUF1 (N19208, N19206);
and AND2 (N19209, N19195, N6612);
nor NOR4 (N19210, N19203, N4355, N16175, N6404);
buf BUF1 (N19211, N19207);
nand NAND4 (N19212, N19210, N4188, N8409, N17988);
xor XOR2 (N19213, N19199, N11070);
nor NOR2 (N19214, N19201, N17268);
nor NOR4 (N19215, N19209, N6028, N4424, N5721);
not NOT1 (N19216, N19214);
nand NAND4 (N19217, N19204, N13578, N4988, N11887);
or OR4 (N19218, N19208, N2696, N9200, N3749);
nor NOR3 (N19219, N19218, N17262, N797);
buf BUF1 (N19220, N19212);
buf BUF1 (N19221, N19217);
buf BUF1 (N19222, N19220);
buf BUF1 (N19223, N19211);
or OR4 (N19224, N19223, N11879, N2988, N16402);
xor XOR2 (N19225, N19224, N16349);
xor XOR2 (N19226, N19225, N14102);
buf BUF1 (N19227, N19226);
buf BUF1 (N19228, N19182);
not NOT1 (N19229, N19213);
and AND3 (N19230, N19215, N16315, N14391);
or OR2 (N19231, N19221, N5204);
xor XOR2 (N19232, N19227, N3808);
or OR4 (N19233, N19216, N19129, N1881, N12331);
nor NOR3 (N19234, N19229, N5639, N2572);
or OR2 (N19235, N19228, N4692);
nand NAND2 (N19236, N19233, N350);
nor NOR2 (N19237, N19234, N17463);
nor NOR2 (N19238, N19235, N15675);
nand NAND4 (N19239, N19230, N3470, N9677, N16291);
not NOT1 (N19240, N19200);
buf BUF1 (N19241, N19236);
buf BUF1 (N19242, N19238);
nand NAND4 (N19243, N19240, N16110, N296, N12769);
buf BUF1 (N19244, N19243);
and AND2 (N19245, N19231, N11510);
not NOT1 (N19246, N19232);
buf BUF1 (N19247, N19222);
xor XOR2 (N19248, N19219, N4919);
nand NAND3 (N19249, N19247, N16746, N14936);
buf BUF1 (N19250, N19239);
and AND2 (N19251, N19241, N6053);
nand NAND2 (N19252, N19244, N14384);
and AND3 (N19253, N19191, N15340, N3945);
or OR3 (N19254, N19253, N16559, N11100);
buf BUF1 (N19255, N19254);
not NOT1 (N19256, N19255);
buf BUF1 (N19257, N19256);
and AND4 (N19258, N19250, N1269, N13156, N1458);
nor NOR4 (N19259, N19258, N13160, N6448, N13197);
xor XOR2 (N19260, N19252, N18149);
nand NAND4 (N19261, N19246, N4428, N1276, N14757);
buf BUF1 (N19262, N19260);
nand NAND3 (N19263, N19237, N4575, N6871);
and AND3 (N19264, N19259, N11046, N13848);
buf BUF1 (N19265, N19245);
nand NAND3 (N19266, N19264, N14039, N14246);
nand NAND3 (N19267, N19261, N3647, N8795);
nand NAND3 (N19268, N19266, N18685, N4218);
nand NAND3 (N19269, N19263, N12602, N1284);
nand NAND4 (N19270, N19268, N3711, N17757, N2997);
not NOT1 (N19271, N19269);
or OR2 (N19272, N19257, N9217);
buf BUF1 (N19273, N19248);
nor NOR3 (N19274, N19251, N2579, N8699);
nand NAND3 (N19275, N19272, N10407, N12995);
buf BUF1 (N19276, N19267);
buf BUF1 (N19277, N19273);
nand NAND4 (N19278, N19275, N4533, N1740, N14766);
or OR4 (N19279, N19242, N14895, N5701, N17303);
nand NAND2 (N19280, N19262, N246);
xor XOR2 (N19281, N19277, N3101);
not NOT1 (N19282, N19271);
xor XOR2 (N19283, N19280, N4656);
or OR2 (N19284, N19279, N433);
or OR2 (N19285, N19283, N202);
and AND4 (N19286, N19285, N7697, N5670, N11508);
or OR4 (N19287, N19270, N4455, N17592, N17830);
nand NAND3 (N19288, N19286, N2058, N935);
not NOT1 (N19289, N19281);
or OR2 (N19290, N19276, N11028);
nand NAND4 (N19291, N19287, N4417, N7715, N7798);
nand NAND4 (N19292, N19284, N13624, N13191, N728);
and AND3 (N19293, N19274, N9192, N7927);
nor NOR4 (N19294, N19265, N14468, N16069, N14786);
nand NAND4 (N19295, N19290, N12571, N8537, N16016);
xor XOR2 (N19296, N19289, N12396);
or OR3 (N19297, N19292, N2749, N14041);
buf BUF1 (N19298, N19278);
buf BUF1 (N19299, N19297);
and AND3 (N19300, N19293, N10707, N7934);
not NOT1 (N19301, N19296);
not NOT1 (N19302, N19298);
and AND4 (N19303, N19300, N14737, N8192, N2438);
buf BUF1 (N19304, N19303);
nand NAND4 (N19305, N19299, N10309, N6930, N6809);
xor XOR2 (N19306, N19295, N11690);
nand NAND3 (N19307, N19302, N11227, N16475);
or OR3 (N19308, N19304, N4213, N8220);
xor XOR2 (N19309, N19282, N12349);
or OR2 (N19310, N19306, N5947);
xor XOR2 (N19311, N19308, N3578);
xor XOR2 (N19312, N19309, N15155);
xor XOR2 (N19313, N19291, N15272);
nand NAND3 (N19314, N19312, N2946, N9862);
or OR2 (N19315, N19313, N13042);
buf BUF1 (N19316, N19310);
nor NOR4 (N19317, N19288, N7792, N15712, N2389);
and AND4 (N19318, N19315, N9904, N18812, N12076);
not NOT1 (N19319, N19316);
nand NAND4 (N19320, N19318, N18911, N7283, N4296);
buf BUF1 (N19321, N19311);
xor XOR2 (N19322, N19294, N5480);
not NOT1 (N19323, N19320);
not NOT1 (N19324, N19321);
or OR2 (N19325, N19249, N11789);
or OR4 (N19326, N19314, N10852, N15493, N893);
xor XOR2 (N19327, N19322, N16251);
or OR4 (N19328, N19307, N14868, N2238, N4076);
nand NAND4 (N19329, N19328, N18908, N13080, N7183);
and AND2 (N19330, N19317, N16368);
xor XOR2 (N19331, N19324, N9846);
or OR3 (N19332, N19331, N4941, N7059);
xor XOR2 (N19333, N19325, N12058);
and AND2 (N19334, N19332, N17456);
or OR3 (N19335, N19329, N4521, N16948);
buf BUF1 (N19336, N19301);
and AND3 (N19337, N19330, N357, N7208);
xor XOR2 (N19338, N19336, N5258);
or OR3 (N19339, N19334, N14412, N8790);
not NOT1 (N19340, N19335);
and AND4 (N19341, N19333, N17658, N8952, N16296);
buf BUF1 (N19342, N19339);
or OR4 (N19343, N19323, N13370, N6437, N12991);
xor XOR2 (N19344, N19327, N3478);
xor XOR2 (N19345, N19340, N5731);
not NOT1 (N19346, N19338);
and AND2 (N19347, N19346, N8474);
nor NOR3 (N19348, N19319, N2816, N12918);
nand NAND4 (N19349, N19344, N1383, N16680, N15188);
xor XOR2 (N19350, N19349, N9269);
xor XOR2 (N19351, N19343, N13507);
or OR2 (N19352, N19348, N16353);
nand NAND2 (N19353, N19347, N5852);
or OR3 (N19354, N19337, N7710, N12405);
not NOT1 (N19355, N19354);
nand NAND2 (N19356, N19355, N15923);
and AND4 (N19357, N19326, N13985, N15507, N12630);
buf BUF1 (N19358, N19350);
or OR4 (N19359, N19342, N11261, N15483, N18569);
not NOT1 (N19360, N19341);
not NOT1 (N19361, N19358);
nand NAND2 (N19362, N19351, N1626);
nor NOR2 (N19363, N19356, N3024);
or OR3 (N19364, N19357, N12994, N17547);
and AND3 (N19365, N19352, N7008, N10471);
buf BUF1 (N19366, N19362);
or OR2 (N19367, N19359, N4654);
xor XOR2 (N19368, N19353, N19185);
nand NAND2 (N19369, N19360, N19352);
nand NAND4 (N19370, N19305, N10979, N14130, N1693);
buf BUF1 (N19371, N19363);
nand NAND3 (N19372, N19345, N7890, N9076);
or OR3 (N19373, N19364, N17384, N4947);
or OR4 (N19374, N19367, N4721, N18919, N16634);
xor XOR2 (N19375, N19361, N12950);
buf BUF1 (N19376, N19375);
buf BUF1 (N19377, N19372);
nor NOR3 (N19378, N19366, N5141, N13000);
not NOT1 (N19379, N19370);
nor NOR4 (N19380, N19377, N12766, N3518, N17455);
xor XOR2 (N19381, N19365, N13383);
and AND2 (N19382, N19369, N7723);
and AND3 (N19383, N19374, N9565, N3829);
not NOT1 (N19384, N19381);
xor XOR2 (N19385, N19384, N11075);
or OR2 (N19386, N19379, N12391);
nor NOR4 (N19387, N19383, N6934, N18649, N4195);
not NOT1 (N19388, N19382);
nor NOR2 (N19389, N19380, N12728);
and AND2 (N19390, N19385, N8371);
buf BUF1 (N19391, N19387);
or OR4 (N19392, N19391, N8884, N14325, N2004);
xor XOR2 (N19393, N19376, N11455);
and AND3 (N19394, N19392, N7436, N3467);
or OR3 (N19395, N19390, N9856, N1221);
nand NAND2 (N19396, N19373, N382);
buf BUF1 (N19397, N19378);
or OR3 (N19398, N19395, N16492, N11799);
xor XOR2 (N19399, N19371, N10399);
or OR3 (N19400, N19386, N9058, N6272);
or OR2 (N19401, N19368, N8002);
or OR4 (N19402, N19393, N5026, N13295, N11135);
xor XOR2 (N19403, N19402, N987);
xor XOR2 (N19404, N19399, N17250);
not NOT1 (N19405, N19398);
nor NOR3 (N19406, N19405, N9637, N9401);
xor XOR2 (N19407, N19394, N8388);
nor NOR4 (N19408, N19396, N10866, N16499, N13027);
and AND2 (N19409, N19403, N4269);
buf BUF1 (N19410, N19388);
nand NAND2 (N19411, N19397, N2664);
nand NAND2 (N19412, N19409, N2173);
not NOT1 (N19413, N19404);
nor NOR4 (N19414, N19400, N18135, N15525, N6712);
nand NAND2 (N19415, N19413, N7074);
and AND4 (N19416, N19401, N7005, N16558, N14430);
xor XOR2 (N19417, N19412, N14582);
xor XOR2 (N19418, N19414, N3902);
or OR2 (N19419, N19416, N16317);
xor XOR2 (N19420, N19389, N2537);
nand NAND4 (N19421, N19417, N6245, N15661, N9599);
buf BUF1 (N19422, N19418);
nor NOR3 (N19423, N19408, N8871, N14394);
and AND4 (N19424, N19420, N9972, N11730, N13033);
not NOT1 (N19425, N19419);
nand NAND2 (N19426, N19410, N185);
nand NAND2 (N19427, N19425, N3573);
nor NOR3 (N19428, N19422, N17645, N18862);
nor NOR4 (N19429, N19424, N9451, N15051, N13852);
not NOT1 (N19430, N19411);
or OR2 (N19431, N19423, N10046);
nand NAND3 (N19432, N19430, N6422, N9430);
or OR4 (N19433, N19407, N15022, N14663, N1516);
or OR3 (N19434, N19432, N10855, N16534);
xor XOR2 (N19435, N19406, N17192);
or OR4 (N19436, N19431, N564, N15579, N17727);
or OR2 (N19437, N19421, N16172);
xor XOR2 (N19438, N19435, N8378);
and AND3 (N19439, N19438, N15210, N6599);
xor XOR2 (N19440, N19428, N143);
and AND3 (N19441, N19437, N11751, N10006);
nor NOR3 (N19442, N19436, N1999, N18647);
buf BUF1 (N19443, N19429);
nand NAND3 (N19444, N19439, N2424, N14670);
nand NAND4 (N19445, N19426, N2488, N15508, N2286);
nand NAND3 (N19446, N19442, N3094, N6975);
xor XOR2 (N19447, N19440, N7025);
or OR4 (N19448, N19445, N17847, N5962, N12505);
nor NOR2 (N19449, N19446, N4412);
or OR2 (N19450, N19433, N5807);
nor NOR2 (N19451, N19443, N1188);
not NOT1 (N19452, N19450);
nand NAND3 (N19453, N19452, N5723, N132);
or OR3 (N19454, N19451, N2207, N200);
xor XOR2 (N19455, N19448, N13967);
and AND3 (N19456, N19427, N15648, N12949);
buf BUF1 (N19457, N19434);
buf BUF1 (N19458, N19454);
or OR4 (N19459, N19444, N11939, N17402, N12676);
xor XOR2 (N19460, N19457, N2023);
and AND3 (N19461, N19447, N14687, N18258);
nand NAND3 (N19462, N19459, N12845, N3234);
not NOT1 (N19463, N19453);
buf BUF1 (N19464, N19456);
xor XOR2 (N19465, N19458, N9585);
xor XOR2 (N19466, N19462, N16664);
not NOT1 (N19467, N19464);
xor XOR2 (N19468, N19466, N14245);
or OR3 (N19469, N19455, N15544, N16353);
and AND2 (N19470, N19460, N16164);
nand NAND2 (N19471, N19465, N3369);
nand NAND2 (N19472, N19470, N2264);
nor NOR4 (N19473, N19469, N7251, N9172, N14335);
and AND2 (N19474, N19415, N13873);
nor NOR3 (N19475, N19449, N10037, N10340);
not NOT1 (N19476, N19461);
xor XOR2 (N19477, N19468, N3022);
or OR4 (N19478, N19475, N18890, N15692, N3189);
nor NOR3 (N19479, N19471, N8162, N6783);
not NOT1 (N19480, N19473);
and AND4 (N19481, N19463, N17789, N13398, N2744);
nor NOR2 (N19482, N19481, N19356);
nand NAND2 (N19483, N19482, N3947);
nand NAND4 (N19484, N19467, N7768, N6621, N6943);
or OR3 (N19485, N19476, N116, N12723);
buf BUF1 (N19486, N19480);
xor XOR2 (N19487, N19441, N1055);
not NOT1 (N19488, N19484);
nand NAND2 (N19489, N19477, N7182);
nor NOR2 (N19490, N19486, N10404);
or OR4 (N19491, N19488, N12142, N11979, N14542);
buf BUF1 (N19492, N19479);
xor XOR2 (N19493, N19490, N11118);
or OR4 (N19494, N19487, N6999, N9573, N16012);
xor XOR2 (N19495, N19491, N8998);
nor NOR2 (N19496, N19494, N742);
not NOT1 (N19497, N19478);
and AND4 (N19498, N19492, N5829, N11797, N9552);
xor XOR2 (N19499, N19485, N9836);
nand NAND2 (N19500, N19483, N15433);
buf BUF1 (N19501, N19496);
nor NOR2 (N19502, N19472, N6033);
buf BUF1 (N19503, N19489);
buf BUF1 (N19504, N19495);
buf BUF1 (N19505, N19504);
nor NOR4 (N19506, N19474, N7418, N18443, N19354);
or OR2 (N19507, N19503, N2964);
nand NAND3 (N19508, N19506, N466, N1364);
buf BUF1 (N19509, N19497);
xor XOR2 (N19510, N19505, N10566);
nor NOR2 (N19511, N19498, N10050);
nor NOR2 (N19512, N19508, N11193);
nor NOR3 (N19513, N19499, N6524, N16157);
buf BUF1 (N19514, N19507);
buf BUF1 (N19515, N19510);
nand NAND3 (N19516, N19513, N16781, N15469);
nor NOR2 (N19517, N19516, N3716);
not NOT1 (N19518, N19514);
nand NAND2 (N19519, N19500, N16410);
and AND4 (N19520, N19501, N2379, N1604, N13144);
and AND3 (N19521, N19502, N3328, N13949);
nand NAND3 (N19522, N19517, N4405, N11297);
and AND2 (N19523, N19509, N10624);
buf BUF1 (N19524, N19521);
xor XOR2 (N19525, N19518, N13574);
buf BUF1 (N19526, N19523);
or OR2 (N19527, N19525, N17936);
and AND4 (N19528, N19519, N11475, N18533, N4770);
nor NOR3 (N19529, N19527, N4574, N15175);
or OR4 (N19530, N19512, N6020, N13413, N747);
buf BUF1 (N19531, N19526);
xor XOR2 (N19532, N19529, N8195);
buf BUF1 (N19533, N19522);
and AND3 (N19534, N19524, N7092, N5289);
and AND3 (N19535, N19528, N1927, N15895);
and AND4 (N19536, N19530, N13617, N11953, N4199);
xor XOR2 (N19537, N19511, N2371);
nand NAND4 (N19538, N19533, N4378, N7737, N1172);
buf BUF1 (N19539, N19520);
buf BUF1 (N19540, N19535);
and AND3 (N19541, N19540, N5971, N1136);
not NOT1 (N19542, N19541);
or OR4 (N19543, N19539, N2365, N3402, N10423);
buf BUF1 (N19544, N19493);
nand NAND2 (N19545, N19531, N18987);
buf BUF1 (N19546, N19536);
nor NOR3 (N19547, N19534, N15297, N7925);
or OR2 (N19548, N19545, N4081);
not NOT1 (N19549, N19542);
xor XOR2 (N19550, N19515, N18493);
nor NOR3 (N19551, N19538, N4914, N4797);
and AND4 (N19552, N19547, N9218, N16601, N13121);
not NOT1 (N19553, N19551);
xor XOR2 (N19554, N19532, N8441);
xor XOR2 (N19555, N19549, N12439);
and AND2 (N19556, N19544, N17877);
and AND4 (N19557, N19555, N13694, N8797, N13874);
nand NAND4 (N19558, N19553, N9444, N499, N18929);
buf BUF1 (N19559, N19543);
nand NAND4 (N19560, N19550, N15843, N5513, N2120);
and AND3 (N19561, N19537, N15727, N2622);
buf BUF1 (N19562, N19559);
nor NOR2 (N19563, N19554, N13931);
nor NOR2 (N19564, N19561, N9484);
and AND2 (N19565, N19563, N18604);
and AND3 (N19566, N19565, N9266, N14904);
nand NAND2 (N19567, N19558, N16783);
and AND4 (N19568, N19564, N8865, N5411, N8026);
not NOT1 (N19569, N19566);
nor NOR3 (N19570, N19556, N13664, N3893);
nand NAND2 (N19571, N19552, N4791);
or OR3 (N19572, N19569, N2420, N7154);
not NOT1 (N19573, N19548);
nand NAND3 (N19574, N19573, N321, N14196);
nand NAND4 (N19575, N19570, N19151, N6896, N1371);
or OR2 (N19576, N19560, N16429);
buf BUF1 (N19577, N19576);
and AND4 (N19578, N19562, N4329, N3290, N18249);
or OR4 (N19579, N19568, N9655, N2351, N7679);
nor NOR2 (N19580, N19546, N17655);
buf BUF1 (N19581, N19579);
not NOT1 (N19582, N19578);
not NOT1 (N19583, N19574);
nor NOR3 (N19584, N19575, N18728, N2065);
buf BUF1 (N19585, N19581);
and AND4 (N19586, N19567, N8870, N15569, N4229);
buf BUF1 (N19587, N19577);
xor XOR2 (N19588, N19583, N4776);
nor NOR4 (N19589, N19585, N11984, N12264, N5303);
nor NOR3 (N19590, N19584, N9353, N10953);
xor XOR2 (N19591, N19571, N5116);
and AND4 (N19592, N19588, N4415, N13179, N13478);
or OR4 (N19593, N19587, N17831, N5082, N12324);
xor XOR2 (N19594, N19593, N12476);
and AND2 (N19595, N19591, N4975);
nand NAND4 (N19596, N19580, N9534, N7713, N10536);
and AND3 (N19597, N19594, N15418, N12285);
nand NAND2 (N19598, N19582, N10687);
buf BUF1 (N19599, N19572);
buf BUF1 (N19600, N19597);
not NOT1 (N19601, N19586);
xor XOR2 (N19602, N19600, N6858);
nor NOR2 (N19603, N19589, N9265);
nor NOR3 (N19604, N19599, N4497, N16279);
nand NAND4 (N19605, N19596, N17938, N4313, N719);
buf BUF1 (N19606, N19557);
xor XOR2 (N19607, N19606, N17724);
nor NOR4 (N19608, N19590, N52, N15108, N6516);
nand NAND3 (N19609, N19595, N8739, N9906);
not NOT1 (N19610, N19592);
or OR4 (N19611, N19605, N994, N2898, N13880);
nand NAND3 (N19612, N19610, N13457, N12883);
xor XOR2 (N19613, N19602, N285);
xor XOR2 (N19614, N19603, N16253);
xor XOR2 (N19615, N19612, N6655);
and AND3 (N19616, N19607, N4251, N18560);
nor NOR4 (N19617, N19604, N19453, N14652, N3276);
and AND3 (N19618, N19598, N4621, N13201);
buf BUF1 (N19619, N19615);
nand NAND2 (N19620, N19608, N19492);
and AND2 (N19621, N19611, N6158);
not NOT1 (N19622, N19601);
and AND2 (N19623, N19614, N15696);
buf BUF1 (N19624, N19617);
and AND4 (N19625, N19620, N10469, N12910, N14371);
and AND3 (N19626, N19609, N4103, N5612);
nand NAND2 (N19627, N19619, N209);
nor NOR3 (N19628, N19618, N15939, N4412);
buf BUF1 (N19629, N19621);
nand NAND2 (N19630, N19616, N733);
nand NAND3 (N19631, N19628, N16355, N6230);
or OR4 (N19632, N19623, N13072, N3491, N2508);
xor XOR2 (N19633, N19625, N4569);
and AND3 (N19634, N19627, N19161, N19344);
not NOT1 (N19635, N19634);
and AND4 (N19636, N19622, N9379, N6901, N15842);
xor XOR2 (N19637, N19635, N2358);
not NOT1 (N19638, N19629);
not NOT1 (N19639, N19637);
nor NOR3 (N19640, N19624, N1164, N7286);
or OR3 (N19641, N19638, N14564, N11577);
and AND2 (N19642, N19636, N2488);
not NOT1 (N19643, N19631);
buf BUF1 (N19644, N19640);
and AND4 (N19645, N19613, N10993, N8246, N2153);
and AND2 (N19646, N19642, N12841);
nand NAND3 (N19647, N19633, N1533, N2995);
or OR2 (N19648, N19645, N3825);
or OR3 (N19649, N19644, N12335, N2831);
buf BUF1 (N19650, N19641);
or OR2 (N19651, N19639, N11616);
nand NAND4 (N19652, N19643, N1975, N8206, N822);
xor XOR2 (N19653, N19648, N2548);
nand NAND4 (N19654, N19653, N15004, N15697, N12617);
xor XOR2 (N19655, N19630, N17702);
not NOT1 (N19656, N19652);
xor XOR2 (N19657, N19650, N18315);
nor NOR2 (N19658, N19654, N7374);
and AND3 (N19659, N19656, N5477, N4321);
nor NOR2 (N19660, N19659, N763);
or OR4 (N19661, N19655, N7987, N16314, N15322);
nor NOR2 (N19662, N19657, N5985);
not NOT1 (N19663, N19662);
or OR3 (N19664, N19646, N6229, N15715);
xor XOR2 (N19665, N19658, N17464);
or OR4 (N19666, N19651, N12335, N14779, N11618);
and AND3 (N19667, N19665, N13973, N9884);
and AND4 (N19668, N19666, N17756, N8995, N2163);
and AND4 (N19669, N19649, N17458, N1986, N228);
buf BUF1 (N19670, N19632);
nor NOR4 (N19671, N19660, N11608, N10597, N2586);
and AND2 (N19672, N19664, N13660);
buf BUF1 (N19673, N19670);
buf BUF1 (N19674, N19668);
nand NAND4 (N19675, N19674, N16518, N12710, N6574);
nor NOR4 (N19676, N19675, N63, N667, N342);
nand NAND4 (N19677, N19672, N7103, N17277, N16221);
nand NAND3 (N19678, N19676, N9244, N3007);
nor NOR2 (N19679, N19663, N7057);
buf BUF1 (N19680, N19626);
nand NAND2 (N19681, N19677, N15591);
xor XOR2 (N19682, N19681, N9389);
xor XOR2 (N19683, N19671, N13855);
buf BUF1 (N19684, N19680);
buf BUF1 (N19685, N19673);
nand NAND2 (N19686, N19683, N8542);
nor NOR4 (N19687, N19684, N10478, N12700, N10469);
or OR3 (N19688, N19687, N9029, N16648);
xor XOR2 (N19689, N19678, N7897);
not NOT1 (N19690, N19682);
nor NOR2 (N19691, N19685, N11947);
nor NOR3 (N19692, N19690, N12766, N15691);
xor XOR2 (N19693, N19669, N6233);
not NOT1 (N19694, N19689);
xor XOR2 (N19695, N19686, N5389);
nand NAND3 (N19696, N19692, N17215, N7203);
not NOT1 (N19697, N19694);
not NOT1 (N19698, N19667);
nor NOR3 (N19699, N19693, N14528, N19180);
xor XOR2 (N19700, N19661, N17821);
buf BUF1 (N19701, N19697);
nand NAND2 (N19702, N19700, N5218);
xor XOR2 (N19703, N19688, N9594);
xor XOR2 (N19704, N19696, N9394);
nor NOR4 (N19705, N19702, N3839, N10476, N3740);
and AND2 (N19706, N19703, N15095);
xor XOR2 (N19707, N19704, N2);
not NOT1 (N19708, N19679);
nand NAND3 (N19709, N19691, N3937, N11088);
nand NAND4 (N19710, N19647, N15740, N2298, N130);
nand NAND3 (N19711, N19710, N10010, N8024);
not NOT1 (N19712, N19699);
or OR4 (N19713, N19709, N10740, N9068, N6836);
not NOT1 (N19714, N19705);
nand NAND2 (N19715, N19712, N15895);
not NOT1 (N19716, N19713);
buf BUF1 (N19717, N19708);
nand NAND4 (N19718, N19698, N11393, N6871, N7896);
not NOT1 (N19719, N19717);
or OR3 (N19720, N19711, N17710, N16118);
xor XOR2 (N19721, N19701, N2074);
nand NAND4 (N19722, N19715, N1322, N9230, N17515);
or OR2 (N19723, N19706, N57);
buf BUF1 (N19724, N19718);
or OR2 (N19725, N19695, N10986);
or OR4 (N19726, N19723, N3733, N3640, N11087);
nand NAND4 (N19727, N19716, N10322, N9093, N7704);
not NOT1 (N19728, N19727);
not NOT1 (N19729, N19726);
nand NAND3 (N19730, N19724, N17489, N16227);
buf BUF1 (N19731, N19714);
xor XOR2 (N19732, N19729, N18096);
not NOT1 (N19733, N19720);
xor XOR2 (N19734, N19722, N2200);
nand NAND3 (N19735, N19731, N15332, N11015);
not NOT1 (N19736, N19728);
xor XOR2 (N19737, N19736, N2385);
nand NAND3 (N19738, N19733, N2711, N13737);
buf BUF1 (N19739, N19735);
or OR2 (N19740, N19738, N1040);
nor NOR3 (N19741, N19734, N5350, N449);
nor NOR4 (N19742, N19739, N16528, N17376, N13593);
buf BUF1 (N19743, N19737);
and AND3 (N19744, N19719, N695, N8900);
or OR4 (N19745, N19741, N15881, N15412, N1954);
not NOT1 (N19746, N19707);
and AND3 (N19747, N19746, N19622, N9165);
xor XOR2 (N19748, N19725, N11547);
nand NAND4 (N19749, N19744, N2124, N3375, N2158);
or OR2 (N19750, N19748, N11568);
nand NAND4 (N19751, N19745, N9615, N6191, N10585);
not NOT1 (N19752, N19751);
or OR4 (N19753, N19732, N7566, N3938, N267);
or OR3 (N19754, N19752, N9629, N7598);
and AND4 (N19755, N19740, N14047, N14566, N1617);
not NOT1 (N19756, N19747);
xor XOR2 (N19757, N19750, N2759);
nor NOR4 (N19758, N19721, N3944, N12726, N2164);
buf BUF1 (N19759, N19754);
xor XOR2 (N19760, N19742, N2998);
or OR3 (N19761, N19757, N14232, N3135);
xor XOR2 (N19762, N19749, N8980);
buf BUF1 (N19763, N19753);
xor XOR2 (N19764, N19759, N4193);
nor NOR2 (N19765, N19762, N15306);
and AND2 (N19766, N19765, N15097);
nand NAND3 (N19767, N19763, N7790, N1060);
nand NAND4 (N19768, N19761, N18469, N12819, N12189);
nor NOR2 (N19769, N19764, N9504);
nor NOR3 (N19770, N19730, N17685, N8913);
nand NAND2 (N19771, N19767, N5971);
and AND2 (N19772, N19769, N3305);
xor XOR2 (N19773, N19758, N19062);
xor XOR2 (N19774, N19755, N18826);
and AND4 (N19775, N19756, N14363, N1292, N18063);
xor XOR2 (N19776, N19771, N13058);
nand NAND2 (N19777, N19773, N8200);
not NOT1 (N19778, N19774);
buf BUF1 (N19779, N19743);
or OR4 (N19780, N19770, N1151, N13213, N12887);
not NOT1 (N19781, N19760);
xor XOR2 (N19782, N19778, N5101);
xor XOR2 (N19783, N19775, N13609);
and AND3 (N19784, N19779, N18246, N108);
nor NOR4 (N19785, N19768, N4146, N11172, N15889);
nor NOR3 (N19786, N19784, N16280, N10196);
or OR4 (N19787, N19782, N616, N7626, N8887);
and AND4 (N19788, N19786, N3115, N3649, N18409);
xor XOR2 (N19789, N19783, N2937);
or OR2 (N19790, N19781, N12634);
nor NOR2 (N19791, N19780, N7522);
buf BUF1 (N19792, N19766);
nand NAND2 (N19793, N19785, N9917);
nand NAND2 (N19794, N19787, N11453);
buf BUF1 (N19795, N19777);
nand NAND3 (N19796, N19788, N1963, N17150);
not NOT1 (N19797, N19792);
or OR3 (N19798, N19797, N13120, N9780);
xor XOR2 (N19799, N19772, N819);
xor XOR2 (N19800, N19799, N16813);
nor NOR2 (N19801, N19798, N3634);
nand NAND4 (N19802, N19801, N17893, N5704, N1609);
not NOT1 (N19803, N19790);
or OR3 (N19804, N19802, N10373, N6028);
nand NAND4 (N19805, N19800, N946, N5610, N16433);
not NOT1 (N19806, N19791);
or OR3 (N19807, N19804, N17366, N10030);
not NOT1 (N19808, N19794);
xor XOR2 (N19809, N19807, N2053);
nor NOR2 (N19810, N19808, N14798);
and AND3 (N19811, N19793, N7107, N957);
nor NOR2 (N19812, N19776, N12553);
not NOT1 (N19813, N19809);
xor XOR2 (N19814, N19812, N10052);
xor XOR2 (N19815, N19805, N12079);
not NOT1 (N19816, N19813);
and AND4 (N19817, N19816, N7645, N17351, N19533);
buf BUF1 (N19818, N19795);
xor XOR2 (N19819, N19803, N15805);
and AND3 (N19820, N19789, N18948, N19495);
and AND4 (N19821, N19815, N8763, N14153, N6489);
nand NAND4 (N19822, N19818, N5584, N10483, N11948);
nor NOR3 (N19823, N19810, N1006, N14071);
or OR3 (N19824, N19823, N14531, N12656);
buf BUF1 (N19825, N19806);
nand NAND3 (N19826, N19819, N9060, N8524);
buf BUF1 (N19827, N19825);
buf BUF1 (N19828, N19820);
buf BUF1 (N19829, N19817);
nand NAND3 (N19830, N19829, N13138, N7210);
and AND4 (N19831, N19828, N4829, N5821, N19012);
nor NOR4 (N19832, N19830, N17098, N519, N434);
or OR2 (N19833, N19814, N4206);
xor XOR2 (N19834, N19811, N7804);
xor XOR2 (N19835, N19821, N17572);
not NOT1 (N19836, N19834);
nand NAND2 (N19837, N19831, N11765);
and AND2 (N19838, N19837, N5384);
nand NAND4 (N19839, N19838, N7084, N8190, N1084);
nand NAND2 (N19840, N19835, N6920);
xor XOR2 (N19841, N19796, N5312);
and AND4 (N19842, N19836, N4081, N13127, N16341);
nor NOR3 (N19843, N19826, N6304, N18916);
and AND2 (N19844, N19841, N6982);
xor XOR2 (N19845, N19842, N8714);
buf BUF1 (N19846, N19845);
buf BUF1 (N19847, N19824);
nor NOR4 (N19848, N19846, N7743, N19395, N8267);
not NOT1 (N19849, N19844);
not NOT1 (N19850, N19843);
or OR2 (N19851, N19850, N4644);
and AND3 (N19852, N19822, N4373, N11776);
buf BUF1 (N19853, N19849);
xor XOR2 (N19854, N19839, N6139);
not NOT1 (N19855, N19853);
and AND3 (N19856, N19827, N15978, N12812);
nand NAND2 (N19857, N19854, N5071);
or OR2 (N19858, N19857, N433);
nor NOR2 (N19859, N19833, N14976);
or OR2 (N19860, N19851, N6869);
xor XOR2 (N19861, N19840, N6624);
and AND4 (N19862, N19855, N17918, N9899, N17048);
and AND2 (N19863, N19859, N828);
not NOT1 (N19864, N19832);
nand NAND3 (N19865, N19861, N7730, N19030);
xor XOR2 (N19866, N19864, N10582);
xor XOR2 (N19867, N19858, N15540);
not NOT1 (N19868, N19848);
not NOT1 (N19869, N19847);
xor XOR2 (N19870, N19856, N12435);
and AND2 (N19871, N19852, N17836);
not NOT1 (N19872, N19869);
nand NAND2 (N19873, N19872, N3486);
buf BUF1 (N19874, N19860);
nand NAND2 (N19875, N19867, N13847);
nand NAND2 (N19876, N19874, N12261);
nand NAND3 (N19877, N19868, N9003, N15681);
and AND3 (N19878, N19871, N14088, N8698);
nand NAND4 (N19879, N19877, N18695, N1421, N14226);
and AND4 (N19880, N19879, N6170, N3155, N5003);
nand NAND4 (N19881, N19866, N11837, N9293, N18390);
not NOT1 (N19882, N19862);
nor NOR2 (N19883, N19873, N4397);
nor NOR3 (N19884, N19881, N8132, N9630);
not NOT1 (N19885, N19870);
and AND2 (N19886, N19880, N12888);
nor NOR4 (N19887, N19883, N13083, N17773, N6797);
not NOT1 (N19888, N19875);
or OR4 (N19889, N19878, N641, N10484, N14637);
and AND2 (N19890, N19882, N11592);
nor NOR3 (N19891, N19865, N17841, N5693);
nand NAND3 (N19892, N19863, N13044, N18843);
buf BUF1 (N19893, N19886);
and AND2 (N19894, N19884, N1115);
and AND3 (N19895, N19888, N10819, N11690);
nor NOR3 (N19896, N19887, N10394, N11185);
and AND2 (N19897, N19894, N4132);
not NOT1 (N19898, N19892);
not NOT1 (N19899, N19893);
and AND3 (N19900, N19899, N9023, N16265);
xor XOR2 (N19901, N19885, N8134);
xor XOR2 (N19902, N19890, N16084);
buf BUF1 (N19903, N19897);
nand NAND2 (N19904, N19901, N13286);
nand NAND2 (N19905, N19898, N9176);
and AND2 (N19906, N19903, N1362);
nand NAND3 (N19907, N19904, N824, N1388);
buf BUF1 (N19908, N19906);
nor NOR2 (N19909, N19876, N4168);
or OR2 (N19910, N19889, N13519);
buf BUF1 (N19911, N19907);
not NOT1 (N19912, N19910);
buf BUF1 (N19913, N19900);
or OR2 (N19914, N19909, N11147);
or OR2 (N19915, N19905, N10948);
buf BUF1 (N19916, N19914);
xor XOR2 (N19917, N19911, N9273);
or OR3 (N19918, N19896, N6736, N10825);
buf BUF1 (N19919, N19902);
nor NOR3 (N19920, N19917, N1016, N17935);
xor XOR2 (N19921, N19915, N3471);
nor NOR2 (N19922, N19921, N17566);
or OR2 (N19923, N19922, N3551);
nand NAND2 (N19924, N19908, N4750);
buf BUF1 (N19925, N19916);
or OR3 (N19926, N19925, N870, N874);
nor NOR4 (N19927, N19919, N3437, N10414, N3879);
or OR2 (N19928, N19918, N10377);
not NOT1 (N19929, N19891);
buf BUF1 (N19930, N19920);
or OR2 (N19931, N19930, N2840);
xor XOR2 (N19932, N19895, N9383);
nor NOR3 (N19933, N19929, N6272, N1552);
xor XOR2 (N19934, N19928, N7164);
xor XOR2 (N19935, N19924, N14408);
xor XOR2 (N19936, N19926, N8020);
and AND2 (N19937, N19923, N12278);
xor XOR2 (N19938, N19936, N19620);
nand NAND2 (N19939, N19927, N14274);
and AND2 (N19940, N19939, N19098);
or OR3 (N19941, N19933, N15038, N9204);
nand NAND4 (N19942, N19938, N18537, N8714, N8103);
or OR2 (N19943, N19941, N11069);
buf BUF1 (N19944, N19940);
or OR3 (N19945, N19932, N1108, N2491);
not NOT1 (N19946, N19944);
nor NOR4 (N19947, N19931, N7768, N9740, N13148);
nand NAND3 (N19948, N19943, N3578, N13150);
or OR2 (N19949, N19946, N18349);
and AND3 (N19950, N19935, N2440, N16765);
buf BUF1 (N19951, N19945);
xor XOR2 (N19952, N19942, N16781);
not NOT1 (N19953, N19948);
nor NOR3 (N19954, N19912, N16128, N5200);
xor XOR2 (N19955, N19953, N12691);
not NOT1 (N19956, N19937);
buf BUF1 (N19957, N19955);
or OR3 (N19958, N19954, N7156, N11752);
xor XOR2 (N19959, N19951, N4378);
and AND4 (N19960, N19947, N12520, N17770, N11292);
nand NAND2 (N19961, N19956, N17941);
nor NOR4 (N19962, N19949, N10434, N19926, N12913);
buf BUF1 (N19963, N19950);
nand NAND4 (N19964, N19952, N4213, N5925, N588);
and AND2 (N19965, N19913, N19380);
nor NOR3 (N19966, N19964, N7838, N17391);
xor XOR2 (N19967, N19959, N9334);
not NOT1 (N19968, N19966);
or OR4 (N19969, N19957, N3255, N798, N3840);
not NOT1 (N19970, N19961);
or OR2 (N19971, N19958, N17745);
nand NAND2 (N19972, N19963, N3834);
or OR3 (N19973, N19965, N3645, N213);
xor XOR2 (N19974, N19973, N5017);
and AND2 (N19975, N19960, N8005);
nand NAND3 (N19976, N19971, N18650, N18998);
nor NOR3 (N19977, N19974, N5610, N14248);
and AND3 (N19978, N19969, N10567, N3342);
nand NAND4 (N19979, N19972, N7538, N341, N7964);
nor NOR4 (N19980, N19975, N4851, N13136, N17521);
buf BUF1 (N19981, N19934);
and AND3 (N19982, N19962, N4241, N18071);
and AND2 (N19983, N19968, N18428);
nand NAND4 (N19984, N19970, N9979, N13014, N16727);
xor XOR2 (N19985, N19981, N15996);
and AND3 (N19986, N19980, N6438, N9487);
and AND4 (N19987, N19983, N19245, N1576, N4912);
and AND2 (N19988, N19977, N688);
and AND2 (N19989, N19979, N8861);
nand NAND4 (N19990, N19985, N15529, N10161, N15729);
not NOT1 (N19991, N19984);
nand NAND4 (N19992, N19976, N475, N4561, N10830);
buf BUF1 (N19993, N19990);
and AND4 (N19994, N19978, N3613, N15304, N16174);
not NOT1 (N19995, N19989);
or OR4 (N19996, N19967, N12139, N13385, N8920);
not NOT1 (N19997, N19992);
nand NAND3 (N19998, N19991, N15893, N4226);
nand NAND3 (N19999, N19982, N14589, N1396);
or OR3 (N20000, N19994, N18854, N11205);
nor NOR3 (N20001, N19997, N19164, N10588);
or OR3 (N20002, N20000, N6117, N13463);
and AND2 (N20003, N19998, N2215);
nor NOR4 (N20004, N19996, N12948, N6117, N16901);
xor XOR2 (N20005, N19987, N1329);
and AND2 (N20006, N20001, N2900);
nand NAND3 (N20007, N19999, N7930, N5681);
and AND4 (N20008, N19993, N16973, N16920, N609);
and AND2 (N20009, N20003, N5343);
and AND2 (N20010, N20004, N8926);
xor XOR2 (N20011, N20009, N14601);
not NOT1 (N20012, N20011);
nand NAND3 (N20013, N20002, N7969, N1094);
buf BUF1 (N20014, N20008);
and AND3 (N20015, N19995, N15876, N5644);
nor NOR2 (N20016, N20006, N4294);
not NOT1 (N20017, N19988);
and AND4 (N20018, N20016, N2612, N16021, N13276);
nor NOR4 (N20019, N20015, N3007, N2923, N235);
and AND3 (N20020, N19986, N19267, N16129);
nor NOR2 (N20021, N20020, N4000);
not NOT1 (N20022, N20007);
buf BUF1 (N20023, N20010);
nor NOR2 (N20024, N20014, N9722);
not NOT1 (N20025, N20018);
not NOT1 (N20026, N20021);
or OR4 (N20027, N20013, N4705, N8242, N12075);
xor XOR2 (N20028, N20005, N16161);
nand NAND4 (N20029, N20026, N9026, N19328, N7001);
not NOT1 (N20030, N20023);
xor XOR2 (N20031, N20030, N1386);
not NOT1 (N20032, N20019);
not NOT1 (N20033, N20024);
xor XOR2 (N20034, N20012, N16469);
not NOT1 (N20035, N20017);
and AND2 (N20036, N20035, N9185);
not NOT1 (N20037, N20025);
or OR4 (N20038, N20022, N16313, N12679, N13456);
not NOT1 (N20039, N20031);
and AND4 (N20040, N20029, N17045, N7641, N1870);
or OR4 (N20041, N20034, N1591, N6249, N18806);
and AND4 (N20042, N20036, N3045, N18029, N6241);
and AND3 (N20043, N20039, N606, N9395);
or OR2 (N20044, N20041, N7409);
nand NAND3 (N20045, N20033, N18672, N14451);
and AND2 (N20046, N20037, N19268);
nand NAND3 (N20047, N20040, N2259, N10483);
nand NAND3 (N20048, N20038, N5647, N6350);
xor XOR2 (N20049, N20045, N3119);
nand NAND2 (N20050, N20032, N1405);
buf BUF1 (N20051, N20043);
buf BUF1 (N20052, N20049);
xor XOR2 (N20053, N20050, N5501);
buf BUF1 (N20054, N20044);
not NOT1 (N20055, N20053);
nand NAND3 (N20056, N20046, N3405, N12214);
nand NAND2 (N20057, N20047, N6864);
buf BUF1 (N20058, N20054);
nor NOR4 (N20059, N20056, N1453, N3924, N351);
xor XOR2 (N20060, N20055, N5944);
and AND4 (N20061, N20058, N11981, N230, N6285);
and AND3 (N20062, N20061, N8984, N1339);
or OR3 (N20063, N20057, N14845, N13051);
xor XOR2 (N20064, N20059, N19267);
or OR4 (N20065, N20048, N15806, N16269, N739);
or OR4 (N20066, N20064, N11918, N4111, N11060);
and AND4 (N20067, N20027, N1621, N12765, N2188);
nor NOR2 (N20068, N20028, N4471);
and AND3 (N20069, N20042, N435, N9364);
or OR4 (N20070, N20068, N13795, N6244, N3805);
or OR4 (N20071, N20069, N1540, N7115, N16127);
not NOT1 (N20072, N20066);
buf BUF1 (N20073, N20052);
nand NAND2 (N20074, N20051, N14117);
not NOT1 (N20075, N20063);
nor NOR4 (N20076, N20071, N7565, N14647, N13202);
not NOT1 (N20077, N20062);
or OR3 (N20078, N20076, N16093, N1281);
nor NOR4 (N20079, N20075, N13145, N9251, N12005);
or OR3 (N20080, N20074, N19657, N8056);
or OR4 (N20081, N20070, N7851, N17720, N6336);
not NOT1 (N20082, N20078);
or OR2 (N20083, N20065, N11047);
or OR4 (N20084, N20081, N6767, N14864, N10054);
and AND3 (N20085, N20083, N12670, N7482);
nand NAND4 (N20086, N20084, N19024, N16684, N17412);
nor NOR3 (N20087, N20082, N764, N44);
and AND4 (N20088, N20080, N5121, N160, N17802);
nand NAND4 (N20089, N20073, N15283, N9569, N4340);
xor XOR2 (N20090, N20085, N2872);
not NOT1 (N20091, N20089);
buf BUF1 (N20092, N20077);
xor XOR2 (N20093, N20086, N3365);
nor NOR3 (N20094, N20079, N11252, N5689);
buf BUF1 (N20095, N20060);
not NOT1 (N20096, N20092);
not NOT1 (N20097, N20095);
not NOT1 (N20098, N20088);
not NOT1 (N20099, N20096);
and AND3 (N20100, N20099, N16330, N1975);
or OR3 (N20101, N20087, N9848, N6922);
and AND3 (N20102, N20091, N2, N6343);
or OR4 (N20103, N20093, N16432, N3431, N8470);
nor NOR4 (N20104, N20067, N15081, N11744, N8424);
nor NOR4 (N20105, N20090, N5374, N116, N3109);
nand NAND4 (N20106, N20072, N11600, N11470, N19611);
not NOT1 (N20107, N20103);
nor NOR4 (N20108, N20105, N2688, N7557, N2197);
nand NAND2 (N20109, N20108, N8232);
not NOT1 (N20110, N20104);
nor NOR3 (N20111, N20109, N18071, N12884);
nor NOR2 (N20112, N20106, N945);
buf BUF1 (N20113, N20098);
nand NAND4 (N20114, N20100, N6720, N281, N4862);
or OR2 (N20115, N20107, N17198);
buf BUF1 (N20116, N20111);
and AND2 (N20117, N20097, N17251);
or OR4 (N20118, N20113, N2211, N4728, N19705);
not NOT1 (N20119, N20118);
buf BUF1 (N20120, N20119);
not NOT1 (N20121, N20112);
xor XOR2 (N20122, N20117, N12357);
nand NAND2 (N20123, N20121, N3552);
nor NOR2 (N20124, N20123, N3108);
nor NOR2 (N20125, N20114, N7051);
buf BUF1 (N20126, N20120);
not NOT1 (N20127, N20102);
not NOT1 (N20128, N20122);
and AND4 (N20129, N20128, N13791, N7990, N6948);
xor XOR2 (N20130, N20094, N19860);
not NOT1 (N20131, N20116);
nand NAND3 (N20132, N20130, N19293, N4701);
or OR2 (N20133, N20131, N10463);
or OR2 (N20134, N20129, N12274);
nor NOR3 (N20135, N20101, N19522, N14727);
or OR3 (N20136, N20132, N123, N16402);
nor NOR2 (N20137, N20125, N16600);
buf BUF1 (N20138, N20115);
or OR2 (N20139, N20124, N19695);
xor XOR2 (N20140, N20126, N2548);
xor XOR2 (N20141, N20133, N3705);
or OR2 (N20142, N20138, N5068);
xor XOR2 (N20143, N20135, N8237);
not NOT1 (N20144, N20141);
nor NOR4 (N20145, N20127, N10343, N12955, N9125);
xor XOR2 (N20146, N20144, N13381);
nand NAND4 (N20147, N20110, N12001, N15316, N10812);
xor XOR2 (N20148, N20140, N3397);
buf BUF1 (N20149, N20136);
xor XOR2 (N20150, N20134, N11739);
xor XOR2 (N20151, N20139, N1531);
and AND2 (N20152, N20148, N15171);
buf BUF1 (N20153, N20143);
not NOT1 (N20154, N20153);
or OR3 (N20155, N20150, N6599, N4650);
xor XOR2 (N20156, N20147, N9755);
or OR4 (N20157, N20156, N15121, N18222, N4395);
xor XOR2 (N20158, N20149, N14721);
nor NOR2 (N20159, N20155, N5303);
or OR3 (N20160, N20152, N13700, N3486);
or OR3 (N20161, N20157, N18051, N11268);
xor XOR2 (N20162, N20137, N15093);
not NOT1 (N20163, N20145);
buf BUF1 (N20164, N20151);
buf BUF1 (N20165, N20163);
or OR4 (N20166, N20160, N587, N6442, N5776);
nand NAND2 (N20167, N20165, N13872);
nand NAND4 (N20168, N20164, N14275, N7473, N16716);
or OR4 (N20169, N20146, N11745, N1188, N7081);
not NOT1 (N20170, N20154);
buf BUF1 (N20171, N20162);
xor XOR2 (N20172, N20170, N9071);
nand NAND2 (N20173, N20167, N9117);
buf BUF1 (N20174, N20159);
nand NAND4 (N20175, N20174, N7387, N6843, N19282);
nor NOR3 (N20176, N20166, N6399, N18538);
nor NOR2 (N20177, N20142, N4443);
not NOT1 (N20178, N20173);
and AND3 (N20179, N20172, N13394, N1315);
nor NOR3 (N20180, N20175, N19934, N16629);
buf BUF1 (N20181, N20171);
and AND3 (N20182, N20158, N7655, N6151);
or OR4 (N20183, N20176, N18656, N7467, N2016);
or OR2 (N20184, N20182, N1774);
not NOT1 (N20185, N20179);
xor XOR2 (N20186, N20184, N3484);
and AND4 (N20187, N20186, N12601, N16135, N7740);
nand NAND4 (N20188, N20161, N2050, N7155, N5613);
and AND2 (N20189, N20188, N1978);
buf BUF1 (N20190, N20183);
and AND2 (N20191, N20181, N9813);
or OR2 (N20192, N20185, N13150);
nor NOR2 (N20193, N20178, N12120);
or OR2 (N20194, N20191, N3804);
not NOT1 (N20195, N20180);
or OR4 (N20196, N20194, N9553, N12877, N18810);
xor XOR2 (N20197, N20193, N8466);
nor NOR4 (N20198, N20187, N9825, N182, N3080);
or OR2 (N20199, N20177, N18018);
and AND4 (N20200, N20197, N4545, N10440, N4783);
and AND2 (N20201, N20198, N11612);
and AND4 (N20202, N20192, N18837, N16900, N800);
or OR4 (N20203, N20199, N5594, N9023, N7421);
nor NOR3 (N20204, N20196, N5965, N18578);
not NOT1 (N20205, N20195);
nand NAND4 (N20206, N20168, N5673, N10989, N7671);
nor NOR2 (N20207, N20203, N17757);
or OR3 (N20208, N20200, N8333, N528);
xor XOR2 (N20209, N20205, N6774);
or OR4 (N20210, N20208, N19638, N19294, N16534);
buf BUF1 (N20211, N20209);
or OR2 (N20212, N20204, N11578);
or OR3 (N20213, N20169, N8779, N15664);
not NOT1 (N20214, N20201);
and AND2 (N20215, N20212, N13118);
nor NOR3 (N20216, N20207, N17990, N182);
nand NAND3 (N20217, N20214, N6410, N9603);
not NOT1 (N20218, N20215);
not NOT1 (N20219, N20190);
buf BUF1 (N20220, N20219);
nand NAND2 (N20221, N20202, N6337);
xor XOR2 (N20222, N20220, N7736);
not NOT1 (N20223, N20213);
or OR3 (N20224, N20223, N7143, N12350);
buf BUF1 (N20225, N20221);
nor NOR2 (N20226, N20206, N10074);
not NOT1 (N20227, N20189);
xor XOR2 (N20228, N20216, N8493);
or OR2 (N20229, N20227, N18240);
buf BUF1 (N20230, N20228);
xor XOR2 (N20231, N20230, N2490);
buf BUF1 (N20232, N20217);
nand NAND3 (N20233, N20232, N19522, N18477);
xor XOR2 (N20234, N20225, N8501);
buf BUF1 (N20235, N20234);
nand NAND3 (N20236, N20211, N19078, N19909);
or OR4 (N20237, N20235, N19471, N1237, N17962);
not NOT1 (N20238, N20236);
or OR4 (N20239, N20210, N5157, N8032, N2373);
nand NAND2 (N20240, N20238, N2016);
and AND4 (N20241, N20224, N4636, N19360, N17028);
and AND2 (N20242, N20233, N4757);
or OR2 (N20243, N20242, N17043);
and AND3 (N20244, N20239, N1689, N3645);
and AND4 (N20245, N20237, N11330, N16051, N11800);
xor XOR2 (N20246, N20229, N18366);
and AND2 (N20247, N20241, N15727);
nand NAND2 (N20248, N20240, N11895);
nor NOR2 (N20249, N20244, N17837);
or OR4 (N20250, N20247, N19031, N19445, N9591);
not NOT1 (N20251, N20248);
xor XOR2 (N20252, N20243, N593);
xor XOR2 (N20253, N20218, N18799);
nor NOR2 (N20254, N20231, N19275);
or OR4 (N20255, N20253, N441, N13697, N15466);
nor NOR2 (N20256, N20250, N7863);
nor NOR4 (N20257, N20246, N6236, N11722, N7604);
buf BUF1 (N20258, N20251);
xor XOR2 (N20259, N20256, N10703);
nand NAND2 (N20260, N20249, N7371);
buf BUF1 (N20261, N20226);
nor NOR3 (N20262, N20255, N17635, N4504);
nor NOR2 (N20263, N20259, N2767);
and AND3 (N20264, N20257, N9680, N5158);
and AND4 (N20265, N20245, N3811, N1178, N9798);
or OR3 (N20266, N20254, N5844, N10157);
not NOT1 (N20267, N20265);
and AND3 (N20268, N20222, N10378, N1611);
buf BUF1 (N20269, N20267);
nand NAND3 (N20270, N20268, N12579, N17303);
and AND3 (N20271, N20263, N3349, N11135);
xor XOR2 (N20272, N20261, N11008);
not NOT1 (N20273, N20264);
buf BUF1 (N20274, N20260);
nor NOR4 (N20275, N20270, N14858, N14114, N16605);
nand NAND4 (N20276, N20271, N3800, N15006, N18907);
xor XOR2 (N20277, N20252, N7306);
or OR3 (N20278, N20277, N7695, N1632);
buf BUF1 (N20279, N20274);
buf BUF1 (N20280, N20262);
nand NAND3 (N20281, N20273, N5019, N1214);
not NOT1 (N20282, N20272);
nor NOR4 (N20283, N20266, N5449, N13509, N9175);
nor NOR3 (N20284, N20283, N43, N2395);
nor NOR2 (N20285, N20276, N10009);
buf BUF1 (N20286, N20278);
xor XOR2 (N20287, N20279, N1064);
nor NOR3 (N20288, N20258, N18046, N16366);
xor XOR2 (N20289, N20269, N19120);
and AND4 (N20290, N20275, N8327, N9161, N14355);
xor XOR2 (N20291, N20282, N3412);
buf BUF1 (N20292, N20291);
or OR4 (N20293, N20290, N3248, N8343, N3897);
nor NOR3 (N20294, N20286, N5025, N17694);
or OR4 (N20295, N20284, N1150, N14062, N8531);
xor XOR2 (N20296, N20293, N3473);
buf BUF1 (N20297, N20280);
xor XOR2 (N20298, N20295, N7884);
nor NOR4 (N20299, N20294, N1433, N15133, N11840);
buf BUF1 (N20300, N20281);
and AND4 (N20301, N20299, N14887, N18838, N11628);
not NOT1 (N20302, N20296);
nor NOR2 (N20303, N20285, N18683);
nand NAND2 (N20304, N20287, N182);
buf BUF1 (N20305, N20302);
nor NOR2 (N20306, N20305, N7258);
nor NOR4 (N20307, N20301, N5627, N9070, N15403);
buf BUF1 (N20308, N20303);
and AND3 (N20309, N20306, N12107, N13521);
or OR2 (N20310, N20300, N1307);
not NOT1 (N20311, N20288);
not NOT1 (N20312, N20309);
buf BUF1 (N20313, N20311);
xor XOR2 (N20314, N20310, N4444);
nor NOR2 (N20315, N20312, N9024);
buf BUF1 (N20316, N20289);
or OR3 (N20317, N20298, N12771, N2887);
and AND3 (N20318, N20292, N12969, N17879);
xor XOR2 (N20319, N20314, N19097);
not NOT1 (N20320, N20319);
and AND2 (N20321, N20297, N4124);
buf BUF1 (N20322, N20316);
nand NAND4 (N20323, N20317, N14336, N4613, N9781);
xor XOR2 (N20324, N20321, N12474);
nor NOR4 (N20325, N20320, N774, N4192, N5241);
xor XOR2 (N20326, N20322, N11195);
xor XOR2 (N20327, N20308, N12157);
nor NOR2 (N20328, N20324, N5657);
buf BUF1 (N20329, N20327);
nor NOR2 (N20330, N20326, N16724);
nand NAND4 (N20331, N20330, N6154, N5607, N20266);
nor NOR2 (N20332, N20329, N14904);
nand NAND2 (N20333, N20307, N19595);
nand NAND3 (N20334, N20325, N3683, N13058);
nor NOR4 (N20335, N20304, N8000, N11405, N13352);
xor XOR2 (N20336, N20328, N12101);
nor NOR4 (N20337, N20332, N13315, N11163, N3963);
and AND2 (N20338, N20334, N2579);
not NOT1 (N20339, N20337);
or OR3 (N20340, N20313, N7592, N14380);
or OR2 (N20341, N20338, N8157);
buf BUF1 (N20342, N20341);
xor XOR2 (N20343, N20339, N13677);
and AND3 (N20344, N20343, N19037, N3329);
buf BUF1 (N20345, N20344);
nand NAND3 (N20346, N20333, N3163, N14524);
xor XOR2 (N20347, N20340, N3629);
or OR3 (N20348, N20315, N18895, N12820);
not NOT1 (N20349, N20348);
or OR2 (N20350, N20345, N18132);
nand NAND4 (N20351, N20350, N17642, N20032, N18924);
not NOT1 (N20352, N20351);
not NOT1 (N20353, N20346);
nand NAND3 (N20354, N20352, N8119, N13207);
buf BUF1 (N20355, N20318);
not NOT1 (N20356, N20331);
buf BUF1 (N20357, N20354);
xor XOR2 (N20358, N20347, N4675);
nand NAND4 (N20359, N20323, N12774, N18128, N12210);
xor XOR2 (N20360, N20353, N2585);
nand NAND2 (N20361, N20360, N18333);
or OR3 (N20362, N20361, N14811, N6115);
and AND3 (N20363, N20335, N17168, N4132);
xor XOR2 (N20364, N20358, N18024);
nor NOR3 (N20365, N20356, N12434, N20082);
nor NOR4 (N20366, N20342, N1907, N13904, N3728);
nor NOR2 (N20367, N20359, N9837);
not NOT1 (N20368, N20363);
xor XOR2 (N20369, N20366, N4868);
nand NAND4 (N20370, N20368, N20103, N1021, N11581);
not NOT1 (N20371, N20336);
buf BUF1 (N20372, N20365);
buf BUF1 (N20373, N20371);
xor XOR2 (N20374, N20355, N10287);
xor XOR2 (N20375, N20370, N11014);
not NOT1 (N20376, N20373);
nand NAND3 (N20377, N20369, N9791, N7077);
xor XOR2 (N20378, N20377, N3359);
not NOT1 (N20379, N20364);
nor NOR4 (N20380, N20372, N283, N4068, N11184);
nor NOR2 (N20381, N20375, N3368);
and AND3 (N20382, N20349, N19147, N12311);
nand NAND4 (N20383, N20380, N7110, N19414, N1899);
nand NAND3 (N20384, N20367, N6462, N5807);
nand NAND3 (N20385, N20376, N9074, N10076);
buf BUF1 (N20386, N20362);
nand NAND2 (N20387, N20378, N10823);
or OR2 (N20388, N20381, N2467);
xor XOR2 (N20389, N20357, N5);
and AND2 (N20390, N20374, N13383);
nand NAND3 (N20391, N20379, N5399, N1903);
and AND4 (N20392, N20388, N9876, N1921, N19857);
not NOT1 (N20393, N20384);
buf BUF1 (N20394, N20392);
or OR3 (N20395, N20394, N13814, N18670);
nand NAND3 (N20396, N20383, N18808, N8003);
xor XOR2 (N20397, N20389, N3240);
or OR2 (N20398, N20396, N13546);
xor XOR2 (N20399, N20393, N10);
not NOT1 (N20400, N20397);
buf BUF1 (N20401, N20398);
and AND3 (N20402, N20387, N16568, N2368);
or OR4 (N20403, N20382, N1760, N5352, N1816);
or OR2 (N20404, N20402, N6832);
not NOT1 (N20405, N20401);
and AND2 (N20406, N20404, N9884);
or OR2 (N20407, N20406, N5635);
buf BUF1 (N20408, N20386);
and AND2 (N20409, N20385, N19218);
nor NOR2 (N20410, N20405, N12011);
nor NOR3 (N20411, N20407, N13137, N2178);
nor NOR4 (N20412, N20411, N7290, N3790, N8905);
xor XOR2 (N20413, N20399, N8027);
nor NOR4 (N20414, N20395, N9248, N12263, N4378);
and AND4 (N20415, N20409, N3329, N589, N2794);
nor NOR2 (N20416, N20415, N10598);
not NOT1 (N20417, N20412);
nand NAND3 (N20418, N20391, N18672, N19091);
and AND4 (N20419, N20403, N3369, N12684, N10941);
nor NOR2 (N20420, N20390, N19304);
or OR3 (N20421, N20413, N6898, N17153);
xor XOR2 (N20422, N20417, N19251);
or OR3 (N20423, N20400, N3393, N8046);
buf BUF1 (N20424, N20420);
buf BUF1 (N20425, N20419);
xor XOR2 (N20426, N20425, N2156);
nand NAND2 (N20427, N20426, N16633);
nand NAND3 (N20428, N20410, N10695, N14888);
nor NOR2 (N20429, N20418, N1126);
not NOT1 (N20430, N20423);
nor NOR4 (N20431, N20429, N3282, N15420, N10496);
buf BUF1 (N20432, N20416);
buf BUF1 (N20433, N20414);
buf BUF1 (N20434, N20421);
nor NOR3 (N20435, N20433, N10258, N7924);
or OR4 (N20436, N20431, N4670, N7746, N14453);
not NOT1 (N20437, N20432);
or OR3 (N20438, N20422, N1084, N4480);
not NOT1 (N20439, N20438);
and AND4 (N20440, N20439, N11816, N16101, N2839);
nor NOR4 (N20441, N20424, N3777, N11739, N8004);
or OR3 (N20442, N20435, N5982, N16144);
xor XOR2 (N20443, N20427, N11050);
xor XOR2 (N20444, N20437, N327);
nand NAND4 (N20445, N20436, N5143, N9278, N11447);
nor NOR3 (N20446, N20443, N5963, N4246);
xor XOR2 (N20447, N20442, N9193);
nand NAND3 (N20448, N20434, N20438, N7035);
nor NOR3 (N20449, N20408, N12454, N17025);
or OR4 (N20450, N20447, N8538, N10167, N12486);
or OR4 (N20451, N20449, N4952, N15055, N15503);
not NOT1 (N20452, N20441);
not NOT1 (N20453, N20445);
nor NOR2 (N20454, N20453, N1822);
xor XOR2 (N20455, N20446, N13211);
and AND4 (N20456, N20448, N4017, N2881, N11690);
not NOT1 (N20457, N20455);
buf BUF1 (N20458, N20430);
not NOT1 (N20459, N20456);
buf BUF1 (N20460, N20458);
buf BUF1 (N20461, N20460);
nand NAND4 (N20462, N20450, N19234, N15374, N18868);
buf BUF1 (N20463, N20451);
or OR4 (N20464, N20461, N19227, N16008, N2854);
or OR2 (N20465, N20452, N20332);
buf BUF1 (N20466, N20440);
nand NAND4 (N20467, N20459, N13227, N20400, N6757);
and AND2 (N20468, N20462, N8896);
buf BUF1 (N20469, N20444);
xor XOR2 (N20470, N20466, N17485);
or OR4 (N20471, N20454, N16070, N14904, N18485);
nor NOR4 (N20472, N20464, N7146, N18368, N9558);
and AND2 (N20473, N20472, N1272);
not NOT1 (N20474, N20467);
or OR2 (N20475, N20469, N6713);
xor XOR2 (N20476, N20473, N2932);
and AND2 (N20477, N20468, N17339);
xor XOR2 (N20478, N20474, N12783);
not NOT1 (N20479, N20476);
nand NAND4 (N20480, N20477, N76, N6675, N10715);
nor NOR4 (N20481, N20470, N3487, N15868, N3302);
xor XOR2 (N20482, N20471, N5128);
and AND3 (N20483, N20481, N16202, N11734);
and AND4 (N20484, N20428, N16616, N19182, N19071);
nor NOR4 (N20485, N20465, N14614, N14653, N8560);
not NOT1 (N20486, N20475);
not NOT1 (N20487, N20482);
xor XOR2 (N20488, N20484, N18719);
nand NAND4 (N20489, N20486, N16260, N945, N17795);
and AND2 (N20490, N20479, N12022);
nor NOR3 (N20491, N20485, N14245, N18458);
nand NAND4 (N20492, N20480, N9853, N9619, N15841);
nor NOR2 (N20493, N20457, N10492);
xor XOR2 (N20494, N20491, N20481);
or OR3 (N20495, N20493, N4620, N6492);
not NOT1 (N20496, N20492);
or OR4 (N20497, N20494, N4590, N4154, N20337);
buf BUF1 (N20498, N20489);
nor NOR2 (N20499, N20487, N17057);
xor XOR2 (N20500, N20483, N16065);
nand NAND2 (N20501, N20495, N4905);
buf BUF1 (N20502, N20496);
or OR4 (N20503, N20478, N13250, N5720, N18919);
nor NOR4 (N20504, N20488, N487, N382, N18372);
or OR4 (N20505, N20503, N2999, N3316, N19716);
or OR2 (N20506, N20463, N1780);
nor NOR3 (N20507, N20502, N7541, N15068);
not NOT1 (N20508, N20504);
buf BUF1 (N20509, N20501);
nor NOR4 (N20510, N20505, N14030, N3457, N12918);
xor XOR2 (N20511, N20508, N6753);
and AND4 (N20512, N20499, N1898, N7950, N9958);
or OR4 (N20513, N20498, N12252, N4953, N8061);
and AND2 (N20514, N20500, N3744);
nor NOR3 (N20515, N20512, N15978, N5654);
not NOT1 (N20516, N20490);
xor XOR2 (N20517, N20509, N18406);
nand NAND4 (N20518, N20506, N19385, N3448, N13123);
buf BUF1 (N20519, N20514);
xor XOR2 (N20520, N20507, N8753);
or OR3 (N20521, N20516, N1545, N15122);
not NOT1 (N20522, N20518);
xor XOR2 (N20523, N20515, N12274);
and AND2 (N20524, N20511, N15510);
nor NOR3 (N20525, N20523, N3370, N11434);
buf BUF1 (N20526, N20520);
and AND3 (N20527, N20525, N11756, N12003);
nand NAND3 (N20528, N20510, N19721, N19215);
or OR3 (N20529, N20521, N5258, N3377);
buf BUF1 (N20530, N20527);
nand NAND3 (N20531, N20529, N18451, N1892);
nand NAND2 (N20532, N20517, N6365);
xor XOR2 (N20533, N20532, N12382);
and AND4 (N20534, N20519, N2195, N10657, N6718);
xor XOR2 (N20535, N20530, N10888);
xor XOR2 (N20536, N20533, N9667);
or OR2 (N20537, N20528, N4038);
or OR3 (N20538, N20497, N15908, N3139);
not NOT1 (N20539, N20538);
not NOT1 (N20540, N20513);
xor XOR2 (N20541, N20537, N8981);
and AND4 (N20542, N20535, N19433, N10531, N17804);
or OR3 (N20543, N20524, N8474, N10228);
and AND3 (N20544, N20531, N19293, N17937);
nor NOR4 (N20545, N20541, N3496, N1758, N7173);
not NOT1 (N20546, N20540);
nor NOR2 (N20547, N20536, N4405);
nor NOR3 (N20548, N20542, N11696, N15589);
nor NOR3 (N20549, N20539, N19452, N6031);
and AND3 (N20550, N20543, N1858, N5955);
not NOT1 (N20551, N20522);
or OR2 (N20552, N20544, N10426);
xor XOR2 (N20553, N20549, N15915);
xor XOR2 (N20554, N20551, N15977);
buf BUF1 (N20555, N20534);
nor NOR3 (N20556, N20547, N11036, N2797);
buf BUF1 (N20557, N20556);
nand NAND2 (N20558, N20555, N1665);
buf BUF1 (N20559, N20550);
buf BUF1 (N20560, N20553);
not NOT1 (N20561, N20552);
not NOT1 (N20562, N20545);
nand NAND4 (N20563, N20562, N16546, N16200, N329);
and AND4 (N20564, N20546, N19706, N3059, N16153);
or OR4 (N20565, N20564, N2868, N17561, N19232);
nor NOR3 (N20566, N20561, N12279, N9027);
or OR3 (N20567, N20557, N167, N7883);
nand NAND3 (N20568, N20565, N16299, N513);
not NOT1 (N20569, N20563);
not NOT1 (N20570, N20554);
xor XOR2 (N20571, N20526, N4432);
and AND2 (N20572, N20570, N18288);
xor XOR2 (N20573, N20566, N14790);
nand NAND4 (N20574, N20571, N14274, N3019, N13991);
and AND3 (N20575, N20558, N4305, N1854);
nor NOR4 (N20576, N20560, N13803, N199, N6209);
or OR3 (N20577, N20568, N3042, N3236);
nand NAND2 (N20578, N20574, N10750);
buf BUF1 (N20579, N20578);
buf BUF1 (N20580, N20572);
or OR3 (N20581, N20580, N13180, N14193);
xor XOR2 (N20582, N20577, N10537);
and AND3 (N20583, N20548, N11491, N13196);
buf BUF1 (N20584, N20569);
nand NAND4 (N20585, N20583, N2129, N15808, N19653);
buf BUF1 (N20586, N20573);
nor NOR3 (N20587, N20585, N4350, N18685);
xor XOR2 (N20588, N20582, N14498);
nand NAND2 (N20589, N20559, N14346);
and AND3 (N20590, N20589, N9553, N3997);
buf BUF1 (N20591, N20584);
nand NAND3 (N20592, N20588, N6237, N10096);
and AND4 (N20593, N20567, N974, N19227, N7955);
xor XOR2 (N20594, N20593, N3608);
nand NAND3 (N20595, N20587, N14163, N19088);
not NOT1 (N20596, N20592);
not NOT1 (N20597, N20586);
nor NOR2 (N20598, N20575, N2185);
or OR4 (N20599, N20598, N16439, N18898, N10711);
nand NAND2 (N20600, N20590, N11065);
xor XOR2 (N20601, N20596, N11354);
buf BUF1 (N20602, N20576);
or OR2 (N20603, N20591, N16819);
xor XOR2 (N20604, N20600, N1239);
nor NOR3 (N20605, N20599, N16736, N6919);
xor XOR2 (N20606, N20603, N10630);
nor NOR4 (N20607, N20606, N12572, N17397, N6187);
or OR4 (N20608, N20581, N20158, N17593, N19526);
or OR3 (N20609, N20602, N16426, N15879);
or OR3 (N20610, N20601, N4737, N13445);
and AND2 (N20611, N20607, N1116);
nor NOR3 (N20612, N20604, N19210, N14225);
not NOT1 (N20613, N20612);
and AND3 (N20614, N20595, N18147, N19130);
and AND3 (N20615, N20605, N7253, N17593);
not NOT1 (N20616, N20579);
and AND3 (N20617, N20616, N6826, N8049);
buf BUF1 (N20618, N20613);
or OR2 (N20619, N20609, N17907);
or OR4 (N20620, N20608, N18552, N19932, N3881);
and AND4 (N20621, N20614, N4842, N16064, N635);
or OR3 (N20622, N20618, N6377, N4523);
buf BUF1 (N20623, N20620);
or OR3 (N20624, N20594, N10005, N9773);
not NOT1 (N20625, N20610);
nor NOR4 (N20626, N20611, N8907, N5836, N8601);
nand NAND4 (N20627, N20625, N12129, N16118, N11076);
not NOT1 (N20628, N20617);
xor XOR2 (N20629, N20615, N9969);
buf BUF1 (N20630, N20626);
or OR3 (N20631, N20621, N10522, N3545);
not NOT1 (N20632, N20627);
and AND2 (N20633, N20629, N11928);
or OR3 (N20634, N20630, N8712, N8058);
nor NOR3 (N20635, N20622, N20388, N15152);
buf BUF1 (N20636, N20635);
nor NOR4 (N20637, N20636, N16303, N19126, N15708);
and AND4 (N20638, N20637, N5630, N17377, N6086);
nand NAND4 (N20639, N20632, N6745, N4681, N8045);
or OR2 (N20640, N20623, N10072);
nand NAND2 (N20641, N20631, N15154);
and AND3 (N20642, N20619, N12649, N12521);
nor NOR2 (N20643, N20624, N2137);
xor XOR2 (N20644, N20641, N8572);
or OR3 (N20645, N20642, N6157, N6421);
nand NAND2 (N20646, N20633, N17038);
buf BUF1 (N20647, N20640);
or OR4 (N20648, N20639, N596, N2356, N2433);
buf BUF1 (N20649, N20628);
buf BUF1 (N20650, N20638);
and AND4 (N20651, N20643, N14617, N17220, N14699);
xor XOR2 (N20652, N20646, N10437);
buf BUF1 (N20653, N20650);
or OR3 (N20654, N20652, N11610, N20582);
buf BUF1 (N20655, N20649);
nor NOR4 (N20656, N20654, N5367, N6964, N4247);
or OR2 (N20657, N20645, N7472);
and AND3 (N20658, N20634, N17845, N14524);
or OR4 (N20659, N20644, N1415, N16174, N11321);
and AND4 (N20660, N20648, N9745, N173, N7262);
not NOT1 (N20661, N20653);
nor NOR2 (N20662, N20656, N5024);
nor NOR3 (N20663, N20662, N5440, N1861);
and AND3 (N20664, N20651, N9051, N15466);
nor NOR3 (N20665, N20660, N18304, N13710);
not NOT1 (N20666, N20655);
nor NOR2 (N20667, N20647, N1032);
buf BUF1 (N20668, N20664);
nand NAND4 (N20669, N20657, N2957, N7352, N12965);
not NOT1 (N20670, N20659);
nor NOR3 (N20671, N20669, N13156, N4815);
nor NOR3 (N20672, N20658, N20306, N16612);
nand NAND4 (N20673, N20668, N6914, N13115, N19371);
not NOT1 (N20674, N20663);
not NOT1 (N20675, N20667);
xor XOR2 (N20676, N20675, N5488);
and AND2 (N20677, N20673, N8230);
xor XOR2 (N20678, N20597, N15205);
not NOT1 (N20679, N20672);
buf BUF1 (N20680, N20676);
nor NOR2 (N20681, N20666, N423);
and AND3 (N20682, N20661, N16819, N13130);
xor XOR2 (N20683, N20678, N17347);
and AND4 (N20684, N20679, N5858, N8788, N9146);
xor XOR2 (N20685, N20680, N13225);
nand NAND3 (N20686, N20685, N1657, N14689);
xor XOR2 (N20687, N20681, N3715);
buf BUF1 (N20688, N20670);
nor NOR3 (N20689, N20665, N16526, N6327);
buf BUF1 (N20690, N20684);
nor NOR3 (N20691, N20687, N7199, N12395);
nand NAND3 (N20692, N20677, N15055, N16688);
and AND4 (N20693, N20688, N8150, N10896, N1446);
nor NOR3 (N20694, N20693, N11911, N18629);
nand NAND2 (N20695, N20689, N6563);
buf BUF1 (N20696, N20683);
buf BUF1 (N20697, N20691);
and AND2 (N20698, N20682, N15125);
or OR2 (N20699, N20695, N19488);
not NOT1 (N20700, N20686);
not NOT1 (N20701, N20692);
nand NAND4 (N20702, N20697, N15658, N19410, N7613);
not NOT1 (N20703, N20698);
buf BUF1 (N20704, N20699);
and AND4 (N20705, N20704, N13829, N10460, N644);
xor XOR2 (N20706, N20696, N1400);
nor NOR3 (N20707, N20674, N5899, N3882);
xor XOR2 (N20708, N20694, N17070);
and AND3 (N20709, N20703, N11986, N14123);
or OR3 (N20710, N20671, N5908, N735);
nor NOR4 (N20711, N20701, N7076, N2940, N18495);
xor XOR2 (N20712, N20690, N20420);
or OR4 (N20713, N20707, N10484, N4063, N12400);
buf BUF1 (N20714, N20711);
and AND3 (N20715, N20706, N20613, N8906);
not NOT1 (N20716, N20713);
xor XOR2 (N20717, N20708, N10695);
buf BUF1 (N20718, N20702);
xor XOR2 (N20719, N20710, N1781);
or OR2 (N20720, N20718, N17890);
xor XOR2 (N20721, N20719, N3038);
and AND3 (N20722, N20712, N360, N18565);
or OR3 (N20723, N20720, N5856, N11639);
nand NAND3 (N20724, N20717, N17421, N9659);
not NOT1 (N20725, N20705);
not NOT1 (N20726, N20723);
or OR3 (N20727, N20724, N15012, N15064);
and AND4 (N20728, N20716, N8143, N778, N2037);
nand NAND3 (N20729, N20728, N6661, N1297);
and AND3 (N20730, N20715, N7673, N3747);
or OR3 (N20731, N20700, N10315, N20595);
and AND3 (N20732, N20731, N9683, N20113);
or OR2 (N20733, N20709, N8085);
nor NOR2 (N20734, N20729, N18472);
and AND2 (N20735, N20714, N19126);
and AND3 (N20736, N20721, N7184, N19168);
nand NAND2 (N20737, N20730, N3918);
buf BUF1 (N20738, N20737);
or OR3 (N20739, N20735, N16474, N19851);
or OR3 (N20740, N20727, N8718, N9714);
nor NOR4 (N20741, N20722, N9207, N18143, N3906);
nand NAND2 (N20742, N20725, N12182);
nor NOR3 (N20743, N20742, N10161, N11289);
buf BUF1 (N20744, N20734);
buf BUF1 (N20745, N20738);
xor XOR2 (N20746, N20732, N15467);
not NOT1 (N20747, N20726);
or OR3 (N20748, N20736, N449, N18674);
nor NOR3 (N20749, N20741, N572, N20090);
xor XOR2 (N20750, N20739, N13993);
nand NAND3 (N20751, N20747, N15028, N4513);
nand NAND3 (N20752, N20746, N14883, N12824);
xor XOR2 (N20753, N20733, N17633);
nand NAND4 (N20754, N20740, N20680, N9753, N17117);
not NOT1 (N20755, N20744);
or OR4 (N20756, N20751, N12559, N6304, N5338);
nand NAND2 (N20757, N20743, N17306);
and AND4 (N20758, N20745, N11327, N6471, N6244);
xor XOR2 (N20759, N20749, N6855);
buf BUF1 (N20760, N20757);
nand NAND4 (N20761, N20759, N2627, N7607, N19025);
nand NAND4 (N20762, N20760, N11474, N8342, N20348);
nor NOR3 (N20763, N20748, N20667, N13534);
nand NAND2 (N20764, N20756, N12656);
nand NAND4 (N20765, N20752, N6033, N9003, N4436);
and AND3 (N20766, N20750, N1285, N17368);
nand NAND4 (N20767, N20758, N14169, N20337, N7649);
or OR2 (N20768, N20764, N16333);
not NOT1 (N20769, N20761);
and AND2 (N20770, N20763, N14190);
buf BUF1 (N20771, N20762);
or OR4 (N20772, N20767, N372, N19075, N5248);
xor XOR2 (N20773, N20770, N9977);
not NOT1 (N20774, N20769);
or OR2 (N20775, N20754, N15603);
buf BUF1 (N20776, N20753);
nand NAND3 (N20777, N20772, N20131, N17646);
and AND2 (N20778, N20773, N15841);
nand NAND2 (N20779, N20771, N3937);
nand NAND2 (N20780, N20755, N3768);
or OR3 (N20781, N20775, N20349, N14746);
nor NOR3 (N20782, N20765, N3600, N7985);
xor XOR2 (N20783, N20777, N16538);
and AND3 (N20784, N20780, N19367, N8550);
not NOT1 (N20785, N20781);
nand NAND3 (N20786, N20783, N1403, N737);
xor XOR2 (N20787, N20778, N11421);
nor NOR2 (N20788, N20766, N10883);
buf BUF1 (N20789, N20786);
xor XOR2 (N20790, N20768, N2809);
or OR2 (N20791, N20785, N17023);
and AND4 (N20792, N20782, N10601, N11013, N1372);
or OR4 (N20793, N20774, N15478, N18315, N18172);
or OR4 (N20794, N20784, N6288, N20605, N19346);
nor NOR3 (N20795, N20776, N19499, N12205);
nand NAND4 (N20796, N20789, N678, N20242, N18131);
and AND4 (N20797, N20793, N3656, N13759, N11750);
or OR4 (N20798, N20796, N8862, N17216, N13083);
xor XOR2 (N20799, N20797, N9416);
nand NAND2 (N20800, N20795, N1381);
nand NAND2 (N20801, N20792, N13549);
nand NAND3 (N20802, N20801, N229, N15931);
xor XOR2 (N20803, N20794, N10292);
nor NOR3 (N20804, N20798, N17326, N1879);
buf BUF1 (N20805, N20799);
and AND2 (N20806, N20788, N10808);
not NOT1 (N20807, N20805);
buf BUF1 (N20808, N20800);
nand NAND2 (N20809, N20806, N4529);
or OR4 (N20810, N20807, N3205, N10741, N17960);
or OR4 (N20811, N20810, N14866, N97, N7464);
and AND3 (N20812, N20779, N17527, N1760);
nand NAND4 (N20813, N20804, N13454, N1176, N1397);
buf BUF1 (N20814, N20802);
xor XOR2 (N20815, N20808, N4724);
nand NAND2 (N20816, N20791, N17757);
nand NAND3 (N20817, N20816, N746, N16787);
xor XOR2 (N20818, N20787, N14458);
nand NAND3 (N20819, N20818, N9225, N14611);
buf BUF1 (N20820, N20817);
buf BUF1 (N20821, N20811);
not NOT1 (N20822, N20790);
nand NAND2 (N20823, N20821, N11643);
nor NOR3 (N20824, N20815, N12840, N16970);
nand NAND2 (N20825, N20814, N1208);
not NOT1 (N20826, N20809);
buf BUF1 (N20827, N20824);
or OR4 (N20828, N20803, N18317, N11702, N17969);
or OR3 (N20829, N20813, N5623, N15697);
not NOT1 (N20830, N20812);
or OR2 (N20831, N20825, N17163);
nand NAND3 (N20832, N20827, N7116, N10088);
and AND4 (N20833, N20823, N1067, N9968, N10916);
and AND3 (N20834, N20820, N7098, N12288);
nand NAND2 (N20835, N20819, N9696);
and AND4 (N20836, N20828, N9991, N8559, N3925);
and AND4 (N20837, N20822, N3116, N6448, N19396);
and AND3 (N20838, N20831, N15702, N6566);
xor XOR2 (N20839, N20832, N18229);
or OR2 (N20840, N20834, N12102);
and AND3 (N20841, N20840, N17810, N4141);
not NOT1 (N20842, N20838);
xor XOR2 (N20843, N20842, N1805);
nor NOR2 (N20844, N20826, N4563);
or OR4 (N20845, N20830, N7216, N17465, N348);
buf BUF1 (N20846, N20837);
and AND2 (N20847, N20844, N10861);
not NOT1 (N20848, N20846);
nor NOR4 (N20849, N20829, N7815, N14257, N2172);
not NOT1 (N20850, N20843);
or OR4 (N20851, N20845, N20310, N18990, N2319);
and AND2 (N20852, N20833, N15493);
xor XOR2 (N20853, N20835, N14700);
or OR4 (N20854, N20849, N7840, N7975, N19953);
xor XOR2 (N20855, N20854, N2481);
xor XOR2 (N20856, N20855, N7615);
buf BUF1 (N20857, N20848);
or OR4 (N20858, N20847, N4485, N13444, N9242);
buf BUF1 (N20859, N20836);
and AND3 (N20860, N20853, N4472, N19982);
not NOT1 (N20861, N20859);
nor NOR2 (N20862, N20861, N1101);
nor NOR2 (N20863, N20841, N12003);
nor NOR2 (N20864, N20839, N17811);
or OR2 (N20865, N20864, N18784);
buf BUF1 (N20866, N20857);
buf BUF1 (N20867, N20866);
buf BUF1 (N20868, N20850);
not NOT1 (N20869, N20867);
and AND4 (N20870, N20856, N16733, N12601, N9027);
buf BUF1 (N20871, N20860);
buf BUF1 (N20872, N20868);
and AND4 (N20873, N20865, N13657, N171, N8149);
nand NAND2 (N20874, N20858, N5546);
or OR3 (N20875, N20872, N12743, N11056);
buf BUF1 (N20876, N20871);
or OR2 (N20877, N20851, N7274);
not NOT1 (N20878, N20873);
nor NOR2 (N20879, N20852, N19270);
buf BUF1 (N20880, N20870);
xor XOR2 (N20881, N20876, N15157);
and AND3 (N20882, N20877, N8375, N10136);
not NOT1 (N20883, N20869);
and AND3 (N20884, N20878, N14336, N18837);
or OR4 (N20885, N20884, N4123, N4583, N8365);
nor NOR2 (N20886, N20885, N13287);
xor XOR2 (N20887, N20880, N12688);
buf BUF1 (N20888, N20879);
or OR2 (N20889, N20862, N15262);
and AND3 (N20890, N20875, N15538, N20070);
xor XOR2 (N20891, N20883, N13130);
nand NAND3 (N20892, N20890, N13500, N6341);
or OR4 (N20893, N20891, N6238, N13223, N9504);
and AND3 (N20894, N20893, N17535, N17349);
and AND3 (N20895, N20889, N14595, N15599);
buf BUF1 (N20896, N20874);
xor XOR2 (N20897, N20892, N11955);
xor XOR2 (N20898, N20894, N15210);
buf BUF1 (N20899, N20863);
buf BUF1 (N20900, N20895);
and AND3 (N20901, N20886, N13326, N2362);
nor NOR4 (N20902, N20900, N16139, N1034, N10830);
xor XOR2 (N20903, N20898, N11395);
and AND2 (N20904, N20902, N3452);
buf BUF1 (N20905, N20881);
nor NOR4 (N20906, N20887, N19312, N7444, N1126);
buf BUF1 (N20907, N20904);
buf BUF1 (N20908, N20882);
xor XOR2 (N20909, N20901, N13261);
or OR3 (N20910, N20908, N6829, N13104);
nor NOR3 (N20911, N20888, N12281, N18968);
nand NAND4 (N20912, N20906, N16351, N9075, N4193);
xor XOR2 (N20913, N20912, N20602);
buf BUF1 (N20914, N20896);
buf BUF1 (N20915, N20899);
buf BUF1 (N20916, N20915);
xor XOR2 (N20917, N20914, N12578);
nor NOR2 (N20918, N20911, N8006);
not NOT1 (N20919, N20913);
and AND3 (N20920, N20919, N20615, N20825);
and AND4 (N20921, N20918, N268, N3779, N16714);
xor XOR2 (N20922, N20897, N485);
not NOT1 (N20923, N20921);
buf BUF1 (N20924, N20909);
not NOT1 (N20925, N20924);
or OR4 (N20926, N20916, N16975, N10688, N4092);
not NOT1 (N20927, N20923);
nor NOR3 (N20928, N20910, N18218, N3665);
nand NAND2 (N20929, N20903, N16921);
or OR3 (N20930, N20907, N2875, N5292);
not NOT1 (N20931, N20922);
or OR4 (N20932, N20931, N20380, N13435, N4356);
buf BUF1 (N20933, N20929);
or OR4 (N20934, N20917, N7664, N952, N2146);
nand NAND3 (N20935, N20926, N5361, N1093);
or OR3 (N20936, N20925, N20013, N18348);
and AND3 (N20937, N20933, N6231, N20846);
nor NOR3 (N20938, N20935, N1646, N1314);
xor XOR2 (N20939, N20937, N4367);
not NOT1 (N20940, N20934);
and AND2 (N20941, N20939, N20836);
and AND2 (N20942, N20927, N4270);
and AND4 (N20943, N20942, N4759, N18687, N3128);
xor XOR2 (N20944, N20943, N7032);
buf BUF1 (N20945, N20941);
or OR4 (N20946, N20932, N15742, N16392, N1205);
or OR3 (N20947, N20920, N5415, N2805);
or OR2 (N20948, N20938, N8801);
or OR2 (N20949, N20945, N13447);
not NOT1 (N20950, N20936);
or OR2 (N20951, N20944, N8641);
nor NOR4 (N20952, N20948, N12652, N147, N13934);
xor XOR2 (N20953, N20951, N16507);
buf BUF1 (N20954, N20940);
buf BUF1 (N20955, N20905);
or OR2 (N20956, N20930, N2777);
or OR4 (N20957, N20954, N15940, N2230, N14767);
buf BUF1 (N20958, N20950);
and AND2 (N20959, N20949, N956);
and AND4 (N20960, N20958, N2253, N4853, N211);
not NOT1 (N20961, N20952);
xor XOR2 (N20962, N20956, N15719);
xor XOR2 (N20963, N20960, N13368);
or OR3 (N20964, N20959, N17575, N544);
or OR4 (N20965, N20955, N10386, N3510, N8781);
xor XOR2 (N20966, N20953, N8941);
nand NAND4 (N20967, N20964, N16839, N11579, N9722);
xor XOR2 (N20968, N20962, N8229);
xor XOR2 (N20969, N20968, N5949);
and AND3 (N20970, N20957, N4142, N142);
buf BUF1 (N20971, N20928);
and AND4 (N20972, N20969, N12782, N2772, N9853);
nand NAND2 (N20973, N20961, N18433);
or OR3 (N20974, N20971, N19529, N18684);
or OR2 (N20975, N20974, N10379);
nor NOR3 (N20976, N20963, N10296, N16909);
buf BUF1 (N20977, N20972);
not NOT1 (N20978, N20966);
nand NAND2 (N20979, N20946, N9203);
and AND3 (N20980, N20976, N19335, N15130);
nand NAND3 (N20981, N20979, N10716, N4422);
xor XOR2 (N20982, N20965, N20274);
and AND3 (N20983, N20981, N12520, N13956);
not NOT1 (N20984, N20975);
not NOT1 (N20985, N20980);
nand NAND2 (N20986, N20967, N18779);
xor XOR2 (N20987, N20977, N9650);
buf BUF1 (N20988, N20987);
nor NOR2 (N20989, N20986, N822);
xor XOR2 (N20990, N20989, N576);
or OR3 (N20991, N20947, N2454, N12152);
or OR4 (N20992, N20982, N6682, N20444, N7791);
nor NOR2 (N20993, N20991, N3958);
nor NOR4 (N20994, N20993, N9043, N16633, N2274);
buf BUF1 (N20995, N20990);
xor XOR2 (N20996, N20973, N13067);
xor XOR2 (N20997, N20984, N14658);
nor NOR4 (N20998, N20996, N1332, N8941, N16136);
nor NOR3 (N20999, N20995, N765, N10718);
xor XOR2 (N21000, N20978, N1394);
not NOT1 (N21001, N20998);
not NOT1 (N21002, N20994);
nand NAND2 (N21003, N20999, N8715);
buf BUF1 (N21004, N20997);
xor XOR2 (N21005, N21001, N11841);
or OR2 (N21006, N21002, N3852);
buf BUF1 (N21007, N21004);
nand NAND4 (N21008, N21006, N18261, N19476, N3314);
not NOT1 (N21009, N21007);
buf BUF1 (N21010, N21005);
not NOT1 (N21011, N20970);
and AND3 (N21012, N20988, N2014, N4563);
nor NOR2 (N21013, N20992, N5125);
and AND4 (N21014, N21013, N6907, N6162, N2721);
nand NAND3 (N21015, N21011, N11330, N13931);
or OR2 (N21016, N21009, N2506);
xor XOR2 (N21017, N21010, N3470);
not NOT1 (N21018, N21017);
nand NAND4 (N21019, N20985, N17853, N20378, N11855);
not NOT1 (N21020, N21008);
nor NOR4 (N21021, N21000, N4200, N18392, N16125);
or OR4 (N21022, N21014, N8523, N10019, N17903);
nor NOR2 (N21023, N20983, N113);
nand NAND2 (N21024, N21019, N9067);
buf BUF1 (N21025, N21024);
and AND3 (N21026, N21023, N16511, N3434);
xor XOR2 (N21027, N21022, N12584);
and AND4 (N21028, N21018, N16221, N10371, N3095);
and AND4 (N21029, N21003, N5010, N11260, N9911);
nor NOR3 (N21030, N21016, N8057, N13658);
xor XOR2 (N21031, N21021, N19825);
nand NAND3 (N21032, N21031, N7036, N5055);
and AND4 (N21033, N21012, N9591, N3793, N17975);
and AND3 (N21034, N21015, N14909, N14869);
nor NOR4 (N21035, N21029, N19387, N7441, N12034);
buf BUF1 (N21036, N21032);
not NOT1 (N21037, N21026);
or OR4 (N21038, N21028, N19456, N13478, N13676);
xor XOR2 (N21039, N21027, N6496);
and AND3 (N21040, N21039, N3370, N9721);
and AND2 (N21041, N21034, N16457);
xor XOR2 (N21042, N21033, N6753);
xor XOR2 (N21043, N21036, N9740);
buf BUF1 (N21044, N21038);
and AND2 (N21045, N21043, N6013);
nor NOR4 (N21046, N21020, N3521, N17146, N13797);
nor NOR2 (N21047, N21040, N8006);
and AND3 (N21048, N21047, N11196, N19250);
or OR2 (N21049, N21030, N1162);
buf BUF1 (N21050, N21048);
or OR2 (N21051, N21045, N20927);
nor NOR2 (N21052, N21042, N9021);
xor XOR2 (N21053, N21049, N20539);
and AND2 (N21054, N21053, N14826);
nand NAND3 (N21055, N21054, N15422, N20212);
not NOT1 (N21056, N21037);
xor XOR2 (N21057, N21044, N9218);
nor NOR3 (N21058, N21052, N13180, N4757);
or OR3 (N21059, N21041, N20038, N18368);
nor NOR2 (N21060, N21056, N16400);
nand NAND2 (N21061, N21046, N20005);
not NOT1 (N21062, N21025);
and AND4 (N21063, N21060, N5862, N2486, N15784);
not NOT1 (N21064, N21051);
nor NOR3 (N21065, N21062, N5946, N9411);
not NOT1 (N21066, N21050);
nand NAND2 (N21067, N21058, N18154);
xor XOR2 (N21068, N21064, N2490);
and AND2 (N21069, N21055, N8175);
not NOT1 (N21070, N21057);
nor NOR2 (N21071, N21065, N5584);
nand NAND4 (N21072, N21067, N19935, N8746, N15937);
or OR3 (N21073, N21061, N4430, N21046);
nor NOR4 (N21074, N21066, N3636, N9878, N3835);
nor NOR4 (N21075, N21068, N16624, N20687, N5484);
nand NAND4 (N21076, N21071, N17795, N6781, N13585);
or OR3 (N21077, N21059, N10516, N1750);
not NOT1 (N21078, N21073);
not NOT1 (N21079, N21069);
buf BUF1 (N21080, N21070);
and AND2 (N21081, N21079, N18066);
not NOT1 (N21082, N21081);
or OR3 (N21083, N21035, N9111, N12430);
not NOT1 (N21084, N21063);
or OR4 (N21085, N21077, N11261, N13392, N3571);
and AND4 (N21086, N21084, N7488, N15728, N1215);
not NOT1 (N21087, N21085);
nor NOR3 (N21088, N21078, N19228, N15984);
nand NAND4 (N21089, N21074, N20719, N11208, N403);
buf BUF1 (N21090, N21082);
or OR2 (N21091, N21090, N11919);
and AND4 (N21092, N21088, N17325, N8196, N3744);
buf BUF1 (N21093, N21080);
buf BUF1 (N21094, N21087);
buf BUF1 (N21095, N21086);
or OR2 (N21096, N21095, N11059);
nor NOR3 (N21097, N21072, N10123, N13042);
nor NOR2 (N21098, N21083, N16411);
nand NAND3 (N21099, N21089, N2166, N1704);
xor XOR2 (N21100, N21094, N1892);
and AND2 (N21101, N21097, N1354);
not NOT1 (N21102, N21101);
nand NAND3 (N21103, N21098, N17772, N5763);
buf BUF1 (N21104, N21103);
nand NAND4 (N21105, N21102, N15280, N14290, N19802);
xor XOR2 (N21106, N21091, N20798);
nor NOR2 (N21107, N21100, N10179);
or OR4 (N21108, N21075, N11297, N8835, N13290);
buf BUF1 (N21109, N21104);
not NOT1 (N21110, N21093);
or OR3 (N21111, N21110, N15327, N14626);
buf BUF1 (N21112, N21076);
nor NOR2 (N21113, N21096, N348);
xor XOR2 (N21114, N21112, N15348);
and AND3 (N21115, N21099, N2672, N2875);
not NOT1 (N21116, N21105);
and AND2 (N21117, N21092, N1828);
nand NAND4 (N21118, N21107, N10190, N3777, N19137);
not NOT1 (N21119, N21111);
not NOT1 (N21120, N21108);
nor NOR2 (N21121, N21118, N7448);
nor NOR3 (N21122, N21115, N18504, N342);
buf BUF1 (N21123, N21122);
xor XOR2 (N21124, N21120, N713);
buf BUF1 (N21125, N21123);
not NOT1 (N21126, N21125);
xor XOR2 (N21127, N21116, N1054);
or OR4 (N21128, N21124, N18778, N2848, N9653);
nand NAND4 (N21129, N21128, N20013, N19844, N17991);
or OR2 (N21130, N21106, N11074);
and AND3 (N21131, N21117, N12835, N15811);
xor XOR2 (N21132, N21113, N11971);
not NOT1 (N21133, N21130);
or OR3 (N21134, N21119, N7925, N16005);
nand NAND4 (N21135, N21114, N4737, N7689, N6514);
nor NOR2 (N21136, N21135, N20964);
or OR4 (N21137, N21133, N18292, N9710, N5159);
nor NOR4 (N21138, N21127, N8100, N18557, N4191);
and AND4 (N21139, N21132, N18369, N11334, N8445);
xor XOR2 (N21140, N21137, N5301);
xor XOR2 (N21141, N21134, N5474);
nand NAND2 (N21142, N21140, N15840);
xor XOR2 (N21143, N21121, N16395);
not NOT1 (N21144, N21136);
not NOT1 (N21145, N21143);
buf BUF1 (N21146, N21142);
not NOT1 (N21147, N21109);
not NOT1 (N21148, N21141);
xor XOR2 (N21149, N21126, N12942);
not NOT1 (N21150, N21139);
nand NAND4 (N21151, N21131, N5531, N13246, N13076);
nand NAND3 (N21152, N21148, N17647, N15176);
nor NOR2 (N21153, N21149, N19209);
xor XOR2 (N21154, N21145, N19487);
or OR2 (N21155, N21153, N10621);
and AND2 (N21156, N21138, N13375);
nor NOR4 (N21157, N21146, N19010, N18459, N1380);
nor NOR4 (N21158, N21156, N7333, N2962, N13653);
nor NOR4 (N21159, N21129, N13528, N8171, N8877);
not NOT1 (N21160, N21144);
buf BUF1 (N21161, N21158);
and AND3 (N21162, N21155, N16848, N11734);
and AND4 (N21163, N21160, N19734, N7150, N14182);
buf BUF1 (N21164, N21154);
buf BUF1 (N21165, N21150);
and AND2 (N21166, N21152, N5098);
not NOT1 (N21167, N21147);
and AND4 (N21168, N21162, N8708, N9301, N15045);
xor XOR2 (N21169, N21163, N10871);
or OR4 (N21170, N21169, N9373, N18109, N9013);
or OR2 (N21171, N21166, N6130);
xor XOR2 (N21172, N21159, N2749);
xor XOR2 (N21173, N21161, N2114);
nor NOR2 (N21174, N21167, N3019);
not NOT1 (N21175, N21171);
buf BUF1 (N21176, N21175);
nor NOR3 (N21177, N21168, N1709, N3331);
not NOT1 (N21178, N21172);
or OR2 (N21179, N21157, N9734);
not NOT1 (N21180, N21176);
nand NAND2 (N21181, N21151, N13266);
xor XOR2 (N21182, N21181, N7435);
xor XOR2 (N21183, N21164, N2944);
nor NOR2 (N21184, N21180, N13869);
nand NAND2 (N21185, N21173, N17906);
buf BUF1 (N21186, N21177);
and AND4 (N21187, N21174, N20754, N411, N3583);
nand NAND4 (N21188, N21178, N9189, N13772, N532);
and AND2 (N21189, N21185, N4963);
not NOT1 (N21190, N21165);
buf BUF1 (N21191, N21190);
buf BUF1 (N21192, N21191);
not NOT1 (N21193, N21183);
or OR3 (N21194, N21182, N5709, N15842);
xor XOR2 (N21195, N21179, N17907);
or OR3 (N21196, N21195, N3308, N15819);
nand NAND2 (N21197, N21170, N16622);
nand NAND2 (N21198, N21184, N7985);
buf BUF1 (N21199, N21187);
buf BUF1 (N21200, N21186);
and AND3 (N21201, N21192, N236, N2935);
nor NOR2 (N21202, N21201, N20325);
buf BUF1 (N21203, N21199);
buf BUF1 (N21204, N21193);
nor NOR3 (N21205, N21203, N14636, N17235);
xor XOR2 (N21206, N21200, N16189);
or OR4 (N21207, N21194, N5293, N16319, N20534);
or OR4 (N21208, N21196, N9895, N13690, N6705);
buf BUF1 (N21209, N21189);
xor XOR2 (N21210, N21209, N18381);
buf BUF1 (N21211, N21204);
nand NAND2 (N21212, N21211, N9106);
and AND3 (N21213, N21205, N9191, N11733);
and AND4 (N21214, N21188, N7131, N16664, N4247);
not NOT1 (N21215, N21206);
or OR4 (N21216, N21207, N3215, N20739, N150);
and AND2 (N21217, N21215, N20827);
and AND3 (N21218, N21198, N11630, N8766);
nor NOR3 (N21219, N21197, N3561, N18707);
and AND4 (N21220, N21219, N138, N16019, N7278);
or OR2 (N21221, N21202, N15190);
or OR3 (N21222, N21212, N12305, N14535);
nor NOR4 (N21223, N21218, N10041, N13985, N13517);
nor NOR4 (N21224, N21217, N1338, N10816, N4430);
nor NOR3 (N21225, N21220, N215, N6846);
not NOT1 (N21226, N21221);
or OR2 (N21227, N21216, N13386);
nor NOR3 (N21228, N21208, N17019, N8285);
not NOT1 (N21229, N21223);
buf BUF1 (N21230, N21228);
and AND3 (N21231, N21226, N6050, N14157);
xor XOR2 (N21232, N21222, N14174);
xor XOR2 (N21233, N21229, N1974);
buf BUF1 (N21234, N21224);
and AND4 (N21235, N21213, N569, N13974, N10527);
nand NAND2 (N21236, N21235, N10942);
or OR2 (N21237, N21227, N15790);
nor NOR4 (N21238, N21210, N9364, N3607, N4110);
buf BUF1 (N21239, N21237);
nand NAND4 (N21240, N21233, N10216, N9004, N498);
xor XOR2 (N21241, N21230, N17979);
or OR3 (N21242, N21238, N17143, N16111);
and AND4 (N21243, N21240, N5560, N7390, N12410);
not NOT1 (N21244, N21241);
nand NAND4 (N21245, N21231, N6331, N16423, N7199);
xor XOR2 (N21246, N21245, N9826);
xor XOR2 (N21247, N21214, N12333);
and AND2 (N21248, N21239, N10115);
nor NOR2 (N21249, N21234, N17550);
or OR3 (N21250, N21249, N11575, N15881);
not NOT1 (N21251, N21242);
or OR2 (N21252, N21248, N2389);
and AND4 (N21253, N21225, N14198, N15956, N10429);
not NOT1 (N21254, N21250);
not NOT1 (N21255, N21253);
and AND3 (N21256, N21252, N3245, N2178);
xor XOR2 (N21257, N21256, N18009);
buf BUF1 (N21258, N21257);
buf BUF1 (N21259, N21255);
nor NOR3 (N21260, N21258, N8838, N15838);
and AND2 (N21261, N21247, N21161);
xor XOR2 (N21262, N21254, N15839);
buf BUF1 (N21263, N21232);
xor XOR2 (N21264, N21243, N5329);
buf BUF1 (N21265, N21261);
xor XOR2 (N21266, N21263, N18436);
xor XOR2 (N21267, N21244, N2295);
xor XOR2 (N21268, N21236, N7611);
and AND4 (N21269, N21246, N4336, N10620, N17594);
xor XOR2 (N21270, N21269, N13988);
not NOT1 (N21271, N21265);
not NOT1 (N21272, N21268);
nor NOR3 (N21273, N21262, N12096, N2482);
not NOT1 (N21274, N21264);
buf BUF1 (N21275, N21273);
nor NOR4 (N21276, N21275, N9931, N17974, N9842);
nor NOR4 (N21277, N21271, N16479, N3552, N20969);
nand NAND3 (N21278, N21266, N17781, N21028);
nor NOR3 (N21279, N21259, N10307, N4173);
buf BUF1 (N21280, N21276);
nor NOR4 (N21281, N21277, N4715, N14102, N7770);
xor XOR2 (N21282, N21272, N14367);
xor XOR2 (N21283, N21278, N17211);
nor NOR4 (N21284, N21251, N1774, N18894, N9498);
buf BUF1 (N21285, N21282);
and AND4 (N21286, N21270, N14339, N3778, N4571);
not NOT1 (N21287, N21279);
or OR3 (N21288, N21285, N11451, N16098);
and AND3 (N21289, N21284, N17081, N8125);
nand NAND4 (N21290, N21267, N18646, N14523, N13066);
and AND3 (N21291, N21288, N588, N11415);
or OR2 (N21292, N21280, N3304);
or OR3 (N21293, N21287, N16961, N17971);
xor XOR2 (N21294, N21292, N9659);
xor XOR2 (N21295, N21260, N6457);
not NOT1 (N21296, N21295);
nor NOR4 (N21297, N21290, N2259, N15718, N13825);
nand NAND3 (N21298, N21289, N7462, N5386);
buf BUF1 (N21299, N21291);
not NOT1 (N21300, N21298);
not NOT1 (N21301, N21293);
and AND2 (N21302, N21300, N18104);
buf BUF1 (N21303, N21286);
nand NAND4 (N21304, N21302, N5212, N10732, N15803);
not NOT1 (N21305, N21304);
buf BUF1 (N21306, N21274);
and AND2 (N21307, N21301, N20290);
not NOT1 (N21308, N21307);
nor NOR3 (N21309, N21281, N5480, N18543);
buf BUF1 (N21310, N21283);
buf BUF1 (N21311, N21296);
or OR4 (N21312, N21309, N4856, N456, N9243);
xor XOR2 (N21313, N21310, N5256);
and AND4 (N21314, N21312, N7786, N8037, N12885);
buf BUF1 (N21315, N21297);
not NOT1 (N21316, N21315);
xor XOR2 (N21317, N21311, N20424);
buf BUF1 (N21318, N21314);
buf BUF1 (N21319, N21317);
or OR2 (N21320, N21318, N15021);
buf BUF1 (N21321, N21305);
and AND3 (N21322, N21306, N20844, N1099);
or OR2 (N21323, N21303, N3603);
buf BUF1 (N21324, N21321);
nor NOR2 (N21325, N21299, N19348);
xor XOR2 (N21326, N21323, N5328);
buf BUF1 (N21327, N21320);
and AND3 (N21328, N21308, N6124, N14535);
nor NOR2 (N21329, N21319, N10379);
and AND2 (N21330, N21294, N3989);
nand NAND2 (N21331, N21322, N15720);
nor NOR2 (N21332, N21324, N18046);
not NOT1 (N21333, N21325);
xor XOR2 (N21334, N21326, N19621);
or OR2 (N21335, N21327, N4943);
or OR3 (N21336, N21334, N13986, N357);
not NOT1 (N21337, N21313);
nand NAND4 (N21338, N21335, N17707, N10208, N13410);
xor XOR2 (N21339, N21329, N9865);
nand NAND3 (N21340, N21337, N10212, N2049);
not NOT1 (N21341, N21333);
buf BUF1 (N21342, N21338);
xor XOR2 (N21343, N21330, N11392);
and AND2 (N21344, N21340, N7817);
nor NOR2 (N21345, N21342, N3373);
or OR4 (N21346, N21328, N17059, N20461, N7320);
nor NOR2 (N21347, N21346, N15692);
or OR3 (N21348, N21344, N14309, N15490);
nor NOR2 (N21349, N21348, N9292);
nand NAND2 (N21350, N21316, N18580);
nor NOR4 (N21351, N21349, N16718, N21242, N8976);
and AND2 (N21352, N21331, N2029);
or OR3 (N21353, N21332, N17188, N5399);
xor XOR2 (N21354, N21350, N16632);
nand NAND3 (N21355, N21353, N9198, N9336);
not NOT1 (N21356, N21339);
nor NOR2 (N21357, N21354, N14119);
not NOT1 (N21358, N21336);
nor NOR4 (N21359, N21358, N17308, N2734, N887);
nor NOR2 (N21360, N21355, N6117);
not NOT1 (N21361, N21352);
buf BUF1 (N21362, N21359);
not NOT1 (N21363, N21341);
nand NAND2 (N21364, N21362, N17757);
and AND3 (N21365, N21361, N12180, N14722);
and AND3 (N21366, N21345, N5291, N4709);
not NOT1 (N21367, N21357);
nor NOR3 (N21368, N21360, N17351, N13464);
nor NOR3 (N21369, N21364, N1423, N10300);
not NOT1 (N21370, N21356);
buf BUF1 (N21371, N21369);
nor NOR4 (N21372, N21363, N18838, N6715, N20294);
nor NOR2 (N21373, N21371, N10182);
not NOT1 (N21374, N21366);
nor NOR3 (N21375, N21351, N17938, N9845);
or OR2 (N21376, N21372, N11007);
nand NAND4 (N21377, N21365, N5224, N16456, N19716);
nand NAND4 (N21378, N21374, N16723, N4066, N9991);
and AND4 (N21379, N21376, N5653, N2984, N16813);
nor NOR3 (N21380, N21370, N2966, N3647);
or OR2 (N21381, N21367, N15557);
or OR3 (N21382, N21377, N3873, N18476);
nand NAND2 (N21383, N21373, N13971);
or OR3 (N21384, N21347, N911, N2684);
and AND4 (N21385, N21368, N13683, N5954, N12338);
nor NOR4 (N21386, N21384, N13434, N13153, N4916);
nand NAND3 (N21387, N21378, N13400, N19099);
or OR3 (N21388, N21385, N21051, N5367);
and AND4 (N21389, N21380, N10989, N3584, N17034);
nor NOR3 (N21390, N21387, N6584, N8530);
and AND4 (N21391, N21379, N1850, N19024, N10175);
buf BUF1 (N21392, N21381);
nand NAND3 (N21393, N21382, N5917, N13553);
or OR2 (N21394, N21383, N924);
buf BUF1 (N21395, N21375);
nor NOR3 (N21396, N21390, N3699, N14633);
not NOT1 (N21397, N21388);
nand NAND3 (N21398, N21394, N8962, N8558);
and AND4 (N21399, N21397, N1471, N8760, N4962);
and AND4 (N21400, N21391, N18230, N14870, N6802);
not NOT1 (N21401, N21389);
xor XOR2 (N21402, N21395, N8421);
not NOT1 (N21403, N21392);
xor XOR2 (N21404, N21398, N20580);
nand NAND3 (N21405, N21396, N672, N7776);
or OR3 (N21406, N21403, N6071, N12924);
or OR3 (N21407, N21393, N290, N13243);
buf BUF1 (N21408, N21343);
nand NAND2 (N21409, N21407, N5676);
not NOT1 (N21410, N21404);
buf BUF1 (N21411, N21399);
nor NOR4 (N21412, N21402, N20223, N17721, N10340);
nor NOR4 (N21413, N21401, N5600, N12456, N14286);
buf BUF1 (N21414, N21408);
buf BUF1 (N21415, N21409);
or OR3 (N21416, N21411, N19001, N17623);
not NOT1 (N21417, N21410);
nor NOR3 (N21418, N21416, N15205, N13667);
buf BUF1 (N21419, N21400);
xor XOR2 (N21420, N21419, N16033);
nand NAND3 (N21421, N21414, N1842, N17339);
not NOT1 (N21422, N21412);
buf BUF1 (N21423, N21415);
not NOT1 (N21424, N21420);
not NOT1 (N21425, N21405);
not NOT1 (N21426, N21421);
nor NOR3 (N21427, N21413, N9547, N19966);
and AND4 (N21428, N21386, N7475, N18431, N1468);
xor XOR2 (N21429, N21423, N4660);
buf BUF1 (N21430, N21425);
not NOT1 (N21431, N21430);
xor XOR2 (N21432, N21427, N20646);
not NOT1 (N21433, N21428);
buf BUF1 (N21434, N21429);
nand NAND2 (N21435, N21406, N7039);
and AND3 (N21436, N21431, N7860, N20583);
xor XOR2 (N21437, N21426, N16461);
xor XOR2 (N21438, N21435, N19404);
nand NAND3 (N21439, N21433, N3397, N1950);
nand NAND2 (N21440, N21437, N603);
not NOT1 (N21441, N21432);
nor NOR2 (N21442, N21438, N14760);
nand NAND4 (N21443, N21439, N15336, N9112, N8379);
not NOT1 (N21444, N21442);
and AND2 (N21445, N21440, N14782);
xor XOR2 (N21446, N21422, N2983);
xor XOR2 (N21447, N21445, N1613);
nand NAND4 (N21448, N21447, N18411, N11611, N3729);
and AND3 (N21449, N21424, N20686, N10862);
not NOT1 (N21450, N21434);
buf BUF1 (N21451, N21449);
and AND3 (N21452, N21448, N6511, N11475);
and AND3 (N21453, N21417, N10113, N8784);
not NOT1 (N21454, N21441);
buf BUF1 (N21455, N21454);
nor NOR4 (N21456, N21452, N13561, N13514, N20663);
buf BUF1 (N21457, N21453);
nor NOR2 (N21458, N21450, N20247);
xor XOR2 (N21459, N21418, N18576);
nor NOR4 (N21460, N21444, N19109, N9941, N9113);
buf BUF1 (N21461, N21455);
buf BUF1 (N21462, N21436);
and AND2 (N21463, N21461, N10994);
nor NOR4 (N21464, N21462, N21163, N19155, N11177);
and AND4 (N21465, N21460, N15677, N11715, N4883);
nor NOR2 (N21466, N21459, N16941);
nor NOR2 (N21467, N21463, N19833);
and AND2 (N21468, N21466, N15281);
nand NAND2 (N21469, N21467, N921);
xor XOR2 (N21470, N21464, N8828);
nand NAND3 (N21471, N21470, N16813, N16195);
nand NAND2 (N21472, N21465, N21457);
and AND2 (N21473, N14057, N8640);
xor XOR2 (N21474, N21473, N3342);
and AND4 (N21475, N21451, N14970, N17209, N6371);
nor NOR2 (N21476, N21469, N12104);
nand NAND2 (N21477, N21456, N13335);
nand NAND4 (N21478, N21468, N40, N1305, N5168);
buf BUF1 (N21479, N21471);
buf BUF1 (N21480, N21443);
nor NOR4 (N21481, N21479, N9975, N8807, N19457);
and AND3 (N21482, N21478, N20905, N13184);
nand NAND4 (N21483, N21481, N3528, N20160, N4907);
not NOT1 (N21484, N21482);
xor XOR2 (N21485, N21446, N4577);
xor XOR2 (N21486, N21474, N12748);
buf BUF1 (N21487, N21484);
xor XOR2 (N21488, N21458, N13009);
and AND4 (N21489, N21476, N21477, N5760, N17372);
xor XOR2 (N21490, N11033, N1837);
buf BUF1 (N21491, N21475);
and AND4 (N21492, N21489, N18227, N12524, N17940);
and AND3 (N21493, N21490, N1562, N13914);
nor NOR3 (N21494, N21493, N16974, N6170);
buf BUF1 (N21495, N21485);
nor NOR3 (N21496, N21492, N14143, N6660);
or OR2 (N21497, N21472, N5570);
buf BUF1 (N21498, N21480);
and AND4 (N21499, N21497, N15333, N19648, N15686);
and AND4 (N21500, N21496, N14518, N8217, N18735);
not NOT1 (N21501, N21488);
buf BUF1 (N21502, N21500);
not NOT1 (N21503, N21498);
nor NOR3 (N21504, N21499, N20469, N19938);
or OR3 (N21505, N21503, N14970, N4080);
xor XOR2 (N21506, N21491, N7858);
or OR4 (N21507, N21487, N18082, N2313, N328);
xor XOR2 (N21508, N21502, N9459);
buf BUF1 (N21509, N21483);
nor NOR3 (N21510, N21501, N2694, N21359);
xor XOR2 (N21511, N21508, N9834);
xor XOR2 (N21512, N21486, N12308);
or OR2 (N21513, N21511, N20757);
nand NAND3 (N21514, N21510, N3315, N18827);
nand NAND3 (N21515, N21504, N5658, N13293);
or OR2 (N21516, N21495, N19147);
buf BUF1 (N21517, N21512);
or OR4 (N21518, N21505, N14205, N7017, N20697);
and AND2 (N21519, N21514, N18150);
nor NOR2 (N21520, N21506, N11623);
not NOT1 (N21521, N21515);
not NOT1 (N21522, N21509);
buf BUF1 (N21523, N21518);
xor XOR2 (N21524, N21521, N11452);
buf BUF1 (N21525, N21523);
xor XOR2 (N21526, N21507, N8414);
and AND3 (N21527, N21522, N20988, N14025);
not NOT1 (N21528, N21516);
or OR4 (N21529, N21517, N5171, N11793, N13741);
xor XOR2 (N21530, N21525, N3363);
buf BUF1 (N21531, N21519);
xor XOR2 (N21532, N21529, N10733);
not NOT1 (N21533, N21530);
and AND4 (N21534, N21532, N2239, N18683, N7141);
xor XOR2 (N21535, N21527, N6075);
buf BUF1 (N21536, N21533);
or OR2 (N21537, N21513, N189);
nand NAND3 (N21538, N21528, N19369, N19281);
not NOT1 (N21539, N21535);
nor NOR4 (N21540, N21539, N8783, N8111, N3848);
nor NOR4 (N21541, N21534, N18954, N619, N16517);
buf BUF1 (N21542, N21531);
or OR2 (N21543, N21494, N11154);
and AND3 (N21544, N21526, N17118, N16482);
buf BUF1 (N21545, N21537);
buf BUF1 (N21546, N21540);
xor XOR2 (N21547, N21543, N11441);
nand NAND3 (N21548, N21546, N16541, N5745);
buf BUF1 (N21549, N21520);
and AND2 (N21550, N21536, N20709);
and AND4 (N21551, N21548, N19510, N1362, N10916);
or OR4 (N21552, N21545, N36, N16495, N17685);
nand NAND3 (N21553, N21551, N10290, N14268);
xor XOR2 (N21554, N21544, N10476);
buf BUF1 (N21555, N21538);
xor XOR2 (N21556, N21555, N6702);
or OR4 (N21557, N21552, N13645, N17755, N3316);
or OR4 (N21558, N21554, N15672, N21322, N14095);
nor NOR2 (N21559, N21542, N6421);
or OR2 (N21560, N21559, N16528);
nand NAND2 (N21561, N21557, N11093);
buf BUF1 (N21562, N21561);
nor NOR2 (N21563, N21562, N16933);
or OR3 (N21564, N21558, N3284, N9320);
not NOT1 (N21565, N21553);
nand NAND3 (N21566, N21524, N4256, N13329);
nor NOR3 (N21567, N21556, N1018, N614);
buf BUF1 (N21568, N21550);
xor XOR2 (N21569, N21563, N21257);
not NOT1 (N21570, N21541);
nand NAND4 (N21571, N21567, N16231, N6432, N1287);
nand NAND2 (N21572, N21547, N3370);
nor NOR4 (N21573, N21568, N11666, N19166, N4615);
xor XOR2 (N21574, N21571, N10909);
and AND3 (N21575, N21572, N12526, N17614);
nand NAND4 (N21576, N21564, N8588, N9432, N19491);
and AND2 (N21577, N21575, N16674);
xor XOR2 (N21578, N21577, N7727);
xor XOR2 (N21579, N21565, N3415);
and AND2 (N21580, N21569, N18695);
not NOT1 (N21581, N21580);
nand NAND3 (N21582, N21574, N16792, N16083);
not NOT1 (N21583, N21579);
xor XOR2 (N21584, N21566, N15269);
not NOT1 (N21585, N21584);
and AND2 (N21586, N21570, N14853);
nand NAND2 (N21587, N21585, N17238);
nand NAND3 (N21588, N21560, N11971, N21466);
nor NOR2 (N21589, N21582, N20590);
xor XOR2 (N21590, N21578, N4521);
xor XOR2 (N21591, N21587, N1167);
nor NOR4 (N21592, N21576, N2312, N20689, N1349);
and AND4 (N21593, N21592, N7174, N12972, N13036);
nor NOR2 (N21594, N21588, N13728);
and AND3 (N21595, N21549, N18807, N20024);
nand NAND2 (N21596, N21595, N6422);
or OR4 (N21597, N21586, N12437, N112, N13096);
nand NAND3 (N21598, N21573, N10848, N12283);
not NOT1 (N21599, N21590);
or OR2 (N21600, N21597, N10109);
nor NOR2 (N21601, N21598, N2397);
or OR2 (N21602, N21589, N14358);
nand NAND4 (N21603, N21581, N17492, N2998, N3807);
nand NAND3 (N21604, N21601, N21003, N20569);
and AND3 (N21605, N21604, N2980, N16918);
nand NAND4 (N21606, N21602, N2619, N2174, N15231);
or OR4 (N21607, N21596, N6345, N15680, N16991);
not NOT1 (N21608, N21593);
buf BUF1 (N21609, N21583);
nand NAND2 (N21610, N21591, N2225);
nor NOR3 (N21611, N21599, N15497, N3764);
and AND3 (N21612, N21594, N11714, N14273);
buf BUF1 (N21613, N21609);
nor NOR2 (N21614, N21603, N19482);
not NOT1 (N21615, N21613);
not NOT1 (N21616, N21612);
or OR3 (N21617, N21608, N7404, N6575);
or OR4 (N21618, N21617, N17867, N18229, N1663);
buf BUF1 (N21619, N21614);
buf BUF1 (N21620, N21615);
nand NAND3 (N21621, N21607, N9608, N12600);
not NOT1 (N21622, N21606);
buf BUF1 (N21623, N21621);
and AND4 (N21624, N21620, N6542, N3817, N19874);
nor NOR4 (N21625, N21616, N18800, N2489, N5557);
or OR3 (N21626, N21625, N1666, N10598);
and AND3 (N21627, N21619, N2733, N6843);
not NOT1 (N21628, N21600);
nand NAND4 (N21629, N21628, N11285, N1314, N6748);
nor NOR3 (N21630, N21605, N14300, N14236);
or OR3 (N21631, N21618, N12011, N6030);
not NOT1 (N21632, N21626);
and AND3 (N21633, N21631, N17332, N550);
nor NOR3 (N21634, N21633, N17206, N6334);
or OR4 (N21635, N21624, N12978, N15480, N7926);
not NOT1 (N21636, N21610);
not NOT1 (N21637, N21635);
or OR3 (N21638, N21636, N17907, N2998);
nand NAND4 (N21639, N21627, N21440, N6276, N15316);
not NOT1 (N21640, N21623);
not NOT1 (N21641, N21622);
not NOT1 (N21642, N21637);
nand NAND4 (N21643, N21639, N17423, N1970, N1270);
buf BUF1 (N21644, N21629);
nor NOR4 (N21645, N21634, N3727, N3920, N13674);
buf BUF1 (N21646, N21645);
nand NAND3 (N21647, N21630, N11495, N5934);
xor XOR2 (N21648, N21641, N18529);
or OR3 (N21649, N21643, N5276, N4264);
and AND4 (N21650, N21647, N10184, N3070, N20554);
and AND2 (N21651, N21648, N226);
and AND2 (N21652, N21646, N6268);
and AND2 (N21653, N21642, N20570);
and AND3 (N21654, N21644, N7814, N19289);
nand NAND4 (N21655, N21652, N11764, N18275, N7543);
or OR4 (N21656, N21650, N5080, N21291, N7597);
or OR2 (N21657, N21640, N2313);
buf BUF1 (N21658, N21657);
nand NAND3 (N21659, N21655, N8525, N9057);
and AND4 (N21660, N21656, N7866, N17118, N12956);
nand NAND3 (N21661, N21653, N8302, N5341);
nor NOR4 (N21662, N21632, N12410, N3405, N19517);
nand NAND4 (N21663, N21651, N10601, N21358, N20550);
not NOT1 (N21664, N21659);
buf BUF1 (N21665, N21663);
xor XOR2 (N21666, N21662, N11461);
buf BUF1 (N21667, N21654);
nor NOR4 (N21668, N21660, N18980, N15104, N950);
nor NOR4 (N21669, N21666, N3639, N13720, N12869);
xor XOR2 (N21670, N21638, N10004);
not NOT1 (N21671, N21664);
nand NAND3 (N21672, N21671, N11688, N6065);
and AND3 (N21673, N21649, N13815, N5620);
nand NAND2 (N21674, N21669, N7549);
or OR4 (N21675, N21670, N5690, N13953, N19800);
not NOT1 (N21676, N21674);
nand NAND3 (N21677, N21667, N1830, N7124);
nor NOR4 (N21678, N21658, N20262, N19584, N20742);
nor NOR4 (N21679, N21661, N11468, N1579, N18616);
not NOT1 (N21680, N21672);
nand NAND3 (N21681, N21679, N12797, N15878);
nand NAND2 (N21682, N21681, N1416);
nor NOR3 (N21683, N21673, N12174, N5278);
and AND2 (N21684, N21683, N20743);
xor XOR2 (N21685, N21675, N12334);
or OR2 (N21686, N21682, N7089);
not NOT1 (N21687, N21678);
buf BUF1 (N21688, N21677);
nor NOR4 (N21689, N21687, N7257, N9578, N17455);
not NOT1 (N21690, N21676);
and AND2 (N21691, N21611, N18274);
or OR2 (N21692, N21685, N12122);
buf BUF1 (N21693, N21680);
not NOT1 (N21694, N21693);
nor NOR2 (N21695, N21665, N16193);
or OR3 (N21696, N21668, N8569, N8764);
xor XOR2 (N21697, N21689, N3261);
buf BUF1 (N21698, N21696);
and AND2 (N21699, N21688, N12204);
nand NAND3 (N21700, N21690, N8027, N8682);
and AND4 (N21701, N21695, N19074, N2856, N8784);
nand NAND3 (N21702, N21686, N987, N18029);
nor NOR4 (N21703, N21691, N14782, N5284, N19380);
buf BUF1 (N21704, N21684);
xor XOR2 (N21705, N21699, N11975);
nand NAND4 (N21706, N21700, N6717, N924, N18103);
xor XOR2 (N21707, N21692, N12455);
nor NOR4 (N21708, N21702, N18888, N4504, N18282);
or OR2 (N21709, N21703, N3732);
or OR4 (N21710, N21707, N6067, N7339, N18922);
or OR3 (N21711, N21697, N6803, N16371);
nand NAND4 (N21712, N21709, N1648, N8815, N6623);
not NOT1 (N21713, N21705);
buf BUF1 (N21714, N21701);
nand NAND4 (N21715, N21711, N5026, N18667, N4332);
xor XOR2 (N21716, N21710, N3933);
or OR4 (N21717, N21708, N10301, N20923, N15801);
not NOT1 (N21718, N21717);
nand NAND2 (N21719, N21713, N20463);
xor XOR2 (N21720, N21715, N4936);
buf BUF1 (N21721, N21704);
buf BUF1 (N21722, N21712);
not NOT1 (N21723, N21698);
not NOT1 (N21724, N21714);
nand NAND3 (N21725, N21694, N21563, N19420);
nor NOR3 (N21726, N21716, N9464, N3799);
and AND4 (N21727, N21706, N7525, N3375, N6719);
nand NAND3 (N21728, N21718, N12919, N9441);
and AND3 (N21729, N21728, N2765, N14673);
or OR2 (N21730, N21720, N11723);
and AND4 (N21731, N21723, N9059, N14487, N17434);
and AND4 (N21732, N21730, N7710, N17906, N4086);
xor XOR2 (N21733, N21729, N15081);
xor XOR2 (N21734, N21724, N13866);
or OR4 (N21735, N21719, N17730, N2158, N1974);
not NOT1 (N21736, N21731);
or OR3 (N21737, N21733, N17327, N10880);
buf BUF1 (N21738, N21736);
nor NOR4 (N21739, N21722, N4850, N13844, N2392);
buf BUF1 (N21740, N21737);
nand NAND2 (N21741, N21734, N5707);
buf BUF1 (N21742, N21732);
xor XOR2 (N21743, N21741, N13305);
and AND4 (N21744, N21726, N4237, N4005, N10360);
or OR2 (N21745, N21742, N11810);
not NOT1 (N21746, N21735);
buf BUF1 (N21747, N21744);
buf BUF1 (N21748, N21740);
or OR3 (N21749, N21739, N12148, N10861);
xor XOR2 (N21750, N21749, N16631);
xor XOR2 (N21751, N21745, N2428);
and AND3 (N21752, N21721, N498, N16715);
or OR4 (N21753, N21748, N4427, N15252, N12524);
or OR2 (N21754, N21751, N16475);
and AND3 (N21755, N21747, N18405, N14935);
nor NOR3 (N21756, N21738, N12320, N13440);
or OR3 (N21757, N21725, N5000, N12957);
and AND4 (N21758, N21746, N6956, N1436, N6805);
nand NAND4 (N21759, N21758, N18366, N15548, N12751);
buf BUF1 (N21760, N21756);
nand NAND2 (N21761, N21727, N416);
or OR2 (N21762, N21755, N20918);
and AND3 (N21763, N21757, N14690, N3045);
not NOT1 (N21764, N21743);
not NOT1 (N21765, N21752);
nand NAND2 (N21766, N21760, N13106);
nor NOR4 (N21767, N21763, N16118, N19797, N12468);
xor XOR2 (N21768, N21767, N1394);
buf BUF1 (N21769, N21750);
not NOT1 (N21770, N21768);
xor XOR2 (N21771, N21770, N11946);
nor NOR2 (N21772, N21769, N14036);
buf BUF1 (N21773, N21759);
buf BUF1 (N21774, N21753);
not NOT1 (N21775, N21761);
buf BUF1 (N21776, N21774);
not NOT1 (N21777, N21754);
and AND3 (N21778, N21762, N1480, N7139);
or OR4 (N21779, N21772, N15524, N13443, N11441);
nor NOR2 (N21780, N21765, N10733);
or OR4 (N21781, N21771, N3875, N114, N11755);
or OR2 (N21782, N21776, N17776);
xor XOR2 (N21783, N21777, N11067);
nand NAND3 (N21784, N21778, N10268, N228);
or OR4 (N21785, N21784, N6315, N2558, N18516);
xor XOR2 (N21786, N21764, N1984);
not NOT1 (N21787, N21780);
not NOT1 (N21788, N21787);
nand NAND3 (N21789, N21782, N16273, N6808);
or OR4 (N21790, N21783, N12249, N7250, N8313);
and AND2 (N21791, N21786, N5625);
buf BUF1 (N21792, N21779);
and AND4 (N21793, N21775, N14697, N21403, N57);
or OR3 (N21794, N21791, N15207, N8063);
nand NAND2 (N21795, N21781, N21671);
not NOT1 (N21796, N21789);
nor NOR3 (N21797, N21796, N9657, N19377);
or OR3 (N21798, N21794, N15790, N18990);
not NOT1 (N21799, N21792);
nor NOR4 (N21800, N21773, N9170, N9003, N20785);
buf BUF1 (N21801, N21797);
buf BUF1 (N21802, N21766);
buf BUF1 (N21803, N21798);
buf BUF1 (N21804, N21800);
nor NOR4 (N21805, N21802, N11268, N16946, N6294);
xor XOR2 (N21806, N21801, N7823);
or OR3 (N21807, N21785, N12002, N11220);
or OR4 (N21808, N21803, N8294, N19852, N17088);
nand NAND3 (N21809, N21793, N2802, N6831);
nor NOR4 (N21810, N21808, N20572, N16992, N13845);
nand NAND4 (N21811, N21795, N12047, N8460, N7420);
xor XOR2 (N21812, N21809, N20077);
or OR3 (N21813, N21807, N314, N20827);
not NOT1 (N21814, N21810);
nand NAND4 (N21815, N21788, N21555, N18765, N21286);
nand NAND3 (N21816, N21805, N20817, N11422);
nand NAND4 (N21817, N21814, N14071, N17521, N20203);
not NOT1 (N21818, N21817);
or OR4 (N21819, N21804, N14773, N12029, N20389);
not NOT1 (N21820, N21790);
xor XOR2 (N21821, N21813, N5415);
xor XOR2 (N21822, N21806, N18089);
or OR2 (N21823, N21818, N16173);
or OR3 (N21824, N21811, N9018, N13967);
not NOT1 (N21825, N21812);
not NOT1 (N21826, N21820);
nand NAND2 (N21827, N21823, N15955);
not NOT1 (N21828, N21816);
nand NAND4 (N21829, N21815, N8868, N2024, N6598);
not NOT1 (N21830, N21829);
or OR4 (N21831, N21799, N13693, N10337, N16496);
buf BUF1 (N21832, N21831);
xor XOR2 (N21833, N21828, N11143);
and AND3 (N21834, N21822, N4870, N10940);
buf BUF1 (N21835, N21819);
xor XOR2 (N21836, N21835, N18087);
xor XOR2 (N21837, N21832, N8524);
not NOT1 (N21838, N21836);
buf BUF1 (N21839, N21837);
and AND2 (N21840, N21830, N9138);
buf BUF1 (N21841, N21839);
not NOT1 (N21842, N21827);
not NOT1 (N21843, N21825);
or OR4 (N21844, N21826, N9166, N10449, N12790);
nor NOR2 (N21845, N21838, N19567);
and AND4 (N21846, N21842, N12665, N15209, N14464);
xor XOR2 (N21847, N21845, N7657);
buf BUF1 (N21848, N21821);
nand NAND2 (N21849, N21840, N164);
nor NOR2 (N21850, N21824, N9649);
not NOT1 (N21851, N21833);
xor XOR2 (N21852, N21846, N11890);
buf BUF1 (N21853, N21843);
or OR4 (N21854, N21849, N6652, N6130, N7427);
nand NAND4 (N21855, N21847, N10129, N16324, N14473);
nand NAND2 (N21856, N21841, N20381);
nor NOR4 (N21857, N21844, N10939, N11977, N6153);
or OR3 (N21858, N21850, N17843, N5713);
buf BUF1 (N21859, N21855);
or OR3 (N21860, N21853, N15985, N18183);
not NOT1 (N21861, N21852);
nand NAND2 (N21862, N21857, N5602);
or OR3 (N21863, N21859, N14467, N11438);
and AND2 (N21864, N21863, N8812);
and AND3 (N21865, N21864, N4853, N17817);
buf BUF1 (N21866, N21854);
nand NAND2 (N21867, N21848, N9185);
not NOT1 (N21868, N21834);
buf BUF1 (N21869, N21865);
xor XOR2 (N21870, N21867, N5677);
and AND4 (N21871, N21856, N14054, N2453, N6549);
or OR4 (N21872, N21851, N19330, N10274, N5120);
xor XOR2 (N21873, N21868, N4331);
and AND3 (N21874, N21873, N34, N823);
xor XOR2 (N21875, N21874, N9780);
and AND4 (N21876, N21862, N14356, N14662, N15318);
xor XOR2 (N21877, N21869, N10114);
buf BUF1 (N21878, N21877);
nor NOR3 (N21879, N21876, N7805, N17970);
and AND4 (N21880, N21879, N4141, N13278, N14026);
nand NAND2 (N21881, N21870, N3683);
and AND4 (N21882, N21881, N15938, N3299, N16961);
buf BUF1 (N21883, N21861);
xor XOR2 (N21884, N21871, N19021);
nand NAND2 (N21885, N21875, N10041);
nor NOR4 (N21886, N21872, N14655, N14955, N7905);
buf BUF1 (N21887, N21885);
xor XOR2 (N21888, N21883, N11505);
and AND3 (N21889, N21858, N18551, N975);
nor NOR3 (N21890, N21884, N5328, N11841);
nand NAND2 (N21891, N21878, N9167);
buf BUF1 (N21892, N21860);
xor XOR2 (N21893, N21888, N7796);
nor NOR2 (N21894, N21889, N2906);
buf BUF1 (N21895, N21866);
and AND2 (N21896, N21882, N13692);
xor XOR2 (N21897, N21896, N7557);
nor NOR3 (N21898, N21886, N20119, N14077);
buf BUF1 (N21899, N21898);
not NOT1 (N21900, N21899);
nand NAND3 (N21901, N21894, N18813, N16018);
not NOT1 (N21902, N21895);
nor NOR3 (N21903, N21902, N21696, N5562);
buf BUF1 (N21904, N21892);
xor XOR2 (N21905, N21893, N7593);
buf BUF1 (N21906, N21891);
nor NOR3 (N21907, N21905, N15314, N5373);
xor XOR2 (N21908, N21890, N19686);
not NOT1 (N21909, N21907);
not NOT1 (N21910, N21880);
and AND4 (N21911, N21901, N16640, N11562, N10218);
buf BUF1 (N21912, N21904);
and AND3 (N21913, N21900, N16662, N9298);
or OR4 (N21914, N21912, N6340, N13567, N10284);
and AND4 (N21915, N21906, N19151, N17617, N3172);
buf BUF1 (N21916, N21915);
not NOT1 (N21917, N21903);
and AND4 (N21918, N21887, N2484, N6030, N13161);
buf BUF1 (N21919, N21910);
not NOT1 (N21920, N21918);
xor XOR2 (N21921, N21917, N6156);
not NOT1 (N21922, N21909);
nand NAND2 (N21923, N21897, N11332);
or OR2 (N21924, N21908, N18450);
not NOT1 (N21925, N21924);
not NOT1 (N21926, N21911);
nand NAND3 (N21927, N21920, N11253, N16986);
not NOT1 (N21928, N21922);
or OR3 (N21929, N21914, N10114, N3299);
or OR3 (N21930, N21923, N20568, N3268);
not NOT1 (N21931, N21926);
buf BUF1 (N21932, N21913);
xor XOR2 (N21933, N21916, N21173);
nand NAND4 (N21934, N21929, N18505, N17209, N6635);
or OR2 (N21935, N21927, N10662);
not NOT1 (N21936, N21919);
xor XOR2 (N21937, N21925, N14116);
buf BUF1 (N21938, N21921);
nand NAND4 (N21939, N21934, N5390, N13921, N4141);
not NOT1 (N21940, N21928);
not NOT1 (N21941, N21937);
buf BUF1 (N21942, N21933);
xor XOR2 (N21943, N21938, N20352);
nand NAND2 (N21944, N21943, N21499);
nand NAND2 (N21945, N21931, N19158);
nor NOR2 (N21946, N21942, N10246);
and AND3 (N21947, N21939, N15319, N881);
nand NAND3 (N21948, N21947, N5311, N431);
or OR2 (N21949, N21944, N2062);
and AND3 (N21950, N21949, N18275, N9205);
buf BUF1 (N21951, N21941);
xor XOR2 (N21952, N21951, N7757);
and AND4 (N21953, N21936, N16908, N876, N14114);
xor XOR2 (N21954, N21930, N8030);
xor XOR2 (N21955, N21948, N8878);
not NOT1 (N21956, N21954);
nor NOR2 (N21957, N21953, N10800);
or OR4 (N21958, N21932, N3204, N14011, N8926);
and AND4 (N21959, N21957, N9775, N20957, N4492);
and AND2 (N21960, N21940, N4217);
buf BUF1 (N21961, N21960);
nand NAND4 (N21962, N21955, N1808, N18039, N1193);
nand NAND4 (N21963, N21961, N612, N14860, N7639);
or OR2 (N21964, N21963, N14515);
and AND4 (N21965, N21962, N11612, N15743, N9807);
nand NAND3 (N21966, N21965, N206, N19167);
not NOT1 (N21967, N21945);
not NOT1 (N21968, N21935);
and AND3 (N21969, N21956, N4954, N17462);
nand NAND4 (N21970, N21950, N15505, N7320, N3872);
buf BUF1 (N21971, N21967);
nor NOR2 (N21972, N21958, N135);
xor XOR2 (N21973, N21971, N9366);
xor XOR2 (N21974, N21970, N18592);
not NOT1 (N21975, N21952);
not NOT1 (N21976, N21975);
not NOT1 (N21977, N21972);
or OR4 (N21978, N21966, N20817, N4677, N7261);
or OR4 (N21979, N21946, N20051, N6851, N5602);
or OR2 (N21980, N21964, N13840);
not NOT1 (N21981, N21978);
nor NOR2 (N21982, N21969, N10562);
nor NOR4 (N21983, N21976, N4050, N17701, N11178);
not NOT1 (N21984, N21977);
xor XOR2 (N21985, N21968, N3616);
xor XOR2 (N21986, N21959, N17753);
and AND2 (N21987, N21982, N1014);
and AND3 (N21988, N21986, N10318, N6748);
nand NAND2 (N21989, N21988, N20974);
and AND4 (N21990, N21981, N10492, N6541, N5132);
not NOT1 (N21991, N21990);
or OR4 (N21992, N21987, N3925, N12885, N4699);
xor XOR2 (N21993, N21974, N17855);
nor NOR4 (N21994, N21989, N10756, N5893, N5437);
not NOT1 (N21995, N21983);
not NOT1 (N21996, N21979);
nand NAND3 (N21997, N21993, N7434, N13710);
not NOT1 (N21998, N21995);
not NOT1 (N21999, N21973);
xor XOR2 (N22000, N21992, N20244);
or OR2 (N22001, N21991, N5635);
buf BUF1 (N22002, N21985);
buf BUF1 (N22003, N21980);
not NOT1 (N22004, N22001);
and AND2 (N22005, N21999, N15286);
nor NOR2 (N22006, N22005, N17639);
not NOT1 (N22007, N22000);
xor XOR2 (N22008, N22006, N9634);
and AND3 (N22009, N21996, N7058, N4143);
not NOT1 (N22010, N21984);
not NOT1 (N22011, N21997);
xor XOR2 (N22012, N21994, N9292);
nor NOR3 (N22013, N22009, N11301, N4273);
xor XOR2 (N22014, N21998, N16736);
nor NOR2 (N22015, N22011, N8726);
nor NOR2 (N22016, N22010, N21008);
nand NAND3 (N22017, N22008, N949, N11758);
xor XOR2 (N22018, N22015, N16579);
nand NAND2 (N22019, N22003, N6781);
nand NAND4 (N22020, N22004, N3394, N9323, N20423);
or OR3 (N22021, N22020, N21042, N4228);
not NOT1 (N22022, N22018);
not NOT1 (N22023, N22012);
and AND3 (N22024, N22013, N2065, N12183);
nand NAND3 (N22025, N22019, N10331, N16571);
and AND2 (N22026, N22017, N2326);
nand NAND4 (N22027, N22025, N17123, N1548, N18127);
nor NOR3 (N22028, N22026, N10077, N15949);
xor XOR2 (N22029, N22028, N10691);
and AND2 (N22030, N22024, N18124);
buf BUF1 (N22031, N22016);
or OR2 (N22032, N22030, N13895);
nand NAND2 (N22033, N22002, N11623);
nand NAND2 (N22034, N22023, N16895);
xor XOR2 (N22035, N22032, N321);
nor NOR2 (N22036, N22022, N5959);
nor NOR3 (N22037, N22035, N14518, N21860);
buf BUF1 (N22038, N22029);
buf BUF1 (N22039, N22021);
nand NAND4 (N22040, N22038, N17058, N3266, N18713);
not NOT1 (N22041, N22037);
xor XOR2 (N22042, N22007, N18613);
nand NAND2 (N22043, N22031, N13898);
nor NOR3 (N22044, N22033, N17971, N20332);
and AND4 (N22045, N22043, N2424, N9289, N4381);
buf BUF1 (N22046, N22036);
nand NAND4 (N22047, N22034, N14778, N221, N3307);
buf BUF1 (N22048, N22044);
nor NOR3 (N22049, N22042, N6833, N3046);
nand NAND4 (N22050, N22045, N4490, N10929, N1939);
buf BUF1 (N22051, N22039);
nor NOR2 (N22052, N22014, N16273);
nand NAND3 (N22053, N22027, N5822, N16382);
buf BUF1 (N22054, N22047);
and AND4 (N22055, N22041, N18989, N6529, N8984);
xor XOR2 (N22056, N22040, N11489);
buf BUF1 (N22057, N22048);
or OR2 (N22058, N22055, N16453);
xor XOR2 (N22059, N22051, N18545);
nor NOR3 (N22060, N22057, N7589, N9537);
buf BUF1 (N22061, N22058);
and AND3 (N22062, N22050, N2584, N7853);
xor XOR2 (N22063, N22049, N18604);
nand NAND2 (N22064, N22059, N20436);
buf BUF1 (N22065, N22054);
xor XOR2 (N22066, N22065, N13019);
xor XOR2 (N22067, N22060, N17493);
nand NAND4 (N22068, N22062, N9672, N18935, N8765);
and AND2 (N22069, N22046, N3821);
xor XOR2 (N22070, N22068, N9855);
nor NOR4 (N22071, N22061, N18802, N11926, N17250);
xor XOR2 (N22072, N22063, N4679);
not NOT1 (N22073, N22069);
nor NOR2 (N22074, N22053, N7854);
and AND3 (N22075, N22072, N12140, N1945);
not NOT1 (N22076, N22066);
nor NOR3 (N22077, N22052, N9841, N18816);
nand NAND4 (N22078, N22074, N9007, N4114, N18213);
nand NAND4 (N22079, N22071, N19673, N3950, N16571);
and AND3 (N22080, N22064, N19417, N4273);
nand NAND3 (N22081, N22070, N4955, N18400);
nor NOR3 (N22082, N22056, N5527, N11858);
nor NOR3 (N22083, N22073, N10703, N11070);
not NOT1 (N22084, N22083);
or OR3 (N22085, N22076, N17886, N14193);
and AND3 (N22086, N22082, N11553, N7373);
and AND2 (N22087, N22084, N9178);
and AND3 (N22088, N22087, N1113, N11736);
or OR2 (N22089, N22075, N5618);
nand NAND3 (N22090, N22067, N13736, N4280);
nand NAND4 (N22091, N22085, N15760, N789, N6047);
buf BUF1 (N22092, N22091);
buf BUF1 (N22093, N22090);
xor XOR2 (N22094, N22077, N12893);
buf BUF1 (N22095, N22093);
nand NAND2 (N22096, N22092, N7700);
xor XOR2 (N22097, N22089, N14781);
not NOT1 (N22098, N22097);
xor XOR2 (N22099, N22095, N9782);
xor XOR2 (N22100, N22080, N161);
xor XOR2 (N22101, N22088, N8247);
and AND4 (N22102, N22096, N8934, N14084, N6709);
nor NOR4 (N22103, N22079, N14387, N12798, N9936);
or OR3 (N22104, N22103, N6075, N6231);
xor XOR2 (N22105, N22100, N1679);
nor NOR4 (N22106, N22099, N11996, N3592, N17199);
or OR4 (N22107, N22102, N17984, N3209, N19007);
not NOT1 (N22108, N22107);
nor NOR4 (N22109, N22081, N9978, N5551, N12588);
and AND3 (N22110, N22105, N17035, N10466);
or OR4 (N22111, N22109, N10552, N14627, N10620);
nor NOR4 (N22112, N22094, N5334, N16598, N2395);
or OR3 (N22113, N22078, N19398, N11059);
nand NAND2 (N22114, N22106, N4775);
not NOT1 (N22115, N22086);
nor NOR2 (N22116, N22110, N18081);
nor NOR4 (N22117, N22108, N13196, N16315, N14301);
nand NAND3 (N22118, N22117, N18885, N15827);
and AND3 (N22119, N22118, N929, N2705);
not NOT1 (N22120, N22101);
not NOT1 (N22121, N22111);
or OR2 (N22122, N22112, N8);
not NOT1 (N22123, N22104);
not NOT1 (N22124, N22122);
xor XOR2 (N22125, N22123, N7163);
nor NOR2 (N22126, N22121, N18515);
not NOT1 (N22127, N22116);
nor NOR4 (N22128, N22126, N3917, N5571, N11585);
not NOT1 (N22129, N22125);
buf BUF1 (N22130, N22124);
buf BUF1 (N22131, N22120);
nand NAND2 (N22132, N22113, N18897);
and AND4 (N22133, N22127, N4715, N1139, N8281);
and AND2 (N22134, N22132, N10789);
and AND2 (N22135, N22133, N5538);
xor XOR2 (N22136, N22115, N17631);
buf BUF1 (N22137, N22130);
nor NOR4 (N22138, N22131, N19702, N7180, N13727);
and AND2 (N22139, N22114, N4296);
buf BUF1 (N22140, N22136);
nand NAND2 (N22141, N22137, N18343);
not NOT1 (N22142, N22128);
and AND2 (N22143, N22119, N4807);
nor NOR2 (N22144, N22140, N1106);
nand NAND4 (N22145, N22098, N1349, N7939, N17031);
nor NOR4 (N22146, N22144, N3497, N9312, N5973);
buf BUF1 (N22147, N22145);
and AND4 (N22148, N22138, N4601, N21201, N1401);
and AND4 (N22149, N22134, N4320, N17299, N2314);
or OR4 (N22150, N22148, N11220, N7409, N21843);
xor XOR2 (N22151, N22141, N13351);
xor XOR2 (N22152, N22139, N21133);
not NOT1 (N22153, N22146);
or OR4 (N22154, N22147, N2861, N20824, N14381);
nor NOR4 (N22155, N22143, N3889, N11653, N21073);
nand NAND2 (N22156, N22129, N16450);
not NOT1 (N22157, N22152);
or OR2 (N22158, N22151, N17813);
xor XOR2 (N22159, N22156, N2831);
nand NAND3 (N22160, N22149, N11314, N14792);
xor XOR2 (N22161, N22135, N10833);
nand NAND3 (N22162, N22158, N3818, N20214);
and AND2 (N22163, N22155, N11799);
xor XOR2 (N22164, N22163, N21545);
nand NAND3 (N22165, N22164, N13324, N9453);
buf BUF1 (N22166, N22150);
xor XOR2 (N22167, N22153, N8863);
or OR3 (N22168, N22159, N1851, N8046);
or OR2 (N22169, N22157, N22100);
nand NAND4 (N22170, N22165, N18813, N9688, N3755);
or OR4 (N22171, N22142, N21966, N14890, N11110);
xor XOR2 (N22172, N22166, N13819);
not NOT1 (N22173, N22172);
nor NOR3 (N22174, N22173, N2232, N17688);
or OR4 (N22175, N22168, N19612, N13809, N19677);
or OR2 (N22176, N22169, N6274);
xor XOR2 (N22177, N22161, N12315);
nor NOR3 (N22178, N22170, N17942, N15263);
and AND4 (N22179, N22160, N21807, N19588, N19527);
buf BUF1 (N22180, N22177);
xor XOR2 (N22181, N22167, N3124);
and AND3 (N22182, N22178, N11197, N5857);
nor NOR2 (N22183, N22174, N4233);
and AND3 (N22184, N22181, N4197, N13646);
or OR3 (N22185, N22179, N10875, N13578);
buf BUF1 (N22186, N22183);
or OR4 (N22187, N22175, N4448, N8224, N1057);
nand NAND4 (N22188, N22154, N16921, N9573, N4113);
xor XOR2 (N22189, N22176, N2724);
or OR3 (N22190, N22180, N21353, N15137);
or OR4 (N22191, N22190, N13480, N9243, N15601);
xor XOR2 (N22192, N22191, N9230);
xor XOR2 (N22193, N22188, N2369);
and AND3 (N22194, N22184, N2266, N20132);
buf BUF1 (N22195, N22192);
and AND2 (N22196, N22195, N5681);
nor NOR4 (N22197, N22189, N14907, N15931, N22040);
nand NAND2 (N22198, N22196, N5966);
buf BUF1 (N22199, N22193);
or OR2 (N22200, N22162, N11932);
nand NAND3 (N22201, N22200, N9221, N2988);
xor XOR2 (N22202, N22199, N8712);
or OR3 (N22203, N22197, N18377, N18639);
or OR2 (N22204, N22203, N14733);
xor XOR2 (N22205, N22198, N20749);
xor XOR2 (N22206, N22205, N6750);
nor NOR3 (N22207, N22201, N19536, N17007);
nand NAND3 (N22208, N22206, N21747, N14236);
nor NOR2 (N22209, N22187, N22106);
not NOT1 (N22210, N22207);
nand NAND3 (N22211, N22204, N19548, N17648);
xor XOR2 (N22212, N22194, N3591);
or OR4 (N22213, N22186, N14062, N20020, N9319);
or OR3 (N22214, N22210, N2515, N8609);
nor NOR4 (N22215, N22182, N8097, N9410, N4543);
buf BUF1 (N22216, N22208);
buf BUF1 (N22217, N22185);
or OR3 (N22218, N22217, N6096, N7652);
nor NOR2 (N22219, N22202, N8193);
nand NAND4 (N22220, N22212, N8120, N8500, N7034);
nor NOR4 (N22221, N22171, N11269, N19095, N15773);
xor XOR2 (N22222, N22209, N1428);
not NOT1 (N22223, N22216);
nand NAND3 (N22224, N22220, N5785, N6405);
nor NOR4 (N22225, N22218, N3844, N17341, N3673);
or OR4 (N22226, N22214, N17275, N11861, N6892);
and AND2 (N22227, N22224, N12778);
not NOT1 (N22228, N22215);
nand NAND2 (N22229, N22226, N13695);
not NOT1 (N22230, N22227);
not NOT1 (N22231, N22223);
nand NAND4 (N22232, N22230, N8574, N9917, N20761);
nor NOR2 (N22233, N22231, N1293);
not NOT1 (N22234, N22228);
and AND3 (N22235, N22221, N2210, N11922);
buf BUF1 (N22236, N22232);
xor XOR2 (N22237, N22229, N2451);
or OR2 (N22238, N22213, N9493);
nor NOR2 (N22239, N22211, N7186);
buf BUF1 (N22240, N22222);
and AND2 (N22241, N22235, N22053);
nand NAND3 (N22242, N22241, N8510, N20190);
buf BUF1 (N22243, N22236);
nor NOR2 (N22244, N22225, N19826);
nand NAND2 (N22245, N22242, N21678);
or OR2 (N22246, N22243, N10151);
or OR3 (N22247, N22234, N7681, N10338);
not NOT1 (N22248, N22247);
nand NAND4 (N22249, N22239, N3154, N14832, N1755);
and AND3 (N22250, N22238, N4527, N18554);
buf BUF1 (N22251, N22249);
nand NAND4 (N22252, N22244, N1019, N1379, N2014);
not NOT1 (N22253, N22219);
and AND3 (N22254, N22237, N5887, N10834);
nand NAND4 (N22255, N22245, N4124, N7120, N15878);
nor NOR3 (N22256, N22253, N16895, N2674);
buf BUF1 (N22257, N22233);
and AND2 (N22258, N22248, N20540);
buf BUF1 (N22259, N22257);
buf BUF1 (N22260, N22252);
nor NOR2 (N22261, N22258, N15221);
or OR2 (N22262, N22256, N14638);
xor XOR2 (N22263, N22255, N16203);
and AND2 (N22264, N22250, N27);
buf BUF1 (N22265, N22259);
not NOT1 (N22266, N22261);
not NOT1 (N22267, N22260);
buf BUF1 (N22268, N22240);
nand NAND3 (N22269, N22268, N1982, N17071);
nor NOR2 (N22270, N22246, N14605);
nor NOR3 (N22271, N22264, N13748, N15811);
and AND3 (N22272, N22270, N18165, N1106);
buf BUF1 (N22273, N22266);
xor XOR2 (N22274, N22254, N9830);
nor NOR2 (N22275, N22272, N17363);
buf BUF1 (N22276, N22265);
nand NAND3 (N22277, N22275, N12983, N173);
nand NAND3 (N22278, N22273, N10265, N9584);
nor NOR4 (N22279, N22251, N21789, N11242, N8590);
nor NOR2 (N22280, N22278, N6483);
or OR3 (N22281, N22277, N18925, N20252);
xor XOR2 (N22282, N22281, N19472);
nor NOR2 (N22283, N22269, N10637);
not NOT1 (N22284, N22282);
buf BUF1 (N22285, N22262);
and AND3 (N22286, N22276, N10311, N6220);
nor NOR2 (N22287, N22274, N21438);
or OR3 (N22288, N22267, N18969, N20544);
or OR2 (N22289, N22279, N13703);
and AND2 (N22290, N22283, N3888);
nand NAND2 (N22291, N22263, N6684);
nand NAND4 (N22292, N22287, N9167, N13801, N7585);
not NOT1 (N22293, N22284);
buf BUF1 (N22294, N22288);
nor NOR4 (N22295, N22271, N10920, N9859, N17236);
and AND2 (N22296, N22286, N4476);
buf BUF1 (N22297, N22293);
nor NOR4 (N22298, N22296, N18841, N607, N427);
buf BUF1 (N22299, N22292);
nor NOR3 (N22300, N22291, N7889, N2465);
not NOT1 (N22301, N22285);
xor XOR2 (N22302, N22301, N4195);
and AND4 (N22303, N22295, N173, N5423, N10461);
buf BUF1 (N22304, N22294);
or OR2 (N22305, N22297, N19985);
xor XOR2 (N22306, N22304, N3633);
or OR2 (N22307, N22290, N18350);
or OR3 (N22308, N22305, N21659, N9261);
xor XOR2 (N22309, N22308, N7663);
or OR4 (N22310, N22306, N21221, N7797, N1156);
and AND3 (N22311, N22302, N9988, N13827);
nor NOR2 (N22312, N22310, N13500);
buf BUF1 (N22313, N22312);
xor XOR2 (N22314, N22313, N11099);
and AND2 (N22315, N22289, N581);
and AND4 (N22316, N22303, N3223, N19653, N3668);
xor XOR2 (N22317, N22309, N1093);
or OR4 (N22318, N22315, N7921, N11910, N12400);
nand NAND3 (N22319, N22300, N20428, N3733);
and AND4 (N22320, N22319, N14649, N20718, N20457);
xor XOR2 (N22321, N22311, N13878);
nor NOR3 (N22322, N22320, N1298, N6809);
nor NOR2 (N22323, N22307, N10653);
and AND3 (N22324, N22299, N3816, N17091);
not NOT1 (N22325, N22280);
and AND3 (N22326, N22317, N7541, N7021);
xor XOR2 (N22327, N22314, N2725);
not NOT1 (N22328, N22325);
nand NAND3 (N22329, N22322, N15496, N8691);
not NOT1 (N22330, N22326);
or OR3 (N22331, N22324, N16110, N2100);
nand NAND3 (N22332, N22321, N21469, N526);
xor XOR2 (N22333, N22323, N3648);
buf BUF1 (N22334, N22316);
and AND3 (N22335, N22327, N738, N14067);
buf BUF1 (N22336, N22332);
nor NOR3 (N22337, N22318, N8706, N6859);
and AND4 (N22338, N22336, N18804, N19311, N16514);
nor NOR2 (N22339, N22328, N18559);
nand NAND4 (N22340, N22331, N21881, N13427, N12427);
buf BUF1 (N22341, N22333);
buf BUF1 (N22342, N22340);
and AND4 (N22343, N22339, N20947, N19467, N8041);
not NOT1 (N22344, N22334);
and AND3 (N22345, N22342, N17133, N18621);
not NOT1 (N22346, N22345);
and AND2 (N22347, N22337, N14154);
nor NOR4 (N22348, N22330, N19195, N2932, N4644);
buf BUF1 (N22349, N22343);
or OR2 (N22350, N22341, N2672);
nor NOR4 (N22351, N22344, N2678, N4213, N16077);
buf BUF1 (N22352, N22347);
and AND3 (N22353, N22348, N5018, N9241);
buf BUF1 (N22354, N22349);
buf BUF1 (N22355, N22338);
xor XOR2 (N22356, N22353, N5686);
not NOT1 (N22357, N22350);
not NOT1 (N22358, N22355);
not NOT1 (N22359, N22356);
buf BUF1 (N22360, N22359);
buf BUF1 (N22361, N22360);
or OR4 (N22362, N22346, N11241, N2216, N1994);
nand NAND2 (N22363, N22298, N10886);
buf BUF1 (N22364, N22362);
xor XOR2 (N22365, N22358, N3381);
not NOT1 (N22366, N22363);
xor XOR2 (N22367, N22351, N17021);
nor NOR2 (N22368, N22357, N20473);
xor XOR2 (N22369, N22329, N3810);
nor NOR3 (N22370, N22367, N21726, N4012);
nand NAND3 (N22371, N22364, N9754, N5911);
and AND2 (N22372, N22371, N20218);
nor NOR2 (N22373, N22354, N13738);
xor XOR2 (N22374, N22361, N8174);
not NOT1 (N22375, N22365);
or OR4 (N22376, N22374, N14558, N6964, N11749);
xor XOR2 (N22377, N22372, N20177);
buf BUF1 (N22378, N22373);
nand NAND2 (N22379, N22378, N13516);
and AND4 (N22380, N22375, N7913, N6218, N11943);
and AND3 (N22381, N22335, N20808, N18558);
or OR2 (N22382, N22379, N16488);
buf BUF1 (N22383, N22369);
nand NAND2 (N22384, N22382, N13584);
nand NAND3 (N22385, N22381, N2005, N20813);
nor NOR4 (N22386, N22352, N8571, N8258, N16313);
buf BUF1 (N22387, N22368);
nor NOR2 (N22388, N22387, N18617);
and AND2 (N22389, N22376, N15576);
nand NAND3 (N22390, N22377, N6664, N18728);
nor NOR4 (N22391, N22388, N8265, N13867, N18827);
nor NOR3 (N22392, N22390, N5747, N17011);
nor NOR4 (N22393, N22386, N2880, N74, N8434);
xor XOR2 (N22394, N22389, N18721);
buf BUF1 (N22395, N22383);
and AND4 (N22396, N22370, N19096, N15563, N7454);
buf BUF1 (N22397, N22392);
xor XOR2 (N22398, N22391, N2020);
nand NAND4 (N22399, N22397, N7243, N17564, N17915);
nand NAND3 (N22400, N22384, N8380, N8657);
nor NOR3 (N22401, N22393, N4386, N15291);
nand NAND4 (N22402, N22398, N20171, N4688, N819);
nor NOR4 (N22403, N22385, N10134, N16458, N2693);
buf BUF1 (N22404, N22402);
and AND4 (N22405, N22395, N15969, N15418, N20607);
and AND4 (N22406, N22403, N1358, N2617, N3104);
not NOT1 (N22407, N22401);
not NOT1 (N22408, N22405);
buf BUF1 (N22409, N22408);
and AND2 (N22410, N22399, N18572);
nor NOR3 (N22411, N22366, N14898, N15304);
or OR2 (N22412, N22406, N6125);
buf BUF1 (N22413, N22407);
or OR4 (N22414, N22409, N11452, N7722, N3358);
xor XOR2 (N22415, N22404, N18506);
and AND2 (N22416, N22410, N15134);
nor NOR2 (N22417, N22411, N6687);
nand NAND2 (N22418, N22413, N9852);
buf BUF1 (N22419, N22412);
and AND3 (N22420, N22416, N8119, N6339);
or OR3 (N22421, N22419, N12571, N16612);
and AND2 (N22422, N22394, N19656);
or OR3 (N22423, N22415, N10161, N16965);
not NOT1 (N22424, N22396);
or OR2 (N22425, N22400, N20719);
or OR4 (N22426, N22417, N2422, N12995, N13058);
not NOT1 (N22427, N22420);
not NOT1 (N22428, N22414);
not NOT1 (N22429, N22425);
and AND4 (N22430, N22421, N7757, N1560, N12421);
or OR4 (N22431, N22428, N10159, N6707, N11307);
buf BUF1 (N22432, N22427);
or OR4 (N22433, N22430, N17392, N19784, N7140);
nand NAND2 (N22434, N22380, N1196);
nor NOR2 (N22435, N22426, N4797);
buf BUF1 (N22436, N22434);
xor XOR2 (N22437, N22436, N19102);
or OR4 (N22438, N22432, N15798, N8191, N2095);
or OR4 (N22439, N22433, N22132, N12684, N14269);
xor XOR2 (N22440, N22438, N14855);
and AND4 (N22441, N22424, N2480, N1459, N614);
and AND4 (N22442, N22418, N10215, N18220, N233);
and AND2 (N22443, N22422, N514);
and AND4 (N22444, N22443, N12232, N11980, N3496);
buf BUF1 (N22445, N22439);
nand NAND4 (N22446, N22442, N16921, N5835, N18398);
nand NAND4 (N22447, N22444, N18947, N3069, N7687);
or OR2 (N22448, N22441, N10162);
or OR3 (N22449, N22446, N15312, N2552);
not NOT1 (N22450, N22447);
xor XOR2 (N22451, N22440, N15096);
and AND2 (N22452, N22437, N18469);
not NOT1 (N22453, N22451);
nor NOR3 (N22454, N22423, N4115, N2848);
xor XOR2 (N22455, N22429, N2756);
and AND3 (N22456, N22450, N19788, N18057);
buf BUF1 (N22457, N22448);
buf BUF1 (N22458, N22455);
not NOT1 (N22459, N22454);
and AND3 (N22460, N22457, N8573, N13396);
buf BUF1 (N22461, N22435);
nand NAND3 (N22462, N22458, N19899, N7157);
not NOT1 (N22463, N22431);
or OR2 (N22464, N22456, N8224);
not NOT1 (N22465, N22460);
not NOT1 (N22466, N22453);
nor NOR3 (N22467, N22452, N55, N10264);
xor XOR2 (N22468, N22445, N15223);
nand NAND4 (N22469, N22467, N5515, N8995, N21347);
and AND3 (N22470, N22461, N6552, N3213);
or OR2 (N22471, N22449, N18861);
nor NOR4 (N22472, N22470, N20759, N20885, N9857);
or OR4 (N22473, N22466, N19063, N4178, N13072);
xor XOR2 (N22474, N22472, N698);
and AND3 (N22475, N22469, N10153, N20054);
or OR2 (N22476, N22474, N7014);
xor XOR2 (N22477, N22473, N13249);
nand NAND3 (N22478, N22459, N18615, N5160);
xor XOR2 (N22479, N22462, N12025);
not NOT1 (N22480, N22477);
buf BUF1 (N22481, N22476);
or OR2 (N22482, N22475, N426);
or OR2 (N22483, N22463, N2969);
not NOT1 (N22484, N22471);
and AND2 (N22485, N22479, N18517);
buf BUF1 (N22486, N22468);
and AND4 (N22487, N22486, N20478, N15616, N9346);
nand NAND2 (N22488, N22484, N6849);
xor XOR2 (N22489, N22483, N17996);
xor XOR2 (N22490, N22480, N5675);
or OR3 (N22491, N22482, N1613, N19536);
nand NAND3 (N22492, N22489, N18018, N2400);
xor XOR2 (N22493, N22488, N3517);
not NOT1 (N22494, N22481);
xor XOR2 (N22495, N22492, N16527);
or OR2 (N22496, N22478, N18836);
not NOT1 (N22497, N22496);
nor NOR2 (N22498, N22490, N9617);
nor NOR3 (N22499, N22487, N18677, N21239);
xor XOR2 (N22500, N22498, N10773);
or OR2 (N22501, N22495, N12196);
xor XOR2 (N22502, N22491, N5536);
xor XOR2 (N22503, N22493, N12166);
nand NAND2 (N22504, N22502, N3625);
not NOT1 (N22505, N22497);
xor XOR2 (N22506, N22494, N5724);
and AND2 (N22507, N22499, N19458);
or OR2 (N22508, N22464, N12571);
and AND2 (N22509, N22508, N5168);
or OR3 (N22510, N22485, N11230, N13466);
or OR3 (N22511, N22510, N11208, N16390);
and AND3 (N22512, N22506, N21074, N5400);
not NOT1 (N22513, N22504);
nand NAND2 (N22514, N22465, N15284);
or OR2 (N22515, N22501, N9820);
xor XOR2 (N22516, N22505, N11335);
or OR2 (N22517, N22514, N7427);
or OR3 (N22518, N22509, N3607, N9342);
not NOT1 (N22519, N22503);
not NOT1 (N22520, N22517);
buf BUF1 (N22521, N22500);
nor NOR4 (N22522, N22516, N13998, N13462, N18892);
xor XOR2 (N22523, N22521, N16001);
nand NAND3 (N22524, N22515, N18626, N16963);
and AND2 (N22525, N22512, N21232);
or OR2 (N22526, N22507, N15437);
xor XOR2 (N22527, N22511, N12197);
nor NOR4 (N22528, N22519, N11903, N3696, N756);
or OR4 (N22529, N22513, N2227, N21838, N9634);
or OR4 (N22530, N22520, N3100, N18729, N4420);
nor NOR4 (N22531, N22524, N7712, N12528, N8596);
not NOT1 (N22532, N22526);
nand NAND2 (N22533, N22523, N8690);
and AND3 (N22534, N22531, N18154, N10621);
or OR2 (N22535, N22528, N12487);
buf BUF1 (N22536, N22527);
nor NOR3 (N22537, N22534, N17030, N16089);
and AND2 (N22538, N22530, N6928);
or OR3 (N22539, N22525, N21546, N6524);
buf BUF1 (N22540, N22518);
buf BUF1 (N22541, N22540);
nand NAND4 (N22542, N22539, N18015, N5809, N21196);
xor XOR2 (N22543, N22532, N5363);
xor XOR2 (N22544, N22538, N13062);
or OR3 (N22545, N22536, N2974, N15574);
nor NOR2 (N22546, N22541, N11335);
not NOT1 (N22547, N22542);
and AND4 (N22548, N22529, N667, N12253, N12375);
nor NOR4 (N22549, N22545, N13914, N12576, N16891);
or OR2 (N22550, N22548, N12345);
nor NOR3 (N22551, N22522, N2595, N2902);
buf BUF1 (N22552, N22546);
nand NAND2 (N22553, N22549, N2113);
xor XOR2 (N22554, N22533, N1075);
buf BUF1 (N22555, N22537);
buf BUF1 (N22556, N22552);
nand NAND2 (N22557, N22553, N11590);
nand NAND2 (N22558, N22557, N17866);
not NOT1 (N22559, N22535);
buf BUF1 (N22560, N22556);
xor XOR2 (N22561, N22550, N2682);
nand NAND2 (N22562, N22561, N1407);
or OR2 (N22563, N22555, N9707);
nand NAND3 (N22564, N22554, N5535, N16406);
or OR3 (N22565, N22551, N12153, N19626);
nand NAND3 (N22566, N22543, N2334, N21887);
nand NAND2 (N22567, N22565, N9132);
or OR3 (N22568, N22566, N22293, N10574);
nand NAND2 (N22569, N22562, N2396);
or OR3 (N22570, N22563, N21604, N11179);
buf BUF1 (N22571, N22544);
not NOT1 (N22572, N22571);
and AND4 (N22573, N22567, N11756, N13322, N17821);
buf BUF1 (N22574, N22547);
or OR2 (N22575, N22559, N14955);
or OR3 (N22576, N22572, N7522, N9240);
or OR3 (N22577, N22560, N6632, N18111);
nor NOR4 (N22578, N22575, N997, N9661, N14282);
nand NAND3 (N22579, N22564, N9437, N6167);
xor XOR2 (N22580, N22579, N20546);
xor XOR2 (N22581, N22569, N6491);
and AND4 (N22582, N22577, N1481, N22076, N21891);
and AND4 (N22583, N22582, N17827, N18674, N4051);
nand NAND4 (N22584, N22574, N10456, N7171, N12637);
nor NOR3 (N22585, N22580, N18174, N4691);
and AND3 (N22586, N22585, N15651, N19827);
nor NOR3 (N22587, N22576, N10020, N1348);
buf BUF1 (N22588, N22586);
nand NAND2 (N22589, N22568, N9886);
and AND2 (N22590, N22589, N8194);
buf BUF1 (N22591, N22558);
not NOT1 (N22592, N22583);
and AND3 (N22593, N22587, N17469, N18242);
xor XOR2 (N22594, N22570, N18645);
xor XOR2 (N22595, N22573, N5755);
or OR3 (N22596, N22591, N16635, N5685);
and AND4 (N22597, N22581, N21065, N2758, N5639);
nor NOR2 (N22598, N22597, N15161);
xor XOR2 (N22599, N22596, N22405);
buf BUF1 (N22600, N22592);
buf BUF1 (N22601, N22600);
nor NOR3 (N22602, N22590, N17351, N2647);
nor NOR2 (N22603, N22593, N22458);
xor XOR2 (N22604, N22584, N15882);
xor XOR2 (N22605, N22595, N5623);
buf BUF1 (N22606, N22588);
xor XOR2 (N22607, N22604, N14089);
not NOT1 (N22608, N22598);
and AND3 (N22609, N22605, N15347, N2974);
or OR2 (N22610, N22603, N21979);
or OR2 (N22611, N22578, N14332);
not NOT1 (N22612, N22606);
nand NAND4 (N22613, N22610, N9645, N3593, N8308);
or OR3 (N22614, N22608, N16954, N5846);
nand NAND2 (N22615, N22594, N17823);
and AND4 (N22616, N22611, N4270, N3139, N1687);
nand NAND3 (N22617, N22599, N2555, N18167);
and AND3 (N22618, N22607, N6518, N5269);
nor NOR4 (N22619, N22615, N5665, N18747, N16666);
not NOT1 (N22620, N22614);
or OR3 (N22621, N22620, N3442, N705);
not NOT1 (N22622, N22609);
nand NAND2 (N22623, N22618, N15553);
not NOT1 (N22624, N22617);
xor XOR2 (N22625, N22619, N14626);
not NOT1 (N22626, N22602);
or OR3 (N22627, N22612, N2575, N14490);
not NOT1 (N22628, N22623);
or OR2 (N22629, N22626, N3889);
and AND3 (N22630, N22624, N6504, N1607);
xor XOR2 (N22631, N22628, N17683);
nand NAND3 (N22632, N22630, N17212, N3177);
nor NOR4 (N22633, N22625, N13622, N14999, N9754);
buf BUF1 (N22634, N22622);
nor NOR3 (N22635, N22627, N5594, N4378);
buf BUF1 (N22636, N22621);
and AND2 (N22637, N22633, N11359);
xor XOR2 (N22638, N22631, N12295);
buf BUF1 (N22639, N22637);
buf BUF1 (N22640, N22638);
nor NOR2 (N22641, N22639, N15033);
not NOT1 (N22642, N22616);
and AND3 (N22643, N22635, N19965, N21706);
or OR3 (N22644, N22642, N16156, N19580);
nand NAND3 (N22645, N22636, N10341, N10887);
buf BUF1 (N22646, N22632);
not NOT1 (N22647, N22641);
and AND2 (N22648, N22645, N16628);
xor XOR2 (N22649, N22613, N9366);
or OR4 (N22650, N22644, N20365, N12690, N12625);
and AND2 (N22651, N22640, N9251);
and AND3 (N22652, N22649, N10985, N13248);
not NOT1 (N22653, N22647);
and AND2 (N22654, N22601, N22173);
xor XOR2 (N22655, N22652, N16401);
or OR2 (N22656, N22634, N3074);
or OR4 (N22657, N22655, N11884, N161, N2742);
xor XOR2 (N22658, N22629, N5959);
or OR2 (N22659, N22651, N618);
nand NAND2 (N22660, N22643, N9234);
nor NOR4 (N22661, N22653, N16107, N18696, N22156);
or OR4 (N22662, N22654, N12028, N9125, N19839);
buf BUF1 (N22663, N22660);
nand NAND2 (N22664, N22659, N20658);
and AND2 (N22665, N22658, N1782);
buf BUF1 (N22666, N22665);
nor NOR3 (N22667, N22661, N10033, N17845);
buf BUF1 (N22668, N22648);
not NOT1 (N22669, N22662);
buf BUF1 (N22670, N22664);
xor XOR2 (N22671, N22663, N13358);
not NOT1 (N22672, N22667);
xor XOR2 (N22673, N22672, N19126);
or OR3 (N22674, N22669, N11434, N7004);
buf BUF1 (N22675, N22650);
and AND3 (N22676, N22674, N20859, N10927);
and AND4 (N22677, N22673, N14499, N6066, N5921);
and AND2 (N22678, N22677, N1712);
and AND2 (N22679, N22670, N13895);
or OR2 (N22680, N22656, N7602);
not NOT1 (N22681, N22668);
xor XOR2 (N22682, N22657, N21977);
not NOT1 (N22683, N22681);
and AND2 (N22684, N22646, N55);
xor XOR2 (N22685, N22683, N7785);
not NOT1 (N22686, N22679);
buf BUF1 (N22687, N22666);
nor NOR2 (N22688, N22686, N12930);
nor NOR3 (N22689, N22675, N1744, N7068);
or OR2 (N22690, N22685, N193);
xor XOR2 (N22691, N22690, N1481);
and AND3 (N22692, N22691, N16376, N21926);
nand NAND3 (N22693, N22688, N3632, N15018);
not NOT1 (N22694, N22689);
xor XOR2 (N22695, N22694, N11220);
not NOT1 (N22696, N22671);
and AND3 (N22697, N22693, N13197, N4842);
xor XOR2 (N22698, N22678, N22205);
or OR3 (N22699, N22696, N3209, N4586);
or OR2 (N22700, N22698, N8284);
not NOT1 (N22701, N22684);
buf BUF1 (N22702, N22699);
not NOT1 (N22703, N22700);
not NOT1 (N22704, N22682);
or OR3 (N22705, N22703, N666, N5299);
nand NAND2 (N22706, N22705, N1163);
not NOT1 (N22707, N22706);
buf BUF1 (N22708, N22707);
or OR3 (N22709, N22695, N12948, N20736);
and AND4 (N22710, N22676, N8174, N4187, N7434);
xor XOR2 (N22711, N22710, N10909);
buf BUF1 (N22712, N22711);
not NOT1 (N22713, N22702);
not NOT1 (N22714, N22713);
nand NAND2 (N22715, N22697, N14054);
xor XOR2 (N22716, N22701, N19935);
xor XOR2 (N22717, N22687, N7969);
xor XOR2 (N22718, N22692, N9401);
nor NOR2 (N22719, N22715, N6616);
or OR4 (N22720, N22709, N13956, N18893, N13827);
or OR3 (N22721, N22718, N20869, N5418);
and AND3 (N22722, N22708, N17384, N9754);
or OR4 (N22723, N22712, N247, N1539, N8537);
xor XOR2 (N22724, N22723, N12952);
buf BUF1 (N22725, N22717);
not NOT1 (N22726, N22722);
buf BUF1 (N22727, N22680);
or OR2 (N22728, N22726, N4327);
or OR2 (N22729, N22714, N11424);
nor NOR4 (N22730, N22724, N2376, N9533, N19273);
or OR4 (N22731, N22716, N11107, N19094, N5284);
or OR4 (N22732, N22719, N19787, N1781, N13030);
xor XOR2 (N22733, N22729, N11592);
xor XOR2 (N22734, N22725, N11775);
nor NOR4 (N22735, N22731, N19329, N20872, N7820);
not NOT1 (N22736, N22730);
and AND3 (N22737, N22736, N1647, N304);
nor NOR3 (N22738, N22728, N5805, N4832);
xor XOR2 (N22739, N22721, N5178);
or OR4 (N22740, N22735, N20862, N14208, N3154);
not NOT1 (N22741, N22737);
and AND4 (N22742, N22740, N12586, N2831, N3707);
and AND4 (N22743, N22733, N13016, N6280, N8660);
and AND3 (N22744, N22704, N9618, N7402);
or OR2 (N22745, N22741, N21640);
buf BUF1 (N22746, N22745);
xor XOR2 (N22747, N22739, N7514);
and AND2 (N22748, N22742, N6933);
and AND3 (N22749, N22732, N10852, N16228);
nor NOR4 (N22750, N22744, N7705, N21930, N12910);
nand NAND2 (N22751, N22747, N7915);
or OR2 (N22752, N22743, N3403);
not NOT1 (N22753, N22720);
xor XOR2 (N22754, N22753, N9754);
not NOT1 (N22755, N22734);
or OR3 (N22756, N22750, N4566, N8647);
not NOT1 (N22757, N22754);
buf BUF1 (N22758, N22755);
and AND2 (N22759, N22758, N2325);
xor XOR2 (N22760, N22748, N14445);
not NOT1 (N22761, N22727);
nor NOR4 (N22762, N22749, N18460, N7766, N14956);
not NOT1 (N22763, N22738);
and AND3 (N22764, N22752, N5194, N3618);
nand NAND2 (N22765, N22763, N2091);
nand NAND3 (N22766, N22761, N7781, N17351);
or OR2 (N22767, N22764, N22700);
buf BUF1 (N22768, N22760);
not NOT1 (N22769, N22766);
nor NOR3 (N22770, N22746, N3014, N11950);
and AND4 (N22771, N22757, N17262, N17117, N12005);
buf BUF1 (N22772, N22756);
nand NAND4 (N22773, N22770, N191, N18779, N413);
xor XOR2 (N22774, N22767, N5622);
xor XOR2 (N22775, N22768, N18117);
not NOT1 (N22776, N22774);
nor NOR4 (N22777, N22765, N10544, N7427, N12986);
buf BUF1 (N22778, N22772);
nand NAND3 (N22779, N22773, N4331, N6484);
not NOT1 (N22780, N22759);
buf BUF1 (N22781, N22778);
nor NOR4 (N22782, N22777, N10334, N1840, N16760);
and AND3 (N22783, N22776, N17774, N3529);
xor XOR2 (N22784, N22771, N13505);
or OR3 (N22785, N22775, N620, N10226);
buf BUF1 (N22786, N22769);
xor XOR2 (N22787, N22784, N13070);
xor XOR2 (N22788, N22786, N21800);
xor XOR2 (N22789, N22780, N6644);
not NOT1 (N22790, N22782);
and AND4 (N22791, N22779, N20730, N2319, N17024);
nand NAND4 (N22792, N22788, N19291, N821, N2547);
xor XOR2 (N22793, N22783, N6412);
and AND4 (N22794, N22762, N3812, N15007, N1778);
not NOT1 (N22795, N22787);
not NOT1 (N22796, N22792);
and AND2 (N22797, N22789, N12463);
buf BUF1 (N22798, N22791);
or OR2 (N22799, N22796, N1573);
not NOT1 (N22800, N22798);
not NOT1 (N22801, N22793);
buf BUF1 (N22802, N22751);
nand NAND3 (N22803, N22795, N20948, N16595);
xor XOR2 (N22804, N22802, N22233);
not NOT1 (N22805, N22801);
not NOT1 (N22806, N22804);
buf BUF1 (N22807, N22805);
or OR4 (N22808, N22797, N6584, N1705, N21428);
xor XOR2 (N22809, N22808, N4006);
nand NAND3 (N22810, N22803, N14175, N15520);
or OR2 (N22811, N22794, N2594);
nand NAND2 (N22812, N22811, N15564);
or OR4 (N22813, N22790, N14529, N13509, N8175);
buf BUF1 (N22814, N22800);
buf BUF1 (N22815, N22814);
or OR4 (N22816, N22785, N4052, N19856, N4700);
and AND2 (N22817, N22799, N5827);
nor NOR4 (N22818, N22810, N14758, N22159, N5148);
and AND3 (N22819, N22818, N4581, N681);
or OR2 (N22820, N22815, N13154);
nor NOR4 (N22821, N22809, N2967, N22255, N5883);
and AND2 (N22822, N22813, N15707);
and AND4 (N22823, N22822, N16998, N6667, N17661);
nand NAND2 (N22824, N22820, N5586);
nor NOR4 (N22825, N22812, N6785, N18676, N9547);
xor XOR2 (N22826, N22821, N20619);
and AND2 (N22827, N22823, N12007);
not NOT1 (N22828, N22827);
and AND3 (N22829, N22806, N16927, N11368);
and AND4 (N22830, N22829, N2018, N6655, N12591);
buf BUF1 (N22831, N22816);
not NOT1 (N22832, N22819);
nor NOR2 (N22833, N22825, N19872);
buf BUF1 (N22834, N22831);
or OR4 (N22835, N22824, N14376, N16467, N2979);
or OR2 (N22836, N22830, N20132);
or OR2 (N22837, N22832, N18960);
or OR3 (N22838, N22807, N5007, N8930);
nand NAND2 (N22839, N22834, N9032);
nand NAND4 (N22840, N22781, N16556, N3601, N10958);
nand NAND3 (N22841, N22836, N19115, N8588);
nand NAND4 (N22842, N22841, N5818, N12740, N12221);
not NOT1 (N22843, N22840);
nor NOR4 (N22844, N22843, N6292, N1404, N9071);
and AND4 (N22845, N22844, N10716, N5899, N16744);
or OR4 (N22846, N22842, N9824, N2079, N18344);
or OR3 (N22847, N22828, N19000, N4010);
or OR3 (N22848, N22837, N8663, N17101);
xor XOR2 (N22849, N22833, N13562);
and AND4 (N22850, N22848, N6433, N8243, N10586);
nor NOR2 (N22851, N22849, N13422);
buf BUF1 (N22852, N22838);
nor NOR4 (N22853, N22845, N14189, N19099, N4658);
nor NOR4 (N22854, N22846, N2906, N21547, N9767);
or OR4 (N22855, N22817, N18461, N390, N1950);
nand NAND4 (N22856, N22854, N4900, N2848, N17124);
nand NAND2 (N22857, N22856, N8598);
xor XOR2 (N22858, N22826, N12015);
buf BUF1 (N22859, N22858);
or OR2 (N22860, N22850, N20249);
nor NOR3 (N22861, N22857, N9046, N15264);
or OR3 (N22862, N22835, N14746, N18471);
not NOT1 (N22863, N22847);
buf BUF1 (N22864, N22863);
buf BUF1 (N22865, N22851);
buf BUF1 (N22866, N22852);
not NOT1 (N22867, N22866);
not NOT1 (N22868, N22864);
nand NAND3 (N22869, N22862, N1717, N9165);
and AND4 (N22870, N22859, N7221, N18764, N16337);
and AND2 (N22871, N22870, N8872);
buf BUF1 (N22872, N22869);
nand NAND3 (N22873, N22853, N12573, N22596);
and AND3 (N22874, N22873, N13877, N16800);
not NOT1 (N22875, N22867);
not NOT1 (N22876, N22855);
not NOT1 (N22877, N22871);
xor XOR2 (N22878, N22865, N20252);
or OR3 (N22879, N22861, N22068, N20668);
xor XOR2 (N22880, N22839, N5879);
buf BUF1 (N22881, N22860);
nand NAND2 (N22882, N22878, N17096);
xor XOR2 (N22883, N22872, N17915);
not NOT1 (N22884, N22881);
buf BUF1 (N22885, N22884);
not NOT1 (N22886, N22880);
xor XOR2 (N22887, N22885, N17651);
buf BUF1 (N22888, N22876);
buf BUF1 (N22889, N22877);
nor NOR3 (N22890, N22868, N11498, N14670);
nand NAND3 (N22891, N22875, N15441, N17317);
nand NAND4 (N22892, N22874, N5670, N8739, N15093);
nand NAND2 (N22893, N22890, N21917);
nand NAND2 (N22894, N22883, N22606);
or OR2 (N22895, N22894, N8428);
buf BUF1 (N22896, N22879);
nor NOR2 (N22897, N22887, N19349);
xor XOR2 (N22898, N22895, N12962);
or OR2 (N22899, N22889, N4569);
buf BUF1 (N22900, N22897);
and AND3 (N22901, N22896, N1681, N14634);
and AND4 (N22902, N22898, N15082, N9091, N22782);
xor XOR2 (N22903, N22901, N5337);
and AND2 (N22904, N22899, N17335);
and AND3 (N22905, N22900, N2188, N3033);
nand NAND3 (N22906, N22891, N22456, N1859);
nand NAND3 (N22907, N22882, N1234, N9457);
not NOT1 (N22908, N22893);
and AND2 (N22909, N22903, N14417);
nand NAND3 (N22910, N22902, N10909, N22595);
nor NOR3 (N22911, N22908, N7968, N13191);
buf BUF1 (N22912, N22907);
nand NAND4 (N22913, N22888, N4301, N1026, N14370);
nand NAND2 (N22914, N22910, N5150);
not NOT1 (N22915, N22909);
xor XOR2 (N22916, N22906, N6570);
not NOT1 (N22917, N22916);
xor XOR2 (N22918, N22912, N15815);
or OR4 (N22919, N22904, N22258, N9594, N6155);
xor XOR2 (N22920, N22886, N5305);
buf BUF1 (N22921, N22892);
or OR2 (N22922, N22915, N5681);
or OR4 (N22923, N22919, N11902, N15894, N9914);
and AND2 (N22924, N22914, N19059);
buf BUF1 (N22925, N22923);
not NOT1 (N22926, N22918);
buf BUF1 (N22927, N22926);
nor NOR3 (N22928, N22913, N13632, N9152);
and AND4 (N22929, N22917, N9913, N17997, N22901);
not NOT1 (N22930, N22924);
or OR4 (N22931, N22925, N5609, N20373, N1920);
nand NAND3 (N22932, N22928, N9081, N2755);
xor XOR2 (N22933, N22927, N8075);
buf BUF1 (N22934, N22921);
or OR4 (N22935, N22922, N2427, N2409, N22031);
nand NAND4 (N22936, N22905, N309, N16286, N16504);
not NOT1 (N22937, N22936);
buf BUF1 (N22938, N22935);
xor XOR2 (N22939, N22929, N4396);
buf BUF1 (N22940, N22939);
and AND2 (N22941, N22932, N2763);
or OR3 (N22942, N22938, N13132, N15783);
and AND3 (N22943, N22920, N4051, N10232);
and AND3 (N22944, N22942, N22026, N13629);
buf BUF1 (N22945, N22941);
not NOT1 (N22946, N22911);
not NOT1 (N22947, N22934);
xor XOR2 (N22948, N22943, N22198);
and AND2 (N22949, N22945, N22070);
buf BUF1 (N22950, N22949);
and AND4 (N22951, N22937, N195, N13768, N6921);
not NOT1 (N22952, N22931);
not NOT1 (N22953, N22940);
and AND4 (N22954, N22946, N3542, N3482, N10965);
nor NOR3 (N22955, N22947, N9950, N15082);
and AND3 (N22956, N22952, N14437, N522);
xor XOR2 (N22957, N22948, N582);
and AND2 (N22958, N22944, N22788);
and AND4 (N22959, N22933, N14558, N11310, N12791);
xor XOR2 (N22960, N22959, N21214);
xor XOR2 (N22961, N22956, N21078);
xor XOR2 (N22962, N22960, N3906);
and AND2 (N22963, N22953, N7479);
xor XOR2 (N22964, N22961, N16500);
or OR3 (N22965, N22955, N6989, N17379);
nor NOR3 (N22966, N22965, N12244, N19261);
xor XOR2 (N22967, N22951, N17539);
nand NAND4 (N22968, N22966, N12513, N2997, N12032);
not NOT1 (N22969, N22954);
and AND3 (N22970, N22950, N19971, N4994);
buf BUF1 (N22971, N22970);
nor NOR3 (N22972, N22964, N7884, N21151);
nand NAND4 (N22973, N22962, N1390, N5019, N9203);
xor XOR2 (N22974, N22972, N5360);
xor XOR2 (N22975, N22968, N18586);
nor NOR3 (N22976, N22967, N8910, N4393);
not NOT1 (N22977, N22930);
or OR4 (N22978, N22975, N1202, N6808, N8083);
and AND3 (N22979, N22974, N7866, N1772);
or OR4 (N22980, N22973, N1086, N19985, N10427);
not NOT1 (N22981, N22958);
buf BUF1 (N22982, N22978);
nor NOR2 (N22983, N22976, N10216);
nand NAND2 (N22984, N22982, N20830);
buf BUF1 (N22985, N22969);
xor XOR2 (N22986, N22981, N3841);
buf BUF1 (N22987, N22977);
or OR3 (N22988, N22980, N16035, N14919);
not NOT1 (N22989, N22986);
buf BUF1 (N22990, N22984);
or OR4 (N22991, N22963, N20157, N3200, N21261);
nor NOR3 (N22992, N22988, N4011, N21169);
or OR3 (N22993, N22983, N1359, N18639);
xor XOR2 (N22994, N22985, N3017);
not NOT1 (N22995, N22991);
and AND4 (N22996, N22994, N19185, N18732, N12333);
nand NAND3 (N22997, N22971, N15452, N4277);
xor XOR2 (N22998, N22979, N5087);
nand NAND2 (N22999, N22997, N20301);
buf BUF1 (N23000, N22996);
nor NOR3 (N23001, N22990, N2348, N11769);
or OR2 (N23002, N22992, N13166);
nor NOR3 (N23003, N22999, N17212, N6541);
nand NAND3 (N23004, N22957, N22558, N11385);
or OR3 (N23005, N22995, N8565, N4993);
nor NOR3 (N23006, N22998, N10910, N15605);
nor NOR2 (N23007, N22993, N11141);
not NOT1 (N23008, N23004);
nor NOR4 (N23009, N22989, N19770, N7984, N15405);
or OR3 (N23010, N23003, N1110, N14645);
not NOT1 (N23011, N23001);
xor XOR2 (N23012, N23005, N20118);
nand NAND4 (N23013, N23010, N15663, N18947, N20830);
nor NOR3 (N23014, N22987, N2921, N19738);
or OR4 (N23015, N23012, N20350, N3976, N11421);
buf BUF1 (N23016, N23007);
or OR4 (N23017, N23008, N14591, N20905, N9244);
xor XOR2 (N23018, N23015, N8767);
or OR2 (N23019, N23018, N14946);
nor NOR4 (N23020, N23009, N231, N11494, N6025);
nand NAND3 (N23021, N23017, N13177, N13558);
and AND4 (N23022, N23021, N7973, N8531, N17593);
nand NAND3 (N23023, N23014, N4215, N2275);
or OR3 (N23024, N23013, N8539, N11928);
buf BUF1 (N23025, N23019);
nor NOR3 (N23026, N23000, N5456, N18886);
nand NAND2 (N23027, N23011, N5231);
nand NAND3 (N23028, N23006, N6368, N12855);
xor XOR2 (N23029, N23023, N15460);
or OR3 (N23030, N23028, N18508, N13389);
buf BUF1 (N23031, N23026);
buf BUF1 (N23032, N23002);
not NOT1 (N23033, N23016);
buf BUF1 (N23034, N23020);
nand NAND3 (N23035, N23031, N14138, N5756);
not NOT1 (N23036, N23029);
nor NOR2 (N23037, N23032, N1148);
nor NOR4 (N23038, N23033, N7340, N615, N16893);
nand NAND4 (N23039, N23036, N21785, N11468, N10411);
not NOT1 (N23040, N23038);
buf BUF1 (N23041, N23025);
not NOT1 (N23042, N23035);
and AND4 (N23043, N23027, N21497, N21115, N1391);
nand NAND3 (N23044, N23040, N6657, N20823);
nand NAND2 (N23045, N23042, N12421);
not NOT1 (N23046, N23037);
and AND3 (N23047, N23044, N13576, N3081);
buf BUF1 (N23048, N23039);
buf BUF1 (N23049, N23041);
not NOT1 (N23050, N23047);
xor XOR2 (N23051, N23043, N15715);
buf BUF1 (N23052, N23049);
nand NAND3 (N23053, N23048, N21287, N12877);
buf BUF1 (N23054, N23053);
nor NOR4 (N23055, N23024, N7951, N1085, N6158);
and AND4 (N23056, N23034, N20227, N2806, N2139);
nor NOR2 (N23057, N23055, N19486);
nand NAND3 (N23058, N23051, N5752, N13459);
nand NAND2 (N23059, N23046, N16021);
nor NOR4 (N23060, N23058, N22133, N1590, N19983);
buf BUF1 (N23061, N23056);
or OR3 (N23062, N23022, N17203, N668);
xor XOR2 (N23063, N23050, N12621);
and AND4 (N23064, N23052, N21762, N10082, N9553);
xor XOR2 (N23065, N23061, N22308);
or OR4 (N23066, N23062, N22523, N2329, N3840);
nand NAND3 (N23067, N23066, N19449, N14926);
nor NOR2 (N23068, N23065, N3543);
nor NOR3 (N23069, N23067, N12672, N197);
or OR3 (N23070, N23059, N19566, N11047);
xor XOR2 (N23071, N23054, N20434);
nand NAND2 (N23072, N23068, N9039);
buf BUF1 (N23073, N23057);
buf BUF1 (N23074, N23069);
buf BUF1 (N23075, N23073);
buf BUF1 (N23076, N23075);
nand NAND2 (N23077, N23072, N6683);
buf BUF1 (N23078, N23070);
or OR4 (N23079, N23063, N16655, N8517, N5599);
nand NAND2 (N23080, N23071, N18107);
buf BUF1 (N23081, N23030);
not NOT1 (N23082, N23064);
nand NAND3 (N23083, N23082, N1142, N1640);
or OR4 (N23084, N23078, N2863, N13697, N8142);
nor NOR4 (N23085, N23083, N9639, N12967, N18631);
or OR3 (N23086, N23081, N2305, N14661);
and AND2 (N23087, N23060, N16171);
buf BUF1 (N23088, N23045);
and AND2 (N23089, N23084, N11836);
and AND2 (N23090, N23089, N10569);
nand NAND3 (N23091, N23087, N3735, N20716);
nand NAND2 (N23092, N23088, N23082);
not NOT1 (N23093, N23086);
buf BUF1 (N23094, N23085);
xor XOR2 (N23095, N23074, N916);
and AND3 (N23096, N23094, N21040, N4121);
not NOT1 (N23097, N23076);
nand NAND4 (N23098, N23092, N1103, N13546, N19696);
nand NAND3 (N23099, N23096, N13467, N8521);
nor NOR4 (N23100, N23079, N23008, N9907, N21028);
not NOT1 (N23101, N23080);
nor NOR2 (N23102, N23077, N1598);
buf BUF1 (N23103, N23093);
nand NAND2 (N23104, N23100, N14779);
buf BUF1 (N23105, N23095);
xor XOR2 (N23106, N23097, N4188);
nand NAND2 (N23107, N23102, N13713);
not NOT1 (N23108, N23106);
not NOT1 (N23109, N23103);
nor NOR4 (N23110, N23101, N14826, N20225, N8842);
not NOT1 (N23111, N23098);
buf BUF1 (N23112, N23111);
nand NAND2 (N23113, N23110, N10367);
xor XOR2 (N23114, N23105, N5458);
buf BUF1 (N23115, N23108);
nand NAND4 (N23116, N23112, N15496, N1268, N455);
buf BUF1 (N23117, N23114);
not NOT1 (N23118, N23099);
or OR4 (N23119, N23117, N14272, N18886, N7558);
nand NAND4 (N23120, N23107, N15010, N17244, N16063);
not NOT1 (N23121, N23116);
and AND3 (N23122, N23090, N13312, N11975);
xor XOR2 (N23123, N23120, N19660);
xor XOR2 (N23124, N23121, N7281);
nand NAND3 (N23125, N23104, N11050, N2647);
or OR4 (N23126, N23109, N21231, N8202, N5470);
and AND2 (N23127, N23126, N3919);
and AND3 (N23128, N23125, N19339, N2030);
nor NOR2 (N23129, N23128, N13451);
and AND2 (N23130, N23127, N19215);
xor XOR2 (N23131, N23122, N21297);
nand NAND2 (N23132, N23119, N8646);
buf BUF1 (N23133, N23091);
not NOT1 (N23134, N23133);
and AND4 (N23135, N23134, N17505, N16944, N18361);
nor NOR2 (N23136, N23129, N13822);
buf BUF1 (N23137, N23136);
nand NAND3 (N23138, N23123, N18712, N8108);
not NOT1 (N23139, N23130);
xor XOR2 (N23140, N23132, N16946);
nor NOR2 (N23141, N23139, N16859);
nand NAND2 (N23142, N23141, N13253);
nand NAND3 (N23143, N23138, N924, N2851);
or OR2 (N23144, N23137, N12125);
nor NOR2 (N23145, N23118, N2949);
and AND2 (N23146, N23140, N17319);
xor XOR2 (N23147, N23131, N638);
not NOT1 (N23148, N23144);
and AND2 (N23149, N23145, N740);
nor NOR3 (N23150, N23143, N6768, N20822);
or OR2 (N23151, N23142, N7398);
not NOT1 (N23152, N23150);
or OR4 (N23153, N23115, N19048, N20169, N113);
nor NOR4 (N23154, N23135, N14985, N3354, N5007);
xor XOR2 (N23155, N23149, N18183);
and AND2 (N23156, N23124, N11578);
xor XOR2 (N23157, N23154, N8052);
and AND2 (N23158, N23151, N2012);
nor NOR4 (N23159, N23113, N9324, N19472, N11117);
or OR4 (N23160, N23157, N3026, N5676, N12523);
or OR3 (N23161, N23148, N1023, N12351);
not NOT1 (N23162, N23158);
not NOT1 (N23163, N23146);
or OR3 (N23164, N23161, N17470, N6485);
or OR3 (N23165, N23164, N4013, N4519);
nor NOR2 (N23166, N23163, N11275);
nand NAND4 (N23167, N23153, N18820, N20868, N11991);
and AND2 (N23168, N23147, N20838);
nor NOR2 (N23169, N23162, N21243);
or OR4 (N23170, N23160, N11267, N7215, N17208);
xor XOR2 (N23171, N23159, N12671);
not NOT1 (N23172, N23168);
nand NAND2 (N23173, N23171, N2895);
buf BUF1 (N23174, N23166);
xor XOR2 (N23175, N23173, N4336);
nor NOR3 (N23176, N23174, N13093, N19012);
not NOT1 (N23177, N23155);
nand NAND3 (N23178, N23165, N11909, N3993);
nand NAND2 (N23179, N23170, N10477);
xor XOR2 (N23180, N23179, N8491);
not NOT1 (N23181, N23152);
or OR4 (N23182, N23156, N22303, N2427, N3659);
nor NOR2 (N23183, N23177, N13059);
not NOT1 (N23184, N23183);
nand NAND2 (N23185, N23176, N20974);
nand NAND2 (N23186, N23181, N18798);
and AND3 (N23187, N23169, N6623, N13372);
not NOT1 (N23188, N23180);
or OR3 (N23189, N23167, N2996, N19995);
not NOT1 (N23190, N23178);
xor XOR2 (N23191, N23190, N18998);
xor XOR2 (N23192, N23182, N21781);
xor XOR2 (N23193, N23172, N9585);
nand NAND2 (N23194, N23175, N5990);
xor XOR2 (N23195, N23194, N6676);
nor NOR4 (N23196, N23184, N7253, N264, N4266);
nand NAND2 (N23197, N23188, N6666);
nand NAND4 (N23198, N23192, N14709, N7026, N19898);
xor XOR2 (N23199, N23193, N15644);
and AND4 (N23200, N23191, N8922, N357, N15977);
nor NOR2 (N23201, N23199, N3829);
not NOT1 (N23202, N23187);
xor XOR2 (N23203, N23196, N22016);
or OR2 (N23204, N23202, N19437);
buf BUF1 (N23205, N23198);
xor XOR2 (N23206, N23200, N16383);
nor NOR4 (N23207, N23204, N10421, N11378, N15795);
xor XOR2 (N23208, N23197, N11377);
nor NOR3 (N23209, N23203, N3907, N18064);
not NOT1 (N23210, N23209);
xor XOR2 (N23211, N23207, N22974);
xor XOR2 (N23212, N23201, N12476);
not NOT1 (N23213, N23195);
xor XOR2 (N23214, N23206, N12798);
buf BUF1 (N23215, N23210);
nor NOR4 (N23216, N23215, N20427, N817, N2895);
not NOT1 (N23217, N23212);
nand NAND2 (N23218, N23205, N7016);
and AND2 (N23219, N23214, N5148);
not NOT1 (N23220, N23211);
and AND3 (N23221, N23217, N6308, N11617);
xor XOR2 (N23222, N23185, N1707);
buf BUF1 (N23223, N23220);
or OR4 (N23224, N23219, N3719, N17157, N2101);
buf BUF1 (N23225, N23218);
buf BUF1 (N23226, N23186);
buf BUF1 (N23227, N23208);
xor XOR2 (N23228, N23224, N1204);
and AND3 (N23229, N23225, N9906, N8064);
nand NAND3 (N23230, N23229, N2288, N20037);
and AND4 (N23231, N23216, N3767, N218, N13168);
nand NAND3 (N23232, N23213, N15449, N5162);
nor NOR3 (N23233, N23189, N1696, N10114);
xor XOR2 (N23234, N23227, N5701);
not NOT1 (N23235, N23233);
and AND4 (N23236, N23232, N3214, N12206, N19228);
not NOT1 (N23237, N23236);
nand NAND4 (N23238, N23222, N12604, N14957, N4955);
or OR2 (N23239, N23226, N14515);
or OR3 (N23240, N23237, N7991, N6266);
nor NOR3 (N23241, N23230, N16967, N5425);
not NOT1 (N23242, N23240);
not NOT1 (N23243, N23241);
nor NOR3 (N23244, N23234, N1307, N21253);
buf BUF1 (N23245, N23235);
not NOT1 (N23246, N23242);
not NOT1 (N23247, N23245);
buf BUF1 (N23248, N23238);
xor XOR2 (N23249, N23221, N2347);
or OR4 (N23250, N23249, N18703, N881, N1764);
and AND4 (N23251, N23223, N2576, N6686, N14723);
nor NOR2 (N23252, N23247, N8609);
nor NOR4 (N23253, N23228, N7749, N14774, N10248);
and AND3 (N23254, N23246, N15018, N23215);
nand NAND4 (N23255, N23253, N14979, N7233, N17669);
nor NOR3 (N23256, N23244, N5313, N8895);
nor NOR4 (N23257, N23252, N2597, N2609, N16875);
xor XOR2 (N23258, N23256, N12311);
and AND2 (N23259, N23239, N7697);
xor XOR2 (N23260, N23254, N18452);
or OR2 (N23261, N23258, N7973);
or OR2 (N23262, N23243, N6381);
buf BUF1 (N23263, N23250);
nand NAND4 (N23264, N23251, N22017, N11327, N4168);
nor NOR3 (N23265, N23263, N22211, N10937);
nor NOR4 (N23266, N23264, N8973, N19167, N15496);
buf BUF1 (N23267, N23255);
not NOT1 (N23268, N23257);
xor XOR2 (N23269, N23248, N16656);
nor NOR2 (N23270, N23261, N14382);
buf BUF1 (N23271, N23260);
nand NAND2 (N23272, N23262, N2367);
xor XOR2 (N23273, N23259, N22440);
nor NOR3 (N23274, N23267, N13263, N11234);
nor NOR3 (N23275, N23266, N9894, N17578);
buf BUF1 (N23276, N23269);
nand NAND3 (N23277, N23274, N1263, N21560);
xor XOR2 (N23278, N23273, N9895);
nand NAND4 (N23279, N23268, N17896, N9634, N11543);
nand NAND4 (N23280, N23272, N750, N6943, N12253);
and AND2 (N23281, N23276, N2251);
or OR2 (N23282, N23270, N13272);
xor XOR2 (N23283, N23271, N2193);
not NOT1 (N23284, N23282);
not NOT1 (N23285, N23231);
nand NAND4 (N23286, N23281, N1095, N7670, N9337);
or OR4 (N23287, N23278, N21870, N7555, N8473);
and AND3 (N23288, N23279, N2212, N23176);
xor XOR2 (N23289, N23275, N14623);
nand NAND3 (N23290, N23286, N17341, N18748);
xor XOR2 (N23291, N23284, N11619);
nor NOR4 (N23292, N23289, N13462, N6614, N10909);
not NOT1 (N23293, N23290);
or OR3 (N23294, N23287, N1145, N1390);
buf BUF1 (N23295, N23283);
xor XOR2 (N23296, N23288, N22568);
not NOT1 (N23297, N23277);
or OR2 (N23298, N23265, N13038);
not NOT1 (N23299, N23295);
or OR3 (N23300, N23285, N5151, N19126);
or OR2 (N23301, N23300, N17454);
and AND2 (N23302, N23297, N2641);
nor NOR3 (N23303, N23293, N16668, N21110);
nand NAND3 (N23304, N23296, N8376, N8121);
nand NAND2 (N23305, N23301, N10542);
and AND2 (N23306, N23304, N11774);
or OR4 (N23307, N23298, N4574, N13025, N14055);
nor NOR4 (N23308, N23307, N19223, N7289, N17712);
or OR2 (N23309, N23280, N20820);
and AND2 (N23310, N23292, N9052);
nor NOR3 (N23311, N23291, N2231, N16953);
nand NAND4 (N23312, N23310, N14638, N8745, N22494);
nor NOR3 (N23313, N23306, N4618, N16440);
or OR2 (N23314, N23305, N22158);
nand NAND4 (N23315, N23299, N16868, N14442, N19885);
not NOT1 (N23316, N23312);
xor XOR2 (N23317, N23309, N14241);
nor NOR2 (N23318, N23302, N9604);
buf BUF1 (N23319, N23318);
and AND2 (N23320, N23317, N6528);
not NOT1 (N23321, N23316);
xor XOR2 (N23322, N23313, N15443);
and AND2 (N23323, N23321, N20733);
nand NAND2 (N23324, N23311, N15925);
or OR4 (N23325, N23294, N6878, N21872, N22626);
nand NAND2 (N23326, N23325, N15351);
buf BUF1 (N23327, N23308);
xor XOR2 (N23328, N23314, N667);
or OR4 (N23329, N23326, N21453, N5790, N329);
nor NOR2 (N23330, N23315, N7627);
not NOT1 (N23331, N23324);
or OR2 (N23332, N23331, N22358);
buf BUF1 (N23333, N23332);
nand NAND2 (N23334, N23319, N7948);
or OR2 (N23335, N23322, N7708);
or OR4 (N23336, N23333, N11981, N14468, N4304);
not NOT1 (N23337, N23320);
not NOT1 (N23338, N23303);
not NOT1 (N23339, N23338);
nor NOR2 (N23340, N23323, N6337);
nand NAND2 (N23341, N23328, N432);
buf BUF1 (N23342, N23339);
buf BUF1 (N23343, N23341);
nor NOR3 (N23344, N23337, N16918, N21097);
or OR3 (N23345, N23340, N5785, N5884);
or OR2 (N23346, N23334, N109);
nand NAND3 (N23347, N23345, N13711, N1315);
buf BUF1 (N23348, N23343);
nor NOR3 (N23349, N23330, N9718, N15923);
buf BUF1 (N23350, N23329);
and AND2 (N23351, N23335, N4851);
or OR2 (N23352, N23327, N3853);
buf BUF1 (N23353, N23349);
xor XOR2 (N23354, N23342, N20853);
xor XOR2 (N23355, N23352, N3650);
buf BUF1 (N23356, N23350);
buf BUF1 (N23357, N23353);
or OR2 (N23358, N23356, N3379);
buf BUF1 (N23359, N23346);
and AND2 (N23360, N23348, N22806);
or OR2 (N23361, N23347, N21358);
xor XOR2 (N23362, N23358, N15436);
or OR2 (N23363, N23359, N10437);
nor NOR2 (N23364, N23360, N19766);
xor XOR2 (N23365, N23357, N11739);
nand NAND4 (N23366, N23336, N18779, N14130, N4238);
nand NAND2 (N23367, N23351, N59);
xor XOR2 (N23368, N23365, N20952);
buf BUF1 (N23369, N23362);
and AND2 (N23370, N23355, N342);
nand NAND4 (N23371, N23344, N23344, N10200, N21168);
xor XOR2 (N23372, N23367, N13974);
and AND3 (N23373, N23366, N9534, N12475);
not NOT1 (N23374, N23373);
or OR4 (N23375, N23363, N16711, N12259, N17393);
and AND2 (N23376, N23370, N10670);
nor NOR4 (N23377, N23371, N6056, N18637, N5084);
nor NOR3 (N23378, N23374, N9586, N18402);
nor NOR4 (N23379, N23368, N18866, N20586, N1297);
buf BUF1 (N23380, N23361);
and AND3 (N23381, N23364, N19702, N1961);
nor NOR3 (N23382, N23376, N881, N6502);
and AND3 (N23383, N23378, N22151, N12035);
and AND2 (N23384, N23375, N397);
nor NOR2 (N23385, N23372, N11838);
nand NAND3 (N23386, N23354, N17586, N3692);
or OR3 (N23387, N23369, N1791, N14653);
nand NAND2 (N23388, N23381, N7321);
not NOT1 (N23389, N23388);
or OR2 (N23390, N23383, N4265);
nand NAND4 (N23391, N23377, N6133, N8647, N9944);
nand NAND2 (N23392, N23379, N19715);
or OR3 (N23393, N23385, N17166, N16203);
nand NAND4 (N23394, N23391, N19144, N2337, N18186);
and AND3 (N23395, N23384, N14501, N19207);
or OR4 (N23396, N23392, N11784, N2734, N15540);
buf BUF1 (N23397, N23386);
nor NOR3 (N23398, N23395, N11806, N11622);
nor NOR4 (N23399, N23398, N10530, N23100, N12293);
nor NOR4 (N23400, N23387, N19531, N16374, N22570);
and AND4 (N23401, N23400, N8202, N7614, N8601);
nand NAND2 (N23402, N23396, N12595);
buf BUF1 (N23403, N23399);
nor NOR4 (N23404, N23394, N19129, N7831, N8537);
and AND2 (N23405, N23404, N15774);
not NOT1 (N23406, N23401);
buf BUF1 (N23407, N23389);
xor XOR2 (N23408, N23393, N16407);
buf BUF1 (N23409, N23390);
nor NOR3 (N23410, N23380, N4118, N6426);
xor XOR2 (N23411, N23397, N19566);
nor NOR3 (N23412, N23403, N8952, N22962);
nor NOR4 (N23413, N23405, N9413, N16405, N7277);
nor NOR3 (N23414, N23382, N15538, N1352);
nor NOR2 (N23415, N23407, N2578);
nor NOR4 (N23416, N23402, N23139, N1608, N5032);
or OR3 (N23417, N23409, N10360, N16028);
nand NAND4 (N23418, N23417, N508, N1637, N407);
nand NAND3 (N23419, N23411, N3668, N5699);
buf BUF1 (N23420, N23412);
not NOT1 (N23421, N23416);
xor XOR2 (N23422, N23415, N16876);
or OR3 (N23423, N23410, N19533, N12843);
nor NOR3 (N23424, N23423, N6582, N6225);
nor NOR2 (N23425, N23406, N21898);
and AND4 (N23426, N23414, N11780, N20807, N6981);
buf BUF1 (N23427, N23426);
nor NOR3 (N23428, N23408, N19391, N15212);
buf BUF1 (N23429, N23419);
not NOT1 (N23430, N23425);
and AND3 (N23431, N23428, N15126, N5955);
xor XOR2 (N23432, N23420, N15601);
not NOT1 (N23433, N23413);
nand NAND3 (N23434, N23429, N23078, N13267);
not NOT1 (N23435, N23430);
nand NAND4 (N23436, N23427, N7188, N22541, N5208);
and AND4 (N23437, N23422, N3994, N12142, N8339);
and AND2 (N23438, N23424, N5590);
xor XOR2 (N23439, N23431, N13500);
or OR2 (N23440, N23434, N10592);
buf BUF1 (N23441, N23421);
not NOT1 (N23442, N23439);
nor NOR4 (N23443, N23432, N16641, N1792, N7391);
xor XOR2 (N23444, N23441, N9314);
nand NAND3 (N23445, N23433, N23065, N7980);
buf BUF1 (N23446, N23444);
or OR3 (N23447, N23440, N11453, N2605);
xor XOR2 (N23448, N23446, N5992);
xor XOR2 (N23449, N23437, N1594);
xor XOR2 (N23450, N23443, N20061);
nand NAND3 (N23451, N23448, N18841, N21406);
or OR3 (N23452, N23435, N17401, N2603);
nor NOR4 (N23453, N23452, N5697, N14818, N20331);
not NOT1 (N23454, N23445);
or OR3 (N23455, N23450, N1400, N2664);
nand NAND2 (N23456, N23449, N19377);
not NOT1 (N23457, N23438);
and AND2 (N23458, N23457, N4381);
nand NAND3 (N23459, N23455, N2819, N20894);
nor NOR4 (N23460, N23451, N2102, N8365, N9302);
nand NAND4 (N23461, N23458, N14772, N12378, N18705);
nor NOR2 (N23462, N23447, N5124);
nor NOR4 (N23463, N23460, N13404, N12138, N5992);
nor NOR2 (N23464, N23463, N11283);
buf BUF1 (N23465, N23459);
or OR4 (N23466, N23462, N10524, N18530, N2567);
xor XOR2 (N23467, N23442, N13242);
nand NAND3 (N23468, N23454, N951, N9826);
or OR2 (N23469, N23453, N13194);
and AND4 (N23470, N23465, N6148, N22771, N22415);
buf BUF1 (N23471, N23436);
and AND2 (N23472, N23418, N12097);
not NOT1 (N23473, N23470);
nor NOR2 (N23474, N23456, N22254);
and AND4 (N23475, N23469, N12134, N7400, N19160);
nor NOR4 (N23476, N23474, N13263, N9284, N14758);
not NOT1 (N23477, N23468);
buf BUF1 (N23478, N23476);
nor NOR4 (N23479, N23472, N8477, N18558, N13670);
not NOT1 (N23480, N23471);
nand NAND4 (N23481, N23479, N7288, N20380, N11863);
and AND3 (N23482, N23466, N9301, N19583);
and AND4 (N23483, N23467, N23394, N1179, N7646);
xor XOR2 (N23484, N23477, N7357);
nor NOR4 (N23485, N23483, N23465, N16141, N21439);
or OR4 (N23486, N23485, N6120, N1691, N21265);
xor XOR2 (N23487, N23486, N21716);
not NOT1 (N23488, N23487);
and AND3 (N23489, N23488, N811, N14041);
and AND4 (N23490, N23489, N2587, N7005, N5764);
nand NAND4 (N23491, N23484, N7842, N9145, N929);
nor NOR3 (N23492, N23461, N22368, N11086);
or OR2 (N23493, N23473, N20838);
buf BUF1 (N23494, N23493);
nor NOR3 (N23495, N23482, N12691, N20322);
nor NOR2 (N23496, N23491, N15231);
and AND4 (N23497, N23494, N12357, N3096, N20967);
buf BUF1 (N23498, N23497);
or OR4 (N23499, N23495, N9585, N9409, N9484);
nor NOR4 (N23500, N23498, N19088, N19558, N3590);
xor XOR2 (N23501, N23490, N11888);
buf BUF1 (N23502, N23496);
nor NOR4 (N23503, N23475, N17510, N15593, N13858);
nor NOR4 (N23504, N23499, N6791, N19895, N17504);
and AND2 (N23505, N23480, N6942);
nor NOR2 (N23506, N23504, N15802);
xor XOR2 (N23507, N23500, N22721);
xor XOR2 (N23508, N23478, N7395);
nor NOR3 (N23509, N23481, N876, N6027);
or OR4 (N23510, N23492, N19795, N22340, N3415);
not NOT1 (N23511, N23502);
xor XOR2 (N23512, N23464, N9824);
or OR2 (N23513, N23512, N12763);
or OR2 (N23514, N23505, N9905);
nand NAND4 (N23515, N23510, N2165, N8749, N14784);
xor XOR2 (N23516, N23515, N6894);
and AND3 (N23517, N23509, N17008, N1273);
or OR3 (N23518, N23506, N8833, N7948);
and AND2 (N23519, N23507, N22786);
not NOT1 (N23520, N23508);
buf BUF1 (N23521, N23514);
nand NAND4 (N23522, N23501, N8969, N11559, N13806);
nor NOR2 (N23523, N23522, N23435);
xor XOR2 (N23524, N23520, N6077);
not NOT1 (N23525, N23517);
or OR2 (N23526, N23511, N16603);
xor XOR2 (N23527, N23503, N23501);
or OR2 (N23528, N23523, N2425);
not NOT1 (N23529, N23513);
buf BUF1 (N23530, N23525);
xor XOR2 (N23531, N23528, N3462);
not NOT1 (N23532, N23521);
nand NAND4 (N23533, N23531, N2235, N15839, N18032);
or OR3 (N23534, N23526, N14486, N15430);
buf BUF1 (N23535, N23524);
buf BUF1 (N23536, N23519);
xor XOR2 (N23537, N23534, N21825);
not NOT1 (N23538, N23537);
not NOT1 (N23539, N23536);
and AND3 (N23540, N23518, N19752, N6765);
nand NAND4 (N23541, N23538, N13287, N17316, N23055);
or OR2 (N23542, N23541, N2260);
xor XOR2 (N23543, N23540, N20004);
not NOT1 (N23544, N23527);
nor NOR2 (N23545, N23544, N17555);
buf BUF1 (N23546, N23533);
nor NOR2 (N23547, N23530, N20740);
buf BUF1 (N23548, N23545);
and AND2 (N23549, N23542, N5139);
nand NAND4 (N23550, N23548, N13086, N2176, N19671);
or OR2 (N23551, N23516, N12072);
or OR4 (N23552, N23543, N14910, N14174, N17426);
nand NAND3 (N23553, N23547, N16312, N13821);
xor XOR2 (N23554, N23539, N23015);
and AND2 (N23555, N23529, N20188);
buf BUF1 (N23556, N23546);
nor NOR2 (N23557, N23532, N13141);
xor XOR2 (N23558, N23554, N22321);
or OR4 (N23559, N23552, N13840, N12905, N19449);
nor NOR4 (N23560, N23557, N4480, N19548, N2553);
not NOT1 (N23561, N23551);
or OR4 (N23562, N23560, N12730, N19315, N3312);
nand NAND2 (N23563, N23555, N5958);
xor XOR2 (N23564, N23550, N575);
nor NOR2 (N23565, N23564, N7901);
xor XOR2 (N23566, N23535, N8495);
or OR4 (N23567, N23563, N7933, N11183, N8555);
and AND4 (N23568, N23558, N15966, N305, N16247);
nor NOR2 (N23569, N23562, N3257);
nor NOR2 (N23570, N23561, N22693);
and AND3 (N23571, N23570, N2221, N11696);
not NOT1 (N23572, N23566);
or OR2 (N23573, N23553, N21124);
or OR3 (N23574, N23549, N1947, N4075);
xor XOR2 (N23575, N23569, N21713);
nor NOR3 (N23576, N23568, N19783, N20259);
and AND4 (N23577, N23556, N5053, N3327, N14991);
nand NAND3 (N23578, N23571, N13050, N10305);
buf BUF1 (N23579, N23572);
or OR4 (N23580, N23576, N6712, N14809, N10279);
and AND3 (N23581, N23559, N5501, N8420);
nand NAND3 (N23582, N23567, N397, N5541);
not NOT1 (N23583, N23574);
not NOT1 (N23584, N23580);
xor XOR2 (N23585, N23577, N16924);
and AND4 (N23586, N23582, N13737, N16442, N3040);
nand NAND4 (N23587, N23583, N11140, N11040, N15680);
nand NAND2 (N23588, N23584, N2255);
xor XOR2 (N23589, N23587, N2783);
xor XOR2 (N23590, N23575, N22974);
nor NOR3 (N23591, N23565, N2720, N624);
not NOT1 (N23592, N23586);
nor NOR4 (N23593, N23585, N3433, N14430, N5007);
buf BUF1 (N23594, N23581);
or OR3 (N23595, N23594, N18648, N19390);
buf BUF1 (N23596, N23595);
nand NAND3 (N23597, N23573, N4386, N18505);
and AND2 (N23598, N23591, N18518);
buf BUF1 (N23599, N23598);
nand NAND3 (N23600, N23596, N22978, N4473);
buf BUF1 (N23601, N23593);
or OR2 (N23602, N23599, N21173);
xor XOR2 (N23603, N23590, N2582);
xor XOR2 (N23604, N23597, N18369);
xor XOR2 (N23605, N23589, N21083);
or OR2 (N23606, N23601, N13612);
xor XOR2 (N23607, N23604, N21015);
buf BUF1 (N23608, N23588);
buf BUF1 (N23609, N23578);
and AND2 (N23610, N23592, N11929);
nor NOR4 (N23611, N23600, N20783, N15589, N4472);
or OR3 (N23612, N23610, N22680, N16248);
nand NAND2 (N23613, N23607, N15410);
xor XOR2 (N23614, N23605, N23225);
xor XOR2 (N23615, N23613, N15267);
nand NAND2 (N23616, N23609, N8432);
nor NOR2 (N23617, N23603, N21187);
nor NOR2 (N23618, N23614, N20078);
or OR4 (N23619, N23612, N4519, N19151, N1768);
and AND4 (N23620, N23611, N5318, N5259, N8488);
buf BUF1 (N23621, N23608);
buf BUF1 (N23622, N23606);
buf BUF1 (N23623, N23622);
not NOT1 (N23624, N23618);
not NOT1 (N23625, N23615);
not NOT1 (N23626, N23624);
xor XOR2 (N23627, N23620, N8163);
not NOT1 (N23628, N23621);
not NOT1 (N23629, N23627);
xor XOR2 (N23630, N23602, N19750);
nand NAND3 (N23631, N23623, N5498, N7943);
nor NOR4 (N23632, N23619, N2092, N11193, N16929);
not NOT1 (N23633, N23617);
nand NAND2 (N23634, N23629, N7420);
buf BUF1 (N23635, N23631);
and AND3 (N23636, N23626, N18967, N10246);
and AND2 (N23637, N23630, N7170);
xor XOR2 (N23638, N23634, N9392);
nor NOR2 (N23639, N23628, N7784);
not NOT1 (N23640, N23638);
and AND4 (N23641, N23640, N16785, N18013, N13132);
xor XOR2 (N23642, N23641, N17626);
nand NAND4 (N23643, N23642, N21062, N11249, N7794);
or OR2 (N23644, N23579, N10869);
or OR3 (N23645, N23635, N22767, N827);
xor XOR2 (N23646, N23636, N8499);
nor NOR3 (N23647, N23639, N14022, N9753);
nand NAND4 (N23648, N23647, N3282, N5252, N18174);
nor NOR3 (N23649, N23637, N11485, N15703);
nor NOR3 (N23650, N23644, N15171, N3471);
or OR2 (N23651, N23645, N16966);
nor NOR2 (N23652, N23643, N16440);
not NOT1 (N23653, N23632);
not NOT1 (N23654, N23653);
nand NAND2 (N23655, N23651, N7204);
nand NAND3 (N23656, N23646, N10665, N15298);
nor NOR2 (N23657, N23650, N8983);
nor NOR3 (N23658, N23652, N9370, N9292);
xor XOR2 (N23659, N23657, N18202);
xor XOR2 (N23660, N23625, N11343);
not NOT1 (N23661, N23656);
or OR4 (N23662, N23616, N17390, N8901, N13534);
xor XOR2 (N23663, N23662, N9994);
nand NAND2 (N23664, N23660, N11165);
not NOT1 (N23665, N23654);
and AND4 (N23666, N23655, N7896, N7400, N10032);
not NOT1 (N23667, N23658);
xor XOR2 (N23668, N23663, N5610);
not NOT1 (N23669, N23633);
xor XOR2 (N23670, N23669, N2364);
buf BUF1 (N23671, N23670);
and AND2 (N23672, N23659, N3339);
and AND3 (N23673, N23672, N5927, N17364);
not NOT1 (N23674, N23673);
and AND2 (N23675, N23664, N16553);
buf BUF1 (N23676, N23674);
xor XOR2 (N23677, N23671, N11826);
not NOT1 (N23678, N23648);
not NOT1 (N23679, N23668);
xor XOR2 (N23680, N23667, N19216);
or OR2 (N23681, N23661, N5741);
not NOT1 (N23682, N23680);
xor XOR2 (N23683, N23665, N7801);
buf BUF1 (N23684, N23683);
nor NOR2 (N23685, N23675, N20191);
nor NOR4 (N23686, N23678, N9750, N20456, N17201);
and AND4 (N23687, N23677, N4028, N13756, N800);
nand NAND4 (N23688, N23687, N5779, N3186, N13148);
not NOT1 (N23689, N23682);
buf BUF1 (N23690, N23688);
nand NAND4 (N23691, N23681, N8391, N6052, N14349);
or OR3 (N23692, N23691, N2332, N7899);
nor NOR3 (N23693, N23690, N15858, N7809);
nand NAND3 (N23694, N23684, N7896, N6515);
nor NOR2 (N23695, N23676, N15459);
or OR3 (N23696, N23649, N2274, N626);
nor NOR3 (N23697, N23679, N1267, N13063);
and AND2 (N23698, N23697, N15488);
xor XOR2 (N23699, N23666, N8632);
not NOT1 (N23700, N23696);
nand NAND3 (N23701, N23685, N15063, N2663);
or OR2 (N23702, N23700, N10675);
nand NAND3 (N23703, N23699, N6882, N14154);
buf BUF1 (N23704, N23701);
nor NOR4 (N23705, N23704, N13882, N3979, N17759);
not NOT1 (N23706, N23702);
or OR2 (N23707, N23686, N20050);
nand NAND4 (N23708, N23698, N3561, N21251, N7028);
xor XOR2 (N23709, N23693, N7146);
buf BUF1 (N23710, N23708);
nand NAND4 (N23711, N23709, N13355, N1774, N7138);
nor NOR4 (N23712, N23692, N13518, N13846, N10587);
buf BUF1 (N23713, N23694);
buf BUF1 (N23714, N23707);
buf BUF1 (N23715, N23710);
xor XOR2 (N23716, N23711, N6115);
or OR4 (N23717, N23715, N9695, N21568, N7729);
nand NAND3 (N23718, N23689, N1238, N9926);
not NOT1 (N23719, N23695);
xor XOR2 (N23720, N23718, N719);
xor XOR2 (N23721, N23703, N11372);
not NOT1 (N23722, N23714);
nor NOR3 (N23723, N23716, N21407, N13624);
nand NAND2 (N23724, N23713, N21999);
nand NAND4 (N23725, N23720, N15630, N4494, N7246);
or OR2 (N23726, N23723, N13419);
nand NAND3 (N23727, N23721, N21622, N5570);
nor NOR3 (N23728, N23725, N10690, N663);
not NOT1 (N23729, N23717);
nand NAND3 (N23730, N23706, N4982, N4151);
nor NOR2 (N23731, N23705, N7729);
nor NOR3 (N23732, N23727, N19811, N8499);
nor NOR2 (N23733, N23722, N17163);
nor NOR4 (N23734, N23724, N23646, N6484, N11811);
not NOT1 (N23735, N23729);
nor NOR2 (N23736, N23726, N975);
buf BUF1 (N23737, N23712);
buf BUF1 (N23738, N23736);
not NOT1 (N23739, N23728);
and AND4 (N23740, N23735, N10206, N11310, N15461);
nor NOR3 (N23741, N23737, N21895, N13153);
buf BUF1 (N23742, N23739);
or OR2 (N23743, N23740, N5705);
xor XOR2 (N23744, N23741, N9456);
buf BUF1 (N23745, N23744);
nand NAND3 (N23746, N23733, N16895, N9028);
not NOT1 (N23747, N23732);
or OR3 (N23748, N23745, N14991, N11869);
nand NAND3 (N23749, N23746, N22946, N17872);
nand NAND4 (N23750, N23731, N14852, N2898, N17276);
nor NOR3 (N23751, N23734, N10319, N6438);
not NOT1 (N23752, N23748);
buf BUF1 (N23753, N23738);
nor NOR4 (N23754, N23750, N11339, N13847, N5121);
not NOT1 (N23755, N23747);
nor NOR4 (N23756, N23730, N1307, N12666, N20943);
not NOT1 (N23757, N23743);
not NOT1 (N23758, N23742);
nand NAND2 (N23759, N23719, N19650);
and AND4 (N23760, N23756, N12692, N21674, N13955);
not NOT1 (N23761, N23755);
and AND2 (N23762, N23761, N2240);
or OR2 (N23763, N23752, N902);
nand NAND3 (N23764, N23753, N7851, N1468);
buf BUF1 (N23765, N23758);
or OR2 (N23766, N23763, N5781);
buf BUF1 (N23767, N23759);
not NOT1 (N23768, N23754);
nor NOR3 (N23769, N23749, N7464, N7529);
nand NAND2 (N23770, N23765, N20621);
nand NAND4 (N23771, N23770, N4352, N19641, N9953);
nor NOR3 (N23772, N23757, N2681, N13661);
xor XOR2 (N23773, N23767, N15644);
not NOT1 (N23774, N23773);
buf BUF1 (N23775, N23774);
nand NAND3 (N23776, N23762, N2512, N23717);
buf BUF1 (N23777, N23775);
not NOT1 (N23778, N23768);
and AND3 (N23779, N23771, N7037, N2416);
xor XOR2 (N23780, N23764, N23338);
or OR2 (N23781, N23751, N8898);
nor NOR2 (N23782, N23779, N8646);
buf BUF1 (N23783, N23778);
not NOT1 (N23784, N23781);
nand NAND2 (N23785, N23784, N14920);
nor NOR2 (N23786, N23766, N9783);
nor NOR4 (N23787, N23769, N21801, N15293, N4308);
buf BUF1 (N23788, N23760);
not NOT1 (N23789, N23787);
or OR4 (N23790, N23789, N473, N15049, N16274);
not NOT1 (N23791, N23780);
and AND3 (N23792, N23788, N9061, N2741);
not NOT1 (N23793, N23790);
not NOT1 (N23794, N23793);
buf BUF1 (N23795, N23791);
xor XOR2 (N23796, N23782, N17069);
and AND2 (N23797, N23794, N23539);
or OR3 (N23798, N23776, N14142, N4553);
xor XOR2 (N23799, N23783, N22394);
or OR4 (N23800, N23772, N18501, N18107, N22098);
and AND2 (N23801, N23798, N4289);
and AND2 (N23802, N23785, N14935);
xor XOR2 (N23803, N23799, N9656);
nor NOR4 (N23804, N23800, N15496, N7157, N8795);
not NOT1 (N23805, N23802);
nand NAND4 (N23806, N23795, N23538, N20259, N18376);
buf BUF1 (N23807, N23777);
nor NOR4 (N23808, N23801, N7122, N5120, N9452);
or OR4 (N23809, N23796, N15624, N20999, N1936);
nor NOR4 (N23810, N23792, N15416, N18647, N6952);
nor NOR3 (N23811, N23806, N22630, N8195);
buf BUF1 (N23812, N23804);
buf BUF1 (N23813, N23811);
or OR3 (N23814, N23810, N4169, N18780);
buf BUF1 (N23815, N23805);
buf BUF1 (N23816, N23812);
not NOT1 (N23817, N23815);
xor XOR2 (N23818, N23803, N7702);
nor NOR3 (N23819, N23809, N2022, N10538);
or OR4 (N23820, N23808, N22170, N23049, N6264);
and AND3 (N23821, N23820, N3614, N20551);
not NOT1 (N23822, N23807);
nand NAND2 (N23823, N23797, N17666);
nand NAND4 (N23824, N23814, N8079, N8568, N14970);
not NOT1 (N23825, N23813);
or OR2 (N23826, N23822, N22544);
nor NOR4 (N23827, N23821, N7614, N6882, N7971);
nand NAND2 (N23828, N23819, N714);
nor NOR4 (N23829, N23786, N12219, N16921, N21573);
or OR3 (N23830, N23818, N12444, N17336);
nor NOR3 (N23831, N23828, N9005, N9696);
nor NOR3 (N23832, N23826, N21398, N11896);
buf BUF1 (N23833, N23829);
buf BUF1 (N23834, N23817);
not NOT1 (N23835, N23827);
not NOT1 (N23836, N23831);
not NOT1 (N23837, N23832);
not NOT1 (N23838, N23825);
and AND3 (N23839, N23816, N15709, N10843);
nand NAND4 (N23840, N23838, N9987, N19717, N12032);
or OR4 (N23841, N23839, N7607, N746, N1034);
or OR2 (N23842, N23824, N478);
and AND2 (N23843, N23842, N21997);
and AND4 (N23844, N23830, N6322, N7318, N10443);
nor NOR3 (N23845, N23841, N3805, N16177);
nand NAND2 (N23846, N23845, N15467);
nor NOR2 (N23847, N23840, N19663);
nor NOR4 (N23848, N23835, N5585, N5886, N1012);
nand NAND3 (N23849, N23834, N88, N6794);
xor XOR2 (N23850, N23846, N12628);
not NOT1 (N23851, N23843);
xor XOR2 (N23852, N23850, N17050);
buf BUF1 (N23853, N23851);
xor XOR2 (N23854, N23852, N768);
buf BUF1 (N23855, N23849);
nor NOR2 (N23856, N23855, N10524);
nor NOR3 (N23857, N23836, N11327, N22469);
or OR4 (N23858, N23857, N17319, N3040, N7009);
nor NOR3 (N23859, N23848, N821, N11889);
nand NAND3 (N23860, N23859, N366, N17207);
buf BUF1 (N23861, N23833);
xor XOR2 (N23862, N23861, N23807);
and AND4 (N23863, N23858, N17522, N3818, N20589);
not NOT1 (N23864, N23863);
nand NAND3 (N23865, N23860, N16988, N22824);
and AND3 (N23866, N23847, N2252, N3008);
or OR3 (N23867, N23864, N19725, N14423);
buf BUF1 (N23868, N23853);
buf BUF1 (N23869, N23867);
buf BUF1 (N23870, N23856);
xor XOR2 (N23871, N23837, N10093);
and AND3 (N23872, N23870, N6516, N5414);
xor XOR2 (N23873, N23823, N662);
and AND3 (N23874, N23871, N4909, N13646);
or OR3 (N23875, N23872, N523, N11920);
not NOT1 (N23876, N23854);
nor NOR2 (N23877, N23866, N15043);
not NOT1 (N23878, N23865);
buf BUF1 (N23879, N23868);
nor NOR2 (N23880, N23877, N9649);
and AND3 (N23881, N23878, N1613, N10166);
and AND2 (N23882, N23862, N23597);
and AND3 (N23883, N23869, N9873, N17194);
or OR4 (N23884, N23874, N17317, N17006, N16268);
and AND2 (N23885, N23879, N8544);
and AND2 (N23886, N23882, N4051);
nor NOR4 (N23887, N23876, N11394, N268, N1852);
or OR3 (N23888, N23844, N11079, N6473);
nand NAND4 (N23889, N23873, N18066, N19829, N22881);
not NOT1 (N23890, N23881);
not NOT1 (N23891, N23885);
xor XOR2 (N23892, N23875, N14582);
nor NOR4 (N23893, N23883, N13659, N15532, N19476);
buf BUF1 (N23894, N23891);
nor NOR4 (N23895, N23886, N23568, N20771, N6067);
not NOT1 (N23896, N23895);
and AND3 (N23897, N23887, N9973, N14424);
buf BUF1 (N23898, N23884);
nand NAND4 (N23899, N23896, N16566, N2729, N16480);
nand NAND3 (N23900, N23893, N8139, N19060);
not NOT1 (N23901, N23897);
xor XOR2 (N23902, N23901, N10038);
and AND2 (N23903, N23898, N23142);
nand NAND3 (N23904, N23902, N623, N7443);
buf BUF1 (N23905, N23899);
or OR2 (N23906, N23888, N3370);
or OR3 (N23907, N23894, N19582, N21061);
xor XOR2 (N23908, N23892, N1112);
nor NOR4 (N23909, N23903, N10937, N23139, N432);
and AND2 (N23910, N23908, N13766);
or OR2 (N23911, N23890, N20435);
not NOT1 (N23912, N23904);
or OR4 (N23913, N23900, N23144, N10947, N4294);
nor NOR4 (N23914, N23906, N4926, N442, N9006);
and AND2 (N23915, N23912, N11900);
and AND4 (N23916, N23914, N17285, N23525, N10551);
or OR4 (N23917, N23911, N17548, N20368, N8869);
xor XOR2 (N23918, N23907, N9529);
buf BUF1 (N23919, N23915);
nor NOR4 (N23920, N23919, N4207, N23179, N8358);
not NOT1 (N23921, N23918);
nor NOR2 (N23922, N23913, N10071);
and AND3 (N23923, N23920, N13449, N10598);
or OR2 (N23924, N23910, N1282);
nand NAND4 (N23925, N23923, N2145, N9001, N6336);
not NOT1 (N23926, N23925);
nand NAND4 (N23927, N23905, N9972, N14482, N10701);
nand NAND2 (N23928, N23909, N7748);
xor XOR2 (N23929, N23922, N18387);
or OR2 (N23930, N23889, N15398);
nand NAND3 (N23931, N23916, N6259, N16775);
buf BUF1 (N23932, N23924);
xor XOR2 (N23933, N23917, N101);
not NOT1 (N23934, N23928);
or OR4 (N23935, N23933, N23384, N23407, N22804);
nand NAND4 (N23936, N23929, N1399, N5185, N22238);
xor XOR2 (N23937, N23931, N14461);
and AND2 (N23938, N23936, N13633);
and AND3 (N23939, N23937, N13896, N23819);
nor NOR2 (N23940, N23930, N7245);
nor NOR2 (N23941, N23935, N129);
nand NAND3 (N23942, N23880, N11845, N12045);
nor NOR2 (N23943, N23940, N10649);
xor XOR2 (N23944, N23943, N18559);
nor NOR2 (N23945, N23934, N2478);
or OR3 (N23946, N23927, N16613, N5544);
and AND3 (N23947, N23932, N11046, N11315);
and AND3 (N23948, N23945, N11541, N15755);
xor XOR2 (N23949, N23948, N10783);
nor NOR4 (N23950, N23949, N12122, N10367, N14176);
xor XOR2 (N23951, N23921, N1327);
and AND2 (N23952, N23947, N10245);
xor XOR2 (N23953, N23939, N6518);
or OR3 (N23954, N23938, N1788, N2556);
nand NAND3 (N23955, N23926, N14988, N22143);
xor XOR2 (N23956, N23955, N23445);
or OR2 (N23957, N23952, N10294);
nand NAND4 (N23958, N23942, N22987, N3033, N14468);
xor XOR2 (N23959, N23954, N662);
nor NOR3 (N23960, N23946, N9646, N21173);
not NOT1 (N23961, N23956);
xor XOR2 (N23962, N23957, N10016);
nor NOR3 (N23963, N23958, N7565, N5800);
nand NAND2 (N23964, N23953, N7482);
and AND2 (N23965, N23959, N1474);
xor XOR2 (N23966, N23960, N4230);
and AND4 (N23967, N23965, N8692, N15315, N20756);
nand NAND4 (N23968, N23967, N13707, N10002, N19633);
nand NAND2 (N23969, N23951, N6264);
nor NOR2 (N23970, N23966, N20287);
nor NOR2 (N23971, N23962, N5067);
not NOT1 (N23972, N23941);
xor XOR2 (N23973, N23970, N23129);
and AND3 (N23974, N23968, N18173, N22231);
xor XOR2 (N23975, N23971, N13636);
nor NOR3 (N23976, N23950, N16285, N2829);
and AND4 (N23977, N23963, N1573, N22248, N5798);
not NOT1 (N23978, N23973);
and AND4 (N23979, N23972, N18067, N23700, N21580);
and AND3 (N23980, N23961, N16739, N18454);
nor NOR2 (N23981, N23980, N20080);
xor XOR2 (N23982, N23975, N19005);
nand NAND3 (N23983, N23977, N23147, N23230);
nand NAND3 (N23984, N23981, N3548, N21561);
buf BUF1 (N23985, N23964);
nor NOR3 (N23986, N23978, N6506, N5800);
nor NOR3 (N23987, N23986, N20406, N22140);
or OR2 (N23988, N23944, N14737);
nor NOR3 (N23989, N23983, N4951, N10709);
xor XOR2 (N23990, N23984, N4581);
and AND3 (N23991, N23988, N4510, N845);
nor NOR3 (N23992, N23976, N11182, N9157);
nand NAND3 (N23993, N23991, N13791, N21516);
nor NOR3 (N23994, N23993, N23574, N16875);
and AND4 (N23995, N23969, N19286, N15183, N5973);
nor NOR4 (N23996, N23990, N7016, N12457, N11427);
buf BUF1 (N23997, N23985);
or OR3 (N23998, N23979, N16829, N19194);
not NOT1 (N23999, N23995);
and AND3 (N24000, N23998, N13246, N12885);
or OR4 (N24001, N24000, N8554, N5149, N20);
xor XOR2 (N24002, N23997, N6511);
and AND2 (N24003, N23999, N20669);
buf BUF1 (N24004, N23989);
not NOT1 (N24005, N24002);
nor NOR4 (N24006, N23987, N16301, N5818, N17953);
buf BUF1 (N24007, N24001);
nand NAND3 (N24008, N24005, N10018, N20790);
buf BUF1 (N24009, N23974);
or OR2 (N24010, N24003, N10162);
xor XOR2 (N24011, N23996, N14628);
buf BUF1 (N24012, N24009);
or OR4 (N24013, N24008, N20097, N19299, N11265);
not NOT1 (N24014, N24010);
nor NOR2 (N24015, N24011, N20692);
not NOT1 (N24016, N23992);
not NOT1 (N24017, N24016);
nor NOR4 (N24018, N24012, N14373, N14771, N16088);
nand NAND4 (N24019, N24018, N10791, N1437, N3001);
buf BUF1 (N24020, N23982);
not NOT1 (N24021, N24004);
nor NOR4 (N24022, N24014, N8590, N12437, N4709);
nor NOR4 (N24023, N24013, N515, N890, N12937);
nor NOR4 (N24024, N24017, N10788, N5804, N18949);
xor XOR2 (N24025, N24020, N8008);
not NOT1 (N24026, N24021);
buf BUF1 (N24027, N24022);
and AND4 (N24028, N23994, N8768, N3222, N4986);
xor XOR2 (N24029, N24025, N23252);
nand NAND3 (N24030, N24019, N16546, N19213);
not NOT1 (N24031, N24015);
or OR3 (N24032, N24029, N13511, N5055);
or OR3 (N24033, N24006, N11757, N15990);
nand NAND4 (N24034, N24033, N21471, N5222, N17128);
nand NAND3 (N24035, N24007, N12673, N22251);
buf BUF1 (N24036, N24031);
or OR2 (N24037, N24024, N17853);
or OR3 (N24038, N24027, N8897, N14826);
xor XOR2 (N24039, N24030, N12184);
buf BUF1 (N24040, N24038);
xor XOR2 (N24041, N24023, N11401);
not NOT1 (N24042, N24037);
or OR4 (N24043, N24026, N21100, N19187, N2205);
buf BUF1 (N24044, N24032);
buf BUF1 (N24045, N24043);
or OR3 (N24046, N24045, N8403, N23817);
or OR4 (N24047, N24041, N1795, N15482, N15166);
nand NAND3 (N24048, N24047, N1692, N8183);
and AND3 (N24049, N24035, N17717, N2721);
buf BUF1 (N24050, N24046);
and AND4 (N24051, N24028, N12835, N22649, N3077);
not NOT1 (N24052, N24036);
and AND2 (N24053, N24052, N9460);
not NOT1 (N24054, N24053);
or OR3 (N24055, N24050, N8626, N17346);
buf BUF1 (N24056, N24044);
not NOT1 (N24057, N24040);
nand NAND4 (N24058, N24042, N6102, N2723, N6220);
or OR4 (N24059, N24051, N14570, N78, N13503);
buf BUF1 (N24060, N24055);
buf BUF1 (N24061, N24058);
xor XOR2 (N24062, N24057, N16981);
nand NAND3 (N24063, N24062, N3293, N19496);
nand NAND2 (N24064, N24048, N9281);
buf BUF1 (N24065, N24063);
buf BUF1 (N24066, N24065);
xor XOR2 (N24067, N24060, N19736);
and AND2 (N24068, N24049, N645);
buf BUF1 (N24069, N24039);
nor NOR3 (N24070, N24066, N1812, N23153);
or OR4 (N24071, N24054, N4367, N18972, N13309);
or OR4 (N24072, N24061, N1439, N6164, N23193);
xor XOR2 (N24073, N24071, N7970);
nor NOR2 (N24074, N24056, N11349);
or OR4 (N24075, N24034, N5848, N2536, N997);
buf BUF1 (N24076, N24075);
nor NOR4 (N24077, N24067, N7904, N9864, N6050);
or OR3 (N24078, N24070, N22337, N3235);
xor XOR2 (N24079, N24064, N1619);
buf BUF1 (N24080, N24068);
nor NOR2 (N24081, N24076, N22290);
not NOT1 (N24082, N24080);
xor XOR2 (N24083, N24074, N5192);
xor XOR2 (N24084, N24059, N7117);
xor XOR2 (N24085, N24073, N20608);
nand NAND3 (N24086, N24072, N752, N15762);
or OR2 (N24087, N24085, N10335);
xor XOR2 (N24088, N24086, N7658);
buf BUF1 (N24089, N24082);
and AND3 (N24090, N24078, N24041, N13800);
not NOT1 (N24091, N24081);
or OR3 (N24092, N24084, N14277, N12120);
buf BUF1 (N24093, N24092);
nor NOR2 (N24094, N24091, N4199);
not NOT1 (N24095, N24077);
and AND4 (N24096, N24089, N9293, N16277, N12779);
nor NOR2 (N24097, N24069, N18085);
xor XOR2 (N24098, N24095, N21719);
buf BUF1 (N24099, N24090);
or OR4 (N24100, N24096, N13444, N662, N5602);
or OR3 (N24101, N24094, N23099, N15219);
nor NOR4 (N24102, N24101, N14823, N11224, N21030);
nor NOR4 (N24103, N24079, N21366, N10978, N15715);
nand NAND3 (N24104, N24083, N6738, N12527);
nand NAND4 (N24105, N24088, N19671, N21262, N13113);
nand NAND3 (N24106, N24098, N17622, N18519);
nor NOR2 (N24107, N24106, N21466);
not NOT1 (N24108, N24093);
or OR2 (N24109, N24104, N18163);
and AND3 (N24110, N24099, N8370, N7312);
nand NAND2 (N24111, N24107, N12472);
and AND3 (N24112, N24110, N17246, N24097);
and AND4 (N24113, N403, N10817, N15635, N19273);
buf BUF1 (N24114, N24108);
not NOT1 (N24115, N24102);
xor XOR2 (N24116, N24112, N6761);
xor XOR2 (N24117, N24100, N3541);
nand NAND2 (N24118, N24114, N2782);
or OR3 (N24119, N24117, N15921, N1876);
buf BUF1 (N24120, N24115);
xor XOR2 (N24121, N24118, N20447);
or OR2 (N24122, N24116, N8694);
xor XOR2 (N24123, N24122, N2803);
not NOT1 (N24124, N24105);
not NOT1 (N24125, N24087);
buf BUF1 (N24126, N24113);
or OR3 (N24127, N24123, N10175, N301);
or OR2 (N24128, N24124, N15303);
buf BUF1 (N24129, N24126);
buf BUF1 (N24130, N24120);
and AND2 (N24131, N24109, N7580);
nand NAND4 (N24132, N24130, N6724, N15257, N5288);
nand NAND4 (N24133, N24129, N3483, N21553, N24067);
not NOT1 (N24134, N24133);
buf BUF1 (N24135, N24132);
or OR2 (N24136, N24121, N11441);
buf BUF1 (N24137, N24125);
buf BUF1 (N24138, N24128);
xor XOR2 (N24139, N24138, N4437);
nand NAND2 (N24140, N24119, N7234);
xor XOR2 (N24141, N24137, N18381);
xor XOR2 (N24142, N24131, N20877);
buf BUF1 (N24143, N24127);
or OR4 (N24144, N24134, N12268, N882, N1517);
nand NAND2 (N24145, N24111, N14998);
nand NAND2 (N24146, N24144, N2134);
nand NAND3 (N24147, N24103, N3149, N23814);
nor NOR3 (N24148, N24135, N22655, N1336);
not NOT1 (N24149, N24143);
and AND3 (N24150, N24139, N11667, N10929);
nor NOR3 (N24151, N24150, N5215, N18036);
xor XOR2 (N24152, N24147, N8823);
not NOT1 (N24153, N24149);
or OR4 (N24154, N24146, N1842, N20995, N20762);
nor NOR4 (N24155, N24154, N10428, N4091, N18919);
buf BUF1 (N24156, N24151);
not NOT1 (N24157, N24156);
or OR3 (N24158, N24148, N14948, N14418);
or OR2 (N24159, N24158, N16250);
or OR2 (N24160, N24159, N17362);
nand NAND3 (N24161, N24136, N20556, N3665);
or OR3 (N24162, N24145, N14696, N3352);
buf BUF1 (N24163, N24162);
buf BUF1 (N24164, N24141);
nor NOR3 (N24165, N24160, N21564, N12286);
or OR2 (N24166, N24165, N448);
or OR4 (N24167, N24140, N273, N1882, N19999);
nor NOR3 (N24168, N24153, N22752, N24048);
buf BUF1 (N24169, N24142);
or OR4 (N24170, N24163, N12782, N1894, N6276);
or OR3 (N24171, N24167, N5439, N13649);
xor XOR2 (N24172, N24155, N2296);
buf BUF1 (N24173, N24169);
or OR4 (N24174, N24171, N18594, N8714, N9809);
not NOT1 (N24175, N24174);
and AND2 (N24176, N24164, N19681);
not NOT1 (N24177, N24161);
nor NOR2 (N24178, N24152, N8188);
buf BUF1 (N24179, N24170);
not NOT1 (N24180, N24177);
or OR2 (N24181, N24157, N20414);
or OR3 (N24182, N24173, N1145, N19936);
buf BUF1 (N24183, N24181);
nor NOR2 (N24184, N24168, N3734);
and AND4 (N24185, N24179, N18553, N13143, N19727);
and AND4 (N24186, N24183, N10488, N7983, N12848);
and AND3 (N24187, N24184, N21537, N11593);
or OR4 (N24188, N24187, N21009, N15321, N10057);
and AND2 (N24189, N24178, N5232);
xor XOR2 (N24190, N24172, N22943);
nor NOR4 (N24191, N24190, N6166, N10643, N19692);
buf BUF1 (N24192, N24186);
nand NAND2 (N24193, N24188, N4613);
xor XOR2 (N24194, N24191, N9621);
and AND3 (N24195, N24193, N12387, N10634);
nor NOR3 (N24196, N24194, N3096, N22050);
xor XOR2 (N24197, N24176, N3545);
xor XOR2 (N24198, N24185, N22930);
nand NAND3 (N24199, N24180, N6493, N6427);
buf BUF1 (N24200, N24198);
nor NOR4 (N24201, N24195, N6193, N11551, N6209);
nand NAND4 (N24202, N24189, N19323, N22473, N18081);
nand NAND3 (N24203, N24182, N148, N6848);
and AND2 (N24204, N24199, N8828);
and AND2 (N24205, N24175, N14731);
and AND3 (N24206, N24205, N5697, N4269);
xor XOR2 (N24207, N24200, N21393);
nand NAND3 (N24208, N24196, N21545, N15299);
or OR3 (N24209, N24207, N20539, N23334);
nand NAND4 (N24210, N24203, N20516, N9577, N4334);
xor XOR2 (N24211, N24210, N6755);
nor NOR2 (N24212, N24206, N9905);
nand NAND4 (N24213, N24204, N21445, N21327, N19197);
or OR2 (N24214, N24208, N23589);
nand NAND4 (N24215, N24213, N5742, N21504, N15796);
xor XOR2 (N24216, N24212, N18946);
and AND3 (N24217, N24166, N6642, N21762);
nor NOR2 (N24218, N24211, N4115);
not NOT1 (N24219, N24218);
buf BUF1 (N24220, N24219);
and AND3 (N24221, N24214, N5925, N13136);
and AND3 (N24222, N24202, N18523, N9973);
and AND4 (N24223, N24197, N15195, N23829, N16596);
or OR3 (N24224, N24217, N4288, N15721);
nor NOR3 (N24225, N24221, N5904, N15449);
xor XOR2 (N24226, N24209, N1077);
not NOT1 (N24227, N24220);
xor XOR2 (N24228, N24224, N1884);
buf BUF1 (N24229, N24192);
and AND4 (N24230, N24227, N3603, N7083, N13387);
nand NAND2 (N24231, N24216, N20791);
nor NOR2 (N24232, N24223, N5575);
nand NAND3 (N24233, N24230, N8077, N16387);
and AND4 (N24234, N24215, N19668, N873, N18707);
nand NAND2 (N24235, N24225, N17713);
not NOT1 (N24236, N24235);
not NOT1 (N24237, N24234);
or OR2 (N24238, N24201, N17666);
buf BUF1 (N24239, N24222);
xor XOR2 (N24240, N24231, N12055);
xor XOR2 (N24241, N24238, N19533);
buf BUF1 (N24242, N24237);
or OR3 (N24243, N24228, N15871, N2869);
xor XOR2 (N24244, N24233, N22796);
and AND3 (N24245, N24229, N8917, N3442);
not NOT1 (N24246, N24232);
or OR2 (N24247, N24236, N3776);
nand NAND3 (N24248, N24246, N6735, N10518);
or OR2 (N24249, N24226, N7036);
and AND2 (N24250, N24248, N9523);
xor XOR2 (N24251, N24243, N17506);
nor NOR2 (N24252, N24249, N12785);
nand NAND4 (N24253, N24252, N17624, N1966, N3618);
buf BUF1 (N24254, N24251);
buf BUF1 (N24255, N24240);
and AND3 (N24256, N24244, N8172, N22152);
buf BUF1 (N24257, N24247);
buf BUF1 (N24258, N24253);
not NOT1 (N24259, N24254);
nor NOR3 (N24260, N24255, N7508, N21210);
xor XOR2 (N24261, N24258, N5672);
nor NOR3 (N24262, N24257, N8097, N21327);
and AND3 (N24263, N24241, N2754, N881);
nand NAND3 (N24264, N24259, N18361, N8613);
not NOT1 (N24265, N24262);
buf BUF1 (N24266, N24239);
nand NAND3 (N24267, N24250, N23749, N7499);
not NOT1 (N24268, N24260);
not NOT1 (N24269, N24261);
nor NOR4 (N24270, N24265, N16059, N11371, N12785);
xor XOR2 (N24271, N24266, N13203);
and AND3 (N24272, N24256, N17715, N6565);
buf BUF1 (N24273, N24270);
buf BUF1 (N24274, N24245);
not NOT1 (N24275, N24264);
xor XOR2 (N24276, N24268, N23794);
and AND3 (N24277, N24272, N4926, N19786);
buf BUF1 (N24278, N24275);
nand NAND3 (N24279, N24271, N22633, N17777);
or OR3 (N24280, N24274, N18748, N14015);
buf BUF1 (N24281, N24269);
xor XOR2 (N24282, N24267, N21456);
or OR3 (N24283, N24273, N11418, N4658);
and AND2 (N24284, N24283, N23588);
or OR3 (N24285, N24278, N8773, N22428);
xor XOR2 (N24286, N24277, N14239);
not NOT1 (N24287, N24263);
buf BUF1 (N24288, N24276);
or OR4 (N24289, N24279, N2476, N21791, N8171);
nor NOR3 (N24290, N24242, N6580, N12599);
nor NOR4 (N24291, N24289, N15781, N8761, N19774);
and AND4 (N24292, N24290, N22966, N4924, N22307);
nand NAND3 (N24293, N24287, N13530, N23116);
xor XOR2 (N24294, N24285, N8766);
not NOT1 (N24295, N24293);
buf BUF1 (N24296, N24294);
and AND3 (N24297, N24291, N22912, N4011);
nand NAND2 (N24298, N24286, N8516);
or OR2 (N24299, N24298, N15028);
not NOT1 (N24300, N24295);
not NOT1 (N24301, N24280);
xor XOR2 (N24302, N24292, N1747);
buf BUF1 (N24303, N24302);
nor NOR3 (N24304, N24284, N5543, N9679);
and AND3 (N24305, N24282, N151, N13690);
or OR3 (N24306, N24305, N10659, N7302);
xor XOR2 (N24307, N24306, N3132);
nand NAND4 (N24308, N24303, N2166, N2941, N6507);
buf BUF1 (N24309, N24304);
nor NOR2 (N24310, N24301, N15436);
not NOT1 (N24311, N24310);
nand NAND4 (N24312, N24308, N22623, N7, N2153);
buf BUF1 (N24313, N24296);
nand NAND3 (N24314, N24281, N20850, N22376);
or OR4 (N24315, N24312, N13064, N19160, N10120);
nor NOR3 (N24316, N24297, N12334, N15323);
or OR2 (N24317, N24316, N2936);
and AND3 (N24318, N24299, N12291, N1468);
or OR4 (N24319, N24315, N3758, N15849, N9817);
buf BUF1 (N24320, N24288);
xor XOR2 (N24321, N24314, N2115);
xor XOR2 (N24322, N24321, N14955);
nor NOR3 (N24323, N24318, N13544, N12355);
or OR4 (N24324, N24311, N10779, N9598, N5393);
and AND4 (N24325, N24319, N6337, N10874, N18303);
buf BUF1 (N24326, N24323);
or OR2 (N24327, N24317, N18798);
not NOT1 (N24328, N24325);
not NOT1 (N24329, N24309);
nor NOR2 (N24330, N24324, N5744);
and AND2 (N24331, N24328, N15846);
not NOT1 (N24332, N24330);
nor NOR2 (N24333, N24313, N8821);
xor XOR2 (N24334, N24332, N5050);
nand NAND2 (N24335, N24320, N22736);
nor NOR3 (N24336, N24333, N17197, N12128);
not NOT1 (N24337, N24331);
not NOT1 (N24338, N24300);
buf BUF1 (N24339, N24338);
nand NAND4 (N24340, N24329, N11688, N23681, N5657);
nand NAND4 (N24341, N24335, N2052, N2099, N7752);
buf BUF1 (N24342, N24307);
not NOT1 (N24343, N24327);
xor XOR2 (N24344, N24337, N12075);
xor XOR2 (N24345, N24322, N5824);
xor XOR2 (N24346, N24343, N15265);
nand NAND2 (N24347, N24326, N10188);
buf BUF1 (N24348, N24336);
and AND3 (N24349, N24347, N14955, N17499);
xor XOR2 (N24350, N24348, N1013);
buf BUF1 (N24351, N24342);
nor NOR4 (N24352, N24350, N22460, N7492, N23314);
nor NOR2 (N24353, N24345, N13265);
not NOT1 (N24354, N24346);
or OR4 (N24355, N24341, N9072, N23857, N16952);
xor XOR2 (N24356, N24355, N16063);
or OR2 (N24357, N24356, N2870);
and AND4 (N24358, N24339, N653, N17347, N7073);
nand NAND2 (N24359, N24354, N20231);
buf BUF1 (N24360, N24340);
xor XOR2 (N24361, N24358, N3013);
and AND2 (N24362, N24334, N24162);
xor XOR2 (N24363, N24357, N6670);
not NOT1 (N24364, N24353);
xor XOR2 (N24365, N24363, N18698);
nand NAND2 (N24366, N24359, N21698);
not NOT1 (N24367, N24365);
or OR2 (N24368, N24352, N12168);
nor NOR2 (N24369, N24364, N7984);
nor NOR3 (N24370, N24349, N22552, N18883);
nand NAND3 (N24371, N24369, N22129, N6257);
nor NOR4 (N24372, N24360, N2187, N7233, N21482);
nand NAND3 (N24373, N24366, N19848, N12410);
xor XOR2 (N24374, N24368, N23976);
or OR2 (N24375, N24367, N7645);
buf BUF1 (N24376, N24351);
or OR2 (N24377, N24373, N6135);
or OR3 (N24378, N24344, N2898, N18867);
or OR3 (N24379, N24376, N11907, N17873);
and AND2 (N24380, N24372, N24165);
xor XOR2 (N24381, N24377, N12708);
nand NAND2 (N24382, N24375, N8615);
not NOT1 (N24383, N24379);
xor XOR2 (N24384, N24378, N22267);
and AND4 (N24385, N24381, N17548, N23654, N4256);
and AND3 (N24386, N24380, N465, N20691);
xor XOR2 (N24387, N24386, N10561);
not NOT1 (N24388, N24362);
or OR3 (N24389, N24385, N8469, N13241);
xor XOR2 (N24390, N24387, N19180);
buf BUF1 (N24391, N24370);
xor XOR2 (N24392, N24383, N23180);
not NOT1 (N24393, N24374);
nor NOR2 (N24394, N24361, N3105);
buf BUF1 (N24395, N24382);
xor XOR2 (N24396, N24371, N14003);
not NOT1 (N24397, N24390);
not NOT1 (N24398, N24396);
not NOT1 (N24399, N24394);
or OR4 (N24400, N24384, N5135, N1677, N12243);
and AND2 (N24401, N24395, N18624);
not NOT1 (N24402, N24392);
nand NAND4 (N24403, N24397, N8059, N13903, N13825);
not NOT1 (N24404, N24391);
nand NAND4 (N24405, N24404, N19301, N6809, N23680);
and AND3 (N24406, N24401, N21527, N6735);
nor NOR4 (N24407, N24405, N22539, N15534, N4154);
and AND3 (N24408, N24402, N22465, N9652);
xor XOR2 (N24409, N24406, N3004);
and AND2 (N24410, N24400, N12541);
not NOT1 (N24411, N24389);
and AND2 (N24412, N24398, N23669);
nand NAND3 (N24413, N24408, N18029, N22340);
nor NOR4 (N24414, N24409, N19883, N24063, N17096);
nor NOR4 (N24415, N24403, N461, N9928, N14966);
and AND2 (N24416, N24393, N8685);
and AND4 (N24417, N24413, N19707, N8264, N13777);
not NOT1 (N24418, N24399);
nor NOR4 (N24419, N24416, N1753, N22177, N6159);
buf BUF1 (N24420, N24414);
or OR3 (N24421, N24417, N19721, N19285);
nor NOR3 (N24422, N24418, N13811, N21428);
or OR2 (N24423, N24421, N22444);
buf BUF1 (N24424, N24411);
nor NOR3 (N24425, N24415, N574, N13909);
or OR2 (N24426, N24419, N13085);
nor NOR4 (N24427, N24412, N2730, N13212, N1221);
xor XOR2 (N24428, N24426, N7344);
and AND2 (N24429, N24427, N21704);
nand NAND3 (N24430, N24407, N15433, N9706);
or OR2 (N24431, N24429, N23023);
and AND2 (N24432, N24425, N14824);
nor NOR2 (N24433, N24431, N12748);
nor NOR3 (N24434, N24430, N2793, N14773);
or OR4 (N24435, N24388, N6698, N2335, N22970);
buf BUF1 (N24436, N24432);
nand NAND3 (N24437, N24420, N3147, N5171);
and AND2 (N24438, N24434, N18500);
buf BUF1 (N24439, N24435);
or OR3 (N24440, N24423, N11233, N4856);
nand NAND2 (N24441, N24422, N9123);
or OR4 (N24442, N24438, N14955, N13118, N4349);
and AND3 (N24443, N24433, N7546, N13833);
buf BUF1 (N24444, N24440);
nand NAND2 (N24445, N24410, N9108);
not NOT1 (N24446, N24437);
nand NAND4 (N24447, N24444, N16751, N22768, N15775);
buf BUF1 (N24448, N24428);
not NOT1 (N24449, N24441);
nand NAND4 (N24450, N24436, N8849, N6653, N15209);
not NOT1 (N24451, N24442);
buf BUF1 (N24452, N24447);
and AND2 (N24453, N24424, N1539);
buf BUF1 (N24454, N24446);
not NOT1 (N24455, N24443);
and AND3 (N24456, N24452, N21775, N21314);
and AND3 (N24457, N24451, N7913, N23557);
and AND2 (N24458, N24445, N14645);
xor XOR2 (N24459, N24449, N24117);
or OR2 (N24460, N24459, N5247);
nand NAND4 (N24461, N24439, N1141, N6662, N16373);
and AND3 (N24462, N24453, N1663, N17147);
buf BUF1 (N24463, N24448);
nand NAND3 (N24464, N24456, N11535, N10157);
not NOT1 (N24465, N24454);
and AND4 (N24466, N24461, N17846, N5906, N16747);
and AND4 (N24467, N24466, N12271, N19274, N22875);
and AND2 (N24468, N24465, N7539);
nor NOR4 (N24469, N24458, N11763, N6309, N856);
nand NAND2 (N24470, N24463, N16670);
xor XOR2 (N24471, N24470, N3796);
or OR4 (N24472, N24468, N16284, N21834, N20644);
buf BUF1 (N24473, N24462);
and AND4 (N24474, N24464, N23463, N170, N19502);
not NOT1 (N24475, N24467);
or OR4 (N24476, N24457, N11454, N22754, N14532);
buf BUF1 (N24477, N24471);
buf BUF1 (N24478, N24455);
xor XOR2 (N24479, N24475, N19877);
buf BUF1 (N24480, N24478);
or OR3 (N24481, N24472, N2072, N14306);
or OR4 (N24482, N24450, N18022, N1918, N4543);
nor NOR3 (N24483, N24480, N2418, N7241);
nor NOR2 (N24484, N24476, N6528);
xor XOR2 (N24485, N24474, N352);
buf BUF1 (N24486, N24477);
nor NOR2 (N24487, N24482, N9196);
not NOT1 (N24488, N24479);
buf BUF1 (N24489, N24460);
or OR2 (N24490, N24489, N19156);
not NOT1 (N24491, N24490);
nand NAND2 (N24492, N24484, N1251);
buf BUF1 (N24493, N24473);
nor NOR2 (N24494, N24485, N19308);
or OR4 (N24495, N24487, N24211, N1065, N16386);
buf BUF1 (N24496, N24488);
or OR4 (N24497, N24469, N9269, N17266, N8851);
or OR2 (N24498, N24494, N7725);
buf BUF1 (N24499, N24492);
or OR3 (N24500, N24496, N17402, N9372);
or OR2 (N24501, N24493, N3461);
or OR4 (N24502, N24501, N13622, N11282, N8738);
xor XOR2 (N24503, N24499, N8979);
not NOT1 (N24504, N24498);
buf BUF1 (N24505, N24503);
or OR3 (N24506, N24500, N2659, N23956);
not NOT1 (N24507, N24502);
and AND2 (N24508, N24505, N9648);
buf BUF1 (N24509, N24483);
not NOT1 (N24510, N24506);
nand NAND4 (N24511, N24507, N23184, N19512, N522);
nand NAND4 (N24512, N24497, N5426, N9145, N24379);
and AND2 (N24513, N24511, N7114);
nor NOR2 (N24514, N24504, N12249);
or OR4 (N24515, N24513, N19992, N6773, N4189);
and AND2 (N24516, N24486, N3431);
not NOT1 (N24517, N24481);
and AND2 (N24518, N24491, N64);
and AND3 (N24519, N24517, N11426, N16628);
xor XOR2 (N24520, N24516, N22587);
nand NAND3 (N24521, N24519, N23315, N17823);
or OR4 (N24522, N24518, N17990, N4767, N7890);
buf BUF1 (N24523, N24510);
nor NOR2 (N24524, N24515, N3130);
or OR2 (N24525, N24508, N6240);
and AND4 (N24526, N24524, N3658, N21468, N1427);
nand NAND2 (N24527, N24521, N6199);
nor NOR2 (N24528, N24527, N5998);
or OR4 (N24529, N24514, N13878, N11336, N2171);
or OR4 (N24530, N24528, N20588, N14834, N8559);
nand NAND2 (N24531, N24529, N842);
nand NAND3 (N24532, N24520, N12734, N18110);
xor XOR2 (N24533, N24522, N21538);
buf BUF1 (N24534, N24532);
xor XOR2 (N24535, N24512, N20719);
or OR2 (N24536, N24523, N12468);
not NOT1 (N24537, N24530);
or OR3 (N24538, N24525, N3989, N359);
buf BUF1 (N24539, N24536);
or OR2 (N24540, N24539, N21784);
buf BUF1 (N24541, N24526);
and AND2 (N24542, N24538, N15111);
not NOT1 (N24543, N24534);
not NOT1 (N24544, N24533);
not NOT1 (N24545, N24495);
or OR4 (N24546, N24540, N14517, N12409, N11283);
not NOT1 (N24547, N24546);
buf BUF1 (N24548, N24544);
and AND3 (N24549, N24531, N19690, N12295);
buf BUF1 (N24550, N24537);
nand NAND2 (N24551, N24543, N14423);
nor NOR2 (N24552, N24547, N17153);
buf BUF1 (N24553, N24535);
or OR3 (N24554, N24509, N21750, N9702);
or OR4 (N24555, N24550, N22379, N19148, N16366);
not NOT1 (N24556, N24553);
xor XOR2 (N24557, N24542, N23179);
buf BUF1 (N24558, N24541);
or OR4 (N24559, N24554, N2829, N16771, N20480);
or OR2 (N24560, N24555, N7302);
xor XOR2 (N24561, N24558, N11622);
nor NOR4 (N24562, N24552, N16073, N5424, N23004);
and AND3 (N24563, N24549, N2277, N18754);
not NOT1 (N24564, N24561);
and AND2 (N24565, N24556, N1349);
not NOT1 (N24566, N24557);
nand NAND2 (N24567, N24560, N18463);
nor NOR4 (N24568, N24567, N7149, N11510, N22760);
buf BUF1 (N24569, N24562);
nand NAND4 (N24570, N24568, N3788, N20056, N5824);
and AND2 (N24571, N24548, N11890);
nand NAND3 (N24572, N24571, N899, N12715);
nand NAND4 (N24573, N24559, N11859, N1703, N13241);
nand NAND2 (N24574, N24564, N22734);
buf BUF1 (N24575, N24572);
and AND2 (N24576, N24566, N21153);
nor NOR3 (N24577, N24569, N23174, N15806);
xor XOR2 (N24578, N24565, N23454);
not NOT1 (N24579, N24570);
nand NAND2 (N24580, N24551, N10827);
xor XOR2 (N24581, N24574, N9391);
nand NAND4 (N24582, N24580, N22448, N7278, N11384);
xor XOR2 (N24583, N24577, N23654);
xor XOR2 (N24584, N24581, N14773);
or OR2 (N24585, N24578, N6474);
not NOT1 (N24586, N24573);
and AND4 (N24587, N24582, N15392, N9121, N23397);
and AND2 (N24588, N24587, N16469);
and AND2 (N24589, N24585, N854);
nand NAND2 (N24590, N24588, N20916);
xor XOR2 (N24591, N24563, N14221);
or OR4 (N24592, N24590, N3672, N5490, N5239);
nand NAND4 (N24593, N24584, N19412, N6744, N20281);
not NOT1 (N24594, N24592);
xor XOR2 (N24595, N24589, N20499);
or OR3 (N24596, N24591, N22423, N13998);
nor NOR3 (N24597, N24575, N23389, N16090);
and AND4 (N24598, N24595, N17364, N1361, N18980);
or OR3 (N24599, N24583, N10964, N20553);
not NOT1 (N24600, N24586);
nand NAND4 (N24601, N24597, N17017, N12584, N5254);
xor XOR2 (N24602, N24545, N9984);
not NOT1 (N24603, N24579);
and AND4 (N24604, N24593, N21092, N2686, N20490);
not NOT1 (N24605, N24600);
nand NAND2 (N24606, N24603, N9201);
buf BUF1 (N24607, N24602);
nand NAND4 (N24608, N24599, N24194, N1956, N3803);
buf BUF1 (N24609, N24604);
or OR3 (N24610, N24605, N10895, N4439);
xor XOR2 (N24611, N24608, N841);
not NOT1 (N24612, N24576);
xor XOR2 (N24613, N24598, N22841);
and AND4 (N24614, N24610, N18629, N9574, N18486);
xor XOR2 (N24615, N24611, N21799);
or OR3 (N24616, N24615, N23939, N651);
xor XOR2 (N24617, N24606, N1732);
and AND2 (N24618, N24609, N18927);
nand NAND3 (N24619, N24614, N12600, N5177);
nor NOR4 (N24620, N24619, N1856, N7792, N23322);
nand NAND3 (N24621, N24601, N11167, N10043);
buf BUF1 (N24622, N24613);
or OR3 (N24623, N24596, N2813, N10759);
buf BUF1 (N24624, N24622);
nor NOR2 (N24625, N24616, N21123);
nor NOR3 (N24626, N24623, N18937, N7684);
nand NAND2 (N24627, N24625, N1469);
and AND4 (N24628, N24612, N20909, N23272, N7472);
nor NOR3 (N24629, N24626, N16457, N6244);
or OR3 (N24630, N24620, N11636, N18592);
and AND3 (N24631, N24621, N21088, N14843);
or OR2 (N24632, N24617, N7376);
nand NAND3 (N24633, N24630, N11414, N19793);
or OR2 (N24634, N24631, N22758);
not NOT1 (N24635, N24632);
and AND3 (N24636, N24607, N15157, N360);
and AND2 (N24637, N24594, N7065);
or OR3 (N24638, N24637, N5558, N3052);
not NOT1 (N24639, N24635);
or OR4 (N24640, N24627, N16891, N14407, N20769);
or OR4 (N24641, N24638, N10833, N8309, N2565);
nor NOR3 (N24642, N24624, N9724, N6581);
xor XOR2 (N24643, N24629, N22490);
nor NOR2 (N24644, N24639, N7616);
or OR3 (N24645, N24628, N13120, N1805);
or OR4 (N24646, N24634, N18304, N5391, N17064);
or OR2 (N24647, N24636, N550);
or OR3 (N24648, N24647, N244, N12577);
nand NAND3 (N24649, N24646, N15571, N435);
not NOT1 (N24650, N24648);
and AND3 (N24651, N24641, N3246, N12423);
nand NAND3 (N24652, N24633, N17795, N2967);
buf BUF1 (N24653, N24651);
buf BUF1 (N24654, N24645);
xor XOR2 (N24655, N24642, N24116);
not NOT1 (N24656, N24644);
nor NOR4 (N24657, N24656, N12724, N2325, N10179);
nor NOR3 (N24658, N24643, N1212, N663);
buf BUF1 (N24659, N24618);
xor XOR2 (N24660, N24653, N20126);
nor NOR2 (N24661, N24650, N15845);
not NOT1 (N24662, N24652);
buf BUF1 (N24663, N24640);
or OR3 (N24664, N24661, N15434, N22928);
or OR3 (N24665, N24654, N11496, N11623);
nor NOR3 (N24666, N24662, N10611, N7863);
nor NOR3 (N24667, N24663, N5344, N20219);
or OR3 (N24668, N24658, N2013, N13421);
and AND4 (N24669, N24666, N3598, N18853, N19825);
nor NOR2 (N24670, N24655, N13756);
not NOT1 (N24671, N24668);
xor XOR2 (N24672, N24659, N16686);
or OR3 (N24673, N24665, N21121, N16258);
xor XOR2 (N24674, N24669, N19657);
not NOT1 (N24675, N24649);
not NOT1 (N24676, N24673);
and AND3 (N24677, N24674, N16898, N6828);
xor XOR2 (N24678, N24675, N20936);
or OR2 (N24679, N24664, N14431);
and AND3 (N24680, N24671, N19079, N16184);
and AND2 (N24681, N24660, N9946);
xor XOR2 (N24682, N24677, N284);
not NOT1 (N24683, N24672);
buf BUF1 (N24684, N24679);
and AND2 (N24685, N24683, N5729);
and AND2 (N24686, N24682, N15842);
not NOT1 (N24687, N24667);
xor XOR2 (N24688, N24687, N22312);
xor XOR2 (N24689, N24688, N2490);
or OR2 (N24690, N24686, N18246);
xor XOR2 (N24691, N24657, N11916);
and AND4 (N24692, N24690, N15607, N4886, N5837);
buf BUF1 (N24693, N24691);
xor XOR2 (N24694, N24692, N20824);
nand NAND4 (N24695, N24681, N18363, N10476, N16515);
nand NAND4 (N24696, N24680, N22239, N13041, N680);
buf BUF1 (N24697, N24696);
nor NOR4 (N24698, N24695, N15028, N22262, N9062);
xor XOR2 (N24699, N24697, N10615);
buf BUF1 (N24700, N24685);
buf BUF1 (N24701, N24689);
and AND2 (N24702, N24676, N8848);
or OR3 (N24703, N24678, N12068, N17792);
or OR4 (N24704, N24670, N3153, N5981, N24310);
or OR2 (N24705, N24700, N20467);
not NOT1 (N24706, N24699);
nor NOR2 (N24707, N24694, N8017);
nand NAND2 (N24708, N24704, N184);
nor NOR3 (N24709, N24684, N1219, N5685);
nor NOR2 (N24710, N24703, N12459);
not NOT1 (N24711, N24707);
and AND4 (N24712, N24693, N126, N15887, N20685);
xor XOR2 (N24713, N24710, N15933);
xor XOR2 (N24714, N24713, N7884);
or OR3 (N24715, N24698, N5037, N23407);
or OR4 (N24716, N24706, N10440, N12698, N19316);
not NOT1 (N24717, N24711);
nand NAND4 (N24718, N24715, N19030, N13385, N10921);
not NOT1 (N24719, N24716);
nor NOR2 (N24720, N24719, N2241);
and AND3 (N24721, N24702, N9894, N21889);
or OR3 (N24722, N24720, N6312, N17127);
nand NAND3 (N24723, N24712, N3095, N22981);
nor NOR4 (N24724, N24708, N93, N5500, N2718);
or OR4 (N24725, N24723, N296, N8390, N19359);
nand NAND2 (N24726, N24709, N7560);
buf BUF1 (N24727, N24705);
or OR3 (N24728, N24724, N21769, N2108);
nor NOR4 (N24729, N24728, N9359, N16982, N4787);
or OR4 (N24730, N24725, N22240, N8833, N24086);
buf BUF1 (N24731, N24721);
or OR3 (N24732, N24722, N10225, N21060);
buf BUF1 (N24733, N24730);
xor XOR2 (N24734, N24727, N8184);
not NOT1 (N24735, N24734);
nor NOR4 (N24736, N24731, N14372, N14686, N12534);
and AND3 (N24737, N24701, N3843, N758);
nand NAND4 (N24738, N24733, N4313, N23457, N14874);
and AND4 (N24739, N24735, N21578, N12462, N4882);
not NOT1 (N24740, N24718);
nand NAND3 (N24741, N24717, N19162, N10012);
nor NOR2 (N24742, N24714, N17435);
nor NOR4 (N24743, N24741, N5827, N10562, N8146);
and AND4 (N24744, N24740, N12292, N17527, N11938);
buf BUF1 (N24745, N24737);
not NOT1 (N24746, N24736);
buf BUF1 (N24747, N24745);
nor NOR4 (N24748, N24726, N8915, N22953, N7698);
or OR3 (N24749, N24738, N8864, N22734);
or OR4 (N24750, N24749, N9383, N19742, N9037);
nand NAND4 (N24751, N24739, N17584, N1826, N6159);
not NOT1 (N24752, N24746);
nand NAND2 (N24753, N24750, N7821);
nand NAND4 (N24754, N24751, N496, N16582, N16459);
xor XOR2 (N24755, N24742, N16320);
buf BUF1 (N24756, N24729);
not NOT1 (N24757, N24755);
and AND3 (N24758, N24743, N6004, N17506);
or OR3 (N24759, N24757, N5757, N10190);
xor XOR2 (N24760, N24759, N3544);
xor XOR2 (N24761, N24752, N13165);
nor NOR4 (N24762, N24754, N22440, N15617, N18917);
nor NOR3 (N24763, N24748, N5476, N17701);
and AND4 (N24764, N24732, N13709, N8035, N15556);
xor XOR2 (N24765, N24760, N5199);
nand NAND4 (N24766, N24753, N12652, N23102, N21537);
nor NOR4 (N24767, N24766, N18699, N10564, N14486);
and AND4 (N24768, N24765, N12427, N21555, N2071);
and AND3 (N24769, N24768, N12200, N6872);
and AND3 (N24770, N24747, N22919, N6360);
or OR2 (N24771, N24761, N16322);
nand NAND2 (N24772, N24764, N22262);
xor XOR2 (N24773, N24771, N1207);
xor XOR2 (N24774, N24770, N8066);
xor XOR2 (N24775, N24763, N13120);
nand NAND4 (N24776, N24775, N2933, N7622, N13255);
and AND2 (N24777, N24758, N2916);
and AND2 (N24778, N24756, N1009);
nand NAND2 (N24779, N24772, N23961);
xor XOR2 (N24780, N24779, N14298);
nand NAND4 (N24781, N24780, N18530, N23441, N8827);
buf BUF1 (N24782, N24767);
or OR3 (N24783, N24776, N865, N10847);
xor XOR2 (N24784, N24774, N12804);
and AND4 (N24785, N24777, N3341, N1078, N4418);
nor NOR4 (N24786, N24783, N2952, N360, N19114);
buf BUF1 (N24787, N24773);
or OR2 (N24788, N24785, N1585);
nor NOR4 (N24789, N24769, N13601, N1453, N12090);
xor XOR2 (N24790, N24781, N4249);
buf BUF1 (N24791, N24787);
xor XOR2 (N24792, N24786, N6653);
not NOT1 (N24793, N24744);
not NOT1 (N24794, N24778);
buf BUF1 (N24795, N24791);
nor NOR4 (N24796, N24762, N18974, N6473, N3691);
buf BUF1 (N24797, N24790);
nand NAND3 (N24798, N24789, N5081, N7326);
nand NAND3 (N24799, N24782, N18680, N12161);
buf BUF1 (N24800, N24795);
or OR2 (N24801, N24788, N13702);
nand NAND3 (N24802, N24796, N21926, N17096);
or OR4 (N24803, N24797, N12083, N8617, N6781);
and AND4 (N24804, N24784, N22564, N14644, N2848);
not NOT1 (N24805, N24792);
and AND3 (N24806, N24794, N1733, N19284);
nand NAND4 (N24807, N24801, N2545, N22866, N18182);
or OR4 (N24808, N24793, N5915, N17992, N18715);
not NOT1 (N24809, N24804);
and AND3 (N24810, N24806, N11967, N2614);
nor NOR3 (N24811, N24800, N24316, N13013);
nor NOR4 (N24812, N24810, N3422, N9746, N10472);
xor XOR2 (N24813, N24812, N18945);
or OR4 (N24814, N24799, N503, N3633, N18824);
or OR2 (N24815, N24807, N1181);
and AND3 (N24816, N24808, N10611, N9171);
xor XOR2 (N24817, N24811, N531);
xor XOR2 (N24818, N24798, N12068);
nand NAND3 (N24819, N24817, N13385, N22118);
or OR2 (N24820, N24803, N4179);
buf BUF1 (N24821, N24813);
nand NAND3 (N24822, N24821, N11482, N5365);
not NOT1 (N24823, N24819);
not NOT1 (N24824, N24815);
xor XOR2 (N24825, N24824, N6716);
or OR2 (N24826, N24814, N3167);
buf BUF1 (N24827, N24802);
xor XOR2 (N24828, N24827, N6233);
buf BUF1 (N24829, N24822);
and AND2 (N24830, N24826, N15684);
or OR2 (N24831, N24823, N4876);
and AND4 (N24832, N24805, N23213, N13006, N7728);
not NOT1 (N24833, N24829);
xor XOR2 (N24834, N24809, N15261);
buf BUF1 (N24835, N24833);
and AND4 (N24836, N24831, N24583, N15884, N4828);
buf BUF1 (N24837, N24828);
or OR3 (N24838, N24816, N7271, N20448);
nor NOR2 (N24839, N24825, N9493);
xor XOR2 (N24840, N24820, N2036);
nor NOR3 (N24841, N24834, N12937, N5476);
nand NAND2 (N24842, N24830, N4286);
nand NAND4 (N24843, N24837, N4448, N19352, N21562);
nor NOR2 (N24844, N24843, N7572);
xor XOR2 (N24845, N24836, N18088);
xor XOR2 (N24846, N24840, N23040);
or OR2 (N24847, N24846, N20126);
buf BUF1 (N24848, N24844);
not NOT1 (N24849, N24835);
not NOT1 (N24850, N24845);
buf BUF1 (N24851, N24839);
nand NAND3 (N24852, N24832, N16674, N11519);
nand NAND4 (N24853, N24838, N15492, N3503, N21645);
not NOT1 (N24854, N24848);
not NOT1 (N24855, N24818);
and AND3 (N24856, N24842, N1221, N1430);
nand NAND2 (N24857, N24847, N7532);
not NOT1 (N24858, N24855);
buf BUF1 (N24859, N24853);
and AND3 (N24860, N24856, N6742, N11893);
nand NAND4 (N24861, N24858, N2015, N4131, N1942);
not NOT1 (N24862, N24861);
nor NOR2 (N24863, N24854, N2411);
xor XOR2 (N24864, N24863, N17419);
xor XOR2 (N24865, N24862, N2669);
or OR4 (N24866, N24849, N2330, N8381, N8632);
nand NAND4 (N24867, N24860, N21211, N4177, N18582);
and AND4 (N24868, N24857, N17085, N8960, N21322);
xor XOR2 (N24869, N24850, N24770);
and AND4 (N24870, N24852, N14593, N12082, N3456);
buf BUF1 (N24871, N24869);
and AND2 (N24872, N24870, N14366);
not NOT1 (N24873, N24871);
and AND2 (N24874, N24868, N6725);
xor XOR2 (N24875, N24841, N16422);
or OR3 (N24876, N24874, N1194, N19096);
or OR4 (N24877, N24875, N8941, N3831, N21061);
or OR3 (N24878, N24865, N3044, N15897);
nor NOR3 (N24879, N24873, N23893, N24424);
buf BUF1 (N24880, N24864);
xor XOR2 (N24881, N24877, N10912);
nand NAND4 (N24882, N24859, N6316, N1109, N20734);
xor XOR2 (N24883, N24879, N8645);
or OR3 (N24884, N24882, N18335, N7656);
and AND2 (N24885, N24881, N13020);
or OR4 (N24886, N24851, N15030, N7895, N10488);
or OR4 (N24887, N24872, N9057, N4108, N20254);
or OR2 (N24888, N24887, N3289);
xor XOR2 (N24889, N24880, N1553);
buf BUF1 (N24890, N24867);
and AND4 (N24891, N24876, N1168, N11434, N2018);
buf BUF1 (N24892, N24890);
and AND3 (N24893, N24884, N23378, N4070);
or OR3 (N24894, N24891, N2262, N15632);
not NOT1 (N24895, N24883);
nand NAND3 (N24896, N24886, N22999, N12082);
nor NOR2 (N24897, N24895, N3798);
and AND2 (N24898, N24897, N24582);
nor NOR2 (N24899, N24889, N15901);
nand NAND4 (N24900, N24885, N14830, N8707, N18996);
buf BUF1 (N24901, N24892);
not NOT1 (N24902, N24901);
buf BUF1 (N24903, N24893);
and AND2 (N24904, N24902, N14680);
xor XOR2 (N24905, N24878, N12011);
and AND3 (N24906, N24905, N17817, N12295);
nor NOR2 (N24907, N24900, N5271);
nor NOR3 (N24908, N24866, N4955, N23951);
buf BUF1 (N24909, N24896);
xor XOR2 (N24910, N24903, N5322);
not NOT1 (N24911, N24904);
buf BUF1 (N24912, N24894);
xor XOR2 (N24913, N24912, N1618);
xor XOR2 (N24914, N24907, N3793);
not NOT1 (N24915, N24914);
xor XOR2 (N24916, N24888, N5003);
or OR2 (N24917, N24915, N3062);
xor XOR2 (N24918, N24909, N4231);
or OR4 (N24919, N24898, N3238, N1769, N9086);
nor NOR3 (N24920, N24913, N9349, N4842);
or OR2 (N24921, N24920, N9861);
nor NOR3 (N24922, N24917, N17385, N13419);
nand NAND4 (N24923, N24916, N2989, N9494, N19159);
not NOT1 (N24924, N24918);
not NOT1 (N24925, N24911);
xor XOR2 (N24926, N24899, N19062);
and AND4 (N24927, N24923, N8728, N22387, N18545);
xor XOR2 (N24928, N24926, N964);
buf BUF1 (N24929, N24906);
nor NOR4 (N24930, N24928, N4747, N4031, N13894);
nand NAND4 (N24931, N24924, N4498, N5841, N17859);
and AND4 (N24932, N24910, N1863, N2512, N16410);
and AND4 (N24933, N24927, N15144, N1802, N18755);
xor XOR2 (N24934, N24929, N21640);
nor NOR3 (N24935, N24922, N6408, N1809);
xor XOR2 (N24936, N24932, N10755);
or OR3 (N24937, N24934, N3529, N13965);
buf BUF1 (N24938, N24933);
xor XOR2 (N24939, N24931, N11735);
nor NOR2 (N24940, N24936, N8229);
nor NOR2 (N24941, N24935, N23239);
nand NAND4 (N24942, N24940, N20095, N14566, N12318);
not NOT1 (N24943, N24937);
or OR2 (N24944, N24939, N15086);
nand NAND3 (N24945, N24941, N13763, N5402);
buf BUF1 (N24946, N24908);
buf BUF1 (N24947, N24921);
xor XOR2 (N24948, N24947, N7026);
or OR2 (N24949, N24942, N14171);
not NOT1 (N24950, N24944);
buf BUF1 (N24951, N24925);
xor XOR2 (N24952, N24938, N6905);
not NOT1 (N24953, N24946);
not NOT1 (N24954, N24951);
xor XOR2 (N24955, N24945, N2636);
or OR2 (N24956, N24930, N8836);
and AND2 (N24957, N24943, N20712);
nor NOR2 (N24958, N24954, N10235);
nand NAND4 (N24959, N24950, N18939, N16569, N18247);
xor XOR2 (N24960, N24948, N3107);
or OR3 (N24961, N24952, N12143, N7586);
not NOT1 (N24962, N24957);
nand NAND4 (N24963, N24949, N22172, N3012, N8676);
xor XOR2 (N24964, N24955, N15549);
nor NOR2 (N24965, N24959, N17335);
nand NAND4 (N24966, N24962, N23947, N14194, N17326);
nand NAND4 (N24967, N24965, N9960, N20442, N22767);
nand NAND2 (N24968, N24956, N18191);
not NOT1 (N24969, N24960);
and AND4 (N24970, N24958, N16683, N1903, N15625);
nor NOR3 (N24971, N24966, N8446, N8888);
not NOT1 (N24972, N24919);
not NOT1 (N24973, N24964);
not NOT1 (N24974, N24972);
buf BUF1 (N24975, N24961);
buf BUF1 (N24976, N24969);
not NOT1 (N24977, N24973);
not NOT1 (N24978, N24976);
or OR4 (N24979, N24970, N1532, N30, N22903);
nand NAND4 (N24980, N24967, N18625, N22651, N16128);
buf BUF1 (N24981, N24980);
buf BUF1 (N24982, N24971);
nor NOR4 (N24983, N24974, N16780, N6698, N4572);
buf BUF1 (N24984, N24968);
buf BUF1 (N24985, N24953);
not NOT1 (N24986, N24982);
buf BUF1 (N24987, N24983);
not NOT1 (N24988, N24984);
not NOT1 (N24989, N24979);
not NOT1 (N24990, N24989);
and AND4 (N24991, N24988, N19090, N22890, N22193);
nor NOR4 (N24992, N24986, N24242, N20066, N21417);
or OR3 (N24993, N24987, N12273, N22572);
and AND2 (N24994, N24993, N17614);
buf BUF1 (N24995, N24992);
buf BUF1 (N24996, N24963);
and AND2 (N24997, N24981, N177);
or OR2 (N24998, N24977, N6899);
xor XOR2 (N24999, N24991, N9657);
buf BUF1 (N25000, N24975);
xor XOR2 (N25001, N24998, N5367);
and AND3 (N25002, N24995, N1866, N6999);
nor NOR2 (N25003, N24996, N12809);
nor NOR3 (N25004, N24997, N16993, N2880);
or OR2 (N25005, N24994, N23706);
buf BUF1 (N25006, N25002);
xor XOR2 (N25007, N24985, N11554);
and AND2 (N25008, N24990, N11157);
nor NOR2 (N25009, N24978, N6893);
not NOT1 (N25010, N25007);
or OR4 (N25011, N25006, N1123, N20441, N17484);
not NOT1 (N25012, N25008);
not NOT1 (N25013, N25004);
and AND4 (N25014, N25013, N10391, N17634, N3049);
not NOT1 (N25015, N25003);
xor XOR2 (N25016, N25011, N15898);
and AND4 (N25017, N25015, N2182, N9749, N17680);
not NOT1 (N25018, N25012);
and AND3 (N25019, N25017, N155, N6999);
buf BUF1 (N25020, N25014);
nand NAND3 (N25021, N25010, N2596, N194);
or OR3 (N25022, N25019, N10488, N23655);
or OR4 (N25023, N24999, N3981, N14080, N4581);
or OR3 (N25024, N25009, N9827, N6524);
xor XOR2 (N25025, N25016, N7384);
and AND2 (N25026, N25000, N6982);
buf BUF1 (N25027, N25020);
or OR3 (N25028, N25024, N10426, N7126);
not NOT1 (N25029, N25018);
not NOT1 (N25030, N25023);
nand NAND2 (N25031, N25025, N13444);
or OR4 (N25032, N25028, N6320, N19977, N11787);
nor NOR2 (N25033, N25032, N9524);
or OR2 (N25034, N25029, N17412);
xor XOR2 (N25035, N25022, N16381);
xor XOR2 (N25036, N25026, N2604);
or OR4 (N25037, N25031, N5383, N11758, N284);
and AND4 (N25038, N25001, N13063, N21253, N10365);
buf BUF1 (N25039, N25037);
buf BUF1 (N25040, N25005);
not NOT1 (N25041, N25035);
xor XOR2 (N25042, N25038, N6076);
not NOT1 (N25043, N25036);
nand NAND2 (N25044, N25030, N15145);
or OR4 (N25045, N25027, N13250, N19682, N17165);
nand NAND3 (N25046, N25044, N14927, N21747);
not NOT1 (N25047, N25034);
or OR2 (N25048, N25021, N732);
xor XOR2 (N25049, N25040, N10003);
or OR2 (N25050, N25046, N8243);
and AND4 (N25051, N25042, N6897, N6648, N14926);
xor XOR2 (N25052, N25041, N5160);
nor NOR3 (N25053, N25048, N12085, N9766);
xor XOR2 (N25054, N25049, N4830);
xor XOR2 (N25055, N25053, N17612);
not NOT1 (N25056, N25052);
nor NOR4 (N25057, N25047, N22798, N9923, N2214);
nor NOR3 (N25058, N25055, N13988, N3657);
buf BUF1 (N25059, N25057);
buf BUF1 (N25060, N25059);
xor XOR2 (N25061, N25056, N19632);
or OR3 (N25062, N25051, N1976, N15146);
not NOT1 (N25063, N25045);
buf BUF1 (N25064, N25060);
or OR4 (N25065, N25054, N11997, N10256, N4297);
or OR2 (N25066, N25039, N6494);
not NOT1 (N25067, N25063);
xor XOR2 (N25068, N25061, N4221);
buf BUF1 (N25069, N25068);
or OR2 (N25070, N25050, N18814);
and AND4 (N25071, N25067, N20362, N16297, N7530);
nand NAND4 (N25072, N25066, N22557, N3054, N17606);
nor NOR4 (N25073, N25071, N11332, N24577, N14824);
not NOT1 (N25074, N25043);
nor NOR4 (N25075, N25072, N6642, N6102, N3955);
buf BUF1 (N25076, N25064);
nand NAND4 (N25077, N25074, N9714, N16635, N10838);
buf BUF1 (N25078, N25076);
nand NAND4 (N25079, N25070, N14524, N12298, N21166);
nand NAND3 (N25080, N25069, N24838, N22251);
xor XOR2 (N25081, N25065, N18995);
or OR2 (N25082, N25033, N446);
nor NOR4 (N25083, N25062, N15735, N23473, N11459);
not NOT1 (N25084, N25081);
not NOT1 (N25085, N25084);
and AND4 (N25086, N25058, N22520, N21707, N16404);
and AND2 (N25087, N25075, N3743);
and AND2 (N25088, N25087, N5540);
xor XOR2 (N25089, N25073, N9116);
nand NAND2 (N25090, N25086, N18974);
nand NAND3 (N25091, N25088, N3527, N21183);
or OR3 (N25092, N25082, N11506, N3312);
or OR4 (N25093, N25091, N4552, N19338, N1732);
not NOT1 (N25094, N25083);
buf BUF1 (N25095, N25079);
nand NAND4 (N25096, N25077, N12624, N738, N19648);
not NOT1 (N25097, N25085);
nor NOR2 (N25098, N25090, N12945);
buf BUF1 (N25099, N25098);
nor NOR4 (N25100, N25093, N15290, N22853, N20701);
not NOT1 (N25101, N25095);
or OR2 (N25102, N25080, N9787);
or OR3 (N25103, N25096, N502, N7374);
xor XOR2 (N25104, N25102, N8494);
nor NOR3 (N25105, N25104, N13253, N12125);
buf BUF1 (N25106, N25099);
or OR3 (N25107, N25105, N4838, N3972);
nand NAND3 (N25108, N25089, N12558, N11186);
nand NAND4 (N25109, N25100, N15142, N14533, N3561);
nand NAND3 (N25110, N25109, N20535, N22706);
and AND4 (N25111, N25094, N5306, N8212, N17925);
and AND2 (N25112, N25107, N7214);
and AND3 (N25113, N25106, N535, N5381);
nor NOR2 (N25114, N25103, N15079);
buf BUF1 (N25115, N25113);
xor XOR2 (N25116, N25097, N8402);
buf BUF1 (N25117, N25111);
or OR3 (N25118, N25078, N6432, N21060);
xor XOR2 (N25119, N25115, N22840);
or OR4 (N25120, N25119, N17188, N5689, N21193);
buf BUF1 (N25121, N25117);
nand NAND4 (N25122, N25121, N12006, N12135, N8486);
nor NOR4 (N25123, N25122, N7095, N17680, N7582);
buf BUF1 (N25124, N25120);
buf BUF1 (N25125, N25110);
not NOT1 (N25126, N25118);
xor XOR2 (N25127, N25112, N274);
and AND2 (N25128, N25108, N13529);
or OR3 (N25129, N25092, N23539, N828);
buf BUF1 (N25130, N25126);
not NOT1 (N25131, N25128);
buf BUF1 (N25132, N25131);
not NOT1 (N25133, N25129);
nor NOR2 (N25134, N25101, N2561);
or OR2 (N25135, N25127, N15720);
nand NAND4 (N25136, N25130, N24497, N250, N7958);
or OR2 (N25137, N25123, N9842);
nor NOR3 (N25138, N25124, N1939, N3368);
nand NAND2 (N25139, N25132, N7859);
buf BUF1 (N25140, N25138);
buf BUF1 (N25141, N25133);
nor NOR3 (N25142, N25140, N20398, N9116);
xor XOR2 (N25143, N25141, N15036);
nand NAND2 (N25144, N25114, N6910);
and AND2 (N25145, N25142, N19060);
not NOT1 (N25146, N25144);
and AND3 (N25147, N25116, N6987, N3348);
nor NOR3 (N25148, N25137, N6092, N12646);
or OR2 (N25149, N25135, N2655);
not NOT1 (N25150, N25134);
or OR3 (N25151, N25136, N1039, N22478);
and AND4 (N25152, N25148, N13553, N23045, N10775);
nor NOR4 (N25153, N25146, N8924, N23115, N2023);
nor NOR4 (N25154, N25151, N19759, N22069, N14849);
or OR4 (N25155, N25150, N21699, N7252, N16887);
and AND3 (N25156, N25139, N22323, N16702);
nor NOR3 (N25157, N25145, N2746, N11);
and AND2 (N25158, N25155, N18878);
or OR2 (N25159, N25149, N21214);
not NOT1 (N25160, N25157);
buf BUF1 (N25161, N25147);
or OR2 (N25162, N25158, N14223);
nand NAND4 (N25163, N25152, N11202, N4223, N12397);
not NOT1 (N25164, N25125);
and AND3 (N25165, N25160, N22831, N21295);
and AND3 (N25166, N25162, N3371, N17004);
nand NAND2 (N25167, N25164, N15025);
and AND2 (N25168, N25166, N23020);
or OR4 (N25169, N25163, N7654, N3195, N14922);
buf BUF1 (N25170, N25168);
and AND4 (N25171, N25154, N24837, N5994, N8085);
xor XOR2 (N25172, N25161, N23123);
or OR3 (N25173, N25159, N15179, N18502);
or OR4 (N25174, N25173, N6425, N15365, N8531);
buf BUF1 (N25175, N25143);
xor XOR2 (N25176, N25170, N24897);
and AND4 (N25177, N25175, N2170, N10733, N22747);
nor NOR3 (N25178, N25174, N24289, N13359);
and AND4 (N25179, N25165, N19147, N5293, N5109);
nor NOR2 (N25180, N25167, N1325);
xor XOR2 (N25181, N25176, N1472);
and AND3 (N25182, N25169, N16581, N13747);
and AND4 (N25183, N25182, N14367, N15509, N18229);
and AND2 (N25184, N25171, N15221);
or OR2 (N25185, N25177, N14850);
not NOT1 (N25186, N25183);
or OR2 (N25187, N25180, N17804);
not NOT1 (N25188, N25156);
not NOT1 (N25189, N25153);
buf BUF1 (N25190, N25189);
buf BUF1 (N25191, N25178);
not NOT1 (N25192, N25190);
nand NAND4 (N25193, N25172, N22692, N13388, N11544);
nor NOR4 (N25194, N25193, N7966, N23323, N5060);
nand NAND2 (N25195, N25186, N5734);
or OR4 (N25196, N25179, N16079, N22329, N8251);
not NOT1 (N25197, N25192);
and AND3 (N25198, N25181, N2336, N9347);
and AND4 (N25199, N25196, N9636, N20308, N22968);
or OR2 (N25200, N25184, N9456);
not NOT1 (N25201, N25187);
xor XOR2 (N25202, N25197, N21869);
nor NOR4 (N25203, N25202, N7255, N5296, N17847);
or OR4 (N25204, N25200, N5652, N145, N6754);
xor XOR2 (N25205, N25194, N25191);
not NOT1 (N25206, N3716);
and AND2 (N25207, N25204, N9228);
buf BUF1 (N25208, N25185);
or OR4 (N25209, N25195, N9911, N13242, N15921);
buf BUF1 (N25210, N25208);
or OR3 (N25211, N25206, N5522, N7908);
or OR4 (N25212, N25209, N9559, N4323, N24048);
not NOT1 (N25213, N25201);
and AND2 (N25214, N25207, N13226);
xor XOR2 (N25215, N25212, N19202);
nand NAND2 (N25216, N25205, N14595);
not NOT1 (N25217, N25199);
nor NOR2 (N25218, N25188, N22148);
buf BUF1 (N25219, N25214);
not NOT1 (N25220, N25218);
buf BUF1 (N25221, N25215);
buf BUF1 (N25222, N25203);
xor XOR2 (N25223, N25210, N15972);
nand NAND3 (N25224, N25217, N16501, N415);
nand NAND3 (N25225, N25222, N11329, N467);
or OR2 (N25226, N25198, N18477);
xor XOR2 (N25227, N25220, N306);
and AND2 (N25228, N25213, N20184);
buf BUF1 (N25229, N25211);
buf BUF1 (N25230, N25227);
buf BUF1 (N25231, N25224);
buf BUF1 (N25232, N25226);
or OR4 (N25233, N25216, N4497, N15538, N524);
buf BUF1 (N25234, N25228);
and AND4 (N25235, N25221, N19525, N21256, N1832);
and AND3 (N25236, N25223, N10149, N16694);
nor NOR3 (N25237, N25233, N20054, N17676);
or OR3 (N25238, N25230, N16670, N20765);
xor XOR2 (N25239, N25234, N5758);
not NOT1 (N25240, N25219);
or OR2 (N25241, N25225, N24930);
xor XOR2 (N25242, N25229, N6442);
buf BUF1 (N25243, N25238);
nor NOR2 (N25244, N25236, N13956);
nor NOR3 (N25245, N25237, N12959, N23798);
nor NOR4 (N25246, N25239, N24491, N12147, N25062);
not NOT1 (N25247, N25242);
nor NOR4 (N25248, N25245, N10259, N20916, N9587);
buf BUF1 (N25249, N25244);
or OR4 (N25250, N25241, N19170, N16348, N5030);
nand NAND4 (N25251, N25240, N23072, N5855, N21576);
not NOT1 (N25252, N25232);
buf BUF1 (N25253, N25243);
and AND3 (N25254, N25235, N18442, N4584);
nand NAND4 (N25255, N25252, N4638, N12286, N8697);
nor NOR3 (N25256, N25246, N12876, N24042);
nand NAND2 (N25257, N25247, N20527);
nand NAND3 (N25258, N25256, N21472, N5744);
xor XOR2 (N25259, N25253, N2885);
buf BUF1 (N25260, N25254);
nor NOR4 (N25261, N25258, N24474, N17952, N13688);
and AND2 (N25262, N25261, N22314);
nand NAND2 (N25263, N25257, N12270);
or OR3 (N25264, N25255, N23616, N15333);
not NOT1 (N25265, N25264);
and AND4 (N25266, N25250, N21035, N21861, N24216);
nand NAND3 (N25267, N25231, N8617, N8075);
or OR2 (N25268, N25262, N7874);
or OR4 (N25269, N25265, N9733, N17840, N22529);
or OR4 (N25270, N25249, N6500, N18075, N5491);
nor NOR3 (N25271, N25248, N8779, N616);
and AND3 (N25272, N25266, N121, N15751);
not NOT1 (N25273, N25260);
or OR3 (N25274, N25273, N10958, N5258);
nand NAND2 (N25275, N25274, N4973);
not NOT1 (N25276, N25268);
not NOT1 (N25277, N25270);
not NOT1 (N25278, N25263);
or OR2 (N25279, N25259, N12610);
nand NAND2 (N25280, N25278, N9455);
not NOT1 (N25281, N25251);
buf BUF1 (N25282, N25280);
nor NOR4 (N25283, N25271, N10363, N5076, N24020);
nand NAND2 (N25284, N25275, N19291);
buf BUF1 (N25285, N25284);
or OR4 (N25286, N25285, N14888, N8355, N16351);
xor XOR2 (N25287, N25269, N3669);
xor XOR2 (N25288, N25281, N18126);
or OR4 (N25289, N25279, N6619, N8706, N8947);
xor XOR2 (N25290, N25282, N11525);
or OR2 (N25291, N25286, N19446);
and AND2 (N25292, N25272, N22714);
or OR3 (N25293, N25289, N3222, N3015);
xor XOR2 (N25294, N25290, N21538);
and AND2 (N25295, N25276, N251);
and AND4 (N25296, N25277, N15910, N13861, N8910);
nand NAND4 (N25297, N25287, N13884, N3377, N938);
not NOT1 (N25298, N25295);
not NOT1 (N25299, N25293);
buf BUF1 (N25300, N25297);
or OR4 (N25301, N25296, N12053, N3133, N2961);
nor NOR4 (N25302, N25291, N20901, N24066, N23033);
xor XOR2 (N25303, N25288, N15859);
nand NAND2 (N25304, N25283, N14727);
buf BUF1 (N25305, N25304);
or OR2 (N25306, N25292, N20101);
and AND3 (N25307, N25298, N17373, N10978);
nor NOR3 (N25308, N25303, N875, N23378);
xor XOR2 (N25309, N25307, N9617);
nand NAND4 (N25310, N25294, N25022, N20002, N24888);
nand NAND3 (N25311, N25301, N5264, N8659);
nand NAND2 (N25312, N25305, N9011);
nor NOR3 (N25313, N25300, N23072, N3976);
and AND4 (N25314, N25267, N3863, N13932, N1115);
not NOT1 (N25315, N25312);
nor NOR3 (N25316, N25315, N21667, N6076);
xor XOR2 (N25317, N25309, N7105);
nand NAND3 (N25318, N25308, N2851, N18168);
buf BUF1 (N25319, N25314);
xor XOR2 (N25320, N25310, N1859);
or OR3 (N25321, N25320, N11911, N16722);
nor NOR2 (N25322, N25302, N14192);
and AND3 (N25323, N25313, N788, N8927);
xor XOR2 (N25324, N25323, N4684);
buf BUF1 (N25325, N25322);
xor XOR2 (N25326, N25311, N17880);
nand NAND2 (N25327, N25318, N16204);
or OR2 (N25328, N25327, N21198);
and AND2 (N25329, N25328, N20470);
nor NOR4 (N25330, N25326, N20042, N25284, N1729);
buf BUF1 (N25331, N25316);
nand NAND2 (N25332, N25331, N2402);
nand NAND3 (N25333, N25321, N19674, N24638);
and AND3 (N25334, N25299, N12888, N748);
xor XOR2 (N25335, N25306, N1567);
nor NOR3 (N25336, N25317, N10745, N2469);
xor XOR2 (N25337, N25336, N21199);
nor NOR4 (N25338, N25337, N16935, N1970, N17134);
nor NOR4 (N25339, N25324, N21640, N12447, N9100);
nor NOR4 (N25340, N25332, N11189, N11324, N24031);
and AND4 (N25341, N25329, N9724, N14141, N18621);
buf BUF1 (N25342, N25333);
xor XOR2 (N25343, N25334, N15672);
xor XOR2 (N25344, N25338, N13251);
and AND3 (N25345, N25319, N21354, N6651);
not NOT1 (N25346, N25343);
not NOT1 (N25347, N25339);
nor NOR3 (N25348, N25346, N2317, N10635);
buf BUF1 (N25349, N25325);
not NOT1 (N25350, N25345);
or OR3 (N25351, N25347, N13733, N1162);
or OR4 (N25352, N25342, N21724, N10934, N12610);
or OR2 (N25353, N25351, N17908);
nor NOR3 (N25354, N25344, N9187, N10861);
nor NOR2 (N25355, N25340, N3835);
or OR3 (N25356, N25349, N2029, N1376);
not NOT1 (N25357, N25355);
and AND3 (N25358, N25356, N2538, N8914);
buf BUF1 (N25359, N25348);
xor XOR2 (N25360, N25352, N23459);
nor NOR2 (N25361, N25360, N23772);
nor NOR3 (N25362, N25361, N8236, N6061);
buf BUF1 (N25363, N25359);
not NOT1 (N25364, N25358);
nand NAND4 (N25365, N25354, N1124, N1623, N15512);
xor XOR2 (N25366, N25335, N18190);
and AND2 (N25367, N25362, N22098);
and AND4 (N25368, N25353, N24551, N3639, N5409);
or OR4 (N25369, N25341, N2845, N23776, N10581);
nand NAND4 (N25370, N25363, N2956, N23880, N1168);
or OR4 (N25371, N25370, N3329, N2841, N24348);
nand NAND2 (N25372, N25368, N10860);
or OR2 (N25373, N25367, N21255);
and AND2 (N25374, N25357, N8847);
and AND4 (N25375, N25373, N3182, N14474, N912);
not NOT1 (N25376, N25371);
buf BUF1 (N25377, N25375);
not NOT1 (N25378, N25376);
not NOT1 (N25379, N25330);
nand NAND4 (N25380, N25378, N19077, N19422, N18938);
nand NAND3 (N25381, N25379, N17320, N18777);
not NOT1 (N25382, N25377);
xor XOR2 (N25383, N25365, N15523);
buf BUF1 (N25384, N25372);
buf BUF1 (N25385, N25366);
or OR3 (N25386, N25364, N19023, N5679);
not NOT1 (N25387, N25381);
nor NOR2 (N25388, N25382, N1743);
or OR4 (N25389, N25380, N11785, N8838, N3849);
nor NOR4 (N25390, N25387, N18663, N23537, N5037);
nor NOR4 (N25391, N25389, N14732, N19281, N23455);
nand NAND2 (N25392, N25384, N5120);
and AND4 (N25393, N25390, N12235, N7736, N9447);
and AND2 (N25394, N25391, N9004);
buf BUF1 (N25395, N25394);
nor NOR3 (N25396, N25386, N14677, N11232);
or OR4 (N25397, N25369, N9371, N17202, N11055);
xor XOR2 (N25398, N25388, N24328);
nand NAND2 (N25399, N25395, N16430);
buf BUF1 (N25400, N25383);
not NOT1 (N25401, N25398);
not NOT1 (N25402, N25393);
or OR4 (N25403, N25397, N21642, N10094, N6691);
or OR2 (N25404, N25402, N16465);
and AND2 (N25405, N25392, N4259);
xor XOR2 (N25406, N25403, N67);
or OR3 (N25407, N25350, N1997, N8783);
xor XOR2 (N25408, N25396, N23293);
nand NAND4 (N25409, N25374, N4340, N2602, N4824);
not NOT1 (N25410, N25407);
nor NOR4 (N25411, N25404, N6501, N25121, N23771);
buf BUF1 (N25412, N25405);
nand NAND2 (N25413, N25401, N21842);
xor XOR2 (N25414, N25409, N11307);
or OR4 (N25415, N25406, N20262, N5485, N14864);
and AND2 (N25416, N25400, N18058);
xor XOR2 (N25417, N25399, N6017);
and AND4 (N25418, N25412, N14815, N2033, N10653);
not NOT1 (N25419, N25413);
or OR4 (N25420, N25385, N20128, N13062, N1974);
not NOT1 (N25421, N25419);
or OR2 (N25422, N25417, N5719);
and AND3 (N25423, N25411, N21028, N6979);
nor NOR3 (N25424, N25414, N20540, N19238);
not NOT1 (N25425, N25422);
nand NAND2 (N25426, N25425, N3329);
xor XOR2 (N25427, N25418, N4242);
not NOT1 (N25428, N25410);
buf BUF1 (N25429, N25420);
and AND4 (N25430, N25415, N5309, N24968, N147);
or OR3 (N25431, N25408, N15100, N4715);
nor NOR3 (N25432, N25428, N19169, N3492);
nand NAND4 (N25433, N25427, N7798, N19646, N22355);
and AND2 (N25434, N25421, N8024);
and AND3 (N25435, N25416, N1074, N21033);
xor XOR2 (N25436, N25429, N20582);
buf BUF1 (N25437, N25423);
not NOT1 (N25438, N25435);
nor NOR3 (N25439, N25434, N18763, N24501);
buf BUF1 (N25440, N25438);
nand NAND3 (N25441, N25430, N23788, N5631);
or OR2 (N25442, N25426, N18449);
and AND2 (N25443, N25436, N7955);
buf BUF1 (N25444, N25424);
nor NOR4 (N25445, N25441, N4783, N4372, N20118);
or OR3 (N25446, N25433, N8530, N1622);
nor NOR3 (N25447, N25445, N15883, N960);
xor XOR2 (N25448, N25446, N17019);
or OR3 (N25449, N25432, N24785, N18947);
and AND3 (N25450, N25448, N16202, N13133);
xor XOR2 (N25451, N25437, N19855);
nor NOR4 (N25452, N25451, N20952, N24129, N18517);
nor NOR2 (N25453, N25440, N11316);
buf BUF1 (N25454, N25449);
or OR3 (N25455, N25444, N23386, N14472);
buf BUF1 (N25456, N25439);
not NOT1 (N25457, N25455);
nor NOR2 (N25458, N25431, N19059);
or OR4 (N25459, N25450, N13050, N15247, N20962);
xor XOR2 (N25460, N25459, N8107);
buf BUF1 (N25461, N25460);
not NOT1 (N25462, N25458);
and AND3 (N25463, N25454, N10569, N12343);
or OR3 (N25464, N25462, N23611, N2274);
buf BUF1 (N25465, N25464);
xor XOR2 (N25466, N25461, N3235);
or OR2 (N25467, N25447, N6556);
and AND2 (N25468, N25467, N5566);
buf BUF1 (N25469, N25457);
or OR4 (N25470, N25468, N12296, N10654, N17508);
nand NAND2 (N25471, N25469, N14290);
and AND4 (N25472, N25463, N15311, N19215, N7342);
and AND2 (N25473, N25442, N11496);
nand NAND2 (N25474, N25471, N11772);
and AND4 (N25475, N25465, N25142, N14801, N512);
not NOT1 (N25476, N25453);
or OR4 (N25477, N25443, N13843, N17138, N6043);
and AND3 (N25478, N25473, N24758, N13036);
nor NOR4 (N25479, N25456, N14725, N4291, N23262);
nand NAND3 (N25480, N25452, N8064, N20356);
buf BUF1 (N25481, N25466);
nor NOR4 (N25482, N25470, N20120, N13810, N9859);
or OR3 (N25483, N25478, N11674, N23792);
nor NOR3 (N25484, N25482, N14946, N21966);
buf BUF1 (N25485, N25484);
buf BUF1 (N25486, N25474);
nor NOR2 (N25487, N25483, N1031);
buf BUF1 (N25488, N25487);
xor XOR2 (N25489, N25479, N18818);
or OR4 (N25490, N25476, N942, N16981, N18102);
and AND4 (N25491, N25477, N13825, N23227, N12543);
nor NOR2 (N25492, N25472, N7259);
and AND3 (N25493, N25475, N19703, N24057);
nand NAND2 (N25494, N25491, N9868);
nor NOR2 (N25495, N25486, N20599);
and AND2 (N25496, N25489, N9875);
xor XOR2 (N25497, N25493, N20107);
nor NOR3 (N25498, N25481, N22612, N7384);
xor XOR2 (N25499, N25496, N3004);
nand NAND3 (N25500, N25495, N24357, N322);
nor NOR2 (N25501, N25488, N15878);
buf BUF1 (N25502, N25480);
nor NOR4 (N25503, N25498, N24348, N21501, N18712);
buf BUF1 (N25504, N25499);
xor XOR2 (N25505, N25501, N12230);
xor XOR2 (N25506, N25502, N2085);
and AND3 (N25507, N25503, N11003, N11796);
buf BUF1 (N25508, N25494);
nor NOR4 (N25509, N25506, N16527, N11015, N13633);
buf BUF1 (N25510, N25492);
and AND2 (N25511, N25509, N24582);
nand NAND4 (N25512, N25507, N16252, N25225, N4615);
nand NAND3 (N25513, N25511, N16667, N24400);
nor NOR3 (N25514, N25505, N20301, N5678);
or OR3 (N25515, N25514, N11073, N23736);
nand NAND4 (N25516, N25508, N24938, N19460, N5124);
or OR2 (N25517, N25515, N22712);
or OR4 (N25518, N25510, N21614, N22059, N19147);
xor XOR2 (N25519, N25516, N679);
or OR4 (N25520, N25512, N25229, N19992, N5088);
buf BUF1 (N25521, N25518);
or OR4 (N25522, N25520, N13124, N1450, N15153);
buf BUF1 (N25523, N25504);
or OR4 (N25524, N25517, N5767, N11372, N5570);
nor NOR4 (N25525, N25522, N1277, N10840, N1065);
not NOT1 (N25526, N25500);
nor NOR2 (N25527, N25523, N21909);
xor XOR2 (N25528, N25490, N20922);
or OR4 (N25529, N25528, N4926, N768, N2733);
or OR4 (N25530, N25513, N11287, N4303, N5190);
buf BUF1 (N25531, N25497);
not NOT1 (N25532, N25524);
or OR3 (N25533, N25531, N18182, N10812);
or OR3 (N25534, N25526, N14656, N25286);
or OR3 (N25535, N25527, N12331, N1356);
nand NAND4 (N25536, N25519, N17795, N7698, N23055);
nor NOR2 (N25537, N25530, N5326);
and AND3 (N25538, N25536, N20789, N23185);
nor NOR4 (N25539, N25529, N9691, N22091, N12078);
buf BUF1 (N25540, N25525);
buf BUF1 (N25541, N25535);
xor XOR2 (N25542, N25538, N12311);
buf BUF1 (N25543, N25541);
not NOT1 (N25544, N25542);
or OR4 (N25545, N25537, N1910, N2583, N7306);
nand NAND3 (N25546, N25543, N2911, N14288);
nor NOR3 (N25547, N25539, N12792, N5226);
or OR4 (N25548, N25540, N13134, N25000, N20849);
nor NOR2 (N25549, N25485, N20530);
nor NOR3 (N25550, N25532, N10686, N3734);
and AND2 (N25551, N25521, N1504);
or OR2 (N25552, N25546, N9696);
nor NOR3 (N25553, N25534, N16941, N21610);
buf BUF1 (N25554, N25552);
or OR3 (N25555, N25554, N10814, N15876);
nor NOR4 (N25556, N25548, N8910, N9637, N2142);
buf BUF1 (N25557, N25545);
nor NOR4 (N25558, N25551, N24085, N7759, N8133);
and AND4 (N25559, N25547, N2087, N143, N17975);
not NOT1 (N25560, N25553);
buf BUF1 (N25561, N25549);
nor NOR4 (N25562, N25544, N1811, N6578, N5963);
buf BUF1 (N25563, N25558);
and AND2 (N25564, N25563, N19877);
nand NAND2 (N25565, N25556, N15619);
buf BUF1 (N25566, N25561);
nand NAND3 (N25567, N25555, N11579, N4445);
and AND3 (N25568, N25550, N12901, N22472);
and AND3 (N25569, N25568, N17694, N21963);
xor XOR2 (N25570, N25562, N12022);
buf BUF1 (N25571, N25570);
and AND4 (N25572, N25566, N11993, N22538, N11959);
or OR2 (N25573, N25571, N23942);
nor NOR2 (N25574, N25565, N9361);
nor NOR3 (N25575, N25557, N18221, N16892);
nand NAND2 (N25576, N25575, N23825);
or OR3 (N25577, N25560, N22007, N10962);
and AND3 (N25578, N25564, N15369, N4099);
nand NAND2 (N25579, N25567, N16484);
and AND2 (N25580, N25577, N899);
nor NOR2 (N25581, N25572, N10327);
buf BUF1 (N25582, N25578);
nand NAND2 (N25583, N25559, N24911);
nand NAND3 (N25584, N25569, N16606, N14517);
not NOT1 (N25585, N25584);
nand NAND2 (N25586, N25574, N24614);
nor NOR4 (N25587, N25579, N11942, N18602, N13626);
xor XOR2 (N25588, N25573, N6614);
nor NOR3 (N25589, N25576, N22077, N8084);
not NOT1 (N25590, N25585);
not NOT1 (N25591, N25587);
xor XOR2 (N25592, N25589, N8417);
xor XOR2 (N25593, N25592, N16688);
and AND2 (N25594, N25590, N25113);
nand NAND2 (N25595, N25593, N22239);
and AND3 (N25596, N25595, N21419, N21064);
xor XOR2 (N25597, N25591, N14930);
not NOT1 (N25598, N25596);
or OR3 (N25599, N25588, N10910, N7171);
and AND4 (N25600, N25533, N2349, N7911, N13094);
or OR2 (N25601, N25594, N24774);
buf BUF1 (N25602, N25581);
not NOT1 (N25603, N25582);
xor XOR2 (N25604, N25598, N11150);
buf BUF1 (N25605, N25597);
xor XOR2 (N25606, N25603, N12574);
nand NAND2 (N25607, N25602, N783);
buf BUF1 (N25608, N25583);
nor NOR3 (N25609, N25606, N16255, N16706);
not NOT1 (N25610, N25604);
buf BUF1 (N25611, N25599);
buf BUF1 (N25612, N25607);
and AND4 (N25613, N25601, N2410, N10164, N23298);
nand NAND2 (N25614, N25612, N12859);
not NOT1 (N25615, N25600);
buf BUF1 (N25616, N25580);
and AND2 (N25617, N25613, N4787);
endmodule