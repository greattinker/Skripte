// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N1618,N1606,N1615,N1599,N1603,N1619,N1611,N1608,N1620,N1621;

buf BUF1 (N22, N11);
buf BUF1 (N23, N20);
xor XOR2 (N24, N10, N9);
xor XOR2 (N25, N7, N20);
or OR4 (N26, N21, N15, N4, N19);
or OR3 (N27, N2, N9, N23);
nor NOR3 (N28, N3, N17, N23);
xor XOR2 (N29, N26, N7);
or OR2 (N30, N21, N10);
and AND3 (N31, N6, N27, N4);
nand NAND4 (N32, N11, N9, N15, N27);
and AND2 (N33, N15, N2);
nor NOR2 (N34, N18, N3);
xor XOR2 (N35, N32, N2);
buf BUF1 (N36, N29);
xor XOR2 (N37, N28, N35);
and AND4 (N38, N36, N31, N15, N30);
xor XOR2 (N39, N25, N9);
nor NOR4 (N40, N11, N25, N39, N37);
buf BUF1 (N41, N14);
or OR4 (N42, N7, N5, N11, N34);
xor XOR2 (N43, N9, N40);
and AND3 (N44, N34, N42, N9);
nand NAND3 (N45, N14, N25, N36);
nand NAND4 (N46, N15, N34, N17, N23);
buf BUF1 (N47, N38);
not NOT1 (N48, N17);
xor XOR2 (N49, N33, N4);
xor XOR2 (N50, N41, N15);
not NOT1 (N51, N43);
nor NOR4 (N52, N48, N27, N17, N42);
nor NOR2 (N53, N52, N23);
nor NOR3 (N54, N45, N27, N35);
not NOT1 (N55, N22);
and AND2 (N56, N53, N36);
and AND2 (N57, N47, N27);
nor NOR4 (N58, N57, N48, N25, N11);
or OR4 (N59, N24, N38, N45, N51);
buf BUF1 (N60, N54);
buf BUF1 (N61, N42);
xor XOR2 (N62, N60, N34);
buf BUF1 (N63, N46);
and AND2 (N64, N49, N32);
buf BUF1 (N65, N44);
nand NAND2 (N66, N62, N23);
nand NAND2 (N67, N56, N9);
buf BUF1 (N68, N66);
or OR4 (N69, N50, N62, N21, N38);
or OR2 (N70, N69, N55);
or OR4 (N71, N56, N56, N3, N54);
not NOT1 (N72, N71);
buf BUF1 (N73, N65);
nand NAND2 (N74, N70, N28);
not NOT1 (N75, N61);
or OR2 (N76, N68, N44);
xor XOR2 (N77, N76, N10);
or OR3 (N78, N59, N20, N60);
nand NAND3 (N79, N78, N77, N36);
nand NAND4 (N80, N31, N72, N22, N30);
and AND3 (N81, N5, N79, N14);
nor NOR3 (N82, N7, N10, N66);
and AND2 (N83, N81, N60);
buf BUF1 (N84, N64);
not NOT1 (N85, N83);
and AND4 (N86, N85, N79, N41, N43);
and AND3 (N87, N67, N10, N63);
buf BUF1 (N88, N84);
xor XOR2 (N89, N42, N42);
xor XOR2 (N90, N74, N16);
xor XOR2 (N91, N58, N17);
xor XOR2 (N92, N80, N29);
nand NAND3 (N93, N92, N60, N28);
and AND3 (N94, N75, N54, N68);
not NOT1 (N95, N91);
and AND2 (N96, N88, N18);
buf BUF1 (N97, N86);
nand NAND3 (N98, N93, N3, N84);
buf BUF1 (N99, N90);
nand NAND3 (N100, N89, N98, N87);
nand NAND4 (N101, N89, N92, N13, N37);
or OR2 (N102, N59, N24);
not NOT1 (N103, N101);
or OR4 (N104, N103, N77, N85, N58);
or OR4 (N105, N95, N38, N83, N67);
xor XOR2 (N106, N82, N23);
buf BUF1 (N107, N73);
nand NAND2 (N108, N100, N58);
nor NOR2 (N109, N108, N6);
nor NOR4 (N110, N99, N6, N40, N50);
not NOT1 (N111, N94);
xor XOR2 (N112, N109, N50);
and AND4 (N113, N102, N100, N20, N46);
xor XOR2 (N114, N110, N69);
nor NOR3 (N115, N104, N1, N49);
xor XOR2 (N116, N96, N67);
or OR4 (N117, N113, N32, N96, N46);
not NOT1 (N118, N116);
xor XOR2 (N119, N118, N12);
not NOT1 (N120, N97);
xor XOR2 (N121, N105, N103);
or OR4 (N122, N120, N46, N15, N117);
not NOT1 (N123, N64);
and AND3 (N124, N106, N67, N7);
or OR2 (N125, N121, N29);
or OR4 (N126, N119, N1, N38, N88);
nand NAND2 (N127, N125, N79);
buf BUF1 (N128, N112);
xor XOR2 (N129, N124, N71);
not NOT1 (N130, N122);
and AND3 (N131, N130, N6, N57);
not NOT1 (N132, N111);
not NOT1 (N133, N129);
nor NOR4 (N134, N128, N101, N54, N100);
and AND2 (N135, N107, N85);
nand NAND3 (N136, N133, N112, N29);
buf BUF1 (N137, N114);
nand NAND4 (N138, N123, N37, N130, N122);
nor NOR2 (N139, N135, N117);
nand NAND3 (N140, N126, N60, N98);
or OR3 (N141, N140, N94, N98);
or OR2 (N142, N137, N126);
xor XOR2 (N143, N115, N139);
not NOT1 (N144, N47);
xor XOR2 (N145, N138, N56);
nand NAND2 (N146, N144, N129);
buf BUF1 (N147, N132);
and AND2 (N148, N134, N67);
xor XOR2 (N149, N145, N101);
buf BUF1 (N150, N136);
nor NOR4 (N151, N131, N145, N144, N34);
buf BUF1 (N152, N147);
nand NAND3 (N153, N146, N53, N70);
or OR3 (N154, N150, N86, N27);
and AND3 (N155, N142, N113, N8);
nor NOR2 (N156, N127, N46);
and AND4 (N157, N156, N53, N143, N36);
nor NOR4 (N158, N130, N108, N60, N2);
or OR3 (N159, N148, N143, N74);
nand NAND4 (N160, N149, N60, N41, N114);
not NOT1 (N161, N154);
and AND3 (N162, N158, N39, N63);
not NOT1 (N163, N155);
buf BUF1 (N164, N152);
nor NOR2 (N165, N160, N20);
and AND3 (N166, N157, N115, N136);
and AND4 (N167, N166, N88, N138, N132);
and AND2 (N168, N153, N161);
or OR3 (N169, N43, N114, N130);
nor NOR4 (N170, N151, N52, N48, N155);
not NOT1 (N171, N164);
nor NOR4 (N172, N169, N144, N14, N108);
nand NAND3 (N173, N159, N50, N28);
and AND4 (N174, N162, N162, N122, N20);
not NOT1 (N175, N173);
and AND2 (N176, N171, N115);
and AND2 (N177, N170, N141);
buf BUF1 (N178, N47);
nor NOR3 (N179, N174, N150, N92);
nand NAND4 (N180, N175, N59, N25, N140);
nor NOR4 (N181, N163, N126, N113, N103);
nand NAND3 (N182, N178, N31, N151);
buf BUF1 (N183, N168);
or OR4 (N184, N177, N15, N25, N154);
nor NOR3 (N185, N180, N154, N86);
not NOT1 (N186, N176);
nor NOR2 (N187, N172, N92);
not NOT1 (N188, N182);
nor NOR4 (N189, N179, N64, N104, N169);
or OR3 (N190, N183, N157, N4);
or OR4 (N191, N184, N52, N40, N85);
not NOT1 (N192, N188);
not NOT1 (N193, N167);
nor NOR3 (N194, N189, N80, N180);
and AND2 (N195, N193, N75);
or OR4 (N196, N181, N152, N163, N112);
buf BUF1 (N197, N196);
or OR2 (N198, N195, N109);
not NOT1 (N199, N194);
nor NOR2 (N200, N165, N58);
nand NAND4 (N201, N198, N64, N23, N44);
nand NAND2 (N202, N190, N19);
xor XOR2 (N203, N186, N142);
or OR2 (N204, N200, N138);
xor XOR2 (N205, N187, N85);
not NOT1 (N206, N191);
not NOT1 (N207, N205);
nor NOR4 (N208, N197, N165, N166, N81);
not NOT1 (N209, N192);
nor NOR2 (N210, N185, N76);
nor NOR3 (N211, N199, N116, N149);
not NOT1 (N212, N207);
not NOT1 (N213, N201);
or OR3 (N214, N208, N150, N44);
xor XOR2 (N215, N203, N212);
xor XOR2 (N216, N5, N97);
buf BUF1 (N217, N206);
xor XOR2 (N218, N213, N12);
buf BUF1 (N219, N211);
or OR2 (N220, N214, N189);
nor NOR2 (N221, N215, N214);
buf BUF1 (N222, N221);
or OR2 (N223, N210, N123);
xor XOR2 (N224, N218, N112);
and AND3 (N225, N223, N9, N66);
and AND3 (N226, N209, N208, N34);
nor NOR2 (N227, N224, N119);
nor NOR2 (N228, N220, N138);
and AND2 (N229, N202, N165);
and AND2 (N230, N219, N130);
nor NOR2 (N231, N216, N70);
not NOT1 (N232, N231);
nor NOR3 (N233, N229, N169, N76);
buf BUF1 (N234, N232);
xor XOR2 (N235, N217, N183);
or OR3 (N236, N227, N75, N123);
nor NOR2 (N237, N226, N150);
and AND2 (N238, N236, N115);
nor NOR2 (N239, N222, N110);
or OR3 (N240, N239, N164, N13);
nor NOR4 (N241, N230, N178, N35, N179);
and AND2 (N242, N228, N232);
xor XOR2 (N243, N242, N99);
not NOT1 (N244, N225);
and AND2 (N245, N244, N17);
xor XOR2 (N246, N234, N231);
xor XOR2 (N247, N204, N87);
or OR4 (N248, N240, N194, N112, N166);
not NOT1 (N249, N241);
or OR4 (N250, N245, N243, N164, N106);
nand NAND3 (N251, N87, N213, N166);
buf BUF1 (N252, N250);
nor NOR2 (N253, N238, N203);
or OR2 (N254, N235, N161);
nand NAND4 (N255, N249, N59, N172, N179);
nand NAND4 (N256, N248, N5, N14, N240);
buf BUF1 (N257, N253);
buf BUF1 (N258, N252);
and AND2 (N259, N257, N12);
nor NOR3 (N260, N237, N104, N253);
not NOT1 (N261, N256);
or OR2 (N262, N260, N154);
nor NOR3 (N263, N254, N113, N144);
xor XOR2 (N264, N246, N233);
nand NAND4 (N265, N156, N257, N129, N227);
or OR2 (N266, N265, N204);
nor NOR4 (N267, N247, N49, N231, N68);
xor XOR2 (N268, N251, N118);
xor XOR2 (N269, N264, N113);
not NOT1 (N270, N268);
nand NAND2 (N271, N267, N19);
nor NOR2 (N272, N271, N43);
or OR3 (N273, N255, N250, N5);
xor XOR2 (N274, N272, N98);
nand NAND2 (N275, N273, N258);
nor NOR2 (N276, N36, N96);
or OR2 (N277, N259, N51);
not NOT1 (N278, N269);
nor NOR2 (N279, N276, N270);
buf BUF1 (N280, N242);
not NOT1 (N281, N266);
nor NOR2 (N282, N281, N64);
xor XOR2 (N283, N274, N12);
or OR2 (N284, N263, N114);
or OR2 (N285, N283, N101);
buf BUF1 (N286, N285);
buf BUF1 (N287, N275);
and AND3 (N288, N261, N239, N144);
buf BUF1 (N289, N279);
or OR2 (N290, N288, N37);
not NOT1 (N291, N287);
buf BUF1 (N292, N286);
not NOT1 (N293, N277);
and AND4 (N294, N280, N139, N94, N33);
and AND2 (N295, N289, N178);
not NOT1 (N296, N295);
xor XOR2 (N297, N291, N215);
and AND2 (N298, N282, N236);
buf BUF1 (N299, N284);
not NOT1 (N300, N278);
and AND4 (N301, N294, N160, N171, N188);
nand NAND4 (N302, N290, N163, N162, N64);
and AND2 (N303, N298, N61);
and AND2 (N304, N262, N46);
and AND3 (N305, N292, N101, N174);
buf BUF1 (N306, N300);
and AND4 (N307, N293, N218, N253, N215);
buf BUF1 (N308, N307);
not NOT1 (N309, N304);
nor NOR3 (N310, N299, N89, N57);
nand NAND2 (N311, N302, N301);
and AND4 (N312, N266, N210, N36, N117);
xor XOR2 (N313, N297, N249);
not NOT1 (N314, N305);
buf BUF1 (N315, N313);
and AND3 (N316, N296, N231, N274);
xor XOR2 (N317, N303, N50);
nor NOR3 (N318, N310, N306, N150);
not NOT1 (N319, N232);
xor XOR2 (N320, N315, N27);
nand NAND4 (N321, N319, N120, N278, N175);
nand NAND2 (N322, N311, N196);
nand NAND4 (N323, N308, N95, N142, N303);
nor NOR2 (N324, N323, N11);
and AND4 (N325, N321, N289, N266, N200);
not NOT1 (N326, N320);
or OR3 (N327, N309, N109, N159);
nand NAND2 (N328, N326, N28);
buf BUF1 (N329, N312);
buf BUF1 (N330, N324);
and AND4 (N331, N325, N79, N129, N104);
or OR2 (N332, N327, N189);
nand NAND4 (N333, N318, N260, N225, N191);
nor NOR2 (N334, N329, N75);
not NOT1 (N335, N314);
and AND4 (N336, N332, N269, N294, N42);
buf BUF1 (N337, N317);
nor NOR4 (N338, N328, N242, N331, N122);
and AND4 (N339, N321, N139, N121, N106);
not NOT1 (N340, N322);
or OR3 (N341, N339, N32, N32);
or OR3 (N342, N335, N338, N253);
and AND4 (N343, N89, N165, N192, N268);
not NOT1 (N344, N342);
nand NAND2 (N345, N343, N12);
nand NAND2 (N346, N336, N231);
nand NAND3 (N347, N341, N88, N226);
nand NAND4 (N348, N334, N273, N216, N2);
or OR3 (N349, N330, N148, N343);
buf BUF1 (N350, N347);
xor XOR2 (N351, N346, N98);
nand NAND3 (N352, N333, N89, N19);
not NOT1 (N353, N340);
nor NOR4 (N354, N351, N324, N351, N247);
nand NAND2 (N355, N345, N236);
not NOT1 (N356, N352);
not NOT1 (N357, N350);
xor XOR2 (N358, N344, N154);
nor NOR2 (N359, N358, N22);
not NOT1 (N360, N357);
not NOT1 (N361, N316);
buf BUF1 (N362, N361);
nand NAND2 (N363, N354, N329);
nand NAND4 (N364, N349, N114, N231, N91);
buf BUF1 (N365, N363);
xor XOR2 (N366, N355, N97);
not NOT1 (N367, N356);
xor XOR2 (N368, N360, N138);
buf BUF1 (N369, N366);
nor NOR2 (N370, N365, N320);
and AND2 (N371, N368, N325);
not NOT1 (N372, N337);
nor NOR3 (N373, N362, N88, N351);
or OR4 (N374, N353, N76, N25, N109);
buf BUF1 (N375, N359);
nand NAND3 (N376, N348, N132, N269);
buf BUF1 (N377, N376);
not NOT1 (N378, N364);
and AND3 (N379, N378, N188, N239);
and AND2 (N380, N370, N237);
buf BUF1 (N381, N379);
or OR3 (N382, N374, N165, N373);
nor NOR4 (N383, N218, N221, N139, N332);
not NOT1 (N384, N380);
or OR2 (N385, N375, N197);
and AND2 (N386, N371, N193);
or OR3 (N387, N384, N213, N332);
nor NOR3 (N388, N381, N113, N101);
not NOT1 (N389, N369);
not NOT1 (N390, N367);
and AND2 (N391, N383, N73);
and AND4 (N392, N386, N313, N91, N324);
xor XOR2 (N393, N392, N334);
buf BUF1 (N394, N391);
nor NOR4 (N395, N393, N108, N106, N285);
xor XOR2 (N396, N382, N362);
xor XOR2 (N397, N389, N176);
buf BUF1 (N398, N385);
not NOT1 (N399, N390);
or OR4 (N400, N397, N136, N303, N215);
not NOT1 (N401, N396);
buf BUF1 (N402, N395);
xor XOR2 (N403, N377, N111);
and AND3 (N404, N403, N347, N197);
nand NAND3 (N405, N394, N98, N120);
or OR3 (N406, N404, N172, N17);
and AND2 (N407, N388, N365);
nor NOR2 (N408, N399, N59);
and AND4 (N409, N372, N226, N146, N78);
nor NOR2 (N410, N405, N241);
buf BUF1 (N411, N401);
nor NOR3 (N412, N406, N150, N298);
and AND4 (N413, N387, N113, N236, N83);
nor NOR3 (N414, N412, N135, N244);
buf BUF1 (N415, N413);
nor NOR3 (N416, N398, N397, N40);
not NOT1 (N417, N400);
or OR3 (N418, N415, N67, N399);
not NOT1 (N419, N418);
and AND3 (N420, N407, N390, N19);
xor XOR2 (N421, N411, N164);
not NOT1 (N422, N414);
or OR4 (N423, N417, N26, N252, N289);
not NOT1 (N424, N423);
xor XOR2 (N425, N402, N159);
and AND3 (N426, N422, N89, N91);
and AND2 (N427, N421, N3);
and AND2 (N428, N416, N44);
not NOT1 (N429, N420);
not NOT1 (N430, N425);
not NOT1 (N431, N419);
and AND4 (N432, N410, N108, N366, N265);
xor XOR2 (N433, N408, N85);
nand NAND3 (N434, N409, N227, N230);
xor XOR2 (N435, N432, N76);
buf BUF1 (N436, N434);
nand NAND4 (N437, N424, N94, N109, N110);
nor NOR4 (N438, N426, N173, N128, N336);
xor XOR2 (N439, N430, N218);
or OR4 (N440, N429, N371, N422, N223);
nand NAND3 (N441, N433, N381, N30);
or OR4 (N442, N440, N406, N200, N152);
xor XOR2 (N443, N441, N143);
nand NAND2 (N444, N438, N229);
buf BUF1 (N445, N437);
and AND2 (N446, N439, N129);
nor NOR4 (N447, N446, N442, N178, N310);
not NOT1 (N448, N125);
not NOT1 (N449, N436);
and AND4 (N450, N443, N132, N74, N422);
nor NOR3 (N451, N435, N147, N183);
not NOT1 (N452, N447);
xor XOR2 (N453, N448, N99);
and AND3 (N454, N453, N440, N300);
buf BUF1 (N455, N449);
xor XOR2 (N456, N431, N19);
or OR4 (N457, N452, N209, N250, N139);
or OR2 (N458, N457, N101);
nor NOR3 (N459, N451, N178, N289);
or OR4 (N460, N454, N101, N207, N38);
xor XOR2 (N461, N456, N27);
xor XOR2 (N462, N427, N82);
nand NAND3 (N463, N462, N227, N228);
nor NOR2 (N464, N460, N146);
buf BUF1 (N465, N464);
xor XOR2 (N466, N465, N87);
nor NOR3 (N467, N458, N164, N12);
or OR3 (N468, N428, N48, N429);
not NOT1 (N469, N444);
not NOT1 (N470, N461);
and AND2 (N471, N467, N99);
and AND4 (N472, N463, N338, N77, N297);
and AND3 (N473, N455, N153, N69);
nand NAND4 (N474, N470, N121, N194, N392);
nor NOR4 (N475, N459, N409, N417, N83);
not NOT1 (N476, N450);
xor XOR2 (N477, N469, N265);
or OR2 (N478, N468, N212);
xor XOR2 (N479, N472, N375);
nand NAND2 (N480, N478, N277);
nand NAND3 (N481, N471, N289, N243);
nor NOR2 (N482, N480, N61);
or OR3 (N483, N473, N146, N84);
or OR3 (N484, N479, N236, N452);
xor XOR2 (N485, N475, N386);
not NOT1 (N486, N477);
buf BUF1 (N487, N486);
and AND3 (N488, N466, N112, N410);
nor NOR4 (N489, N488, N173, N344, N219);
buf BUF1 (N490, N485);
not NOT1 (N491, N481);
xor XOR2 (N492, N490, N149);
xor XOR2 (N493, N492, N309);
nor NOR3 (N494, N482, N91, N48);
nor NOR3 (N495, N474, N421, N174);
nor NOR3 (N496, N484, N254, N381);
and AND4 (N497, N493, N74, N389, N151);
not NOT1 (N498, N491);
and AND2 (N499, N494, N72);
or OR2 (N500, N497, N51);
nor NOR2 (N501, N499, N115);
buf BUF1 (N502, N495);
nor NOR4 (N503, N501, N167, N4, N200);
and AND4 (N504, N503, N205, N359, N273);
or OR3 (N505, N445, N121, N112);
nor NOR3 (N506, N487, N375, N50);
nor NOR4 (N507, N483, N88, N441, N88);
xor XOR2 (N508, N496, N34);
xor XOR2 (N509, N504, N253);
or OR2 (N510, N509, N233);
buf BUF1 (N511, N502);
xor XOR2 (N512, N506, N60);
or OR4 (N513, N500, N116, N9, N248);
nor NOR2 (N514, N508, N310);
or OR3 (N515, N511, N293, N8);
not NOT1 (N516, N515);
nand NAND3 (N517, N498, N410, N341);
or OR2 (N518, N476, N469);
and AND3 (N519, N505, N318, N238);
nor NOR2 (N520, N507, N1);
and AND2 (N521, N514, N210);
buf BUF1 (N522, N519);
buf BUF1 (N523, N510);
not NOT1 (N524, N516);
nand NAND4 (N525, N524, N470, N87, N78);
and AND4 (N526, N517, N115, N413, N505);
nor NOR4 (N527, N522, N425, N249, N25);
or OR4 (N528, N526, N149, N390, N394);
nor NOR3 (N529, N512, N414, N109);
xor XOR2 (N530, N520, N511);
and AND3 (N531, N530, N481, N521);
nand NAND2 (N532, N465, N258);
buf BUF1 (N533, N513);
buf BUF1 (N534, N518);
nor NOR2 (N535, N531, N287);
buf BUF1 (N536, N525);
and AND4 (N537, N533, N21, N244, N469);
xor XOR2 (N538, N536, N154);
nand NAND2 (N539, N527, N354);
or OR2 (N540, N534, N160);
or OR2 (N541, N540, N363);
nand NAND4 (N542, N535, N95, N80, N497);
nor NOR3 (N543, N532, N431, N319);
not NOT1 (N544, N528);
nand NAND2 (N545, N541, N141);
xor XOR2 (N546, N544, N316);
xor XOR2 (N547, N523, N489);
nor NOR4 (N548, N448, N19, N126, N220);
nor NOR2 (N549, N539, N135);
and AND4 (N550, N538, N85, N244, N3);
and AND4 (N551, N537, N245, N438, N212);
or OR3 (N552, N550, N94, N89);
not NOT1 (N553, N551);
nand NAND3 (N554, N546, N223, N374);
nor NOR4 (N555, N545, N474, N169, N554);
buf BUF1 (N556, N297);
nor NOR3 (N557, N543, N205, N257);
nor NOR3 (N558, N552, N495, N341);
and AND4 (N559, N549, N91, N531, N459);
xor XOR2 (N560, N556, N297);
and AND3 (N561, N529, N299, N435);
or OR3 (N562, N547, N52, N85);
nand NAND3 (N563, N548, N92, N509);
xor XOR2 (N564, N558, N525);
nand NAND2 (N565, N542, N297);
xor XOR2 (N566, N562, N261);
and AND4 (N567, N561, N183, N358, N343);
not NOT1 (N568, N557);
and AND3 (N569, N553, N259, N368);
and AND4 (N570, N559, N108, N3, N86);
nor NOR3 (N571, N560, N339, N31);
xor XOR2 (N572, N563, N250);
not NOT1 (N573, N568);
nand NAND3 (N574, N571, N463, N341);
xor XOR2 (N575, N567, N549);
xor XOR2 (N576, N572, N171);
or OR2 (N577, N566, N36);
nor NOR2 (N578, N565, N363);
buf BUF1 (N579, N569);
xor XOR2 (N580, N578, N523);
nor NOR3 (N581, N576, N547, N193);
and AND4 (N582, N581, N407, N384, N166);
nor NOR2 (N583, N564, N514);
buf BUF1 (N584, N580);
buf BUF1 (N585, N577);
xor XOR2 (N586, N585, N89);
buf BUF1 (N587, N582);
xor XOR2 (N588, N574, N484);
nand NAND4 (N589, N587, N540, N472, N300);
xor XOR2 (N590, N588, N139);
xor XOR2 (N591, N579, N204);
xor XOR2 (N592, N575, N559);
xor XOR2 (N593, N589, N262);
nand NAND3 (N594, N593, N272, N466);
not NOT1 (N595, N590);
or OR3 (N596, N584, N249, N120);
or OR2 (N597, N583, N218);
nor NOR4 (N598, N597, N546, N306, N450);
nand NAND2 (N599, N598, N566);
not NOT1 (N600, N591);
not NOT1 (N601, N570);
buf BUF1 (N602, N586);
nand NAND2 (N603, N555, N295);
not NOT1 (N604, N595);
nor NOR2 (N605, N596, N226);
nor NOR2 (N606, N602, N245);
xor XOR2 (N607, N599, N604);
xor XOR2 (N608, N181, N528);
buf BUF1 (N609, N601);
xor XOR2 (N610, N606, N406);
or OR4 (N611, N608, N538, N24, N570);
or OR3 (N612, N605, N165, N570);
nor NOR2 (N613, N609, N97);
nor NOR2 (N614, N573, N312);
nand NAND3 (N615, N610, N425, N512);
xor XOR2 (N616, N611, N568);
nand NAND3 (N617, N614, N3, N387);
nand NAND2 (N618, N617, N27);
or OR4 (N619, N616, N71, N430, N50);
nand NAND2 (N620, N612, N82);
or OR3 (N621, N607, N409, N447);
nor NOR2 (N622, N594, N144);
nor NOR2 (N623, N619, N335);
not NOT1 (N624, N600);
nand NAND4 (N625, N613, N355, N623, N606);
nor NOR4 (N626, N163, N449, N352, N220);
and AND4 (N627, N622, N346, N221, N581);
buf BUF1 (N628, N615);
and AND4 (N629, N620, N131, N255, N368);
xor XOR2 (N630, N603, N581);
not NOT1 (N631, N625);
not NOT1 (N632, N621);
nor NOR2 (N633, N631, N397);
nor NOR4 (N634, N624, N480, N454, N234);
nor NOR4 (N635, N627, N326, N398, N173);
nand NAND3 (N636, N629, N107, N600);
nor NOR4 (N637, N618, N271, N275, N305);
and AND2 (N638, N592, N41);
buf BUF1 (N639, N628);
nor NOR3 (N640, N632, N169, N30);
nand NAND4 (N641, N634, N580, N90, N390);
buf BUF1 (N642, N638);
and AND4 (N643, N642, N26, N366, N35);
buf BUF1 (N644, N633);
not NOT1 (N645, N641);
not NOT1 (N646, N626);
and AND2 (N647, N639, N24);
nand NAND3 (N648, N630, N415, N199);
xor XOR2 (N649, N644, N311);
buf BUF1 (N650, N643);
buf BUF1 (N651, N646);
and AND2 (N652, N648, N363);
buf BUF1 (N653, N645);
not NOT1 (N654, N652);
xor XOR2 (N655, N635, N436);
not NOT1 (N656, N653);
buf BUF1 (N657, N649);
buf BUF1 (N658, N651);
nand NAND3 (N659, N650, N264, N342);
xor XOR2 (N660, N658, N83);
nand NAND3 (N661, N659, N407, N425);
and AND2 (N662, N640, N506);
xor XOR2 (N663, N647, N652);
or OR2 (N664, N662, N78);
not NOT1 (N665, N663);
xor XOR2 (N666, N660, N325);
xor XOR2 (N667, N661, N506);
and AND2 (N668, N667, N205);
not NOT1 (N669, N654);
buf BUF1 (N670, N636);
nand NAND4 (N671, N656, N276, N540, N26);
nor NOR3 (N672, N669, N112, N472);
and AND4 (N673, N672, N116, N66, N270);
buf BUF1 (N674, N673);
nand NAND4 (N675, N665, N53, N44, N232);
or OR3 (N676, N668, N292, N65);
nand NAND4 (N677, N670, N447, N30, N304);
nor NOR2 (N678, N671, N615);
nor NOR2 (N679, N655, N451);
and AND2 (N680, N679, N92);
nor NOR3 (N681, N674, N520, N264);
nor NOR3 (N682, N657, N435, N681);
xor XOR2 (N683, N303, N388);
xor XOR2 (N684, N637, N96);
and AND3 (N685, N664, N26, N562);
and AND3 (N686, N678, N344, N377);
nor NOR4 (N687, N684, N10, N205, N10);
buf BUF1 (N688, N686);
and AND4 (N689, N683, N395, N226, N642);
buf BUF1 (N690, N676);
or OR3 (N691, N687, N384, N279);
nor NOR2 (N692, N689, N38);
or OR4 (N693, N677, N557, N246, N678);
or OR2 (N694, N666, N6);
and AND3 (N695, N688, N161, N477);
xor XOR2 (N696, N692, N243);
not NOT1 (N697, N691);
xor XOR2 (N698, N682, N380);
buf BUF1 (N699, N698);
buf BUF1 (N700, N695);
buf BUF1 (N701, N693);
and AND3 (N702, N690, N512, N118);
or OR3 (N703, N699, N475, N86);
and AND3 (N704, N696, N679, N645);
xor XOR2 (N705, N680, N77);
xor XOR2 (N706, N694, N510);
or OR2 (N707, N701, N91);
nor NOR3 (N708, N703, N628, N474);
xor XOR2 (N709, N700, N209);
not NOT1 (N710, N705);
nand NAND3 (N711, N702, N43, N83);
buf BUF1 (N712, N707);
buf BUF1 (N713, N712);
nor NOR3 (N714, N685, N608, N711);
not NOT1 (N715, N368);
and AND3 (N716, N714, N196, N213);
buf BUF1 (N717, N697);
not NOT1 (N718, N717);
xor XOR2 (N719, N718, N138);
nor NOR2 (N720, N675, N157);
xor XOR2 (N721, N706, N565);
or OR2 (N722, N713, N327);
nor NOR4 (N723, N709, N34, N187, N611);
and AND4 (N724, N719, N651, N241, N537);
xor XOR2 (N725, N716, N651);
buf BUF1 (N726, N715);
buf BUF1 (N727, N723);
or OR4 (N728, N704, N222, N88, N227);
xor XOR2 (N729, N710, N182);
buf BUF1 (N730, N722);
buf BUF1 (N731, N725);
and AND3 (N732, N708, N327, N32);
not NOT1 (N733, N720);
nand NAND4 (N734, N732, N610, N720, N644);
xor XOR2 (N735, N731, N454);
not NOT1 (N736, N726);
xor XOR2 (N737, N724, N59);
xor XOR2 (N738, N734, N67);
nand NAND2 (N739, N721, N447);
xor XOR2 (N740, N733, N426);
not NOT1 (N741, N735);
nand NAND3 (N742, N739, N229, N238);
not NOT1 (N743, N736);
nand NAND2 (N744, N743, N156);
or OR4 (N745, N741, N42, N191, N347);
xor XOR2 (N746, N745, N506);
xor XOR2 (N747, N737, N102);
xor XOR2 (N748, N729, N681);
or OR3 (N749, N740, N302, N261);
nor NOR4 (N750, N746, N741, N362, N718);
buf BUF1 (N751, N742);
not NOT1 (N752, N751);
nor NOR3 (N753, N738, N104, N500);
nand NAND3 (N754, N747, N548, N410);
and AND4 (N755, N749, N485, N215, N102);
nor NOR4 (N756, N750, N434, N305, N280);
not NOT1 (N757, N727);
xor XOR2 (N758, N744, N237);
and AND2 (N759, N754, N264);
xor XOR2 (N760, N728, N204);
nand NAND4 (N761, N760, N387, N17, N339);
or OR3 (N762, N748, N234, N146);
xor XOR2 (N763, N759, N233);
buf BUF1 (N764, N757);
not NOT1 (N765, N762);
nand NAND4 (N766, N756, N615, N125, N299);
nor NOR4 (N767, N761, N139, N433, N762);
nand NAND4 (N768, N766, N388, N7, N483);
buf BUF1 (N769, N730);
not NOT1 (N770, N764);
nor NOR3 (N771, N765, N49, N391);
nand NAND4 (N772, N770, N743, N161, N484);
or OR2 (N773, N755, N417);
and AND3 (N774, N771, N140, N247);
nand NAND2 (N775, N772, N701);
xor XOR2 (N776, N753, N380);
and AND4 (N777, N773, N251, N142, N190);
xor XOR2 (N778, N775, N607);
and AND4 (N779, N774, N443, N453, N340);
and AND3 (N780, N767, N264, N719);
buf BUF1 (N781, N758);
or OR2 (N782, N779, N538);
nor NOR2 (N783, N781, N703);
and AND4 (N784, N778, N746, N529, N493);
nor NOR2 (N785, N782, N718);
nor NOR2 (N786, N768, N225);
not NOT1 (N787, N780);
or OR2 (N788, N786, N577);
buf BUF1 (N789, N784);
nor NOR2 (N790, N769, N330);
or OR4 (N791, N787, N29, N93, N72);
not NOT1 (N792, N777);
and AND2 (N793, N789, N569);
nand NAND4 (N794, N792, N423, N237, N481);
nor NOR3 (N795, N776, N74, N288);
and AND2 (N796, N752, N291);
and AND3 (N797, N795, N53, N231);
xor XOR2 (N798, N797, N265);
and AND2 (N799, N798, N442);
buf BUF1 (N800, N790);
or OR4 (N801, N799, N220, N411, N662);
xor XOR2 (N802, N785, N531);
nor NOR3 (N803, N788, N415, N756);
xor XOR2 (N804, N793, N561);
nand NAND3 (N805, N803, N444, N656);
nor NOR4 (N806, N791, N386, N277, N211);
xor XOR2 (N807, N763, N325);
or OR4 (N808, N794, N557, N97, N424);
and AND4 (N809, N796, N711, N363, N27);
or OR4 (N810, N802, N294, N213, N619);
xor XOR2 (N811, N805, N220);
and AND4 (N812, N808, N700, N555, N769);
nand NAND2 (N813, N810, N714);
nor NOR2 (N814, N806, N115);
nor NOR3 (N815, N811, N211, N248);
not NOT1 (N816, N812);
and AND3 (N817, N800, N800, N768);
xor XOR2 (N818, N807, N679);
and AND2 (N819, N815, N586);
xor XOR2 (N820, N818, N412);
buf BUF1 (N821, N817);
xor XOR2 (N822, N809, N73);
not NOT1 (N823, N804);
not NOT1 (N824, N823);
nand NAND2 (N825, N813, N231);
nor NOR3 (N826, N816, N659, N384);
nor NOR2 (N827, N801, N46);
xor XOR2 (N828, N820, N748);
and AND4 (N829, N828, N1, N34, N260);
buf BUF1 (N830, N814);
nand NAND2 (N831, N829, N320);
buf BUF1 (N832, N830);
nor NOR3 (N833, N826, N371, N492);
nand NAND2 (N834, N833, N517);
and AND2 (N835, N825, N23);
or OR2 (N836, N831, N119);
xor XOR2 (N837, N835, N527);
nand NAND3 (N838, N824, N266, N364);
nor NOR4 (N839, N783, N578, N555, N713);
or OR4 (N840, N838, N269, N301, N737);
nor NOR3 (N841, N834, N519, N258);
not NOT1 (N842, N819);
not NOT1 (N843, N832);
nor NOR3 (N844, N822, N406, N663);
xor XOR2 (N845, N842, N653);
and AND2 (N846, N827, N5);
nand NAND4 (N847, N836, N461, N783, N149);
nor NOR3 (N848, N821, N593, N734);
buf BUF1 (N849, N847);
nand NAND4 (N850, N841, N213, N846, N568);
and AND2 (N851, N137, N37);
nand NAND3 (N852, N848, N318, N150);
xor XOR2 (N853, N845, N388);
or OR2 (N854, N844, N212);
nor NOR2 (N855, N839, N673);
or OR2 (N856, N852, N190);
xor XOR2 (N857, N855, N287);
or OR2 (N858, N843, N750);
buf BUF1 (N859, N856);
or OR2 (N860, N858, N112);
xor XOR2 (N861, N854, N646);
and AND4 (N862, N859, N675, N60, N172);
and AND3 (N863, N837, N27, N704);
xor XOR2 (N864, N850, N519);
not NOT1 (N865, N857);
buf BUF1 (N866, N865);
or OR4 (N867, N853, N341, N761, N203);
nand NAND3 (N868, N866, N674, N93);
nand NAND2 (N869, N867, N569);
or OR2 (N870, N849, N333);
or OR4 (N871, N864, N187, N664, N506);
nor NOR2 (N872, N851, N194);
not NOT1 (N873, N861);
nand NAND3 (N874, N868, N336, N471);
not NOT1 (N875, N871);
nor NOR2 (N876, N862, N358);
or OR2 (N877, N875, N321);
not NOT1 (N878, N860);
and AND4 (N879, N869, N662, N462, N683);
nor NOR2 (N880, N872, N389);
nor NOR4 (N881, N880, N374, N309, N562);
xor XOR2 (N882, N876, N159);
or OR4 (N883, N863, N746, N838, N404);
or OR4 (N884, N882, N61, N275, N238);
nor NOR2 (N885, N881, N573);
nor NOR4 (N886, N884, N547, N320, N581);
xor XOR2 (N887, N873, N873);
buf BUF1 (N888, N886);
buf BUF1 (N889, N887);
buf BUF1 (N890, N877);
nor NOR4 (N891, N879, N433, N758, N507);
or OR2 (N892, N883, N321);
xor XOR2 (N893, N888, N307);
buf BUF1 (N894, N891);
and AND2 (N895, N874, N93);
nand NAND4 (N896, N870, N342, N490, N490);
not NOT1 (N897, N894);
xor XOR2 (N898, N896, N94);
buf BUF1 (N899, N898);
buf BUF1 (N900, N897);
and AND2 (N901, N890, N761);
not NOT1 (N902, N901);
xor XOR2 (N903, N899, N786);
xor XOR2 (N904, N878, N44);
xor XOR2 (N905, N892, N646);
nor NOR4 (N906, N903, N501, N561, N822);
not NOT1 (N907, N905);
nand NAND3 (N908, N893, N454, N13);
not NOT1 (N909, N900);
nor NOR3 (N910, N889, N286, N311);
and AND2 (N911, N840, N503);
xor XOR2 (N912, N911, N679);
nor NOR2 (N913, N895, N286);
nand NAND2 (N914, N906, N104);
and AND2 (N915, N904, N281);
nor NOR2 (N916, N913, N327);
buf BUF1 (N917, N916);
not NOT1 (N918, N915);
buf BUF1 (N919, N918);
and AND4 (N920, N885, N55, N388, N13);
buf BUF1 (N921, N920);
not NOT1 (N922, N912);
not NOT1 (N923, N921);
nor NOR3 (N924, N907, N796, N708);
nand NAND2 (N925, N922, N567);
xor XOR2 (N926, N909, N524);
and AND3 (N927, N910, N155, N892);
not NOT1 (N928, N908);
nor NOR3 (N929, N928, N872, N309);
and AND4 (N930, N919, N296, N521, N123);
xor XOR2 (N931, N929, N205);
nand NAND2 (N932, N902, N143);
buf BUF1 (N933, N924);
not NOT1 (N934, N931);
xor XOR2 (N935, N923, N275);
or OR4 (N936, N933, N68, N469, N689);
or OR2 (N937, N927, N705);
not NOT1 (N938, N935);
or OR4 (N939, N925, N285, N824, N561);
buf BUF1 (N940, N926);
xor XOR2 (N941, N930, N323);
not NOT1 (N942, N938);
nor NOR4 (N943, N914, N748, N833, N88);
or OR4 (N944, N917, N73, N902, N364);
not NOT1 (N945, N932);
xor XOR2 (N946, N937, N790);
or OR2 (N947, N945, N226);
and AND2 (N948, N943, N375);
or OR4 (N949, N934, N578, N931, N825);
not NOT1 (N950, N940);
not NOT1 (N951, N949);
nor NOR3 (N952, N948, N888, N847);
not NOT1 (N953, N950);
not NOT1 (N954, N941);
not NOT1 (N955, N952);
not NOT1 (N956, N947);
nand NAND2 (N957, N946, N107);
or OR3 (N958, N955, N538, N111);
not NOT1 (N959, N956);
xor XOR2 (N960, N936, N524);
nor NOR3 (N961, N953, N234, N548);
and AND2 (N962, N942, N296);
buf BUF1 (N963, N957);
and AND4 (N964, N944, N610, N491, N260);
not NOT1 (N965, N958);
buf BUF1 (N966, N961);
or OR2 (N967, N962, N273);
nor NOR3 (N968, N967, N628, N932);
nand NAND4 (N969, N960, N618, N895, N163);
nand NAND4 (N970, N964, N840, N455, N684);
or OR2 (N971, N939, N820);
not NOT1 (N972, N963);
not NOT1 (N973, N954);
and AND3 (N974, N959, N739, N396);
not NOT1 (N975, N969);
nand NAND3 (N976, N970, N846, N144);
nand NAND3 (N977, N975, N918, N446);
not NOT1 (N978, N951);
and AND2 (N979, N978, N159);
xor XOR2 (N980, N965, N666);
xor XOR2 (N981, N968, N106);
or OR2 (N982, N980, N488);
or OR3 (N983, N976, N442, N485);
nor NOR2 (N984, N983, N363);
not NOT1 (N985, N979);
and AND4 (N986, N966, N358, N350, N955);
nand NAND2 (N987, N986, N176);
xor XOR2 (N988, N985, N109);
nand NAND2 (N989, N974, N879);
or OR4 (N990, N973, N739, N51, N339);
buf BUF1 (N991, N971);
and AND2 (N992, N981, N866);
xor XOR2 (N993, N987, N219);
nand NAND3 (N994, N984, N115, N367);
buf BUF1 (N995, N972);
and AND4 (N996, N989, N601, N653, N869);
or OR4 (N997, N993, N49, N879, N192);
nor NOR3 (N998, N995, N498, N27);
or OR2 (N999, N998, N646);
not NOT1 (N1000, N996);
nand NAND3 (N1001, N982, N111, N931);
buf BUF1 (N1002, N977);
nand NAND2 (N1003, N1000, N258);
and AND4 (N1004, N997, N905, N385, N532);
buf BUF1 (N1005, N988);
and AND4 (N1006, N1002, N140, N493, N975);
or OR3 (N1007, N1004, N128, N648);
nand NAND4 (N1008, N1001, N699, N978, N102);
nor NOR4 (N1009, N1003, N203, N222, N265);
not NOT1 (N1010, N1007);
buf BUF1 (N1011, N1006);
not NOT1 (N1012, N1008);
buf BUF1 (N1013, N994);
buf BUF1 (N1014, N991);
nand NAND3 (N1015, N990, N416, N88);
nor NOR2 (N1016, N1015, N653);
nand NAND4 (N1017, N999, N107, N542, N36);
nand NAND2 (N1018, N1010, N63);
nor NOR2 (N1019, N1017, N623);
and AND4 (N1020, N1009, N185, N744, N916);
and AND4 (N1021, N992, N53, N207, N317);
or OR2 (N1022, N1011, N288);
and AND3 (N1023, N1005, N170, N539);
and AND4 (N1024, N1023, N90, N217, N1018);
xor XOR2 (N1025, N9, N553);
buf BUF1 (N1026, N1019);
not NOT1 (N1027, N1022);
nor NOR3 (N1028, N1016, N703, N939);
not NOT1 (N1029, N1014);
and AND3 (N1030, N1025, N377, N29);
nand NAND4 (N1031, N1029, N460, N115, N50);
not NOT1 (N1032, N1031);
not NOT1 (N1033, N1030);
nand NAND3 (N1034, N1027, N831, N99);
or OR3 (N1035, N1021, N857, N127);
not NOT1 (N1036, N1034);
not NOT1 (N1037, N1026);
not NOT1 (N1038, N1013);
and AND2 (N1039, N1024, N973);
buf BUF1 (N1040, N1039);
or OR2 (N1041, N1020, N70);
buf BUF1 (N1042, N1041);
and AND2 (N1043, N1036, N101);
not NOT1 (N1044, N1033);
and AND3 (N1045, N1035, N718, N129);
xor XOR2 (N1046, N1044, N775);
or OR2 (N1047, N1042, N435);
not NOT1 (N1048, N1032);
nand NAND2 (N1049, N1038, N857);
buf BUF1 (N1050, N1040);
not NOT1 (N1051, N1012);
or OR3 (N1052, N1045, N927, N170);
nand NAND2 (N1053, N1049, N855);
nand NAND4 (N1054, N1028, N480, N1032, N446);
and AND4 (N1055, N1037, N1008, N421, N560);
or OR3 (N1056, N1050, N163, N977);
and AND4 (N1057, N1046, N557, N479, N628);
or OR2 (N1058, N1054, N1033);
and AND4 (N1059, N1055, N688, N869, N674);
not NOT1 (N1060, N1052);
or OR2 (N1061, N1053, N462);
buf BUF1 (N1062, N1047);
nor NOR4 (N1063, N1048, N141, N1004, N427);
or OR2 (N1064, N1062, N97);
buf BUF1 (N1065, N1064);
nor NOR2 (N1066, N1061, N857);
buf BUF1 (N1067, N1043);
xor XOR2 (N1068, N1067, N656);
not NOT1 (N1069, N1063);
nor NOR2 (N1070, N1051, N746);
not NOT1 (N1071, N1056);
nand NAND3 (N1072, N1069, N338, N733);
or OR4 (N1073, N1065, N960, N843, N538);
xor XOR2 (N1074, N1068, N334);
xor XOR2 (N1075, N1059, N612);
or OR2 (N1076, N1071, N301);
nand NAND2 (N1077, N1076, N363);
buf BUF1 (N1078, N1072);
nand NAND4 (N1079, N1073, N1002, N606, N182);
and AND2 (N1080, N1074, N962);
xor XOR2 (N1081, N1058, N213);
nor NOR3 (N1082, N1077, N771, N1060);
buf BUF1 (N1083, N1002);
nor NOR4 (N1084, N1080, N345, N754, N682);
and AND2 (N1085, N1078, N416);
nand NAND4 (N1086, N1079, N235, N607, N569);
nand NAND2 (N1087, N1085, N323);
not NOT1 (N1088, N1087);
and AND2 (N1089, N1057, N835);
xor XOR2 (N1090, N1066, N290);
nand NAND3 (N1091, N1089, N323, N995);
or OR3 (N1092, N1081, N775, N972);
nor NOR3 (N1093, N1075, N175, N928);
or OR4 (N1094, N1092, N742, N437, N960);
or OR3 (N1095, N1094, N976, N962);
xor XOR2 (N1096, N1084, N469);
buf BUF1 (N1097, N1088);
buf BUF1 (N1098, N1070);
buf BUF1 (N1099, N1090);
not NOT1 (N1100, N1095);
or OR3 (N1101, N1096, N103, N613);
not NOT1 (N1102, N1086);
buf BUF1 (N1103, N1099);
not NOT1 (N1104, N1091);
nand NAND2 (N1105, N1103, N342);
and AND3 (N1106, N1097, N878, N191);
buf BUF1 (N1107, N1093);
nor NOR3 (N1108, N1106, N623, N185);
nor NOR4 (N1109, N1098, N1107, N370, N896);
nand NAND3 (N1110, N233, N77, N570);
or OR2 (N1111, N1108, N614);
nand NAND3 (N1112, N1101, N124, N294);
xor XOR2 (N1113, N1105, N698);
xor XOR2 (N1114, N1109, N187);
and AND3 (N1115, N1110, N1079, N995);
nand NAND3 (N1116, N1104, N22, N572);
not NOT1 (N1117, N1083);
nand NAND4 (N1118, N1111, N828, N972, N4);
and AND4 (N1119, N1115, N775, N102, N299);
nand NAND2 (N1120, N1118, N858);
xor XOR2 (N1121, N1117, N166);
and AND3 (N1122, N1116, N765, N321);
buf BUF1 (N1123, N1102);
and AND2 (N1124, N1122, N251);
nor NOR3 (N1125, N1119, N526, N418);
nand NAND4 (N1126, N1125, N476, N328, N79);
or OR4 (N1127, N1100, N1118, N135, N622);
nor NOR2 (N1128, N1112, N1095);
xor XOR2 (N1129, N1128, N248);
nand NAND4 (N1130, N1114, N688, N971, N31);
and AND4 (N1131, N1126, N194, N834, N385);
or OR4 (N1132, N1131, N189, N567, N605);
nand NAND4 (N1133, N1123, N1022, N981, N685);
or OR4 (N1134, N1120, N812, N1092, N14);
nand NAND2 (N1135, N1129, N1021);
nand NAND3 (N1136, N1132, N121, N751);
not NOT1 (N1137, N1136);
buf BUF1 (N1138, N1130);
xor XOR2 (N1139, N1124, N248);
buf BUF1 (N1140, N1134);
nor NOR3 (N1141, N1139, N352, N312);
not NOT1 (N1142, N1082);
nand NAND2 (N1143, N1135, N629);
nor NOR4 (N1144, N1121, N1025, N117, N260);
buf BUF1 (N1145, N1141);
and AND2 (N1146, N1133, N60);
xor XOR2 (N1147, N1113, N178);
not NOT1 (N1148, N1144);
not NOT1 (N1149, N1145);
nand NAND3 (N1150, N1127, N1049, N701);
xor XOR2 (N1151, N1150, N106);
buf BUF1 (N1152, N1149);
buf BUF1 (N1153, N1138);
nor NOR2 (N1154, N1137, N32);
nand NAND4 (N1155, N1151, N1083, N680, N299);
or OR2 (N1156, N1153, N272);
nand NAND2 (N1157, N1147, N901);
buf BUF1 (N1158, N1157);
buf BUF1 (N1159, N1146);
not NOT1 (N1160, N1159);
or OR4 (N1161, N1140, N47, N537, N681);
nor NOR3 (N1162, N1142, N764, N630);
or OR3 (N1163, N1152, N859, N586);
and AND2 (N1164, N1148, N173);
not NOT1 (N1165, N1158);
or OR2 (N1166, N1154, N108);
or OR3 (N1167, N1164, N286, N646);
not NOT1 (N1168, N1155);
not NOT1 (N1169, N1143);
nand NAND4 (N1170, N1168, N406, N981, N1101);
nand NAND4 (N1171, N1163, N685, N114, N901);
buf BUF1 (N1172, N1165);
or OR3 (N1173, N1160, N457, N799);
and AND2 (N1174, N1161, N667);
or OR4 (N1175, N1162, N961, N990, N372);
or OR2 (N1176, N1166, N561);
buf BUF1 (N1177, N1170);
nand NAND2 (N1178, N1176, N164);
and AND3 (N1179, N1177, N1105, N820);
nor NOR2 (N1180, N1175, N144);
nand NAND2 (N1181, N1178, N1125);
not NOT1 (N1182, N1172);
nor NOR4 (N1183, N1173, N946, N813, N823);
nor NOR2 (N1184, N1167, N384);
buf BUF1 (N1185, N1174);
not NOT1 (N1186, N1156);
and AND3 (N1187, N1180, N514, N656);
not NOT1 (N1188, N1186);
nor NOR4 (N1189, N1171, N1150, N440, N886);
nand NAND4 (N1190, N1182, N104, N824, N1179);
nor NOR3 (N1191, N827, N621, N640);
xor XOR2 (N1192, N1190, N904);
and AND4 (N1193, N1187, N403, N1021, N893);
and AND4 (N1194, N1191, N464, N533, N722);
xor XOR2 (N1195, N1193, N1030);
nor NOR2 (N1196, N1194, N373);
and AND3 (N1197, N1189, N235, N176);
nand NAND4 (N1198, N1192, N991, N546, N840);
buf BUF1 (N1199, N1181);
or OR4 (N1200, N1199, N884, N246, N856);
nor NOR2 (N1201, N1200, N778);
or OR2 (N1202, N1185, N698);
xor XOR2 (N1203, N1195, N823);
nand NAND2 (N1204, N1184, N930);
or OR4 (N1205, N1204, N951, N824, N75);
nor NOR2 (N1206, N1188, N912);
nor NOR2 (N1207, N1205, N1200);
or OR4 (N1208, N1169, N1042, N39, N17);
buf BUF1 (N1209, N1183);
not NOT1 (N1210, N1198);
or OR3 (N1211, N1202, N1050, N1049);
nand NAND4 (N1212, N1203, N644, N859, N315);
nor NOR2 (N1213, N1211, N640);
nor NOR2 (N1214, N1209, N733);
and AND3 (N1215, N1213, N601, N190);
not NOT1 (N1216, N1210);
nor NOR2 (N1217, N1212, N58);
nand NAND3 (N1218, N1217, N472, N706);
and AND4 (N1219, N1207, N840, N1141, N824);
nor NOR2 (N1220, N1215, N1163);
xor XOR2 (N1221, N1220, N1028);
buf BUF1 (N1222, N1196);
buf BUF1 (N1223, N1218);
buf BUF1 (N1224, N1221);
buf BUF1 (N1225, N1214);
and AND4 (N1226, N1206, N520, N257, N760);
buf BUF1 (N1227, N1197);
or OR4 (N1228, N1227, N957, N641, N775);
nor NOR2 (N1229, N1201, N234);
nor NOR2 (N1230, N1216, N255);
not NOT1 (N1231, N1226);
nand NAND2 (N1232, N1230, N876);
or OR4 (N1233, N1228, N845, N103, N351);
nand NAND3 (N1234, N1232, N671, N254);
or OR4 (N1235, N1231, N563, N383, N261);
nor NOR2 (N1236, N1222, N1217);
or OR3 (N1237, N1223, N145, N1118);
or OR2 (N1238, N1237, N317);
not NOT1 (N1239, N1224);
buf BUF1 (N1240, N1233);
buf BUF1 (N1241, N1234);
not NOT1 (N1242, N1229);
xor XOR2 (N1243, N1241, N193);
and AND3 (N1244, N1208, N1207, N287);
and AND3 (N1245, N1242, N1130, N345);
nor NOR2 (N1246, N1245, N324);
and AND2 (N1247, N1219, N961);
nor NOR4 (N1248, N1247, N953, N448, N805);
not NOT1 (N1249, N1235);
nand NAND2 (N1250, N1248, N1098);
and AND2 (N1251, N1239, N63);
nand NAND4 (N1252, N1246, N453, N684, N84);
nor NOR3 (N1253, N1250, N481, N608);
not NOT1 (N1254, N1238);
nand NAND3 (N1255, N1240, N905, N1228);
buf BUF1 (N1256, N1253);
buf BUF1 (N1257, N1243);
xor XOR2 (N1258, N1244, N882);
not NOT1 (N1259, N1256);
nand NAND2 (N1260, N1259, N1136);
xor XOR2 (N1261, N1225, N962);
not NOT1 (N1262, N1254);
or OR2 (N1263, N1252, N1016);
or OR4 (N1264, N1260, N1156, N49, N1134);
xor XOR2 (N1265, N1263, N39);
or OR2 (N1266, N1249, N478);
nor NOR3 (N1267, N1258, N376, N610);
xor XOR2 (N1268, N1255, N987);
buf BUF1 (N1269, N1261);
or OR2 (N1270, N1236, N967);
nor NOR2 (N1271, N1257, N1021);
not NOT1 (N1272, N1251);
xor XOR2 (N1273, N1264, N840);
nand NAND3 (N1274, N1272, N211, N1150);
buf BUF1 (N1275, N1274);
or OR3 (N1276, N1262, N1173, N853);
and AND4 (N1277, N1266, N828, N784, N212);
xor XOR2 (N1278, N1270, N163);
nand NAND3 (N1279, N1267, N786, N473);
and AND4 (N1280, N1269, N865, N870, N346);
buf BUF1 (N1281, N1279);
nor NOR3 (N1282, N1275, N1141, N668);
and AND2 (N1283, N1281, N3);
buf BUF1 (N1284, N1280);
buf BUF1 (N1285, N1265);
buf BUF1 (N1286, N1282);
nand NAND2 (N1287, N1277, N1046);
nand NAND3 (N1288, N1283, N110, N806);
and AND2 (N1289, N1271, N758);
and AND2 (N1290, N1288, N172);
nand NAND3 (N1291, N1284, N834, N12);
nand NAND3 (N1292, N1290, N1157, N201);
and AND3 (N1293, N1291, N881, N117);
nand NAND3 (N1294, N1293, N15, N680);
buf BUF1 (N1295, N1273);
not NOT1 (N1296, N1276);
or OR3 (N1297, N1289, N1101, N666);
nor NOR2 (N1298, N1296, N11);
buf BUF1 (N1299, N1268);
or OR2 (N1300, N1287, N275);
xor XOR2 (N1301, N1299, N479);
nor NOR4 (N1302, N1285, N876, N177, N17);
and AND3 (N1303, N1278, N682, N425);
not NOT1 (N1304, N1292);
or OR2 (N1305, N1286, N544);
and AND2 (N1306, N1295, N697);
nand NAND2 (N1307, N1302, N401);
or OR3 (N1308, N1304, N366, N229);
buf BUF1 (N1309, N1308);
nand NAND3 (N1310, N1298, N828, N947);
and AND2 (N1311, N1300, N49);
and AND3 (N1312, N1311, N407, N876);
and AND2 (N1313, N1309, N345);
nor NOR2 (N1314, N1312, N504);
xor XOR2 (N1315, N1306, N77);
buf BUF1 (N1316, N1307);
buf BUF1 (N1317, N1301);
buf BUF1 (N1318, N1314);
not NOT1 (N1319, N1294);
not NOT1 (N1320, N1315);
or OR4 (N1321, N1310, N656, N1030, N668);
not NOT1 (N1322, N1305);
and AND2 (N1323, N1317, N338);
and AND4 (N1324, N1319, N234, N35, N822);
or OR2 (N1325, N1297, N855);
not NOT1 (N1326, N1324);
xor XOR2 (N1327, N1303, N1026);
not NOT1 (N1328, N1321);
nor NOR2 (N1329, N1316, N84);
not NOT1 (N1330, N1329);
xor XOR2 (N1331, N1326, N1256);
or OR2 (N1332, N1331, N1058);
not NOT1 (N1333, N1327);
buf BUF1 (N1334, N1325);
nor NOR3 (N1335, N1328, N440, N676);
not NOT1 (N1336, N1333);
nor NOR3 (N1337, N1318, N290, N1228);
buf BUF1 (N1338, N1332);
nor NOR3 (N1339, N1323, N591, N1121);
nor NOR2 (N1340, N1334, N1049);
and AND2 (N1341, N1340, N1290);
not NOT1 (N1342, N1320);
or OR3 (N1343, N1342, N667, N394);
or OR4 (N1344, N1322, N1284, N396, N1247);
xor XOR2 (N1345, N1338, N742);
not NOT1 (N1346, N1343);
not NOT1 (N1347, N1341);
nor NOR4 (N1348, N1347, N67, N1238, N1000);
and AND2 (N1349, N1330, N682);
xor XOR2 (N1350, N1339, N492);
nor NOR3 (N1351, N1335, N679, N305);
or OR4 (N1352, N1345, N591, N128, N1101);
xor XOR2 (N1353, N1349, N489);
buf BUF1 (N1354, N1352);
nand NAND2 (N1355, N1313, N179);
and AND2 (N1356, N1346, N1191);
and AND2 (N1357, N1350, N1175);
not NOT1 (N1358, N1357);
nand NAND2 (N1359, N1356, N1341);
nor NOR2 (N1360, N1353, N268);
buf BUF1 (N1361, N1344);
nand NAND3 (N1362, N1348, N549, N1010);
buf BUF1 (N1363, N1354);
nand NAND2 (N1364, N1351, N1067);
nand NAND2 (N1365, N1358, N1313);
not NOT1 (N1366, N1336);
and AND3 (N1367, N1355, N639, N374);
xor XOR2 (N1368, N1359, N568);
and AND3 (N1369, N1360, N168, N757);
not NOT1 (N1370, N1367);
buf BUF1 (N1371, N1370);
and AND4 (N1372, N1368, N822, N1133, N1055);
or OR3 (N1373, N1364, N820, N1304);
nand NAND3 (N1374, N1362, N250, N738);
or OR3 (N1375, N1363, N933, N676);
not NOT1 (N1376, N1365);
buf BUF1 (N1377, N1372);
and AND4 (N1378, N1373, N790, N1361, N317);
nor NOR4 (N1379, N638, N597, N669, N508);
and AND3 (N1380, N1374, N1005, N286);
and AND4 (N1381, N1371, N1076, N277, N1182);
xor XOR2 (N1382, N1376, N949);
nor NOR2 (N1383, N1375, N744);
and AND3 (N1384, N1380, N1065, N144);
nand NAND3 (N1385, N1379, N1071, N27);
buf BUF1 (N1386, N1384);
buf BUF1 (N1387, N1383);
not NOT1 (N1388, N1385);
nor NOR4 (N1389, N1378, N1295, N504, N767);
nor NOR3 (N1390, N1377, N1367, N193);
not NOT1 (N1391, N1381);
not NOT1 (N1392, N1387);
and AND3 (N1393, N1386, N896, N975);
xor XOR2 (N1394, N1382, N1053);
and AND2 (N1395, N1391, N1102);
nand NAND3 (N1396, N1369, N910, N286);
or OR2 (N1397, N1366, N487);
nand NAND2 (N1398, N1390, N608);
nand NAND2 (N1399, N1398, N875);
nand NAND4 (N1400, N1397, N275, N1012, N105);
not NOT1 (N1401, N1395);
not NOT1 (N1402, N1388);
and AND2 (N1403, N1401, N360);
or OR2 (N1404, N1394, N207);
nand NAND2 (N1405, N1399, N725);
nor NOR2 (N1406, N1403, N1245);
nand NAND4 (N1407, N1405, N1397, N585, N241);
and AND2 (N1408, N1393, N1178);
buf BUF1 (N1409, N1389);
and AND2 (N1410, N1392, N273);
not NOT1 (N1411, N1406);
buf BUF1 (N1412, N1400);
or OR4 (N1413, N1411, N950, N443, N35);
buf BUF1 (N1414, N1409);
buf BUF1 (N1415, N1404);
and AND4 (N1416, N1414, N505, N987, N1246);
not NOT1 (N1417, N1410);
not NOT1 (N1418, N1413);
nand NAND3 (N1419, N1418, N1344, N320);
not NOT1 (N1420, N1402);
buf BUF1 (N1421, N1416);
and AND3 (N1422, N1417, N623, N7);
nand NAND2 (N1423, N1412, N25);
nand NAND2 (N1424, N1337, N1145);
nand NAND4 (N1425, N1420, N1227, N1283, N1419);
nor NOR4 (N1426, N55, N1348, N405, N211);
nor NOR2 (N1427, N1421, N694);
not NOT1 (N1428, N1423);
nor NOR4 (N1429, N1428, N1114, N168, N372);
or OR2 (N1430, N1408, N1139);
nor NOR3 (N1431, N1396, N326, N1090);
xor XOR2 (N1432, N1424, N438);
or OR2 (N1433, N1425, N666);
and AND2 (N1434, N1427, N698);
nor NOR4 (N1435, N1422, N9, N167, N1050);
or OR3 (N1436, N1435, N476, N536);
and AND3 (N1437, N1432, N424, N527);
nand NAND3 (N1438, N1436, N72, N582);
and AND2 (N1439, N1437, N578);
or OR3 (N1440, N1439, N130, N144);
or OR3 (N1441, N1438, N698, N1375);
nand NAND4 (N1442, N1433, N304, N45, N74);
nor NOR3 (N1443, N1407, N435, N955);
buf BUF1 (N1444, N1441);
not NOT1 (N1445, N1444);
or OR3 (N1446, N1415, N168, N383);
xor XOR2 (N1447, N1434, N560);
or OR3 (N1448, N1447, N1037, N571);
and AND4 (N1449, N1448, N559, N1359, N797);
xor XOR2 (N1450, N1430, N1182);
xor XOR2 (N1451, N1443, N900);
and AND2 (N1452, N1445, N346);
or OR3 (N1453, N1440, N1062, N1227);
not NOT1 (N1454, N1452);
xor XOR2 (N1455, N1431, N649);
buf BUF1 (N1456, N1455);
and AND4 (N1457, N1451, N852, N608, N95);
xor XOR2 (N1458, N1450, N267);
nor NOR2 (N1459, N1446, N209);
buf BUF1 (N1460, N1458);
nand NAND4 (N1461, N1426, N663, N992, N149);
buf BUF1 (N1462, N1460);
and AND4 (N1463, N1454, N585, N1364, N818);
or OR3 (N1464, N1456, N414, N986);
not NOT1 (N1465, N1449);
or OR2 (N1466, N1461, N194);
and AND4 (N1467, N1465, N208, N172, N77);
not NOT1 (N1468, N1429);
nor NOR4 (N1469, N1464, N1, N948, N182);
or OR4 (N1470, N1467, N441, N288, N180);
not NOT1 (N1471, N1463);
nand NAND3 (N1472, N1466, N874, N202);
not NOT1 (N1473, N1471);
and AND2 (N1474, N1459, N652);
xor XOR2 (N1475, N1442, N349);
not NOT1 (N1476, N1470);
or OR4 (N1477, N1462, N285, N243, N48);
nor NOR4 (N1478, N1453, N449, N974, N46);
and AND3 (N1479, N1474, N73, N483);
and AND3 (N1480, N1468, N934, N8);
and AND2 (N1481, N1469, N691);
nand NAND3 (N1482, N1472, N1344, N523);
nand NAND2 (N1483, N1480, N518);
xor XOR2 (N1484, N1482, N836);
nor NOR3 (N1485, N1479, N974, N832);
buf BUF1 (N1486, N1484);
nand NAND2 (N1487, N1457, N376);
and AND4 (N1488, N1475, N1024, N525, N626);
not NOT1 (N1489, N1485);
xor XOR2 (N1490, N1476, N601);
nand NAND3 (N1491, N1486, N601, N912);
buf BUF1 (N1492, N1483);
nor NOR3 (N1493, N1481, N1351, N1143);
xor XOR2 (N1494, N1491, N1058);
not NOT1 (N1495, N1477);
and AND4 (N1496, N1473, N1229, N435, N911);
nor NOR4 (N1497, N1493, N362, N596, N467);
not NOT1 (N1498, N1489);
nor NOR2 (N1499, N1495, N1369);
xor XOR2 (N1500, N1488, N1319);
nor NOR4 (N1501, N1490, N1458, N384, N323);
xor XOR2 (N1502, N1500, N42);
and AND4 (N1503, N1496, N1277, N418, N1465);
buf BUF1 (N1504, N1487);
xor XOR2 (N1505, N1492, N21);
and AND3 (N1506, N1505, N1236, N1461);
nor NOR4 (N1507, N1503, N516, N973, N383);
nor NOR2 (N1508, N1506, N732);
xor XOR2 (N1509, N1494, N1417);
nand NAND3 (N1510, N1502, N743, N1116);
buf BUF1 (N1511, N1499);
buf BUF1 (N1512, N1509);
nor NOR2 (N1513, N1511, N821);
nor NOR2 (N1514, N1497, N805);
or OR4 (N1515, N1514, N48, N1332, N1509);
or OR4 (N1516, N1510, N452, N998, N376);
nand NAND3 (N1517, N1513, N1112, N664);
nand NAND3 (N1518, N1504, N1409, N437);
or OR3 (N1519, N1518, N1372, N83);
buf BUF1 (N1520, N1508);
and AND4 (N1521, N1519, N1008, N1396, N927);
or OR3 (N1522, N1478, N381, N395);
not NOT1 (N1523, N1498);
not NOT1 (N1524, N1523);
not NOT1 (N1525, N1501);
nor NOR2 (N1526, N1524, N1035);
buf BUF1 (N1527, N1522);
xor XOR2 (N1528, N1527, N428);
not NOT1 (N1529, N1526);
or OR4 (N1530, N1512, N1291, N622, N1347);
nand NAND2 (N1531, N1528, N63);
not NOT1 (N1532, N1516);
nor NOR4 (N1533, N1521, N766, N506, N798);
nor NOR3 (N1534, N1520, N983, N36);
or OR4 (N1535, N1530, N1085, N318, N976);
nor NOR2 (N1536, N1515, N631);
xor XOR2 (N1537, N1532, N1515);
xor XOR2 (N1538, N1535, N405);
not NOT1 (N1539, N1529);
nor NOR3 (N1540, N1537, N1499, N994);
and AND2 (N1541, N1525, N537);
or OR4 (N1542, N1517, N991, N899, N1196);
buf BUF1 (N1543, N1531);
or OR4 (N1544, N1541, N102, N1100, N1227);
buf BUF1 (N1545, N1533);
nand NAND2 (N1546, N1534, N643);
nor NOR2 (N1547, N1543, N1346);
and AND2 (N1548, N1539, N1298);
nand NAND3 (N1549, N1544, N1406, N1169);
buf BUF1 (N1550, N1546);
or OR4 (N1551, N1550, N1489, N486, N988);
nand NAND4 (N1552, N1549, N870, N1137, N860);
buf BUF1 (N1553, N1551);
nand NAND4 (N1554, N1552, N80, N630, N535);
nor NOR3 (N1555, N1548, N295, N254);
not NOT1 (N1556, N1540);
nand NAND3 (N1557, N1545, N1250, N1227);
buf BUF1 (N1558, N1507);
nor NOR3 (N1559, N1555, N298, N1116);
nand NAND4 (N1560, N1558, N483, N1401, N57);
nor NOR3 (N1561, N1547, N626, N1558);
buf BUF1 (N1562, N1560);
not NOT1 (N1563, N1554);
nor NOR2 (N1564, N1538, N1327);
not NOT1 (N1565, N1556);
xor XOR2 (N1566, N1553, N1546);
and AND2 (N1567, N1536, N20);
nand NAND2 (N1568, N1557, N525);
not NOT1 (N1569, N1567);
buf BUF1 (N1570, N1565);
xor XOR2 (N1571, N1561, N1512);
or OR3 (N1572, N1562, N599, N1196);
nor NOR2 (N1573, N1571, N1030);
nor NOR2 (N1574, N1566, N1153);
xor XOR2 (N1575, N1574, N702);
xor XOR2 (N1576, N1542, N1285);
xor XOR2 (N1577, N1569, N63);
not NOT1 (N1578, N1575);
nor NOR3 (N1579, N1559, N195, N1327);
xor XOR2 (N1580, N1576, N136);
xor XOR2 (N1581, N1577, N554);
nor NOR3 (N1582, N1579, N140, N1114);
not NOT1 (N1583, N1563);
xor XOR2 (N1584, N1582, N1154);
buf BUF1 (N1585, N1568);
not NOT1 (N1586, N1581);
xor XOR2 (N1587, N1564, N1461);
not NOT1 (N1588, N1584);
nand NAND2 (N1589, N1572, N48);
nand NAND3 (N1590, N1586, N754, N990);
xor XOR2 (N1591, N1570, N764);
xor XOR2 (N1592, N1588, N1136);
and AND3 (N1593, N1585, N517, N438);
nand NAND2 (N1594, N1592, N882);
nand NAND3 (N1595, N1589, N1579, N28);
buf BUF1 (N1596, N1578);
xor XOR2 (N1597, N1587, N1397);
buf BUF1 (N1598, N1596);
or OR4 (N1599, N1590, N1507, N643, N890);
nand NAND2 (N1600, N1583, N675);
or OR4 (N1601, N1600, N248, N1392, N648);
or OR2 (N1602, N1573, N74);
nand NAND4 (N1603, N1598, N547, N1411, N18);
nand NAND2 (N1604, N1595, N1127);
or OR2 (N1605, N1593, N63);
and AND4 (N1606, N1580, N901, N260, N1580);
not NOT1 (N1607, N1604);
nand NAND3 (N1608, N1607, N852, N1203);
and AND2 (N1609, N1591, N1286);
nor NOR4 (N1610, N1609, N899, N1424, N376);
buf BUF1 (N1611, N1601);
not NOT1 (N1612, N1605);
and AND2 (N1613, N1597, N1297);
or OR3 (N1614, N1610, N943, N123);
nor NOR2 (N1615, N1614, N750);
nand NAND4 (N1616, N1594, N607, N1585, N1020);
and AND3 (N1617, N1612, N860, N1602);
nand NAND4 (N1618, N478, N1374, N408, N1041);
nand NAND4 (N1619, N1616, N847, N549, N865);
and AND4 (N1620, N1613, N684, N1128, N1617);
buf BUF1 (N1621, N207);
endmodule