// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;

output N4023,N4005,N4004,N4022,N4019,N4011,N4021,N4017,N4003,N4024;

or OR2 (N25, N23, N5);
buf BUF1 (N26, N19);
nor NOR4 (N27, N17, N16, N12, N4);
not NOT1 (N28, N12);
and AND3 (N29, N16, N9, N13);
nand NAND2 (N30, N13, N23);
nor NOR2 (N31, N25, N4);
not NOT1 (N32, N27);
nor NOR4 (N33, N27, N24, N30, N2);
and AND2 (N34, N29, N18);
buf BUF1 (N35, N3);
xor XOR2 (N36, N3, N10);
nand NAND2 (N37, N4, N13);
buf BUF1 (N38, N22);
nand NAND2 (N39, N33, N19);
or OR2 (N40, N35, N3);
buf BUF1 (N41, N37);
or OR4 (N42, N40, N11, N35, N41);
not NOT1 (N43, N26);
xor XOR2 (N44, N2, N1);
xor XOR2 (N45, N44, N36);
nor NOR2 (N46, N34, N4);
nor NOR3 (N47, N8, N10, N2);
buf BUF1 (N48, N38);
nor NOR4 (N49, N45, N34, N45, N41);
xor XOR2 (N50, N49, N5);
not NOT1 (N51, N32);
not NOT1 (N52, N28);
not NOT1 (N53, N42);
nand NAND2 (N54, N39, N18);
xor XOR2 (N55, N52, N34);
xor XOR2 (N56, N47, N24);
buf BUF1 (N57, N46);
xor XOR2 (N58, N50, N31);
nor NOR3 (N59, N13, N47, N23);
and AND4 (N60, N59, N30, N54, N20);
nand NAND2 (N61, N52, N14);
and AND3 (N62, N58, N34, N38);
not NOT1 (N63, N61);
xor XOR2 (N64, N63, N47);
and AND4 (N65, N64, N10, N37, N39);
nand NAND4 (N66, N56, N10, N31, N14);
not NOT1 (N67, N60);
buf BUF1 (N68, N55);
nand NAND3 (N69, N68, N20, N67);
and AND2 (N70, N53, N61);
or OR4 (N71, N3, N64, N54, N60);
xor XOR2 (N72, N57, N36);
not NOT1 (N73, N62);
and AND3 (N74, N51, N12, N43);
buf BUF1 (N75, N50);
or OR2 (N76, N70, N4);
and AND4 (N77, N74, N18, N10, N14);
nor NOR3 (N78, N73, N6, N15);
nand NAND4 (N79, N71, N34, N37, N33);
nor NOR2 (N80, N78, N12);
xor XOR2 (N81, N75, N61);
xor XOR2 (N82, N48, N13);
not NOT1 (N83, N66);
nand NAND2 (N84, N82, N33);
or OR3 (N85, N81, N25, N47);
nor NOR3 (N86, N83, N6, N53);
or OR4 (N87, N79, N64, N27, N76);
xor XOR2 (N88, N60, N35);
nor NOR4 (N89, N84, N9, N44, N78);
nand NAND3 (N90, N89, N37, N85);
or OR4 (N91, N26, N80, N37, N90);
buf BUF1 (N92, N63);
or OR4 (N93, N36, N63, N69, N70);
xor XOR2 (N94, N92, N4);
not NOT1 (N95, N37);
not NOT1 (N96, N77);
not NOT1 (N97, N72);
or OR4 (N98, N97, N35, N81, N92);
nor NOR4 (N99, N93, N89, N6, N53);
nand NAND2 (N100, N96, N9);
buf BUF1 (N101, N99);
xor XOR2 (N102, N65, N16);
and AND3 (N103, N95, N51, N4);
buf BUF1 (N104, N102);
buf BUF1 (N105, N86);
nand NAND4 (N106, N88, N81, N102, N9);
xor XOR2 (N107, N94, N26);
not NOT1 (N108, N103);
nand NAND3 (N109, N106, N97, N79);
buf BUF1 (N110, N107);
nand NAND3 (N111, N105, N89, N3);
and AND4 (N112, N100, N39, N15, N68);
buf BUF1 (N113, N109);
and AND3 (N114, N87, N93, N107);
nor NOR2 (N115, N101, N108);
xor XOR2 (N116, N27, N80);
not NOT1 (N117, N115);
and AND2 (N118, N112, N102);
or OR4 (N119, N116, N101, N99, N111);
xor XOR2 (N120, N36, N54);
nand NAND3 (N121, N114, N46, N103);
and AND2 (N122, N110, N121);
xor XOR2 (N123, N19, N77);
xor XOR2 (N124, N122, N38);
nor NOR3 (N125, N119, N37, N58);
xor XOR2 (N126, N104, N81);
buf BUF1 (N127, N113);
or OR4 (N128, N127, N51, N40, N66);
and AND3 (N129, N128, N100, N23);
not NOT1 (N130, N120);
nand NAND4 (N131, N91, N86, N108, N124);
xor XOR2 (N132, N77, N80);
xor XOR2 (N133, N118, N89);
nor NOR3 (N134, N123, N77, N83);
buf BUF1 (N135, N131);
nand NAND4 (N136, N130, N57, N48, N9);
or OR2 (N137, N126, N34);
and AND2 (N138, N135, N25);
buf BUF1 (N139, N125);
nand NAND3 (N140, N117, N127, N31);
and AND4 (N141, N138, N88, N54, N13);
not NOT1 (N142, N132);
or OR3 (N143, N98, N24, N48);
nor NOR4 (N144, N133, N137, N82, N24);
not NOT1 (N145, N132);
nor NOR3 (N146, N139, N63, N33);
or OR4 (N147, N146, N141, N8, N132);
xor XOR2 (N148, N70, N113);
nand NAND3 (N149, N144, N95, N64);
nor NOR2 (N150, N136, N75);
nor NOR4 (N151, N142, N72, N146, N4);
nand NAND3 (N152, N148, N48, N69);
or OR3 (N153, N152, N147, N67);
and AND2 (N154, N76, N152);
or OR4 (N155, N151, N137, N46, N119);
xor XOR2 (N156, N154, N146);
not NOT1 (N157, N143);
not NOT1 (N158, N145);
xor XOR2 (N159, N153, N67);
buf BUF1 (N160, N134);
nand NAND3 (N161, N159, N77, N67);
xor XOR2 (N162, N157, N47);
buf BUF1 (N163, N156);
and AND2 (N164, N155, N70);
or OR2 (N165, N140, N156);
xor XOR2 (N166, N165, N24);
xor XOR2 (N167, N162, N136);
and AND3 (N168, N166, N56, N141);
not NOT1 (N169, N158);
or OR2 (N170, N167, N60);
nand NAND4 (N171, N160, N47, N139, N62);
not NOT1 (N172, N171);
buf BUF1 (N173, N149);
and AND4 (N174, N161, N77, N55, N110);
not NOT1 (N175, N150);
nand NAND4 (N176, N129, N131, N155, N95);
or OR4 (N177, N173, N99, N135, N143);
buf BUF1 (N178, N175);
or OR4 (N179, N178, N63, N85, N174);
and AND3 (N180, N69, N148, N49);
nand NAND3 (N181, N176, N110, N103);
or OR3 (N182, N180, N34, N64);
buf BUF1 (N183, N182);
nor NOR4 (N184, N168, N34, N124, N58);
xor XOR2 (N185, N177, N73);
and AND4 (N186, N181, N163, N50, N42);
or OR2 (N187, N142, N84);
buf BUF1 (N188, N179);
nand NAND4 (N189, N186, N130, N83, N115);
and AND2 (N190, N172, N131);
xor XOR2 (N191, N188, N63);
nor NOR2 (N192, N184, N25);
buf BUF1 (N193, N170);
or OR3 (N194, N169, N120, N177);
nand NAND2 (N195, N183, N58);
or OR2 (N196, N193, N112);
nand NAND2 (N197, N192, N57);
not NOT1 (N198, N194);
xor XOR2 (N199, N189, N4);
not NOT1 (N200, N196);
or OR2 (N201, N187, N49);
and AND3 (N202, N198, N62, N38);
buf BUF1 (N203, N185);
buf BUF1 (N204, N202);
not NOT1 (N205, N201);
buf BUF1 (N206, N200);
nor NOR2 (N207, N164, N90);
nand NAND2 (N208, N204, N78);
and AND4 (N209, N199, N33, N203, N172);
nand NAND4 (N210, N108, N55, N166, N68);
xor XOR2 (N211, N205, N128);
xor XOR2 (N212, N207, N27);
or OR2 (N213, N197, N76);
nand NAND3 (N214, N213, N204, N138);
nand NAND2 (N215, N191, N18);
nand NAND2 (N216, N190, N118);
nand NAND4 (N217, N206, N28, N11, N216);
and AND4 (N218, N185, N34, N209, N162);
xor XOR2 (N219, N169, N28);
nor NOR4 (N220, N195, N110, N206, N44);
and AND4 (N221, N212, N73, N65, N34);
or OR3 (N222, N221, N130, N161);
nor NOR3 (N223, N215, N22, N27);
or OR2 (N224, N219, N54);
xor XOR2 (N225, N214, N74);
not NOT1 (N226, N217);
buf BUF1 (N227, N218);
buf BUF1 (N228, N211);
buf BUF1 (N229, N223);
and AND4 (N230, N224, N179, N198, N223);
xor XOR2 (N231, N226, N103);
or OR3 (N232, N231, N174, N169);
and AND2 (N233, N228, N221);
not NOT1 (N234, N232);
or OR4 (N235, N225, N172, N196, N3);
nand NAND4 (N236, N233, N212, N193, N132);
or OR2 (N237, N229, N35);
not NOT1 (N238, N227);
buf BUF1 (N239, N237);
nand NAND4 (N240, N239, N21, N82, N45);
nor NOR2 (N241, N236, N4);
nor NOR3 (N242, N238, N60, N101);
nand NAND4 (N243, N241, N41, N183, N16);
not NOT1 (N244, N230);
nor NOR3 (N245, N240, N59, N18);
nor NOR3 (N246, N208, N205, N7);
buf BUF1 (N247, N245);
nor NOR2 (N248, N220, N73);
not NOT1 (N249, N234);
buf BUF1 (N250, N222);
nand NAND4 (N251, N210, N95, N242, N210);
buf BUF1 (N252, N91);
nand NAND4 (N253, N252, N23, N44, N2);
nand NAND2 (N254, N243, N192);
buf BUF1 (N255, N248);
nor NOR2 (N256, N247, N236);
nand NAND3 (N257, N251, N61, N205);
nand NAND2 (N258, N254, N176);
and AND2 (N259, N249, N245);
nand NAND4 (N260, N256, N100, N241, N19);
nand NAND4 (N261, N259, N111, N244, N21);
nor NOR3 (N262, N38, N231, N138);
buf BUF1 (N263, N261);
nor NOR3 (N264, N263, N213, N37);
nor NOR4 (N265, N235, N182, N173, N162);
buf BUF1 (N266, N253);
buf BUF1 (N267, N262);
nand NAND2 (N268, N267, N226);
nand NAND2 (N269, N260, N204);
nand NAND4 (N270, N264, N97, N236, N211);
and AND2 (N271, N270, N92);
xor XOR2 (N272, N268, N15);
nand NAND2 (N273, N272, N111);
nand NAND4 (N274, N271, N99, N125, N230);
nor NOR3 (N275, N266, N192, N260);
buf BUF1 (N276, N258);
nand NAND4 (N277, N257, N276, N163, N245);
nand NAND2 (N278, N172, N226);
nand NAND4 (N279, N265, N55, N260, N165);
and AND2 (N280, N274, N175);
nand NAND4 (N281, N275, N174, N136, N144);
xor XOR2 (N282, N246, N102);
or OR2 (N283, N280, N215);
nand NAND4 (N284, N283, N49, N244, N63);
buf BUF1 (N285, N281);
or OR4 (N286, N250, N125, N263, N256);
or OR3 (N287, N285, N266, N21);
not NOT1 (N288, N284);
not NOT1 (N289, N255);
xor XOR2 (N290, N286, N263);
and AND2 (N291, N290, N123);
or OR2 (N292, N269, N165);
nor NOR2 (N293, N273, N231);
buf BUF1 (N294, N278);
buf BUF1 (N295, N277);
and AND3 (N296, N287, N2, N192);
xor XOR2 (N297, N282, N243);
not NOT1 (N298, N289);
nand NAND3 (N299, N292, N173, N68);
xor XOR2 (N300, N294, N291);
or OR2 (N301, N242, N294);
not NOT1 (N302, N298);
nor NOR2 (N303, N301, N213);
and AND4 (N304, N279, N33, N220, N215);
xor XOR2 (N305, N296, N163);
not NOT1 (N306, N293);
xor XOR2 (N307, N288, N29);
nand NAND2 (N308, N295, N201);
nand NAND4 (N309, N308, N100, N124, N30);
xor XOR2 (N310, N309, N158);
nand NAND2 (N311, N303, N199);
nand NAND4 (N312, N310, N164, N65, N36);
nand NAND4 (N313, N300, N52, N178, N93);
not NOT1 (N314, N302);
nor NOR2 (N315, N299, N287);
nand NAND4 (N316, N311, N183, N240, N303);
not NOT1 (N317, N315);
or OR3 (N318, N314, N173, N259);
nor NOR4 (N319, N313, N43, N212, N313);
buf BUF1 (N320, N319);
and AND4 (N321, N307, N46, N85, N263);
nor NOR4 (N322, N318, N49, N55, N320);
nand NAND4 (N323, N280, N212, N108, N37);
nand NAND2 (N324, N317, N224);
and AND4 (N325, N304, N205, N295, N278);
buf BUF1 (N326, N312);
or OR3 (N327, N316, N263, N143);
nand NAND3 (N328, N327, N215, N302);
buf BUF1 (N329, N322);
nand NAND2 (N330, N323, N58);
or OR3 (N331, N305, N316, N131);
xor XOR2 (N332, N329, N6);
xor XOR2 (N333, N325, N90);
or OR3 (N334, N332, N195, N102);
nor NOR4 (N335, N331, N303, N319, N74);
nand NAND2 (N336, N326, N54);
nand NAND4 (N337, N297, N155, N19, N129);
and AND3 (N338, N306, N31, N209);
xor XOR2 (N339, N333, N295);
nor NOR3 (N340, N338, N19, N292);
and AND3 (N341, N330, N129, N267);
xor XOR2 (N342, N341, N126);
buf BUF1 (N343, N321);
xor XOR2 (N344, N343, N71);
or OR4 (N345, N342, N23, N143, N62);
nand NAND2 (N346, N335, N246);
nand NAND4 (N347, N345, N62, N295, N180);
xor XOR2 (N348, N324, N300);
xor XOR2 (N349, N334, N114);
xor XOR2 (N350, N339, N58);
xor XOR2 (N351, N346, N121);
nor NOR2 (N352, N337, N284);
and AND3 (N353, N347, N95, N15);
and AND4 (N354, N348, N240, N65, N7);
nand NAND2 (N355, N336, N324);
or OR4 (N356, N352, N123, N293, N133);
or OR2 (N357, N350, N32);
or OR4 (N358, N353, N44, N241, N346);
and AND4 (N359, N355, N208, N304, N83);
or OR2 (N360, N357, N95);
xor XOR2 (N361, N328, N128);
and AND3 (N362, N360, N139, N252);
buf BUF1 (N363, N349);
not NOT1 (N364, N361);
not NOT1 (N365, N363);
not NOT1 (N366, N340);
and AND4 (N367, N358, N207, N137, N186);
not NOT1 (N368, N356);
or OR4 (N369, N368, N32, N71, N2);
nor NOR2 (N370, N369, N51);
not NOT1 (N371, N366);
buf BUF1 (N372, N354);
buf BUF1 (N373, N370);
or OR3 (N374, N364, N89, N66);
or OR2 (N375, N371, N82);
not NOT1 (N376, N344);
and AND3 (N377, N373, N76, N165);
xor XOR2 (N378, N351, N87);
nand NAND2 (N379, N377, N81);
or OR2 (N380, N379, N115);
nand NAND2 (N381, N372, N337);
or OR3 (N382, N375, N129, N299);
not NOT1 (N383, N374);
xor XOR2 (N384, N382, N146);
buf BUF1 (N385, N362);
nor NOR2 (N386, N359, N242);
xor XOR2 (N387, N367, N147);
nor NOR2 (N388, N386, N194);
not NOT1 (N389, N365);
xor XOR2 (N390, N376, N208);
xor XOR2 (N391, N388, N67);
nand NAND3 (N392, N380, N316, N361);
or OR4 (N393, N384, N383, N50, N175);
nand NAND4 (N394, N195, N279, N25, N16);
or OR3 (N395, N392, N4, N254);
nand NAND4 (N396, N385, N10, N215, N230);
or OR3 (N397, N396, N123, N354);
nor NOR3 (N398, N395, N66, N322);
buf BUF1 (N399, N397);
xor XOR2 (N400, N393, N289);
xor XOR2 (N401, N378, N180);
buf BUF1 (N402, N390);
buf BUF1 (N403, N402);
nor NOR3 (N404, N400, N132, N146);
nor NOR4 (N405, N391, N59, N315, N357);
xor XOR2 (N406, N394, N286);
xor XOR2 (N407, N404, N208);
or OR2 (N408, N399, N121);
not NOT1 (N409, N398);
buf BUF1 (N410, N389);
or OR4 (N411, N408, N211, N174, N293);
not NOT1 (N412, N401);
xor XOR2 (N413, N387, N316);
or OR3 (N414, N407, N96, N122);
nand NAND2 (N415, N409, N304);
and AND3 (N416, N403, N91, N116);
nor NOR3 (N417, N416, N270, N270);
or OR3 (N418, N412, N189, N258);
or OR4 (N419, N411, N46, N194, N267);
buf BUF1 (N420, N417);
or OR4 (N421, N405, N67, N273, N38);
not NOT1 (N422, N419);
nor NOR3 (N423, N413, N283, N147);
buf BUF1 (N424, N418);
not NOT1 (N425, N414);
buf BUF1 (N426, N406);
buf BUF1 (N427, N415);
nand NAND2 (N428, N425, N171);
nand NAND4 (N429, N424, N285, N76, N238);
or OR4 (N430, N421, N198, N317, N114);
or OR4 (N431, N430, N151, N99, N53);
not NOT1 (N432, N420);
or OR4 (N433, N427, N144, N142, N120);
and AND3 (N434, N432, N100, N60);
xor XOR2 (N435, N428, N153);
nand NAND4 (N436, N410, N113, N254, N377);
buf BUF1 (N437, N431);
xor XOR2 (N438, N434, N338);
buf BUF1 (N439, N422);
or OR2 (N440, N429, N158);
xor XOR2 (N441, N433, N433);
buf BUF1 (N442, N437);
or OR4 (N443, N423, N415, N266, N347);
not NOT1 (N444, N440);
xor XOR2 (N445, N444, N354);
buf BUF1 (N446, N441);
and AND2 (N447, N438, N95);
or OR2 (N448, N442, N241);
not NOT1 (N449, N447);
not NOT1 (N450, N436);
and AND3 (N451, N443, N100, N48);
xor XOR2 (N452, N450, N287);
nor NOR4 (N453, N435, N157, N203, N230);
nand NAND4 (N454, N452, N65, N145, N170);
nand NAND4 (N455, N439, N279, N188, N340);
nand NAND4 (N456, N381, N201, N277, N387);
nor NOR3 (N457, N445, N271, N14);
nor NOR2 (N458, N451, N262);
xor XOR2 (N459, N446, N88);
buf BUF1 (N460, N448);
nor NOR3 (N461, N449, N99, N13);
buf BUF1 (N462, N456);
nor NOR4 (N463, N459, N196, N400, N288);
or OR3 (N464, N426, N52, N274);
nand NAND2 (N465, N463, N276);
not NOT1 (N466, N453);
xor XOR2 (N467, N465, N206);
not NOT1 (N468, N464);
buf BUF1 (N469, N468);
buf BUF1 (N470, N466);
and AND3 (N471, N461, N334, N279);
xor XOR2 (N472, N460, N469);
nor NOR4 (N473, N259, N98, N79, N240);
or OR4 (N474, N462, N317, N140, N221);
or OR4 (N475, N471, N185, N219, N295);
or OR3 (N476, N455, N156, N172);
nor NOR2 (N477, N475, N26);
xor XOR2 (N478, N474, N474);
nor NOR2 (N479, N458, N63);
nor NOR2 (N480, N478, N6);
xor XOR2 (N481, N457, N74);
nor NOR3 (N482, N473, N6, N241);
and AND3 (N483, N454, N147, N428);
xor XOR2 (N484, N470, N146);
nor NOR4 (N485, N481, N37, N246, N272);
and AND4 (N486, N472, N331, N404, N376);
buf BUF1 (N487, N477);
or OR3 (N488, N476, N232, N187);
and AND4 (N489, N485, N211, N375, N226);
buf BUF1 (N490, N479);
buf BUF1 (N491, N489);
nand NAND3 (N492, N467, N302, N201);
or OR4 (N493, N480, N322, N443, N187);
buf BUF1 (N494, N492);
xor XOR2 (N495, N483, N218);
or OR3 (N496, N490, N293, N271);
xor XOR2 (N497, N496, N442);
buf BUF1 (N498, N484);
xor XOR2 (N499, N493, N210);
xor XOR2 (N500, N491, N152);
nand NAND2 (N501, N497, N477);
buf BUF1 (N502, N499);
and AND4 (N503, N488, N388, N233, N305);
xor XOR2 (N504, N482, N150);
and AND4 (N505, N495, N280, N193, N162);
nor NOR2 (N506, N494, N491);
buf BUF1 (N507, N498);
xor XOR2 (N508, N504, N223);
or OR2 (N509, N501, N20);
or OR2 (N510, N487, N215);
xor XOR2 (N511, N509, N364);
nand NAND2 (N512, N502, N150);
buf BUF1 (N513, N507);
nand NAND3 (N514, N508, N313, N212);
xor XOR2 (N515, N511, N360);
xor XOR2 (N516, N510, N119);
not NOT1 (N517, N513);
buf BUF1 (N518, N500);
or OR4 (N519, N517, N307, N32, N281);
buf BUF1 (N520, N516);
or OR4 (N521, N503, N362, N45, N44);
nor NOR2 (N522, N512, N25);
or OR3 (N523, N486, N72, N286);
nor NOR2 (N524, N505, N52);
nor NOR2 (N525, N518, N95);
xor XOR2 (N526, N514, N506);
nor NOR4 (N527, N512, N190, N324, N358);
not NOT1 (N528, N527);
xor XOR2 (N529, N522, N17);
buf BUF1 (N530, N524);
nand NAND4 (N531, N528, N385, N432, N480);
not NOT1 (N532, N530);
and AND3 (N533, N526, N510, N441);
nor NOR4 (N534, N521, N199, N493, N354);
nor NOR4 (N535, N533, N54, N457, N290);
and AND2 (N536, N519, N511);
nor NOR2 (N537, N536, N529);
nor NOR3 (N538, N514, N31, N476);
xor XOR2 (N539, N534, N389);
or OR4 (N540, N520, N357, N234, N486);
not NOT1 (N541, N538);
nand NAND2 (N542, N525, N242);
nor NOR2 (N543, N531, N445);
not NOT1 (N544, N543);
xor XOR2 (N545, N535, N291);
and AND3 (N546, N515, N543, N472);
nand NAND2 (N547, N537, N57);
not NOT1 (N548, N542);
nand NAND2 (N549, N541, N454);
not NOT1 (N550, N544);
xor XOR2 (N551, N546, N231);
and AND4 (N552, N532, N465, N396, N143);
buf BUF1 (N553, N523);
xor XOR2 (N554, N550, N24);
nand NAND3 (N555, N539, N14, N299);
nand NAND3 (N556, N549, N384, N394);
xor XOR2 (N557, N540, N531);
or OR3 (N558, N551, N487, N392);
xor XOR2 (N559, N554, N489);
buf BUF1 (N560, N553);
nor NOR4 (N561, N557, N523, N21, N465);
xor XOR2 (N562, N547, N226);
not NOT1 (N563, N561);
buf BUF1 (N564, N556);
xor XOR2 (N565, N548, N247);
or OR4 (N566, N565, N74, N380, N409);
xor XOR2 (N567, N558, N149);
not NOT1 (N568, N564);
nor NOR2 (N569, N567, N156);
buf BUF1 (N570, N568);
nor NOR3 (N571, N555, N94, N539);
buf BUF1 (N572, N570);
nor NOR4 (N573, N552, N394, N122, N7);
buf BUF1 (N574, N545);
and AND2 (N575, N562, N314);
nor NOR3 (N576, N563, N155, N484);
and AND2 (N577, N576, N39);
not NOT1 (N578, N572);
or OR3 (N579, N571, N32, N380);
and AND4 (N580, N575, N239, N201, N529);
buf BUF1 (N581, N569);
not NOT1 (N582, N581);
or OR3 (N583, N580, N513, N2);
nand NAND2 (N584, N573, N508);
buf BUF1 (N585, N582);
or OR2 (N586, N585, N423);
xor XOR2 (N587, N583, N125);
nor NOR4 (N588, N566, N96, N225, N533);
and AND2 (N589, N578, N465);
buf BUF1 (N590, N589);
buf BUF1 (N591, N588);
nor NOR3 (N592, N587, N440, N375);
and AND3 (N593, N590, N547, N381);
nor NOR3 (N594, N559, N132, N144);
and AND4 (N595, N591, N214, N151, N465);
nand NAND2 (N596, N577, N554);
nor NOR3 (N597, N560, N435, N391);
nor NOR4 (N598, N594, N459, N549, N223);
or OR3 (N599, N598, N380, N391);
not NOT1 (N600, N596);
or OR3 (N601, N584, N134, N507);
xor XOR2 (N602, N593, N528);
buf BUF1 (N603, N574);
nor NOR4 (N604, N586, N528, N207, N163);
nor NOR3 (N605, N600, N15, N28);
nand NAND2 (N606, N601, N78);
not NOT1 (N607, N606);
nor NOR4 (N608, N597, N552, N285, N591);
buf BUF1 (N609, N603);
buf BUF1 (N610, N579);
and AND3 (N611, N609, N458, N232);
xor XOR2 (N612, N595, N209);
and AND2 (N613, N610, N3);
not NOT1 (N614, N608);
or OR4 (N615, N604, N569, N275, N485);
nand NAND2 (N616, N607, N465);
nand NAND2 (N617, N592, N44);
buf BUF1 (N618, N613);
nor NOR3 (N619, N617, N88, N280);
xor XOR2 (N620, N612, N227);
or OR3 (N621, N618, N501, N434);
buf BUF1 (N622, N615);
not NOT1 (N623, N620);
xor XOR2 (N624, N602, N87);
and AND2 (N625, N605, N343);
buf BUF1 (N626, N621);
or OR4 (N627, N624, N130, N323, N610);
nor NOR4 (N628, N627, N3, N43, N73);
xor XOR2 (N629, N622, N420);
buf BUF1 (N630, N628);
xor XOR2 (N631, N611, N33);
buf BUF1 (N632, N623);
nor NOR4 (N633, N625, N584, N617, N533);
xor XOR2 (N634, N619, N349);
nor NOR3 (N635, N616, N630, N385);
xor XOR2 (N636, N504, N141);
not NOT1 (N637, N626);
not NOT1 (N638, N629);
nor NOR3 (N639, N614, N257, N30);
or OR3 (N640, N631, N66, N592);
or OR4 (N641, N638, N85, N534, N600);
nor NOR3 (N642, N632, N428, N576);
nand NAND4 (N643, N634, N565, N164, N158);
xor XOR2 (N644, N642, N140);
and AND3 (N645, N641, N18, N310);
xor XOR2 (N646, N643, N364);
nor NOR4 (N647, N637, N363, N377, N472);
xor XOR2 (N648, N635, N207);
xor XOR2 (N649, N647, N97);
and AND4 (N650, N636, N97, N91, N422);
and AND4 (N651, N648, N619, N612, N627);
buf BUF1 (N652, N650);
nor NOR3 (N653, N640, N84, N169);
and AND3 (N654, N599, N94, N216);
not NOT1 (N655, N649);
and AND4 (N656, N639, N298, N204, N326);
nor NOR2 (N657, N653, N85);
nand NAND3 (N658, N655, N224, N29);
and AND4 (N659, N633, N382, N319, N64);
buf BUF1 (N660, N659);
buf BUF1 (N661, N652);
not NOT1 (N662, N658);
xor XOR2 (N663, N651, N170);
and AND2 (N664, N645, N637);
and AND3 (N665, N646, N632, N382);
and AND3 (N666, N665, N602, N525);
or OR3 (N667, N660, N453, N343);
nand NAND3 (N668, N664, N139, N398);
not NOT1 (N669, N657);
xor XOR2 (N670, N662, N203);
xor XOR2 (N671, N644, N521);
nor NOR4 (N672, N663, N195, N125, N432);
nand NAND2 (N673, N668, N170);
nor NOR3 (N674, N656, N442, N520);
not NOT1 (N675, N672);
or OR3 (N676, N671, N603, N500);
not NOT1 (N677, N669);
nand NAND2 (N678, N674, N368);
or OR3 (N679, N678, N361, N94);
not NOT1 (N680, N661);
or OR4 (N681, N654, N403, N89, N544);
xor XOR2 (N682, N676, N658);
not NOT1 (N683, N682);
nand NAND3 (N684, N673, N61, N19);
not NOT1 (N685, N675);
buf BUF1 (N686, N667);
nor NOR3 (N687, N686, N212, N471);
not NOT1 (N688, N666);
not NOT1 (N689, N683);
xor XOR2 (N690, N670, N393);
buf BUF1 (N691, N687);
or OR3 (N692, N677, N491, N34);
buf BUF1 (N693, N680);
not NOT1 (N694, N679);
not NOT1 (N695, N688);
not NOT1 (N696, N684);
not NOT1 (N697, N694);
and AND4 (N698, N695, N253, N576, N654);
buf BUF1 (N699, N681);
nand NAND4 (N700, N689, N423, N322, N666);
not NOT1 (N701, N692);
not NOT1 (N702, N691);
not NOT1 (N703, N701);
not NOT1 (N704, N696);
xor XOR2 (N705, N700, N168);
nand NAND4 (N706, N699, N150, N544, N565);
or OR3 (N707, N685, N303, N623);
and AND4 (N708, N690, N37, N662, N549);
xor XOR2 (N709, N697, N338);
not NOT1 (N710, N698);
xor XOR2 (N711, N703, N54);
xor XOR2 (N712, N711, N564);
buf BUF1 (N713, N704);
xor XOR2 (N714, N707, N192);
nor NOR2 (N715, N706, N711);
nor NOR3 (N716, N710, N226, N141);
nand NAND2 (N717, N693, N669);
and AND2 (N718, N713, N251);
and AND2 (N719, N705, N255);
buf BUF1 (N720, N712);
and AND2 (N721, N716, N576);
nor NOR2 (N722, N721, N186);
nor NOR3 (N723, N715, N678, N234);
not NOT1 (N724, N720);
or OR2 (N725, N724, N595);
and AND4 (N726, N708, N172, N206, N679);
not NOT1 (N727, N726);
buf BUF1 (N728, N723);
xor XOR2 (N729, N718, N484);
buf BUF1 (N730, N725);
not NOT1 (N731, N717);
and AND4 (N732, N722, N59, N140, N173);
not NOT1 (N733, N729);
not NOT1 (N734, N732);
buf BUF1 (N735, N730);
not NOT1 (N736, N733);
xor XOR2 (N737, N736, N251);
or OR4 (N738, N709, N443, N683, N319);
not NOT1 (N739, N702);
or OR2 (N740, N734, N182);
or OR2 (N741, N731, N242);
xor XOR2 (N742, N737, N257);
and AND2 (N743, N739, N690);
buf BUF1 (N744, N743);
nand NAND2 (N745, N735, N73);
not NOT1 (N746, N740);
buf BUF1 (N747, N741);
xor XOR2 (N748, N742, N690);
nor NOR4 (N749, N746, N632, N526, N258);
nand NAND2 (N750, N745, N198);
buf BUF1 (N751, N750);
or OR3 (N752, N744, N370, N286);
not NOT1 (N753, N751);
not NOT1 (N754, N719);
nor NOR2 (N755, N752, N696);
or OR2 (N756, N755, N665);
buf BUF1 (N757, N738);
not NOT1 (N758, N714);
not NOT1 (N759, N758);
nand NAND3 (N760, N756, N602, N513);
not NOT1 (N761, N760);
and AND4 (N762, N727, N761, N732, N143);
xor XOR2 (N763, N731, N608);
xor XOR2 (N764, N762, N560);
and AND3 (N765, N753, N30, N547);
not NOT1 (N766, N757);
not NOT1 (N767, N765);
not NOT1 (N768, N749);
not NOT1 (N769, N767);
nand NAND2 (N770, N769, N92);
buf BUF1 (N771, N747);
nand NAND3 (N772, N766, N120, N226);
or OR3 (N773, N772, N461, N97);
xor XOR2 (N774, N771, N648);
not NOT1 (N775, N728);
nor NOR2 (N776, N754, N342);
nor NOR2 (N777, N763, N441);
not NOT1 (N778, N775);
or OR3 (N779, N748, N627, N560);
nand NAND2 (N780, N774, N43);
nor NOR4 (N781, N780, N117, N453, N382);
not NOT1 (N782, N773);
nor NOR4 (N783, N779, N167, N518, N45);
nand NAND4 (N784, N764, N143, N92, N191);
xor XOR2 (N785, N778, N527);
nand NAND3 (N786, N781, N740, N276);
nor NOR4 (N787, N782, N676, N694, N73);
nor NOR4 (N788, N785, N157, N484, N40);
nor NOR2 (N789, N768, N465);
or OR3 (N790, N789, N717, N98);
and AND2 (N791, N788, N367);
and AND3 (N792, N759, N635, N239);
buf BUF1 (N793, N786);
xor XOR2 (N794, N793, N170);
and AND2 (N795, N783, N575);
and AND4 (N796, N795, N639, N180, N778);
not NOT1 (N797, N784);
nand NAND2 (N798, N797, N581);
xor XOR2 (N799, N777, N445);
buf BUF1 (N800, N776);
and AND2 (N801, N796, N251);
and AND2 (N802, N770, N237);
or OR3 (N803, N799, N672, N131);
buf BUF1 (N804, N787);
not NOT1 (N805, N804);
or OR2 (N806, N791, N400);
buf BUF1 (N807, N798);
buf BUF1 (N808, N803);
buf BUF1 (N809, N806);
and AND2 (N810, N790, N441);
nor NOR2 (N811, N802, N15);
nand NAND2 (N812, N805, N589);
xor XOR2 (N813, N809, N650);
nor NOR2 (N814, N811, N431);
nand NAND2 (N815, N808, N775);
nand NAND4 (N816, N800, N485, N578, N77);
xor XOR2 (N817, N794, N743);
or OR2 (N818, N815, N178);
and AND3 (N819, N810, N392, N505);
or OR3 (N820, N818, N508, N255);
not NOT1 (N821, N813);
nand NAND2 (N822, N801, N632);
not NOT1 (N823, N819);
nand NAND3 (N824, N807, N431, N441);
nand NAND2 (N825, N820, N134);
nor NOR3 (N826, N812, N726, N480);
and AND2 (N827, N822, N539);
buf BUF1 (N828, N823);
not NOT1 (N829, N821);
xor XOR2 (N830, N825, N114);
buf BUF1 (N831, N829);
or OR3 (N832, N792, N823, N792);
nor NOR2 (N833, N824, N806);
nor NOR3 (N834, N831, N143, N691);
buf BUF1 (N835, N832);
xor XOR2 (N836, N827, N162);
not NOT1 (N837, N834);
not NOT1 (N838, N814);
and AND2 (N839, N838, N388);
xor XOR2 (N840, N837, N687);
not NOT1 (N841, N836);
or OR4 (N842, N833, N144, N839, N322);
and AND3 (N843, N499, N48, N226);
nand NAND4 (N844, N840, N267, N115, N219);
nor NOR3 (N845, N844, N801, N304);
buf BUF1 (N846, N828);
nor NOR4 (N847, N835, N367, N728, N723);
not NOT1 (N848, N830);
nor NOR2 (N849, N846, N573);
not NOT1 (N850, N848);
buf BUF1 (N851, N845);
xor XOR2 (N852, N841, N483);
buf BUF1 (N853, N817);
nor NOR4 (N854, N816, N771, N393, N513);
not NOT1 (N855, N853);
buf BUF1 (N856, N854);
nor NOR4 (N857, N855, N655, N427, N63);
or OR4 (N858, N850, N467, N186, N857);
nor NOR4 (N859, N114, N514, N700, N144);
nor NOR3 (N860, N849, N85, N348);
and AND4 (N861, N859, N579, N533, N533);
and AND3 (N862, N826, N93, N227);
xor XOR2 (N863, N842, N456);
buf BUF1 (N864, N856);
not NOT1 (N865, N847);
or OR4 (N866, N858, N242, N710, N605);
buf BUF1 (N867, N843);
xor XOR2 (N868, N862, N168);
not NOT1 (N869, N863);
nor NOR3 (N870, N851, N554, N103);
and AND3 (N871, N864, N739, N648);
not NOT1 (N872, N869);
or OR4 (N873, N860, N356, N350, N158);
buf BUF1 (N874, N871);
nand NAND3 (N875, N865, N361, N453);
buf BUF1 (N876, N852);
nor NOR3 (N877, N870, N863, N315);
nand NAND3 (N878, N868, N483, N810);
nand NAND2 (N879, N874, N674);
and AND2 (N880, N867, N696);
and AND2 (N881, N861, N251);
nor NOR4 (N882, N872, N313, N276, N566);
xor XOR2 (N883, N875, N372);
not NOT1 (N884, N866);
not NOT1 (N885, N880);
not NOT1 (N886, N877);
and AND2 (N887, N878, N245);
or OR3 (N888, N884, N13, N720);
buf BUF1 (N889, N876);
buf BUF1 (N890, N881);
nand NAND2 (N891, N883, N417);
and AND2 (N892, N873, N597);
nor NOR3 (N893, N885, N237, N148);
nand NAND4 (N894, N891, N520, N557, N648);
xor XOR2 (N895, N890, N571);
not NOT1 (N896, N879);
xor XOR2 (N897, N896, N60);
nand NAND2 (N898, N892, N297);
or OR3 (N899, N898, N158, N665);
nand NAND3 (N900, N887, N556, N511);
or OR3 (N901, N899, N592, N547);
xor XOR2 (N902, N893, N354);
nand NAND4 (N903, N897, N204, N873, N70);
not NOT1 (N904, N894);
buf BUF1 (N905, N900);
and AND3 (N906, N904, N337, N313);
nand NAND2 (N907, N902, N597);
nand NAND3 (N908, N882, N528, N10);
or OR4 (N909, N895, N449, N467, N107);
not NOT1 (N910, N905);
nand NAND3 (N911, N901, N29, N353);
nor NOR2 (N912, N909, N697);
and AND4 (N913, N903, N34, N526, N880);
nor NOR3 (N914, N910, N716, N261);
not NOT1 (N915, N913);
buf BUF1 (N916, N906);
not NOT1 (N917, N914);
buf BUF1 (N918, N912);
nand NAND4 (N919, N917, N149, N540, N268);
or OR4 (N920, N918, N572, N90, N121);
buf BUF1 (N921, N911);
nand NAND4 (N922, N907, N533, N310, N608);
xor XOR2 (N923, N889, N419);
xor XOR2 (N924, N923, N793);
or OR3 (N925, N924, N521, N208);
nor NOR3 (N926, N916, N514, N433);
or OR2 (N927, N886, N687);
or OR2 (N928, N915, N641);
buf BUF1 (N929, N920);
nor NOR2 (N930, N888, N800);
or OR3 (N931, N921, N163, N604);
or OR2 (N932, N908, N113);
xor XOR2 (N933, N928, N754);
or OR2 (N934, N919, N695);
not NOT1 (N935, N934);
buf BUF1 (N936, N932);
not NOT1 (N937, N931);
nor NOR2 (N938, N935, N912);
nor NOR2 (N939, N925, N696);
nand NAND3 (N940, N929, N129, N111);
nand NAND2 (N941, N939, N390);
nand NAND3 (N942, N941, N704, N100);
and AND4 (N943, N926, N857, N539, N118);
not NOT1 (N944, N936);
or OR2 (N945, N938, N773);
buf BUF1 (N946, N922);
not NOT1 (N947, N946);
xor XOR2 (N948, N945, N342);
not NOT1 (N949, N943);
or OR4 (N950, N942, N513, N946, N935);
nand NAND2 (N951, N950, N22);
buf BUF1 (N952, N947);
nand NAND3 (N953, N933, N521, N181);
buf BUF1 (N954, N948);
xor XOR2 (N955, N927, N248);
and AND2 (N956, N951, N515);
nand NAND4 (N957, N955, N379, N500, N590);
nor NOR3 (N958, N954, N473, N498);
buf BUF1 (N959, N953);
not NOT1 (N960, N930);
xor XOR2 (N961, N944, N325);
xor XOR2 (N962, N937, N511);
and AND3 (N963, N957, N430, N820);
xor XOR2 (N964, N963, N673);
or OR3 (N965, N958, N879, N933);
xor XOR2 (N966, N961, N203);
nor NOR2 (N967, N965, N150);
nand NAND3 (N968, N940, N522, N350);
nor NOR4 (N969, N966, N828, N948, N819);
nor NOR2 (N970, N967, N601);
not NOT1 (N971, N964);
or OR4 (N972, N952, N164, N836, N361);
xor XOR2 (N973, N969, N619);
and AND2 (N974, N972, N69);
nor NOR4 (N975, N959, N579, N845, N402);
nor NOR3 (N976, N949, N379, N506);
not NOT1 (N977, N960);
xor XOR2 (N978, N975, N164);
buf BUF1 (N979, N977);
nand NAND2 (N980, N973, N501);
xor XOR2 (N981, N974, N156);
nor NOR2 (N982, N976, N403);
xor XOR2 (N983, N978, N767);
xor XOR2 (N984, N983, N471);
xor XOR2 (N985, N971, N975);
nand NAND4 (N986, N962, N756, N875, N874);
nand NAND3 (N987, N984, N407, N483);
or OR3 (N988, N968, N40, N837);
and AND4 (N989, N985, N547, N316, N516);
nor NOR3 (N990, N987, N93, N541);
nand NAND2 (N991, N981, N492);
nor NOR2 (N992, N970, N434);
nor NOR2 (N993, N989, N544);
nor NOR3 (N994, N980, N189, N738);
nor NOR4 (N995, N993, N298, N573, N635);
buf BUF1 (N996, N979);
and AND4 (N997, N991, N454, N608, N421);
xor XOR2 (N998, N995, N762);
xor XOR2 (N999, N994, N44);
buf BUF1 (N1000, N998);
or OR3 (N1001, N997, N78, N749);
nand NAND4 (N1002, N990, N589, N448, N829);
not NOT1 (N1003, N982);
and AND4 (N1004, N1002, N273, N270, N606);
or OR2 (N1005, N956, N609);
not NOT1 (N1006, N1004);
xor XOR2 (N1007, N999, N368);
not NOT1 (N1008, N996);
nand NAND4 (N1009, N1001, N635, N786, N697);
nand NAND2 (N1010, N1003, N559);
xor XOR2 (N1011, N992, N705);
not NOT1 (N1012, N1007);
nor NOR2 (N1013, N1010, N400);
and AND2 (N1014, N1011, N992);
and AND4 (N1015, N1014, N408, N864, N870);
nor NOR4 (N1016, N1015, N370, N845, N44);
nand NAND3 (N1017, N1006, N120, N95);
buf BUF1 (N1018, N1005);
nand NAND2 (N1019, N988, N565);
buf BUF1 (N1020, N1009);
xor XOR2 (N1021, N1008, N176);
nor NOR2 (N1022, N1021, N153);
and AND4 (N1023, N1017, N576, N72, N133);
not NOT1 (N1024, N1019);
nand NAND3 (N1025, N1024, N684, N157);
not NOT1 (N1026, N986);
or OR2 (N1027, N1026, N193);
nor NOR4 (N1028, N1000, N32, N712, N691);
or OR2 (N1029, N1012, N593);
not NOT1 (N1030, N1022);
and AND3 (N1031, N1018, N390, N478);
or OR3 (N1032, N1025, N1000, N580);
or OR3 (N1033, N1028, N819, N96);
nor NOR4 (N1034, N1030, N580, N798, N566);
buf BUF1 (N1035, N1016);
xor XOR2 (N1036, N1013, N114);
not NOT1 (N1037, N1036);
and AND2 (N1038, N1032, N398);
nor NOR4 (N1039, N1023, N857, N330, N120);
or OR4 (N1040, N1034, N628, N359, N298);
nor NOR4 (N1041, N1039, N220, N169, N18);
not NOT1 (N1042, N1041);
nor NOR4 (N1043, N1020, N215, N824, N48);
nor NOR3 (N1044, N1029, N763, N306);
and AND3 (N1045, N1043, N599, N1009);
not NOT1 (N1046, N1027);
or OR2 (N1047, N1037, N528);
buf BUF1 (N1048, N1040);
and AND4 (N1049, N1047, N983, N22, N807);
nor NOR4 (N1050, N1033, N386, N401, N322);
nand NAND3 (N1051, N1046, N992, N960);
xor XOR2 (N1052, N1044, N304);
nor NOR2 (N1053, N1042, N297);
xor XOR2 (N1054, N1045, N693);
not NOT1 (N1055, N1050);
buf BUF1 (N1056, N1031);
nor NOR2 (N1057, N1055, N752);
not NOT1 (N1058, N1052);
nand NAND3 (N1059, N1049, N230, N29);
xor XOR2 (N1060, N1053, N189);
and AND4 (N1061, N1057, N452, N925, N803);
xor XOR2 (N1062, N1059, N953);
xor XOR2 (N1063, N1060, N160);
buf BUF1 (N1064, N1062);
and AND3 (N1065, N1054, N1033, N656);
or OR4 (N1066, N1048, N66, N359, N643);
or OR3 (N1067, N1064, N949, N466);
buf BUF1 (N1068, N1061);
and AND3 (N1069, N1038, N41, N209);
not NOT1 (N1070, N1066);
xor XOR2 (N1071, N1065, N903);
or OR3 (N1072, N1056, N827, N738);
not NOT1 (N1073, N1035);
nor NOR3 (N1074, N1068, N642, N581);
or OR3 (N1075, N1074, N10, N1020);
or OR2 (N1076, N1073, N301);
and AND3 (N1077, N1058, N882, N825);
buf BUF1 (N1078, N1077);
xor XOR2 (N1079, N1071, N821);
and AND2 (N1080, N1075, N956);
nand NAND2 (N1081, N1072, N352);
nor NOR4 (N1082, N1076, N125, N317, N32);
xor XOR2 (N1083, N1082, N710);
buf BUF1 (N1084, N1080);
or OR2 (N1085, N1067, N553);
not NOT1 (N1086, N1083);
nand NAND4 (N1087, N1081, N788, N944, N179);
nor NOR3 (N1088, N1070, N112, N881);
and AND2 (N1089, N1087, N500);
nand NAND4 (N1090, N1051, N1048, N28, N16);
or OR3 (N1091, N1084, N267, N118);
or OR3 (N1092, N1091, N586, N760);
and AND2 (N1093, N1079, N96);
buf BUF1 (N1094, N1090);
or OR2 (N1095, N1092, N686);
not NOT1 (N1096, N1094);
xor XOR2 (N1097, N1086, N1064);
and AND3 (N1098, N1096, N376, N650);
and AND2 (N1099, N1095, N284);
buf BUF1 (N1100, N1089);
buf BUF1 (N1101, N1088);
nor NOR3 (N1102, N1093, N855, N605);
not NOT1 (N1103, N1063);
and AND2 (N1104, N1078, N885);
nor NOR3 (N1105, N1104, N749, N106);
or OR4 (N1106, N1098, N652, N182, N763);
not NOT1 (N1107, N1101);
buf BUF1 (N1108, N1102);
buf BUF1 (N1109, N1100);
or OR3 (N1110, N1099, N153, N601);
nand NAND4 (N1111, N1109, N881, N349, N501);
buf BUF1 (N1112, N1097);
xor XOR2 (N1113, N1069, N763);
xor XOR2 (N1114, N1085, N357);
buf BUF1 (N1115, N1106);
and AND2 (N1116, N1103, N722);
and AND4 (N1117, N1105, N954, N879, N243);
nand NAND3 (N1118, N1117, N97, N777);
nand NAND2 (N1119, N1107, N180);
nand NAND2 (N1120, N1119, N621);
and AND3 (N1121, N1116, N303, N429);
and AND2 (N1122, N1110, N824);
xor XOR2 (N1123, N1120, N963);
not NOT1 (N1124, N1123);
xor XOR2 (N1125, N1108, N33);
xor XOR2 (N1126, N1124, N952);
nor NOR2 (N1127, N1125, N591);
and AND3 (N1128, N1115, N306, N545);
not NOT1 (N1129, N1121);
and AND3 (N1130, N1111, N319, N1074);
buf BUF1 (N1131, N1129);
nand NAND2 (N1132, N1118, N683);
and AND2 (N1133, N1112, N589);
nor NOR4 (N1134, N1131, N400, N604, N1043);
buf BUF1 (N1135, N1127);
or OR4 (N1136, N1135, N538, N1062, N490);
and AND2 (N1137, N1133, N279);
nand NAND4 (N1138, N1126, N768, N243, N873);
buf BUF1 (N1139, N1122);
not NOT1 (N1140, N1134);
nor NOR2 (N1141, N1140, N1081);
nand NAND2 (N1142, N1114, N32);
nor NOR2 (N1143, N1142, N1101);
not NOT1 (N1144, N1139);
not NOT1 (N1145, N1144);
nand NAND3 (N1146, N1128, N911, N206);
xor XOR2 (N1147, N1132, N241);
buf BUF1 (N1148, N1145);
buf BUF1 (N1149, N1141);
nand NAND4 (N1150, N1146, N270, N1039, N230);
xor XOR2 (N1151, N1113, N529);
nand NAND2 (N1152, N1147, N88);
buf BUF1 (N1153, N1137);
not NOT1 (N1154, N1136);
or OR2 (N1155, N1152, N822);
nor NOR4 (N1156, N1153, N855, N841, N442);
not NOT1 (N1157, N1148);
and AND3 (N1158, N1150, N997, N216);
buf BUF1 (N1159, N1130);
nor NOR4 (N1160, N1143, N714, N124, N103);
not NOT1 (N1161, N1155);
nor NOR3 (N1162, N1156, N655, N785);
not NOT1 (N1163, N1154);
nor NOR2 (N1164, N1151, N211);
and AND2 (N1165, N1161, N432);
xor XOR2 (N1166, N1159, N200);
nand NAND2 (N1167, N1158, N965);
or OR2 (N1168, N1167, N307);
and AND2 (N1169, N1138, N664);
nor NOR3 (N1170, N1166, N365, N1045);
nor NOR2 (N1171, N1165, N1158);
or OR4 (N1172, N1169, N231, N203, N444);
and AND3 (N1173, N1162, N555, N659);
xor XOR2 (N1174, N1171, N957);
xor XOR2 (N1175, N1172, N560);
not NOT1 (N1176, N1157);
or OR4 (N1177, N1173, N326, N779, N715);
buf BUF1 (N1178, N1160);
nor NOR3 (N1179, N1149, N363, N815);
xor XOR2 (N1180, N1175, N542);
buf BUF1 (N1181, N1176);
buf BUF1 (N1182, N1179);
nand NAND4 (N1183, N1180, N295, N549, N553);
buf BUF1 (N1184, N1182);
nor NOR4 (N1185, N1170, N846, N913, N526);
buf BUF1 (N1186, N1174);
not NOT1 (N1187, N1177);
or OR3 (N1188, N1186, N155, N522);
and AND3 (N1189, N1168, N684, N1032);
xor XOR2 (N1190, N1164, N194);
nor NOR3 (N1191, N1184, N506, N892);
xor XOR2 (N1192, N1183, N286);
or OR3 (N1193, N1181, N898, N214);
and AND2 (N1194, N1193, N734);
or OR3 (N1195, N1191, N549, N853);
xor XOR2 (N1196, N1195, N247);
or OR2 (N1197, N1163, N804);
nand NAND4 (N1198, N1188, N1058, N238, N542);
nor NOR3 (N1199, N1189, N327, N1103);
or OR2 (N1200, N1187, N475);
or OR4 (N1201, N1194, N5, N382, N244);
nor NOR2 (N1202, N1201, N511);
or OR3 (N1203, N1178, N537, N130);
and AND4 (N1204, N1203, N312, N883, N176);
and AND3 (N1205, N1197, N671, N1033);
not NOT1 (N1206, N1205);
buf BUF1 (N1207, N1202);
not NOT1 (N1208, N1199);
buf BUF1 (N1209, N1208);
xor XOR2 (N1210, N1206, N854);
xor XOR2 (N1211, N1185, N134);
xor XOR2 (N1212, N1207, N871);
and AND3 (N1213, N1190, N1153, N1210);
not NOT1 (N1214, N451);
nand NAND3 (N1215, N1200, N25, N735);
nand NAND4 (N1216, N1192, N745, N328, N242);
and AND2 (N1217, N1209, N939);
xor XOR2 (N1218, N1198, N1189);
not NOT1 (N1219, N1196);
xor XOR2 (N1220, N1214, N312);
xor XOR2 (N1221, N1217, N328);
nor NOR3 (N1222, N1216, N517, N949);
and AND4 (N1223, N1212, N775, N264, N347);
nor NOR2 (N1224, N1211, N353);
not NOT1 (N1225, N1222);
nand NAND2 (N1226, N1221, N222);
or OR3 (N1227, N1225, N693, N262);
nand NAND2 (N1228, N1223, N482);
and AND2 (N1229, N1215, N931);
not NOT1 (N1230, N1213);
not NOT1 (N1231, N1218);
or OR2 (N1232, N1229, N1049);
xor XOR2 (N1233, N1230, N249);
not NOT1 (N1234, N1233);
not NOT1 (N1235, N1227);
or OR4 (N1236, N1231, N1128, N697, N602);
nor NOR2 (N1237, N1234, N616);
not NOT1 (N1238, N1204);
nand NAND3 (N1239, N1238, N192, N1204);
nand NAND2 (N1240, N1237, N1165);
nor NOR4 (N1241, N1236, N357, N499, N455);
not NOT1 (N1242, N1235);
nand NAND4 (N1243, N1241, N1025, N1135, N851);
and AND3 (N1244, N1228, N725, N169);
not NOT1 (N1245, N1220);
xor XOR2 (N1246, N1224, N136);
xor XOR2 (N1247, N1239, N193);
nand NAND2 (N1248, N1243, N864);
nand NAND4 (N1249, N1232, N601, N621, N1244);
or OR3 (N1250, N283, N1049, N1223);
and AND3 (N1251, N1248, N1045, N739);
nor NOR4 (N1252, N1242, N974, N785, N196);
nand NAND3 (N1253, N1240, N381, N866);
xor XOR2 (N1254, N1246, N192);
or OR3 (N1255, N1253, N952, N739);
buf BUF1 (N1256, N1245);
nor NOR4 (N1257, N1249, N504, N544, N825);
nor NOR3 (N1258, N1254, N756, N848);
xor XOR2 (N1259, N1247, N622);
buf BUF1 (N1260, N1252);
nor NOR3 (N1261, N1257, N561, N893);
nor NOR3 (N1262, N1226, N185, N568);
and AND3 (N1263, N1255, N236, N1240);
and AND4 (N1264, N1251, N304, N1064, N146);
nor NOR3 (N1265, N1219, N16, N1147);
nand NAND2 (N1266, N1265, N137);
buf BUF1 (N1267, N1256);
nand NAND3 (N1268, N1258, N850, N82);
not NOT1 (N1269, N1259);
buf BUF1 (N1270, N1267);
not NOT1 (N1271, N1268);
buf BUF1 (N1272, N1250);
xor XOR2 (N1273, N1262, N890);
or OR3 (N1274, N1271, N719, N546);
and AND2 (N1275, N1260, N455);
not NOT1 (N1276, N1263);
xor XOR2 (N1277, N1269, N151);
and AND3 (N1278, N1272, N115, N119);
nor NOR2 (N1279, N1276, N331);
xor XOR2 (N1280, N1264, N266);
xor XOR2 (N1281, N1279, N780);
not NOT1 (N1282, N1266);
xor XOR2 (N1283, N1273, N1177);
not NOT1 (N1284, N1283);
xor XOR2 (N1285, N1284, N743);
nand NAND4 (N1286, N1282, N20, N909, N505);
xor XOR2 (N1287, N1261, N593);
nand NAND4 (N1288, N1274, N487, N209, N285);
nand NAND4 (N1289, N1277, N314, N1141, N974);
and AND2 (N1290, N1280, N933);
nor NOR2 (N1291, N1288, N287);
nor NOR2 (N1292, N1289, N32);
buf BUF1 (N1293, N1292);
not NOT1 (N1294, N1275);
buf BUF1 (N1295, N1287);
nor NOR3 (N1296, N1295, N973, N919);
nor NOR2 (N1297, N1270, N579);
and AND2 (N1298, N1281, N1010);
buf BUF1 (N1299, N1297);
xor XOR2 (N1300, N1286, N906);
buf BUF1 (N1301, N1290);
or OR2 (N1302, N1301, N20);
not NOT1 (N1303, N1285);
not NOT1 (N1304, N1298);
xor XOR2 (N1305, N1300, N1114);
not NOT1 (N1306, N1291);
buf BUF1 (N1307, N1293);
buf BUF1 (N1308, N1302);
or OR4 (N1309, N1299, N519, N338, N844);
not NOT1 (N1310, N1306);
and AND3 (N1311, N1296, N1181, N9);
or OR3 (N1312, N1307, N304, N449);
xor XOR2 (N1313, N1309, N1085);
or OR2 (N1314, N1304, N943);
nand NAND3 (N1315, N1312, N721, N409);
nand NAND4 (N1316, N1278, N1120, N1237, N150);
nor NOR2 (N1317, N1316, N275);
xor XOR2 (N1318, N1313, N1072);
or OR2 (N1319, N1317, N1238);
buf BUF1 (N1320, N1308);
nor NOR4 (N1321, N1320, N983, N602, N515);
and AND3 (N1322, N1319, N110, N1038);
not NOT1 (N1323, N1294);
or OR4 (N1324, N1322, N750, N935, N246);
not NOT1 (N1325, N1310);
xor XOR2 (N1326, N1305, N342);
buf BUF1 (N1327, N1318);
or OR4 (N1328, N1325, N680, N248, N54);
xor XOR2 (N1329, N1323, N1313);
or OR3 (N1330, N1321, N1116, N541);
not NOT1 (N1331, N1328);
xor XOR2 (N1332, N1327, N568);
nand NAND3 (N1333, N1329, N427, N278);
nand NAND2 (N1334, N1315, N1051);
buf BUF1 (N1335, N1332);
nor NOR3 (N1336, N1311, N733, N96);
and AND3 (N1337, N1331, N389, N66);
nor NOR3 (N1338, N1324, N1134, N1019);
or OR3 (N1339, N1336, N1305, N999);
nand NAND3 (N1340, N1337, N787, N309);
nand NAND3 (N1341, N1340, N1091, N562);
xor XOR2 (N1342, N1338, N437);
xor XOR2 (N1343, N1335, N914);
buf BUF1 (N1344, N1341);
not NOT1 (N1345, N1343);
nand NAND3 (N1346, N1330, N592, N765);
nor NOR2 (N1347, N1339, N97);
buf BUF1 (N1348, N1342);
nor NOR2 (N1349, N1348, N319);
nor NOR3 (N1350, N1345, N758, N146);
not NOT1 (N1351, N1303);
xor XOR2 (N1352, N1347, N1015);
and AND2 (N1353, N1350, N1178);
or OR3 (N1354, N1346, N508, N76);
xor XOR2 (N1355, N1344, N398);
nor NOR3 (N1356, N1352, N1149, N963);
nand NAND2 (N1357, N1353, N517);
nand NAND4 (N1358, N1333, N1353, N764, N364);
or OR2 (N1359, N1326, N638);
xor XOR2 (N1360, N1356, N240);
nand NAND2 (N1361, N1357, N1135);
not NOT1 (N1362, N1355);
buf BUF1 (N1363, N1361);
not NOT1 (N1364, N1363);
not NOT1 (N1365, N1351);
or OR2 (N1366, N1360, N431);
and AND4 (N1367, N1314, N413, N278, N865);
not NOT1 (N1368, N1349);
or OR2 (N1369, N1334, N1181);
and AND2 (N1370, N1364, N439);
not NOT1 (N1371, N1359);
nand NAND2 (N1372, N1358, N1300);
and AND4 (N1373, N1370, N405, N1090, N947);
not NOT1 (N1374, N1373);
and AND3 (N1375, N1366, N952, N148);
buf BUF1 (N1376, N1375);
buf BUF1 (N1377, N1371);
nor NOR4 (N1378, N1369, N164, N388, N65);
xor XOR2 (N1379, N1354, N739);
or OR4 (N1380, N1367, N1019, N32, N379);
xor XOR2 (N1381, N1362, N822);
nand NAND3 (N1382, N1365, N1216, N599);
nand NAND4 (N1383, N1368, N253, N898, N103);
not NOT1 (N1384, N1380);
nor NOR3 (N1385, N1382, N1335, N1055);
xor XOR2 (N1386, N1378, N1150);
xor XOR2 (N1387, N1381, N771);
buf BUF1 (N1388, N1385);
buf BUF1 (N1389, N1384);
or OR4 (N1390, N1374, N238, N377, N1328);
nor NOR2 (N1391, N1388, N307);
xor XOR2 (N1392, N1376, N3);
not NOT1 (N1393, N1392);
xor XOR2 (N1394, N1389, N798);
nand NAND2 (N1395, N1372, N520);
or OR3 (N1396, N1393, N351, N76);
nand NAND2 (N1397, N1395, N988);
nor NOR4 (N1398, N1387, N705, N714, N1194);
and AND2 (N1399, N1390, N643);
not NOT1 (N1400, N1377);
and AND3 (N1401, N1383, N803, N115);
nor NOR4 (N1402, N1399, N1097, N263, N335);
nor NOR2 (N1403, N1398, N752);
or OR4 (N1404, N1386, N477, N42, N396);
or OR3 (N1405, N1401, N86, N606);
and AND3 (N1406, N1397, N130, N874);
and AND3 (N1407, N1379, N183, N1180);
xor XOR2 (N1408, N1404, N918);
and AND2 (N1409, N1396, N352);
nor NOR4 (N1410, N1403, N181, N1038, N1166);
nand NAND4 (N1411, N1409, N572, N895, N1035);
nor NOR2 (N1412, N1400, N75);
xor XOR2 (N1413, N1407, N797);
xor XOR2 (N1414, N1405, N443);
not NOT1 (N1415, N1410);
xor XOR2 (N1416, N1415, N318);
buf BUF1 (N1417, N1411);
or OR4 (N1418, N1391, N1145, N1131, N685);
nor NOR2 (N1419, N1412, N1250);
and AND3 (N1420, N1413, N161, N614);
and AND4 (N1421, N1394, N986, N665, N616);
buf BUF1 (N1422, N1421);
buf BUF1 (N1423, N1416);
nand NAND3 (N1424, N1402, N326, N369);
not NOT1 (N1425, N1420);
and AND4 (N1426, N1423, N112, N1215, N528);
not NOT1 (N1427, N1406);
nand NAND3 (N1428, N1417, N1181, N553);
or OR3 (N1429, N1425, N336, N1022);
xor XOR2 (N1430, N1418, N1213);
not NOT1 (N1431, N1426);
and AND2 (N1432, N1422, N814);
xor XOR2 (N1433, N1414, N729);
and AND4 (N1434, N1432, N771, N1043, N509);
buf BUF1 (N1435, N1429);
xor XOR2 (N1436, N1424, N1347);
and AND4 (N1437, N1431, N1048, N207, N1249);
nand NAND2 (N1438, N1427, N307);
or OR3 (N1439, N1437, N1084, N1014);
and AND4 (N1440, N1419, N1023, N1194, N941);
nand NAND4 (N1441, N1434, N845, N662, N332);
nor NOR3 (N1442, N1436, N671, N1431);
not NOT1 (N1443, N1441);
nor NOR3 (N1444, N1443, N241, N213);
not NOT1 (N1445, N1439);
or OR4 (N1446, N1445, N1337, N491, N1053);
not NOT1 (N1447, N1408);
and AND3 (N1448, N1433, N466, N700);
not NOT1 (N1449, N1435);
and AND4 (N1450, N1448, N753, N796, N300);
xor XOR2 (N1451, N1444, N1218);
buf BUF1 (N1452, N1440);
buf BUF1 (N1453, N1446);
not NOT1 (N1454, N1442);
nor NOR3 (N1455, N1451, N286, N1438);
nand NAND2 (N1456, N1317, N540);
or OR3 (N1457, N1455, N370, N454);
and AND2 (N1458, N1447, N429);
nor NOR3 (N1459, N1453, N297, N157);
nor NOR2 (N1460, N1452, N305);
buf BUF1 (N1461, N1449);
nand NAND2 (N1462, N1461, N149);
nor NOR2 (N1463, N1460, N888);
nor NOR3 (N1464, N1463, N1265, N1245);
and AND4 (N1465, N1457, N704, N1427, N760);
nor NOR3 (N1466, N1462, N812, N690);
nand NAND3 (N1467, N1464, N11, N1019);
buf BUF1 (N1468, N1465);
or OR3 (N1469, N1458, N566, N690);
and AND3 (N1470, N1454, N170, N1372);
and AND3 (N1471, N1466, N341, N1039);
buf BUF1 (N1472, N1428);
and AND4 (N1473, N1471, N1077, N135, N316);
nor NOR2 (N1474, N1473, N281);
and AND3 (N1475, N1474, N567, N1078);
nand NAND4 (N1476, N1472, N1215, N1307, N815);
buf BUF1 (N1477, N1467);
xor XOR2 (N1478, N1430, N376);
nor NOR3 (N1479, N1459, N1043, N769);
or OR4 (N1480, N1456, N420, N802, N1237);
buf BUF1 (N1481, N1478);
or OR2 (N1482, N1480, N431);
buf BUF1 (N1483, N1470);
not NOT1 (N1484, N1479);
xor XOR2 (N1485, N1477, N430);
nor NOR3 (N1486, N1484, N1084, N1018);
or OR3 (N1487, N1450, N345, N1103);
and AND4 (N1488, N1486, N1031, N1102, N57);
xor XOR2 (N1489, N1469, N1176);
nand NAND3 (N1490, N1476, N1243, N907);
buf BUF1 (N1491, N1485);
nand NAND3 (N1492, N1491, N18, N433);
and AND2 (N1493, N1481, N564);
and AND2 (N1494, N1488, N1351);
xor XOR2 (N1495, N1493, N338);
and AND4 (N1496, N1492, N581, N699, N258);
and AND4 (N1497, N1489, N92, N572, N586);
nor NOR4 (N1498, N1496, N472, N1133, N389);
nand NAND4 (N1499, N1475, N844, N1409, N236);
buf BUF1 (N1500, N1499);
xor XOR2 (N1501, N1483, N1143);
not NOT1 (N1502, N1494);
not NOT1 (N1503, N1500);
xor XOR2 (N1504, N1497, N672);
and AND3 (N1505, N1495, N1269, N781);
xor XOR2 (N1506, N1502, N211);
xor XOR2 (N1507, N1468, N1036);
buf BUF1 (N1508, N1503);
nor NOR2 (N1509, N1482, N1308);
nand NAND2 (N1510, N1504, N1053);
nand NAND2 (N1511, N1510, N74);
or OR3 (N1512, N1511, N460, N1311);
not NOT1 (N1513, N1487);
or OR2 (N1514, N1508, N703);
xor XOR2 (N1515, N1505, N487);
nor NOR2 (N1516, N1515, N1234);
buf BUF1 (N1517, N1512);
nand NAND2 (N1518, N1501, N833);
nand NAND2 (N1519, N1516, N655);
xor XOR2 (N1520, N1507, N1233);
buf BUF1 (N1521, N1509);
xor XOR2 (N1522, N1514, N1001);
and AND4 (N1523, N1521, N1058, N363, N22);
and AND3 (N1524, N1506, N1047, N820);
not NOT1 (N1525, N1522);
nor NOR2 (N1526, N1524, N73);
and AND4 (N1527, N1518, N746, N836, N89);
buf BUF1 (N1528, N1520);
nor NOR2 (N1529, N1525, N193);
xor XOR2 (N1530, N1528, N236);
buf BUF1 (N1531, N1526);
nor NOR4 (N1532, N1531, N282, N907, N126);
or OR4 (N1533, N1523, N1284, N1233, N95);
or OR3 (N1534, N1513, N552, N593);
and AND2 (N1535, N1517, N1452);
or OR3 (N1536, N1527, N1203, N1219);
buf BUF1 (N1537, N1533);
nand NAND3 (N1538, N1537, N519, N1275);
nand NAND4 (N1539, N1490, N930, N112, N1294);
nand NAND3 (N1540, N1539, N1538, N144);
nor NOR4 (N1541, N676, N439, N911, N323);
nor NOR2 (N1542, N1519, N367);
or OR4 (N1543, N1542, N1116, N1274, N152);
not NOT1 (N1544, N1540);
buf BUF1 (N1545, N1535);
or OR2 (N1546, N1532, N175);
not NOT1 (N1547, N1530);
not NOT1 (N1548, N1546);
nand NAND4 (N1549, N1544, N263, N252, N588);
and AND3 (N1550, N1541, N802, N222);
nand NAND3 (N1551, N1536, N508, N177);
or OR3 (N1552, N1534, N1334, N214);
xor XOR2 (N1553, N1498, N561);
or OR3 (N1554, N1553, N482, N1316);
nor NOR3 (N1555, N1545, N861, N503);
nor NOR2 (N1556, N1551, N1165);
not NOT1 (N1557, N1547);
buf BUF1 (N1558, N1557);
xor XOR2 (N1559, N1529, N1233);
nor NOR3 (N1560, N1556, N655, N168);
buf BUF1 (N1561, N1560);
or OR2 (N1562, N1559, N1154);
not NOT1 (N1563, N1552);
xor XOR2 (N1564, N1563, N873);
nand NAND4 (N1565, N1550, N322, N829, N214);
nand NAND3 (N1566, N1558, N1518, N1142);
nor NOR3 (N1567, N1566, N998, N1385);
xor XOR2 (N1568, N1543, N1532);
nor NOR2 (N1569, N1555, N619);
or OR2 (N1570, N1549, N1078);
xor XOR2 (N1571, N1570, N96);
xor XOR2 (N1572, N1567, N444);
xor XOR2 (N1573, N1572, N982);
and AND2 (N1574, N1562, N409);
nand NAND3 (N1575, N1569, N1222, N1293);
buf BUF1 (N1576, N1561);
nand NAND4 (N1577, N1564, N554, N670, N1000);
or OR2 (N1578, N1577, N723);
buf BUF1 (N1579, N1565);
not NOT1 (N1580, N1574);
and AND3 (N1581, N1571, N358, N891);
or OR3 (N1582, N1548, N1114, N226);
buf BUF1 (N1583, N1579);
xor XOR2 (N1584, N1575, N133);
not NOT1 (N1585, N1580);
xor XOR2 (N1586, N1584, N737);
and AND4 (N1587, N1583, N555, N404, N1086);
and AND3 (N1588, N1585, N1023, N197);
nand NAND4 (N1589, N1554, N1130, N1095, N1137);
buf BUF1 (N1590, N1573);
or OR4 (N1591, N1576, N27, N882, N1293);
not NOT1 (N1592, N1568);
nor NOR4 (N1593, N1581, N799, N31, N385);
buf BUF1 (N1594, N1588);
xor XOR2 (N1595, N1578, N664);
not NOT1 (N1596, N1589);
buf BUF1 (N1597, N1587);
nand NAND2 (N1598, N1595, N396);
or OR2 (N1599, N1592, N1487);
xor XOR2 (N1600, N1598, N488);
and AND2 (N1601, N1594, N1233);
nor NOR4 (N1602, N1597, N151, N328, N423);
buf BUF1 (N1603, N1599);
buf BUF1 (N1604, N1590);
nor NOR4 (N1605, N1591, N921, N235, N1039);
not NOT1 (N1606, N1582);
buf BUF1 (N1607, N1601);
nand NAND3 (N1608, N1602, N1348, N186);
buf BUF1 (N1609, N1586);
buf BUF1 (N1610, N1600);
and AND2 (N1611, N1605, N678);
xor XOR2 (N1612, N1604, N1110);
nor NOR2 (N1613, N1611, N663);
buf BUF1 (N1614, N1596);
or OR3 (N1615, N1608, N206, N1416);
nand NAND3 (N1616, N1610, N326, N368);
nand NAND2 (N1617, N1607, N673);
xor XOR2 (N1618, N1615, N343);
buf BUF1 (N1619, N1603);
and AND2 (N1620, N1609, N471);
xor XOR2 (N1621, N1614, N1508);
buf BUF1 (N1622, N1613);
buf BUF1 (N1623, N1620);
not NOT1 (N1624, N1617);
buf BUF1 (N1625, N1618);
nor NOR3 (N1626, N1622, N225, N662);
nand NAND4 (N1627, N1625, N1154, N1108, N61);
nand NAND4 (N1628, N1606, N1179, N1364, N772);
buf BUF1 (N1629, N1627);
xor XOR2 (N1630, N1612, N6);
buf BUF1 (N1631, N1616);
not NOT1 (N1632, N1630);
xor XOR2 (N1633, N1629, N1164);
nand NAND3 (N1634, N1593, N210, N577);
and AND3 (N1635, N1624, N1328, N1318);
nor NOR3 (N1636, N1619, N505, N1261);
nand NAND3 (N1637, N1632, N333, N1513);
and AND4 (N1638, N1634, N1038, N419, N701);
nand NAND2 (N1639, N1621, N1308);
nor NOR4 (N1640, N1639, N8, N1513, N1013);
or OR2 (N1641, N1633, N64);
nor NOR3 (N1642, N1626, N547, N1484);
buf BUF1 (N1643, N1641);
or OR4 (N1644, N1638, N981, N1107, N1407);
buf BUF1 (N1645, N1636);
nor NOR3 (N1646, N1643, N416, N1604);
and AND2 (N1647, N1640, N120);
xor XOR2 (N1648, N1628, N67);
xor XOR2 (N1649, N1642, N1398);
not NOT1 (N1650, N1648);
or OR3 (N1651, N1631, N655, N741);
buf BUF1 (N1652, N1635);
or OR4 (N1653, N1649, N1032, N207, N287);
not NOT1 (N1654, N1644);
buf BUF1 (N1655, N1654);
nand NAND4 (N1656, N1623, N581, N1614, N50);
xor XOR2 (N1657, N1637, N1432);
and AND2 (N1658, N1646, N749);
and AND2 (N1659, N1656, N689);
and AND3 (N1660, N1655, N632, N1175);
not NOT1 (N1661, N1645);
nand NAND2 (N1662, N1651, N721);
and AND3 (N1663, N1660, N117, N1316);
nor NOR4 (N1664, N1661, N388, N10, N1417);
nand NAND3 (N1665, N1650, N736, N270);
nand NAND4 (N1666, N1665, N1577, N1289, N411);
nor NOR2 (N1667, N1647, N511);
nand NAND4 (N1668, N1657, N1586, N664, N645);
nand NAND2 (N1669, N1658, N388);
nand NAND3 (N1670, N1664, N1326, N1636);
nor NOR2 (N1671, N1667, N979);
nor NOR3 (N1672, N1669, N48, N375);
and AND3 (N1673, N1662, N296, N1194);
and AND2 (N1674, N1670, N635);
not NOT1 (N1675, N1668);
nor NOR2 (N1676, N1675, N660);
or OR4 (N1677, N1659, N929, N1187, N1077);
xor XOR2 (N1678, N1673, N299);
or OR3 (N1679, N1678, N582, N233);
nor NOR3 (N1680, N1676, N699, N974);
and AND3 (N1681, N1666, N1067, N1610);
xor XOR2 (N1682, N1672, N335);
buf BUF1 (N1683, N1652);
or OR3 (N1684, N1680, N1260, N228);
or OR2 (N1685, N1674, N1132);
nor NOR4 (N1686, N1679, N767, N860, N1055);
nor NOR3 (N1687, N1683, N883, N238);
and AND2 (N1688, N1682, N1575);
buf BUF1 (N1689, N1653);
and AND3 (N1690, N1681, N586, N187);
and AND2 (N1691, N1686, N183);
nor NOR3 (N1692, N1677, N180, N1085);
nand NAND2 (N1693, N1688, N198);
not NOT1 (N1694, N1685);
xor XOR2 (N1695, N1693, N136);
and AND3 (N1696, N1687, N1177, N657);
and AND2 (N1697, N1696, N819);
xor XOR2 (N1698, N1694, N765);
not NOT1 (N1699, N1697);
nand NAND2 (N1700, N1663, N559);
not NOT1 (N1701, N1692);
not NOT1 (N1702, N1700);
and AND3 (N1703, N1698, N1388, N838);
not NOT1 (N1704, N1695);
nor NOR3 (N1705, N1701, N1575, N1279);
xor XOR2 (N1706, N1690, N903);
nor NOR3 (N1707, N1684, N1692, N1027);
and AND3 (N1708, N1702, N480, N1072);
buf BUF1 (N1709, N1707);
xor XOR2 (N1710, N1689, N1653);
xor XOR2 (N1711, N1671, N1164);
and AND2 (N1712, N1706, N148);
or OR4 (N1713, N1704, N89, N401, N1541);
and AND3 (N1714, N1691, N1483, N1614);
or OR2 (N1715, N1710, N632);
xor XOR2 (N1716, N1699, N289);
buf BUF1 (N1717, N1716);
nand NAND2 (N1718, N1713, N334);
buf BUF1 (N1719, N1718);
and AND3 (N1720, N1711, N498, N588);
buf BUF1 (N1721, N1703);
and AND3 (N1722, N1714, N584, N1465);
or OR4 (N1723, N1709, N1722, N19, N709);
xor XOR2 (N1724, N49, N1494);
or OR2 (N1725, N1708, N492);
nand NAND2 (N1726, N1719, N284);
and AND2 (N1727, N1721, N866);
xor XOR2 (N1728, N1723, N187);
or OR3 (N1729, N1705, N138, N384);
or OR3 (N1730, N1720, N606, N1610);
not NOT1 (N1731, N1724);
nand NAND2 (N1732, N1717, N1096);
and AND2 (N1733, N1726, N956);
and AND2 (N1734, N1727, N1541);
or OR4 (N1735, N1730, N1149, N1056, N726);
nor NOR2 (N1736, N1733, N1295);
and AND2 (N1737, N1736, N416);
not NOT1 (N1738, N1735);
or OR2 (N1739, N1738, N835);
or OR3 (N1740, N1731, N1102, N733);
buf BUF1 (N1741, N1725);
nor NOR2 (N1742, N1740, N643);
nand NAND3 (N1743, N1734, N472, N1225);
buf BUF1 (N1744, N1741);
buf BUF1 (N1745, N1732);
nor NOR4 (N1746, N1745, N1242, N707, N550);
and AND2 (N1747, N1739, N303);
not NOT1 (N1748, N1728);
xor XOR2 (N1749, N1742, N771);
not NOT1 (N1750, N1744);
or OR4 (N1751, N1750, N879, N680, N980);
buf BUF1 (N1752, N1748);
not NOT1 (N1753, N1715);
nor NOR4 (N1754, N1729, N775, N98, N1659);
nand NAND2 (N1755, N1752, N1017);
xor XOR2 (N1756, N1747, N1690);
nor NOR2 (N1757, N1746, N1568);
and AND4 (N1758, N1754, N1223, N1517, N445);
or OR2 (N1759, N1712, N854);
or OR3 (N1760, N1757, N603, N694);
nor NOR3 (N1761, N1751, N430, N846);
nor NOR4 (N1762, N1759, N1050, N953, N494);
nor NOR2 (N1763, N1760, N65);
or OR2 (N1764, N1758, N1408);
not NOT1 (N1765, N1737);
nor NOR2 (N1766, N1764, N299);
not NOT1 (N1767, N1755);
nor NOR2 (N1768, N1749, N1233);
nand NAND4 (N1769, N1761, N1513, N496, N595);
nor NOR2 (N1770, N1766, N1592);
not NOT1 (N1771, N1743);
not NOT1 (N1772, N1770);
and AND3 (N1773, N1762, N1315, N295);
nand NAND2 (N1774, N1753, N558);
nor NOR3 (N1775, N1769, N1761, N454);
nor NOR3 (N1776, N1765, N886, N1461);
nand NAND2 (N1777, N1768, N1698);
buf BUF1 (N1778, N1773);
not NOT1 (N1779, N1775);
or OR4 (N1780, N1756, N1649, N519, N808);
or OR3 (N1781, N1779, N705, N583);
and AND3 (N1782, N1777, N1646, N1631);
not NOT1 (N1783, N1767);
buf BUF1 (N1784, N1783);
not NOT1 (N1785, N1781);
and AND2 (N1786, N1785, N1775);
buf BUF1 (N1787, N1778);
buf BUF1 (N1788, N1784);
not NOT1 (N1789, N1788);
nor NOR4 (N1790, N1763, N277, N1395, N1239);
xor XOR2 (N1791, N1776, N708);
not NOT1 (N1792, N1782);
or OR3 (N1793, N1787, N1439, N1192);
not NOT1 (N1794, N1786);
or OR4 (N1795, N1794, N1228, N478, N1348);
not NOT1 (N1796, N1795);
or OR4 (N1797, N1774, N1035, N1090, N720);
buf BUF1 (N1798, N1789);
nor NOR4 (N1799, N1790, N791, N1216, N1701);
xor XOR2 (N1800, N1798, N1264);
xor XOR2 (N1801, N1780, N1758);
or OR4 (N1802, N1792, N589, N1151, N180);
not NOT1 (N1803, N1797);
and AND2 (N1804, N1803, N1789);
nor NOR2 (N1805, N1793, N1103);
not NOT1 (N1806, N1800);
buf BUF1 (N1807, N1791);
not NOT1 (N1808, N1796);
or OR3 (N1809, N1808, N163, N720);
and AND2 (N1810, N1805, N1618);
buf BUF1 (N1811, N1801);
or OR4 (N1812, N1811, N607, N403, N285);
or OR2 (N1813, N1806, N127);
or OR2 (N1814, N1802, N972);
buf BUF1 (N1815, N1807);
not NOT1 (N1816, N1771);
xor XOR2 (N1817, N1812, N461);
nor NOR3 (N1818, N1813, N551, N1083);
nor NOR4 (N1819, N1817, N581, N287, N474);
nand NAND3 (N1820, N1810, N1571, N977);
xor XOR2 (N1821, N1820, N767);
nor NOR3 (N1822, N1818, N243, N945);
xor XOR2 (N1823, N1814, N445);
and AND3 (N1824, N1809, N772, N1585);
not NOT1 (N1825, N1824);
or OR3 (N1826, N1799, N619, N1621);
and AND4 (N1827, N1772, N1010, N1754, N80);
xor XOR2 (N1828, N1821, N603);
nor NOR4 (N1829, N1804, N661, N566, N864);
nand NAND4 (N1830, N1822, N169, N1166, N1362);
nand NAND3 (N1831, N1825, N1295, N305);
xor XOR2 (N1832, N1816, N1705);
not NOT1 (N1833, N1826);
xor XOR2 (N1834, N1828, N1635);
buf BUF1 (N1835, N1834);
and AND3 (N1836, N1827, N722, N1141);
nor NOR2 (N1837, N1823, N1140);
and AND4 (N1838, N1829, N500, N316, N1294);
nor NOR3 (N1839, N1832, N679, N285);
buf BUF1 (N1840, N1838);
nand NAND3 (N1841, N1833, N1527, N362);
and AND4 (N1842, N1841, N816, N1106, N1526);
and AND4 (N1843, N1842, N954, N368, N1813);
xor XOR2 (N1844, N1837, N261);
nand NAND2 (N1845, N1836, N580);
xor XOR2 (N1846, N1815, N959);
or OR3 (N1847, N1819, N324, N852);
buf BUF1 (N1848, N1844);
buf BUF1 (N1849, N1831);
nor NOR2 (N1850, N1835, N226);
and AND4 (N1851, N1840, N271, N118, N289);
and AND2 (N1852, N1850, N1279);
not NOT1 (N1853, N1847);
or OR2 (N1854, N1846, N1308);
nand NAND3 (N1855, N1845, N445, N1030);
not NOT1 (N1856, N1843);
nand NAND2 (N1857, N1856, N1645);
nand NAND2 (N1858, N1852, N652);
not NOT1 (N1859, N1858);
and AND3 (N1860, N1830, N1002, N64);
nor NOR2 (N1861, N1855, N1179);
and AND4 (N1862, N1859, N1627, N1581, N1392);
nand NAND4 (N1863, N1854, N788, N1082, N1249);
and AND3 (N1864, N1862, N156, N464);
and AND3 (N1865, N1849, N133, N918);
nor NOR2 (N1866, N1851, N228);
or OR4 (N1867, N1857, N1678, N1406, N855);
nor NOR2 (N1868, N1864, N1832);
not NOT1 (N1869, N1848);
or OR3 (N1870, N1860, N244, N1780);
nor NOR2 (N1871, N1866, N1679);
xor XOR2 (N1872, N1839, N925);
buf BUF1 (N1873, N1865);
buf BUF1 (N1874, N1870);
and AND4 (N1875, N1867, N532, N344, N1044);
or OR2 (N1876, N1871, N1781);
or OR2 (N1877, N1853, N1645);
or OR4 (N1878, N1868, N1462, N827, N996);
xor XOR2 (N1879, N1863, N577);
or OR3 (N1880, N1872, N652, N1669);
nand NAND3 (N1881, N1879, N394, N73);
and AND2 (N1882, N1861, N754);
buf BUF1 (N1883, N1873);
buf BUF1 (N1884, N1874);
nand NAND4 (N1885, N1883, N1290, N787, N435);
not NOT1 (N1886, N1875);
not NOT1 (N1887, N1885);
and AND2 (N1888, N1877, N1726);
and AND4 (N1889, N1887, N256, N1078, N402);
xor XOR2 (N1890, N1878, N558);
and AND2 (N1891, N1888, N1183);
buf BUF1 (N1892, N1876);
xor XOR2 (N1893, N1882, N1074);
and AND4 (N1894, N1884, N1746, N1106, N1354);
not NOT1 (N1895, N1881);
or OR2 (N1896, N1880, N1474);
nand NAND4 (N1897, N1886, N1287, N1483, N997);
xor XOR2 (N1898, N1895, N131);
nor NOR2 (N1899, N1890, N716);
and AND4 (N1900, N1897, N1249, N1231, N1421);
not NOT1 (N1901, N1899);
or OR3 (N1902, N1869, N28, N211);
or OR4 (N1903, N1894, N1477, N1794, N1442);
nor NOR2 (N1904, N1898, N1391);
or OR2 (N1905, N1904, N1201);
and AND3 (N1906, N1902, N2, N462);
buf BUF1 (N1907, N1893);
xor XOR2 (N1908, N1896, N284);
nor NOR2 (N1909, N1907, N780);
not NOT1 (N1910, N1906);
and AND3 (N1911, N1905, N1575, N1745);
not NOT1 (N1912, N1901);
nand NAND3 (N1913, N1900, N684, N34);
buf BUF1 (N1914, N1889);
buf BUF1 (N1915, N1909);
buf BUF1 (N1916, N1910);
not NOT1 (N1917, N1914);
and AND2 (N1918, N1908, N1319);
nor NOR3 (N1919, N1918, N1354, N121);
and AND2 (N1920, N1917, N871);
nand NAND4 (N1921, N1903, N1534, N995, N1463);
not NOT1 (N1922, N1892);
nand NAND4 (N1923, N1911, N147, N1532, N94);
nor NOR2 (N1924, N1920, N1105);
and AND4 (N1925, N1915, N646, N616, N879);
or OR3 (N1926, N1922, N1566, N401);
nand NAND3 (N1927, N1923, N1766, N495);
nor NOR2 (N1928, N1921, N1622);
buf BUF1 (N1929, N1891);
xor XOR2 (N1930, N1913, N1349);
xor XOR2 (N1931, N1926, N1024);
buf BUF1 (N1932, N1930);
nand NAND3 (N1933, N1925, N1007, N1096);
nand NAND2 (N1934, N1927, N118);
buf BUF1 (N1935, N1929);
buf BUF1 (N1936, N1935);
nor NOR3 (N1937, N1934, N1650, N847);
or OR4 (N1938, N1924, N810, N1043, N970);
buf BUF1 (N1939, N1912);
not NOT1 (N1940, N1938);
nand NAND4 (N1941, N1931, N94, N449, N579);
or OR4 (N1942, N1939, N1229, N449, N540);
not NOT1 (N1943, N1937);
not NOT1 (N1944, N1940);
and AND3 (N1945, N1936, N1001, N1196);
buf BUF1 (N1946, N1945);
xor XOR2 (N1947, N1928, N1247);
not NOT1 (N1948, N1933);
xor XOR2 (N1949, N1919, N1260);
nand NAND3 (N1950, N1947, N1156, N802);
buf BUF1 (N1951, N1946);
and AND2 (N1952, N1932, N1686);
nand NAND3 (N1953, N1916, N1452, N1837);
and AND4 (N1954, N1949, N1374, N1520, N793);
and AND4 (N1955, N1954, N939, N1764, N1924);
xor XOR2 (N1956, N1950, N1160);
not NOT1 (N1957, N1953);
or OR4 (N1958, N1956, N980, N843, N1248);
xor XOR2 (N1959, N1952, N1421);
nor NOR4 (N1960, N1957, N1413, N49, N1203);
nand NAND2 (N1961, N1941, N686);
xor XOR2 (N1962, N1948, N743);
not NOT1 (N1963, N1943);
nand NAND3 (N1964, N1955, N1741, N1305);
and AND3 (N1965, N1961, N1805, N1550);
xor XOR2 (N1966, N1951, N595);
not NOT1 (N1967, N1962);
nor NOR2 (N1968, N1964, N1408);
nor NOR3 (N1969, N1959, N682, N1538);
and AND2 (N1970, N1944, N1363);
not NOT1 (N1971, N1942);
or OR4 (N1972, N1969, N480, N1174, N339);
xor XOR2 (N1973, N1972, N605);
not NOT1 (N1974, N1960);
nand NAND2 (N1975, N1963, N1277);
or OR3 (N1976, N1967, N1406, N741);
xor XOR2 (N1977, N1971, N1326);
and AND3 (N1978, N1965, N674, N716);
xor XOR2 (N1979, N1975, N793);
xor XOR2 (N1980, N1978, N304);
buf BUF1 (N1981, N1979);
not NOT1 (N1982, N1976);
buf BUF1 (N1983, N1958);
xor XOR2 (N1984, N1980, N1421);
nor NOR2 (N1985, N1984, N1362);
not NOT1 (N1986, N1985);
buf BUF1 (N1987, N1977);
buf BUF1 (N1988, N1973);
nand NAND2 (N1989, N1970, N654);
or OR3 (N1990, N1989, N1875, N1912);
or OR2 (N1991, N1988, N1329);
xor XOR2 (N1992, N1987, N531);
buf BUF1 (N1993, N1981);
buf BUF1 (N1994, N1982);
nand NAND4 (N1995, N1974, N522, N851, N478);
and AND4 (N1996, N1968, N567, N652, N501);
buf BUF1 (N1997, N1993);
buf BUF1 (N1998, N1995);
or OR3 (N1999, N1991, N1770, N815);
and AND3 (N2000, N1966, N258, N24);
buf BUF1 (N2001, N1990);
buf BUF1 (N2002, N1994);
buf BUF1 (N2003, N1983);
not NOT1 (N2004, N2001);
and AND2 (N2005, N1996, N1632);
nand NAND4 (N2006, N1986, N899, N1068, N884);
and AND4 (N2007, N1998, N1234, N1308, N1509);
buf BUF1 (N2008, N1999);
buf BUF1 (N2009, N2008);
or OR3 (N2010, N2006, N2005, N1538);
or OR2 (N2011, N831, N196);
buf BUF1 (N2012, N1997);
not NOT1 (N2013, N2012);
nand NAND2 (N2014, N2007, N1981);
and AND3 (N2015, N1992, N1562, N1841);
and AND3 (N2016, N2002, N740, N1968);
and AND4 (N2017, N2000, N85, N1267, N713);
or OR3 (N2018, N2011, N1544, N110);
nand NAND3 (N2019, N2013, N1925, N1280);
and AND3 (N2020, N2009, N1437, N1771);
nand NAND3 (N2021, N2004, N1405, N416);
buf BUF1 (N2022, N2003);
not NOT1 (N2023, N2018);
and AND4 (N2024, N2017, N163, N1737, N1140);
nand NAND3 (N2025, N2023, N1725, N1169);
xor XOR2 (N2026, N2019, N448);
nor NOR2 (N2027, N2022, N1013);
nand NAND4 (N2028, N2014, N699, N1863, N546);
nand NAND2 (N2029, N2020, N1350);
xor XOR2 (N2030, N2015, N1822);
and AND3 (N2031, N2016, N1650, N1219);
nand NAND3 (N2032, N2024, N1394, N498);
or OR3 (N2033, N2029, N630, N1907);
nand NAND3 (N2034, N2025, N12, N289);
xor XOR2 (N2035, N2027, N535);
not NOT1 (N2036, N2033);
nor NOR4 (N2037, N2031, N1041, N593, N487);
or OR4 (N2038, N2021, N2003, N973, N948);
xor XOR2 (N2039, N2010, N693);
not NOT1 (N2040, N2035);
nor NOR2 (N2041, N2030, N1095);
nand NAND3 (N2042, N2034, N1185, N318);
nand NAND4 (N2043, N2038, N1862, N933, N1436);
nand NAND2 (N2044, N2041, N528);
nand NAND2 (N2045, N2043, N926);
and AND4 (N2046, N2045, N714, N590, N170);
xor XOR2 (N2047, N2037, N1278);
nor NOR3 (N2048, N2036, N117, N129);
buf BUF1 (N2049, N2028);
not NOT1 (N2050, N2040);
nor NOR3 (N2051, N2044, N846, N108);
nand NAND3 (N2052, N2049, N1968, N1321);
nand NAND4 (N2053, N2047, N1300, N277, N1197);
xor XOR2 (N2054, N2052, N1124);
buf BUF1 (N2055, N2046);
not NOT1 (N2056, N2048);
xor XOR2 (N2057, N2042, N1349);
not NOT1 (N2058, N2055);
and AND2 (N2059, N2057, N1785);
not NOT1 (N2060, N2051);
buf BUF1 (N2061, N2026);
and AND3 (N2062, N2053, N645, N177);
and AND4 (N2063, N2056, N1779, N1188, N1741);
nand NAND4 (N2064, N2060, N680, N1808, N1681);
buf BUF1 (N2065, N2062);
xor XOR2 (N2066, N2064, N1419);
buf BUF1 (N2067, N2061);
nor NOR2 (N2068, N2059, N777);
nor NOR2 (N2069, N2050, N476);
not NOT1 (N2070, N2054);
nor NOR4 (N2071, N2058, N1009, N1929, N1870);
or OR2 (N2072, N2068, N86);
not NOT1 (N2073, N2039);
buf BUF1 (N2074, N2032);
and AND2 (N2075, N2073, N1297);
nand NAND3 (N2076, N2069, N58, N1900);
xor XOR2 (N2077, N2063, N1130);
not NOT1 (N2078, N2075);
xor XOR2 (N2079, N2074, N1682);
nor NOR2 (N2080, N2078, N675);
xor XOR2 (N2081, N2077, N1343);
xor XOR2 (N2082, N2081, N1902);
xor XOR2 (N2083, N2071, N286);
nand NAND4 (N2084, N2083, N822, N235, N1441);
nor NOR3 (N2085, N2076, N1380, N70);
not NOT1 (N2086, N2079);
xor XOR2 (N2087, N2072, N146);
or OR3 (N2088, N2087, N489, N1087);
or OR4 (N2089, N2080, N750, N1351, N139);
nand NAND3 (N2090, N2070, N1549, N778);
buf BUF1 (N2091, N2066);
xor XOR2 (N2092, N2065, N2078);
not NOT1 (N2093, N2089);
nand NAND4 (N2094, N2082, N1301, N1993, N971);
nor NOR4 (N2095, N2088, N2075, N1666, N1567);
buf BUF1 (N2096, N2093);
not NOT1 (N2097, N2086);
not NOT1 (N2098, N2085);
and AND4 (N2099, N2084, N1033, N222, N1863);
xor XOR2 (N2100, N2099, N1739);
buf BUF1 (N2101, N2067);
xor XOR2 (N2102, N2091, N690);
nor NOR3 (N2103, N2097, N837, N1702);
buf BUF1 (N2104, N2095);
buf BUF1 (N2105, N2103);
buf BUF1 (N2106, N2105);
not NOT1 (N2107, N2102);
and AND2 (N2108, N2101, N830);
buf BUF1 (N2109, N2092);
buf BUF1 (N2110, N2108);
or OR2 (N2111, N2104, N676);
nand NAND3 (N2112, N2110, N1157, N498);
not NOT1 (N2113, N2094);
buf BUF1 (N2114, N2109);
nand NAND2 (N2115, N2100, N1916);
nand NAND4 (N2116, N2112, N1676, N517, N1900);
nand NAND4 (N2117, N2098, N2083, N1645, N713);
buf BUF1 (N2118, N2117);
or OR3 (N2119, N2106, N277, N155);
not NOT1 (N2120, N2115);
nand NAND3 (N2121, N2090, N1904, N762);
or OR2 (N2122, N2107, N1537);
nor NOR2 (N2123, N2119, N1021);
nor NOR4 (N2124, N2111, N712, N1553, N1459);
nor NOR4 (N2125, N2121, N1678, N1594, N1305);
or OR4 (N2126, N2120, N1621, N1177, N1664);
and AND3 (N2127, N2122, N2107, N37);
and AND2 (N2128, N2125, N1411);
xor XOR2 (N2129, N2114, N303);
not NOT1 (N2130, N2096);
or OR4 (N2131, N2123, N1293, N1216, N1063);
not NOT1 (N2132, N2118);
buf BUF1 (N2133, N2127);
xor XOR2 (N2134, N2124, N331);
buf BUF1 (N2135, N2132);
nor NOR4 (N2136, N2131, N188, N1281, N353);
buf BUF1 (N2137, N2129);
xor XOR2 (N2138, N2116, N1091);
nor NOR2 (N2139, N2136, N846);
nand NAND2 (N2140, N2138, N98);
nor NOR3 (N2141, N2126, N958, N1076);
or OR4 (N2142, N2134, N240, N1067, N836);
nand NAND4 (N2143, N2137, N346, N673, N200);
buf BUF1 (N2144, N2135);
not NOT1 (N2145, N2141);
nor NOR3 (N2146, N2113, N1626, N303);
and AND2 (N2147, N2142, N314);
nand NAND3 (N2148, N2133, N999, N1160);
nor NOR4 (N2149, N2140, N259, N1699, N1054);
nor NOR2 (N2150, N2139, N1239);
or OR4 (N2151, N2148, N1367, N1591, N1866);
nand NAND2 (N2152, N2145, N173);
buf BUF1 (N2153, N2143);
nor NOR4 (N2154, N2150, N1289, N898, N1431);
xor XOR2 (N2155, N2147, N1299);
and AND2 (N2156, N2152, N1405);
not NOT1 (N2157, N2156);
buf BUF1 (N2158, N2144);
and AND2 (N2159, N2146, N112);
nand NAND3 (N2160, N2155, N1635, N683);
or OR3 (N2161, N2151, N1819, N637);
nor NOR3 (N2162, N2130, N116, N311);
nor NOR2 (N2163, N2162, N933);
buf BUF1 (N2164, N2153);
xor XOR2 (N2165, N2128, N2019);
not NOT1 (N2166, N2163);
buf BUF1 (N2167, N2154);
or OR2 (N2168, N2149, N362);
and AND4 (N2169, N2165, N1711, N229, N1365);
nand NAND2 (N2170, N2166, N971);
nor NOR2 (N2171, N2157, N844);
or OR2 (N2172, N2158, N838);
and AND4 (N2173, N2164, N1208, N1535, N66);
buf BUF1 (N2174, N2168);
xor XOR2 (N2175, N2170, N1523);
nor NOR4 (N2176, N2173, N1385, N1259, N1893);
nand NAND2 (N2177, N2171, N800);
or OR3 (N2178, N2172, N71, N542);
not NOT1 (N2179, N2167);
xor XOR2 (N2180, N2177, N1719);
buf BUF1 (N2181, N2161);
and AND4 (N2182, N2159, N1830, N1214, N848);
xor XOR2 (N2183, N2176, N350);
buf BUF1 (N2184, N2178);
nand NAND4 (N2185, N2179, N1747, N1631, N231);
buf BUF1 (N2186, N2180);
nor NOR4 (N2187, N2175, N1048, N1406, N246);
nand NAND3 (N2188, N2187, N415, N1881);
xor XOR2 (N2189, N2181, N1824);
or OR2 (N2190, N2184, N948);
or OR4 (N2191, N2185, N491, N43, N2132);
xor XOR2 (N2192, N2189, N1346);
xor XOR2 (N2193, N2160, N1421);
nand NAND3 (N2194, N2182, N669, N477);
xor XOR2 (N2195, N2191, N2134);
or OR2 (N2196, N2195, N1110);
xor XOR2 (N2197, N2190, N214);
or OR3 (N2198, N2197, N915, N1075);
not NOT1 (N2199, N2196);
nor NOR4 (N2200, N2199, N1882, N958, N715);
xor XOR2 (N2201, N2186, N1633);
buf BUF1 (N2202, N2188);
xor XOR2 (N2203, N2169, N1752);
xor XOR2 (N2204, N2198, N908);
nand NAND2 (N2205, N2174, N1359);
buf BUF1 (N2206, N2194);
nand NAND2 (N2207, N2203, N1549);
nand NAND2 (N2208, N2183, N1153);
not NOT1 (N2209, N2202);
xor XOR2 (N2210, N2204, N1381);
nand NAND4 (N2211, N2207, N170, N1563, N1760);
nor NOR4 (N2212, N2210, N1175, N1638, N1512);
buf BUF1 (N2213, N2208);
nor NOR4 (N2214, N2213, N2103, N2102, N2109);
nand NAND3 (N2215, N2200, N1970, N538);
buf BUF1 (N2216, N2205);
nor NOR3 (N2217, N2192, N725, N1082);
xor XOR2 (N2218, N2217, N1790);
xor XOR2 (N2219, N2215, N104);
not NOT1 (N2220, N2218);
nand NAND4 (N2221, N2211, N1243, N470, N372);
or OR2 (N2222, N2209, N2009);
nand NAND2 (N2223, N2221, N1912);
nor NOR4 (N2224, N2220, N528, N75, N1244);
and AND3 (N2225, N2212, N530, N655);
or OR2 (N2226, N2206, N2077);
and AND4 (N2227, N2201, N35, N2134, N1115);
nand NAND2 (N2228, N2216, N1483);
and AND4 (N2229, N2226, N1297, N1485, N1781);
and AND3 (N2230, N2193, N971, N799);
not NOT1 (N2231, N2214);
or OR2 (N2232, N2231, N1468);
xor XOR2 (N2233, N2223, N2093);
xor XOR2 (N2234, N2228, N967);
buf BUF1 (N2235, N2230);
buf BUF1 (N2236, N2227);
buf BUF1 (N2237, N2233);
nor NOR3 (N2238, N2232, N1764, N1054);
buf BUF1 (N2239, N2224);
and AND4 (N2240, N2222, N2097, N938, N1461);
or OR3 (N2241, N2236, N2110, N1593);
nand NAND4 (N2242, N2241, N2215, N437, N473);
nor NOR3 (N2243, N2229, N2062, N1740);
nand NAND2 (N2244, N2238, N902);
buf BUF1 (N2245, N2239);
xor XOR2 (N2246, N2245, N534);
xor XOR2 (N2247, N2243, N1477);
not NOT1 (N2248, N2240);
not NOT1 (N2249, N2248);
or OR4 (N2250, N2249, N153, N2238, N827);
not NOT1 (N2251, N2235);
not NOT1 (N2252, N2247);
not NOT1 (N2253, N2244);
buf BUF1 (N2254, N2225);
and AND3 (N2255, N2219, N552, N738);
and AND2 (N2256, N2234, N1444);
nand NAND4 (N2257, N2242, N1804, N1429, N2033);
nor NOR4 (N2258, N2255, N551, N2135, N679);
not NOT1 (N2259, N2250);
not NOT1 (N2260, N2254);
not NOT1 (N2261, N2259);
xor XOR2 (N2262, N2260, N711);
not NOT1 (N2263, N2256);
or OR2 (N2264, N2261, N1012);
xor XOR2 (N2265, N2263, N271);
nand NAND3 (N2266, N2251, N804, N216);
or OR4 (N2267, N2266, N122, N1222, N401);
buf BUF1 (N2268, N2267);
buf BUF1 (N2269, N2268);
not NOT1 (N2270, N2258);
buf BUF1 (N2271, N2246);
buf BUF1 (N2272, N2264);
xor XOR2 (N2273, N2265, N956);
nor NOR2 (N2274, N2262, N1585);
nand NAND3 (N2275, N2274, N1173, N1404);
not NOT1 (N2276, N2237);
buf BUF1 (N2277, N2253);
or OR3 (N2278, N2277, N1691, N1690);
nand NAND2 (N2279, N2269, N676);
nand NAND4 (N2280, N2272, N1639, N1050, N946);
xor XOR2 (N2281, N2270, N511);
and AND3 (N2282, N2281, N1558, N833);
and AND3 (N2283, N2282, N328, N1602);
not NOT1 (N2284, N2252);
not NOT1 (N2285, N2278);
buf BUF1 (N2286, N2285);
buf BUF1 (N2287, N2257);
buf BUF1 (N2288, N2275);
and AND4 (N2289, N2276, N177, N861, N1760);
or OR4 (N2290, N2283, N1779, N1004, N284);
or OR3 (N2291, N2288, N2045, N731);
or OR4 (N2292, N2287, N2014, N859, N918);
or OR2 (N2293, N2290, N2203);
nor NOR3 (N2294, N2271, N1762, N2029);
nor NOR4 (N2295, N2292, N751, N1701, N657);
not NOT1 (N2296, N2293);
buf BUF1 (N2297, N2273);
xor XOR2 (N2298, N2294, N957);
nand NAND2 (N2299, N2297, N812);
or OR4 (N2300, N2289, N648, N1788, N1008);
or OR4 (N2301, N2279, N474, N768, N1764);
and AND2 (N2302, N2295, N2295);
not NOT1 (N2303, N2284);
not NOT1 (N2304, N2280);
not NOT1 (N2305, N2300);
or OR3 (N2306, N2298, N906, N1570);
and AND4 (N2307, N2305, N542, N1897, N1514);
nor NOR3 (N2308, N2304, N1099, N613);
xor XOR2 (N2309, N2307, N938);
and AND4 (N2310, N2296, N1539, N2176, N1594);
and AND4 (N2311, N2303, N562, N1616, N1556);
nor NOR4 (N2312, N2308, N692, N394, N274);
not NOT1 (N2313, N2286);
nor NOR4 (N2314, N2310, N1481, N256, N1621);
or OR3 (N2315, N2301, N1392, N1542);
not NOT1 (N2316, N2311);
nor NOR2 (N2317, N2315, N1067);
buf BUF1 (N2318, N2299);
or OR4 (N2319, N2317, N1275, N1483, N235);
and AND4 (N2320, N2312, N1358, N1128, N213);
nor NOR4 (N2321, N2318, N1300, N1668, N1341);
xor XOR2 (N2322, N2321, N1995);
nor NOR2 (N2323, N2291, N852);
not NOT1 (N2324, N2309);
nand NAND4 (N2325, N2306, N1617, N1627, N37);
nor NOR4 (N2326, N2319, N2064, N1554, N1778);
not NOT1 (N2327, N2316);
nand NAND2 (N2328, N2325, N875);
and AND2 (N2329, N2322, N932);
nor NOR2 (N2330, N2302, N186);
buf BUF1 (N2331, N2314);
or OR3 (N2332, N2329, N1338, N2271);
nand NAND2 (N2333, N2313, N2283);
or OR2 (N2334, N2331, N2275);
or OR3 (N2335, N2334, N679, N705);
nor NOR2 (N2336, N2335, N15);
or OR4 (N2337, N2327, N983, N1099, N1437);
nand NAND4 (N2338, N2326, N985, N386, N1357);
or OR4 (N2339, N2330, N313, N988, N2335);
nand NAND2 (N2340, N2324, N633);
buf BUF1 (N2341, N2320);
or OR3 (N2342, N2328, N763, N1663);
buf BUF1 (N2343, N2333);
not NOT1 (N2344, N2332);
buf BUF1 (N2345, N2340);
xor XOR2 (N2346, N2337, N1007);
nor NOR4 (N2347, N2339, N749, N43, N292);
nor NOR4 (N2348, N2338, N1108, N1468, N364);
and AND2 (N2349, N2323, N1282);
or OR4 (N2350, N2346, N1529, N521, N2105);
not NOT1 (N2351, N2342);
nand NAND4 (N2352, N2348, N1216, N2006, N780);
xor XOR2 (N2353, N2350, N17);
or OR3 (N2354, N2341, N458, N220);
and AND4 (N2355, N2352, N1614, N567, N158);
or OR4 (N2356, N2336, N602, N689, N734);
not NOT1 (N2357, N2345);
or OR3 (N2358, N2357, N2143, N879);
nand NAND3 (N2359, N2347, N451, N2335);
not NOT1 (N2360, N2343);
nor NOR4 (N2361, N2358, N1791, N1011, N2217);
xor XOR2 (N2362, N2356, N984);
not NOT1 (N2363, N2344);
nand NAND3 (N2364, N2351, N445, N2332);
xor XOR2 (N2365, N2359, N2253);
nand NAND2 (N2366, N2360, N249);
xor XOR2 (N2367, N2362, N1353);
or OR3 (N2368, N2365, N1008, N361);
and AND3 (N2369, N2363, N1859, N1991);
xor XOR2 (N2370, N2354, N478);
xor XOR2 (N2371, N2366, N542);
nor NOR3 (N2372, N2371, N419, N1651);
xor XOR2 (N2373, N2369, N2331);
and AND2 (N2374, N2353, N439);
nor NOR3 (N2375, N2370, N14, N831);
or OR3 (N2376, N2375, N1832, N832);
not NOT1 (N2377, N2372);
or OR3 (N2378, N2368, N2058, N235);
nand NAND2 (N2379, N2377, N1639);
or OR3 (N2380, N2373, N721, N1731);
buf BUF1 (N2381, N2361);
nand NAND4 (N2382, N2367, N808, N784, N1905);
not NOT1 (N2383, N2380);
xor XOR2 (N2384, N2382, N595);
nor NOR4 (N2385, N2355, N886, N254, N1511);
or OR4 (N2386, N2384, N1369, N117, N846);
nor NOR2 (N2387, N2383, N800);
or OR3 (N2388, N2364, N1973, N1317);
and AND4 (N2389, N2386, N852, N688, N1526);
nand NAND4 (N2390, N2376, N1539, N316, N355);
or OR2 (N2391, N2381, N1089);
xor XOR2 (N2392, N2388, N646);
and AND4 (N2393, N2349, N465, N76, N834);
nand NAND2 (N2394, N2379, N641);
nor NOR4 (N2395, N2393, N1999, N1704, N103);
nor NOR3 (N2396, N2387, N2130, N76);
or OR3 (N2397, N2391, N42, N1446);
not NOT1 (N2398, N2385);
not NOT1 (N2399, N2394);
xor XOR2 (N2400, N2374, N1707);
nor NOR2 (N2401, N2395, N746);
or OR4 (N2402, N2398, N619, N1694, N2095);
nand NAND2 (N2403, N2400, N329);
nand NAND2 (N2404, N2392, N1087);
nor NOR2 (N2405, N2390, N177);
xor XOR2 (N2406, N2403, N942);
and AND2 (N2407, N2406, N50);
or OR4 (N2408, N2389, N1517, N580, N2377);
nand NAND3 (N2409, N2402, N2097, N256);
or OR3 (N2410, N2401, N1632, N273);
buf BUF1 (N2411, N2410);
and AND4 (N2412, N2404, N1450, N687, N998);
not NOT1 (N2413, N2378);
not NOT1 (N2414, N2411);
nor NOR4 (N2415, N2399, N1187, N1532, N915);
xor XOR2 (N2416, N2409, N446);
nand NAND4 (N2417, N2397, N1812, N2029, N1240);
xor XOR2 (N2418, N2413, N1278);
buf BUF1 (N2419, N2408);
nand NAND2 (N2420, N2412, N1435);
buf BUF1 (N2421, N2414);
nor NOR4 (N2422, N2405, N548, N407, N1541);
xor XOR2 (N2423, N2407, N947);
nor NOR4 (N2424, N2423, N1840, N361, N157);
not NOT1 (N2425, N2396);
and AND3 (N2426, N2417, N1955, N1402);
not NOT1 (N2427, N2421);
not NOT1 (N2428, N2427);
buf BUF1 (N2429, N2422);
xor XOR2 (N2430, N2429, N139);
buf BUF1 (N2431, N2430);
nor NOR3 (N2432, N2428, N2425, N402);
not NOT1 (N2433, N1553);
not NOT1 (N2434, N2416);
nand NAND2 (N2435, N2434, N961);
buf BUF1 (N2436, N2431);
xor XOR2 (N2437, N2419, N677);
not NOT1 (N2438, N2435);
and AND2 (N2439, N2418, N755);
and AND4 (N2440, N2437, N1778, N1523, N1663);
nor NOR4 (N2441, N2424, N1729, N311, N1640);
nor NOR4 (N2442, N2438, N1858, N861, N1512);
not NOT1 (N2443, N2426);
buf BUF1 (N2444, N2443);
and AND4 (N2445, N2415, N1377, N826, N1163);
nor NOR2 (N2446, N2441, N510);
or OR3 (N2447, N2433, N919, N517);
nor NOR2 (N2448, N2420, N750);
not NOT1 (N2449, N2442);
or OR3 (N2450, N2445, N1701, N1994);
or OR2 (N2451, N2440, N803);
not NOT1 (N2452, N2448);
buf BUF1 (N2453, N2450);
or OR3 (N2454, N2444, N105, N257);
xor XOR2 (N2455, N2452, N2169);
not NOT1 (N2456, N2455);
or OR4 (N2457, N2451, N2071, N1021, N1277);
nand NAND2 (N2458, N2432, N2107);
nor NOR3 (N2459, N2456, N2325, N2379);
nor NOR4 (N2460, N2446, N2266, N1457, N2008);
buf BUF1 (N2461, N2458);
xor XOR2 (N2462, N2449, N1554);
nor NOR3 (N2463, N2436, N1311, N1096);
nor NOR2 (N2464, N2453, N451);
nand NAND4 (N2465, N2454, N2454, N2310, N795);
xor XOR2 (N2466, N2465, N421);
xor XOR2 (N2467, N2447, N183);
or OR3 (N2468, N2461, N2327, N2275);
or OR3 (N2469, N2463, N1158, N1342);
nand NAND4 (N2470, N2439, N2405, N945, N2090);
nor NOR2 (N2471, N2466, N906);
nand NAND3 (N2472, N2457, N338, N670);
xor XOR2 (N2473, N2470, N2326);
buf BUF1 (N2474, N2472);
buf BUF1 (N2475, N2474);
buf BUF1 (N2476, N2467);
and AND3 (N2477, N2476, N31, N2443);
and AND2 (N2478, N2475, N1860);
xor XOR2 (N2479, N2478, N1271);
nor NOR3 (N2480, N2464, N2179, N2066);
buf BUF1 (N2481, N2468);
nand NAND4 (N2482, N2479, N1701, N1039, N154);
nand NAND2 (N2483, N2473, N2094);
nor NOR3 (N2484, N2471, N1428, N898);
nand NAND4 (N2485, N2477, N1177, N2306, N827);
nor NOR4 (N2486, N2484, N25, N578, N1298);
nand NAND4 (N2487, N2481, N80, N2286, N2289);
nor NOR4 (N2488, N2480, N340, N1543, N1122);
nand NAND2 (N2489, N2488, N1033);
not NOT1 (N2490, N2486);
nand NAND4 (N2491, N2483, N1420, N2215, N73);
or OR2 (N2492, N2489, N1931);
buf BUF1 (N2493, N2482);
nor NOR4 (N2494, N2469, N905, N6, N309);
not NOT1 (N2495, N2459);
or OR4 (N2496, N2491, N2121, N236, N2344);
buf BUF1 (N2497, N2487);
or OR4 (N2498, N2496, N1744, N2144, N1470);
and AND2 (N2499, N2492, N1743);
nor NOR4 (N2500, N2498, N1329, N2200, N739);
or OR2 (N2501, N2499, N1211);
nor NOR3 (N2502, N2494, N1034, N1741);
xor XOR2 (N2503, N2462, N1287);
buf BUF1 (N2504, N2490);
nor NOR4 (N2505, N2493, N1111, N1033, N99);
not NOT1 (N2506, N2500);
and AND3 (N2507, N2505, N284, N174);
not NOT1 (N2508, N2506);
nor NOR3 (N2509, N2507, N650, N532);
not NOT1 (N2510, N2497);
not NOT1 (N2511, N2502);
not NOT1 (N2512, N2508);
xor XOR2 (N2513, N2509, N1656);
or OR3 (N2514, N2503, N1504, N2170);
and AND4 (N2515, N2460, N1793, N1115, N1823);
buf BUF1 (N2516, N2514);
nand NAND2 (N2517, N2510, N1971);
buf BUF1 (N2518, N2516);
nor NOR4 (N2519, N2495, N539, N1802, N1619);
nand NAND2 (N2520, N2515, N1492);
not NOT1 (N2521, N2518);
buf BUF1 (N2522, N2520);
nand NAND2 (N2523, N2513, N192);
xor XOR2 (N2524, N2522, N45);
not NOT1 (N2525, N2523);
xor XOR2 (N2526, N2524, N2091);
or OR2 (N2527, N2519, N897);
or OR2 (N2528, N2526, N221);
xor XOR2 (N2529, N2521, N1424);
nand NAND4 (N2530, N2501, N1841, N2281, N2477);
nand NAND2 (N2531, N2504, N198);
and AND4 (N2532, N2525, N2014, N2082, N1552);
not NOT1 (N2533, N2511);
not NOT1 (N2534, N2532);
nand NAND2 (N2535, N2517, N1321);
not NOT1 (N2536, N2529);
buf BUF1 (N2537, N2533);
nand NAND3 (N2538, N2534, N1364, N815);
xor XOR2 (N2539, N2512, N629);
not NOT1 (N2540, N2535);
or OR3 (N2541, N2540, N821, N737);
not NOT1 (N2542, N2538);
not NOT1 (N2543, N2531);
or OR3 (N2544, N2530, N184, N582);
nor NOR4 (N2545, N2543, N2059, N1231, N1178);
xor XOR2 (N2546, N2537, N631);
and AND2 (N2547, N2541, N1680);
or OR3 (N2548, N2545, N1858, N281);
not NOT1 (N2549, N2527);
nand NAND2 (N2550, N2536, N1106);
nor NOR3 (N2551, N2548, N2273, N508);
xor XOR2 (N2552, N2528, N1943);
not NOT1 (N2553, N2552);
or OR4 (N2554, N2553, N850, N1132, N2173);
nor NOR3 (N2555, N2554, N743, N509);
or OR4 (N2556, N2551, N428, N772, N1271);
nand NAND4 (N2557, N2546, N1128, N995, N1711);
buf BUF1 (N2558, N2539);
nor NOR2 (N2559, N2550, N404);
and AND2 (N2560, N2556, N1626);
buf BUF1 (N2561, N2544);
nand NAND4 (N2562, N2542, N2321, N2238, N361);
xor XOR2 (N2563, N2560, N2005);
nor NOR2 (N2564, N2561, N793);
xor XOR2 (N2565, N2485, N2316);
xor XOR2 (N2566, N2565, N2264);
and AND2 (N2567, N2555, N211);
and AND2 (N2568, N2562, N1364);
and AND3 (N2569, N2564, N2540, N1505);
and AND4 (N2570, N2549, N989, N1928, N2155);
xor XOR2 (N2571, N2547, N2099);
xor XOR2 (N2572, N2558, N466);
nand NAND4 (N2573, N2568, N2407, N2528, N348);
not NOT1 (N2574, N2563);
buf BUF1 (N2575, N2574);
buf BUF1 (N2576, N2573);
xor XOR2 (N2577, N2557, N1782);
and AND2 (N2578, N2577, N269);
nand NAND2 (N2579, N2570, N1084);
buf BUF1 (N2580, N2575);
or OR3 (N2581, N2559, N254, N1580);
nor NOR4 (N2582, N2580, N1328, N1810, N509);
nand NAND4 (N2583, N2582, N743, N2492, N1786);
not NOT1 (N2584, N2581);
and AND2 (N2585, N2583, N576);
nor NOR3 (N2586, N2572, N2454, N177);
not NOT1 (N2587, N2567);
and AND4 (N2588, N2578, N2476, N91, N1179);
not NOT1 (N2589, N2571);
nand NAND3 (N2590, N2586, N2088, N1562);
nor NOR2 (N2591, N2587, N612);
or OR3 (N2592, N2590, N864, N312);
buf BUF1 (N2593, N2569);
nor NOR2 (N2594, N2588, N900);
not NOT1 (N2595, N2566);
or OR2 (N2596, N2585, N1139);
and AND4 (N2597, N2595, N2566, N1103, N572);
and AND4 (N2598, N2593, N1727, N229, N1849);
xor XOR2 (N2599, N2594, N408);
nand NAND2 (N2600, N2596, N2211);
not NOT1 (N2601, N2589);
and AND3 (N2602, N2592, N408, N468);
xor XOR2 (N2603, N2599, N2271);
not NOT1 (N2604, N2584);
not NOT1 (N2605, N2579);
buf BUF1 (N2606, N2597);
xor XOR2 (N2607, N2603, N1591);
or OR4 (N2608, N2605, N158, N185, N1051);
buf BUF1 (N2609, N2600);
not NOT1 (N2610, N2604);
xor XOR2 (N2611, N2602, N1894);
and AND3 (N2612, N2610, N2228, N445);
nor NOR4 (N2613, N2591, N767, N2113, N1015);
and AND4 (N2614, N2598, N1402, N1952, N2267);
or OR3 (N2615, N2607, N1919, N1035);
not NOT1 (N2616, N2612);
nor NOR3 (N2617, N2616, N358, N1524);
not NOT1 (N2618, N2615);
nor NOR3 (N2619, N2611, N2435, N2282);
not NOT1 (N2620, N2608);
not NOT1 (N2621, N2576);
xor XOR2 (N2622, N2620, N1455);
and AND2 (N2623, N2621, N2390);
and AND4 (N2624, N2606, N1754, N524, N290);
buf BUF1 (N2625, N2614);
and AND4 (N2626, N2625, N2310, N2276, N1920);
and AND2 (N2627, N2623, N251);
nand NAND3 (N2628, N2617, N1015, N1757);
nor NOR3 (N2629, N2626, N2002, N1619);
nand NAND4 (N2630, N2628, N2129, N1634, N629);
buf BUF1 (N2631, N2627);
buf BUF1 (N2632, N2630);
xor XOR2 (N2633, N2631, N2161);
or OR4 (N2634, N2619, N1283, N1138, N213);
or OR4 (N2635, N2613, N729, N48, N2069);
or OR4 (N2636, N2632, N299, N403, N2333);
xor XOR2 (N2637, N2601, N2393);
or OR2 (N2638, N2636, N2176);
xor XOR2 (N2639, N2637, N1094);
nand NAND4 (N2640, N2624, N790, N315, N2388);
buf BUF1 (N2641, N2609);
not NOT1 (N2642, N2640);
nand NAND4 (N2643, N2642, N47, N1184, N1099);
buf BUF1 (N2644, N2643);
xor XOR2 (N2645, N2644, N994);
xor XOR2 (N2646, N2618, N1860);
not NOT1 (N2647, N2638);
nand NAND4 (N2648, N2641, N715, N129, N1607);
and AND4 (N2649, N2645, N458, N2180, N858);
not NOT1 (N2650, N2648);
nand NAND4 (N2651, N2647, N573, N583, N1769);
or OR2 (N2652, N2633, N1526);
or OR4 (N2653, N2639, N2042, N376, N96);
xor XOR2 (N2654, N2635, N838);
or OR4 (N2655, N2634, N1794, N609, N1798);
nor NOR3 (N2656, N2629, N340, N2182);
nand NAND2 (N2657, N2656, N329);
or OR4 (N2658, N2657, N1189, N825, N571);
nand NAND2 (N2659, N2654, N2083);
xor XOR2 (N2660, N2649, N971);
and AND3 (N2661, N2660, N591, N1973);
nand NAND4 (N2662, N2652, N1981, N105, N2645);
and AND2 (N2663, N2650, N1547);
and AND3 (N2664, N2646, N1112, N604);
not NOT1 (N2665, N2664);
not NOT1 (N2666, N2662);
buf BUF1 (N2667, N2659);
or OR3 (N2668, N2663, N2415, N1541);
nor NOR3 (N2669, N2661, N301, N507);
nor NOR3 (N2670, N2653, N2526, N693);
or OR2 (N2671, N2670, N695);
nand NAND4 (N2672, N2669, N727, N1916, N1757);
buf BUF1 (N2673, N2666);
not NOT1 (N2674, N2668);
nor NOR3 (N2675, N2673, N2662, N2316);
xor XOR2 (N2676, N2672, N1485);
or OR2 (N2677, N2651, N2025);
nand NAND3 (N2678, N2665, N2153, N2157);
buf BUF1 (N2679, N2678);
buf BUF1 (N2680, N2676);
buf BUF1 (N2681, N2675);
and AND4 (N2682, N2680, N94, N2070, N2387);
nand NAND2 (N2683, N2622, N1535);
nor NOR3 (N2684, N2679, N2627, N1020);
xor XOR2 (N2685, N2677, N1747);
xor XOR2 (N2686, N2683, N2290);
or OR3 (N2687, N2684, N970, N694);
not NOT1 (N2688, N2681);
or OR4 (N2689, N2655, N1058, N1453, N216);
or OR3 (N2690, N2688, N773, N198);
and AND4 (N2691, N2687, N1560, N2402, N1114);
and AND4 (N2692, N2690, N36, N1807, N1435);
buf BUF1 (N2693, N2686);
nor NOR4 (N2694, N2674, N1251, N918, N999);
nand NAND4 (N2695, N2682, N2082, N1979, N2610);
nor NOR2 (N2696, N2692, N2628);
xor XOR2 (N2697, N2685, N43);
or OR4 (N2698, N2691, N2399, N664, N746);
or OR2 (N2699, N2698, N394);
and AND3 (N2700, N2699, N1067, N2069);
xor XOR2 (N2701, N2695, N1577);
or OR2 (N2702, N2671, N503);
buf BUF1 (N2703, N2700);
and AND2 (N2704, N2693, N2091);
nor NOR3 (N2705, N2704, N1514, N385);
nor NOR3 (N2706, N2667, N403, N2341);
nor NOR3 (N2707, N2694, N1330, N2080);
nand NAND2 (N2708, N2689, N496);
nor NOR2 (N2709, N2706, N1549);
xor XOR2 (N2710, N2707, N128);
or OR4 (N2711, N2708, N361, N964, N1135);
buf BUF1 (N2712, N2711);
or OR4 (N2713, N2710, N753, N1942, N932);
xor XOR2 (N2714, N2697, N993);
nand NAND3 (N2715, N2709, N656, N275);
nand NAND2 (N2716, N2714, N736);
xor XOR2 (N2717, N2701, N1623);
and AND4 (N2718, N2705, N242, N2180, N2222);
xor XOR2 (N2719, N2696, N1899);
or OR2 (N2720, N2702, N837);
not NOT1 (N2721, N2716);
and AND3 (N2722, N2703, N411, N2084);
or OR4 (N2723, N2712, N1724, N1079, N1240);
nor NOR4 (N2724, N2715, N575, N2402, N427);
and AND4 (N2725, N2724, N1216, N1263, N197);
buf BUF1 (N2726, N2721);
nor NOR4 (N2727, N2726, N2062, N114, N1318);
nor NOR4 (N2728, N2723, N528, N473, N1332);
not NOT1 (N2729, N2725);
buf BUF1 (N2730, N2658);
or OR3 (N2731, N2718, N1199, N2222);
xor XOR2 (N2732, N2730, N2329);
nor NOR2 (N2733, N2722, N861);
not NOT1 (N2734, N2733);
nor NOR2 (N2735, N2713, N61);
buf BUF1 (N2736, N2727);
xor XOR2 (N2737, N2731, N2393);
nor NOR3 (N2738, N2729, N2631, N318);
and AND2 (N2739, N2737, N1885);
nand NAND3 (N2740, N2736, N1022, N1265);
and AND3 (N2741, N2738, N775, N1774);
buf BUF1 (N2742, N2734);
nand NAND2 (N2743, N2739, N2546);
not NOT1 (N2744, N2743);
buf BUF1 (N2745, N2744);
not NOT1 (N2746, N2720);
not NOT1 (N2747, N2717);
or OR4 (N2748, N2719, N234, N2014, N1808);
and AND2 (N2749, N2728, N749);
or OR3 (N2750, N2732, N1278, N1871);
and AND4 (N2751, N2750, N1733, N724, N1451);
buf BUF1 (N2752, N2751);
not NOT1 (N2753, N2747);
nand NAND3 (N2754, N2752, N2666, N236);
nand NAND3 (N2755, N2748, N1565, N2570);
xor XOR2 (N2756, N2749, N300);
nand NAND3 (N2757, N2740, N2417, N1219);
buf BUF1 (N2758, N2741);
xor XOR2 (N2759, N2745, N2419);
not NOT1 (N2760, N2746);
xor XOR2 (N2761, N2742, N2583);
not NOT1 (N2762, N2757);
nand NAND4 (N2763, N2754, N2225, N1760, N2577);
xor XOR2 (N2764, N2755, N427);
and AND2 (N2765, N2763, N2442);
xor XOR2 (N2766, N2765, N532);
not NOT1 (N2767, N2756);
or OR3 (N2768, N2735, N1032, N990);
nor NOR4 (N2769, N2753, N752, N1267, N796);
not NOT1 (N2770, N2760);
nor NOR3 (N2771, N2770, N1959, N2665);
not NOT1 (N2772, N2771);
nor NOR2 (N2773, N2766, N703);
nand NAND4 (N2774, N2768, N1497, N595, N514);
buf BUF1 (N2775, N2761);
not NOT1 (N2776, N2767);
buf BUF1 (N2777, N2764);
nor NOR3 (N2778, N2772, N750, N884);
nand NAND4 (N2779, N2773, N1615, N2338, N771);
and AND3 (N2780, N2779, N1564, N1498);
nand NAND2 (N2781, N2759, N1499);
nand NAND2 (N2782, N2762, N321);
not NOT1 (N2783, N2782);
nand NAND4 (N2784, N2758, N1269, N2345, N2643);
xor XOR2 (N2785, N2774, N1102);
and AND4 (N2786, N2783, N595, N384, N1101);
nand NAND3 (N2787, N2769, N2629, N169);
xor XOR2 (N2788, N2775, N1233);
and AND2 (N2789, N2780, N1240);
nand NAND3 (N2790, N2786, N1258, N2723);
and AND4 (N2791, N2788, N1779, N2077, N2268);
or OR3 (N2792, N2778, N1230, N703);
or OR3 (N2793, N2781, N1101, N27);
or OR2 (N2794, N2776, N1930);
nand NAND3 (N2795, N2791, N177, N2531);
buf BUF1 (N2796, N2790);
not NOT1 (N2797, N2784);
not NOT1 (N2798, N2785);
and AND2 (N2799, N2792, N1661);
or OR3 (N2800, N2794, N71, N198);
buf BUF1 (N2801, N2795);
not NOT1 (N2802, N2793);
or OR4 (N2803, N2777, N1354, N181, N423);
nand NAND3 (N2804, N2789, N2203, N739);
xor XOR2 (N2805, N2798, N872);
xor XOR2 (N2806, N2802, N1285);
buf BUF1 (N2807, N2806);
xor XOR2 (N2808, N2797, N1161);
not NOT1 (N2809, N2808);
or OR4 (N2810, N2807, N1742, N345, N2014);
or OR2 (N2811, N2804, N2715);
and AND2 (N2812, N2803, N750);
xor XOR2 (N2813, N2812, N795);
and AND4 (N2814, N2813, N2234, N524, N1149);
and AND2 (N2815, N2800, N197);
and AND4 (N2816, N2787, N2030, N1692, N564);
not NOT1 (N2817, N2809);
and AND3 (N2818, N2810, N2454, N1263);
nor NOR3 (N2819, N2805, N2814, N2089);
and AND3 (N2820, N1845, N1585, N1893);
not NOT1 (N2821, N2801);
not NOT1 (N2822, N2819);
nor NOR3 (N2823, N2799, N696, N771);
or OR4 (N2824, N2815, N2696, N1982, N579);
nand NAND3 (N2825, N2818, N1230, N264);
buf BUF1 (N2826, N2821);
and AND2 (N2827, N2826, N32);
nand NAND4 (N2828, N2824, N1405, N958, N1689);
not NOT1 (N2829, N2811);
and AND4 (N2830, N2816, N1268, N1113, N2308);
nand NAND4 (N2831, N2822, N753, N642, N1366);
buf BUF1 (N2832, N2830);
or OR3 (N2833, N2823, N2569, N1037);
or OR4 (N2834, N2829, N1636, N317, N574);
nor NOR3 (N2835, N2834, N2061, N352);
or OR3 (N2836, N2828, N2581, N2441);
not NOT1 (N2837, N2832);
and AND2 (N2838, N2820, N2106);
buf BUF1 (N2839, N2827);
or OR3 (N2840, N2817, N1787, N2131);
and AND3 (N2841, N2840, N2637, N1263);
xor XOR2 (N2842, N2796, N1178);
not NOT1 (N2843, N2836);
buf BUF1 (N2844, N2838);
or OR3 (N2845, N2839, N652, N1610);
nor NOR3 (N2846, N2845, N2740, N792);
and AND2 (N2847, N2831, N45);
and AND4 (N2848, N2841, N699, N2129, N193);
xor XOR2 (N2849, N2837, N1055);
not NOT1 (N2850, N2842);
nand NAND2 (N2851, N2846, N1067);
or OR2 (N2852, N2825, N243);
nand NAND2 (N2853, N2847, N1672);
xor XOR2 (N2854, N2849, N562);
nand NAND4 (N2855, N2833, N1654, N2102, N2691);
nand NAND2 (N2856, N2855, N1852);
nand NAND4 (N2857, N2852, N1900, N2834, N2020);
or OR2 (N2858, N2850, N2094);
or OR3 (N2859, N2858, N1320, N2594);
not NOT1 (N2860, N2857);
buf BUF1 (N2861, N2860);
not NOT1 (N2862, N2859);
and AND4 (N2863, N2861, N1812, N204, N2059);
nor NOR3 (N2864, N2835, N2532, N593);
nor NOR4 (N2865, N2844, N2738, N174, N2709);
or OR4 (N2866, N2864, N832, N1604, N1229);
not NOT1 (N2867, N2863);
buf BUF1 (N2868, N2843);
nor NOR2 (N2869, N2851, N2410);
nand NAND3 (N2870, N2854, N1553, N1439);
nor NOR2 (N2871, N2865, N232);
and AND4 (N2872, N2870, N1907, N1981, N1448);
buf BUF1 (N2873, N2862);
nand NAND4 (N2874, N2867, N978, N1723, N751);
buf BUF1 (N2875, N2874);
buf BUF1 (N2876, N2848);
nor NOR3 (N2877, N2869, N2607, N2620);
and AND3 (N2878, N2877, N1245, N1518);
or OR3 (N2879, N2868, N163, N1138);
nor NOR2 (N2880, N2873, N2651);
and AND3 (N2881, N2879, N22, N2360);
nor NOR4 (N2882, N2853, N1327, N545, N325);
and AND2 (N2883, N2878, N2317);
or OR3 (N2884, N2875, N1845, N604);
nor NOR4 (N2885, N2876, N2720, N1979, N1820);
and AND3 (N2886, N2884, N953, N940);
nand NAND4 (N2887, N2883, N2136, N559, N373);
not NOT1 (N2888, N2856);
not NOT1 (N2889, N2880);
buf BUF1 (N2890, N2882);
nand NAND4 (N2891, N2887, N2867, N1554, N2415);
buf BUF1 (N2892, N2872);
and AND2 (N2893, N2885, N349);
nand NAND4 (N2894, N2891, N1596, N2676, N1120);
and AND3 (N2895, N2894, N1236, N1654);
or OR4 (N2896, N2886, N2694, N2317, N914);
nor NOR2 (N2897, N2866, N1756);
nor NOR3 (N2898, N2890, N2435, N1510);
nand NAND4 (N2899, N2881, N598, N604, N1365);
nor NOR2 (N2900, N2871, N1731);
not NOT1 (N2901, N2888);
or OR4 (N2902, N2901, N178, N2886, N1376);
or OR4 (N2903, N2896, N2878, N2509, N1466);
or OR4 (N2904, N2889, N2390, N1593, N2617);
nor NOR2 (N2905, N2893, N2481);
nand NAND3 (N2906, N2903, N651, N1254);
buf BUF1 (N2907, N2906);
and AND3 (N2908, N2899, N1321, N1441);
xor XOR2 (N2909, N2907, N998);
and AND3 (N2910, N2900, N1852, N1012);
or OR2 (N2911, N2908, N636);
nand NAND3 (N2912, N2897, N576, N248);
nor NOR3 (N2913, N2911, N932, N2643);
buf BUF1 (N2914, N2895);
nand NAND2 (N2915, N2910, N1200);
nor NOR4 (N2916, N2905, N1808, N696, N2310);
and AND2 (N2917, N2904, N1356);
nor NOR4 (N2918, N2915, N1183, N2048, N1643);
not NOT1 (N2919, N2892);
buf BUF1 (N2920, N2898);
buf BUF1 (N2921, N2914);
not NOT1 (N2922, N2918);
not NOT1 (N2923, N2909);
and AND3 (N2924, N2902, N86, N656);
and AND4 (N2925, N2923, N377, N2114, N539);
not NOT1 (N2926, N2920);
not NOT1 (N2927, N2925);
xor XOR2 (N2928, N2912, N2736);
or OR4 (N2929, N2917, N668, N1638, N1164);
nor NOR2 (N2930, N2929, N2698);
not NOT1 (N2931, N2916);
and AND4 (N2932, N2928, N2543, N2487, N2169);
or OR2 (N2933, N2927, N1566);
xor XOR2 (N2934, N2919, N68);
and AND4 (N2935, N2932, N1631, N1245, N2709);
and AND2 (N2936, N2922, N547);
nand NAND2 (N2937, N2921, N2891);
not NOT1 (N2938, N2937);
or OR3 (N2939, N2933, N2704, N1942);
nor NOR3 (N2940, N2930, N2873, N1620);
nor NOR4 (N2941, N2924, N442, N2670, N1520);
xor XOR2 (N2942, N2940, N1454);
buf BUF1 (N2943, N2935);
buf BUF1 (N2944, N2942);
nor NOR4 (N2945, N2936, N2675, N1528, N354);
buf BUF1 (N2946, N2943);
and AND4 (N2947, N2946, N1936, N2280, N443);
xor XOR2 (N2948, N2938, N642);
buf BUF1 (N2949, N2948);
not NOT1 (N2950, N2941);
or OR3 (N2951, N2944, N1873, N619);
not NOT1 (N2952, N2951);
xor XOR2 (N2953, N2950, N843);
nand NAND4 (N2954, N2945, N1034, N902, N1970);
not NOT1 (N2955, N2954);
and AND4 (N2956, N2953, N416, N2132, N1316);
buf BUF1 (N2957, N2939);
nor NOR4 (N2958, N2931, N1924, N96, N2846);
nor NOR2 (N2959, N2957, N2933);
xor XOR2 (N2960, N2947, N1623);
nor NOR3 (N2961, N2926, N2496, N678);
nor NOR4 (N2962, N2960, N2900, N2267, N2722);
xor XOR2 (N2963, N2956, N1347);
or OR4 (N2964, N2952, N1772, N247, N143);
xor XOR2 (N2965, N2961, N2657);
and AND3 (N2966, N2955, N1203, N1524);
nor NOR3 (N2967, N2913, N2674, N2207);
nor NOR3 (N2968, N2965, N1010, N246);
not NOT1 (N2969, N2964);
and AND4 (N2970, N2934, N2386, N708, N2934);
and AND2 (N2971, N2962, N2611);
xor XOR2 (N2972, N2959, N403);
nand NAND2 (N2973, N2966, N1581);
or OR2 (N2974, N2970, N1172);
nor NOR3 (N2975, N2974, N1475, N550);
or OR3 (N2976, N2949, N1878, N1975);
and AND4 (N2977, N2963, N821, N1495, N2935);
or OR3 (N2978, N2973, N1480, N1375);
xor XOR2 (N2979, N2977, N1189);
nor NOR4 (N2980, N2968, N2761, N1998, N1196);
and AND3 (N2981, N2969, N1167, N406);
and AND2 (N2982, N2976, N1322);
not NOT1 (N2983, N2975);
xor XOR2 (N2984, N2981, N348);
not NOT1 (N2985, N2978);
not NOT1 (N2986, N2980);
buf BUF1 (N2987, N2971);
nand NAND4 (N2988, N2983, N1425, N1928, N1089);
nand NAND2 (N2989, N2984, N1844);
or OR4 (N2990, N2985, N1642, N1409, N180);
not NOT1 (N2991, N2990);
nor NOR4 (N2992, N2988, N1905, N2782, N558);
nor NOR3 (N2993, N2991, N54, N1179);
buf BUF1 (N2994, N2987);
nand NAND2 (N2995, N2986, N1624);
not NOT1 (N2996, N2967);
nor NOR2 (N2997, N2958, N102);
nor NOR2 (N2998, N2982, N1319);
nor NOR4 (N2999, N2992, N1781, N2161, N56);
nor NOR4 (N3000, N2979, N2398, N2782, N731);
nor NOR4 (N3001, N2997, N2184, N8, N110);
nor NOR2 (N3002, N3001, N1858);
not NOT1 (N3003, N2993);
nor NOR2 (N3004, N2989, N174);
nand NAND2 (N3005, N3000, N614);
or OR2 (N3006, N3004, N423);
and AND4 (N3007, N3002, N411, N395, N2149);
nand NAND2 (N3008, N3006, N587);
xor XOR2 (N3009, N2995, N1117);
buf BUF1 (N3010, N3009);
and AND3 (N3011, N2999, N1032, N1383);
and AND3 (N3012, N2996, N88, N2740);
not NOT1 (N3013, N3012);
and AND3 (N3014, N2994, N2970, N1333);
not NOT1 (N3015, N2998);
buf BUF1 (N3016, N3005);
or OR4 (N3017, N3003, N376, N1668, N2525);
buf BUF1 (N3018, N3013);
nor NOR2 (N3019, N3015, N2473);
nand NAND2 (N3020, N3014, N539);
not NOT1 (N3021, N3008);
nand NAND4 (N3022, N3017, N2089, N528, N2780);
not NOT1 (N3023, N3011);
nor NOR2 (N3024, N3021, N1959);
xor XOR2 (N3025, N3016, N243);
nor NOR3 (N3026, N3024, N1869, N1128);
nor NOR2 (N3027, N3022, N923);
nor NOR4 (N3028, N3010, N1154, N633, N449);
nand NAND3 (N3029, N3019, N1885, N734);
nor NOR2 (N3030, N3023, N2954);
or OR2 (N3031, N3025, N1666);
not NOT1 (N3032, N3027);
and AND4 (N3033, N3020, N1258, N1690, N2679);
and AND4 (N3034, N3007, N299, N1474, N1960);
nand NAND4 (N3035, N3031, N527, N536, N748);
not NOT1 (N3036, N2972);
nand NAND3 (N3037, N3029, N1532, N922);
not NOT1 (N3038, N3037);
not NOT1 (N3039, N3030);
buf BUF1 (N3040, N3036);
and AND2 (N3041, N3034, N2876);
buf BUF1 (N3042, N3033);
xor XOR2 (N3043, N3040, N3024);
nor NOR3 (N3044, N3028, N174, N318);
nor NOR4 (N3045, N3041, N1701, N2824, N2149);
nand NAND4 (N3046, N3026, N2262, N1870, N2008);
not NOT1 (N3047, N3038);
nor NOR3 (N3048, N3047, N1862, N2359);
and AND4 (N3049, N3044, N1902, N2157, N918);
nor NOR3 (N3050, N3043, N813, N2096);
or OR2 (N3051, N3032, N2589);
nand NAND3 (N3052, N3018, N2882, N1751);
and AND4 (N3053, N3050, N1921, N195, N1668);
xor XOR2 (N3054, N3035, N936);
nand NAND2 (N3055, N3051, N1158);
and AND4 (N3056, N3042, N2396, N397, N187);
nand NAND3 (N3057, N3039, N2009, N2946);
nor NOR2 (N3058, N3052, N58);
not NOT1 (N3059, N3045);
buf BUF1 (N3060, N3048);
buf BUF1 (N3061, N3054);
not NOT1 (N3062, N3055);
nor NOR3 (N3063, N3049, N1357, N1875);
xor XOR2 (N3064, N3058, N2073);
nand NAND4 (N3065, N3062, N2984, N2417, N235);
buf BUF1 (N3066, N3057);
xor XOR2 (N3067, N3063, N1534);
nand NAND4 (N3068, N3066, N1815, N372, N512);
or OR4 (N3069, N3046, N734, N2031, N2902);
and AND3 (N3070, N3067, N2751, N1714);
nor NOR3 (N3071, N3053, N883, N1892);
nand NAND4 (N3072, N3056, N878, N372, N1778);
not NOT1 (N3073, N3059);
or OR4 (N3074, N3070, N153, N1671, N38);
buf BUF1 (N3075, N3068);
nor NOR2 (N3076, N3072, N1268);
buf BUF1 (N3077, N3071);
nor NOR3 (N3078, N3077, N2263, N1826);
nand NAND4 (N3079, N3075, N2883, N2521, N1522);
nand NAND3 (N3080, N3064, N2665, N430);
buf BUF1 (N3081, N3080);
or OR3 (N3082, N3078, N2287, N1397);
xor XOR2 (N3083, N3076, N3074);
not NOT1 (N3084, N2549);
nand NAND4 (N3085, N3073, N2472, N686, N2144);
buf BUF1 (N3086, N3079);
xor XOR2 (N3087, N3081, N1300);
nand NAND4 (N3088, N3060, N2777, N2330, N1983);
xor XOR2 (N3089, N3087, N2913);
not NOT1 (N3090, N3085);
and AND2 (N3091, N3061, N2441);
xor XOR2 (N3092, N3091, N2626);
or OR2 (N3093, N3083, N2449);
xor XOR2 (N3094, N3069, N1816);
nor NOR2 (N3095, N3086, N549);
buf BUF1 (N3096, N3089);
buf BUF1 (N3097, N3090);
nand NAND2 (N3098, N3082, N213);
xor XOR2 (N3099, N3095, N411);
not NOT1 (N3100, N3099);
nor NOR4 (N3101, N3093, N2304, N1756, N713);
not NOT1 (N3102, N3097);
nand NAND4 (N3103, N3101, N752, N832, N1499);
buf BUF1 (N3104, N3096);
and AND2 (N3105, N3098, N2540);
or OR4 (N3106, N3100, N2126, N2352, N2006);
xor XOR2 (N3107, N3104, N388);
nand NAND4 (N3108, N3094, N1875, N2846, N291);
or OR4 (N3109, N3108, N66, N2234, N1530);
nor NOR3 (N3110, N3084, N1585, N333);
nor NOR4 (N3111, N3109, N2501, N2698, N2085);
or OR4 (N3112, N3107, N765, N2021, N2804);
nor NOR3 (N3113, N3106, N2588, N46);
nor NOR3 (N3114, N3113, N2364, N214);
nand NAND3 (N3115, N3112, N2290, N1170);
xor XOR2 (N3116, N3088, N1253);
xor XOR2 (N3117, N3116, N2253);
nand NAND3 (N3118, N3065, N1210, N3020);
and AND3 (N3119, N3103, N1399, N518);
nor NOR4 (N3120, N3118, N2863, N2383, N1084);
and AND3 (N3121, N3092, N199, N897);
not NOT1 (N3122, N3119);
and AND4 (N3123, N3111, N1659, N477, N808);
and AND2 (N3124, N3115, N12);
xor XOR2 (N3125, N3102, N2589);
or OR4 (N3126, N3125, N1137, N299, N1866);
or OR3 (N3127, N3114, N2424, N2956);
or OR3 (N3128, N3117, N554, N2735);
nand NAND4 (N3129, N3128, N940, N1371, N2089);
xor XOR2 (N3130, N3121, N119);
or OR3 (N3131, N3126, N647, N255);
xor XOR2 (N3132, N3122, N1749);
or OR4 (N3133, N3132, N307, N1836, N2145);
nand NAND4 (N3134, N3120, N2967, N1235, N2204);
buf BUF1 (N3135, N3127);
nand NAND2 (N3136, N3129, N2088);
or OR2 (N3137, N3136, N688);
nor NOR2 (N3138, N3110, N1145);
xor XOR2 (N3139, N3130, N2563);
xor XOR2 (N3140, N3135, N1457);
xor XOR2 (N3141, N3124, N875);
nand NAND2 (N3142, N3131, N2808);
or OR4 (N3143, N3123, N553, N949, N2774);
nand NAND2 (N3144, N3143, N1515);
not NOT1 (N3145, N3142);
buf BUF1 (N3146, N3134);
xor XOR2 (N3147, N3138, N1273);
or OR2 (N3148, N3139, N1678);
nand NAND4 (N3149, N3147, N2302, N421, N2937);
and AND2 (N3150, N3140, N2486);
or OR2 (N3151, N3145, N2563);
nand NAND2 (N3152, N3133, N2788);
buf BUF1 (N3153, N3148);
nand NAND2 (N3154, N3137, N543);
buf BUF1 (N3155, N3105);
xor XOR2 (N3156, N3151, N900);
not NOT1 (N3157, N3156);
buf BUF1 (N3158, N3153);
buf BUF1 (N3159, N3141);
nand NAND3 (N3160, N3144, N1547, N3074);
not NOT1 (N3161, N3158);
and AND4 (N3162, N3152, N2416, N1684, N2438);
not NOT1 (N3163, N3159);
not NOT1 (N3164, N3162);
xor XOR2 (N3165, N3161, N1351);
buf BUF1 (N3166, N3155);
or OR3 (N3167, N3165, N2825, N1500);
nand NAND4 (N3168, N3166, N730, N1214, N2254);
buf BUF1 (N3169, N3168);
or OR3 (N3170, N3167, N2453, N1530);
xor XOR2 (N3171, N3154, N2676);
or OR3 (N3172, N3169, N1676, N2404);
or OR4 (N3173, N3157, N864, N141, N935);
nor NOR3 (N3174, N3172, N2786, N20);
nor NOR2 (N3175, N3173, N3160);
nor NOR3 (N3176, N2440, N1227, N388);
or OR3 (N3177, N3174, N1048, N768);
nand NAND4 (N3178, N3163, N3160, N1655, N519);
xor XOR2 (N3179, N3146, N1569);
or OR2 (N3180, N3164, N2902);
nand NAND3 (N3181, N3180, N836, N310);
xor XOR2 (N3182, N3150, N278);
not NOT1 (N3183, N3170);
and AND4 (N3184, N3171, N1937, N519, N1423);
and AND3 (N3185, N3175, N814, N734);
and AND4 (N3186, N3182, N2310, N2429, N1531);
or OR3 (N3187, N3181, N2987, N2694);
nor NOR4 (N3188, N3176, N3116, N2693, N349);
or OR3 (N3189, N3186, N1343, N1258);
nor NOR2 (N3190, N3184, N746);
nand NAND2 (N3191, N3179, N69);
or OR3 (N3192, N3191, N2208, N1644);
and AND2 (N3193, N3189, N954);
buf BUF1 (N3194, N3178);
buf BUF1 (N3195, N3193);
and AND3 (N3196, N3188, N1912, N2645);
nor NOR3 (N3197, N3194, N1651, N474);
and AND3 (N3198, N3190, N1999, N2843);
or OR4 (N3199, N3196, N153, N2333, N2804);
xor XOR2 (N3200, N3149, N733);
nand NAND2 (N3201, N3183, N1886);
not NOT1 (N3202, N3185);
not NOT1 (N3203, N3198);
or OR3 (N3204, N3197, N2254, N2814);
nor NOR2 (N3205, N3202, N814);
not NOT1 (N3206, N3204);
nand NAND3 (N3207, N3195, N615, N1906);
xor XOR2 (N3208, N3207, N2971);
or OR3 (N3209, N3199, N3113, N2929);
and AND2 (N3210, N3205, N1433);
xor XOR2 (N3211, N3201, N1349);
nor NOR2 (N3212, N3177, N872);
or OR2 (N3213, N3203, N2904);
xor XOR2 (N3214, N3212, N3050);
nand NAND4 (N3215, N3211, N2993, N275, N1303);
nor NOR3 (N3216, N3206, N689, N2001);
nand NAND3 (N3217, N3209, N1224, N1668);
xor XOR2 (N3218, N3200, N347);
xor XOR2 (N3219, N3192, N2193);
or OR2 (N3220, N3187, N2312);
xor XOR2 (N3221, N3210, N2967);
nand NAND2 (N3222, N3217, N785);
and AND2 (N3223, N3222, N2982);
buf BUF1 (N3224, N3219);
not NOT1 (N3225, N3224);
and AND2 (N3226, N3218, N2908);
nor NOR3 (N3227, N3216, N1339, N3157);
nand NAND4 (N3228, N3225, N1594, N2500, N1873);
xor XOR2 (N3229, N3220, N358);
buf BUF1 (N3230, N3223);
xor XOR2 (N3231, N3213, N1806);
nand NAND2 (N3232, N3231, N1365);
nand NAND4 (N3233, N3208, N1711, N421, N2960);
nor NOR4 (N3234, N3233, N971, N2572, N1501);
nor NOR3 (N3235, N3227, N2719, N3023);
buf BUF1 (N3236, N3235);
xor XOR2 (N3237, N3230, N627);
nor NOR2 (N3238, N3232, N1121);
nand NAND3 (N3239, N3221, N84, N3070);
or OR2 (N3240, N3237, N113);
or OR4 (N3241, N3215, N611, N2404, N317);
or OR4 (N3242, N3234, N1594, N2638, N2139);
or OR2 (N3243, N3228, N2807);
buf BUF1 (N3244, N3238);
buf BUF1 (N3245, N3244);
and AND3 (N3246, N3236, N2255, N250);
and AND2 (N3247, N3226, N2297);
and AND2 (N3248, N3242, N2907);
or OR2 (N3249, N3240, N101);
or OR4 (N3250, N3241, N215, N2566, N2061);
buf BUF1 (N3251, N3250);
nand NAND4 (N3252, N3246, N892, N2477, N1279);
nand NAND3 (N3253, N3239, N2869, N3136);
or OR3 (N3254, N3253, N1545, N3116);
and AND4 (N3255, N3247, N3070, N2989, N2174);
xor XOR2 (N3256, N3229, N29);
xor XOR2 (N3257, N3251, N51);
buf BUF1 (N3258, N3249);
and AND2 (N3259, N3257, N40);
buf BUF1 (N3260, N3254);
or OR3 (N3261, N3256, N2493, N882);
xor XOR2 (N3262, N3245, N449);
and AND2 (N3263, N3252, N1542);
or OR2 (N3264, N3258, N2163);
not NOT1 (N3265, N3259);
and AND2 (N3266, N3214, N712);
nand NAND3 (N3267, N3255, N1532, N3230);
nor NOR3 (N3268, N3263, N1825, N737);
not NOT1 (N3269, N3261);
nand NAND2 (N3270, N3248, N2556);
nor NOR4 (N3271, N3266, N1006, N2039, N32);
or OR3 (N3272, N3270, N390, N175);
and AND2 (N3273, N3264, N2062);
buf BUF1 (N3274, N3269);
nor NOR2 (N3275, N3268, N557);
nor NOR4 (N3276, N3275, N2809, N646, N709);
and AND4 (N3277, N3276, N446, N1339, N2302);
nor NOR4 (N3278, N3273, N647, N963, N1377);
nand NAND4 (N3279, N3243, N441, N938, N1538);
nand NAND3 (N3280, N3277, N2306, N800);
xor XOR2 (N3281, N3265, N97);
nand NAND4 (N3282, N3281, N1367, N2137, N2854);
not NOT1 (N3283, N3274);
buf BUF1 (N3284, N3271);
nand NAND2 (N3285, N3262, N823);
buf BUF1 (N3286, N3282);
xor XOR2 (N3287, N3279, N2798);
not NOT1 (N3288, N3285);
nor NOR3 (N3289, N3267, N3071, N1962);
or OR3 (N3290, N3289, N1370, N2872);
buf BUF1 (N3291, N3272);
buf BUF1 (N3292, N3278);
nand NAND3 (N3293, N3260, N1018, N555);
nand NAND4 (N3294, N3288, N2294, N3004, N2460);
buf BUF1 (N3295, N3283);
xor XOR2 (N3296, N3280, N448);
not NOT1 (N3297, N3296);
nand NAND3 (N3298, N3286, N930, N729);
nand NAND4 (N3299, N3295, N2270, N3196, N2525);
not NOT1 (N3300, N3297);
buf BUF1 (N3301, N3292);
and AND4 (N3302, N3301, N1488, N669, N3289);
not NOT1 (N3303, N3284);
and AND3 (N3304, N3293, N1806, N3264);
buf BUF1 (N3305, N3300);
or OR4 (N3306, N3305, N2094, N1138, N3005);
not NOT1 (N3307, N3291);
nor NOR3 (N3308, N3302, N2830, N1835);
or OR2 (N3309, N3304, N1355);
and AND3 (N3310, N3306, N2242, N3163);
buf BUF1 (N3311, N3307);
or OR3 (N3312, N3290, N1428, N943);
not NOT1 (N3313, N3310);
or OR4 (N3314, N3308, N1073, N233, N2839);
not NOT1 (N3315, N3311);
nor NOR3 (N3316, N3315, N1896, N515);
not NOT1 (N3317, N3314);
or OR3 (N3318, N3317, N1898, N3287);
or OR4 (N3319, N264, N242, N2473, N1105);
xor XOR2 (N3320, N3313, N2270);
nor NOR3 (N3321, N3294, N1471, N961);
xor XOR2 (N3322, N3309, N3091);
buf BUF1 (N3323, N3316);
buf BUF1 (N3324, N3319);
and AND4 (N3325, N3318, N2332, N965, N2263);
xor XOR2 (N3326, N3303, N3178);
buf BUF1 (N3327, N3320);
xor XOR2 (N3328, N3321, N837);
not NOT1 (N3329, N3312);
buf BUF1 (N3330, N3327);
buf BUF1 (N3331, N3330);
buf BUF1 (N3332, N3323);
nand NAND3 (N3333, N3326, N3201, N225);
xor XOR2 (N3334, N3322, N982);
and AND4 (N3335, N3325, N1078, N1392, N3268);
xor XOR2 (N3336, N3331, N50);
xor XOR2 (N3337, N3299, N2675);
buf BUF1 (N3338, N3333);
xor XOR2 (N3339, N3338, N2854);
or OR3 (N3340, N3298, N598, N2533);
or OR3 (N3341, N3334, N605, N3154);
not NOT1 (N3342, N3335);
nand NAND4 (N3343, N3342, N398, N1158, N3086);
nand NAND3 (N3344, N3332, N2041, N1968);
nor NOR2 (N3345, N3343, N313);
not NOT1 (N3346, N3345);
buf BUF1 (N3347, N3329);
nand NAND3 (N3348, N3347, N2696, N1432);
not NOT1 (N3349, N3339);
and AND3 (N3350, N3324, N1384, N1746);
or OR2 (N3351, N3328, N3036);
and AND3 (N3352, N3351, N558, N371);
nor NOR4 (N3353, N3350, N1063, N610, N2734);
nand NAND3 (N3354, N3340, N680, N2367);
not NOT1 (N3355, N3353);
or OR3 (N3356, N3354, N1267, N1357);
nand NAND3 (N3357, N3336, N1114, N1518);
and AND3 (N3358, N3349, N577, N397);
xor XOR2 (N3359, N3344, N79);
or OR4 (N3360, N3355, N1116, N3024, N1534);
not NOT1 (N3361, N3357);
not NOT1 (N3362, N3348);
buf BUF1 (N3363, N3356);
xor XOR2 (N3364, N3346, N122);
xor XOR2 (N3365, N3360, N1299);
nor NOR2 (N3366, N3365, N1551);
or OR2 (N3367, N3337, N2063);
not NOT1 (N3368, N3362);
xor XOR2 (N3369, N3358, N1227);
buf BUF1 (N3370, N3369);
not NOT1 (N3371, N3366);
and AND2 (N3372, N3341, N238);
not NOT1 (N3373, N3359);
not NOT1 (N3374, N3370);
xor XOR2 (N3375, N3361, N2806);
nor NOR2 (N3376, N3375, N870);
and AND2 (N3377, N3376, N624);
nor NOR3 (N3378, N3371, N1450, N94);
buf BUF1 (N3379, N3363);
or OR3 (N3380, N3373, N1387, N1096);
nor NOR3 (N3381, N3367, N2738, N2151);
xor XOR2 (N3382, N3374, N1910);
and AND4 (N3383, N3380, N1736, N1342, N1249);
not NOT1 (N3384, N3368);
not NOT1 (N3385, N3377);
xor XOR2 (N3386, N3385, N896);
nand NAND2 (N3387, N3379, N2608);
xor XOR2 (N3388, N3383, N1239);
buf BUF1 (N3389, N3382);
buf BUF1 (N3390, N3389);
xor XOR2 (N3391, N3386, N2971);
not NOT1 (N3392, N3352);
not NOT1 (N3393, N3372);
not NOT1 (N3394, N3388);
buf BUF1 (N3395, N3364);
nand NAND3 (N3396, N3392, N1169, N713);
not NOT1 (N3397, N3381);
nand NAND4 (N3398, N3384, N281, N2405, N1693);
and AND3 (N3399, N3387, N1218, N225);
xor XOR2 (N3400, N3395, N941);
not NOT1 (N3401, N3396);
nand NAND4 (N3402, N3393, N439, N1610, N341);
xor XOR2 (N3403, N3401, N2542);
and AND2 (N3404, N3402, N1315);
nor NOR4 (N3405, N3390, N2974, N3006, N2580);
buf BUF1 (N3406, N3405);
nand NAND2 (N3407, N3398, N565);
not NOT1 (N3408, N3400);
nor NOR3 (N3409, N3397, N3377, N2793);
and AND3 (N3410, N3409, N453, N588);
buf BUF1 (N3411, N3391);
nand NAND3 (N3412, N3408, N3052, N1110);
or OR4 (N3413, N3394, N1126, N112, N420);
xor XOR2 (N3414, N3413, N2795);
not NOT1 (N3415, N3414);
xor XOR2 (N3416, N3403, N2993);
or OR4 (N3417, N3412, N21, N540, N575);
xor XOR2 (N3418, N3399, N3146);
nand NAND4 (N3419, N3407, N266, N392, N548);
xor XOR2 (N3420, N3415, N433);
not NOT1 (N3421, N3418);
xor XOR2 (N3422, N3419, N969);
and AND3 (N3423, N3420, N1484, N2001);
buf BUF1 (N3424, N3421);
and AND4 (N3425, N3406, N3268, N1370, N1013);
nor NOR4 (N3426, N3404, N416, N1465, N567);
xor XOR2 (N3427, N3378, N1164);
not NOT1 (N3428, N3425);
nor NOR2 (N3429, N3417, N1536);
nand NAND3 (N3430, N3428, N658, N1702);
not NOT1 (N3431, N3422);
and AND3 (N3432, N3416, N553, N3325);
xor XOR2 (N3433, N3410, N5);
buf BUF1 (N3434, N3432);
not NOT1 (N3435, N3423);
buf BUF1 (N3436, N3430);
not NOT1 (N3437, N3424);
nor NOR3 (N3438, N3426, N2152, N2754);
nand NAND4 (N3439, N3431, N834, N1331, N1642);
xor XOR2 (N3440, N3433, N1697);
xor XOR2 (N3441, N3438, N1161);
nand NAND2 (N3442, N3441, N1730);
or OR3 (N3443, N3429, N1724, N426);
or OR4 (N3444, N3411, N415, N1583, N980);
buf BUF1 (N3445, N3443);
not NOT1 (N3446, N3440);
buf BUF1 (N3447, N3434);
or OR4 (N3448, N3427, N1282, N3042, N2302);
and AND4 (N3449, N3444, N1692, N1694, N2312);
and AND4 (N3450, N3448, N1171, N1274, N728);
not NOT1 (N3451, N3435);
nand NAND2 (N3452, N3439, N563);
not NOT1 (N3453, N3445);
not NOT1 (N3454, N3451);
not NOT1 (N3455, N3442);
not NOT1 (N3456, N3455);
buf BUF1 (N3457, N3452);
or OR2 (N3458, N3456, N40);
not NOT1 (N3459, N3449);
and AND4 (N3460, N3453, N1176, N3388, N2708);
or OR4 (N3461, N3460, N2072, N1906, N2514);
xor XOR2 (N3462, N3447, N1299);
or OR4 (N3463, N3457, N287, N3027, N592);
xor XOR2 (N3464, N3463, N791);
nor NOR4 (N3465, N3436, N2189, N1505, N1826);
buf BUF1 (N3466, N3461);
not NOT1 (N3467, N3462);
xor XOR2 (N3468, N3446, N827);
nor NOR3 (N3469, N3454, N2628, N3148);
or OR3 (N3470, N3450, N2311, N2192);
buf BUF1 (N3471, N3465);
xor XOR2 (N3472, N3471, N1489);
xor XOR2 (N3473, N3437, N674);
and AND4 (N3474, N3458, N1711, N1292, N2822);
buf BUF1 (N3475, N3472);
buf BUF1 (N3476, N3467);
not NOT1 (N3477, N3470);
or OR4 (N3478, N3468, N2390, N2615, N2106);
buf BUF1 (N3479, N3464);
nand NAND2 (N3480, N3466, N261);
not NOT1 (N3481, N3477);
not NOT1 (N3482, N3474);
buf BUF1 (N3483, N3475);
buf BUF1 (N3484, N3480);
nand NAND3 (N3485, N3469, N1571, N3202);
and AND3 (N3486, N3481, N482, N12);
not NOT1 (N3487, N3483);
nor NOR3 (N3488, N3485, N496, N1394);
xor XOR2 (N3489, N3479, N3475);
and AND2 (N3490, N3476, N316);
and AND4 (N3491, N3484, N990, N200, N405);
nand NAND2 (N3492, N3487, N360);
and AND3 (N3493, N3489, N132, N220);
nand NAND4 (N3494, N3478, N2549, N2489, N3415);
and AND2 (N3495, N3486, N3328);
not NOT1 (N3496, N3459);
nor NOR3 (N3497, N3492, N1133, N1713);
and AND3 (N3498, N3488, N1902, N1742);
buf BUF1 (N3499, N3473);
xor XOR2 (N3500, N3490, N1946);
and AND3 (N3501, N3494, N688, N3092);
nor NOR2 (N3502, N3499, N212);
or OR2 (N3503, N3493, N2210);
xor XOR2 (N3504, N3482, N306);
xor XOR2 (N3505, N3498, N2640);
nor NOR4 (N3506, N3505, N2892, N1902, N3242);
or OR2 (N3507, N3503, N2665);
not NOT1 (N3508, N3502);
and AND2 (N3509, N3506, N1100);
xor XOR2 (N3510, N3496, N2983);
and AND2 (N3511, N3507, N3455);
xor XOR2 (N3512, N3509, N256);
buf BUF1 (N3513, N3508);
xor XOR2 (N3514, N3501, N2155);
nand NAND4 (N3515, N3497, N2737, N767, N2123);
not NOT1 (N3516, N3514);
nor NOR4 (N3517, N3515, N2448, N1501, N3427);
not NOT1 (N3518, N3510);
and AND3 (N3519, N3518, N2535, N476);
nand NAND4 (N3520, N3504, N2763, N2105, N2776);
nor NOR2 (N3521, N3520, N2750);
not NOT1 (N3522, N3500);
and AND2 (N3523, N3517, N798);
or OR2 (N3524, N3511, N2251);
not NOT1 (N3525, N3491);
not NOT1 (N3526, N3523);
nand NAND3 (N3527, N3522, N2973, N3389);
and AND3 (N3528, N3512, N1694, N2498);
or OR2 (N3529, N3528, N1894);
nand NAND3 (N3530, N3521, N3108, N888);
xor XOR2 (N3531, N3524, N730);
buf BUF1 (N3532, N3513);
nand NAND4 (N3533, N3525, N2330, N2386, N63);
nor NOR2 (N3534, N3495, N2499);
nor NOR2 (N3535, N3519, N1405);
or OR3 (N3536, N3530, N163, N2401);
and AND3 (N3537, N3533, N3276, N1257);
and AND3 (N3538, N3534, N2230, N1869);
nor NOR4 (N3539, N3527, N1131, N1, N33);
xor XOR2 (N3540, N3535, N2170);
and AND2 (N3541, N3532, N2278);
or OR4 (N3542, N3540, N2430, N2078, N1508);
not NOT1 (N3543, N3516);
nor NOR4 (N3544, N3538, N2257, N1461, N3430);
or OR4 (N3545, N3541, N2082, N74, N520);
buf BUF1 (N3546, N3542);
buf BUF1 (N3547, N3526);
not NOT1 (N3548, N3531);
nor NOR3 (N3549, N3539, N3080, N1888);
not NOT1 (N3550, N3529);
and AND4 (N3551, N3550, N1329, N2899, N241);
not NOT1 (N3552, N3549);
buf BUF1 (N3553, N3546);
buf BUF1 (N3554, N3545);
or OR4 (N3555, N3547, N3492, N2369, N1961);
or OR4 (N3556, N3537, N2368, N852, N3539);
or OR2 (N3557, N3544, N1559);
nor NOR3 (N3558, N3553, N360, N2859);
not NOT1 (N3559, N3556);
buf BUF1 (N3560, N3543);
nor NOR3 (N3561, N3554, N209, N3223);
buf BUF1 (N3562, N3551);
buf BUF1 (N3563, N3552);
or OR4 (N3564, N3555, N2938, N1948, N611);
and AND4 (N3565, N3536, N644, N3350, N1977);
and AND3 (N3566, N3558, N1323, N1411);
and AND4 (N3567, N3561, N300, N2771, N2635);
nor NOR2 (N3568, N3560, N288);
or OR2 (N3569, N3565, N650);
or OR3 (N3570, N3562, N1466, N3440);
and AND4 (N3571, N3566, N1074, N2292, N1626);
xor XOR2 (N3572, N3567, N2085);
or OR2 (N3573, N3564, N2318);
xor XOR2 (N3574, N3573, N1210);
nor NOR3 (N3575, N3548, N692, N661);
nor NOR2 (N3576, N3572, N1325);
not NOT1 (N3577, N3568);
nor NOR4 (N3578, N3569, N1923, N3200, N2416);
nor NOR3 (N3579, N3563, N747, N2487);
nand NAND4 (N3580, N3576, N1997, N2391, N1288);
xor XOR2 (N3581, N3578, N351);
buf BUF1 (N3582, N3575);
nand NAND2 (N3583, N3559, N3020);
xor XOR2 (N3584, N3571, N3115);
not NOT1 (N3585, N3570);
not NOT1 (N3586, N3557);
not NOT1 (N3587, N3574);
nor NOR2 (N3588, N3577, N3001);
or OR2 (N3589, N3588, N3303);
nand NAND3 (N3590, N3584, N3099, N2382);
and AND3 (N3591, N3582, N2627, N2279);
buf BUF1 (N3592, N3586);
nand NAND4 (N3593, N3579, N3162, N1133, N1321);
xor XOR2 (N3594, N3591, N1288);
buf BUF1 (N3595, N3580);
or OR3 (N3596, N3595, N1586, N1317);
and AND3 (N3597, N3583, N266, N1832);
nand NAND3 (N3598, N3594, N1639, N1818);
nor NOR3 (N3599, N3581, N3058, N3237);
buf BUF1 (N3600, N3589);
nand NAND3 (N3601, N3597, N1466, N2555);
nor NOR2 (N3602, N3593, N2672);
and AND4 (N3603, N3587, N1343, N3012, N3344);
buf BUF1 (N3604, N3600);
or OR3 (N3605, N3604, N3515, N2957);
not NOT1 (N3606, N3601);
or OR4 (N3607, N3596, N2177, N1799, N640);
xor XOR2 (N3608, N3599, N1197);
not NOT1 (N3609, N3608);
and AND2 (N3610, N3607, N884);
nand NAND3 (N3611, N3592, N2048, N2761);
xor XOR2 (N3612, N3598, N54);
or OR3 (N3613, N3606, N3560, N1380);
and AND4 (N3614, N3603, N2083, N2414, N1082);
buf BUF1 (N3615, N3613);
and AND2 (N3616, N3602, N3409);
not NOT1 (N3617, N3612);
not NOT1 (N3618, N3614);
not NOT1 (N3619, N3610);
not NOT1 (N3620, N3616);
nor NOR3 (N3621, N3618, N511, N2663);
nor NOR4 (N3622, N3619, N1261, N3559, N1786);
xor XOR2 (N3623, N3590, N2915);
or OR2 (N3624, N3623, N3174);
not NOT1 (N3625, N3622);
xor XOR2 (N3626, N3609, N989);
buf BUF1 (N3627, N3611);
nand NAND2 (N3628, N3627, N75);
nor NOR3 (N3629, N3626, N1136, N2681);
and AND3 (N3630, N3628, N1320, N2220);
nand NAND3 (N3631, N3617, N2442, N491);
nand NAND3 (N3632, N3621, N2018, N450);
nand NAND2 (N3633, N3605, N1054);
xor XOR2 (N3634, N3620, N1457);
xor XOR2 (N3635, N3629, N407);
and AND3 (N3636, N3633, N1447, N1990);
xor XOR2 (N3637, N3631, N555);
and AND2 (N3638, N3615, N1061);
nor NOR3 (N3639, N3635, N1891, N2818);
buf BUF1 (N3640, N3625);
nand NAND4 (N3641, N3634, N304, N2550, N3637);
xor XOR2 (N3642, N3076, N3499);
nand NAND3 (N3643, N3640, N116, N3327);
and AND4 (N3644, N3642, N980, N2267, N2858);
xor XOR2 (N3645, N3638, N2632);
or OR3 (N3646, N3641, N2198, N117);
or OR2 (N3647, N3585, N3460);
xor XOR2 (N3648, N3643, N1853);
and AND2 (N3649, N3648, N36);
xor XOR2 (N3650, N3646, N678);
buf BUF1 (N3651, N3645);
nand NAND4 (N3652, N3649, N65, N566, N74);
or OR4 (N3653, N3632, N3243, N2070, N2907);
xor XOR2 (N3654, N3636, N689);
xor XOR2 (N3655, N3652, N1953);
nand NAND2 (N3656, N3644, N690);
buf BUF1 (N3657, N3653);
nor NOR3 (N3658, N3624, N1669, N209);
xor XOR2 (N3659, N3656, N1862);
nor NOR4 (N3660, N3658, N645, N1223, N2137);
nor NOR3 (N3661, N3651, N666, N1695);
nand NAND4 (N3662, N3647, N5, N3190, N3047);
xor XOR2 (N3663, N3661, N2023);
xor XOR2 (N3664, N3657, N3181);
or OR3 (N3665, N3664, N2580, N3524);
not NOT1 (N3666, N3663);
buf BUF1 (N3667, N3630);
nor NOR4 (N3668, N3666, N3629, N3304, N2775);
and AND2 (N3669, N3659, N2636);
and AND4 (N3670, N3667, N3300, N2051, N3068);
not NOT1 (N3671, N3660);
buf BUF1 (N3672, N3655);
nor NOR3 (N3673, N3669, N3133, N1225);
not NOT1 (N3674, N3671);
xor XOR2 (N3675, N3673, N2317);
nand NAND3 (N3676, N3639, N1276, N3305);
not NOT1 (N3677, N3676);
nand NAND2 (N3678, N3665, N922);
not NOT1 (N3679, N3650);
nand NAND3 (N3680, N3654, N770, N811);
buf BUF1 (N3681, N3662);
buf BUF1 (N3682, N3668);
and AND4 (N3683, N3675, N1675, N259, N2422);
or OR3 (N3684, N3679, N963, N281);
buf BUF1 (N3685, N3672);
not NOT1 (N3686, N3683);
nor NOR2 (N3687, N3677, N1489);
xor XOR2 (N3688, N3681, N119);
not NOT1 (N3689, N3688);
nor NOR4 (N3690, N3687, N398, N554, N49);
buf BUF1 (N3691, N3674);
and AND4 (N3692, N3684, N3271, N2485, N605);
or OR2 (N3693, N3692, N2831);
or OR3 (N3694, N3690, N693, N543);
nor NOR4 (N3695, N3678, N474, N926, N3311);
buf BUF1 (N3696, N3689);
nor NOR4 (N3697, N3685, N1314, N3467, N266);
not NOT1 (N3698, N3691);
nor NOR2 (N3699, N3670, N2246);
buf BUF1 (N3700, N3699);
nor NOR2 (N3701, N3698, N1687);
and AND3 (N3702, N3697, N108, N1266);
buf BUF1 (N3703, N3700);
nor NOR3 (N3704, N3702, N3499, N2902);
not NOT1 (N3705, N3682);
nor NOR4 (N3706, N3703, N2047, N2143, N1603);
not NOT1 (N3707, N3701);
nand NAND3 (N3708, N3693, N1264, N1349);
nor NOR2 (N3709, N3705, N3095);
not NOT1 (N3710, N3706);
nand NAND3 (N3711, N3707, N3269, N1103);
nand NAND2 (N3712, N3686, N2857);
and AND3 (N3713, N3711, N1313, N3126);
nor NOR3 (N3714, N3713, N992, N1290);
or OR3 (N3715, N3710, N3451, N2764);
not NOT1 (N3716, N3680);
xor XOR2 (N3717, N3709, N3292);
nor NOR2 (N3718, N3717, N2427);
and AND2 (N3719, N3714, N2910);
or OR3 (N3720, N3694, N2718, N3643);
not NOT1 (N3721, N3718);
nand NAND3 (N3722, N3708, N583, N1511);
not NOT1 (N3723, N3720);
nand NAND2 (N3724, N3716, N3481);
nand NAND3 (N3725, N3696, N663, N2065);
and AND3 (N3726, N3721, N2985, N2030);
nor NOR4 (N3727, N3715, N3655, N2538, N3208);
xor XOR2 (N3728, N3727, N2821);
nand NAND4 (N3729, N3704, N591, N896, N3672);
buf BUF1 (N3730, N3719);
nand NAND4 (N3731, N3726, N1760, N214, N2383);
buf BUF1 (N3732, N3722);
xor XOR2 (N3733, N3723, N1789);
buf BUF1 (N3734, N3729);
nor NOR4 (N3735, N3712, N1780, N2584, N1507);
nor NOR2 (N3736, N3731, N2690);
or OR4 (N3737, N3724, N1570, N1892, N1834);
or OR3 (N3738, N3732, N2361, N2840);
xor XOR2 (N3739, N3695, N2071);
not NOT1 (N3740, N3738);
or OR2 (N3741, N3735, N1042);
or OR3 (N3742, N3728, N1249, N724);
or OR3 (N3743, N3736, N3689, N3675);
or OR2 (N3744, N3740, N474);
not NOT1 (N3745, N3741);
nor NOR3 (N3746, N3744, N3642, N1108);
buf BUF1 (N3747, N3725);
and AND2 (N3748, N3739, N1136);
nand NAND2 (N3749, N3742, N2094);
not NOT1 (N3750, N3733);
and AND2 (N3751, N3745, N1909);
nor NOR2 (N3752, N3750, N2187);
buf BUF1 (N3753, N3747);
or OR4 (N3754, N3753, N3480, N1012, N3560);
and AND3 (N3755, N3730, N3411, N3541);
xor XOR2 (N3756, N3743, N2689);
or OR3 (N3757, N3734, N2456, N2712);
xor XOR2 (N3758, N3756, N3519);
nor NOR3 (N3759, N3749, N1514, N346);
not NOT1 (N3760, N3752);
and AND2 (N3761, N3759, N2161);
xor XOR2 (N3762, N3760, N3668);
and AND4 (N3763, N3761, N1229, N605, N735);
not NOT1 (N3764, N3746);
and AND2 (N3765, N3762, N1147);
buf BUF1 (N3766, N3755);
or OR3 (N3767, N3764, N1036, N456);
and AND3 (N3768, N3751, N574, N602);
buf BUF1 (N3769, N3754);
not NOT1 (N3770, N3748);
and AND4 (N3771, N3758, N3405, N1281, N1760);
xor XOR2 (N3772, N3763, N1879);
buf BUF1 (N3773, N3737);
buf BUF1 (N3774, N3773);
xor XOR2 (N3775, N3774, N1034);
nand NAND3 (N3776, N3769, N1517, N1623);
not NOT1 (N3777, N3766);
nor NOR3 (N3778, N3777, N567, N2237);
and AND2 (N3779, N3765, N61);
nor NOR4 (N3780, N3767, N1105, N1763, N613);
not NOT1 (N3781, N3771);
xor XOR2 (N3782, N3770, N693);
not NOT1 (N3783, N3776);
buf BUF1 (N3784, N3779);
nor NOR3 (N3785, N3780, N1337, N351);
or OR4 (N3786, N3775, N105, N1747, N2017);
nor NOR2 (N3787, N3785, N3552);
and AND3 (N3788, N3782, N2692, N343);
buf BUF1 (N3789, N3784);
buf BUF1 (N3790, N3783);
or OR4 (N3791, N3757, N3440, N1230, N1986);
or OR4 (N3792, N3768, N3419, N1932, N1885);
not NOT1 (N3793, N3789);
not NOT1 (N3794, N3786);
buf BUF1 (N3795, N3787);
nor NOR4 (N3796, N3795, N2474, N1274, N2706);
and AND4 (N3797, N3778, N3171, N237, N2837);
xor XOR2 (N3798, N3781, N2952);
xor XOR2 (N3799, N3797, N2993);
buf BUF1 (N3800, N3790);
nand NAND2 (N3801, N3798, N1701);
xor XOR2 (N3802, N3788, N897);
buf BUF1 (N3803, N3794);
buf BUF1 (N3804, N3800);
xor XOR2 (N3805, N3804, N105);
or OR3 (N3806, N3791, N1097, N2165);
not NOT1 (N3807, N3792);
nor NOR4 (N3808, N3805, N2104, N23, N2263);
nor NOR2 (N3809, N3806, N1390);
or OR2 (N3810, N3803, N925);
nand NAND2 (N3811, N3799, N3490);
nand NAND4 (N3812, N3796, N834, N2272, N1243);
nand NAND3 (N3813, N3807, N1085, N3175);
or OR3 (N3814, N3802, N3004, N1040);
nor NOR3 (N3815, N3801, N3379, N314);
xor XOR2 (N3816, N3813, N540);
buf BUF1 (N3817, N3812);
nand NAND4 (N3818, N3811, N3400, N845, N1330);
buf BUF1 (N3819, N3817);
buf BUF1 (N3820, N3793);
xor XOR2 (N3821, N3772, N1461);
buf BUF1 (N3822, N3809);
buf BUF1 (N3823, N3810);
buf BUF1 (N3824, N3815);
buf BUF1 (N3825, N3818);
xor XOR2 (N3826, N3819, N771);
not NOT1 (N3827, N3823);
buf BUF1 (N3828, N3816);
xor XOR2 (N3829, N3814, N2390);
and AND2 (N3830, N3826, N76);
or OR3 (N3831, N3821, N1811, N2916);
not NOT1 (N3832, N3822);
nor NOR3 (N3833, N3825, N3026, N1925);
buf BUF1 (N3834, N3820);
and AND3 (N3835, N3828, N612, N1223);
and AND2 (N3836, N3827, N3504);
not NOT1 (N3837, N3834);
buf BUF1 (N3838, N3835);
buf BUF1 (N3839, N3830);
xor XOR2 (N3840, N3832, N944);
nor NOR4 (N3841, N3808, N1843, N945, N930);
nor NOR2 (N3842, N3840, N2976);
nor NOR2 (N3843, N3841, N2789);
and AND2 (N3844, N3839, N2210);
and AND2 (N3845, N3833, N2326);
not NOT1 (N3846, N3836);
xor XOR2 (N3847, N3837, N1002);
or OR3 (N3848, N3824, N2492, N3303);
nor NOR3 (N3849, N3848, N1758, N3678);
buf BUF1 (N3850, N3845);
nor NOR2 (N3851, N3846, N2632);
and AND4 (N3852, N3850, N2829, N1037, N121);
nand NAND4 (N3853, N3847, N335, N2498, N519);
not NOT1 (N3854, N3838);
and AND3 (N3855, N3854, N883, N2412);
xor XOR2 (N3856, N3855, N1758);
not NOT1 (N3857, N3853);
and AND2 (N3858, N3831, N1902);
or OR4 (N3859, N3851, N527, N3591, N1502);
not NOT1 (N3860, N3842);
not NOT1 (N3861, N3857);
and AND3 (N3862, N3860, N706, N1238);
nand NAND4 (N3863, N3844, N49, N1591, N3327);
nor NOR4 (N3864, N3861, N3435, N1227, N729);
nor NOR2 (N3865, N3852, N1696);
not NOT1 (N3866, N3859);
nand NAND4 (N3867, N3863, N2518, N141, N1395);
and AND2 (N3868, N3867, N2905);
nor NOR3 (N3869, N3849, N2184, N3594);
not NOT1 (N3870, N3865);
nor NOR3 (N3871, N3870, N410, N274);
and AND2 (N3872, N3858, N3678);
xor XOR2 (N3873, N3856, N2498);
buf BUF1 (N3874, N3864);
or OR4 (N3875, N3829, N2178, N3030, N3710);
nor NOR3 (N3876, N3868, N321, N2035);
xor XOR2 (N3877, N3872, N1545);
nand NAND3 (N3878, N3874, N390, N3757);
and AND4 (N3879, N3869, N1002, N958, N3333);
and AND3 (N3880, N3866, N3058, N2924);
nor NOR2 (N3881, N3875, N2813);
nand NAND4 (N3882, N3880, N2893, N1567, N736);
nor NOR2 (N3883, N3878, N2531);
nand NAND2 (N3884, N3876, N2084);
nand NAND3 (N3885, N3862, N211, N1135);
buf BUF1 (N3886, N3877);
nor NOR4 (N3887, N3884, N2487, N3601, N3619);
and AND2 (N3888, N3886, N2077);
buf BUF1 (N3889, N3883);
and AND4 (N3890, N3889, N1890, N3536, N2789);
not NOT1 (N3891, N3885);
or OR4 (N3892, N3888, N94, N2490, N903);
nand NAND4 (N3893, N3871, N1616, N2753, N504);
nor NOR4 (N3894, N3881, N1241, N926, N474);
or OR3 (N3895, N3879, N1677, N1699);
nand NAND4 (N3896, N3882, N2595, N3585, N2089);
buf BUF1 (N3897, N3890);
not NOT1 (N3898, N3891);
and AND2 (N3899, N3843, N1123);
and AND3 (N3900, N3897, N2871, N2260);
not NOT1 (N3901, N3899);
not NOT1 (N3902, N3895);
and AND3 (N3903, N3902, N2024, N1324);
buf BUF1 (N3904, N3892);
and AND2 (N3905, N3903, N1938);
nand NAND4 (N3906, N3893, N1131, N1270, N2201);
xor XOR2 (N3907, N3901, N2357);
buf BUF1 (N3908, N3900);
or OR4 (N3909, N3908, N3497, N3646, N2965);
nand NAND4 (N3910, N3904, N507, N2430, N2559);
buf BUF1 (N3911, N3894);
or OR4 (N3912, N3898, N3068, N2204, N1356);
and AND3 (N3913, N3873, N1021, N3854);
nor NOR3 (N3914, N3905, N1477, N3861);
nand NAND2 (N3915, N3907, N2544);
and AND4 (N3916, N3910, N1472, N3493, N3385);
nor NOR4 (N3917, N3914, N3898, N2050, N3262);
and AND4 (N3918, N3906, N3823, N2591, N1688);
nor NOR3 (N3919, N3917, N1722, N683);
nand NAND4 (N3920, N3909, N3343, N562, N1797);
nand NAND2 (N3921, N3913, N1699);
buf BUF1 (N3922, N3920);
or OR3 (N3923, N3912, N1714, N3664);
nor NOR3 (N3924, N3919, N3291, N2030);
and AND3 (N3925, N3916, N2552, N391);
nor NOR4 (N3926, N3918, N1041, N499, N2175);
xor XOR2 (N3927, N3915, N3611);
not NOT1 (N3928, N3896);
buf BUF1 (N3929, N3887);
nor NOR4 (N3930, N3922, N2907, N1532, N450);
nand NAND2 (N3931, N3921, N3819);
buf BUF1 (N3932, N3929);
and AND4 (N3933, N3924, N695, N1663, N1463);
nand NAND3 (N3934, N3931, N1862, N542);
buf BUF1 (N3935, N3930);
not NOT1 (N3936, N3928);
or OR3 (N3937, N3935, N2602, N82);
nor NOR4 (N3938, N3936, N3837, N3022, N628);
nand NAND3 (N3939, N3938, N2916, N1938);
and AND3 (N3940, N3939, N1562, N2839);
xor XOR2 (N3941, N3932, N3156);
nor NOR3 (N3942, N3925, N3218, N3526);
nor NOR3 (N3943, N3923, N1512, N1347);
xor XOR2 (N3944, N3927, N1955);
or OR3 (N3945, N3943, N2210, N6);
nor NOR4 (N3946, N3942, N74, N3216, N3666);
and AND3 (N3947, N3926, N2, N772);
xor XOR2 (N3948, N3937, N3339);
not NOT1 (N3949, N3941);
or OR4 (N3950, N3911, N191, N2617, N3571);
xor XOR2 (N3951, N3948, N3764);
nand NAND3 (N3952, N3945, N409, N1412);
buf BUF1 (N3953, N3952);
or OR3 (N3954, N3950, N3019, N3488);
nor NOR2 (N3955, N3954, N3855);
xor XOR2 (N3956, N3953, N3669);
buf BUF1 (N3957, N3934);
buf BUF1 (N3958, N3956);
and AND3 (N3959, N3957, N2465, N2273);
or OR3 (N3960, N3955, N1145, N242);
xor XOR2 (N3961, N3960, N3207);
nand NAND2 (N3962, N3961, N1768);
nor NOR3 (N3963, N3946, N700, N3769);
and AND3 (N3964, N3944, N1958, N1646);
nor NOR4 (N3965, N3951, N3695, N3466, N2514);
nand NAND4 (N3966, N3964, N3110, N2979, N219);
buf BUF1 (N3967, N3933);
not NOT1 (N3968, N3958);
nor NOR4 (N3969, N3965, N3250, N1707, N1796);
buf BUF1 (N3970, N3949);
not NOT1 (N3971, N3962);
nor NOR3 (N3972, N3963, N1605, N2630);
buf BUF1 (N3973, N3959);
xor XOR2 (N3974, N3972, N2464);
not NOT1 (N3975, N3969);
nand NAND4 (N3976, N3966, N3692, N2041, N3327);
nor NOR2 (N3977, N3967, N2706);
nand NAND4 (N3978, N3968, N1416, N826, N1589);
xor XOR2 (N3979, N3976, N2140);
buf BUF1 (N3980, N3947);
not NOT1 (N3981, N3979);
not NOT1 (N3982, N3980);
nor NOR3 (N3983, N3940, N3265, N2182);
buf BUF1 (N3984, N3982);
buf BUF1 (N3985, N3978);
not NOT1 (N3986, N3971);
or OR4 (N3987, N3974, N2987, N1165, N1236);
xor XOR2 (N3988, N3984, N93);
xor XOR2 (N3989, N3970, N3858);
or OR2 (N3990, N3988, N2320);
and AND4 (N3991, N3981, N313, N264, N3933);
nand NAND2 (N3992, N3991, N2965);
and AND4 (N3993, N3983, N2614, N1958, N1777);
xor XOR2 (N3994, N3985, N1212);
buf BUF1 (N3995, N3987);
not NOT1 (N3996, N3975);
or OR3 (N3997, N3977, N3795, N2414);
or OR4 (N3998, N3990, N1491, N94, N2553);
nor NOR3 (N3999, N3973, N3004, N699);
xor XOR2 (N4000, N3993, N2360);
buf BUF1 (N4001, N3995);
nand NAND3 (N4002, N4001, N566, N3717);
not NOT1 (N4003, N3999);
nor NOR4 (N4004, N4000, N461, N1352, N3829);
xor XOR2 (N4005, N3997, N3941);
or OR4 (N4006, N3996, N1548, N1342, N3846);
nor NOR3 (N4007, N3989, N3192, N3269);
not NOT1 (N4008, N3986);
nand NAND3 (N4009, N3998, N555, N3856);
nor NOR4 (N4010, N4006, N1530, N1024, N1412);
xor XOR2 (N4011, N3994, N2587);
not NOT1 (N4012, N4010);
nand NAND4 (N4013, N4002, N3097, N1363, N1411);
xor XOR2 (N4014, N3992, N1645);
or OR4 (N4015, N4007, N3281, N560, N1528);
nand NAND4 (N4016, N4015, N3603, N3978, N2506);
not NOT1 (N4017, N4009);
buf BUF1 (N4018, N4014);
or OR2 (N4019, N4008, N1574);
and AND4 (N4020, N4018, N2975, N989, N2391);
or OR3 (N4021, N4012, N897, N1770);
nand NAND4 (N4022, N4016, N3683, N3530, N3868);
and AND3 (N4023, N4013, N2342, N2499);
nor NOR2 (N4024, N4020, N2110);
endmodule