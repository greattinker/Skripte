// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N16009,N16018,N16017,N16014,N16008,N16012,N16015,N16019,N15995,N16020;

nor NOR4 (N21, N2, N15, N14, N12);
not NOT1 (N22, N8);
nor NOR2 (N23, N19, N11);
and AND3 (N24, N5, N12, N19);
or OR4 (N25, N1, N3, N4, N19);
and AND3 (N26, N16, N7, N22);
xor XOR2 (N27, N6, N22);
nor NOR4 (N28, N3, N24, N9, N25);
or OR2 (N29, N4, N19);
nand NAND2 (N30, N15, N10);
nor NOR2 (N31, N8, N30);
or OR3 (N32, N4, N23, N26);
nand NAND4 (N33, N13, N26, N9, N32);
nand NAND4 (N34, N16, N5, N10, N12);
nand NAND3 (N35, N1, N3, N11);
and AND3 (N36, N2, N13, N33);
buf BUF1 (N37, N7);
not NOT1 (N38, N33);
buf BUF1 (N39, N28);
xor XOR2 (N40, N21, N19);
not NOT1 (N41, N40);
nand NAND4 (N42, N27, N31, N19, N16);
nor NOR4 (N43, N35, N24, N19, N7);
or OR2 (N44, N6, N21);
nor NOR4 (N45, N29, N27, N41, N2);
xor XOR2 (N46, N24, N20);
xor XOR2 (N47, N46, N40);
nor NOR2 (N48, N36, N33);
not NOT1 (N49, N44);
xor XOR2 (N50, N43, N5);
or OR3 (N51, N45, N32, N9);
not NOT1 (N52, N37);
and AND2 (N53, N47, N6);
nand NAND3 (N54, N52, N26, N16);
nor NOR4 (N55, N39, N4, N53, N6);
nor NOR3 (N56, N46, N47, N8);
xor XOR2 (N57, N51, N50);
nand NAND2 (N58, N34, N4);
not NOT1 (N59, N19);
nand NAND2 (N60, N55, N4);
not NOT1 (N61, N42);
nand NAND2 (N62, N59, N20);
xor XOR2 (N63, N60, N39);
xor XOR2 (N64, N63, N31);
nand NAND4 (N65, N48, N25, N28, N60);
not NOT1 (N66, N61);
buf BUF1 (N67, N65);
and AND2 (N68, N67, N58);
and AND3 (N69, N10, N58, N11);
nor NOR2 (N70, N56, N35);
and AND3 (N71, N70, N61, N26);
or OR2 (N72, N49, N22);
or OR3 (N73, N38, N56, N19);
nand NAND3 (N74, N66, N72, N46);
buf BUF1 (N75, N20);
buf BUF1 (N76, N68);
and AND3 (N77, N54, N34, N40);
buf BUF1 (N78, N69);
nand NAND2 (N79, N71, N71);
buf BUF1 (N80, N75);
xor XOR2 (N81, N62, N30);
buf BUF1 (N82, N81);
not NOT1 (N83, N79);
nand NAND4 (N84, N76, N45, N82, N71);
nand NAND2 (N85, N83, N82);
nor NOR3 (N86, N52, N47, N35);
and AND4 (N87, N73, N37, N19, N10);
not NOT1 (N88, N87);
xor XOR2 (N89, N88, N84);
and AND3 (N90, N33, N17, N49);
buf BUF1 (N91, N85);
xor XOR2 (N92, N64, N65);
not NOT1 (N93, N78);
xor XOR2 (N94, N77, N25);
buf BUF1 (N95, N90);
and AND4 (N96, N95, N47, N75, N54);
nor NOR3 (N97, N89, N64, N58);
nor NOR2 (N98, N91, N52);
not NOT1 (N99, N98);
nor NOR2 (N100, N99, N31);
xor XOR2 (N101, N97, N36);
not NOT1 (N102, N57);
nand NAND3 (N103, N96, N79, N53);
not NOT1 (N104, N94);
nand NAND3 (N105, N92, N42, N3);
nand NAND2 (N106, N102, N46);
not NOT1 (N107, N74);
not NOT1 (N108, N86);
nor NOR3 (N109, N108, N16, N67);
or OR2 (N110, N104, N57);
or OR3 (N111, N110, N28, N67);
not NOT1 (N112, N100);
and AND3 (N113, N93, N111, N96);
nand NAND4 (N114, N26, N37, N53, N42);
buf BUF1 (N115, N103);
nand NAND3 (N116, N112, N105, N88);
xor XOR2 (N117, N13, N83);
xor XOR2 (N118, N101, N79);
or OR3 (N119, N107, N112, N104);
buf BUF1 (N120, N80);
and AND3 (N121, N119, N41, N34);
xor XOR2 (N122, N116, N117);
nand NAND4 (N123, N13, N47, N25, N112);
nor NOR4 (N124, N120, N42, N86, N79);
nor NOR4 (N125, N109, N124, N97, N116);
nor NOR4 (N126, N8, N65, N25, N20);
or OR3 (N127, N125, N106, N24);
nand NAND3 (N128, N35, N25, N13);
not NOT1 (N129, N123);
xor XOR2 (N130, N128, N22);
or OR2 (N131, N126, N29);
not NOT1 (N132, N130);
nand NAND3 (N133, N115, N93, N37);
and AND4 (N134, N127, N5, N101, N59);
xor XOR2 (N135, N133, N127);
or OR4 (N136, N129, N108, N82, N70);
nand NAND2 (N137, N121, N119);
xor XOR2 (N138, N122, N67);
not NOT1 (N139, N132);
buf BUF1 (N140, N114);
not NOT1 (N141, N131);
nor NOR3 (N142, N118, N16, N122);
nor NOR2 (N143, N113, N142);
nand NAND4 (N144, N115, N107, N141, N6);
or OR4 (N145, N43, N40, N19, N2);
nand NAND4 (N146, N136, N18, N139, N116);
or OR2 (N147, N143, N55);
and AND2 (N148, N71, N129);
nor NOR2 (N149, N146, N126);
not NOT1 (N150, N137);
or OR4 (N151, N145, N81, N26, N133);
not NOT1 (N152, N149);
nand NAND3 (N153, N144, N93, N129);
or OR4 (N154, N140, N72, N84, N76);
xor XOR2 (N155, N151, N8);
nand NAND2 (N156, N153, N147);
and AND2 (N157, N142, N42);
xor XOR2 (N158, N154, N138);
not NOT1 (N159, N112);
nor NOR3 (N160, N159, N31, N12);
not NOT1 (N161, N150);
and AND4 (N162, N156, N108, N48, N41);
not NOT1 (N163, N155);
or OR3 (N164, N148, N116, N84);
not NOT1 (N165, N162);
or OR3 (N166, N163, N23, N111);
buf BUF1 (N167, N161);
nor NOR4 (N168, N166, N46, N164, N71);
nand NAND4 (N169, N2, N142, N24, N127);
buf BUF1 (N170, N160);
xor XOR2 (N171, N157, N1);
or OR2 (N172, N168, N64);
buf BUF1 (N173, N172);
not NOT1 (N174, N173);
xor XOR2 (N175, N135, N54);
buf BUF1 (N176, N171);
nand NAND2 (N177, N170, N2);
xor XOR2 (N178, N177, N136);
buf BUF1 (N179, N169);
nand NAND3 (N180, N174, N9, N14);
nand NAND3 (N181, N152, N105, N166);
and AND4 (N182, N165, N108, N5, N115);
nand NAND2 (N183, N182, N132);
xor XOR2 (N184, N158, N99);
and AND4 (N185, N176, N117, N29, N179);
and AND3 (N186, N73, N72, N73);
xor XOR2 (N187, N180, N138);
and AND4 (N188, N187, N171, N42, N111);
nor NOR4 (N189, N134, N61, N54, N147);
nor NOR4 (N190, N178, N130, N44, N150);
buf BUF1 (N191, N186);
xor XOR2 (N192, N190, N95);
and AND4 (N193, N192, N152, N98, N125);
nand NAND3 (N194, N184, N183, N119);
not NOT1 (N195, N132);
not NOT1 (N196, N175);
nor NOR2 (N197, N188, N47);
nor NOR4 (N198, N193, N115, N5, N155);
buf BUF1 (N199, N191);
nor NOR3 (N200, N196, N40, N22);
nand NAND3 (N201, N199, N83, N120);
buf BUF1 (N202, N200);
and AND3 (N203, N198, N133, N46);
nor NOR3 (N204, N194, N135, N37);
not NOT1 (N205, N181);
not NOT1 (N206, N205);
or OR3 (N207, N185, N62, N69);
xor XOR2 (N208, N203, N44);
buf BUF1 (N209, N197);
nor NOR4 (N210, N167, N9, N59, N183);
not NOT1 (N211, N209);
nand NAND2 (N212, N206, N97);
buf BUF1 (N213, N202);
xor XOR2 (N214, N211, N52);
or OR2 (N215, N210, N107);
not NOT1 (N216, N195);
buf BUF1 (N217, N207);
nor NOR2 (N218, N217, N145);
xor XOR2 (N219, N216, N128);
nor NOR2 (N220, N201, N207);
nand NAND4 (N221, N220, N205, N162, N190);
buf BUF1 (N222, N214);
nor NOR2 (N223, N204, N87);
buf BUF1 (N224, N219);
and AND3 (N225, N189, N72, N102);
nor NOR4 (N226, N212, N73, N195, N94);
xor XOR2 (N227, N223, N183);
and AND3 (N228, N208, N113, N171);
not NOT1 (N229, N225);
not NOT1 (N230, N228);
not NOT1 (N231, N227);
xor XOR2 (N232, N226, N7);
xor XOR2 (N233, N230, N10);
not NOT1 (N234, N231);
buf BUF1 (N235, N213);
buf BUF1 (N236, N215);
nor NOR3 (N237, N222, N196, N85);
and AND3 (N238, N232, N107, N208);
nor NOR4 (N239, N234, N41, N124, N16);
nor NOR3 (N240, N218, N11, N58);
or OR4 (N241, N240, N234, N177, N169);
not NOT1 (N242, N237);
and AND4 (N243, N233, N233, N192, N163);
xor XOR2 (N244, N236, N3);
nand NAND2 (N245, N224, N51);
buf BUF1 (N246, N241);
or OR2 (N247, N239, N210);
nand NAND3 (N248, N242, N114, N72);
and AND4 (N249, N235, N38, N34, N153);
xor XOR2 (N250, N246, N105);
and AND2 (N251, N247, N239);
not NOT1 (N252, N251);
buf BUF1 (N253, N229);
or OR4 (N254, N249, N51, N234, N127);
or OR4 (N255, N248, N224, N244, N149);
or OR3 (N256, N2, N86, N147);
and AND2 (N257, N243, N66);
xor XOR2 (N258, N221, N82);
nor NOR3 (N259, N252, N40, N144);
not NOT1 (N260, N245);
nand NAND4 (N261, N258, N245, N88, N155);
nor NOR3 (N262, N260, N42, N143);
or OR3 (N263, N254, N183, N66);
not NOT1 (N264, N263);
nor NOR4 (N265, N255, N54, N86, N169);
xor XOR2 (N266, N256, N22);
not NOT1 (N267, N257);
nand NAND4 (N268, N238, N149, N201, N251);
not NOT1 (N269, N267);
buf BUF1 (N270, N264);
or OR2 (N271, N266, N101);
not NOT1 (N272, N271);
not NOT1 (N273, N253);
buf BUF1 (N274, N250);
buf BUF1 (N275, N269);
nand NAND4 (N276, N272, N18, N186, N50);
and AND3 (N277, N268, N180, N125);
or OR4 (N278, N277, N159, N225, N127);
xor XOR2 (N279, N274, N193);
nor NOR4 (N280, N279, N81, N28, N83);
xor XOR2 (N281, N273, N113);
or OR3 (N282, N270, N118, N209);
nand NAND3 (N283, N259, N141, N129);
and AND3 (N284, N261, N183, N199);
buf BUF1 (N285, N282);
or OR2 (N286, N285, N147);
xor XOR2 (N287, N284, N121);
xor XOR2 (N288, N278, N97);
or OR3 (N289, N276, N160, N144);
and AND3 (N290, N281, N289, N254);
nor NOR4 (N291, N242, N95, N80, N170);
xor XOR2 (N292, N265, N272);
nand NAND4 (N293, N288, N233, N79, N183);
buf BUF1 (N294, N283);
or OR2 (N295, N291, N198);
nor NOR2 (N296, N290, N238);
not NOT1 (N297, N293);
buf BUF1 (N298, N296);
nand NAND2 (N299, N298, N276);
or OR4 (N300, N299, N224, N122, N12);
buf BUF1 (N301, N275);
xor XOR2 (N302, N294, N183);
xor XOR2 (N303, N301, N18);
nor NOR3 (N304, N280, N123, N117);
or OR2 (N305, N287, N222);
nor NOR3 (N306, N302, N124, N26);
xor XOR2 (N307, N262, N32);
or OR2 (N308, N305, N163);
or OR4 (N309, N308, N193, N68, N97);
nor NOR2 (N310, N306, N239);
xor XOR2 (N311, N286, N239);
or OR2 (N312, N307, N85);
nand NAND2 (N313, N297, N114);
nand NAND4 (N314, N313, N305, N292, N226);
or OR4 (N315, N254, N136, N249, N261);
xor XOR2 (N316, N309, N72);
or OR3 (N317, N312, N163, N176);
not NOT1 (N318, N303);
nand NAND3 (N319, N310, N266, N173);
nor NOR3 (N320, N295, N167, N187);
xor XOR2 (N321, N317, N210);
and AND3 (N322, N314, N164, N243);
nor NOR2 (N323, N319, N298);
nor NOR2 (N324, N318, N300);
or OR3 (N325, N89, N39, N101);
or OR4 (N326, N321, N158, N263, N35);
nand NAND4 (N327, N315, N271, N298, N261);
buf BUF1 (N328, N327);
nor NOR3 (N329, N328, N201, N55);
or OR3 (N330, N324, N21, N89);
not NOT1 (N331, N311);
not NOT1 (N332, N330);
nand NAND2 (N333, N320, N248);
buf BUF1 (N334, N322);
not NOT1 (N335, N334);
nand NAND2 (N336, N325, N194);
or OR3 (N337, N316, N277, N64);
not NOT1 (N338, N336);
xor XOR2 (N339, N304, N113);
or OR2 (N340, N332, N164);
nor NOR2 (N341, N339, N180);
buf BUF1 (N342, N323);
nor NOR3 (N343, N337, N131, N248);
xor XOR2 (N344, N329, N277);
or OR3 (N345, N335, N30, N85);
and AND3 (N346, N342, N57, N117);
xor XOR2 (N347, N345, N120);
nor NOR3 (N348, N326, N105, N36);
nand NAND3 (N349, N343, N213, N307);
not NOT1 (N350, N349);
nand NAND3 (N351, N348, N225, N246);
nor NOR4 (N352, N351, N136, N65, N306);
not NOT1 (N353, N352);
or OR3 (N354, N331, N164, N10);
not NOT1 (N355, N354);
nor NOR4 (N356, N340, N123, N54, N26);
and AND4 (N357, N338, N120, N59, N134);
nand NAND3 (N358, N355, N183, N67);
nor NOR4 (N359, N356, N82, N27, N110);
nand NAND2 (N360, N357, N37);
buf BUF1 (N361, N360);
or OR2 (N362, N341, N203);
not NOT1 (N363, N350);
nor NOR4 (N364, N347, N234, N114, N338);
nor NOR4 (N365, N362, N332, N265, N190);
buf BUF1 (N366, N346);
nor NOR3 (N367, N361, N272, N39);
buf BUF1 (N368, N365);
xor XOR2 (N369, N367, N284);
nor NOR3 (N370, N353, N238, N258);
nand NAND2 (N371, N369, N278);
or OR4 (N372, N358, N169, N366, N140);
and AND4 (N373, N133, N299, N225, N145);
nand NAND2 (N374, N333, N285);
xor XOR2 (N375, N370, N98);
buf BUF1 (N376, N364);
not NOT1 (N377, N374);
xor XOR2 (N378, N373, N74);
and AND2 (N379, N377, N23);
or OR3 (N380, N379, N78, N324);
not NOT1 (N381, N380);
nand NAND3 (N382, N372, N346, N370);
buf BUF1 (N383, N371);
nor NOR3 (N384, N382, N92, N182);
nand NAND3 (N385, N375, N280, N218);
and AND2 (N386, N344, N81);
xor XOR2 (N387, N383, N205);
buf BUF1 (N388, N363);
or OR2 (N389, N381, N379);
or OR3 (N390, N385, N256, N217);
or OR4 (N391, N388, N85, N166, N338);
not NOT1 (N392, N384);
not NOT1 (N393, N386);
buf BUF1 (N394, N378);
and AND3 (N395, N394, N186, N385);
or OR3 (N396, N390, N197, N225);
nor NOR3 (N397, N395, N193, N104);
nor NOR4 (N398, N397, N381, N240, N20);
nor NOR3 (N399, N392, N176, N275);
buf BUF1 (N400, N376);
buf BUF1 (N401, N396);
buf BUF1 (N402, N391);
and AND3 (N403, N402, N238, N365);
not NOT1 (N404, N403);
nor NOR2 (N405, N404, N4);
nand NAND2 (N406, N387, N23);
not NOT1 (N407, N359);
nor NOR4 (N408, N401, N244, N177, N256);
buf BUF1 (N409, N405);
nand NAND3 (N410, N399, N172, N209);
and AND2 (N411, N368, N193);
nand NAND4 (N412, N398, N344, N133, N306);
nand NAND3 (N413, N409, N212, N338);
buf BUF1 (N414, N393);
nand NAND2 (N415, N413, N282);
and AND4 (N416, N414, N62, N70, N120);
or OR4 (N417, N415, N108, N21, N212);
buf BUF1 (N418, N407);
not NOT1 (N419, N418);
or OR2 (N420, N419, N390);
xor XOR2 (N421, N408, N225);
nor NOR3 (N422, N410, N54, N40);
buf BUF1 (N423, N416);
buf BUF1 (N424, N422);
xor XOR2 (N425, N417, N189);
buf BUF1 (N426, N421);
nand NAND3 (N427, N424, N145, N118);
and AND2 (N428, N425, N231);
xor XOR2 (N429, N406, N181);
or OR3 (N430, N428, N126, N74);
nand NAND4 (N431, N427, N272, N48, N179);
not NOT1 (N432, N412);
buf BUF1 (N433, N432);
not NOT1 (N434, N411);
nand NAND2 (N435, N429, N402);
not NOT1 (N436, N426);
nand NAND3 (N437, N420, N251, N211);
and AND4 (N438, N423, N3, N260, N247);
nand NAND2 (N439, N430, N136);
buf BUF1 (N440, N433);
and AND4 (N441, N435, N316, N37, N99);
nand NAND4 (N442, N431, N229, N360, N15);
xor XOR2 (N443, N439, N103);
not NOT1 (N444, N437);
and AND2 (N445, N438, N285);
nand NAND2 (N446, N441, N11);
and AND3 (N447, N443, N340, N153);
and AND3 (N448, N447, N431, N173);
nor NOR3 (N449, N442, N255, N399);
buf BUF1 (N450, N446);
xor XOR2 (N451, N450, N416);
nand NAND3 (N452, N440, N146, N171);
nor NOR2 (N453, N434, N366);
nand NAND4 (N454, N400, N435, N230, N6);
or OR4 (N455, N449, N342, N225, N184);
buf BUF1 (N456, N455);
nand NAND2 (N457, N454, N34);
or OR4 (N458, N444, N420, N37, N237);
xor XOR2 (N459, N458, N120);
nand NAND3 (N460, N457, N173, N422);
not NOT1 (N461, N445);
xor XOR2 (N462, N451, N426);
nor NOR2 (N463, N461, N94);
nor NOR3 (N464, N436, N11, N55);
buf BUF1 (N465, N389);
not NOT1 (N466, N459);
nor NOR3 (N467, N452, N341, N310);
and AND3 (N468, N453, N414, N14);
buf BUF1 (N469, N468);
not NOT1 (N470, N469);
not NOT1 (N471, N464);
buf BUF1 (N472, N462);
nor NOR2 (N473, N465, N281);
or OR3 (N474, N467, N299, N114);
and AND2 (N475, N470, N459);
buf BUF1 (N476, N460);
nand NAND3 (N477, N474, N264, N152);
xor XOR2 (N478, N448, N59);
and AND2 (N479, N463, N267);
not NOT1 (N480, N456);
xor XOR2 (N481, N476, N444);
and AND4 (N482, N478, N335, N171, N473);
buf BUF1 (N483, N421);
not NOT1 (N484, N480);
nand NAND3 (N485, N472, N362, N123);
or OR4 (N486, N484, N183, N74, N397);
not NOT1 (N487, N482);
not NOT1 (N488, N485);
nand NAND3 (N489, N466, N294, N268);
not NOT1 (N490, N475);
buf BUF1 (N491, N486);
and AND4 (N492, N481, N211, N175, N11);
buf BUF1 (N493, N492);
nor NOR4 (N494, N490, N69, N364, N429);
or OR4 (N495, N488, N170, N467, N161);
nand NAND4 (N496, N494, N52, N137, N225);
xor XOR2 (N497, N477, N2);
or OR2 (N498, N471, N471);
nor NOR2 (N499, N496, N196);
buf BUF1 (N500, N487);
and AND4 (N501, N497, N134, N361, N181);
not NOT1 (N502, N501);
nor NOR3 (N503, N491, N248, N473);
and AND3 (N504, N500, N258, N404);
or OR2 (N505, N483, N483);
buf BUF1 (N506, N495);
not NOT1 (N507, N499);
and AND4 (N508, N505, N52, N436, N157);
xor XOR2 (N509, N493, N237);
nor NOR4 (N510, N489, N444, N116, N484);
buf BUF1 (N511, N506);
and AND2 (N512, N508, N262);
buf BUF1 (N513, N509);
buf BUF1 (N514, N510);
nor NOR4 (N515, N507, N507, N225, N442);
and AND3 (N516, N504, N4, N373);
or OR3 (N517, N511, N69, N249);
buf BUF1 (N518, N503);
buf BUF1 (N519, N516);
or OR2 (N520, N502, N431);
and AND3 (N521, N520, N516, N154);
nor NOR4 (N522, N514, N293, N484, N172);
xor XOR2 (N523, N522, N324);
xor XOR2 (N524, N479, N85);
and AND4 (N525, N523, N426, N440, N306);
or OR3 (N526, N513, N228, N161);
or OR4 (N527, N517, N284, N354, N235);
nand NAND2 (N528, N525, N54);
or OR3 (N529, N526, N349, N356);
buf BUF1 (N530, N527);
nor NOR2 (N531, N512, N58);
xor XOR2 (N532, N518, N183);
buf BUF1 (N533, N524);
xor XOR2 (N534, N530, N280);
xor XOR2 (N535, N533, N126);
nand NAND3 (N536, N532, N4, N424);
and AND2 (N537, N535, N291);
nor NOR4 (N538, N536, N47, N41, N355);
not NOT1 (N539, N515);
xor XOR2 (N540, N538, N503);
and AND3 (N541, N534, N463, N398);
nor NOR4 (N542, N528, N343, N383, N223);
buf BUF1 (N543, N529);
xor XOR2 (N544, N498, N255);
not NOT1 (N545, N537);
and AND2 (N546, N542, N38);
or OR3 (N547, N541, N373, N63);
and AND4 (N548, N519, N171, N87, N167);
xor XOR2 (N549, N545, N507);
nand NAND4 (N550, N521, N156, N122, N436);
nand NAND3 (N551, N548, N430, N200);
buf BUF1 (N552, N544);
or OR3 (N553, N543, N46, N474);
nand NAND4 (N554, N531, N513, N503, N408);
not NOT1 (N555, N553);
and AND4 (N556, N550, N454, N282, N493);
xor XOR2 (N557, N546, N452);
or OR2 (N558, N549, N526);
or OR3 (N559, N540, N140, N191);
and AND2 (N560, N539, N355);
and AND4 (N561, N554, N355, N335, N54);
buf BUF1 (N562, N561);
buf BUF1 (N563, N557);
and AND3 (N564, N555, N14, N163);
nor NOR2 (N565, N547, N405);
xor XOR2 (N566, N556, N178);
xor XOR2 (N567, N566, N375);
or OR4 (N568, N558, N358, N203, N510);
xor XOR2 (N569, N560, N85);
nand NAND4 (N570, N563, N539, N97, N315);
and AND2 (N571, N564, N175);
nand NAND3 (N572, N552, N422, N114);
buf BUF1 (N573, N570);
nor NOR4 (N574, N565, N188, N380, N547);
buf BUF1 (N575, N567);
not NOT1 (N576, N568);
xor XOR2 (N577, N572, N249);
or OR3 (N578, N574, N407, N47);
buf BUF1 (N579, N576);
nor NOR4 (N580, N569, N489, N370, N6);
xor XOR2 (N581, N579, N474);
not NOT1 (N582, N577);
buf BUF1 (N583, N551);
or OR4 (N584, N581, N402, N42, N292);
nand NAND4 (N585, N578, N356, N305, N545);
not NOT1 (N586, N571);
nor NOR4 (N587, N582, N359, N29, N18);
not NOT1 (N588, N585);
buf BUF1 (N589, N586);
xor XOR2 (N590, N583, N270);
xor XOR2 (N591, N575, N367);
nand NAND2 (N592, N588, N495);
nor NOR3 (N593, N562, N375, N221);
or OR4 (N594, N580, N457, N271, N436);
nand NAND3 (N595, N590, N77, N484);
nor NOR2 (N596, N595, N199);
and AND2 (N597, N591, N592);
nand NAND2 (N598, N407, N371);
nand NAND3 (N599, N573, N189, N514);
nand NAND3 (N600, N559, N6, N462);
nand NAND3 (N601, N597, N271, N453);
buf BUF1 (N602, N587);
xor XOR2 (N603, N584, N107);
nand NAND4 (N604, N599, N141, N39, N166);
or OR3 (N605, N600, N120, N596);
and AND2 (N606, N9, N59);
xor XOR2 (N607, N593, N471);
not NOT1 (N608, N594);
or OR3 (N609, N604, N460, N516);
not NOT1 (N610, N598);
nand NAND4 (N611, N602, N512, N231, N370);
and AND2 (N612, N611, N385);
nand NAND2 (N613, N608, N474);
or OR4 (N614, N603, N255, N176, N519);
not NOT1 (N615, N605);
nand NAND4 (N616, N589, N470, N383, N556);
buf BUF1 (N617, N610);
not NOT1 (N618, N609);
not NOT1 (N619, N618);
or OR4 (N620, N612, N20, N75, N21);
nor NOR2 (N621, N614, N223);
or OR3 (N622, N616, N146, N313);
xor XOR2 (N623, N620, N170);
nor NOR4 (N624, N617, N201, N400, N594);
and AND4 (N625, N621, N178, N392, N27);
or OR3 (N626, N613, N91, N369);
or OR4 (N627, N607, N403, N281, N588);
buf BUF1 (N628, N624);
not NOT1 (N629, N606);
xor XOR2 (N630, N629, N452);
buf BUF1 (N631, N622);
and AND2 (N632, N626, N399);
and AND3 (N633, N623, N512, N234);
nor NOR3 (N634, N632, N452, N552);
nor NOR3 (N635, N634, N516, N257);
and AND4 (N636, N635, N324, N228, N221);
xor XOR2 (N637, N615, N602);
xor XOR2 (N638, N601, N119);
buf BUF1 (N639, N638);
nor NOR3 (N640, N630, N162, N287);
not NOT1 (N641, N631);
buf BUF1 (N642, N627);
not NOT1 (N643, N637);
xor XOR2 (N644, N625, N8);
xor XOR2 (N645, N633, N209);
nor NOR2 (N646, N639, N172);
not NOT1 (N647, N646);
or OR4 (N648, N636, N76, N400, N632);
xor XOR2 (N649, N648, N204);
or OR4 (N650, N619, N325, N53, N395);
and AND2 (N651, N649, N635);
and AND2 (N652, N647, N404);
or OR4 (N653, N640, N247, N555, N218);
not NOT1 (N654, N644);
nand NAND4 (N655, N654, N292, N376, N549);
buf BUF1 (N656, N655);
or OR4 (N657, N653, N187, N349, N301);
and AND3 (N658, N656, N113, N76);
nand NAND4 (N659, N642, N258, N296, N468);
or OR4 (N660, N651, N24, N176, N262);
not NOT1 (N661, N659);
nand NAND2 (N662, N628, N456);
buf BUF1 (N663, N658);
and AND3 (N664, N645, N532, N207);
or OR3 (N665, N661, N88, N646);
xor XOR2 (N666, N665, N33);
xor XOR2 (N667, N662, N636);
nand NAND3 (N668, N652, N510, N282);
nand NAND2 (N669, N657, N506);
not NOT1 (N670, N663);
and AND2 (N671, N650, N24);
xor XOR2 (N672, N668, N576);
nor NOR2 (N673, N672, N437);
not NOT1 (N674, N670);
not NOT1 (N675, N660);
buf BUF1 (N676, N666);
nand NAND2 (N677, N669, N161);
nor NOR2 (N678, N641, N42);
nor NOR3 (N679, N667, N375, N607);
buf BUF1 (N680, N671);
buf BUF1 (N681, N679);
and AND2 (N682, N677, N587);
and AND4 (N683, N680, N639, N80, N377);
or OR4 (N684, N676, N201, N526, N568);
buf BUF1 (N685, N681);
buf BUF1 (N686, N674);
and AND2 (N687, N673, N246);
or OR3 (N688, N683, N117, N308);
and AND2 (N689, N687, N613);
nor NOR4 (N690, N689, N426, N329, N494);
not NOT1 (N691, N664);
nor NOR4 (N692, N691, N365, N134, N628);
nor NOR2 (N693, N688, N442);
and AND4 (N694, N675, N388, N60, N346);
xor XOR2 (N695, N682, N468);
nor NOR3 (N696, N678, N278, N396);
xor XOR2 (N697, N695, N311);
xor XOR2 (N698, N697, N568);
nor NOR3 (N699, N694, N296, N110);
nand NAND2 (N700, N643, N269);
or OR3 (N701, N700, N307, N536);
not NOT1 (N702, N685);
and AND4 (N703, N698, N236, N187, N531);
xor XOR2 (N704, N696, N580);
buf BUF1 (N705, N699);
not NOT1 (N706, N702);
xor XOR2 (N707, N706, N687);
or OR2 (N708, N707, N101);
and AND3 (N709, N684, N550, N542);
nor NOR4 (N710, N690, N414, N143, N268);
nand NAND4 (N711, N705, N318, N55, N368);
xor XOR2 (N712, N692, N415);
xor XOR2 (N713, N712, N136);
nand NAND4 (N714, N710, N268, N569, N113);
not NOT1 (N715, N701);
nor NOR2 (N716, N708, N118);
or OR3 (N717, N686, N34, N343);
nor NOR2 (N718, N704, N312);
nor NOR4 (N719, N713, N184, N110, N342);
nand NAND3 (N720, N709, N595, N108);
buf BUF1 (N721, N716);
nand NAND3 (N722, N714, N356, N21);
not NOT1 (N723, N721);
buf BUF1 (N724, N718);
nor NOR4 (N725, N693, N170, N686, N311);
not NOT1 (N726, N711);
and AND4 (N727, N723, N725, N101, N67);
and AND3 (N728, N587, N140, N329);
xor XOR2 (N729, N727, N223);
buf BUF1 (N730, N728);
not NOT1 (N731, N720);
nand NAND3 (N732, N717, N133, N252);
and AND2 (N733, N715, N419);
not NOT1 (N734, N730);
buf BUF1 (N735, N703);
nand NAND4 (N736, N726, N230, N586, N175);
nand NAND2 (N737, N733, N264);
nand NAND3 (N738, N722, N189, N160);
buf BUF1 (N739, N737);
buf BUF1 (N740, N729);
nor NOR3 (N741, N734, N277, N398);
or OR3 (N742, N738, N242, N599);
nor NOR3 (N743, N735, N594, N254);
or OR3 (N744, N732, N386, N265);
or OR4 (N745, N724, N626, N253, N311);
nor NOR4 (N746, N740, N46, N16, N25);
nor NOR4 (N747, N739, N621, N267, N70);
not NOT1 (N748, N744);
and AND4 (N749, N748, N325, N253, N199);
xor XOR2 (N750, N736, N328);
buf BUF1 (N751, N741);
not NOT1 (N752, N746);
and AND4 (N753, N745, N674, N473, N467);
or OR2 (N754, N742, N605);
xor XOR2 (N755, N753, N539);
or OR2 (N756, N755, N252);
or OR3 (N757, N752, N261, N123);
nand NAND2 (N758, N747, N745);
buf BUF1 (N759, N758);
nand NAND2 (N760, N757, N303);
not NOT1 (N761, N719);
or OR4 (N762, N759, N415, N557, N598);
and AND2 (N763, N756, N567);
nand NAND2 (N764, N749, N376);
buf BUF1 (N765, N761);
buf BUF1 (N766, N754);
not NOT1 (N767, N765);
and AND2 (N768, N763, N742);
nand NAND3 (N769, N764, N554, N43);
not NOT1 (N770, N750);
not NOT1 (N771, N768);
xor XOR2 (N772, N731, N624);
buf BUF1 (N773, N770);
nand NAND3 (N774, N767, N333, N102);
nand NAND3 (N775, N766, N298, N309);
buf BUF1 (N776, N772);
nand NAND2 (N777, N762, N233);
xor XOR2 (N778, N760, N621);
or OR4 (N779, N743, N77, N301, N382);
nor NOR3 (N780, N751, N101, N631);
buf BUF1 (N781, N780);
not NOT1 (N782, N778);
buf BUF1 (N783, N782);
or OR4 (N784, N777, N777, N443, N329);
nand NAND3 (N785, N776, N481, N70);
nor NOR4 (N786, N779, N167, N562, N457);
buf BUF1 (N787, N769);
nor NOR2 (N788, N771, N564);
or OR3 (N789, N783, N393, N451);
nor NOR4 (N790, N789, N321, N54, N374);
buf BUF1 (N791, N790);
nand NAND2 (N792, N787, N721);
and AND2 (N793, N786, N555);
not NOT1 (N794, N773);
buf BUF1 (N795, N793);
nand NAND2 (N796, N785, N577);
nand NAND2 (N797, N794, N384);
xor XOR2 (N798, N784, N60);
buf BUF1 (N799, N798);
buf BUF1 (N800, N791);
and AND3 (N801, N797, N571, N447);
not NOT1 (N802, N792);
not NOT1 (N803, N774);
xor XOR2 (N804, N801, N771);
not NOT1 (N805, N795);
not NOT1 (N806, N788);
not NOT1 (N807, N803);
not NOT1 (N808, N805);
nand NAND3 (N809, N807, N94, N108);
xor XOR2 (N810, N775, N235);
xor XOR2 (N811, N809, N383);
xor XOR2 (N812, N810, N438);
and AND2 (N813, N812, N312);
nor NOR2 (N814, N800, N714);
and AND4 (N815, N802, N258, N80, N733);
nand NAND3 (N816, N799, N733, N692);
or OR3 (N817, N808, N117, N768);
nor NOR3 (N818, N781, N315, N702);
nor NOR2 (N819, N796, N146);
xor XOR2 (N820, N814, N168);
or OR2 (N821, N813, N189);
or OR2 (N822, N811, N712);
and AND2 (N823, N822, N708);
nor NOR2 (N824, N821, N765);
xor XOR2 (N825, N818, N703);
nand NAND4 (N826, N817, N702, N455, N542);
nor NOR2 (N827, N806, N58);
and AND4 (N828, N826, N324, N106, N504);
and AND4 (N829, N824, N605, N690, N770);
nor NOR3 (N830, N827, N551, N423);
or OR3 (N831, N820, N370, N677);
and AND4 (N832, N816, N10, N482, N14);
buf BUF1 (N833, N823);
xor XOR2 (N834, N830, N605);
nand NAND4 (N835, N831, N687, N167, N377);
buf BUF1 (N836, N833);
and AND4 (N837, N829, N785, N420, N497);
xor XOR2 (N838, N836, N530);
and AND2 (N839, N804, N339);
not NOT1 (N840, N835);
nand NAND4 (N841, N839, N203, N760, N18);
xor XOR2 (N842, N828, N422);
nor NOR2 (N843, N842, N321);
not NOT1 (N844, N832);
nand NAND4 (N845, N825, N782, N181, N593);
xor XOR2 (N846, N843, N216);
xor XOR2 (N847, N815, N497);
buf BUF1 (N848, N847);
xor XOR2 (N849, N837, N592);
not NOT1 (N850, N849);
xor XOR2 (N851, N850, N567);
and AND2 (N852, N819, N671);
or OR2 (N853, N844, N640);
or OR2 (N854, N846, N853);
nor NOR4 (N855, N852, N386, N103, N327);
nand NAND2 (N856, N675, N748);
buf BUF1 (N857, N848);
or OR2 (N858, N854, N485);
buf BUF1 (N859, N840);
nor NOR2 (N860, N838, N316);
xor XOR2 (N861, N855, N569);
or OR2 (N862, N861, N141);
and AND3 (N863, N859, N861, N836);
nand NAND2 (N864, N858, N850);
nand NAND4 (N865, N857, N135, N592, N591);
or OR4 (N866, N865, N186, N65, N823);
xor XOR2 (N867, N856, N50);
and AND3 (N868, N867, N430, N143);
buf BUF1 (N869, N862);
buf BUF1 (N870, N841);
or OR3 (N871, N863, N35, N186);
or OR3 (N872, N870, N402, N644);
or OR3 (N873, N864, N30, N496);
not NOT1 (N874, N845);
xor XOR2 (N875, N866, N297);
and AND4 (N876, N873, N150, N750, N862);
nand NAND3 (N877, N874, N44, N14);
xor XOR2 (N878, N877, N816);
nor NOR4 (N879, N878, N253, N564, N829);
nor NOR4 (N880, N834, N497, N861, N500);
not NOT1 (N881, N860);
nor NOR4 (N882, N872, N803, N755, N442);
nor NOR3 (N883, N871, N663, N594);
nand NAND2 (N884, N851, N230);
xor XOR2 (N885, N868, N212);
nor NOR4 (N886, N883, N91, N814, N294);
xor XOR2 (N887, N884, N658);
nor NOR4 (N888, N886, N823, N493, N867);
or OR3 (N889, N876, N688, N153);
nand NAND2 (N890, N888, N748);
or OR3 (N891, N881, N262, N489);
nor NOR2 (N892, N869, N494);
and AND4 (N893, N882, N222, N695, N526);
nand NAND4 (N894, N890, N403, N313, N303);
and AND3 (N895, N892, N511, N352);
buf BUF1 (N896, N894);
nor NOR3 (N897, N887, N829, N463);
not NOT1 (N898, N891);
not NOT1 (N899, N880);
nor NOR3 (N900, N893, N466, N852);
or OR3 (N901, N889, N605, N72);
or OR3 (N902, N875, N791, N500);
or OR3 (N903, N885, N545, N888);
nor NOR3 (N904, N898, N586, N466);
nor NOR3 (N905, N879, N397, N512);
not NOT1 (N906, N904);
xor XOR2 (N907, N899, N157);
nand NAND4 (N908, N901, N125, N844, N645);
nand NAND4 (N909, N896, N477, N815, N453);
nor NOR4 (N910, N897, N254, N438, N657);
and AND2 (N911, N900, N118);
nor NOR4 (N912, N911, N698, N227, N593);
buf BUF1 (N913, N910);
buf BUF1 (N914, N913);
xor XOR2 (N915, N895, N356);
nor NOR4 (N916, N912, N144, N412, N655);
xor XOR2 (N917, N908, N787);
not NOT1 (N918, N903);
not NOT1 (N919, N902);
buf BUF1 (N920, N909);
nand NAND3 (N921, N917, N820, N613);
nor NOR4 (N922, N907, N687, N124, N702);
nor NOR4 (N923, N906, N336, N905, N776);
nand NAND3 (N924, N153, N223, N230);
nand NAND3 (N925, N915, N374, N560);
xor XOR2 (N926, N919, N200);
buf BUF1 (N927, N916);
xor XOR2 (N928, N925, N332);
or OR3 (N929, N928, N84, N911);
and AND3 (N930, N914, N929, N692);
and AND2 (N931, N254, N912);
nor NOR3 (N932, N922, N558, N356);
buf BUF1 (N933, N923);
or OR2 (N934, N920, N721);
not NOT1 (N935, N934);
nand NAND4 (N936, N924, N847, N549, N666);
nand NAND3 (N937, N933, N19, N394);
not NOT1 (N938, N937);
not NOT1 (N939, N921);
or OR2 (N940, N931, N140);
and AND4 (N941, N935, N586, N249, N861);
not NOT1 (N942, N932);
xor XOR2 (N943, N940, N849);
buf BUF1 (N944, N938);
or OR4 (N945, N936, N727, N889, N623);
not NOT1 (N946, N918);
xor XOR2 (N947, N943, N25);
or OR2 (N948, N941, N856);
nor NOR3 (N949, N948, N37, N941);
and AND2 (N950, N942, N581);
nand NAND4 (N951, N930, N936, N591, N700);
nor NOR2 (N952, N949, N705);
or OR3 (N953, N951, N324, N294);
and AND2 (N954, N947, N398);
xor XOR2 (N955, N954, N397);
buf BUF1 (N956, N945);
buf BUF1 (N957, N955);
and AND4 (N958, N927, N96, N363, N673);
nand NAND4 (N959, N958, N729, N474, N869);
not NOT1 (N960, N950);
xor XOR2 (N961, N960, N424);
xor XOR2 (N962, N957, N627);
nor NOR2 (N963, N961, N878);
not NOT1 (N964, N959);
nor NOR4 (N965, N964, N872, N325, N124);
and AND2 (N966, N946, N256);
xor XOR2 (N967, N953, N850);
buf BUF1 (N968, N966);
buf BUF1 (N969, N956);
buf BUF1 (N970, N926);
or OR3 (N971, N962, N793, N643);
nand NAND2 (N972, N939, N581);
nor NOR2 (N973, N952, N373);
and AND3 (N974, N972, N923, N645);
not NOT1 (N975, N971);
nor NOR3 (N976, N963, N420, N125);
xor XOR2 (N977, N965, N875);
not NOT1 (N978, N976);
xor XOR2 (N979, N978, N819);
xor XOR2 (N980, N975, N123);
or OR4 (N981, N980, N435, N339, N114);
nor NOR4 (N982, N968, N505, N240, N224);
nor NOR2 (N983, N979, N4);
buf BUF1 (N984, N981);
nand NAND2 (N985, N977, N706);
not NOT1 (N986, N973);
nand NAND2 (N987, N984, N496);
xor XOR2 (N988, N985, N643);
xor XOR2 (N989, N986, N387);
or OR2 (N990, N982, N659);
buf BUF1 (N991, N983);
nand NAND4 (N992, N974, N571, N905, N31);
xor XOR2 (N993, N969, N574);
nand NAND3 (N994, N991, N920, N929);
or OR2 (N995, N970, N533);
nand NAND4 (N996, N990, N748, N131, N601);
or OR2 (N997, N996, N639);
nor NOR2 (N998, N989, N65);
or OR4 (N999, N988, N198, N464, N180);
not NOT1 (N1000, N993);
not NOT1 (N1001, N967);
nand NAND4 (N1002, N992, N483, N803, N369);
nor NOR4 (N1003, N998, N514, N962, N40);
not NOT1 (N1004, N944);
nand NAND4 (N1005, N997, N997, N639, N446);
xor XOR2 (N1006, N1004, N145);
nand NAND4 (N1007, N1000, N751, N362, N448);
or OR2 (N1008, N994, N87);
not NOT1 (N1009, N995);
or OR4 (N1010, N1007, N483, N786, N125);
and AND2 (N1011, N1009, N69);
xor XOR2 (N1012, N1003, N572);
not NOT1 (N1013, N1010);
and AND4 (N1014, N987, N431, N408, N669);
nand NAND2 (N1015, N1014, N384);
buf BUF1 (N1016, N1012);
or OR3 (N1017, N1008, N975, N897);
or OR4 (N1018, N1011, N290, N465, N714);
nand NAND3 (N1019, N1016, N552, N733);
buf BUF1 (N1020, N1017);
not NOT1 (N1021, N1006);
xor XOR2 (N1022, N1018, N955);
xor XOR2 (N1023, N1001, N545);
nor NOR4 (N1024, N1020, N604, N33, N97);
or OR2 (N1025, N1021, N581);
nor NOR3 (N1026, N1023, N101, N268);
or OR4 (N1027, N999, N195, N707, N637);
buf BUF1 (N1028, N1022);
xor XOR2 (N1029, N1019, N691);
or OR3 (N1030, N1025, N188, N1010);
and AND3 (N1031, N1029, N855, N115);
xor XOR2 (N1032, N1027, N938);
and AND3 (N1033, N1002, N311, N599);
buf BUF1 (N1034, N1028);
buf BUF1 (N1035, N1031);
or OR2 (N1036, N1033, N140);
and AND2 (N1037, N1030, N635);
nor NOR4 (N1038, N1015, N398, N232, N684);
and AND4 (N1039, N1036, N686, N652, N869);
and AND3 (N1040, N1039, N56, N912);
nand NAND3 (N1041, N1034, N645, N532);
xor XOR2 (N1042, N1037, N205);
nand NAND4 (N1043, N1035, N48, N771, N861);
not NOT1 (N1044, N1024);
xor XOR2 (N1045, N1042, N461);
or OR4 (N1046, N1041, N143, N363, N174);
nor NOR2 (N1047, N1044, N218);
nand NAND3 (N1048, N1026, N374, N868);
xor XOR2 (N1049, N1038, N985);
not NOT1 (N1050, N1046);
buf BUF1 (N1051, N1005);
not NOT1 (N1052, N1043);
and AND2 (N1053, N1051, N208);
not NOT1 (N1054, N1013);
nand NAND2 (N1055, N1049, N167);
nand NAND4 (N1056, N1053, N349, N345, N746);
and AND4 (N1057, N1040, N867, N380, N4);
not NOT1 (N1058, N1050);
nor NOR3 (N1059, N1056, N859, N321);
buf BUF1 (N1060, N1055);
or OR4 (N1061, N1059, N297, N583, N974);
or OR3 (N1062, N1057, N256, N281);
nand NAND3 (N1063, N1060, N812, N285);
nor NOR2 (N1064, N1047, N74);
not NOT1 (N1065, N1061);
buf BUF1 (N1066, N1058);
and AND2 (N1067, N1048, N181);
and AND2 (N1068, N1052, N156);
nand NAND3 (N1069, N1066, N1052, N380);
and AND4 (N1070, N1054, N795, N313, N1061);
not NOT1 (N1071, N1065);
buf BUF1 (N1072, N1045);
buf BUF1 (N1073, N1069);
and AND2 (N1074, N1062, N863);
xor XOR2 (N1075, N1064, N905);
not NOT1 (N1076, N1063);
nor NOR4 (N1077, N1070, N424, N697, N640);
nor NOR2 (N1078, N1077, N243);
and AND2 (N1079, N1075, N793);
nor NOR4 (N1080, N1032, N611, N160, N999);
buf BUF1 (N1081, N1067);
nor NOR2 (N1082, N1072, N877);
xor XOR2 (N1083, N1076, N598);
or OR2 (N1084, N1074, N102);
buf BUF1 (N1085, N1071);
xor XOR2 (N1086, N1083, N320);
or OR2 (N1087, N1086, N975);
not NOT1 (N1088, N1078);
and AND4 (N1089, N1081, N120, N671, N925);
buf BUF1 (N1090, N1082);
nor NOR2 (N1091, N1085, N949);
and AND2 (N1092, N1090, N75);
nor NOR4 (N1093, N1080, N4, N962, N495);
nand NAND2 (N1094, N1093, N318);
nor NOR4 (N1095, N1084, N718, N944, N585);
nor NOR2 (N1096, N1092, N537);
not NOT1 (N1097, N1073);
and AND3 (N1098, N1088, N972, N698);
nand NAND2 (N1099, N1095, N928);
nand NAND3 (N1100, N1091, N595, N386);
nor NOR2 (N1101, N1099, N841);
buf BUF1 (N1102, N1097);
not NOT1 (N1103, N1098);
xor XOR2 (N1104, N1068, N1038);
xor XOR2 (N1105, N1087, N12);
not NOT1 (N1106, N1096);
xor XOR2 (N1107, N1079, N205);
buf BUF1 (N1108, N1089);
xor XOR2 (N1109, N1094, N95);
or OR3 (N1110, N1106, N109, N151);
or OR2 (N1111, N1102, N862);
or OR3 (N1112, N1107, N20, N67);
nor NOR3 (N1113, N1105, N663, N678);
and AND3 (N1114, N1101, N544, N855);
not NOT1 (N1115, N1111);
and AND4 (N1116, N1110, N604, N20, N628);
buf BUF1 (N1117, N1116);
buf BUF1 (N1118, N1100);
and AND3 (N1119, N1104, N297, N79);
nand NAND3 (N1120, N1119, N583, N886);
nor NOR2 (N1121, N1114, N678);
or OR2 (N1122, N1117, N666);
and AND3 (N1123, N1118, N1017, N20);
not NOT1 (N1124, N1103);
or OR4 (N1125, N1123, N461, N165, N926);
nor NOR2 (N1126, N1112, N154);
nor NOR3 (N1127, N1121, N325, N555);
and AND3 (N1128, N1109, N145, N510);
nor NOR2 (N1129, N1113, N1118);
and AND4 (N1130, N1120, N664, N363, N605);
nand NAND2 (N1131, N1130, N645);
not NOT1 (N1132, N1128);
nand NAND2 (N1133, N1131, N1013);
nand NAND2 (N1134, N1132, N1120);
nand NAND3 (N1135, N1124, N878, N1042);
not NOT1 (N1136, N1115);
nand NAND4 (N1137, N1134, N644, N1113, N997);
nor NOR3 (N1138, N1136, N324, N670);
xor XOR2 (N1139, N1133, N854);
nor NOR4 (N1140, N1127, N574, N197, N613);
xor XOR2 (N1141, N1125, N972);
or OR2 (N1142, N1141, N555);
not NOT1 (N1143, N1140);
or OR4 (N1144, N1135, N160, N749, N543);
not NOT1 (N1145, N1126);
and AND2 (N1146, N1108, N621);
nor NOR2 (N1147, N1143, N871);
and AND3 (N1148, N1138, N428, N1131);
not NOT1 (N1149, N1146);
not NOT1 (N1150, N1139);
or OR2 (N1151, N1137, N965);
and AND4 (N1152, N1122, N1028, N36, N745);
nand NAND2 (N1153, N1150, N224);
and AND4 (N1154, N1142, N499, N714, N116);
and AND4 (N1155, N1149, N633, N454, N942);
buf BUF1 (N1156, N1155);
nor NOR4 (N1157, N1152, N559, N1150, N600);
xor XOR2 (N1158, N1148, N330);
xor XOR2 (N1159, N1145, N502);
nor NOR4 (N1160, N1158, N531, N361, N263);
or OR2 (N1161, N1156, N777);
nand NAND2 (N1162, N1129, N707);
and AND2 (N1163, N1144, N139);
and AND2 (N1164, N1153, N339);
nor NOR4 (N1165, N1157, N690, N663, N819);
not NOT1 (N1166, N1159);
nor NOR4 (N1167, N1165, N789, N1125, N177);
nand NAND3 (N1168, N1164, N136, N387);
not NOT1 (N1169, N1163);
nand NAND4 (N1170, N1169, N605, N444, N945);
not NOT1 (N1171, N1170);
or OR3 (N1172, N1166, N193, N982);
nand NAND4 (N1173, N1171, N78, N729, N349);
nor NOR3 (N1174, N1161, N678, N400);
or OR3 (N1175, N1151, N779, N539);
nand NAND2 (N1176, N1168, N447);
or OR2 (N1177, N1173, N413);
buf BUF1 (N1178, N1154);
nand NAND2 (N1179, N1162, N54);
and AND4 (N1180, N1172, N586, N93, N942);
xor XOR2 (N1181, N1160, N25);
buf BUF1 (N1182, N1174);
not NOT1 (N1183, N1180);
xor XOR2 (N1184, N1176, N254);
nand NAND3 (N1185, N1182, N870, N481);
nor NOR3 (N1186, N1184, N325, N936);
xor XOR2 (N1187, N1185, N131);
nand NAND4 (N1188, N1167, N300, N568, N1147);
and AND2 (N1189, N983, N341);
nor NOR3 (N1190, N1178, N244, N676);
nand NAND4 (N1191, N1181, N713, N861, N594);
not NOT1 (N1192, N1186);
or OR3 (N1193, N1179, N555, N276);
buf BUF1 (N1194, N1192);
or OR4 (N1195, N1175, N711, N1031, N324);
nor NOR4 (N1196, N1195, N10, N485, N215);
nand NAND2 (N1197, N1193, N680);
and AND2 (N1198, N1187, N85);
not NOT1 (N1199, N1177);
not NOT1 (N1200, N1188);
buf BUF1 (N1201, N1198);
and AND4 (N1202, N1196, N1171, N547, N199);
not NOT1 (N1203, N1189);
or OR2 (N1204, N1199, N113);
not NOT1 (N1205, N1191);
not NOT1 (N1206, N1200);
and AND4 (N1207, N1202, N822, N987, N1011);
not NOT1 (N1208, N1201);
nand NAND4 (N1209, N1183, N981, N992, N303);
and AND3 (N1210, N1208, N399, N84);
xor XOR2 (N1211, N1205, N352);
nand NAND4 (N1212, N1203, N389, N629, N1046);
or OR2 (N1213, N1207, N155);
nand NAND4 (N1214, N1194, N580, N44, N578);
nor NOR3 (N1215, N1206, N469, N987);
buf BUF1 (N1216, N1213);
buf BUF1 (N1217, N1215);
nand NAND2 (N1218, N1190, N1076);
and AND3 (N1219, N1210, N103, N725);
not NOT1 (N1220, N1219);
not NOT1 (N1221, N1217);
nor NOR4 (N1222, N1204, N861, N917, N428);
nor NOR3 (N1223, N1220, N342, N488);
not NOT1 (N1224, N1209);
not NOT1 (N1225, N1218);
not NOT1 (N1226, N1197);
buf BUF1 (N1227, N1222);
buf BUF1 (N1228, N1227);
or OR2 (N1229, N1224, N463);
buf BUF1 (N1230, N1229);
or OR4 (N1231, N1216, N1180, N407, N1129);
xor XOR2 (N1232, N1225, N1206);
nor NOR4 (N1233, N1212, N95, N1193, N678);
xor XOR2 (N1234, N1226, N803);
buf BUF1 (N1235, N1228);
or OR4 (N1236, N1221, N243, N125, N799);
buf BUF1 (N1237, N1235);
and AND2 (N1238, N1214, N1016);
nand NAND2 (N1239, N1231, N285);
and AND4 (N1240, N1232, N1111, N1197, N282);
nand NAND3 (N1241, N1238, N934, N973);
buf BUF1 (N1242, N1236);
nand NAND2 (N1243, N1234, N34);
nor NOR3 (N1244, N1237, N653, N163);
nor NOR3 (N1245, N1223, N1235, N157);
or OR4 (N1246, N1240, N975, N821, N351);
and AND3 (N1247, N1242, N241, N586);
buf BUF1 (N1248, N1211);
buf BUF1 (N1249, N1248);
or OR2 (N1250, N1246, N885);
or OR4 (N1251, N1243, N1105, N1233, N154);
not NOT1 (N1252, N480);
or OR2 (N1253, N1251, N532);
and AND3 (N1254, N1250, N392, N357);
and AND3 (N1255, N1253, N785, N166);
and AND4 (N1256, N1230, N209, N606, N717);
or OR3 (N1257, N1247, N271, N688);
not NOT1 (N1258, N1244);
nand NAND2 (N1259, N1252, N168);
nand NAND4 (N1260, N1241, N277, N1152, N1182);
and AND3 (N1261, N1259, N425, N408);
or OR2 (N1262, N1254, N1003);
not NOT1 (N1263, N1257);
buf BUF1 (N1264, N1261);
or OR3 (N1265, N1258, N969, N752);
and AND4 (N1266, N1255, N644, N898, N812);
or OR3 (N1267, N1260, N1087, N272);
nor NOR4 (N1268, N1262, N237, N961, N24);
and AND3 (N1269, N1249, N649, N995);
not NOT1 (N1270, N1265);
or OR2 (N1271, N1266, N1154);
not NOT1 (N1272, N1267);
xor XOR2 (N1273, N1272, N515);
buf BUF1 (N1274, N1264);
or OR3 (N1275, N1273, N973, N946);
nand NAND2 (N1276, N1268, N435);
and AND2 (N1277, N1271, N750);
and AND2 (N1278, N1239, N1224);
xor XOR2 (N1279, N1245, N1214);
or OR4 (N1280, N1279, N884, N822, N264);
or OR4 (N1281, N1263, N688, N359, N1240);
nand NAND4 (N1282, N1278, N470, N313, N905);
buf BUF1 (N1283, N1280);
nand NAND3 (N1284, N1282, N844, N540);
nor NOR3 (N1285, N1270, N1149, N1208);
nand NAND2 (N1286, N1275, N20);
nand NAND2 (N1287, N1269, N170);
or OR2 (N1288, N1281, N190);
nand NAND4 (N1289, N1284, N245, N616, N340);
or OR3 (N1290, N1277, N539, N1269);
or OR4 (N1291, N1289, N1083, N1092, N550);
not NOT1 (N1292, N1283);
and AND3 (N1293, N1290, N154, N114);
xor XOR2 (N1294, N1256, N133);
or OR2 (N1295, N1291, N227);
not NOT1 (N1296, N1292);
and AND3 (N1297, N1288, N1198, N703);
buf BUF1 (N1298, N1293);
or OR4 (N1299, N1285, N717, N1151, N867);
nor NOR3 (N1300, N1287, N103, N455);
not NOT1 (N1301, N1294);
or OR3 (N1302, N1298, N201, N1215);
and AND3 (N1303, N1276, N757, N583);
buf BUF1 (N1304, N1296);
nand NAND3 (N1305, N1303, N921, N81);
and AND3 (N1306, N1274, N112, N702);
nor NOR2 (N1307, N1297, N38);
nor NOR4 (N1308, N1301, N1270, N1261, N1299);
nor NOR2 (N1309, N73, N1099);
not NOT1 (N1310, N1307);
and AND4 (N1311, N1300, N1138, N180, N373);
nor NOR3 (N1312, N1286, N760, N480);
xor XOR2 (N1313, N1308, N1251);
nand NAND2 (N1314, N1311, N1094);
buf BUF1 (N1315, N1314);
nor NOR3 (N1316, N1315, N1051, N139);
or OR4 (N1317, N1304, N558, N259, N1198);
nand NAND3 (N1318, N1313, N774, N646);
buf BUF1 (N1319, N1305);
xor XOR2 (N1320, N1306, N861);
and AND3 (N1321, N1316, N115, N991);
or OR2 (N1322, N1302, N806);
xor XOR2 (N1323, N1319, N566);
nand NAND2 (N1324, N1322, N659);
not NOT1 (N1325, N1321);
nor NOR2 (N1326, N1310, N957);
nand NAND3 (N1327, N1325, N743, N402);
xor XOR2 (N1328, N1327, N253);
and AND4 (N1329, N1317, N84, N553, N258);
and AND2 (N1330, N1328, N558);
buf BUF1 (N1331, N1323);
not NOT1 (N1332, N1330);
or OR4 (N1333, N1329, N709, N990, N699);
not NOT1 (N1334, N1332);
or OR3 (N1335, N1324, N1227, N120);
nor NOR3 (N1336, N1326, N798, N271);
xor XOR2 (N1337, N1334, N929);
xor XOR2 (N1338, N1312, N666);
nand NAND3 (N1339, N1318, N412, N1272);
not NOT1 (N1340, N1309);
not NOT1 (N1341, N1337);
buf BUF1 (N1342, N1339);
or OR4 (N1343, N1336, N970, N663, N871);
or OR3 (N1344, N1295, N1214, N975);
nor NOR3 (N1345, N1320, N1100, N389);
buf BUF1 (N1346, N1335);
nor NOR3 (N1347, N1331, N1305, N1093);
nand NAND4 (N1348, N1344, N39, N887, N1338);
or OR4 (N1349, N11, N150, N1095, N176);
not NOT1 (N1350, N1333);
nand NAND2 (N1351, N1341, N1013);
and AND2 (N1352, N1351, N478);
buf BUF1 (N1353, N1352);
not NOT1 (N1354, N1350);
or OR4 (N1355, N1346, N904, N380, N662);
xor XOR2 (N1356, N1353, N139);
or OR3 (N1357, N1356, N1033, N359);
nor NOR3 (N1358, N1348, N1062, N78);
not NOT1 (N1359, N1343);
xor XOR2 (N1360, N1357, N648);
or OR2 (N1361, N1360, N111);
not NOT1 (N1362, N1355);
buf BUF1 (N1363, N1347);
nor NOR3 (N1364, N1358, N435, N229);
nor NOR4 (N1365, N1359, N1293, N654, N813);
nor NOR4 (N1366, N1349, N162, N897, N1348);
and AND3 (N1367, N1362, N122, N232);
nor NOR2 (N1368, N1364, N1077);
xor XOR2 (N1369, N1368, N1057);
nor NOR4 (N1370, N1369, N326, N1, N1070);
nor NOR4 (N1371, N1367, N606, N37, N320);
not NOT1 (N1372, N1342);
and AND3 (N1373, N1354, N1308, N204);
or OR2 (N1374, N1340, N462);
xor XOR2 (N1375, N1374, N871);
nor NOR2 (N1376, N1372, N717);
not NOT1 (N1377, N1376);
buf BUF1 (N1378, N1345);
xor XOR2 (N1379, N1371, N190);
nor NOR3 (N1380, N1361, N312, N1139);
buf BUF1 (N1381, N1365);
or OR3 (N1382, N1373, N375, N837);
xor XOR2 (N1383, N1363, N1149);
nand NAND2 (N1384, N1380, N579);
buf BUF1 (N1385, N1379);
or OR3 (N1386, N1381, N1293, N893);
nor NOR3 (N1387, N1370, N1354, N364);
or OR3 (N1388, N1382, N765, N869);
and AND4 (N1389, N1388, N17, N949, N989);
nor NOR4 (N1390, N1375, N585, N971, N954);
buf BUF1 (N1391, N1377);
and AND2 (N1392, N1385, N342);
not NOT1 (N1393, N1384);
and AND3 (N1394, N1391, N183, N1142);
xor XOR2 (N1395, N1393, N1350);
or OR4 (N1396, N1387, N242, N332, N925);
buf BUF1 (N1397, N1386);
not NOT1 (N1398, N1366);
buf BUF1 (N1399, N1397);
xor XOR2 (N1400, N1394, N259);
nand NAND4 (N1401, N1383, N1177, N716, N332);
and AND2 (N1402, N1401, N124);
nor NOR2 (N1403, N1395, N782);
not NOT1 (N1404, N1398);
nand NAND2 (N1405, N1402, N30);
and AND2 (N1406, N1390, N898);
and AND4 (N1407, N1404, N445, N118, N1237);
or OR2 (N1408, N1396, N1121);
buf BUF1 (N1409, N1407);
xor XOR2 (N1410, N1408, N142);
and AND3 (N1411, N1400, N446, N1258);
buf BUF1 (N1412, N1411);
and AND4 (N1413, N1389, N321, N1209, N22);
buf BUF1 (N1414, N1409);
buf BUF1 (N1415, N1410);
xor XOR2 (N1416, N1403, N850);
nor NOR3 (N1417, N1399, N953, N1382);
and AND3 (N1418, N1406, N318, N925);
not NOT1 (N1419, N1378);
not NOT1 (N1420, N1419);
xor XOR2 (N1421, N1417, N818);
and AND4 (N1422, N1418, N1299, N1380, N441);
nand NAND4 (N1423, N1405, N774, N951, N930);
nand NAND4 (N1424, N1414, N675, N1128, N783);
nand NAND3 (N1425, N1392, N1040, N198);
nor NOR2 (N1426, N1423, N546);
nor NOR4 (N1427, N1424, N1003, N937, N924);
nand NAND2 (N1428, N1425, N986);
or OR2 (N1429, N1413, N458);
not NOT1 (N1430, N1428);
and AND4 (N1431, N1429, N635, N1205, N865);
not NOT1 (N1432, N1422);
xor XOR2 (N1433, N1420, N956);
nor NOR2 (N1434, N1416, N1103);
not NOT1 (N1435, N1421);
xor XOR2 (N1436, N1412, N712);
and AND2 (N1437, N1427, N990);
nor NOR4 (N1438, N1426, N235, N4, N269);
and AND2 (N1439, N1431, N402);
xor XOR2 (N1440, N1437, N182);
xor XOR2 (N1441, N1433, N1188);
xor XOR2 (N1442, N1440, N362);
and AND3 (N1443, N1430, N1186, N1238);
or OR4 (N1444, N1438, N711, N1397, N583);
or OR3 (N1445, N1432, N445, N773);
xor XOR2 (N1446, N1442, N502);
nor NOR2 (N1447, N1415, N270);
and AND3 (N1448, N1435, N1025, N324);
not NOT1 (N1449, N1436);
nand NAND3 (N1450, N1444, N855, N742);
nor NOR3 (N1451, N1441, N647, N406);
not NOT1 (N1452, N1449);
not NOT1 (N1453, N1447);
buf BUF1 (N1454, N1443);
buf BUF1 (N1455, N1448);
buf BUF1 (N1456, N1451);
buf BUF1 (N1457, N1445);
nor NOR2 (N1458, N1446, N34);
xor XOR2 (N1459, N1434, N1343);
nor NOR3 (N1460, N1458, N1033, N237);
nor NOR2 (N1461, N1455, N555);
nor NOR3 (N1462, N1439, N1068, N357);
not NOT1 (N1463, N1454);
nor NOR3 (N1464, N1457, N806, N675);
nand NAND3 (N1465, N1452, N555, N469);
nand NAND3 (N1466, N1459, N379, N484);
nor NOR2 (N1467, N1464, N473);
not NOT1 (N1468, N1450);
not NOT1 (N1469, N1460);
nand NAND2 (N1470, N1465, N479);
and AND4 (N1471, N1461, N1355, N1455, N566);
buf BUF1 (N1472, N1462);
xor XOR2 (N1473, N1469, N623);
xor XOR2 (N1474, N1471, N1167);
nor NOR2 (N1475, N1466, N641);
nand NAND4 (N1476, N1468, N1414, N1017, N376);
nor NOR4 (N1477, N1473, N1469, N458, N1222);
nor NOR3 (N1478, N1456, N1021, N217);
not NOT1 (N1479, N1472);
and AND4 (N1480, N1478, N674, N885, N30);
nand NAND4 (N1481, N1475, N1002, N1085, N171);
nor NOR3 (N1482, N1453, N241, N317);
nand NAND3 (N1483, N1476, N1267, N518);
nand NAND4 (N1484, N1467, N865, N353, N1102);
nand NAND4 (N1485, N1480, N513, N980, N1300);
nor NOR2 (N1486, N1477, N1136);
or OR4 (N1487, N1474, N1202, N911, N45);
nor NOR3 (N1488, N1483, N1370, N786);
not NOT1 (N1489, N1463);
or OR4 (N1490, N1481, N1103, N118, N893);
and AND2 (N1491, N1487, N459);
not NOT1 (N1492, N1488);
or OR4 (N1493, N1479, N425, N1255, N920);
xor XOR2 (N1494, N1485, N1239);
or OR3 (N1495, N1494, N961, N106);
not NOT1 (N1496, N1484);
nor NOR3 (N1497, N1482, N1199, N776);
buf BUF1 (N1498, N1496);
not NOT1 (N1499, N1489);
xor XOR2 (N1500, N1498, N679);
and AND3 (N1501, N1492, N862, N1102);
xor XOR2 (N1502, N1493, N218);
buf BUF1 (N1503, N1500);
or OR2 (N1504, N1486, N770);
or OR4 (N1505, N1495, N203, N274, N336);
nor NOR4 (N1506, N1504, N29, N967, N262);
nand NAND4 (N1507, N1497, N956, N1143, N271);
nor NOR4 (N1508, N1505, N742, N747, N1380);
xor XOR2 (N1509, N1503, N36);
nor NOR3 (N1510, N1507, N174, N1148);
nor NOR2 (N1511, N1491, N754);
or OR2 (N1512, N1510, N977);
or OR4 (N1513, N1508, N18, N139, N1317);
not NOT1 (N1514, N1509);
and AND4 (N1515, N1501, N1230, N944, N1497);
and AND2 (N1516, N1506, N1081);
nand NAND4 (N1517, N1511, N855, N1192, N905);
not NOT1 (N1518, N1502);
xor XOR2 (N1519, N1499, N660);
nand NAND2 (N1520, N1519, N1451);
nor NOR3 (N1521, N1514, N522, N1382);
or OR3 (N1522, N1516, N1055, N1175);
not NOT1 (N1523, N1517);
xor XOR2 (N1524, N1523, N1052);
nor NOR3 (N1525, N1520, N584, N1312);
not NOT1 (N1526, N1518);
not NOT1 (N1527, N1512);
or OR2 (N1528, N1513, N655);
buf BUF1 (N1529, N1522);
and AND3 (N1530, N1470, N1008, N103);
xor XOR2 (N1531, N1530, N1427);
xor XOR2 (N1532, N1524, N125);
not NOT1 (N1533, N1526);
nand NAND3 (N1534, N1531, N1300, N529);
or OR2 (N1535, N1528, N770);
and AND4 (N1536, N1533, N74, N755, N1032);
nand NAND4 (N1537, N1515, N1445, N420, N224);
or OR4 (N1538, N1534, N94, N591, N870);
buf BUF1 (N1539, N1536);
xor XOR2 (N1540, N1525, N677);
or OR4 (N1541, N1490, N535, N1081, N322);
not NOT1 (N1542, N1535);
or OR2 (N1543, N1532, N917);
xor XOR2 (N1544, N1539, N464);
nand NAND2 (N1545, N1521, N628);
nor NOR2 (N1546, N1540, N744);
not NOT1 (N1547, N1543);
nor NOR3 (N1548, N1527, N748, N1415);
or OR2 (N1549, N1538, N1287);
buf BUF1 (N1550, N1545);
or OR2 (N1551, N1547, N1126);
buf BUF1 (N1552, N1550);
nor NOR2 (N1553, N1552, N5);
nor NOR2 (N1554, N1546, N238);
and AND4 (N1555, N1541, N956, N1145, N372);
buf BUF1 (N1556, N1555);
nand NAND4 (N1557, N1542, N805, N134, N1206);
or OR2 (N1558, N1549, N740);
buf BUF1 (N1559, N1537);
or OR3 (N1560, N1548, N1212, N330);
or OR2 (N1561, N1556, N325);
buf BUF1 (N1562, N1544);
buf BUF1 (N1563, N1559);
nor NOR4 (N1564, N1551, N1385, N756, N187);
xor XOR2 (N1565, N1529, N766);
nor NOR4 (N1566, N1565, N803, N919, N1367);
and AND2 (N1567, N1561, N537);
or OR3 (N1568, N1566, N458, N163);
not NOT1 (N1569, N1567);
or OR2 (N1570, N1568, N163);
and AND4 (N1571, N1564, N635, N267, N227);
xor XOR2 (N1572, N1554, N1039);
buf BUF1 (N1573, N1553);
not NOT1 (N1574, N1571);
nand NAND2 (N1575, N1557, N890);
buf BUF1 (N1576, N1572);
or OR4 (N1577, N1563, N1083, N215, N1276);
and AND2 (N1578, N1560, N3);
nor NOR4 (N1579, N1574, N74, N1554, N1235);
nor NOR2 (N1580, N1575, N1213);
xor XOR2 (N1581, N1573, N1433);
buf BUF1 (N1582, N1576);
or OR3 (N1583, N1578, N733, N1088);
xor XOR2 (N1584, N1558, N1561);
nand NAND4 (N1585, N1584, N836, N414, N380);
xor XOR2 (N1586, N1583, N11);
and AND2 (N1587, N1569, N1548);
nor NOR3 (N1588, N1579, N1384, N1117);
nand NAND4 (N1589, N1562, N1443, N1514, N83);
nand NAND4 (N1590, N1589, N1338, N761, N1282);
or OR3 (N1591, N1577, N250, N817);
xor XOR2 (N1592, N1587, N434);
buf BUF1 (N1593, N1582);
nor NOR3 (N1594, N1580, N356, N1360);
not NOT1 (N1595, N1593);
xor XOR2 (N1596, N1581, N215);
nor NOR3 (N1597, N1586, N240, N824);
nor NOR4 (N1598, N1591, N663, N360, N1103);
or OR3 (N1599, N1598, N478, N72);
or OR2 (N1600, N1570, N872);
xor XOR2 (N1601, N1585, N875);
xor XOR2 (N1602, N1594, N291);
nor NOR3 (N1603, N1601, N981, N643);
buf BUF1 (N1604, N1596);
xor XOR2 (N1605, N1604, N212);
nand NAND2 (N1606, N1600, N539);
nor NOR2 (N1607, N1590, N1108);
or OR3 (N1608, N1603, N243, N818);
nor NOR2 (N1609, N1602, N1523);
nand NAND2 (N1610, N1588, N686);
or OR3 (N1611, N1597, N1297, N469);
and AND3 (N1612, N1599, N288, N340);
nand NAND2 (N1613, N1607, N1424);
and AND2 (N1614, N1605, N18);
or OR3 (N1615, N1592, N96, N399);
xor XOR2 (N1616, N1615, N173);
or OR3 (N1617, N1614, N652, N347);
nand NAND3 (N1618, N1611, N608, N1138);
not NOT1 (N1619, N1608);
or OR4 (N1620, N1609, N329, N1102, N882);
nand NAND3 (N1621, N1618, N1324, N1110);
nor NOR3 (N1622, N1595, N239, N20);
and AND4 (N1623, N1613, N1559, N1031, N1577);
not NOT1 (N1624, N1617);
not NOT1 (N1625, N1606);
xor XOR2 (N1626, N1622, N668);
or OR3 (N1627, N1624, N1234, N744);
xor XOR2 (N1628, N1616, N642);
nand NAND4 (N1629, N1628, N691, N997, N1326);
and AND3 (N1630, N1620, N227, N1626);
not NOT1 (N1631, N732);
and AND3 (N1632, N1623, N551, N2);
or OR4 (N1633, N1629, N91, N751, N1194);
nand NAND3 (N1634, N1612, N1326, N1146);
and AND4 (N1635, N1630, N584, N317, N1172);
buf BUF1 (N1636, N1619);
xor XOR2 (N1637, N1610, N199);
and AND3 (N1638, N1635, N766, N1495);
xor XOR2 (N1639, N1637, N838);
nor NOR4 (N1640, N1633, N837, N298, N1483);
nand NAND4 (N1641, N1621, N965, N1266, N1090);
xor XOR2 (N1642, N1631, N1089);
and AND3 (N1643, N1639, N817, N20);
and AND2 (N1644, N1642, N1152);
buf BUF1 (N1645, N1627);
xor XOR2 (N1646, N1645, N1503);
buf BUF1 (N1647, N1625);
nand NAND3 (N1648, N1646, N246, N1273);
xor XOR2 (N1649, N1634, N163);
xor XOR2 (N1650, N1640, N1440);
nand NAND4 (N1651, N1644, N180, N267, N710);
or OR2 (N1652, N1648, N123);
xor XOR2 (N1653, N1647, N297);
buf BUF1 (N1654, N1636);
nor NOR3 (N1655, N1653, N217, N1403);
and AND2 (N1656, N1649, N549);
xor XOR2 (N1657, N1651, N255);
nand NAND4 (N1658, N1657, N793, N229, N210);
xor XOR2 (N1659, N1643, N745);
xor XOR2 (N1660, N1650, N1655);
buf BUF1 (N1661, N906);
not NOT1 (N1662, N1652);
buf BUF1 (N1663, N1662);
nor NOR3 (N1664, N1660, N1607, N237);
xor XOR2 (N1665, N1641, N103);
or OR2 (N1666, N1661, N242);
xor XOR2 (N1667, N1638, N1108);
not NOT1 (N1668, N1632);
not NOT1 (N1669, N1659);
and AND2 (N1670, N1658, N757);
xor XOR2 (N1671, N1667, N948);
not NOT1 (N1672, N1663);
nor NOR4 (N1673, N1666, N1193, N259, N226);
nor NOR4 (N1674, N1672, N719, N1588, N581);
nand NAND4 (N1675, N1670, N1404, N489, N734);
or OR3 (N1676, N1669, N153, N1098);
not NOT1 (N1677, N1654);
buf BUF1 (N1678, N1677);
and AND4 (N1679, N1674, N1619, N983, N786);
not NOT1 (N1680, N1664);
and AND4 (N1681, N1656, N405, N583, N278);
xor XOR2 (N1682, N1675, N1673);
nand NAND2 (N1683, N1278, N544);
xor XOR2 (N1684, N1671, N835);
nand NAND2 (N1685, N1665, N1675);
xor XOR2 (N1686, N1680, N1125);
buf BUF1 (N1687, N1681);
buf BUF1 (N1688, N1686);
nor NOR4 (N1689, N1668, N780, N1614, N394);
and AND3 (N1690, N1685, N1190, N38);
buf BUF1 (N1691, N1683);
xor XOR2 (N1692, N1689, N914);
not NOT1 (N1693, N1687);
or OR4 (N1694, N1693, N1099, N1408, N646);
nand NAND2 (N1695, N1684, N334);
nand NAND2 (N1696, N1688, N565);
buf BUF1 (N1697, N1678);
xor XOR2 (N1698, N1695, N47);
xor XOR2 (N1699, N1682, N1228);
buf BUF1 (N1700, N1676);
or OR2 (N1701, N1691, N879);
not NOT1 (N1702, N1698);
and AND4 (N1703, N1694, N759, N1142, N920);
nand NAND3 (N1704, N1696, N1135, N1590);
nor NOR4 (N1705, N1703, N543, N774, N323);
not NOT1 (N1706, N1704);
nor NOR4 (N1707, N1706, N203, N1473, N1012);
and AND3 (N1708, N1707, N1455, N921);
or OR2 (N1709, N1690, N1533);
buf BUF1 (N1710, N1709);
xor XOR2 (N1711, N1710, N1383);
and AND3 (N1712, N1700, N1469, N1647);
and AND3 (N1713, N1708, N333, N1349);
buf BUF1 (N1714, N1679);
nor NOR3 (N1715, N1701, N1608, N92);
xor XOR2 (N1716, N1712, N729);
buf BUF1 (N1717, N1715);
xor XOR2 (N1718, N1705, N774);
xor XOR2 (N1719, N1697, N1061);
nor NOR4 (N1720, N1692, N331, N234, N644);
buf BUF1 (N1721, N1711);
nor NOR4 (N1722, N1718, N528, N356, N765);
xor XOR2 (N1723, N1716, N1669);
xor XOR2 (N1724, N1719, N111);
nor NOR2 (N1725, N1721, N595);
or OR2 (N1726, N1724, N731);
buf BUF1 (N1727, N1725);
and AND4 (N1728, N1699, N376, N31, N60);
buf BUF1 (N1729, N1713);
or OR4 (N1730, N1720, N126, N485, N1254);
or OR4 (N1731, N1730, N1342, N596, N1264);
xor XOR2 (N1732, N1723, N395);
nor NOR2 (N1733, N1702, N1181);
not NOT1 (N1734, N1726);
and AND2 (N1735, N1729, N1557);
buf BUF1 (N1736, N1731);
xor XOR2 (N1737, N1733, N104);
nand NAND2 (N1738, N1722, N1080);
nand NAND2 (N1739, N1728, N1214);
and AND3 (N1740, N1727, N771, N1576);
xor XOR2 (N1741, N1738, N755);
nor NOR2 (N1742, N1734, N357);
not NOT1 (N1743, N1736);
nor NOR4 (N1744, N1742, N1742, N323, N254);
or OR3 (N1745, N1737, N703, N806);
and AND2 (N1746, N1732, N247);
xor XOR2 (N1747, N1717, N1553);
and AND4 (N1748, N1747, N163, N741, N1259);
not NOT1 (N1749, N1741);
buf BUF1 (N1750, N1743);
nand NAND2 (N1751, N1714, N185);
nor NOR3 (N1752, N1735, N1102, N773);
nor NOR3 (N1753, N1745, N846, N941);
nand NAND3 (N1754, N1740, N803, N1140);
nand NAND2 (N1755, N1750, N1283);
nand NAND3 (N1756, N1749, N1720, N577);
or OR2 (N1757, N1756, N317);
nor NOR3 (N1758, N1751, N380, N1506);
nor NOR3 (N1759, N1758, N1413, N1555);
nand NAND2 (N1760, N1752, N902);
xor XOR2 (N1761, N1760, N328);
buf BUF1 (N1762, N1748);
not NOT1 (N1763, N1755);
and AND4 (N1764, N1759, N441, N1598, N739);
nand NAND4 (N1765, N1753, N1107, N377, N403);
not NOT1 (N1766, N1761);
nor NOR3 (N1767, N1764, N1732, N611);
not NOT1 (N1768, N1762);
nand NAND3 (N1769, N1754, N940, N1704);
nand NAND3 (N1770, N1746, N1235, N52);
buf BUF1 (N1771, N1769);
and AND2 (N1772, N1739, N873);
or OR3 (N1773, N1768, N95, N1511);
nand NAND2 (N1774, N1772, N370);
nor NOR4 (N1775, N1771, N128, N53, N1711);
xor XOR2 (N1776, N1766, N834);
buf BUF1 (N1777, N1763);
not NOT1 (N1778, N1777);
buf BUF1 (N1779, N1778);
nor NOR4 (N1780, N1774, N274, N591, N563);
nor NOR4 (N1781, N1776, N119, N313, N660);
or OR2 (N1782, N1757, N56);
buf BUF1 (N1783, N1782);
not NOT1 (N1784, N1781);
buf BUF1 (N1785, N1783);
nor NOR2 (N1786, N1780, N1588);
xor XOR2 (N1787, N1784, N1689);
nand NAND4 (N1788, N1779, N37, N880, N332);
nand NAND2 (N1789, N1785, N1342);
or OR2 (N1790, N1765, N1688);
nor NOR4 (N1791, N1773, N483, N903, N1372);
nand NAND2 (N1792, N1791, N723);
or OR4 (N1793, N1790, N609, N1247, N1773);
nand NAND4 (N1794, N1788, N1370, N517, N305);
nand NAND2 (N1795, N1794, N698);
or OR3 (N1796, N1775, N1495, N635);
nor NOR4 (N1797, N1795, N9, N657, N547);
nor NOR4 (N1798, N1796, N168, N251, N189);
nor NOR4 (N1799, N1793, N1394, N103, N942);
buf BUF1 (N1800, N1792);
not NOT1 (N1801, N1789);
or OR4 (N1802, N1801, N292, N227, N276);
not NOT1 (N1803, N1798);
and AND4 (N1804, N1799, N133, N1332, N1625);
buf BUF1 (N1805, N1797);
xor XOR2 (N1806, N1800, N768);
and AND3 (N1807, N1804, N310, N1722);
nand NAND2 (N1808, N1767, N1297);
not NOT1 (N1809, N1786);
or OR3 (N1810, N1787, N851, N1128);
and AND4 (N1811, N1802, N1094, N529, N317);
buf BUF1 (N1812, N1770);
and AND2 (N1813, N1803, N1412);
xor XOR2 (N1814, N1744, N121);
nand NAND3 (N1815, N1812, N225, N1673);
and AND2 (N1816, N1811, N43);
buf BUF1 (N1817, N1810);
nor NOR3 (N1818, N1816, N1360, N1618);
xor XOR2 (N1819, N1805, N590);
or OR2 (N1820, N1815, N318);
nand NAND4 (N1821, N1809, N1768, N1393, N1630);
or OR3 (N1822, N1813, N353, N1201);
nand NAND4 (N1823, N1819, N413, N1595, N1112);
xor XOR2 (N1824, N1823, N597);
xor XOR2 (N1825, N1808, N196);
nand NAND3 (N1826, N1817, N733, N141);
xor XOR2 (N1827, N1820, N715);
xor XOR2 (N1828, N1826, N269);
nor NOR4 (N1829, N1827, N653, N1307, N196);
not NOT1 (N1830, N1821);
not NOT1 (N1831, N1814);
nand NAND3 (N1832, N1829, N191, N41);
buf BUF1 (N1833, N1824);
not NOT1 (N1834, N1833);
and AND3 (N1835, N1828, N931, N217);
buf BUF1 (N1836, N1818);
not NOT1 (N1837, N1822);
not NOT1 (N1838, N1825);
or OR2 (N1839, N1806, N854);
or OR3 (N1840, N1807, N946, N17);
or OR2 (N1841, N1838, N1594);
nand NAND3 (N1842, N1830, N1635, N1813);
not NOT1 (N1843, N1839);
and AND2 (N1844, N1837, N1215);
or OR2 (N1845, N1841, N72);
nand NAND3 (N1846, N1836, N712, N61);
nor NOR4 (N1847, N1845, N267, N1522, N1620);
not NOT1 (N1848, N1831);
nor NOR2 (N1849, N1847, N1666);
nor NOR4 (N1850, N1849, N1030, N667, N891);
not NOT1 (N1851, N1846);
and AND2 (N1852, N1844, N1599);
nand NAND2 (N1853, N1848, N1621);
or OR3 (N1854, N1843, N1680, N190);
nor NOR3 (N1855, N1834, N377, N1428);
not NOT1 (N1856, N1835);
not NOT1 (N1857, N1852);
not NOT1 (N1858, N1850);
xor XOR2 (N1859, N1842, N1262);
or OR2 (N1860, N1858, N151);
or OR2 (N1861, N1856, N722);
not NOT1 (N1862, N1853);
or OR4 (N1863, N1861, N88, N1259, N235);
or OR2 (N1864, N1862, N488);
nor NOR4 (N1865, N1855, N1722, N710, N1450);
and AND2 (N1866, N1840, N1503);
buf BUF1 (N1867, N1860);
nor NOR3 (N1868, N1867, N1631, N1750);
buf BUF1 (N1869, N1832);
and AND4 (N1870, N1857, N567, N521, N1723);
buf BUF1 (N1871, N1863);
nor NOR3 (N1872, N1870, N1653, N1673);
nor NOR4 (N1873, N1865, N537, N1612, N1523);
xor XOR2 (N1874, N1851, N18);
nand NAND2 (N1875, N1871, N987);
and AND4 (N1876, N1869, N675, N1069, N1726);
buf BUF1 (N1877, N1875);
nor NOR2 (N1878, N1873, N1310);
buf BUF1 (N1879, N1854);
xor XOR2 (N1880, N1879, N588);
nand NAND3 (N1881, N1872, N1000, N388);
buf BUF1 (N1882, N1864);
not NOT1 (N1883, N1868);
not NOT1 (N1884, N1866);
nand NAND2 (N1885, N1882, N262);
not NOT1 (N1886, N1885);
buf BUF1 (N1887, N1878);
not NOT1 (N1888, N1887);
xor XOR2 (N1889, N1876, N1784);
not NOT1 (N1890, N1881);
and AND2 (N1891, N1888, N1503);
buf BUF1 (N1892, N1874);
nor NOR3 (N1893, N1891, N119, N1179);
xor XOR2 (N1894, N1890, N165);
not NOT1 (N1895, N1892);
nand NAND4 (N1896, N1859, N1862, N1101, N182);
nor NOR2 (N1897, N1893, N1641);
and AND4 (N1898, N1897, N1481, N1391, N1027);
and AND2 (N1899, N1880, N1543);
and AND4 (N1900, N1895, N657, N926, N1441);
buf BUF1 (N1901, N1886);
not NOT1 (N1902, N1894);
and AND4 (N1903, N1884, N1293, N1388, N1437);
nor NOR4 (N1904, N1898, N413, N1713, N114);
buf BUF1 (N1905, N1901);
not NOT1 (N1906, N1896);
or OR2 (N1907, N1902, N217);
buf BUF1 (N1908, N1900);
and AND3 (N1909, N1883, N706, N528);
not NOT1 (N1910, N1877);
and AND4 (N1911, N1908, N1417, N658, N169);
buf BUF1 (N1912, N1906);
nand NAND3 (N1913, N1912, N980, N906);
buf BUF1 (N1914, N1910);
and AND2 (N1915, N1914, N463);
or OR2 (N1916, N1907, N800);
nor NOR4 (N1917, N1903, N128, N1488, N1665);
not NOT1 (N1918, N1915);
nand NAND2 (N1919, N1899, N1335);
nand NAND3 (N1920, N1909, N199, N1438);
not NOT1 (N1921, N1917);
xor XOR2 (N1922, N1889, N118);
nor NOR2 (N1923, N1922, N889);
xor XOR2 (N1924, N1921, N1549);
or OR2 (N1925, N1916, N1620);
and AND3 (N1926, N1925, N1873, N1876);
and AND3 (N1927, N1913, N784, N1198);
not NOT1 (N1928, N1926);
and AND2 (N1929, N1911, N171);
nor NOR4 (N1930, N1918, N1109, N1419, N246);
buf BUF1 (N1931, N1905);
and AND4 (N1932, N1920, N1921, N1885, N1396);
nand NAND2 (N1933, N1919, N1026);
and AND2 (N1934, N1904, N984);
xor XOR2 (N1935, N1924, N1593);
buf BUF1 (N1936, N1934);
and AND2 (N1937, N1930, N268);
xor XOR2 (N1938, N1927, N791);
and AND2 (N1939, N1931, N1142);
not NOT1 (N1940, N1937);
xor XOR2 (N1941, N1923, N789);
nor NOR2 (N1942, N1939, N499);
not NOT1 (N1943, N1935);
not NOT1 (N1944, N1929);
nand NAND2 (N1945, N1938, N1796);
nor NOR4 (N1946, N1942, N445, N693, N1725);
nand NAND4 (N1947, N1936, N1830, N413, N508);
not NOT1 (N1948, N1928);
xor XOR2 (N1949, N1932, N822);
or OR3 (N1950, N1948, N1332, N335);
nor NOR2 (N1951, N1940, N1594);
nor NOR4 (N1952, N1941, N834, N472, N1079);
xor XOR2 (N1953, N1945, N1894);
buf BUF1 (N1954, N1933);
buf BUF1 (N1955, N1950);
buf BUF1 (N1956, N1944);
or OR3 (N1957, N1956, N252, N581);
xor XOR2 (N1958, N1953, N131);
xor XOR2 (N1959, N1952, N83);
xor XOR2 (N1960, N1943, N1918);
not NOT1 (N1961, N1959);
nor NOR2 (N1962, N1954, N1448);
and AND4 (N1963, N1946, N336, N369, N1277);
not NOT1 (N1964, N1949);
not NOT1 (N1965, N1961);
xor XOR2 (N1966, N1947, N1079);
xor XOR2 (N1967, N1965, N353);
xor XOR2 (N1968, N1962, N505);
or OR3 (N1969, N1966, N1592, N321);
nand NAND3 (N1970, N1964, N800, N1923);
and AND4 (N1971, N1968, N1679, N1764, N1527);
not NOT1 (N1972, N1951);
xor XOR2 (N1973, N1969, N1024);
or OR2 (N1974, N1957, N1848);
not NOT1 (N1975, N1973);
not NOT1 (N1976, N1971);
nand NAND4 (N1977, N1955, N213, N1347, N746);
nand NAND2 (N1978, N1975, N1397);
xor XOR2 (N1979, N1960, N764);
and AND3 (N1980, N1967, N1231, N741);
not NOT1 (N1981, N1978);
nand NAND3 (N1982, N1981, N85, N1483);
buf BUF1 (N1983, N1963);
buf BUF1 (N1984, N1976);
nand NAND4 (N1985, N1979, N80, N1041, N38);
and AND2 (N1986, N1972, N1816);
or OR3 (N1987, N1984, N676, N933);
nand NAND4 (N1988, N1977, N1802, N79, N631);
xor XOR2 (N1989, N1985, N276);
buf BUF1 (N1990, N1989);
and AND3 (N1991, N1970, N1305, N299);
or OR2 (N1992, N1988, N457);
not NOT1 (N1993, N1991);
nor NOR2 (N1994, N1986, N1149);
nand NAND4 (N1995, N1990, N632, N69, N1188);
or OR4 (N1996, N1992, N149, N709, N1391);
xor XOR2 (N1997, N1987, N1093);
and AND3 (N1998, N1958, N182, N914);
buf BUF1 (N1999, N1994);
not NOT1 (N2000, N1997);
nor NOR3 (N2001, N1996, N1111, N676);
nor NOR2 (N2002, N2000, N1058);
nor NOR2 (N2003, N1974, N47);
or OR3 (N2004, N1983, N297, N209);
buf BUF1 (N2005, N1980);
and AND3 (N2006, N2005, N909, N573);
not NOT1 (N2007, N2002);
nand NAND2 (N2008, N1995, N1508);
xor XOR2 (N2009, N2008, N772);
nor NOR4 (N2010, N2009, N1563, N1858, N1042);
xor XOR2 (N2011, N1999, N738);
buf BUF1 (N2012, N1982);
nand NAND3 (N2013, N2006, N991, N1970);
xor XOR2 (N2014, N2003, N1625);
xor XOR2 (N2015, N2004, N1599);
nor NOR2 (N2016, N2010, N778);
xor XOR2 (N2017, N2007, N913);
not NOT1 (N2018, N2011);
nor NOR3 (N2019, N2015, N1989, N1861);
and AND3 (N2020, N2001, N1725, N908);
and AND4 (N2021, N2016, N215, N1868, N539);
xor XOR2 (N2022, N2014, N1788);
nand NAND3 (N2023, N2022, N557, N1187);
nand NAND3 (N2024, N2017, N126, N657);
nor NOR2 (N2025, N2012, N784);
and AND4 (N2026, N2019, N311, N2000, N207);
buf BUF1 (N2027, N1998);
xor XOR2 (N2028, N2020, N919);
xor XOR2 (N2029, N2028, N717);
not NOT1 (N2030, N2025);
nand NAND4 (N2031, N2027, N1923, N18, N741);
xor XOR2 (N2032, N2031, N1529);
xor XOR2 (N2033, N1993, N56);
or OR4 (N2034, N2013, N1504, N1697, N1737);
buf BUF1 (N2035, N2030);
buf BUF1 (N2036, N2018);
nor NOR4 (N2037, N2035, N749, N809, N489);
and AND4 (N2038, N2034, N746, N1123, N892);
xor XOR2 (N2039, N2024, N963);
buf BUF1 (N2040, N2032);
xor XOR2 (N2041, N2038, N1400);
and AND2 (N2042, N2023, N245);
buf BUF1 (N2043, N2039);
nand NAND3 (N2044, N2026, N101, N1794);
and AND4 (N2045, N2044, N1483, N1862, N1700);
nand NAND4 (N2046, N2040, N489, N356, N466);
not NOT1 (N2047, N2033);
buf BUF1 (N2048, N2045);
nor NOR3 (N2049, N2037, N1184, N1153);
or OR2 (N2050, N2043, N646);
not NOT1 (N2051, N2042);
nor NOR4 (N2052, N2048, N892, N591, N1108);
or OR2 (N2053, N2049, N127);
and AND2 (N2054, N2021, N1682);
and AND3 (N2055, N2050, N287, N1578);
xor XOR2 (N2056, N2052, N337);
xor XOR2 (N2057, N2053, N1542);
or OR4 (N2058, N2054, N795, N964, N61);
or OR3 (N2059, N2041, N1759, N250);
and AND2 (N2060, N2051, N961);
and AND2 (N2061, N2060, N631);
not NOT1 (N2062, N2036);
buf BUF1 (N2063, N2055);
not NOT1 (N2064, N2047);
or OR4 (N2065, N2062, N1201, N404, N1323);
nand NAND4 (N2066, N2059, N1369, N1019, N1807);
nand NAND2 (N2067, N2064, N701);
or OR3 (N2068, N2058, N518, N263);
nor NOR2 (N2069, N2046, N165);
and AND4 (N2070, N2067, N963, N356, N136);
nand NAND4 (N2071, N2070, N732, N575, N1803);
xor XOR2 (N2072, N2071, N1806);
or OR3 (N2073, N2057, N1711, N814);
nor NOR3 (N2074, N2063, N535, N1028);
not NOT1 (N2075, N2073);
not NOT1 (N2076, N2056);
not NOT1 (N2077, N2029);
and AND2 (N2078, N2066, N1652);
and AND4 (N2079, N2075, N396, N1596, N1456);
xor XOR2 (N2080, N2079, N775);
nor NOR4 (N2081, N2061, N2071, N2025, N1675);
nor NOR2 (N2082, N2074, N419);
xor XOR2 (N2083, N2080, N402);
not NOT1 (N2084, N2081);
nand NAND4 (N2085, N2083, N641, N1253, N346);
not NOT1 (N2086, N2068);
nand NAND3 (N2087, N2065, N1467, N937);
not NOT1 (N2088, N2087);
and AND2 (N2089, N2082, N1761);
or OR2 (N2090, N2077, N606);
buf BUF1 (N2091, N2090);
and AND2 (N2092, N2084, N456);
or OR4 (N2093, N2078, N254, N371, N1618);
nor NOR3 (N2094, N2092, N780, N262);
not NOT1 (N2095, N2094);
not NOT1 (N2096, N2093);
xor XOR2 (N2097, N2069, N1433);
xor XOR2 (N2098, N2088, N606);
or OR3 (N2099, N2097, N1633, N319);
nand NAND2 (N2100, N2089, N1751);
nor NOR4 (N2101, N2099, N482, N1380, N1661);
nor NOR4 (N2102, N2095, N1849, N218, N227);
or OR3 (N2103, N2100, N44, N1012);
nor NOR4 (N2104, N2096, N1339, N1191, N670);
nand NAND2 (N2105, N2086, N1999);
nor NOR4 (N2106, N2105, N1211, N1981, N845);
nor NOR2 (N2107, N2103, N176);
or OR2 (N2108, N2101, N997);
nor NOR4 (N2109, N2098, N1127, N606, N1996);
nor NOR3 (N2110, N2072, N332, N468);
and AND2 (N2111, N2091, N1138);
xor XOR2 (N2112, N2108, N325);
and AND2 (N2113, N2110, N1355);
nand NAND4 (N2114, N2113, N1790, N523, N1542);
xor XOR2 (N2115, N2104, N1585);
nor NOR3 (N2116, N2107, N1828, N1357);
buf BUF1 (N2117, N2112);
buf BUF1 (N2118, N2102);
xor XOR2 (N2119, N2076, N972);
nor NOR4 (N2120, N2114, N938, N82, N477);
nor NOR4 (N2121, N2085, N2026, N1395, N533);
nand NAND4 (N2122, N2119, N1118, N1737, N19);
nand NAND2 (N2123, N2118, N465);
not NOT1 (N2124, N2111);
nor NOR2 (N2125, N2117, N251);
or OR2 (N2126, N2109, N1445);
not NOT1 (N2127, N2115);
xor XOR2 (N2128, N2116, N1501);
nor NOR2 (N2129, N2121, N1555);
and AND2 (N2130, N2122, N2049);
xor XOR2 (N2131, N2124, N1500);
not NOT1 (N2132, N2106);
nand NAND3 (N2133, N2128, N1202, N210);
and AND3 (N2134, N2123, N1640, N1492);
not NOT1 (N2135, N2134);
buf BUF1 (N2136, N2127);
nor NOR4 (N2137, N2136, N1417, N1414, N1177);
and AND3 (N2138, N2120, N1171, N715);
or OR3 (N2139, N2133, N1771, N1541);
and AND2 (N2140, N2126, N1530);
and AND2 (N2141, N2138, N1003);
xor XOR2 (N2142, N2140, N1149);
nand NAND4 (N2143, N2142, N944, N883, N1020);
nand NAND4 (N2144, N2129, N750, N1721, N200);
or OR4 (N2145, N2131, N1141, N1789, N848);
nor NOR3 (N2146, N2143, N1086, N2021);
xor XOR2 (N2147, N2135, N1357);
xor XOR2 (N2148, N2146, N1459);
nor NOR4 (N2149, N2145, N81, N484, N884);
and AND4 (N2150, N2139, N1843, N1766, N256);
nand NAND3 (N2151, N2148, N482, N1474);
xor XOR2 (N2152, N2147, N1218);
or OR3 (N2153, N2130, N939, N1911);
not NOT1 (N2154, N2132);
or OR4 (N2155, N2149, N855, N1570, N1765);
or OR3 (N2156, N2141, N1863, N1293);
xor XOR2 (N2157, N2137, N1781);
or OR2 (N2158, N2125, N1958);
nand NAND3 (N2159, N2153, N568, N2104);
nand NAND3 (N2160, N2155, N464, N1987);
buf BUF1 (N2161, N2160);
or OR2 (N2162, N2152, N235);
buf BUF1 (N2163, N2151);
not NOT1 (N2164, N2162);
or OR4 (N2165, N2157, N1109, N1406, N1446);
and AND2 (N2166, N2144, N485);
buf BUF1 (N2167, N2161);
buf BUF1 (N2168, N2164);
not NOT1 (N2169, N2156);
and AND4 (N2170, N2166, N1892, N900, N489);
xor XOR2 (N2171, N2150, N1803);
nor NOR3 (N2172, N2154, N200, N2025);
not NOT1 (N2173, N2171);
and AND2 (N2174, N2173, N506);
and AND4 (N2175, N2168, N1736, N401, N778);
xor XOR2 (N2176, N2159, N1965);
nand NAND3 (N2177, N2167, N60, N1481);
nor NOR2 (N2178, N2174, N1492);
nand NAND4 (N2179, N2178, N2101, N1028, N1875);
xor XOR2 (N2180, N2172, N759);
and AND4 (N2181, N2163, N1713, N94, N2110);
nor NOR4 (N2182, N2176, N2155, N80, N242);
nand NAND4 (N2183, N2158, N177, N393, N489);
buf BUF1 (N2184, N2181);
buf BUF1 (N2185, N2165);
nand NAND2 (N2186, N2175, N934);
nand NAND3 (N2187, N2184, N417, N1679);
nand NAND3 (N2188, N2187, N832, N2099);
not NOT1 (N2189, N2170);
xor XOR2 (N2190, N2182, N644);
not NOT1 (N2191, N2180);
buf BUF1 (N2192, N2183);
xor XOR2 (N2193, N2185, N436);
nand NAND2 (N2194, N2193, N1414);
not NOT1 (N2195, N2192);
and AND4 (N2196, N2179, N218, N1851, N1634);
or OR3 (N2197, N2191, N852, N1886);
nand NAND2 (N2198, N2197, N705);
not NOT1 (N2199, N2169);
nor NOR3 (N2200, N2189, N1737, N1879);
nand NAND4 (N2201, N2190, N1211, N1558, N2012);
and AND3 (N2202, N2198, N164, N664);
buf BUF1 (N2203, N2202);
xor XOR2 (N2204, N2199, N1613);
xor XOR2 (N2205, N2195, N117);
not NOT1 (N2206, N2201);
buf BUF1 (N2207, N2196);
nor NOR3 (N2208, N2186, N2154, N1766);
buf BUF1 (N2209, N2205);
nand NAND4 (N2210, N2204, N1766, N666, N193);
buf BUF1 (N2211, N2210);
not NOT1 (N2212, N2207);
xor XOR2 (N2213, N2209, N1753);
buf BUF1 (N2214, N2200);
buf BUF1 (N2215, N2188);
nor NOR3 (N2216, N2211, N1134, N1350);
and AND4 (N2217, N2206, N975, N1575, N46);
or OR3 (N2218, N2203, N908, N1887);
and AND3 (N2219, N2208, N691, N1170);
not NOT1 (N2220, N2216);
or OR4 (N2221, N2218, N1663, N669, N1844);
xor XOR2 (N2222, N2194, N510);
xor XOR2 (N2223, N2220, N1862);
nand NAND3 (N2224, N2177, N1588, N962);
nand NAND3 (N2225, N2214, N959, N709);
not NOT1 (N2226, N2224);
or OR2 (N2227, N2225, N999);
and AND3 (N2228, N2213, N1954, N1570);
and AND3 (N2229, N2226, N2083, N1707);
and AND4 (N2230, N2212, N388, N880, N478);
nor NOR2 (N2231, N2229, N41);
xor XOR2 (N2232, N2227, N2155);
or OR3 (N2233, N2217, N2057, N994);
nor NOR3 (N2234, N2230, N685, N996);
xor XOR2 (N2235, N2221, N616);
buf BUF1 (N2236, N2228);
and AND4 (N2237, N2219, N815, N2087, N759);
nor NOR4 (N2238, N2223, N154, N1880, N962);
buf BUF1 (N2239, N2237);
not NOT1 (N2240, N2231);
not NOT1 (N2241, N2235);
xor XOR2 (N2242, N2238, N44);
buf BUF1 (N2243, N2240);
nand NAND4 (N2244, N2241, N30, N1209, N2105);
nand NAND2 (N2245, N2243, N301);
and AND3 (N2246, N2232, N1654, N1914);
or OR2 (N2247, N2242, N1597);
nor NOR3 (N2248, N2245, N1129, N1376);
or OR2 (N2249, N2247, N1768);
not NOT1 (N2250, N2244);
buf BUF1 (N2251, N2236);
nor NOR4 (N2252, N2233, N1968, N1564, N1824);
buf BUF1 (N2253, N2252);
buf BUF1 (N2254, N2250);
xor XOR2 (N2255, N2248, N1136);
nor NOR4 (N2256, N2246, N534, N1600, N210);
or OR4 (N2257, N2256, N877, N602, N244);
and AND3 (N2258, N2255, N1830, N2038);
or OR3 (N2259, N2234, N1062, N32);
xor XOR2 (N2260, N2249, N396);
not NOT1 (N2261, N2257);
and AND4 (N2262, N2253, N729, N268, N2024);
xor XOR2 (N2263, N2262, N683);
nand NAND4 (N2264, N2254, N372, N1499, N2079);
xor XOR2 (N2265, N2259, N2141);
buf BUF1 (N2266, N2258);
not NOT1 (N2267, N2222);
and AND2 (N2268, N2264, N561);
xor XOR2 (N2269, N2268, N2004);
not NOT1 (N2270, N2215);
or OR3 (N2271, N2267, N1367, N1171);
not NOT1 (N2272, N2260);
xor XOR2 (N2273, N2263, N1269);
nand NAND4 (N2274, N2271, N751, N534, N1078);
and AND2 (N2275, N2272, N167);
buf BUF1 (N2276, N2274);
buf BUF1 (N2277, N2273);
buf BUF1 (N2278, N2275);
buf BUF1 (N2279, N2265);
and AND3 (N2280, N2279, N2032, N2057);
nor NOR3 (N2281, N2280, N1824, N630);
or OR3 (N2282, N2278, N232, N1955);
buf BUF1 (N2283, N2281);
and AND2 (N2284, N2239, N494);
or OR4 (N2285, N2269, N934, N700, N475);
nand NAND2 (N2286, N2284, N2189);
nand NAND2 (N2287, N2285, N2130);
xor XOR2 (N2288, N2261, N1554);
nor NOR2 (N2289, N2282, N2268);
nand NAND2 (N2290, N2283, N858);
nor NOR4 (N2291, N2286, N988, N800, N2217);
nor NOR4 (N2292, N2276, N1069, N2208, N2005);
buf BUF1 (N2293, N2266);
xor XOR2 (N2294, N2277, N1271);
nor NOR3 (N2295, N2290, N870, N1319);
and AND2 (N2296, N2287, N1617);
buf BUF1 (N2297, N2270);
and AND4 (N2298, N2292, N1616, N188, N202);
nor NOR4 (N2299, N2289, N222, N1062, N1936);
not NOT1 (N2300, N2298);
nand NAND2 (N2301, N2295, N47);
and AND3 (N2302, N2293, N566, N1494);
buf BUF1 (N2303, N2297);
and AND4 (N2304, N2251, N1054, N955, N833);
xor XOR2 (N2305, N2296, N1465);
or OR2 (N2306, N2299, N129);
buf BUF1 (N2307, N2306);
or OR2 (N2308, N2288, N1832);
and AND4 (N2309, N2303, N1929, N2222, N629);
not NOT1 (N2310, N2309);
and AND3 (N2311, N2307, N1447, N327);
nor NOR3 (N2312, N2301, N2302, N1316);
nand NAND4 (N2313, N2149, N229, N396, N1382);
not NOT1 (N2314, N2310);
not NOT1 (N2315, N2304);
not NOT1 (N2316, N2315);
or OR3 (N2317, N2316, N426, N799);
and AND3 (N2318, N2300, N1683, N1295);
xor XOR2 (N2319, N2311, N444);
not NOT1 (N2320, N2313);
xor XOR2 (N2321, N2317, N713);
and AND2 (N2322, N2305, N1938);
buf BUF1 (N2323, N2322);
buf BUF1 (N2324, N2320);
nor NOR4 (N2325, N2308, N629, N1323, N1016);
and AND3 (N2326, N2294, N1048, N992);
or OR2 (N2327, N2323, N54);
or OR3 (N2328, N2321, N2071, N1618);
and AND2 (N2329, N2291, N917);
nor NOR2 (N2330, N2326, N80);
or OR3 (N2331, N2329, N560, N1848);
buf BUF1 (N2332, N2328);
nand NAND4 (N2333, N2312, N2180, N550, N2090);
buf BUF1 (N2334, N2319);
not NOT1 (N2335, N2331);
and AND4 (N2336, N2324, N1675, N2197, N591);
or OR2 (N2337, N2336, N1339);
or OR4 (N2338, N2327, N1813, N240, N574);
xor XOR2 (N2339, N2332, N1370);
xor XOR2 (N2340, N2314, N2312);
buf BUF1 (N2341, N2340);
or OR4 (N2342, N2330, N1625, N1958, N977);
nand NAND2 (N2343, N2335, N1279);
nand NAND4 (N2344, N2343, N890, N318, N1549);
nand NAND3 (N2345, N2342, N820, N956);
xor XOR2 (N2346, N2325, N1716);
buf BUF1 (N2347, N2318);
and AND2 (N2348, N2341, N2177);
nand NAND2 (N2349, N2334, N1438);
nor NOR4 (N2350, N2344, N1959, N1493, N876);
or OR3 (N2351, N2333, N1791, N964);
nand NAND3 (N2352, N2347, N544, N668);
buf BUF1 (N2353, N2337);
not NOT1 (N2354, N2350);
xor XOR2 (N2355, N2352, N2229);
or OR3 (N2356, N2338, N951, N242);
nand NAND4 (N2357, N2356, N1393, N748, N1184);
nor NOR2 (N2358, N2351, N2132);
nor NOR4 (N2359, N2354, N2283, N1590, N694);
nor NOR3 (N2360, N2355, N525, N163);
nand NAND2 (N2361, N2353, N1206);
xor XOR2 (N2362, N2345, N2211);
and AND4 (N2363, N2359, N488, N722, N1275);
xor XOR2 (N2364, N2363, N1411);
nor NOR4 (N2365, N2357, N628, N1934, N2233);
or OR4 (N2366, N2362, N1712, N677, N816);
nand NAND4 (N2367, N2364, N451, N717, N886);
buf BUF1 (N2368, N2346);
or OR2 (N2369, N2349, N1005);
or OR3 (N2370, N2368, N2358, N840);
not NOT1 (N2371, N147);
xor XOR2 (N2372, N2365, N470);
and AND2 (N2373, N2371, N823);
nor NOR2 (N2374, N2370, N801);
nand NAND2 (N2375, N2339, N1410);
or OR4 (N2376, N2348, N1370, N1992, N2327);
xor XOR2 (N2377, N2376, N184);
nand NAND4 (N2378, N2375, N1390, N313, N241);
nand NAND3 (N2379, N2372, N2293, N1489);
or OR2 (N2380, N2367, N302);
nor NOR4 (N2381, N2380, N924, N428, N708);
not NOT1 (N2382, N2378);
or OR3 (N2383, N2369, N2147, N308);
nor NOR2 (N2384, N2366, N367);
nand NAND4 (N2385, N2381, N1197, N2116, N1814);
nand NAND4 (N2386, N2379, N1621, N1329, N1455);
xor XOR2 (N2387, N2361, N2246);
not NOT1 (N2388, N2374);
buf BUF1 (N2389, N2386);
not NOT1 (N2390, N2389);
and AND3 (N2391, N2387, N1732, N2362);
xor XOR2 (N2392, N2373, N2082);
or OR2 (N2393, N2385, N647);
or OR4 (N2394, N2392, N2134, N160, N1523);
nor NOR3 (N2395, N2377, N451, N397);
buf BUF1 (N2396, N2360);
nor NOR4 (N2397, N2395, N2089, N1122, N1893);
and AND2 (N2398, N2396, N1649);
or OR4 (N2399, N2390, N1368, N1777, N1928);
buf BUF1 (N2400, N2399);
buf BUF1 (N2401, N2393);
xor XOR2 (N2402, N2383, N578);
xor XOR2 (N2403, N2384, N2055);
or OR4 (N2404, N2394, N1811, N1029, N1111);
nand NAND3 (N2405, N2388, N1431, N2077);
nand NAND2 (N2406, N2398, N152);
or OR3 (N2407, N2403, N1083, N1708);
and AND4 (N2408, N2382, N1363, N1596, N1286);
xor XOR2 (N2409, N2397, N414);
xor XOR2 (N2410, N2391, N488);
xor XOR2 (N2411, N2407, N1737);
and AND3 (N2412, N2411, N1706, N1047);
nor NOR2 (N2413, N2408, N1928);
and AND4 (N2414, N2400, N105, N534, N1634);
xor XOR2 (N2415, N2409, N745);
xor XOR2 (N2416, N2402, N1655);
not NOT1 (N2417, N2404);
or OR4 (N2418, N2415, N563, N1826, N827);
nand NAND4 (N2419, N2401, N16, N1615, N2127);
nand NAND2 (N2420, N2416, N2114);
not NOT1 (N2421, N2406);
buf BUF1 (N2422, N2405);
and AND4 (N2423, N2413, N1660, N290, N897);
and AND2 (N2424, N2421, N324);
not NOT1 (N2425, N2419);
nor NOR4 (N2426, N2410, N1012, N853, N1709);
or OR3 (N2427, N2422, N1108, N1705);
or OR3 (N2428, N2424, N2378, N1295);
nand NAND2 (N2429, N2418, N998);
nand NAND2 (N2430, N2420, N453);
or OR3 (N2431, N2417, N1221, N1756);
not NOT1 (N2432, N2430);
buf BUF1 (N2433, N2427);
nor NOR2 (N2434, N2414, N2130);
xor XOR2 (N2435, N2428, N667);
and AND2 (N2436, N2425, N2062);
nor NOR2 (N2437, N2426, N671);
xor XOR2 (N2438, N2429, N1134);
nand NAND4 (N2439, N2435, N300, N68, N1135);
or OR2 (N2440, N2423, N124);
or OR2 (N2441, N2432, N572);
not NOT1 (N2442, N2438);
buf BUF1 (N2443, N2431);
nand NAND2 (N2444, N2437, N1175);
xor XOR2 (N2445, N2434, N2239);
xor XOR2 (N2446, N2445, N578);
nor NOR3 (N2447, N2440, N2188, N319);
nor NOR4 (N2448, N2441, N1868, N2168, N198);
nor NOR2 (N2449, N2439, N368);
or OR2 (N2450, N2443, N219);
xor XOR2 (N2451, N2444, N1347);
or OR3 (N2452, N2436, N62, N1720);
xor XOR2 (N2453, N2433, N1519);
xor XOR2 (N2454, N2450, N2270);
xor XOR2 (N2455, N2451, N1030);
and AND3 (N2456, N2448, N2283, N2368);
nand NAND4 (N2457, N2453, N99, N1421, N2352);
nor NOR4 (N2458, N2457, N128, N2303, N1221);
or OR4 (N2459, N2412, N1684, N2156, N1137);
nand NAND2 (N2460, N2446, N605);
xor XOR2 (N2461, N2442, N2244);
xor XOR2 (N2462, N2461, N2442);
nand NAND2 (N2463, N2455, N866);
or OR3 (N2464, N2449, N1887, N20);
buf BUF1 (N2465, N2456);
and AND2 (N2466, N2465, N625);
buf BUF1 (N2467, N2462);
buf BUF1 (N2468, N2447);
nor NOR3 (N2469, N2460, N2062, N1588);
nor NOR2 (N2470, N2469, N1330);
nor NOR4 (N2471, N2454, N98, N560, N1280);
and AND2 (N2472, N2470, N1547);
buf BUF1 (N2473, N2467);
or OR2 (N2474, N2459, N1779);
nand NAND4 (N2475, N2458, N472, N99, N2015);
buf BUF1 (N2476, N2471);
xor XOR2 (N2477, N2452, N926);
nor NOR2 (N2478, N2464, N823);
nand NAND2 (N2479, N2474, N1646);
nor NOR4 (N2480, N2463, N632, N1310, N1849);
xor XOR2 (N2481, N2476, N870);
and AND3 (N2482, N2480, N603, N2035);
buf BUF1 (N2483, N2468);
xor XOR2 (N2484, N2483, N2003);
nand NAND2 (N2485, N2473, N1962);
nor NOR3 (N2486, N2484, N696, N76);
buf BUF1 (N2487, N2479);
and AND4 (N2488, N2478, N26, N1894, N2372);
nand NAND4 (N2489, N2487, N1108, N2168, N1572);
nor NOR2 (N2490, N2488, N46);
or OR2 (N2491, N2466, N2381);
xor XOR2 (N2492, N2486, N1089);
xor XOR2 (N2493, N2472, N1922);
nor NOR4 (N2494, N2492, N2383, N1126, N206);
xor XOR2 (N2495, N2475, N1722);
or OR3 (N2496, N2482, N75, N2495);
or OR4 (N2497, N1959, N999, N1186, N1998);
nand NAND3 (N2498, N2485, N1504, N541);
and AND3 (N2499, N2497, N1752, N763);
nor NOR3 (N2500, N2491, N891, N1554);
not NOT1 (N2501, N2490);
xor XOR2 (N2502, N2489, N2443);
xor XOR2 (N2503, N2481, N634);
not NOT1 (N2504, N2493);
and AND3 (N2505, N2496, N1518, N139);
nand NAND4 (N2506, N2477, N1710, N2021, N1062);
xor XOR2 (N2507, N2498, N583);
xor XOR2 (N2508, N2500, N2354);
xor XOR2 (N2509, N2502, N1485);
not NOT1 (N2510, N2494);
xor XOR2 (N2511, N2499, N973);
and AND2 (N2512, N2503, N1168);
or OR3 (N2513, N2501, N329, N222);
nor NOR2 (N2514, N2512, N1192);
nor NOR3 (N2515, N2505, N146, N968);
buf BUF1 (N2516, N2504);
and AND4 (N2517, N2514, N1872, N1282, N348);
not NOT1 (N2518, N2508);
and AND2 (N2519, N2518, N806);
and AND3 (N2520, N2515, N838, N84);
buf BUF1 (N2521, N2520);
or OR2 (N2522, N2509, N1255);
or OR4 (N2523, N2510, N516, N2306, N676);
not NOT1 (N2524, N2522);
nor NOR4 (N2525, N2521, N1240, N1666, N2522);
nand NAND2 (N2526, N2523, N1657);
not NOT1 (N2527, N2511);
not NOT1 (N2528, N2516);
and AND4 (N2529, N2528, N338, N666, N2005);
and AND2 (N2530, N2517, N734);
or OR2 (N2531, N2506, N2422);
nand NAND4 (N2532, N2525, N241, N2022, N1250);
not NOT1 (N2533, N2507);
buf BUF1 (N2534, N2524);
nor NOR2 (N2535, N2519, N1471);
buf BUF1 (N2536, N2532);
nor NOR2 (N2537, N2529, N445);
xor XOR2 (N2538, N2527, N677);
xor XOR2 (N2539, N2535, N2328);
not NOT1 (N2540, N2534);
or OR3 (N2541, N2530, N2023, N811);
xor XOR2 (N2542, N2538, N1094);
or OR4 (N2543, N2531, N1652, N1009, N2025);
not NOT1 (N2544, N2526);
buf BUF1 (N2545, N2513);
xor XOR2 (N2546, N2544, N1159);
nor NOR3 (N2547, N2536, N335, N1822);
xor XOR2 (N2548, N2533, N234);
and AND2 (N2549, N2548, N1925);
nor NOR4 (N2550, N2539, N2255, N2321, N342);
xor XOR2 (N2551, N2547, N1331);
xor XOR2 (N2552, N2549, N392);
xor XOR2 (N2553, N2551, N243);
nand NAND4 (N2554, N2542, N2474, N2013, N1676);
buf BUF1 (N2555, N2541);
or OR4 (N2556, N2550, N2406, N2022, N1835);
buf BUF1 (N2557, N2537);
xor XOR2 (N2558, N2554, N1639);
xor XOR2 (N2559, N2556, N1707);
not NOT1 (N2560, N2558);
not NOT1 (N2561, N2553);
nand NAND4 (N2562, N2557, N1719, N1295, N2080);
xor XOR2 (N2563, N2540, N1563);
nand NAND3 (N2564, N2545, N1307, N2233);
xor XOR2 (N2565, N2546, N2423);
not NOT1 (N2566, N2562);
or OR2 (N2567, N2559, N1674);
not NOT1 (N2568, N2564);
xor XOR2 (N2569, N2563, N1524);
nor NOR3 (N2570, N2561, N2469, N422);
buf BUF1 (N2571, N2543);
nor NOR4 (N2572, N2567, N1489, N909, N2029);
not NOT1 (N2573, N2568);
xor XOR2 (N2574, N2560, N258);
buf BUF1 (N2575, N2574);
buf BUF1 (N2576, N2552);
or OR2 (N2577, N2572, N1437);
xor XOR2 (N2578, N2573, N389);
nand NAND4 (N2579, N2577, N587, N443, N2194);
and AND2 (N2580, N2576, N1692);
nand NAND3 (N2581, N2566, N778, N401);
not NOT1 (N2582, N2578);
or OR3 (N2583, N2575, N2343, N1774);
nor NOR3 (N2584, N2565, N75, N547);
xor XOR2 (N2585, N2582, N1245);
or OR3 (N2586, N2571, N323, N1050);
not NOT1 (N2587, N2580);
nand NAND4 (N2588, N2555, N2255, N2170, N1736);
nor NOR2 (N2589, N2588, N1031);
not NOT1 (N2590, N2589);
buf BUF1 (N2591, N2579);
xor XOR2 (N2592, N2581, N2078);
nand NAND2 (N2593, N2583, N1646);
buf BUF1 (N2594, N2587);
nor NOR4 (N2595, N2584, N2586, N1206, N301);
not NOT1 (N2596, N1713);
not NOT1 (N2597, N2585);
and AND2 (N2598, N2596, N1816);
xor XOR2 (N2599, N2591, N212);
xor XOR2 (N2600, N2599, N494);
nand NAND4 (N2601, N2569, N2305, N2120, N2564);
and AND3 (N2602, N2601, N882, N934);
nor NOR3 (N2603, N2597, N563, N2211);
buf BUF1 (N2604, N2600);
buf BUF1 (N2605, N2595);
buf BUF1 (N2606, N2598);
nand NAND4 (N2607, N2605, N1492, N1834, N2595);
buf BUF1 (N2608, N2594);
nand NAND2 (N2609, N2608, N1712);
xor XOR2 (N2610, N2606, N1734);
buf BUF1 (N2611, N2593);
xor XOR2 (N2612, N2603, N1302);
not NOT1 (N2613, N2609);
xor XOR2 (N2614, N2610, N245);
not NOT1 (N2615, N2570);
and AND2 (N2616, N2604, N2049);
buf BUF1 (N2617, N2614);
not NOT1 (N2618, N2612);
and AND4 (N2619, N2616, N2251, N1826, N1087);
buf BUF1 (N2620, N2613);
or OR2 (N2621, N2617, N1346);
nand NAND4 (N2622, N2621, N2529, N1282, N1191);
nand NAND2 (N2623, N2607, N65);
nand NAND2 (N2624, N2590, N966);
or OR3 (N2625, N2619, N1757, N1822);
nor NOR4 (N2626, N2622, N1029, N2285, N848);
nand NAND3 (N2627, N2623, N1398, N2537);
nand NAND2 (N2628, N2602, N488);
buf BUF1 (N2629, N2624);
buf BUF1 (N2630, N2627);
nand NAND4 (N2631, N2615, N820, N2214, N2103);
or OR2 (N2632, N2618, N451);
nor NOR2 (N2633, N2632, N1656);
nor NOR2 (N2634, N2611, N2227);
and AND4 (N2635, N2592, N549, N1879, N125);
or OR3 (N2636, N2628, N1794, N424);
xor XOR2 (N2637, N2626, N1812);
or OR4 (N2638, N2620, N1054, N292, N195);
buf BUF1 (N2639, N2629);
xor XOR2 (N2640, N2636, N2290);
buf BUF1 (N2641, N2638);
not NOT1 (N2642, N2640);
and AND2 (N2643, N2630, N1667);
and AND2 (N2644, N2631, N544);
nand NAND4 (N2645, N2625, N1840, N1711, N1242);
buf BUF1 (N2646, N2644);
or OR3 (N2647, N2641, N2521, N1549);
not NOT1 (N2648, N2645);
not NOT1 (N2649, N2633);
nor NOR4 (N2650, N2642, N1108, N2243, N10);
xor XOR2 (N2651, N2647, N2549);
or OR3 (N2652, N2639, N1649, N799);
xor XOR2 (N2653, N2648, N1302);
nand NAND4 (N2654, N2646, N2010, N1226, N2095);
nand NAND4 (N2655, N2649, N1351, N503, N1756);
not NOT1 (N2656, N2650);
buf BUF1 (N2657, N2637);
nor NOR3 (N2658, N2651, N60, N2238);
not NOT1 (N2659, N2656);
xor XOR2 (N2660, N2652, N1030);
xor XOR2 (N2661, N2660, N555);
or OR2 (N2662, N2635, N1227);
and AND3 (N2663, N2643, N841, N803);
not NOT1 (N2664, N2661);
nand NAND4 (N2665, N2662, N2063, N1532, N758);
buf BUF1 (N2666, N2657);
nor NOR3 (N2667, N2653, N335, N443);
nor NOR4 (N2668, N2655, N1790, N1306, N530);
not NOT1 (N2669, N2664);
nor NOR4 (N2670, N2634, N1699, N2561, N2527);
nand NAND2 (N2671, N2667, N1223);
or OR2 (N2672, N2671, N2099);
and AND2 (N2673, N2668, N739);
not NOT1 (N2674, N2663);
nor NOR2 (N2675, N2670, N582);
not NOT1 (N2676, N2659);
nand NAND3 (N2677, N2675, N1304, N2349);
nand NAND4 (N2678, N2665, N2580, N1943, N2128);
or OR4 (N2679, N2677, N772, N1004, N2069);
or OR2 (N2680, N2666, N765);
nand NAND3 (N2681, N2673, N487, N2528);
buf BUF1 (N2682, N2674);
or OR4 (N2683, N2682, N1621, N2588, N910);
nand NAND3 (N2684, N2672, N240, N882);
nor NOR3 (N2685, N2658, N1758, N583);
nand NAND4 (N2686, N2676, N228, N60, N2651);
not NOT1 (N2687, N2678);
buf BUF1 (N2688, N2679);
and AND3 (N2689, N2683, N2013, N70);
nand NAND4 (N2690, N2669, N5, N1898, N639);
xor XOR2 (N2691, N2680, N1325);
and AND4 (N2692, N2685, N58, N674, N1014);
xor XOR2 (N2693, N2691, N1100);
and AND3 (N2694, N2689, N2151, N2117);
nand NAND3 (N2695, N2692, N834, N2285);
buf BUF1 (N2696, N2688);
nand NAND3 (N2697, N2654, N2115, N2006);
or OR2 (N2698, N2697, N1287);
or OR2 (N2699, N2696, N2234);
buf BUF1 (N2700, N2681);
nor NOR4 (N2701, N2699, N1205, N662, N73);
xor XOR2 (N2702, N2684, N1782);
xor XOR2 (N2703, N2698, N1696);
and AND2 (N2704, N2690, N455);
nor NOR4 (N2705, N2695, N1658, N330, N531);
nor NOR2 (N2706, N2705, N1205);
not NOT1 (N2707, N2694);
and AND4 (N2708, N2701, N2469, N223, N251);
nor NOR3 (N2709, N2702, N280, N1824);
buf BUF1 (N2710, N2709);
nand NAND3 (N2711, N2693, N1165, N1442);
nor NOR4 (N2712, N2710, N829, N2116, N624);
nor NOR3 (N2713, N2704, N1437, N1819);
or OR4 (N2714, N2713, N892, N83, N2166);
nor NOR2 (N2715, N2686, N1406);
nand NAND3 (N2716, N2712, N2431, N2283);
and AND2 (N2717, N2708, N1181);
or OR3 (N2718, N2716, N1851, N156);
not NOT1 (N2719, N2718);
xor XOR2 (N2720, N2719, N476);
nor NOR3 (N2721, N2714, N182, N230);
buf BUF1 (N2722, N2711);
xor XOR2 (N2723, N2706, N371);
nor NOR3 (N2724, N2700, N532, N1136);
nand NAND2 (N2725, N2687, N2156);
xor XOR2 (N2726, N2715, N2582);
not NOT1 (N2727, N2717);
not NOT1 (N2728, N2720);
nand NAND3 (N2729, N2725, N1879, N768);
nand NAND3 (N2730, N2723, N1725, N1560);
xor XOR2 (N2731, N2727, N601);
buf BUF1 (N2732, N2721);
xor XOR2 (N2733, N2731, N76);
buf BUF1 (N2734, N2733);
and AND4 (N2735, N2728, N401, N682, N2375);
nor NOR2 (N2736, N2730, N11);
nor NOR4 (N2737, N2724, N667, N2665, N2027);
or OR4 (N2738, N2722, N1241, N1618, N2053);
buf BUF1 (N2739, N2732);
xor XOR2 (N2740, N2737, N1309);
buf BUF1 (N2741, N2736);
and AND4 (N2742, N2734, N1678, N39, N1048);
xor XOR2 (N2743, N2707, N1250);
or OR4 (N2744, N2729, N788, N439, N1663);
or OR3 (N2745, N2741, N1033, N1669);
nand NAND4 (N2746, N2745, N547, N906, N1279);
not NOT1 (N2747, N2703);
not NOT1 (N2748, N2738);
or OR2 (N2749, N2740, N1498);
and AND3 (N2750, N2743, N946, N141);
and AND2 (N2751, N2735, N1841);
not NOT1 (N2752, N2751);
nor NOR2 (N2753, N2742, N2032);
and AND4 (N2754, N2752, N1864, N435, N1237);
nand NAND4 (N2755, N2726, N2467, N635, N704);
or OR3 (N2756, N2755, N1664, N1166);
or OR2 (N2757, N2744, N2721);
nand NAND2 (N2758, N2739, N1836);
nand NAND4 (N2759, N2748, N1089, N1489, N289);
nor NOR2 (N2760, N2754, N401);
and AND2 (N2761, N2747, N1280);
not NOT1 (N2762, N2753);
or OR4 (N2763, N2762, N2066, N1413, N2272);
xor XOR2 (N2764, N2750, N600);
and AND3 (N2765, N2759, N1936, N477);
not NOT1 (N2766, N2757);
nor NOR3 (N2767, N2764, N2391, N2026);
and AND4 (N2768, N2756, N963, N520, N162);
or OR3 (N2769, N2768, N130, N629);
or OR2 (N2770, N2766, N366);
nor NOR3 (N2771, N2767, N451, N1853);
or OR4 (N2772, N2763, N1162, N2485, N1573);
buf BUF1 (N2773, N2758);
buf BUF1 (N2774, N2772);
xor XOR2 (N2775, N2773, N985);
buf BUF1 (N2776, N2775);
xor XOR2 (N2777, N2776, N2577);
or OR4 (N2778, N2760, N1444, N2044, N452);
nand NAND4 (N2779, N2765, N696, N492, N2681);
xor XOR2 (N2780, N2749, N1838);
buf BUF1 (N2781, N2774);
and AND2 (N2782, N2746, N1962);
and AND3 (N2783, N2778, N598, N1408);
and AND4 (N2784, N2783, N938, N87, N2723);
or OR3 (N2785, N2771, N871, N1136);
nand NAND2 (N2786, N2770, N1269);
buf BUF1 (N2787, N2777);
or OR2 (N2788, N2761, N36);
nor NOR3 (N2789, N2787, N2132, N718);
and AND2 (N2790, N2789, N1813);
nand NAND3 (N2791, N2788, N2210, N2682);
nor NOR3 (N2792, N2790, N34, N2049);
nand NAND4 (N2793, N2780, N1404, N38, N2441);
and AND4 (N2794, N2792, N837, N1101, N433);
or OR2 (N2795, N2791, N351);
buf BUF1 (N2796, N2784);
not NOT1 (N2797, N2785);
xor XOR2 (N2798, N2786, N556);
and AND4 (N2799, N2769, N992, N1930, N1023);
or OR3 (N2800, N2799, N2766, N114);
buf BUF1 (N2801, N2794);
nand NAND4 (N2802, N2793, N324, N2348, N1385);
or OR4 (N2803, N2797, N2577, N919, N68);
not NOT1 (N2804, N2798);
xor XOR2 (N2805, N2802, N2293);
nor NOR3 (N2806, N2782, N1643, N482);
and AND4 (N2807, N2805, N335, N2170, N1189);
and AND4 (N2808, N2801, N1997, N2123, N141);
not NOT1 (N2809, N2804);
xor XOR2 (N2810, N2795, N145);
nand NAND2 (N2811, N2809, N1962);
nand NAND3 (N2812, N2800, N2521, N1287);
or OR3 (N2813, N2796, N1106, N919);
nor NOR3 (N2814, N2813, N2037, N83);
not NOT1 (N2815, N2811);
nor NOR3 (N2816, N2812, N770, N1090);
not NOT1 (N2817, N2810);
not NOT1 (N2818, N2815);
buf BUF1 (N2819, N2808);
nor NOR2 (N2820, N2806, N1389);
buf BUF1 (N2821, N2817);
nand NAND2 (N2822, N2820, N2048);
nand NAND3 (N2823, N2803, N886, N2664);
xor XOR2 (N2824, N2814, N2101);
and AND2 (N2825, N2819, N1605);
xor XOR2 (N2826, N2807, N2259);
nor NOR4 (N2827, N2824, N1183, N1681, N616);
nor NOR2 (N2828, N2816, N1387);
or OR4 (N2829, N2821, N2641, N216, N1293);
nor NOR3 (N2830, N2779, N1677, N1940);
xor XOR2 (N2831, N2823, N1763);
not NOT1 (N2832, N2830);
not NOT1 (N2833, N2781);
buf BUF1 (N2834, N2826);
nand NAND3 (N2835, N2834, N2285, N1491);
not NOT1 (N2836, N2827);
and AND2 (N2837, N2832, N410);
not NOT1 (N2838, N2836);
nand NAND2 (N2839, N2831, N2405);
xor XOR2 (N2840, N2835, N1719);
not NOT1 (N2841, N2839);
buf BUF1 (N2842, N2838);
buf BUF1 (N2843, N2829);
buf BUF1 (N2844, N2837);
and AND3 (N2845, N2840, N209, N1332);
nand NAND4 (N2846, N2828, N402, N2755, N1024);
and AND3 (N2847, N2822, N130, N698);
or OR4 (N2848, N2818, N1472, N2361, N1368);
nand NAND4 (N2849, N2825, N1655, N2282, N691);
nand NAND4 (N2850, N2848, N1139, N881, N296);
and AND2 (N2851, N2847, N1994);
nor NOR3 (N2852, N2846, N1720, N434);
xor XOR2 (N2853, N2842, N369);
nor NOR3 (N2854, N2841, N61, N2364);
or OR2 (N2855, N2845, N476);
or OR2 (N2856, N2844, N1767);
xor XOR2 (N2857, N2854, N92);
not NOT1 (N2858, N2843);
or OR4 (N2859, N2856, N458, N1955, N671);
not NOT1 (N2860, N2833);
xor XOR2 (N2861, N2849, N1670);
not NOT1 (N2862, N2851);
and AND2 (N2863, N2857, N1642);
not NOT1 (N2864, N2852);
nor NOR4 (N2865, N2860, N105, N1670, N1764);
or OR3 (N2866, N2862, N2114, N1609);
and AND3 (N2867, N2866, N775, N563);
not NOT1 (N2868, N2863);
nand NAND4 (N2869, N2859, N2096, N342, N69);
buf BUF1 (N2870, N2853);
not NOT1 (N2871, N2861);
buf BUF1 (N2872, N2865);
nor NOR3 (N2873, N2858, N1387, N23);
not NOT1 (N2874, N2869);
xor XOR2 (N2875, N2872, N2337);
xor XOR2 (N2876, N2864, N1285);
buf BUF1 (N2877, N2867);
not NOT1 (N2878, N2874);
nand NAND4 (N2879, N2878, N772, N2563, N1035);
nor NOR3 (N2880, N2855, N1655, N2183);
or OR3 (N2881, N2873, N1309, N919);
not NOT1 (N2882, N2880);
and AND2 (N2883, N2875, N2684);
and AND4 (N2884, N2870, N2337, N2623, N339);
nand NAND2 (N2885, N2850, N2801);
nand NAND4 (N2886, N2871, N2236, N1158, N29);
or OR4 (N2887, N2882, N1174, N1459, N2037);
nor NOR3 (N2888, N2881, N2395, N1695);
not NOT1 (N2889, N2879);
or OR2 (N2890, N2876, N2816);
not NOT1 (N2891, N2888);
xor XOR2 (N2892, N2885, N1875);
or OR4 (N2893, N2877, N69, N606, N1980);
nor NOR3 (N2894, N2883, N1771, N1738);
buf BUF1 (N2895, N2893);
not NOT1 (N2896, N2895);
nor NOR4 (N2897, N2892, N2660, N2204, N2495);
xor XOR2 (N2898, N2894, N1949);
or OR3 (N2899, N2890, N1116, N2014);
or OR4 (N2900, N2897, N1894, N1430, N1750);
or OR2 (N2901, N2900, N2044);
buf BUF1 (N2902, N2901);
buf BUF1 (N2903, N2899);
buf BUF1 (N2904, N2891);
buf BUF1 (N2905, N2904);
buf BUF1 (N2906, N2887);
and AND2 (N2907, N2886, N1902);
nor NOR2 (N2908, N2903, N2358);
or OR3 (N2909, N2889, N996, N1307);
or OR3 (N2910, N2906, N1933, N466);
and AND2 (N2911, N2907, N955);
xor XOR2 (N2912, N2884, N270);
buf BUF1 (N2913, N2898);
or OR4 (N2914, N2912, N1988, N2014, N1774);
buf BUF1 (N2915, N2902);
and AND3 (N2916, N2905, N1177, N859);
buf BUF1 (N2917, N2911);
or OR2 (N2918, N2896, N729);
or OR4 (N2919, N2913, N2744, N917, N2693);
or OR3 (N2920, N2918, N1851, N1751);
or OR2 (N2921, N2909, N323);
and AND2 (N2922, N2919, N848);
nand NAND2 (N2923, N2914, N1116);
xor XOR2 (N2924, N2921, N782);
not NOT1 (N2925, N2923);
and AND2 (N2926, N2920, N2230);
nand NAND2 (N2927, N2917, N689);
nor NOR4 (N2928, N2924, N1908, N2020, N2214);
xor XOR2 (N2929, N2868, N2568);
nor NOR2 (N2930, N2929, N2049);
or OR4 (N2931, N2925, N1377, N892, N2342);
and AND4 (N2932, N2908, N831, N1812, N1324);
and AND2 (N2933, N2932, N2843);
not NOT1 (N2934, N2927);
xor XOR2 (N2935, N2928, N21);
nor NOR4 (N2936, N2933, N2616, N2797, N1452);
nand NAND3 (N2937, N2916, N52, N2202);
xor XOR2 (N2938, N2915, N2063);
xor XOR2 (N2939, N2931, N1661);
not NOT1 (N2940, N2922);
nand NAND2 (N2941, N2935, N1592);
buf BUF1 (N2942, N2937);
nor NOR3 (N2943, N2939, N2249, N301);
not NOT1 (N2944, N2941);
and AND3 (N2945, N2926, N1693, N154);
nand NAND2 (N2946, N2930, N2259);
nor NOR4 (N2947, N2938, N2344, N2807, N2429);
buf BUF1 (N2948, N2910);
or OR2 (N2949, N2947, N180);
and AND2 (N2950, N2944, N2884);
nand NAND2 (N2951, N2934, N1984);
not NOT1 (N2952, N2940);
nand NAND2 (N2953, N2948, N1486);
or OR4 (N2954, N2946, N2628, N1310, N139);
nand NAND4 (N2955, N2936, N918, N1359, N1301);
nand NAND4 (N2956, N2950, N794, N1394, N278);
buf BUF1 (N2957, N2955);
buf BUF1 (N2958, N2954);
xor XOR2 (N2959, N2945, N382);
or OR4 (N2960, N2953, N1090, N957, N158);
not NOT1 (N2961, N2956);
buf BUF1 (N2962, N2961);
nand NAND2 (N2963, N2959, N1543);
nor NOR2 (N2964, N2958, N658);
not NOT1 (N2965, N2952);
nor NOR2 (N2966, N2942, N1762);
or OR3 (N2967, N2962, N1630, N1863);
nand NAND4 (N2968, N2963, N1330, N1414, N2131);
not NOT1 (N2969, N2968);
nor NOR3 (N2970, N2969, N2858, N1548);
or OR4 (N2971, N2965, N2763, N719, N1487);
or OR2 (N2972, N2964, N635);
xor XOR2 (N2973, N2970, N1271);
xor XOR2 (N2974, N2973, N2927);
not NOT1 (N2975, N2967);
and AND4 (N2976, N2943, N1366, N2286, N1353);
nand NAND3 (N2977, N2960, N829, N324);
nand NAND3 (N2978, N2957, N1832, N1327);
buf BUF1 (N2979, N2977);
and AND4 (N2980, N2975, N394, N565, N1953);
and AND4 (N2981, N2980, N327, N2267, N1597);
or OR4 (N2982, N2981, N2799, N2904, N1145);
xor XOR2 (N2983, N2976, N2722);
nor NOR4 (N2984, N2979, N1054, N2916, N1193);
or OR2 (N2985, N2972, N365);
or OR2 (N2986, N2966, N512);
and AND4 (N2987, N2974, N197, N155, N60);
nor NOR4 (N2988, N2983, N788, N729, N1299);
nand NAND4 (N2989, N2986, N514, N2037, N1645);
buf BUF1 (N2990, N2949);
nor NOR3 (N2991, N2990, N2389, N1007);
or OR2 (N2992, N2971, N187);
nor NOR3 (N2993, N2987, N2619, N146);
buf BUF1 (N2994, N2978);
nand NAND2 (N2995, N2951, N408);
or OR4 (N2996, N2984, N2063, N972, N881);
nand NAND3 (N2997, N2993, N23, N1107);
xor XOR2 (N2998, N2985, N2199);
buf BUF1 (N2999, N2998);
xor XOR2 (N3000, N2988, N1789);
not NOT1 (N3001, N2982);
and AND4 (N3002, N2991, N125, N364, N935);
xor XOR2 (N3003, N2994, N688);
xor XOR2 (N3004, N2989, N967);
or OR4 (N3005, N2996, N2529, N2354, N820);
nand NAND4 (N3006, N2992, N2516, N2746, N585);
xor XOR2 (N3007, N3006, N72);
not NOT1 (N3008, N2997);
buf BUF1 (N3009, N3000);
not NOT1 (N3010, N2995);
and AND4 (N3011, N3007, N1412, N99, N157);
xor XOR2 (N3012, N3010, N283);
xor XOR2 (N3013, N2999, N2135);
xor XOR2 (N3014, N3011, N2327);
and AND2 (N3015, N3005, N688);
or OR3 (N3016, N3014, N740, N2967);
and AND3 (N3017, N3001, N1868, N1709);
or OR4 (N3018, N3015, N2756, N567, N1680);
or OR2 (N3019, N3002, N567);
xor XOR2 (N3020, N3018, N2486);
buf BUF1 (N3021, N3003);
and AND4 (N3022, N3008, N1726, N2755, N1356);
not NOT1 (N3023, N3019);
not NOT1 (N3024, N3013);
buf BUF1 (N3025, N3004);
buf BUF1 (N3026, N3023);
or OR2 (N3027, N3021, N1417);
buf BUF1 (N3028, N3026);
and AND4 (N3029, N3016, N1973, N2586, N2256);
xor XOR2 (N3030, N3028, N2739);
not NOT1 (N3031, N3012);
nand NAND3 (N3032, N3029, N891, N1243);
buf BUF1 (N3033, N3017);
not NOT1 (N3034, N3020);
nand NAND4 (N3035, N3033, N1002, N168, N1578);
and AND3 (N3036, N3032, N773, N2210);
xor XOR2 (N3037, N3035, N1688);
or OR2 (N3038, N3031, N765);
and AND2 (N3039, N3037, N1232);
not NOT1 (N3040, N3039);
or OR4 (N3041, N3038, N111, N2804, N528);
nand NAND2 (N3042, N3040, N1312);
nand NAND4 (N3043, N3022, N2962, N2349, N2460);
nand NAND2 (N3044, N3042, N393);
xor XOR2 (N3045, N3044, N198);
and AND3 (N3046, N3043, N2922, N859);
nor NOR3 (N3047, N3034, N32, N1016);
nand NAND4 (N3048, N3047, N45, N1453, N1944);
xor XOR2 (N3049, N3048, N1037);
buf BUF1 (N3050, N3024);
and AND2 (N3051, N3046, N629);
nand NAND4 (N3052, N3041, N182, N2889, N396);
or OR3 (N3053, N3050, N2838, N746);
nand NAND2 (N3054, N3049, N1336);
and AND3 (N3055, N3054, N816, N1086);
nand NAND4 (N3056, N3009, N162, N247, N1503);
and AND4 (N3057, N3055, N167, N140, N2310);
and AND3 (N3058, N3057, N300, N348);
xor XOR2 (N3059, N3045, N2322);
xor XOR2 (N3060, N3036, N3);
nor NOR3 (N3061, N3060, N2628, N842);
xor XOR2 (N3062, N3051, N1284);
not NOT1 (N3063, N3062);
or OR3 (N3064, N3053, N873, N2387);
and AND4 (N3065, N3061, N1427, N3, N2542);
not NOT1 (N3066, N3065);
xor XOR2 (N3067, N3063, N173);
xor XOR2 (N3068, N3056, N1936);
nor NOR3 (N3069, N3064, N363, N3006);
or OR3 (N3070, N3069, N807, N2815);
not NOT1 (N3071, N3027);
nor NOR4 (N3072, N3059, N1549, N2312, N1344);
nor NOR4 (N3073, N3066, N935, N2931, N1243);
nor NOR3 (N3074, N3068, N1997, N2359);
xor XOR2 (N3075, N3030, N3055);
not NOT1 (N3076, N3074);
xor XOR2 (N3077, N3072, N931);
not NOT1 (N3078, N3070);
nand NAND2 (N3079, N3077, N1932);
nand NAND3 (N3080, N3078, N2791, N1844);
nor NOR2 (N3081, N3058, N243);
nand NAND2 (N3082, N3076, N2195);
xor XOR2 (N3083, N3052, N935);
not NOT1 (N3084, N3079);
nor NOR4 (N3085, N3073, N2631, N1290, N1477);
and AND3 (N3086, N3084, N431, N1919);
or OR3 (N3087, N3083, N2062, N1608);
not NOT1 (N3088, N3087);
buf BUF1 (N3089, N3088);
nand NAND3 (N3090, N3025, N1448, N403);
nor NOR3 (N3091, N3067, N1891, N694);
and AND4 (N3092, N3089, N915, N2648, N891);
nand NAND4 (N3093, N3090, N1037, N299, N1578);
nor NOR4 (N3094, N3082, N2006, N1503, N525);
buf BUF1 (N3095, N3086);
buf BUF1 (N3096, N3093);
not NOT1 (N3097, N3094);
buf BUF1 (N3098, N3080);
nor NOR2 (N3099, N3098, N192);
or OR3 (N3100, N3097, N2075, N2165);
xor XOR2 (N3101, N3075, N1221);
and AND4 (N3102, N3092, N2768, N1890, N514);
buf BUF1 (N3103, N3099);
nor NOR4 (N3104, N3095, N1868, N1955, N621);
buf BUF1 (N3105, N3102);
not NOT1 (N3106, N3081);
nand NAND4 (N3107, N3100, N221, N312, N817);
nand NAND4 (N3108, N3101, N87, N828, N804);
and AND3 (N3109, N3096, N522, N974);
nor NOR3 (N3110, N3085, N2405, N2195);
not NOT1 (N3111, N3107);
nor NOR2 (N3112, N3110, N237);
xor XOR2 (N3113, N3105, N2302);
buf BUF1 (N3114, N3071);
buf BUF1 (N3115, N3111);
buf BUF1 (N3116, N3113);
xor XOR2 (N3117, N3112, N1326);
nand NAND3 (N3118, N3116, N2763, N2199);
buf BUF1 (N3119, N3106);
nand NAND2 (N3120, N3108, N3096);
not NOT1 (N3121, N3114);
nor NOR3 (N3122, N3120, N1807, N1333);
and AND4 (N3123, N3103, N430, N89, N143);
xor XOR2 (N3124, N3118, N2906);
nand NAND2 (N3125, N3109, N1611);
and AND4 (N3126, N3091, N194, N1368, N1572);
nand NAND4 (N3127, N3123, N1757, N1128, N2048);
or OR3 (N3128, N3122, N1162, N1634);
buf BUF1 (N3129, N3125);
or OR2 (N3130, N3121, N1612);
not NOT1 (N3131, N3130);
xor XOR2 (N3132, N3104, N1493);
xor XOR2 (N3133, N3119, N3081);
not NOT1 (N3134, N3117);
xor XOR2 (N3135, N3133, N675);
not NOT1 (N3136, N3127);
xor XOR2 (N3137, N3131, N375);
xor XOR2 (N3138, N3136, N364);
buf BUF1 (N3139, N3134);
and AND2 (N3140, N3115, N1897);
xor XOR2 (N3141, N3124, N2463);
or OR2 (N3142, N3132, N2050);
or OR2 (N3143, N3141, N2135);
not NOT1 (N3144, N3139);
and AND4 (N3145, N3138, N441, N943, N2698);
nand NAND3 (N3146, N3145, N2859, N2942);
nor NOR3 (N3147, N3140, N1259, N1239);
buf BUF1 (N3148, N3142);
buf BUF1 (N3149, N3137);
and AND4 (N3150, N3148, N1819, N2795, N2446);
and AND3 (N3151, N3150, N711, N1554);
nor NOR2 (N3152, N3149, N1207);
xor XOR2 (N3153, N3146, N2745);
or OR2 (N3154, N3126, N1798);
xor XOR2 (N3155, N3147, N157);
and AND4 (N3156, N3128, N1335, N1260, N2177);
or OR4 (N3157, N3135, N2751, N95, N420);
or OR2 (N3158, N3153, N746);
xor XOR2 (N3159, N3156, N2824);
buf BUF1 (N3160, N3152);
or OR3 (N3161, N3157, N925, N2623);
and AND4 (N3162, N3129, N648, N2244, N453);
not NOT1 (N3163, N3143);
nand NAND4 (N3164, N3151, N2889, N2655, N2278);
not NOT1 (N3165, N3162);
and AND4 (N3166, N3159, N3154, N1883, N2568);
or OR4 (N3167, N2376, N1313, N2971, N166);
nor NOR3 (N3168, N3144, N174, N1893);
nand NAND3 (N3169, N3165, N184, N657);
not NOT1 (N3170, N3166);
nand NAND4 (N3171, N3160, N1760, N1356, N943);
or OR4 (N3172, N3164, N695, N177, N2222);
not NOT1 (N3173, N3167);
nor NOR2 (N3174, N3170, N2375);
and AND3 (N3175, N3173, N1459, N1888);
buf BUF1 (N3176, N3163);
or OR3 (N3177, N3175, N439, N2495);
not NOT1 (N3178, N3172);
xor XOR2 (N3179, N3168, N845);
xor XOR2 (N3180, N3158, N2471);
or OR3 (N3181, N3179, N2598, N3169);
xor XOR2 (N3182, N2648, N754);
xor XOR2 (N3183, N3171, N3131);
or OR3 (N3184, N3182, N902, N1026);
nand NAND3 (N3185, N3177, N19, N2802);
xor XOR2 (N3186, N3181, N3132);
nand NAND4 (N3187, N3161, N729, N2258, N1610);
nor NOR4 (N3188, N3155, N2260, N602, N2925);
nor NOR4 (N3189, N3178, N199, N1000, N983);
or OR3 (N3190, N3184, N910, N3149);
nor NOR2 (N3191, N3186, N2679);
nor NOR2 (N3192, N3176, N1893);
xor XOR2 (N3193, N3187, N1648);
and AND4 (N3194, N3190, N2014, N1836, N1135);
buf BUF1 (N3195, N3185);
xor XOR2 (N3196, N3192, N1777);
buf BUF1 (N3197, N3193);
not NOT1 (N3198, N3188);
not NOT1 (N3199, N3180);
buf BUF1 (N3200, N3189);
xor XOR2 (N3201, N3194, N3126);
or OR2 (N3202, N3174, N2151);
not NOT1 (N3203, N3183);
xor XOR2 (N3204, N3191, N2959);
not NOT1 (N3205, N3196);
not NOT1 (N3206, N3195);
nor NOR2 (N3207, N3200, N1096);
and AND4 (N3208, N3197, N1920, N324, N2613);
xor XOR2 (N3209, N3207, N30);
or OR3 (N3210, N3204, N487, N3179);
nor NOR4 (N3211, N3208, N2979, N2219, N919);
and AND2 (N3212, N3211, N842);
nand NAND4 (N3213, N3199, N486, N276, N2763);
nand NAND3 (N3214, N3209, N2488, N230);
and AND4 (N3215, N3201, N775, N2458, N3062);
not NOT1 (N3216, N3206);
nor NOR3 (N3217, N3205, N459, N2767);
buf BUF1 (N3218, N3212);
nor NOR3 (N3219, N3215, N1377, N2006);
buf BUF1 (N3220, N3218);
and AND4 (N3221, N3214, N641, N485, N2059);
or OR4 (N3222, N3217, N1623, N2150, N2545);
nor NOR2 (N3223, N3202, N2393);
or OR2 (N3224, N3220, N2197);
buf BUF1 (N3225, N3216);
or OR3 (N3226, N3219, N254, N2699);
nand NAND4 (N3227, N3198, N2494, N759, N292);
not NOT1 (N3228, N3213);
and AND3 (N3229, N3221, N2553, N2687);
nand NAND2 (N3230, N3224, N610);
buf BUF1 (N3231, N3210);
and AND4 (N3232, N3226, N713, N1916, N354);
or OR3 (N3233, N3229, N236, N1354);
and AND4 (N3234, N3225, N674, N1678, N2474);
xor XOR2 (N3235, N3228, N841);
or OR4 (N3236, N3235, N2445, N1670, N2186);
not NOT1 (N3237, N3203);
or OR3 (N3238, N3223, N931, N1333);
nor NOR3 (N3239, N3227, N1700, N1820);
xor XOR2 (N3240, N3231, N2808);
or OR3 (N3241, N3233, N2030, N2248);
not NOT1 (N3242, N3240);
nand NAND4 (N3243, N3222, N1600, N2101, N87);
or OR2 (N3244, N3243, N2642);
xor XOR2 (N3245, N3244, N1565);
xor XOR2 (N3246, N3245, N2942);
xor XOR2 (N3247, N3237, N2221);
buf BUF1 (N3248, N3232);
xor XOR2 (N3249, N3246, N653);
nor NOR4 (N3250, N3249, N2745, N3058, N603);
nand NAND3 (N3251, N3234, N1370, N373);
nand NAND2 (N3252, N3238, N2403);
nand NAND3 (N3253, N3252, N1014, N1746);
xor XOR2 (N3254, N3241, N3138);
or OR3 (N3255, N3251, N1760, N1787);
or OR4 (N3256, N3253, N1526, N199, N1158);
nor NOR2 (N3257, N3256, N295);
nor NOR3 (N3258, N3254, N3099, N2601);
xor XOR2 (N3259, N3248, N2882);
buf BUF1 (N3260, N3247);
and AND4 (N3261, N3236, N752, N1073, N1322);
buf BUF1 (N3262, N3255);
or OR4 (N3263, N3261, N135, N2661, N3115);
and AND4 (N3264, N3260, N1949, N1386, N233);
xor XOR2 (N3265, N3259, N1244);
or OR3 (N3266, N3258, N2265, N295);
nand NAND4 (N3267, N3257, N2576, N2170, N101);
buf BUF1 (N3268, N3265);
or OR3 (N3269, N3230, N2303, N2035);
xor XOR2 (N3270, N3263, N2595);
and AND2 (N3271, N3269, N1965);
not NOT1 (N3272, N3271);
not NOT1 (N3273, N3250);
not NOT1 (N3274, N3239);
buf BUF1 (N3275, N3274);
buf BUF1 (N3276, N3270);
or OR3 (N3277, N3275, N1633, N936);
buf BUF1 (N3278, N3262);
or OR3 (N3279, N3266, N490, N3083);
nand NAND4 (N3280, N3273, N1343, N184, N651);
xor XOR2 (N3281, N3277, N2237);
not NOT1 (N3282, N3267);
nand NAND4 (N3283, N3281, N339, N2466, N993);
nand NAND4 (N3284, N3282, N2816, N3112, N968);
not NOT1 (N3285, N3268);
nor NOR2 (N3286, N3279, N296);
buf BUF1 (N3287, N3284);
xor XOR2 (N3288, N3264, N2388);
or OR3 (N3289, N3272, N3064, N750);
xor XOR2 (N3290, N3278, N227);
not NOT1 (N3291, N3286);
not NOT1 (N3292, N3285);
nor NOR4 (N3293, N3292, N1892, N1342, N712);
nand NAND2 (N3294, N3283, N1723);
nand NAND4 (N3295, N3291, N1532, N77, N2848);
buf BUF1 (N3296, N3289);
nor NOR2 (N3297, N3288, N329);
and AND3 (N3298, N3297, N1945, N123);
buf BUF1 (N3299, N3294);
or OR3 (N3300, N3298, N2853, N209);
and AND2 (N3301, N3295, N322);
and AND4 (N3302, N3287, N1426, N2352, N1488);
not NOT1 (N3303, N3301);
nand NAND2 (N3304, N3300, N2340);
xor XOR2 (N3305, N3290, N3206);
nand NAND4 (N3306, N3304, N1582, N2954, N3102);
nand NAND2 (N3307, N3293, N982);
xor XOR2 (N3308, N3302, N1201);
xor XOR2 (N3309, N3307, N1339);
and AND4 (N3310, N3299, N2562, N360, N2150);
not NOT1 (N3311, N3306);
or OR3 (N3312, N3242, N2322, N676);
or OR2 (N3313, N3311, N3207);
nand NAND3 (N3314, N3296, N1769, N1549);
nor NOR4 (N3315, N3305, N458, N3156, N2603);
nand NAND4 (N3316, N3313, N127, N482, N346);
and AND3 (N3317, N3316, N1125, N2432);
not NOT1 (N3318, N3303);
buf BUF1 (N3319, N3309);
and AND4 (N3320, N3312, N2213, N1747, N841);
nand NAND4 (N3321, N3318, N1687, N2123, N2034);
buf BUF1 (N3322, N3321);
or OR3 (N3323, N3308, N3267, N445);
not NOT1 (N3324, N3310);
not NOT1 (N3325, N3280);
nor NOR4 (N3326, N3319, N2951, N3177, N1871);
buf BUF1 (N3327, N3322);
nor NOR2 (N3328, N3314, N553);
xor XOR2 (N3329, N3328, N564);
buf BUF1 (N3330, N3323);
or OR2 (N3331, N3325, N2775);
and AND4 (N3332, N3315, N1900, N1701, N1932);
and AND2 (N3333, N3326, N340);
not NOT1 (N3334, N3327);
xor XOR2 (N3335, N3330, N1623);
not NOT1 (N3336, N3334);
not NOT1 (N3337, N3331);
and AND2 (N3338, N3317, N1313);
and AND3 (N3339, N3276, N730, N785);
not NOT1 (N3340, N3329);
or OR2 (N3341, N3335, N2534);
not NOT1 (N3342, N3320);
and AND3 (N3343, N3341, N1869, N1043);
nand NAND4 (N3344, N3340, N2097, N1063, N2264);
or OR2 (N3345, N3339, N3168);
and AND4 (N3346, N3338, N2460, N1318, N2396);
not NOT1 (N3347, N3345);
not NOT1 (N3348, N3346);
buf BUF1 (N3349, N3324);
buf BUF1 (N3350, N3336);
not NOT1 (N3351, N3349);
buf BUF1 (N3352, N3351);
xor XOR2 (N3353, N3352, N1994);
not NOT1 (N3354, N3350);
not NOT1 (N3355, N3342);
nand NAND4 (N3356, N3348, N3135, N1406, N2008);
buf BUF1 (N3357, N3333);
not NOT1 (N3358, N3347);
not NOT1 (N3359, N3353);
xor XOR2 (N3360, N3359, N3181);
or OR2 (N3361, N3358, N2415);
and AND2 (N3362, N3354, N2218);
and AND4 (N3363, N3356, N1600, N1581, N67);
or OR2 (N3364, N3357, N3251);
and AND3 (N3365, N3337, N3247, N2586);
buf BUF1 (N3366, N3365);
nor NOR3 (N3367, N3344, N1750, N2640);
buf BUF1 (N3368, N3363);
nor NOR4 (N3369, N3362, N475, N2444, N2328);
buf BUF1 (N3370, N3369);
nor NOR4 (N3371, N3343, N28, N1062, N2474);
not NOT1 (N3372, N3355);
nor NOR2 (N3373, N3360, N3296);
xor XOR2 (N3374, N3372, N172);
xor XOR2 (N3375, N3368, N2440);
buf BUF1 (N3376, N3366);
xor XOR2 (N3377, N3371, N1005);
nor NOR2 (N3378, N3367, N2688);
buf BUF1 (N3379, N3332);
nand NAND4 (N3380, N3370, N843, N1024, N478);
xor XOR2 (N3381, N3380, N1807);
and AND4 (N3382, N3378, N1515, N1631, N1082);
nor NOR4 (N3383, N3381, N842, N961, N568);
nor NOR4 (N3384, N3364, N159, N655, N1247);
buf BUF1 (N3385, N3384);
nand NAND3 (N3386, N3385, N2221, N1421);
and AND2 (N3387, N3386, N3191);
buf BUF1 (N3388, N3377);
xor XOR2 (N3389, N3361, N783);
xor XOR2 (N3390, N3388, N6);
and AND4 (N3391, N3375, N3333, N289, N2374);
buf BUF1 (N3392, N3376);
and AND4 (N3393, N3374, N553, N2800, N2426);
xor XOR2 (N3394, N3383, N2295);
nor NOR2 (N3395, N3391, N849);
xor XOR2 (N3396, N3392, N2739);
or OR3 (N3397, N3382, N1960, N1379);
or OR3 (N3398, N3379, N1854, N472);
and AND3 (N3399, N3390, N2211, N1470);
or OR4 (N3400, N3394, N1323, N897, N2370);
nor NOR2 (N3401, N3397, N127);
and AND3 (N3402, N3387, N2350, N532);
not NOT1 (N3403, N3400);
not NOT1 (N3404, N3402);
nand NAND2 (N3405, N3396, N3137);
nor NOR2 (N3406, N3389, N262);
and AND3 (N3407, N3406, N1988, N49);
nor NOR3 (N3408, N3405, N2429, N2957);
nor NOR3 (N3409, N3398, N172, N2030);
not NOT1 (N3410, N3395);
or OR3 (N3411, N3373, N215, N3234);
and AND2 (N3412, N3393, N1560);
or OR2 (N3413, N3403, N2870);
xor XOR2 (N3414, N3409, N3313);
and AND4 (N3415, N3414, N2165, N486, N700);
nand NAND3 (N3416, N3415, N2102, N1088);
nand NAND2 (N3417, N3412, N2371);
and AND4 (N3418, N3410, N808, N584, N2210);
or OR3 (N3419, N3401, N2136, N1182);
nand NAND2 (N3420, N3417, N175);
not NOT1 (N3421, N3418);
or OR3 (N3422, N3407, N423, N1785);
nand NAND2 (N3423, N3421, N1920);
xor XOR2 (N3424, N3416, N814);
or OR2 (N3425, N3399, N1368);
or OR4 (N3426, N3424, N2542, N1048, N2167);
nand NAND2 (N3427, N3425, N2221);
not NOT1 (N3428, N3426);
xor XOR2 (N3429, N3404, N57);
nand NAND4 (N3430, N3429, N1803, N2, N2217);
buf BUF1 (N3431, N3413);
not NOT1 (N3432, N3408);
nor NOR4 (N3433, N3428, N1397, N1228, N3178);
nand NAND3 (N3434, N3433, N2997, N2743);
and AND3 (N3435, N3432, N151, N2932);
xor XOR2 (N3436, N3427, N2205);
xor XOR2 (N3437, N3431, N2360);
nor NOR4 (N3438, N3437, N1854, N1291, N2812);
nand NAND2 (N3439, N3438, N2163);
or OR2 (N3440, N3423, N3099);
not NOT1 (N3441, N3440);
xor XOR2 (N3442, N3422, N2476);
nand NAND2 (N3443, N3435, N2587);
and AND2 (N3444, N3442, N1478);
not NOT1 (N3445, N3411);
buf BUF1 (N3446, N3444);
and AND4 (N3447, N3439, N1380, N1116, N695);
or OR2 (N3448, N3430, N2124);
or OR3 (N3449, N3434, N1944, N96);
nand NAND4 (N3450, N3445, N1705, N3009, N3282);
buf BUF1 (N3451, N3448);
and AND2 (N3452, N3450, N1775);
nor NOR3 (N3453, N3446, N3003, N1912);
nand NAND4 (N3454, N3436, N839, N2972, N3331);
buf BUF1 (N3455, N3447);
and AND4 (N3456, N3420, N922, N2591, N923);
and AND3 (N3457, N3443, N2350, N594);
xor XOR2 (N3458, N3452, N2006);
nor NOR4 (N3459, N3441, N3108, N2119, N206);
not NOT1 (N3460, N3457);
nor NOR3 (N3461, N3453, N2082, N73);
xor XOR2 (N3462, N3455, N2409);
xor XOR2 (N3463, N3419, N1458);
nand NAND3 (N3464, N3458, N2108, N2515);
nand NAND3 (N3465, N3451, N3456, N3008);
not NOT1 (N3466, N387);
xor XOR2 (N3467, N3459, N755);
and AND2 (N3468, N3460, N548);
xor XOR2 (N3469, N3449, N3461);
nand NAND4 (N3470, N3328, N2907, N660, N981);
nor NOR3 (N3471, N3464, N2157, N1201);
or OR3 (N3472, N3467, N1101, N719);
nand NAND3 (N3473, N3470, N2635, N2096);
xor XOR2 (N3474, N3454, N682);
xor XOR2 (N3475, N3465, N1026);
nor NOR2 (N3476, N3474, N361);
not NOT1 (N3477, N3462);
or OR2 (N3478, N3475, N825);
nand NAND3 (N3479, N3466, N1990, N1900);
buf BUF1 (N3480, N3479);
buf BUF1 (N3481, N3476);
nand NAND3 (N3482, N3463, N2309, N477);
and AND4 (N3483, N3471, N2851, N263, N69);
and AND2 (N3484, N3480, N742);
buf BUF1 (N3485, N3483);
or OR4 (N3486, N3469, N958, N2042, N1919);
not NOT1 (N3487, N3482);
not NOT1 (N3488, N3477);
xor XOR2 (N3489, N3472, N2781);
or OR4 (N3490, N3468, N192, N2511, N3457);
or OR3 (N3491, N3486, N1350, N1867);
nand NAND4 (N3492, N3489, N2410, N3332, N3040);
xor XOR2 (N3493, N3490, N2549);
buf BUF1 (N3494, N3492);
nand NAND4 (N3495, N3478, N3373, N811, N369);
xor XOR2 (N3496, N3491, N2765);
and AND2 (N3497, N3481, N2862);
not NOT1 (N3498, N3494);
not NOT1 (N3499, N3484);
nor NOR4 (N3500, N3496, N2283, N1940, N2365);
nand NAND2 (N3501, N3487, N1880);
and AND3 (N3502, N3493, N1328, N51);
nor NOR4 (N3503, N3497, N1336, N2455, N1471);
buf BUF1 (N3504, N3501);
xor XOR2 (N3505, N3500, N499);
nor NOR2 (N3506, N3498, N3168);
or OR2 (N3507, N3473, N2073);
nand NAND3 (N3508, N3485, N578, N59);
nor NOR2 (N3509, N3495, N1312);
buf BUF1 (N3510, N3509);
or OR2 (N3511, N3508, N2936);
nor NOR2 (N3512, N3507, N958);
xor XOR2 (N3513, N3502, N47);
or OR2 (N3514, N3511, N2157);
nand NAND4 (N3515, N3499, N2493, N805, N2711);
or OR2 (N3516, N3505, N2953);
xor XOR2 (N3517, N3512, N2419);
buf BUF1 (N3518, N3514);
buf BUF1 (N3519, N3518);
xor XOR2 (N3520, N3488, N1964);
not NOT1 (N3521, N3513);
xor XOR2 (N3522, N3521, N3278);
nor NOR3 (N3523, N3504, N2529, N1007);
and AND3 (N3524, N3523, N2987, N1262);
not NOT1 (N3525, N3519);
buf BUF1 (N3526, N3510);
and AND4 (N3527, N3503, N1760, N3411, N2166);
or OR2 (N3528, N3506, N1802);
nor NOR2 (N3529, N3525, N2237);
and AND4 (N3530, N3520, N1407, N375, N2113);
not NOT1 (N3531, N3516);
buf BUF1 (N3532, N3529);
and AND3 (N3533, N3531, N666, N1855);
xor XOR2 (N3534, N3517, N1165);
nand NAND2 (N3535, N3522, N3094);
nor NOR4 (N3536, N3524, N2614, N1464, N1758);
nor NOR4 (N3537, N3515, N131, N3126, N1364);
not NOT1 (N3538, N3532);
nor NOR2 (N3539, N3538, N1940);
nor NOR2 (N3540, N3534, N313);
and AND2 (N3541, N3533, N3180);
or OR2 (N3542, N3540, N172);
buf BUF1 (N3543, N3539);
or OR4 (N3544, N3528, N3336, N2724, N1027);
nor NOR3 (N3545, N3542, N3416, N284);
nand NAND2 (N3546, N3541, N140);
nor NOR3 (N3547, N3543, N498, N361);
and AND4 (N3548, N3535, N756, N1816, N237);
not NOT1 (N3549, N3526);
nand NAND3 (N3550, N3530, N818, N475);
buf BUF1 (N3551, N3545);
buf BUF1 (N3552, N3547);
and AND2 (N3553, N3552, N2999);
or OR4 (N3554, N3551, N1945, N1303, N1832);
or OR2 (N3555, N3550, N512);
nor NOR4 (N3556, N3548, N3466, N837, N3416);
nor NOR3 (N3557, N3536, N2331, N1158);
nor NOR2 (N3558, N3553, N1531);
not NOT1 (N3559, N3554);
nor NOR4 (N3560, N3556, N1210, N2853, N1182);
xor XOR2 (N3561, N3537, N1244);
nand NAND4 (N3562, N3549, N2851, N2840, N1194);
or OR2 (N3563, N3546, N106);
buf BUF1 (N3564, N3563);
and AND3 (N3565, N3557, N666, N2155);
not NOT1 (N3566, N3561);
and AND4 (N3567, N3564, N2128, N2990, N1479);
nand NAND2 (N3568, N3544, N2834);
or OR2 (N3569, N3567, N1704);
not NOT1 (N3570, N3555);
nand NAND3 (N3571, N3570, N2040, N3299);
not NOT1 (N3572, N3527);
and AND2 (N3573, N3568, N3560);
buf BUF1 (N3574, N1282);
not NOT1 (N3575, N3573);
or OR4 (N3576, N3565, N750, N208, N1325);
xor XOR2 (N3577, N3575, N2601);
buf BUF1 (N3578, N3577);
or OR3 (N3579, N3572, N1019, N3160);
or OR3 (N3580, N3566, N2921, N332);
and AND4 (N3581, N3571, N3489, N1631, N694);
buf BUF1 (N3582, N3562);
or OR4 (N3583, N3558, N938, N2078, N2672);
or OR2 (N3584, N3559, N3474);
buf BUF1 (N3585, N3582);
nor NOR2 (N3586, N3579, N679);
or OR4 (N3587, N3578, N771, N226, N3304);
not NOT1 (N3588, N3587);
xor XOR2 (N3589, N3581, N2914);
and AND3 (N3590, N3589, N288, N302);
nand NAND3 (N3591, N3569, N1864, N1716);
and AND2 (N3592, N3576, N1093);
and AND2 (N3593, N3592, N3323);
xor XOR2 (N3594, N3585, N1056);
or OR2 (N3595, N3590, N1833);
buf BUF1 (N3596, N3594);
not NOT1 (N3597, N3588);
or OR2 (N3598, N3574, N3579);
xor XOR2 (N3599, N3596, N2442);
or OR3 (N3600, N3583, N198, N580);
xor XOR2 (N3601, N3600, N2756);
not NOT1 (N3602, N3591);
nor NOR2 (N3603, N3601, N2605);
or OR2 (N3604, N3595, N1811);
not NOT1 (N3605, N3598);
not NOT1 (N3606, N3603);
buf BUF1 (N3607, N3597);
buf BUF1 (N3608, N3580);
buf BUF1 (N3609, N3602);
nand NAND2 (N3610, N3599, N2087);
xor XOR2 (N3611, N3610, N683);
nor NOR2 (N3612, N3593, N3426);
nand NAND2 (N3613, N3611, N2657);
not NOT1 (N3614, N3606);
buf BUF1 (N3615, N3584);
nor NOR3 (N3616, N3609, N1944, N1035);
and AND3 (N3617, N3586, N2368, N3023);
not NOT1 (N3618, N3608);
nand NAND3 (N3619, N3615, N1514, N3346);
xor XOR2 (N3620, N3604, N3605);
buf BUF1 (N3621, N3152);
not NOT1 (N3622, N3614);
nand NAND3 (N3623, N3619, N1014, N3401);
buf BUF1 (N3624, N3612);
nor NOR2 (N3625, N3624, N10);
nor NOR2 (N3626, N3621, N1567);
not NOT1 (N3627, N3626);
xor XOR2 (N3628, N3622, N3072);
and AND3 (N3629, N3627, N1852, N652);
nand NAND2 (N3630, N3618, N126);
xor XOR2 (N3631, N3620, N3172);
and AND3 (N3632, N3630, N3347, N524);
xor XOR2 (N3633, N3625, N1838);
nand NAND4 (N3634, N3631, N3380, N1933, N2652);
and AND2 (N3635, N3617, N2170);
or OR3 (N3636, N3616, N2492, N2903);
nor NOR4 (N3637, N3636, N999, N2134, N492);
xor XOR2 (N3638, N3629, N1735);
or OR3 (N3639, N3633, N2488, N3561);
xor XOR2 (N3640, N3623, N1864);
nand NAND4 (N3641, N3607, N2728, N359, N2734);
buf BUF1 (N3642, N3632);
or OR3 (N3643, N3635, N3139, N1257);
buf BUF1 (N3644, N3639);
and AND2 (N3645, N3640, N347);
or OR2 (N3646, N3628, N2777);
or OR3 (N3647, N3638, N1360, N909);
nand NAND2 (N3648, N3647, N3012);
nand NAND2 (N3649, N3644, N1589);
not NOT1 (N3650, N3613);
and AND2 (N3651, N3646, N911);
or OR4 (N3652, N3637, N3110, N850, N2154);
buf BUF1 (N3653, N3643);
buf BUF1 (N3654, N3649);
xor XOR2 (N3655, N3653, N2355);
xor XOR2 (N3656, N3651, N430);
nand NAND3 (N3657, N3641, N3060, N1514);
not NOT1 (N3658, N3650);
buf BUF1 (N3659, N3634);
and AND4 (N3660, N3648, N645, N3176, N2154);
nor NOR3 (N3661, N3658, N2104, N3312);
not NOT1 (N3662, N3656);
and AND4 (N3663, N3662, N2850, N341, N11);
or OR3 (N3664, N3655, N2984, N770);
and AND4 (N3665, N3657, N2941, N3631, N2943);
nor NOR3 (N3666, N3654, N2292, N3604);
and AND2 (N3667, N3665, N1371);
and AND4 (N3668, N3667, N1505, N2076, N3181);
xor XOR2 (N3669, N3668, N1098);
nand NAND3 (N3670, N3669, N2967, N3251);
nand NAND2 (N3671, N3645, N1855);
or OR2 (N3672, N3670, N533);
buf BUF1 (N3673, N3659);
or OR3 (N3674, N3672, N2352, N3311);
nand NAND3 (N3675, N3660, N34, N971);
nand NAND2 (N3676, N3652, N1802);
nor NOR2 (N3677, N3671, N468);
and AND3 (N3678, N3666, N70, N1204);
or OR3 (N3679, N3676, N954, N156);
and AND2 (N3680, N3674, N540);
nand NAND3 (N3681, N3661, N201, N728);
nand NAND4 (N3682, N3678, N37, N271, N1410);
not NOT1 (N3683, N3673);
nand NAND4 (N3684, N3675, N3243, N1578, N1361);
or OR2 (N3685, N3679, N2437);
nor NOR2 (N3686, N3683, N1119);
xor XOR2 (N3687, N3663, N119);
nand NAND3 (N3688, N3664, N1676, N130);
or OR3 (N3689, N3686, N2676, N1138);
nor NOR3 (N3690, N3688, N2237, N1704);
and AND3 (N3691, N3682, N2524, N2254);
or OR3 (N3692, N3685, N439, N2008);
buf BUF1 (N3693, N3691);
and AND2 (N3694, N3693, N3507);
and AND2 (N3695, N3684, N874);
xor XOR2 (N3696, N3680, N386);
not NOT1 (N3697, N3677);
nand NAND2 (N3698, N3692, N3341);
or OR4 (N3699, N3695, N2164, N1876, N1378);
or OR3 (N3700, N3687, N1858, N649);
xor XOR2 (N3701, N3700, N3672);
xor XOR2 (N3702, N3689, N1111);
buf BUF1 (N3703, N3697);
buf BUF1 (N3704, N3701);
not NOT1 (N3705, N3694);
xor XOR2 (N3706, N3642, N1298);
xor XOR2 (N3707, N3699, N1814);
or OR2 (N3708, N3702, N1799);
not NOT1 (N3709, N3696);
or OR3 (N3710, N3704, N1324, N2057);
or OR4 (N3711, N3705, N356, N89, N293);
or OR2 (N3712, N3698, N3244);
nor NOR4 (N3713, N3707, N1277, N1168, N2030);
or OR2 (N3714, N3713, N2424);
not NOT1 (N3715, N3714);
and AND3 (N3716, N3706, N2504, N664);
not NOT1 (N3717, N3690);
not NOT1 (N3718, N3711);
nand NAND4 (N3719, N3712, N934, N161, N102);
or OR3 (N3720, N3710, N758, N2273);
not NOT1 (N3721, N3717);
nor NOR3 (N3722, N3716, N2076, N2024);
or OR2 (N3723, N3715, N2324);
buf BUF1 (N3724, N3722);
nand NAND4 (N3725, N3709, N3201, N254, N1801);
or OR2 (N3726, N3718, N3150);
buf BUF1 (N3727, N3725);
nand NAND4 (N3728, N3724, N2078, N287, N3532);
and AND4 (N3729, N3726, N2624, N3384, N2845);
not NOT1 (N3730, N3729);
nor NOR4 (N3731, N3703, N1213, N1394, N124);
nand NAND2 (N3732, N3731, N186);
and AND2 (N3733, N3732, N1578);
nor NOR3 (N3734, N3719, N3158, N2342);
xor XOR2 (N3735, N3730, N3268);
buf BUF1 (N3736, N3734);
xor XOR2 (N3737, N3681, N1712);
nand NAND3 (N3738, N3733, N340, N707);
nand NAND2 (N3739, N3736, N1030);
not NOT1 (N3740, N3728);
xor XOR2 (N3741, N3708, N2984);
not NOT1 (N3742, N3738);
or OR4 (N3743, N3739, N553, N2066, N2117);
nand NAND2 (N3744, N3727, N1692);
and AND2 (N3745, N3720, N3173);
and AND3 (N3746, N3737, N1306, N93);
and AND4 (N3747, N3723, N82, N731, N1622);
and AND2 (N3748, N3740, N1289);
and AND3 (N3749, N3743, N2728, N3551);
xor XOR2 (N3750, N3744, N3348);
or OR3 (N3751, N3749, N1952, N1829);
and AND3 (N3752, N3748, N2016, N1325);
and AND3 (N3753, N3752, N676, N2881);
nor NOR2 (N3754, N3753, N2830);
and AND2 (N3755, N3741, N162);
xor XOR2 (N3756, N3750, N2502);
nand NAND4 (N3757, N3747, N2167, N985, N2434);
nand NAND4 (N3758, N3757, N1742, N301, N1286);
nand NAND2 (N3759, N3745, N1992);
nor NOR2 (N3760, N3754, N2724);
or OR4 (N3761, N3751, N374, N237, N2151);
not NOT1 (N3762, N3760);
nor NOR4 (N3763, N3756, N3485, N3020, N2354);
nor NOR3 (N3764, N3758, N3613, N3723);
buf BUF1 (N3765, N3764);
not NOT1 (N3766, N3759);
or OR4 (N3767, N3742, N1980, N541, N3624);
xor XOR2 (N3768, N3765, N1131);
not NOT1 (N3769, N3746);
nor NOR3 (N3770, N3768, N393, N825);
buf BUF1 (N3771, N3762);
not NOT1 (N3772, N3767);
nand NAND2 (N3773, N3770, N347);
nand NAND3 (N3774, N3761, N829, N382);
buf BUF1 (N3775, N3721);
or OR3 (N3776, N3769, N2794, N531);
nand NAND3 (N3777, N3771, N657, N636);
not NOT1 (N3778, N3777);
buf BUF1 (N3779, N3778);
or OR3 (N3780, N3766, N463, N2009);
buf BUF1 (N3781, N3775);
nand NAND2 (N3782, N3755, N3514);
nand NAND3 (N3783, N3780, N2822, N1123);
and AND2 (N3784, N3772, N584);
not NOT1 (N3785, N3776);
and AND3 (N3786, N3782, N1270, N184);
not NOT1 (N3787, N3763);
or OR2 (N3788, N3783, N2483);
nor NOR2 (N3789, N3781, N3382);
buf BUF1 (N3790, N3787);
buf BUF1 (N3791, N3784);
or OR4 (N3792, N3774, N998, N256, N2247);
or OR3 (N3793, N3735, N1334, N968);
nand NAND3 (N3794, N3790, N1467, N3502);
and AND3 (N3795, N3773, N3714, N129);
or OR2 (N3796, N3785, N2323);
and AND2 (N3797, N3789, N910);
nand NAND4 (N3798, N3795, N372, N2505, N3258);
buf BUF1 (N3799, N3791);
buf BUF1 (N3800, N3796);
buf BUF1 (N3801, N3800);
xor XOR2 (N3802, N3801, N2730);
or OR2 (N3803, N3793, N1204);
nor NOR3 (N3804, N3779, N1115, N316);
xor XOR2 (N3805, N3797, N2085);
not NOT1 (N3806, N3794);
and AND2 (N3807, N3802, N1324);
or OR4 (N3808, N3799, N2228, N825, N926);
nand NAND2 (N3809, N3808, N2857);
nand NAND3 (N3810, N3788, N1455, N2827);
xor XOR2 (N3811, N3809, N2195);
nand NAND3 (N3812, N3804, N1719, N3697);
xor XOR2 (N3813, N3786, N1220);
not NOT1 (N3814, N3807);
and AND4 (N3815, N3803, N3087, N3083, N2499);
nand NAND3 (N3816, N3811, N1279, N3169);
nand NAND3 (N3817, N3816, N2379, N724);
nand NAND3 (N3818, N3812, N3732, N2534);
or OR4 (N3819, N3792, N2546, N633, N798);
buf BUF1 (N3820, N3806);
and AND4 (N3821, N3798, N2384, N3521, N461);
not NOT1 (N3822, N3818);
buf BUF1 (N3823, N3810);
not NOT1 (N3824, N3822);
xor XOR2 (N3825, N3813, N2746);
xor XOR2 (N3826, N3823, N395);
xor XOR2 (N3827, N3805, N2218);
xor XOR2 (N3828, N3821, N2261);
not NOT1 (N3829, N3817);
buf BUF1 (N3830, N3829);
not NOT1 (N3831, N3828);
and AND4 (N3832, N3830, N1691, N2452, N1895);
or OR4 (N3833, N3826, N3739, N826, N813);
and AND3 (N3834, N3814, N2058, N2487);
nand NAND3 (N3835, N3824, N1486, N3204);
xor XOR2 (N3836, N3820, N159);
nor NOR3 (N3837, N3819, N2730, N3491);
or OR2 (N3838, N3831, N2230);
or OR2 (N3839, N3837, N3607);
nor NOR3 (N3840, N3838, N546, N2650);
xor XOR2 (N3841, N3825, N3585);
nor NOR4 (N3842, N3815, N1023, N765, N1277);
xor XOR2 (N3843, N3840, N3564);
buf BUF1 (N3844, N3833);
nand NAND4 (N3845, N3835, N2069, N3515, N3355);
and AND2 (N3846, N3834, N3266);
buf BUF1 (N3847, N3841);
xor XOR2 (N3848, N3832, N1479);
nor NOR2 (N3849, N3842, N1693);
xor XOR2 (N3850, N3839, N3065);
or OR2 (N3851, N3844, N3006);
xor XOR2 (N3852, N3847, N633);
not NOT1 (N3853, N3852);
nor NOR4 (N3854, N3853, N994, N3145, N2363);
buf BUF1 (N3855, N3849);
not NOT1 (N3856, N3827);
and AND3 (N3857, N3854, N2939, N506);
not NOT1 (N3858, N3850);
and AND2 (N3859, N3836, N1603);
not NOT1 (N3860, N3855);
xor XOR2 (N3861, N3860, N2591);
buf BUF1 (N3862, N3845);
not NOT1 (N3863, N3861);
nand NAND2 (N3864, N3846, N3284);
or OR3 (N3865, N3859, N1598, N3308);
xor XOR2 (N3866, N3864, N1240);
buf BUF1 (N3867, N3848);
xor XOR2 (N3868, N3863, N501);
or OR3 (N3869, N3851, N122, N1748);
and AND3 (N3870, N3865, N119, N1172);
nand NAND3 (N3871, N3857, N3120, N1948);
buf BUF1 (N3872, N3871);
or OR3 (N3873, N3866, N1971, N79);
or OR4 (N3874, N3843, N1137, N1644, N3747);
nor NOR3 (N3875, N3874, N2043, N1182);
or OR2 (N3876, N3869, N418);
xor XOR2 (N3877, N3862, N821);
xor XOR2 (N3878, N3873, N3543);
nand NAND2 (N3879, N3870, N3064);
nand NAND4 (N3880, N3878, N2811, N72, N2011);
nor NOR2 (N3881, N3867, N3802);
nand NAND2 (N3882, N3880, N2317);
buf BUF1 (N3883, N3868);
nand NAND3 (N3884, N3875, N9, N2224);
buf BUF1 (N3885, N3883);
not NOT1 (N3886, N3858);
xor XOR2 (N3887, N3882, N2803);
or OR3 (N3888, N3886, N3617, N392);
not NOT1 (N3889, N3872);
not NOT1 (N3890, N3887);
nor NOR4 (N3891, N3856, N3376, N1080, N2922);
nor NOR2 (N3892, N3891, N1371);
or OR3 (N3893, N3884, N3644, N2930);
buf BUF1 (N3894, N3890);
nor NOR2 (N3895, N3892, N3091);
not NOT1 (N3896, N3881);
or OR3 (N3897, N3889, N745, N3144);
xor XOR2 (N3898, N3885, N2718);
xor XOR2 (N3899, N3897, N2425);
buf BUF1 (N3900, N3894);
xor XOR2 (N3901, N3899, N1644);
xor XOR2 (N3902, N3898, N1108);
buf BUF1 (N3903, N3893);
not NOT1 (N3904, N3888);
and AND2 (N3905, N3904, N2730);
or OR2 (N3906, N3896, N787);
xor XOR2 (N3907, N3905, N451);
buf BUF1 (N3908, N3900);
xor XOR2 (N3909, N3879, N1601);
or OR4 (N3910, N3908, N2043, N3308, N2519);
nor NOR3 (N3911, N3876, N222, N3780);
nor NOR4 (N3912, N3910, N1880, N543, N1946);
nor NOR4 (N3913, N3909, N3429, N1309, N3005);
or OR2 (N3914, N3901, N1956);
nor NOR2 (N3915, N3912, N1034);
nand NAND2 (N3916, N3907, N1708);
or OR2 (N3917, N3911, N2233);
buf BUF1 (N3918, N3877);
not NOT1 (N3919, N3918);
not NOT1 (N3920, N3906);
or OR4 (N3921, N3915, N1359, N2120, N902);
buf BUF1 (N3922, N3914);
and AND3 (N3923, N3922, N2842, N2912);
xor XOR2 (N3924, N3916, N2185);
nor NOR4 (N3925, N3920, N2794, N3204, N258);
and AND2 (N3926, N3921, N2572);
buf BUF1 (N3927, N3902);
buf BUF1 (N3928, N3925);
not NOT1 (N3929, N3928);
xor XOR2 (N3930, N3923, N66);
nand NAND4 (N3931, N3919, N3001, N2849, N664);
and AND4 (N3932, N3929, N732, N1561, N2170);
nor NOR2 (N3933, N3913, N300);
not NOT1 (N3934, N3930);
and AND4 (N3935, N3926, N970, N808, N2939);
and AND4 (N3936, N3935, N441, N3543, N1328);
or OR2 (N3937, N3931, N1707);
and AND2 (N3938, N3924, N1507);
buf BUF1 (N3939, N3938);
nor NOR4 (N3940, N3933, N1955, N2016, N1102);
nand NAND4 (N3941, N3936, N3806, N3076, N2944);
not NOT1 (N3942, N3927);
not NOT1 (N3943, N3939);
and AND2 (N3944, N3917, N583);
nand NAND3 (N3945, N3895, N1992, N249);
nand NAND3 (N3946, N3944, N2855, N1174);
xor XOR2 (N3947, N3945, N3011);
nand NAND3 (N3948, N3932, N474, N3695);
and AND3 (N3949, N3943, N2919, N2969);
or OR2 (N3950, N3934, N3336);
and AND3 (N3951, N3948, N1048, N2836);
or OR2 (N3952, N3949, N902);
buf BUF1 (N3953, N3937);
or OR3 (N3954, N3946, N2788, N741);
and AND4 (N3955, N3951, N3364, N3679, N2733);
not NOT1 (N3956, N3955);
buf BUF1 (N3957, N3952);
nand NAND3 (N3958, N3953, N3357, N237);
and AND2 (N3959, N3954, N329);
not NOT1 (N3960, N3950);
xor XOR2 (N3961, N3941, N2751);
buf BUF1 (N3962, N3940);
and AND2 (N3963, N3960, N705);
not NOT1 (N3964, N3947);
xor XOR2 (N3965, N3964, N3638);
nand NAND4 (N3966, N3959, N796, N829, N2270);
or OR3 (N3967, N3903, N679, N421);
buf BUF1 (N3968, N3958);
and AND3 (N3969, N3963, N1381, N1931);
nand NAND4 (N3970, N3962, N1540, N1592, N460);
not NOT1 (N3971, N3957);
nor NOR3 (N3972, N3942, N3671, N2815);
not NOT1 (N3973, N3970);
or OR3 (N3974, N3969, N541, N1515);
and AND4 (N3975, N3971, N3408, N3510, N1316);
xor XOR2 (N3976, N3968, N3038);
buf BUF1 (N3977, N3973);
and AND4 (N3978, N3966, N1594, N490, N3294);
xor XOR2 (N3979, N3978, N94);
buf BUF1 (N3980, N3965);
and AND3 (N3981, N3979, N3476, N1200);
nand NAND4 (N3982, N3967, N2982, N1685, N311);
or OR3 (N3983, N3961, N1555, N1189);
and AND3 (N3984, N3976, N1951, N3010);
and AND3 (N3985, N3980, N2369, N3594);
buf BUF1 (N3986, N3974);
not NOT1 (N3987, N3984);
and AND2 (N3988, N3987, N994);
or OR2 (N3989, N3986, N433);
or OR3 (N3990, N3975, N1868, N1489);
and AND3 (N3991, N3985, N3536, N582);
nand NAND2 (N3992, N3981, N2758);
nor NOR3 (N3993, N3983, N3540, N930);
nor NOR2 (N3994, N3990, N1965);
buf BUF1 (N3995, N3956);
and AND4 (N3996, N3992, N2924, N3204, N460);
or OR2 (N3997, N3996, N589);
xor XOR2 (N3998, N3993, N2630);
xor XOR2 (N3999, N3998, N1583);
nand NAND3 (N4000, N3972, N1120, N1939);
nand NAND4 (N4001, N3997, N2757, N1166, N2331);
not NOT1 (N4002, N4000);
or OR4 (N4003, N3995, N313, N3359, N2983);
not NOT1 (N4004, N4002);
not NOT1 (N4005, N3988);
or OR4 (N4006, N3982, N2506, N3089, N1951);
nand NAND3 (N4007, N4003, N3403, N1438);
not NOT1 (N4008, N3977);
and AND3 (N4009, N3991, N2420, N3803);
nor NOR2 (N4010, N4005, N2024);
xor XOR2 (N4011, N4009, N253);
and AND2 (N4012, N4004, N2122);
nand NAND4 (N4013, N3999, N2522, N2216, N2437);
not NOT1 (N4014, N4012);
buf BUF1 (N4015, N4006);
and AND2 (N4016, N3989, N2879);
nor NOR4 (N4017, N4011, N551, N284, N2907);
nor NOR3 (N4018, N4007, N3288, N3236);
nor NOR2 (N4019, N4017, N2495);
buf BUF1 (N4020, N3994);
nand NAND4 (N4021, N4019, N1124, N3102, N1623);
or OR3 (N4022, N4021, N1945, N1138);
and AND4 (N4023, N4013, N561, N2195, N1943);
nor NOR3 (N4024, N4001, N1454, N3624);
and AND3 (N4025, N4015, N2651, N1480);
not NOT1 (N4026, N4016);
nor NOR4 (N4027, N4020, N3660, N580, N726);
or OR4 (N4028, N4027, N2781, N1626, N236);
nor NOR3 (N4029, N4010, N2166, N2351);
not NOT1 (N4030, N4026);
nor NOR2 (N4031, N4018, N3878);
nand NAND4 (N4032, N4022, N1203, N1223, N1484);
not NOT1 (N4033, N4031);
buf BUF1 (N4034, N4023);
nand NAND4 (N4035, N4025, N616, N79, N3677);
and AND4 (N4036, N4024, N2259, N1826, N690);
or OR2 (N4037, N4030, N1058);
and AND4 (N4038, N4037, N3508, N1761, N2265);
and AND2 (N4039, N4038, N2309);
xor XOR2 (N4040, N4032, N243);
and AND2 (N4041, N4029, N1130);
or OR3 (N4042, N4040, N1666, N1229);
not NOT1 (N4043, N4042);
and AND4 (N4044, N4033, N2563, N1048, N1299);
and AND2 (N4045, N4014, N1818);
and AND2 (N4046, N4035, N2382);
xor XOR2 (N4047, N4046, N3725);
nor NOR3 (N4048, N4047, N1828, N3033);
xor XOR2 (N4049, N4043, N2639);
buf BUF1 (N4050, N4034);
xor XOR2 (N4051, N4028, N2631);
and AND2 (N4052, N4048, N447);
nand NAND2 (N4053, N4008, N2626);
or OR2 (N4054, N4045, N23);
nand NAND2 (N4055, N4036, N3922);
nor NOR2 (N4056, N4055, N3928);
not NOT1 (N4057, N4039);
and AND3 (N4058, N4053, N619, N1429);
nor NOR4 (N4059, N4052, N883, N4052, N1377);
and AND2 (N4060, N4044, N1510);
nand NAND4 (N4061, N4049, N1513, N3409, N940);
not NOT1 (N4062, N4060);
not NOT1 (N4063, N4050);
nand NAND3 (N4064, N4062, N3782, N1664);
nor NOR2 (N4065, N4064, N3922);
nor NOR3 (N4066, N4059, N1652, N1064);
nand NAND4 (N4067, N4041, N1085, N742, N700);
nand NAND4 (N4068, N4051, N1794, N3118, N1228);
nand NAND3 (N4069, N4066, N3275, N476);
xor XOR2 (N4070, N4065, N309);
or OR3 (N4071, N4061, N2400, N1088);
not NOT1 (N4072, N4068);
nand NAND2 (N4073, N4067, N2433);
xor XOR2 (N4074, N4069, N249);
buf BUF1 (N4075, N4072);
not NOT1 (N4076, N4063);
nor NOR2 (N4077, N4057, N2123);
not NOT1 (N4078, N4070);
or OR3 (N4079, N4073, N3348, N1112);
xor XOR2 (N4080, N4058, N2656);
nor NOR2 (N4081, N4079, N234);
or OR3 (N4082, N4080, N1100, N577);
and AND4 (N4083, N4082, N1262, N464, N892);
nand NAND3 (N4084, N4078, N519, N754);
and AND2 (N4085, N4056, N957);
nand NAND4 (N4086, N4085, N2840, N2134, N1393);
nand NAND2 (N4087, N4054, N1712);
and AND4 (N4088, N4071, N4039, N170, N2830);
nand NAND2 (N4089, N4086, N3909);
and AND2 (N4090, N4081, N2060);
and AND3 (N4091, N4075, N3415, N2053);
not NOT1 (N4092, N4074);
and AND4 (N4093, N4092, N2396, N2486, N382);
buf BUF1 (N4094, N4077);
nand NAND2 (N4095, N4083, N1022);
or OR4 (N4096, N4076, N2406, N2947, N1157);
or OR2 (N4097, N4087, N185);
buf BUF1 (N4098, N4094);
not NOT1 (N4099, N4091);
and AND4 (N4100, N4096, N2701, N2031, N1928);
or OR4 (N4101, N4093, N1484, N3752, N1415);
not NOT1 (N4102, N4097);
or OR3 (N4103, N4090, N2339, N1602);
not NOT1 (N4104, N4103);
or OR3 (N4105, N4095, N2052, N3101);
nor NOR4 (N4106, N4099, N779, N3534, N3718);
nand NAND3 (N4107, N4101, N1961, N3243);
buf BUF1 (N4108, N4088);
or OR2 (N4109, N4100, N3181);
and AND4 (N4110, N4102, N761, N1615, N1591);
or OR3 (N4111, N4098, N1469, N1904);
or OR3 (N4112, N4110, N1811, N1323);
xor XOR2 (N4113, N4108, N1503);
buf BUF1 (N4114, N4104);
xor XOR2 (N4115, N4109, N1031);
nand NAND4 (N4116, N4105, N641, N1844, N941);
nor NOR4 (N4117, N4084, N1030, N2702, N2490);
nand NAND2 (N4118, N4107, N4100);
nand NAND2 (N4119, N4106, N488);
nand NAND3 (N4120, N4112, N1342, N1913);
nor NOR3 (N4121, N4113, N3761, N2223);
xor XOR2 (N4122, N4121, N2448);
and AND4 (N4123, N4115, N3867, N3583, N242);
or OR3 (N4124, N4114, N2896, N1079);
and AND3 (N4125, N4116, N633, N2033);
xor XOR2 (N4126, N4123, N3873);
or OR4 (N4127, N4111, N3740, N506, N708);
nor NOR4 (N4128, N4119, N3924, N464, N3060);
buf BUF1 (N4129, N4126);
nand NAND2 (N4130, N4128, N829);
nand NAND3 (N4131, N4117, N4079, N208);
and AND4 (N4132, N4118, N1890, N3925, N3458);
and AND3 (N4133, N4122, N875, N3328);
or OR2 (N4134, N4133, N3047);
nor NOR2 (N4135, N4127, N1659);
xor XOR2 (N4136, N4132, N2391);
not NOT1 (N4137, N4129);
and AND4 (N4138, N4136, N1528, N4135, N3004);
nor NOR4 (N4139, N1477, N3473, N144, N3704);
buf BUF1 (N4140, N4089);
nor NOR2 (N4141, N4138, N2936);
nor NOR3 (N4142, N4141, N2486, N1154);
not NOT1 (N4143, N4142);
and AND3 (N4144, N4139, N1072, N2193);
or OR3 (N4145, N4140, N950, N146);
buf BUF1 (N4146, N4130);
nand NAND2 (N4147, N4124, N2436);
xor XOR2 (N4148, N4147, N2861);
buf BUF1 (N4149, N4134);
buf BUF1 (N4150, N4148);
or OR3 (N4151, N4150, N1189, N3819);
nand NAND2 (N4152, N4131, N236);
nand NAND2 (N4153, N4144, N1000);
buf BUF1 (N4154, N4146);
nor NOR4 (N4155, N4149, N711, N25, N1878);
or OR2 (N4156, N4153, N1248);
nor NOR3 (N4157, N4152, N3767, N3396);
buf BUF1 (N4158, N4125);
xor XOR2 (N4159, N4120, N3026);
nand NAND3 (N4160, N4145, N2670, N2388);
buf BUF1 (N4161, N4154);
xor XOR2 (N4162, N4158, N2380);
and AND3 (N4163, N4137, N2757, N492);
not NOT1 (N4164, N4156);
not NOT1 (N4165, N4164);
and AND3 (N4166, N4143, N2628, N686);
nand NAND4 (N4167, N4161, N1425, N1766, N2771);
and AND3 (N4168, N4160, N849, N1967);
not NOT1 (N4169, N4168);
and AND2 (N4170, N4163, N3852);
nor NOR3 (N4171, N4169, N3465, N2618);
nand NAND2 (N4172, N4159, N3048);
nand NAND4 (N4173, N4172, N44, N3585, N4067);
or OR4 (N4174, N4171, N3139, N2555, N3867);
and AND3 (N4175, N4162, N737, N2337);
buf BUF1 (N4176, N4170);
nor NOR4 (N4177, N4165, N241, N749, N837);
or OR4 (N4178, N4167, N2286, N893, N2997);
and AND4 (N4179, N4177, N685, N736, N3361);
nand NAND2 (N4180, N4151, N3647);
and AND2 (N4181, N4180, N1850);
xor XOR2 (N4182, N4166, N4171);
and AND3 (N4183, N4173, N1357, N2311);
xor XOR2 (N4184, N4178, N23);
not NOT1 (N4185, N4174);
not NOT1 (N4186, N4157);
buf BUF1 (N4187, N4155);
and AND4 (N4188, N4183, N920, N680, N3409);
buf BUF1 (N4189, N4187);
nor NOR2 (N4190, N4189, N1968);
and AND2 (N4191, N4179, N2222);
nor NOR3 (N4192, N4175, N17, N2950);
buf BUF1 (N4193, N4188);
buf BUF1 (N4194, N4190);
nor NOR2 (N4195, N4181, N588);
xor XOR2 (N4196, N4191, N2955);
nor NOR2 (N4197, N4196, N2204);
or OR2 (N4198, N4193, N3160);
buf BUF1 (N4199, N4197);
xor XOR2 (N4200, N4176, N2559);
xor XOR2 (N4201, N4194, N2025);
nor NOR4 (N4202, N4182, N1389, N1084, N1450);
or OR2 (N4203, N4200, N69);
or OR4 (N4204, N4195, N4180, N3921, N97);
not NOT1 (N4205, N4201);
xor XOR2 (N4206, N4202, N3998);
nor NOR4 (N4207, N4184, N3294, N1977, N3355);
nand NAND4 (N4208, N4206, N1472, N869, N3226);
nand NAND2 (N4209, N4208, N2817);
or OR2 (N4210, N4185, N2118);
or OR2 (N4211, N4210, N2395);
not NOT1 (N4212, N4199);
xor XOR2 (N4213, N4203, N1988);
and AND3 (N4214, N4204, N439, N1813);
or OR2 (N4215, N4211, N3493);
nand NAND4 (N4216, N4214, N2440, N2253, N2236);
and AND3 (N4217, N4205, N3642, N273);
or OR3 (N4218, N4207, N4107, N827);
nand NAND4 (N4219, N4216, N2435, N1940, N1443);
buf BUF1 (N4220, N4209);
nand NAND2 (N4221, N4212, N3318);
not NOT1 (N4222, N4221);
not NOT1 (N4223, N4218);
buf BUF1 (N4224, N4192);
buf BUF1 (N4225, N4220);
or OR4 (N4226, N4219, N257, N2403, N3588);
or OR2 (N4227, N4223, N188);
xor XOR2 (N4228, N4225, N1586);
and AND4 (N4229, N4228, N517, N628, N3403);
buf BUF1 (N4230, N4198);
buf BUF1 (N4231, N4222);
not NOT1 (N4232, N4230);
or OR3 (N4233, N4224, N2855, N1099);
and AND3 (N4234, N4215, N1792, N2121);
nand NAND4 (N4235, N4227, N2954, N3101, N3696);
and AND3 (N4236, N4229, N1111, N1590);
buf BUF1 (N4237, N4236);
nor NOR3 (N4238, N4237, N3407, N1302);
xor XOR2 (N4239, N4217, N610);
and AND3 (N4240, N4232, N930, N2645);
buf BUF1 (N4241, N4186);
nand NAND3 (N4242, N4226, N3001, N36);
not NOT1 (N4243, N4213);
nor NOR2 (N4244, N4242, N2016);
nor NOR3 (N4245, N4244, N4065, N588);
nand NAND4 (N4246, N4235, N2714, N3134, N1845);
not NOT1 (N4247, N4234);
nor NOR4 (N4248, N4247, N709, N1438, N3624);
not NOT1 (N4249, N4231);
buf BUF1 (N4250, N4246);
or OR2 (N4251, N4241, N1508);
buf BUF1 (N4252, N4251);
or OR2 (N4253, N4248, N1029);
and AND3 (N4254, N4249, N3000, N2715);
and AND3 (N4255, N4245, N1273, N1753);
nor NOR3 (N4256, N4255, N2022, N3247);
or OR3 (N4257, N4250, N4041, N3406);
not NOT1 (N4258, N4240);
not NOT1 (N4259, N4243);
nand NAND2 (N4260, N4252, N272);
xor XOR2 (N4261, N4257, N918);
nand NAND2 (N4262, N4239, N2137);
not NOT1 (N4263, N4259);
and AND4 (N4264, N4233, N1195, N1187, N3454);
xor XOR2 (N4265, N4264, N3942);
nor NOR2 (N4266, N4258, N664);
and AND3 (N4267, N4238, N696, N2690);
not NOT1 (N4268, N4266);
and AND4 (N4269, N4261, N1749, N4159, N22);
and AND4 (N4270, N4267, N2812, N3332, N3459);
buf BUF1 (N4271, N4256);
nand NAND3 (N4272, N4260, N596, N3073);
and AND2 (N4273, N4271, N1400);
nor NOR2 (N4274, N4263, N2748);
nor NOR4 (N4275, N4274, N2607, N3806, N3340);
xor XOR2 (N4276, N4262, N2329);
or OR3 (N4277, N4269, N3817, N502);
buf BUF1 (N4278, N4275);
not NOT1 (N4279, N4270);
nor NOR4 (N4280, N4268, N3728, N3498, N2603);
or OR3 (N4281, N4273, N3264, N6);
buf BUF1 (N4282, N4253);
and AND2 (N4283, N4278, N801);
not NOT1 (N4284, N4281);
nand NAND3 (N4285, N4282, N295, N3003);
nand NAND4 (N4286, N4277, N481, N1903, N1955);
or OR4 (N4287, N4283, N4255, N3886, N561);
buf BUF1 (N4288, N4284);
not NOT1 (N4289, N4288);
and AND3 (N4290, N4272, N17, N1602);
buf BUF1 (N4291, N4287);
xor XOR2 (N4292, N4280, N120);
not NOT1 (N4293, N4286);
nand NAND4 (N4294, N4254, N3922, N80, N2193);
nand NAND3 (N4295, N4292, N623, N693);
not NOT1 (N4296, N4265);
xor XOR2 (N4297, N4295, N3992);
nor NOR2 (N4298, N4294, N307);
nand NAND3 (N4299, N4289, N2262, N2074);
xor XOR2 (N4300, N4293, N3504);
buf BUF1 (N4301, N4297);
and AND4 (N4302, N4300, N2253, N2360, N1068);
and AND2 (N4303, N4302, N2786);
not NOT1 (N4304, N4279);
buf BUF1 (N4305, N4290);
nor NOR2 (N4306, N4299, N1153);
and AND3 (N4307, N4306, N4013, N2458);
or OR3 (N4308, N4291, N3956, N174);
and AND2 (N4309, N4304, N3947);
nor NOR2 (N4310, N4285, N1965);
or OR4 (N4311, N4276, N3128, N3293, N2800);
buf BUF1 (N4312, N4307);
not NOT1 (N4313, N4298);
xor XOR2 (N4314, N4308, N3113);
buf BUF1 (N4315, N4311);
not NOT1 (N4316, N4314);
buf BUF1 (N4317, N4316);
buf BUF1 (N4318, N4312);
or OR4 (N4319, N4309, N3674, N2570, N1707);
and AND4 (N4320, N4318, N925, N2307, N3788);
not NOT1 (N4321, N4303);
buf BUF1 (N4322, N4305);
xor XOR2 (N4323, N4315, N3565);
not NOT1 (N4324, N4320);
buf BUF1 (N4325, N4296);
buf BUF1 (N4326, N4323);
nand NAND4 (N4327, N4319, N4034, N3535, N63);
or OR2 (N4328, N4324, N3284);
xor XOR2 (N4329, N4325, N2866);
and AND4 (N4330, N4317, N4193, N3334, N2250);
nand NAND3 (N4331, N4301, N310, N927);
not NOT1 (N4332, N4310);
not NOT1 (N4333, N4331);
nand NAND2 (N4334, N4332, N1964);
and AND4 (N4335, N4328, N1381, N1463, N2991);
buf BUF1 (N4336, N4327);
and AND3 (N4337, N4335, N1682, N3692);
not NOT1 (N4338, N4333);
buf BUF1 (N4339, N4322);
and AND4 (N4340, N4326, N2528, N876, N984);
or OR2 (N4341, N4334, N2552);
not NOT1 (N4342, N4340);
or OR3 (N4343, N4337, N383, N3909);
and AND4 (N4344, N4341, N921, N2317, N1067);
buf BUF1 (N4345, N4343);
xor XOR2 (N4346, N4313, N1950);
buf BUF1 (N4347, N4336);
not NOT1 (N4348, N4342);
not NOT1 (N4349, N4321);
nor NOR3 (N4350, N4329, N1900, N1391);
buf BUF1 (N4351, N4344);
xor XOR2 (N4352, N4338, N2702);
and AND2 (N4353, N4349, N487);
xor XOR2 (N4354, N4350, N587);
not NOT1 (N4355, N4351);
and AND3 (N4356, N4353, N1976, N1108);
or OR2 (N4357, N4352, N2538);
not NOT1 (N4358, N4345);
and AND2 (N4359, N4330, N424);
nand NAND2 (N4360, N4347, N1775);
nor NOR4 (N4361, N4355, N918, N512, N4062);
or OR2 (N4362, N4359, N2612);
and AND4 (N4363, N4356, N3632, N2153, N2605);
buf BUF1 (N4364, N4357);
and AND2 (N4365, N4360, N4007);
or OR3 (N4366, N4348, N1366, N3396);
nor NOR3 (N4367, N4366, N1915, N1974);
buf BUF1 (N4368, N4364);
and AND3 (N4369, N4368, N1545, N1430);
buf BUF1 (N4370, N4369);
buf BUF1 (N4371, N4362);
xor XOR2 (N4372, N4365, N4016);
xor XOR2 (N4373, N4339, N539);
nor NOR3 (N4374, N4370, N3321, N3571);
xor XOR2 (N4375, N4373, N3964);
not NOT1 (N4376, N4372);
nand NAND3 (N4377, N4361, N3230, N225);
not NOT1 (N4378, N4376);
not NOT1 (N4379, N4375);
xor XOR2 (N4380, N4371, N2915);
buf BUF1 (N4381, N4374);
not NOT1 (N4382, N4367);
nor NOR3 (N4383, N4363, N318, N3570);
nand NAND2 (N4384, N4379, N1059);
nand NAND3 (N4385, N4381, N697, N1685);
buf BUF1 (N4386, N4385);
xor XOR2 (N4387, N4354, N3289);
nor NOR3 (N4388, N4358, N3611, N221);
xor XOR2 (N4389, N4380, N265);
or OR4 (N4390, N4387, N948, N2366, N167);
xor XOR2 (N4391, N4388, N4236);
xor XOR2 (N4392, N4382, N412);
or OR3 (N4393, N4346, N397, N2455);
and AND4 (N4394, N4378, N3956, N2467, N4040);
not NOT1 (N4395, N4393);
xor XOR2 (N4396, N4394, N2703);
or OR3 (N4397, N4386, N1765, N2171);
xor XOR2 (N4398, N4377, N320);
not NOT1 (N4399, N4383);
nand NAND4 (N4400, N4396, N2417, N4100, N580);
or OR4 (N4401, N4389, N483, N563, N1491);
and AND4 (N4402, N4391, N3245, N2193, N2758);
xor XOR2 (N4403, N4395, N3213);
not NOT1 (N4404, N4392);
buf BUF1 (N4405, N4402);
not NOT1 (N4406, N4390);
nand NAND3 (N4407, N4403, N1861, N588);
and AND2 (N4408, N4404, N621);
not NOT1 (N4409, N4405);
buf BUF1 (N4410, N4406);
or OR4 (N4411, N4384, N2823, N2180, N1917);
nand NAND4 (N4412, N4407, N2405, N2470, N2385);
nor NOR4 (N4413, N4399, N1383, N1328, N498);
not NOT1 (N4414, N4413);
xor XOR2 (N4415, N4409, N4233);
xor XOR2 (N4416, N4411, N2149);
and AND2 (N4417, N4408, N2886);
nand NAND2 (N4418, N4397, N1649);
nand NAND2 (N4419, N4400, N1101);
or OR4 (N4420, N4398, N3882, N428, N3961);
xor XOR2 (N4421, N4418, N2951);
not NOT1 (N4422, N4414);
buf BUF1 (N4423, N4416);
and AND3 (N4424, N4415, N2386, N794);
or OR4 (N4425, N4401, N625, N2881, N3468);
or OR3 (N4426, N4417, N1545, N2807);
buf BUF1 (N4427, N4425);
xor XOR2 (N4428, N4412, N641);
nor NOR4 (N4429, N4426, N2332, N25, N1707);
not NOT1 (N4430, N4423);
xor XOR2 (N4431, N4421, N3002);
nor NOR3 (N4432, N4431, N302, N2508);
and AND3 (N4433, N4420, N3940, N618);
and AND3 (N4434, N4419, N586, N89);
not NOT1 (N4435, N4433);
and AND3 (N4436, N4428, N3936, N171);
and AND4 (N4437, N4410, N537, N139, N982);
buf BUF1 (N4438, N4430);
or OR2 (N4439, N4434, N2609);
or OR4 (N4440, N4436, N4283, N408, N3826);
not NOT1 (N4441, N4424);
and AND3 (N4442, N4440, N1004, N3675);
nor NOR3 (N4443, N4429, N1368, N1534);
buf BUF1 (N4444, N4427);
xor XOR2 (N4445, N4437, N3178);
nor NOR3 (N4446, N4435, N3630, N1895);
xor XOR2 (N4447, N4446, N1410);
buf BUF1 (N4448, N4438);
buf BUF1 (N4449, N4432);
nand NAND3 (N4450, N4447, N87, N1424);
not NOT1 (N4451, N4450);
or OR2 (N4452, N4444, N3729);
and AND3 (N4453, N4439, N2707, N2243);
and AND2 (N4454, N4453, N3683);
nand NAND2 (N4455, N4451, N4109);
xor XOR2 (N4456, N4442, N2387);
or OR2 (N4457, N4449, N2820);
buf BUF1 (N4458, N4445);
not NOT1 (N4459, N4452);
or OR2 (N4460, N4458, N2389);
and AND3 (N4461, N4457, N2846, N248);
xor XOR2 (N4462, N4460, N3307);
not NOT1 (N4463, N4443);
nor NOR2 (N4464, N4462, N2276);
and AND3 (N4465, N4456, N2758, N3651);
not NOT1 (N4466, N4454);
nand NAND3 (N4467, N4455, N2604, N1924);
or OR4 (N4468, N4448, N1411, N3768, N2431);
buf BUF1 (N4469, N4468);
nand NAND4 (N4470, N4467, N1425, N3437, N4451);
not NOT1 (N4471, N4441);
nand NAND3 (N4472, N4469, N3559, N2087);
nor NOR2 (N4473, N4472, N3605);
not NOT1 (N4474, N4465);
or OR3 (N4475, N4459, N2039, N1350);
not NOT1 (N4476, N4473);
or OR3 (N4477, N4463, N3986, N1828);
xor XOR2 (N4478, N4464, N192);
nand NAND3 (N4479, N4471, N3594, N166);
nor NOR4 (N4480, N4466, N2879, N509, N360);
nand NAND3 (N4481, N4478, N1245, N334);
nand NAND3 (N4482, N4470, N795, N1014);
nand NAND4 (N4483, N4476, N399, N332, N3936);
nor NOR4 (N4484, N4482, N2946, N2759, N2957);
nand NAND4 (N4485, N4474, N481, N3236, N129);
not NOT1 (N4486, N4485);
nand NAND2 (N4487, N4475, N2822);
or OR4 (N4488, N4484, N3870, N3979, N285);
not NOT1 (N4489, N4486);
not NOT1 (N4490, N4461);
nor NOR4 (N4491, N4487, N2689, N4453, N4479);
not NOT1 (N4492, N3547);
xor XOR2 (N4493, N4490, N2290);
nand NAND2 (N4494, N4489, N3677);
nor NOR4 (N4495, N4492, N1888, N3120, N4449);
nand NAND3 (N4496, N4480, N3211, N3503);
xor XOR2 (N4497, N4494, N978);
buf BUF1 (N4498, N4493);
and AND4 (N4499, N4497, N4487, N655, N2101);
nor NOR3 (N4500, N4496, N3816, N3210);
nand NAND4 (N4501, N4500, N872, N2545, N2239);
nor NOR3 (N4502, N4499, N2036, N3811);
and AND2 (N4503, N4488, N1557);
xor XOR2 (N4504, N4477, N3491);
buf BUF1 (N4505, N4481);
not NOT1 (N4506, N4505);
nor NOR4 (N4507, N4422, N779, N3541, N2371);
or OR2 (N4508, N4501, N718);
not NOT1 (N4509, N4506);
nor NOR3 (N4510, N4504, N371, N3000);
and AND2 (N4511, N4507, N256);
not NOT1 (N4512, N4511);
xor XOR2 (N4513, N4483, N486);
and AND4 (N4514, N4498, N4195, N4058, N2653);
or OR2 (N4515, N4508, N3310);
buf BUF1 (N4516, N4503);
or OR2 (N4517, N4512, N2082);
or OR4 (N4518, N4509, N464, N3323, N1603);
xor XOR2 (N4519, N4502, N463);
nor NOR2 (N4520, N4519, N695);
and AND4 (N4521, N4513, N610, N174, N3658);
xor XOR2 (N4522, N4515, N2092);
nand NAND2 (N4523, N4491, N2420);
not NOT1 (N4524, N4517);
xor XOR2 (N4525, N4514, N3816);
xor XOR2 (N4526, N4520, N2483);
nand NAND2 (N4527, N4522, N3814);
xor XOR2 (N4528, N4495, N885);
or OR2 (N4529, N4510, N3357);
not NOT1 (N4530, N4528);
not NOT1 (N4531, N4518);
nor NOR4 (N4532, N4526, N4525, N1637, N199);
nor NOR4 (N4533, N3845, N944, N268, N2279);
buf BUF1 (N4534, N4527);
not NOT1 (N4535, N4530);
and AND2 (N4536, N4521, N3348);
buf BUF1 (N4537, N4535);
not NOT1 (N4538, N4537);
and AND2 (N4539, N4516, N4226);
nand NAND4 (N4540, N4536, N3719, N1035, N3403);
or OR3 (N4541, N4540, N674, N2955);
xor XOR2 (N4542, N4533, N1543);
buf BUF1 (N4543, N4531);
and AND4 (N4544, N4534, N2072, N1094, N3537);
not NOT1 (N4545, N4538);
or OR3 (N4546, N4545, N3721, N2995);
nor NOR2 (N4547, N4543, N707);
nand NAND2 (N4548, N4523, N4494);
xor XOR2 (N4549, N4541, N1388);
nand NAND3 (N4550, N4546, N2005, N1887);
xor XOR2 (N4551, N4542, N3777);
nand NAND3 (N4552, N4548, N4413, N2517);
xor XOR2 (N4553, N4539, N2309);
or OR3 (N4554, N4524, N3041, N2803);
nor NOR2 (N4555, N4554, N2878);
nand NAND4 (N4556, N4555, N3856, N4126, N1580);
buf BUF1 (N4557, N4550);
or OR2 (N4558, N4547, N1103);
buf BUF1 (N4559, N4552);
nand NAND3 (N4560, N4553, N1378, N1198);
and AND4 (N4561, N4557, N4403, N2661, N1454);
or OR3 (N4562, N4556, N2671, N3945);
xor XOR2 (N4563, N4561, N4545);
and AND4 (N4564, N4549, N1523, N1876, N685);
nand NAND4 (N4565, N4529, N337, N2534, N4406);
not NOT1 (N4566, N4560);
nand NAND2 (N4567, N4562, N2819);
nor NOR2 (N4568, N4567, N2353);
buf BUF1 (N4569, N4559);
buf BUF1 (N4570, N4551);
xor XOR2 (N4571, N4565, N501);
and AND4 (N4572, N4558, N1223, N2530, N2639);
nand NAND4 (N4573, N4569, N964, N1612, N530);
or OR2 (N4574, N4571, N101);
not NOT1 (N4575, N4574);
nor NOR2 (N4576, N4568, N220);
nor NOR3 (N4577, N4575, N8, N3100);
nor NOR3 (N4578, N4564, N1274, N117);
and AND3 (N4579, N4578, N2496, N2501);
or OR3 (N4580, N4566, N4356, N2157);
buf BUF1 (N4581, N4576);
nand NAND2 (N4582, N4570, N3512);
nand NAND2 (N4583, N4577, N1128);
not NOT1 (N4584, N4532);
buf BUF1 (N4585, N4583);
not NOT1 (N4586, N4582);
nand NAND2 (N4587, N4585, N357);
xor XOR2 (N4588, N4544, N14);
or OR4 (N4589, N4573, N3856, N3834, N2037);
buf BUF1 (N4590, N4563);
not NOT1 (N4591, N4584);
and AND2 (N4592, N4586, N3624);
nand NAND4 (N4593, N4572, N2778, N4300, N604);
not NOT1 (N4594, N4591);
and AND2 (N4595, N4580, N4084);
not NOT1 (N4596, N4587);
and AND2 (N4597, N4592, N3089);
nand NAND2 (N4598, N4594, N1224);
not NOT1 (N4599, N4579);
xor XOR2 (N4600, N4581, N4263);
xor XOR2 (N4601, N4599, N2568);
nor NOR4 (N4602, N4589, N1450, N4071, N3429);
nor NOR2 (N4603, N4593, N2884);
or OR3 (N4604, N4597, N1656, N4567);
not NOT1 (N4605, N4604);
xor XOR2 (N4606, N4600, N1850);
xor XOR2 (N4607, N4596, N1900);
and AND4 (N4608, N4601, N1547, N2679, N119);
buf BUF1 (N4609, N4606);
xor XOR2 (N4610, N4602, N3366);
and AND3 (N4611, N4598, N1602, N2356);
buf BUF1 (N4612, N4611);
nor NOR4 (N4613, N4590, N539, N2804, N2662);
nand NAND2 (N4614, N4605, N2659);
nand NAND2 (N4615, N4612, N226);
or OR4 (N4616, N4610, N2536, N906, N50);
or OR4 (N4617, N4595, N2297, N3874, N2856);
and AND3 (N4618, N4614, N3440, N610);
or OR4 (N4619, N4609, N4060, N1448, N25);
nor NOR3 (N4620, N4617, N3300, N2673);
nor NOR3 (N4621, N4607, N388, N3969);
or OR3 (N4622, N4619, N2736, N1051);
nand NAND3 (N4623, N4608, N1818, N3567);
buf BUF1 (N4624, N4615);
nor NOR2 (N4625, N4620, N3810);
nand NAND2 (N4626, N4623, N4521);
not NOT1 (N4627, N4621);
and AND4 (N4628, N4613, N2504, N2856, N3442);
buf BUF1 (N4629, N4625);
nand NAND2 (N4630, N4622, N2808);
nand NAND4 (N4631, N4588, N3686, N1008, N116);
not NOT1 (N4632, N4618);
nor NOR4 (N4633, N4630, N867, N4469, N3581);
or OR4 (N4634, N4631, N1015, N2663, N3381);
buf BUF1 (N4635, N4632);
xor XOR2 (N4636, N4603, N1425);
or OR2 (N4637, N4626, N4619);
not NOT1 (N4638, N4637);
and AND3 (N4639, N4635, N1084, N2113);
nand NAND4 (N4640, N4634, N2671, N3306, N2172);
buf BUF1 (N4641, N4633);
and AND3 (N4642, N4636, N3863, N410);
xor XOR2 (N4643, N4640, N4396);
and AND3 (N4644, N4639, N673, N176);
or OR2 (N4645, N4616, N381);
xor XOR2 (N4646, N4643, N3966);
and AND3 (N4647, N4629, N844, N2116);
xor XOR2 (N4648, N4642, N2877);
not NOT1 (N4649, N4648);
xor XOR2 (N4650, N4628, N201);
not NOT1 (N4651, N4645);
not NOT1 (N4652, N4644);
or OR3 (N4653, N4624, N3471, N639);
xor XOR2 (N4654, N4651, N1765);
nor NOR3 (N4655, N4654, N358, N1956);
not NOT1 (N4656, N4652);
not NOT1 (N4657, N4650);
not NOT1 (N4658, N4649);
buf BUF1 (N4659, N4627);
nor NOR3 (N4660, N4646, N3447, N670);
not NOT1 (N4661, N4657);
buf BUF1 (N4662, N4655);
and AND3 (N4663, N4661, N4534, N3085);
nor NOR4 (N4664, N4638, N2325, N2036, N274);
nor NOR3 (N4665, N4647, N1199, N1983);
nor NOR3 (N4666, N4658, N2085, N2814);
buf BUF1 (N4667, N4663);
or OR4 (N4668, N4653, N4578, N4193, N2398);
not NOT1 (N4669, N4664);
not NOT1 (N4670, N4669);
not NOT1 (N4671, N4662);
and AND2 (N4672, N4659, N3108);
xor XOR2 (N4673, N4666, N3967);
xor XOR2 (N4674, N4670, N2228);
nand NAND3 (N4675, N4641, N2538, N3941);
not NOT1 (N4676, N4660);
buf BUF1 (N4677, N4665);
buf BUF1 (N4678, N4675);
or OR3 (N4679, N4677, N278, N4255);
or OR3 (N4680, N4656, N18, N4277);
not NOT1 (N4681, N4672);
and AND2 (N4682, N4674, N3625);
xor XOR2 (N4683, N4676, N1342);
xor XOR2 (N4684, N4668, N4293);
buf BUF1 (N4685, N4682);
xor XOR2 (N4686, N4684, N3367);
nand NAND3 (N4687, N4681, N1017, N460);
or OR3 (N4688, N4667, N3140, N1189);
nor NOR3 (N4689, N4685, N2216, N2677);
xor XOR2 (N4690, N4673, N3157);
not NOT1 (N4691, N4688);
or OR4 (N4692, N4680, N2217, N3455, N1663);
and AND4 (N4693, N4686, N2348, N227, N2412);
buf BUF1 (N4694, N4691);
not NOT1 (N4695, N4689);
or OR3 (N4696, N4678, N1636, N2172);
buf BUF1 (N4697, N4696);
nand NAND4 (N4698, N4694, N991, N3496, N2000);
buf BUF1 (N4699, N4692);
buf BUF1 (N4700, N4683);
nand NAND4 (N4701, N4690, N2977, N1714, N2758);
nor NOR4 (N4702, N4695, N512, N1826, N701);
and AND2 (N4703, N4693, N370);
xor XOR2 (N4704, N4671, N1139);
not NOT1 (N4705, N4697);
nand NAND3 (N4706, N4702, N4465, N222);
not NOT1 (N4707, N4704);
and AND4 (N4708, N4700, N1984, N112, N3743);
nor NOR2 (N4709, N4698, N4422);
nor NOR3 (N4710, N4705, N3026, N4406);
and AND3 (N4711, N4709, N4084, N733);
nand NAND2 (N4712, N4710, N1176);
not NOT1 (N4713, N4701);
not NOT1 (N4714, N4713);
nor NOR2 (N4715, N4699, N3488);
xor XOR2 (N4716, N4711, N4326);
buf BUF1 (N4717, N4712);
and AND3 (N4718, N4687, N4144, N4222);
not NOT1 (N4719, N4679);
nand NAND2 (N4720, N4717, N2825);
or OR3 (N4721, N4719, N2215, N3969);
xor XOR2 (N4722, N4708, N3417);
and AND2 (N4723, N4714, N1676);
not NOT1 (N4724, N4716);
nand NAND3 (N4725, N4706, N4570, N702);
not NOT1 (N4726, N4715);
not NOT1 (N4727, N4718);
not NOT1 (N4728, N4703);
buf BUF1 (N4729, N4728);
and AND4 (N4730, N4721, N139, N1847, N1232);
nor NOR2 (N4731, N4722, N703);
nand NAND4 (N4732, N4724, N2844, N4229, N1451);
and AND3 (N4733, N4732, N2966, N3417);
buf BUF1 (N4734, N4729);
and AND3 (N4735, N4723, N605, N519);
nand NAND3 (N4736, N4725, N2611, N4287);
buf BUF1 (N4737, N4733);
or OR2 (N4738, N4726, N3232);
not NOT1 (N4739, N4707);
not NOT1 (N4740, N4736);
nor NOR3 (N4741, N4730, N2878, N926);
and AND4 (N4742, N4739, N4189, N2770, N4511);
and AND3 (N4743, N4742, N1928, N1446);
not NOT1 (N4744, N4738);
xor XOR2 (N4745, N4731, N2363);
nor NOR4 (N4746, N4743, N4098, N3915, N1117);
and AND3 (N4747, N4746, N3460, N2402);
nand NAND3 (N4748, N4734, N786, N3900);
nor NOR3 (N4749, N4745, N3098, N2289);
nand NAND4 (N4750, N4744, N4415, N1495, N222);
not NOT1 (N4751, N4749);
xor XOR2 (N4752, N4751, N1519);
nand NAND3 (N4753, N4737, N831, N2742);
nor NOR4 (N4754, N4752, N4563, N610, N4477);
not NOT1 (N4755, N4740);
nand NAND3 (N4756, N4741, N2441, N1043);
and AND3 (N4757, N4747, N418, N4274);
and AND3 (N4758, N4727, N2618, N3625);
nor NOR3 (N4759, N4754, N1475, N676);
or OR4 (N4760, N4720, N2330, N2525, N2885);
or OR3 (N4761, N4760, N4346, N3941);
nand NAND4 (N4762, N4748, N3020, N2622, N3242);
buf BUF1 (N4763, N4755);
and AND2 (N4764, N4758, N2679);
nand NAND3 (N4765, N4756, N2460, N4099);
not NOT1 (N4766, N4750);
or OR3 (N4767, N4757, N4449, N830);
buf BUF1 (N4768, N4767);
or OR3 (N4769, N4766, N2539, N2536);
xor XOR2 (N4770, N4765, N2560);
and AND4 (N4771, N4769, N1318, N224, N1202);
nand NAND2 (N4772, N4753, N4645);
and AND4 (N4773, N4762, N2307, N2579, N38);
and AND3 (N4774, N4771, N4355, N313);
nand NAND3 (N4775, N4772, N2865, N2661);
nand NAND3 (N4776, N4768, N3783, N670);
and AND4 (N4777, N4770, N1364, N4580, N1606);
nor NOR4 (N4778, N4735, N1101, N3170, N3158);
buf BUF1 (N4779, N4774);
not NOT1 (N4780, N4775);
buf BUF1 (N4781, N4777);
xor XOR2 (N4782, N4759, N188);
nand NAND2 (N4783, N4780, N870);
buf BUF1 (N4784, N4783);
buf BUF1 (N4785, N4776);
or OR4 (N4786, N4779, N1727, N2862, N2512);
buf BUF1 (N4787, N4778);
or OR3 (N4788, N4787, N2124, N291);
nand NAND2 (N4789, N4764, N4121);
xor XOR2 (N4790, N4788, N3775);
buf BUF1 (N4791, N4773);
and AND2 (N4792, N4784, N307);
buf BUF1 (N4793, N4782);
or OR4 (N4794, N4790, N1055, N3976, N2797);
xor XOR2 (N4795, N4761, N652);
not NOT1 (N4796, N4763);
not NOT1 (N4797, N4789);
buf BUF1 (N4798, N4795);
nor NOR4 (N4799, N4797, N3741, N260, N3758);
xor XOR2 (N4800, N4798, N4356);
and AND3 (N4801, N4800, N2451, N3488);
and AND4 (N4802, N4793, N2544, N4478, N145);
nor NOR2 (N4803, N4802, N3312);
or OR4 (N4804, N4801, N949, N1796, N4501);
nand NAND2 (N4805, N4792, N1084);
or OR4 (N4806, N4781, N4288, N956, N4415);
or OR4 (N4807, N4791, N2567, N4572, N2875);
buf BUF1 (N4808, N4803);
not NOT1 (N4809, N4785);
and AND3 (N4810, N4808, N2866, N3406);
nand NAND4 (N4811, N4804, N2133, N2517, N2905);
nand NAND3 (N4812, N4786, N1598, N1484);
xor XOR2 (N4813, N4796, N1741);
buf BUF1 (N4814, N4807);
not NOT1 (N4815, N4812);
not NOT1 (N4816, N4813);
buf BUF1 (N4817, N4816);
nand NAND4 (N4818, N4814, N4121, N2870, N3298);
not NOT1 (N4819, N4818);
not NOT1 (N4820, N4815);
or OR4 (N4821, N4809, N3151, N1118, N3516);
or OR4 (N4822, N4819, N812, N2235, N660);
nor NOR2 (N4823, N4794, N2046);
buf BUF1 (N4824, N4823);
nand NAND3 (N4825, N4799, N2328, N2056);
not NOT1 (N4826, N4822);
nand NAND4 (N4827, N4820, N1111, N4359, N1294);
buf BUF1 (N4828, N4821);
buf BUF1 (N4829, N4824);
buf BUF1 (N4830, N4817);
xor XOR2 (N4831, N4805, N1841);
not NOT1 (N4832, N4825);
nor NOR2 (N4833, N4810, N3818);
not NOT1 (N4834, N4830);
nand NAND3 (N4835, N4832, N2043, N68);
not NOT1 (N4836, N4834);
nand NAND2 (N4837, N4833, N2344);
and AND3 (N4838, N4831, N2815, N3959);
nor NOR3 (N4839, N4837, N3461, N3362);
and AND4 (N4840, N4811, N340, N2058, N1167);
nand NAND2 (N4841, N4838, N275);
buf BUF1 (N4842, N4826);
or OR2 (N4843, N4840, N1708);
nand NAND2 (N4844, N4843, N2238);
not NOT1 (N4845, N4827);
xor XOR2 (N4846, N4842, N1193);
and AND2 (N4847, N4835, N4614);
buf BUF1 (N4848, N4828);
xor XOR2 (N4849, N4846, N1182);
and AND2 (N4850, N4806, N2817);
buf BUF1 (N4851, N4841);
xor XOR2 (N4852, N4847, N1868);
not NOT1 (N4853, N4829);
not NOT1 (N4854, N4839);
or OR4 (N4855, N4845, N3818, N3737, N2566);
not NOT1 (N4856, N4844);
nand NAND2 (N4857, N4836, N4812);
buf BUF1 (N4858, N4855);
nor NOR2 (N4859, N4853, N738);
xor XOR2 (N4860, N4850, N4006);
xor XOR2 (N4861, N4848, N4633);
nand NAND4 (N4862, N4849, N1227, N1960, N2753);
buf BUF1 (N4863, N4851);
or OR4 (N4864, N4857, N884, N413, N4693);
nand NAND3 (N4865, N4863, N1208, N1001);
nand NAND4 (N4866, N4861, N3656, N1083, N3518);
not NOT1 (N4867, N4856);
nand NAND4 (N4868, N4854, N1640, N3441, N3640);
xor XOR2 (N4869, N4859, N3399);
and AND3 (N4870, N4858, N2434, N1194);
nand NAND2 (N4871, N4852, N2860);
not NOT1 (N4872, N4865);
buf BUF1 (N4873, N4866);
nand NAND3 (N4874, N4872, N3912, N604);
buf BUF1 (N4875, N4864);
xor XOR2 (N4876, N4873, N4166);
nand NAND2 (N4877, N4871, N1717);
xor XOR2 (N4878, N4874, N2426);
buf BUF1 (N4879, N4860);
and AND4 (N4880, N4868, N1849, N3986, N101);
nor NOR2 (N4881, N4879, N304);
buf BUF1 (N4882, N4877);
xor XOR2 (N4883, N4869, N3517);
nor NOR4 (N4884, N4867, N1385, N2025, N3722);
and AND3 (N4885, N4883, N4531, N3947);
nand NAND2 (N4886, N4885, N4241);
buf BUF1 (N4887, N4882);
not NOT1 (N4888, N4884);
nand NAND4 (N4889, N4881, N4664, N967, N1318);
or OR2 (N4890, N4880, N3588);
buf BUF1 (N4891, N4876);
not NOT1 (N4892, N4887);
nor NOR3 (N4893, N4878, N844, N2606);
buf BUF1 (N4894, N4888);
and AND3 (N4895, N4889, N591, N3332);
not NOT1 (N4896, N4893);
buf BUF1 (N4897, N4891);
or OR3 (N4898, N4892, N4284, N1862);
or OR3 (N4899, N4896, N3165, N2345);
xor XOR2 (N4900, N4894, N1299);
nand NAND3 (N4901, N4900, N3454, N1175);
xor XOR2 (N4902, N4901, N3790);
nand NAND4 (N4903, N4895, N2794, N1391, N698);
and AND2 (N4904, N4875, N3628);
buf BUF1 (N4905, N4902);
buf BUF1 (N4906, N4886);
not NOT1 (N4907, N4898);
or OR2 (N4908, N4897, N2677);
buf BUF1 (N4909, N4907);
nand NAND2 (N4910, N4905, N4141);
nor NOR4 (N4911, N4910, N3380, N4509, N1776);
and AND4 (N4912, N4911, N1646, N4383, N1586);
and AND2 (N4913, N4909, N3622);
nor NOR4 (N4914, N4904, N2315, N1531, N3992);
or OR3 (N4915, N4870, N732, N886);
and AND2 (N4916, N4890, N2283);
nand NAND2 (N4917, N4912, N1287);
and AND3 (N4918, N4908, N4285, N489);
not NOT1 (N4919, N4915);
not NOT1 (N4920, N4903);
buf BUF1 (N4921, N4917);
and AND2 (N4922, N4916, N4241);
xor XOR2 (N4923, N4918, N4067);
buf BUF1 (N4924, N4921);
nor NOR2 (N4925, N4906, N3149);
xor XOR2 (N4926, N4913, N2659);
xor XOR2 (N4927, N4923, N3655);
nor NOR4 (N4928, N4862, N143, N4875, N4823);
buf BUF1 (N4929, N4919);
nor NOR2 (N4930, N4922, N1541);
xor XOR2 (N4931, N4920, N2781);
xor XOR2 (N4932, N4926, N2389);
nor NOR2 (N4933, N4925, N3036);
not NOT1 (N4934, N4929);
xor XOR2 (N4935, N4914, N3120);
not NOT1 (N4936, N4930);
not NOT1 (N4937, N4933);
nand NAND2 (N4938, N4936, N1248);
and AND2 (N4939, N4931, N3179);
xor XOR2 (N4940, N4927, N2715);
and AND3 (N4941, N4940, N477, N4865);
buf BUF1 (N4942, N4938);
and AND3 (N4943, N4924, N2668, N4356);
not NOT1 (N4944, N4935);
xor XOR2 (N4945, N4937, N3851);
or OR2 (N4946, N4939, N3616);
and AND3 (N4947, N4945, N4881, N470);
buf BUF1 (N4948, N4947);
or OR3 (N4949, N4934, N1206, N590);
nand NAND2 (N4950, N4944, N3484);
nand NAND2 (N4951, N4941, N612);
nor NOR2 (N4952, N4948, N1966);
or OR4 (N4953, N4899, N420, N3960, N2672);
or OR2 (N4954, N4953, N2029);
xor XOR2 (N4955, N4946, N3046);
nand NAND4 (N4956, N4932, N3490, N512, N1631);
or OR3 (N4957, N4942, N3481, N1412);
not NOT1 (N4958, N4949);
nand NAND4 (N4959, N4952, N1159, N4245, N367);
and AND2 (N4960, N4956, N2721);
and AND3 (N4961, N4955, N622, N79);
xor XOR2 (N4962, N4960, N1106);
or OR4 (N4963, N4951, N4407, N2009, N289);
buf BUF1 (N4964, N4963);
not NOT1 (N4965, N4964);
nor NOR4 (N4966, N4959, N1876, N2777, N4492);
nand NAND3 (N4967, N4957, N2106, N4632);
nor NOR4 (N4968, N4954, N1069, N2579, N4264);
nor NOR4 (N4969, N4950, N931, N3369, N2194);
and AND2 (N4970, N4962, N3465);
buf BUF1 (N4971, N4965);
nor NOR3 (N4972, N4961, N3158, N1023);
xor XOR2 (N4973, N4966, N677);
and AND2 (N4974, N4972, N1539);
and AND3 (N4975, N4943, N2062, N571);
xor XOR2 (N4976, N4969, N695);
nand NAND3 (N4977, N4968, N3067, N1552);
not NOT1 (N4978, N4973);
buf BUF1 (N4979, N4975);
xor XOR2 (N4980, N4976, N1163);
or OR3 (N4981, N4971, N889, N3473);
xor XOR2 (N4982, N4958, N4941);
buf BUF1 (N4983, N4981);
nand NAND3 (N4984, N4970, N4431, N3349);
nor NOR4 (N4985, N4979, N3875, N4498, N3609);
nand NAND4 (N4986, N4984, N4571, N2708, N3561);
nand NAND4 (N4987, N4977, N2856, N91, N191);
nor NOR3 (N4988, N4982, N4869, N3780);
nor NOR4 (N4989, N4983, N1941, N4132, N3290);
nor NOR2 (N4990, N4928, N1678);
xor XOR2 (N4991, N4990, N3993);
nor NOR4 (N4992, N4974, N3649, N4058, N2076);
xor XOR2 (N4993, N4980, N1336);
nor NOR3 (N4994, N4987, N1637, N2050);
nand NAND2 (N4995, N4986, N3518);
or OR2 (N4996, N4967, N4279);
or OR2 (N4997, N4978, N2661);
xor XOR2 (N4998, N4996, N4252);
and AND4 (N4999, N4992, N4208, N785, N2382);
and AND2 (N5000, N4993, N3205);
not NOT1 (N5001, N4997);
xor XOR2 (N5002, N4985, N369);
and AND4 (N5003, N4988, N1210, N4233, N3437);
and AND3 (N5004, N5003, N616, N1525);
xor XOR2 (N5005, N4994, N2110);
xor XOR2 (N5006, N4998, N1236);
nor NOR3 (N5007, N5000, N4681, N2867);
xor XOR2 (N5008, N5004, N4128);
nor NOR4 (N5009, N5002, N1459, N1043, N3621);
xor XOR2 (N5010, N5008, N4958);
not NOT1 (N5011, N4995);
xor XOR2 (N5012, N5001, N781);
buf BUF1 (N5013, N5010);
nor NOR3 (N5014, N5012, N4353, N142);
xor XOR2 (N5015, N4999, N1383);
nand NAND3 (N5016, N5013, N4175, N3140);
xor XOR2 (N5017, N5015, N180);
buf BUF1 (N5018, N5014);
or OR3 (N5019, N5007, N3857, N222);
not NOT1 (N5020, N5005);
nand NAND2 (N5021, N4989, N2863);
not NOT1 (N5022, N5006);
nor NOR3 (N5023, N5020, N1542, N3354);
buf BUF1 (N5024, N5016);
nor NOR2 (N5025, N4991, N1237);
nor NOR4 (N5026, N5024, N692, N4458, N1139);
nand NAND3 (N5027, N5011, N3911, N111);
not NOT1 (N5028, N5025);
xor XOR2 (N5029, N5021, N2159);
buf BUF1 (N5030, N5017);
or OR4 (N5031, N5019, N3532, N2787, N2383);
nor NOR3 (N5032, N5009, N1458, N4497);
or OR2 (N5033, N5031, N2820);
buf BUF1 (N5034, N5018);
xor XOR2 (N5035, N5029, N672);
nand NAND2 (N5036, N5030, N2122);
or OR2 (N5037, N5023, N3229);
and AND3 (N5038, N5026, N3820, N448);
buf BUF1 (N5039, N5028);
xor XOR2 (N5040, N5034, N4359);
nor NOR4 (N5041, N5036, N117, N834, N418);
buf BUF1 (N5042, N5027);
not NOT1 (N5043, N5039);
xor XOR2 (N5044, N5040, N241);
and AND2 (N5045, N5033, N3770);
or OR3 (N5046, N5042, N2781, N3866);
buf BUF1 (N5047, N5038);
buf BUF1 (N5048, N5035);
buf BUF1 (N5049, N5044);
buf BUF1 (N5050, N5037);
nor NOR3 (N5051, N5032, N869, N4543);
or OR3 (N5052, N5051, N3916, N276);
and AND4 (N5053, N5047, N2071, N1387, N2556);
not NOT1 (N5054, N5043);
not NOT1 (N5055, N5050);
and AND3 (N5056, N5052, N4484, N3603);
or OR4 (N5057, N5022, N708, N3760, N1453);
xor XOR2 (N5058, N5053, N4967);
nor NOR4 (N5059, N5046, N3715, N2771, N3385);
xor XOR2 (N5060, N5048, N3806);
not NOT1 (N5061, N5059);
and AND3 (N5062, N5058, N4968, N3747);
or OR3 (N5063, N5049, N620, N4878);
nor NOR3 (N5064, N5057, N4948, N1920);
buf BUF1 (N5065, N5041);
and AND3 (N5066, N5065, N3352, N4632);
and AND2 (N5067, N5063, N1343);
or OR2 (N5068, N5064, N4366);
buf BUF1 (N5069, N5060);
not NOT1 (N5070, N5045);
or OR2 (N5071, N5067, N410);
and AND3 (N5072, N5062, N2374, N1618);
xor XOR2 (N5073, N5072, N2265);
and AND4 (N5074, N5056, N428, N614, N2593);
and AND4 (N5075, N5066, N4189, N4903, N3284);
not NOT1 (N5076, N5061);
not NOT1 (N5077, N5055);
or OR4 (N5078, N5070, N2196, N4050, N1386);
not NOT1 (N5079, N5069);
nor NOR3 (N5080, N5071, N3728, N4164);
and AND4 (N5081, N5076, N4844, N2436, N2691);
nand NAND3 (N5082, N5081, N4779, N424);
nor NOR3 (N5083, N5078, N2769, N63);
nor NOR3 (N5084, N5068, N122, N2544);
xor XOR2 (N5085, N5075, N3610);
and AND2 (N5086, N5074, N3096);
xor XOR2 (N5087, N5079, N4399);
and AND4 (N5088, N5087, N2757, N37, N429);
or OR3 (N5089, N5080, N2970, N3513);
nand NAND4 (N5090, N5089, N1509, N4284, N1808);
xor XOR2 (N5091, N5088, N623);
buf BUF1 (N5092, N5090);
or OR4 (N5093, N5077, N496, N4070, N1922);
and AND2 (N5094, N5082, N3120);
buf BUF1 (N5095, N5086);
nor NOR2 (N5096, N5094, N1586);
not NOT1 (N5097, N5095);
not NOT1 (N5098, N5092);
nand NAND2 (N5099, N5073, N3466);
buf BUF1 (N5100, N5084);
nor NOR3 (N5101, N5083, N2025, N2783);
and AND3 (N5102, N5054, N3239, N4971);
and AND3 (N5103, N5091, N4131, N4262);
xor XOR2 (N5104, N5085, N3558);
not NOT1 (N5105, N5103);
or OR3 (N5106, N5102, N1672, N4230);
or OR4 (N5107, N5098, N3602, N1465, N4727);
xor XOR2 (N5108, N5096, N2191);
or OR4 (N5109, N5099, N3846, N135, N2296);
nand NAND2 (N5110, N5100, N4567);
not NOT1 (N5111, N5101);
nand NAND2 (N5112, N5111, N1759);
xor XOR2 (N5113, N5109, N299);
and AND3 (N5114, N5097, N4589, N448);
or OR4 (N5115, N5106, N2592, N2918, N1397);
and AND2 (N5116, N5112, N666);
not NOT1 (N5117, N5113);
xor XOR2 (N5118, N5117, N1280);
or OR2 (N5119, N5114, N2860);
not NOT1 (N5120, N5118);
and AND4 (N5121, N5104, N1723, N1216, N4650);
nand NAND3 (N5122, N5107, N1059, N3422);
buf BUF1 (N5123, N5115);
xor XOR2 (N5124, N5105, N4414);
buf BUF1 (N5125, N5124);
or OR4 (N5126, N5123, N2026, N2741, N2413);
nand NAND3 (N5127, N5126, N3746, N3977);
and AND3 (N5128, N5122, N2293, N2210);
xor XOR2 (N5129, N5116, N3149);
nor NOR2 (N5130, N5119, N3804);
or OR2 (N5131, N5128, N2189);
or OR2 (N5132, N5120, N3243);
xor XOR2 (N5133, N5131, N1358);
or OR4 (N5134, N5108, N3171, N1040, N458);
not NOT1 (N5135, N5129);
nand NAND4 (N5136, N5134, N3328, N1088, N157);
buf BUF1 (N5137, N5132);
or OR2 (N5138, N5125, N1738);
xor XOR2 (N5139, N5130, N2964);
and AND2 (N5140, N5133, N4508);
nor NOR3 (N5141, N5135, N2829, N991);
nor NOR2 (N5142, N5136, N1282);
or OR4 (N5143, N5121, N1800, N4575, N2426);
xor XOR2 (N5144, N5139, N3109);
buf BUF1 (N5145, N5137);
xor XOR2 (N5146, N5140, N3044);
xor XOR2 (N5147, N5141, N204);
xor XOR2 (N5148, N5142, N2502);
xor XOR2 (N5149, N5147, N4152);
or OR2 (N5150, N5110, N560);
buf BUF1 (N5151, N5143);
xor XOR2 (N5152, N5138, N3216);
nand NAND2 (N5153, N5145, N1219);
nand NAND2 (N5154, N5151, N2593);
nand NAND2 (N5155, N5148, N617);
buf BUF1 (N5156, N5150);
nand NAND2 (N5157, N5144, N4715);
not NOT1 (N5158, N5154);
not NOT1 (N5159, N5158);
nor NOR3 (N5160, N5152, N4834, N2846);
buf BUF1 (N5161, N5153);
xor XOR2 (N5162, N5160, N2980);
not NOT1 (N5163, N5156);
not NOT1 (N5164, N5155);
nand NAND2 (N5165, N5127, N5141);
buf BUF1 (N5166, N5159);
xor XOR2 (N5167, N5093, N2714);
xor XOR2 (N5168, N5166, N4040);
nor NOR4 (N5169, N5164, N2027, N4714, N2383);
buf BUF1 (N5170, N5162);
and AND4 (N5171, N5165, N3399, N3402, N911);
and AND2 (N5172, N5163, N165);
nand NAND3 (N5173, N5171, N4868, N4702);
buf BUF1 (N5174, N5167);
nor NOR4 (N5175, N5149, N3065, N5064, N4459);
buf BUF1 (N5176, N5161);
xor XOR2 (N5177, N5168, N2516);
nor NOR4 (N5178, N5176, N1179, N448, N4621);
or OR3 (N5179, N5178, N1416, N2440);
nor NOR3 (N5180, N5175, N1362, N3224);
not NOT1 (N5181, N5180);
xor XOR2 (N5182, N5173, N4732);
not NOT1 (N5183, N5174);
buf BUF1 (N5184, N5181);
nand NAND2 (N5185, N5169, N3930);
nand NAND3 (N5186, N5157, N1634, N2019);
xor XOR2 (N5187, N5186, N1817);
xor XOR2 (N5188, N5146, N1041);
buf BUF1 (N5189, N5177);
nor NOR2 (N5190, N5185, N3115);
nand NAND4 (N5191, N5182, N3960, N383, N2015);
buf BUF1 (N5192, N5187);
not NOT1 (N5193, N5188);
xor XOR2 (N5194, N5183, N3016);
or OR3 (N5195, N5192, N2708, N2198);
buf BUF1 (N5196, N5170);
buf BUF1 (N5197, N5184);
or OR2 (N5198, N5172, N4836);
and AND2 (N5199, N5198, N3028);
or OR3 (N5200, N5189, N3077, N86);
or OR4 (N5201, N5190, N1095, N562, N28);
or OR3 (N5202, N5194, N3554, N2826);
and AND2 (N5203, N5179, N5163);
xor XOR2 (N5204, N5201, N2288);
or OR2 (N5205, N5204, N3501);
and AND2 (N5206, N5203, N1016);
nand NAND2 (N5207, N5199, N3633);
buf BUF1 (N5208, N5207);
nor NOR3 (N5209, N5202, N149, N1941);
or OR4 (N5210, N5193, N4863, N4856, N5068);
nand NAND4 (N5211, N5206, N5196, N4431, N3516);
buf BUF1 (N5212, N672);
not NOT1 (N5213, N5208);
buf BUF1 (N5214, N5213);
nand NAND2 (N5215, N5214, N157);
buf BUF1 (N5216, N5197);
and AND3 (N5217, N5195, N74, N5119);
or OR3 (N5218, N5216, N579, N1747);
xor XOR2 (N5219, N5205, N4202);
and AND3 (N5220, N5212, N1872, N4575);
and AND2 (N5221, N5191, N2030);
xor XOR2 (N5222, N5217, N4756);
and AND3 (N5223, N5210, N677, N2608);
nand NAND4 (N5224, N5209, N708, N1767, N2422);
xor XOR2 (N5225, N5222, N2808);
xor XOR2 (N5226, N5218, N2340);
xor XOR2 (N5227, N5223, N69);
nor NOR4 (N5228, N5221, N2228, N3074, N1185);
not NOT1 (N5229, N5227);
buf BUF1 (N5230, N5225);
or OR2 (N5231, N5230, N4100);
buf BUF1 (N5232, N5215);
nor NOR2 (N5233, N5219, N2404);
or OR4 (N5234, N5200, N4213, N1705, N3158);
xor XOR2 (N5235, N5233, N3140);
not NOT1 (N5236, N5226);
not NOT1 (N5237, N5228);
nor NOR3 (N5238, N5237, N4435, N4172);
buf BUF1 (N5239, N5231);
xor XOR2 (N5240, N5211, N90);
and AND4 (N5241, N5236, N3326, N459, N3949);
buf BUF1 (N5242, N5229);
or OR4 (N5243, N5240, N2295, N1558, N4147);
nand NAND2 (N5244, N5235, N1297);
not NOT1 (N5245, N5242);
xor XOR2 (N5246, N5244, N2270);
buf BUF1 (N5247, N5224);
or OR3 (N5248, N5239, N3852, N1762);
not NOT1 (N5249, N5245);
and AND3 (N5250, N5238, N5224, N1838);
not NOT1 (N5251, N5249);
buf BUF1 (N5252, N5234);
not NOT1 (N5253, N5247);
and AND2 (N5254, N5252, N2632);
nor NOR3 (N5255, N5254, N61, N183);
and AND3 (N5256, N5251, N4396, N1545);
buf BUF1 (N5257, N5253);
or OR4 (N5258, N5246, N2447, N792, N1597);
not NOT1 (N5259, N5220);
nand NAND3 (N5260, N5243, N5088, N3606);
buf BUF1 (N5261, N5259);
not NOT1 (N5262, N5241);
not NOT1 (N5263, N5258);
buf BUF1 (N5264, N5263);
nor NOR4 (N5265, N5262, N2546, N2351, N5171);
or OR2 (N5266, N5248, N1210);
buf BUF1 (N5267, N5266);
nor NOR3 (N5268, N5267, N2015, N4906);
and AND4 (N5269, N5232, N4835, N3768, N2420);
not NOT1 (N5270, N5264);
or OR2 (N5271, N5257, N4091);
nand NAND3 (N5272, N5250, N1935, N2834);
nor NOR3 (N5273, N5272, N1918, N1573);
and AND4 (N5274, N5265, N1888, N2148, N1644);
buf BUF1 (N5275, N5270);
xor XOR2 (N5276, N5274, N3437);
nor NOR2 (N5277, N5269, N1509);
buf BUF1 (N5278, N5273);
and AND4 (N5279, N5276, N119, N5054, N89);
and AND4 (N5280, N5278, N2281, N745, N4103);
nor NOR2 (N5281, N5256, N4005);
not NOT1 (N5282, N5271);
nand NAND4 (N5283, N5277, N2966, N2514, N3723);
or OR4 (N5284, N5280, N3915, N924, N731);
buf BUF1 (N5285, N5275);
nor NOR4 (N5286, N5282, N737, N4714, N5141);
or OR2 (N5287, N5279, N1668);
or OR2 (N5288, N5287, N428);
not NOT1 (N5289, N5285);
nor NOR2 (N5290, N5261, N3589);
nand NAND4 (N5291, N5281, N1091, N988, N1854);
and AND3 (N5292, N5284, N5045, N4662);
nor NOR3 (N5293, N5290, N2634, N1772);
buf BUF1 (N5294, N5283);
and AND2 (N5295, N5268, N4435);
not NOT1 (N5296, N5295);
and AND4 (N5297, N5291, N1044, N967, N84);
buf BUF1 (N5298, N5288);
nor NOR3 (N5299, N5298, N4591, N349);
nor NOR4 (N5300, N5292, N4559, N167, N3390);
nor NOR4 (N5301, N5300, N3118, N2419, N5253);
or OR3 (N5302, N5286, N4989, N1314);
not NOT1 (N5303, N5294);
xor XOR2 (N5304, N5296, N1548);
xor XOR2 (N5305, N5301, N3408);
xor XOR2 (N5306, N5293, N427);
nor NOR2 (N5307, N5299, N2377);
or OR3 (N5308, N5307, N155, N1521);
not NOT1 (N5309, N5255);
and AND3 (N5310, N5309, N1867, N2513);
or OR3 (N5311, N5310, N902, N1465);
nor NOR4 (N5312, N5297, N3793, N557, N4912);
or OR4 (N5313, N5306, N1118, N2081, N748);
or OR4 (N5314, N5308, N1604, N3437, N2543);
not NOT1 (N5315, N5260);
xor XOR2 (N5316, N5313, N3131);
nor NOR3 (N5317, N5305, N1303, N1579);
and AND4 (N5318, N5316, N5066, N1168, N5276);
and AND4 (N5319, N5315, N1153, N460, N2548);
nand NAND2 (N5320, N5312, N5190);
nor NOR4 (N5321, N5289, N30, N3421, N2444);
nor NOR3 (N5322, N5302, N1046, N589);
not NOT1 (N5323, N5319);
or OR4 (N5324, N5320, N4220, N1357, N3069);
and AND2 (N5325, N5321, N2290);
or OR2 (N5326, N5304, N148);
buf BUF1 (N5327, N5323);
not NOT1 (N5328, N5324);
nand NAND2 (N5329, N5328, N1381);
nand NAND2 (N5330, N5314, N3010);
buf BUF1 (N5331, N5326);
nand NAND4 (N5332, N5325, N178, N2322, N2760);
nor NOR3 (N5333, N5311, N3474, N4964);
nor NOR2 (N5334, N5329, N585);
nand NAND4 (N5335, N5317, N3662, N2866, N1663);
xor XOR2 (N5336, N5335, N3932);
buf BUF1 (N5337, N5303);
and AND4 (N5338, N5336, N498, N2621, N2001);
not NOT1 (N5339, N5330);
nand NAND3 (N5340, N5332, N1765, N4373);
or OR3 (N5341, N5334, N5166, N3466);
not NOT1 (N5342, N5338);
buf BUF1 (N5343, N5341);
buf BUF1 (N5344, N5342);
buf BUF1 (N5345, N5327);
not NOT1 (N5346, N5331);
and AND2 (N5347, N5322, N920);
buf BUF1 (N5348, N5345);
nand NAND3 (N5349, N5343, N2346, N4690);
buf BUF1 (N5350, N5333);
not NOT1 (N5351, N5348);
nor NOR2 (N5352, N5347, N23);
not NOT1 (N5353, N5339);
not NOT1 (N5354, N5349);
not NOT1 (N5355, N5337);
nand NAND3 (N5356, N5355, N342, N259);
nand NAND4 (N5357, N5344, N1859, N2575, N79);
buf BUF1 (N5358, N5354);
buf BUF1 (N5359, N5340);
xor XOR2 (N5360, N5350, N2220);
and AND3 (N5361, N5351, N4055, N4440);
and AND2 (N5362, N5346, N4711);
buf BUF1 (N5363, N5356);
nor NOR2 (N5364, N5362, N4403);
buf BUF1 (N5365, N5363);
and AND3 (N5366, N5360, N3873, N4057);
nand NAND2 (N5367, N5361, N1156);
buf BUF1 (N5368, N5366);
or OR4 (N5369, N5357, N418, N169, N3269);
xor XOR2 (N5370, N5318, N468);
not NOT1 (N5371, N5353);
not NOT1 (N5372, N5364);
not NOT1 (N5373, N5352);
nand NAND2 (N5374, N5371, N3580);
xor XOR2 (N5375, N5374, N206);
or OR2 (N5376, N5370, N1070);
or OR4 (N5377, N5365, N3180, N4515, N4270);
xor XOR2 (N5378, N5376, N2355);
not NOT1 (N5379, N5372);
buf BUF1 (N5380, N5378);
not NOT1 (N5381, N5358);
or OR3 (N5382, N5368, N753, N5363);
buf BUF1 (N5383, N5373);
and AND2 (N5384, N5377, N287);
and AND2 (N5385, N5384, N627);
not NOT1 (N5386, N5381);
nand NAND3 (N5387, N5383, N3805, N4077);
buf BUF1 (N5388, N5386);
nand NAND3 (N5389, N5369, N3031, N1714);
xor XOR2 (N5390, N5359, N1028);
nor NOR2 (N5391, N5375, N320);
nor NOR3 (N5392, N5380, N2987, N3718);
buf BUF1 (N5393, N5389);
or OR2 (N5394, N5388, N1783);
nand NAND3 (N5395, N5379, N5282, N2486);
nand NAND3 (N5396, N5367, N1654, N4517);
nand NAND2 (N5397, N5385, N5017);
xor XOR2 (N5398, N5387, N3168);
and AND2 (N5399, N5394, N1224);
or OR2 (N5400, N5395, N2106);
or OR3 (N5401, N5399, N3998, N3174);
nand NAND2 (N5402, N5382, N2460);
nor NOR3 (N5403, N5396, N976, N3950);
buf BUF1 (N5404, N5401);
nand NAND3 (N5405, N5390, N4932, N948);
nor NOR3 (N5406, N5391, N2774, N3525);
xor XOR2 (N5407, N5403, N2322);
nor NOR4 (N5408, N5398, N1903, N3207, N3623);
buf BUF1 (N5409, N5408);
buf BUF1 (N5410, N5409);
and AND3 (N5411, N5405, N819, N2773);
xor XOR2 (N5412, N5410, N2219);
nand NAND2 (N5413, N5411, N4091);
xor XOR2 (N5414, N5397, N4725);
or OR3 (N5415, N5414, N2518, N3421);
not NOT1 (N5416, N5412);
and AND3 (N5417, N5404, N495, N2330);
nand NAND2 (N5418, N5416, N4578);
and AND3 (N5419, N5407, N655, N3754);
nor NOR4 (N5420, N5406, N2012, N5173, N1435);
or OR3 (N5421, N5400, N5245, N2348);
or OR4 (N5422, N5418, N2973, N855, N4524);
nand NAND2 (N5423, N5413, N4414);
or OR3 (N5424, N5421, N28, N2960);
and AND2 (N5425, N5417, N60);
buf BUF1 (N5426, N5422);
or OR4 (N5427, N5426, N1192, N1033, N4439);
nor NOR2 (N5428, N5425, N2588);
nor NOR2 (N5429, N5392, N3729);
nor NOR4 (N5430, N5420, N1899, N3310, N300);
buf BUF1 (N5431, N5393);
and AND3 (N5432, N5424, N2596, N4634);
or OR4 (N5433, N5429, N5081, N1588, N3720);
xor XOR2 (N5434, N5432, N1728);
nor NOR4 (N5435, N5423, N4776, N12, N3512);
nor NOR2 (N5436, N5433, N3082);
xor XOR2 (N5437, N5427, N383);
xor XOR2 (N5438, N5428, N3123);
and AND3 (N5439, N5438, N1030, N1557);
not NOT1 (N5440, N5430);
buf BUF1 (N5441, N5402);
or OR3 (N5442, N5441, N4786, N4027);
not NOT1 (N5443, N5442);
or OR2 (N5444, N5435, N608);
xor XOR2 (N5445, N5419, N4787);
buf BUF1 (N5446, N5443);
xor XOR2 (N5447, N5440, N2508);
nand NAND3 (N5448, N5447, N2099, N834);
nand NAND3 (N5449, N5445, N3167, N1087);
xor XOR2 (N5450, N5434, N419);
or OR2 (N5451, N5437, N3295);
nand NAND2 (N5452, N5439, N13);
and AND4 (N5453, N5449, N1140, N3883, N4964);
or OR2 (N5454, N5446, N4546);
not NOT1 (N5455, N5454);
xor XOR2 (N5456, N5431, N4390);
nor NOR3 (N5457, N5452, N306, N4320);
not NOT1 (N5458, N5453);
buf BUF1 (N5459, N5450);
buf BUF1 (N5460, N5455);
nor NOR2 (N5461, N5444, N1918);
or OR4 (N5462, N5461, N2452, N514, N3401);
nand NAND4 (N5463, N5451, N3064, N4506, N867);
buf BUF1 (N5464, N5415);
not NOT1 (N5465, N5463);
not NOT1 (N5466, N5464);
not NOT1 (N5467, N5456);
or OR2 (N5468, N5467, N2026);
nor NOR4 (N5469, N5462, N4987, N3173, N2980);
nand NAND3 (N5470, N5466, N3148, N3705);
or OR2 (N5471, N5465, N756);
nand NAND3 (N5472, N5470, N534, N620);
nor NOR3 (N5473, N5472, N4717, N688);
or OR2 (N5474, N5468, N1502);
not NOT1 (N5475, N5457);
nor NOR2 (N5476, N5471, N4534);
xor XOR2 (N5477, N5436, N4801);
xor XOR2 (N5478, N5476, N2584);
or OR4 (N5479, N5460, N4280, N298, N968);
xor XOR2 (N5480, N5473, N2734);
nor NOR3 (N5481, N5475, N1716, N3725);
and AND4 (N5482, N5459, N466, N3492, N2433);
nor NOR2 (N5483, N5480, N2235);
xor XOR2 (N5484, N5477, N1566);
not NOT1 (N5485, N5481);
xor XOR2 (N5486, N5479, N2854);
and AND4 (N5487, N5469, N2474, N4184, N3043);
nand NAND2 (N5488, N5483, N3681);
or OR3 (N5489, N5482, N569, N1565);
buf BUF1 (N5490, N5487);
buf BUF1 (N5491, N5478);
nor NOR3 (N5492, N5474, N4985, N887);
or OR3 (N5493, N5484, N613, N3859);
or OR3 (N5494, N5488, N4260, N2672);
xor XOR2 (N5495, N5493, N929);
or OR2 (N5496, N5485, N5125);
nor NOR2 (N5497, N5448, N3450);
or OR2 (N5498, N5486, N1810);
or OR2 (N5499, N5489, N4522);
xor XOR2 (N5500, N5458, N2829);
buf BUF1 (N5501, N5491);
and AND3 (N5502, N5499, N4987, N2533);
xor XOR2 (N5503, N5497, N3304);
buf BUF1 (N5504, N5494);
buf BUF1 (N5505, N5504);
and AND4 (N5506, N5502, N4282, N3187, N2630);
not NOT1 (N5507, N5495);
nand NAND3 (N5508, N5507, N3504, N3584);
buf BUF1 (N5509, N5508);
xor XOR2 (N5510, N5500, N3815);
nor NOR4 (N5511, N5509, N907, N827, N2928);
and AND4 (N5512, N5506, N5093, N82, N3910);
and AND2 (N5513, N5492, N1706);
xor XOR2 (N5514, N5498, N370);
and AND4 (N5515, N5511, N478, N2110, N3575);
or OR2 (N5516, N5503, N2501);
buf BUF1 (N5517, N5512);
nor NOR2 (N5518, N5514, N4069);
nor NOR2 (N5519, N5518, N1430);
xor XOR2 (N5520, N5496, N5249);
not NOT1 (N5521, N5515);
nand NAND2 (N5522, N5521, N914);
or OR2 (N5523, N5510, N1876);
not NOT1 (N5524, N5519);
xor XOR2 (N5525, N5523, N5220);
nor NOR3 (N5526, N5490, N5027, N1905);
and AND2 (N5527, N5513, N3639);
xor XOR2 (N5528, N5526, N1554);
or OR4 (N5529, N5528, N3973, N2320, N368);
buf BUF1 (N5530, N5505);
and AND3 (N5531, N5527, N878, N1953);
xor XOR2 (N5532, N5524, N1714);
nand NAND4 (N5533, N5529, N1331, N3628, N1105);
xor XOR2 (N5534, N5525, N5310);
xor XOR2 (N5535, N5522, N4424);
or OR2 (N5536, N5535, N2266);
not NOT1 (N5537, N5536);
not NOT1 (N5538, N5537);
not NOT1 (N5539, N5501);
not NOT1 (N5540, N5516);
nand NAND3 (N5541, N5533, N132, N770);
or OR3 (N5542, N5540, N661, N167);
xor XOR2 (N5543, N5531, N843);
not NOT1 (N5544, N5517);
xor XOR2 (N5545, N5520, N4958);
or OR2 (N5546, N5542, N2400);
and AND2 (N5547, N5539, N114);
xor XOR2 (N5548, N5546, N2150);
not NOT1 (N5549, N5541);
buf BUF1 (N5550, N5534);
xor XOR2 (N5551, N5550, N4729);
not NOT1 (N5552, N5545);
xor XOR2 (N5553, N5552, N4479);
nand NAND3 (N5554, N5532, N1203, N852);
and AND2 (N5555, N5530, N661);
nand NAND3 (N5556, N5543, N3842, N1760);
and AND3 (N5557, N5544, N5261, N4000);
not NOT1 (N5558, N5556);
nor NOR2 (N5559, N5558, N4476);
and AND2 (N5560, N5538, N1550);
and AND3 (N5561, N5553, N3134, N2732);
or OR4 (N5562, N5547, N2733, N5358, N5034);
not NOT1 (N5563, N5554);
nand NAND4 (N5564, N5549, N2831, N1969, N1273);
nor NOR2 (N5565, N5551, N1605);
xor XOR2 (N5566, N5565, N4024);
buf BUF1 (N5567, N5561);
or OR2 (N5568, N5566, N161);
or OR2 (N5569, N5568, N3140);
nand NAND4 (N5570, N5569, N842, N2296, N1684);
nor NOR2 (N5571, N5559, N5347);
and AND2 (N5572, N5562, N3380);
nor NOR4 (N5573, N5555, N1457, N4528, N622);
xor XOR2 (N5574, N5563, N4073);
not NOT1 (N5575, N5567);
nor NOR3 (N5576, N5564, N1586, N4251);
nor NOR2 (N5577, N5573, N4382);
and AND4 (N5578, N5577, N2032, N2303, N5508);
buf BUF1 (N5579, N5576);
not NOT1 (N5580, N5578);
or OR3 (N5581, N5560, N5372, N2134);
not NOT1 (N5582, N5579);
buf BUF1 (N5583, N5548);
xor XOR2 (N5584, N5575, N3162);
xor XOR2 (N5585, N5583, N1410);
or OR3 (N5586, N5584, N5162, N757);
buf BUF1 (N5587, N5582);
not NOT1 (N5588, N5572);
not NOT1 (N5589, N5571);
not NOT1 (N5590, N5574);
buf BUF1 (N5591, N5586);
buf BUF1 (N5592, N5587);
not NOT1 (N5593, N5590);
nand NAND4 (N5594, N5585, N5021, N2603, N3890);
xor XOR2 (N5595, N5591, N5587);
nand NAND2 (N5596, N5588, N3048);
nand NAND2 (N5597, N5596, N1147);
buf BUF1 (N5598, N5593);
buf BUF1 (N5599, N5581);
buf BUF1 (N5600, N5595);
nand NAND2 (N5601, N5589, N5588);
xor XOR2 (N5602, N5600, N632);
nor NOR4 (N5603, N5580, N387, N2728, N1716);
xor XOR2 (N5604, N5599, N1295);
and AND4 (N5605, N5592, N5546, N3645, N2089);
nand NAND2 (N5606, N5597, N1099);
nor NOR2 (N5607, N5605, N881);
nand NAND4 (N5608, N5598, N3422, N416, N5372);
or OR3 (N5609, N5557, N2665, N696);
buf BUF1 (N5610, N5608);
and AND2 (N5611, N5570, N3060);
or OR2 (N5612, N5604, N3893);
nor NOR2 (N5613, N5594, N979);
not NOT1 (N5614, N5607);
and AND4 (N5615, N5610, N359, N1256, N2924);
or OR3 (N5616, N5614, N4534, N2620);
xor XOR2 (N5617, N5606, N389);
and AND2 (N5618, N5603, N872);
not NOT1 (N5619, N5601);
or OR2 (N5620, N5609, N801);
and AND3 (N5621, N5617, N4920, N1603);
xor XOR2 (N5622, N5616, N3713);
xor XOR2 (N5623, N5615, N4489);
buf BUF1 (N5624, N5618);
xor XOR2 (N5625, N5612, N2440);
not NOT1 (N5626, N5623);
nand NAND2 (N5627, N5626, N1914);
nand NAND2 (N5628, N5619, N4155);
not NOT1 (N5629, N5602);
not NOT1 (N5630, N5622);
not NOT1 (N5631, N5627);
nand NAND4 (N5632, N5620, N2435, N739, N5188);
xor XOR2 (N5633, N5613, N2534);
or OR3 (N5634, N5624, N5137, N3672);
nand NAND2 (N5635, N5631, N1113);
nand NAND4 (N5636, N5632, N3577, N716, N4859);
buf BUF1 (N5637, N5621);
nand NAND3 (N5638, N5630, N4891, N3011);
buf BUF1 (N5639, N5638);
not NOT1 (N5640, N5633);
or OR2 (N5641, N5611, N4489);
nor NOR2 (N5642, N5640, N4362);
nor NOR3 (N5643, N5636, N2692, N5560);
buf BUF1 (N5644, N5642);
and AND4 (N5645, N5641, N2834, N2662, N1687);
nand NAND4 (N5646, N5637, N3741, N5318, N4699);
nor NOR4 (N5647, N5629, N4873, N1109, N2775);
or OR4 (N5648, N5634, N4860, N5151, N3081);
and AND4 (N5649, N5635, N3555, N4010, N2172);
xor XOR2 (N5650, N5625, N813);
nor NOR2 (N5651, N5646, N963);
nand NAND4 (N5652, N5644, N3940, N3991, N4618);
and AND3 (N5653, N5650, N1978, N2752);
or OR4 (N5654, N5653, N2309, N2531, N4183);
nor NOR2 (N5655, N5651, N2579);
nor NOR3 (N5656, N5654, N492, N2949);
and AND4 (N5657, N5645, N2934, N4220, N2460);
nand NAND2 (N5658, N5649, N4425);
or OR3 (N5659, N5656, N405, N967);
or OR4 (N5660, N5648, N4115, N2724, N5518);
and AND2 (N5661, N5639, N1149);
not NOT1 (N5662, N5661);
buf BUF1 (N5663, N5659);
xor XOR2 (N5664, N5655, N425);
xor XOR2 (N5665, N5657, N4875);
and AND2 (N5666, N5658, N4053);
xor XOR2 (N5667, N5628, N3679);
nor NOR4 (N5668, N5665, N84, N4329, N1271);
buf BUF1 (N5669, N5667);
or OR4 (N5670, N5647, N650, N1098, N3195);
or OR3 (N5671, N5643, N3597, N354);
or OR3 (N5672, N5670, N3662, N2823);
nor NOR2 (N5673, N5668, N5110);
nand NAND2 (N5674, N5663, N2382);
buf BUF1 (N5675, N5666);
xor XOR2 (N5676, N5660, N4140);
or OR4 (N5677, N5669, N4390, N4338, N2793);
xor XOR2 (N5678, N5672, N2110);
nor NOR2 (N5679, N5678, N3089);
or OR4 (N5680, N5677, N1642, N575, N710);
xor XOR2 (N5681, N5652, N1081);
nor NOR2 (N5682, N5674, N1278);
nor NOR3 (N5683, N5676, N3249, N1162);
or OR2 (N5684, N5664, N693);
or OR2 (N5685, N5682, N1319);
not NOT1 (N5686, N5683);
and AND4 (N5687, N5673, N5426, N2858, N534);
or OR2 (N5688, N5662, N1899);
nand NAND4 (N5689, N5684, N396, N3133, N2821);
not NOT1 (N5690, N5671);
or OR4 (N5691, N5679, N4537, N1362, N5468);
not NOT1 (N5692, N5675);
or OR4 (N5693, N5685, N4806, N5089, N985);
nand NAND2 (N5694, N5687, N2581);
xor XOR2 (N5695, N5691, N5419);
or OR4 (N5696, N5690, N5170, N5540, N3115);
nand NAND2 (N5697, N5688, N3751);
nor NOR4 (N5698, N5680, N728, N3705, N5589);
buf BUF1 (N5699, N5692);
and AND2 (N5700, N5693, N396);
nor NOR3 (N5701, N5697, N4040, N3825);
xor XOR2 (N5702, N5701, N4619);
and AND3 (N5703, N5700, N1191, N197);
nand NAND3 (N5704, N5698, N4333, N3131);
and AND2 (N5705, N5686, N723);
and AND3 (N5706, N5696, N2946, N2162);
nor NOR3 (N5707, N5705, N513, N1728);
or OR4 (N5708, N5699, N203, N3324, N4874);
and AND4 (N5709, N5702, N5225, N522, N2019);
or OR3 (N5710, N5694, N4731, N2182);
nand NAND4 (N5711, N5703, N670, N5456, N2448);
xor XOR2 (N5712, N5706, N2181);
not NOT1 (N5713, N5712);
xor XOR2 (N5714, N5708, N5576);
not NOT1 (N5715, N5714);
nand NAND4 (N5716, N5713, N4798, N2542, N3760);
xor XOR2 (N5717, N5704, N3242);
or OR4 (N5718, N5689, N186, N1619, N1556);
buf BUF1 (N5719, N5710);
nand NAND3 (N5720, N5716, N3298, N1695);
xor XOR2 (N5721, N5695, N1408);
buf BUF1 (N5722, N5721);
xor XOR2 (N5723, N5715, N4518);
buf BUF1 (N5724, N5717);
nor NOR2 (N5725, N5720, N2300);
xor XOR2 (N5726, N5718, N3260);
nand NAND3 (N5727, N5719, N5501, N4177);
nor NOR2 (N5728, N5727, N1957);
buf BUF1 (N5729, N5728);
buf BUF1 (N5730, N5711);
xor XOR2 (N5731, N5709, N1018);
or OR4 (N5732, N5723, N504, N3825, N3895);
not NOT1 (N5733, N5707);
buf BUF1 (N5734, N5733);
or OR2 (N5735, N5731, N4135);
xor XOR2 (N5736, N5722, N4766);
xor XOR2 (N5737, N5735, N4051);
and AND4 (N5738, N5729, N1801, N1043, N1781);
nor NOR3 (N5739, N5732, N3943, N4875);
buf BUF1 (N5740, N5725);
or OR4 (N5741, N5739, N1738, N608, N3318);
and AND3 (N5742, N5736, N856, N2777);
nor NOR4 (N5743, N5681, N2820, N5657, N2767);
and AND2 (N5744, N5730, N2231);
or OR3 (N5745, N5743, N3946, N1551);
and AND3 (N5746, N5745, N5339, N503);
not NOT1 (N5747, N5726);
and AND2 (N5748, N5747, N2699);
or OR3 (N5749, N5738, N996, N3973);
xor XOR2 (N5750, N5724, N1875);
xor XOR2 (N5751, N5744, N4575);
not NOT1 (N5752, N5740);
or OR2 (N5753, N5749, N1150);
nand NAND2 (N5754, N5750, N3873);
and AND3 (N5755, N5737, N506, N3393);
not NOT1 (N5756, N5754);
not NOT1 (N5757, N5748);
buf BUF1 (N5758, N5734);
buf BUF1 (N5759, N5752);
nor NOR2 (N5760, N5757, N270);
not NOT1 (N5761, N5742);
not NOT1 (N5762, N5760);
xor XOR2 (N5763, N5746, N196);
nand NAND4 (N5764, N5751, N4130, N2714, N4981);
nand NAND2 (N5765, N5763, N1109);
nand NAND2 (N5766, N5762, N2265);
xor XOR2 (N5767, N5756, N3999);
xor XOR2 (N5768, N5755, N3338);
xor XOR2 (N5769, N5758, N4727);
nand NAND2 (N5770, N5765, N1371);
nand NAND4 (N5771, N5761, N4393, N431, N2721);
nor NOR2 (N5772, N5771, N30);
buf BUF1 (N5773, N5769);
buf BUF1 (N5774, N5741);
nand NAND2 (N5775, N5759, N4799);
or OR3 (N5776, N5774, N5038, N362);
buf BUF1 (N5777, N5772);
xor XOR2 (N5778, N5776, N5485);
xor XOR2 (N5779, N5764, N460);
or OR2 (N5780, N5770, N1359);
buf BUF1 (N5781, N5780);
xor XOR2 (N5782, N5775, N5728);
buf BUF1 (N5783, N5778);
buf BUF1 (N5784, N5753);
xor XOR2 (N5785, N5781, N3739);
or OR4 (N5786, N5773, N866, N330, N5112);
and AND3 (N5787, N5786, N734, N2283);
nor NOR3 (N5788, N5768, N4491, N2828);
nor NOR4 (N5789, N5783, N1786, N2833, N2888);
and AND3 (N5790, N5766, N3992, N4814);
buf BUF1 (N5791, N5790);
or OR2 (N5792, N5789, N3088);
buf BUF1 (N5793, N5787);
or OR2 (N5794, N5792, N4397);
buf BUF1 (N5795, N5785);
not NOT1 (N5796, N5794);
xor XOR2 (N5797, N5788, N4759);
xor XOR2 (N5798, N5795, N3611);
not NOT1 (N5799, N5796);
not NOT1 (N5800, N5799);
buf BUF1 (N5801, N5797);
nand NAND3 (N5802, N5793, N441, N1539);
or OR2 (N5803, N5801, N1856);
not NOT1 (N5804, N5779);
xor XOR2 (N5805, N5802, N575);
not NOT1 (N5806, N5791);
nor NOR3 (N5807, N5784, N547, N1838);
not NOT1 (N5808, N5803);
nand NAND2 (N5809, N5777, N64);
and AND3 (N5810, N5806, N1575, N4512);
xor XOR2 (N5811, N5804, N3912);
nor NOR2 (N5812, N5810, N396);
and AND4 (N5813, N5800, N5325, N8, N3616);
nor NOR3 (N5814, N5809, N242, N1244);
buf BUF1 (N5815, N5813);
buf BUF1 (N5816, N5782);
nor NOR4 (N5817, N5815, N2455, N1692, N3057);
buf BUF1 (N5818, N5807);
nand NAND3 (N5819, N5814, N3331, N2143);
or OR2 (N5820, N5818, N5487);
nor NOR2 (N5821, N5812, N5122);
or OR3 (N5822, N5767, N5509, N4453);
or OR4 (N5823, N5805, N3646, N5585, N4259);
buf BUF1 (N5824, N5823);
or OR3 (N5825, N5822, N1991, N2836);
and AND3 (N5826, N5824, N203, N1852);
or OR2 (N5827, N5819, N36);
xor XOR2 (N5828, N5827, N4142);
nand NAND2 (N5829, N5811, N1219);
buf BUF1 (N5830, N5825);
and AND3 (N5831, N5816, N2244, N4571);
not NOT1 (N5832, N5820);
or OR4 (N5833, N5826, N857, N5275, N2380);
nand NAND4 (N5834, N5833, N475, N883, N5570);
and AND4 (N5835, N5834, N3169, N5466, N1684);
nand NAND2 (N5836, N5817, N1312);
nand NAND4 (N5837, N5808, N840, N155, N2496);
xor XOR2 (N5838, N5835, N299);
nand NAND4 (N5839, N5832, N855, N1479, N2808);
buf BUF1 (N5840, N5798);
nand NAND2 (N5841, N5829, N1992);
and AND2 (N5842, N5841, N1301);
or OR2 (N5843, N5836, N4136);
nor NOR2 (N5844, N5840, N5509);
nor NOR2 (N5845, N5843, N165);
buf BUF1 (N5846, N5839);
nand NAND4 (N5847, N5821, N3195, N521, N1294);
nand NAND2 (N5848, N5845, N4038);
not NOT1 (N5849, N5842);
nor NOR2 (N5850, N5831, N1718);
and AND2 (N5851, N5830, N4468);
not NOT1 (N5852, N5838);
not NOT1 (N5853, N5850);
xor XOR2 (N5854, N5844, N2479);
nor NOR2 (N5855, N5848, N2638);
or OR2 (N5856, N5828, N5378);
not NOT1 (N5857, N5855);
nor NOR3 (N5858, N5854, N361, N2411);
xor XOR2 (N5859, N5837, N5317);
nand NAND3 (N5860, N5849, N604, N834);
not NOT1 (N5861, N5846);
nand NAND2 (N5862, N5856, N1606);
not NOT1 (N5863, N5847);
or OR2 (N5864, N5852, N2298);
not NOT1 (N5865, N5858);
nor NOR4 (N5866, N5862, N3079, N939, N232);
xor XOR2 (N5867, N5851, N5305);
nand NAND2 (N5868, N5861, N1806);
nor NOR2 (N5869, N5860, N675);
not NOT1 (N5870, N5857);
and AND3 (N5871, N5865, N4262, N4971);
xor XOR2 (N5872, N5859, N72);
buf BUF1 (N5873, N5870);
nor NOR2 (N5874, N5864, N3829);
nand NAND4 (N5875, N5863, N1091, N3813, N3371);
or OR4 (N5876, N5872, N4493, N3495, N1491);
or OR2 (N5877, N5874, N1315);
nor NOR2 (N5878, N5871, N20);
nor NOR4 (N5879, N5868, N717, N4826, N1243);
nor NOR2 (N5880, N5853, N4467);
nand NAND3 (N5881, N5869, N1893, N5580);
nor NOR3 (N5882, N5879, N2901, N5677);
nand NAND2 (N5883, N5875, N4815);
buf BUF1 (N5884, N5881);
nand NAND4 (N5885, N5882, N4281, N4923, N2240);
buf BUF1 (N5886, N5883);
nand NAND4 (N5887, N5867, N5797, N5566, N831);
nor NOR2 (N5888, N5877, N2855);
nor NOR3 (N5889, N5866, N1158, N2870);
nor NOR2 (N5890, N5886, N5170);
buf BUF1 (N5891, N5873);
not NOT1 (N5892, N5887);
and AND3 (N5893, N5878, N3789, N3973);
or OR2 (N5894, N5888, N1314);
nand NAND3 (N5895, N5885, N1454, N4863);
nor NOR2 (N5896, N5891, N5175);
and AND2 (N5897, N5876, N1193);
not NOT1 (N5898, N5897);
not NOT1 (N5899, N5880);
nand NAND3 (N5900, N5894, N4827, N4527);
not NOT1 (N5901, N5895);
nor NOR4 (N5902, N5892, N2366, N605, N610);
nor NOR3 (N5903, N5899, N5723, N5355);
xor XOR2 (N5904, N5896, N1818);
nand NAND4 (N5905, N5893, N4243, N2204, N5747);
not NOT1 (N5906, N5898);
xor XOR2 (N5907, N5906, N749);
nor NOR4 (N5908, N5884, N5125, N1711, N5718);
and AND2 (N5909, N5901, N4546);
and AND3 (N5910, N5889, N1636, N5668);
xor XOR2 (N5911, N5903, N4736);
and AND2 (N5912, N5908, N3784);
or OR4 (N5913, N5905, N5212, N3909, N3369);
xor XOR2 (N5914, N5904, N5460);
not NOT1 (N5915, N5912);
xor XOR2 (N5916, N5890, N3512);
xor XOR2 (N5917, N5902, N2973);
or OR3 (N5918, N5900, N254, N5480);
not NOT1 (N5919, N5907);
and AND3 (N5920, N5914, N2332, N4350);
or OR2 (N5921, N5919, N3605);
and AND3 (N5922, N5916, N114, N2513);
xor XOR2 (N5923, N5909, N1576);
or OR2 (N5924, N5910, N3150);
not NOT1 (N5925, N5918);
buf BUF1 (N5926, N5925);
buf BUF1 (N5927, N5921);
nor NOR2 (N5928, N5927, N5432);
buf BUF1 (N5929, N5923);
or OR3 (N5930, N5929, N4907, N380);
not NOT1 (N5931, N5926);
nor NOR2 (N5932, N5917, N4881);
and AND3 (N5933, N5922, N1048, N3041);
not NOT1 (N5934, N5920);
nand NAND4 (N5935, N5934, N1303, N5571, N1257);
nand NAND2 (N5936, N5924, N1459);
nand NAND3 (N5937, N5932, N359, N2216);
buf BUF1 (N5938, N5931);
buf BUF1 (N5939, N5913);
nand NAND2 (N5940, N5915, N3587);
nand NAND4 (N5941, N5939, N1948, N4964, N1553);
nor NOR4 (N5942, N5941, N2354, N2715, N5326);
or OR2 (N5943, N5930, N4257);
nor NOR3 (N5944, N5937, N5649, N1817);
not NOT1 (N5945, N5911);
xor XOR2 (N5946, N5938, N1740);
buf BUF1 (N5947, N5946);
or OR4 (N5948, N5933, N3489, N3818, N3370);
buf BUF1 (N5949, N5945);
and AND2 (N5950, N5936, N4745);
buf BUF1 (N5951, N5935);
and AND4 (N5952, N5950, N2577, N61, N2513);
nand NAND2 (N5953, N5928, N377);
buf BUF1 (N5954, N5952);
or OR3 (N5955, N5943, N550, N3824);
nand NAND3 (N5956, N5944, N1831, N4458);
and AND3 (N5957, N5948, N4584, N4993);
nand NAND3 (N5958, N5942, N1775, N5735);
nand NAND2 (N5959, N5955, N5624);
nand NAND2 (N5960, N5954, N3170);
and AND2 (N5961, N5951, N2424);
nor NOR2 (N5962, N5961, N1747);
nor NOR2 (N5963, N5958, N1650);
buf BUF1 (N5964, N5959);
xor XOR2 (N5965, N5947, N598);
nor NOR3 (N5966, N5965, N2436, N4759);
and AND3 (N5967, N5956, N1536, N536);
xor XOR2 (N5968, N5962, N1331);
and AND4 (N5969, N5940, N2459, N4582, N4488);
or OR4 (N5970, N5966, N948, N5499, N5338);
and AND3 (N5971, N5960, N2744, N5761);
or OR2 (N5972, N5957, N1632);
buf BUF1 (N5973, N5970);
or OR4 (N5974, N5973, N2722, N2870, N1885);
xor XOR2 (N5975, N5969, N2508);
not NOT1 (N5976, N5975);
buf BUF1 (N5977, N5953);
and AND3 (N5978, N5964, N1864, N2778);
not NOT1 (N5979, N5972);
or OR3 (N5980, N5978, N1687, N4567);
and AND4 (N5981, N5977, N4884, N102, N111);
buf BUF1 (N5982, N5981);
nand NAND4 (N5983, N5967, N3935, N2838, N3154);
not NOT1 (N5984, N5980);
nor NOR4 (N5985, N5971, N1371, N1460, N5340);
nand NAND3 (N5986, N5968, N1510, N2314);
not NOT1 (N5987, N5984);
and AND2 (N5988, N5985, N4080);
not NOT1 (N5989, N5986);
buf BUF1 (N5990, N5976);
not NOT1 (N5991, N5974);
and AND4 (N5992, N5949, N2964, N5692, N3005);
or OR4 (N5993, N5983, N513, N4337, N5206);
and AND3 (N5994, N5963, N2261, N5219);
nor NOR2 (N5995, N5990, N5993);
buf BUF1 (N5996, N4318);
nor NOR4 (N5997, N5987, N1189, N5208, N4932);
or OR2 (N5998, N5991, N637);
xor XOR2 (N5999, N5996, N1658);
buf BUF1 (N6000, N5982);
nor NOR2 (N6001, N6000, N2743);
nand NAND3 (N6002, N6001, N3522, N5195);
not NOT1 (N6003, N5992);
nor NOR3 (N6004, N5997, N207, N1586);
xor XOR2 (N6005, N5999, N5506);
buf BUF1 (N6006, N5995);
nand NAND4 (N6007, N6004, N5398, N4388, N1964);
not NOT1 (N6008, N5994);
buf BUF1 (N6009, N6007);
buf BUF1 (N6010, N6009);
nor NOR4 (N6011, N6003, N3422, N2694, N4402);
buf BUF1 (N6012, N6010);
nand NAND3 (N6013, N6005, N1795, N5119);
nand NAND4 (N6014, N6012, N31, N1086, N182);
and AND4 (N6015, N5979, N5861, N5579, N4449);
nand NAND4 (N6016, N6011, N1984, N5038, N3474);
nor NOR4 (N6017, N6014, N2768, N4189, N5983);
nand NAND2 (N6018, N6013, N434);
not NOT1 (N6019, N6008);
and AND2 (N6020, N6015, N3036);
nand NAND4 (N6021, N6020, N1287, N1752, N4827);
xor XOR2 (N6022, N5988, N1691);
not NOT1 (N6023, N6021);
not NOT1 (N6024, N5998);
or OR3 (N6025, N6019, N115, N1368);
not NOT1 (N6026, N6016);
nor NOR2 (N6027, N6024, N3490);
buf BUF1 (N6028, N6002);
nand NAND2 (N6029, N6022, N1119);
nand NAND4 (N6030, N6027, N4387, N5866, N5483);
xor XOR2 (N6031, N6028, N899);
nand NAND2 (N6032, N6023, N460);
and AND2 (N6033, N6029, N5435);
and AND2 (N6034, N6017, N1714);
xor XOR2 (N6035, N6026, N5791);
xor XOR2 (N6036, N6033, N1150);
not NOT1 (N6037, N6018);
xor XOR2 (N6038, N6035, N2491);
xor XOR2 (N6039, N6038, N778);
xor XOR2 (N6040, N6034, N3610);
not NOT1 (N6041, N6032);
xor XOR2 (N6042, N6025, N3904);
and AND4 (N6043, N6039, N4650, N5323, N1931);
and AND2 (N6044, N6043, N5280);
buf BUF1 (N6045, N6006);
xor XOR2 (N6046, N6031, N5702);
and AND4 (N6047, N6046, N4999, N3654, N5027);
or OR3 (N6048, N6037, N1753, N1899);
nor NOR3 (N6049, N6044, N512, N322);
or OR4 (N6050, N6045, N817, N3605, N3718);
or OR3 (N6051, N5989, N5560, N2665);
nor NOR3 (N6052, N6041, N1220, N1252);
xor XOR2 (N6053, N6036, N3086);
and AND3 (N6054, N6042, N2338, N2676);
buf BUF1 (N6055, N6040);
not NOT1 (N6056, N6049);
not NOT1 (N6057, N6051);
and AND4 (N6058, N6052, N1025, N4210, N2862);
or OR2 (N6059, N6030, N3065);
or OR3 (N6060, N6054, N4255, N1940);
not NOT1 (N6061, N6050);
nor NOR4 (N6062, N6048, N736, N2355, N5389);
buf BUF1 (N6063, N6056);
xor XOR2 (N6064, N6055, N4341);
xor XOR2 (N6065, N6063, N3982);
not NOT1 (N6066, N6058);
or OR2 (N6067, N6064, N3776);
or OR4 (N6068, N6062, N267, N4191, N1391);
xor XOR2 (N6069, N6057, N6065);
buf BUF1 (N6070, N2368);
or OR4 (N6071, N6067, N2878, N4420, N5456);
buf BUF1 (N6072, N6061);
xor XOR2 (N6073, N6071, N2025);
or OR3 (N6074, N6066, N3783, N5539);
and AND4 (N6075, N6073, N1182, N1170, N4182);
or OR3 (N6076, N6069, N772, N405);
or OR3 (N6077, N6074, N2233, N3581);
xor XOR2 (N6078, N6053, N1723);
buf BUF1 (N6079, N6076);
and AND2 (N6080, N6077, N3000);
nor NOR2 (N6081, N6059, N1978);
nand NAND2 (N6082, N6078, N2750);
nor NOR3 (N6083, N6080, N2132, N1843);
not NOT1 (N6084, N6068);
and AND3 (N6085, N6082, N5943, N3863);
and AND4 (N6086, N6084, N2677, N1186, N5944);
and AND2 (N6087, N6079, N4336);
xor XOR2 (N6088, N6087, N517);
and AND2 (N6089, N6070, N5749);
not NOT1 (N6090, N6075);
not NOT1 (N6091, N6090);
nor NOR4 (N6092, N6081, N6019, N996, N6001);
not NOT1 (N6093, N6083);
nor NOR3 (N6094, N6047, N3943, N285);
nand NAND4 (N6095, N6060, N2332, N3370, N4291);
and AND2 (N6096, N6093, N2633);
not NOT1 (N6097, N6089);
and AND3 (N6098, N6085, N5728, N6087);
xor XOR2 (N6099, N6096, N3526);
buf BUF1 (N6100, N6088);
xor XOR2 (N6101, N6072, N310);
or OR2 (N6102, N6099, N2377);
nor NOR3 (N6103, N6094, N4455, N2178);
buf BUF1 (N6104, N6092);
or OR2 (N6105, N6104, N4395);
not NOT1 (N6106, N6105);
not NOT1 (N6107, N6098);
and AND3 (N6108, N6086, N1551, N1435);
not NOT1 (N6109, N6095);
nor NOR2 (N6110, N6108, N201);
not NOT1 (N6111, N6106);
nor NOR4 (N6112, N6097, N3437, N1298, N2511);
xor XOR2 (N6113, N6109, N2247);
nand NAND4 (N6114, N6107, N1990, N618, N4846);
and AND4 (N6115, N6101, N3493, N5092, N884);
or OR3 (N6116, N6112, N4012, N3201);
buf BUF1 (N6117, N6115);
nand NAND2 (N6118, N6116, N5271);
buf BUF1 (N6119, N6100);
xor XOR2 (N6120, N6118, N5905);
buf BUF1 (N6121, N6102);
not NOT1 (N6122, N6113);
or OR2 (N6123, N6114, N3986);
nand NAND3 (N6124, N6122, N1721, N266);
or OR3 (N6125, N6111, N5428, N5084);
and AND3 (N6126, N6119, N4864, N664);
buf BUF1 (N6127, N6124);
or OR3 (N6128, N6127, N3193, N2399);
xor XOR2 (N6129, N6121, N4285);
or OR4 (N6130, N6110, N5446, N1538, N2616);
and AND4 (N6131, N6117, N4208, N4964, N5656);
xor XOR2 (N6132, N6103, N2387);
buf BUF1 (N6133, N6125);
and AND2 (N6134, N6091, N1974);
buf BUF1 (N6135, N6133);
buf BUF1 (N6136, N6131);
nor NOR2 (N6137, N6132, N1694);
buf BUF1 (N6138, N6137);
nor NOR3 (N6139, N6134, N1826, N3594);
nand NAND2 (N6140, N6139, N3216);
buf BUF1 (N6141, N6130);
not NOT1 (N6142, N6120);
nand NAND2 (N6143, N6141, N2090);
not NOT1 (N6144, N6140);
buf BUF1 (N6145, N6138);
nand NAND3 (N6146, N6135, N863, N882);
buf BUF1 (N6147, N6123);
xor XOR2 (N6148, N6144, N3912);
nand NAND3 (N6149, N6143, N4837, N1115);
buf BUF1 (N6150, N6126);
not NOT1 (N6151, N6150);
xor XOR2 (N6152, N6142, N4434);
and AND3 (N6153, N6145, N1922, N2997);
and AND3 (N6154, N6148, N5552, N5667);
buf BUF1 (N6155, N6153);
nand NAND4 (N6156, N6146, N527, N1941, N3475);
xor XOR2 (N6157, N6147, N3531);
nand NAND4 (N6158, N6154, N3886, N5276, N685);
not NOT1 (N6159, N6151);
xor XOR2 (N6160, N6157, N3668);
nor NOR4 (N6161, N6152, N195, N1933, N5656);
nand NAND2 (N6162, N6160, N319);
and AND3 (N6163, N6149, N2190, N5479);
or OR2 (N6164, N6161, N4755);
not NOT1 (N6165, N6163);
nand NAND4 (N6166, N6158, N5109, N4970, N1326);
not NOT1 (N6167, N6159);
nor NOR4 (N6168, N6128, N4455, N286, N5440);
nand NAND4 (N6169, N6164, N5123, N1647, N3097);
xor XOR2 (N6170, N6166, N578);
not NOT1 (N6171, N6129);
xor XOR2 (N6172, N6155, N179);
nor NOR4 (N6173, N6156, N5507, N4153, N2918);
nor NOR4 (N6174, N6169, N616, N2725, N2560);
buf BUF1 (N6175, N6173);
xor XOR2 (N6176, N6162, N3294);
xor XOR2 (N6177, N6167, N579);
not NOT1 (N6178, N6170);
buf BUF1 (N6179, N6176);
xor XOR2 (N6180, N6171, N5521);
not NOT1 (N6181, N6172);
nor NOR2 (N6182, N6177, N3482);
nor NOR2 (N6183, N6168, N1994);
not NOT1 (N6184, N6136);
buf BUF1 (N6185, N6180);
and AND2 (N6186, N6179, N425);
not NOT1 (N6187, N6186);
nor NOR2 (N6188, N6175, N347);
buf BUF1 (N6189, N6165);
not NOT1 (N6190, N6181);
nand NAND3 (N6191, N6182, N3628, N3432);
nand NAND3 (N6192, N6178, N689, N3591);
nand NAND2 (N6193, N6185, N154);
buf BUF1 (N6194, N6187);
buf BUF1 (N6195, N6190);
nor NOR3 (N6196, N6183, N3664, N4600);
xor XOR2 (N6197, N6193, N6040);
buf BUF1 (N6198, N6194);
and AND2 (N6199, N6198, N1341);
buf BUF1 (N6200, N6191);
not NOT1 (N6201, N6189);
not NOT1 (N6202, N6197);
buf BUF1 (N6203, N6188);
buf BUF1 (N6204, N6203);
and AND2 (N6205, N6202, N979);
and AND4 (N6206, N6195, N2718, N926, N3069);
nor NOR3 (N6207, N6204, N3026, N5924);
buf BUF1 (N6208, N6207);
xor XOR2 (N6209, N6200, N1477);
or OR3 (N6210, N6206, N3417, N1255);
not NOT1 (N6211, N6174);
and AND2 (N6212, N6208, N4624);
nor NOR3 (N6213, N6209, N4279, N5469);
and AND2 (N6214, N6211, N1649);
xor XOR2 (N6215, N6201, N2997);
xor XOR2 (N6216, N6184, N5945);
nand NAND3 (N6217, N6214, N4746, N1495);
not NOT1 (N6218, N6217);
nand NAND3 (N6219, N6215, N2802, N598);
nand NAND2 (N6220, N6213, N3364);
nor NOR4 (N6221, N6199, N2905, N2365, N4036);
xor XOR2 (N6222, N6218, N4556);
xor XOR2 (N6223, N6196, N1977);
not NOT1 (N6224, N6221);
or OR3 (N6225, N6223, N3020, N2244);
and AND3 (N6226, N6216, N2380, N2162);
xor XOR2 (N6227, N6222, N2192);
and AND4 (N6228, N6220, N2353, N4974, N1071);
xor XOR2 (N6229, N6225, N3695);
and AND2 (N6230, N6226, N3429);
or OR3 (N6231, N6192, N784, N507);
not NOT1 (N6232, N6205);
nand NAND2 (N6233, N6230, N449);
xor XOR2 (N6234, N6224, N5564);
and AND3 (N6235, N6234, N1753, N3765);
and AND2 (N6236, N6210, N5423);
buf BUF1 (N6237, N6231);
buf BUF1 (N6238, N6235);
and AND2 (N6239, N6228, N2317);
not NOT1 (N6240, N6236);
not NOT1 (N6241, N6219);
nand NAND4 (N6242, N6240, N5246, N4063, N1468);
xor XOR2 (N6243, N6237, N3027);
nand NAND2 (N6244, N6239, N4551);
and AND4 (N6245, N6232, N2073, N4157, N3576);
buf BUF1 (N6246, N6245);
not NOT1 (N6247, N6229);
nand NAND2 (N6248, N6233, N3879);
nand NAND2 (N6249, N6247, N970);
not NOT1 (N6250, N6212);
or OR2 (N6251, N6227, N730);
buf BUF1 (N6252, N6244);
xor XOR2 (N6253, N6241, N2004);
not NOT1 (N6254, N6248);
not NOT1 (N6255, N6246);
nor NOR2 (N6256, N6249, N4913);
nor NOR4 (N6257, N6238, N71, N1783, N2609);
or OR3 (N6258, N6256, N5561, N4221);
or OR2 (N6259, N6257, N964);
nor NOR2 (N6260, N6255, N1203);
nand NAND3 (N6261, N6254, N1875, N2589);
nand NAND4 (N6262, N6243, N4267, N4590, N4509);
or OR4 (N6263, N6242, N2120, N121, N2311);
buf BUF1 (N6264, N6251);
nor NOR4 (N6265, N6250, N939, N6012, N1465);
and AND4 (N6266, N6262, N882, N5541, N5947);
nor NOR3 (N6267, N6266, N398, N1901);
buf BUF1 (N6268, N6259);
and AND3 (N6269, N6263, N2513, N3024);
nand NAND2 (N6270, N6258, N2487);
not NOT1 (N6271, N6269);
xor XOR2 (N6272, N6265, N19);
xor XOR2 (N6273, N6261, N3158);
nor NOR3 (N6274, N6267, N4359, N638);
or OR2 (N6275, N6271, N2749);
buf BUF1 (N6276, N6252);
not NOT1 (N6277, N6272);
and AND2 (N6278, N6260, N1769);
not NOT1 (N6279, N6276);
buf BUF1 (N6280, N6273);
not NOT1 (N6281, N6270);
not NOT1 (N6282, N6277);
and AND4 (N6283, N6264, N46, N720, N6146);
nand NAND4 (N6284, N6278, N4308, N5204, N5135);
nor NOR4 (N6285, N6281, N5644, N4366, N1106);
nand NAND3 (N6286, N6279, N4993, N5621);
buf BUF1 (N6287, N6253);
not NOT1 (N6288, N6280);
nor NOR3 (N6289, N6286, N4819, N598);
or OR4 (N6290, N6289, N4145, N3731, N3468);
nand NAND4 (N6291, N6274, N2569, N3851, N3959);
xor XOR2 (N6292, N6290, N2855);
nor NOR2 (N6293, N6268, N3086);
and AND2 (N6294, N6284, N269);
nand NAND3 (N6295, N6291, N2223, N2912);
and AND3 (N6296, N6294, N6181, N1723);
not NOT1 (N6297, N6282);
nand NAND4 (N6298, N6297, N4198, N1299, N3726);
xor XOR2 (N6299, N6293, N4050);
nor NOR3 (N6300, N6287, N1271, N6096);
not NOT1 (N6301, N6296);
xor XOR2 (N6302, N6288, N401);
nand NAND4 (N6303, N6275, N4040, N6109, N5205);
nor NOR3 (N6304, N6285, N5440, N5427);
and AND2 (N6305, N6292, N1022);
buf BUF1 (N6306, N6283);
and AND3 (N6307, N6305, N798, N397);
and AND4 (N6308, N6307, N3638, N3216, N970);
not NOT1 (N6309, N6298);
not NOT1 (N6310, N6306);
or OR3 (N6311, N6304, N1561, N1594);
buf BUF1 (N6312, N6295);
xor XOR2 (N6313, N6303, N2526);
nand NAND2 (N6314, N6311, N5379);
not NOT1 (N6315, N6312);
or OR2 (N6316, N6310, N1977);
xor XOR2 (N6317, N6302, N4870);
and AND3 (N6318, N6301, N1530, N2809);
nand NAND2 (N6319, N6299, N2104);
not NOT1 (N6320, N6300);
not NOT1 (N6321, N6320);
nand NAND2 (N6322, N6321, N3513);
xor XOR2 (N6323, N6322, N3554);
and AND2 (N6324, N6323, N1800);
or OR2 (N6325, N6315, N3603);
or OR4 (N6326, N6313, N4274, N1529, N6101);
nor NOR4 (N6327, N6326, N4092, N6036, N1722);
or OR2 (N6328, N6327, N4403);
and AND4 (N6329, N6317, N4051, N1161, N1161);
and AND2 (N6330, N6309, N1519);
and AND2 (N6331, N6319, N4791);
buf BUF1 (N6332, N6314);
not NOT1 (N6333, N6332);
or OR2 (N6334, N6331, N1679);
not NOT1 (N6335, N6325);
not NOT1 (N6336, N6333);
nor NOR3 (N6337, N6334, N5078, N2899);
and AND2 (N6338, N6316, N433);
buf BUF1 (N6339, N6335);
not NOT1 (N6340, N6339);
or OR4 (N6341, N6340, N5404, N5459, N1697);
buf BUF1 (N6342, N6337);
or OR3 (N6343, N6330, N6168, N3830);
nor NOR2 (N6344, N6342, N4611);
nor NOR3 (N6345, N6329, N4910, N1973);
nand NAND3 (N6346, N6345, N5440, N3025);
and AND4 (N6347, N6341, N5876, N825, N4502);
buf BUF1 (N6348, N6343);
or OR4 (N6349, N6308, N630, N958, N4135);
and AND4 (N6350, N6336, N2815, N3471, N2117);
not NOT1 (N6351, N6350);
nor NOR3 (N6352, N6348, N1512, N5898);
nand NAND2 (N6353, N6349, N1820);
and AND4 (N6354, N6352, N3372, N5885, N3336);
xor XOR2 (N6355, N6353, N3024);
buf BUF1 (N6356, N6324);
xor XOR2 (N6357, N6346, N4120);
and AND3 (N6358, N6354, N3216, N2827);
xor XOR2 (N6359, N6347, N3873);
nor NOR3 (N6360, N6356, N4808, N4852);
not NOT1 (N6361, N6328);
buf BUF1 (N6362, N6351);
buf BUF1 (N6363, N6344);
xor XOR2 (N6364, N6362, N3126);
buf BUF1 (N6365, N6363);
or OR2 (N6366, N6355, N2669);
or OR2 (N6367, N6364, N5878);
or OR2 (N6368, N6357, N2350);
nor NOR4 (N6369, N6367, N4136, N489, N2618);
xor XOR2 (N6370, N6365, N1596);
not NOT1 (N6371, N6318);
nand NAND4 (N6372, N6338, N4790, N1146, N3488);
and AND3 (N6373, N6361, N2767, N4443);
nor NOR3 (N6374, N6369, N3863, N171);
xor XOR2 (N6375, N6372, N2688);
not NOT1 (N6376, N6371);
not NOT1 (N6377, N6368);
nand NAND4 (N6378, N6374, N2163, N589, N335);
or OR3 (N6379, N6376, N2467, N3726);
nand NAND4 (N6380, N6379, N1613, N4495, N2850);
nand NAND4 (N6381, N6360, N5045, N1574, N6126);
buf BUF1 (N6382, N6373);
not NOT1 (N6383, N6370);
nand NAND4 (N6384, N6377, N3846, N600, N3365);
nor NOR2 (N6385, N6375, N5591);
or OR2 (N6386, N6359, N2419);
not NOT1 (N6387, N6385);
buf BUF1 (N6388, N6381);
and AND3 (N6389, N6386, N1715, N6036);
nand NAND4 (N6390, N6358, N597, N4085, N5875);
and AND4 (N6391, N6387, N4826, N6290, N5634);
or OR4 (N6392, N6383, N912, N1099, N3686);
and AND3 (N6393, N6382, N2677, N4549);
xor XOR2 (N6394, N6366, N2797);
nand NAND4 (N6395, N6392, N2245, N5906, N5039);
not NOT1 (N6396, N6389);
not NOT1 (N6397, N6394);
xor XOR2 (N6398, N6380, N3630);
or OR3 (N6399, N6393, N2254, N6105);
buf BUF1 (N6400, N6396);
nand NAND2 (N6401, N6378, N1290);
or OR2 (N6402, N6390, N5990);
nor NOR4 (N6403, N6395, N3261, N2576, N5937);
nand NAND3 (N6404, N6388, N3900, N323);
not NOT1 (N6405, N6400);
and AND2 (N6406, N6391, N3196);
and AND3 (N6407, N6406, N4895, N1923);
xor XOR2 (N6408, N6407, N689);
and AND2 (N6409, N6408, N5062);
not NOT1 (N6410, N6404);
or OR2 (N6411, N6398, N5170);
nor NOR2 (N6412, N6397, N1047);
or OR2 (N6413, N6409, N1619);
and AND2 (N6414, N6403, N2687);
and AND4 (N6415, N6405, N5736, N6044, N4501);
not NOT1 (N6416, N6410);
buf BUF1 (N6417, N6412);
buf BUF1 (N6418, N6414);
buf BUF1 (N6419, N6384);
or OR2 (N6420, N6416, N674);
not NOT1 (N6421, N6402);
xor XOR2 (N6422, N6415, N4540);
xor XOR2 (N6423, N6420, N3041);
xor XOR2 (N6424, N6417, N3261);
nor NOR4 (N6425, N6418, N5451, N4478, N5612);
nor NOR2 (N6426, N6425, N2230);
and AND2 (N6427, N6424, N3359);
nor NOR4 (N6428, N6413, N5289, N2200, N89);
or OR4 (N6429, N6428, N1982, N349, N4274);
buf BUF1 (N6430, N6429);
xor XOR2 (N6431, N6430, N4977);
or OR2 (N6432, N6427, N4131);
buf BUF1 (N6433, N6421);
or OR3 (N6434, N6432, N3329, N1388);
or OR2 (N6435, N6423, N3268);
not NOT1 (N6436, N6419);
xor XOR2 (N6437, N6434, N2813);
not NOT1 (N6438, N6411);
xor XOR2 (N6439, N6433, N2980);
or OR3 (N6440, N6426, N5550, N3956);
xor XOR2 (N6441, N6440, N3019);
buf BUF1 (N6442, N6441);
buf BUF1 (N6443, N6401);
and AND3 (N6444, N6438, N3575, N3748);
not NOT1 (N6445, N6422);
xor XOR2 (N6446, N6439, N2832);
buf BUF1 (N6447, N6437);
nand NAND2 (N6448, N6435, N2842);
and AND4 (N6449, N6448, N3110, N5552, N2557);
not NOT1 (N6450, N6444);
xor XOR2 (N6451, N6450, N5187);
not NOT1 (N6452, N6431);
nor NOR3 (N6453, N6443, N4621, N4663);
nand NAND3 (N6454, N6445, N790, N3433);
not NOT1 (N6455, N6436);
xor XOR2 (N6456, N6399, N1352);
nor NOR2 (N6457, N6454, N834);
xor XOR2 (N6458, N6446, N2001);
buf BUF1 (N6459, N6453);
or OR4 (N6460, N6456, N2415, N112, N652);
or OR2 (N6461, N6460, N4294);
or OR2 (N6462, N6459, N4202);
or OR4 (N6463, N6461, N1899, N4658, N3772);
not NOT1 (N6464, N6458);
not NOT1 (N6465, N6463);
not NOT1 (N6466, N6442);
nand NAND2 (N6467, N6464, N101);
nand NAND2 (N6468, N6447, N533);
or OR3 (N6469, N6455, N5600, N5085);
buf BUF1 (N6470, N6462);
or OR3 (N6471, N6466, N715, N2067);
and AND4 (N6472, N6469, N1815, N2, N4523);
and AND4 (N6473, N6471, N5684, N3594, N597);
nor NOR2 (N6474, N6470, N2105);
or OR2 (N6475, N6457, N4125);
not NOT1 (N6476, N6473);
nand NAND4 (N6477, N6452, N3628, N5127, N664);
not NOT1 (N6478, N6472);
nand NAND3 (N6479, N6474, N1146, N2553);
xor XOR2 (N6480, N6478, N2829);
or OR3 (N6481, N6449, N592, N4409);
not NOT1 (N6482, N6475);
or OR4 (N6483, N6465, N5865, N945, N5741);
not NOT1 (N6484, N6451);
or OR4 (N6485, N6484, N848, N4323, N3548);
and AND2 (N6486, N6480, N5022);
not NOT1 (N6487, N6482);
nand NAND3 (N6488, N6477, N3233, N5195);
xor XOR2 (N6489, N6467, N5168);
nand NAND2 (N6490, N6483, N2363);
or OR4 (N6491, N6487, N1609, N3317, N2828);
or OR2 (N6492, N6479, N4424);
and AND3 (N6493, N6476, N5970, N3435);
nand NAND3 (N6494, N6485, N1272, N2347);
and AND2 (N6495, N6486, N4789);
buf BUF1 (N6496, N6481);
nor NOR4 (N6497, N6492, N3609, N2503, N1984);
nor NOR4 (N6498, N6489, N6488, N5671, N712);
nor NOR4 (N6499, N516, N122, N6395, N4646);
nor NOR3 (N6500, N6499, N413, N5461);
and AND2 (N6501, N6493, N2018);
and AND3 (N6502, N6498, N1896, N3611);
buf BUF1 (N6503, N6491);
nand NAND2 (N6504, N6496, N5377);
or OR4 (N6505, N6490, N4277, N2575, N1046);
and AND3 (N6506, N6504, N2088, N4680);
buf BUF1 (N6507, N6495);
nor NOR2 (N6508, N6502, N3817);
or OR4 (N6509, N6497, N332, N2537, N6012);
and AND4 (N6510, N6506, N243, N2996, N2921);
nand NAND2 (N6511, N6509, N498);
not NOT1 (N6512, N6505);
buf BUF1 (N6513, N6468);
nand NAND4 (N6514, N6511, N6070, N3562, N3038);
or OR4 (N6515, N6500, N1258, N6403, N1420);
nand NAND3 (N6516, N6494, N3035, N789);
xor XOR2 (N6517, N6516, N2000);
nand NAND2 (N6518, N6512, N5733);
buf BUF1 (N6519, N6518);
nor NOR3 (N6520, N6513, N5382, N4924);
nand NAND4 (N6521, N6503, N827, N1868, N167);
or OR3 (N6522, N6510, N1488, N4316);
or OR2 (N6523, N6515, N6336);
not NOT1 (N6524, N6523);
and AND3 (N6525, N6517, N4756, N1217);
nand NAND4 (N6526, N6525, N4521, N226, N1485);
buf BUF1 (N6527, N6514);
buf BUF1 (N6528, N6508);
nor NOR2 (N6529, N6524, N1569);
nand NAND4 (N6530, N6521, N4136, N3775, N5454);
and AND4 (N6531, N6507, N946, N242, N174);
nor NOR4 (N6532, N6501, N1716, N1685, N702);
and AND4 (N6533, N6530, N5159, N1461, N2236);
not NOT1 (N6534, N6527);
and AND2 (N6535, N6526, N512);
buf BUF1 (N6536, N6533);
not NOT1 (N6537, N6522);
nand NAND4 (N6538, N6519, N56, N4550, N826);
buf BUF1 (N6539, N6537);
buf BUF1 (N6540, N6539);
or OR2 (N6541, N6528, N730);
and AND4 (N6542, N6529, N1119, N4904, N5018);
or OR3 (N6543, N6532, N894, N3376);
buf BUF1 (N6544, N6541);
nor NOR4 (N6545, N6531, N3630, N1284, N1231);
not NOT1 (N6546, N6542);
and AND3 (N6547, N6544, N322, N4593);
nor NOR2 (N6548, N6520, N5256);
and AND2 (N6549, N6535, N6362);
and AND3 (N6550, N6548, N2307, N460);
buf BUF1 (N6551, N6538);
nor NOR2 (N6552, N6549, N926);
buf BUF1 (N6553, N6551);
xor XOR2 (N6554, N6543, N2113);
and AND3 (N6555, N6552, N3292, N2469);
nor NOR4 (N6556, N6534, N2160, N352, N4471);
or OR3 (N6557, N6545, N412, N4561);
and AND3 (N6558, N6550, N6328, N2754);
xor XOR2 (N6559, N6558, N828);
nand NAND4 (N6560, N6559, N4013, N3171, N6177);
and AND2 (N6561, N6540, N445);
nor NOR2 (N6562, N6555, N3745);
or OR4 (N6563, N6557, N5838, N4067, N4381);
or OR2 (N6564, N6562, N3621);
or OR3 (N6565, N6560, N1545, N4243);
not NOT1 (N6566, N6553);
buf BUF1 (N6567, N6561);
buf BUF1 (N6568, N6565);
nand NAND4 (N6569, N6547, N3141, N2449, N5586);
buf BUF1 (N6570, N6556);
or OR2 (N6571, N6536, N1103);
and AND3 (N6572, N6571, N4845, N3290);
buf BUF1 (N6573, N6566);
or OR4 (N6574, N6572, N6322, N2074, N1369);
nor NOR3 (N6575, N6554, N2379, N4653);
nor NOR2 (N6576, N6575, N2356);
or OR2 (N6577, N6573, N1734);
or OR3 (N6578, N6568, N4852, N4243);
or OR3 (N6579, N6563, N4552, N4304);
or OR4 (N6580, N6570, N5424, N1758, N2474);
or OR2 (N6581, N6564, N113);
nor NOR2 (N6582, N6580, N3501);
not NOT1 (N6583, N6576);
or OR3 (N6584, N6546, N1625, N2187);
not NOT1 (N6585, N6567);
buf BUF1 (N6586, N6578);
or OR2 (N6587, N6574, N1234);
buf BUF1 (N6588, N6587);
not NOT1 (N6589, N6577);
nand NAND2 (N6590, N6589, N4216);
buf BUF1 (N6591, N6582);
nor NOR3 (N6592, N6586, N5660, N5978);
or OR4 (N6593, N6583, N2331, N4214, N1508);
and AND3 (N6594, N6581, N3965, N3559);
nor NOR2 (N6595, N6579, N2098);
not NOT1 (N6596, N6588);
xor XOR2 (N6597, N6585, N5037);
and AND3 (N6598, N6591, N4460, N491);
nor NOR3 (N6599, N6590, N2207, N4188);
and AND4 (N6600, N6596, N3471, N2718, N2116);
and AND2 (N6601, N6592, N3974);
nor NOR4 (N6602, N6598, N2260, N2386, N5117);
not NOT1 (N6603, N6584);
xor XOR2 (N6604, N6601, N1988);
and AND4 (N6605, N6603, N6043, N4493, N6121);
buf BUF1 (N6606, N6595);
nand NAND4 (N6607, N6597, N2998, N1772, N6426);
and AND4 (N6608, N6594, N128, N2645, N385);
or OR2 (N6609, N6569, N6479);
xor XOR2 (N6610, N6606, N3759);
and AND2 (N6611, N6602, N1670);
buf BUF1 (N6612, N6609);
nand NAND3 (N6613, N6605, N357, N1894);
not NOT1 (N6614, N6610);
buf BUF1 (N6615, N6599);
nand NAND3 (N6616, N6614, N4665, N4100);
and AND2 (N6617, N6600, N380);
xor XOR2 (N6618, N6608, N5090);
xor XOR2 (N6619, N6607, N4151);
nand NAND4 (N6620, N6611, N1284, N2174, N3000);
or OR4 (N6621, N6613, N2189, N3674, N2200);
and AND2 (N6622, N6616, N3933);
or OR4 (N6623, N6615, N835, N2467, N1740);
nand NAND2 (N6624, N6618, N2152);
nor NOR2 (N6625, N6624, N4547);
xor XOR2 (N6626, N6622, N1255);
xor XOR2 (N6627, N6593, N6141);
nor NOR2 (N6628, N6617, N4577);
nand NAND4 (N6629, N6628, N4712, N1053, N1911);
buf BUF1 (N6630, N6623);
nor NOR4 (N6631, N6620, N1376, N6150, N6211);
or OR4 (N6632, N6630, N4605, N4726, N998);
xor XOR2 (N6633, N6631, N5860);
and AND4 (N6634, N6632, N5763, N5728, N1545);
not NOT1 (N6635, N6612);
not NOT1 (N6636, N6621);
and AND3 (N6637, N6633, N2996, N3750);
buf BUF1 (N6638, N6626);
xor XOR2 (N6639, N6604, N4702);
buf BUF1 (N6640, N6619);
xor XOR2 (N6641, N6625, N1982);
nand NAND2 (N6642, N6639, N3139);
or OR4 (N6643, N6640, N701, N756, N429);
xor XOR2 (N6644, N6636, N6574);
not NOT1 (N6645, N6634);
and AND4 (N6646, N6642, N4971, N5526, N878);
xor XOR2 (N6647, N6645, N3888);
not NOT1 (N6648, N6647);
nor NOR4 (N6649, N6648, N6016, N3979, N4791);
buf BUF1 (N6650, N6629);
nor NOR2 (N6651, N6646, N5436);
buf BUF1 (N6652, N6650);
xor XOR2 (N6653, N6651, N2159);
and AND2 (N6654, N6643, N2112);
not NOT1 (N6655, N6637);
not NOT1 (N6656, N6652);
or OR3 (N6657, N6641, N4522, N6458);
nand NAND4 (N6658, N6644, N4125, N2454, N617);
not NOT1 (N6659, N6638);
buf BUF1 (N6660, N6659);
or OR4 (N6661, N6654, N3572, N2880, N2919);
buf BUF1 (N6662, N6656);
and AND4 (N6663, N6653, N1796, N4608, N473);
nor NOR3 (N6664, N6658, N6118, N4306);
nor NOR2 (N6665, N6661, N5763);
buf BUF1 (N6666, N6663);
nand NAND2 (N6667, N6662, N3977);
xor XOR2 (N6668, N6664, N4600);
and AND2 (N6669, N6668, N1263);
and AND2 (N6670, N6666, N3895);
xor XOR2 (N6671, N6649, N6341);
and AND2 (N6672, N6669, N3445);
xor XOR2 (N6673, N6655, N5340);
nand NAND4 (N6674, N6670, N3943, N2481, N5384);
xor XOR2 (N6675, N6627, N3371);
and AND2 (N6676, N6660, N968);
and AND4 (N6677, N6675, N4860, N5218, N4496);
not NOT1 (N6678, N6667);
buf BUF1 (N6679, N6657);
nand NAND4 (N6680, N6674, N4159, N1915, N275);
not NOT1 (N6681, N6676);
and AND3 (N6682, N6635, N6640, N6419);
or OR3 (N6683, N6672, N5333, N4348);
nor NOR2 (N6684, N6671, N3564);
or OR2 (N6685, N6680, N4641);
or OR2 (N6686, N6684, N2948);
nand NAND2 (N6687, N6673, N965);
nor NOR4 (N6688, N6679, N355, N3989, N50);
nand NAND4 (N6689, N6688, N3034, N1212, N5296);
or OR4 (N6690, N6681, N6037, N3100, N4805);
buf BUF1 (N6691, N6682);
nand NAND2 (N6692, N6686, N3808);
or OR4 (N6693, N6665, N2559, N2141, N781);
and AND2 (N6694, N6677, N5688);
xor XOR2 (N6695, N6693, N5203);
nand NAND4 (N6696, N6689, N3582, N5450, N3458);
or OR3 (N6697, N6683, N6320, N4441);
xor XOR2 (N6698, N6690, N1472);
or OR4 (N6699, N6695, N3967, N5092, N6455);
buf BUF1 (N6700, N6698);
or OR3 (N6701, N6694, N2119, N4015);
nor NOR2 (N6702, N6678, N6397);
nor NOR2 (N6703, N6696, N2827);
buf BUF1 (N6704, N6685);
nor NOR2 (N6705, N6699, N3958);
or OR4 (N6706, N6691, N467, N1785, N2288);
nor NOR3 (N6707, N6703, N1103, N3586);
or OR4 (N6708, N6692, N5413, N999, N1768);
nor NOR2 (N6709, N6697, N681);
nand NAND3 (N6710, N6700, N2765, N4841);
buf BUF1 (N6711, N6705);
nor NOR2 (N6712, N6704, N5894);
nand NAND3 (N6713, N6702, N1513, N6377);
xor XOR2 (N6714, N6701, N5027);
buf BUF1 (N6715, N6709);
nand NAND4 (N6716, N6707, N6537, N1020, N2070);
buf BUF1 (N6717, N6711);
and AND4 (N6718, N6715, N6526, N1552, N5182);
xor XOR2 (N6719, N6712, N6067);
nand NAND3 (N6720, N6706, N1123, N1262);
nor NOR3 (N6721, N6718, N1140, N3967);
or OR4 (N6722, N6719, N3220, N5179, N3062);
or OR3 (N6723, N6687, N691, N5359);
and AND4 (N6724, N6723, N4591, N2097, N1955);
not NOT1 (N6725, N6717);
buf BUF1 (N6726, N6710);
buf BUF1 (N6727, N6726);
or OR2 (N6728, N6721, N424);
or OR3 (N6729, N6727, N326, N422);
nor NOR2 (N6730, N6724, N4293);
or OR3 (N6731, N6716, N4526, N3790);
and AND3 (N6732, N6731, N2166, N4162);
nor NOR2 (N6733, N6720, N2020);
or OR3 (N6734, N6722, N3488, N5747);
nand NAND4 (N6735, N6732, N3971, N4701, N5712);
and AND3 (N6736, N6730, N858, N3293);
or OR2 (N6737, N6725, N969);
nor NOR4 (N6738, N6714, N1540, N308, N979);
nor NOR4 (N6739, N6708, N6326, N3152, N127);
and AND4 (N6740, N6739, N6196, N1200, N6656);
buf BUF1 (N6741, N6740);
nor NOR3 (N6742, N6741, N1155, N1564);
and AND4 (N6743, N6713, N2816, N6246, N5626);
buf BUF1 (N6744, N6735);
or OR4 (N6745, N6736, N1608, N5166, N594);
nand NAND4 (N6746, N6737, N1402, N3433, N2219);
or OR3 (N6747, N6743, N378, N1838);
nand NAND2 (N6748, N6729, N5090);
nand NAND4 (N6749, N6738, N1407, N3253, N1854);
xor XOR2 (N6750, N6745, N3463);
buf BUF1 (N6751, N6748);
nor NOR2 (N6752, N6733, N5450);
nand NAND2 (N6753, N6752, N3378);
or OR3 (N6754, N6746, N2554, N3489);
xor XOR2 (N6755, N6742, N6048);
not NOT1 (N6756, N6749);
xor XOR2 (N6757, N6747, N3486);
or OR2 (N6758, N6750, N4191);
or OR4 (N6759, N6751, N2078, N4590, N99);
and AND3 (N6760, N6759, N5955, N4094);
nand NAND2 (N6761, N6760, N9);
xor XOR2 (N6762, N6761, N6027);
xor XOR2 (N6763, N6758, N4996);
xor XOR2 (N6764, N6753, N2016);
nand NAND4 (N6765, N6728, N6056, N2784, N4491);
buf BUF1 (N6766, N6765);
or OR2 (N6767, N6762, N226);
not NOT1 (N6768, N6754);
nand NAND2 (N6769, N6755, N5983);
or OR2 (N6770, N6766, N2462);
buf BUF1 (N6771, N6764);
nor NOR4 (N6772, N6769, N2362, N2533, N4923);
or OR2 (N6773, N6767, N3050);
nor NOR2 (N6774, N6770, N6350);
and AND2 (N6775, N6757, N86);
or OR2 (N6776, N6773, N6068);
or OR2 (N6777, N6734, N876);
not NOT1 (N6778, N6772);
or OR2 (N6779, N6771, N1827);
buf BUF1 (N6780, N6778);
buf BUF1 (N6781, N6775);
buf BUF1 (N6782, N6756);
nand NAND4 (N6783, N6780, N1036, N6470, N3614);
xor XOR2 (N6784, N6779, N381);
nand NAND2 (N6785, N6782, N6589);
nand NAND4 (N6786, N6763, N1488, N6137, N149);
xor XOR2 (N6787, N6783, N115);
or OR4 (N6788, N6784, N3563, N1024, N3722);
and AND3 (N6789, N6787, N2998, N2698);
nand NAND3 (N6790, N6788, N1296, N4173);
not NOT1 (N6791, N6768);
and AND3 (N6792, N6781, N6773, N5258);
not NOT1 (N6793, N6776);
xor XOR2 (N6794, N6793, N870);
and AND2 (N6795, N6786, N4746);
not NOT1 (N6796, N6774);
and AND2 (N6797, N6744, N4948);
not NOT1 (N6798, N6777);
nor NOR4 (N6799, N6797, N2109, N582, N5422);
not NOT1 (N6800, N6796);
or OR3 (N6801, N6792, N4088, N4986);
nand NAND3 (N6802, N6795, N4786, N6514);
not NOT1 (N6803, N6794);
buf BUF1 (N6804, N6798);
nor NOR4 (N6805, N6789, N6091, N1514, N5992);
xor XOR2 (N6806, N6799, N5109);
and AND3 (N6807, N6800, N5758, N6252);
nor NOR4 (N6808, N6791, N3394, N3081, N2018);
or OR4 (N6809, N6790, N648, N5430, N131);
nand NAND3 (N6810, N6805, N5604, N4735);
nand NAND4 (N6811, N6803, N4933, N3906, N335);
not NOT1 (N6812, N6801);
nor NOR4 (N6813, N6808, N1174, N1207, N382);
xor XOR2 (N6814, N6809, N3620);
nand NAND4 (N6815, N6804, N2281, N2052, N566);
nor NOR3 (N6816, N6811, N4392, N6593);
buf BUF1 (N6817, N6802);
xor XOR2 (N6818, N6807, N508);
buf BUF1 (N6819, N6785);
not NOT1 (N6820, N6810);
nor NOR2 (N6821, N6813, N1694);
xor XOR2 (N6822, N6817, N6821);
or OR3 (N6823, N608, N1675, N4801);
buf BUF1 (N6824, N6814);
nor NOR2 (N6825, N6822, N1123);
nor NOR3 (N6826, N6815, N2287, N4155);
not NOT1 (N6827, N6819);
and AND2 (N6828, N6818, N3184);
or OR4 (N6829, N6826, N3254, N4723, N5938);
xor XOR2 (N6830, N6827, N5001);
and AND2 (N6831, N6824, N6428);
and AND2 (N6832, N6829, N5776);
nor NOR3 (N6833, N6820, N788, N4195);
nor NOR2 (N6834, N6816, N1833);
and AND2 (N6835, N6834, N828);
nand NAND4 (N6836, N6812, N1201, N3542, N1366);
buf BUF1 (N6837, N6828);
buf BUF1 (N6838, N6833);
and AND3 (N6839, N6832, N5444, N2569);
and AND3 (N6840, N6806, N968, N4267);
or OR3 (N6841, N6835, N1989, N354);
buf BUF1 (N6842, N6836);
nor NOR3 (N6843, N6842, N256, N3242);
and AND4 (N6844, N6825, N1726, N3479, N2671);
not NOT1 (N6845, N6830);
or OR2 (N6846, N6841, N1572);
buf BUF1 (N6847, N6831);
xor XOR2 (N6848, N6843, N6720);
and AND3 (N6849, N6823, N1374, N4534);
or OR2 (N6850, N6837, N3359);
nor NOR2 (N6851, N6844, N4080);
or OR4 (N6852, N6840, N4424, N899, N6663);
nor NOR3 (N6853, N6852, N5666, N5829);
nor NOR3 (N6854, N6847, N3928, N2263);
and AND3 (N6855, N6838, N5728, N2772);
buf BUF1 (N6856, N6855);
nor NOR2 (N6857, N6846, N3177);
buf BUF1 (N6858, N6845);
nor NOR4 (N6859, N6848, N4748, N2135, N5617);
xor XOR2 (N6860, N6853, N4422);
or OR2 (N6861, N6856, N760);
or OR3 (N6862, N6851, N268, N1306);
and AND4 (N6863, N6850, N5841, N3433, N4796);
and AND4 (N6864, N6862, N254, N3175, N4039);
not NOT1 (N6865, N6839);
xor XOR2 (N6866, N6857, N2470);
or OR4 (N6867, N6864, N550, N6812, N216);
buf BUF1 (N6868, N6866);
and AND2 (N6869, N6861, N1290);
or OR3 (N6870, N6849, N4796, N4014);
nor NOR2 (N6871, N6870, N5666);
nand NAND3 (N6872, N6869, N4301, N6832);
nand NAND4 (N6873, N6858, N351, N6237, N6283);
xor XOR2 (N6874, N6854, N6550);
buf BUF1 (N6875, N6872);
xor XOR2 (N6876, N6859, N1629);
buf BUF1 (N6877, N6871);
and AND2 (N6878, N6877, N5757);
and AND2 (N6879, N6860, N1040);
nor NOR3 (N6880, N6867, N1426, N699);
xor XOR2 (N6881, N6863, N5000);
not NOT1 (N6882, N6874);
not NOT1 (N6883, N6876);
and AND3 (N6884, N6865, N3796, N2824);
not NOT1 (N6885, N6878);
nor NOR2 (N6886, N6880, N1506);
not NOT1 (N6887, N6886);
and AND4 (N6888, N6885, N4480, N6518, N6495);
nor NOR4 (N6889, N6888, N1654, N641, N1459);
not NOT1 (N6890, N6883);
nand NAND2 (N6891, N6887, N5082);
or OR3 (N6892, N6891, N4370, N6645);
not NOT1 (N6893, N6868);
or OR3 (N6894, N6881, N338, N601);
nor NOR2 (N6895, N6882, N5422);
not NOT1 (N6896, N6884);
or OR3 (N6897, N6896, N763, N2052);
buf BUF1 (N6898, N6873);
buf BUF1 (N6899, N6889);
or OR2 (N6900, N6898, N594);
xor XOR2 (N6901, N6894, N2716);
xor XOR2 (N6902, N6899, N3526);
and AND3 (N6903, N6893, N1353, N1468);
or OR2 (N6904, N6892, N5179);
not NOT1 (N6905, N6900);
nor NOR4 (N6906, N6905, N925, N4316, N1741);
not NOT1 (N6907, N6895);
not NOT1 (N6908, N6890);
xor XOR2 (N6909, N6902, N2344);
xor XOR2 (N6910, N6908, N6827);
nor NOR4 (N6911, N6904, N4180, N5255, N3420);
nor NOR2 (N6912, N6909, N1855);
not NOT1 (N6913, N6903);
not NOT1 (N6914, N6910);
or OR3 (N6915, N6913, N4434, N5647);
nand NAND3 (N6916, N6906, N4293, N4704);
or OR3 (N6917, N6879, N6258, N3532);
nor NOR2 (N6918, N6912, N6393);
or OR4 (N6919, N6917, N1227, N3013, N3280);
and AND3 (N6920, N6919, N6800, N286);
nand NAND3 (N6921, N6914, N6476, N273);
nor NOR2 (N6922, N6901, N5008);
and AND2 (N6923, N6921, N6880);
not NOT1 (N6924, N6875);
or OR3 (N6925, N6915, N2653, N1816);
xor XOR2 (N6926, N6920, N3606);
nor NOR3 (N6927, N6916, N2969, N2378);
nor NOR3 (N6928, N6897, N1112, N3465);
nor NOR4 (N6929, N6924, N5499, N6113, N2170);
buf BUF1 (N6930, N6923);
buf BUF1 (N6931, N6927);
or OR2 (N6932, N6907, N153);
buf BUF1 (N6933, N6911);
or OR3 (N6934, N6925, N4818, N5230);
not NOT1 (N6935, N6929);
nor NOR4 (N6936, N6933, N3723, N6698, N6450);
xor XOR2 (N6937, N6936, N3428);
or OR4 (N6938, N6928, N4655, N2243, N4245);
nor NOR3 (N6939, N6937, N6469, N2543);
buf BUF1 (N6940, N6935);
nand NAND2 (N6941, N6932, N4376);
not NOT1 (N6942, N6934);
xor XOR2 (N6943, N6930, N6224);
buf BUF1 (N6944, N6931);
xor XOR2 (N6945, N6938, N5312);
buf BUF1 (N6946, N6918);
not NOT1 (N6947, N6926);
xor XOR2 (N6948, N6922, N6696);
or OR2 (N6949, N6939, N1254);
buf BUF1 (N6950, N6945);
buf BUF1 (N6951, N6941);
xor XOR2 (N6952, N6948, N4842);
not NOT1 (N6953, N6946);
xor XOR2 (N6954, N6942, N6885);
buf BUF1 (N6955, N6944);
nor NOR4 (N6956, N6952, N4831, N724, N5075);
and AND3 (N6957, N6954, N6868, N6785);
nor NOR4 (N6958, N6955, N6436, N2545, N2363);
buf BUF1 (N6959, N6957);
nor NOR2 (N6960, N6950, N4458);
not NOT1 (N6961, N6949);
xor XOR2 (N6962, N6958, N470);
or OR4 (N6963, N6959, N4764, N446, N44);
xor XOR2 (N6964, N6956, N950);
nor NOR3 (N6965, N6943, N4452, N2641);
and AND3 (N6966, N6961, N6766, N3902);
nand NAND2 (N6967, N6966, N2410);
buf BUF1 (N6968, N6962);
nand NAND4 (N6969, N6965, N3838, N6856, N1911);
not NOT1 (N6970, N6967);
xor XOR2 (N6971, N6964, N1368);
nand NAND4 (N6972, N6969, N3550, N710, N1443);
and AND3 (N6973, N6947, N1775, N6229);
xor XOR2 (N6974, N6971, N2918);
and AND2 (N6975, N6973, N5049);
xor XOR2 (N6976, N6963, N2728);
xor XOR2 (N6977, N6953, N3885);
buf BUF1 (N6978, N6940);
nand NAND3 (N6979, N6975, N3979, N6);
buf BUF1 (N6980, N6976);
xor XOR2 (N6981, N6951, N2104);
buf BUF1 (N6982, N6980);
and AND3 (N6983, N6977, N3748, N2383);
or OR2 (N6984, N6982, N5636);
and AND4 (N6985, N6960, N1644, N525, N4657);
buf BUF1 (N6986, N6970);
or OR4 (N6987, N6972, N3248, N1058, N1638);
nor NOR3 (N6988, N6983, N2533, N841);
and AND4 (N6989, N6987, N5117, N4351, N6934);
not NOT1 (N6990, N6986);
or OR4 (N6991, N6985, N2919, N6294, N6399);
nor NOR3 (N6992, N6974, N3840, N972);
nor NOR4 (N6993, N6981, N6371, N6335, N359);
not NOT1 (N6994, N6978);
and AND4 (N6995, N6994, N4285, N6205, N2858);
buf BUF1 (N6996, N6993);
nor NOR2 (N6997, N6995, N300);
xor XOR2 (N6998, N6988, N4288);
buf BUF1 (N6999, N6991);
buf BUF1 (N7000, N6997);
not NOT1 (N7001, N6984);
or OR4 (N7002, N6998, N34, N3278, N340);
xor XOR2 (N7003, N6979, N2365);
not NOT1 (N7004, N6968);
or OR2 (N7005, N7002, N1910);
and AND2 (N7006, N6999, N5971);
or OR2 (N7007, N7005, N2478);
and AND4 (N7008, N6989, N85, N4688, N5104);
xor XOR2 (N7009, N7007, N6793);
or OR4 (N7010, N7001, N4019, N1921, N3828);
or OR2 (N7011, N7009, N4426);
not NOT1 (N7012, N7000);
not NOT1 (N7013, N7004);
nand NAND2 (N7014, N7008, N4103);
or OR3 (N7015, N6992, N5074, N6716);
not NOT1 (N7016, N7012);
and AND4 (N7017, N6996, N6497, N5339, N2948);
not NOT1 (N7018, N7011);
and AND4 (N7019, N6990, N4558, N5731, N1547);
xor XOR2 (N7020, N7013, N6895);
not NOT1 (N7021, N7018);
nand NAND3 (N7022, N7003, N145, N5750);
or OR2 (N7023, N7010, N3176);
not NOT1 (N7024, N7015);
xor XOR2 (N7025, N7016, N3547);
and AND2 (N7026, N7014, N3520);
not NOT1 (N7027, N7025);
buf BUF1 (N7028, N7022);
or OR4 (N7029, N7020, N3097, N4120, N163);
and AND2 (N7030, N7019, N403);
not NOT1 (N7031, N7024);
buf BUF1 (N7032, N7023);
nand NAND4 (N7033, N7027, N1213, N2251, N3709);
not NOT1 (N7034, N7030);
or OR4 (N7035, N7028, N4982, N6921, N3525);
buf BUF1 (N7036, N7035);
and AND3 (N7037, N7032, N6479, N2026);
buf BUF1 (N7038, N7021);
nor NOR4 (N7039, N7036, N471, N414, N1110);
nand NAND2 (N7040, N7034, N5081);
not NOT1 (N7041, N7037);
xor XOR2 (N7042, N7006, N2554);
nor NOR4 (N7043, N7042, N7004, N3081, N6615);
not NOT1 (N7044, N7043);
and AND4 (N7045, N7038, N6685, N3907, N6395);
nor NOR4 (N7046, N7033, N3330, N4423, N4674);
not NOT1 (N7047, N7044);
or OR2 (N7048, N7046, N5681);
buf BUF1 (N7049, N7045);
and AND2 (N7050, N7049, N4565);
or OR4 (N7051, N7048, N1168, N451, N270);
nor NOR2 (N7052, N7026, N502);
nor NOR4 (N7053, N7039, N1636, N285, N2436);
not NOT1 (N7054, N7050);
buf BUF1 (N7055, N7029);
nand NAND4 (N7056, N7041, N3100, N6855, N3162);
not NOT1 (N7057, N7056);
nand NAND3 (N7058, N7053, N1041, N5215);
and AND4 (N7059, N7055, N3915, N3632, N3766);
nand NAND4 (N7060, N7052, N637, N824, N6348);
buf BUF1 (N7061, N7059);
nor NOR2 (N7062, N7017, N6505);
not NOT1 (N7063, N7054);
nor NOR4 (N7064, N7060, N2141, N846, N2063);
or OR3 (N7065, N7063, N3395, N870);
nor NOR2 (N7066, N7051, N274);
xor XOR2 (N7067, N7058, N4678);
nand NAND2 (N7068, N7031, N2393);
nand NAND2 (N7069, N7068, N4025);
xor XOR2 (N7070, N7047, N414);
xor XOR2 (N7071, N7069, N2748);
buf BUF1 (N7072, N7064);
nand NAND2 (N7073, N7072, N3479);
and AND4 (N7074, N7062, N4353, N5188, N1662);
xor XOR2 (N7075, N7074, N3230);
nor NOR3 (N7076, N7073, N2940, N4252);
nand NAND2 (N7077, N7057, N6846);
or OR4 (N7078, N7071, N3877, N2092, N6160);
or OR4 (N7079, N7040, N2732, N5267, N1111);
and AND4 (N7080, N7079, N117, N3478, N63);
nand NAND2 (N7081, N7067, N5849);
nand NAND2 (N7082, N7061, N1642);
nand NAND4 (N7083, N7082, N5822, N6935, N5027);
buf BUF1 (N7084, N7065);
and AND4 (N7085, N7076, N6158, N4701, N577);
and AND4 (N7086, N7078, N2600, N3898, N353);
xor XOR2 (N7087, N7083, N5668);
buf BUF1 (N7088, N7070);
or OR3 (N7089, N7077, N4164, N1355);
and AND3 (N7090, N7075, N6072, N1873);
xor XOR2 (N7091, N7084, N379);
nand NAND2 (N7092, N7085, N5627);
not NOT1 (N7093, N7087);
not NOT1 (N7094, N7080);
xor XOR2 (N7095, N7092, N6768);
and AND3 (N7096, N7091, N3521, N2509);
buf BUF1 (N7097, N7086);
or OR4 (N7098, N7095, N5763, N4809, N4002);
or OR4 (N7099, N7094, N4160, N5367, N1035);
and AND4 (N7100, N7099, N3431, N2322, N456);
or OR2 (N7101, N7089, N5774);
nand NAND2 (N7102, N7066, N3004);
and AND4 (N7103, N7093, N4448, N912, N4095);
xor XOR2 (N7104, N7088, N3205);
buf BUF1 (N7105, N7104);
buf BUF1 (N7106, N7096);
and AND2 (N7107, N7097, N2810);
buf BUF1 (N7108, N7103);
buf BUF1 (N7109, N7106);
not NOT1 (N7110, N7107);
xor XOR2 (N7111, N7098, N1279);
not NOT1 (N7112, N7101);
or OR4 (N7113, N7100, N4500, N6910, N2721);
xor XOR2 (N7114, N7112, N554);
or OR2 (N7115, N7102, N1995);
or OR3 (N7116, N7111, N5894, N2478);
nor NOR3 (N7117, N7105, N4445, N4041);
and AND3 (N7118, N7113, N1740, N6590);
nor NOR3 (N7119, N7110, N4225, N966);
and AND3 (N7120, N7090, N3323, N4573);
or OR3 (N7121, N7120, N4470, N1002);
or OR2 (N7122, N7081, N5208);
or OR4 (N7123, N7108, N6496, N6359, N2258);
xor XOR2 (N7124, N7116, N1036);
xor XOR2 (N7125, N7121, N2399);
nand NAND2 (N7126, N7124, N1842);
xor XOR2 (N7127, N7117, N583);
or OR4 (N7128, N7119, N5362, N1545, N4334);
and AND3 (N7129, N7114, N4882, N481);
and AND4 (N7130, N7109, N4054, N2522, N4530);
nand NAND4 (N7131, N7125, N4914, N5714, N4691);
not NOT1 (N7132, N7118);
xor XOR2 (N7133, N7126, N6636);
nor NOR3 (N7134, N7131, N2181, N893);
xor XOR2 (N7135, N7122, N6437);
nand NAND2 (N7136, N7128, N2729);
and AND4 (N7137, N7129, N3771, N5624, N3895);
or OR4 (N7138, N7133, N1725, N2926, N2223);
xor XOR2 (N7139, N7135, N4806);
nor NOR4 (N7140, N7115, N5074, N2277, N2507);
nand NAND2 (N7141, N7137, N6615);
not NOT1 (N7142, N7127);
or OR3 (N7143, N7140, N3170, N6237);
and AND4 (N7144, N7139, N6541, N4092, N5527);
buf BUF1 (N7145, N7132);
buf BUF1 (N7146, N7134);
and AND4 (N7147, N7123, N91, N1911, N546);
nand NAND4 (N7148, N7146, N2113, N3148, N7054);
not NOT1 (N7149, N7147);
or OR3 (N7150, N7142, N3126, N4379);
or OR2 (N7151, N7136, N5225);
nor NOR3 (N7152, N7150, N6133, N1630);
xor XOR2 (N7153, N7148, N4586);
not NOT1 (N7154, N7138);
or OR2 (N7155, N7143, N153);
nor NOR4 (N7156, N7144, N3450, N785, N4460);
or OR4 (N7157, N7156, N7133, N3334, N394);
not NOT1 (N7158, N7157);
buf BUF1 (N7159, N7152);
nand NAND2 (N7160, N7130, N122);
and AND2 (N7161, N7158, N3692);
nand NAND4 (N7162, N7145, N6810, N1576, N1089);
nand NAND4 (N7163, N7161, N4689, N1858, N5772);
nor NOR3 (N7164, N7149, N5686, N6064);
nand NAND3 (N7165, N7160, N1827, N4907);
nand NAND2 (N7166, N7162, N2428);
buf BUF1 (N7167, N7154);
not NOT1 (N7168, N7155);
xor XOR2 (N7169, N7153, N151);
nor NOR2 (N7170, N7159, N3046);
nor NOR2 (N7171, N7151, N5411);
nand NAND4 (N7172, N7165, N5853, N1989, N6441);
nor NOR3 (N7173, N7141, N6055, N3977);
or OR2 (N7174, N7167, N4018);
not NOT1 (N7175, N7170);
not NOT1 (N7176, N7163);
nand NAND4 (N7177, N7176, N1944, N483, N2098);
nand NAND3 (N7178, N7171, N4676, N4962);
buf BUF1 (N7179, N7168);
xor XOR2 (N7180, N7169, N711);
not NOT1 (N7181, N7178);
nand NAND4 (N7182, N7179, N386, N2953, N3571);
buf BUF1 (N7183, N7181);
nor NOR4 (N7184, N7180, N5446, N1291, N6477);
buf BUF1 (N7185, N7182);
xor XOR2 (N7186, N7164, N5025);
or OR4 (N7187, N7184, N181, N902, N5683);
not NOT1 (N7188, N7172);
xor XOR2 (N7189, N7173, N4959);
or OR4 (N7190, N7183, N5355, N5754, N679);
nand NAND4 (N7191, N7185, N665, N2416, N6365);
and AND4 (N7192, N7166, N2974, N5399, N1770);
nand NAND2 (N7193, N7189, N940);
buf BUF1 (N7194, N7191);
not NOT1 (N7195, N7190);
nand NAND3 (N7196, N7193, N6356, N7039);
and AND3 (N7197, N7195, N930, N2602);
nor NOR3 (N7198, N7192, N5996, N4817);
nor NOR4 (N7199, N7194, N3059, N586, N7187);
buf BUF1 (N7200, N3187);
buf BUF1 (N7201, N7198);
and AND4 (N7202, N7175, N279, N6336, N2605);
xor XOR2 (N7203, N7177, N6029);
buf BUF1 (N7204, N7202);
buf BUF1 (N7205, N7203);
buf BUF1 (N7206, N7201);
nand NAND2 (N7207, N7205, N3187);
not NOT1 (N7208, N7199);
or OR4 (N7209, N7200, N794, N4279, N2002);
buf BUF1 (N7210, N7174);
xor XOR2 (N7211, N7209, N772);
nor NOR2 (N7212, N7208, N30);
buf BUF1 (N7213, N7196);
or OR4 (N7214, N7212, N2359, N3828, N1017);
buf BUF1 (N7215, N7214);
nor NOR2 (N7216, N7210, N6357);
and AND3 (N7217, N7216, N3692, N193);
nor NOR3 (N7218, N7206, N5503, N1048);
buf BUF1 (N7219, N7186);
xor XOR2 (N7220, N7218, N4318);
buf BUF1 (N7221, N7220);
xor XOR2 (N7222, N7204, N1573);
or OR2 (N7223, N7188, N4825);
nor NOR2 (N7224, N7222, N6018);
nand NAND2 (N7225, N7219, N6497);
or OR2 (N7226, N7207, N5863);
or OR2 (N7227, N7217, N825);
xor XOR2 (N7228, N7197, N5249);
xor XOR2 (N7229, N7223, N1941);
nand NAND3 (N7230, N7213, N6217, N1347);
not NOT1 (N7231, N7225);
or OR4 (N7232, N7224, N1205, N1377, N5800);
xor XOR2 (N7233, N7215, N1595);
xor XOR2 (N7234, N7221, N3489);
nor NOR4 (N7235, N7226, N1764, N2073, N1412);
buf BUF1 (N7236, N7211);
or OR2 (N7237, N7236, N579);
nor NOR2 (N7238, N7233, N6640);
nor NOR3 (N7239, N7234, N2886, N1504);
not NOT1 (N7240, N7239);
nand NAND4 (N7241, N7238, N4110, N4421, N6703);
nand NAND4 (N7242, N7228, N558, N3900, N3715);
or OR3 (N7243, N7241, N4294, N5730);
xor XOR2 (N7244, N7237, N2619);
or OR4 (N7245, N7231, N6870, N2347, N1212);
nand NAND2 (N7246, N7229, N5624);
nand NAND4 (N7247, N7245, N1496, N3321, N6502);
or OR3 (N7248, N7244, N5973, N5674);
nor NOR4 (N7249, N7235, N3994, N6313, N4516);
xor XOR2 (N7250, N7232, N547);
not NOT1 (N7251, N7248);
and AND2 (N7252, N7227, N6149);
and AND2 (N7253, N7246, N3562);
buf BUF1 (N7254, N7249);
or OR4 (N7255, N7250, N5305, N6076, N6573);
buf BUF1 (N7256, N7230);
nor NOR3 (N7257, N7243, N1173, N2195);
xor XOR2 (N7258, N7240, N1788);
xor XOR2 (N7259, N7242, N1859);
nor NOR2 (N7260, N7256, N5021);
nor NOR4 (N7261, N7257, N945, N3021, N1727);
or OR2 (N7262, N7260, N5664);
nor NOR4 (N7263, N7251, N600, N3409, N1435);
buf BUF1 (N7264, N7258);
not NOT1 (N7265, N7253);
xor XOR2 (N7266, N7265, N6484);
and AND2 (N7267, N7254, N216);
or OR4 (N7268, N7259, N3361, N7231, N4201);
and AND4 (N7269, N7255, N6951, N6434, N966);
buf BUF1 (N7270, N7269);
and AND2 (N7271, N7252, N5705);
and AND2 (N7272, N7268, N4265);
buf BUF1 (N7273, N7270);
buf BUF1 (N7274, N7247);
xor XOR2 (N7275, N7266, N5183);
xor XOR2 (N7276, N7267, N2834);
not NOT1 (N7277, N7271);
xor XOR2 (N7278, N7263, N6889);
and AND2 (N7279, N7275, N677);
nand NAND4 (N7280, N7274, N2904, N7272, N4140);
nor NOR3 (N7281, N6293, N4151, N1787);
buf BUF1 (N7282, N7276);
nand NAND3 (N7283, N7277, N3909, N257);
nand NAND2 (N7284, N7281, N4494);
and AND2 (N7285, N7261, N3004);
buf BUF1 (N7286, N7283);
and AND2 (N7287, N7285, N6897);
nor NOR2 (N7288, N7278, N7164);
xor XOR2 (N7289, N7262, N3714);
xor XOR2 (N7290, N7288, N2427);
nand NAND4 (N7291, N7279, N6348, N321, N5101);
or OR4 (N7292, N7291, N5564, N425, N5904);
nor NOR3 (N7293, N7287, N7067, N6893);
nand NAND4 (N7294, N7282, N2145, N5831, N4927);
and AND4 (N7295, N7273, N4197, N3364, N1131);
buf BUF1 (N7296, N7280);
nand NAND2 (N7297, N7264, N93);
or OR4 (N7298, N7295, N6200, N2463, N1079);
not NOT1 (N7299, N7284);
nand NAND4 (N7300, N7299, N1691, N212, N4095);
nand NAND4 (N7301, N7289, N6056, N7172, N3481);
and AND2 (N7302, N7301, N628);
buf BUF1 (N7303, N7298);
buf BUF1 (N7304, N7294);
and AND4 (N7305, N7297, N1240, N7196, N962);
xor XOR2 (N7306, N7300, N3806);
buf BUF1 (N7307, N7296);
and AND4 (N7308, N7290, N1450, N6869, N1839);
nand NAND4 (N7309, N7286, N2837, N1503, N2517);
buf BUF1 (N7310, N7304);
buf BUF1 (N7311, N7309);
xor XOR2 (N7312, N7302, N5470);
nor NOR2 (N7313, N7310, N6002);
xor XOR2 (N7314, N7292, N5240);
and AND3 (N7315, N7313, N4662, N3200);
buf BUF1 (N7316, N7315);
or OR2 (N7317, N7305, N627);
nand NAND4 (N7318, N7311, N4379, N121, N689);
buf BUF1 (N7319, N7293);
or OR4 (N7320, N7317, N1465, N2397, N2786);
and AND3 (N7321, N7308, N7255, N4614);
nand NAND4 (N7322, N7314, N6504, N1784, N6109);
and AND4 (N7323, N7321, N6016, N5296, N3623);
nand NAND3 (N7324, N7319, N6888, N5968);
not NOT1 (N7325, N7316);
not NOT1 (N7326, N7323);
nor NOR3 (N7327, N7325, N1385, N3662);
and AND3 (N7328, N7318, N3027, N3601);
or OR3 (N7329, N7324, N4511, N6085);
nand NAND4 (N7330, N7303, N1145, N2698, N4730);
or OR4 (N7331, N7330, N2239, N1957, N6316);
or OR2 (N7332, N7331, N2799);
not NOT1 (N7333, N7320);
or OR3 (N7334, N7329, N4621, N989);
or OR3 (N7335, N7328, N4187, N3234);
nor NOR3 (N7336, N7333, N856, N2093);
or OR2 (N7337, N7327, N2030);
not NOT1 (N7338, N7336);
and AND2 (N7339, N7334, N6900);
nor NOR2 (N7340, N7337, N6599);
and AND2 (N7341, N7338, N4348);
and AND2 (N7342, N7332, N5528);
nand NAND3 (N7343, N7307, N5047, N4597);
not NOT1 (N7344, N7343);
and AND3 (N7345, N7322, N6652, N368);
nor NOR2 (N7346, N7335, N644);
not NOT1 (N7347, N7341);
nand NAND2 (N7348, N7347, N4102);
xor XOR2 (N7349, N7346, N3470);
buf BUF1 (N7350, N7344);
and AND4 (N7351, N7345, N5197, N5367, N1138);
or OR3 (N7352, N7340, N5018, N2619);
nor NOR4 (N7353, N7339, N963, N5964, N2708);
nor NOR3 (N7354, N7306, N3454, N7245);
not NOT1 (N7355, N7312);
nand NAND4 (N7356, N7349, N54, N2104, N1041);
not NOT1 (N7357, N7348);
not NOT1 (N7358, N7351);
nand NAND3 (N7359, N7354, N356, N544);
or OR2 (N7360, N7356, N710);
nor NOR2 (N7361, N7360, N7359);
buf BUF1 (N7362, N3851);
or OR3 (N7363, N7358, N2209, N5336);
nor NOR3 (N7364, N7355, N559, N4097);
not NOT1 (N7365, N7342);
nand NAND4 (N7366, N7353, N1120, N5267, N4564);
not NOT1 (N7367, N7326);
nand NAND3 (N7368, N7357, N3021, N3118);
buf BUF1 (N7369, N7352);
xor XOR2 (N7370, N7350, N4438);
or OR3 (N7371, N7361, N3661, N6947);
nand NAND2 (N7372, N7371, N1238);
not NOT1 (N7373, N7370);
not NOT1 (N7374, N7367);
not NOT1 (N7375, N7365);
xor XOR2 (N7376, N7363, N1909);
nand NAND3 (N7377, N7366, N5671, N1429);
buf BUF1 (N7378, N7362);
buf BUF1 (N7379, N7376);
not NOT1 (N7380, N7372);
buf BUF1 (N7381, N7368);
and AND4 (N7382, N7380, N4068, N6348, N418);
xor XOR2 (N7383, N7375, N6338);
buf BUF1 (N7384, N7381);
xor XOR2 (N7385, N7374, N804);
nand NAND4 (N7386, N7369, N7032, N5856, N93);
not NOT1 (N7387, N7384);
xor XOR2 (N7388, N7379, N5040);
xor XOR2 (N7389, N7383, N4256);
buf BUF1 (N7390, N7378);
and AND3 (N7391, N7389, N932, N5775);
or OR4 (N7392, N7386, N1214, N6715, N335);
not NOT1 (N7393, N7391);
xor XOR2 (N7394, N7392, N2156);
buf BUF1 (N7395, N7385);
and AND3 (N7396, N7364, N7344, N6392);
or OR4 (N7397, N7396, N5615, N3532, N5368);
nand NAND4 (N7398, N7394, N1909, N4922, N4311);
xor XOR2 (N7399, N7387, N2372);
or OR3 (N7400, N7397, N3365, N6233);
nand NAND3 (N7401, N7393, N246, N2839);
buf BUF1 (N7402, N7373);
or OR2 (N7403, N7390, N1378);
xor XOR2 (N7404, N7395, N5526);
or OR3 (N7405, N7382, N3198, N1804);
xor XOR2 (N7406, N7401, N557);
or OR4 (N7407, N7377, N103, N6543, N5478);
nand NAND4 (N7408, N7399, N1092, N6714, N5875);
buf BUF1 (N7409, N7405);
or OR2 (N7410, N7398, N5598);
xor XOR2 (N7411, N7410, N6611);
or OR3 (N7412, N7403, N3698, N638);
and AND3 (N7413, N7407, N6240, N3434);
not NOT1 (N7414, N7388);
not NOT1 (N7415, N7413);
xor XOR2 (N7416, N7411, N758);
and AND4 (N7417, N7415, N1782, N5952, N219);
or OR2 (N7418, N7417, N2404);
or OR3 (N7419, N7404, N7053, N5189);
not NOT1 (N7420, N7409);
and AND3 (N7421, N7400, N6659, N5607);
and AND3 (N7422, N7418, N7135, N690);
nor NOR2 (N7423, N7421, N1542);
xor XOR2 (N7424, N7422, N927);
xor XOR2 (N7425, N7406, N7019);
and AND4 (N7426, N7416, N4410, N6197, N7314);
not NOT1 (N7427, N7408);
buf BUF1 (N7428, N7424);
buf BUF1 (N7429, N7425);
xor XOR2 (N7430, N7423, N3196);
and AND4 (N7431, N7428, N2251, N1413, N4400);
buf BUF1 (N7432, N7427);
nand NAND4 (N7433, N7402, N3706, N1256, N1072);
nor NOR4 (N7434, N7414, N229, N4241, N2256);
nand NAND4 (N7435, N7433, N1032, N4485, N3999);
nor NOR3 (N7436, N7430, N2267, N5920);
xor XOR2 (N7437, N7436, N3521);
xor XOR2 (N7438, N7431, N1904);
or OR4 (N7439, N7438, N7206, N3027, N5982);
nand NAND4 (N7440, N7439, N479, N4969, N188);
and AND3 (N7441, N7435, N1371, N5065);
not NOT1 (N7442, N7437);
buf BUF1 (N7443, N7429);
nand NAND3 (N7444, N7412, N6982, N2527);
not NOT1 (N7445, N7432);
or OR2 (N7446, N7443, N1468);
or OR4 (N7447, N7419, N5728, N146, N913);
not NOT1 (N7448, N7440);
xor XOR2 (N7449, N7426, N5725);
or OR4 (N7450, N7434, N3321, N5427, N4937);
and AND3 (N7451, N7446, N5727, N3078);
buf BUF1 (N7452, N7441);
not NOT1 (N7453, N7449);
and AND3 (N7454, N7442, N6400, N3038);
xor XOR2 (N7455, N7447, N6518);
xor XOR2 (N7456, N7450, N666);
not NOT1 (N7457, N7445);
xor XOR2 (N7458, N7452, N572);
nand NAND2 (N7459, N7451, N4895);
not NOT1 (N7460, N7448);
and AND3 (N7461, N7420, N915, N332);
and AND3 (N7462, N7461, N4786, N5984);
xor XOR2 (N7463, N7457, N2564);
or OR4 (N7464, N7463, N4825, N1799, N1548);
not NOT1 (N7465, N7458);
not NOT1 (N7466, N7460);
or OR3 (N7467, N7456, N609, N5207);
or OR2 (N7468, N7465, N968);
buf BUF1 (N7469, N7453);
buf BUF1 (N7470, N7469);
nand NAND3 (N7471, N7466, N1558, N2341);
nor NOR2 (N7472, N7462, N4204);
buf BUF1 (N7473, N7471);
buf BUF1 (N7474, N7473);
xor XOR2 (N7475, N7444, N3344);
and AND3 (N7476, N7470, N1478, N1318);
or OR4 (N7477, N7472, N5598, N2810, N4463);
nor NOR2 (N7478, N7459, N293);
buf BUF1 (N7479, N7477);
xor XOR2 (N7480, N7464, N54);
not NOT1 (N7481, N7480);
buf BUF1 (N7482, N7454);
or OR3 (N7483, N7476, N373, N6374);
and AND3 (N7484, N7478, N2218, N2538);
and AND2 (N7485, N7474, N6774);
xor XOR2 (N7486, N7467, N5490);
nor NOR4 (N7487, N7479, N3872, N809, N1241);
or OR4 (N7488, N7481, N1307, N2302, N6001);
or OR4 (N7489, N7475, N2910, N751, N6351);
nor NOR3 (N7490, N7485, N388, N3843);
and AND4 (N7491, N7483, N5505, N5767, N3217);
or OR4 (N7492, N7490, N427, N2561, N463);
nor NOR3 (N7493, N7484, N1465, N6140);
nand NAND4 (N7494, N7482, N2563, N1879, N4190);
nor NOR3 (N7495, N7489, N4106, N6681);
or OR4 (N7496, N7486, N1229, N6059, N550);
not NOT1 (N7497, N7492);
not NOT1 (N7498, N7495);
xor XOR2 (N7499, N7468, N615);
not NOT1 (N7500, N7488);
xor XOR2 (N7501, N7499, N6919);
nor NOR2 (N7502, N7496, N2993);
or OR4 (N7503, N7498, N6693, N5276, N2871);
xor XOR2 (N7504, N7494, N1007);
buf BUF1 (N7505, N7504);
nor NOR2 (N7506, N7493, N6654);
buf BUF1 (N7507, N7455);
xor XOR2 (N7508, N7502, N4688);
nor NOR3 (N7509, N7505, N1700, N4382);
buf BUF1 (N7510, N7487);
nor NOR2 (N7511, N7503, N5857);
not NOT1 (N7512, N7497);
or OR2 (N7513, N7507, N5900);
not NOT1 (N7514, N7500);
xor XOR2 (N7515, N7509, N5970);
nand NAND2 (N7516, N7511, N3767);
not NOT1 (N7517, N7516);
and AND3 (N7518, N7513, N6504, N6954);
not NOT1 (N7519, N7506);
and AND3 (N7520, N7508, N7157, N6770);
not NOT1 (N7521, N7501);
not NOT1 (N7522, N7521);
nor NOR3 (N7523, N7520, N5050, N7063);
nor NOR2 (N7524, N7517, N6349);
and AND3 (N7525, N7515, N3568, N6422);
xor XOR2 (N7526, N7491, N7173);
and AND3 (N7527, N7524, N1829, N6400);
buf BUF1 (N7528, N7525);
buf BUF1 (N7529, N7527);
not NOT1 (N7530, N7522);
xor XOR2 (N7531, N7510, N1485);
buf BUF1 (N7532, N7514);
not NOT1 (N7533, N7528);
or OR3 (N7534, N7523, N1005, N1286);
and AND3 (N7535, N7532, N7499, N2297);
nand NAND3 (N7536, N7512, N6347, N7097);
not NOT1 (N7537, N7534);
nand NAND4 (N7538, N7533, N6523, N787, N4063);
xor XOR2 (N7539, N7537, N3026);
or OR3 (N7540, N7519, N6829, N5787);
nor NOR2 (N7541, N7539, N5553);
nand NAND3 (N7542, N7541, N2487, N2768);
and AND3 (N7543, N7529, N2289, N4118);
buf BUF1 (N7544, N7526);
nor NOR2 (N7545, N7518, N141);
or OR2 (N7546, N7545, N6507);
buf BUF1 (N7547, N7531);
nand NAND2 (N7548, N7543, N159);
xor XOR2 (N7549, N7535, N4376);
buf BUF1 (N7550, N7538);
xor XOR2 (N7551, N7546, N105);
xor XOR2 (N7552, N7542, N3788);
nand NAND3 (N7553, N7547, N2317, N6616);
and AND4 (N7554, N7540, N1334, N3809, N5722);
nor NOR3 (N7555, N7552, N1067, N360);
buf BUF1 (N7556, N7544);
and AND2 (N7557, N7551, N2753);
nand NAND3 (N7558, N7548, N2232, N902);
nor NOR2 (N7559, N7555, N1047);
not NOT1 (N7560, N7559);
nor NOR4 (N7561, N7553, N2273, N1603, N3054);
or OR3 (N7562, N7550, N1355, N2318);
or OR2 (N7563, N7562, N5228);
or OR4 (N7564, N7554, N3432, N4962, N5139);
and AND3 (N7565, N7563, N7003, N5240);
and AND4 (N7566, N7556, N5436, N5637, N5319);
buf BUF1 (N7567, N7549);
or OR4 (N7568, N7564, N5627, N3920, N7283);
buf BUF1 (N7569, N7566);
xor XOR2 (N7570, N7565, N4261);
nand NAND3 (N7571, N7530, N3638, N1900);
or OR2 (N7572, N7571, N5182);
not NOT1 (N7573, N7560);
nand NAND3 (N7574, N7567, N1355, N1943);
buf BUF1 (N7575, N7536);
xor XOR2 (N7576, N7573, N157);
or OR2 (N7577, N7570, N4762);
or OR4 (N7578, N7561, N3573, N2306, N1727);
buf BUF1 (N7579, N7568);
and AND2 (N7580, N7576, N4181);
not NOT1 (N7581, N7569);
nand NAND2 (N7582, N7577, N7536);
not NOT1 (N7583, N7579);
nand NAND4 (N7584, N7583, N1785, N7446, N571);
buf BUF1 (N7585, N7580);
nor NOR4 (N7586, N7575, N2401, N2444, N6840);
nand NAND3 (N7587, N7578, N5523, N1993);
not NOT1 (N7588, N7585);
buf BUF1 (N7589, N7588);
not NOT1 (N7590, N7586);
not NOT1 (N7591, N7581);
nand NAND4 (N7592, N7582, N2335, N1675, N4039);
buf BUF1 (N7593, N7557);
nor NOR4 (N7594, N7592, N2573, N5488, N1689);
or OR4 (N7595, N7593, N195, N581, N2476);
and AND4 (N7596, N7574, N4563, N4751, N450);
and AND4 (N7597, N7595, N6681, N1791, N7008);
and AND3 (N7598, N7590, N6416, N231);
or OR3 (N7599, N7572, N6106, N5160);
buf BUF1 (N7600, N7598);
and AND2 (N7601, N7597, N4674);
nor NOR4 (N7602, N7589, N929, N651, N2328);
not NOT1 (N7603, N7601);
nand NAND4 (N7604, N7594, N6944, N6097, N7198);
buf BUF1 (N7605, N7596);
xor XOR2 (N7606, N7584, N7562);
nand NAND4 (N7607, N7603, N2253, N660, N3066);
buf BUF1 (N7608, N7558);
not NOT1 (N7609, N7606);
xor XOR2 (N7610, N7607, N6305);
nor NOR2 (N7611, N7608, N746);
nor NOR2 (N7612, N7600, N6675);
or OR2 (N7613, N7611, N5869);
or OR4 (N7614, N7605, N7563, N4460, N1409);
and AND4 (N7615, N7587, N2683, N720, N345);
or OR3 (N7616, N7602, N2673, N4517);
nand NAND3 (N7617, N7613, N1433, N1593);
or OR3 (N7618, N7599, N1194, N6179);
buf BUF1 (N7619, N7612);
nor NOR2 (N7620, N7604, N978);
and AND2 (N7621, N7591, N3871);
or OR2 (N7622, N7621, N4103);
not NOT1 (N7623, N7609);
or OR4 (N7624, N7614, N6618, N676, N3605);
buf BUF1 (N7625, N7623);
xor XOR2 (N7626, N7610, N5444);
nor NOR3 (N7627, N7622, N4087, N4617);
buf BUF1 (N7628, N7627);
or OR4 (N7629, N7616, N512, N6299, N7421);
xor XOR2 (N7630, N7629, N2899);
nand NAND4 (N7631, N7630, N6692, N5613, N2217);
xor XOR2 (N7632, N7625, N6237);
or OR3 (N7633, N7626, N6235, N3731);
not NOT1 (N7634, N7628);
not NOT1 (N7635, N7620);
nand NAND3 (N7636, N7631, N1653, N5479);
buf BUF1 (N7637, N7633);
buf BUF1 (N7638, N7636);
nor NOR2 (N7639, N7619, N1445);
nand NAND2 (N7640, N7618, N88);
and AND3 (N7641, N7640, N3250, N1744);
xor XOR2 (N7642, N7638, N6329);
nor NOR4 (N7643, N7634, N5060, N5866, N7315);
and AND4 (N7644, N7615, N942, N3891, N2563);
buf BUF1 (N7645, N7644);
nor NOR4 (N7646, N7643, N1808, N3001, N1028);
or OR2 (N7647, N7617, N6586);
nand NAND2 (N7648, N7647, N3076);
not NOT1 (N7649, N7641);
xor XOR2 (N7650, N7635, N6361);
or OR2 (N7651, N7639, N4613);
and AND2 (N7652, N7650, N6345);
xor XOR2 (N7653, N7637, N5959);
xor XOR2 (N7654, N7645, N1615);
buf BUF1 (N7655, N7648);
nand NAND4 (N7656, N7624, N738, N6270, N3790);
xor XOR2 (N7657, N7632, N6000);
not NOT1 (N7658, N7652);
nand NAND4 (N7659, N7642, N1264, N1576, N5982);
nor NOR2 (N7660, N7649, N6515);
or OR3 (N7661, N7656, N5997, N2454);
nand NAND3 (N7662, N7653, N3800, N7281);
xor XOR2 (N7663, N7658, N6935);
and AND2 (N7664, N7662, N5334);
or OR3 (N7665, N7661, N6935, N4058);
or OR2 (N7666, N7665, N4274);
and AND2 (N7667, N7663, N896);
nand NAND4 (N7668, N7664, N3935, N1679, N130);
xor XOR2 (N7669, N7654, N350);
or OR2 (N7670, N7657, N5868);
or OR3 (N7671, N7670, N5689, N6480);
buf BUF1 (N7672, N7667);
buf BUF1 (N7673, N7651);
and AND4 (N7674, N7673, N3579, N3436, N4528);
xor XOR2 (N7675, N7668, N2913);
and AND3 (N7676, N7646, N4984, N6359);
xor XOR2 (N7677, N7655, N2785);
nand NAND2 (N7678, N7666, N5154);
xor XOR2 (N7679, N7677, N227);
nor NOR2 (N7680, N7672, N1729);
or OR4 (N7681, N7675, N4670, N5162, N1219);
or OR3 (N7682, N7669, N3406, N231);
or OR4 (N7683, N7660, N1427, N5378, N4432);
buf BUF1 (N7684, N7678);
xor XOR2 (N7685, N7681, N7621);
xor XOR2 (N7686, N7684, N7591);
nor NOR3 (N7687, N7686, N5891, N3746);
and AND2 (N7688, N7671, N724);
not NOT1 (N7689, N7683);
xor XOR2 (N7690, N7680, N191);
xor XOR2 (N7691, N7659, N158);
not NOT1 (N7692, N7676);
not NOT1 (N7693, N7688);
nand NAND3 (N7694, N7692, N3102, N4976);
not NOT1 (N7695, N7693);
not NOT1 (N7696, N7679);
nor NOR4 (N7697, N7691, N4858, N6736, N6568);
xor XOR2 (N7698, N7695, N987);
and AND2 (N7699, N7698, N6855);
buf BUF1 (N7700, N7674);
or OR2 (N7701, N7700, N1564);
or OR4 (N7702, N7696, N5115, N2591, N2005);
or OR2 (N7703, N7701, N2308);
xor XOR2 (N7704, N7703, N7261);
nor NOR4 (N7705, N7689, N3256, N214, N6631);
nor NOR3 (N7706, N7690, N181, N6624);
xor XOR2 (N7707, N7706, N7497);
buf BUF1 (N7708, N7697);
nor NOR4 (N7709, N7702, N6671, N5326, N6320);
nor NOR4 (N7710, N7708, N5039, N1598, N6603);
xor XOR2 (N7711, N7699, N4302);
nand NAND4 (N7712, N7704, N7486, N4606, N4115);
or OR4 (N7713, N7710, N7180, N5586, N1032);
and AND3 (N7714, N7687, N1602, N6454);
nor NOR2 (N7715, N7714, N5929);
or OR2 (N7716, N7705, N893);
nor NOR3 (N7717, N7712, N5234, N4697);
or OR3 (N7718, N7682, N343, N2389);
buf BUF1 (N7719, N7718);
nor NOR2 (N7720, N7715, N910);
not NOT1 (N7721, N7713);
and AND2 (N7722, N7721, N5651);
or OR4 (N7723, N7707, N6615, N1026, N2161);
and AND3 (N7724, N7709, N5626, N6044);
xor XOR2 (N7725, N7719, N332);
xor XOR2 (N7726, N7722, N5710);
nand NAND3 (N7727, N7717, N5145, N3234);
xor XOR2 (N7728, N7720, N1859);
buf BUF1 (N7729, N7725);
and AND2 (N7730, N7694, N7690);
and AND4 (N7731, N7724, N2268, N66, N1606);
nand NAND2 (N7732, N7731, N5404);
or OR3 (N7733, N7727, N4138, N268);
nand NAND2 (N7734, N7729, N4098);
xor XOR2 (N7735, N7716, N4629);
xor XOR2 (N7736, N7733, N2986);
or OR4 (N7737, N7732, N5128, N1663, N1685);
and AND2 (N7738, N7734, N2061);
not NOT1 (N7739, N7723);
xor XOR2 (N7740, N7685, N7147);
buf BUF1 (N7741, N7711);
nor NOR2 (N7742, N7735, N76);
nand NAND2 (N7743, N7742, N6316);
nand NAND3 (N7744, N7740, N4296, N2159);
or OR3 (N7745, N7743, N2129, N2036);
and AND4 (N7746, N7739, N1491, N7099, N3824);
or OR2 (N7747, N7741, N2685);
or OR2 (N7748, N7746, N7240);
not NOT1 (N7749, N7728);
or OR2 (N7750, N7736, N1209);
and AND4 (N7751, N7726, N4416, N1199, N4844);
nand NAND3 (N7752, N7738, N2723, N2601);
nand NAND2 (N7753, N7751, N7337);
nand NAND2 (N7754, N7752, N6167);
or OR4 (N7755, N7750, N1023, N3951, N1300);
nor NOR3 (N7756, N7745, N4048, N4275);
not NOT1 (N7757, N7748);
buf BUF1 (N7758, N7754);
xor XOR2 (N7759, N7755, N7393);
nor NOR2 (N7760, N7753, N6742);
buf BUF1 (N7761, N7758);
not NOT1 (N7762, N7747);
nor NOR4 (N7763, N7749, N5176, N6067, N5965);
nand NAND2 (N7764, N7757, N6811);
or OR4 (N7765, N7763, N1807, N5622, N3588);
buf BUF1 (N7766, N7760);
or OR2 (N7767, N7744, N873);
xor XOR2 (N7768, N7756, N5646);
nor NOR4 (N7769, N7766, N194, N2162, N1304);
nand NAND4 (N7770, N7730, N2389, N1317, N1540);
nand NAND2 (N7771, N7765, N7249);
xor XOR2 (N7772, N7771, N3338);
xor XOR2 (N7773, N7764, N7190);
buf BUF1 (N7774, N7768);
xor XOR2 (N7775, N7762, N7369);
nand NAND2 (N7776, N7770, N4547);
nor NOR4 (N7777, N7737, N4435, N994, N4624);
or OR3 (N7778, N7769, N3523, N3254);
and AND4 (N7779, N7777, N3228, N1678, N7664);
xor XOR2 (N7780, N7775, N2495);
nor NOR2 (N7781, N7779, N7121);
xor XOR2 (N7782, N7774, N651);
and AND2 (N7783, N7767, N2541);
and AND4 (N7784, N7761, N4306, N1513, N4346);
or OR4 (N7785, N7759, N1831, N6690, N1113);
nor NOR3 (N7786, N7780, N7285, N7710);
nor NOR2 (N7787, N7772, N2074);
nor NOR4 (N7788, N7782, N1453, N3078, N5069);
buf BUF1 (N7789, N7784);
or OR3 (N7790, N7788, N929, N6752);
not NOT1 (N7791, N7789);
xor XOR2 (N7792, N7773, N6788);
and AND4 (N7793, N7787, N2783, N3319, N1598);
nand NAND2 (N7794, N7778, N2375);
buf BUF1 (N7795, N7792);
nand NAND4 (N7796, N7791, N1721, N6203, N7646);
xor XOR2 (N7797, N7794, N4319);
nand NAND2 (N7798, N7796, N1576);
nand NAND4 (N7799, N7790, N1048, N1617, N5897);
buf BUF1 (N7800, N7799);
and AND2 (N7801, N7781, N5055);
and AND2 (N7802, N7786, N5343);
not NOT1 (N7803, N7776);
nor NOR4 (N7804, N7798, N5008, N7075, N5846);
xor XOR2 (N7805, N7797, N3419);
xor XOR2 (N7806, N7795, N4990);
nand NAND4 (N7807, N7801, N4230, N686, N7164);
buf BUF1 (N7808, N7805);
buf BUF1 (N7809, N7802);
not NOT1 (N7810, N7809);
not NOT1 (N7811, N7806);
nor NOR4 (N7812, N7803, N5323, N2405, N3102);
buf BUF1 (N7813, N7800);
nor NOR3 (N7814, N7785, N4705, N7683);
xor XOR2 (N7815, N7804, N1312);
buf BUF1 (N7816, N7783);
buf BUF1 (N7817, N7808);
xor XOR2 (N7818, N7811, N3930);
buf BUF1 (N7819, N7793);
buf BUF1 (N7820, N7817);
and AND3 (N7821, N7819, N4404, N3380);
xor XOR2 (N7822, N7814, N1865);
and AND4 (N7823, N7821, N881, N4470, N3044);
buf BUF1 (N7824, N7812);
buf BUF1 (N7825, N7810);
or OR2 (N7826, N7824, N1437);
and AND4 (N7827, N7816, N1867, N5634, N1303);
not NOT1 (N7828, N7815);
buf BUF1 (N7829, N7820);
nor NOR4 (N7830, N7827, N5187, N4204, N726);
nor NOR4 (N7831, N7825, N2747, N822, N2691);
nor NOR4 (N7832, N7826, N6979, N3557, N2768);
nand NAND2 (N7833, N7807, N7328);
buf BUF1 (N7834, N7813);
not NOT1 (N7835, N7818);
xor XOR2 (N7836, N7831, N5526);
and AND3 (N7837, N7836, N578, N410);
nand NAND4 (N7838, N7829, N1762, N2936, N2829);
and AND4 (N7839, N7834, N813, N3675, N348);
nand NAND4 (N7840, N7830, N4076, N4026, N323);
nor NOR2 (N7841, N7837, N2673);
nand NAND3 (N7842, N7840, N3942, N3474);
nand NAND2 (N7843, N7838, N5072);
nand NAND3 (N7844, N7841, N2752, N2443);
nand NAND3 (N7845, N7828, N2420, N4699);
and AND2 (N7846, N7822, N6232);
not NOT1 (N7847, N7839);
nor NOR2 (N7848, N7846, N5129);
nor NOR3 (N7849, N7848, N1077, N1636);
nand NAND3 (N7850, N7845, N7767, N1489);
nor NOR4 (N7851, N7835, N170, N3113, N3323);
xor XOR2 (N7852, N7844, N737);
nor NOR2 (N7853, N7832, N2815);
or OR3 (N7854, N7849, N6198, N2927);
not NOT1 (N7855, N7847);
and AND3 (N7856, N7833, N615, N1723);
not NOT1 (N7857, N7854);
nand NAND3 (N7858, N7857, N2693, N5002);
or OR2 (N7859, N7855, N7326);
nor NOR3 (N7860, N7859, N5867, N1230);
or OR3 (N7861, N7860, N2572, N2737);
and AND2 (N7862, N7853, N1599);
or OR3 (N7863, N7851, N4314, N3850);
not NOT1 (N7864, N7862);
xor XOR2 (N7865, N7856, N2363);
and AND2 (N7866, N7861, N2135);
not NOT1 (N7867, N7864);
or OR3 (N7868, N7858, N4647, N5806);
buf BUF1 (N7869, N7852);
xor XOR2 (N7870, N7867, N6725);
buf BUF1 (N7871, N7868);
nor NOR2 (N7872, N7843, N2686);
and AND3 (N7873, N7869, N6314, N7688);
buf BUF1 (N7874, N7873);
buf BUF1 (N7875, N7872);
and AND3 (N7876, N7865, N3285, N5308);
nor NOR4 (N7877, N7842, N778, N3080, N3208);
not NOT1 (N7878, N7870);
nor NOR4 (N7879, N7878, N2103, N163, N2521);
nor NOR3 (N7880, N7877, N5020, N3378);
not NOT1 (N7881, N7866);
nand NAND2 (N7882, N7879, N2228);
xor XOR2 (N7883, N7871, N7084);
or OR2 (N7884, N7863, N338);
xor XOR2 (N7885, N7883, N1017);
nor NOR3 (N7886, N7884, N7681, N7148);
buf BUF1 (N7887, N7886);
xor XOR2 (N7888, N7875, N1464);
nor NOR2 (N7889, N7880, N2221);
or OR3 (N7890, N7888, N7102, N1897);
buf BUF1 (N7891, N7881);
nor NOR2 (N7892, N7891, N6421);
nand NAND4 (N7893, N7874, N1835, N1269, N3383);
or OR2 (N7894, N7893, N7166);
nand NAND3 (N7895, N7890, N4796, N5422);
nor NOR3 (N7896, N7876, N7271, N6723);
buf BUF1 (N7897, N7882);
xor XOR2 (N7898, N7887, N5379);
buf BUF1 (N7899, N7823);
or OR3 (N7900, N7894, N3793, N5723);
and AND4 (N7901, N7895, N4831, N616, N5418);
nand NAND4 (N7902, N7885, N253, N4239, N7822);
and AND3 (N7903, N7901, N3602, N7417);
or OR4 (N7904, N7896, N406, N7881, N4593);
and AND2 (N7905, N7897, N7359);
nand NAND2 (N7906, N7902, N3890);
xor XOR2 (N7907, N7905, N2953);
and AND4 (N7908, N7907, N5549, N3475, N6333);
buf BUF1 (N7909, N7892);
and AND2 (N7910, N7906, N4852);
nand NAND2 (N7911, N7903, N5616);
xor XOR2 (N7912, N7850, N1640);
and AND4 (N7913, N7912, N4252, N7767, N2375);
xor XOR2 (N7914, N7904, N7451);
nand NAND3 (N7915, N7909, N6532, N1757);
and AND3 (N7916, N7915, N6842, N3604);
nand NAND2 (N7917, N7911, N6032);
nor NOR4 (N7918, N7916, N868, N4579, N7289);
nor NOR2 (N7919, N7913, N1969);
and AND2 (N7920, N7908, N2914);
and AND4 (N7921, N7917, N5309, N6679, N1049);
or OR4 (N7922, N7889, N7459, N272, N1511);
not NOT1 (N7923, N7919);
not NOT1 (N7924, N7922);
and AND3 (N7925, N7920, N5554, N7691);
not NOT1 (N7926, N7921);
nand NAND3 (N7927, N7925, N481, N2020);
nand NAND4 (N7928, N7900, N4494, N7659, N2181);
buf BUF1 (N7929, N7926);
nand NAND2 (N7930, N7898, N4517);
xor XOR2 (N7931, N7918, N7286);
nand NAND3 (N7932, N7914, N2756, N4730);
nor NOR3 (N7933, N7931, N603, N5588);
nor NOR3 (N7934, N7910, N2690, N2298);
and AND3 (N7935, N7899, N4036, N7734);
not NOT1 (N7936, N7924);
not NOT1 (N7937, N7936);
not NOT1 (N7938, N7929);
buf BUF1 (N7939, N7923);
nand NAND3 (N7940, N7927, N716, N4891);
nand NAND3 (N7941, N7928, N2436, N1410);
xor XOR2 (N7942, N7932, N6016);
nand NAND3 (N7943, N7941, N6249, N2879);
nand NAND3 (N7944, N7939, N7233, N5960);
and AND3 (N7945, N7938, N1972, N575);
not NOT1 (N7946, N7930);
not NOT1 (N7947, N7935);
buf BUF1 (N7948, N7945);
nand NAND2 (N7949, N7948, N1238);
not NOT1 (N7950, N7937);
buf BUF1 (N7951, N7934);
and AND2 (N7952, N7944, N5870);
and AND4 (N7953, N7949, N7826, N2674, N6426);
xor XOR2 (N7954, N7951, N2519);
not NOT1 (N7955, N7942);
nor NOR4 (N7956, N7947, N5554, N5874, N432);
and AND4 (N7957, N7952, N1837, N2437, N5680);
or OR2 (N7958, N7943, N5939);
not NOT1 (N7959, N7950);
not NOT1 (N7960, N7956);
buf BUF1 (N7961, N7960);
and AND2 (N7962, N7961, N49);
buf BUF1 (N7963, N7955);
or OR4 (N7964, N7953, N1887, N4146, N4009);
nor NOR2 (N7965, N7958, N23);
and AND3 (N7966, N7957, N7938, N3142);
not NOT1 (N7967, N7959);
buf BUF1 (N7968, N7962);
buf BUF1 (N7969, N7968);
buf BUF1 (N7970, N7966);
and AND3 (N7971, N7940, N7143, N3733);
or OR3 (N7972, N7954, N6725, N7556);
xor XOR2 (N7973, N7965, N1820);
buf BUF1 (N7974, N7973);
nand NAND4 (N7975, N7964, N975, N1403, N3100);
nor NOR2 (N7976, N7974, N6998);
nor NOR2 (N7977, N7963, N36);
buf BUF1 (N7978, N7970);
buf BUF1 (N7979, N7977);
buf BUF1 (N7980, N7933);
not NOT1 (N7981, N7967);
nor NOR3 (N7982, N7946, N5686, N3839);
buf BUF1 (N7983, N7975);
nand NAND2 (N7984, N7982, N7031);
not NOT1 (N7985, N7976);
buf BUF1 (N7986, N7980);
or OR2 (N7987, N7969, N7964);
nand NAND4 (N7988, N7983, N1940, N6571, N5137);
nor NOR4 (N7989, N7986, N6945, N6135, N6791);
and AND2 (N7990, N7978, N2110);
or OR2 (N7991, N7985, N2955);
buf BUF1 (N7992, N7971);
or OR2 (N7993, N7979, N6502);
nand NAND2 (N7994, N7988, N1313);
nand NAND4 (N7995, N7994, N5306, N1774, N1310);
xor XOR2 (N7996, N7984, N1995);
nand NAND4 (N7997, N7995, N3661, N2883, N4646);
not NOT1 (N7998, N7987);
and AND2 (N7999, N7998, N7492);
nand NAND2 (N8000, N7997, N6791);
nor NOR3 (N8001, N7989, N5059, N845);
nor NOR2 (N8002, N7992, N7834);
and AND4 (N8003, N8001, N795, N4146, N4043);
and AND4 (N8004, N7991, N3241, N1774, N5771);
or OR4 (N8005, N7996, N2723, N2041, N5581);
nand NAND2 (N8006, N7972, N3901);
or OR4 (N8007, N7981, N302, N1050, N3786);
nand NAND4 (N8008, N7993, N3707, N1819, N6483);
nor NOR4 (N8009, N8006, N5931, N1115, N4690);
nand NAND2 (N8010, N8004, N5968);
nand NAND3 (N8011, N8000, N5598, N687);
and AND3 (N8012, N8009, N5060, N6651);
not NOT1 (N8013, N7999);
not NOT1 (N8014, N8005);
not NOT1 (N8015, N7990);
nor NOR2 (N8016, N8011, N4446);
nor NOR3 (N8017, N8014, N114, N5711);
nand NAND4 (N8018, N8008, N5338, N7191, N2048);
nand NAND4 (N8019, N8016, N357, N3016, N645);
or OR3 (N8020, N8018, N7758, N4608);
xor XOR2 (N8021, N8020, N1566);
xor XOR2 (N8022, N8019, N7285);
nor NOR2 (N8023, N8017, N350);
or OR2 (N8024, N8022, N312);
buf BUF1 (N8025, N8010);
xor XOR2 (N8026, N8015, N2690);
buf BUF1 (N8027, N8013);
and AND3 (N8028, N8027, N6754, N3746);
not NOT1 (N8029, N8028);
not NOT1 (N8030, N8003);
nor NOR3 (N8031, N8024, N3983, N3968);
and AND2 (N8032, N8002, N2832);
and AND3 (N8033, N8032, N4658, N7856);
not NOT1 (N8034, N8031);
or OR3 (N8035, N8007, N363, N542);
buf BUF1 (N8036, N8021);
or OR3 (N8037, N8025, N2816, N1044);
buf BUF1 (N8038, N8012);
and AND3 (N8039, N8029, N7036, N4472);
or OR2 (N8040, N8026, N3722);
and AND2 (N8041, N8039, N7765);
xor XOR2 (N8042, N8038, N3364);
nor NOR4 (N8043, N8035, N4109, N6104, N4132);
or OR3 (N8044, N8034, N3891, N1125);
nor NOR2 (N8045, N8040, N2521);
nand NAND4 (N8046, N8023, N7057, N1612, N3259);
or OR4 (N8047, N8033, N5086, N1891, N5537);
not NOT1 (N8048, N8045);
not NOT1 (N8049, N8036);
xor XOR2 (N8050, N8037, N6108);
nor NOR3 (N8051, N8044, N6971, N4829);
nor NOR4 (N8052, N8048, N3465, N4543, N7233);
buf BUF1 (N8053, N8050);
buf BUF1 (N8054, N8042);
buf BUF1 (N8055, N8053);
and AND2 (N8056, N8055, N7898);
xor XOR2 (N8057, N8041, N5485);
and AND4 (N8058, N8052, N801, N1779, N4290);
buf BUF1 (N8059, N8046);
and AND3 (N8060, N8049, N535, N3476);
not NOT1 (N8061, N8057);
and AND3 (N8062, N8059, N2499, N996);
xor XOR2 (N8063, N8060, N2288);
and AND3 (N8064, N8056, N6206, N4642);
and AND4 (N8065, N8062, N7193, N1384, N2006);
and AND2 (N8066, N8063, N3319);
nor NOR4 (N8067, N8054, N6868, N5468, N4075);
buf BUF1 (N8068, N8064);
and AND4 (N8069, N8068, N3189, N7100, N2715);
buf BUF1 (N8070, N8030);
not NOT1 (N8071, N8058);
and AND4 (N8072, N8047, N7130, N2096, N1400);
xor XOR2 (N8073, N8069, N6718);
not NOT1 (N8074, N8071);
nand NAND4 (N8075, N8043, N1974, N282, N746);
xor XOR2 (N8076, N8075, N5141);
xor XOR2 (N8077, N8065, N7219);
not NOT1 (N8078, N8076);
or OR3 (N8079, N8061, N1532, N5290);
xor XOR2 (N8080, N8072, N3273);
xor XOR2 (N8081, N8079, N4301);
and AND3 (N8082, N8066, N974, N3605);
or OR3 (N8083, N8073, N6164, N14);
not NOT1 (N8084, N8082);
buf BUF1 (N8085, N8077);
buf BUF1 (N8086, N8081);
nor NOR4 (N8087, N8078, N5429, N4051, N1453);
or OR4 (N8088, N8074, N5540, N2380, N3697);
not NOT1 (N8089, N8084);
buf BUF1 (N8090, N8080);
and AND3 (N8091, N8087, N7445, N2100);
and AND3 (N8092, N8067, N1362, N7819);
not NOT1 (N8093, N8091);
or OR2 (N8094, N8093, N3204);
not NOT1 (N8095, N8086);
nand NAND3 (N8096, N8085, N990, N3189);
and AND4 (N8097, N8090, N2671, N247, N1629);
or OR3 (N8098, N8083, N3756, N7110);
or OR4 (N8099, N8098, N3733, N5457, N5650);
and AND4 (N8100, N8051, N5199, N7240, N4965);
nand NAND4 (N8101, N8095, N6313, N2123, N7761);
nand NAND2 (N8102, N8096, N3085);
xor XOR2 (N8103, N8088, N2235);
nand NAND3 (N8104, N8089, N4070, N8048);
not NOT1 (N8105, N8097);
not NOT1 (N8106, N8100);
buf BUF1 (N8107, N8106);
or OR4 (N8108, N8094, N2317, N2992, N1009);
xor XOR2 (N8109, N8102, N3202);
and AND2 (N8110, N8109, N4983);
not NOT1 (N8111, N8110);
or OR4 (N8112, N8111, N2921, N5210, N3798);
nor NOR2 (N8113, N8112, N6535);
nand NAND2 (N8114, N8092, N3800);
nor NOR2 (N8115, N8113, N3187);
and AND3 (N8116, N8070, N2658, N4064);
and AND3 (N8117, N8108, N1919, N6169);
or OR3 (N8118, N8116, N3686, N2252);
and AND3 (N8119, N8105, N4019, N6835);
nor NOR2 (N8120, N8119, N2943);
buf BUF1 (N8121, N8101);
buf BUF1 (N8122, N8118);
not NOT1 (N8123, N8104);
nor NOR2 (N8124, N8122, N6938);
not NOT1 (N8125, N8114);
buf BUF1 (N8126, N8099);
not NOT1 (N8127, N8123);
or OR4 (N8128, N8121, N2696, N485, N2386);
nor NOR3 (N8129, N8125, N4753, N8001);
nand NAND2 (N8130, N8103, N2234);
not NOT1 (N8131, N8107);
or OR4 (N8132, N8127, N3561, N6860, N596);
nor NOR3 (N8133, N8132, N5961, N6221);
nand NAND4 (N8134, N8130, N1447, N4131, N2460);
nor NOR4 (N8135, N8133, N5755, N6915, N6265);
xor XOR2 (N8136, N8120, N7423);
buf BUF1 (N8137, N8126);
nand NAND4 (N8138, N8134, N1828, N7506, N8016);
and AND4 (N8139, N8138, N1157, N2187, N6831);
nand NAND4 (N8140, N8124, N5281, N2213, N3290);
and AND2 (N8141, N8139, N1924);
not NOT1 (N8142, N8128);
not NOT1 (N8143, N8140);
buf BUF1 (N8144, N8115);
and AND4 (N8145, N8144, N3298, N4910, N2939);
and AND4 (N8146, N8129, N1172, N7889, N6098);
buf BUF1 (N8147, N8145);
buf BUF1 (N8148, N8142);
nor NOR3 (N8149, N8137, N1246, N3411);
nand NAND2 (N8150, N8131, N5217);
nand NAND2 (N8151, N8146, N7632);
nand NAND4 (N8152, N8117, N3917, N7168, N722);
buf BUF1 (N8153, N8151);
not NOT1 (N8154, N8141);
not NOT1 (N8155, N8154);
not NOT1 (N8156, N8143);
nand NAND4 (N8157, N8149, N575, N688, N7810);
and AND2 (N8158, N8157, N5848);
or OR3 (N8159, N8158, N7283, N3215);
not NOT1 (N8160, N8150);
nor NOR2 (N8161, N8159, N2271);
not NOT1 (N8162, N8135);
xor XOR2 (N8163, N8153, N7607);
buf BUF1 (N8164, N8136);
nor NOR2 (N8165, N8147, N5386);
nand NAND3 (N8166, N8160, N2140, N4127);
nand NAND2 (N8167, N8164, N4202);
nor NOR4 (N8168, N8162, N3026, N2969, N3649);
xor XOR2 (N8169, N8166, N7210);
and AND4 (N8170, N8155, N7601, N1108, N7078);
not NOT1 (N8171, N8165);
or OR4 (N8172, N8168, N5174, N1810, N7412);
not NOT1 (N8173, N8167);
not NOT1 (N8174, N8148);
nor NOR4 (N8175, N8156, N5424, N7002, N4128);
xor XOR2 (N8176, N8161, N2981);
nand NAND2 (N8177, N8170, N434);
not NOT1 (N8178, N8152);
or OR4 (N8179, N8178, N7391, N4918, N988);
nor NOR2 (N8180, N8174, N3963);
nor NOR2 (N8181, N8163, N540);
buf BUF1 (N8182, N8173);
buf BUF1 (N8183, N8169);
or OR3 (N8184, N8180, N5849, N446);
xor XOR2 (N8185, N8179, N6167);
buf BUF1 (N8186, N8175);
or OR3 (N8187, N8177, N7875, N2771);
buf BUF1 (N8188, N8185);
nand NAND4 (N8189, N8186, N1362, N3554, N4618);
buf BUF1 (N8190, N8184);
nor NOR3 (N8191, N8172, N103, N3101);
not NOT1 (N8192, N8187);
not NOT1 (N8193, N8191);
nand NAND4 (N8194, N8176, N704, N7886, N4268);
xor XOR2 (N8195, N8190, N3008);
buf BUF1 (N8196, N8188);
or OR4 (N8197, N8195, N1578, N4989, N4945);
or OR3 (N8198, N8196, N2061, N7933);
not NOT1 (N8199, N8198);
not NOT1 (N8200, N8194);
buf BUF1 (N8201, N8192);
xor XOR2 (N8202, N8183, N4607);
and AND4 (N8203, N8181, N1281, N4749, N3018);
nor NOR2 (N8204, N8202, N5195);
nor NOR4 (N8205, N8199, N4745, N5441, N3346);
not NOT1 (N8206, N8204);
nand NAND4 (N8207, N8200, N1080, N5095, N195);
or OR3 (N8208, N8207, N2918, N4883);
or OR3 (N8209, N8208, N3276, N168);
or OR2 (N8210, N8193, N4005);
xor XOR2 (N8211, N8205, N882);
nor NOR4 (N8212, N8201, N4521, N1256, N7198);
xor XOR2 (N8213, N8206, N1661);
xor XOR2 (N8214, N8189, N7322);
xor XOR2 (N8215, N8211, N1498);
or OR2 (N8216, N8215, N6999);
nand NAND3 (N8217, N8210, N789, N5822);
or OR2 (N8218, N8212, N2486);
buf BUF1 (N8219, N8209);
not NOT1 (N8220, N8182);
nand NAND2 (N8221, N8203, N6094);
nand NAND3 (N8222, N8217, N3926, N6822);
and AND4 (N8223, N8221, N4700, N1629, N6443);
or OR3 (N8224, N8213, N7397, N4556);
nor NOR4 (N8225, N8219, N5408, N5688, N4652);
not NOT1 (N8226, N8171);
nand NAND3 (N8227, N8226, N7206, N7809);
xor XOR2 (N8228, N8214, N6268);
nor NOR2 (N8229, N8228, N3204);
not NOT1 (N8230, N8227);
nor NOR2 (N8231, N8197, N3047);
buf BUF1 (N8232, N8229);
xor XOR2 (N8233, N8231, N4651);
and AND4 (N8234, N8216, N7915, N8016, N2672);
not NOT1 (N8235, N8225);
xor XOR2 (N8236, N8222, N2835);
xor XOR2 (N8237, N8236, N1971);
xor XOR2 (N8238, N8237, N7906);
nor NOR2 (N8239, N8223, N7210);
nor NOR3 (N8240, N8218, N670, N1938);
xor XOR2 (N8241, N8233, N2212);
and AND2 (N8242, N8235, N6654);
buf BUF1 (N8243, N8230);
xor XOR2 (N8244, N8232, N7855);
nand NAND2 (N8245, N8244, N2861);
not NOT1 (N8246, N8242);
buf BUF1 (N8247, N8245);
buf BUF1 (N8248, N8240);
xor XOR2 (N8249, N8224, N960);
xor XOR2 (N8250, N8246, N257);
or OR3 (N8251, N8248, N3930, N6025);
not NOT1 (N8252, N8239);
or OR4 (N8253, N8234, N5139, N7249, N1526);
nor NOR2 (N8254, N8247, N2921);
buf BUF1 (N8255, N8254);
nand NAND3 (N8256, N8249, N8012, N4460);
and AND4 (N8257, N8251, N35, N3696, N4282);
not NOT1 (N8258, N8257);
and AND4 (N8259, N8243, N308, N8251, N3037);
and AND4 (N8260, N8255, N7225, N652, N4626);
or OR4 (N8261, N8220, N2053, N5495, N708);
xor XOR2 (N8262, N8253, N1675);
nor NOR2 (N8263, N8241, N5761);
not NOT1 (N8264, N8238);
nor NOR2 (N8265, N8250, N1085);
nand NAND3 (N8266, N8260, N6302, N453);
or OR3 (N8267, N8264, N3431, N1391);
buf BUF1 (N8268, N8259);
xor XOR2 (N8269, N8267, N3430);
and AND3 (N8270, N8258, N2785, N3721);
xor XOR2 (N8271, N8252, N7109);
buf BUF1 (N8272, N8265);
buf BUF1 (N8273, N8261);
nor NOR3 (N8274, N8268, N1752, N5015);
and AND2 (N8275, N8263, N3646);
nand NAND3 (N8276, N8272, N5541, N4340);
and AND3 (N8277, N8276, N7414, N491);
not NOT1 (N8278, N8273);
or OR4 (N8279, N8275, N5814, N5293, N5484);
nand NAND2 (N8280, N8271, N6883);
or OR2 (N8281, N8266, N1120);
and AND3 (N8282, N8277, N3025, N1132);
nand NAND4 (N8283, N8278, N5152, N6375, N4568);
not NOT1 (N8284, N8279);
xor XOR2 (N8285, N8280, N7582);
and AND2 (N8286, N8285, N2406);
xor XOR2 (N8287, N8256, N3334);
buf BUF1 (N8288, N8270);
xor XOR2 (N8289, N8288, N2685);
nand NAND3 (N8290, N8287, N1857, N5583);
xor XOR2 (N8291, N8283, N3621);
or OR4 (N8292, N8262, N2454, N1168, N2176);
buf BUF1 (N8293, N8292);
or OR2 (N8294, N8282, N7529);
xor XOR2 (N8295, N8293, N5084);
buf BUF1 (N8296, N8295);
xor XOR2 (N8297, N8296, N546);
and AND4 (N8298, N8291, N8061, N5747, N3029);
and AND4 (N8299, N8289, N1494, N1614, N7715);
not NOT1 (N8300, N8284);
nand NAND3 (N8301, N8281, N231, N2951);
nor NOR2 (N8302, N8274, N3850);
nand NAND4 (N8303, N8300, N4228, N5980, N3819);
nand NAND2 (N8304, N8269, N2560);
nor NOR3 (N8305, N8303, N5769, N5928);
nor NOR2 (N8306, N8304, N1456);
and AND4 (N8307, N8301, N509, N4824, N6026);
nor NOR4 (N8308, N8307, N7845, N1153, N1950);
nand NAND2 (N8309, N8294, N6639);
or OR3 (N8310, N8306, N4020, N5096);
nand NAND3 (N8311, N8299, N7380, N6413);
nor NOR4 (N8312, N8297, N5389, N8024, N2073);
not NOT1 (N8313, N8309);
and AND4 (N8314, N8290, N518, N792, N1398);
not NOT1 (N8315, N8298);
xor XOR2 (N8316, N8311, N2147);
buf BUF1 (N8317, N8316);
not NOT1 (N8318, N8312);
nor NOR2 (N8319, N8310, N921);
nand NAND4 (N8320, N8313, N3894, N3509, N3657);
xor XOR2 (N8321, N8314, N6506);
and AND3 (N8322, N8305, N1692, N651);
and AND2 (N8323, N8321, N1110);
buf BUF1 (N8324, N8308);
or OR3 (N8325, N8319, N8302, N3791);
not NOT1 (N8326, N7917);
buf BUF1 (N8327, N8322);
or OR2 (N8328, N8326, N3898);
and AND2 (N8329, N8315, N1490);
buf BUF1 (N8330, N8325);
and AND4 (N8331, N8318, N2587, N3728, N318);
xor XOR2 (N8332, N8286, N7680);
nand NAND2 (N8333, N8330, N3759);
nor NOR4 (N8334, N8324, N990, N3046, N5838);
xor XOR2 (N8335, N8323, N2203);
or OR2 (N8336, N8328, N4655);
not NOT1 (N8337, N8334);
and AND4 (N8338, N8337, N5620, N3752, N4115);
buf BUF1 (N8339, N8335);
nand NAND3 (N8340, N8329, N1743, N4318);
nand NAND3 (N8341, N8333, N2787, N6920);
nand NAND3 (N8342, N8339, N5291, N1100);
buf BUF1 (N8343, N8338);
and AND2 (N8344, N8336, N5222);
not NOT1 (N8345, N8341);
buf BUF1 (N8346, N8320);
buf BUF1 (N8347, N8340);
nor NOR2 (N8348, N8346, N2600);
xor XOR2 (N8349, N8332, N6704);
xor XOR2 (N8350, N8349, N3804);
and AND2 (N8351, N8343, N2088);
nand NAND4 (N8352, N8348, N33, N1658, N899);
buf BUF1 (N8353, N8351);
xor XOR2 (N8354, N8350, N5209);
xor XOR2 (N8355, N8354, N1062);
xor XOR2 (N8356, N8352, N3386);
buf BUF1 (N8357, N8327);
not NOT1 (N8358, N8347);
nand NAND2 (N8359, N8355, N1311);
nand NAND3 (N8360, N8358, N7430, N5208);
nor NOR3 (N8361, N8356, N2252, N6811);
buf BUF1 (N8362, N8361);
not NOT1 (N8363, N8331);
buf BUF1 (N8364, N8360);
or OR4 (N8365, N8344, N7231, N3494, N3542);
nor NOR3 (N8366, N8359, N5063, N2318);
nand NAND2 (N8367, N8366, N5343);
xor XOR2 (N8368, N8317, N7028);
xor XOR2 (N8369, N8345, N5673);
or OR2 (N8370, N8369, N6837);
not NOT1 (N8371, N8367);
buf BUF1 (N8372, N8371);
not NOT1 (N8373, N8368);
and AND3 (N8374, N8364, N8215, N5126);
xor XOR2 (N8375, N8372, N3132);
nor NOR3 (N8376, N8370, N4741, N2792);
buf BUF1 (N8377, N8363);
nor NOR2 (N8378, N8375, N2119);
xor XOR2 (N8379, N8342, N221);
buf BUF1 (N8380, N8378);
nor NOR3 (N8381, N8376, N2159, N1413);
buf BUF1 (N8382, N8373);
xor XOR2 (N8383, N8379, N4022);
or OR4 (N8384, N8374, N2235, N912, N5823);
or OR3 (N8385, N8383, N4908, N4878);
or OR2 (N8386, N8357, N4283);
nor NOR3 (N8387, N8386, N2823, N3313);
buf BUF1 (N8388, N8377);
nand NAND4 (N8389, N8385, N6261, N4811, N3721);
not NOT1 (N8390, N8382);
or OR2 (N8391, N8362, N7857);
nand NAND2 (N8392, N8389, N567);
not NOT1 (N8393, N8353);
buf BUF1 (N8394, N8387);
xor XOR2 (N8395, N8391, N7483);
and AND3 (N8396, N8380, N8279, N3422);
xor XOR2 (N8397, N8388, N485);
not NOT1 (N8398, N8365);
xor XOR2 (N8399, N8384, N4878);
not NOT1 (N8400, N8396);
not NOT1 (N8401, N8393);
nor NOR2 (N8402, N8394, N6010);
buf BUF1 (N8403, N8397);
nor NOR4 (N8404, N8381, N4125, N1233, N3980);
xor XOR2 (N8405, N8401, N5448);
and AND3 (N8406, N8402, N5610, N4024);
nor NOR4 (N8407, N8395, N7647, N3547, N7127);
nand NAND2 (N8408, N8405, N4746);
nor NOR2 (N8409, N8398, N3797);
nor NOR2 (N8410, N8392, N114);
not NOT1 (N8411, N8406);
buf BUF1 (N8412, N8400);
nand NAND2 (N8413, N8390, N5447);
and AND3 (N8414, N8403, N6145, N1367);
not NOT1 (N8415, N8399);
not NOT1 (N8416, N8412);
or OR3 (N8417, N8415, N1553, N1615);
not NOT1 (N8418, N8414);
or OR4 (N8419, N8409, N475, N5251, N1880);
buf BUF1 (N8420, N8413);
or OR4 (N8421, N8416, N3589, N4467, N2525);
nand NAND3 (N8422, N8411, N415, N5345);
buf BUF1 (N8423, N8410);
xor XOR2 (N8424, N8421, N6753);
not NOT1 (N8425, N8407);
not NOT1 (N8426, N8404);
xor XOR2 (N8427, N8422, N8117);
or OR2 (N8428, N8427, N6263);
xor XOR2 (N8429, N8420, N25);
or OR2 (N8430, N8424, N4296);
xor XOR2 (N8431, N8425, N3365);
buf BUF1 (N8432, N8419);
xor XOR2 (N8433, N8418, N4695);
nor NOR3 (N8434, N8431, N1347, N4092);
and AND4 (N8435, N8432, N1611, N2264, N3007);
or OR2 (N8436, N8423, N6885);
nand NAND3 (N8437, N8430, N3051, N960);
and AND2 (N8438, N8429, N4087);
and AND2 (N8439, N8435, N3021);
xor XOR2 (N8440, N8426, N5098);
buf BUF1 (N8441, N8434);
not NOT1 (N8442, N8437);
nor NOR3 (N8443, N8436, N3600, N2734);
and AND4 (N8444, N8428, N30, N5942, N8208);
or OR4 (N8445, N8433, N6854, N5652, N458);
or OR2 (N8446, N8417, N3519);
not NOT1 (N8447, N8438);
nand NAND2 (N8448, N8442, N1535);
not NOT1 (N8449, N8448);
and AND3 (N8450, N8447, N2428, N2249);
xor XOR2 (N8451, N8444, N2558);
nor NOR3 (N8452, N8445, N6544, N1019);
not NOT1 (N8453, N8452);
buf BUF1 (N8454, N8408);
and AND4 (N8455, N8443, N3519, N5051, N2730);
and AND4 (N8456, N8441, N6609, N5356, N1931);
or OR4 (N8457, N8446, N7518, N1258, N6788);
nor NOR4 (N8458, N8439, N7652, N3983, N201);
xor XOR2 (N8459, N8453, N5070);
nand NAND4 (N8460, N8454, N514, N4656, N314);
buf BUF1 (N8461, N8449);
and AND3 (N8462, N8461, N8399, N1348);
and AND2 (N8463, N8460, N473);
xor XOR2 (N8464, N8459, N5168);
or OR2 (N8465, N8463, N7982);
nand NAND2 (N8466, N8464, N6920);
xor XOR2 (N8467, N8440, N7456);
or OR2 (N8468, N8465, N594);
nand NAND3 (N8469, N8457, N697, N5698);
or OR3 (N8470, N8469, N2631, N1670);
xor XOR2 (N8471, N8467, N3680);
buf BUF1 (N8472, N8451);
buf BUF1 (N8473, N8455);
nor NOR3 (N8474, N8456, N4991, N681);
and AND2 (N8475, N8473, N977);
xor XOR2 (N8476, N8462, N3422);
nor NOR4 (N8477, N8470, N7664, N1227, N2103);
xor XOR2 (N8478, N8476, N3065);
buf BUF1 (N8479, N8468);
nand NAND2 (N8480, N8458, N6289);
xor XOR2 (N8481, N8450, N5408);
or OR4 (N8482, N8480, N1832, N325, N5554);
not NOT1 (N8483, N8474);
and AND2 (N8484, N8475, N465);
xor XOR2 (N8485, N8482, N4843);
nand NAND3 (N8486, N8479, N7320, N329);
nand NAND4 (N8487, N8471, N693, N8317, N4994);
nor NOR2 (N8488, N8477, N7305);
buf BUF1 (N8489, N8472);
nor NOR3 (N8490, N8485, N5130, N3263);
xor XOR2 (N8491, N8486, N1519);
or OR2 (N8492, N8481, N2162);
or OR2 (N8493, N8487, N1413);
buf BUF1 (N8494, N8466);
or OR2 (N8495, N8489, N3927);
or OR3 (N8496, N8484, N7600, N6786);
and AND2 (N8497, N8488, N4033);
xor XOR2 (N8498, N8496, N4016);
nor NOR2 (N8499, N8493, N2829);
nor NOR4 (N8500, N8494, N4565, N1635, N5689);
nor NOR4 (N8501, N8491, N6703, N2032, N2256);
xor XOR2 (N8502, N8501, N4383);
or OR2 (N8503, N8478, N5846);
not NOT1 (N8504, N8498);
xor XOR2 (N8505, N8503, N7869);
nand NAND3 (N8506, N8500, N6202, N2192);
or OR2 (N8507, N8502, N836);
not NOT1 (N8508, N8495);
nor NOR3 (N8509, N8505, N5603, N7634);
and AND3 (N8510, N8490, N4892, N4709);
nand NAND4 (N8511, N8492, N3197, N6960, N2526);
not NOT1 (N8512, N8497);
xor XOR2 (N8513, N8506, N7487);
or OR2 (N8514, N8507, N2037);
and AND2 (N8515, N8509, N8089);
or OR2 (N8516, N8512, N2314);
not NOT1 (N8517, N8508);
xor XOR2 (N8518, N8511, N8002);
or OR4 (N8519, N8515, N1699, N4838, N3980);
nand NAND4 (N8520, N8519, N1374, N8121, N2627);
not NOT1 (N8521, N8517);
nor NOR3 (N8522, N8513, N289, N3567);
nand NAND4 (N8523, N8521, N6037, N7957, N4221);
nand NAND4 (N8524, N8516, N4661, N847, N1254);
not NOT1 (N8525, N8510);
nor NOR2 (N8526, N8514, N1742);
nor NOR2 (N8527, N8523, N1139);
nor NOR3 (N8528, N8524, N3749, N2298);
or OR4 (N8529, N8525, N4440, N6060, N8456);
nor NOR3 (N8530, N8529, N1092, N7440);
nor NOR3 (N8531, N8528, N306, N1338);
nand NAND4 (N8532, N8483, N3720, N3866, N2945);
nor NOR2 (N8533, N8530, N5614);
nand NAND4 (N8534, N8499, N3934, N8452, N7);
not NOT1 (N8535, N8533);
nand NAND4 (N8536, N8535, N899, N5633, N6760);
not NOT1 (N8537, N8536);
nor NOR3 (N8538, N8520, N3315, N7460);
buf BUF1 (N8539, N8518);
xor XOR2 (N8540, N8527, N3110);
nand NAND2 (N8541, N8522, N5304);
nand NAND2 (N8542, N8540, N2979);
nand NAND2 (N8543, N8542, N7181);
nor NOR3 (N8544, N8531, N1018, N4966);
xor XOR2 (N8545, N8537, N3519);
not NOT1 (N8546, N8526);
not NOT1 (N8547, N8532);
nand NAND4 (N8548, N8544, N7430, N7172, N956);
and AND3 (N8549, N8539, N7656, N1613);
not NOT1 (N8550, N8546);
or OR4 (N8551, N8550, N3685, N3923, N3188);
nor NOR3 (N8552, N8541, N4726, N1003);
nor NOR3 (N8553, N8504, N119, N5292);
not NOT1 (N8554, N8552);
xor XOR2 (N8555, N8534, N7385);
not NOT1 (N8556, N8553);
or OR4 (N8557, N8554, N1256, N6655, N2456);
nor NOR2 (N8558, N8557, N1418);
xor XOR2 (N8559, N8545, N2842);
xor XOR2 (N8560, N8538, N1528);
and AND4 (N8561, N8543, N3049, N879, N6304);
buf BUF1 (N8562, N8551);
and AND4 (N8563, N8559, N6695, N3963, N7591);
xor XOR2 (N8564, N8561, N522);
nor NOR4 (N8565, N8562, N5491, N6020, N1112);
not NOT1 (N8566, N8548);
or OR4 (N8567, N8556, N5266, N6029, N3014);
nor NOR2 (N8568, N8560, N8123);
and AND3 (N8569, N8564, N7809, N1486);
and AND2 (N8570, N8555, N932);
nor NOR2 (N8571, N8570, N3779);
and AND3 (N8572, N8547, N7487, N4040);
or OR3 (N8573, N8572, N3782, N7472);
nor NOR4 (N8574, N8568, N4982, N4748, N218);
nand NAND4 (N8575, N8558, N7171, N71, N6093);
and AND2 (N8576, N8549, N7873);
nor NOR2 (N8577, N8567, N1420);
not NOT1 (N8578, N8574);
nand NAND3 (N8579, N8577, N5945, N6954);
or OR3 (N8580, N8578, N577, N8433);
buf BUF1 (N8581, N8566);
xor XOR2 (N8582, N8571, N7596);
nor NOR2 (N8583, N8569, N7240);
buf BUF1 (N8584, N8563);
or OR2 (N8585, N8573, N6204);
nor NOR4 (N8586, N8576, N5448, N7018, N3208);
and AND4 (N8587, N8582, N3069, N4636, N8266);
or OR3 (N8588, N8579, N5717, N4935);
buf BUF1 (N8589, N8586);
nand NAND3 (N8590, N8584, N3456, N8501);
or OR3 (N8591, N8583, N3727, N1883);
buf BUF1 (N8592, N8575);
nand NAND3 (N8593, N8587, N481, N6432);
or OR2 (N8594, N8591, N7298);
or OR3 (N8595, N8581, N2530, N2307);
and AND2 (N8596, N8594, N7142);
buf BUF1 (N8597, N8592);
and AND3 (N8598, N8597, N3209, N160);
nand NAND3 (N8599, N8590, N6645, N4937);
and AND3 (N8600, N8593, N1222, N1483);
nand NAND3 (N8601, N8595, N735, N6271);
xor XOR2 (N8602, N8588, N5258);
buf BUF1 (N8603, N8565);
and AND2 (N8604, N8589, N6910);
nor NOR3 (N8605, N8585, N1396, N6810);
not NOT1 (N8606, N8599);
nor NOR2 (N8607, N8598, N8553);
or OR2 (N8608, N8602, N6964);
nand NAND2 (N8609, N8600, N1470);
nand NAND4 (N8610, N8604, N7205, N3491, N2874);
nor NOR2 (N8611, N8580, N6058);
or OR2 (N8612, N8601, N8377);
not NOT1 (N8613, N8606);
nor NOR2 (N8614, N8608, N7033);
or OR4 (N8615, N8612, N7006, N8190, N5170);
not NOT1 (N8616, N8614);
nand NAND4 (N8617, N8615, N1608, N7979, N6736);
not NOT1 (N8618, N8607);
not NOT1 (N8619, N8603);
not NOT1 (N8620, N8613);
not NOT1 (N8621, N8619);
or OR4 (N8622, N8618, N8372, N2404, N996);
and AND4 (N8623, N8616, N2366, N667, N4227);
nand NAND3 (N8624, N8622, N1338, N2552);
nor NOR4 (N8625, N8611, N5074, N8623, N370);
nor NOR4 (N8626, N1879, N3972, N6566, N6305);
and AND3 (N8627, N8620, N76, N6443);
nand NAND4 (N8628, N8621, N2255, N2955, N832);
or OR3 (N8629, N8609, N7940, N100);
nand NAND2 (N8630, N8605, N805);
or OR4 (N8631, N8610, N2114, N7033, N61);
nand NAND4 (N8632, N8617, N1334, N8173, N704);
nor NOR3 (N8633, N8631, N3265, N5497);
nand NAND4 (N8634, N8596, N865, N52, N4878);
and AND3 (N8635, N8628, N3712, N713);
or OR3 (N8636, N8633, N6370, N1237);
nand NAND2 (N8637, N8624, N7637);
or OR4 (N8638, N8635, N7061, N8139, N3265);
nand NAND3 (N8639, N8626, N5610, N2329);
and AND3 (N8640, N8636, N1725, N8513);
or OR2 (N8641, N8634, N7925);
and AND4 (N8642, N8637, N1459, N2220, N1680);
not NOT1 (N8643, N8627);
not NOT1 (N8644, N8642);
not NOT1 (N8645, N8629);
xor XOR2 (N8646, N8638, N5185);
or OR2 (N8647, N8640, N2296);
or OR4 (N8648, N8645, N5649, N7901, N612);
not NOT1 (N8649, N8643);
xor XOR2 (N8650, N8625, N7312);
buf BUF1 (N8651, N8649);
nor NOR3 (N8652, N8630, N6950, N7489);
nand NAND3 (N8653, N8639, N6553, N3494);
and AND3 (N8654, N8648, N3057, N749);
xor XOR2 (N8655, N8644, N8448);
nor NOR4 (N8656, N8650, N2894, N7980, N2482);
nor NOR3 (N8657, N8656, N5408, N7258);
and AND4 (N8658, N8641, N170, N1667, N1889);
or OR4 (N8659, N8655, N1380, N806, N5818);
and AND3 (N8660, N8654, N7858, N1912);
and AND4 (N8661, N8651, N2004, N1072, N3211);
xor XOR2 (N8662, N8658, N8370);
or OR2 (N8663, N8657, N4259);
xor XOR2 (N8664, N8660, N8354);
or OR3 (N8665, N8647, N7360, N5675);
xor XOR2 (N8666, N8646, N1300);
or OR2 (N8667, N8661, N4660);
and AND4 (N8668, N8652, N3602, N2468, N3500);
nand NAND4 (N8669, N8665, N16, N2482, N7238);
xor XOR2 (N8670, N8653, N6730);
nor NOR2 (N8671, N8663, N3495);
and AND4 (N8672, N8671, N342, N1209, N2338);
or OR2 (N8673, N8632, N3055);
nand NAND2 (N8674, N8662, N4652);
buf BUF1 (N8675, N8669);
xor XOR2 (N8676, N8667, N1745);
xor XOR2 (N8677, N8670, N3911);
or OR3 (N8678, N8666, N4246, N7108);
nor NOR3 (N8679, N8676, N2648, N8069);
and AND2 (N8680, N8673, N505);
buf BUF1 (N8681, N8672);
buf BUF1 (N8682, N8675);
buf BUF1 (N8683, N8680);
xor XOR2 (N8684, N8679, N4362);
not NOT1 (N8685, N8681);
not NOT1 (N8686, N8674);
xor XOR2 (N8687, N8677, N5432);
nand NAND4 (N8688, N8685, N8530, N8070, N149);
nor NOR2 (N8689, N8668, N6602);
and AND4 (N8690, N8683, N3032, N2509, N1620);
not NOT1 (N8691, N8684);
not NOT1 (N8692, N8688);
nor NOR2 (N8693, N8689, N3513);
nor NOR4 (N8694, N8693, N4075, N6048, N2546);
xor XOR2 (N8695, N8691, N5326);
buf BUF1 (N8696, N8692);
nand NAND2 (N8697, N8686, N180);
nand NAND3 (N8698, N8659, N1446, N895);
and AND3 (N8699, N8695, N3682, N3774);
and AND3 (N8700, N8694, N7496, N7213);
buf BUF1 (N8701, N8687);
or OR3 (N8702, N8664, N6429, N4711);
buf BUF1 (N8703, N8696);
buf BUF1 (N8704, N8701);
buf BUF1 (N8705, N8700);
and AND4 (N8706, N8698, N7834, N2366, N3008);
xor XOR2 (N8707, N8678, N565);
and AND4 (N8708, N8697, N4012, N1325, N8283);
nand NAND2 (N8709, N8682, N2917);
buf BUF1 (N8710, N8705);
buf BUF1 (N8711, N8704);
xor XOR2 (N8712, N8709, N2278);
and AND4 (N8713, N8708, N5336, N1188, N8447);
buf BUF1 (N8714, N8713);
not NOT1 (N8715, N8711);
xor XOR2 (N8716, N8699, N2993);
or OR4 (N8717, N8706, N1352, N4260, N134);
or OR3 (N8718, N8690, N245, N8492);
buf BUF1 (N8719, N8715);
buf BUF1 (N8720, N8716);
nor NOR4 (N8721, N8717, N6340, N6973, N7750);
nor NOR3 (N8722, N8707, N1182, N580);
xor XOR2 (N8723, N8714, N6054);
not NOT1 (N8724, N8703);
buf BUF1 (N8725, N8702);
nor NOR2 (N8726, N8720, N7233);
not NOT1 (N8727, N8726);
nand NAND3 (N8728, N8719, N4153, N182);
or OR4 (N8729, N8712, N4081, N7676, N4537);
xor XOR2 (N8730, N8724, N4607);
xor XOR2 (N8731, N8723, N4166);
and AND2 (N8732, N8725, N2282);
nand NAND3 (N8733, N8721, N3573, N3972);
or OR4 (N8734, N8710, N5045, N2006, N3098);
and AND3 (N8735, N8734, N2177, N1613);
xor XOR2 (N8736, N8731, N8605);
nand NAND4 (N8737, N8722, N3497, N4859, N910);
xor XOR2 (N8738, N8732, N1022);
or OR3 (N8739, N8738, N1508, N1414);
not NOT1 (N8740, N8737);
xor XOR2 (N8741, N8736, N8159);
and AND2 (N8742, N8741, N5281);
and AND2 (N8743, N8735, N1450);
or OR4 (N8744, N8733, N123, N7785, N3316);
nand NAND4 (N8745, N8742, N5332, N2195, N224);
and AND3 (N8746, N8718, N6159, N3173);
or OR3 (N8747, N8727, N5156, N4154);
buf BUF1 (N8748, N8728);
xor XOR2 (N8749, N8739, N4171);
buf BUF1 (N8750, N8744);
not NOT1 (N8751, N8740);
and AND2 (N8752, N8747, N5592);
xor XOR2 (N8753, N8743, N8329);
or OR2 (N8754, N8730, N2730);
nand NAND2 (N8755, N8754, N6800);
nand NAND3 (N8756, N8748, N3724, N3095);
not NOT1 (N8757, N8752);
and AND4 (N8758, N8729, N3910, N1595, N5464);
nor NOR2 (N8759, N8758, N8627);
and AND2 (N8760, N8750, N2808);
nand NAND4 (N8761, N8745, N5337, N7039, N5988);
buf BUF1 (N8762, N8759);
xor XOR2 (N8763, N8761, N7864);
or OR3 (N8764, N8763, N8623, N7933);
xor XOR2 (N8765, N8755, N1942);
xor XOR2 (N8766, N8753, N2984);
xor XOR2 (N8767, N8751, N6810);
and AND4 (N8768, N8762, N5657, N2178, N1731);
xor XOR2 (N8769, N8746, N5279);
nand NAND4 (N8770, N8769, N2573, N1208, N1362);
buf BUF1 (N8771, N8768);
buf BUF1 (N8772, N8765);
or OR4 (N8773, N8772, N7262, N4316, N8745);
nand NAND2 (N8774, N8767, N1068);
nor NOR2 (N8775, N8760, N788);
or OR2 (N8776, N8775, N677);
nor NOR3 (N8777, N8776, N4152, N2469);
nand NAND3 (N8778, N8757, N6257, N8129);
xor XOR2 (N8779, N8773, N3874);
buf BUF1 (N8780, N8749);
or OR4 (N8781, N8770, N6835, N250, N1533);
nor NOR4 (N8782, N8764, N2397, N8319, N4745);
buf BUF1 (N8783, N8782);
buf BUF1 (N8784, N8779);
nand NAND2 (N8785, N8756, N4702);
and AND4 (N8786, N8781, N1042, N2872, N4913);
and AND2 (N8787, N8777, N7996);
nor NOR2 (N8788, N8784, N1746);
nor NOR2 (N8789, N8786, N5689);
buf BUF1 (N8790, N8783);
xor XOR2 (N8791, N8774, N4487);
or OR2 (N8792, N8778, N145);
not NOT1 (N8793, N8787);
and AND2 (N8794, N8789, N2354);
nor NOR4 (N8795, N8785, N1596, N5904, N796);
nand NAND4 (N8796, N8792, N6594, N4508, N5765);
nand NAND3 (N8797, N8780, N5908, N6983);
not NOT1 (N8798, N8797);
nand NAND2 (N8799, N8788, N3321);
buf BUF1 (N8800, N8790);
nor NOR3 (N8801, N8791, N3271, N5028);
nand NAND3 (N8802, N8766, N1872, N8718);
and AND3 (N8803, N8798, N7269, N2598);
not NOT1 (N8804, N8771);
not NOT1 (N8805, N8800);
not NOT1 (N8806, N8795);
not NOT1 (N8807, N8803);
buf BUF1 (N8808, N8804);
and AND2 (N8809, N8801, N3541);
buf BUF1 (N8810, N8796);
not NOT1 (N8811, N8794);
buf BUF1 (N8812, N8799);
nand NAND2 (N8813, N8805, N4136);
or OR3 (N8814, N8802, N7189, N3993);
nor NOR2 (N8815, N8813, N8191);
xor XOR2 (N8816, N8809, N8517);
nor NOR2 (N8817, N8815, N3535);
buf BUF1 (N8818, N8793);
nand NAND3 (N8819, N8806, N4322, N7525);
xor XOR2 (N8820, N8812, N5371);
buf BUF1 (N8821, N8819);
xor XOR2 (N8822, N8807, N2412);
and AND3 (N8823, N8808, N8667, N4068);
and AND3 (N8824, N8821, N6911, N2986);
buf BUF1 (N8825, N8820);
xor XOR2 (N8826, N8817, N8204);
nand NAND2 (N8827, N8816, N8756);
or OR4 (N8828, N8825, N4111, N1871, N36);
xor XOR2 (N8829, N8814, N2672);
nand NAND3 (N8830, N8824, N5374, N6156);
nand NAND4 (N8831, N8811, N5074, N7504, N3271);
nand NAND4 (N8832, N8826, N1736, N3069, N1317);
buf BUF1 (N8833, N8827);
xor XOR2 (N8834, N8822, N944);
buf BUF1 (N8835, N8818);
not NOT1 (N8836, N8810);
or OR2 (N8837, N8832, N6067);
or OR3 (N8838, N8833, N8067, N1835);
xor XOR2 (N8839, N8836, N6856);
not NOT1 (N8840, N8828);
xor XOR2 (N8841, N8837, N2975);
buf BUF1 (N8842, N8838);
nor NOR4 (N8843, N8840, N6937, N6515, N2644);
nor NOR3 (N8844, N8835, N1296, N2516);
nor NOR4 (N8845, N8834, N5196, N5583, N5656);
buf BUF1 (N8846, N8842);
or OR2 (N8847, N8846, N5261);
nand NAND2 (N8848, N8829, N6381);
buf BUF1 (N8849, N8830);
nand NAND4 (N8850, N8845, N3529, N8276, N4155);
and AND3 (N8851, N8849, N4273, N1534);
buf BUF1 (N8852, N8839);
buf BUF1 (N8853, N8847);
and AND3 (N8854, N8841, N3864, N5652);
or OR3 (N8855, N8844, N6997, N5410);
nor NOR2 (N8856, N8843, N5386);
and AND3 (N8857, N8853, N6910, N979);
nor NOR4 (N8858, N8856, N8769, N4123, N4790);
or OR3 (N8859, N8852, N150, N746);
and AND4 (N8860, N8859, N6090, N5746, N328);
or OR3 (N8861, N8823, N1161, N1727);
nand NAND3 (N8862, N8848, N5650, N8855);
xor XOR2 (N8863, N1697, N5288);
or OR3 (N8864, N8863, N7983, N5859);
not NOT1 (N8865, N8858);
and AND2 (N8866, N8865, N4411);
nor NOR3 (N8867, N8857, N3487, N7077);
nor NOR3 (N8868, N8861, N3814, N6725);
xor XOR2 (N8869, N8867, N2715);
or OR2 (N8870, N8869, N3153);
nor NOR2 (N8871, N8866, N7339);
nand NAND3 (N8872, N8862, N5740, N742);
and AND3 (N8873, N8850, N843, N3853);
and AND4 (N8874, N8871, N1294, N7088, N4094);
nor NOR4 (N8875, N8860, N2264, N3053, N4559);
or OR2 (N8876, N8873, N7325);
nor NOR4 (N8877, N8872, N3425, N8234, N263);
nor NOR4 (N8878, N8876, N7804, N878, N1967);
nor NOR3 (N8879, N8870, N5772, N7642);
and AND4 (N8880, N8879, N2641, N7892, N1626);
nand NAND3 (N8881, N8851, N6950, N5047);
and AND4 (N8882, N8880, N447, N7264, N4330);
nor NOR4 (N8883, N8875, N8163, N3907, N5367);
nand NAND3 (N8884, N8854, N6908, N5578);
or OR3 (N8885, N8878, N6857, N6484);
and AND4 (N8886, N8881, N5934, N5040, N5549);
and AND3 (N8887, N8886, N4034, N408);
nor NOR3 (N8888, N8884, N8486, N5333);
or OR3 (N8889, N8831, N1271, N2093);
not NOT1 (N8890, N8883);
and AND3 (N8891, N8877, N7643, N4619);
xor XOR2 (N8892, N8890, N7415);
nor NOR4 (N8893, N8888, N8124, N8741, N938);
nand NAND3 (N8894, N8864, N2884, N4403);
and AND3 (N8895, N8874, N8174, N1626);
or OR4 (N8896, N8885, N3604, N2465, N6401);
or OR2 (N8897, N8895, N859);
nand NAND2 (N8898, N8891, N5033);
and AND4 (N8899, N8896, N5987, N3900, N6328);
nand NAND2 (N8900, N8889, N5997);
not NOT1 (N8901, N8897);
and AND3 (N8902, N8899, N8332, N3602);
nor NOR3 (N8903, N8882, N2480, N3478);
and AND3 (N8904, N8868, N84, N5839);
nor NOR2 (N8905, N8894, N3249);
xor XOR2 (N8906, N8902, N8146);
nand NAND3 (N8907, N8901, N8356, N5450);
xor XOR2 (N8908, N8906, N3878);
buf BUF1 (N8909, N8907);
not NOT1 (N8910, N8905);
nand NAND2 (N8911, N8909, N7401);
or OR3 (N8912, N8910, N2488, N4346);
xor XOR2 (N8913, N8904, N7152);
not NOT1 (N8914, N8900);
xor XOR2 (N8915, N8913, N7238);
nand NAND2 (N8916, N8911, N8344);
and AND4 (N8917, N8912, N4091, N4116, N3007);
nand NAND2 (N8918, N8916, N2933);
nor NOR4 (N8919, N8917, N483, N5786, N7678);
or OR3 (N8920, N8887, N3988, N2225);
and AND3 (N8921, N8908, N7041, N4453);
xor XOR2 (N8922, N8920, N5270);
not NOT1 (N8923, N8915);
xor XOR2 (N8924, N8898, N564);
xor XOR2 (N8925, N8922, N1212);
nor NOR3 (N8926, N8924, N7939, N7827);
nand NAND3 (N8927, N8925, N2444, N7235);
and AND3 (N8928, N8921, N4327, N3629);
nand NAND4 (N8929, N8927, N3190, N1951, N6473);
and AND4 (N8930, N8923, N4153, N3112, N5811);
nor NOR4 (N8931, N8930, N3736, N3160, N8490);
and AND4 (N8932, N8914, N5121, N803, N4617);
and AND3 (N8933, N8929, N8513, N7925);
xor XOR2 (N8934, N8918, N5133);
nand NAND2 (N8935, N8893, N7344);
buf BUF1 (N8936, N8903);
buf BUF1 (N8937, N8926);
buf BUF1 (N8938, N8919);
nor NOR2 (N8939, N8937, N6963);
nand NAND3 (N8940, N8933, N5165, N8672);
nand NAND4 (N8941, N8928, N7309, N8549, N8468);
nand NAND3 (N8942, N8892, N5217, N1077);
buf BUF1 (N8943, N8942);
not NOT1 (N8944, N8943);
xor XOR2 (N8945, N8941, N3160);
or OR2 (N8946, N8940, N1975);
nand NAND3 (N8947, N8936, N7434, N7283);
nor NOR2 (N8948, N8938, N5695);
and AND3 (N8949, N8931, N8257, N5066);
nand NAND2 (N8950, N8948, N6517);
buf BUF1 (N8951, N8950);
xor XOR2 (N8952, N8951, N712);
or OR2 (N8953, N8935, N6845);
not NOT1 (N8954, N8932);
or OR3 (N8955, N8947, N343, N2815);
and AND2 (N8956, N8955, N7370);
or OR2 (N8957, N8939, N1925);
xor XOR2 (N8958, N8957, N3889);
nand NAND4 (N8959, N8958, N141, N1744, N2498);
and AND3 (N8960, N8953, N5213, N4136);
xor XOR2 (N8961, N8949, N2738);
nor NOR4 (N8962, N8959, N2137, N254, N4439);
nand NAND3 (N8963, N8956, N8533, N1721);
xor XOR2 (N8964, N8961, N2473);
nand NAND3 (N8965, N8946, N2623, N7764);
nand NAND2 (N8966, N8963, N6440);
nor NOR3 (N8967, N8944, N6171, N1660);
xor XOR2 (N8968, N8934, N133);
not NOT1 (N8969, N8960);
not NOT1 (N8970, N8965);
not NOT1 (N8971, N8964);
buf BUF1 (N8972, N8952);
nand NAND3 (N8973, N8954, N1148, N6408);
or OR2 (N8974, N8968, N5883);
buf BUF1 (N8975, N8967);
not NOT1 (N8976, N8945);
buf BUF1 (N8977, N8969);
nand NAND3 (N8978, N8973, N8207, N4517);
and AND2 (N8979, N8976, N8768);
and AND2 (N8980, N8974, N4120);
buf BUF1 (N8981, N8978);
or OR4 (N8982, N8971, N7480, N8013, N3137);
and AND3 (N8983, N8981, N6341, N7230);
nand NAND4 (N8984, N8972, N464, N2723, N3756);
and AND3 (N8985, N8962, N1457, N6501);
buf BUF1 (N8986, N8980);
xor XOR2 (N8987, N8970, N2242);
or OR2 (N8988, N8983, N3438);
or OR2 (N8989, N8975, N1508);
not NOT1 (N8990, N8989);
or OR3 (N8991, N8982, N3328, N5312);
nand NAND3 (N8992, N8987, N2046, N2079);
or OR4 (N8993, N8966, N4182, N6155, N5960);
buf BUF1 (N8994, N8990);
and AND4 (N8995, N8992, N7770, N2922, N1190);
xor XOR2 (N8996, N8984, N4872);
and AND4 (N8997, N8986, N6451, N1061, N4216);
not NOT1 (N8998, N8977);
and AND4 (N8999, N8985, N594, N8840, N3579);
and AND3 (N9000, N8998, N8202, N6217);
and AND4 (N9001, N8995, N5592, N4274, N2937);
or OR4 (N9002, N8991, N6560, N3151, N1494);
nor NOR4 (N9003, N9002, N8682, N782, N7162);
nand NAND3 (N9004, N9003, N6783, N4722);
nor NOR4 (N9005, N8996, N8401, N6917, N4266);
and AND3 (N9006, N8997, N4938, N1236);
xor XOR2 (N9007, N8979, N2062);
nor NOR4 (N9008, N8999, N3104, N4381, N1525);
or OR2 (N9009, N9005, N2742);
and AND2 (N9010, N8988, N4942);
nor NOR3 (N9011, N9001, N6439, N5425);
nand NAND2 (N9012, N8994, N5142);
and AND4 (N9013, N9008, N8869, N192, N648);
xor XOR2 (N9014, N9006, N5453);
nand NAND4 (N9015, N9000, N4166, N1668, N6138);
or OR2 (N9016, N8993, N5879);
xor XOR2 (N9017, N9009, N2588);
buf BUF1 (N9018, N9016);
and AND3 (N9019, N9017, N6896, N7191);
nor NOR4 (N9020, N9012, N3950, N7506, N7408);
nor NOR4 (N9021, N9015, N4706, N7479, N4859);
buf BUF1 (N9022, N9007);
nor NOR4 (N9023, N9011, N2545, N7794, N6931);
nor NOR4 (N9024, N9023, N3956, N1115, N5887);
nand NAND2 (N9025, N9018, N1079);
and AND2 (N9026, N9013, N4987);
nor NOR3 (N9027, N9004, N6893, N2377);
not NOT1 (N9028, N9014);
and AND3 (N9029, N9025, N8852, N5698);
nor NOR3 (N9030, N9024, N1446, N5346);
xor XOR2 (N9031, N9026, N2963);
not NOT1 (N9032, N9022);
nor NOR2 (N9033, N9019, N8926);
not NOT1 (N9034, N9027);
nand NAND4 (N9035, N9034, N8456, N6952, N3291);
xor XOR2 (N9036, N9010, N8635);
xor XOR2 (N9037, N9033, N4913);
or OR3 (N9038, N9029, N1965, N5679);
buf BUF1 (N9039, N9021);
or OR3 (N9040, N9035, N8979, N4257);
and AND3 (N9041, N9037, N3145, N7815);
nor NOR4 (N9042, N9028, N5778, N8617, N654);
and AND3 (N9043, N9020, N4598, N7735);
nand NAND4 (N9044, N9040, N5353, N8963, N5513);
not NOT1 (N9045, N9031);
nand NAND2 (N9046, N9043, N1385);
and AND2 (N9047, N9046, N489);
not NOT1 (N9048, N9041);
nand NAND3 (N9049, N9047, N4351, N1756);
nor NOR4 (N9050, N9048, N984, N6956, N4683);
nand NAND2 (N9051, N9039, N5033);
nand NAND4 (N9052, N9038, N7103, N5578, N2663);
buf BUF1 (N9053, N9042);
nor NOR2 (N9054, N9030, N4897);
nand NAND2 (N9055, N9051, N7946);
nor NOR2 (N9056, N9032, N6897);
nor NOR4 (N9057, N9056, N815, N5537, N4757);
nor NOR4 (N9058, N9053, N4018, N3316, N1438);
and AND2 (N9059, N9045, N2892);
buf BUF1 (N9060, N9055);
xor XOR2 (N9061, N9057, N5814);
nand NAND4 (N9062, N9036, N835, N5011, N3497);
not NOT1 (N9063, N9060);
or OR2 (N9064, N9054, N6618);
nor NOR4 (N9065, N9062, N7127, N3505, N823);
buf BUF1 (N9066, N9059);
nand NAND2 (N9067, N9058, N7862);
buf BUF1 (N9068, N9063);
or OR4 (N9069, N9052, N5630, N1879, N1691);
not NOT1 (N9070, N9068);
not NOT1 (N9071, N9044);
xor XOR2 (N9072, N9071, N7826);
and AND4 (N9073, N9050, N5592, N4539, N8281);
or OR4 (N9074, N9069, N4693, N7239, N5800);
xor XOR2 (N9075, N9061, N1768);
not NOT1 (N9076, N9066);
nand NAND3 (N9077, N9075, N4974, N4842);
and AND3 (N9078, N9076, N7698, N3657);
nand NAND2 (N9079, N9067, N3623);
buf BUF1 (N9080, N9077);
and AND4 (N9081, N9073, N3356, N3171, N356);
buf BUF1 (N9082, N9070);
or OR4 (N9083, N9065, N8529, N7169, N4371);
or OR4 (N9084, N9083, N3380, N6950, N1843);
buf BUF1 (N9085, N9081);
or OR3 (N9086, N9085, N3322, N4484);
nand NAND4 (N9087, N9078, N5779, N8913, N18);
not NOT1 (N9088, N9049);
and AND2 (N9089, N9080, N5866);
nand NAND4 (N9090, N9079, N7483, N692, N7116);
xor XOR2 (N9091, N9086, N2260);
xor XOR2 (N9092, N9087, N5936);
not NOT1 (N9093, N9064);
and AND3 (N9094, N9091, N641, N3709);
not NOT1 (N9095, N9082);
xor XOR2 (N9096, N9092, N6844);
and AND3 (N9097, N9096, N373, N7339);
buf BUF1 (N9098, N9095);
or OR4 (N9099, N9084, N5231, N4580, N5181);
xor XOR2 (N9100, N9074, N2176);
not NOT1 (N9101, N9099);
buf BUF1 (N9102, N9088);
buf BUF1 (N9103, N9101);
nand NAND4 (N9104, N9093, N4916, N4135, N4798);
nand NAND2 (N9105, N9072, N1044);
not NOT1 (N9106, N9100);
and AND2 (N9107, N9105, N2923);
buf BUF1 (N9108, N9103);
nand NAND4 (N9109, N9094, N7724, N8917, N1406);
or OR2 (N9110, N9089, N5032);
buf BUF1 (N9111, N9098);
nor NOR3 (N9112, N9106, N7183, N7894);
nor NOR4 (N9113, N9111, N1159, N1886, N4893);
and AND3 (N9114, N9110, N9002, N2503);
nor NOR3 (N9115, N9108, N7503, N6517);
buf BUF1 (N9116, N9109);
nor NOR3 (N9117, N9112, N4899, N1172);
and AND2 (N9118, N9107, N8848);
xor XOR2 (N9119, N9090, N8493);
not NOT1 (N9120, N9119);
or OR3 (N9121, N9102, N4419, N8318);
not NOT1 (N9122, N9117);
nor NOR2 (N9123, N9118, N6430);
xor XOR2 (N9124, N9114, N1641);
buf BUF1 (N9125, N9122);
and AND2 (N9126, N9116, N2369);
buf BUF1 (N9127, N9115);
xor XOR2 (N9128, N9126, N4840);
or OR3 (N9129, N9127, N3042, N4598);
nor NOR3 (N9130, N9113, N3288, N6856);
and AND2 (N9131, N9128, N7516);
nor NOR2 (N9132, N9125, N6906);
nor NOR4 (N9133, N9123, N6318, N1727, N8668);
xor XOR2 (N9134, N9097, N8527);
or OR2 (N9135, N9134, N43);
nor NOR3 (N9136, N9135, N3888, N4038);
nand NAND4 (N9137, N9129, N4632, N975, N3289);
nor NOR4 (N9138, N9132, N2640, N136, N5488);
nand NAND4 (N9139, N9130, N2283, N1852, N5499);
or OR3 (N9140, N9139, N5010, N2249);
and AND4 (N9141, N9140, N3221, N4883, N3948);
xor XOR2 (N9142, N9131, N8409);
not NOT1 (N9143, N9121);
or OR4 (N9144, N9120, N4352, N7252, N701);
not NOT1 (N9145, N9143);
not NOT1 (N9146, N9124);
buf BUF1 (N9147, N9133);
and AND3 (N9148, N9137, N5512, N8881);
not NOT1 (N9149, N9142);
and AND4 (N9150, N9145, N2651, N2158, N8713);
nand NAND4 (N9151, N9146, N8070, N4076, N581);
xor XOR2 (N9152, N9136, N2027);
buf BUF1 (N9153, N9152);
and AND2 (N9154, N9149, N3818);
buf BUF1 (N9155, N9154);
nand NAND2 (N9156, N9150, N1286);
buf BUF1 (N9157, N9156);
nand NAND2 (N9158, N9148, N6513);
buf BUF1 (N9159, N9157);
and AND2 (N9160, N9155, N460);
or OR4 (N9161, N9151, N702, N7050, N1816);
nand NAND3 (N9162, N9159, N7510, N1756);
not NOT1 (N9163, N9160);
buf BUF1 (N9164, N9163);
or OR4 (N9165, N9161, N8595, N3507, N9100);
xor XOR2 (N9166, N9158, N4465);
or OR3 (N9167, N9141, N5400, N7696);
xor XOR2 (N9168, N9167, N6580);
xor XOR2 (N9169, N9144, N8450);
not NOT1 (N9170, N9153);
buf BUF1 (N9171, N9169);
xor XOR2 (N9172, N9104, N5);
or OR4 (N9173, N9147, N8094, N7469, N1871);
nand NAND2 (N9174, N9172, N3501);
buf BUF1 (N9175, N9164);
not NOT1 (N9176, N9138);
or OR2 (N9177, N9173, N3122);
nor NOR3 (N9178, N9166, N6564, N3144);
not NOT1 (N9179, N9175);
or OR3 (N9180, N9165, N2864, N3054);
buf BUF1 (N9181, N9170);
or OR2 (N9182, N9180, N5813);
buf BUF1 (N9183, N9182);
and AND4 (N9184, N9162, N6127, N7218, N511);
or OR3 (N9185, N9184, N3299, N3633);
and AND3 (N9186, N9183, N3933, N6257);
xor XOR2 (N9187, N9185, N4325);
and AND4 (N9188, N9174, N4967, N8678, N1112);
buf BUF1 (N9189, N9171);
xor XOR2 (N9190, N9189, N4571);
nor NOR2 (N9191, N9179, N3757);
buf BUF1 (N9192, N9177);
buf BUF1 (N9193, N9190);
not NOT1 (N9194, N9176);
and AND4 (N9195, N9193, N1003, N6987, N8230);
xor XOR2 (N9196, N9188, N8658);
nor NOR3 (N9197, N9192, N753, N5513);
or OR3 (N9198, N9186, N1717, N4124);
not NOT1 (N9199, N9187);
xor XOR2 (N9200, N9191, N6726);
xor XOR2 (N9201, N9181, N5218);
and AND3 (N9202, N9197, N6745, N41);
xor XOR2 (N9203, N9178, N8319);
and AND4 (N9204, N9200, N1559, N121, N4051);
and AND4 (N9205, N9195, N3675, N8066, N1998);
and AND3 (N9206, N9201, N2054, N2213);
nand NAND2 (N9207, N9202, N7800);
or OR3 (N9208, N9205, N426, N3567);
buf BUF1 (N9209, N9199);
nor NOR3 (N9210, N9196, N5950, N6472);
and AND3 (N9211, N9209, N8686, N4122);
buf BUF1 (N9212, N9207);
buf BUF1 (N9213, N9212);
not NOT1 (N9214, N9213);
nor NOR4 (N9215, N9194, N9001, N3599, N7453);
or OR2 (N9216, N9204, N7043);
nand NAND2 (N9217, N9168, N8783);
not NOT1 (N9218, N9216);
nor NOR4 (N9219, N9203, N2720, N5027, N779);
buf BUF1 (N9220, N9198);
nand NAND4 (N9221, N9210, N1891, N1671, N7073);
or OR3 (N9222, N9221, N361, N7499);
nor NOR3 (N9223, N9215, N6913, N4614);
xor XOR2 (N9224, N9208, N6033);
and AND3 (N9225, N9222, N4396, N7787);
xor XOR2 (N9226, N9214, N2461);
or OR4 (N9227, N9206, N7485, N3227, N8595);
nor NOR3 (N9228, N9226, N3972, N165);
or OR2 (N9229, N9219, N1642);
nand NAND4 (N9230, N9227, N5060, N4152, N2891);
nor NOR4 (N9231, N9217, N8252, N1976, N3479);
nand NAND2 (N9232, N9223, N5663);
nor NOR4 (N9233, N9231, N8952, N9116, N7333);
and AND4 (N9234, N9233, N6137, N5163, N4435);
buf BUF1 (N9235, N9220);
buf BUF1 (N9236, N9230);
not NOT1 (N9237, N9228);
xor XOR2 (N9238, N9211, N8650);
nor NOR2 (N9239, N9224, N5595);
nor NOR3 (N9240, N9229, N1311, N8794);
or OR4 (N9241, N9234, N7534, N938, N6110);
not NOT1 (N9242, N9218);
nand NAND2 (N9243, N9242, N5577);
buf BUF1 (N9244, N9236);
or OR3 (N9245, N9239, N1969, N1683);
nor NOR2 (N9246, N9225, N169);
and AND4 (N9247, N9246, N4069, N7185, N5771);
or OR2 (N9248, N9243, N9062);
or OR3 (N9249, N9241, N3124, N9019);
buf BUF1 (N9250, N9244);
nand NAND3 (N9251, N9247, N3831, N4104);
nor NOR4 (N9252, N9235, N4438, N5573, N8344);
buf BUF1 (N9253, N9251);
and AND2 (N9254, N9245, N5246);
nor NOR2 (N9255, N9249, N5971);
not NOT1 (N9256, N9250);
nor NOR3 (N9257, N9232, N2899, N4904);
not NOT1 (N9258, N9254);
nor NOR4 (N9259, N9253, N8516, N4685, N4045);
nor NOR2 (N9260, N9237, N159);
nor NOR4 (N9261, N9255, N8127, N2531, N2509);
and AND2 (N9262, N9256, N3383);
and AND2 (N9263, N9238, N2044);
buf BUF1 (N9264, N9248);
buf BUF1 (N9265, N9257);
or OR2 (N9266, N9261, N1376);
buf BUF1 (N9267, N9265);
nor NOR2 (N9268, N9266, N1229);
nand NAND3 (N9269, N9267, N3064, N2751);
not NOT1 (N9270, N9260);
xor XOR2 (N9271, N9259, N8713);
or OR4 (N9272, N9252, N8919, N983, N8176);
and AND3 (N9273, N9262, N1103, N4099);
xor XOR2 (N9274, N9269, N1374);
or OR3 (N9275, N9240, N8206, N856);
nor NOR2 (N9276, N9264, N1536);
nand NAND4 (N9277, N9268, N5335, N2126, N2321);
buf BUF1 (N9278, N9273);
and AND2 (N9279, N9258, N39);
not NOT1 (N9280, N9272);
or OR3 (N9281, N9277, N7547, N4870);
buf BUF1 (N9282, N9271);
buf BUF1 (N9283, N9282);
and AND4 (N9284, N9263, N7420, N5426, N6814);
nand NAND3 (N9285, N9270, N1170, N7438);
not NOT1 (N9286, N9280);
buf BUF1 (N9287, N9284);
buf BUF1 (N9288, N9281);
nor NOR3 (N9289, N9275, N2102, N85);
and AND2 (N9290, N9274, N1067);
or OR2 (N9291, N9289, N4862);
nand NAND2 (N9292, N9278, N7300);
nand NAND4 (N9293, N9292, N1685, N7191, N7766);
and AND3 (N9294, N9290, N276, N8868);
buf BUF1 (N9295, N9283);
and AND4 (N9296, N9285, N564, N9126, N5783);
and AND2 (N9297, N9279, N7802);
nor NOR2 (N9298, N9286, N5343);
nand NAND2 (N9299, N9296, N8686);
nor NOR3 (N9300, N9294, N2420, N174);
buf BUF1 (N9301, N9295);
buf BUF1 (N9302, N9291);
nand NAND3 (N9303, N9288, N2650, N209);
and AND4 (N9304, N9287, N6844, N14, N8154);
xor XOR2 (N9305, N9304, N18);
not NOT1 (N9306, N9293);
nor NOR4 (N9307, N9298, N6785, N1517, N6551);
not NOT1 (N9308, N9303);
and AND2 (N9309, N9306, N2876);
nand NAND4 (N9310, N9308, N8713, N1085, N2310);
or OR2 (N9311, N9302, N4246);
or OR2 (N9312, N9276, N8390);
nand NAND2 (N9313, N9300, N1297);
nand NAND4 (N9314, N9301, N1562, N4231, N7607);
or OR2 (N9315, N9309, N6455);
not NOT1 (N9316, N9315);
xor XOR2 (N9317, N9310, N262);
not NOT1 (N9318, N9313);
not NOT1 (N9319, N9299);
not NOT1 (N9320, N9305);
and AND2 (N9321, N9307, N6423);
not NOT1 (N9322, N9320);
not NOT1 (N9323, N9321);
and AND2 (N9324, N9297, N555);
xor XOR2 (N9325, N9314, N8574);
not NOT1 (N9326, N9312);
or OR3 (N9327, N9325, N1135, N8325);
nand NAND2 (N9328, N9326, N5759);
not NOT1 (N9329, N9323);
or OR3 (N9330, N9328, N5098, N9041);
nand NAND3 (N9331, N9330, N8495, N276);
not NOT1 (N9332, N9318);
not NOT1 (N9333, N9311);
not NOT1 (N9334, N9333);
or OR3 (N9335, N9324, N1736, N1329);
not NOT1 (N9336, N9335);
buf BUF1 (N9337, N9319);
or OR3 (N9338, N9334, N889, N9217);
buf BUF1 (N9339, N9322);
and AND3 (N9340, N9336, N9234, N4303);
buf BUF1 (N9341, N9339);
nand NAND2 (N9342, N9332, N9174);
xor XOR2 (N9343, N9337, N153);
xor XOR2 (N9344, N9316, N7408);
or OR2 (N9345, N9338, N1162);
not NOT1 (N9346, N9317);
and AND4 (N9347, N9342, N5192, N1754, N3041);
and AND3 (N9348, N9347, N8494, N6808);
and AND4 (N9349, N9345, N2680, N5340, N7176);
buf BUF1 (N9350, N9346);
and AND2 (N9351, N9341, N373);
xor XOR2 (N9352, N9327, N2236);
nor NOR2 (N9353, N9352, N747);
or OR3 (N9354, N9344, N6524, N1574);
buf BUF1 (N9355, N9343);
nand NAND2 (N9356, N9331, N127);
and AND2 (N9357, N9353, N5065);
and AND4 (N9358, N9340, N5623, N7801, N3291);
or OR4 (N9359, N9349, N6228, N6344, N8716);
and AND2 (N9360, N9350, N4028);
nand NAND4 (N9361, N9348, N1215, N5657, N3278);
nor NOR2 (N9362, N9356, N1473);
buf BUF1 (N9363, N9360);
or OR3 (N9364, N9329, N2502, N8811);
buf BUF1 (N9365, N9354);
buf BUF1 (N9366, N9358);
nand NAND4 (N9367, N9355, N4213, N4951, N6654);
or OR3 (N9368, N9362, N3013, N4057);
or OR2 (N9369, N9368, N4855);
and AND3 (N9370, N9369, N947, N157);
xor XOR2 (N9371, N9370, N5755);
nor NOR2 (N9372, N9371, N2442);
xor XOR2 (N9373, N9357, N9018);
xor XOR2 (N9374, N9365, N5599);
or OR2 (N9375, N9363, N5881);
not NOT1 (N9376, N9359);
nor NOR3 (N9377, N9373, N6194, N3120);
nor NOR3 (N9378, N9372, N1593, N602);
or OR3 (N9379, N9376, N6483, N2918);
nor NOR3 (N9380, N9377, N73, N8797);
buf BUF1 (N9381, N9379);
nand NAND3 (N9382, N9374, N2923, N3688);
nand NAND3 (N9383, N9375, N8957, N8159);
nor NOR4 (N9384, N9383, N7889, N7104, N7931);
or OR2 (N9385, N9361, N6865);
xor XOR2 (N9386, N9351, N9023);
nand NAND4 (N9387, N9385, N7031, N6620, N9290);
and AND2 (N9388, N9378, N8054);
buf BUF1 (N9389, N9382);
nor NOR3 (N9390, N9367, N1628, N9342);
not NOT1 (N9391, N9386);
xor XOR2 (N9392, N9390, N4542);
nand NAND2 (N9393, N9387, N7568);
nor NOR2 (N9394, N9381, N5234);
or OR4 (N9395, N9392, N8487, N481, N773);
nand NAND2 (N9396, N9394, N2696);
or OR3 (N9397, N9396, N9240, N474);
nor NOR3 (N9398, N9393, N2542, N7642);
xor XOR2 (N9399, N9366, N8901);
xor XOR2 (N9400, N9391, N7404);
and AND3 (N9401, N9388, N2210, N742);
not NOT1 (N9402, N9400);
nand NAND2 (N9403, N9395, N1000);
and AND4 (N9404, N9401, N1200, N8228, N5907);
nor NOR4 (N9405, N9389, N1406, N5220, N4542);
or OR2 (N9406, N9398, N7595);
xor XOR2 (N9407, N9384, N3239);
and AND2 (N9408, N9364, N5417);
nand NAND3 (N9409, N9404, N4634, N7698);
xor XOR2 (N9410, N9403, N6169);
nor NOR2 (N9411, N9402, N5834);
and AND4 (N9412, N9409, N2290, N1058, N5633);
and AND4 (N9413, N9408, N2353, N3108, N7065);
xor XOR2 (N9414, N9399, N7533);
nand NAND4 (N9415, N9380, N8498, N3856, N9340);
not NOT1 (N9416, N9411);
nor NOR2 (N9417, N9405, N8850);
nand NAND4 (N9418, N9416, N8552, N272, N8956);
nand NAND2 (N9419, N9413, N5781);
not NOT1 (N9420, N9417);
and AND4 (N9421, N9412, N6603, N8912, N3982);
nor NOR3 (N9422, N9419, N348, N5320);
nor NOR3 (N9423, N9406, N3124, N8111);
buf BUF1 (N9424, N9422);
buf BUF1 (N9425, N9410);
buf BUF1 (N9426, N9423);
nand NAND2 (N9427, N9424, N2363);
xor XOR2 (N9428, N9397, N1937);
xor XOR2 (N9429, N9428, N6057);
or OR4 (N9430, N9429, N4328, N2409, N4042);
or OR3 (N9431, N9426, N1628, N277);
and AND3 (N9432, N9420, N7573, N1085);
and AND3 (N9433, N9431, N1402, N7032);
and AND2 (N9434, N9430, N7010);
nand NAND3 (N9435, N9415, N7754, N5333);
and AND4 (N9436, N9434, N711, N9334, N1806);
nor NOR3 (N9437, N9418, N950, N6639);
nor NOR4 (N9438, N9421, N3874, N8668, N1323);
buf BUF1 (N9439, N9436);
not NOT1 (N9440, N9414);
not NOT1 (N9441, N9439);
not NOT1 (N9442, N9433);
not NOT1 (N9443, N9441);
or OR4 (N9444, N9425, N6926, N9361, N8230);
or OR4 (N9445, N9407, N7862, N5999, N4293);
xor XOR2 (N9446, N9442, N1276);
buf BUF1 (N9447, N9446);
buf BUF1 (N9448, N9435);
buf BUF1 (N9449, N9444);
xor XOR2 (N9450, N9448, N8572);
nand NAND3 (N9451, N9449, N7197, N6082);
xor XOR2 (N9452, N9443, N5975);
and AND4 (N9453, N9445, N1689, N3891, N5345);
not NOT1 (N9454, N9453);
nor NOR3 (N9455, N9447, N1119, N6735);
xor XOR2 (N9456, N9427, N7818);
not NOT1 (N9457, N9440);
nand NAND2 (N9458, N9457, N7719);
nand NAND4 (N9459, N9432, N3656, N9080, N8582);
nand NAND3 (N9460, N9438, N1568, N7294);
nand NAND4 (N9461, N9437, N817, N954, N5194);
nand NAND2 (N9462, N9461, N2904);
and AND4 (N9463, N9462, N1701, N3115, N7907);
nor NOR2 (N9464, N9451, N3227);
and AND4 (N9465, N9450, N6437, N5737, N1408);
or OR3 (N9466, N9463, N3561, N5526);
buf BUF1 (N9467, N9452);
not NOT1 (N9468, N9454);
buf BUF1 (N9469, N9456);
and AND4 (N9470, N9465, N6173, N3697, N3012);
xor XOR2 (N9471, N9464, N9030);
and AND3 (N9472, N9467, N9125, N86);
and AND2 (N9473, N9468, N509);
or OR3 (N9474, N9466, N2717, N554);
nor NOR2 (N9475, N9458, N1259);
nor NOR4 (N9476, N9475, N3990, N6433, N4926);
nand NAND3 (N9477, N9474, N7909, N3599);
nand NAND3 (N9478, N9470, N8569, N2568);
buf BUF1 (N9479, N9459);
or OR4 (N9480, N9471, N8743, N7420, N6146);
xor XOR2 (N9481, N9469, N2426);
buf BUF1 (N9482, N9455);
nand NAND3 (N9483, N9477, N8341, N182);
nand NAND4 (N9484, N9482, N472, N8276, N3182);
nor NOR3 (N9485, N9473, N6032, N1910);
buf BUF1 (N9486, N9479);
buf BUF1 (N9487, N9480);
xor XOR2 (N9488, N9483, N3932);
xor XOR2 (N9489, N9485, N1492);
nand NAND2 (N9490, N9472, N3206);
and AND2 (N9491, N9490, N9077);
xor XOR2 (N9492, N9491, N2294);
not NOT1 (N9493, N9492);
not NOT1 (N9494, N9481);
xor XOR2 (N9495, N9493, N874);
nand NAND2 (N9496, N9495, N5384);
buf BUF1 (N9497, N9476);
nor NOR4 (N9498, N9497, N8082, N9111, N1717);
xor XOR2 (N9499, N9496, N5377);
not NOT1 (N9500, N9499);
and AND3 (N9501, N9478, N2528, N1936);
or OR2 (N9502, N9501, N1638);
and AND2 (N9503, N9500, N4885);
xor XOR2 (N9504, N9488, N7217);
buf BUF1 (N9505, N9489);
nand NAND2 (N9506, N9484, N5036);
nor NOR2 (N9507, N9504, N4826);
xor XOR2 (N9508, N9506, N2069);
buf BUF1 (N9509, N9487);
buf BUF1 (N9510, N9486);
buf BUF1 (N9511, N9498);
nand NAND3 (N9512, N9511, N8675, N1156);
nor NOR4 (N9513, N9508, N7350, N1825, N6441);
or OR2 (N9514, N9494, N7115);
nand NAND4 (N9515, N9507, N8698, N3950, N541);
nand NAND3 (N9516, N9505, N6057, N9395);
and AND3 (N9517, N9513, N198, N4382);
nor NOR2 (N9518, N9514, N4807);
buf BUF1 (N9519, N9503);
and AND2 (N9520, N9510, N3434);
or OR4 (N9521, N9502, N7841, N8867, N4666);
nor NOR3 (N9522, N9520, N3390, N7843);
xor XOR2 (N9523, N9521, N1015);
and AND2 (N9524, N9517, N1938);
not NOT1 (N9525, N9523);
xor XOR2 (N9526, N9519, N7909);
and AND2 (N9527, N9526, N7682);
or OR4 (N9528, N9512, N5859, N1786, N5931);
and AND2 (N9529, N9460, N7768);
nand NAND3 (N9530, N9524, N1784, N40);
and AND3 (N9531, N9509, N2374, N7743);
or OR2 (N9532, N9531, N3963);
nand NAND3 (N9533, N9525, N2396, N524);
and AND2 (N9534, N9522, N7830);
nor NOR4 (N9535, N9515, N3271, N3514, N4369);
nand NAND2 (N9536, N9527, N8964);
nand NAND4 (N9537, N9532, N1781, N8373, N235);
not NOT1 (N9538, N9530);
or OR4 (N9539, N9535, N1451, N7020, N6552);
nand NAND2 (N9540, N9538, N3505);
nor NOR3 (N9541, N9528, N7715, N123);
xor XOR2 (N9542, N9518, N9028);
xor XOR2 (N9543, N9534, N7564);
and AND3 (N9544, N9516, N3032, N1492);
nand NAND3 (N9545, N9537, N1510, N2779);
or OR3 (N9546, N9545, N8293, N582);
nand NAND2 (N9547, N9540, N2060);
xor XOR2 (N9548, N9542, N2050);
xor XOR2 (N9549, N9544, N458);
xor XOR2 (N9550, N9533, N7538);
not NOT1 (N9551, N9536);
nand NAND2 (N9552, N9548, N4817);
not NOT1 (N9553, N9546);
buf BUF1 (N9554, N9543);
nor NOR4 (N9555, N9539, N8447, N5883, N4319);
and AND4 (N9556, N9551, N2101, N3609, N3685);
nand NAND2 (N9557, N9552, N6649);
xor XOR2 (N9558, N9541, N8289);
and AND3 (N9559, N9547, N5944, N1826);
not NOT1 (N9560, N9550);
and AND2 (N9561, N9529, N290);
or OR3 (N9562, N9554, N7177, N713);
nand NAND2 (N9563, N9561, N7214);
or OR4 (N9564, N9549, N7303, N5961, N5180);
buf BUF1 (N9565, N9560);
not NOT1 (N9566, N9557);
and AND4 (N9567, N9566, N2665, N8344, N1711);
and AND2 (N9568, N9555, N971);
and AND3 (N9569, N9565, N4599, N7427);
xor XOR2 (N9570, N9567, N1949);
buf BUF1 (N9571, N9556);
nand NAND3 (N9572, N9571, N999, N8069);
nor NOR2 (N9573, N9562, N2037);
or OR2 (N9574, N9572, N3462);
not NOT1 (N9575, N9559);
xor XOR2 (N9576, N9570, N5452);
not NOT1 (N9577, N9568);
and AND4 (N9578, N9558, N5884, N365, N1326);
not NOT1 (N9579, N9577);
not NOT1 (N9580, N9563);
or OR4 (N9581, N9575, N7336, N3255, N420);
xor XOR2 (N9582, N9579, N298);
xor XOR2 (N9583, N9580, N7856);
or OR3 (N9584, N9574, N5776, N4842);
buf BUF1 (N9585, N9573);
buf BUF1 (N9586, N9585);
buf BUF1 (N9587, N9586);
nor NOR2 (N9588, N9553, N7040);
nand NAND2 (N9589, N9581, N8815);
not NOT1 (N9590, N9564);
xor XOR2 (N9591, N9582, N5197);
not NOT1 (N9592, N9584);
xor XOR2 (N9593, N9589, N3420);
buf BUF1 (N9594, N9588);
xor XOR2 (N9595, N9591, N3946);
and AND2 (N9596, N9595, N7979);
xor XOR2 (N9597, N9578, N5575);
xor XOR2 (N9598, N9597, N8598);
not NOT1 (N9599, N9569);
not NOT1 (N9600, N9596);
xor XOR2 (N9601, N9587, N200);
nor NOR4 (N9602, N9593, N45, N4198, N8168);
or OR2 (N9603, N9590, N4018);
nand NAND2 (N9604, N9592, N5281);
and AND4 (N9605, N9604, N4386, N3828, N7938);
not NOT1 (N9606, N9602);
nor NOR3 (N9607, N9583, N4299, N5593);
nor NOR4 (N9608, N9606, N4725, N2019, N4489);
nand NAND4 (N9609, N9603, N9378, N95, N5220);
and AND3 (N9610, N9601, N4063, N8492);
xor XOR2 (N9611, N9576, N6038);
xor XOR2 (N9612, N9609, N3996);
or OR2 (N9613, N9607, N649);
buf BUF1 (N9614, N9612);
xor XOR2 (N9615, N9611, N5710);
buf BUF1 (N9616, N9615);
not NOT1 (N9617, N9605);
or OR4 (N9618, N9599, N5861, N1934, N8756);
nand NAND4 (N9619, N9598, N9417, N392, N3128);
and AND2 (N9620, N9600, N6475);
and AND2 (N9621, N9610, N6840);
and AND3 (N9622, N9608, N1795, N3844);
or OR3 (N9623, N9614, N2848, N811);
nand NAND4 (N9624, N9622, N8554, N9189, N1694);
and AND4 (N9625, N9613, N711, N421, N1852);
buf BUF1 (N9626, N9623);
nor NOR4 (N9627, N9625, N6974, N7317, N5246);
nor NOR4 (N9628, N9619, N2260, N819, N4273);
buf BUF1 (N9629, N9616);
or OR4 (N9630, N9626, N5609, N2890, N6912);
buf BUF1 (N9631, N9621);
and AND4 (N9632, N9620, N4568, N5734, N627);
xor XOR2 (N9633, N9629, N2506);
buf BUF1 (N9634, N9618);
xor XOR2 (N9635, N9633, N1881);
and AND2 (N9636, N9617, N8401);
nor NOR4 (N9637, N9594, N9051, N5935, N1037);
nor NOR3 (N9638, N9635, N253, N1822);
not NOT1 (N9639, N9630);
nor NOR3 (N9640, N9624, N1682, N746);
nand NAND3 (N9641, N9632, N9065, N8567);
or OR4 (N9642, N9639, N4841, N4202, N4105);
buf BUF1 (N9643, N9641);
or OR4 (N9644, N9627, N6896, N3281, N1581);
or OR3 (N9645, N9642, N8079, N3579);
and AND2 (N9646, N9628, N298);
or OR2 (N9647, N9631, N8985);
nor NOR3 (N9648, N9637, N6298, N9616);
nor NOR4 (N9649, N9634, N5648, N6365, N7250);
and AND3 (N9650, N9640, N9455, N7971);
nor NOR2 (N9651, N9647, N8298);
not NOT1 (N9652, N9638);
and AND2 (N9653, N9648, N7901);
or OR2 (N9654, N9650, N2019);
nand NAND4 (N9655, N9636, N784, N1141, N2579);
xor XOR2 (N9656, N9655, N1657);
buf BUF1 (N9657, N9654);
xor XOR2 (N9658, N9653, N1715);
not NOT1 (N9659, N9646);
not NOT1 (N9660, N9657);
buf BUF1 (N9661, N9659);
buf BUF1 (N9662, N9645);
and AND4 (N9663, N9643, N7853, N4882, N3656);
and AND3 (N9664, N9658, N7318, N5103);
or OR2 (N9665, N9660, N8825);
nor NOR2 (N9666, N9662, N6564);
not NOT1 (N9667, N9656);
xor XOR2 (N9668, N9649, N1557);
xor XOR2 (N9669, N9664, N6374);
or OR4 (N9670, N9666, N5599, N9618, N9143);
or OR4 (N9671, N9652, N488, N9568, N2015);
xor XOR2 (N9672, N9669, N4301);
not NOT1 (N9673, N9667);
nor NOR3 (N9674, N9665, N1382, N7888);
not NOT1 (N9675, N9668);
xor XOR2 (N9676, N9675, N3326);
or OR3 (N9677, N9671, N1855, N7346);
nor NOR4 (N9678, N9676, N5349, N167, N3809);
not NOT1 (N9679, N9677);
and AND3 (N9680, N9661, N1252, N1456);
and AND4 (N9681, N9678, N8644, N3518, N3124);
xor XOR2 (N9682, N9679, N8807);
buf BUF1 (N9683, N9681);
nand NAND2 (N9684, N9663, N6376);
and AND4 (N9685, N9680, N8295, N4578, N9176);
nand NAND3 (N9686, N9684, N6330, N4004);
nand NAND2 (N9687, N9682, N3065);
xor XOR2 (N9688, N9687, N929);
or OR4 (N9689, N9688, N6381, N4439, N9393);
buf BUF1 (N9690, N9689);
and AND3 (N9691, N9670, N7595, N9612);
nand NAND4 (N9692, N9673, N4546, N1623, N1923);
xor XOR2 (N9693, N9651, N4099);
xor XOR2 (N9694, N9686, N9281);
buf BUF1 (N9695, N9693);
and AND3 (N9696, N9691, N8879, N8277);
xor XOR2 (N9697, N9685, N7273);
xor XOR2 (N9698, N9683, N6203);
buf BUF1 (N9699, N9692);
nor NOR4 (N9700, N9674, N1757, N5574, N8085);
not NOT1 (N9701, N9698);
nand NAND4 (N9702, N9699, N7612, N2612, N1481);
xor XOR2 (N9703, N9702, N5389);
nor NOR2 (N9704, N9690, N3552);
not NOT1 (N9705, N9672);
nand NAND2 (N9706, N9697, N6532);
nor NOR3 (N9707, N9700, N990, N3260);
xor XOR2 (N9708, N9694, N1289);
not NOT1 (N9709, N9696);
xor XOR2 (N9710, N9703, N2046);
xor XOR2 (N9711, N9701, N5174);
or OR4 (N9712, N9706, N3030, N3403, N4947);
or OR3 (N9713, N9710, N8762, N9375);
not NOT1 (N9714, N9708);
not NOT1 (N9715, N9709);
not NOT1 (N9716, N9712);
and AND2 (N9717, N9716, N6874);
nor NOR4 (N9718, N9717, N8050, N5496, N4658);
nand NAND4 (N9719, N9704, N5853, N6055, N5800);
not NOT1 (N9720, N9714);
buf BUF1 (N9721, N9707);
nand NAND4 (N9722, N9715, N1605, N2084, N6798);
and AND3 (N9723, N9644, N3620, N4040);
and AND3 (N9724, N9705, N2328, N3707);
buf BUF1 (N9725, N9721);
not NOT1 (N9726, N9711);
nor NOR2 (N9727, N9723, N8703);
buf BUF1 (N9728, N9718);
and AND2 (N9729, N9722, N4607);
and AND4 (N9730, N9724, N765, N7059, N6545);
not NOT1 (N9731, N9725);
not NOT1 (N9732, N9730);
or OR2 (N9733, N9720, N3363);
nand NAND3 (N9734, N9719, N8823, N5391);
or OR3 (N9735, N9728, N574, N6962);
or OR3 (N9736, N9727, N7676, N8897);
not NOT1 (N9737, N9695);
or OR3 (N9738, N9731, N242, N6729);
nand NAND3 (N9739, N9713, N6718, N632);
xor XOR2 (N9740, N9732, N9321);
not NOT1 (N9741, N9736);
nand NAND2 (N9742, N9735, N1488);
and AND3 (N9743, N9737, N3326, N4834);
nor NOR2 (N9744, N9739, N3981);
not NOT1 (N9745, N9734);
and AND2 (N9746, N9742, N5774);
nor NOR2 (N9747, N9746, N5526);
buf BUF1 (N9748, N9747);
not NOT1 (N9749, N9729);
buf BUF1 (N9750, N9745);
not NOT1 (N9751, N9738);
buf BUF1 (N9752, N9741);
nand NAND2 (N9753, N9751, N808);
not NOT1 (N9754, N9749);
buf BUF1 (N9755, N9743);
not NOT1 (N9756, N9740);
not NOT1 (N9757, N9726);
xor XOR2 (N9758, N9752, N4319);
xor XOR2 (N9759, N9756, N2772);
and AND2 (N9760, N9753, N3272);
buf BUF1 (N9761, N9755);
not NOT1 (N9762, N9758);
and AND3 (N9763, N9750, N182, N8293);
not NOT1 (N9764, N9748);
and AND3 (N9765, N9761, N2836, N3924);
not NOT1 (N9766, N9754);
xor XOR2 (N9767, N9733, N1600);
not NOT1 (N9768, N9767);
nand NAND4 (N9769, N9768, N3528, N2582, N2318);
xor XOR2 (N9770, N9759, N9420);
xor XOR2 (N9771, N9757, N6613);
nand NAND4 (N9772, N9760, N1491, N4353, N1881);
nand NAND4 (N9773, N9769, N4144, N5119, N2975);
nor NOR4 (N9774, N9763, N1743, N5442, N6740);
xor XOR2 (N9775, N9744, N5294);
nor NOR2 (N9776, N9774, N1334);
and AND4 (N9777, N9776, N4049, N4075, N1973);
nand NAND2 (N9778, N9764, N8134);
nor NOR4 (N9779, N9775, N2323, N1915, N1199);
buf BUF1 (N9780, N9779);
buf BUF1 (N9781, N9777);
or OR2 (N9782, N9771, N7708);
or OR2 (N9783, N9781, N5384);
and AND2 (N9784, N9766, N8982);
not NOT1 (N9785, N9772);
and AND4 (N9786, N9784, N610, N1671, N2662);
nor NOR3 (N9787, N9783, N8359, N4875);
nor NOR4 (N9788, N9780, N962, N228, N4333);
or OR2 (N9789, N9773, N2678);
xor XOR2 (N9790, N9786, N1066);
not NOT1 (N9791, N9790);
xor XOR2 (N9792, N9782, N3041);
xor XOR2 (N9793, N9791, N9342);
not NOT1 (N9794, N9785);
buf BUF1 (N9795, N9794);
or OR3 (N9796, N9762, N3297, N6082);
nor NOR4 (N9797, N9792, N769, N8104, N3844);
buf BUF1 (N9798, N9788);
and AND2 (N9799, N9789, N9261);
buf BUF1 (N9800, N9765);
xor XOR2 (N9801, N9800, N146);
nor NOR2 (N9802, N9778, N729);
and AND3 (N9803, N9795, N5493, N3974);
or OR2 (N9804, N9787, N3025);
not NOT1 (N9805, N9804);
and AND2 (N9806, N9801, N8562);
xor XOR2 (N9807, N9796, N2974);
buf BUF1 (N9808, N9806);
nor NOR3 (N9809, N9793, N621, N9735);
nor NOR3 (N9810, N9770, N1044, N5622);
nand NAND3 (N9811, N9799, N3681, N8096);
nor NOR4 (N9812, N9797, N2718, N3405, N9354);
buf BUF1 (N9813, N9805);
not NOT1 (N9814, N9811);
not NOT1 (N9815, N9814);
and AND2 (N9816, N9808, N8123);
and AND4 (N9817, N9813, N9643, N8400, N4044);
nand NAND4 (N9818, N9803, N4587, N3965, N161);
nor NOR2 (N9819, N9812, N9199);
buf BUF1 (N9820, N9818);
nor NOR2 (N9821, N9809, N5559);
or OR2 (N9822, N9810, N2430);
nor NOR3 (N9823, N9802, N5072, N4214);
nand NAND2 (N9824, N9815, N874);
or OR3 (N9825, N9816, N5940, N5686);
not NOT1 (N9826, N9798);
nor NOR4 (N9827, N9825, N3396, N3996, N1203);
and AND4 (N9828, N9824, N7320, N5596, N9603);
buf BUF1 (N9829, N9822);
buf BUF1 (N9830, N9817);
nor NOR4 (N9831, N9820, N3371, N7273, N4228);
buf BUF1 (N9832, N9807);
or OR2 (N9833, N9819, N7461);
nor NOR2 (N9834, N9828, N4451);
nand NAND4 (N9835, N9831, N2558, N2689, N5596);
and AND4 (N9836, N9821, N8899, N3125, N4519);
or OR2 (N9837, N9823, N7070);
or OR3 (N9838, N9833, N5945, N5466);
or OR3 (N9839, N9838, N9701, N1478);
xor XOR2 (N9840, N9835, N8358);
or OR3 (N9841, N9834, N9285, N7137);
xor XOR2 (N9842, N9837, N1053);
xor XOR2 (N9843, N9826, N8782);
not NOT1 (N9844, N9843);
xor XOR2 (N9845, N9839, N3992);
or OR3 (N9846, N9842, N1370, N4072);
or OR3 (N9847, N9841, N8490, N4532);
not NOT1 (N9848, N9832);
nand NAND4 (N9849, N9847, N7071, N4168, N6666);
and AND3 (N9850, N9849, N5626, N8952);
xor XOR2 (N9851, N9844, N5985);
or OR3 (N9852, N9851, N8314, N4515);
or OR3 (N9853, N9850, N6785, N4283);
or OR3 (N9854, N9845, N7740, N5577);
and AND3 (N9855, N9854, N401, N3538);
or OR4 (N9856, N9827, N6654, N4148, N5264);
nand NAND4 (N9857, N9829, N2052, N5103, N7687);
and AND2 (N9858, N9856, N1527);
nor NOR4 (N9859, N9857, N3084, N4893, N2036);
not NOT1 (N9860, N9853);
nand NAND3 (N9861, N9855, N7911, N2648);
or OR2 (N9862, N9836, N8022);
nand NAND3 (N9863, N9860, N6510, N6166);
nand NAND2 (N9864, N9846, N5147);
xor XOR2 (N9865, N9864, N234);
or OR3 (N9866, N9830, N4778, N3537);
nor NOR2 (N9867, N9848, N7105);
xor XOR2 (N9868, N9859, N6357);
nor NOR4 (N9869, N9861, N3391, N383, N6897);
and AND2 (N9870, N9863, N176);
xor XOR2 (N9871, N9840, N9851);
xor XOR2 (N9872, N9868, N2930);
nor NOR4 (N9873, N9870, N2219, N236, N6707);
nor NOR4 (N9874, N9867, N3501, N9086, N2174);
xor XOR2 (N9875, N9873, N6396);
nand NAND4 (N9876, N9871, N3113, N7766, N1591);
and AND2 (N9877, N9866, N9829);
nand NAND3 (N9878, N9862, N6271, N6276);
nor NOR4 (N9879, N9872, N6746, N1227, N1018);
or OR3 (N9880, N9877, N8827, N996);
buf BUF1 (N9881, N9858);
buf BUF1 (N9882, N9878);
not NOT1 (N9883, N9852);
xor XOR2 (N9884, N9876, N8896);
buf BUF1 (N9885, N9874);
and AND3 (N9886, N9869, N7795, N1220);
not NOT1 (N9887, N9865);
buf BUF1 (N9888, N9879);
or OR3 (N9889, N9888, N74, N9657);
or OR3 (N9890, N9883, N6536, N8314);
buf BUF1 (N9891, N9881);
not NOT1 (N9892, N9889);
and AND4 (N9893, N9890, N432, N2070, N7882);
buf BUF1 (N9894, N9893);
xor XOR2 (N9895, N9875, N6321);
nand NAND4 (N9896, N9887, N2716, N1488, N2517);
not NOT1 (N9897, N9896);
or OR2 (N9898, N9892, N2192);
buf BUF1 (N9899, N9886);
buf BUF1 (N9900, N9885);
xor XOR2 (N9901, N9884, N270);
nand NAND3 (N9902, N9901, N411, N7621);
and AND3 (N9903, N9899, N6578, N7419);
and AND3 (N9904, N9894, N8517, N6621);
or OR4 (N9905, N9882, N7557, N1987, N5358);
buf BUF1 (N9906, N9905);
buf BUF1 (N9907, N9904);
xor XOR2 (N9908, N9903, N289);
not NOT1 (N9909, N9898);
not NOT1 (N9910, N9880);
nor NOR2 (N9911, N9902, N4309);
nand NAND3 (N9912, N9909, N2062, N3969);
or OR2 (N9913, N9906, N3515);
xor XOR2 (N9914, N9891, N6720);
xor XOR2 (N9915, N9907, N6244);
xor XOR2 (N9916, N9895, N4888);
not NOT1 (N9917, N9897);
and AND2 (N9918, N9912, N8273);
not NOT1 (N9919, N9910);
xor XOR2 (N9920, N9911, N4033);
nor NOR4 (N9921, N9920, N9646, N9060, N4770);
nand NAND3 (N9922, N9913, N7942, N5088);
and AND4 (N9923, N9921, N4285, N8456, N1778);
not NOT1 (N9924, N9919);
xor XOR2 (N9925, N9923, N4870);
or OR3 (N9926, N9916, N8655, N4776);
or OR4 (N9927, N9914, N1532, N1500, N9635);
not NOT1 (N9928, N9900);
xor XOR2 (N9929, N9917, N9897);
buf BUF1 (N9930, N9922);
not NOT1 (N9931, N9926);
not NOT1 (N9932, N9930);
and AND2 (N9933, N9932, N6079);
nand NAND2 (N9934, N9925, N1947);
not NOT1 (N9935, N9924);
xor XOR2 (N9936, N9935, N6992);
xor XOR2 (N9937, N9931, N4556);
or OR4 (N9938, N9908, N1731, N8495, N2732);
not NOT1 (N9939, N9936);
nor NOR3 (N9940, N9937, N4314, N8501);
nand NAND2 (N9941, N9929, N2792);
buf BUF1 (N9942, N9939);
nand NAND2 (N9943, N9934, N5075);
xor XOR2 (N9944, N9942, N6385);
nand NAND2 (N9945, N9943, N6923);
buf BUF1 (N9946, N9945);
or OR3 (N9947, N9941, N1423, N947);
or OR4 (N9948, N9946, N8768, N488, N8738);
nor NOR3 (N9949, N9927, N1148, N5432);
not NOT1 (N9950, N9918);
not NOT1 (N9951, N9915);
xor XOR2 (N9952, N9949, N3989);
not NOT1 (N9953, N9951);
and AND3 (N9954, N9933, N6305, N3283);
xor XOR2 (N9955, N9954, N7623);
nor NOR4 (N9956, N9947, N7955, N6717, N4470);
or OR4 (N9957, N9952, N5123, N3966, N1801);
or OR2 (N9958, N9956, N595);
or OR3 (N9959, N9938, N2212, N867);
nor NOR3 (N9960, N9957, N1717, N3839);
nand NAND4 (N9961, N9959, N7830, N9106, N9241);
nor NOR3 (N9962, N9944, N8256, N2690);
buf BUF1 (N9963, N9960);
and AND3 (N9964, N9950, N195, N598);
or OR4 (N9965, N9962, N7153, N730, N8410);
nand NAND2 (N9966, N9955, N376);
nor NOR2 (N9967, N9948, N4422);
nor NOR4 (N9968, N9966, N8043, N7091, N5455);
not NOT1 (N9969, N9968);
or OR4 (N9970, N9961, N7482, N762, N6384);
buf BUF1 (N9971, N9965);
nor NOR3 (N9972, N9940, N4336, N3313);
not NOT1 (N9973, N9967);
and AND4 (N9974, N9953, N4002, N7612, N6545);
xor XOR2 (N9975, N9972, N215);
buf BUF1 (N9976, N9964);
not NOT1 (N9977, N9963);
nand NAND3 (N9978, N9969, N8977, N566);
xor XOR2 (N9979, N9971, N4467);
buf BUF1 (N9980, N9979);
xor XOR2 (N9981, N9958, N8954);
nand NAND3 (N9982, N9975, N9073, N6275);
xor XOR2 (N9983, N9973, N3066);
nor NOR4 (N9984, N9983, N3390, N3491, N8667);
xor XOR2 (N9985, N9984, N3726);
xor XOR2 (N9986, N9976, N748);
or OR3 (N9987, N9970, N2732, N5136);
not NOT1 (N9988, N9987);
nor NOR4 (N9989, N9974, N6733, N5026, N1158);
and AND3 (N9990, N9985, N9252, N609);
nand NAND4 (N9991, N9981, N8633, N498, N2482);
nor NOR3 (N9992, N9989, N8164, N8852);
buf BUF1 (N9993, N9986);
or OR3 (N9994, N9990, N9528, N6507);
buf BUF1 (N9995, N9977);
nor NOR4 (N9996, N9995, N2826, N7368, N5462);
xor XOR2 (N9997, N9993, N2555);
or OR4 (N9998, N9992, N5690, N1528, N8117);
and AND3 (N9999, N9978, N9718, N1867);
not NOT1 (N10000, N9998);
not NOT1 (N10001, N9982);
buf BUF1 (N10002, N9988);
or OR2 (N10003, N10002, N9523);
buf BUF1 (N10004, N9997);
or OR4 (N10005, N9994, N4003, N1218, N6514);
nor NOR4 (N10006, N10005, N1926, N4990, N428);
xor XOR2 (N10007, N9999, N4420);
not NOT1 (N10008, N9928);
or OR3 (N10009, N10003, N1076, N923);
and AND2 (N10010, N10004, N2270);
or OR2 (N10011, N9991, N9695);
buf BUF1 (N10012, N10010);
nor NOR4 (N10013, N9996, N3191, N3794, N285);
nor NOR4 (N10014, N10007, N9024, N8057, N3361);
and AND4 (N10015, N10009, N1630, N8882, N1232);
xor XOR2 (N10016, N10015, N9998);
buf BUF1 (N10017, N10014);
not NOT1 (N10018, N10008);
buf BUF1 (N10019, N10017);
buf BUF1 (N10020, N10018);
and AND2 (N10021, N10000, N4227);
not NOT1 (N10022, N10006);
and AND3 (N10023, N10019, N6254, N6224);
and AND2 (N10024, N10011, N6311);
buf BUF1 (N10025, N10020);
and AND4 (N10026, N10012, N9143, N6793, N6654);
buf BUF1 (N10027, N10025);
not NOT1 (N10028, N10021);
nor NOR4 (N10029, N10026, N4015, N7002, N557);
nand NAND3 (N10030, N10027, N3419, N5818);
or OR3 (N10031, N10030, N2368, N1588);
buf BUF1 (N10032, N10022);
and AND2 (N10033, N10001, N8616);
nand NAND2 (N10034, N10032, N320);
or OR2 (N10035, N10034, N9567);
not NOT1 (N10036, N10013);
nand NAND4 (N10037, N10028, N3884, N8861, N8136);
and AND3 (N10038, N9980, N7633, N5911);
not NOT1 (N10039, N10036);
or OR4 (N10040, N10038, N6029, N5119, N213);
xor XOR2 (N10041, N10016, N9544);
and AND3 (N10042, N10033, N3253, N8829);
nand NAND3 (N10043, N10037, N6641, N2482);
nand NAND2 (N10044, N10039, N2879);
not NOT1 (N10045, N10040);
or OR2 (N10046, N10045, N8795);
not NOT1 (N10047, N10042);
and AND2 (N10048, N10029, N9386);
buf BUF1 (N10049, N10047);
and AND2 (N10050, N10048, N4678);
nand NAND3 (N10051, N10043, N9464, N7158);
nand NAND2 (N10052, N10046, N4449);
buf BUF1 (N10053, N10041);
xor XOR2 (N10054, N10023, N9084);
nand NAND2 (N10055, N10053, N1526);
and AND4 (N10056, N10054, N5343, N10004, N2554);
or OR2 (N10057, N10049, N4205);
not NOT1 (N10058, N10051);
nand NAND2 (N10059, N10050, N3393);
and AND3 (N10060, N10056, N9240, N1202);
buf BUF1 (N10061, N10031);
xor XOR2 (N10062, N10061, N8265);
and AND4 (N10063, N10052, N3697, N1282, N1607);
nand NAND3 (N10064, N10044, N4137, N2889);
and AND4 (N10065, N10057, N7507, N2760, N5414);
not NOT1 (N10066, N10055);
nand NAND4 (N10067, N10064, N8447, N3346, N3216);
not NOT1 (N10068, N10059);
nor NOR3 (N10069, N10068, N4997, N2583);
not NOT1 (N10070, N10067);
not NOT1 (N10071, N10070);
xor XOR2 (N10072, N10069, N2750);
xor XOR2 (N10073, N10035, N5457);
not NOT1 (N10074, N10065);
xor XOR2 (N10075, N10073, N5123);
or OR3 (N10076, N10060, N6797, N1953);
nand NAND3 (N10077, N10058, N708, N2073);
nand NAND2 (N10078, N10074, N8387);
nand NAND4 (N10079, N10063, N9874, N7626, N9494);
not NOT1 (N10080, N10062);
xor XOR2 (N10081, N10075, N7512);
xor XOR2 (N10082, N10078, N7009);
xor XOR2 (N10083, N10077, N258);
not NOT1 (N10084, N10071);
or OR4 (N10085, N10066, N8019, N481, N9484);
xor XOR2 (N10086, N10081, N4712);
xor XOR2 (N10087, N10084, N7440);
nor NOR4 (N10088, N10085, N4703, N74, N8633);
not NOT1 (N10089, N10080);
nand NAND3 (N10090, N10082, N5735, N2870);
xor XOR2 (N10091, N10089, N1452);
or OR3 (N10092, N10076, N9847, N1927);
nand NAND4 (N10093, N10079, N7298, N6610, N3415);
not NOT1 (N10094, N10088);
or OR3 (N10095, N10072, N2828, N421);
or OR2 (N10096, N10086, N1362);
and AND4 (N10097, N10094, N7568, N3296, N4447);
nor NOR4 (N10098, N10095, N9403, N7413, N6672);
buf BUF1 (N10099, N10096);
nor NOR4 (N10100, N10092, N9888, N769, N5505);
nand NAND3 (N10101, N10091, N3888, N1818);
nor NOR4 (N10102, N10083, N1020, N7644, N8397);
nor NOR4 (N10103, N10087, N7794, N5602, N9489);
or OR2 (N10104, N10101, N1676);
buf BUF1 (N10105, N10103);
buf BUF1 (N10106, N10100);
nand NAND2 (N10107, N10105, N7442);
or OR4 (N10108, N10107, N2562, N7733, N3137);
xor XOR2 (N10109, N10090, N5279);
xor XOR2 (N10110, N10106, N5277);
xor XOR2 (N10111, N10109, N9716);
buf BUF1 (N10112, N10110);
not NOT1 (N10113, N10024);
nor NOR4 (N10114, N10102, N6059, N9602, N6579);
not NOT1 (N10115, N10093);
not NOT1 (N10116, N10115);
xor XOR2 (N10117, N10098, N8003);
xor XOR2 (N10118, N10097, N2594);
not NOT1 (N10119, N10114);
nand NAND2 (N10120, N10117, N3033);
not NOT1 (N10121, N10118);
xor XOR2 (N10122, N10119, N7379);
and AND3 (N10123, N10108, N4265, N9264);
buf BUF1 (N10124, N10104);
nor NOR2 (N10125, N10123, N8240);
nand NAND4 (N10126, N10112, N1993, N10117, N8902);
nor NOR4 (N10127, N10126, N313, N9328, N668);
or OR2 (N10128, N10120, N9531);
or OR4 (N10129, N10121, N1477, N5200, N5459);
nand NAND4 (N10130, N10128, N6724, N4665, N4600);
or OR4 (N10131, N10124, N8556, N1060, N2235);
or OR3 (N10132, N10130, N2624, N9563);
buf BUF1 (N10133, N10131);
not NOT1 (N10134, N10127);
nor NOR3 (N10135, N10129, N6569, N4337);
nor NOR2 (N10136, N10113, N4132);
nor NOR2 (N10137, N10136, N5064);
buf BUF1 (N10138, N10135);
xor XOR2 (N10139, N10099, N2333);
nor NOR4 (N10140, N10116, N9130, N3621, N4122);
or OR4 (N10141, N10134, N9208, N5105, N2971);
nor NOR3 (N10142, N10133, N9816, N1655);
nor NOR4 (N10143, N10111, N7916, N9127, N2148);
xor XOR2 (N10144, N10141, N6495);
nand NAND3 (N10145, N10125, N5291, N8452);
not NOT1 (N10146, N10138);
nand NAND4 (N10147, N10122, N2419, N3375, N3925);
nor NOR2 (N10148, N10146, N2951);
nand NAND4 (N10149, N10137, N9411, N4274, N7273);
not NOT1 (N10150, N10143);
xor XOR2 (N10151, N10145, N202);
xor XOR2 (N10152, N10140, N3824);
not NOT1 (N10153, N10147);
nor NOR4 (N10154, N10148, N7827, N4723, N4706);
xor XOR2 (N10155, N10139, N3945);
buf BUF1 (N10156, N10149);
not NOT1 (N10157, N10154);
or OR2 (N10158, N10144, N6509);
or OR4 (N10159, N10156, N7387, N1028, N6122);
not NOT1 (N10160, N10159);
nand NAND3 (N10161, N10153, N552, N8794);
nor NOR2 (N10162, N10161, N3855);
nor NOR3 (N10163, N10158, N7822, N1973);
nor NOR3 (N10164, N10142, N443, N1831);
buf BUF1 (N10165, N10155);
nand NAND4 (N10166, N10165, N906, N8993, N8933);
and AND2 (N10167, N10157, N8206);
and AND2 (N10168, N10163, N8725);
or OR3 (N10169, N10166, N8254, N5994);
xor XOR2 (N10170, N10151, N4897);
and AND3 (N10171, N10132, N3088, N5692);
nand NAND3 (N10172, N10167, N8647, N1047);
and AND3 (N10173, N10170, N3474, N9718);
buf BUF1 (N10174, N10171);
or OR3 (N10175, N10172, N4798, N8533);
xor XOR2 (N10176, N10175, N8013);
nand NAND3 (N10177, N10160, N9879, N28);
nand NAND2 (N10178, N10150, N10044);
buf BUF1 (N10179, N10162);
or OR2 (N10180, N10177, N6482);
and AND4 (N10181, N10176, N1390, N1150, N3158);
nor NOR4 (N10182, N10168, N8211, N2967, N3532);
xor XOR2 (N10183, N10174, N6465);
or OR4 (N10184, N10164, N1482, N7508, N5971);
buf BUF1 (N10185, N10173);
nor NOR4 (N10186, N10185, N4071, N3511, N247);
not NOT1 (N10187, N10186);
not NOT1 (N10188, N10178);
nand NAND4 (N10189, N10180, N1642, N9653, N1321);
or OR2 (N10190, N10182, N12);
buf BUF1 (N10191, N10184);
nand NAND3 (N10192, N10187, N9465, N6372);
not NOT1 (N10193, N10179);
not NOT1 (N10194, N10188);
not NOT1 (N10195, N10181);
nand NAND3 (N10196, N10195, N3520, N7681);
nand NAND4 (N10197, N10169, N568, N1308, N1551);
xor XOR2 (N10198, N10190, N9714);
and AND3 (N10199, N10192, N7152, N3191);
not NOT1 (N10200, N10183);
xor XOR2 (N10201, N10200, N1798);
and AND4 (N10202, N10201, N5577, N5495, N10068);
nor NOR3 (N10203, N10199, N9524, N2873);
nand NAND3 (N10204, N10197, N4283, N2800);
nand NAND3 (N10205, N10193, N3219, N2978);
nor NOR4 (N10206, N10204, N9970, N7927, N902);
nand NAND3 (N10207, N10189, N10145, N7995);
or OR3 (N10208, N10198, N3220, N6140);
xor XOR2 (N10209, N10202, N1031);
nor NOR4 (N10210, N10152, N51, N5278, N2574);
nor NOR3 (N10211, N10203, N2534, N4963);
buf BUF1 (N10212, N10191);
buf BUF1 (N10213, N10207);
buf BUF1 (N10214, N10213);
nand NAND2 (N10215, N10205, N7748);
nor NOR3 (N10216, N10212, N2712, N30);
not NOT1 (N10217, N10209);
not NOT1 (N10218, N10214);
not NOT1 (N10219, N10218);
buf BUF1 (N10220, N10208);
or OR4 (N10221, N10219, N6586, N9258, N8635);
nor NOR2 (N10222, N10194, N8040);
or OR2 (N10223, N10221, N10012);
nand NAND2 (N10224, N10217, N6923);
and AND2 (N10225, N10224, N3401);
nor NOR3 (N10226, N10206, N4616, N8201);
and AND4 (N10227, N10223, N8390, N9976, N10194);
and AND2 (N10228, N10211, N8677);
and AND2 (N10229, N10227, N2272);
buf BUF1 (N10230, N10220);
nand NAND3 (N10231, N10216, N232, N5842);
not NOT1 (N10232, N10229);
and AND4 (N10233, N10226, N5215, N4231, N4036);
buf BUF1 (N10234, N10232);
or OR2 (N10235, N10228, N1490);
nand NAND4 (N10236, N10215, N2424, N1667, N4214);
or OR4 (N10237, N10210, N6572, N10031, N7659);
nand NAND4 (N10238, N10235, N9081, N9494, N3986);
not NOT1 (N10239, N10231);
buf BUF1 (N10240, N10239);
buf BUF1 (N10241, N10230);
nand NAND4 (N10242, N10225, N10221, N5611, N3929);
or OR4 (N10243, N10242, N10011, N7203, N4424);
nor NOR2 (N10244, N10196, N4676);
xor XOR2 (N10245, N10237, N2044);
nand NAND2 (N10246, N10238, N5939);
buf BUF1 (N10247, N10234);
xor XOR2 (N10248, N10241, N9528);
or OR2 (N10249, N10244, N6232);
nand NAND2 (N10250, N10249, N5671);
and AND3 (N10251, N10246, N9089, N3898);
not NOT1 (N10252, N10233);
buf BUF1 (N10253, N10247);
buf BUF1 (N10254, N10250);
and AND2 (N10255, N10254, N7635);
or OR3 (N10256, N10245, N13, N1356);
nor NOR2 (N10257, N10252, N9048);
or OR3 (N10258, N10257, N8561, N3662);
xor XOR2 (N10259, N10248, N4579);
nor NOR2 (N10260, N10243, N1993);
or OR2 (N10261, N10260, N3052);
or OR3 (N10262, N10222, N4137, N494);
and AND2 (N10263, N10236, N4157);
and AND4 (N10264, N10251, N3836, N2780, N2440);
nor NOR3 (N10265, N10262, N9944, N2913);
buf BUF1 (N10266, N10264);
nand NAND4 (N10267, N10240, N3358, N5866, N7964);
nor NOR3 (N10268, N10267, N7760, N2937);
nor NOR3 (N10269, N10255, N6668, N4661);
and AND2 (N10270, N10263, N1737);
or OR3 (N10271, N10266, N7164, N2582);
and AND3 (N10272, N10256, N9203, N2044);
xor XOR2 (N10273, N10258, N1845);
buf BUF1 (N10274, N10269);
nand NAND4 (N10275, N10261, N675, N9173, N5906);
or OR3 (N10276, N10253, N4713, N8549);
nand NAND2 (N10277, N10268, N8140);
buf BUF1 (N10278, N10272);
and AND2 (N10279, N10277, N1107);
or OR4 (N10280, N10278, N6130, N857, N6908);
or OR2 (N10281, N10270, N2641);
xor XOR2 (N10282, N10273, N4834);
and AND4 (N10283, N10275, N9812, N4207, N9579);
buf BUF1 (N10284, N10274);
xor XOR2 (N10285, N10265, N7708);
not NOT1 (N10286, N10284);
or OR2 (N10287, N10279, N10006);
not NOT1 (N10288, N10280);
not NOT1 (N10289, N10285);
nand NAND2 (N10290, N10286, N7912);
buf BUF1 (N10291, N10282);
and AND3 (N10292, N10288, N1969, N7001);
or OR3 (N10293, N10289, N7204, N439);
buf BUF1 (N10294, N10292);
buf BUF1 (N10295, N10281);
buf BUF1 (N10296, N10271);
not NOT1 (N10297, N10287);
not NOT1 (N10298, N10297);
or OR4 (N10299, N10293, N4065, N6334, N5755);
and AND2 (N10300, N10276, N2255);
or OR2 (N10301, N10300, N1357);
buf BUF1 (N10302, N10290);
and AND4 (N10303, N10295, N4690, N1458, N7689);
buf BUF1 (N10304, N10283);
buf BUF1 (N10305, N10301);
nand NAND2 (N10306, N10294, N6565);
or OR2 (N10307, N10259, N3117);
nand NAND4 (N10308, N10306, N8384, N3979, N4272);
not NOT1 (N10309, N10296);
nand NAND2 (N10310, N10305, N4060);
and AND2 (N10311, N10307, N7775);
buf BUF1 (N10312, N10310);
buf BUF1 (N10313, N10302);
and AND4 (N10314, N10298, N8508, N7664, N402);
nand NAND2 (N10315, N10311, N5367);
and AND2 (N10316, N10308, N7614);
xor XOR2 (N10317, N10304, N3135);
xor XOR2 (N10318, N10291, N4937);
nor NOR2 (N10319, N10312, N3197);
not NOT1 (N10320, N10313);
nor NOR2 (N10321, N10315, N5150);
buf BUF1 (N10322, N10319);
nand NAND3 (N10323, N10314, N769, N2051);
nor NOR2 (N10324, N10321, N7661);
and AND4 (N10325, N10303, N6312, N5861, N6785);
not NOT1 (N10326, N10316);
not NOT1 (N10327, N10320);
not NOT1 (N10328, N10325);
or OR2 (N10329, N10324, N2771);
nor NOR3 (N10330, N10317, N8621, N417);
xor XOR2 (N10331, N10327, N2714);
nand NAND2 (N10332, N10309, N5863);
and AND3 (N10333, N10332, N6461, N9295);
nor NOR2 (N10334, N10322, N3325);
nor NOR3 (N10335, N10330, N8707, N4036);
not NOT1 (N10336, N10323);
or OR4 (N10337, N10334, N2594, N3521, N8910);
not NOT1 (N10338, N10333);
or OR3 (N10339, N10328, N1320, N877);
nor NOR4 (N10340, N10338, N3252, N7340, N6038);
nand NAND2 (N10341, N10340, N3315);
not NOT1 (N10342, N10339);
not NOT1 (N10343, N10331);
nand NAND4 (N10344, N10299, N7827, N2747, N1662);
buf BUF1 (N10345, N10342);
not NOT1 (N10346, N10337);
nor NOR4 (N10347, N10326, N1369, N861, N5105);
not NOT1 (N10348, N10336);
buf BUF1 (N10349, N10343);
or OR3 (N10350, N10335, N7395, N6059);
nand NAND2 (N10351, N10318, N426);
nand NAND4 (N10352, N10348, N8615, N3482, N9662);
xor XOR2 (N10353, N10346, N2304);
and AND2 (N10354, N10353, N8667);
buf BUF1 (N10355, N10354);
not NOT1 (N10356, N10341);
xor XOR2 (N10357, N10345, N28);
xor XOR2 (N10358, N10347, N8851);
not NOT1 (N10359, N10356);
nand NAND4 (N10360, N10350, N3739, N6218, N2710);
buf BUF1 (N10361, N10359);
nand NAND3 (N10362, N10357, N6402, N9207);
xor XOR2 (N10363, N10360, N118);
nor NOR3 (N10364, N10329, N10259, N10255);
buf BUF1 (N10365, N10344);
not NOT1 (N10366, N10349);
or OR4 (N10367, N10358, N9802, N8621, N6866);
nor NOR4 (N10368, N10351, N1994, N426, N4077);
not NOT1 (N10369, N10367);
and AND4 (N10370, N10363, N3675, N4945, N462);
or OR2 (N10371, N10352, N8039);
xor XOR2 (N10372, N10369, N4010);
or OR3 (N10373, N10361, N3647, N8209);
not NOT1 (N10374, N10372);
xor XOR2 (N10375, N10366, N717);
or OR2 (N10376, N10368, N1844);
nand NAND4 (N10377, N10374, N766, N6713, N9381);
nand NAND2 (N10378, N10373, N5438);
or OR3 (N10379, N10365, N596, N1983);
not NOT1 (N10380, N10376);
nor NOR2 (N10381, N10378, N9172);
and AND4 (N10382, N10377, N5495, N7197, N2084);
or OR2 (N10383, N10364, N3615);
nand NAND4 (N10384, N10370, N1985, N2907, N9918);
not NOT1 (N10385, N10384);
or OR2 (N10386, N10362, N10327);
buf BUF1 (N10387, N10383);
and AND4 (N10388, N10355, N2748, N887, N664);
buf BUF1 (N10389, N10385);
or OR3 (N10390, N10371, N6146, N1774);
or OR2 (N10391, N10381, N7769);
xor XOR2 (N10392, N10380, N8194);
not NOT1 (N10393, N10392);
and AND4 (N10394, N10379, N6333, N9435, N5361);
buf BUF1 (N10395, N10382);
xor XOR2 (N10396, N10395, N794);
xor XOR2 (N10397, N10388, N6355);
xor XOR2 (N10398, N10389, N1235);
xor XOR2 (N10399, N10386, N5083);
nor NOR4 (N10400, N10391, N8610, N880, N9953);
nand NAND4 (N10401, N10398, N1592, N5334, N5519);
not NOT1 (N10402, N10375);
buf BUF1 (N10403, N10397);
or OR4 (N10404, N10390, N6206, N2965, N84);
buf BUF1 (N10405, N10393);
not NOT1 (N10406, N10399);
buf BUF1 (N10407, N10400);
not NOT1 (N10408, N10403);
xor XOR2 (N10409, N10404, N8252);
xor XOR2 (N10410, N10387, N3013);
xor XOR2 (N10411, N10402, N1796);
and AND2 (N10412, N10396, N8810);
buf BUF1 (N10413, N10409);
not NOT1 (N10414, N10405);
nor NOR2 (N10415, N10412, N5952);
xor XOR2 (N10416, N10414, N7612);
xor XOR2 (N10417, N10394, N4430);
and AND4 (N10418, N10415, N3059, N2267, N9313);
and AND3 (N10419, N10408, N8789, N7151);
and AND2 (N10420, N10407, N5170);
nand NAND2 (N10421, N10401, N1827);
xor XOR2 (N10422, N10410, N8579);
xor XOR2 (N10423, N10421, N4048);
nand NAND2 (N10424, N10423, N7668);
nand NAND3 (N10425, N10417, N6802, N3670);
buf BUF1 (N10426, N10419);
and AND3 (N10427, N10425, N2911, N2531);
not NOT1 (N10428, N10426);
and AND3 (N10429, N10413, N8556, N5981);
or OR2 (N10430, N10422, N2152);
nand NAND2 (N10431, N10428, N3385);
and AND3 (N10432, N10427, N7441, N2855);
or OR2 (N10433, N10420, N10114);
nand NAND4 (N10434, N10433, N10337, N1670, N3257);
nand NAND4 (N10435, N10430, N1839, N6760, N897);
and AND4 (N10436, N10432, N8881, N7797, N7360);
and AND3 (N10437, N10406, N507, N919);
and AND2 (N10438, N10434, N8444);
buf BUF1 (N10439, N10416);
and AND3 (N10440, N10429, N3182, N528);
nor NOR4 (N10441, N10440, N3605, N9865, N2611);
or OR4 (N10442, N10438, N7682, N9965, N4984);
nor NOR3 (N10443, N10418, N9784, N9316);
xor XOR2 (N10444, N10436, N5622);
or OR4 (N10445, N10441, N3250, N8966, N4773);
xor XOR2 (N10446, N10442, N5265);
or OR3 (N10447, N10445, N2533, N5917);
xor XOR2 (N10448, N10411, N4705);
not NOT1 (N10449, N10443);
buf BUF1 (N10450, N10444);
nor NOR4 (N10451, N10447, N9410, N1645, N6337);
and AND3 (N10452, N10446, N2770, N7409);
or OR3 (N10453, N10449, N7575, N7492);
and AND2 (N10454, N10431, N4417);
xor XOR2 (N10455, N10450, N9842);
nor NOR3 (N10456, N10452, N3430, N9907);
or OR4 (N10457, N10435, N4381, N7219, N7415);
nor NOR3 (N10458, N10454, N6983, N265);
nand NAND3 (N10459, N10439, N7767, N9356);
or OR4 (N10460, N10455, N87, N10095, N5737);
nand NAND4 (N10461, N10460, N2462, N5403, N793);
nand NAND4 (N10462, N10456, N6748, N3079, N4059);
and AND2 (N10463, N10459, N8338);
or OR2 (N10464, N10458, N4368);
not NOT1 (N10465, N10463);
nand NAND3 (N10466, N10437, N911, N6975);
buf BUF1 (N10467, N10462);
or OR3 (N10468, N10453, N9481, N222);
xor XOR2 (N10469, N10451, N1615);
nand NAND2 (N10470, N10465, N9809);
or OR4 (N10471, N10424, N4598, N6797, N6280);
and AND4 (N10472, N10471, N8656, N2354, N6313);
xor XOR2 (N10473, N10448, N6162);
buf BUF1 (N10474, N10461);
not NOT1 (N10475, N10467);
nand NAND4 (N10476, N10470, N6965, N2601, N3179);
not NOT1 (N10477, N10457);
not NOT1 (N10478, N10468);
nor NOR4 (N10479, N10473, N4201, N3387, N9364);
nand NAND2 (N10480, N10464, N5369);
not NOT1 (N10481, N10474);
and AND2 (N10482, N10479, N9863);
xor XOR2 (N10483, N10482, N4145);
nand NAND2 (N10484, N10478, N8473);
and AND4 (N10485, N10476, N2826, N5455, N10391);
nor NOR3 (N10486, N10485, N5034, N1477);
or OR4 (N10487, N10483, N4302, N8506, N8062);
buf BUF1 (N10488, N10486);
or OR4 (N10489, N10466, N8313, N6397, N5341);
nand NAND4 (N10490, N10469, N8085, N9508, N7714);
nor NOR2 (N10491, N10487, N4394);
and AND2 (N10492, N10488, N8445);
or OR2 (N10493, N10480, N9691);
xor XOR2 (N10494, N10484, N7874);
nand NAND3 (N10495, N10490, N3796, N1622);
nand NAND4 (N10496, N10472, N6642, N8781, N3878);
buf BUF1 (N10497, N10496);
not NOT1 (N10498, N10489);
not NOT1 (N10499, N10492);
buf BUF1 (N10500, N10481);
not NOT1 (N10501, N10500);
nand NAND4 (N10502, N10495, N1917, N7183, N5518);
nor NOR2 (N10503, N10494, N5615);
and AND4 (N10504, N10502, N1130, N9414, N34);
buf BUF1 (N10505, N10497);
nor NOR3 (N10506, N10493, N6298, N1143);
or OR3 (N10507, N10498, N9998, N3892);
nor NOR4 (N10508, N10491, N10123, N5873, N7381);
not NOT1 (N10509, N10503);
not NOT1 (N10510, N10477);
nor NOR2 (N10511, N10508, N10346);
or OR4 (N10512, N10475, N5574, N688, N10004);
not NOT1 (N10513, N10507);
xor XOR2 (N10514, N10511, N7896);
buf BUF1 (N10515, N10506);
buf BUF1 (N10516, N10504);
buf BUF1 (N10517, N10515);
buf BUF1 (N10518, N10514);
nand NAND4 (N10519, N10516, N8629, N6157, N9096);
and AND2 (N10520, N10499, N6902);
xor XOR2 (N10521, N10519, N9298);
or OR4 (N10522, N10513, N9327, N764, N4278);
and AND3 (N10523, N10509, N5211, N3005);
and AND3 (N10524, N10522, N4148, N6814);
xor XOR2 (N10525, N10501, N9188);
or OR4 (N10526, N10512, N2862, N1599, N3614);
xor XOR2 (N10527, N10524, N9193);
xor XOR2 (N10528, N10521, N6495);
or OR2 (N10529, N10505, N10361);
nor NOR3 (N10530, N10520, N5511, N2141);
not NOT1 (N10531, N10529);
not NOT1 (N10532, N10527);
or OR3 (N10533, N10523, N2041, N7982);
xor XOR2 (N10534, N10525, N4492);
buf BUF1 (N10535, N10526);
nor NOR4 (N10536, N10530, N10264, N1446, N6458);
buf BUF1 (N10537, N10536);
nor NOR3 (N10538, N10531, N6545, N3092);
and AND2 (N10539, N10535, N9021);
nand NAND4 (N10540, N10538, N1698, N673, N7807);
xor XOR2 (N10541, N10510, N6342);
buf BUF1 (N10542, N10534);
and AND3 (N10543, N10542, N10389, N5789);
nor NOR3 (N10544, N10518, N8066, N271);
nand NAND2 (N10545, N10533, N5275);
and AND4 (N10546, N10543, N3489, N6925, N5799);
or OR2 (N10547, N10541, N8689);
nand NAND2 (N10548, N10547, N5056);
buf BUF1 (N10549, N10540);
not NOT1 (N10550, N10549);
not NOT1 (N10551, N10537);
buf BUF1 (N10552, N10544);
not NOT1 (N10553, N10552);
or OR4 (N10554, N10550, N3098, N8387, N9179);
not NOT1 (N10555, N10517);
nand NAND3 (N10556, N10539, N1963, N5391);
buf BUF1 (N10557, N10556);
buf BUF1 (N10558, N10546);
nand NAND2 (N10559, N10554, N2958);
or OR4 (N10560, N10532, N3240, N7962, N5902);
xor XOR2 (N10561, N10559, N6839);
buf BUF1 (N10562, N10545);
buf BUF1 (N10563, N10555);
nor NOR4 (N10564, N10561, N3033, N9521, N10310);
buf BUF1 (N10565, N10558);
and AND2 (N10566, N10560, N2564);
nand NAND3 (N10567, N10551, N10075, N1267);
nor NOR2 (N10568, N10564, N5318);
or OR4 (N10569, N10557, N2935, N1451, N8093);
nand NAND4 (N10570, N10563, N4140, N5445, N4656);
nor NOR3 (N10571, N10569, N6948, N5493);
xor XOR2 (N10572, N10553, N5350);
nand NAND3 (N10573, N10567, N1702, N6017);
nand NAND4 (N10574, N10568, N5308, N5624, N8761);
and AND4 (N10575, N10566, N4693, N4424, N5444);
nand NAND3 (N10576, N10562, N727, N10020);
or OR3 (N10577, N10571, N7272, N7115);
nand NAND3 (N10578, N10577, N10537, N3974);
buf BUF1 (N10579, N10573);
xor XOR2 (N10580, N10528, N3010);
or OR4 (N10581, N10575, N2376, N4770, N1602);
nor NOR4 (N10582, N10579, N10278, N2659, N8862);
not NOT1 (N10583, N10574);
nand NAND2 (N10584, N10583, N9916);
and AND3 (N10585, N10572, N376, N9930);
not NOT1 (N10586, N10580);
buf BUF1 (N10587, N10565);
buf BUF1 (N10588, N10587);
nor NOR3 (N10589, N10585, N5433, N6637);
not NOT1 (N10590, N10581);
not NOT1 (N10591, N10590);
xor XOR2 (N10592, N10584, N8389);
buf BUF1 (N10593, N10582);
or OR4 (N10594, N10589, N3841, N68, N1352);
not NOT1 (N10595, N10593);
or OR3 (N10596, N10570, N5960, N6938);
nand NAND4 (N10597, N10595, N6787, N4275, N7548);
xor XOR2 (N10598, N10596, N8852);
nand NAND4 (N10599, N10588, N10507, N6082, N1953);
nand NAND4 (N10600, N10578, N7694, N1857, N4702);
or OR3 (N10601, N10576, N7939, N6137);
and AND4 (N10602, N10597, N7375, N7062, N1222);
or OR2 (N10603, N10598, N4122);
xor XOR2 (N10604, N10594, N5046);
or OR3 (N10605, N10548, N49, N5394);
nand NAND4 (N10606, N10602, N2278, N9748, N1861);
buf BUF1 (N10607, N10603);
xor XOR2 (N10608, N10600, N5095);
nor NOR4 (N10609, N10591, N6689, N413, N8125);
nand NAND2 (N10610, N10605, N9545);
not NOT1 (N10611, N10606);
xor XOR2 (N10612, N10611, N5185);
nor NOR2 (N10613, N10601, N10106);
nor NOR4 (N10614, N10610, N7966, N641, N3952);
xor XOR2 (N10615, N10592, N2665);
not NOT1 (N10616, N10604);
nor NOR4 (N10617, N10607, N7877, N3446, N7529);
xor XOR2 (N10618, N10616, N6147);
nand NAND2 (N10619, N10618, N421);
nor NOR3 (N10620, N10619, N7534, N4095);
and AND4 (N10621, N10615, N9025, N695, N7090);
xor XOR2 (N10622, N10617, N4427);
buf BUF1 (N10623, N10620);
nor NOR2 (N10624, N10599, N1866);
or OR2 (N10625, N10624, N4655);
or OR3 (N10626, N10623, N2461, N1159);
or OR3 (N10627, N10586, N8195, N565);
xor XOR2 (N10628, N10627, N10367);
buf BUF1 (N10629, N10621);
or OR3 (N10630, N10622, N128, N4364);
or OR3 (N10631, N10613, N156, N7534);
buf BUF1 (N10632, N10629);
nand NAND2 (N10633, N10614, N3648);
not NOT1 (N10634, N10609);
xor XOR2 (N10635, N10612, N3024);
not NOT1 (N10636, N10633);
nor NOR3 (N10637, N10626, N9549, N7488);
nand NAND3 (N10638, N10632, N3619, N7810);
or OR2 (N10639, N10630, N4525);
not NOT1 (N10640, N10637);
xor XOR2 (N10641, N10631, N1974);
buf BUF1 (N10642, N10634);
or OR3 (N10643, N10628, N5459, N5129);
buf BUF1 (N10644, N10608);
nor NOR3 (N10645, N10640, N2408, N8139);
or OR4 (N10646, N10643, N3091, N7560, N4995);
nand NAND3 (N10647, N10625, N9104, N10433);
xor XOR2 (N10648, N10642, N1334);
not NOT1 (N10649, N10641);
not NOT1 (N10650, N10638);
nor NOR4 (N10651, N10650, N5492, N7202, N1819);
nand NAND3 (N10652, N10651, N3304, N9733);
not NOT1 (N10653, N10646);
or OR3 (N10654, N10648, N5922, N8985);
nand NAND4 (N10655, N10654, N6909, N4561, N468);
buf BUF1 (N10656, N10649);
and AND3 (N10657, N10656, N9895, N7960);
nand NAND3 (N10658, N10644, N5677, N3177);
buf BUF1 (N10659, N10636);
not NOT1 (N10660, N10657);
or OR4 (N10661, N10645, N1461, N2778, N4567);
xor XOR2 (N10662, N10652, N1396);
nor NOR4 (N10663, N10635, N2644, N1198, N3109);
xor XOR2 (N10664, N10661, N7045);
buf BUF1 (N10665, N10658);
or OR3 (N10666, N10653, N3867, N8432);
xor XOR2 (N10667, N10665, N8292);
nand NAND2 (N10668, N10655, N1216);
nor NOR2 (N10669, N10668, N1870);
nor NOR2 (N10670, N10664, N6586);
nand NAND2 (N10671, N10647, N5636);
xor XOR2 (N10672, N10639, N3332);
xor XOR2 (N10673, N10671, N2124);
xor XOR2 (N10674, N10662, N974);
xor XOR2 (N10675, N10673, N3738);
or OR4 (N10676, N10667, N1168, N6777, N6163);
and AND3 (N10677, N10659, N2698, N6744);
not NOT1 (N10678, N10672);
or OR2 (N10679, N10670, N10604);
nor NOR4 (N10680, N10666, N9803, N8550, N10126);
and AND4 (N10681, N10677, N5023, N7775, N483);
xor XOR2 (N10682, N10679, N8598);
or OR2 (N10683, N10675, N9072);
not NOT1 (N10684, N10669);
and AND2 (N10685, N10663, N2070);
or OR4 (N10686, N10680, N3783, N4475, N6323);
or OR3 (N10687, N10686, N1791, N7231);
or OR3 (N10688, N10678, N622, N5545);
nand NAND3 (N10689, N10684, N9802, N330);
or OR2 (N10690, N10681, N2408);
or OR2 (N10691, N10685, N9953);
or OR2 (N10692, N10690, N645);
nor NOR4 (N10693, N10660, N2970, N4768, N3150);
nand NAND4 (N10694, N10683, N4341, N83, N3149);
nand NAND4 (N10695, N10688, N3638, N7084, N10560);
and AND2 (N10696, N10691, N2423);
xor XOR2 (N10697, N10695, N501);
nand NAND3 (N10698, N10674, N4857, N7790);
buf BUF1 (N10699, N10676);
nand NAND3 (N10700, N10687, N3254, N1453);
buf BUF1 (N10701, N10696);
xor XOR2 (N10702, N10693, N6171);
or OR3 (N10703, N10694, N2188, N5236);
or OR3 (N10704, N10689, N9968, N2420);
not NOT1 (N10705, N10700);
or OR2 (N10706, N10701, N8068);
and AND2 (N10707, N10692, N1865);
and AND2 (N10708, N10702, N7619);
nand NAND2 (N10709, N10699, N5072);
xor XOR2 (N10710, N10708, N10583);
xor XOR2 (N10711, N10697, N10148);
nor NOR3 (N10712, N10698, N6334, N9505);
nand NAND3 (N10713, N10703, N9023, N8546);
nor NOR4 (N10714, N10709, N645, N1670, N9581);
nand NAND4 (N10715, N10710, N6521, N2539, N6399);
and AND4 (N10716, N10715, N10047, N9330, N4142);
nand NAND4 (N10717, N10705, N1657, N4218, N6616);
nand NAND4 (N10718, N10717, N7948, N308, N5306);
buf BUF1 (N10719, N10713);
nor NOR4 (N10720, N10716, N607, N3796, N4734);
or OR3 (N10721, N10718, N3487, N3540);
and AND4 (N10722, N10682, N4352, N7775, N2105);
xor XOR2 (N10723, N10712, N1230);
xor XOR2 (N10724, N10723, N8379);
or OR4 (N10725, N10706, N6394, N6125, N6138);
xor XOR2 (N10726, N10719, N9364);
or OR2 (N10727, N10725, N6458);
nor NOR3 (N10728, N10707, N3514, N1738);
or OR3 (N10729, N10724, N6561, N308);
or OR2 (N10730, N10714, N2344);
and AND4 (N10731, N10704, N108, N10141, N9381);
not NOT1 (N10732, N10722);
xor XOR2 (N10733, N10731, N7253);
nor NOR3 (N10734, N10727, N1405, N10616);
buf BUF1 (N10735, N10734);
nor NOR3 (N10736, N10732, N8025, N8325);
xor XOR2 (N10737, N10733, N7649);
or OR4 (N10738, N10726, N10017, N1911, N9207);
buf BUF1 (N10739, N10736);
nor NOR3 (N10740, N10735, N8588, N2659);
buf BUF1 (N10741, N10729);
nand NAND2 (N10742, N10711, N4028);
nand NAND2 (N10743, N10742, N8486);
or OR4 (N10744, N10738, N861, N8469, N6795);
or OR4 (N10745, N10744, N4282, N6872, N5561);
buf BUF1 (N10746, N10745);
nand NAND3 (N10747, N10740, N5194, N6159);
nor NOR3 (N10748, N10739, N5540, N3617);
not NOT1 (N10749, N10730);
nor NOR2 (N10750, N10748, N9448);
and AND2 (N10751, N10737, N5534);
xor XOR2 (N10752, N10728, N3171);
nand NAND2 (N10753, N10746, N10162);
xor XOR2 (N10754, N10753, N1847);
buf BUF1 (N10755, N10750);
xor XOR2 (N10756, N10755, N5263);
buf BUF1 (N10757, N10743);
nand NAND3 (N10758, N10756, N8016, N5477);
not NOT1 (N10759, N10751);
nor NOR2 (N10760, N10754, N844);
or OR2 (N10761, N10720, N1235);
or OR3 (N10762, N10757, N1317, N6743);
and AND3 (N10763, N10749, N4612, N1035);
and AND3 (N10764, N10760, N3391, N2697);
xor XOR2 (N10765, N10762, N4514);
and AND2 (N10766, N10741, N6031);
and AND3 (N10767, N10747, N2953, N5054);
nor NOR2 (N10768, N10767, N5981);
or OR3 (N10769, N10766, N5218, N1207);
nor NOR2 (N10770, N10761, N9139);
not NOT1 (N10771, N10752);
or OR3 (N10772, N10769, N6766, N2521);
nor NOR2 (N10773, N10759, N9177);
buf BUF1 (N10774, N10758);
and AND3 (N10775, N10774, N6204, N5961);
nor NOR3 (N10776, N10770, N7026, N8628);
or OR4 (N10777, N10765, N8403, N1350, N3999);
not NOT1 (N10778, N10768);
and AND4 (N10779, N10764, N2941, N2209, N3876);
not NOT1 (N10780, N10776);
xor XOR2 (N10781, N10763, N8410);
and AND3 (N10782, N10771, N8306, N7748);
and AND2 (N10783, N10779, N3592);
xor XOR2 (N10784, N10721, N373);
xor XOR2 (N10785, N10780, N3097);
not NOT1 (N10786, N10777);
buf BUF1 (N10787, N10786);
nor NOR2 (N10788, N10782, N4732);
nor NOR3 (N10789, N10781, N2293, N3090);
nand NAND2 (N10790, N10783, N8520);
xor XOR2 (N10791, N10784, N9541);
nor NOR4 (N10792, N10773, N1176, N3376, N4104);
or OR4 (N10793, N10792, N7066, N436, N3967);
xor XOR2 (N10794, N10790, N8732);
buf BUF1 (N10795, N10793);
xor XOR2 (N10796, N10795, N2773);
and AND2 (N10797, N10787, N3033);
xor XOR2 (N10798, N10796, N3171);
xor XOR2 (N10799, N10798, N2409);
xor XOR2 (N10800, N10797, N10044);
buf BUF1 (N10801, N10800);
not NOT1 (N10802, N10794);
not NOT1 (N10803, N10778);
nor NOR2 (N10804, N10785, N563);
nand NAND2 (N10805, N10788, N9536);
not NOT1 (N10806, N10802);
buf BUF1 (N10807, N10772);
nor NOR4 (N10808, N10805, N505, N5309, N9981);
or OR3 (N10809, N10791, N822, N5113);
and AND3 (N10810, N10789, N8791, N6637);
nand NAND4 (N10811, N10803, N7115, N5370, N2375);
or OR2 (N10812, N10806, N10166);
or OR2 (N10813, N10811, N8186);
not NOT1 (N10814, N10807);
and AND2 (N10815, N10814, N8134);
xor XOR2 (N10816, N10801, N9338);
xor XOR2 (N10817, N10815, N8392);
nor NOR2 (N10818, N10808, N6668);
xor XOR2 (N10819, N10804, N7014);
not NOT1 (N10820, N10819);
xor XOR2 (N10821, N10809, N8803);
nor NOR4 (N10822, N10816, N1285, N8912, N10133);
xor XOR2 (N10823, N10820, N6564);
or OR4 (N10824, N10823, N9089, N6948, N10198);
or OR4 (N10825, N10824, N5668, N9639, N1042);
or OR4 (N10826, N10822, N3029, N9502, N9334);
and AND4 (N10827, N10810, N5036, N3437, N7466);
xor XOR2 (N10828, N10827, N7522);
buf BUF1 (N10829, N10812);
xor XOR2 (N10830, N10829, N9132);
not NOT1 (N10831, N10828);
buf BUF1 (N10832, N10799);
not NOT1 (N10833, N10813);
nor NOR3 (N10834, N10826, N4842, N3363);
buf BUF1 (N10835, N10831);
nand NAND3 (N10836, N10833, N7759, N539);
not NOT1 (N10837, N10834);
and AND4 (N10838, N10821, N9825, N933, N524);
xor XOR2 (N10839, N10836, N5107);
buf BUF1 (N10840, N10838);
or OR2 (N10841, N10825, N9638);
not NOT1 (N10842, N10830);
nor NOR2 (N10843, N10839, N1899);
not NOT1 (N10844, N10840);
and AND2 (N10845, N10841, N8486);
or OR3 (N10846, N10817, N7639, N2832);
buf BUF1 (N10847, N10842);
not NOT1 (N10848, N10844);
nand NAND4 (N10849, N10832, N8760, N7998, N3758);
nand NAND3 (N10850, N10847, N1529, N9107);
xor XOR2 (N10851, N10849, N6283);
and AND4 (N10852, N10851, N4912, N6016, N8558);
buf BUF1 (N10853, N10848);
buf BUF1 (N10854, N10818);
and AND2 (N10855, N10853, N4327);
or OR3 (N10856, N10843, N4598, N2447);
nor NOR4 (N10857, N10850, N7474, N2915, N8590);
nand NAND4 (N10858, N10837, N3167, N9494, N1592);
xor XOR2 (N10859, N10835, N1399);
buf BUF1 (N10860, N10845);
buf BUF1 (N10861, N10854);
xor XOR2 (N10862, N10861, N7399);
xor XOR2 (N10863, N10859, N4293);
or OR2 (N10864, N10858, N8992);
or OR4 (N10865, N10855, N5034, N6297, N9211);
buf BUF1 (N10866, N10775);
buf BUF1 (N10867, N10865);
nor NOR3 (N10868, N10864, N7877, N1760);
nand NAND3 (N10869, N10867, N7687, N8347);
buf BUF1 (N10870, N10862);
not NOT1 (N10871, N10863);
buf BUF1 (N10872, N10856);
and AND4 (N10873, N10852, N8194, N2114, N7072);
xor XOR2 (N10874, N10846, N8751);
or OR2 (N10875, N10874, N2735);
or OR2 (N10876, N10860, N4980);
and AND3 (N10877, N10869, N4565, N5743);
xor XOR2 (N10878, N10875, N2329);
and AND2 (N10879, N10876, N7330);
buf BUF1 (N10880, N10871);
buf BUF1 (N10881, N10877);
nand NAND4 (N10882, N10872, N3115, N8363, N5478);
nor NOR4 (N10883, N10873, N10089, N7306, N2977);
not NOT1 (N10884, N10870);
and AND2 (N10885, N10881, N6587);
or OR3 (N10886, N10880, N3618, N3226);
and AND4 (N10887, N10868, N7038, N310, N1629);
not NOT1 (N10888, N10883);
xor XOR2 (N10889, N10866, N8626);
nand NAND2 (N10890, N10857, N10027);
buf BUF1 (N10891, N10887);
nand NAND3 (N10892, N10878, N3854, N788);
xor XOR2 (N10893, N10882, N4658);
nand NAND3 (N10894, N10891, N4916, N633);
buf BUF1 (N10895, N10884);
nand NAND3 (N10896, N10894, N3126, N4991);
xor XOR2 (N10897, N10879, N6910);
nand NAND4 (N10898, N10893, N6673, N4867, N9226);
nand NAND3 (N10899, N10888, N3344, N2315);
nor NOR2 (N10900, N10899, N10673);
not NOT1 (N10901, N10898);
buf BUF1 (N10902, N10885);
and AND3 (N10903, N10890, N4784, N449);
or OR2 (N10904, N10900, N5374);
not NOT1 (N10905, N10886);
xor XOR2 (N10906, N10902, N205);
or OR2 (N10907, N10903, N4148);
nor NOR3 (N10908, N10889, N2113, N3270);
or OR3 (N10909, N10907, N7987, N101);
and AND2 (N10910, N10909, N8485);
and AND2 (N10911, N10892, N1814);
buf BUF1 (N10912, N10904);
not NOT1 (N10913, N10912);
or OR4 (N10914, N10895, N193, N8420, N10749);
nand NAND2 (N10915, N10914, N4682);
xor XOR2 (N10916, N10908, N519);
xor XOR2 (N10917, N10915, N3424);
xor XOR2 (N10918, N10906, N965);
nor NOR4 (N10919, N10917, N4308, N3159, N8281);
and AND3 (N10920, N10919, N10435, N9120);
and AND2 (N10921, N10918, N9811);
nand NAND4 (N10922, N10896, N6237, N5110, N6831);
not NOT1 (N10923, N10916);
nor NOR2 (N10924, N10897, N6346);
xor XOR2 (N10925, N10910, N5052);
nor NOR2 (N10926, N10924, N9360);
or OR2 (N10927, N10905, N1095);
not NOT1 (N10928, N10926);
xor XOR2 (N10929, N10901, N3478);
nor NOR2 (N10930, N10921, N8867);
buf BUF1 (N10931, N10930);
xor XOR2 (N10932, N10929, N6221);
and AND4 (N10933, N10920, N4763, N7490, N1996);
buf BUF1 (N10934, N10927);
nor NOR2 (N10935, N10934, N400);
nor NOR4 (N10936, N10928, N3204, N2579, N2223);
xor XOR2 (N10937, N10932, N10095);
and AND3 (N10938, N10922, N8509, N2809);
buf BUF1 (N10939, N10938);
and AND4 (N10940, N10931, N9421, N8264, N3190);
nand NAND4 (N10941, N10935, N1783, N558, N6973);
or OR2 (N10942, N10936, N2415);
nand NAND3 (N10943, N10925, N9978, N3630);
xor XOR2 (N10944, N10937, N5481);
nand NAND2 (N10945, N10923, N4282);
or OR3 (N10946, N10940, N10515, N2017);
and AND2 (N10947, N10945, N5047);
buf BUF1 (N10948, N10943);
xor XOR2 (N10949, N10913, N1002);
xor XOR2 (N10950, N10947, N2630);
and AND4 (N10951, N10941, N10222, N4416, N1870);
not NOT1 (N10952, N10944);
nor NOR3 (N10953, N10933, N10048, N5814);
or OR2 (N10954, N10950, N4977);
xor XOR2 (N10955, N10954, N5489);
or OR2 (N10956, N10949, N2435);
nor NOR4 (N10957, N10939, N3115, N9275, N1496);
or OR3 (N10958, N10955, N2813, N101);
or OR2 (N10959, N10948, N9927);
nor NOR4 (N10960, N10953, N9869, N1017, N1023);
buf BUF1 (N10961, N10951);
nand NAND2 (N10962, N10911, N8236);
or OR3 (N10963, N10961, N1505, N4759);
nor NOR3 (N10964, N10960, N2698, N2798);
and AND4 (N10965, N10956, N1077, N1444, N4566);
not NOT1 (N10966, N10958);
buf BUF1 (N10967, N10942);
or OR3 (N10968, N10964, N5661, N7833);
not NOT1 (N10969, N10966);
or OR4 (N10970, N10967, N2113, N5750, N2815);
xor XOR2 (N10971, N10952, N3807);
xor XOR2 (N10972, N10963, N5503);
xor XOR2 (N10973, N10959, N4015);
nand NAND4 (N10974, N10973, N4326, N6745, N10153);
nor NOR4 (N10975, N10946, N9278, N9358, N5326);
or OR2 (N10976, N10970, N6208);
and AND4 (N10977, N10972, N8162, N5905, N5369);
nand NAND3 (N10978, N10962, N3387, N2564);
not NOT1 (N10979, N10978);
nor NOR2 (N10980, N10975, N3093);
and AND3 (N10981, N10976, N10970, N4172);
or OR2 (N10982, N10957, N9828);
and AND4 (N10983, N10980, N2160, N1475, N3255);
not NOT1 (N10984, N10982);
xor XOR2 (N10985, N10979, N7223);
and AND3 (N10986, N10965, N9332, N7525);
buf BUF1 (N10987, N10974);
or OR4 (N10988, N10971, N1365, N10910, N10573);
and AND2 (N10989, N10988, N7859);
and AND2 (N10990, N10984, N2598);
buf BUF1 (N10991, N10986);
or OR3 (N10992, N10987, N7981, N9222);
nand NAND2 (N10993, N10992, N2130);
nand NAND3 (N10994, N10991, N1319, N10859);
or OR4 (N10995, N10989, N23, N1573, N5293);
or OR3 (N10996, N10977, N7534, N5191);
nand NAND3 (N10997, N10990, N7191, N9404);
nand NAND3 (N10998, N10996, N3237, N4829);
xor XOR2 (N10999, N10985, N8872);
or OR4 (N11000, N10993, N2435, N8915, N4466);
xor XOR2 (N11001, N10998, N8101);
nor NOR2 (N11002, N10969, N3705);
and AND4 (N11003, N10999, N2142, N8990, N4756);
not NOT1 (N11004, N11002);
nor NOR3 (N11005, N11003, N2533, N4503);
xor XOR2 (N11006, N10995, N3367);
and AND2 (N11007, N10997, N9291);
or OR4 (N11008, N11000, N8064, N10328, N1976);
nand NAND2 (N11009, N11008, N2124);
nor NOR3 (N11010, N11005, N1929, N5527);
not NOT1 (N11011, N10994);
or OR3 (N11012, N11001, N6121, N10910);
or OR2 (N11013, N10968, N724);
xor XOR2 (N11014, N11009, N9231);
buf BUF1 (N11015, N11012);
nor NOR3 (N11016, N11011, N6018, N926);
nor NOR4 (N11017, N11013, N3373, N1170, N7466);
or OR3 (N11018, N11007, N4098, N6145);
or OR3 (N11019, N11017, N4417, N8124);
buf BUF1 (N11020, N11018);
nor NOR2 (N11021, N10981, N9590);
buf BUF1 (N11022, N11016);
buf BUF1 (N11023, N11022);
not NOT1 (N11024, N10983);
nand NAND3 (N11025, N11006, N7334, N6716);
buf BUF1 (N11026, N11021);
nand NAND3 (N11027, N11010, N1566, N3429);
and AND4 (N11028, N11024, N644, N1944, N4737);
and AND4 (N11029, N11023, N3132, N7041, N7299);
xor XOR2 (N11030, N11028, N1224);
xor XOR2 (N11031, N11026, N8714);
buf BUF1 (N11032, N11029);
or OR4 (N11033, N11027, N8762, N1295, N8965);
nor NOR2 (N11034, N11031, N5181);
buf BUF1 (N11035, N11034);
not NOT1 (N11036, N11004);
xor XOR2 (N11037, N11019, N907);
nor NOR4 (N11038, N11020, N5490, N8780, N7952);
and AND2 (N11039, N11036, N10786);
buf BUF1 (N11040, N11035);
buf BUF1 (N11041, N11037);
nor NOR2 (N11042, N11014, N4061);
and AND4 (N11043, N11025, N8679, N762, N2929);
buf BUF1 (N11044, N11042);
or OR2 (N11045, N11043, N7974);
nor NOR3 (N11046, N11041, N634, N3318);
and AND4 (N11047, N11038, N305, N10349, N4032);
nand NAND3 (N11048, N11047, N744, N9467);
nand NAND3 (N11049, N11044, N2872, N9398);
nor NOR2 (N11050, N11032, N4121);
not NOT1 (N11051, N11049);
and AND4 (N11052, N11033, N1830, N725, N3510);
buf BUF1 (N11053, N11048);
not NOT1 (N11054, N11051);
nand NAND4 (N11055, N11039, N10365, N5104, N2339);
buf BUF1 (N11056, N11046);
xor XOR2 (N11057, N11030, N1741);
buf BUF1 (N11058, N11057);
buf BUF1 (N11059, N11050);
nand NAND4 (N11060, N11059, N5158, N7883, N6612);
or OR3 (N11061, N11055, N307, N9394);
not NOT1 (N11062, N11040);
nor NOR3 (N11063, N11061, N7454, N1948);
nor NOR4 (N11064, N11063, N516, N881, N10445);
not NOT1 (N11065, N11053);
nor NOR2 (N11066, N11045, N10576);
nor NOR4 (N11067, N11064, N2361, N9804, N2090);
xor XOR2 (N11068, N11065, N9545);
xor XOR2 (N11069, N11060, N7391);
and AND4 (N11070, N11068, N5259, N3651, N5923);
and AND2 (N11071, N11062, N10953);
buf BUF1 (N11072, N11056);
nor NOR2 (N11073, N11015, N6688);
nand NAND3 (N11074, N11072, N4721, N9866);
buf BUF1 (N11075, N11069);
nor NOR4 (N11076, N11070, N2115, N1732, N9210);
buf BUF1 (N11077, N11076);
or OR4 (N11078, N11058, N4287, N6170, N10908);
not NOT1 (N11079, N11052);
nand NAND3 (N11080, N11066, N3031, N7995);
not NOT1 (N11081, N11077);
nor NOR3 (N11082, N11079, N6661, N7221);
not NOT1 (N11083, N11075);
nand NAND4 (N11084, N11081, N3360, N7867, N9026);
or OR3 (N11085, N11073, N9393, N6444);
or OR2 (N11086, N11054, N8703);
or OR4 (N11087, N11067, N5277, N1614, N8980);
nand NAND4 (N11088, N11083, N7832, N4781, N8352);
xor XOR2 (N11089, N11080, N1638);
not NOT1 (N11090, N11089);
or OR4 (N11091, N11074, N7434, N1455, N1361);
nor NOR2 (N11092, N11086, N3516);
not NOT1 (N11093, N11091);
buf BUF1 (N11094, N11085);
buf BUF1 (N11095, N11093);
nand NAND3 (N11096, N11087, N7648, N8551);
buf BUF1 (N11097, N11092);
nor NOR3 (N11098, N11096, N3247, N1764);
not NOT1 (N11099, N11094);
buf BUF1 (N11100, N11090);
xor XOR2 (N11101, N11100, N6575);
buf BUF1 (N11102, N11101);
nand NAND4 (N11103, N11088, N541, N8324, N10762);
buf BUF1 (N11104, N11103);
not NOT1 (N11105, N11071);
buf BUF1 (N11106, N11105);
nor NOR3 (N11107, N11097, N2352, N9975);
xor XOR2 (N11108, N11107, N8421);
xor XOR2 (N11109, N11102, N8556);
buf BUF1 (N11110, N11095);
nor NOR3 (N11111, N11078, N1052, N4633);
and AND2 (N11112, N11104, N1704);
and AND3 (N11113, N11098, N8139, N2874);
nand NAND2 (N11114, N11084, N6747);
or OR3 (N11115, N11082, N385, N895);
xor XOR2 (N11116, N11110, N161);
or OR4 (N11117, N11099, N9246, N1641, N8399);
not NOT1 (N11118, N11109);
nand NAND4 (N11119, N11116, N2593, N5993, N3047);
nand NAND4 (N11120, N11111, N6096, N3841, N6806);
and AND3 (N11121, N11117, N1677, N9100);
buf BUF1 (N11122, N11119);
or OR4 (N11123, N11114, N5738, N4707, N5273);
nand NAND3 (N11124, N11115, N2193, N6609);
or OR3 (N11125, N11121, N11004, N2942);
or OR3 (N11126, N11112, N10198, N6427);
buf BUF1 (N11127, N11108);
nand NAND4 (N11128, N11118, N10642, N7565, N1810);
nand NAND4 (N11129, N11125, N4085, N3805, N9459);
xor XOR2 (N11130, N11106, N6250);
and AND4 (N11131, N11124, N9074, N9965, N1089);
or OR3 (N11132, N11130, N1055, N10585);
not NOT1 (N11133, N11129);
nand NAND3 (N11134, N11128, N5067, N8719);
nand NAND3 (N11135, N11133, N2925, N6651);
nor NOR2 (N11136, N11127, N881);
not NOT1 (N11137, N11120);
nand NAND3 (N11138, N11135, N170, N414);
xor XOR2 (N11139, N11132, N2365);
buf BUF1 (N11140, N11137);
nand NAND3 (N11141, N11139, N4944, N3888);
not NOT1 (N11142, N11122);
nand NAND4 (N11143, N11134, N5229, N3258, N1956);
and AND2 (N11144, N11113, N8657);
buf BUF1 (N11145, N11136);
not NOT1 (N11146, N11123);
or OR3 (N11147, N11142, N9840, N6796);
or OR2 (N11148, N11131, N158);
not NOT1 (N11149, N11126);
buf BUF1 (N11150, N11140);
not NOT1 (N11151, N11147);
nand NAND2 (N11152, N11143, N7192);
xor XOR2 (N11153, N11144, N2792);
nand NAND4 (N11154, N11146, N2821, N4215, N2238);
nand NAND2 (N11155, N11141, N1943);
buf BUF1 (N11156, N11149);
nand NAND4 (N11157, N11148, N2560, N11143, N4349);
nand NAND4 (N11158, N11153, N886, N10194, N8460);
nand NAND2 (N11159, N11154, N6111);
nor NOR3 (N11160, N11152, N5451, N3992);
buf BUF1 (N11161, N11150);
nand NAND3 (N11162, N11157, N6341, N7495);
buf BUF1 (N11163, N11162);
buf BUF1 (N11164, N11156);
or OR2 (N11165, N11158, N7010);
buf BUF1 (N11166, N11155);
nand NAND2 (N11167, N11160, N4860);
xor XOR2 (N11168, N11151, N85);
or OR3 (N11169, N11167, N8925, N791);
or OR4 (N11170, N11163, N288, N6117, N2379);
not NOT1 (N11171, N11166);
nor NOR2 (N11172, N11159, N10218);
xor XOR2 (N11173, N11161, N10267);
and AND4 (N11174, N11173, N7979, N798, N5164);
not NOT1 (N11175, N11164);
nand NAND3 (N11176, N11165, N1571, N4613);
buf BUF1 (N11177, N11145);
xor XOR2 (N11178, N11170, N3889);
not NOT1 (N11179, N11169);
not NOT1 (N11180, N11168);
and AND2 (N11181, N11172, N4630);
nand NAND3 (N11182, N11174, N9673, N10925);
nand NAND2 (N11183, N11179, N6260);
nand NAND2 (N11184, N11175, N9043);
not NOT1 (N11185, N11176);
not NOT1 (N11186, N11181);
and AND4 (N11187, N11178, N10208, N5383, N7601);
not NOT1 (N11188, N11138);
not NOT1 (N11189, N11185);
or OR2 (N11190, N11187, N2310);
and AND2 (N11191, N11190, N3831);
or OR4 (N11192, N11188, N11168, N6701, N8947);
or OR3 (N11193, N11177, N5500, N4236);
or OR2 (N11194, N11183, N2862);
and AND4 (N11195, N11189, N9877, N2675, N11187);
buf BUF1 (N11196, N11192);
buf BUF1 (N11197, N11182);
xor XOR2 (N11198, N11171, N2281);
nor NOR2 (N11199, N11184, N1520);
nand NAND3 (N11200, N11195, N2993, N1995);
nor NOR4 (N11201, N11199, N2858, N5295, N10666);
nor NOR2 (N11202, N11196, N8989);
buf BUF1 (N11203, N11180);
not NOT1 (N11204, N11193);
buf BUF1 (N11205, N11197);
not NOT1 (N11206, N11191);
nor NOR3 (N11207, N11202, N96, N9943);
nand NAND2 (N11208, N11205, N7977);
buf BUF1 (N11209, N11200);
and AND2 (N11210, N11186, N4156);
buf BUF1 (N11211, N11206);
nor NOR4 (N11212, N11201, N5304, N7412, N7692);
xor XOR2 (N11213, N11204, N9563);
nand NAND4 (N11214, N11210, N9195, N6098, N10124);
or OR2 (N11215, N11198, N9435);
nand NAND4 (N11216, N11215, N5113, N8789, N4054);
nor NOR4 (N11217, N11212, N8974, N3326, N2033);
nand NAND2 (N11218, N11209, N889);
not NOT1 (N11219, N11217);
xor XOR2 (N11220, N11213, N5689);
not NOT1 (N11221, N11218);
and AND2 (N11222, N11216, N8986);
buf BUF1 (N11223, N11194);
nand NAND2 (N11224, N11223, N2385);
xor XOR2 (N11225, N11214, N326);
and AND3 (N11226, N11203, N7909, N7844);
nor NOR3 (N11227, N11225, N7554, N1016);
buf BUF1 (N11228, N11211);
nand NAND4 (N11229, N11221, N10259, N7228, N6160);
buf BUF1 (N11230, N11208);
buf BUF1 (N11231, N11222);
nand NAND3 (N11232, N11220, N6566, N2908);
nand NAND2 (N11233, N11227, N394);
and AND4 (N11234, N11231, N6273, N9531, N9327);
nand NAND3 (N11235, N11233, N6611, N2254);
not NOT1 (N11236, N11230);
nor NOR4 (N11237, N11234, N6204, N487, N5788);
not NOT1 (N11238, N11219);
and AND2 (N11239, N11236, N7509);
xor XOR2 (N11240, N11237, N1766);
nor NOR2 (N11241, N11228, N6402);
and AND2 (N11242, N11240, N1856);
not NOT1 (N11243, N11226);
not NOT1 (N11244, N11241);
or OR4 (N11245, N11235, N10940, N7083, N4074);
buf BUF1 (N11246, N11207);
not NOT1 (N11247, N11242);
and AND3 (N11248, N11232, N10276, N2699);
buf BUF1 (N11249, N11238);
and AND3 (N11250, N11245, N6115, N1189);
or OR4 (N11251, N11229, N7190, N9700, N9669);
xor XOR2 (N11252, N11251, N11028);
and AND2 (N11253, N11248, N1966);
xor XOR2 (N11254, N11239, N5705);
xor XOR2 (N11255, N11224, N4853);
xor XOR2 (N11256, N11254, N3466);
xor XOR2 (N11257, N11250, N9475);
xor XOR2 (N11258, N11257, N4969);
not NOT1 (N11259, N11255);
nor NOR3 (N11260, N11252, N10307, N8291);
nand NAND4 (N11261, N11258, N10115, N3071, N76);
nand NAND4 (N11262, N11243, N394, N9629, N6261);
xor XOR2 (N11263, N11260, N8989);
buf BUF1 (N11264, N11247);
nand NAND3 (N11265, N11259, N8299, N10882);
not NOT1 (N11266, N11246);
buf BUF1 (N11267, N11265);
xor XOR2 (N11268, N11263, N8086);
and AND4 (N11269, N11261, N3555, N6010, N821);
nand NAND2 (N11270, N11264, N7928);
nor NOR4 (N11271, N11267, N2544, N101, N9508);
or OR4 (N11272, N11270, N3556, N3295, N3279);
and AND3 (N11273, N11269, N4109, N4380);
nor NOR2 (N11274, N11268, N9437);
nor NOR3 (N11275, N11249, N9123, N8373);
not NOT1 (N11276, N11253);
or OR4 (N11277, N11271, N1677, N868, N1437);
buf BUF1 (N11278, N11274);
and AND3 (N11279, N11278, N1594, N5621);
buf BUF1 (N11280, N11279);
xor XOR2 (N11281, N11277, N3703);
and AND3 (N11282, N11275, N1942, N4944);
nand NAND2 (N11283, N11272, N10157);
or OR3 (N11284, N11282, N8492, N1062);
buf BUF1 (N11285, N11256);
or OR2 (N11286, N11266, N1308);
nor NOR4 (N11287, N11280, N10250, N7899, N3763);
and AND4 (N11288, N11284, N6684, N3322, N8700);
xor XOR2 (N11289, N11281, N1194);
not NOT1 (N11290, N11273);
xor XOR2 (N11291, N11286, N10797);
not NOT1 (N11292, N11290);
buf BUF1 (N11293, N11292);
nor NOR4 (N11294, N11244, N3920, N3670, N838);
or OR4 (N11295, N11276, N5177, N8253, N5625);
buf BUF1 (N11296, N11291);
not NOT1 (N11297, N11294);
nand NAND3 (N11298, N11288, N1155, N8067);
nand NAND3 (N11299, N11289, N1372, N3990);
nor NOR3 (N11300, N11283, N1528, N7685);
buf BUF1 (N11301, N11262);
and AND2 (N11302, N11300, N8730);
nor NOR4 (N11303, N11296, N9749, N7158, N3269);
nand NAND3 (N11304, N11297, N1171, N629);
nand NAND3 (N11305, N11295, N6094, N1939);
nand NAND2 (N11306, N11305, N1738);
and AND2 (N11307, N11301, N4894);
xor XOR2 (N11308, N11304, N6537);
not NOT1 (N11309, N11293);
nand NAND4 (N11310, N11306, N7698, N2523, N2841);
nand NAND3 (N11311, N11308, N1932, N5978);
nand NAND4 (N11312, N11287, N7500, N3311, N5068);
nand NAND3 (N11313, N11309, N2937, N3025);
nand NAND2 (N11314, N11312, N394);
nor NOR2 (N11315, N11307, N1400);
not NOT1 (N11316, N11311);
and AND3 (N11317, N11315, N1304, N10588);
nand NAND4 (N11318, N11317, N4502, N8714, N7643);
not NOT1 (N11319, N11310);
not NOT1 (N11320, N11319);
xor XOR2 (N11321, N11316, N1114);
not NOT1 (N11322, N11298);
and AND2 (N11323, N11314, N8426);
nand NAND4 (N11324, N11320, N835, N1388, N8985);
nand NAND2 (N11325, N11322, N9720);
buf BUF1 (N11326, N11285);
and AND2 (N11327, N11299, N910);
nor NOR4 (N11328, N11325, N6002, N2928, N2156);
not NOT1 (N11329, N11313);
or OR4 (N11330, N11303, N6661, N4382, N3612);
buf BUF1 (N11331, N11323);
nand NAND2 (N11332, N11302, N1991);
or OR2 (N11333, N11331, N9476);
nand NAND2 (N11334, N11327, N7001);
buf BUF1 (N11335, N11328);
and AND2 (N11336, N11318, N2324);
nand NAND2 (N11337, N11333, N3753);
nor NOR3 (N11338, N11324, N3618, N10883);
buf BUF1 (N11339, N11326);
or OR3 (N11340, N11338, N1473, N9508);
not NOT1 (N11341, N11334);
not NOT1 (N11342, N11332);
or OR3 (N11343, N11335, N616, N10088);
or OR3 (N11344, N11343, N7904, N461);
not NOT1 (N11345, N11344);
nand NAND3 (N11346, N11342, N6316, N10097);
and AND2 (N11347, N11346, N3428);
xor XOR2 (N11348, N11345, N2766);
not NOT1 (N11349, N11336);
buf BUF1 (N11350, N11340);
and AND4 (N11351, N11341, N6023, N5526, N42);
nor NOR2 (N11352, N11348, N8615);
not NOT1 (N11353, N11329);
or OR2 (N11354, N11353, N8196);
nand NAND3 (N11355, N11354, N2255, N1507);
buf BUF1 (N11356, N11339);
buf BUF1 (N11357, N11321);
nand NAND3 (N11358, N11349, N3866, N7404);
xor XOR2 (N11359, N11355, N10033);
not NOT1 (N11360, N11350);
or OR2 (N11361, N11347, N6824);
xor XOR2 (N11362, N11356, N2458);
buf BUF1 (N11363, N11337);
nor NOR2 (N11364, N11362, N944);
nand NAND4 (N11365, N11363, N10641, N10279, N8076);
nand NAND2 (N11366, N11360, N6389);
not NOT1 (N11367, N11359);
not NOT1 (N11368, N11366);
nand NAND3 (N11369, N11357, N6896, N3350);
nand NAND2 (N11370, N11358, N6745);
and AND3 (N11371, N11361, N2040, N2711);
xor XOR2 (N11372, N11368, N2289);
xor XOR2 (N11373, N11365, N2028);
nand NAND2 (N11374, N11352, N6177);
or OR2 (N11375, N11351, N5917);
nand NAND2 (N11376, N11370, N4244);
not NOT1 (N11377, N11369);
not NOT1 (N11378, N11375);
and AND2 (N11379, N11372, N3751);
or OR4 (N11380, N11373, N6846, N3862, N4367);
not NOT1 (N11381, N11364);
and AND3 (N11382, N11330, N9339, N10048);
or OR2 (N11383, N11378, N3166);
and AND4 (N11384, N11374, N5146, N3966, N10938);
nand NAND4 (N11385, N11371, N6814, N10685, N4755);
nand NAND4 (N11386, N11385, N7626, N517, N2900);
nand NAND4 (N11387, N11367, N3714, N8158, N9398);
nor NOR4 (N11388, N11380, N9255, N2038, N4783);
nor NOR3 (N11389, N11384, N9633, N10384);
buf BUF1 (N11390, N11389);
nand NAND3 (N11391, N11383, N8457, N7481);
nor NOR3 (N11392, N11391, N2369, N4005);
or OR4 (N11393, N11387, N2092, N5062, N133);
or OR2 (N11394, N11390, N2827);
and AND2 (N11395, N11386, N7764);
nor NOR3 (N11396, N11379, N1814, N7963);
nor NOR4 (N11397, N11394, N3216, N4705, N1773);
or OR3 (N11398, N11392, N9289, N902);
xor XOR2 (N11399, N11396, N10763);
nor NOR4 (N11400, N11398, N10329, N6332, N8394);
or OR3 (N11401, N11388, N8415, N10472);
nor NOR2 (N11402, N11377, N9427);
and AND4 (N11403, N11401, N7786, N8373, N10605);
nand NAND3 (N11404, N11400, N9031, N7910);
and AND2 (N11405, N11382, N10507);
or OR4 (N11406, N11393, N7910, N5198, N8029);
not NOT1 (N11407, N11376);
or OR4 (N11408, N11402, N7450, N4982, N3502);
and AND4 (N11409, N11397, N7565, N3533, N3981);
nor NOR2 (N11410, N11404, N2128);
xor XOR2 (N11411, N11399, N887);
nor NOR4 (N11412, N11403, N3574, N4459, N5609);
xor XOR2 (N11413, N11410, N4789);
or OR4 (N11414, N11395, N7764, N11011, N4550);
and AND3 (N11415, N11411, N6750, N8767);
nand NAND4 (N11416, N11413, N7329, N11250, N9053);
nor NOR2 (N11417, N11381, N2774);
buf BUF1 (N11418, N11417);
buf BUF1 (N11419, N11414);
nor NOR3 (N11420, N11406, N4939, N8260);
and AND3 (N11421, N11415, N652, N6129);
nand NAND2 (N11422, N11420, N2489);
or OR3 (N11423, N11418, N2548, N1909);
nor NOR3 (N11424, N11422, N7080, N1059);
buf BUF1 (N11425, N11423);
or OR4 (N11426, N11419, N4298, N7811, N8227);
and AND3 (N11427, N11409, N8304, N2643);
or OR3 (N11428, N11425, N927, N5780);
or OR2 (N11429, N11427, N5126);
and AND3 (N11430, N11412, N7842, N8854);
xor XOR2 (N11431, N11421, N7656);
and AND4 (N11432, N11408, N6777, N6154, N2369);
nand NAND2 (N11433, N11416, N4881);
or OR4 (N11434, N11428, N9424, N7261, N3768);
not NOT1 (N11435, N11432);
buf BUF1 (N11436, N11429);
nor NOR2 (N11437, N11433, N8171);
or OR3 (N11438, N11437, N6788, N3481);
not NOT1 (N11439, N11407);
nand NAND3 (N11440, N11405, N7702, N742);
nor NOR2 (N11441, N11435, N2383);
xor XOR2 (N11442, N11439, N2646);
and AND4 (N11443, N11431, N4550, N3842, N2798);
nor NOR3 (N11444, N11430, N2116, N9983);
nor NOR2 (N11445, N11440, N16);
and AND4 (N11446, N11444, N2980, N9999, N5177);
or OR4 (N11447, N11443, N853, N734, N2500);
nor NOR3 (N11448, N11426, N3322, N8519);
xor XOR2 (N11449, N11424, N7189);
nand NAND3 (N11450, N11434, N7196, N10503);
or OR3 (N11451, N11441, N10550, N10679);
nor NOR3 (N11452, N11446, N7068, N11339);
buf BUF1 (N11453, N11447);
xor XOR2 (N11454, N11452, N8061);
nand NAND2 (N11455, N11438, N1217);
or OR3 (N11456, N11450, N4116, N5124);
buf BUF1 (N11457, N11455);
xor XOR2 (N11458, N11456, N7672);
not NOT1 (N11459, N11451);
not NOT1 (N11460, N11442);
and AND4 (N11461, N11436, N2826, N592, N9918);
buf BUF1 (N11462, N11454);
nor NOR3 (N11463, N11461, N2946, N7196);
xor XOR2 (N11464, N11463, N9938);
buf BUF1 (N11465, N11464);
and AND3 (N11466, N11457, N7725, N3507);
nand NAND3 (N11467, N11465, N9888, N2531);
or OR4 (N11468, N11445, N5647, N2905, N9502);
buf BUF1 (N11469, N11449);
nor NOR2 (N11470, N11469, N2806);
nand NAND2 (N11471, N11467, N1236);
and AND4 (N11472, N11448, N5477, N4332, N10589);
xor XOR2 (N11473, N11459, N6611);
and AND2 (N11474, N11460, N2584);
nand NAND3 (N11475, N11472, N3865, N9900);
buf BUF1 (N11476, N11473);
xor XOR2 (N11477, N11462, N2204);
xor XOR2 (N11478, N11470, N3385);
xor XOR2 (N11479, N11478, N947);
not NOT1 (N11480, N11475);
buf BUF1 (N11481, N11453);
nor NOR3 (N11482, N11466, N3024, N5244);
or OR3 (N11483, N11477, N9960, N8337);
not NOT1 (N11484, N11483);
and AND3 (N11485, N11484, N11022, N376);
not NOT1 (N11486, N11468);
buf BUF1 (N11487, N11458);
nor NOR3 (N11488, N11486, N7051, N5602);
nand NAND2 (N11489, N11480, N672);
and AND3 (N11490, N11481, N10571, N5090);
xor XOR2 (N11491, N11485, N7881);
or OR3 (N11492, N11488, N923, N3864);
nor NOR2 (N11493, N11490, N7719);
not NOT1 (N11494, N11479);
nor NOR2 (N11495, N11493, N6896);
or OR2 (N11496, N11489, N10554);
not NOT1 (N11497, N11496);
or OR2 (N11498, N11492, N6366);
not NOT1 (N11499, N11495);
buf BUF1 (N11500, N11482);
not NOT1 (N11501, N11491);
and AND4 (N11502, N11471, N8895, N668, N7151);
not NOT1 (N11503, N11498);
buf BUF1 (N11504, N11487);
nand NAND3 (N11505, N11474, N6613, N6383);
xor XOR2 (N11506, N11501, N11106);
buf BUF1 (N11507, N11506);
nand NAND3 (N11508, N11497, N3631, N190);
or OR4 (N11509, N11505, N6950, N7998, N2524);
nand NAND2 (N11510, N11499, N9712);
xor XOR2 (N11511, N11502, N5278);
not NOT1 (N11512, N11509);
not NOT1 (N11513, N11503);
nor NOR3 (N11514, N11504, N2495, N2332);
xor XOR2 (N11515, N11508, N3416);
nor NOR3 (N11516, N11494, N9973, N8434);
or OR3 (N11517, N11500, N7517, N11148);
and AND2 (N11518, N11510, N9123);
xor XOR2 (N11519, N11518, N8584);
nand NAND2 (N11520, N11515, N4224);
not NOT1 (N11521, N11516);
nand NAND2 (N11522, N11511, N6186);
and AND2 (N11523, N11521, N8678);
and AND4 (N11524, N11513, N6426, N4615, N3316);
xor XOR2 (N11525, N11524, N10670);
and AND4 (N11526, N11514, N3735, N9530, N237);
nand NAND4 (N11527, N11523, N4897, N3573, N6793);
not NOT1 (N11528, N11522);
nor NOR3 (N11529, N11476, N8383, N7417);
and AND4 (N11530, N11512, N2875, N736, N2046);
buf BUF1 (N11531, N11526);
xor XOR2 (N11532, N11519, N4787);
buf BUF1 (N11533, N11507);
nor NOR2 (N11534, N11530, N9865);
or OR4 (N11535, N11520, N6879, N7864, N3654);
or OR4 (N11536, N11531, N8246, N2093, N5463);
nor NOR3 (N11537, N11529, N10068, N1514);
buf BUF1 (N11538, N11534);
not NOT1 (N11539, N11525);
xor XOR2 (N11540, N11538, N8817);
and AND3 (N11541, N11535, N1798, N4983);
nor NOR2 (N11542, N11536, N866);
nand NAND4 (N11543, N11533, N10260, N2297, N8554);
nor NOR2 (N11544, N11540, N2153);
not NOT1 (N11545, N11528);
nor NOR2 (N11546, N11545, N2752);
not NOT1 (N11547, N11537);
not NOT1 (N11548, N11547);
nor NOR2 (N11549, N11539, N3167);
nor NOR2 (N11550, N11546, N11129);
nand NAND2 (N11551, N11527, N9046);
nor NOR3 (N11552, N11542, N2639, N1775);
nor NOR2 (N11553, N11544, N2043);
nor NOR4 (N11554, N11552, N9880, N3610, N3316);
nor NOR4 (N11555, N11532, N10025, N5409, N9938);
nor NOR4 (N11556, N11549, N9299, N10092, N1162);
and AND4 (N11557, N11548, N6360, N10791, N3210);
buf BUF1 (N11558, N11556);
or OR2 (N11559, N11550, N5908);
nor NOR2 (N11560, N11543, N9812);
nor NOR4 (N11561, N11553, N3102, N5232, N5804);
buf BUF1 (N11562, N11517);
and AND2 (N11563, N11560, N3223);
nand NAND2 (N11564, N11558, N9942);
or OR3 (N11565, N11559, N3141, N5365);
not NOT1 (N11566, N11563);
or OR3 (N11567, N11566, N3632, N4644);
nand NAND4 (N11568, N11565, N11298, N2949, N10199);
nor NOR4 (N11569, N11567, N2332, N8382, N3276);
or OR2 (N11570, N11562, N5514);
or OR2 (N11571, N11568, N737);
nand NAND3 (N11572, N11564, N11411, N8985);
xor XOR2 (N11573, N11541, N7966);
xor XOR2 (N11574, N11561, N840);
nor NOR4 (N11575, N11557, N7077, N6193, N1676);
xor XOR2 (N11576, N11570, N453);
nand NAND4 (N11577, N11571, N2529, N9315, N946);
nand NAND2 (N11578, N11574, N1879);
xor XOR2 (N11579, N11577, N1497);
xor XOR2 (N11580, N11576, N1069);
or OR2 (N11581, N11572, N4363);
nand NAND4 (N11582, N11554, N5426, N8825, N3463);
nor NOR3 (N11583, N11573, N8699, N1940);
not NOT1 (N11584, N11582);
or OR4 (N11585, N11584, N276, N10192, N1595);
xor XOR2 (N11586, N11555, N3360);
nor NOR3 (N11587, N11569, N11362, N6414);
buf BUF1 (N11588, N11581);
nand NAND3 (N11589, N11579, N7355, N2683);
buf BUF1 (N11590, N11578);
nor NOR2 (N11591, N11575, N969);
and AND2 (N11592, N11586, N6730);
or OR2 (N11593, N11591, N9482);
xor XOR2 (N11594, N11593, N586);
or OR4 (N11595, N11587, N7914, N837, N4320);
xor XOR2 (N11596, N11585, N8160);
or OR2 (N11597, N11589, N9858);
and AND3 (N11598, N11595, N2180, N8530);
nor NOR4 (N11599, N11596, N6413, N1765, N9505);
or OR2 (N11600, N11598, N9138);
xor XOR2 (N11601, N11594, N5022);
xor XOR2 (N11602, N11592, N9901);
not NOT1 (N11603, N11600);
nor NOR4 (N11604, N11580, N8351, N6258, N2832);
buf BUF1 (N11605, N11603);
and AND3 (N11606, N11602, N7296, N2363);
nand NAND2 (N11607, N11605, N5910);
nor NOR2 (N11608, N11599, N5083);
nand NAND2 (N11609, N11606, N3774);
xor XOR2 (N11610, N11609, N6507);
buf BUF1 (N11611, N11597);
nand NAND4 (N11612, N11608, N1873, N5923, N2095);
buf BUF1 (N11613, N11588);
xor XOR2 (N11614, N11610, N7167);
or OR4 (N11615, N11551, N9023, N5475, N2362);
and AND3 (N11616, N11601, N5627, N8696);
and AND2 (N11617, N11615, N416);
nor NOR3 (N11618, N11617, N2582, N5368);
and AND4 (N11619, N11618, N9477, N334, N1106);
nor NOR4 (N11620, N11613, N9192, N3144, N2336);
not NOT1 (N11621, N11604);
or OR4 (N11622, N11612, N9076, N695, N4853);
nand NAND2 (N11623, N11590, N2245);
nand NAND3 (N11624, N11623, N850, N297);
and AND3 (N11625, N11619, N6483, N399);
and AND2 (N11626, N11583, N4444);
or OR2 (N11627, N11622, N10807);
buf BUF1 (N11628, N11626);
xor XOR2 (N11629, N11628, N10121);
or OR4 (N11630, N11616, N4675, N10930, N7738);
or OR4 (N11631, N11630, N7848, N5459, N1327);
buf BUF1 (N11632, N11614);
not NOT1 (N11633, N11611);
buf BUF1 (N11634, N11620);
xor XOR2 (N11635, N11607, N5815);
buf BUF1 (N11636, N11621);
nor NOR4 (N11637, N11625, N7885, N259, N1136);
buf BUF1 (N11638, N11629);
and AND3 (N11639, N11634, N254, N8066);
xor XOR2 (N11640, N11636, N4719);
nand NAND2 (N11641, N11639, N1048);
nor NOR4 (N11642, N11641, N8324, N11113, N9512);
nor NOR3 (N11643, N11632, N2544, N2434);
and AND2 (N11644, N11638, N3969);
buf BUF1 (N11645, N11637);
not NOT1 (N11646, N11642);
buf BUF1 (N11647, N11627);
nand NAND4 (N11648, N11633, N6, N5703, N3383);
nand NAND4 (N11649, N11631, N11611, N2335, N5697);
nor NOR3 (N11650, N11643, N6492, N5236);
nand NAND4 (N11651, N11645, N6039, N6791, N8430);
buf BUF1 (N11652, N11649);
and AND2 (N11653, N11651, N3746);
buf BUF1 (N11654, N11647);
and AND4 (N11655, N11646, N8093, N8238, N5759);
not NOT1 (N11656, N11644);
and AND3 (N11657, N11656, N10745, N7967);
nand NAND4 (N11658, N11650, N6701, N5422, N1713);
xor XOR2 (N11659, N11652, N7934);
nand NAND4 (N11660, N11654, N858, N1713, N925);
xor XOR2 (N11661, N11658, N10936);
buf BUF1 (N11662, N11657);
and AND4 (N11663, N11635, N3248, N1693, N11102);
nor NOR3 (N11664, N11663, N2943, N6247);
and AND2 (N11665, N11640, N8013);
not NOT1 (N11666, N11648);
or OR2 (N11667, N11664, N2761);
xor XOR2 (N11668, N11624, N37);
and AND4 (N11669, N11662, N8022, N11051, N6170);
nor NOR2 (N11670, N11665, N6156);
buf BUF1 (N11671, N11661);
nor NOR4 (N11672, N11669, N8026, N8600, N2673);
xor XOR2 (N11673, N11672, N10090);
and AND4 (N11674, N11673, N8184, N4454, N6176);
xor XOR2 (N11675, N11667, N1316);
or OR2 (N11676, N11653, N3346);
nand NAND2 (N11677, N11674, N9352);
nor NOR2 (N11678, N11676, N933);
and AND2 (N11679, N11678, N8786);
nand NAND2 (N11680, N11677, N10253);
buf BUF1 (N11681, N11666);
not NOT1 (N11682, N11659);
nand NAND4 (N11683, N11670, N10695, N8229, N367);
xor XOR2 (N11684, N11668, N4697);
or OR3 (N11685, N11660, N9738, N8550);
nand NAND4 (N11686, N11683, N8739, N7868, N9057);
xor XOR2 (N11687, N11679, N6890);
buf BUF1 (N11688, N11687);
buf BUF1 (N11689, N11681);
xor XOR2 (N11690, N11675, N9215);
nand NAND4 (N11691, N11671, N6526, N508, N7870);
nand NAND3 (N11692, N11682, N7882, N6048);
and AND2 (N11693, N11688, N10958);
or OR3 (N11694, N11680, N3203, N10798);
and AND4 (N11695, N11686, N5393, N8765, N11199);
or OR4 (N11696, N11690, N6983, N6616, N3695);
or OR4 (N11697, N11684, N8887, N5072, N10982);
buf BUF1 (N11698, N11697);
nand NAND4 (N11699, N11692, N7909, N8560, N5780);
xor XOR2 (N11700, N11695, N2490);
buf BUF1 (N11701, N11655);
or OR2 (N11702, N11693, N5600);
xor XOR2 (N11703, N11699, N11201);
xor XOR2 (N11704, N11698, N10077);
buf BUF1 (N11705, N11702);
not NOT1 (N11706, N11694);
nor NOR3 (N11707, N11691, N10345, N3027);
not NOT1 (N11708, N11704);
or OR2 (N11709, N11703, N5855);
not NOT1 (N11710, N11706);
xor XOR2 (N11711, N11709, N10132);
not NOT1 (N11712, N11708);
and AND2 (N11713, N11685, N2624);
nand NAND3 (N11714, N11705, N3268, N1648);
buf BUF1 (N11715, N11707);
nand NAND4 (N11716, N11714, N9729, N4068, N1075);
and AND4 (N11717, N11701, N9364, N2801, N1441);
nor NOR4 (N11718, N11689, N2613, N7873, N187);
nand NAND3 (N11719, N11716, N9624, N4707);
nand NAND3 (N11720, N11719, N10638, N11175);
and AND3 (N11721, N11717, N9232, N966);
or OR2 (N11722, N11715, N3546);
nand NAND4 (N11723, N11720, N6711, N4907, N1364);
or OR4 (N11724, N11712, N9498, N10887, N1093);
nor NOR4 (N11725, N11711, N10749, N9788, N8082);
and AND4 (N11726, N11700, N7632, N7252, N9301);
nand NAND4 (N11727, N11724, N5469, N6494, N10522);
nor NOR4 (N11728, N11710, N5047, N4888, N6334);
not NOT1 (N11729, N11722);
not NOT1 (N11730, N11713);
buf BUF1 (N11731, N11696);
xor XOR2 (N11732, N11729, N9859);
nand NAND3 (N11733, N11732, N8734, N2310);
buf BUF1 (N11734, N11721);
and AND4 (N11735, N11718, N2849, N3925, N4207);
nand NAND2 (N11736, N11731, N3597);
or OR2 (N11737, N11726, N8406);
not NOT1 (N11738, N11727);
or OR4 (N11739, N11733, N870, N6695, N2355);
nor NOR4 (N11740, N11730, N7454, N2903, N158);
buf BUF1 (N11741, N11735);
nor NOR4 (N11742, N11740, N5896, N5198, N3959);
xor XOR2 (N11743, N11738, N491);
nand NAND2 (N11744, N11723, N1743);
nor NOR4 (N11745, N11737, N4712, N8965, N8953);
xor XOR2 (N11746, N11734, N9057);
buf BUF1 (N11747, N11743);
xor XOR2 (N11748, N11741, N11299);
and AND4 (N11749, N11745, N7634, N3684, N2641);
nor NOR4 (N11750, N11746, N10525, N2508, N8179);
or OR3 (N11751, N11749, N3408, N4429);
and AND2 (N11752, N11728, N7159);
or OR3 (N11753, N11747, N3348, N10713);
buf BUF1 (N11754, N11742);
not NOT1 (N11755, N11753);
and AND3 (N11756, N11748, N7098, N9683);
xor XOR2 (N11757, N11736, N1375);
nand NAND2 (N11758, N11755, N10819);
or OR3 (N11759, N11744, N2303, N7205);
buf BUF1 (N11760, N11739);
and AND4 (N11761, N11754, N6428, N2824, N1400);
not NOT1 (N11762, N11758);
buf BUF1 (N11763, N11725);
buf BUF1 (N11764, N11760);
not NOT1 (N11765, N11764);
xor XOR2 (N11766, N11756, N8551);
nor NOR2 (N11767, N11766, N9461);
xor XOR2 (N11768, N11757, N3017);
and AND2 (N11769, N11759, N6850);
buf BUF1 (N11770, N11762);
nor NOR4 (N11771, N11750, N8766, N9295, N1389);
and AND3 (N11772, N11752, N10720, N3564);
not NOT1 (N11773, N11763);
and AND3 (N11774, N11751, N246, N5015);
nand NAND4 (N11775, N11773, N711, N9185, N4181);
buf BUF1 (N11776, N11765);
buf BUF1 (N11777, N11774);
nor NOR3 (N11778, N11776, N5955, N193);
and AND2 (N11779, N11775, N8272);
nand NAND4 (N11780, N11778, N10149, N8364, N2005);
xor XOR2 (N11781, N11769, N3569);
xor XOR2 (N11782, N11781, N4005);
and AND3 (N11783, N11761, N4769, N6783);
not NOT1 (N11784, N11782);
and AND2 (N11785, N11783, N11440);
or OR3 (N11786, N11784, N4695, N8234);
nand NAND2 (N11787, N11780, N9143);
nand NAND4 (N11788, N11768, N3790, N11523, N9891);
xor XOR2 (N11789, N11779, N10191);
nand NAND3 (N11790, N11786, N5221, N8699);
buf BUF1 (N11791, N11771);
buf BUF1 (N11792, N11790);
xor XOR2 (N11793, N11770, N6371);
nand NAND3 (N11794, N11777, N3044, N420);
nor NOR3 (N11795, N11787, N2375, N9998);
or OR2 (N11796, N11785, N7051);
nand NAND2 (N11797, N11793, N9643);
or OR4 (N11798, N11795, N6793, N7536, N4528);
not NOT1 (N11799, N11789);
buf BUF1 (N11800, N11788);
buf BUF1 (N11801, N11767);
nor NOR2 (N11802, N11798, N4865);
xor XOR2 (N11803, N11772, N3941);
not NOT1 (N11804, N11801);
nand NAND4 (N11805, N11796, N4416, N1435, N4811);
nand NAND2 (N11806, N11794, N717);
nand NAND4 (N11807, N11792, N5168, N6747, N5700);
and AND2 (N11808, N11804, N10557);
buf BUF1 (N11809, N11791);
nor NOR2 (N11810, N11802, N5734);
and AND2 (N11811, N11809, N2236);
and AND2 (N11812, N11807, N6175);
nand NAND3 (N11813, N11800, N6221, N1878);
buf BUF1 (N11814, N11812);
and AND2 (N11815, N11803, N6939);
or OR2 (N11816, N11811, N4411);
nor NOR2 (N11817, N11813, N9303);
buf BUF1 (N11818, N11810);
buf BUF1 (N11819, N11815);
nand NAND3 (N11820, N11806, N5707, N11766);
and AND2 (N11821, N11818, N6907);
buf BUF1 (N11822, N11805);
or OR2 (N11823, N11799, N10263);
xor XOR2 (N11824, N11822, N7053);
buf BUF1 (N11825, N11824);
or OR2 (N11826, N11816, N67);
not NOT1 (N11827, N11808);
not NOT1 (N11828, N11825);
or OR3 (N11829, N11797, N6518, N10787);
or OR3 (N11830, N11823, N1538, N4384);
xor XOR2 (N11831, N11828, N9890);
nor NOR2 (N11832, N11814, N10624);
buf BUF1 (N11833, N11832);
buf BUF1 (N11834, N11833);
nor NOR4 (N11835, N11817, N11315, N6735, N7382);
buf BUF1 (N11836, N11830);
or OR4 (N11837, N11827, N9332, N10780, N2926);
nor NOR3 (N11838, N11819, N5418, N1977);
xor XOR2 (N11839, N11836, N713);
or OR3 (N11840, N11829, N11363, N10687);
or OR4 (N11841, N11820, N914, N10313, N10651);
and AND4 (N11842, N11840, N53, N5294, N10131);
or OR4 (N11843, N11837, N884, N9226, N9299);
not NOT1 (N11844, N11843);
not NOT1 (N11845, N11842);
nand NAND4 (N11846, N11841, N3070, N9077, N672);
not NOT1 (N11847, N11831);
not NOT1 (N11848, N11845);
nand NAND3 (N11849, N11835, N998, N9618);
buf BUF1 (N11850, N11846);
nor NOR2 (N11851, N11848, N3884);
xor XOR2 (N11852, N11844, N5202);
nor NOR3 (N11853, N11849, N4893, N3059);
xor XOR2 (N11854, N11838, N1445);
and AND4 (N11855, N11847, N11165, N3155, N3285);
xor XOR2 (N11856, N11839, N8931);
nand NAND3 (N11857, N11855, N1896, N7284);
nor NOR4 (N11858, N11821, N8768, N8082, N11268);
or OR3 (N11859, N11854, N10490, N2316);
xor XOR2 (N11860, N11859, N5513);
xor XOR2 (N11861, N11853, N7405);
buf BUF1 (N11862, N11851);
xor XOR2 (N11863, N11850, N3981);
and AND2 (N11864, N11856, N6143);
or OR4 (N11865, N11826, N7023, N6863, N6785);
nand NAND2 (N11866, N11865, N9297);
nand NAND3 (N11867, N11862, N7900, N2121);
xor XOR2 (N11868, N11866, N2552);
or OR2 (N11869, N11834, N11831);
and AND4 (N11870, N11858, N9979, N6477, N6884);
nor NOR3 (N11871, N11869, N5728, N5671);
buf BUF1 (N11872, N11870);
xor XOR2 (N11873, N11857, N1897);
nand NAND2 (N11874, N11868, N2261);
and AND4 (N11875, N11872, N4174, N11370, N3674);
xor XOR2 (N11876, N11871, N8461);
xor XOR2 (N11877, N11874, N5173);
nand NAND4 (N11878, N11860, N2302, N6873, N191);
xor XOR2 (N11879, N11863, N8675);
and AND4 (N11880, N11864, N746, N10481, N10537);
buf BUF1 (N11881, N11879);
and AND2 (N11882, N11852, N6929);
and AND4 (N11883, N11873, N3745, N227, N601);
xor XOR2 (N11884, N11881, N10620);
not NOT1 (N11885, N11861);
buf BUF1 (N11886, N11884);
and AND4 (N11887, N11878, N4630, N7536, N9588);
buf BUF1 (N11888, N11886);
or OR4 (N11889, N11880, N507, N8803, N8433);
or OR3 (N11890, N11888, N9098, N4597);
nand NAND3 (N11891, N11889, N2079, N9318);
not NOT1 (N11892, N11891);
xor XOR2 (N11893, N11877, N11501);
buf BUF1 (N11894, N11882);
buf BUF1 (N11895, N11875);
not NOT1 (N11896, N11894);
nand NAND4 (N11897, N11890, N1941, N1850, N6076);
not NOT1 (N11898, N11892);
nor NOR3 (N11899, N11897, N138, N4195);
buf BUF1 (N11900, N11899);
buf BUF1 (N11901, N11900);
buf BUF1 (N11902, N11896);
nand NAND4 (N11903, N11883, N10336, N5334, N9511);
and AND2 (N11904, N11895, N7849);
xor XOR2 (N11905, N11876, N414);
buf BUF1 (N11906, N11902);
and AND2 (N11907, N11904, N3702);
and AND3 (N11908, N11901, N10590, N670);
nor NOR2 (N11909, N11885, N7808);
or OR4 (N11910, N11898, N2033, N8363, N6872);
nor NOR3 (N11911, N11909, N2597, N4970);
buf BUF1 (N11912, N11867);
xor XOR2 (N11913, N11911, N9399);
buf BUF1 (N11914, N11912);
nand NAND3 (N11915, N11914, N1093, N9120);
xor XOR2 (N11916, N11905, N4823);
nor NOR3 (N11917, N11906, N6083, N2124);
or OR4 (N11918, N11913, N8849, N7670, N2212);
xor XOR2 (N11919, N11916, N11060);
nand NAND3 (N11920, N11910, N11252, N2573);
xor XOR2 (N11921, N11915, N2603);
nor NOR4 (N11922, N11917, N5936, N7938, N3899);
nand NAND3 (N11923, N11919, N7731, N1174);
nor NOR2 (N11924, N11923, N2102);
nand NAND4 (N11925, N11921, N3323, N3976, N8791);
not NOT1 (N11926, N11918);
nand NAND2 (N11927, N11925, N4469);
buf BUF1 (N11928, N11907);
xor XOR2 (N11929, N11926, N8757);
not NOT1 (N11930, N11929);
not NOT1 (N11931, N11908);
buf BUF1 (N11932, N11922);
nand NAND4 (N11933, N11893, N2342, N7755, N327);
nor NOR4 (N11934, N11930, N104, N2160, N1772);
and AND3 (N11935, N11934, N9416, N4374);
or OR3 (N11936, N11927, N10177, N5063);
nor NOR3 (N11937, N11935, N3914, N3063);
and AND3 (N11938, N11903, N4092, N62);
or OR3 (N11939, N11937, N3927, N10328);
or OR2 (N11940, N11920, N3734);
xor XOR2 (N11941, N11938, N9661);
nor NOR3 (N11942, N11931, N10358, N10628);
not NOT1 (N11943, N11924);
nor NOR2 (N11944, N11943, N8418);
buf BUF1 (N11945, N11928);
nor NOR2 (N11946, N11944, N1938);
not NOT1 (N11947, N11941);
or OR4 (N11948, N11936, N6426, N6366, N2978);
xor XOR2 (N11949, N11940, N6091);
or OR3 (N11950, N11932, N4932, N6112);
not NOT1 (N11951, N11949);
xor XOR2 (N11952, N11939, N3338);
xor XOR2 (N11953, N11946, N9950);
nor NOR3 (N11954, N11952, N10122, N1118);
not NOT1 (N11955, N11951);
nor NOR2 (N11956, N11948, N6138);
or OR4 (N11957, N11887, N9019, N7605, N9616);
not NOT1 (N11958, N11942);
buf BUF1 (N11959, N11945);
nand NAND3 (N11960, N11947, N4191, N1027);
nand NAND4 (N11961, N11954, N10804, N8293, N5273);
or OR3 (N11962, N11957, N2249, N1548);
nand NAND2 (N11963, N11950, N10992);
buf BUF1 (N11964, N11955);
or OR4 (N11965, N11960, N2848, N5398, N6699);
and AND2 (N11966, N11933, N3614);
nand NAND4 (N11967, N11965, N11359, N1175, N5935);
nor NOR4 (N11968, N11964, N8006, N11586, N479);
or OR4 (N11969, N11958, N2661, N11264, N8887);
xor XOR2 (N11970, N11966, N5044);
nand NAND2 (N11971, N11969, N8037);
not NOT1 (N11972, N11968);
or OR3 (N11973, N11961, N8369, N2650);
or OR2 (N11974, N11972, N4198);
and AND3 (N11975, N11953, N8265, N11056);
or OR2 (N11976, N11975, N5953);
or OR2 (N11977, N11967, N8672);
xor XOR2 (N11978, N11977, N6986);
nor NOR4 (N11979, N11973, N1423, N11332, N1741);
nor NOR3 (N11980, N11962, N2571, N10977);
buf BUF1 (N11981, N11974);
or OR2 (N11982, N11971, N11355);
buf BUF1 (N11983, N11956);
nor NOR2 (N11984, N11978, N6752);
not NOT1 (N11985, N11981);
or OR4 (N11986, N11980, N1744, N5325, N1760);
xor XOR2 (N11987, N11985, N8593);
and AND4 (N11988, N11983, N10202, N5175, N7932);
nand NAND3 (N11989, N11987, N189, N2336);
or OR4 (N11990, N11988, N7174, N6905, N9894);
nand NAND4 (N11991, N11963, N2685, N4709, N11532);
nor NOR4 (N11992, N11991, N11391, N1989, N6108);
or OR2 (N11993, N11990, N561);
not NOT1 (N11994, N11984);
or OR4 (N11995, N11992, N965, N10352, N3486);
and AND2 (N11996, N11993, N6558);
not NOT1 (N11997, N11986);
buf BUF1 (N11998, N11995);
xor XOR2 (N11999, N11996, N8885);
nor NOR3 (N12000, N11989, N11550, N9844);
buf BUF1 (N12001, N11998);
nand NAND4 (N12002, N11970, N9388, N3948, N1047);
xor XOR2 (N12003, N11959, N1449);
and AND2 (N12004, N11999, N8751);
nand NAND3 (N12005, N11994, N10522, N11960);
xor XOR2 (N12006, N11979, N9026);
and AND2 (N12007, N12002, N8078);
not NOT1 (N12008, N12004);
not NOT1 (N12009, N11982);
and AND3 (N12010, N12005, N4430, N11300);
and AND4 (N12011, N12001, N10509, N9000, N10676);
buf BUF1 (N12012, N12006);
nor NOR2 (N12013, N12010, N1545);
nor NOR3 (N12014, N11997, N11929, N8940);
nand NAND4 (N12015, N11976, N5743, N10126, N5198);
or OR2 (N12016, N12014, N10249);
not NOT1 (N12017, N12000);
nand NAND4 (N12018, N12013, N9234, N3569, N2464);
nand NAND4 (N12019, N12009, N2845, N6139, N5049);
not NOT1 (N12020, N12007);
or OR2 (N12021, N12017, N3435);
and AND3 (N12022, N12016, N8893, N3148);
buf BUF1 (N12023, N12011);
nand NAND4 (N12024, N12022, N7938, N6132, N4495);
or OR3 (N12025, N12019, N631, N1017);
or OR2 (N12026, N12018, N5315);
nor NOR2 (N12027, N12003, N5347);
or OR4 (N12028, N12012, N3640, N10440, N1964);
xor XOR2 (N12029, N12028, N6160);
or OR2 (N12030, N12020, N10879);
xor XOR2 (N12031, N12029, N8227);
or OR4 (N12032, N12031, N10917, N9007, N2765);
and AND2 (N12033, N12025, N8925);
not NOT1 (N12034, N12032);
and AND4 (N12035, N12034, N7365, N3382, N8363);
not NOT1 (N12036, N12008);
buf BUF1 (N12037, N12021);
xor XOR2 (N12038, N12035, N8703);
not NOT1 (N12039, N12023);
buf BUF1 (N12040, N12030);
nand NAND2 (N12041, N12033, N7762);
or OR3 (N12042, N12041, N5236, N7880);
buf BUF1 (N12043, N12026);
xor XOR2 (N12044, N12042, N3284);
xor XOR2 (N12045, N12039, N11673);
nor NOR4 (N12046, N12043, N11426, N3820, N2679);
buf BUF1 (N12047, N12027);
or OR4 (N12048, N12040, N7618, N184, N6153);
not NOT1 (N12049, N12038);
xor XOR2 (N12050, N12037, N10399);
nor NOR4 (N12051, N12047, N8455, N3163, N8519);
or OR3 (N12052, N12051, N1421, N10759);
and AND3 (N12053, N12036, N9660, N1963);
buf BUF1 (N12054, N12024);
xor XOR2 (N12055, N12052, N8658);
nand NAND4 (N12056, N12055, N2112, N10176, N8465);
or OR3 (N12057, N12045, N5915, N10174);
nand NAND2 (N12058, N12048, N5580);
or OR4 (N12059, N12056, N974, N3610, N9581);
or OR4 (N12060, N12054, N5268, N6677, N701);
nand NAND3 (N12061, N12053, N8335, N3061);
xor XOR2 (N12062, N12049, N632);
or OR3 (N12063, N12046, N7371, N10395);
nand NAND3 (N12064, N12050, N9965, N4775);
or OR4 (N12065, N12063, N2836, N8719, N3250);
buf BUF1 (N12066, N12058);
nand NAND4 (N12067, N12044, N9858, N10011, N3753);
and AND4 (N12068, N12066, N3458, N7004, N4090);
not NOT1 (N12069, N12062);
not NOT1 (N12070, N12061);
nor NOR2 (N12071, N12067, N3273);
nor NOR3 (N12072, N12059, N9372, N2820);
not NOT1 (N12073, N12068);
nor NOR4 (N12074, N12057, N11852, N10857, N8985);
nand NAND4 (N12075, N12074, N5394, N7763, N6277);
nand NAND2 (N12076, N12060, N11955);
and AND4 (N12077, N12076, N1268, N3196, N2627);
nor NOR2 (N12078, N12069, N10977);
not NOT1 (N12079, N12073);
or OR4 (N12080, N12070, N9298, N2926, N6412);
nand NAND2 (N12081, N12078, N5432);
xor XOR2 (N12082, N12064, N9727);
nor NOR4 (N12083, N12077, N5491, N11430, N5553);
or OR2 (N12084, N12015, N7295);
not NOT1 (N12085, N12065);
and AND2 (N12086, N12071, N7561);
nand NAND4 (N12087, N12085, N6627, N11898, N10891);
buf BUF1 (N12088, N12082);
not NOT1 (N12089, N12087);
not NOT1 (N12090, N12080);
and AND4 (N12091, N12090, N9907, N10611, N10086);
nor NOR2 (N12092, N12091, N6061);
nor NOR3 (N12093, N12084, N4206, N8736);
not NOT1 (N12094, N12088);
nand NAND4 (N12095, N12083, N7946, N11091, N126);
buf BUF1 (N12096, N12081);
nor NOR2 (N12097, N12089, N1659);
xor XOR2 (N12098, N12097, N4820);
xor XOR2 (N12099, N12086, N4203);
buf BUF1 (N12100, N12079);
nand NAND3 (N12101, N12100, N4914, N5616);
buf BUF1 (N12102, N12098);
and AND3 (N12103, N12075, N11773, N10184);
buf BUF1 (N12104, N12099);
or OR3 (N12105, N12095, N9732, N3216);
nor NOR2 (N12106, N12105, N3364);
buf BUF1 (N12107, N12093);
and AND3 (N12108, N12103, N5709, N796);
nor NOR3 (N12109, N12094, N466, N4264);
buf BUF1 (N12110, N12072);
xor XOR2 (N12111, N12101, N11106);
buf BUF1 (N12112, N12104);
and AND4 (N12113, N12110, N11815, N11353, N6583);
nand NAND3 (N12114, N12111, N4192, N5220);
buf BUF1 (N12115, N12108);
and AND2 (N12116, N12107, N4694);
not NOT1 (N12117, N12109);
xor XOR2 (N12118, N12102, N698);
not NOT1 (N12119, N12114);
and AND4 (N12120, N12115, N2906, N1769, N4646);
nor NOR4 (N12121, N12119, N5964, N1989, N7456);
and AND3 (N12122, N12117, N8345, N1799);
nor NOR3 (N12123, N12096, N11798, N884);
buf BUF1 (N12124, N12120);
xor XOR2 (N12125, N12121, N2935);
xor XOR2 (N12126, N12092, N9620);
and AND3 (N12127, N12116, N454, N1647);
or OR3 (N12128, N12125, N2659, N437);
nand NAND2 (N12129, N12123, N5237);
and AND4 (N12130, N12128, N9179, N1836, N6438);
buf BUF1 (N12131, N12129);
buf BUF1 (N12132, N12130);
or OR2 (N12133, N12124, N5587);
buf BUF1 (N12134, N12112);
nand NAND2 (N12135, N12118, N3809);
nand NAND4 (N12136, N12106, N3649, N8541, N1158);
nor NOR3 (N12137, N12113, N953, N4941);
not NOT1 (N12138, N12135);
nor NOR3 (N12139, N12131, N7618, N4669);
nor NOR3 (N12140, N12133, N4780, N3672);
nand NAND3 (N12141, N12137, N1143, N11559);
xor XOR2 (N12142, N12141, N18);
or OR4 (N12143, N12127, N11210, N8388, N9765);
nor NOR4 (N12144, N12140, N10809, N9229, N1062);
nand NAND2 (N12145, N12132, N5000);
and AND2 (N12146, N12122, N12140);
nor NOR3 (N12147, N12145, N6295, N3200);
nand NAND3 (N12148, N12144, N8525, N7983);
buf BUF1 (N12149, N12148);
not NOT1 (N12150, N12143);
or OR4 (N12151, N12150, N8204, N10981, N5687);
nor NOR4 (N12152, N12142, N1851, N3426, N7307);
or OR2 (N12153, N12147, N11408);
nand NAND4 (N12154, N12134, N9585, N8888, N5425);
nor NOR2 (N12155, N12126, N10324);
or OR2 (N12156, N12136, N8878);
buf BUF1 (N12157, N12149);
xor XOR2 (N12158, N12157, N8461);
or OR2 (N12159, N12153, N12053);
not NOT1 (N12160, N12155);
xor XOR2 (N12161, N12152, N9268);
not NOT1 (N12162, N12161);
not NOT1 (N12163, N12146);
not NOT1 (N12164, N12163);
and AND3 (N12165, N12160, N7963, N1921);
buf BUF1 (N12166, N12159);
xor XOR2 (N12167, N12165, N4152);
and AND4 (N12168, N12154, N4368, N2855, N6517);
not NOT1 (N12169, N12158);
not NOT1 (N12170, N12166);
nand NAND3 (N12171, N12169, N4045, N9652);
nor NOR3 (N12172, N12156, N3395, N11386);
not NOT1 (N12173, N12170);
xor XOR2 (N12174, N12167, N4054);
nand NAND4 (N12175, N12164, N990, N11372, N4937);
not NOT1 (N12176, N12168);
buf BUF1 (N12177, N12162);
and AND3 (N12178, N12173, N7459, N5651);
buf BUF1 (N12179, N12139);
or OR4 (N12180, N12178, N9602, N7655, N7812);
not NOT1 (N12181, N12180);
nand NAND3 (N12182, N12176, N4250, N6924);
nand NAND2 (N12183, N12171, N7217);
not NOT1 (N12184, N12182);
nor NOR4 (N12185, N12183, N2436, N10751, N3717);
or OR2 (N12186, N12174, N6413);
not NOT1 (N12187, N12172);
buf BUF1 (N12188, N12187);
nand NAND3 (N12189, N12188, N9632, N111);
and AND4 (N12190, N12186, N9870, N536, N4066);
or OR2 (N12191, N12177, N227);
buf BUF1 (N12192, N12138);
nor NOR4 (N12193, N12175, N10055, N11882, N3467);
not NOT1 (N12194, N12185);
and AND2 (N12195, N12191, N6652);
not NOT1 (N12196, N12179);
nor NOR2 (N12197, N12195, N3714);
nand NAND2 (N12198, N12190, N3074);
not NOT1 (N12199, N12192);
and AND2 (N12200, N12196, N5165);
buf BUF1 (N12201, N12193);
nor NOR2 (N12202, N12151, N6788);
buf BUF1 (N12203, N12200);
nand NAND3 (N12204, N12203, N6500, N6576);
or OR4 (N12205, N12184, N6690, N10233, N10753);
and AND4 (N12206, N12197, N1359, N7772, N11015);
nand NAND3 (N12207, N12194, N9852, N6955);
not NOT1 (N12208, N12202);
buf BUF1 (N12209, N12207);
xor XOR2 (N12210, N12181, N3142);
nor NOR3 (N12211, N12205, N7995, N5718);
buf BUF1 (N12212, N12210);
not NOT1 (N12213, N12189);
nor NOR3 (N12214, N12209, N2270, N492);
nor NOR4 (N12215, N12214, N11824, N8216, N5578);
or OR3 (N12216, N12201, N12053, N9657);
buf BUF1 (N12217, N12199);
buf BUF1 (N12218, N12204);
not NOT1 (N12219, N12216);
buf BUF1 (N12220, N12218);
not NOT1 (N12221, N12208);
buf BUF1 (N12222, N12213);
or OR4 (N12223, N12211, N9921, N4388, N1837);
xor XOR2 (N12224, N12206, N2137);
and AND2 (N12225, N12223, N4656);
not NOT1 (N12226, N12219);
nor NOR4 (N12227, N12222, N2679, N2721, N5567);
xor XOR2 (N12228, N12217, N11712);
not NOT1 (N12229, N12226);
not NOT1 (N12230, N12221);
and AND3 (N12231, N12215, N11293, N8567);
or OR3 (N12232, N12229, N6806, N2738);
nand NAND3 (N12233, N12228, N9606, N333);
and AND3 (N12234, N12231, N1444, N8028);
buf BUF1 (N12235, N12234);
xor XOR2 (N12236, N12198, N2707);
xor XOR2 (N12237, N12230, N12077);
or OR4 (N12238, N12224, N10507, N7823, N8685);
not NOT1 (N12239, N12212);
nand NAND4 (N12240, N12237, N6536, N6865, N5163);
or OR4 (N12241, N12233, N8771, N8086, N7891);
xor XOR2 (N12242, N12235, N7940);
buf BUF1 (N12243, N12220);
not NOT1 (N12244, N12225);
nor NOR3 (N12245, N12243, N6762, N9103);
or OR3 (N12246, N12239, N4087, N8154);
xor XOR2 (N12247, N12246, N8088);
nor NOR3 (N12248, N12238, N6168, N8729);
and AND2 (N12249, N12247, N5508);
nor NOR3 (N12250, N12232, N3101, N10699);
xor XOR2 (N12251, N12242, N10555);
xor XOR2 (N12252, N12227, N2675);
or OR3 (N12253, N12244, N5928, N192);
not NOT1 (N12254, N12250);
or OR2 (N12255, N12241, N6336);
buf BUF1 (N12256, N12240);
nor NOR2 (N12257, N12252, N2611);
xor XOR2 (N12258, N12254, N2766);
and AND4 (N12259, N12258, N1787, N10500, N2606);
buf BUF1 (N12260, N12253);
nor NOR4 (N12261, N12255, N10115, N4421, N11920);
nor NOR4 (N12262, N12249, N7828, N2492, N7580);
nor NOR3 (N12263, N12236, N4405, N9999);
nor NOR4 (N12264, N12263, N1200, N4, N8752);
or OR3 (N12265, N12257, N7834, N8843);
nand NAND2 (N12266, N12261, N6820);
and AND2 (N12267, N12248, N9664);
nand NAND3 (N12268, N12245, N9202, N412);
xor XOR2 (N12269, N12264, N78);
nand NAND3 (N12270, N12265, N3049, N12227);
xor XOR2 (N12271, N12256, N3277);
xor XOR2 (N12272, N12266, N3044);
and AND2 (N12273, N12267, N7922);
not NOT1 (N12274, N12268);
nand NAND3 (N12275, N12274, N8869, N1375);
and AND3 (N12276, N12275, N9536, N8739);
and AND2 (N12277, N12276, N11280);
nor NOR4 (N12278, N12270, N149, N7669, N5968);
nand NAND4 (N12279, N12259, N1349, N9749, N12078);
or OR3 (N12280, N12279, N3098, N11000);
buf BUF1 (N12281, N12262);
not NOT1 (N12282, N12277);
and AND2 (N12283, N12282, N1464);
buf BUF1 (N12284, N12271);
or OR3 (N12285, N12269, N7288, N10265);
not NOT1 (N12286, N12283);
nor NOR4 (N12287, N12280, N3647, N5820, N6800);
nand NAND3 (N12288, N12281, N4094, N3695);
xor XOR2 (N12289, N12273, N6954);
xor XOR2 (N12290, N12287, N6369);
or OR2 (N12291, N12290, N2387);
or OR3 (N12292, N12285, N3150, N5326);
not NOT1 (N12293, N12286);
xor XOR2 (N12294, N12272, N8318);
nor NOR4 (N12295, N12260, N7714, N643, N211);
buf BUF1 (N12296, N12291);
nor NOR4 (N12297, N12296, N4905, N6657, N3463);
not NOT1 (N12298, N12284);
not NOT1 (N12299, N12292);
xor XOR2 (N12300, N12299, N9443);
nor NOR4 (N12301, N12294, N4043, N1546, N6582);
xor XOR2 (N12302, N12300, N10300);
not NOT1 (N12303, N12293);
xor XOR2 (N12304, N12301, N1952);
nor NOR2 (N12305, N12297, N6730);
not NOT1 (N12306, N12303);
and AND3 (N12307, N12288, N2829, N5077);
or OR3 (N12308, N12302, N3037, N8298);
nor NOR4 (N12309, N12305, N2935, N4455, N9086);
or OR4 (N12310, N12298, N6331, N4447, N4586);
nand NAND3 (N12311, N12310, N10083, N3920);
or OR4 (N12312, N12278, N7956, N6478, N9431);
not NOT1 (N12313, N12304);
not NOT1 (N12314, N12307);
nand NAND2 (N12315, N12312, N7574);
xor XOR2 (N12316, N12251, N9189);
and AND4 (N12317, N12309, N11565, N5055, N3780);
xor XOR2 (N12318, N12317, N5706);
xor XOR2 (N12319, N12289, N10469);
not NOT1 (N12320, N12316);
nor NOR3 (N12321, N12311, N7703, N5876);
xor XOR2 (N12322, N12295, N7147);
or OR4 (N12323, N12322, N8243, N6725, N2737);
or OR2 (N12324, N12306, N7910);
nand NAND4 (N12325, N12314, N5080, N3544, N5137);
buf BUF1 (N12326, N12325);
and AND4 (N12327, N12320, N4931, N6413, N3275);
nand NAND3 (N12328, N12318, N7728, N5229);
nor NOR3 (N12329, N12326, N1706, N2966);
buf BUF1 (N12330, N12313);
nor NOR4 (N12331, N12328, N11068, N5735, N5520);
xor XOR2 (N12332, N12315, N21);
not NOT1 (N12333, N12323);
xor XOR2 (N12334, N12308, N3637);
not NOT1 (N12335, N12321);
xor XOR2 (N12336, N12335, N6916);
or OR3 (N12337, N12333, N3286, N1078);
nor NOR4 (N12338, N12329, N7961, N3359, N7780);
buf BUF1 (N12339, N12331);
xor XOR2 (N12340, N12330, N3822);
nor NOR4 (N12341, N12339, N3489, N5940, N7834);
not NOT1 (N12342, N12327);
or OR2 (N12343, N12338, N8673);
nor NOR3 (N12344, N12319, N9737, N11502);
nor NOR2 (N12345, N12340, N7841);
nor NOR2 (N12346, N12334, N4047);
not NOT1 (N12347, N12341);
nor NOR3 (N12348, N12347, N9821, N4062);
xor XOR2 (N12349, N12346, N2621);
nand NAND3 (N12350, N12337, N11115, N239);
or OR3 (N12351, N12348, N1791, N7761);
and AND3 (N12352, N12344, N8810, N12021);
not NOT1 (N12353, N12350);
and AND3 (N12354, N12342, N3207, N4289);
or OR3 (N12355, N12332, N6048, N7010);
buf BUF1 (N12356, N12345);
nor NOR4 (N12357, N12353, N2727, N6860, N6109);
nand NAND3 (N12358, N12352, N3555, N9398);
xor XOR2 (N12359, N12357, N11447);
and AND4 (N12360, N12349, N16, N8604, N2402);
nand NAND2 (N12361, N12336, N2740);
nor NOR2 (N12362, N12324, N10719);
buf BUF1 (N12363, N12354);
and AND4 (N12364, N12361, N1654, N2461, N9127);
and AND2 (N12365, N12351, N9727);
and AND3 (N12366, N12360, N10179, N6139);
or OR2 (N12367, N12366, N6873);
xor XOR2 (N12368, N12362, N2917);
nor NOR3 (N12369, N12364, N1058, N11185);
or OR3 (N12370, N12359, N11871, N8330);
nor NOR2 (N12371, N12343, N8161);
nand NAND4 (N12372, N12363, N6933, N9715, N8966);
buf BUF1 (N12373, N12358);
or OR4 (N12374, N12370, N1572, N2262, N6949);
nor NOR3 (N12375, N12372, N3803, N1592);
and AND2 (N12376, N12374, N997);
xor XOR2 (N12377, N12356, N419);
or OR2 (N12378, N12377, N9157);
or OR4 (N12379, N12365, N8594, N7096, N2497);
nand NAND2 (N12380, N12355, N11395);
nor NOR3 (N12381, N12373, N8414, N7570);
nor NOR4 (N12382, N12368, N11690, N2981, N7368);
not NOT1 (N12383, N12382);
xor XOR2 (N12384, N12371, N8040);
nand NAND4 (N12385, N12383, N2090, N11088, N6882);
and AND3 (N12386, N12369, N5754, N2826);
and AND2 (N12387, N12379, N3045);
nand NAND2 (N12388, N12385, N9999);
nand NAND2 (N12389, N12375, N10158);
nor NOR4 (N12390, N12367, N10613, N10624, N1971);
and AND3 (N12391, N12376, N11905, N7209);
buf BUF1 (N12392, N12391);
buf BUF1 (N12393, N12389);
and AND4 (N12394, N12387, N8162, N6560, N2023);
or OR2 (N12395, N12394, N6629);
and AND4 (N12396, N12390, N2521, N4199, N11707);
xor XOR2 (N12397, N12388, N1613);
or OR3 (N12398, N12384, N12377, N5289);
or OR4 (N12399, N12381, N7381, N8530, N6037);
nand NAND2 (N12400, N12396, N11198);
xor XOR2 (N12401, N12393, N8512);
buf BUF1 (N12402, N12399);
nand NAND2 (N12403, N12386, N7938);
xor XOR2 (N12404, N12402, N9104);
buf BUF1 (N12405, N12395);
nand NAND4 (N12406, N12401, N752, N8817, N4852);
nand NAND3 (N12407, N12406, N11463, N2345);
buf BUF1 (N12408, N12407);
not NOT1 (N12409, N12392);
buf BUF1 (N12410, N12378);
nand NAND3 (N12411, N12405, N1513, N6374);
or OR3 (N12412, N12397, N11922, N3630);
and AND4 (N12413, N12408, N1636, N11948, N5398);
nand NAND3 (N12414, N12410, N4754, N2386);
nor NOR4 (N12415, N12398, N11289, N5599, N8155);
nand NAND4 (N12416, N12413, N11121, N11370, N6969);
and AND2 (N12417, N12403, N3412);
nand NAND4 (N12418, N12412, N9919, N12063, N4589);
or OR3 (N12419, N12416, N10224, N368);
xor XOR2 (N12420, N12414, N11507);
nand NAND3 (N12421, N12380, N8959, N3843);
nor NOR3 (N12422, N12419, N8958, N3509);
nand NAND4 (N12423, N12409, N5293, N1533, N4265);
xor XOR2 (N12424, N12421, N5964);
or OR2 (N12425, N12417, N3940);
not NOT1 (N12426, N12424);
nand NAND3 (N12427, N12400, N7580, N11967);
or OR3 (N12428, N12404, N7960, N9700);
nor NOR2 (N12429, N12411, N10118);
or OR4 (N12430, N12418, N9449, N6170, N2567);
nand NAND3 (N12431, N12422, N9152, N5566);
and AND2 (N12432, N12428, N4257);
and AND4 (N12433, N12415, N6534, N6252, N11266);
and AND2 (N12434, N12429, N11619);
nand NAND3 (N12435, N12425, N10357, N1453);
and AND3 (N12436, N12427, N1692, N7024);
nand NAND4 (N12437, N12436, N10303, N5559, N5876);
buf BUF1 (N12438, N12434);
not NOT1 (N12439, N12431);
or OR3 (N12440, N12439, N2008, N6221);
or OR2 (N12441, N12437, N6943);
not NOT1 (N12442, N12438);
nand NAND3 (N12443, N12441, N7932, N4017);
or OR3 (N12444, N12442, N4157, N9541);
buf BUF1 (N12445, N12433);
nor NOR3 (N12446, N12426, N7096, N218);
nor NOR3 (N12447, N12423, N4822, N3516);
nor NOR3 (N12448, N12444, N11465, N904);
nor NOR3 (N12449, N12420, N2161, N2587);
nand NAND3 (N12450, N12446, N2426, N9136);
or OR2 (N12451, N12447, N3217);
xor XOR2 (N12452, N12443, N5849);
or OR4 (N12453, N12449, N12317, N10742, N193);
and AND2 (N12454, N12435, N3499);
and AND2 (N12455, N12430, N3239);
nand NAND4 (N12456, N12455, N6069, N4856, N4741);
xor XOR2 (N12457, N12454, N9685);
buf BUF1 (N12458, N12440);
and AND2 (N12459, N12453, N7667);
nor NOR2 (N12460, N12432, N283);
xor XOR2 (N12461, N12456, N9405);
or OR3 (N12462, N12457, N7729, N6675);
and AND4 (N12463, N12451, N4778, N5857, N11715);
or OR3 (N12464, N12445, N6402, N7614);
buf BUF1 (N12465, N12458);
xor XOR2 (N12466, N12464, N343);
and AND4 (N12467, N12461, N5558, N2484, N6570);
or OR2 (N12468, N12459, N6408);
not NOT1 (N12469, N12448);
not NOT1 (N12470, N12469);
xor XOR2 (N12471, N12466, N7470);
not NOT1 (N12472, N12463);
and AND3 (N12473, N12470, N2151, N2641);
not NOT1 (N12474, N12452);
and AND4 (N12475, N12450, N5215, N6777, N6734);
and AND3 (N12476, N12472, N1983, N1236);
or OR2 (N12477, N12475, N2451);
or OR3 (N12478, N12471, N1116, N2611);
or OR3 (N12479, N12477, N3270, N10374);
and AND3 (N12480, N12460, N10224, N8961);
nor NOR4 (N12481, N12465, N9246, N10205, N8070);
buf BUF1 (N12482, N12462);
nand NAND3 (N12483, N12467, N4670, N3336);
buf BUF1 (N12484, N12473);
xor XOR2 (N12485, N12479, N4829);
xor XOR2 (N12486, N12468, N10415);
and AND2 (N12487, N12482, N5684);
nor NOR3 (N12488, N12486, N1122, N8744);
nand NAND4 (N12489, N12487, N817, N9714, N971);
buf BUF1 (N12490, N12476);
nor NOR4 (N12491, N12484, N222, N2074, N2857);
or OR3 (N12492, N12478, N4034, N10100);
not NOT1 (N12493, N12489);
nand NAND2 (N12494, N12481, N5613);
nand NAND3 (N12495, N12493, N8680, N10014);
or OR2 (N12496, N12483, N8798);
or OR2 (N12497, N12494, N2122);
not NOT1 (N12498, N12497);
not NOT1 (N12499, N12496);
and AND2 (N12500, N12498, N503);
not NOT1 (N12501, N12474);
not NOT1 (N12502, N12490);
buf BUF1 (N12503, N12480);
buf BUF1 (N12504, N12500);
nor NOR3 (N12505, N12499, N7492, N8074);
nand NAND2 (N12506, N12504, N10958);
or OR2 (N12507, N12492, N10226);
buf BUF1 (N12508, N12488);
buf BUF1 (N12509, N12495);
xor XOR2 (N12510, N12485, N7753);
buf BUF1 (N12511, N12491);
or OR4 (N12512, N12507, N5144, N9713, N8774);
xor XOR2 (N12513, N12510, N6376);
not NOT1 (N12514, N12512);
nor NOR2 (N12515, N12503, N12212);
buf BUF1 (N12516, N12514);
buf BUF1 (N12517, N12516);
or OR2 (N12518, N12506, N8031);
buf BUF1 (N12519, N12513);
and AND3 (N12520, N12502, N12125, N4637);
nor NOR4 (N12521, N12518, N8951, N3194, N9170);
not NOT1 (N12522, N12505);
buf BUF1 (N12523, N12520);
xor XOR2 (N12524, N12517, N12430);
buf BUF1 (N12525, N12522);
buf BUF1 (N12526, N12521);
or OR3 (N12527, N12509, N12097, N11378);
nor NOR3 (N12528, N12508, N6412, N6913);
or OR2 (N12529, N12525, N5612);
nand NAND4 (N12530, N12501, N4136, N7748, N2901);
or OR3 (N12531, N12519, N3720, N11283);
buf BUF1 (N12532, N12528);
nor NOR3 (N12533, N12529, N2993, N8023);
nor NOR3 (N12534, N12533, N11125, N9162);
xor XOR2 (N12535, N12511, N4053);
and AND2 (N12536, N12531, N2644);
buf BUF1 (N12537, N12524);
not NOT1 (N12538, N12523);
not NOT1 (N12539, N12527);
nor NOR3 (N12540, N12530, N5153, N11114);
buf BUF1 (N12541, N12540);
xor XOR2 (N12542, N12515, N2993);
or OR2 (N12543, N12538, N6402);
not NOT1 (N12544, N12542);
buf BUF1 (N12545, N12543);
buf BUF1 (N12546, N12541);
buf BUF1 (N12547, N12544);
and AND3 (N12548, N12539, N9627, N1837);
nand NAND3 (N12549, N12526, N6534, N11186);
nor NOR3 (N12550, N12546, N3475, N9568);
and AND3 (N12551, N12547, N1789, N7914);
nand NAND2 (N12552, N12535, N5474);
buf BUF1 (N12553, N12550);
and AND3 (N12554, N12532, N12457, N12172);
nand NAND2 (N12555, N12554, N3174);
xor XOR2 (N12556, N12549, N10431);
nor NOR3 (N12557, N12553, N11668, N7594);
not NOT1 (N12558, N12548);
buf BUF1 (N12559, N12537);
or OR4 (N12560, N12558, N6314, N10689, N10746);
and AND3 (N12561, N12559, N12190, N6916);
or OR4 (N12562, N12551, N3293, N2595, N578);
or OR2 (N12563, N12555, N3290);
or OR4 (N12564, N12563, N95, N8617, N5497);
nand NAND4 (N12565, N12556, N2692, N2054, N5439);
or OR4 (N12566, N12536, N12522, N5397, N4325);
or OR4 (N12567, N12561, N7383, N10541, N1436);
or OR3 (N12568, N12545, N6402, N1092);
not NOT1 (N12569, N12566);
buf BUF1 (N12570, N12534);
nor NOR4 (N12571, N12552, N5967, N3424, N5729);
not NOT1 (N12572, N12557);
and AND2 (N12573, N12567, N510);
nand NAND3 (N12574, N12570, N6360, N2455);
buf BUF1 (N12575, N12569);
nor NOR3 (N12576, N12568, N12227, N259);
xor XOR2 (N12577, N12571, N8832);
not NOT1 (N12578, N12573);
buf BUF1 (N12579, N12578);
nor NOR4 (N12580, N12576, N5164, N134, N7245);
nand NAND2 (N12581, N12562, N1246);
nand NAND4 (N12582, N12581, N961, N1461, N8685);
buf BUF1 (N12583, N12579);
or OR2 (N12584, N12577, N593);
xor XOR2 (N12585, N12565, N3202);
or OR3 (N12586, N12585, N328, N10100);
and AND2 (N12587, N12564, N1413);
and AND4 (N12588, N12584, N4637, N1031, N5195);
or OR3 (N12589, N12574, N2299, N3976);
xor XOR2 (N12590, N12589, N6875);
or OR4 (N12591, N12580, N11054, N12428, N8761);
nor NOR3 (N12592, N12591, N8016, N5286);
xor XOR2 (N12593, N12560, N9106);
and AND3 (N12594, N12586, N5178, N3630);
not NOT1 (N12595, N12587);
nand NAND3 (N12596, N12592, N5289, N10426);
xor XOR2 (N12597, N12594, N11146);
or OR2 (N12598, N12572, N1941);
not NOT1 (N12599, N12598);
xor XOR2 (N12600, N12593, N8558);
nor NOR4 (N12601, N12588, N3223, N6349, N6158);
nor NOR2 (N12602, N12600, N2181);
buf BUF1 (N12603, N12590);
not NOT1 (N12604, N12595);
buf BUF1 (N12605, N12603);
nor NOR4 (N12606, N12582, N9530, N988, N2034);
buf BUF1 (N12607, N12606);
not NOT1 (N12608, N12607);
buf BUF1 (N12609, N12608);
and AND4 (N12610, N12597, N7950, N7953, N7936);
and AND4 (N12611, N12609, N222, N9562, N215);
or OR3 (N12612, N12611, N9810, N5867);
and AND4 (N12613, N12610, N9880, N6809, N5537);
buf BUF1 (N12614, N12602);
or OR2 (N12615, N12604, N5970);
not NOT1 (N12616, N12612);
and AND2 (N12617, N12605, N9266);
buf BUF1 (N12618, N12583);
nand NAND4 (N12619, N12613, N9412, N8645, N1541);
buf BUF1 (N12620, N12618);
nand NAND3 (N12621, N12614, N8601, N2030);
not NOT1 (N12622, N12615);
nor NOR4 (N12623, N12601, N8053, N10746, N8356);
buf BUF1 (N12624, N12575);
not NOT1 (N12625, N12596);
or OR4 (N12626, N12619, N3179, N8298, N8763);
xor XOR2 (N12627, N12626, N5052);
nor NOR4 (N12628, N12617, N12586, N755, N6935);
buf BUF1 (N12629, N12625);
or OR2 (N12630, N12623, N11792);
nor NOR4 (N12631, N12620, N96, N6558, N4280);
nor NOR2 (N12632, N12630, N11626);
and AND4 (N12633, N12599, N11786, N1029, N9482);
nand NAND2 (N12634, N12616, N10825);
not NOT1 (N12635, N12622);
nor NOR3 (N12636, N12628, N9818, N12303);
nand NAND4 (N12637, N12621, N4515, N8899, N8679);
nand NAND4 (N12638, N12631, N10929, N9774, N5032);
nand NAND2 (N12639, N12634, N9262);
nand NAND2 (N12640, N12624, N11000);
not NOT1 (N12641, N12639);
buf BUF1 (N12642, N12636);
nand NAND2 (N12643, N12632, N12332);
nand NAND4 (N12644, N12629, N1927, N10698, N4862);
not NOT1 (N12645, N12640);
xor XOR2 (N12646, N12643, N5265);
and AND4 (N12647, N12641, N1844, N8106, N11904);
not NOT1 (N12648, N12627);
not NOT1 (N12649, N12647);
not NOT1 (N12650, N12644);
xor XOR2 (N12651, N12637, N11364);
nand NAND4 (N12652, N12651, N8165, N7711, N3203);
nand NAND3 (N12653, N12650, N844, N8666);
nor NOR3 (N12654, N12653, N641, N6224);
or OR4 (N12655, N12652, N3825, N6488, N5021);
and AND4 (N12656, N12645, N4982, N5425, N11616);
nor NOR4 (N12657, N12642, N6991, N12334, N2227);
xor XOR2 (N12658, N12657, N3335);
buf BUF1 (N12659, N12638);
and AND2 (N12660, N12655, N3294);
xor XOR2 (N12661, N12649, N5243);
buf BUF1 (N12662, N12660);
buf BUF1 (N12663, N12661);
or OR3 (N12664, N12663, N2386, N8131);
buf BUF1 (N12665, N12654);
buf BUF1 (N12666, N12664);
and AND3 (N12667, N12635, N5505, N2492);
and AND2 (N12668, N12662, N7233);
and AND3 (N12669, N12646, N7590, N8770);
or OR2 (N12670, N12659, N7312);
or OR3 (N12671, N12666, N3217, N137);
buf BUF1 (N12672, N12669);
buf BUF1 (N12673, N12670);
buf BUF1 (N12674, N12658);
xor XOR2 (N12675, N12648, N5239);
xor XOR2 (N12676, N12673, N1660);
not NOT1 (N12677, N12668);
nor NOR2 (N12678, N12676, N7964);
and AND3 (N12679, N12665, N7707, N6971);
nand NAND2 (N12680, N12678, N344);
nand NAND4 (N12681, N12677, N5634, N1735, N12224);
nand NAND4 (N12682, N12633, N587, N912, N4340);
and AND3 (N12683, N12680, N130, N11463);
not NOT1 (N12684, N12681);
or OR2 (N12685, N12679, N12669);
buf BUF1 (N12686, N12672);
nand NAND3 (N12687, N12684, N11951, N4115);
xor XOR2 (N12688, N12683, N2799);
and AND2 (N12689, N12687, N1535);
nor NOR2 (N12690, N12689, N7545);
nor NOR2 (N12691, N12675, N4099);
buf BUF1 (N12692, N12674);
not NOT1 (N12693, N12667);
nor NOR2 (N12694, N12690, N6702);
not NOT1 (N12695, N12682);
or OR2 (N12696, N12693, N9567);
nand NAND2 (N12697, N12696, N8621);
and AND4 (N12698, N12697, N7811, N6598, N9322);
and AND2 (N12699, N12685, N2310);
nand NAND2 (N12700, N12688, N1308);
xor XOR2 (N12701, N12699, N10514);
and AND3 (N12702, N12694, N5090, N1878);
or OR2 (N12703, N12698, N1525);
buf BUF1 (N12704, N12691);
not NOT1 (N12705, N12695);
or OR3 (N12706, N12701, N9995, N11587);
buf BUF1 (N12707, N12656);
nand NAND4 (N12708, N12671, N9138, N8234, N8197);
nand NAND2 (N12709, N12700, N5465);
or OR3 (N12710, N12706, N2622, N5311);
not NOT1 (N12711, N12709);
buf BUF1 (N12712, N12711);
not NOT1 (N12713, N12686);
not NOT1 (N12714, N12713);
nand NAND2 (N12715, N12712, N11005);
and AND3 (N12716, N12702, N497, N5744);
or OR3 (N12717, N12708, N2643, N5200);
xor XOR2 (N12718, N12707, N1708);
nor NOR4 (N12719, N12704, N3039, N6632, N9272);
xor XOR2 (N12720, N12717, N8597);
buf BUF1 (N12721, N12705);
and AND3 (N12722, N12710, N1028, N5066);
nor NOR3 (N12723, N12720, N7009, N4491);
xor XOR2 (N12724, N12722, N4573);
and AND3 (N12725, N12703, N3, N12328);
buf BUF1 (N12726, N12716);
buf BUF1 (N12727, N12718);
not NOT1 (N12728, N12721);
and AND2 (N12729, N12724, N1729);
or OR4 (N12730, N12728, N7358, N6741, N1697);
and AND3 (N12731, N12725, N3490, N5525);
xor XOR2 (N12732, N12731, N8699);
buf BUF1 (N12733, N12729);
and AND2 (N12734, N12692, N3179);
not NOT1 (N12735, N12727);
nor NOR2 (N12736, N12726, N11245);
xor XOR2 (N12737, N12723, N10263);
nor NOR4 (N12738, N12734, N4060, N3302, N11878);
not NOT1 (N12739, N12735);
xor XOR2 (N12740, N12738, N386);
nor NOR4 (N12741, N12715, N8745, N11650, N573);
or OR2 (N12742, N12719, N994);
xor XOR2 (N12743, N12730, N10312);
and AND2 (N12744, N12733, N10497);
nand NAND2 (N12745, N12732, N836);
and AND3 (N12746, N12739, N10202, N10451);
xor XOR2 (N12747, N12746, N3897);
buf BUF1 (N12748, N12740);
nand NAND2 (N12749, N12714, N3711);
not NOT1 (N12750, N12743);
buf BUF1 (N12751, N12747);
not NOT1 (N12752, N12745);
and AND3 (N12753, N12751, N2317, N6248);
and AND2 (N12754, N12744, N8027);
buf BUF1 (N12755, N12749);
nor NOR4 (N12756, N12753, N5046, N12434, N659);
nand NAND2 (N12757, N12736, N7295);
buf BUF1 (N12758, N12741);
not NOT1 (N12759, N12756);
buf BUF1 (N12760, N12737);
and AND2 (N12761, N12742, N6675);
and AND4 (N12762, N12759, N2541, N7479, N9784);
nor NOR2 (N12763, N12755, N742);
buf BUF1 (N12764, N12754);
nor NOR3 (N12765, N12762, N2704, N6829);
xor XOR2 (N12766, N12761, N8999);
nor NOR4 (N12767, N12748, N10073, N9316, N9088);
xor XOR2 (N12768, N12757, N9344);
buf BUF1 (N12769, N12752);
or OR4 (N12770, N12766, N11474, N674, N2314);
nand NAND4 (N12771, N12767, N12132, N9841, N2374);
xor XOR2 (N12772, N12768, N499);
and AND2 (N12773, N12750, N6245);
buf BUF1 (N12774, N12760);
buf BUF1 (N12775, N12772);
nor NOR4 (N12776, N12764, N309, N11223, N4377);
not NOT1 (N12777, N12765);
nor NOR2 (N12778, N12771, N9850);
nor NOR4 (N12779, N12775, N8756, N5283, N1835);
nor NOR4 (N12780, N12774, N8673, N3902, N8075);
buf BUF1 (N12781, N12770);
buf BUF1 (N12782, N12763);
and AND3 (N12783, N12776, N12188, N8355);
buf BUF1 (N12784, N12777);
xor XOR2 (N12785, N12784, N1849);
buf BUF1 (N12786, N12769);
not NOT1 (N12787, N12782);
buf BUF1 (N12788, N12780);
not NOT1 (N12789, N12783);
and AND3 (N12790, N12786, N8979, N10950);
or OR3 (N12791, N12785, N9451, N1277);
nand NAND4 (N12792, N12791, N7860, N5156, N12134);
and AND4 (N12793, N12779, N12452, N9293, N1853);
or OR2 (N12794, N12789, N12064);
nor NOR3 (N12795, N12792, N6707, N7379);
xor XOR2 (N12796, N12788, N7222);
or OR2 (N12797, N12796, N6342);
buf BUF1 (N12798, N12794);
and AND4 (N12799, N12795, N8048, N7505, N11585);
nor NOR4 (N12800, N12778, N6186, N11314, N3501);
nor NOR3 (N12801, N12773, N714, N8201);
nand NAND3 (N12802, N12799, N4556, N2170);
nor NOR3 (N12803, N12781, N2014, N4422);
buf BUF1 (N12804, N12802);
and AND4 (N12805, N12797, N10550, N3763, N3793);
and AND4 (N12806, N12758, N2225, N4926, N5424);
nand NAND4 (N12807, N12804, N11777, N4631, N3489);
nor NOR4 (N12808, N12806, N845, N7734, N10019);
nand NAND2 (N12809, N12800, N10655);
not NOT1 (N12810, N12801);
nor NOR2 (N12811, N12807, N9180);
and AND3 (N12812, N12808, N912, N11177);
not NOT1 (N12813, N12805);
xor XOR2 (N12814, N12787, N1135);
xor XOR2 (N12815, N12798, N11817);
not NOT1 (N12816, N12815);
buf BUF1 (N12817, N12810);
xor XOR2 (N12818, N12814, N3868);
xor XOR2 (N12819, N12817, N10943);
buf BUF1 (N12820, N12803);
not NOT1 (N12821, N12816);
or OR4 (N12822, N12790, N1776, N3588, N11435);
xor XOR2 (N12823, N12822, N11561);
nand NAND4 (N12824, N12821, N9388, N12226, N6073);
or OR3 (N12825, N12809, N6532, N2414);
buf BUF1 (N12826, N12818);
not NOT1 (N12827, N12825);
nor NOR3 (N12828, N12811, N11918, N2214);
not NOT1 (N12829, N12793);
xor XOR2 (N12830, N12820, N3593);
xor XOR2 (N12831, N12823, N12403);
buf BUF1 (N12832, N12828);
and AND2 (N12833, N12832, N149);
nand NAND4 (N12834, N12812, N9222, N3746, N8673);
buf BUF1 (N12835, N12830);
nand NAND4 (N12836, N12833, N754, N6981, N11571);
and AND3 (N12837, N12834, N8781, N11526);
buf BUF1 (N12838, N12819);
buf BUF1 (N12839, N12831);
xor XOR2 (N12840, N12838, N6133);
nand NAND2 (N12841, N12837, N5370);
xor XOR2 (N12842, N12839, N4334);
and AND2 (N12843, N12826, N8482);
or OR3 (N12844, N12827, N10070, N101);
not NOT1 (N12845, N12840);
and AND4 (N12846, N12824, N11442, N9876, N12722);
xor XOR2 (N12847, N12836, N1175);
or OR2 (N12848, N12841, N6973);
not NOT1 (N12849, N12844);
not NOT1 (N12850, N12845);
xor XOR2 (N12851, N12813, N3208);
not NOT1 (N12852, N12848);
nand NAND4 (N12853, N12846, N77, N10150, N1177);
or OR4 (N12854, N12835, N511, N9865, N1943);
buf BUF1 (N12855, N12853);
xor XOR2 (N12856, N12829, N8236);
xor XOR2 (N12857, N12851, N136);
or OR2 (N12858, N12843, N8357);
or OR2 (N12859, N12847, N9510);
or OR3 (N12860, N12852, N10775, N5536);
and AND2 (N12861, N12854, N780);
not NOT1 (N12862, N12860);
and AND3 (N12863, N12842, N4409, N4494);
or OR3 (N12864, N12855, N9763, N6776);
nand NAND4 (N12865, N12858, N11005, N1205, N8095);
or OR2 (N12866, N12863, N4489);
and AND3 (N12867, N12861, N11621, N9807);
buf BUF1 (N12868, N12857);
buf BUF1 (N12869, N12862);
xor XOR2 (N12870, N12865, N10416);
buf BUF1 (N12871, N12869);
not NOT1 (N12872, N12864);
xor XOR2 (N12873, N12867, N10227);
nor NOR4 (N12874, N12870, N6384, N1766, N3276);
not NOT1 (N12875, N12872);
and AND4 (N12876, N12866, N1818, N9648, N456);
not NOT1 (N12877, N12849);
xor XOR2 (N12878, N12877, N7686);
or OR2 (N12879, N12856, N8391);
and AND4 (N12880, N12876, N3285, N10909, N2781);
and AND4 (N12881, N12868, N9473, N8106, N1887);
and AND3 (N12882, N12874, N6392, N9496);
buf BUF1 (N12883, N12850);
nor NOR4 (N12884, N12879, N6467, N4340, N316);
nor NOR4 (N12885, N12881, N9788, N2461, N5621);
not NOT1 (N12886, N12882);
nand NAND4 (N12887, N12880, N7563, N62, N8197);
xor XOR2 (N12888, N12885, N7876);
and AND4 (N12889, N12859, N5150, N3515, N12424);
not NOT1 (N12890, N12887);
not NOT1 (N12891, N12884);
nor NOR2 (N12892, N12891, N2321);
xor XOR2 (N12893, N12875, N7760);
nand NAND3 (N12894, N12883, N2335, N9644);
or OR2 (N12895, N12893, N6576);
and AND3 (N12896, N12894, N9454, N4114);
buf BUF1 (N12897, N12896);
xor XOR2 (N12898, N12889, N11662);
xor XOR2 (N12899, N12890, N59);
nor NOR2 (N12900, N12878, N7475);
buf BUF1 (N12901, N12895);
not NOT1 (N12902, N12899);
and AND3 (N12903, N12871, N6602, N4299);
buf BUF1 (N12904, N12888);
nor NOR4 (N12905, N12901, N4476, N7795, N1469);
and AND4 (N12906, N12904, N10973, N5528, N7946);
and AND2 (N12907, N12897, N1853);
nand NAND3 (N12908, N12902, N5658, N4020);
xor XOR2 (N12909, N12898, N8222);
not NOT1 (N12910, N12905);
or OR2 (N12911, N12900, N3607);
nor NOR3 (N12912, N12909, N3993, N1011);
nand NAND2 (N12913, N12907, N3408);
buf BUF1 (N12914, N12912);
nand NAND3 (N12915, N12914, N3359, N1485);
nor NOR4 (N12916, N12906, N7296, N2094, N4073);
buf BUF1 (N12917, N12908);
buf BUF1 (N12918, N12916);
not NOT1 (N12919, N12903);
or OR3 (N12920, N12892, N10767, N11803);
nand NAND4 (N12921, N12910, N2520, N2684, N3550);
nand NAND3 (N12922, N12921, N10617, N8229);
buf BUF1 (N12923, N12873);
or OR4 (N12924, N12923, N4570, N7652, N3396);
nand NAND2 (N12925, N12911, N5682);
nand NAND2 (N12926, N12913, N2713);
xor XOR2 (N12927, N12926, N8027);
xor XOR2 (N12928, N12924, N6623);
nand NAND3 (N12929, N12927, N3608, N11608);
buf BUF1 (N12930, N12918);
not NOT1 (N12931, N12928);
and AND2 (N12932, N12915, N4308);
nand NAND2 (N12933, N12917, N10960);
and AND3 (N12934, N12919, N6836, N12037);
and AND4 (N12935, N12934, N7909, N6594, N4474);
nand NAND3 (N12936, N12925, N12014, N3171);
buf BUF1 (N12937, N12922);
or OR4 (N12938, N12933, N3232, N4224, N6162);
or OR3 (N12939, N12938, N712, N6422);
buf BUF1 (N12940, N12931);
and AND3 (N12941, N12920, N3620, N4267);
not NOT1 (N12942, N12935);
nor NOR3 (N12943, N12936, N10224, N6584);
nand NAND4 (N12944, N12932, N7732, N8094, N1573);
buf BUF1 (N12945, N12929);
nand NAND3 (N12946, N12945, N7687, N9072);
xor XOR2 (N12947, N12943, N11813);
not NOT1 (N12948, N12937);
nand NAND2 (N12949, N12948, N2902);
not NOT1 (N12950, N12944);
or OR3 (N12951, N12949, N486, N6479);
or OR4 (N12952, N12947, N10653, N971, N8519);
not NOT1 (N12953, N12952);
and AND3 (N12954, N12951, N11759, N8695);
nand NAND3 (N12955, N12940, N650, N5418);
buf BUF1 (N12956, N12930);
not NOT1 (N12957, N12939);
buf BUF1 (N12958, N12956);
buf BUF1 (N12959, N12955);
buf BUF1 (N12960, N12886);
nor NOR2 (N12961, N12950, N9139);
and AND4 (N12962, N12942, N3989, N5698, N10147);
or OR2 (N12963, N12959, N898);
not NOT1 (N12964, N12958);
or OR2 (N12965, N12946, N3011);
xor XOR2 (N12966, N12964, N5793);
and AND3 (N12967, N12963, N4097, N6261);
buf BUF1 (N12968, N12957);
xor XOR2 (N12969, N12967, N9332);
nor NOR2 (N12970, N12966, N12451);
not NOT1 (N12971, N12961);
xor XOR2 (N12972, N12970, N120);
or OR4 (N12973, N12960, N9184, N7834, N3887);
xor XOR2 (N12974, N12973, N1277);
and AND2 (N12975, N12972, N12466);
or OR2 (N12976, N12968, N7731);
xor XOR2 (N12977, N12941, N3723);
xor XOR2 (N12978, N12971, N12284);
xor XOR2 (N12979, N12965, N2129);
or OR3 (N12980, N12969, N6577, N9384);
or OR3 (N12981, N12977, N2751, N4326);
nor NOR4 (N12982, N12974, N9173, N6577, N10134);
buf BUF1 (N12983, N12976);
or OR3 (N12984, N12981, N9433, N11951);
nand NAND3 (N12985, N12980, N7371, N428);
not NOT1 (N12986, N12954);
or OR3 (N12987, N12985, N12570, N937);
or OR4 (N12988, N12986, N8859, N1928, N5779);
nand NAND4 (N12989, N12975, N4373, N10176, N5988);
nor NOR2 (N12990, N12953, N3395);
nor NOR3 (N12991, N12990, N5707, N7523);
nand NAND3 (N12992, N12982, N834, N11717);
nand NAND3 (N12993, N12979, N5317, N11625);
nor NOR3 (N12994, N12993, N443, N1283);
nand NAND4 (N12995, N12978, N6349, N2256, N12448);
and AND4 (N12996, N12984, N359, N554, N3755);
nand NAND4 (N12997, N12989, N8856, N12224, N273);
and AND3 (N12998, N12962, N5255, N11667);
buf BUF1 (N12999, N12987);
xor XOR2 (N13000, N12995, N827);
xor XOR2 (N13001, N12983, N12002);
and AND4 (N13002, N12988, N11407, N9742, N6261);
not NOT1 (N13003, N13000);
not NOT1 (N13004, N12997);
nor NOR3 (N13005, N12991, N7620, N12346);
nand NAND3 (N13006, N12996, N1454, N11475);
xor XOR2 (N13007, N12998, N2158);
not NOT1 (N13008, N13002);
xor XOR2 (N13009, N13007, N5694);
not NOT1 (N13010, N13008);
not NOT1 (N13011, N12992);
nand NAND2 (N13012, N12999, N2729);
xor XOR2 (N13013, N12994, N6536);
xor XOR2 (N13014, N13004, N4386);
nor NOR3 (N13015, N13013, N12426, N6383);
buf BUF1 (N13016, N13006);
or OR2 (N13017, N13015, N2892);
or OR3 (N13018, N13010, N2072, N7063);
nor NOR3 (N13019, N13005, N11831, N4647);
nand NAND3 (N13020, N13001, N9324, N12428);
buf BUF1 (N13021, N13014);
or OR4 (N13022, N13019, N12674, N102, N10058);
and AND2 (N13023, N13018, N5558);
nand NAND2 (N13024, N13021, N2631);
and AND2 (N13025, N13022, N4247);
or OR4 (N13026, N13024, N10973, N4363, N6040);
and AND2 (N13027, N13009, N11670);
not NOT1 (N13028, N13012);
not NOT1 (N13029, N13025);
xor XOR2 (N13030, N13028, N2109);
nor NOR2 (N13031, N13030, N5250);
xor XOR2 (N13032, N13020, N10649);
and AND3 (N13033, N13032, N10077, N12774);
or OR4 (N13034, N13003, N6044, N1173, N2083);
nand NAND3 (N13035, N13027, N10565, N7264);
or OR3 (N13036, N13033, N5596, N6305);
buf BUF1 (N13037, N13023);
nand NAND4 (N13038, N13031, N7955, N9939, N3629);
nand NAND2 (N13039, N13016, N9641);
or OR4 (N13040, N13011, N2179, N5148, N2675);
buf BUF1 (N13041, N13038);
and AND3 (N13042, N13040, N5400, N12200);
xor XOR2 (N13043, N13029, N8196);
xor XOR2 (N13044, N13036, N471);
xor XOR2 (N13045, N13043, N3618);
not NOT1 (N13046, N13039);
nand NAND2 (N13047, N13034, N5326);
xor XOR2 (N13048, N13046, N5730);
or OR2 (N13049, N13042, N7163);
and AND4 (N13050, N13041, N3589, N6712, N11266);
and AND4 (N13051, N13048, N4916, N10841, N10308);
buf BUF1 (N13052, N13017);
buf BUF1 (N13053, N13052);
not NOT1 (N13054, N13037);
buf BUF1 (N13055, N13054);
nand NAND2 (N13056, N13045, N1859);
not NOT1 (N13057, N13049);
or OR3 (N13058, N13057, N8374, N9985);
and AND3 (N13059, N13055, N2897, N9270);
or OR2 (N13060, N13058, N8899);
nor NOR2 (N13061, N13053, N9571);
buf BUF1 (N13062, N13026);
not NOT1 (N13063, N13050);
xor XOR2 (N13064, N13063, N7142);
buf BUF1 (N13065, N13035);
not NOT1 (N13066, N13047);
xor XOR2 (N13067, N13059, N7870);
buf BUF1 (N13068, N13060);
nand NAND3 (N13069, N13051, N12047, N11616);
and AND2 (N13070, N13068, N5016);
xor XOR2 (N13071, N13056, N12070);
xor XOR2 (N13072, N13064, N9724);
buf BUF1 (N13073, N13070);
nand NAND3 (N13074, N13065, N10960, N3296);
and AND2 (N13075, N13062, N11590);
nand NAND4 (N13076, N13074, N8417, N8931, N392);
or OR3 (N13077, N13069, N1067, N11331);
or OR3 (N13078, N13077, N5080, N2224);
not NOT1 (N13079, N13061);
or OR2 (N13080, N13072, N11123);
or OR2 (N13081, N13066, N2900);
xor XOR2 (N13082, N13079, N9633);
xor XOR2 (N13083, N13071, N3807);
not NOT1 (N13084, N13082);
buf BUF1 (N13085, N13081);
and AND4 (N13086, N13083, N7621, N12434, N1458);
not NOT1 (N13087, N13067);
and AND2 (N13088, N13080, N7492);
or OR3 (N13089, N13086, N9472, N4443);
or OR3 (N13090, N13084, N8706, N4803);
or OR2 (N13091, N13078, N1913);
and AND4 (N13092, N13075, N2935, N12900, N1014);
xor XOR2 (N13093, N13090, N752);
and AND4 (N13094, N13085, N827, N6, N7443);
not NOT1 (N13095, N13088);
nand NAND4 (N13096, N13076, N7425, N9671, N10537);
nand NAND3 (N13097, N13087, N3311, N4625);
nand NAND2 (N13098, N13095, N3669);
xor XOR2 (N13099, N13097, N2765);
nand NAND2 (N13100, N13091, N9235);
xor XOR2 (N13101, N13044, N4202);
and AND2 (N13102, N13092, N3068);
or OR4 (N13103, N13101, N3339, N2804, N1505);
xor XOR2 (N13104, N13103, N9723);
and AND4 (N13105, N13094, N3294, N9467, N12938);
buf BUF1 (N13106, N13099);
not NOT1 (N13107, N13093);
buf BUF1 (N13108, N13107);
xor XOR2 (N13109, N13105, N3312);
not NOT1 (N13110, N13109);
not NOT1 (N13111, N13073);
xor XOR2 (N13112, N13111, N347);
xor XOR2 (N13113, N13106, N9260);
xor XOR2 (N13114, N13108, N593);
not NOT1 (N13115, N13112);
xor XOR2 (N13116, N13100, N1442);
or OR3 (N13117, N13116, N10323, N11567);
buf BUF1 (N13118, N13115);
buf BUF1 (N13119, N13098);
nand NAND3 (N13120, N13119, N5899, N7938);
or OR2 (N13121, N13113, N10978);
and AND3 (N13122, N13118, N9494, N8576);
nor NOR3 (N13123, N13114, N13033, N762);
not NOT1 (N13124, N13117);
xor XOR2 (N13125, N13096, N4778);
and AND2 (N13126, N13104, N4667);
nor NOR4 (N13127, N13124, N6417, N9947, N704);
not NOT1 (N13128, N13121);
nand NAND3 (N13129, N13122, N5882, N7447);
nor NOR3 (N13130, N13102, N6293, N9822);
and AND4 (N13131, N13128, N10963, N1791, N2220);
buf BUF1 (N13132, N13125);
nor NOR4 (N13133, N13131, N3643, N1247, N5908);
nand NAND2 (N13134, N13123, N5789);
xor XOR2 (N13135, N13126, N7217);
nand NAND4 (N13136, N13135, N4526, N12931, N12990);
nor NOR4 (N13137, N13089, N7565, N9473, N11420);
buf BUF1 (N13138, N13127);
xor XOR2 (N13139, N13138, N2403);
or OR4 (N13140, N13120, N9697, N2132, N7255);
nor NOR2 (N13141, N13140, N8152);
nor NOR3 (N13142, N13134, N7344, N2840);
and AND3 (N13143, N13136, N3096, N3931);
nor NOR2 (N13144, N13137, N5399);
not NOT1 (N13145, N13130);
nor NOR3 (N13146, N13145, N6258, N9662);
xor XOR2 (N13147, N13142, N7953);
xor XOR2 (N13148, N13144, N12813);
not NOT1 (N13149, N13139);
or OR3 (N13150, N13147, N7790, N2488);
nor NOR2 (N13151, N13141, N389);
or OR3 (N13152, N13129, N6032, N294);
nor NOR2 (N13153, N13148, N12995);
nand NAND2 (N13154, N13110, N10473);
not NOT1 (N13155, N13143);
or OR3 (N13156, N13149, N13029, N7657);
not NOT1 (N13157, N13153);
or OR2 (N13158, N13152, N11607);
and AND4 (N13159, N13156, N8425, N12898, N5355);
not NOT1 (N13160, N13150);
not NOT1 (N13161, N13160);
nor NOR3 (N13162, N13161, N10996, N7933);
not NOT1 (N13163, N13146);
and AND4 (N13164, N13157, N8953, N12722, N10698);
nand NAND2 (N13165, N13151, N6662);
and AND2 (N13166, N13132, N9066);
not NOT1 (N13167, N13159);
not NOT1 (N13168, N13133);
not NOT1 (N13169, N13166);
and AND2 (N13170, N13165, N11206);
nand NAND2 (N13171, N13168, N11694);
not NOT1 (N13172, N13154);
not NOT1 (N13173, N13155);
nor NOR3 (N13174, N13172, N11290, N9601);
not NOT1 (N13175, N13163);
not NOT1 (N13176, N13170);
or OR2 (N13177, N13162, N11493);
xor XOR2 (N13178, N13164, N12951);
or OR2 (N13179, N13169, N592);
nand NAND4 (N13180, N13175, N384, N4556, N1639);
xor XOR2 (N13181, N13176, N6940);
nor NOR2 (N13182, N13167, N9407);
not NOT1 (N13183, N13182);
nand NAND2 (N13184, N13181, N9431);
buf BUF1 (N13185, N13177);
nand NAND2 (N13186, N13178, N11453);
buf BUF1 (N13187, N13158);
nand NAND2 (N13188, N13174, N5722);
xor XOR2 (N13189, N13171, N1467);
nor NOR2 (N13190, N13187, N11336);
nand NAND3 (N13191, N13188, N5043, N620);
nand NAND2 (N13192, N13180, N2959);
nor NOR3 (N13193, N13189, N2539, N4642);
not NOT1 (N13194, N13193);
not NOT1 (N13195, N13179);
nand NAND3 (N13196, N13192, N8421, N1686);
nor NOR2 (N13197, N13185, N11914);
nand NAND2 (N13198, N13194, N12502);
and AND2 (N13199, N13198, N11252);
not NOT1 (N13200, N13186);
and AND3 (N13201, N13199, N9769, N6109);
nor NOR2 (N13202, N13195, N11731);
nand NAND4 (N13203, N13202, N12413, N10532, N5841);
nor NOR3 (N13204, N13203, N11710, N5756);
xor XOR2 (N13205, N13201, N5473);
nor NOR2 (N13206, N13205, N5239);
and AND4 (N13207, N13184, N1550, N476, N12123);
buf BUF1 (N13208, N13206);
nand NAND3 (N13209, N13208, N8405, N10139);
and AND3 (N13210, N13173, N5893, N444);
nand NAND2 (N13211, N13200, N7068);
nand NAND4 (N13212, N13190, N365, N5735, N2617);
xor XOR2 (N13213, N13196, N2966);
nor NOR3 (N13214, N13211, N512, N3619);
xor XOR2 (N13215, N13210, N12961);
nor NOR4 (N13216, N13207, N6191, N1219, N10214);
xor XOR2 (N13217, N13215, N8753);
and AND2 (N13218, N13183, N10391);
xor XOR2 (N13219, N13213, N2636);
xor XOR2 (N13220, N13209, N401);
not NOT1 (N13221, N13212);
and AND4 (N13222, N13217, N1578, N1297, N6484);
nor NOR2 (N13223, N13214, N6970);
and AND2 (N13224, N13218, N2122);
not NOT1 (N13225, N13204);
buf BUF1 (N13226, N13222);
not NOT1 (N13227, N13226);
not NOT1 (N13228, N13224);
and AND4 (N13229, N13191, N579, N12784, N9264);
and AND2 (N13230, N13220, N11233);
not NOT1 (N13231, N13227);
nor NOR4 (N13232, N13230, N4585, N815, N12138);
or OR2 (N13233, N13219, N258);
buf BUF1 (N13234, N13233);
buf BUF1 (N13235, N13234);
or OR3 (N13236, N13231, N4264, N6785);
not NOT1 (N13237, N13236);
xor XOR2 (N13238, N13216, N6936);
nand NAND4 (N13239, N13232, N6185, N10585, N3586);
xor XOR2 (N13240, N13237, N3793);
and AND3 (N13241, N13235, N3781, N3741);
and AND2 (N13242, N13229, N11033);
xor XOR2 (N13243, N13241, N12880);
not NOT1 (N13244, N13239);
and AND4 (N13245, N13244, N8291, N1476, N1700);
nor NOR4 (N13246, N13242, N6455, N4195, N1095);
nand NAND2 (N13247, N13246, N2644);
buf BUF1 (N13248, N13228);
buf BUF1 (N13249, N13247);
nor NOR2 (N13250, N13221, N47);
buf BUF1 (N13251, N13197);
buf BUF1 (N13252, N13251);
nor NOR4 (N13253, N13250, N11673, N10467, N1522);
and AND3 (N13254, N13243, N2657, N51);
xor XOR2 (N13255, N13253, N2074);
and AND4 (N13256, N13252, N4843, N10959, N6880);
nand NAND2 (N13257, N13254, N5551);
or OR2 (N13258, N13256, N3690);
nor NOR4 (N13259, N13258, N7682, N11506, N7152);
and AND4 (N13260, N13223, N1039, N434, N10154);
nor NOR2 (N13261, N13259, N9478);
nand NAND2 (N13262, N13260, N9197);
not NOT1 (N13263, N13261);
xor XOR2 (N13264, N13248, N1331);
nand NAND2 (N13265, N13257, N8836);
xor XOR2 (N13266, N13238, N2741);
xor XOR2 (N13267, N13249, N13234);
nand NAND4 (N13268, N13265, N4842, N9745, N6568);
xor XOR2 (N13269, N13264, N2181);
and AND3 (N13270, N13269, N2002, N8258);
not NOT1 (N13271, N13245);
buf BUF1 (N13272, N13255);
not NOT1 (N13273, N13271);
nand NAND2 (N13274, N13267, N10947);
xor XOR2 (N13275, N13272, N6249);
nand NAND3 (N13276, N13240, N8382, N150);
buf BUF1 (N13277, N13274);
or OR2 (N13278, N13276, N11062);
nand NAND3 (N13279, N13277, N286, N981);
nand NAND4 (N13280, N13266, N7055, N7340, N3616);
xor XOR2 (N13281, N13268, N4185);
xor XOR2 (N13282, N13225, N3279);
nor NOR4 (N13283, N13270, N9983, N11580, N8138);
not NOT1 (N13284, N13283);
xor XOR2 (N13285, N13279, N1543);
buf BUF1 (N13286, N13281);
xor XOR2 (N13287, N13262, N8949);
not NOT1 (N13288, N13282);
buf BUF1 (N13289, N13285);
nor NOR4 (N13290, N13286, N2199, N2303, N5171);
or OR2 (N13291, N13284, N2347);
nor NOR2 (N13292, N13280, N2384);
xor XOR2 (N13293, N13278, N557);
and AND4 (N13294, N13287, N9519, N948, N6873);
xor XOR2 (N13295, N13291, N1590);
and AND3 (N13296, N13263, N1151, N11063);
nor NOR3 (N13297, N13275, N2099, N5225);
buf BUF1 (N13298, N13296);
not NOT1 (N13299, N13298);
and AND2 (N13300, N13293, N4562);
nor NOR3 (N13301, N13299, N7356, N2642);
buf BUF1 (N13302, N13297);
and AND3 (N13303, N13302, N12146, N3632);
nor NOR3 (N13304, N13292, N9184, N1150);
not NOT1 (N13305, N13289);
buf BUF1 (N13306, N13301);
nor NOR2 (N13307, N13288, N12405);
buf BUF1 (N13308, N13306);
xor XOR2 (N13309, N13300, N13094);
not NOT1 (N13310, N13294);
not NOT1 (N13311, N13290);
or OR4 (N13312, N13304, N3049, N4644, N10809);
and AND3 (N13313, N13309, N8489, N9871);
xor XOR2 (N13314, N13295, N319);
nand NAND4 (N13315, N13303, N1312, N4283, N11766);
nand NAND3 (N13316, N13315, N7483, N12009);
buf BUF1 (N13317, N13312);
and AND4 (N13318, N13317, N6319, N3918, N7218);
nor NOR3 (N13319, N13316, N6966, N12640);
xor XOR2 (N13320, N13311, N6584);
buf BUF1 (N13321, N13318);
xor XOR2 (N13322, N13305, N10227);
xor XOR2 (N13323, N13320, N6462);
nand NAND3 (N13324, N13321, N4152, N8590);
buf BUF1 (N13325, N13323);
nand NAND4 (N13326, N13324, N4319, N1578, N11588);
or OR2 (N13327, N13313, N12570);
not NOT1 (N13328, N13319);
nand NAND4 (N13329, N13307, N1486, N5863, N12352);
buf BUF1 (N13330, N13329);
nand NAND4 (N13331, N13308, N3720, N13057, N4772);
nand NAND2 (N13332, N13327, N12800);
nand NAND3 (N13333, N13326, N10530, N10531);
and AND2 (N13334, N13273, N6269);
and AND2 (N13335, N13325, N1409);
or OR3 (N13336, N13332, N3215, N11603);
and AND4 (N13337, N13331, N266, N6275, N10185);
or OR4 (N13338, N13328, N12070, N12890, N4163);
buf BUF1 (N13339, N13322);
xor XOR2 (N13340, N13335, N7907);
or OR3 (N13341, N13333, N7614, N6122);
and AND3 (N13342, N13341, N6142, N1862);
buf BUF1 (N13343, N13330);
and AND2 (N13344, N13310, N969);
xor XOR2 (N13345, N13336, N5006);
buf BUF1 (N13346, N13334);
buf BUF1 (N13347, N13314);
not NOT1 (N13348, N13339);
buf BUF1 (N13349, N13346);
not NOT1 (N13350, N13349);
nand NAND2 (N13351, N13342, N10920);
and AND4 (N13352, N13338, N3749, N5348, N12603);
nand NAND3 (N13353, N13343, N1899, N6142);
buf BUF1 (N13354, N13344);
not NOT1 (N13355, N13352);
buf BUF1 (N13356, N13350);
or OR2 (N13357, N13345, N1769);
and AND4 (N13358, N13340, N1527, N6971, N11624);
and AND2 (N13359, N13351, N5638);
xor XOR2 (N13360, N13353, N13304);
and AND3 (N13361, N13348, N2842, N4379);
not NOT1 (N13362, N13357);
nor NOR2 (N13363, N13361, N3811);
nand NAND2 (N13364, N13356, N4719);
buf BUF1 (N13365, N13337);
or OR3 (N13366, N13347, N5855, N12145);
buf BUF1 (N13367, N13355);
nor NOR3 (N13368, N13364, N10191, N6316);
nor NOR2 (N13369, N13363, N12286);
not NOT1 (N13370, N13368);
nand NAND4 (N13371, N13370, N720, N9113, N242);
xor XOR2 (N13372, N13362, N9836);
and AND4 (N13373, N13354, N9225, N1954, N647);
and AND2 (N13374, N13358, N5819);
and AND4 (N13375, N13367, N12696, N11160, N5430);
nand NAND4 (N13376, N13360, N12851, N5474, N6558);
not NOT1 (N13377, N13373);
buf BUF1 (N13378, N13369);
xor XOR2 (N13379, N13374, N12221);
buf BUF1 (N13380, N13372);
and AND3 (N13381, N13377, N10641, N778);
buf BUF1 (N13382, N13375);
and AND2 (N13383, N13365, N9578);
nor NOR2 (N13384, N13380, N12904);
and AND4 (N13385, N13378, N9392, N2799, N284);
and AND4 (N13386, N13384, N9465, N9137, N4198);
buf BUF1 (N13387, N13383);
nor NOR4 (N13388, N13387, N2107, N10369, N5921);
xor XOR2 (N13389, N13376, N13016);
nand NAND2 (N13390, N13371, N513);
nand NAND2 (N13391, N13390, N11655);
or OR3 (N13392, N13366, N611, N4323);
xor XOR2 (N13393, N13388, N1674);
nor NOR4 (N13394, N13386, N12629, N147, N10058);
xor XOR2 (N13395, N13379, N9154);
and AND3 (N13396, N13392, N11798, N2657);
or OR2 (N13397, N13385, N10793);
buf BUF1 (N13398, N13359);
buf BUF1 (N13399, N13397);
and AND4 (N13400, N13394, N11764, N3430, N4640);
xor XOR2 (N13401, N13395, N9493);
nand NAND3 (N13402, N13398, N5607, N3783);
not NOT1 (N13403, N13401);
nand NAND4 (N13404, N13391, N8532, N584, N9542);
not NOT1 (N13405, N13403);
not NOT1 (N13406, N13404);
not NOT1 (N13407, N13399);
and AND2 (N13408, N13402, N9960);
not NOT1 (N13409, N13407);
and AND4 (N13410, N13393, N1515, N10161, N13060);
or OR2 (N13411, N13382, N8353);
buf BUF1 (N13412, N13405);
xor XOR2 (N13413, N13400, N6613);
nand NAND2 (N13414, N13408, N7209);
and AND2 (N13415, N13409, N460);
nand NAND4 (N13416, N13414, N721, N11301, N9658);
xor XOR2 (N13417, N13406, N367);
buf BUF1 (N13418, N13410);
and AND4 (N13419, N13413, N2513, N5737, N1918);
not NOT1 (N13420, N13389);
nor NOR3 (N13421, N13419, N13100, N6966);
xor XOR2 (N13422, N13411, N10869);
or OR3 (N13423, N13412, N8874, N12658);
nor NOR3 (N13424, N13396, N13260, N7672);
nor NOR2 (N13425, N13381, N7588);
xor XOR2 (N13426, N13418, N3118);
or OR2 (N13427, N13425, N5074);
and AND2 (N13428, N13422, N12160);
nor NOR3 (N13429, N13416, N5455, N339);
nand NAND2 (N13430, N13415, N9297);
buf BUF1 (N13431, N13417);
nand NAND3 (N13432, N13430, N11901, N9528);
nor NOR3 (N13433, N13426, N2467, N8923);
and AND3 (N13434, N13431, N11386, N665);
and AND4 (N13435, N13423, N1283, N5058, N7134);
xor XOR2 (N13436, N13432, N8246);
not NOT1 (N13437, N13421);
not NOT1 (N13438, N13434);
not NOT1 (N13439, N13435);
or OR4 (N13440, N13436, N2043, N4591, N12712);
buf BUF1 (N13441, N13429);
or OR4 (N13442, N13440, N9909, N11678, N9700);
xor XOR2 (N13443, N13437, N7178);
nand NAND3 (N13444, N13428, N12179, N10551);
nand NAND3 (N13445, N13433, N6892, N273);
and AND3 (N13446, N13441, N4144, N13311);
and AND3 (N13447, N13442, N209, N1910);
nand NAND3 (N13448, N13446, N5195, N1010);
nand NAND3 (N13449, N13445, N1044, N8173);
and AND3 (N13450, N13444, N9503, N10474);
nor NOR3 (N13451, N13450, N6414, N8743);
and AND4 (N13452, N13449, N11393, N6822, N5731);
not NOT1 (N13453, N13452);
nand NAND3 (N13454, N13443, N12459, N2261);
xor XOR2 (N13455, N13454, N3587);
buf BUF1 (N13456, N13453);
xor XOR2 (N13457, N13438, N5140);
buf BUF1 (N13458, N13451);
xor XOR2 (N13459, N13456, N6634);
nor NOR2 (N13460, N13427, N8556);
xor XOR2 (N13461, N13420, N5730);
nor NOR4 (N13462, N13459, N9991, N11215, N11422);
nor NOR4 (N13463, N13460, N6561, N2429, N13093);
not NOT1 (N13464, N13462);
nand NAND3 (N13465, N13424, N10566, N2311);
xor XOR2 (N13466, N13465, N1210);
buf BUF1 (N13467, N13466);
nor NOR2 (N13468, N13439, N10895);
xor XOR2 (N13469, N13458, N3893);
or OR3 (N13470, N13468, N12504, N1097);
nor NOR4 (N13471, N13467, N2598, N7940, N12205);
xor XOR2 (N13472, N13448, N4964);
not NOT1 (N13473, N13457);
xor XOR2 (N13474, N13464, N13420);
nand NAND4 (N13475, N13471, N6351, N10307, N1011);
xor XOR2 (N13476, N13470, N1540);
and AND2 (N13477, N13455, N276);
and AND2 (N13478, N13474, N880);
nor NOR2 (N13479, N13472, N10086);
xor XOR2 (N13480, N13473, N10271);
and AND2 (N13481, N13475, N13443);
or OR4 (N13482, N13463, N4940, N8414, N2394);
nand NAND2 (N13483, N13481, N2211);
nand NAND4 (N13484, N13479, N7857, N6570, N6422);
or OR3 (N13485, N13482, N11543, N11020);
buf BUF1 (N13486, N13461);
nand NAND3 (N13487, N13486, N10394, N11314);
or OR3 (N13488, N13483, N2475, N6232);
nor NOR3 (N13489, N13469, N6882, N2528);
nor NOR4 (N13490, N13478, N8584, N2442, N1813);
nand NAND4 (N13491, N13476, N13230, N2042, N3240);
nor NOR2 (N13492, N13487, N6953);
xor XOR2 (N13493, N13484, N5886);
nand NAND2 (N13494, N13489, N1311);
and AND2 (N13495, N13447, N10258);
or OR4 (N13496, N13488, N8256, N3788, N11779);
and AND2 (N13497, N13493, N5024);
and AND2 (N13498, N13477, N1631);
nor NOR2 (N13499, N13494, N3830);
buf BUF1 (N13500, N13496);
or OR3 (N13501, N13490, N7182, N2918);
or OR2 (N13502, N13491, N9205);
buf BUF1 (N13503, N13495);
buf BUF1 (N13504, N13480);
and AND2 (N13505, N13502, N2758);
buf BUF1 (N13506, N13503);
xor XOR2 (N13507, N13500, N11459);
nor NOR3 (N13508, N13499, N11233, N12465);
or OR4 (N13509, N13492, N7942, N1767, N12803);
buf BUF1 (N13510, N13501);
buf BUF1 (N13511, N13507);
nand NAND3 (N13512, N13497, N10091, N13071);
or OR3 (N13513, N13511, N6090, N5418);
nand NAND4 (N13514, N13504, N3924, N4806, N6207);
and AND2 (N13515, N13508, N9081);
and AND4 (N13516, N13515, N1735, N8086, N6435);
xor XOR2 (N13517, N13485, N8474);
nand NAND2 (N13518, N13506, N3308);
xor XOR2 (N13519, N13510, N9364);
buf BUF1 (N13520, N13516);
or OR3 (N13521, N13512, N7288, N1063);
not NOT1 (N13522, N13505);
not NOT1 (N13523, N13521);
nand NAND4 (N13524, N13498, N6133, N1645, N8327);
and AND2 (N13525, N13524, N4755);
nand NAND3 (N13526, N13513, N1110, N10310);
not NOT1 (N13527, N13514);
and AND4 (N13528, N13523, N6505, N5320, N1470);
nor NOR2 (N13529, N13522, N6598);
buf BUF1 (N13530, N13528);
and AND2 (N13531, N13517, N10633);
or OR3 (N13532, N13525, N10275, N4014);
buf BUF1 (N13533, N13526);
xor XOR2 (N13534, N13529, N4234);
nand NAND2 (N13535, N13533, N13027);
not NOT1 (N13536, N13518);
or OR2 (N13537, N13509, N8198);
nor NOR3 (N13538, N13520, N3425, N2745);
or OR2 (N13539, N13537, N9144);
and AND3 (N13540, N13536, N7451, N3945);
or OR2 (N13541, N13530, N4037);
or OR2 (N13542, N13527, N10568);
or OR2 (N13543, N13532, N1697);
nor NOR4 (N13544, N13540, N3978, N8940, N5050);
nand NAND2 (N13545, N13542, N9946);
nand NAND4 (N13546, N13531, N7746, N2182, N3876);
and AND2 (N13547, N13539, N880);
and AND4 (N13548, N13519, N11838, N13094, N7759);
not NOT1 (N13549, N13541);
and AND3 (N13550, N13535, N8948, N13453);
not NOT1 (N13551, N13548);
or OR4 (N13552, N13547, N5212, N148, N13008);
nand NAND2 (N13553, N13534, N7014);
not NOT1 (N13554, N13550);
xor XOR2 (N13555, N13546, N10282);
not NOT1 (N13556, N13555);
xor XOR2 (N13557, N13553, N4008);
and AND3 (N13558, N13544, N12256, N2198);
xor XOR2 (N13559, N13538, N9226);
buf BUF1 (N13560, N13543);
nand NAND4 (N13561, N13558, N9765, N1987, N11489);
buf BUF1 (N13562, N13557);
and AND3 (N13563, N13549, N12805, N10453);
nor NOR2 (N13564, N13563, N872);
nor NOR2 (N13565, N13556, N2374);
buf BUF1 (N13566, N13562);
and AND4 (N13567, N13554, N9233, N4664, N10666);
or OR3 (N13568, N13552, N9557, N4403);
buf BUF1 (N13569, N13551);
or OR3 (N13570, N13567, N3913, N3082);
nor NOR3 (N13571, N13569, N10540, N12223);
xor XOR2 (N13572, N13545, N6571);
nand NAND4 (N13573, N13571, N8345, N7974, N4467);
buf BUF1 (N13574, N13570);
or OR3 (N13575, N13560, N5117, N1014);
xor XOR2 (N13576, N13566, N5736);
nand NAND2 (N13577, N13565, N4044);
buf BUF1 (N13578, N13572);
or OR3 (N13579, N13568, N7534, N1723);
xor XOR2 (N13580, N13559, N1824);
nand NAND4 (N13581, N13573, N278, N5761, N1121);
or OR2 (N13582, N13564, N11603);
xor XOR2 (N13583, N13581, N11547);
nor NOR2 (N13584, N13582, N2582);
nand NAND3 (N13585, N13576, N10591, N10947);
or OR4 (N13586, N13574, N4430, N6895, N172);
xor XOR2 (N13587, N13585, N5968);
xor XOR2 (N13588, N13580, N4380);
nand NAND4 (N13589, N13584, N6675, N10373, N2322);
xor XOR2 (N13590, N13578, N6763);
nand NAND3 (N13591, N13589, N5419, N8691);
nand NAND4 (N13592, N13590, N8055, N2379, N8268);
nor NOR3 (N13593, N13575, N8052, N2157);
xor XOR2 (N13594, N13586, N11289);
and AND3 (N13595, N13593, N9818, N13046);
nand NAND2 (N13596, N13592, N1613);
not NOT1 (N13597, N13579);
nor NOR2 (N13598, N13583, N11796);
or OR2 (N13599, N13594, N10287);
nand NAND4 (N13600, N13596, N11100, N7127, N7269);
and AND2 (N13601, N13598, N11179);
buf BUF1 (N13602, N13601);
or OR3 (N13603, N13577, N11244, N3769);
buf BUF1 (N13604, N13591);
and AND2 (N13605, N13588, N9081);
nor NOR3 (N13606, N13604, N8056, N6683);
or OR4 (N13607, N13600, N11128, N1389, N5481);
and AND4 (N13608, N13606, N13380, N5978, N5654);
buf BUF1 (N13609, N13605);
buf BUF1 (N13610, N13561);
not NOT1 (N13611, N13609);
xor XOR2 (N13612, N13608, N970);
not NOT1 (N13613, N13612);
nand NAND3 (N13614, N13587, N10223, N7834);
buf BUF1 (N13615, N13614);
or OR4 (N13616, N13611, N6860, N9668, N12450);
and AND4 (N13617, N13603, N10453, N9916, N10390);
buf BUF1 (N13618, N13613);
not NOT1 (N13619, N13595);
buf BUF1 (N13620, N13597);
buf BUF1 (N13621, N13607);
nor NOR3 (N13622, N13618, N12274, N5446);
nor NOR4 (N13623, N13615, N10525, N4952, N9380);
nand NAND3 (N13624, N13619, N7610, N2974);
or OR3 (N13625, N13623, N7193, N5220);
xor XOR2 (N13626, N13622, N6993);
nor NOR2 (N13627, N13610, N6142);
and AND4 (N13628, N13620, N11629, N7557, N10673);
not NOT1 (N13629, N13617);
xor XOR2 (N13630, N13626, N11631);
and AND4 (N13631, N13625, N7743, N9950, N5279);
nor NOR3 (N13632, N13621, N3643, N4142);
nand NAND3 (N13633, N13602, N183, N11694);
not NOT1 (N13634, N13627);
or OR4 (N13635, N13633, N8127, N2526, N3188);
or OR4 (N13636, N13616, N3299, N4333, N2526);
not NOT1 (N13637, N13599);
xor XOR2 (N13638, N13635, N12693);
and AND2 (N13639, N13634, N8602);
and AND2 (N13640, N13629, N2270);
buf BUF1 (N13641, N13638);
buf BUF1 (N13642, N13624);
nand NAND3 (N13643, N13628, N4556, N4164);
and AND4 (N13644, N13641, N2427, N3083, N3234);
buf BUF1 (N13645, N13636);
or OR3 (N13646, N13632, N9016, N13318);
xor XOR2 (N13647, N13637, N5136);
and AND3 (N13648, N13644, N7110, N7323);
and AND2 (N13649, N13630, N8420);
nand NAND2 (N13650, N13645, N6732);
nor NOR3 (N13651, N13643, N4718, N1380);
nor NOR3 (N13652, N13631, N2460, N7580);
nand NAND3 (N13653, N13646, N8304, N9423);
not NOT1 (N13654, N13648);
xor XOR2 (N13655, N13654, N8966);
nand NAND4 (N13656, N13639, N1065, N7001, N8967);
nor NOR2 (N13657, N13640, N10373);
nand NAND2 (N13658, N13656, N12926);
nand NAND3 (N13659, N13655, N10494, N13468);
xor XOR2 (N13660, N13653, N4645);
or OR2 (N13661, N13660, N11103);
buf BUF1 (N13662, N13658);
nand NAND4 (N13663, N13662, N11421, N1276, N11730);
or OR4 (N13664, N13659, N650, N10388, N2693);
and AND3 (N13665, N13652, N517, N4966);
or OR4 (N13666, N13663, N3725, N6180, N8934);
and AND3 (N13667, N13666, N11077, N21);
xor XOR2 (N13668, N13657, N9462);
not NOT1 (N13669, N13668);
buf BUF1 (N13670, N13661);
or OR3 (N13671, N13669, N12454, N13040);
buf BUF1 (N13672, N13665);
or OR2 (N13673, N13664, N12374);
nand NAND4 (N13674, N13672, N2675, N7817, N1162);
buf BUF1 (N13675, N13674);
and AND2 (N13676, N13651, N9787);
not NOT1 (N13677, N13675);
and AND3 (N13678, N13667, N9641, N2259);
or OR3 (N13679, N13647, N3856, N923);
xor XOR2 (N13680, N13677, N6123);
or OR2 (N13681, N13670, N6486);
nand NAND4 (N13682, N13676, N6403, N10519, N13615);
not NOT1 (N13683, N13671);
or OR2 (N13684, N13649, N799);
or OR3 (N13685, N13642, N7674, N261);
or OR2 (N13686, N13685, N6063);
buf BUF1 (N13687, N13678);
xor XOR2 (N13688, N13686, N11390);
nor NOR3 (N13689, N13650, N10816, N2078);
buf BUF1 (N13690, N13679);
xor XOR2 (N13691, N13680, N13654);
buf BUF1 (N13692, N13691);
nand NAND3 (N13693, N13681, N9662, N2307);
and AND2 (N13694, N13684, N6155);
xor XOR2 (N13695, N13688, N549);
xor XOR2 (N13696, N13687, N2427);
or OR3 (N13697, N13689, N3214, N7503);
nand NAND2 (N13698, N13690, N666);
nor NOR2 (N13699, N13692, N13142);
not NOT1 (N13700, N13698);
and AND4 (N13701, N13697, N9857, N1235, N5209);
or OR3 (N13702, N13699, N6067, N11907);
nor NOR3 (N13703, N13696, N4348, N3436);
buf BUF1 (N13704, N13703);
nand NAND2 (N13705, N13704, N10982);
xor XOR2 (N13706, N13695, N13639);
nand NAND4 (N13707, N13705, N3983, N3279, N3729);
not NOT1 (N13708, N13702);
buf BUF1 (N13709, N13694);
buf BUF1 (N13710, N13707);
nor NOR4 (N13711, N13701, N9035, N11194, N12657);
nor NOR3 (N13712, N13693, N9385, N8059);
and AND2 (N13713, N13682, N11605);
xor XOR2 (N13714, N13712, N4193);
or OR3 (N13715, N13673, N4062, N7089);
nor NOR2 (N13716, N13711, N12599);
nor NOR4 (N13717, N13716, N4596, N1368, N6467);
xor XOR2 (N13718, N13706, N6122);
and AND4 (N13719, N13714, N5504, N1614, N10703);
not NOT1 (N13720, N13709);
not NOT1 (N13721, N13708);
nor NOR4 (N13722, N13700, N8143, N11059, N9138);
not NOT1 (N13723, N13715);
not NOT1 (N13724, N13718);
xor XOR2 (N13725, N13713, N3023);
and AND2 (N13726, N13717, N3218);
buf BUF1 (N13727, N13721);
and AND3 (N13728, N13683, N8409, N12132);
buf BUF1 (N13729, N13719);
or OR2 (N13730, N13720, N2161);
nor NOR4 (N13731, N13710, N5329, N1252, N9991);
and AND4 (N13732, N13727, N1020, N11153, N1265);
not NOT1 (N13733, N13722);
not NOT1 (N13734, N13730);
xor XOR2 (N13735, N13723, N2298);
nor NOR2 (N13736, N13726, N4690);
and AND3 (N13737, N13728, N12680, N2435);
buf BUF1 (N13738, N13724);
nor NOR4 (N13739, N13737, N12626, N3975, N2837);
nor NOR4 (N13740, N13733, N12220, N10333, N12828);
and AND3 (N13741, N13738, N10432, N8816);
xor XOR2 (N13742, N13731, N11129);
xor XOR2 (N13743, N13725, N12096);
xor XOR2 (N13744, N13734, N10258);
not NOT1 (N13745, N13735);
or OR4 (N13746, N13744, N3269, N8113, N3166);
buf BUF1 (N13747, N13732);
not NOT1 (N13748, N13729);
nand NAND4 (N13749, N13736, N3845, N3591, N3306);
xor XOR2 (N13750, N13739, N13316);
buf BUF1 (N13751, N13750);
nor NOR2 (N13752, N13748, N3848);
and AND3 (N13753, N13747, N10948, N3564);
or OR3 (N13754, N13751, N8752, N2508);
or OR2 (N13755, N13754, N3868);
nand NAND4 (N13756, N13749, N2513, N8507, N10413);
and AND3 (N13757, N13756, N10880, N11891);
not NOT1 (N13758, N13755);
nor NOR4 (N13759, N13741, N5214, N9567, N10056);
not NOT1 (N13760, N13745);
xor XOR2 (N13761, N13753, N5481);
nand NAND3 (N13762, N13761, N7835, N12250);
and AND4 (N13763, N13758, N6886, N13647, N7557);
and AND3 (N13764, N13762, N12494, N6864);
or OR4 (N13765, N13746, N13066, N10895, N11426);
xor XOR2 (N13766, N13764, N5707);
and AND2 (N13767, N13740, N12838);
buf BUF1 (N13768, N13767);
nand NAND3 (N13769, N13742, N2070, N5332);
buf BUF1 (N13770, N13759);
nor NOR3 (N13771, N13765, N8883, N7492);
not NOT1 (N13772, N13770);
xor XOR2 (N13773, N13763, N13220);
xor XOR2 (N13774, N13771, N4025);
not NOT1 (N13775, N13769);
buf BUF1 (N13776, N13766);
nand NAND4 (N13777, N13743, N12918, N13760, N12193);
or OR4 (N13778, N1074, N1602, N10231, N819);
buf BUF1 (N13779, N13752);
nor NOR3 (N13780, N13777, N10323, N4605);
nand NAND3 (N13781, N13778, N12535, N13158);
or OR4 (N13782, N13775, N10822, N12483, N11295);
buf BUF1 (N13783, N13768);
xor XOR2 (N13784, N13773, N13665);
and AND2 (N13785, N13782, N6101);
xor XOR2 (N13786, N13784, N12161);
nor NOR2 (N13787, N13783, N2675);
buf BUF1 (N13788, N13776);
nand NAND4 (N13789, N13781, N8331, N5752, N5309);
nand NAND4 (N13790, N13780, N3311, N10005, N2928);
nor NOR4 (N13791, N13789, N870, N462, N2758);
and AND3 (N13792, N13791, N9003, N149);
xor XOR2 (N13793, N13786, N11171);
and AND3 (N13794, N13793, N12486, N13321);
buf BUF1 (N13795, N13787);
and AND3 (N13796, N13792, N1142, N5056);
nand NAND2 (N13797, N13757, N10058);
or OR4 (N13798, N13772, N6014, N816, N989);
and AND2 (N13799, N13788, N1879);
not NOT1 (N13800, N13779);
and AND2 (N13801, N13798, N10051);
or OR2 (N13802, N13785, N9185);
not NOT1 (N13803, N13802);
or OR4 (N13804, N13790, N813, N10445, N12666);
xor XOR2 (N13805, N13803, N13321);
xor XOR2 (N13806, N13796, N7671);
and AND3 (N13807, N13805, N13203, N11720);
nand NAND2 (N13808, N13804, N6767);
or OR4 (N13809, N13801, N5637, N4200, N1390);
nand NAND2 (N13810, N13808, N1591);
nand NAND2 (N13811, N13795, N6532);
and AND4 (N13812, N13810, N12613, N4246, N9365);
xor XOR2 (N13813, N13811, N5077);
not NOT1 (N13814, N13809);
or OR2 (N13815, N13774, N2574);
nand NAND2 (N13816, N13806, N5667);
or OR4 (N13817, N13814, N12868, N7609, N4157);
not NOT1 (N13818, N13815);
buf BUF1 (N13819, N13807);
buf BUF1 (N13820, N13799);
nand NAND3 (N13821, N13812, N13635, N5839);
not NOT1 (N13822, N13820);
xor XOR2 (N13823, N13797, N4058);
and AND4 (N13824, N13818, N7384, N6873, N5629);
or OR2 (N13825, N13821, N4170);
or OR2 (N13826, N13823, N5624);
nor NOR3 (N13827, N13824, N5573, N3909);
buf BUF1 (N13828, N13825);
not NOT1 (N13829, N13819);
nor NOR3 (N13830, N13813, N3845, N2671);
nor NOR4 (N13831, N13826, N3730, N4220, N12561);
buf BUF1 (N13832, N13794);
and AND2 (N13833, N13800, N1928);
not NOT1 (N13834, N13816);
or OR2 (N13835, N13831, N11082);
xor XOR2 (N13836, N13817, N3610);
not NOT1 (N13837, N13822);
xor XOR2 (N13838, N13836, N2179);
xor XOR2 (N13839, N13829, N4168);
nor NOR2 (N13840, N13834, N2011);
xor XOR2 (N13841, N13828, N6313);
or OR2 (N13842, N13827, N13821);
or OR4 (N13843, N13838, N4148, N4264, N9748);
and AND2 (N13844, N13837, N9647);
xor XOR2 (N13845, N13843, N10762);
or OR4 (N13846, N13830, N8313, N9114, N13207);
and AND4 (N13847, N13833, N5296, N669, N9401);
and AND4 (N13848, N13845, N2176, N11038, N9429);
xor XOR2 (N13849, N13844, N189);
and AND3 (N13850, N13847, N3454, N3887);
and AND4 (N13851, N13835, N1358, N5514, N13449);
nand NAND4 (N13852, N13839, N6324, N8381, N9607);
not NOT1 (N13853, N13832);
nand NAND4 (N13854, N13851, N10371, N3409, N13278);
buf BUF1 (N13855, N13842);
xor XOR2 (N13856, N13852, N9455);
or OR3 (N13857, N13841, N6733, N2416);
nand NAND2 (N13858, N13856, N8365);
xor XOR2 (N13859, N13855, N10360);
buf BUF1 (N13860, N13850);
buf BUF1 (N13861, N13859);
or OR4 (N13862, N13848, N13464, N5982, N978);
and AND2 (N13863, N13861, N3454);
or OR3 (N13864, N13858, N13319, N4860);
nand NAND4 (N13865, N13849, N6528, N8699, N7635);
xor XOR2 (N13866, N13865, N8343);
nor NOR2 (N13867, N13857, N5559);
nor NOR2 (N13868, N13863, N11245);
xor XOR2 (N13869, N13868, N7787);
or OR3 (N13870, N13860, N3433, N3009);
buf BUF1 (N13871, N13867);
and AND4 (N13872, N13864, N11629, N4296, N696);
nand NAND4 (N13873, N13840, N12555, N1048, N10466);
not NOT1 (N13874, N13870);
nand NAND3 (N13875, N13873, N12311, N3080);
xor XOR2 (N13876, N13866, N6133);
buf BUF1 (N13877, N13846);
not NOT1 (N13878, N13854);
buf BUF1 (N13879, N13872);
buf BUF1 (N13880, N13853);
nand NAND2 (N13881, N13874, N9638);
or OR3 (N13882, N13876, N6258, N6128);
nand NAND2 (N13883, N13875, N1197);
xor XOR2 (N13884, N13882, N6496);
nor NOR4 (N13885, N13878, N9629, N2401, N4318);
or OR3 (N13886, N13877, N5075, N6487);
buf BUF1 (N13887, N13885);
nor NOR3 (N13888, N13879, N5424, N7973);
xor XOR2 (N13889, N13886, N10132);
nand NAND2 (N13890, N13869, N12441);
xor XOR2 (N13891, N13890, N10736);
buf BUF1 (N13892, N13881);
xor XOR2 (N13893, N13871, N4435);
not NOT1 (N13894, N13883);
and AND2 (N13895, N13880, N10142);
and AND2 (N13896, N13895, N4297);
and AND2 (N13897, N13887, N8782);
or OR2 (N13898, N13893, N12470);
xor XOR2 (N13899, N13894, N11);
nor NOR3 (N13900, N13896, N12174, N3652);
nor NOR3 (N13901, N13891, N11245, N13365);
not NOT1 (N13902, N13889);
nor NOR4 (N13903, N13897, N10604, N4182, N10539);
or OR4 (N13904, N13902, N10288, N4523, N12333);
or OR2 (N13905, N13899, N8971);
and AND3 (N13906, N13892, N3909, N10378);
buf BUF1 (N13907, N13906);
nand NAND2 (N13908, N13901, N3251);
nand NAND4 (N13909, N13908, N6465, N12645, N4918);
buf BUF1 (N13910, N13903);
and AND2 (N13911, N13900, N3255);
or OR4 (N13912, N13898, N3457, N11379, N2446);
and AND2 (N13913, N13862, N5773);
and AND2 (N13914, N13909, N6706);
xor XOR2 (N13915, N13912, N12148);
or OR3 (N13916, N13911, N2942, N7032);
nor NOR2 (N13917, N13888, N5570);
nand NAND4 (N13918, N13907, N12761, N12504, N7825);
xor XOR2 (N13919, N13884, N12942);
not NOT1 (N13920, N13910);
xor XOR2 (N13921, N13918, N871);
or OR4 (N13922, N13915, N10261, N4316, N8631);
or OR2 (N13923, N13916, N6157);
nand NAND2 (N13924, N13905, N2453);
nor NOR3 (N13925, N13919, N7007, N9926);
not NOT1 (N13926, N13921);
xor XOR2 (N13927, N13925, N5751);
and AND3 (N13928, N13924, N9630, N13786);
or OR2 (N13929, N13914, N9780);
xor XOR2 (N13930, N13926, N246);
nand NAND4 (N13931, N13917, N8985, N784, N6704);
nor NOR3 (N13932, N13930, N3445, N9158);
not NOT1 (N13933, N13927);
xor XOR2 (N13934, N13904, N13757);
xor XOR2 (N13935, N13928, N2642);
nand NAND3 (N13936, N13913, N5925, N13872);
nor NOR4 (N13937, N13932, N12823, N1903, N11599);
and AND3 (N13938, N13934, N12487, N3463);
and AND4 (N13939, N13931, N2966, N13158, N3055);
buf BUF1 (N13940, N13923);
nor NOR4 (N13941, N13933, N9106, N7671, N4482);
xor XOR2 (N13942, N13941, N13421);
buf BUF1 (N13943, N13936);
and AND4 (N13944, N13920, N7186, N12592, N2767);
nand NAND3 (N13945, N13943, N11748, N9267);
buf BUF1 (N13946, N13945);
xor XOR2 (N13947, N13937, N10506);
xor XOR2 (N13948, N13946, N5491);
or OR3 (N13949, N13939, N2058, N6042);
or OR3 (N13950, N13922, N3853, N194);
or OR4 (N13951, N13949, N4239, N9800, N5250);
not NOT1 (N13952, N13947);
and AND3 (N13953, N13952, N3053, N7829);
nor NOR2 (N13954, N13942, N2377);
nor NOR4 (N13955, N13935, N6061, N5528, N10267);
nand NAND3 (N13956, N13944, N2564, N3264);
nor NOR3 (N13957, N13948, N6537, N6209);
nor NOR4 (N13958, N13929, N12948, N1746, N13801);
or OR4 (N13959, N13953, N4353, N12440, N652);
nand NAND4 (N13960, N13955, N5042, N3246, N4156);
nand NAND3 (N13961, N13957, N11403, N3847);
buf BUF1 (N13962, N13950);
not NOT1 (N13963, N13960);
buf BUF1 (N13964, N13938);
xor XOR2 (N13965, N13964, N5889);
and AND4 (N13966, N13961, N5980, N3250, N3105);
buf BUF1 (N13967, N13940);
xor XOR2 (N13968, N13962, N7284);
buf BUF1 (N13969, N13954);
not NOT1 (N13970, N13967);
buf BUF1 (N13971, N13958);
nor NOR4 (N13972, N13963, N3151, N1501, N10303);
not NOT1 (N13973, N13966);
buf BUF1 (N13974, N13968);
nand NAND4 (N13975, N13974, N11073, N3430, N3925);
and AND4 (N13976, N13956, N13457, N5801, N74);
and AND4 (N13977, N13975, N10738, N9057, N10640);
or OR2 (N13978, N13971, N223);
or OR4 (N13979, N13972, N9333, N5214, N10165);
xor XOR2 (N13980, N13976, N2955);
nor NOR2 (N13981, N13980, N4515);
nor NOR2 (N13982, N13977, N1375);
and AND3 (N13983, N13965, N4106, N12038);
nor NOR2 (N13984, N13978, N1594);
nand NAND2 (N13985, N13969, N11757);
buf BUF1 (N13986, N13983);
not NOT1 (N13987, N13973);
and AND3 (N13988, N13951, N1669, N4712);
or OR2 (N13989, N13959, N6349);
and AND3 (N13990, N13987, N8977, N13588);
or OR3 (N13991, N13990, N8524, N9427);
nor NOR2 (N13992, N13991, N12412);
nand NAND4 (N13993, N13985, N6476, N5366, N3321);
not NOT1 (N13994, N13988);
not NOT1 (N13995, N13992);
xor XOR2 (N13996, N13982, N9311);
nand NAND4 (N13997, N13994, N2415, N6734, N4230);
nand NAND2 (N13998, N13981, N4458);
and AND3 (N13999, N13995, N5673, N2733);
nor NOR2 (N14000, N13979, N5126);
xor XOR2 (N14001, N13989, N13769);
and AND4 (N14002, N13986, N8415, N13062, N5897);
nand NAND4 (N14003, N14000, N7199, N10109, N429);
not NOT1 (N14004, N13993);
xor XOR2 (N14005, N14004, N9833);
buf BUF1 (N14006, N14002);
not NOT1 (N14007, N13999);
not NOT1 (N14008, N14005);
and AND4 (N14009, N14006, N5771, N4926, N7068);
not NOT1 (N14010, N13970);
or OR3 (N14011, N13984, N6789, N6051);
nor NOR4 (N14012, N14001, N6140, N4867, N10346);
xor XOR2 (N14013, N14008, N1955);
not NOT1 (N14014, N14007);
nor NOR4 (N14015, N13997, N1507, N13846, N12728);
nor NOR4 (N14016, N14011, N1256, N2441, N12971);
and AND4 (N14017, N13996, N5675, N10981, N8049);
or OR3 (N14018, N14012, N5100, N2037);
and AND2 (N14019, N14016, N12644);
not NOT1 (N14020, N14019);
nand NAND4 (N14021, N14010, N12279, N6899, N1607);
buf BUF1 (N14022, N14013);
buf BUF1 (N14023, N14020);
nand NAND3 (N14024, N14021, N6277, N9874);
xor XOR2 (N14025, N14023, N2449);
buf BUF1 (N14026, N14018);
or OR3 (N14027, N14003, N2506, N660);
and AND4 (N14028, N14027, N11074, N6194, N9719);
or OR2 (N14029, N13998, N3350);
and AND2 (N14030, N14022, N10059);
nor NOR4 (N14031, N14014, N829, N6000, N10363);
nor NOR2 (N14032, N14031, N1302);
nor NOR2 (N14033, N14032, N10570);
nand NAND2 (N14034, N14033, N5450);
buf BUF1 (N14035, N14015);
xor XOR2 (N14036, N14035, N7966);
nor NOR4 (N14037, N14029, N10774, N5149, N1591);
xor XOR2 (N14038, N14024, N13704);
nand NAND4 (N14039, N14030, N1408, N4857, N11771);
nor NOR3 (N14040, N14026, N12781, N6859);
xor XOR2 (N14041, N14040, N12922);
not NOT1 (N14042, N14037);
nand NAND2 (N14043, N14034, N2312);
and AND3 (N14044, N14009, N12340, N4896);
xor XOR2 (N14045, N14043, N11169);
xor XOR2 (N14046, N14045, N9226);
buf BUF1 (N14047, N14039);
nor NOR2 (N14048, N14025, N13667);
and AND4 (N14049, N14047, N10010, N13621, N728);
nand NAND2 (N14050, N14046, N12512);
buf BUF1 (N14051, N14036);
and AND2 (N14052, N14049, N4934);
and AND3 (N14053, N14028, N11546, N1814);
not NOT1 (N14054, N14042);
not NOT1 (N14055, N14041);
buf BUF1 (N14056, N14052);
xor XOR2 (N14057, N14038, N1610);
and AND2 (N14058, N14054, N8211);
buf BUF1 (N14059, N14057);
nand NAND3 (N14060, N14056, N3039, N3968);
not NOT1 (N14061, N14055);
or OR3 (N14062, N14053, N13146, N9159);
not NOT1 (N14063, N14060);
buf BUF1 (N14064, N14061);
nand NAND4 (N14065, N14048, N6816, N12715, N114);
nand NAND4 (N14066, N14058, N8983, N838, N1119);
not NOT1 (N14067, N14044);
not NOT1 (N14068, N14051);
nand NAND2 (N14069, N14063, N3028);
not NOT1 (N14070, N14065);
and AND3 (N14071, N14062, N10122, N9695);
buf BUF1 (N14072, N14017);
or OR3 (N14073, N14071, N11878, N10125);
not NOT1 (N14074, N14070);
nor NOR3 (N14075, N14073, N11142, N6187);
nand NAND2 (N14076, N14066, N9076);
xor XOR2 (N14077, N14074, N7423);
xor XOR2 (N14078, N14077, N11083);
xor XOR2 (N14079, N14069, N8529);
nor NOR2 (N14080, N14068, N6247);
buf BUF1 (N14081, N14050);
nand NAND4 (N14082, N14059, N2705, N9736, N6943);
nor NOR4 (N14083, N14078, N1924, N5178, N5900);
and AND2 (N14084, N14067, N11850);
and AND3 (N14085, N14064, N9950, N5884);
xor XOR2 (N14086, N14083, N8302);
nor NOR3 (N14087, N14085, N9924, N10251);
and AND3 (N14088, N14086, N11175, N12809);
nor NOR3 (N14089, N14082, N10298, N8201);
nor NOR3 (N14090, N14076, N12837, N7898);
buf BUF1 (N14091, N14088);
xor XOR2 (N14092, N14079, N11005);
buf BUF1 (N14093, N14081);
nand NAND4 (N14094, N14080, N7568, N3716, N12561);
nor NOR2 (N14095, N14087, N7272);
or OR3 (N14096, N14084, N6186, N3851);
not NOT1 (N14097, N14096);
xor XOR2 (N14098, N14090, N4625);
nand NAND3 (N14099, N14092, N6627, N3944);
not NOT1 (N14100, N14072);
or OR3 (N14101, N14075, N11788, N12852);
not NOT1 (N14102, N14097);
nand NAND4 (N14103, N14098, N8052, N13364, N3051);
not NOT1 (N14104, N14095);
or OR4 (N14105, N14089, N2310, N2932, N7319);
nor NOR2 (N14106, N14093, N13075);
xor XOR2 (N14107, N14101, N5523);
xor XOR2 (N14108, N14103, N3453);
xor XOR2 (N14109, N14106, N12087);
and AND3 (N14110, N14099, N11166, N9942);
not NOT1 (N14111, N14107);
not NOT1 (N14112, N14105);
not NOT1 (N14113, N14112);
xor XOR2 (N14114, N14102, N13893);
xor XOR2 (N14115, N14094, N10061);
xor XOR2 (N14116, N14115, N9540);
not NOT1 (N14117, N14114);
not NOT1 (N14118, N14091);
buf BUF1 (N14119, N14104);
xor XOR2 (N14120, N14119, N649);
nor NOR2 (N14121, N14110, N11734);
and AND4 (N14122, N14117, N12692, N4222, N5672);
and AND2 (N14123, N14111, N8698);
buf BUF1 (N14124, N14113);
nand NAND2 (N14125, N14123, N12161);
buf BUF1 (N14126, N14108);
buf BUF1 (N14127, N14126);
nor NOR2 (N14128, N14116, N2913);
xor XOR2 (N14129, N14120, N11572);
buf BUF1 (N14130, N14128);
not NOT1 (N14131, N14118);
nand NAND2 (N14132, N14124, N11598);
nand NAND2 (N14133, N14131, N7421);
xor XOR2 (N14134, N14109, N13923);
nor NOR2 (N14135, N14129, N7187);
or OR3 (N14136, N14133, N4505, N2823);
buf BUF1 (N14137, N14134);
and AND4 (N14138, N14130, N2235, N2251, N747);
buf BUF1 (N14139, N14127);
nor NOR2 (N14140, N14139, N4642);
buf BUF1 (N14141, N14138);
nand NAND4 (N14142, N14122, N11124, N10814, N5161);
not NOT1 (N14143, N14141);
nor NOR2 (N14144, N14135, N7583);
and AND4 (N14145, N14142, N7081, N12970, N5080);
buf BUF1 (N14146, N14136);
not NOT1 (N14147, N14143);
nand NAND3 (N14148, N14121, N4669, N53);
nand NAND4 (N14149, N14132, N2820, N11425, N8969);
not NOT1 (N14150, N14149);
buf BUF1 (N14151, N14137);
not NOT1 (N14152, N14144);
or OR3 (N14153, N14125, N10981, N11202);
nor NOR4 (N14154, N14140, N7851, N2027, N3447);
xor XOR2 (N14155, N14147, N6887);
not NOT1 (N14156, N14153);
not NOT1 (N14157, N14146);
or OR3 (N14158, N14100, N8412, N11613);
buf BUF1 (N14159, N14158);
and AND2 (N14160, N14151, N357);
xor XOR2 (N14161, N14157, N9198);
and AND2 (N14162, N14152, N8580);
buf BUF1 (N14163, N14159);
buf BUF1 (N14164, N14161);
nand NAND4 (N14165, N14145, N13517, N5055, N2030);
buf BUF1 (N14166, N14154);
buf BUF1 (N14167, N14163);
buf BUF1 (N14168, N14148);
nand NAND4 (N14169, N14166, N2770, N12716, N12720);
or OR3 (N14170, N14162, N12053, N7920);
xor XOR2 (N14171, N14155, N7575);
and AND4 (N14172, N14167, N10155, N9979, N11055);
xor XOR2 (N14173, N14165, N1438);
buf BUF1 (N14174, N14164);
nand NAND3 (N14175, N14168, N13863, N8048);
buf BUF1 (N14176, N14160);
xor XOR2 (N14177, N14175, N8556);
not NOT1 (N14178, N14173);
not NOT1 (N14179, N14169);
not NOT1 (N14180, N14172);
buf BUF1 (N14181, N14171);
or OR2 (N14182, N14170, N2179);
nor NOR2 (N14183, N14180, N12507);
xor XOR2 (N14184, N14183, N3798);
buf BUF1 (N14185, N14179);
not NOT1 (N14186, N14182);
nor NOR4 (N14187, N14174, N6231, N3511, N2148);
buf BUF1 (N14188, N14185);
or OR2 (N14189, N14150, N2767);
and AND2 (N14190, N14188, N2215);
and AND3 (N14191, N14178, N9375, N6858);
buf BUF1 (N14192, N14176);
nand NAND3 (N14193, N14184, N5214, N9156);
buf BUF1 (N14194, N14189);
buf BUF1 (N14195, N14193);
buf BUF1 (N14196, N14195);
or OR3 (N14197, N14156, N6745, N8365);
not NOT1 (N14198, N14196);
xor XOR2 (N14199, N14190, N3154);
xor XOR2 (N14200, N14197, N4230);
nand NAND2 (N14201, N14186, N3409);
nor NOR2 (N14202, N14199, N7387);
or OR3 (N14203, N14201, N1910, N9423);
buf BUF1 (N14204, N14200);
xor XOR2 (N14205, N14191, N6485);
nand NAND4 (N14206, N14203, N4358, N11859, N2087);
nand NAND3 (N14207, N14192, N13740, N13191);
not NOT1 (N14208, N14202);
and AND4 (N14209, N14198, N4167, N11239, N12185);
or OR4 (N14210, N14208, N2604, N12311, N1770);
not NOT1 (N14211, N14194);
nor NOR4 (N14212, N14177, N3984, N6266, N4291);
buf BUF1 (N14213, N14207);
nor NOR3 (N14214, N14206, N11303, N3320);
and AND2 (N14215, N14211, N9845);
or OR4 (N14216, N14205, N10826, N14119, N4262);
xor XOR2 (N14217, N14215, N4989);
or OR2 (N14218, N14209, N5439);
nor NOR2 (N14219, N14216, N9544);
buf BUF1 (N14220, N14212);
nor NOR4 (N14221, N14181, N6880, N2026, N358);
and AND2 (N14222, N14213, N25);
xor XOR2 (N14223, N14210, N7964);
not NOT1 (N14224, N14214);
or OR3 (N14225, N14220, N3146, N1742);
or OR2 (N14226, N14219, N12621);
and AND2 (N14227, N14204, N6197);
buf BUF1 (N14228, N14217);
buf BUF1 (N14229, N14218);
nand NAND2 (N14230, N14222, N2808);
xor XOR2 (N14231, N14226, N502);
xor XOR2 (N14232, N14187, N6207);
and AND2 (N14233, N14232, N3124);
and AND2 (N14234, N14228, N13845);
xor XOR2 (N14235, N14221, N1395);
or OR3 (N14236, N14227, N8435, N7268);
nor NOR4 (N14237, N14223, N4025, N1577, N9648);
and AND4 (N14238, N14225, N9077, N11568, N8595);
nand NAND3 (N14239, N14237, N8407, N11188);
nor NOR2 (N14240, N14238, N11133);
xor XOR2 (N14241, N14234, N7646);
not NOT1 (N14242, N14239);
xor XOR2 (N14243, N14241, N4788);
xor XOR2 (N14244, N14230, N11733);
nor NOR2 (N14245, N14242, N4712);
and AND3 (N14246, N14229, N9119, N13041);
xor XOR2 (N14247, N14236, N3065);
nor NOR4 (N14248, N14245, N13398, N1478, N5893);
xor XOR2 (N14249, N14244, N8063);
buf BUF1 (N14250, N14224);
not NOT1 (N14251, N14248);
or OR2 (N14252, N14240, N11410);
not NOT1 (N14253, N14251);
buf BUF1 (N14254, N14233);
nand NAND3 (N14255, N14250, N10739, N10173);
nand NAND3 (N14256, N14255, N5764, N5221);
or OR2 (N14257, N14252, N14236);
xor XOR2 (N14258, N14249, N7110);
buf BUF1 (N14259, N14257);
nand NAND3 (N14260, N14256, N3470, N9370);
nor NOR2 (N14261, N14258, N5878);
and AND2 (N14262, N14246, N1387);
and AND4 (N14263, N14243, N5352, N9675, N10628);
nor NOR4 (N14264, N14231, N5111, N13964, N9439);
or OR4 (N14265, N14247, N5980, N7513, N2531);
nor NOR3 (N14266, N14253, N4992, N11717);
and AND4 (N14267, N14235, N1878, N4027, N8966);
nor NOR4 (N14268, N14254, N9990, N8730, N6798);
and AND2 (N14269, N14261, N11698);
or OR3 (N14270, N14260, N6802, N2273);
and AND4 (N14271, N14263, N2218, N1915, N2993);
and AND3 (N14272, N14270, N12339, N7321);
nand NAND3 (N14273, N14259, N1007, N12084);
buf BUF1 (N14274, N14267);
nor NOR3 (N14275, N14269, N14220, N3871);
buf BUF1 (N14276, N14262);
and AND3 (N14277, N14272, N143, N7400);
nor NOR3 (N14278, N14274, N10458, N5437);
and AND3 (N14279, N14271, N9396, N299);
nand NAND3 (N14280, N14265, N12805, N8529);
not NOT1 (N14281, N14278);
and AND2 (N14282, N14277, N6974);
nor NOR3 (N14283, N14273, N6262, N8679);
buf BUF1 (N14284, N14276);
nand NAND4 (N14285, N14284, N7777, N12704, N6776);
buf BUF1 (N14286, N14266);
not NOT1 (N14287, N14264);
and AND2 (N14288, N14268, N1117);
xor XOR2 (N14289, N14288, N12324);
xor XOR2 (N14290, N14282, N6354);
xor XOR2 (N14291, N14287, N6023);
xor XOR2 (N14292, N14285, N3415);
nand NAND3 (N14293, N14275, N7579, N234);
or OR2 (N14294, N14289, N11380);
xor XOR2 (N14295, N14291, N9478);
nand NAND2 (N14296, N14286, N10770);
and AND3 (N14297, N14295, N12611, N1186);
nor NOR2 (N14298, N14296, N11994);
buf BUF1 (N14299, N14283);
nand NAND4 (N14300, N14299, N7578, N11516, N9798);
xor XOR2 (N14301, N14300, N8215);
or OR4 (N14302, N14297, N7003, N1033, N13290);
buf BUF1 (N14303, N14298);
and AND3 (N14304, N14279, N4643, N13448);
and AND3 (N14305, N14294, N12880, N1631);
or OR3 (N14306, N14302, N11265, N6242);
or OR2 (N14307, N14292, N3694);
xor XOR2 (N14308, N14293, N7285);
not NOT1 (N14309, N14280);
buf BUF1 (N14310, N14290);
nand NAND2 (N14311, N14301, N13243);
and AND4 (N14312, N14311, N7325, N4461, N10544);
and AND2 (N14313, N14306, N4363);
or OR2 (N14314, N14312, N6247);
or OR4 (N14315, N14313, N2178, N10629, N1029);
xor XOR2 (N14316, N14305, N4497);
buf BUF1 (N14317, N14308);
nor NOR4 (N14318, N14309, N11959, N8171, N11027);
xor XOR2 (N14319, N14316, N8179);
not NOT1 (N14320, N14281);
and AND2 (N14321, N14310, N9140);
nand NAND4 (N14322, N14314, N5571, N8205, N1343);
not NOT1 (N14323, N14304);
xor XOR2 (N14324, N14317, N4389);
or OR2 (N14325, N14303, N984);
or OR3 (N14326, N14324, N1931, N3052);
or OR2 (N14327, N14307, N10941);
not NOT1 (N14328, N14325);
not NOT1 (N14329, N14322);
nand NAND4 (N14330, N14315, N7622, N12912, N4388);
not NOT1 (N14331, N14326);
or OR2 (N14332, N14320, N7365);
buf BUF1 (N14333, N14330);
or OR2 (N14334, N14327, N420);
buf BUF1 (N14335, N14323);
not NOT1 (N14336, N14333);
xor XOR2 (N14337, N14318, N1355);
nand NAND3 (N14338, N14337, N6021, N12529);
not NOT1 (N14339, N14332);
or OR2 (N14340, N14321, N10831);
not NOT1 (N14341, N14334);
or OR3 (N14342, N14340, N8910, N2788);
nand NAND2 (N14343, N14342, N8312);
xor XOR2 (N14344, N14336, N11742);
nand NAND4 (N14345, N14338, N5762, N10569, N3726);
nor NOR4 (N14346, N14319, N12534, N7733, N10254);
and AND3 (N14347, N14343, N3635, N2439);
not NOT1 (N14348, N14344);
not NOT1 (N14349, N14341);
nor NOR3 (N14350, N14349, N13286, N8484);
not NOT1 (N14351, N14335);
nand NAND2 (N14352, N14345, N10664);
and AND2 (N14353, N14339, N13738);
xor XOR2 (N14354, N14348, N2610);
not NOT1 (N14355, N14350);
xor XOR2 (N14356, N14331, N13153);
or OR4 (N14357, N14346, N691, N13859, N14349);
buf BUF1 (N14358, N14353);
not NOT1 (N14359, N14329);
xor XOR2 (N14360, N14358, N4855);
buf BUF1 (N14361, N14359);
nor NOR4 (N14362, N14328, N8781, N72, N6075);
or OR3 (N14363, N14360, N2249, N798);
not NOT1 (N14364, N14356);
nor NOR2 (N14365, N14362, N14297);
nand NAND4 (N14366, N14351, N6948, N971, N10133);
or OR4 (N14367, N14355, N9325, N8072, N5195);
xor XOR2 (N14368, N14354, N12720);
nand NAND3 (N14369, N14364, N8646, N2879);
nand NAND2 (N14370, N14365, N13915);
or OR3 (N14371, N14347, N11756, N992);
not NOT1 (N14372, N14368);
nor NOR2 (N14373, N14367, N3336);
xor XOR2 (N14374, N14363, N7999);
nor NOR4 (N14375, N14372, N6203, N9029, N1271);
not NOT1 (N14376, N14361);
buf BUF1 (N14377, N14352);
nor NOR2 (N14378, N14373, N12467);
buf BUF1 (N14379, N14374);
nand NAND3 (N14380, N14366, N7237, N65);
buf BUF1 (N14381, N14380);
or OR4 (N14382, N14376, N9088, N106, N13752);
not NOT1 (N14383, N14378);
buf BUF1 (N14384, N14369);
xor XOR2 (N14385, N14370, N9453);
nor NOR2 (N14386, N14381, N10667);
xor XOR2 (N14387, N14377, N12368);
xor XOR2 (N14388, N14385, N2247);
nor NOR2 (N14389, N14383, N94);
and AND4 (N14390, N14375, N2196, N13622, N8346);
not NOT1 (N14391, N14388);
or OR3 (N14392, N14379, N13828, N4637);
not NOT1 (N14393, N14391);
nor NOR2 (N14394, N14357, N11939);
xor XOR2 (N14395, N14382, N4485);
or OR2 (N14396, N14392, N13685);
and AND2 (N14397, N14393, N8454);
xor XOR2 (N14398, N14384, N3728);
xor XOR2 (N14399, N14398, N1439);
not NOT1 (N14400, N14386);
or OR4 (N14401, N14394, N10381, N1680, N5052);
buf BUF1 (N14402, N14371);
xor XOR2 (N14403, N14396, N12336);
nor NOR4 (N14404, N14401, N7166, N5671, N4177);
or OR4 (N14405, N14395, N8503, N11807, N1039);
buf BUF1 (N14406, N14402);
and AND3 (N14407, N14400, N13858, N5458);
nand NAND3 (N14408, N14407, N7165, N10212);
xor XOR2 (N14409, N14397, N14112);
and AND2 (N14410, N14399, N6730);
xor XOR2 (N14411, N14406, N10975);
nand NAND2 (N14412, N14408, N6982);
nand NAND3 (N14413, N14412, N7115, N2646);
nor NOR4 (N14414, N14404, N3699, N8491, N6954);
xor XOR2 (N14415, N14405, N6709);
nand NAND3 (N14416, N14410, N6530, N7900);
nand NAND2 (N14417, N14414, N9969);
nor NOR4 (N14418, N14389, N8725, N6742, N10528);
or OR2 (N14419, N14409, N6986);
not NOT1 (N14420, N14419);
nand NAND2 (N14421, N14413, N11804);
not NOT1 (N14422, N14416);
not NOT1 (N14423, N14422);
nand NAND3 (N14424, N14417, N6767, N11232);
nor NOR3 (N14425, N14415, N13781, N12717);
nor NOR3 (N14426, N14387, N12787, N9977);
buf BUF1 (N14427, N14403);
or OR2 (N14428, N14390, N1667);
and AND3 (N14429, N14420, N7050, N4698);
not NOT1 (N14430, N14411);
buf BUF1 (N14431, N14418);
buf BUF1 (N14432, N14427);
and AND3 (N14433, N14429, N11094, N3979);
nor NOR4 (N14434, N14421, N12144, N13025, N7826);
nor NOR3 (N14435, N14423, N6505, N8769);
not NOT1 (N14436, N14428);
not NOT1 (N14437, N14431);
nor NOR4 (N14438, N14426, N3428, N9526, N882);
xor XOR2 (N14439, N14432, N4835);
not NOT1 (N14440, N14424);
nand NAND2 (N14441, N14434, N5021);
nand NAND2 (N14442, N14435, N3323);
buf BUF1 (N14443, N14440);
and AND2 (N14444, N14430, N1278);
buf BUF1 (N14445, N14425);
or OR2 (N14446, N14438, N3034);
and AND2 (N14447, N14445, N2635);
buf BUF1 (N14448, N14443);
not NOT1 (N14449, N14433);
not NOT1 (N14450, N14448);
or OR3 (N14451, N14449, N652, N9968);
or OR2 (N14452, N14442, N2853);
and AND2 (N14453, N14450, N7778);
nand NAND3 (N14454, N14441, N7525, N13485);
xor XOR2 (N14455, N14439, N694);
nor NOR4 (N14456, N14437, N5767, N3066, N7068);
or OR3 (N14457, N14451, N13426, N14350);
buf BUF1 (N14458, N14444);
nand NAND4 (N14459, N14458, N12361, N12007, N7364);
xor XOR2 (N14460, N14436, N2732);
not NOT1 (N14461, N14459);
buf BUF1 (N14462, N14453);
nand NAND4 (N14463, N14460, N6811, N6671, N13088);
not NOT1 (N14464, N14461);
or OR3 (N14465, N14447, N3468, N4061);
not NOT1 (N14466, N14462);
xor XOR2 (N14467, N14452, N73);
xor XOR2 (N14468, N14466, N13281);
or OR3 (N14469, N14454, N5263, N2052);
nor NOR4 (N14470, N14456, N13506, N10512, N7527);
nor NOR2 (N14471, N14468, N11043);
or OR2 (N14472, N14463, N13289);
not NOT1 (N14473, N14465);
buf BUF1 (N14474, N14455);
or OR2 (N14475, N14473, N12325);
buf BUF1 (N14476, N14469);
not NOT1 (N14477, N14467);
nand NAND2 (N14478, N14471, N11459);
buf BUF1 (N14479, N14477);
nor NOR2 (N14480, N14470, N2056);
and AND2 (N14481, N14476, N10020);
xor XOR2 (N14482, N14481, N1355);
not NOT1 (N14483, N14475);
nor NOR2 (N14484, N14479, N10550);
and AND4 (N14485, N14478, N13727, N8496, N9698);
nor NOR4 (N14486, N14485, N5902, N12157, N8762);
nor NOR3 (N14487, N14472, N4738, N3296);
buf BUF1 (N14488, N14484);
nor NOR3 (N14489, N14486, N1744, N6577);
nor NOR3 (N14490, N14457, N5344, N8486);
buf BUF1 (N14491, N14488);
nor NOR3 (N14492, N14489, N7829, N818);
buf BUF1 (N14493, N14464);
nor NOR4 (N14494, N14493, N10055, N10285, N13216);
and AND2 (N14495, N14480, N9417);
xor XOR2 (N14496, N14483, N1818);
not NOT1 (N14497, N14487);
and AND2 (N14498, N14495, N12555);
not NOT1 (N14499, N14496);
nor NOR3 (N14500, N14494, N813, N7112);
nor NOR3 (N14501, N14490, N10325, N280);
buf BUF1 (N14502, N14498);
buf BUF1 (N14503, N14502);
xor XOR2 (N14504, N14482, N11399);
or OR3 (N14505, N14492, N375, N657);
nor NOR3 (N14506, N14446, N11091, N8629);
and AND4 (N14507, N14491, N4680, N495, N6789);
nand NAND2 (N14508, N14501, N13102);
nor NOR4 (N14509, N14497, N8844, N11760, N12470);
xor XOR2 (N14510, N14507, N11558);
nand NAND2 (N14511, N14508, N14306);
or OR2 (N14512, N14510, N9149);
and AND2 (N14513, N14505, N9738);
nand NAND2 (N14514, N14500, N10149);
not NOT1 (N14515, N14511);
nor NOR4 (N14516, N14514, N342, N5912, N6130);
and AND4 (N14517, N14474, N8678, N14331, N14183);
and AND3 (N14518, N14504, N6184, N12696);
and AND4 (N14519, N14517, N10107, N12516, N831);
not NOT1 (N14520, N14512);
nor NOR2 (N14521, N14518, N11876);
buf BUF1 (N14522, N14509);
or OR4 (N14523, N14503, N10100, N9559, N1162);
not NOT1 (N14524, N14513);
and AND4 (N14525, N14522, N10135, N130, N2673);
nand NAND2 (N14526, N14516, N3720);
not NOT1 (N14527, N14515);
xor XOR2 (N14528, N14506, N8465);
not NOT1 (N14529, N14523);
and AND3 (N14530, N14519, N9775, N7877);
not NOT1 (N14531, N14526);
and AND4 (N14532, N14499, N2832, N6135, N96);
nor NOR4 (N14533, N14520, N7010, N13071, N12281);
nand NAND4 (N14534, N14530, N10345, N11978, N9083);
nor NOR3 (N14535, N14529, N12340, N9795);
nor NOR4 (N14536, N14525, N7340, N12599, N13503);
nor NOR3 (N14537, N14527, N14260, N12867);
not NOT1 (N14538, N14524);
xor XOR2 (N14539, N14532, N7148);
not NOT1 (N14540, N14521);
not NOT1 (N14541, N14535);
buf BUF1 (N14542, N14534);
nor NOR3 (N14543, N14541, N11716, N1221);
nor NOR4 (N14544, N14536, N1373, N10050, N2406);
buf BUF1 (N14545, N14540);
not NOT1 (N14546, N14544);
not NOT1 (N14547, N14531);
buf BUF1 (N14548, N14528);
and AND2 (N14549, N14543, N13783);
xor XOR2 (N14550, N14547, N2926);
and AND3 (N14551, N14548, N13243, N5924);
and AND2 (N14552, N14551, N7867);
or OR2 (N14553, N14538, N6762);
buf BUF1 (N14554, N14552);
buf BUF1 (N14555, N14542);
nor NOR4 (N14556, N14550, N5880, N8222, N7501);
and AND4 (N14557, N14553, N603, N5863, N555);
buf BUF1 (N14558, N14545);
nor NOR3 (N14559, N14549, N10984, N14122);
nor NOR3 (N14560, N14558, N10049, N11436);
nor NOR3 (N14561, N14557, N12465, N1419);
nor NOR3 (N14562, N14561, N11291, N6228);
or OR3 (N14563, N14533, N127, N3743);
or OR3 (N14564, N14555, N7352, N10948);
xor XOR2 (N14565, N14537, N9755);
xor XOR2 (N14566, N14564, N6401);
nor NOR3 (N14567, N14565, N12016, N1060);
xor XOR2 (N14568, N14562, N6158);
and AND2 (N14569, N14568, N12652);
nor NOR4 (N14570, N14563, N6722, N3026, N9484);
nand NAND2 (N14571, N14546, N12922);
nand NAND2 (N14572, N14571, N4209);
nand NAND2 (N14573, N14556, N8357);
nand NAND4 (N14574, N14572, N4570, N2345, N11430);
not NOT1 (N14575, N14554);
nand NAND2 (N14576, N14574, N3286);
and AND2 (N14577, N14539, N8815);
and AND2 (N14578, N14569, N12736);
xor XOR2 (N14579, N14566, N6383);
xor XOR2 (N14580, N14567, N96);
or OR4 (N14581, N14570, N3282, N7782, N2267);
nand NAND3 (N14582, N14576, N7482, N9588);
and AND4 (N14583, N14575, N10091, N11973, N10637);
xor XOR2 (N14584, N14583, N980);
nor NOR2 (N14585, N14580, N7023);
nor NOR3 (N14586, N14573, N6489, N7371);
xor XOR2 (N14587, N14578, N11157);
not NOT1 (N14588, N14585);
xor XOR2 (N14589, N14584, N4477);
nor NOR4 (N14590, N14589, N14393, N4621, N5527);
buf BUF1 (N14591, N14590);
or OR4 (N14592, N14559, N7891, N3192, N4750);
or OR2 (N14593, N14579, N1274);
not NOT1 (N14594, N14587);
not NOT1 (N14595, N14586);
xor XOR2 (N14596, N14591, N4983);
and AND2 (N14597, N14592, N12615);
nand NAND3 (N14598, N14582, N833, N5909);
nor NOR2 (N14599, N14581, N13071);
and AND3 (N14600, N14596, N4626, N4328);
nand NAND4 (N14601, N14597, N2205, N9344, N8101);
buf BUF1 (N14602, N14601);
not NOT1 (N14603, N14588);
xor XOR2 (N14604, N14599, N10463);
buf BUF1 (N14605, N14603);
nor NOR3 (N14606, N14600, N8472, N4268);
xor XOR2 (N14607, N14594, N8033);
nand NAND3 (N14608, N14577, N9735, N11954);
nor NOR4 (N14609, N14595, N2100, N1388, N6993);
or OR2 (N14610, N14602, N728);
nand NAND2 (N14611, N14606, N9357);
and AND4 (N14612, N14611, N14090, N283, N6793);
not NOT1 (N14613, N14609);
not NOT1 (N14614, N14608);
and AND2 (N14615, N14605, N292);
nand NAND2 (N14616, N14614, N14290);
xor XOR2 (N14617, N14607, N516);
not NOT1 (N14618, N14610);
buf BUF1 (N14619, N14612);
not NOT1 (N14620, N14615);
not NOT1 (N14621, N14604);
nor NOR2 (N14622, N14617, N3582);
or OR4 (N14623, N14560, N11065, N3549, N11694);
not NOT1 (N14624, N14593);
nand NAND2 (N14625, N14598, N2719);
not NOT1 (N14626, N14620);
and AND4 (N14627, N14625, N7708, N6943, N13530);
nand NAND4 (N14628, N14621, N6210, N594, N11277);
buf BUF1 (N14629, N14616);
xor XOR2 (N14630, N14618, N1172);
or OR4 (N14631, N14622, N4244, N8123, N2284);
and AND3 (N14632, N14629, N6014, N3029);
not NOT1 (N14633, N14632);
nand NAND3 (N14634, N14623, N1503, N7341);
nand NAND3 (N14635, N14634, N8244, N8794);
nand NAND4 (N14636, N14619, N4867, N7016, N12601);
nand NAND3 (N14637, N14613, N11571, N10183);
xor XOR2 (N14638, N14636, N6892);
and AND4 (N14639, N14630, N2862, N4411, N6591);
nand NAND2 (N14640, N14626, N1931);
or OR3 (N14641, N14631, N2013, N8704);
nor NOR2 (N14642, N14638, N3750);
xor XOR2 (N14643, N14633, N3209);
buf BUF1 (N14644, N14627);
not NOT1 (N14645, N14642);
or OR2 (N14646, N14641, N1135);
nand NAND3 (N14647, N14644, N10166, N12085);
and AND3 (N14648, N14637, N12142, N10144);
nand NAND2 (N14649, N14645, N2056);
buf BUF1 (N14650, N14649);
nand NAND4 (N14651, N14647, N7818, N2797, N14561);
nand NAND3 (N14652, N14635, N4959, N10238);
buf BUF1 (N14653, N14643);
buf BUF1 (N14654, N14628);
and AND2 (N14655, N14648, N1203);
buf BUF1 (N14656, N14651);
nor NOR4 (N14657, N14656, N1405, N9952, N5305);
xor XOR2 (N14658, N14654, N727);
buf BUF1 (N14659, N14652);
nand NAND2 (N14660, N14650, N6709);
nand NAND2 (N14661, N14639, N9278);
not NOT1 (N14662, N14660);
buf BUF1 (N14663, N14653);
xor XOR2 (N14664, N14659, N4588);
nor NOR2 (N14665, N14661, N3449);
or OR4 (N14666, N14663, N1272, N12515, N4609);
nor NOR3 (N14667, N14640, N2724, N3381);
not NOT1 (N14668, N14646);
or OR2 (N14669, N14662, N5205);
and AND2 (N14670, N14668, N3811);
buf BUF1 (N14671, N14655);
or OR4 (N14672, N14665, N4215, N13972, N7351);
nor NOR3 (N14673, N14671, N9194, N121);
nor NOR4 (N14674, N14670, N7184, N3025, N13623);
nor NOR2 (N14675, N14669, N10708);
nand NAND3 (N14676, N14667, N428, N5065);
xor XOR2 (N14677, N14673, N4023);
buf BUF1 (N14678, N14677);
and AND2 (N14679, N14672, N6897);
or OR3 (N14680, N14674, N3574, N12651);
and AND3 (N14681, N14678, N6714, N5359);
buf BUF1 (N14682, N14676);
not NOT1 (N14683, N14681);
and AND4 (N14684, N14664, N6158, N2648, N7435);
nand NAND4 (N14685, N14657, N8204, N13619, N9915);
buf BUF1 (N14686, N14683);
xor XOR2 (N14687, N14685, N13093);
nand NAND2 (N14688, N14687, N10347);
or OR4 (N14689, N14680, N1665, N4987, N8079);
nand NAND4 (N14690, N14688, N9543, N9012, N2322);
nor NOR2 (N14691, N14666, N3429);
nor NOR3 (N14692, N14658, N4643, N5513);
and AND4 (N14693, N14682, N6410, N3699, N9426);
or OR3 (N14694, N14686, N7227, N13592);
nor NOR4 (N14695, N14684, N8980, N7811, N14595);
nand NAND4 (N14696, N14690, N7200, N4867, N9395);
not NOT1 (N14697, N14675);
not NOT1 (N14698, N14696);
and AND4 (N14699, N14697, N7450, N3062, N4076);
xor XOR2 (N14700, N14694, N8453);
nand NAND4 (N14701, N14624, N2381, N2224, N13542);
nor NOR4 (N14702, N14693, N11033, N10734, N11267);
buf BUF1 (N14703, N14699);
buf BUF1 (N14704, N14679);
or OR3 (N14705, N14698, N3638, N5121);
not NOT1 (N14706, N14691);
nor NOR2 (N14707, N14702, N8491);
nor NOR3 (N14708, N14703, N13633, N3631);
and AND3 (N14709, N14689, N13513, N6804);
nand NAND2 (N14710, N14701, N9416);
nand NAND4 (N14711, N14700, N7083, N3010, N3000);
buf BUF1 (N14712, N14708);
or OR2 (N14713, N14692, N7609);
nand NAND4 (N14714, N14712, N8409, N13947, N5350);
or OR4 (N14715, N14705, N5649, N10989, N1011);
nand NAND4 (N14716, N14715, N1315, N11156, N14521);
nor NOR4 (N14717, N14707, N14418, N7683, N6113);
and AND3 (N14718, N14713, N4065, N10764);
xor XOR2 (N14719, N14704, N9256);
xor XOR2 (N14720, N14710, N10621);
and AND4 (N14721, N14719, N5564, N1373, N8655);
xor XOR2 (N14722, N14721, N2794);
nor NOR2 (N14723, N14709, N2011);
or OR3 (N14724, N14706, N5187, N4290);
nor NOR2 (N14725, N14720, N1626);
nor NOR4 (N14726, N14695, N3010, N8359, N9805);
not NOT1 (N14727, N14714);
xor XOR2 (N14728, N14723, N3106);
nor NOR3 (N14729, N14711, N12701, N3917);
and AND2 (N14730, N14724, N6105);
and AND3 (N14731, N14716, N7190, N9835);
not NOT1 (N14732, N14718);
and AND2 (N14733, N14731, N11601);
and AND2 (N14734, N14729, N3895);
or OR3 (N14735, N14725, N6507, N7642);
not NOT1 (N14736, N14727);
nand NAND2 (N14737, N14733, N1613);
nand NAND2 (N14738, N14736, N6084);
nor NOR2 (N14739, N14726, N8075);
buf BUF1 (N14740, N14730);
nor NOR4 (N14741, N14734, N4117, N5587, N8546);
nor NOR3 (N14742, N14722, N2896, N11156);
nand NAND3 (N14743, N14742, N14203, N12225);
not NOT1 (N14744, N14728);
not NOT1 (N14745, N14732);
buf BUF1 (N14746, N14743);
buf BUF1 (N14747, N14746);
nand NAND2 (N14748, N14744, N9750);
nand NAND3 (N14749, N14717, N10826, N4907);
nor NOR3 (N14750, N14739, N10399, N7018);
xor XOR2 (N14751, N14737, N8376);
or OR4 (N14752, N14751, N4361, N9121, N10302);
nand NAND4 (N14753, N14747, N7772, N3408, N14239);
xor XOR2 (N14754, N14753, N4426);
not NOT1 (N14755, N14748);
not NOT1 (N14756, N14741);
buf BUF1 (N14757, N14738);
not NOT1 (N14758, N14740);
not NOT1 (N14759, N14755);
and AND3 (N14760, N14754, N13230, N8013);
or OR2 (N14761, N14745, N8710);
not NOT1 (N14762, N14735);
nor NOR3 (N14763, N14749, N12361, N7705);
not NOT1 (N14764, N14762);
not NOT1 (N14765, N14752);
buf BUF1 (N14766, N14765);
nor NOR4 (N14767, N14760, N8914, N3744, N1528);
xor XOR2 (N14768, N14758, N14202);
buf BUF1 (N14769, N14763);
or OR4 (N14770, N14761, N10335, N3741, N13091);
not NOT1 (N14771, N14757);
or OR4 (N14772, N14768, N2946, N12723, N9580);
or OR4 (N14773, N14769, N6689, N7151, N13087);
nor NOR2 (N14774, N14771, N2816);
not NOT1 (N14775, N14759);
not NOT1 (N14776, N14756);
xor XOR2 (N14777, N14770, N13492);
not NOT1 (N14778, N14774);
not NOT1 (N14779, N14776);
nor NOR4 (N14780, N14773, N12790, N12887, N12801);
xor XOR2 (N14781, N14764, N8484);
xor XOR2 (N14782, N14780, N11028);
or OR2 (N14783, N14778, N5547);
nand NAND2 (N14784, N14766, N4044);
nor NOR3 (N14785, N14767, N3693, N2847);
or OR3 (N14786, N14777, N5543, N12349);
not NOT1 (N14787, N14786);
not NOT1 (N14788, N14781);
xor XOR2 (N14789, N14779, N14756);
buf BUF1 (N14790, N14787);
nand NAND2 (N14791, N14782, N14348);
and AND2 (N14792, N14790, N7954);
and AND3 (N14793, N14784, N6293, N12998);
and AND4 (N14794, N14775, N6980, N8634, N3422);
nand NAND3 (N14795, N14792, N4624, N4862);
and AND4 (N14796, N14794, N599, N1406, N4940);
not NOT1 (N14797, N14783);
xor XOR2 (N14798, N14750, N7726);
and AND2 (N14799, N14785, N3286);
and AND4 (N14800, N14796, N7764, N7105, N12721);
nand NAND2 (N14801, N14800, N11574);
or OR4 (N14802, N14795, N4498, N2961, N3257);
and AND2 (N14803, N14789, N6955);
and AND3 (N14804, N14791, N5581, N5878);
buf BUF1 (N14805, N14803);
and AND3 (N14806, N14793, N11385, N13122);
or OR2 (N14807, N14797, N12675);
buf BUF1 (N14808, N14798);
nand NAND2 (N14809, N14802, N639);
buf BUF1 (N14810, N14804);
or OR4 (N14811, N14801, N5001, N3251, N13922);
nand NAND4 (N14812, N14807, N1739, N8639, N1350);
or OR4 (N14813, N14799, N12258, N11043, N4760);
or OR4 (N14814, N14788, N13685, N3963, N4778);
nand NAND4 (N14815, N14805, N11243, N8774, N9447);
and AND2 (N14816, N14815, N5530);
and AND4 (N14817, N14772, N12856, N11903, N14392);
or OR4 (N14818, N14811, N495, N13841, N2615);
buf BUF1 (N14819, N14814);
and AND3 (N14820, N14812, N11313, N5275);
buf BUF1 (N14821, N14808);
not NOT1 (N14822, N14809);
buf BUF1 (N14823, N14821);
nor NOR3 (N14824, N14823, N5596, N11721);
buf BUF1 (N14825, N14824);
nor NOR4 (N14826, N14820, N8996, N12138, N12507);
buf BUF1 (N14827, N14817);
or OR3 (N14828, N14818, N8306, N2535);
not NOT1 (N14829, N14826);
buf BUF1 (N14830, N14828);
and AND3 (N14831, N14830, N1598, N850);
nor NOR2 (N14832, N14819, N10212);
nor NOR2 (N14833, N14810, N1422);
nand NAND3 (N14834, N14833, N806, N3906);
or OR4 (N14835, N14806, N11976, N4056, N4698);
buf BUF1 (N14836, N14834);
xor XOR2 (N14837, N14831, N6144);
xor XOR2 (N14838, N14829, N1799);
not NOT1 (N14839, N14837);
nor NOR3 (N14840, N14836, N5102, N8356);
nor NOR2 (N14841, N14840, N12407);
and AND4 (N14842, N14825, N2056, N11361, N2487);
or OR4 (N14843, N14816, N14367, N11436, N4238);
nand NAND2 (N14844, N14843, N5947);
nor NOR3 (N14845, N14841, N10424, N13958);
buf BUF1 (N14846, N14838);
xor XOR2 (N14847, N14827, N982);
buf BUF1 (N14848, N14835);
buf BUF1 (N14849, N14845);
not NOT1 (N14850, N14822);
and AND3 (N14851, N14849, N4091, N5446);
and AND4 (N14852, N14850, N2309, N8011, N314);
nor NOR2 (N14853, N14848, N837);
nor NOR4 (N14854, N14853, N5017, N9443, N4449);
and AND3 (N14855, N14844, N1836, N12526);
or OR2 (N14856, N14852, N10956);
nand NAND3 (N14857, N14839, N8654, N3583);
buf BUF1 (N14858, N14856);
nor NOR4 (N14859, N14851, N5509, N7860, N8406);
buf BUF1 (N14860, N14842);
or OR4 (N14861, N14832, N13347, N6927, N380);
nand NAND2 (N14862, N14859, N1989);
xor XOR2 (N14863, N14861, N13082);
and AND3 (N14864, N14847, N12551, N5087);
or OR2 (N14865, N14846, N4750);
xor XOR2 (N14866, N14813, N14466);
or OR4 (N14867, N14865, N8064, N8420, N6362);
xor XOR2 (N14868, N14858, N10913);
buf BUF1 (N14869, N14864);
nand NAND4 (N14870, N14857, N1739, N6009, N13911);
and AND4 (N14871, N14855, N9150, N10153, N3220);
or OR3 (N14872, N14863, N12948, N3088);
xor XOR2 (N14873, N14866, N14350);
nand NAND2 (N14874, N14870, N13258);
xor XOR2 (N14875, N14872, N635);
xor XOR2 (N14876, N14862, N6281);
nor NOR3 (N14877, N14876, N9287, N814);
buf BUF1 (N14878, N14874);
or OR3 (N14879, N14878, N3313, N9912);
buf BUF1 (N14880, N14875);
nor NOR2 (N14881, N14860, N13397);
and AND4 (N14882, N14880, N4100, N4953, N5014);
not NOT1 (N14883, N14873);
not NOT1 (N14884, N14867);
buf BUF1 (N14885, N14868);
nor NOR4 (N14886, N14854, N4118, N4482, N2724);
or OR4 (N14887, N14885, N11586, N9141, N7704);
buf BUF1 (N14888, N14884);
xor XOR2 (N14889, N14882, N2602);
or OR4 (N14890, N14881, N7974, N2749, N141);
xor XOR2 (N14891, N14887, N6119);
and AND4 (N14892, N14891, N11018, N6598, N6892);
not NOT1 (N14893, N14869);
and AND2 (N14894, N14879, N9844);
nor NOR2 (N14895, N14889, N13677);
nor NOR4 (N14896, N14890, N5514, N12270, N3582);
xor XOR2 (N14897, N14888, N4242);
not NOT1 (N14898, N14894);
buf BUF1 (N14899, N14898);
nor NOR4 (N14900, N14893, N4937, N6836, N1242);
not NOT1 (N14901, N14895);
and AND2 (N14902, N14897, N12352);
not NOT1 (N14903, N14899);
xor XOR2 (N14904, N14886, N13648);
not NOT1 (N14905, N14892);
buf BUF1 (N14906, N14871);
or OR2 (N14907, N14877, N9499);
nor NOR2 (N14908, N14905, N11423);
or OR2 (N14909, N14883, N5356);
buf BUF1 (N14910, N14902);
nand NAND2 (N14911, N14903, N2672);
not NOT1 (N14912, N14907);
or OR4 (N14913, N14909, N10385, N10451, N14910);
nand NAND3 (N14914, N9247, N9738, N9311);
nand NAND4 (N14915, N14911, N2654, N13199, N2186);
xor XOR2 (N14916, N14896, N2963);
nand NAND2 (N14917, N14900, N8868);
buf BUF1 (N14918, N14914);
not NOT1 (N14919, N14901);
nor NOR3 (N14920, N14918, N6837, N13712);
xor XOR2 (N14921, N14915, N2625);
nor NOR2 (N14922, N14908, N2424);
nand NAND2 (N14923, N14916, N13676);
not NOT1 (N14924, N14923);
or OR2 (N14925, N14906, N986);
and AND4 (N14926, N14912, N2379, N9063, N11090);
not NOT1 (N14927, N14925);
nand NAND2 (N14928, N14924, N11606);
nand NAND2 (N14929, N14917, N9896);
or OR4 (N14930, N14928, N1991, N9756, N11059);
buf BUF1 (N14931, N14922);
buf BUF1 (N14932, N14920);
xor XOR2 (N14933, N14913, N3056);
buf BUF1 (N14934, N14929);
not NOT1 (N14935, N14904);
and AND4 (N14936, N14930, N6689, N1133, N7405);
and AND4 (N14937, N14934, N5825, N3598, N13678);
and AND2 (N14938, N14932, N9357);
or OR4 (N14939, N14936, N11926, N3450, N10407);
not NOT1 (N14940, N14926);
xor XOR2 (N14941, N14940, N13982);
xor XOR2 (N14942, N14931, N3059);
not NOT1 (N14943, N14942);
nor NOR4 (N14944, N14919, N1397, N1375, N3265);
or OR2 (N14945, N14939, N2420);
xor XOR2 (N14946, N14921, N9154);
nor NOR4 (N14947, N14944, N13405, N4200, N11262);
xor XOR2 (N14948, N14933, N14277);
buf BUF1 (N14949, N14947);
buf BUF1 (N14950, N14948);
nor NOR3 (N14951, N14945, N14778, N9024);
nor NOR4 (N14952, N14946, N11956, N12307, N9200);
nor NOR2 (N14953, N14938, N3303);
nor NOR2 (N14954, N14941, N8483);
not NOT1 (N14955, N14950);
buf BUF1 (N14956, N14937);
buf BUF1 (N14957, N14935);
xor XOR2 (N14958, N14949, N10063);
and AND3 (N14959, N14953, N849, N10661);
nand NAND2 (N14960, N14956, N14075);
and AND3 (N14961, N14955, N6927, N12932);
not NOT1 (N14962, N14952);
or OR4 (N14963, N14960, N10455, N5071, N36);
buf BUF1 (N14964, N14961);
nor NOR4 (N14965, N14959, N12523, N2774, N7116);
nand NAND2 (N14966, N14964, N707);
nand NAND2 (N14967, N14965, N9385);
not NOT1 (N14968, N14958);
not NOT1 (N14969, N14954);
nor NOR2 (N14970, N14969, N8398);
xor XOR2 (N14971, N14963, N6401);
or OR2 (N14972, N14970, N3186);
not NOT1 (N14973, N14968);
not NOT1 (N14974, N14951);
or OR3 (N14975, N14957, N9910, N12817);
and AND2 (N14976, N14966, N13177);
nand NAND3 (N14977, N14943, N14137, N6636);
or OR2 (N14978, N14967, N4673);
and AND4 (N14979, N14971, N2972, N6313, N14628);
and AND4 (N14980, N14927, N13901, N9279, N6769);
buf BUF1 (N14981, N14974);
and AND3 (N14982, N14975, N12168, N9859);
nor NOR4 (N14983, N14981, N964, N1422, N550);
xor XOR2 (N14984, N14979, N10352);
not NOT1 (N14985, N14984);
xor XOR2 (N14986, N14973, N14883);
xor XOR2 (N14987, N14983, N8231);
nor NOR3 (N14988, N14986, N1073, N7499);
or OR3 (N14989, N14962, N14178, N10608);
or OR3 (N14990, N14978, N13686, N11222);
nand NAND2 (N14991, N14976, N2297);
xor XOR2 (N14992, N14989, N7583);
nand NAND4 (N14993, N14988, N922, N1220, N5350);
xor XOR2 (N14994, N14972, N7028);
nor NOR2 (N14995, N14993, N682);
nand NAND2 (N14996, N14985, N11178);
xor XOR2 (N14997, N14982, N6685);
and AND4 (N14998, N14980, N3673, N2492, N1909);
xor XOR2 (N14999, N14990, N7154);
xor XOR2 (N15000, N14998, N1312);
or OR2 (N15001, N15000, N13471);
not NOT1 (N15002, N14994);
nand NAND2 (N15003, N14987, N3314);
not NOT1 (N15004, N14992);
buf BUF1 (N15005, N14999);
xor XOR2 (N15006, N15001, N12763);
or OR3 (N15007, N14997, N7527, N6967);
or OR3 (N15008, N15007, N2698, N12854);
nand NAND4 (N15009, N15006, N1726, N12889, N2692);
not NOT1 (N15010, N15009);
xor XOR2 (N15011, N14991, N8045);
nand NAND4 (N15012, N15004, N14046, N11284, N7980);
buf BUF1 (N15013, N15012);
not NOT1 (N15014, N14995);
nor NOR3 (N15015, N15013, N6479, N2054);
xor XOR2 (N15016, N14996, N11572);
and AND4 (N15017, N15015, N8782, N12566, N7741);
nor NOR4 (N15018, N15002, N10881, N14429, N3857);
nand NAND4 (N15019, N15018, N1047, N1286, N8055);
buf BUF1 (N15020, N15019);
xor XOR2 (N15021, N15003, N2167);
or OR3 (N15022, N15017, N2064, N12511);
not NOT1 (N15023, N15008);
or OR4 (N15024, N14977, N7976, N8468, N3923);
buf BUF1 (N15025, N15022);
or OR3 (N15026, N15025, N2275, N12429);
xor XOR2 (N15027, N15021, N12158);
buf BUF1 (N15028, N15016);
or OR3 (N15029, N15011, N1818, N8874);
nand NAND3 (N15030, N15023, N14782, N14492);
not NOT1 (N15031, N15014);
and AND4 (N15032, N15026, N4620, N2313, N1581);
and AND4 (N15033, N15032, N6517, N13962, N9918);
and AND4 (N15034, N15020, N9833, N3988, N14777);
and AND2 (N15035, N15034, N10906);
buf BUF1 (N15036, N15029);
not NOT1 (N15037, N15033);
or OR4 (N15038, N15037, N9727, N14338, N13323);
nor NOR2 (N15039, N15010, N10371);
buf BUF1 (N15040, N15030);
not NOT1 (N15041, N15028);
xor XOR2 (N15042, N15036, N9148);
buf BUF1 (N15043, N15005);
and AND4 (N15044, N15024, N9350, N1871, N13114);
buf BUF1 (N15045, N15043);
nor NOR3 (N15046, N15031, N13513, N6624);
buf BUF1 (N15047, N15044);
nand NAND3 (N15048, N15041, N6171, N5885);
nor NOR2 (N15049, N15046, N8105);
nand NAND3 (N15050, N15027, N9283, N8905);
or OR2 (N15051, N15039, N9058);
nand NAND2 (N15052, N15047, N13957);
buf BUF1 (N15053, N15048);
or OR4 (N15054, N15038, N11871, N6930, N8135);
nor NOR4 (N15055, N15052, N13368, N11528, N6400);
not NOT1 (N15056, N15049);
xor XOR2 (N15057, N15051, N1952);
buf BUF1 (N15058, N15050);
nor NOR4 (N15059, N15055, N6917, N173, N12877);
buf BUF1 (N15060, N15057);
nand NAND4 (N15061, N15042, N1785, N7022, N5078);
xor XOR2 (N15062, N15056, N6803);
buf BUF1 (N15063, N15053);
nand NAND4 (N15064, N15059, N14643, N1837, N14971);
nand NAND3 (N15065, N15062, N8775, N5501);
or OR3 (N15066, N15063, N7198, N7629);
xor XOR2 (N15067, N15035, N957);
buf BUF1 (N15068, N15040);
and AND2 (N15069, N15060, N11149);
and AND3 (N15070, N15054, N310, N9570);
nand NAND2 (N15071, N15061, N11403);
xor XOR2 (N15072, N15071, N5670);
buf BUF1 (N15073, N15067);
nand NAND4 (N15074, N15064, N6473, N3031, N12932);
and AND4 (N15075, N15065, N2853, N10356, N13050);
or OR2 (N15076, N15058, N5228);
nand NAND3 (N15077, N15075, N14345, N5689);
nor NOR4 (N15078, N15069, N3163, N7492, N13210);
not NOT1 (N15079, N15072);
nand NAND4 (N15080, N15074, N5740, N1594, N7040);
buf BUF1 (N15081, N15076);
nand NAND2 (N15082, N15066, N14164);
nor NOR4 (N15083, N15077, N1211, N10125, N3451);
or OR3 (N15084, N15045, N10138, N11363);
xor XOR2 (N15085, N15083, N8217);
or OR4 (N15086, N15084, N12006, N3354, N424);
xor XOR2 (N15087, N15081, N2798);
nor NOR2 (N15088, N15079, N4268);
or OR4 (N15089, N15070, N213, N10825, N5895);
xor XOR2 (N15090, N15089, N14703);
not NOT1 (N15091, N15087);
and AND3 (N15092, N15080, N6546, N1053);
and AND3 (N15093, N15085, N12136, N3375);
buf BUF1 (N15094, N15088);
buf BUF1 (N15095, N15086);
nand NAND3 (N15096, N15095, N6788, N11163);
xor XOR2 (N15097, N15091, N8041);
buf BUF1 (N15098, N15082);
not NOT1 (N15099, N15073);
not NOT1 (N15100, N15090);
nand NAND4 (N15101, N15078, N4370, N10249, N5399);
buf BUF1 (N15102, N15101);
or OR2 (N15103, N15099, N2762);
nand NAND2 (N15104, N15094, N11803);
xor XOR2 (N15105, N15098, N11409);
buf BUF1 (N15106, N15097);
nor NOR4 (N15107, N15106, N10815, N2907, N4138);
or OR4 (N15108, N15068, N9523, N7052, N10778);
xor XOR2 (N15109, N15092, N1921);
not NOT1 (N15110, N15109);
buf BUF1 (N15111, N15105);
or OR2 (N15112, N15110, N8346);
buf BUF1 (N15113, N15100);
buf BUF1 (N15114, N15112);
buf BUF1 (N15115, N15103);
xor XOR2 (N15116, N15114, N14014);
nor NOR4 (N15117, N15113, N10143, N8885, N15003);
xor XOR2 (N15118, N15093, N2353);
or OR4 (N15119, N15102, N11192, N2604, N15054);
nand NAND2 (N15120, N15116, N3415);
xor XOR2 (N15121, N15115, N2962);
nor NOR4 (N15122, N15111, N5119, N14043, N1576);
nand NAND3 (N15123, N15118, N2588, N4014);
nand NAND2 (N15124, N15096, N12769);
nand NAND2 (N15125, N15120, N2067);
buf BUF1 (N15126, N15124);
xor XOR2 (N15127, N15108, N8814);
nand NAND2 (N15128, N15127, N6983);
nand NAND3 (N15129, N15107, N5233, N14955);
and AND3 (N15130, N15121, N13569, N14611);
and AND3 (N15131, N15117, N13447, N10643);
nor NOR2 (N15132, N15125, N3084);
and AND3 (N15133, N15130, N1226, N15008);
buf BUF1 (N15134, N15119);
and AND3 (N15135, N15129, N5590, N10866);
nand NAND3 (N15136, N15135, N12757, N5418);
nor NOR3 (N15137, N15104, N1320, N5773);
buf BUF1 (N15138, N15123);
nand NAND2 (N15139, N15131, N4072);
xor XOR2 (N15140, N15134, N12255);
not NOT1 (N15141, N15138);
or OR4 (N15142, N15132, N5371, N4350, N7372);
nand NAND3 (N15143, N15141, N938, N5444);
or OR4 (N15144, N15136, N6626, N10594, N5401);
nand NAND3 (N15145, N15144, N8666, N14942);
not NOT1 (N15146, N15140);
and AND2 (N15147, N15143, N9117);
xor XOR2 (N15148, N15133, N37);
xor XOR2 (N15149, N15126, N13836);
nor NOR2 (N15150, N15149, N8636);
and AND2 (N15151, N15150, N11465);
not NOT1 (N15152, N15151);
buf BUF1 (N15153, N15146);
nor NOR2 (N15154, N15122, N12673);
and AND4 (N15155, N15139, N13813, N7102, N13296);
nand NAND2 (N15156, N15155, N18);
buf BUF1 (N15157, N15148);
nand NAND3 (N15158, N15128, N12174, N13672);
nor NOR4 (N15159, N15145, N308, N1301, N1541);
and AND3 (N15160, N15142, N11696, N3650);
nand NAND2 (N15161, N15152, N5796);
xor XOR2 (N15162, N15160, N7502);
nand NAND2 (N15163, N15154, N12426);
and AND4 (N15164, N15157, N7373, N13246, N12081);
nor NOR3 (N15165, N15156, N376, N4236);
nor NOR4 (N15166, N15162, N14954, N12670, N1559);
nor NOR2 (N15167, N15153, N2086);
not NOT1 (N15168, N15167);
buf BUF1 (N15169, N15166);
not NOT1 (N15170, N15165);
and AND2 (N15171, N15169, N3603);
nor NOR3 (N15172, N15164, N9874, N12724);
not NOT1 (N15173, N15158);
buf BUF1 (N15174, N15171);
or OR4 (N15175, N15174, N1978, N2593, N4098);
buf BUF1 (N15176, N15172);
or OR3 (N15177, N15168, N7796, N2089);
and AND4 (N15178, N15147, N2162, N8961, N11449);
nand NAND2 (N15179, N15177, N10409);
nand NAND2 (N15180, N15176, N9191);
not NOT1 (N15181, N15161);
buf BUF1 (N15182, N15175);
or OR2 (N15183, N15137, N3920);
nand NAND4 (N15184, N15170, N4333, N10586, N768);
xor XOR2 (N15185, N15182, N9250);
buf BUF1 (N15186, N15180);
buf BUF1 (N15187, N15185);
buf BUF1 (N15188, N15179);
xor XOR2 (N15189, N15184, N8030);
and AND3 (N15190, N15181, N13049, N9608);
or OR4 (N15191, N15183, N12676, N4537, N14118);
nor NOR2 (N15192, N15191, N6492);
nand NAND3 (N15193, N15159, N13017, N10100);
not NOT1 (N15194, N15189);
nor NOR4 (N15195, N15186, N1141, N9728, N7848);
nor NOR4 (N15196, N15187, N10619, N3220, N14784);
nand NAND4 (N15197, N15195, N2149, N6033, N8109);
and AND4 (N15198, N15178, N12763, N6981, N10249);
not NOT1 (N15199, N15196);
nand NAND4 (N15200, N15190, N4396, N2032, N4307);
or OR2 (N15201, N15199, N7278);
or OR3 (N15202, N15201, N1587, N12999);
or OR3 (N15203, N15194, N5337, N6459);
nand NAND3 (N15204, N15173, N13401, N5474);
nor NOR4 (N15205, N15188, N10245, N6045, N9389);
nand NAND4 (N15206, N15203, N3221, N3478, N8175);
nor NOR2 (N15207, N15192, N1205);
or OR4 (N15208, N15193, N2038, N2611, N9274);
xor XOR2 (N15209, N15163, N14190);
nand NAND4 (N15210, N15205, N5561, N11824, N7413);
and AND2 (N15211, N15198, N6289);
not NOT1 (N15212, N15207);
xor XOR2 (N15213, N15208, N5694);
or OR2 (N15214, N15213, N14649);
or OR2 (N15215, N15214, N11579);
and AND4 (N15216, N15211, N10918, N4056, N12724);
nor NOR3 (N15217, N15200, N14712, N10526);
not NOT1 (N15218, N15212);
nand NAND2 (N15219, N15210, N12831);
and AND3 (N15220, N15216, N11694, N7846);
and AND3 (N15221, N15215, N1605, N2734);
buf BUF1 (N15222, N15206);
nor NOR2 (N15223, N15218, N14321);
buf BUF1 (N15224, N15209);
nand NAND2 (N15225, N15222, N13915);
or OR2 (N15226, N15225, N10630);
buf BUF1 (N15227, N15204);
buf BUF1 (N15228, N15221);
nor NOR2 (N15229, N15197, N8892);
or OR3 (N15230, N15224, N929, N12914);
or OR4 (N15231, N15223, N14916, N6566, N14175);
buf BUF1 (N15232, N15202);
xor XOR2 (N15233, N15219, N4579);
nor NOR3 (N15234, N15226, N9889, N5963);
or OR4 (N15235, N15231, N8369, N1332, N894);
nor NOR3 (N15236, N15220, N6101, N5564);
xor XOR2 (N15237, N15236, N1596);
not NOT1 (N15238, N15217);
not NOT1 (N15239, N15228);
buf BUF1 (N15240, N15238);
not NOT1 (N15241, N15239);
or OR3 (N15242, N15233, N3220, N2920);
and AND3 (N15243, N15234, N6978, N10592);
not NOT1 (N15244, N15242);
xor XOR2 (N15245, N15243, N6491);
nor NOR4 (N15246, N15229, N1152, N2147, N56);
and AND3 (N15247, N15240, N13875, N6016);
nor NOR4 (N15248, N15244, N12061, N7233, N2638);
xor XOR2 (N15249, N15235, N1194);
not NOT1 (N15250, N15246);
or OR2 (N15251, N15237, N6144);
nor NOR4 (N15252, N15230, N9719, N4885, N9795);
nor NOR3 (N15253, N15227, N1785, N7902);
nor NOR4 (N15254, N15245, N6345, N11821, N7793);
or OR4 (N15255, N15248, N14665, N9807, N11575);
or OR3 (N15256, N15253, N8338, N9936);
or OR2 (N15257, N15249, N5999);
buf BUF1 (N15258, N15241);
nor NOR2 (N15259, N15257, N11961);
xor XOR2 (N15260, N15250, N7578);
or OR2 (N15261, N15232, N5239);
nor NOR3 (N15262, N15259, N10954, N13402);
buf BUF1 (N15263, N15251);
buf BUF1 (N15264, N15254);
or OR3 (N15265, N15263, N3402, N1012);
nor NOR2 (N15266, N15260, N2235);
buf BUF1 (N15267, N15255);
not NOT1 (N15268, N15252);
or OR2 (N15269, N15247, N7037);
nor NOR2 (N15270, N15268, N9403);
buf BUF1 (N15271, N15261);
or OR3 (N15272, N15266, N5474, N12088);
nor NOR2 (N15273, N15256, N5611);
nor NOR2 (N15274, N15265, N1783);
and AND3 (N15275, N15274, N8606, N15206);
nor NOR2 (N15276, N15272, N14778);
nand NAND3 (N15277, N15273, N2640, N11537);
nor NOR4 (N15278, N15275, N1143, N12340, N10239);
buf BUF1 (N15279, N15270);
xor XOR2 (N15280, N15264, N4584);
buf BUF1 (N15281, N15267);
or OR2 (N15282, N15262, N6938);
and AND2 (N15283, N15279, N8463);
buf BUF1 (N15284, N15277);
nand NAND2 (N15285, N15283, N14673);
or OR4 (N15286, N15282, N11283, N1432, N13761);
not NOT1 (N15287, N15284);
and AND2 (N15288, N15281, N6675);
or OR2 (N15289, N15286, N2351);
xor XOR2 (N15290, N15285, N10248);
xor XOR2 (N15291, N15271, N2002);
buf BUF1 (N15292, N15258);
not NOT1 (N15293, N15291);
or OR4 (N15294, N15280, N8995, N7885, N12332);
nor NOR3 (N15295, N15292, N5075, N6642);
not NOT1 (N15296, N15295);
not NOT1 (N15297, N15289);
buf BUF1 (N15298, N15293);
and AND3 (N15299, N15297, N10385, N10466);
and AND4 (N15300, N15299, N13680, N10988, N6617);
buf BUF1 (N15301, N15276);
or OR3 (N15302, N15269, N3957, N9064);
nor NOR3 (N15303, N15290, N15048, N12884);
and AND2 (N15304, N15296, N10569);
xor XOR2 (N15305, N15298, N13433);
or OR2 (N15306, N15303, N14775);
or OR3 (N15307, N15278, N12563, N13020);
not NOT1 (N15308, N15302);
buf BUF1 (N15309, N15304);
and AND4 (N15310, N15306, N9754, N10279, N12907);
or OR2 (N15311, N15294, N7534);
buf BUF1 (N15312, N15310);
nand NAND4 (N15313, N15288, N3275, N8195, N7166);
or OR3 (N15314, N15313, N3618, N5775);
nor NOR3 (N15315, N15308, N8972, N9145);
and AND3 (N15316, N15307, N3937, N9924);
or OR2 (N15317, N15311, N373);
nand NAND2 (N15318, N15287, N8639);
buf BUF1 (N15319, N15318);
xor XOR2 (N15320, N15317, N13192);
buf BUF1 (N15321, N15301);
and AND2 (N15322, N15321, N4872);
nor NOR2 (N15323, N15322, N4615);
or OR3 (N15324, N15309, N14206, N3554);
or OR4 (N15325, N15305, N1110, N9563, N4400);
nand NAND2 (N15326, N15323, N3344);
nand NAND3 (N15327, N15324, N8287, N6995);
or OR4 (N15328, N15327, N14918, N15155, N1616);
and AND4 (N15329, N15316, N3454, N6397, N1564);
not NOT1 (N15330, N15312);
or OR2 (N15331, N15315, N3441);
not NOT1 (N15332, N15300);
and AND3 (N15333, N15319, N2653, N14266);
not NOT1 (N15334, N15320);
not NOT1 (N15335, N15328);
nor NOR4 (N15336, N15335, N8444, N10039, N14585);
and AND4 (N15337, N15332, N6018, N2049, N6199);
xor XOR2 (N15338, N15333, N227);
nor NOR4 (N15339, N15330, N13046, N2679, N3359);
buf BUF1 (N15340, N15314);
nor NOR4 (N15341, N15336, N2414, N9682, N11927);
xor XOR2 (N15342, N15341, N6888);
xor XOR2 (N15343, N15339, N13549);
and AND2 (N15344, N15340, N748);
buf BUF1 (N15345, N15342);
not NOT1 (N15346, N15343);
xor XOR2 (N15347, N15331, N4770);
nor NOR4 (N15348, N15346, N9595, N3632, N6459);
xor XOR2 (N15349, N15347, N14937);
nor NOR2 (N15350, N15326, N10685);
nor NOR2 (N15351, N15334, N7806);
nor NOR3 (N15352, N15338, N14156, N3745);
nor NOR3 (N15353, N15337, N10257, N8308);
xor XOR2 (N15354, N15352, N12758);
nand NAND3 (N15355, N15351, N2270, N10036);
or OR4 (N15356, N15344, N3617, N10190, N3611);
xor XOR2 (N15357, N15356, N12367);
xor XOR2 (N15358, N15350, N13097);
nor NOR4 (N15359, N15358, N11587, N2236, N4242);
xor XOR2 (N15360, N15359, N14072);
xor XOR2 (N15361, N15357, N1888);
and AND4 (N15362, N15361, N1516, N3109, N14193);
not NOT1 (N15363, N15362);
nand NAND4 (N15364, N15325, N6950, N5606, N12171);
or OR2 (N15365, N15353, N10532);
nor NOR3 (N15366, N15345, N6306, N13182);
xor XOR2 (N15367, N15366, N7009);
nand NAND2 (N15368, N15348, N12280);
or OR3 (N15369, N15354, N7670, N6123);
buf BUF1 (N15370, N15369);
or OR2 (N15371, N15367, N10009);
or OR4 (N15372, N15329, N7757, N3861, N8772);
or OR2 (N15373, N15349, N1451);
xor XOR2 (N15374, N15360, N11204);
or OR4 (N15375, N15372, N10575, N4784, N10384);
not NOT1 (N15376, N15374);
nand NAND2 (N15377, N15365, N4150);
xor XOR2 (N15378, N15377, N1702);
and AND2 (N15379, N15371, N12454);
nand NAND4 (N15380, N15378, N7193, N5616, N2032);
or OR3 (N15381, N15379, N7674, N8237);
xor XOR2 (N15382, N15370, N3883);
not NOT1 (N15383, N15355);
nand NAND2 (N15384, N15364, N2971);
nor NOR4 (N15385, N15373, N2708, N13823, N12045);
buf BUF1 (N15386, N15363);
buf BUF1 (N15387, N15381);
not NOT1 (N15388, N15376);
nor NOR2 (N15389, N15380, N4792);
and AND4 (N15390, N15388, N9214, N5586, N356);
or OR2 (N15391, N15382, N15262);
or OR2 (N15392, N15389, N9237);
nand NAND4 (N15393, N15387, N8455, N4690, N14334);
not NOT1 (N15394, N15386);
and AND4 (N15395, N15393, N9514, N13570, N14050);
nor NOR3 (N15396, N15385, N14069, N3904);
or OR3 (N15397, N15396, N6857, N9159);
xor XOR2 (N15398, N15390, N9693);
nand NAND3 (N15399, N15368, N11975, N14623);
or OR2 (N15400, N15399, N12275);
xor XOR2 (N15401, N15391, N14503);
xor XOR2 (N15402, N15395, N15292);
buf BUF1 (N15403, N15384);
buf BUF1 (N15404, N15392);
xor XOR2 (N15405, N15400, N2177);
not NOT1 (N15406, N15403);
buf BUF1 (N15407, N15404);
buf BUF1 (N15408, N15407);
or OR2 (N15409, N15402, N7618);
nand NAND4 (N15410, N15375, N10593, N12048, N1776);
or OR2 (N15411, N15409, N5190);
not NOT1 (N15412, N15410);
buf BUF1 (N15413, N15397);
xor XOR2 (N15414, N15394, N12962);
xor XOR2 (N15415, N15383, N987);
not NOT1 (N15416, N15405);
nand NAND4 (N15417, N15398, N6667, N12048, N2587);
buf BUF1 (N15418, N15406);
and AND2 (N15419, N15401, N8198);
xor XOR2 (N15420, N15418, N12606);
nor NOR4 (N15421, N15417, N7156, N3334, N14896);
nor NOR4 (N15422, N15414, N13404, N1992, N7590);
buf BUF1 (N15423, N15408);
and AND4 (N15424, N15415, N10533, N11584, N9750);
buf BUF1 (N15425, N15413);
not NOT1 (N15426, N15423);
and AND3 (N15427, N15426, N14011, N5648);
buf BUF1 (N15428, N15412);
not NOT1 (N15429, N15424);
nand NAND4 (N15430, N15420, N1161, N11598, N2726);
not NOT1 (N15431, N15425);
xor XOR2 (N15432, N15429, N5829);
nand NAND3 (N15433, N15431, N7991, N9009);
nand NAND2 (N15434, N15432, N14535);
nand NAND3 (N15435, N15430, N4388, N12972);
xor XOR2 (N15436, N15427, N11279);
not NOT1 (N15437, N15416);
and AND2 (N15438, N15433, N6307);
not NOT1 (N15439, N15422);
and AND3 (N15440, N15436, N12737, N9115);
xor XOR2 (N15441, N15438, N8572);
or OR4 (N15442, N15421, N11521, N11091, N2447);
xor XOR2 (N15443, N15419, N4567);
or OR4 (N15444, N15428, N7114, N10205, N1145);
or OR2 (N15445, N15411, N6536);
not NOT1 (N15446, N15444);
nor NOR3 (N15447, N15446, N6176, N1057);
xor XOR2 (N15448, N15447, N10609);
xor XOR2 (N15449, N15437, N13672);
buf BUF1 (N15450, N15435);
or OR3 (N15451, N15445, N12677, N10552);
not NOT1 (N15452, N15434);
xor XOR2 (N15453, N15442, N3487);
nor NOR4 (N15454, N15450, N12744, N8183, N8937);
buf BUF1 (N15455, N15452);
buf BUF1 (N15456, N15448);
and AND2 (N15457, N15454, N5794);
nand NAND4 (N15458, N15449, N12213, N12321, N13164);
not NOT1 (N15459, N15451);
or OR2 (N15460, N15439, N8781);
or OR4 (N15461, N15458, N11830, N8055, N3076);
xor XOR2 (N15462, N15441, N12507);
xor XOR2 (N15463, N15456, N5908);
or OR3 (N15464, N15457, N10823, N7397);
or OR3 (N15465, N15463, N5835, N11012);
and AND2 (N15466, N15443, N3326);
nand NAND4 (N15467, N15460, N14083, N7595, N6534);
and AND4 (N15468, N15453, N12380, N14039, N711);
nand NAND2 (N15469, N15468, N9662);
buf BUF1 (N15470, N15459);
or OR4 (N15471, N15462, N13226, N2694, N14223);
and AND3 (N15472, N15440, N2788, N8848);
not NOT1 (N15473, N15464);
or OR2 (N15474, N15467, N9973);
nor NOR4 (N15475, N15469, N10973, N2555, N14462);
buf BUF1 (N15476, N15472);
xor XOR2 (N15477, N15455, N13596);
xor XOR2 (N15478, N15474, N495);
nor NOR4 (N15479, N15471, N5437, N13263, N3037);
buf BUF1 (N15480, N15477);
xor XOR2 (N15481, N15478, N6690);
nor NOR4 (N15482, N15465, N540, N13531, N10905);
not NOT1 (N15483, N15473);
or OR2 (N15484, N15475, N1435);
xor XOR2 (N15485, N15466, N5519);
buf BUF1 (N15486, N15479);
not NOT1 (N15487, N15470);
and AND3 (N15488, N15483, N1544, N5250);
or OR2 (N15489, N15484, N1161);
buf BUF1 (N15490, N15481);
not NOT1 (N15491, N15486);
buf BUF1 (N15492, N15476);
nor NOR3 (N15493, N15487, N12443, N9643);
nand NAND3 (N15494, N15489, N12563, N13861);
nor NOR4 (N15495, N15488, N4510, N13792, N1529);
nand NAND3 (N15496, N15493, N9448, N5703);
nor NOR4 (N15497, N15490, N6287, N3531, N2289);
nor NOR2 (N15498, N15497, N11359);
xor XOR2 (N15499, N15498, N13458);
nor NOR3 (N15500, N15485, N9313, N2937);
not NOT1 (N15501, N15495);
nand NAND2 (N15502, N15461, N12305);
not NOT1 (N15503, N15494);
buf BUF1 (N15504, N15491);
buf BUF1 (N15505, N15482);
and AND2 (N15506, N15496, N8661);
not NOT1 (N15507, N15480);
not NOT1 (N15508, N15503);
not NOT1 (N15509, N15508);
not NOT1 (N15510, N15505);
not NOT1 (N15511, N15504);
nor NOR2 (N15512, N15501, N112);
nand NAND4 (N15513, N15507, N7278, N14812, N14341);
buf BUF1 (N15514, N15509);
not NOT1 (N15515, N15512);
xor XOR2 (N15516, N15510, N14018);
buf BUF1 (N15517, N15500);
not NOT1 (N15518, N15515);
nor NOR4 (N15519, N15492, N9393, N10525, N6155);
nor NOR4 (N15520, N15506, N2295, N504, N5909);
nand NAND3 (N15521, N15517, N13567, N12567);
and AND3 (N15522, N15521, N1571, N2429);
and AND2 (N15523, N15511, N2348);
nor NOR3 (N15524, N15499, N7003, N6593);
and AND4 (N15525, N15518, N9680, N2851, N7801);
or OR2 (N15526, N15502, N11752);
and AND3 (N15527, N15514, N2395, N4812);
and AND2 (N15528, N15525, N7401);
nor NOR4 (N15529, N15522, N2522, N2206, N13138);
and AND4 (N15530, N15528, N9437, N3801, N10042);
buf BUF1 (N15531, N15530);
or OR4 (N15532, N15527, N9183, N9345, N10813);
nand NAND3 (N15533, N15519, N3606, N5684);
or OR3 (N15534, N15524, N2423, N1789);
nor NOR2 (N15535, N15513, N14504);
xor XOR2 (N15536, N15535, N1900);
nor NOR2 (N15537, N15533, N11274);
xor XOR2 (N15538, N15534, N13553);
buf BUF1 (N15539, N15531);
nand NAND2 (N15540, N15538, N10333);
nor NOR3 (N15541, N15536, N13814, N7438);
nor NOR3 (N15542, N15540, N11305, N13486);
and AND2 (N15543, N15537, N1836);
buf BUF1 (N15544, N15523);
or OR2 (N15545, N15529, N5605);
buf BUF1 (N15546, N15543);
nor NOR2 (N15547, N15539, N11922);
xor XOR2 (N15548, N15541, N4621);
nand NAND4 (N15549, N15520, N8600, N10586, N6422);
not NOT1 (N15550, N15544);
and AND4 (N15551, N15516, N5249, N3375, N13594);
or OR2 (N15552, N15532, N13824);
nand NAND2 (N15553, N15545, N7791);
xor XOR2 (N15554, N15542, N10522);
buf BUF1 (N15555, N15554);
nand NAND3 (N15556, N15553, N3023, N2099);
and AND4 (N15557, N15551, N646, N13699, N12255);
or OR2 (N15558, N15549, N11509);
buf BUF1 (N15559, N15546);
nor NOR3 (N15560, N15547, N11225, N8344);
and AND3 (N15561, N15555, N9253, N2485);
not NOT1 (N15562, N15550);
or OR4 (N15563, N15526, N7962, N3703, N9554);
nand NAND2 (N15564, N15560, N2322);
and AND4 (N15565, N15563, N13245, N7976, N14589);
not NOT1 (N15566, N15548);
and AND4 (N15567, N15562, N1001, N725, N11693);
and AND2 (N15568, N15558, N4791);
not NOT1 (N15569, N15559);
and AND2 (N15570, N15557, N3674);
not NOT1 (N15571, N15568);
and AND2 (N15572, N15569, N6249);
and AND4 (N15573, N15570, N7329, N86, N8157);
not NOT1 (N15574, N15573);
nor NOR4 (N15575, N15574, N11635, N8101, N797);
nor NOR3 (N15576, N15552, N2150, N13192);
buf BUF1 (N15577, N15571);
buf BUF1 (N15578, N15576);
xor XOR2 (N15579, N15561, N9036);
not NOT1 (N15580, N15556);
buf BUF1 (N15581, N15565);
and AND2 (N15582, N15577, N3309);
nor NOR3 (N15583, N15572, N15285, N15033);
xor XOR2 (N15584, N15581, N4526);
xor XOR2 (N15585, N15582, N6362);
nor NOR3 (N15586, N15584, N10592, N4627);
nor NOR4 (N15587, N15566, N12902, N1860, N5515);
buf BUF1 (N15588, N15579);
nand NAND2 (N15589, N15587, N10956);
not NOT1 (N15590, N15583);
not NOT1 (N15591, N15564);
nor NOR3 (N15592, N15586, N2595, N13925);
nor NOR3 (N15593, N15580, N13637, N14991);
and AND3 (N15594, N15588, N11574, N15070);
not NOT1 (N15595, N15589);
xor XOR2 (N15596, N15575, N5692);
xor XOR2 (N15597, N15590, N7963);
or OR3 (N15598, N15595, N12797, N9120);
and AND2 (N15599, N15596, N12111);
xor XOR2 (N15600, N15592, N12942);
or OR4 (N15601, N15578, N10142, N13431, N13252);
xor XOR2 (N15602, N15598, N13209);
nand NAND4 (N15603, N15594, N5118, N3422, N3968);
xor XOR2 (N15604, N15602, N7858);
nand NAND3 (N15605, N15585, N11572, N1284);
nor NOR4 (N15606, N15603, N7988, N8034, N694);
and AND2 (N15607, N15601, N11171);
nand NAND2 (N15608, N15607, N7327);
not NOT1 (N15609, N15608);
xor XOR2 (N15610, N15605, N4739);
and AND2 (N15611, N15567, N10051);
and AND2 (N15612, N15591, N1343);
nor NOR2 (N15613, N15604, N2629);
and AND2 (N15614, N15593, N2498);
and AND2 (N15615, N15613, N3597);
nand NAND2 (N15616, N15600, N8378);
or OR2 (N15617, N15606, N14463);
nand NAND3 (N15618, N15612, N3201, N11010);
xor XOR2 (N15619, N15597, N8840);
not NOT1 (N15620, N15610);
xor XOR2 (N15621, N15616, N15479);
not NOT1 (N15622, N15620);
nor NOR3 (N15623, N15599, N1068, N14187);
nor NOR2 (N15624, N15615, N13765);
or OR3 (N15625, N15622, N4529, N14469);
nand NAND3 (N15626, N15623, N4827, N4082);
xor XOR2 (N15627, N15621, N642);
not NOT1 (N15628, N15619);
nand NAND4 (N15629, N15609, N5146, N8515, N11436);
and AND4 (N15630, N15614, N8261, N8598, N5631);
or OR4 (N15631, N15626, N326, N1271, N12403);
and AND2 (N15632, N15628, N6869);
or OR3 (N15633, N15629, N8401, N3940);
and AND4 (N15634, N15618, N15609, N5494, N10783);
not NOT1 (N15635, N15611);
buf BUF1 (N15636, N15624);
and AND2 (N15637, N15617, N7792);
or OR4 (N15638, N15631, N10204, N1005, N11074);
buf BUF1 (N15639, N15627);
or OR2 (N15640, N15625, N12066);
or OR2 (N15641, N15633, N10035);
buf BUF1 (N15642, N15641);
or OR4 (N15643, N15639, N6154, N9803, N749);
not NOT1 (N15644, N15630);
and AND4 (N15645, N15636, N10777, N9318, N5607);
and AND2 (N15646, N15643, N2779);
not NOT1 (N15647, N15640);
buf BUF1 (N15648, N15632);
and AND2 (N15649, N15638, N10293);
buf BUF1 (N15650, N15637);
xor XOR2 (N15651, N15646, N13271);
nor NOR4 (N15652, N15645, N14261, N3986, N10225);
buf BUF1 (N15653, N15635);
xor XOR2 (N15654, N15652, N5539);
xor XOR2 (N15655, N15642, N12725);
buf BUF1 (N15656, N15647);
nor NOR3 (N15657, N15656, N6740, N8829);
nor NOR3 (N15658, N15644, N12168, N6097);
xor XOR2 (N15659, N15649, N4822);
nor NOR3 (N15660, N15655, N4419, N13759);
buf BUF1 (N15661, N15658);
nand NAND3 (N15662, N15634, N5819, N234);
or OR2 (N15663, N15662, N11754);
not NOT1 (N15664, N15663);
or OR3 (N15665, N15661, N14763, N7076);
and AND2 (N15666, N15664, N6720);
or OR2 (N15667, N15659, N5624);
not NOT1 (N15668, N15665);
and AND3 (N15669, N15660, N14107, N14384);
nand NAND3 (N15670, N15651, N6254, N14575);
nor NOR4 (N15671, N15648, N11239, N8282, N15375);
or OR4 (N15672, N15657, N152, N9538, N8366);
and AND4 (N15673, N15653, N14075, N2724, N8256);
or OR2 (N15674, N15670, N8645);
xor XOR2 (N15675, N15672, N1940);
buf BUF1 (N15676, N15667);
nand NAND2 (N15677, N15668, N11648);
and AND3 (N15678, N15673, N11326, N11399);
xor XOR2 (N15679, N15666, N4475);
nand NAND2 (N15680, N15674, N1725);
nand NAND3 (N15681, N15669, N5825, N5256);
not NOT1 (N15682, N15681);
nor NOR4 (N15683, N15675, N15157, N4360, N11580);
not NOT1 (N15684, N15650);
xor XOR2 (N15685, N15683, N1705);
nand NAND2 (N15686, N15685, N10642);
buf BUF1 (N15687, N15654);
not NOT1 (N15688, N15679);
buf BUF1 (N15689, N15676);
or OR3 (N15690, N15682, N14819, N9727);
and AND4 (N15691, N15680, N14014, N11484, N6847);
buf BUF1 (N15692, N15678);
and AND2 (N15693, N15686, N4467);
xor XOR2 (N15694, N15692, N8671);
nand NAND4 (N15695, N15677, N8528, N4611, N13936);
nor NOR2 (N15696, N15684, N8357);
xor XOR2 (N15697, N15691, N6528);
and AND3 (N15698, N15687, N3090, N5704);
or OR3 (N15699, N15671, N1306, N8964);
and AND2 (N15700, N15696, N2585);
and AND2 (N15701, N15690, N10948);
and AND4 (N15702, N15697, N14941, N4579, N9218);
not NOT1 (N15703, N15693);
nor NOR3 (N15704, N15700, N4004, N4010);
and AND2 (N15705, N15703, N3961);
or OR4 (N15706, N15695, N10614, N10679, N9404);
nor NOR3 (N15707, N15702, N14250, N2069);
nand NAND2 (N15708, N15707, N1927);
or OR2 (N15709, N15701, N3670);
xor XOR2 (N15710, N15704, N12198);
not NOT1 (N15711, N15698);
nor NOR4 (N15712, N15689, N7170, N3058, N1353);
nand NAND4 (N15713, N15711, N11798, N15609, N3400);
or OR2 (N15714, N15710, N6631);
nand NAND2 (N15715, N15688, N109);
xor XOR2 (N15716, N15706, N10633);
or OR2 (N15717, N15716, N926);
nor NOR2 (N15718, N15712, N7610);
nand NAND4 (N15719, N15694, N12977, N2036, N1204);
xor XOR2 (N15720, N15699, N2645);
and AND4 (N15721, N15718, N6874, N9083, N11261);
buf BUF1 (N15722, N15717);
or OR4 (N15723, N15714, N7918, N9625, N5168);
buf BUF1 (N15724, N15715);
or OR2 (N15725, N15705, N2483);
nor NOR2 (N15726, N15724, N15617);
not NOT1 (N15727, N15725);
xor XOR2 (N15728, N15723, N13539);
xor XOR2 (N15729, N15721, N1603);
and AND4 (N15730, N15727, N3886, N6755, N5243);
xor XOR2 (N15731, N15713, N4799);
not NOT1 (N15732, N15720);
xor XOR2 (N15733, N15722, N15347);
nor NOR4 (N15734, N15709, N8819, N8578, N11104);
or OR3 (N15735, N15729, N2779, N14931);
or OR4 (N15736, N15735, N8435, N5749, N12538);
buf BUF1 (N15737, N15731);
nand NAND2 (N15738, N15733, N557);
nor NOR2 (N15739, N15726, N2411);
or OR3 (N15740, N15736, N3669, N5140);
xor XOR2 (N15741, N15728, N9532);
and AND2 (N15742, N15738, N2600);
not NOT1 (N15743, N15732);
or OR2 (N15744, N15719, N10926);
or OR3 (N15745, N15734, N4139, N15734);
nand NAND4 (N15746, N15708, N14039, N15197, N12620);
or OR2 (N15747, N15746, N3225);
or OR3 (N15748, N15739, N11723, N3280);
buf BUF1 (N15749, N15740);
buf BUF1 (N15750, N15742);
nand NAND4 (N15751, N15744, N10799, N9622, N12103);
not NOT1 (N15752, N15743);
or OR4 (N15753, N15751, N10589, N13073, N9130);
nand NAND4 (N15754, N15737, N12368, N1526, N7402);
nand NAND3 (N15755, N15749, N6992, N13115);
and AND4 (N15756, N15750, N1070, N1407, N15020);
buf BUF1 (N15757, N15730);
not NOT1 (N15758, N15754);
nor NOR3 (N15759, N15757, N7699, N14208);
nor NOR3 (N15760, N15741, N9408, N5273);
buf BUF1 (N15761, N15759);
nand NAND2 (N15762, N15748, N8607);
nor NOR2 (N15763, N15755, N12747);
nor NOR2 (N15764, N15756, N6941);
or OR4 (N15765, N15762, N6107, N7295, N12820);
nor NOR4 (N15766, N15763, N7369, N12874, N10656);
buf BUF1 (N15767, N15745);
and AND2 (N15768, N15753, N6099);
nor NOR3 (N15769, N15752, N6629, N15069);
not NOT1 (N15770, N15765);
xor XOR2 (N15771, N15760, N2917);
buf BUF1 (N15772, N15758);
nor NOR4 (N15773, N15766, N4358, N6113, N9674);
buf BUF1 (N15774, N15769);
buf BUF1 (N15775, N15774);
xor XOR2 (N15776, N15772, N6614);
or OR2 (N15777, N15764, N14186);
buf BUF1 (N15778, N15776);
xor XOR2 (N15779, N15775, N14135);
nor NOR3 (N15780, N15770, N5692, N7961);
nor NOR2 (N15781, N15747, N2161);
xor XOR2 (N15782, N15768, N808);
or OR3 (N15783, N15780, N11987, N8842);
and AND2 (N15784, N15782, N6365);
xor XOR2 (N15785, N15781, N3781);
and AND2 (N15786, N15784, N7049);
buf BUF1 (N15787, N15761);
nor NOR2 (N15788, N15785, N14599);
not NOT1 (N15789, N15779);
not NOT1 (N15790, N15789);
xor XOR2 (N15791, N15773, N12342);
buf BUF1 (N15792, N15767);
nor NOR2 (N15793, N15792, N8660);
and AND2 (N15794, N15778, N1327);
nand NAND2 (N15795, N15794, N8344);
buf BUF1 (N15796, N15795);
nand NAND4 (N15797, N15771, N15530, N11112, N7658);
xor XOR2 (N15798, N15777, N15640);
not NOT1 (N15799, N15791);
or OR3 (N15800, N15786, N10304, N216);
not NOT1 (N15801, N15798);
or OR4 (N15802, N15797, N11975, N11139, N15708);
nand NAND4 (N15803, N15796, N10232, N6636, N2264);
nor NOR2 (N15804, N15801, N5298);
not NOT1 (N15805, N15803);
nand NAND2 (N15806, N15804, N14349);
nor NOR3 (N15807, N15783, N13159, N2550);
not NOT1 (N15808, N15787);
not NOT1 (N15809, N15788);
xor XOR2 (N15810, N15800, N5863);
not NOT1 (N15811, N15799);
not NOT1 (N15812, N15806);
nor NOR4 (N15813, N15805, N2092, N1694, N3343);
and AND3 (N15814, N15813, N2512, N4567);
xor XOR2 (N15815, N15809, N12409);
nand NAND3 (N15816, N15812, N11102, N11567);
and AND2 (N15817, N15808, N6025);
xor XOR2 (N15818, N15817, N7893);
or OR3 (N15819, N15810, N3555, N7294);
or OR3 (N15820, N15815, N7907, N13832);
nor NOR3 (N15821, N15819, N7883, N4473);
xor XOR2 (N15822, N15802, N3888);
and AND4 (N15823, N15793, N2284, N1361, N4310);
nand NAND3 (N15824, N15820, N1875, N12886);
not NOT1 (N15825, N15818);
and AND4 (N15826, N15821, N13255, N8695, N11731);
buf BUF1 (N15827, N15825);
not NOT1 (N15828, N15807);
nand NAND3 (N15829, N15828, N14731, N2159);
or OR3 (N15830, N15790, N14965, N8945);
or OR2 (N15831, N15814, N14407);
xor XOR2 (N15832, N15829, N6572);
nor NOR4 (N15833, N15822, N8072, N1166, N14030);
and AND4 (N15834, N15824, N13200, N2792, N9236);
or OR2 (N15835, N15834, N12295);
nor NOR4 (N15836, N15831, N2513, N14312, N12293);
or OR3 (N15837, N15816, N2608, N4937);
or OR3 (N15838, N15826, N12289, N12571);
nor NOR2 (N15839, N15835, N6209);
nor NOR4 (N15840, N15838, N14754, N14113, N3224);
buf BUF1 (N15841, N15839);
or OR3 (N15842, N15811, N12548, N4689);
or OR4 (N15843, N15827, N4137, N922, N11017);
and AND4 (N15844, N15842, N3956, N14729, N13997);
or OR4 (N15845, N15840, N4068, N12892, N3726);
not NOT1 (N15846, N15844);
not NOT1 (N15847, N15836);
nor NOR3 (N15848, N15837, N8895, N1958);
xor XOR2 (N15849, N15845, N9662);
xor XOR2 (N15850, N15848, N7883);
and AND3 (N15851, N15833, N9700, N4766);
xor XOR2 (N15852, N15832, N5366);
xor XOR2 (N15853, N15843, N1689);
xor XOR2 (N15854, N15846, N3552);
xor XOR2 (N15855, N15823, N13574);
or OR2 (N15856, N15852, N7648);
nand NAND2 (N15857, N15854, N5856);
nor NOR3 (N15858, N15857, N257, N9898);
nand NAND2 (N15859, N15849, N3506);
or OR2 (N15860, N15841, N14526);
nand NAND3 (N15861, N15851, N689, N12707);
nor NOR2 (N15862, N15858, N4889);
and AND2 (N15863, N15847, N1950);
not NOT1 (N15864, N15856);
xor XOR2 (N15865, N15853, N15476);
nor NOR4 (N15866, N15865, N14081, N3535, N13744);
and AND4 (N15867, N15830, N3015, N10339, N6666);
buf BUF1 (N15868, N15860);
not NOT1 (N15869, N15868);
xor XOR2 (N15870, N15864, N555);
nor NOR3 (N15871, N15867, N15681, N6868);
xor XOR2 (N15872, N15855, N2009);
nand NAND3 (N15873, N15861, N388, N8710);
xor XOR2 (N15874, N15862, N587);
nor NOR3 (N15875, N15863, N7265, N1085);
nor NOR2 (N15876, N15875, N4702);
or OR2 (N15877, N15870, N15610);
or OR4 (N15878, N15850, N15597, N2716, N11402);
or OR2 (N15879, N15877, N10142);
nor NOR3 (N15880, N15873, N13247, N1392);
or OR2 (N15881, N15859, N349);
buf BUF1 (N15882, N15874);
not NOT1 (N15883, N15878);
or OR3 (N15884, N15881, N1820, N15382);
nor NOR4 (N15885, N15872, N6014, N3557, N12337);
nor NOR4 (N15886, N15885, N6665, N6649, N828);
not NOT1 (N15887, N15880);
not NOT1 (N15888, N15886);
nand NAND2 (N15889, N15879, N6750);
or OR2 (N15890, N15882, N1711);
buf BUF1 (N15891, N15866);
or OR4 (N15892, N15871, N3434, N9137, N5848);
nand NAND3 (N15893, N15883, N15503, N12010);
xor XOR2 (N15894, N15892, N881);
nor NOR3 (N15895, N15894, N13008, N1352);
and AND4 (N15896, N15889, N5744, N8580, N9344);
nand NAND2 (N15897, N15888, N14255);
not NOT1 (N15898, N15891);
or OR3 (N15899, N15876, N10155, N9869);
buf BUF1 (N15900, N15893);
buf BUF1 (N15901, N15898);
and AND2 (N15902, N15884, N15863);
nor NOR2 (N15903, N15899, N3235);
not NOT1 (N15904, N15901);
and AND2 (N15905, N15869, N10);
not NOT1 (N15906, N15897);
xor XOR2 (N15907, N15887, N1037);
or OR2 (N15908, N15906, N7533);
not NOT1 (N15909, N15890);
and AND2 (N15910, N15900, N11763);
and AND3 (N15911, N15905, N2237, N10649);
and AND2 (N15912, N15907, N14192);
or OR3 (N15913, N15912, N15666, N806);
nor NOR3 (N15914, N15908, N13861, N3943);
nand NAND4 (N15915, N15895, N4418, N303, N11962);
and AND3 (N15916, N15914, N1717, N5918);
nor NOR3 (N15917, N15902, N31, N10300);
not NOT1 (N15918, N15909);
not NOT1 (N15919, N15904);
and AND3 (N15920, N15917, N8957, N14672);
nand NAND2 (N15921, N15915, N9454);
or OR2 (N15922, N15913, N1861);
not NOT1 (N15923, N15922);
xor XOR2 (N15924, N15918, N7213);
xor XOR2 (N15925, N15910, N13603);
or OR2 (N15926, N15903, N10312);
buf BUF1 (N15927, N15926);
not NOT1 (N15928, N15927);
and AND4 (N15929, N15925, N833, N1985, N6705);
nor NOR3 (N15930, N15911, N4662, N905);
buf BUF1 (N15931, N15920);
and AND3 (N15932, N15916, N4078, N3459);
buf BUF1 (N15933, N15923);
not NOT1 (N15934, N15928);
and AND2 (N15935, N15931, N7319);
not NOT1 (N15936, N15921);
or OR2 (N15937, N15933, N15527);
or OR4 (N15938, N15937, N12767, N11912, N5543);
buf BUF1 (N15939, N15929);
xor XOR2 (N15940, N15896, N8134);
buf BUF1 (N15941, N15938);
buf BUF1 (N15942, N15941);
or OR3 (N15943, N15935, N1740, N7678);
buf BUF1 (N15944, N15939);
and AND3 (N15945, N15919, N2367, N15579);
not NOT1 (N15946, N15930);
or OR2 (N15947, N15942, N5397);
nor NOR3 (N15948, N15934, N11420, N4875);
xor XOR2 (N15949, N15945, N10343);
buf BUF1 (N15950, N15940);
not NOT1 (N15951, N15949);
not NOT1 (N15952, N15943);
buf BUF1 (N15953, N15948);
buf BUF1 (N15954, N15947);
and AND2 (N15955, N15944, N9445);
and AND3 (N15956, N15954, N12917, N9083);
nor NOR4 (N15957, N15952, N15287, N7684, N12385);
xor XOR2 (N15958, N15950, N5314);
buf BUF1 (N15959, N15932);
nand NAND3 (N15960, N15951, N2593, N15626);
nor NOR3 (N15961, N15956, N6834, N3859);
buf BUF1 (N15962, N15946);
nand NAND3 (N15963, N15958, N15578, N7607);
nand NAND2 (N15964, N15962, N12409);
xor XOR2 (N15965, N15961, N1899);
xor XOR2 (N15966, N15963, N744);
or OR4 (N15967, N15966, N981, N12607, N13917);
nor NOR3 (N15968, N15960, N7071, N4574);
nand NAND3 (N15969, N15959, N8242, N12235);
xor XOR2 (N15970, N15969, N2160);
and AND4 (N15971, N15936, N15801, N5806, N12478);
nand NAND3 (N15972, N15970, N2732, N1499);
or OR4 (N15973, N15965, N13220, N60, N13300);
nand NAND2 (N15974, N15924, N9165);
nand NAND3 (N15975, N15974, N14421, N11296);
buf BUF1 (N15976, N15968);
nor NOR2 (N15977, N15955, N4766);
nand NAND2 (N15978, N15953, N13226);
nor NOR3 (N15979, N15972, N10320, N8498);
nor NOR3 (N15980, N15967, N3240, N12380);
and AND4 (N15981, N15978, N4003, N5784, N368);
buf BUF1 (N15982, N15957);
buf BUF1 (N15983, N15973);
not NOT1 (N15984, N15975);
or OR3 (N15985, N15964, N8103, N7820);
or OR4 (N15986, N15977, N1723, N7249, N8102);
or OR3 (N15987, N15976, N9613, N14546);
not NOT1 (N15988, N15981);
buf BUF1 (N15989, N15984);
nor NOR2 (N15990, N15979, N13147);
xor XOR2 (N15991, N15990, N5563);
buf BUF1 (N15992, N15989);
buf BUF1 (N15993, N15982);
or OR4 (N15994, N15992, N2974, N4999, N12560);
nand NAND2 (N15995, N15991, N1521);
xor XOR2 (N15996, N15988, N2104);
or OR4 (N15997, N15986, N5824, N11053, N8971);
or OR2 (N15998, N15987, N11395);
not NOT1 (N15999, N15996);
or OR2 (N16000, N15980, N10200);
nor NOR3 (N16001, N15983, N14201, N3019);
buf BUF1 (N16002, N15998);
xor XOR2 (N16003, N15985, N10603);
not NOT1 (N16004, N15997);
nor NOR4 (N16005, N15993, N13295, N6802, N1860);
nor NOR3 (N16006, N16000, N9977, N14411);
xor XOR2 (N16007, N16001, N2809);
or OR2 (N16008, N16005, N2706);
buf BUF1 (N16009, N16007);
or OR3 (N16010, N16004, N3546, N13358);
buf BUF1 (N16011, N16002);
xor XOR2 (N16012, N15999, N9137);
not NOT1 (N16013, N15994);
buf BUF1 (N16014, N16006);
nor NOR3 (N16015, N16010, N866, N8091);
nand NAND2 (N16016, N16011, N6463);
not NOT1 (N16017, N16013);
buf BUF1 (N16018, N16003);
not NOT1 (N16019, N15971);
buf BUF1 (N16020, N16016);
endmodule