// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N25611,N25604,N25607,N25616,N25619,N25618,N25608,N25595,N25617,N25620;

or OR4 (N21, N18, N16, N9, N1);
not NOT1 (N22, N2);
nor NOR2 (N23, N11, N15);
or OR3 (N24, N23, N2, N12);
xor XOR2 (N25, N16, N1);
nand NAND4 (N26, N14, N16, N17, N17);
or OR3 (N27, N3, N22, N21);
nor NOR3 (N28, N17, N26, N4);
nand NAND2 (N29, N17, N16);
buf BUF1 (N30, N22);
not NOT1 (N31, N18);
nor NOR3 (N32, N20, N17, N9);
not NOT1 (N33, N21);
not NOT1 (N34, N6);
nand NAND2 (N35, N25, N27);
xor XOR2 (N36, N27, N29);
and AND2 (N37, N33, N4);
nor NOR2 (N38, N35, N11);
not NOT1 (N39, N24);
buf BUF1 (N40, N31);
and AND3 (N41, N32, N5, N9);
not NOT1 (N42, N20);
or OR2 (N43, N34, N21);
and AND2 (N44, N36, N40);
or OR4 (N45, N27, N22, N3, N8);
nor NOR2 (N46, N38, N18);
xor XOR2 (N47, N42, N38);
nand NAND4 (N48, N37, N15, N33, N14);
and AND2 (N49, N48, N20);
or OR2 (N50, N28, N13);
and AND4 (N51, N39, N31, N49, N37);
buf BUF1 (N52, N1);
buf BUF1 (N53, N43);
buf BUF1 (N54, N45);
and AND4 (N55, N54, N1, N26, N28);
nand NAND4 (N56, N47, N15, N26, N8);
not NOT1 (N57, N52);
nand NAND3 (N58, N51, N24, N56);
and AND4 (N59, N49, N15, N13, N39);
and AND4 (N60, N44, N57, N53, N41);
nand NAND2 (N61, N19, N21);
nor NOR3 (N62, N2, N13, N44);
buf BUF1 (N63, N23);
not NOT1 (N64, N61);
xor XOR2 (N65, N46, N16);
xor XOR2 (N66, N55, N47);
nand NAND4 (N67, N58, N28, N37, N52);
or OR3 (N68, N59, N12, N40);
buf BUF1 (N69, N30);
nor NOR3 (N70, N66, N25, N68);
xor XOR2 (N71, N7, N39);
xor XOR2 (N72, N62, N8);
xor XOR2 (N73, N63, N63);
nor NOR4 (N74, N71, N29, N46, N18);
nand NAND3 (N75, N70, N20, N4);
not NOT1 (N76, N72);
buf BUF1 (N77, N65);
nor NOR3 (N78, N74, N56, N7);
nand NAND3 (N79, N76, N44, N10);
buf BUF1 (N80, N64);
nand NAND2 (N81, N67, N13);
and AND3 (N82, N79, N46, N77);
nand NAND4 (N83, N17, N15, N24, N79);
and AND2 (N84, N80, N10);
xor XOR2 (N85, N84, N72);
nand NAND2 (N86, N69, N25);
not NOT1 (N87, N81);
or OR2 (N88, N83, N4);
and AND4 (N89, N85, N19, N27, N21);
not NOT1 (N90, N75);
nor NOR3 (N91, N88, N21, N27);
not NOT1 (N92, N89);
xor XOR2 (N93, N60, N8);
not NOT1 (N94, N86);
buf BUF1 (N95, N90);
and AND2 (N96, N91, N49);
nor NOR4 (N97, N94, N41, N8, N93);
buf BUF1 (N98, N75);
nor NOR3 (N99, N87, N90, N40);
nor NOR2 (N100, N95, N59);
not NOT1 (N101, N97);
nand NAND4 (N102, N50, N62, N45, N40);
xor XOR2 (N103, N99, N13);
xor XOR2 (N104, N101, N13);
and AND2 (N105, N96, N90);
not NOT1 (N106, N100);
and AND2 (N107, N98, N80);
xor XOR2 (N108, N103, N78);
buf BUF1 (N109, N46);
and AND4 (N110, N108, N15, N31, N93);
and AND2 (N111, N102, N10);
xor XOR2 (N112, N109, N92);
nor NOR2 (N113, N104, N50);
buf BUF1 (N114, N67);
nor NOR4 (N115, N73, N54, N75, N58);
buf BUF1 (N116, N111);
not NOT1 (N117, N107);
or OR2 (N118, N115, N111);
nand NAND4 (N119, N116, N102, N60, N43);
nor NOR2 (N120, N118, N58);
nand NAND2 (N121, N110, N40);
and AND3 (N122, N112, N12, N31);
and AND3 (N123, N114, N53, N19);
nand NAND3 (N124, N105, N14, N62);
not NOT1 (N125, N117);
buf BUF1 (N126, N122);
buf BUF1 (N127, N126);
not NOT1 (N128, N113);
not NOT1 (N129, N124);
and AND3 (N130, N121, N109, N92);
and AND4 (N131, N106, N54, N126, N25);
xor XOR2 (N132, N130, N48);
xor XOR2 (N133, N127, N57);
nand NAND4 (N134, N119, N104, N31, N14);
or OR4 (N135, N131, N106, N21, N36);
buf BUF1 (N136, N134);
nand NAND2 (N137, N120, N52);
and AND2 (N138, N129, N100);
or OR3 (N139, N136, N43, N24);
nor NOR4 (N140, N133, N99, N77, N26);
xor XOR2 (N141, N128, N33);
nor NOR2 (N142, N140, N42);
nand NAND2 (N143, N82, N7);
xor XOR2 (N144, N141, N9);
not NOT1 (N145, N132);
buf BUF1 (N146, N144);
and AND3 (N147, N143, N8, N60);
nand NAND2 (N148, N137, N128);
nor NOR2 (N149, N145, N7);
and AND2 (N150, N123, N17);
and AND4 (N151, N146, N134, N11, N56);
buf BUF1 (N152, N138);
and AND4 (N153, N148, N50, N61, N76);
buf BUF1 (N154, N153);
or OR3 (N155, N125, N71, N132);
or OR2 (N156, N150, N25);
or OR4 (N157, N152, N13, N97, N129);
xor XOR2 (N158, N156, N143);
and AND3 (N159, N158, N152, N78);
or OR2 (N160, N151, N132);
or OR2 (N161, N142, N141);
nor NOR4 (N162, N135, N82, N41, N46);
and AND2 (N163, N162, N117);
and AND3 (N164, N154, N53, N131);
nand NAND2 (N165, N163, N66);
xor XOR2 (N166, N164, N93);
nor NOR4 (N167, N166, N95, N29, N159);
and AND3 (N168, N150, N131, N128);
and AND2 (N169, N165, N63);
buf BUF1 (N170, N157);
not NOT1 (N171, N160);
and AND3 (N172, N149, N117, N95);
buf BUF1 (N173, N171);
nand NAND4 (N174, N139, N14, N128, N14);
nor NOR4 (N175, N173, N89, N143, N151);
and AND3 (N176, N172, N52, N13);
xor XOR2 (N177, N161, N80);
nand NAND4 (N178, N177, N161, N165, N26);
and AND3 (N179, N175, N137, N50);
nand NAND2 (N180, N167, N39);
and AND3 (N181, N178, N146, N129);
and AND2 (N182, N180, N77);
or OR4 (N183, N176, N66, N50, N137);
xor XOR2 (N184, N174, N46);
nor NOR2 (N185, N183, N104);
and AND4 (N186, N184, N52, N25, N2);
or OR2 (N187, N170, N91);
nand NAND4 (N188, N187, N34, N146, N118);
or OR4 (N189, N182, N124, N82, N68);
not NOT1 (N190, N181);
or OR2 (N191, N189, N146);
buf BUF1 (N192, N168);
and AND2 (N193, N186, N163);
xor XOR2 (N194, N169, N144);
buf BUF1 (N195, N147);
and AND2 (N196, N185, N193);
and AND4 (N197, N2, N138, N112, N143);
xor XOR2 (N198, N197, N180);
or OR2 (N199, N198, N174);
buf BUF1 (N200, N179);
and AND3 (N201, N188, N131, N165);
buf BUF1 (N202, N195);
buf BUF1 (N203, N202);
not NOT1 (N204, N200);
or OR2 (N205, N190, N46);
or OR3 (N206, N205, N1, N14);
or OR3 (N207, N194, N15, N177);
nand NAND4 (N208, N203, N149, N119, N152);
xor XOR2 (N209, N155, N129);
and AND2 (N210, N196, N159);
buf BUF1 (N211, N191);
nor NOR2 (N212, N207, N72);
and AND2 (N213, N192, N105);
and AND2 (N214, N201, N205);
not NOT1 (N215, N199);
xor XOR2 (N216, N214, N170);
and AND2 (N217, N212, N92);
buf BUF1 (N218, N204);
not NOT1 (N219, N210);
xor XOR2 (N220, N209, N35);
xor XOR2 (N221, N220, N191);
and AND2 (N222, N215, N17);
not NOT1 (N223, N208);
nor NOR3 (N224, N219, N144, N177);
nor NOR2 (N225, N224, N14);
nand NAND3 (N226, N218, N197, N114);
nand NAND4 (N227, N221, N162, N11, N177);
and AND2 (N228, N216, N187);
nand NAND4 (N229, N217, N5, N53, N185);
or OR4 (N230, N213, N198, N179, N30);
xor XOR2 (N231, N229, N20);
buf BUF1 (N232, N223);
and AND3 (N233, N225, N192, N17);
nor NOR4 (N234, N233, N154, N150, N5);
buf BUF1 (N235, N227);
or OR3 (N236, N222, N3, N67);
nand NAND4 (N237, N234, N195, N236, N121);
or OR2 (N238, N33, N184);
nor NOR2 (N239, N228, N179);
nor NOR2 (N240, N230, N216);
xor XOR2 (N241, N239, N67);
or OR4 (N242, N231, N208, N52, N178);
xor XOR2 (N243, N237, N51);
or OR3 (N244, N211, N73, N193);
nor NOR3 (N245, N238, N171, N152);
not NOT1 (N246, N243);
and AND3 (N247, N245, N236, N234);
and AND2 (N248, N247, N167);
nand NAND4 (N249, N242, N235, N14, N58);
not NOT1 (N250, N12);
buf BUF1 (N251, N249);
nor NOR4 (N252, N246, N30, N131, N180);
nand NAND2 (N253, N232, N139);
not NOT1 (N254, N248);
nand NAND4 (N255, N250, N74, N26, N35);
and AND2 (N256, N255, N160);
xor XOR2 (N257, N256, N47);
xor XOR2 (N258, N254, N55);
not NOT1 (N259, N252);
or OR4 (N260, N253, N111, N62, N219);
nor NOR4 (N261, N251, N122, N19, N78);
or OR4 (N262, N259, N194, N139, N224);
not NOT1 (N263, N241);
buf BUF1 (N264, N262);
nor NOR3 (N265, N226, N253, N213);
and AND3 (N266, N260, N240, N245);
nor NOR3 (N267, N163, N133, N109);
or OR2 (N268, N258, N153);
buf BUF1 (N269, N268);
nand NAND3 (N270, N264, N158, N8);
and AND4 (N271, N261, N184, N56, N219);
nor NOR3 (N272, N270, N20, N59);
nor NOR4 (N273, N266, N231, N229, N53);
buf BUF1 (N274, N265);
or OR4 (N275, N257, N265, N133, N243);
nor NOR2 (N276, N273, N268);
nand NAND2 (N277, N275, N169);
nor NOR2 (N278, N274, N81);
nor NOR2 (N279, N276, N165);
not NOT1 (N280, N263);
and AND2 (N281, N206, N7);
or OR2 (N282, N280, N68);
and AND3 (N283, N277, N34, N199);
nand NAND4 (N284, N271, N256, N200, N60);
not NOT1 (N285, N279);
not NOT1 (N286, N267);
xor XOR2 (N287, N282, N245);
not NOT1 (N288, N244);
nand NAND3 (N289, N287, N138, N31);
buf BUF1 (N290, N283);
nor NOR3 (N291, N284, N225, N235);
xor XOR2 (N292, N272, N171);
and AND2 (N293, N269, N210);
or OR4 (N294, N288, N19, N207, N146);
xor XOR2 (N295, N286, N281);
xor XOR2 (N296, N231, N33);
not NOT1 (N297, N291);
nand NAND2 (N298, N297, N40);
nand NAND4 (N299, N292, N283, N41, N120);
and AND4 (N300, N278, N163, N298, N51);
xor XOR2 (N301, N236, N42);
not NOT1 (N302, N293);
not NOT1 (N303, N301);
xor XOR2 (N304, N300, N105);
not NOT1 (N305, N290);
nor NOR3 (N306, N289, N294, N4);
and AND2 (N307, N156, N46);
nand NAND4 (N308, N303, N34, N263, N162);
or OR4 (N309, N307, N141, N202, N191);
xor XOR2 (N310, N299, N139);
buf BUF1 (N311, N308);
or OR3 (N312, N305, N83, N239);
or OR4 (N313, N285, N266, N140, N211);
not NOT1 (N314, N302);
not NOT1 (N315, N309);
buf BUF1 (N316, N314);
buf BUF1 (N317, N312);
nand NAND3 (N318, N295, N124, N47);
nand NAND4 (N319, N316, N225, N245, N211);
or OR2 (N320, N306, N8);
nor NOR4 (N321, N315, N126, N153, N48);
nor NOR3 (N322, N321, N123, N286);
nand NAND3 (N323, N317, N235, N201);
nand NAND4 (N324, N311, N247, N255, N260);
not NOT1 (N325, N304);
buf BUF1 (N326, N325);
xor XOR2 (N327, N313, N263);
or OR3 (N328, N323, N142, N264);
or OR4 (N329, N310, N266, N237, N169);
buf BUF1 (N330, N329);
buf BUF1 (N331, N318);
nor NOR3 (N332, N331, N215, N273);
and AND3 (N333, N319, N69, N100);
xor XOR2 (N334, N327, N47);
xor XOR2 (N335, N333, N331);
or OR4 (N336, N326, N51, N5, N176);
nor NOR4 (N337, N334, N136, N153, N95);
nor NOR3 (N338, N336, N266, N269);
and AND4 (N339, N322, N190, N110, N8);
xor XOR2 (N340, N330, N315);
nand NAND4 (N341, N338, N88, N238, N73);
not NOT1 (N342, N296);
or OR4 (N343, N332, N15, N110, N302);
and AND2 (N344, N320, N36);
buf BUF1 (N345, N342);
nand NAND2 (N346, N335, N301);
nor NOR3 (N347, N324, N6, N114);
nand NAND4 (N348, N345, N17, N118, N218);
buf BUF1 (N349, N341);
nor NOR2 (N350, N344, N79);
nor NOR3 (N351, N337, N231, N125);
nand NAND4 (N352, N340, N80, N239, N136);
not NOT1 (N353, N343);
buf BUF1 (N354, N328);
or OR2 (N355, N351, N82);
or OR4 (N356, N349, N9, N168, N129);
nor NOR4 (N357, N339, N65, N269, N206);
nand NAND3 (N358, N355, N265, N324);
not NOT1 (N359, N347);
and AND4 (N360, N353, N130, N13, N10);
xor XOR2 (N361, N356, N203);
nand NAND4 (N362, N346, N3, N300, N194);
and AND2 (N363, N358, N141);
or OR2 (N364, N363, N112);
or OR2 (N365, N359, N330);
or OR3 (N366, N362, N166, N94);
xor XOR2 (N367, N361, N39);
or OR4 (N368, N357, N350, N49, N278);
and AND3 (N369, N127, N9, N173);
buf BUF1 (N370, N369);
or OR4 (N371, N370, N342, N212, N121);
xor XOR2 (N372, N367, N71);
and AND4 (N373, N364, N55, N253, N173);
not NOT1 (N374, N348);
and AND4 (N375, N371, N207, N322, N92);
not NOT1 (N376, N368);
not NOT1 (N377, N372);
nand NAND4 (N378, N354, N237, N26, N167);
nand NAND3 (N379, N366, N71, N184);
nand NAND4 (N380, N374, N139, N55, N37);
nor NOR2 (N381, N352, N225);
nor NOR2 (N382, N376, N227);
not NOT1 (N383, N380);
and AND3 (N384, N383, N128, N67);
nor NOR2 (N385, N373, N375);
nand NAND3 (N386, N111, N345, N344);
buf BUF1 (N387, N365);
buf BUF1 (N388, N381);
buf BUF1 (N389, N384);
nor NOR4 (N390, N382, N34, N236, N105);
buf BUF1 (N391, N360);
nor NOR2 (N392, N388, N272);
or OR4 (N393, N387, N42, N231, N49);
or OR2 (N394, N378, N179);
and AND4 (N395, N386, N330, N22, N217);
and AND3 (N396, N379, N234, N237);
xor XOR2 (N397, N377, N99);
or OR3 (N398, N390, N245, N72);
and AND2 (N399, N397, N56);
not NOT1 (N400, N392);
or OR2 (N401, N395, N86);
xor XOR2 (N402, N398, N13);
and AND3 (N403, N401, N42, N353);
xor XOR2 (N404, N394, N182);
nor NOR4 (N405, N389, N113, N101, N236);
xor XOR2 (N406, N400, N78);
buf BUF1 (N407, N391);
or OR2 (N408, N403, N61);
not NOT1 (N409, N408);
buf BUF1 (N410, N404);
and AND4 (N411, N410, N362, N48, N338);
nand NAND4 (N412, N409, N256, N287, N31);
xor XOR2 (N413, N385, N275);
not NOT1 (N414, N402);
xor XOR2 (N415, N407, N245);
and AND3 (N416, N399, N305, N316);
and AND4 (N417, N411, N67, N391, N124);
nand NAND2 (N418, N414, N225);
not NOT1 (N419, N412);
or OR2 (N420, N416, N281);
nand NAND4 (N421, N417, N297, N52, N316);
or OR2 (N422, N413, N37);
buf BUF1 (N423, N422);
xor XOR2 (N424, N396, N293);
or OR2 (N425, N418, N272);
not NOT1 (N426, N420);
nor NOR4 (N427, N426, N164, N338, N398);
or OR3 (N428, N423, N194, N59);
not NOT1 (N429, N421);
buf BUF1 (N430, N419);
nor NOR4 (N431, N427, N254, N397, N344);
xor XOR2 (N432, N424, N16);
or OR2 (N433, N425, N239);
or OR4 (N434, N432, N136, N109, N156);
nand NAND3 (N435, N405, N164, N55);
or OR3 (N436, N429, N341, N181);
not NOT1 (N437, N434);
nor NOR4 (N438, N430, N240, N407, N409);
not NOT1 (N439, N433);
not NOT1 (N440, N415);
and AND2 (N441, N438, N2);
or OR3 (N442, N440, N296, N36);
buf BUF1 (N443, N439);
buf BUF1 (N444, N441);
xor XOR2 (N445, N444, N189);
nand NAND2 (N446, N443, N259);
nand NAND3 (N447, N431, N142, N401);
not NOT1 (N448, N435);
buf BUF1 (N449, N437);
or OR3 (N450, N446, N342, N402);
xor XOR2 (N451, N406, N96);
not NOT1 (N452, N449);
and AND4 (N453, N445, N123, N266, N289);
or OR3 (N454, N447, N391, N85);
and AND4 (N455, N448, N334, N10, N117);
and AND3 (N456, N442, N79, N328);
nand NAND4 (N457, N455, N124, N437, N20);
not NOT1 (N458, N450);
buf BUF1 (N459, N393);
xor XOR2 (N460, N436, N220);
xor XOR2 (N461, N456, N459);
not NOT1 (N462, N137);
nand NAND3 (N463, N460, N134, N227);
not NOT1 (N464, N428);
xor XOR2 (N465, N453, N240);
xor XOR2 (N466, N462, N33);
buf BUF1 (N467, N461);
and AND3 (N468, N465, N98, N202);
xor XOR2 (N469, N457, N85);
nor NOR3 (N470, N467, N163, N228);
or OR3 (N471, N470, N355, N335);
or OR3 (N472, N463, N178, N431);
or OR2 (N473, N472, N313);
not NOT1 (N474, N468);
and AND4 (N475, N451, N82, N115, N356);
and AND3 (N476, N452, N427, N466);
buf BUF1 (N477, N69);
buf BUF1 (N478, N469);
nor NOR3 (N479, N471, N428, N3);
buf BUF1 (N480, N478);
xor XOR2 (N481, N479, N226);
and AND2 (N482, N474, N341);
or OR3 (N483, N454, N238, N307);
or OR3 (N484, N476, N283, N13);
xor XOR2 (N485, N481, N16);
nand NAND4 (N486, N475, N411, N69, N232);
nor NOR2 (N487, N485, N148);
xor XOR2 (N488, N464, N451);
xor XOR2 (N489, N488, N382);
nor NOR2 (N490, N487, N475);
or OR2 (N491, N458, N290);
and AND2 (N492, N489, N129);
xor XOR2 (N493, N483, N416);
not NOT1 (N494, N491);
nand NAND3 (N495, N490, N56, N72);
xor XOR2 (N496, N484, N207);
buf BUF1 (N497, N477);
and AND2 (N498, N494, N70);
not NOT1 (N499, N493);
buf BUF1 (N500, N495);
xor XOR2 (N501, N499, N352);
nand NAND4 (N502, N496, N470, N155, N167);
not NOT1 (N503, N500);
xor XOR2 (N504, N503, N84);
not NOT1 (N505, N492);
not NOT1 (N506, N482);
or OR3 (N507, N502, N471, N94);
not NOT1 (N508, N507);
and AND2 (N509, N480, N86);
or OR2 (N510, N486, N59);
buf BUF1 (N511, N510);
xor XOR2 (N512, N498, N128);
and AND4 (N513, N509, N469, N333, N19);
and AND3 (N514, N513, N254, N366);
xor XOR2 (N515, N497, N204);
and AND2 (N516, N511, N29);
nor NOR4 (N517, N508, N414, N416, N173);
or OR3 (N518, N473, N325, N208);
xor XOR2 (N519, N505, N373);
nand NAND3 (N520, N504, N382, N114);
and AND4 (N521, N506, N362, N511, N457);
not NOT1 (N522, N521);
xor XOR2 (N523, N515, N333);
nand NAND4 (N524, N523, N310, N362, N209);
nor NOR2 (N525, N516, N452);
and AND2 (N526, N518, N229);
or OR3 (N527, N517, N337, N339);
nor NOR2 (N528, N514, N158);
not NOT1 (N529, N512);
xor XOR2 (N530, N525, N425);
and AND3 (N531, N527, N301, N62);
or OR2 (N532, N531, N132);
nor NOR4 (N533, N524, N62, N310, N95);
and AND2 (N534, N529, N432);
and AND4 (N535, N501, N125, N47, N381);
nor NOR2 (N536, N528, N127);
nand NAND2 (N537, N535, N363);
not NOT1 (N538, N533);
and AND2 (N539, N530, N79);
nor NOR2 (N540, N536, N393);
and AND2 (N541, N539, N158);
xor XOR2 (N542, N522, N498);
and AND3 (N543, N526, N481, N406);
xor XOR2 (N544, N520, N506);
not NOT1 (N545, N534);
xor XOR2 (N546, N541, N510);
nor NOR4 (N547, N544, N336, N545, N98);
buf BUF1 (N548, N526);
xor XOR2 (N549, N546, N95);
buf BUF1 (N550, N538);
not NOT1 (N551, N519);
buf BUF1 (N552, N537);
xor XOR2 (N553, N540, N543);
not NOT1 (N554, N173);
not NOT1 (N555, N550);
not NOT1 (N556, N542);
nand NAND2 (N557, N551, N480);
nor NOR2 (N558, N557, N343);
not NOT1 (N559, N553);
xor XOR2 (N560, N532, N22);
nor NOR4 (N561, N552, N382, N151, N260);
buf BUF1 (N562, N556);
and AND4 (N563, N558, N300, N62, N350);
or OR4 (N564, N548, N75, N234, N388);
xor XOR2 (N565, N549, N424);
or OR2 (N566, N561, N454);
not NOT1 (N567, N560);
or OR4 (N568, N562, N556, N521, N215);
nand NAND3 (N569, N568, N66, N258);
buf BUF1 (N570, N555);
and AND4 (N571, N569, N19, N377, N375);
or OR2 (N572, N559, N156);
nand NAND2 (N573, N563, N571);
buf BUF1 (N574, N442);
buf BUF1 (N575, N572);
or OR3 (N576, N554, N270, N132);
not NOT1 (N577, N575);
not NOT1 (N578, N573);
buf BUF1 (N579, N578);
nor NOR3 (N580, N567, N68, N473);
nor NOR4 (N581, N566, N467, N306, N160);
nand NAND4 (N582, N579, N225, N58, N392);
buf BUF1 (N583, N576);
and AND3 (N584, N581, N504, N365);
or OR4 (N585, N584, N20, N28, N505);
buf BUF1 (N586, N574);
xor XOR2 (N587, N547, N112);
buf BUF1 (N588, N564);
nor NOR2 (N589, N582, N37);
nor NOR4 (N590, N588, N432, N144, N244);
not NOT1 (N591, N577);
not NOT1 (N592, N580);
or OR4 (N593, N589, N325, N120, N392);
nor NOR3 (N594, N592, N139, N260);
and AND2 (N595, N591, N563);
buf BUF1 (N596, N595);
and AND3 (N597, N570, N56, N197);
xor XOR2 (N598, N594, N292);
xor XOR2 (N599, N565, N446);
and AND2 (N600, N597, N336);
not NOT1 (N601, N599);
nand NAND3 (N602, N583, N217, N241);
nor NOR4 (N603, N598, N367, N59, N129);
and AND2 (N604, N596, N373);
xor XOR2 (N605, N587, N531);
and AND4 (N606, N593, N237, N575, N42);
nand NAND4 (N607, N590, N534, N194, N348);
or OR4 (N608, N585, N586, N551, N356);
xor XOR2 (N609, N454, N200);
xor XOR2 (N610, N608, N345);
not NOT1 (N611, N610);
xor XOR2 (N612, N604, N384);
nand NAND2 (N613, N605, N231);
nand NAND4 (N614, N600, N613, N399, N136);
xor XOR2 (N615, N79, N315);
or OR4 (N616, N603, N228, N66, N306);
not NOT1 (N617, N616);
nand NAND4 (N618, N606, N259, N177, N4);
nand NAND2 (N619, N611, N561);
not NOT1 (N620, N612);
and AND3 (N621, N609, N462, N175);
and AND4 (N622, N621, N542, N465, N62);
buf BUF1 (N623, N601);
xor XOR2 (N624, N615, N454);
not NOT1 (N625, N614);
xor XOR2 (N626, N602, N161);
or OR2 (N627, N619, N557);
not NOT1 (N628, N607);
or OR3 (N629, N627, N401, N531);
nand NAND4 (N630, N629, N568, N577, N335);
nand NAND4 (N631, N624, N443, N351, N189);
buf BUF1 (N632, N628);
not NOT1 (N633, N632);
or OR3 (N634, N630, N589, N152);
and AND4 (N635, N633, N176, N521, N530);
and AND3 (N636, N625, N176, N364);
nand NAND4 (N637, N636, N86, N67, N240);
buf BUF1 (N638, N623);
buf BUF1 (N639, N622);
or OR2 (N640, N618, N584);
nor NOR2 (N641, N631, N238);
and AND4 (N642, N640, N23, N596, N194);
and AND2 (N643, N642, N215);
xor XOR2 (N644, N643, N30);
xor XOR2 (N645, N620, N77);
or OR4 (N646, N617, N233, N342, N56);
buf BUF1 (N647, N634);
xor XOR2 (N648, N638, N378);
xor XOR2 (N649, N626, N533);
buf BUF1 (N650, N637);
nor NOR2 (N651, N648, N87);
and AND4 (N652, N646, N89, N23, N549);
and AND2 (N653, N641, N273);
not NOT1 (N654, N645);
nand NAND3 (N655, N649, N636, N285);
or OR2 (N656, N651, N364);
not NOT1 (N657, N654);
nor NOR2 (N658, N635, N483);
nand NAND4 (N659, N644, N491, N523, N221);
xor XOR2 (N660, N657, N569);
or OR3 (N661, N656, N517, N306);
or OR2 (N662, N652, N133);
xor XOR2 (N663, N647, N290);
or OR3 (N664, N660, N544, N470);
not NOT1 (N665, N664);
nor NOR2 (N666, N658, N429);
nor NOR3 (N667, N666, N405, N497);
or OR3 (N668, N662, N504, N601);
xor XOR2 (N669, N655, N465);
nor NOR4 (N670, N668, N203, N27, N25);
nand NAND3 (N671, N663, N604, N470);
and AND2 (N672, N639, N451);
nor NOR3 (N673, N667, N549, N463);
or OR3 (N674, N653, N654, N502);
nand NAND4 (N675, N672, N271, N405, N431);
and AND3 (N676, N674, N66, N142);
xor XOR2 (N677, N659, N540);
and AND3 (N678, N669, N294, N634);
xor XOR2 (N679, N661, N175);
nor NOR3 (N680, N673, N512, N463);
and AND4 (N681, N679, N134, N313, N343);
and AND2 (N682, N650, N257);
and AND3 (N683, N678, N94, N504);
or OR4 (N684, N677, N145, N491, N258);
nand NAND2 (N685, N683, N253);
or OR2 (N686, N671, N412);
nand NAND4 (N687, N680, N398, N166, N647);
xor XOR2 (N688, N685, N325);
xor XOR2 (N689, N675, N370);
nand NAND4 (N690, N670, N196, N130, N464);
or OR4 (N691, N687, N154, N140, N477);
or OR2 (N692, N682, N582);
buf BUF1 (N693, N689);
nor NOR4 (N694, N691, N555, N25, N176);
xor XOR2 (N695, N676, N540);
buf BUF1 (N696, N684);
nand NAND4 (N697, N665, N79, N576, N387);
xor XOR2 (N698, N681, N320);
xor XOR2 (N699, N696, N653);
xor XOR2 (N700, N697, N233);
buf BUF1 (N701, N690);
xor XOR2 (N702, N700, N599);
nand NAND4 (N703, N701, N669, N316, N106);
buf BUF1 (N704, N694);
nor NOR4 (N705, N704, N2, N457, N294);
or OR3 (N706, N702, N355, N671);
buf BUF1 (N707, N693);
buf BUF1 (N708, N698);
buf BUF1 (N709, N699);
nor NOR3 (N710, N708, N32, N662);
and AND4 (N711, N688, N43, N518, N410);
nand NAND3 (N712, N705, N159, N94);
not NOT1 (N713, N711);
nor NOR3 (N714, N707, N210, N5);
nor NOR2 (N715, N710, N5);
nor NOR2 (N716, N695, N699);
and AND4 (N717, N706, N643, N355, N480);
nor NOR4 (N718, N713, N169, N280, N681);
nand NAND4 (N719, N718, N346, N239, N374);
xor XOR2 (N720, N686, N324);
or OR2 (N721, N712, N68);
and AND3 (N722, N692, N511, N50);
or OR3 (N723, N722, N171, N97);
xor XOR2 (N724, N716, N674);
nor NOR4 (N725, N709, N568, N172, N73);
or OR3 (N726, N725, N109, N38);
buf BUF1 (N727, N723);
nor NOR2 (N728, N717, N653);
not NOT1 (N729, N719);
and AND3 (N730, N729, N590, N283);
xor XOR2 (N731, N721, N430);
nand NAND4 (N732, N703, N715, N644, N106);
nand NAND4 (N733, N298, N232, N409, N276);
or OR2 (N734, N714, N580);
xor XOR2 (N735, N731, N174);
buf BUF1 (N736, N732);
nand NAND4 (N737, N730, N75, N530, N389);
not NOT1 (N738, N720);
buf BUF1 (N739, N738);
not NOT1 (N740, N736);
not NOT1 (N741, N734);
and AND2 (N742, N739, N451);
xor XOR2 (N743, N724, N302);
not NOT1 (N744, N733);
nor NOR2 (N745, N740, N87);
xor XOR2 (N746, N728, N647);
xor XOR2 (N747, N741, N623);
nor NOR4 (N748, N742, N33, N143, N219);
xor XOR2 (N749, N748, N605);
and AND2 (N750, N744, N6);
and AND4 (N751, N735, N347, N171, N600);
xor XOR2 (N752, N727, N371);
buf BUF1 (N753, N747);
buf BUF1 (N754, N753);
nand NAND4 (N755, N749, N491, N596, N438);
nor NOR4 (N756, N752, N250, N427, N135);
not NOT1 (N757, N754);
buf BUF1 (N758, N746);
and AND2 (N759, N755, N703);
not NOT1 (N760, N758);
not NOT1 (N761, N760);
xor XOR2 (N762, N761, N25);
nor NOR3 (N763, N726, N219, N445);
not NOT1 (N764, N762);
and AND2 (N765, N759, N302);
or OR2 (N766, N745, N529);
or OR4 (N767, N766, N164, N571, N157);
buf BUF1 (N768, N750);
nand NAND2 (N769, N768, N187);
and AND2 (N770, N756, N751);
and AND2 (N771, N520, N553);
nor NOR3 (N772, N737, N761, N98);
nor NOR4 (N773, N771, N48, N761, N409);
nor NOR4 (N774, N743, N653, N722, N624);
nand NAND2 (N775, N772, N739);
nor NOR3 (N776, N757, N774, N232);
not NOT1 (N777, N186);
and AND2 (N778, N777, N544);
nor NOR4 (N779, N764, N639, N54, N734);
nor NOR4 (N780, N763, N608, N294, N403);
nor NOR4 (N781, N765, N177, N2, N512);
or OR4 (N782, N780, N146, N187, N139);
xor XOR2 (N783, N779, N749);
and AND4 (N784, N767, N158, N298, N580);
xor XOR2 (N785, N775, N661);
xor XOR2 (N786, N778, N86);
not NOT1 (N787, N770);
not NOT1 (N788, N787);
not NOT1 (N789, N773);
and AND4 (N790, N769, N374, N514, N200);
xor XOR2 (N791, N789, N536);
nand NAND4 (N792, N784, N705, N475, N730);
xor XOR2 (N793, N788, N212);
xor XOR2 (N794, N782, N135);
not NOT1 (N795, N794);
xor XOR2 (N796, N790, N596);
buf BUF1 (N797, N776);
nand NAND4 (N798, N785, N280, N487, N188);
nor NOR2 (N799, N781, N408);
buf BUF1 (N800, N792);
xor XOR2 (N801, N800, N531);
buf BUF1 (N802, N791);
not NOT1 (N803, N795);
buf BUF1 (N804, N801);
not NOT1 (N805, N799);
nor NOR2 (N806, N793, N399);
nor NOR4 (N807, N783, N469, N629, N566);
or OR3 (N808, N797, N448, N734);
not NOT1 (N809, N806);
xor XOR2 (N810, N803, N147);
xor XOR2 (N811, N796, N326);
xor XOR2 (N812, N807, N761);
buf BUF1 (N813, N798);
xor XOR2 (N814, N802, N117);
and AND2 (N815, N809, N148);
not NOT1 (N816, N811);
not NOT1 (N817, N815);
not NOT1 (N818, N813);
buf BUF1 (N819, N810);
or OR4 (N820, N804, N640, N356, N562);
and AND2 (N821, N812, N696);
not NOT1 (N822, N817);
and AND2 (N823, N818, N535);
not NOT1 (N824, N816);
buf BUF1 (N825, N814);
buf BUF1 (N826, N822);
xor XOR2 (N827, N825, N329);
or OR4 (N828, N826, N421, N324, N483);
xor XOR2 (N829, N808, N525);
nor NOR4 (N830, N786, N660, N582, N183);
nand NAND3 (N831, N805, N465, N325);
xor XOR2 (N832, N821, N218);
buf BUF1 (N833, N819);
or OR2 (N834, N828, N369);
xor XOR2 (N835, N830, N214);
or OR2 (N836, N820, N48);
xor XOR2 (N837, N829, N386);
and AND4 (N838, N832, N525, N33, N302);
nor NOR2 (N839, N835, N835);
nor NOR3 (N840, N833, N115, N700);
or OR2 (N841, N824, N623);
not NOT1 (N842, N838);
or OR4 (N843, N836, N348, N467, N473);
xor XOR2 (N844, N839, N324);
nand NAND3 (N845, N840, N516, N437);
nor NOR4 (N846, N834, N130, N827, N484);
not NOT1 (N847, N229);
or OR4 (N848, N837, N232, N559, N694);
nor NOR2 (N849, N823, N623);
nand NAND2 (N850, N831, N668);
nand NAND3 (N851, N843, N6, N534);
or OR4 (N852, N847, N754, N284, N767);
or OR2 (N853, N841, N29);
xor XOR2 (N854, N842, N128);
and AND2 (N855, N848, N14);
buf BUF1 (N856, N854);
and AND3 (N857, N846, N302, N411);
buf BUF1 (N858, N845);
nor NOR3 (N859, N851, N840, N706);
and AND2 (N860, N849, N674);
nand NAND4 (N861, N855, N805, N4, N756);
not NOT1 (N862, N853);
or OR3 (N863, N850, N594, N18);
or OR4 (N864, N861, N681, N451, N314);
and AND3 (N865, N852, N34, N471);
buf BUF1 (N866, N863);
not NOT1 (N867, N866);
buf BUF1 (N868, N856);
not NOT1 (N869, N865);
not NOT1 (N870, N859);
or OR4 (N871, N870, N136, N475, N258);
nand NAND3 (N872, N858, N860, N85);
and AND2 (N873, N505, N421);
xor XOR2 (N874, N857, N656);
and AND2 (N875, N872, N632);
and AND4 (N876, N864, N682, N222, N103);
nor NOR2 (N877, N876, N45);
not NOT1 (N878, N874);
buf BUF1 (N879, N877);
nand NAND4 (N880, N878, N304, N624, N355);
nor NOR2 (N881, N873, N549);
xor XOR2 (N882, N875, N615);
not NOT1 (N883, N862);
or OR4 (N884, N883, N453, N684, N77);
not NOT1 (N885, N882);
xor XOR2 (N886, N885, N569);
buf BUF1 (N887, N867);
nand NAND2 (N888, N869, N648);
nor NOR3 (N889, N879, N878, N685);
buf BUF1 (N890, N884);
nand NAND3 (N891, N844, N804, N688);
or OR2 (N892, N880, N201);
and AND3 (N893, N881, N302, N823);
xor XOR2 (N894, N887, N47);
or OR3 (N895, N886, N741, N166);
not NOT1 (N896, N868);
buf BUF1 (N897, N892);
buf BUF1 (N898, N889);
buf BUF1 (N899, N896);
nor NOR4 (N900, N897, N527, N18, N441);
and AND4 (N901, N898, N823, N39, N213);
buf BUF1 (N902, N891);
xor XOR2 (N903, N871, N623);
and AND4 (N904, N900, N810, N798, N755);
buf BUF1 (N905, N902);
xor XOR2 (N906, N905, N87);
and AND2 (N907, N901, N343);
or OR3 (N908, N906, N818, N808);
nor NOR3 (N909, N888, N765, N688);
xor XOR2 (N910, N894, N788);
xor XOR2 (N911, N893, N290);
buf BUF1 (N912, N890);
or OR4 (N913, N909, N736, N730, N112);
buf BUF1 (N914, N899);
nor NOR4 (N915, N903, N89, N914, N81);
nor NOR3 (N916, N30, N173, N548);
nand NAND4 (N917, N916, N384, N786, N452);
and AND3 (N918, N904, N821, N345);
and AND2 (N919, N910, N381);
nor NOR3 (N920, N911, N878, N912);
xor XOR2 (N921, N223, N6);
nand NAND4 (N922, N895, N365, N251, N695);
buf BUF1 (N923, N908);
or OR3 (N924, N922, N873, N261);
nand NAND2 (N925, N918, N762);
not NOT1 (N926, N921);
not NOT1 (N927, N907);
and AND4 (N928, N915, N728, N487, N719);
nand NAND4 (N929, N926, N76, N245, N66);
not NOT1 (N930, N920);
xor XOR2 (N931, N924, N439);
not NOT1 (N932, N927);
or OR2 (N933, N931, N170);
and AND3 (N934, N923, N876, N893);
and AND3 (N935, N913, N124, N417);
and AND3 (N936, N935, N888, N164);
and AND4 (N937, N933, N390, N278, N559);
or OR3 (N938, N930, N52, N71);
or OR3 (N939, N919, N556, N720);
buf BUF1 (N940, N917);
nor NOR3 (N941, N925, N824, N239);
and AND3 (N942, N929, N200, N448);
and AND2 (N943, N936, N255);
or OR4 (N944, N943, N293, N600, N608);
nor NOR3 (N945, N941, N72, N903);
buf BUF1 (N946, N945);
and AND3 (N947, N939, N46, N249);
nor NOR3 (N948, N937, N555, N399);
xor XOR2 (N949, N944, N837);
not NOT1 (N950, N948);
xor XOR2 (N951, N947, N701);
nor NOR4 (N952, N951, N343, N629, N263);
xor XOR2 (N953, N928, N590);
buf BUF1 (N954, N932);
and AND4 (N955, N934, N96, N901, N400);
nand NAND3 (N956, N954, N414, N142);
not NOT1 (N957, N938);
nor NOR4 (N958, N942, N790, N117, N794);
nand NAND3 (N959, N949, N885, N716);
or OR4 (N960, N955, N482, N216, N860);
nor NOR3 (N961, N959, N735, N886);
xor XOR2 (N962, N956, N432);
nor NOR2 (N963, N946, N81);
or OR4 (N964, N962, N798, N396, N5);
and AND2 (N965, N940, N51);
or OR3 (N966, N961, N285, N772);
not NOT1 (N967, N950);
xor XOR2 (N968, N953, N112);
and AND2 (N969, N966, N215);
and AND3 (N970, N967, N917, N76);
nor NOR4 (N971, N968, N804, N565, N60);
or OR3 (N972, N952, N81, N137);
and AND3 (N973, N958, N889, N620);
buf BUF1 (N974, N965);
buf BUF1 (N975, N964);
xor XOR2 (N976, N973, N704);
buf BUF1 (N977, N969);
nand NAND2 (N978, N960, N291);
xor XOR2 (N979, N975, N644);
nand NAND4 (N980, N957, N48, N401, N363);
or OR4 (N981, N977, N769, N628, N745);
nor NOR3 (N982, N980, N74, N557);
nand NAND4 (N983, N976, N77, N57, N784);
buf BUF1 (N984, N982);
nand NAND2 (N985, N981, N8);
and AND4 (N986, N970, N232, N790, N726);
nor NOR4 (N987, N983, N256, N396, N56);
nor NOR4 (N988, N985, N612, N433, N593);
buf BUF1 (N989, N988);
not NOT1 (N990, N987);
buf BUF1 (N991, N974);
buf BUF1 (N992, N984);
buf BUF1 (N993, N989);
nand NAND2 (N994, N990, N19);
buf BUF1 (N995, N994);
and AND4 (N996, N979, N587, N168, N405);
and AND2 (N997, N972, N761);
or OR2 (N998, N986, N377);
and AND2 (N999, N992, N943);
not NOT1 (N1000, N971);
nor NOR4 (N1001, N978, N313, N412, N376);
buf BUF1 (N1002, N991);
nor NOR2 (N1003, N1000, N584);
or OR3 (N1004, N999, N142, N40);
nor NOR3 (N1005, N993, N160, N223);
nor NOR4 (N1006, N998, N626, N986, N577);
and AND3 (N1007, N997, N730, N167);
nand NAND3 (N1008, N1006, N344, N925);
xor XOR2 (N1009, N1004, N45);
nand NAND2 (N1010, N1005, N548);
buf BUF1 (N1011, N1007);
nand NAND3 (N1012, N963, N169, N541);
nor NOR2 (N1013, N1009, N245);
xor XOR2 (N1014, N1012, N671);
xor XOR2 (N1015, N996, N466);
nor NOR4 (N1016, N1010, N898, N751, N558);
not NOT1 (N1017, N1003);
not NOT1 (N1018, N1016);
buf BUF1 (N1019, N1018);
and AND3 (N1020, N1019, N217, N455);
or OR4 (N1021, N1008, N508, N979, N36);
nand NAND3 (N1022, N1021, N855, N441);
nor NOR4 (N1023, N1015, N9, N4, N863);
nor NOR4 (N1024, N1001, N939, N458, N356);
xor XOR2 (N1025, N1022, N907);
or OR3 (N1026, N1002, N703, N799);
or OR2 (N1027, N1014, N202);
nor NOR2 (N1028, N1017, N800);
or OR3 (N1029, N1020, N599, N327);
and AND4 (N1030, N1013, N568, N516, N68);
buf BUF1 (N1031, N1024);
nor NOR2 (N1032, N1028, N923);
nor NOR3 (N1033, N1032, N908, N811);
or OR3 (N1034, N1026, N395, N53);
buf BUF1 (N1035, N1030);
buf BUF1 (N1036, N1025);
and AND2 (N1037, N1031, N673);
not NOT1 (N1038, N1033);
not NOT1 (N1039, N995);
not NOT1 (N1040, N1038);
not NOT1 (N1041, N1034);
nand NAND2 (N1042, N1029, N65);
not NOT1 (N1043, N1027);
or OR2 (N1044, N1023, N764);
or OR4 (N1045, N1041, N10, N221, N522);
or OR3 (N1046, N1036, N993, N70);
and AND3 (N1047, N1045, N412, N400);
nor NOR2 (N1048, N1040, N957);
xor XOR2 (N1049, N1042, N666);
and AND4 (N1050, N1048, N335, N31, N714);
nand NAND4 (N1051, N1035, N397, N469, N757);
nand NAND4 (N1052, N1043, N545, N289, N848);
xor XOR2 (N1053, N1046, N190);
or OR2 (N1054, N1050, N563);
nand NAND3 (N1055, N1052, N222, N61);
or OR2 (N1056, N1049, N137);
buf BUF1 (N1057, N1011);
xor XOR2 (N1058, N1039, N397);
nand NAND3 (N1059, N1037, N367, N901);
and AND2 (N1060, N1051, N739);
not NOT1 (N1061, N1060);
or OR3 (N1062, N1058, N239, N849);
nand NAND3 (N1063, N1057, N434, N929);
or OR3 (N1064, N1056, N18, N155);
buf BUF1 (N1065, N1047);
xor XOR2 (N1066, N1063, N404);
and AND2 (N1067, N1064, N145);
and AND3 (N1068, N1044, N427, N950);
nand NAND3 (N1069, N1065, N203, N657);
or OR2 (N1070, N1061, N401);
or OR4 (N1071, N1055, N189, N199, N898);
not NOT1 (N1072, N1054);
buf BUF1 (N1073, N1069);
or OR4 (N1074, N1053, N879, N795, N1014);
nand NAND4 (N1075, N1068, N618, N570, N222);
or OR2 (N1076, N1072, N483);
xor XOR2 (N1077, N1066, N424);
and AND2 (N1078, N1073, N626);
and AND4 (N1079, N1070, N230, N107, N601);
xor XOR2 (N1080, N1075, N491);
not NOT1 (N1081, N1071);
and AND2 (N1082, N1076, N449);
not NOT1 (N1083, N1059);
or OR4 (N1084, N1079, N257, N880, N360);
not NOT1 (N1085, N1062);
or OR3 (N1086, N1084, N223, N95);
or OR2 (N1087, N1080, N240);
not NOT1 (N1088, N1078);
or OR3 (N1089, N1083, N480, N665);
and AND3 (N1090, N1088, N18, N336);
nand NAND2 (N1091, N1090, N82);
not NOT1 (N1092, N1074);
buf BUF1 (N1093, N1091);
nand NAND3 (N1094, N1085, N916, N125);
not NOT1 (N1095, N1082);
nand NAND3 (N1096, N1086, N1051, N346);
buf BUF1 (N1097, N1089);
nor NOR2 (N1098, N1095, N717);
buf BUF1 (N1099, N1097);
xor XOR2 (N1100, N1099, N483);
nand NAND2 (N1101, N1092, N543);
nand NAND3 (N1102, N1100, N1049, N196);
nor NOR2 (N1103, N1094, N639);
nand NAND3 (N1104, N1096, N875, N620);
nor NOR2 (N1105, N1103, N801);
buf BUF1 (N1106, N1098);
buf BUF1 (N1107, N1101);
buf BUF1 (N1108, N1105);
or OR3 (N1109, N1102, N737, N543);
xor XOR2 (N1110, N1087, N404);
and AND4 (N1111, N1104, N1058, N142, N635);
xor XOR2 (N1112, N1109, N491);
nand NAND2 (N1113, N1112, N1079);
and AND3 (N1114, N1067, N866, N769);
xor XOR2 (N1115, N1113, N221);
nor NOR2 (N1116, N1110, N373);
or OR2 (N1117, N1111, N1112);
or OR3 (N1118, N1107, N499, N223);
nor NOR2 (N1119, N1114, N344);
nand NAND2 (N1120, N1119, N176);
xor XOR2 (N1121, N1117, N167);
nand NAND3 (N1122, N1116, N801, N921);
xor XOR2 (N1123, N1106, N163);
xor XOR2 (N1124, N1093, N378);
or OR2 (N1125, N1115, N807);
nor NOR4 (N1126, N1121, N872, N531, N339);
not NOT1 (N1127, N1126);
xor XOR2 (N1128, N1081, N501);
xor XOR2 (N1129, N1127, N372);
or OR2 (N1130, N1120, N898);
nand NAND3 (N1131, N1122, N900, N76);
and AND4 (N1132, N1125, N523, N430, N1031);
and AND2 (N1133, N1132, N1058);
buf BUF1 (N1134, N1131);
nor NOR2 (N1135, N1077, N509);
xor XOR2 (N1136, N1130, N281);
or OR2 (N1137, N1135, N275);
xor XOR2 (N1138, N1108, N269);
nor NOR2 (N1139, N1123, N1005);
xor XOR2 (N1140, N1137, N503);
or OR4 (N1141, N1140, N40, N297, N248);
xor XOR2 (N1142, N1133, N775);
nand NAND2 (N1143, N1141, N203);
xor XOR2 (N1144, N1139, N565);
or OR3 (N1145, N1142, N631, N611);
xor XOR2 (N1146, N1138, N989);
or OR4 (N1147, N1124, N668, N558, N528);
nor NOR4 (N1148, N1146, N1026, N945, N751);
not NOT1 (N1149, N1143);
or OR2 (N1150, N1134, N106);
nand NAND4 (N1151, N1118, N1037, N103, N876);
not NOT1 (N1152, N1129);
nor NOR3 (N1153, N1128, N771, N860);
buf BUF1 (N1154, N1151);
and AND3 (N1155, N1150, N474, N944);
nor NOR3 (N1156, N1154, N495, N873);
nor NOR4 (N1157, N1136, N244, N750, N690);
or OR4 (N1158, N1148, N959, N700, N946);
xor XOR2 (N1159, N1158, N773);
and AND2 (N1160, N1147, N928);
xor XOR2 (N1161, N1145, N891);
nand NAND3 (N1162, N1155, N755, N857);
buf BUF1 (N1163, N1153);
not NOT1 (N1164, N1160);
and AND3 (N1165, N1162, N746, N860);
or OR2 (N1166, N1159, N519);
or OR4 (N1167, N1166, N86, N1133, N587);
not NOT1 (N1168, N1149);
buf BUF1 (N1169, N1144);
buf BUF1 (N1170, N1167);
nand NAND3 (N1171, N1163, N351, N21);
not NOT1 (N1172, N1169);
nand NAND3 (N1173, N1164, N43, N735);
or OR4 (N1174, N1157, N316, N382, N303);
not NOT1 (N1175, N1172);
buf BUF1 (N1176, N1156);
or OR4 (N1177, N1171, N999, N1161, N287);
xor XOR2 (N1178, N160, N983);
not NOT1 (N1179, N1173);
nand NAND3 (N1180, N1175, N6, N315);
nand NAND3 (N1181, N1180, N96, N550);
or OR3 (N1182, N1178, N243, N295);
nand NAND2 (N1183, N1182, N740);
xor XOR2 (N1184, N1165, N469);
and AND2 (N1185, N1168, N75);
and AND2 (N1186, N1183, N660);
buf BUF1 (N1187, N1181);
or OR3 (N1188, N1184, N418, N202);
buf BUF1 (N1189, N1177);
or OR3 (N1190, N1170, N801, N763);
xor XOR2 (N1191, N1152, N578);
nor NOR4 (N1192, N1189, N224, N122, N478);
nand NAND3 (N1193, N1179, N664, N319);
buf BUF1 (N1194, N1176);
buf BUF1 (N1195, N1185);
nand NAND2 (N1196, N1186, N1039);
and AND2 (N1197, N1192, N48);
xor XOR2 (N1198, N1197, N1080);
or OR4 (N1199, N1174, N578, N310, N521);
nor NOR4 (N1200, N1199, N1118, N1050, N375);
or OR3 (N1201, N1188, N980, N298);
nand NAND3 (N1202, N1193, N741, N1087);
or OR3 (N1203, N1187, N638, N1077);
xor XOR2 (N1204, N1201, N408);
xor XOR2 (N1205, N1200, N842);
nand NAND2 (N1206, N1196, N540);
xor XOR2 (N1207, N1206, N1102);
not NOT1 (N1208, N1191);
and AND4 (N1209, N1207, N1020, N517, N371);
not NOT1 (N1210, N1208);
nor NOR2 (N1211, N1194, N831);
or OR2 (N1212, N1198, N390);
buf BUF1 (N1213, N1212);
not NOT1 (N1214, N1211);
not NOT1 (N1215, N1190);
nor NOR3 (N1216, N1205, N1063, N180);
nand NAND2 (N1217, N1216, N782);
buf BUF1 (N1218, N1214);
nor NOR4 (N1219, N1195, N636, N381, N928);
buf BUF1 (N1220, N1213);
not NOT1 (N1221, N1209);
or OR3 (N1222, N1218, N22, N563);
nor NOR2 (N1223, N1204, N1179);
and AND2 (N1224, N1210, N153);
not NOT1 (N1225, N1223);
nand NAND4 (N1226, N1220, N103, N736, N1163);
and AND2 (N1227, N1222, N553);
and AND2 (N1228, N1215, N728);
buf BUF1 (N1229, N1217);
not NOT1 (N1230, N1226);
or OR2 (N1231, N1228, N147);
nand NAND2 (N1232, N1224, N1108);
nor NOR2 (N1233, N1221, N802);
nor NOR2 (N1234, N1230, N1143);
not NOT1 (N1235, N1229);
xor XOR2 (N1236, N1203, N146);
nor NOR2 (N1237, N1233, N545);
buf BUF1 (N1238, N1232);
not NOT1 (N1239, N1219);
or OR3 (N1240, N1227, N1142, N955);
nand NAND4 (N1241, N1235, N1013, N398, N922);
or OR2 (N1242, N1239, N1159);
not NOT1 (N1243, N1202);
buf BUF1 (N1244, N1231);
and AND4 (N1245, N1242, N110, N1233, N715);
not NOT1 (N1246, N1245);
nand NAND4 (N1247, N1238, N506, N504, N1112);
buf BUF1 (N1248, N1247);
or OR3 (N1249, N1243, N808, N999);
nor NOR3 (N1250, N1246, N273, N968);
not NOT1 (N1251, N1237);
nor NOR2 (N1252, N1249, N336);
nor NOR4 (N1253, N1251, N1057, N763, N985);
not NOT1 (N1254, N1241);
not NOT1 (N1255, N1248);
nor NOR4 (N1256, N1225, N690, N1038, N790);
nor NOR3 (N1257, N1252, N560, N389);
not NOT1 (N1258, N1236);
not NOT1 (N1259, N1253);
or OR2 (N1260, N1250, N456);
xor XOR2 (N1261, N1254, N346);
or OR2 (N1262, N1258, N419);
nand NAND4 (N1263, N1256, N1069, N1150, N724);
nor NOR3 (N1264, N1255, N91, N938);
xor XOR2 (N1265, N1264, N919);
and AND4 (N1266, N1240, N961, N317, N414);
not NOT1 (N1267, N1265);
buf BUF1 (N1268, N1259);
buf BUF1 (N1269, N1261);
not NOT1 (N1270, N1268);
buf BUF1 (N1271, N1266);
and AND2 (N1272, N1257, N720);
xor XOR2 (N1273, N1263, N373);
nand NAND4 (N1274, N1244, N1006, N71, N225);
nand NAND4 (N1275, N1273, N672, N71, N1069);
and AND2 (N1276, N1271, N909);
nand NAND3 (N1277, N1270, N68, N700);
xor XOR2 (N1278, N1274, N655);
and AND4 (N1279, N1267, N249, N44, N211);
buf BUF1 (N1280, N1277);
nand NAND3 (N1281, N1278, N283, N958);
or OR4 (N1282, N1262, N169, N574, N413);
or OR2 (N1283, N1234, N348);
xor XOR2 (N1284, N1276, N1202);
xor XOR2 (N1285, N1283, N234);
and AND3 (N1286, N1279, N523, N292);
xor XOR2 (N1287, N1272, N954);
not NOT1 (N1288, N1275);
not NOT1 (N1289, N1280);
not NOT1 (N1290, N1285);
xor XOR2 (N1291, N1269, N94);
xor XOR2 (N1292, N1281, N1046);
buf BUF1 (N1293, N1282);
and AND2 (N1294, N1289, N896);
not NOT1 (N1295, N1287);
nor NOR4 (N1296, N1293, N1157, N1239, N766);
nand NAND2 (N1297, N1260, N5);
not NOT1 (N1298, N1286);
buf BUF1 (N1299, N1284);
buf BUF1 (N1300, N1292);
and AND3 (N1301, N1290, N181, N612);
nand NAND2 (N1302, N1295, N255);
buf BUF1 (N1303, N1300);
xor XOR2 (N1304, N1302, N801);
buf BUF1 (N1305, N1303);
nor NOR2 (N1306, N1304, N811);
buf BUF1 (N1307, N1301);
xor XOR2 (N1308, N1299, N527);
nand NAND3 (N1309, N1298, N1124, N833);
nand NAND2 (N1310, N1294, N307);
nor NOR3 (N1311, N1307, N814, N1075);
not NOT1 (N1312, N1308);
not NOT1 (N1313, N1306);
nor NOR3 (N1314, N1291, N870, N1043);
not NOT1 (N1315, N1309);
and AND4 (N1316, N1313, N695, N904, N770);
xor XOR2 (N1317, N1305, N30);
buf BUF1 (N1318, N1316);
and AND3 (N1319, N1311, N123, N122);
xor XOR2 (N1320, N1312, N495);
and AND4 (N1321, N1314, N1172, N711, N327);
nor NOR2 (N1322, N1288, N154);
xor XOR2 (N1323, N1310, N647);
and AND3 (N1324, N1322, N70, N128);
buf BUF1 (N1325, N1296);
nor NOR2 (N1326, N1323, N614);
not NOT1 (N1327, N1319);
and AND3 (N1328, N1297, N1048, N1305);
nor NOR2 (N1329, N1325, N997);
nand NAND4 (N1330, N1326, N342, N148, N637);
xor XOR2 (N1331, N1327, N138);
or OR2 (N1332, N1328, N268);
nor NOR2 (N1333, N1318, N1240);
buf BUF1 (N1334, N1332);
buf BUF1 (N1335, N1331);
buf BUF1 (N1336, N1335);
and AND2 (N1337, N1315, N688);
and AND4 (N1338, N1334, N939, N781, N776);
or OR4 (N1339, N1329, N1195, N474, N4);
or OR2 (N1340, N1338, N1219);
not NOT1 (N1341, N1324);
buf BUF1 (N1342, N1341);
and AND3 (N1343, N1339, N1247, N1172);
not NOT1 (N1344, N1336);
nor NOR2 (N1345, N1320, N1165);
nand NAND3 (N1346, N1333, N294, N266);
xor XOR2 (N1347, N1340, N1242);
not NOT1 (N1348, N1321);
nor NOR4 (N1349, N1342, N473, N1231, N655);
buf BUF1 (N1350, N1349);
buf BUF1 (N1351, N1350);
and AND4 (N1352, N1347, N887, N1287, N1257);
and AND4 (N1353, N1348, N1171, N15, N388);
nor NOR2 (N1354, N1337, N213);
and AND3 (N1355, N1353, N1286, N649);
not NOT1 (N1356, N1346);
or OR4 (N1357, N1345, N451, N636, N332);
buf BUF1 (N1358, N1351);
not NOT1 (N1359, N1344);
nand NAND2 (N1360, N1354, N792);
xor XOR2 (N1361, N1343, N1261);
nand NAND3 (N1362, N1360, N579, N1066);
nand NAND2 (N1363, N1361, N207);
nand NAND4 (N1364, N1362, N529, N263, N780);
buf BUF1 (N1365, N1359);
nand NAND3 (N1366, N1356, N240, N462);
buf BUF1 (N1367, N1330);
xor XOR2 (N1368, N1364, N902);
or OR2 (N1369, N1357, N1194);
xor XOR2 (N1370, N1365, N1347);
nor NOR4 (N1371, N1366, N1241, N464, N570);
and AND3 (N1372, N1352, N10, N1208);
xor XOR2 (N1373, N1355, N1363);
buf BUF1 (N1374, N133);
nand NAND4 (N1375, N1371, N646, N1133, N1076);
nand NAND3 (N1376, N1374, N748, N552);
or OR2 (N1377, N1370, N1008);
nand NAND4 (N1378, N1369, N334, N1167, N473);
nand NAND2 (N1379, N1376, N11);
not NOT1 (N1380, N1378);
buf BUF1 (N1381, N1367);
nand NAND4 (N1382, N1372, N207, N145, N273);
nor NOR2 (N1383, N1317, N514);
xor XOR2 (N1384, N1368, N226);
xor XOR2 (N1385, N1382, N862);
xor XOR2 (N1386, N1358, N129);
and AND3 (N1387, N1377, N1317, N895);
not NOT1 (N1388, N1383);
and AND4 (N1389, N1375, N8, N1164, N836);
nor NOR3 (N1390, N1379, N550, N346);
nor NOR3 (N1391, N1380, N1244, N576);
or OR2 (N1392, N1388, N624);
nand NAND4 (N1393, N1385, N4, N77, N760);
nor NOR3 (N1394, N1391, N832, N264);
nor NOR2 (N1395, N1390, N807);
and AND4 (N1396, N1392, N953, N890, N193);
not NOT1 (N1397, N1373);
not NOT1 (N1398, N1381);
xor XOR2 (N1399, N1396, N52);
nand NAND3 (N1400, N1398, N313, N6);
and AND4 (N1401, N1393, N616, N125, N930);
buf BUF1 (N1402, N1400);
not NOT1 (N1403, N1384);
xor XOR2 (N1404, N1402, N1120);
nor NOR3 (N1405, N1399, N108, N740);
buf BUF1 (N1406, N1386);
or OR2 (N1407, N1406, N720);
not NOT1 (N1408, N1389);
buf BUF1 (N1409, N1401);
or OR4 (N1410, N1408, N577, N440, N950);
not NOT1 (N1411, N1410);
or OR3 (N1412, N1394, N42, N1040);
nand NAND4 (N1413, N1407, N623, N131, N130);
buf BUF1 (N1414, N1403);
or OR4 (N1415, N1395, N891, N1275, N178);
buf BUF1 (N1416, N1409);
buf BUF1 (N1417, N1416);
and AND4 (N1418, N1417, N805, N1049, N1092);
or OR4 (N1419, N1404, N71, N789, N484);
nor NOR2 (N1420, N1412, N579);
buf BUF1 (N1421, N1415);
not NOT1 (N1422, N1397);
and AND2 (N1423, N1387, N990);
xor XOR2 (N1424, N1421, N640);
or OR4 (N1425, N1414, N1183, N850, N1204);
or OR4 (N1426, N1419, N354, N1167, N796);
buf BUF1 (N1427, N1426);
and AND2 (N1428, N1418, N1257);
buf BUF1 (N1429, N1428);
not NOT1 (N1430, N1411);
and AND4 (N1431, N1429, N436, N1159, N330);
buf BUF1 (N1432, N1431);
or OR3 (N1433, N1405, N373, N842);
or OR4 (N1434, N1425, N126, N1382, N1389);
not NOT1 (N1435, N1430);
xor XOR2 (N1436, N1435, N782);
nor NOR2 (N1437, N1423, N798);
and AND4 (N1438, N1434, N803, N336, N1344);
xor XOR2 (N1439, N1437, N934);
nor NOR3 (N1440, N1438, N1430, N175);
xor XOR2 (N1441, N1436, N808);
nand NAND2 (N1442, N1427, N1122);
buf BUF1 (N1443, N1432);
buf BUF1 (N1444, N1422);
xor XOR2 (N1445, N1443, N735);
not NOT1 (N1446, N1442);
or OR3 (N1447, N1445, N439, N557);
or OR3 (N1448, N1446, N1032, N310);
buf BUF1 (N1449, N1413);
nor NOR2 (N1450, N1449, N130);
nand NAND3 (N1451, N1433, N850, N665);
or OR4 (N1452, N1451, N317, N650, N588);
or OR3 (N1453, N1448, N1295, N682);
xor XOR2 (N1454, N1440, N481);
buf BUF1 (N1455, N1452);
and AND4 (N1456, N1439, N1086, N547, N255);
not NOT1 (N1457, N1424);
nor NOR3 (N1458, N1457, N502, N860);
buf BUF1 (N1459, N1458);
xor XOR2 (N1460, N1455, N415);
buf BUF1 (N1461, N1456);
nor NOR3 (N1462, N1461, N220, N1005);
nand NAND2 (N1463, N1441, N715);
xor XOR2 (N1464, N1453, N416);
buf BUF1 (N1465, N1420);
nor NOR4 (N1466, N1462, N887, N166, N1134);
or OR3 (N1467, N1454, N1415, N416);
or OR3 (N1468, N1465, N609, N460);
buf BUF1 (N1469, N1466);
or OR3 (N1470, N1450, N835, N535);
not NOT1 (N1471, N1468);
xor XOR2 (N1472, N1467, N192);
nor NOR4 (N1473, N1470, N145, N69, N703);
and AND4 (N1474, N1444, N1380, N101, N827);
not NOT1 (N1475, N1463);
not NOT1 (N1476, N1475);
nand NAND3 (N1477, N1472, N205, N419);
or OR4 (N1478, N1447, N596, N83, N747);
not NOT1 (N1479, N1477);
nand NAND2 (N1480, N1464, N552);
nand NAND4 (N1481, N1476, N1406, N194, N195);
xor XOR2 (N1482, N1459, N79);
and AND2 (N1483, N1471, N929);
nor NOR4 (N1484, N1474, N1409, N496, N244);
and AND4 (N1485, N1479, N1029, N1115, N1003);
not NOT1 (N1486, N1478);
or OR2 (N1487, N1469, N1454);
nand NAND4 (N1488, N1487, N322, N1432, N1175);
not NOT1 (N1489, N1486);
nand NAND2 (N1490, N1483, N1198);
buf BUF1 (N1491, N1489);
not NOT1 (N1492, N1491);
and AND3 (N1493, N1490, N105, N11);
not NOT1 (N1494, N1488);
buf BUF1 (N1495, N1492);
not NOT1 (N1496, N1482);
not NOT1 (N1497, N1494);
not NOT1 (N1498, N1481);
not NOT1 (N1499, N1484);
and AND3 (N1500, N1496, N1470, N1332);
buf BUF1 (N1501, N1485);
or OR4 (N1502, N1495, N292, N1207, N599);
xor XOR2 (N1503, N1473, N726);
and AND2 (N1504, N1480, N906);
or OR3 (N1505, N1493, N554, N1235);
nand NAND2 (N1506, N1500, N108);
nor NOR3 (N1507, N1502, N221, N1495);
nand NAND4 (N1508, N1504, N263, N216, N1387);
and AND2 (N1509, N1507, N211);
nor NOR2 (N1510, N1499, N87);
buf BUF1 (N1511, N1460);
nor NOR3 (N1512, N1511, N288, N1333);
nand NAND2 (N1513, N1512, N1493);
not NOT1 (N1514, N1503);
nor NOR4 (N1515, N1513, N220, N381, N141);
and AND2 (N1516, N1501, N706);
not NOT1 (N1517, N1508);
not NOT1 (N1518, N1498);
xor XOR2 (N1519, N1514, N745);
nor NOR3 (N1520, N1510, N98, N1351);
and AND4 (N1521, N1497, N725, N536, N1012);
buf BUF1 (N1522, N1518);
not NOT1 (N1523, N1515);
not NOT1 (N1524, N1521);
nand NAND4 (N1525, N1506, N1088, N239, N714);
or OR4 (N1526, N1505, N1465, N5, N1422);
nor NOR2 (N1527, N1509, N951);
nand NAND2 (N1528, N1522, N1181);
not NOT1 (N1529, N1524);
buf BUF1 (N1530, N1529);
nor NOR2 (N1531, N1527, N1096);
not NOT1 (N1532, N1526);
nor NOR3 (N1533, N1531, N680, N849);
and AND2 (N1534, N1530, N251);
nor NOR3 (N1535, N1534, N481, N388);
not NOT1 (N1536, N1517);
xor XOR2 (N1537, N1520, N1034);
nor NOR3 (N1538, N1532, N1326, N931);
buf BUF1 (N1539, N1535);
not NOT1 (N1540, N1538);
xor XOR2 (N1541, N1523, N960);
or OR4 (N1542, N1541, N776, N767, N827);
buf BUF1 (N1543, N1516);
and AND4 (N1544, N1537, N1515, N182, N1061);
xor XOR2 (N1545, N1543, N621);
xor XOR2 (N1546, N1544, N340);
or OR3 (N1547, N1525, N1000, N868);
and AND3 (N1548, N1528, N204, N1460);
or OR2 (N1549, N1547, N123);
or OR3 (N1550, N1519, N446, N575);
and AND2 (N1551, N1533, N1534);
and AND2 (N1552, N1548, N231);
not NOT1 (N1553, N1546);
nor NOR4 (N1554, N1545, N1248, N30, N1437);
nor NOR3 (N1555, N1553, N185, N776);
and AND4 (N1556, N1551, N1550, N281, N1207);
and AND2 (N1557, N82, N69);
and AND3 (N1558, N1542, N525, N259);
and AND3 (N1559, N1555, N798, N1480);
nor NOR3 (N1560, N1558, N1160, N251);
nand NAND4 (N1561, N1540, N816, N1327, N886);
or OR3 (N1562, N1559, N1018, N529);
xor XOR2 (N1563, N1552, N852);
nand NAND3 (N1564, N1539, N1378, N1109);
xor XOR2 (N1565, N1536, N1546);
xor XOR2 (N1566, N1563, N1126);
nand NAND3 (N1567, N1554, N933, N298);
not NOT1 (N1568, N1566);
nand NAND4 (N1569, N1567, N374, N12, N17);
buf BUF1 (N1570, N1560);
nor NOR4 (N1571, N1568, N1056, N1438, N1372);
xor XOR2 (N1572, N1549, N949);
xor XOR2 (N1573, N1564, N939);
xor XOR2 (N1574, N1573, N197);
xor XOR2 (N1575, N1556, N1169);
or OR2 (N1576, N1575, N1189);
not NOT1 (N1577, N1561);
buf BUF1 (N1578, N1557);
or OR2 (N1579, N1576, N402);
nand NAND3 (N1580, N1574, N895, N756);
not NOT1 (N1581, N1580);
nor NOR4 (N1582, N1577, N1161, N541, N400);
buf BUF1 (N1583, N1570);
buf BUF1 (N1584, N1562);
and AND3 (N1585, N1584, N340, N949);
and AND4 (N1586, N1572, N1097, N160, N1485);
or OR2 (N1587, N1585, N1028);
nor NOR2 (N1588, N1565, N1533);
not NOT1 (N1589, N1581);
nor NOR3 (N1590, N1578, N220, N1558);
or OR2 (N1591, N1569, N303);
nand NAND2 (N1592, N1589, N266);
nand NAND4 (N1593, N1586, N957, N183, N1422);
and AND4 (N1594, N1571, N658, N24, N1077);
nor NOR2 (N1595, N1587, N191);
and AND3 (N1596, N1583, N608, N887);
nor NOR3 (N1597, N1595, N488, N1283);
nor NOR2 (N1598, N1588, N270);
not NOT1 (N1599, N1596);
or OR2 (N1600, N1590, N519);
xor XOR2 (N1601, N1591, N213);
and AND3 (N1602, N1594, N916, N278);
not NOT1 (N1603, N1598);
not NOT1 (N1604, N1582);
nor NOR4 (N1605, N1579, N1300, N148, N726);
and AND4 (N1606, N1604, N1032, N1314, N191);
or OR4 (N1607, N1605, N58, N361, N61);
buf BUF1 (N1608, N1593);
buf BUF1 (N1609, N1602);
nor NOR4 (N1610, N1603, N778, N1243, N543);
and AND3 (N1611, N1609, N304, N1192);
not NOT1 (N1612, N1610);
nor NOR4 (N1613, N1592, N579, N175, N299);
buf BUF1 (N1614, N1611);
not NOT1 (N1615, N1600);
nand NAND3 (N1616, N1601, N519, N1492);
and AND4 (N1617, N1614, N956, N363, N1122);
xor XOR2 (N1618, N1597, N1485);
nor NOR3 (N1619, N1612, N1431, N519);
nand NAND3 (N1620, N1606, N900, N723);
nand NAND3 (N1621, N1608, N991, N725);
or OR4 (N1622, N1619, N570, N1268, N1037);
buf BUF1 (N1623, N1615);
xor XOR2 (N1624, N1622, N679);
or OR2 (N1625, N1623, N573);
and AND4 (N1626, N1613, N971, N239, N1468);
or OR2 (N1627, N1617, N946);
and AND3 (N1628, N1618, N1239, N590);
xor XOR2 (N1629, N1621, N770);
xor XOR2 (N1630, N1620, N1063);
buf BUF1 (N1631, N1628);
buf BUF1 (N1632, N1629);
nand NAND4 (N1633, N1631, N1437, N117, N1303);
nand NAND4 (N1634, N1625, N1335, N1281, N527);
buf BUF1 (N1635, N1624);
buf BUF1 (N1636, N1616);
buf BUF1 (N1637, N1634);
nand NAND4 (N1638, N1627, N834, N1455, N667);
or OR4 (N1639, N1626, N68, N1216, N43);
buf BUF1 (N1640, N1630);
nand NAND3 (N1641, N1640, N175, N268);
nor NOR3 (N1642, N1633, N769, N689);
and AND4 (N1643, N1637, N1449, N724, N469);
nand NAND2 (N1644, N1632, N1148);
and AND2 (N1645, N1599, N781);
not NOT1 (N1646, N1607);
nor NOR3 (N1647, N1644, N674, N1474);
nor NOR2 (N1648, N1647, N1576);
nor NOR4 (N1649, N1642, N790, N613, N1195);
xor XOR2 (N1650, N1636, N780);
xor XOR2 (N1651, N1639, N1458);
buf BUF1 (N1652, N1650);
and AND4 (N1653, N1651, N86, N1493, N822);
nand NAND3 (N1654, N1638, N38, N1368);
or OR4 (N1655, N1649, N352, N715, N1177);
buf BUF1 (N1656, N1652);
and AND4 (N1657, N1656, N522, N388, N88);
buf BUF1 (N1658, N1643);
xor XOR2 (N1659, N1653, N1118);
or OR3 (N1660, N1645, N117, N1005);
xor XOR2 (N1661, N1660, N1086);
not NOT1 (N1662, N1657);
buf BUF1 (N1663, N1635);
xor XOR2 (N1664, N1655, N858);
or OR3 (N1665, N1646, N661, N223);
xor XOR2 (N1666, N1659, N294);
nor NOR3 (N1667, N1641, N1511, N653);
and AND4 (N1668, N1665, N1488, N518, N814);
nand NAND4 (N1669, N1664, N176, N1379, N1463);
nor NOR3 (N1670, N1666, N811, N1006);
or OR2 (N1671, N1667, N615);
nor NOR4 (N1672, N1661, N120, N45, N409);
buf BUF1 (N1673, N1670);
or OR2 (N1674, N1672, N189);
xor XOR2 (N1675, N1663, N619);
nand NAND3 (N1676, N1668, N1121, N1629);
buf BUF1 (N1677, N1669);
buf BUF1 (N1678, N1676);
or OR4 (N1679, N1648, N498, N808, N1497);
nand NAND3 (N1680, N1674, N311, N695);
nand NAND2 (N1681, N1671, N262);
nor NOR2 (N1682, N1680, N1190);
nand NAND2 (N1683, N1678, N1064);
not NOT1 (N1684, N1677);
nor NOR3 (N1685, N1684, N848, N1358);
buf BUF1 (N1686, N1658);
and AND2 (N1687, N1685, N1221);
and AND4 (N1688, N1683, N619, N1219, N813);
and AND3 (N1689, N1654, N42, N747);
buf BUF1 (N1690, N1686);
nand NAND3 (N1691, N1662, N785, N1492);
nor NOR3 (N1692, N1679, N1664, N1072);
buf BUF1 (N1693, N1690);
xor XOR2 (N1694, N1682, N663);
not NOT1 (N1695, N1693);
not NOT1 (N1696, N1691);
not NOT1 (N1697, N1695);
buf BUF1 (N1698, N1694);
or OR2 (N1699, N1698, N877);
nand NAND3 (N1700, N1699, N1667, N1533);
xor XOR2 (N1701, N1688, N328);
buf BUF1 (N1702, N1687);
or OR2 (N1703, N1673, N1477);
and AND3 (N1704, N1703, N1663, N933);
nor NOR3 (N1705, N1697, N390, N1346);
nand NAND2 (N1706, N1705, N483);
nor NOR4 (N1707, N1696, N1547, N1232, N1015);
nor NOR2 (N1708, N1681, N1204);
nand NAND3 (N1709, N1702, N933, N920);
xor XOR2 (N1710, N1700, N1392);
or OR4 (N1711, N1692, N514, N139, N572);
or OR2 (N1712, N1711, N1063);
buf BUF1 (N1713, N1707);
xor XOR2 (N1714, N1708, N47);
or OR4 (N1715, N1704, N335, N544, N1275);
xor XOR2 (N1716, N1709, N84);
and AND3 (N1717, N1713, N1148, N834);
not NOT1 (N1718, N1715);
or OR2 (N1719, N1706, N1217);
and AND4 (N1720, N1712, N4, N446, N795);
buf BUF1 (N1721, N1675);
nor NOR4 (N1722, N1720, N331, N1613, N874);
not NOT1 (N1723, N1710);
buf BUF1 (N1724, N1689);
nor NOR3 (N1725, N1723, N690, N467);
buf BUF1 (N1726, N1719);
not NOT1 (N1727, N1701);
nand NAND2 (N1728, N1727, N950);
buf BUF1 (N1729, N1717);
buf BUF1 (N1730, N1724);
buf BUF1 (N1731, N1726);
buf BUF1 (N1732, N1718);
xor XOR2 (N1733, N1722, N217);
and AND3 (N1734, N1729, N769, N1101);
not NOT1 (N1735, N1725);
or OR2 (N1736, N1730, N136);
nand NAND2 (N1737, N1734, N416);
not NOT1 (N1738, N1721);
or OR3 (N1739, N1735, N991, N1407);
and AND3 (N1740, N1714, N1613, N1674);
nor NOR2 (N1741, N1732, N372);
xor XOR2 (N1742, N1737, N1302);
buf BUF1 (N1743, N1742);
buf BUF1 (N1744, N1716);
or OR4 (N1745, N1741, N1273, N527, N755);
xor XOR2 (N1746, N1739, N1023);
not NOT1 (N1747, N1733);
or OR4 (N1748, N1747, N1742, N918, N571);
not NOT1 (N1749, N1731);
not NOT1 (N1750, N1749);
nand NAND3 (N1751, N1745, N1445, N910);
and AND3 (N1752, N1744, N317, N352);
xor XOR2 (N1753, N1746, N324);
buf BUF1 (N1754, N1750);
and AND3 (N1755, N1753, N133, N977);
nand NAND4 (N1756, N1748, N1253, N1426, N464);
and AND2 (N1757, N1740, N1189);
not NOT1 (N1758, N1757);
and AND4 (N1759, N1754, N458, N1239, N167);
nor NOR3 (N1760, N1738, N1472, N1694);
or OR3 (N1761, N1758, N710, N1330);
nand NAND3 (N1762, N1751, N952, N570);
buf BUF1 (N1763, N1756);
and AND2 (N1764, N1763, N1759);
and AND2 (N1765, N1340, N1598);
and AND4 (N1766, N1765, N1607, N298, N313);
buf BUF1 (N1767, N1755);
and AND2 (N1768, N1761, N1439);
xor XOR2 (N1769, N1760, N9);
nand NAND4 (N1770, N1768, N1652, N267, N21);
or OR2 (N1771, N1752, N1653);
nand NAND2 (N1772, N1766, N196);
and AND4 (N1773, N1736, N1690, N1282, N982);
not NOT1 (N1774, N1769);
nand NAND4 (N1775, N1771, N158, N1027, N1198);
and AND4 (N1776, N1772, N1630, N886, N61);
not NOT1 (N1777, N1774);
buf BUF1 (N1778, N1767);
buf BUF1 (N1779, N1775);
xor XOR2 (N1780, N1779, N1564);
or OR2 (N1781, N1764, N374);
and AND2 (N1782, N1762, N15);
nor NOR3 (N1783, N1780, N795, N1627);
and AND4 (N1784, N1743, N356, N1415, N947);
and AND3 (N1785, N1784, N1170, N431);
buf BUF1 (N1786, N1782);
not NOT1 (N1787, N1781);
buf BUF1 (N1788, N1728);
nand NAND4 (N1789, N1770, N1741, N1047, N109);
or OR4 (N1790, N1787, N1429, N105, N491);
not NOT1 (N1791, N1777);
nand NAND2 (N1792, N1788, N1529);
nand NAND2 (N1793, N1789, N728);
xor XOR2 (N1794, N1785, N289);
or OR4 (N1795, N1792, N371, N679, N704);
nor NOR4 (N1796, N1773, N49, N1272, N1512);
or OR4 (N1797, N1776, N1093, N820, N1081);
buf BUF1 (N1798, N1783);
nor NOR4 (N1799, N1795, N1692, N1434, N96);
or OR4 (N1800, N1794, N558, N1368, N190);
or OR4 (N1801, N1793, N624, N1005, N425);
nand NAND3 (N1802, N1796, N1086, N1637);
nand NAND2 (N1803, N1801, N690);
and AND3 (N1804, N1778, N343, N834);
or OR3 (N1805, N1799, N1110, N1195);
not NOT1 (N1806, N1800);
and AND4 (N1807, N1802, N758, N1096, N1179);
xor XOR2 (N1808, N1804, N1507);
or OR2 (N1809, N1791, N57);
and AND3 (N1810, N1805, N945, N906);
buf BUF1 (N1811, N1807);
not NOT1 (N1812, N1808);
xor XOR2 (N1813, N1803, N605);
and AND3 (N1814, N1809, N1763, N205);
or OR4 (N1815, N1786, N1729, N1480, N1075);
nor NOR3 (N1816, N1814, N1553, N1516);
or OR2 (N1817, N1812, N1370);
or OR2 (N1818, N1811, N1049);
nor NOR3 (N1819, N1790, N1549, N1704);
or OR3 (N1820, N1813, N149, N1442);
and AND2 (N1821, N1815, N379);
or OR2 (N1822, N1816, N259);
nor NOR4 (N1823, N1810, N146, N1572, N755);
and AND3 (N1824, N1798, N1397, N36);
or OR4 (N1825, N1821, N1772, N869, N1652);
nor NOR3 (N1826, N1818, N689, N739);
nand NAND3 (N1827, N1823, N1255, N845);
xor XOR2 (N1828, N1797, N609);
nand NAND2 (N1829, N1820, N23);
and AND4 (N1830, N1817, N1100, N901, N984);
xor XOR2 (N1831, N1819, N1317);
and AND3 (N1832, N1831, N1659, N668);
not NOT1 (N1833, N1830);
and AND4 (N1834, N1828, N424, N101, N1520);
and AND4 (N1835, N1822, N732, N354, N298);
nor NOR3 (N1836, N1806, N1075, N1003);
or OR2 (N1837, N1825, N241);
not NOT1 (N1838, N1826);
and AND4 (N1839, N1834, N16, N119, N1320);
not NOT1 (N1840, N1833);
or OR4 (N1841, N1829, N219, N1462, N1551);
and AND4 (N1842, N1837, N1393, N1370, N319);
or OR3 (N1843, N1840, N1408, N1396);
nor NOR3 (N1844, N1824, N1193, N1246);
xor XOR2 (N1845, N1836, N282);
buf BUF1 (N1846, N1841);
not NOT1 (N1847, N1845);
not NOT1 (N1848, N1842);
not NOT1 (N1849, N1835);
buf BUF1 (N1850, N1839);
buf BUF1 (N1851, N1832);
nor NOR3 (N1852, N1846, N857, N1704);
xor XOR2 (N1853, N1850, N1750);
and AND2 (N1854, N1848, N1017);
not NOT1 (N1855, N1838);
and AND2 (N1856, N1853, N1020);
or OR3 (N1857, N1847, N914, N33);
or OR2 (N1858, N1857, N406);
or OR4 (N1859, N1827, N1095, N719, N769);
buf BUF1 (N1860, N1849);
and AND2 (N1861, N1860, N968);
nand NAND3 (N1862, N1859, N218, N1496);
or OR4 (N1863, N1858, N240, N1118, N769);
and AND3 (N1864, N1862, N582, N393);
not NOT1 (N1865, N1844);
or OR3 (N1866, N1856, N1628, N491);
buf BUF1 (N1867, N1864);
nor NOR4 (N1868, N1863, N692, N1763, N1518);
nor NOR4 (N1869, N1867, N952, N1241, N558);
buf BUF1 (N1870, N1854);
xor XOR2 (N1871, N1861, N1208);
and AND3 (N1872, N1869, N340, N775);
and AND3 (N1873, N1866, N1084, N356);
buf BUF1 (N1874, N1873);
or OR4 (N1875, N1851, N995, N1232, N1642);
nand NAND2 (N1876, N1855, N1516);
nor NOR4 (N1877, N1852, N55, N293, N1600);
and AND4 (N1878, N1865, N923, N187, N667);
nand NAND4 (N1879, N1878, N259, N1624, N107);
or OR2 (N1880, N1879, N1687);
not NOT1 (N1881, N1875);
nor NOR3 (N1882, N1880, N1332, N1049);
nand NAND3 (N1883, N1877, N1460, N1863);
not NOT1 (N1884, N1870);
and AND4 (N1885, N1874, N80, N1348, N1256);
and AND2 (N1886, N1868, N934);
buf BUF1 (N1887, N1885);
nand NAND2 (N1888, N1884, N1261);
not NOT1 (N1889, N1882);
nand NAND4 (N1890, N1876, N268, N1001, N1631);
or OR3 (N1891, N1872, N575, N1328);
and AND3 (N1892, N1887, N1709, N214);
and AND4 (N1893, N1883, N1004, N1672, N256);
and AND2 (N1894, N1893, N1858);
xor XOR2 (N1895, N1894, N1779);
nor NOR2 (N1896, N1843, N486);
nor NOR2 (N1897, N1888, N262);
xor XOR2 (N1898, N1892, N1248);
and AND4 (N1899, N1895, N346, N1627, N313);
nor NOR2 (N1900, N1890, N490);
nor NOR4 (N1901, N1897, N223, N1813, N457);
and AND3 (N1902, N1901, N43, N51);
nor NOR4 (N1903, N1896, N1381, N490, N852);
not NOT1 (N1904, N1871);
buf BUF1 (N1905, N1889);
nand NAND3 (N1906, N1900, N1309, N747);
and AND2 (N1907, N1905, N1818);
not NOT1 (N1908, N1903);
not NOT1 (N1909, N1906);
and AND3 (N1910, N1908, N1193, N525);
buf BUF1 (N1911, N1904);
and AND2 (N1912, N1898, N1608);
or OR2 (N1913, N1907, N349);
and AND2 (N1914, N1881, N1284);
and AND3 (N1915, N1886, N883, N287);
buf BUF1 (N1916, N1899);
xor XOR2 (N1917, N1914, N238);
or OR2 (N1918, N1911, N435);
not NOT1 (N1919, N1913);
or OR2 (N1920, N1912, N1893);
or OR4 (N1921, N1909, N516, N1337, N19);
xor XOR2 (N1922, N1891, N1889);
buf BUF1 (N1923, N1917);
nor NOR3 (N1924, N1902, N1272, N1851);
nor NOR3 (N1925, N1910, N404, N94);
nand NAND4 (N1926, N1923, N1405, N461, N1275);
buf BUF1 (N1927, N1916);
not NOT1 (N1928, N1925);
nor NOR4 (N1929, N1921, N1790, N1140, N1153);
or OR2 (N1930, N1927, N959);
buf BUF1 (N1931, N1919);
xor XOR2 (N1932, N1915, N1301);
and AND3 (N1933, N1932, N1768, N780);
or OR4 (N1934, N1928, N422, N1368, N169);
xor XOR2 (N1935, N1920, N1190);
and AND3 (N1936, N1930, N197, N1734);
xor XOR2 (N1937, N1918, N1612);
xor XOR2 (N1938, N1936, N49);
nor NOR2 (N1939, N1929, N694);
buf BUF1 (N1940, N1924);
nand NAND3 (N1941, N1937, N1440, N546);
and AND2 (N1942, N1931, N1479);
or OR3 (N1943, N1926, N907, N794);
or OR4 (N1944, N1933, N489, N1834, N262);
or OR3 (N1945, N1942, N489, N985);
and AND2 (N1946, N1945, N1513);
or OR4 (N1947, N1944, N1128, N1164, N861);
not NOT1 (N1948, N1935);
and AND4 (N1949, N1943, N755, N1093, N443);
buf BUF1 (N1950, N1947);
xor XOR2 (N1951, N1922, N277);
and AND3 (N1952, N1946, N106, N1138);
not NOT1 (N1953, N1948);
and AND2 (N1954, N1949, N1796);
not NOT1 (N1955, N1950);
nand NAND4 (N1956, N1938, N908, N31, N412);
not NOT1 (N1957, N1953);
not NOT1 (N1958, N1951);
nor NOR2 (N1959, N1957, N1290);
xor XOR2 (N1960, N1954, N1333);
nand NAND3 (N1961, N1940, N1118, N1597);
nand NAND4 (N1962, N1955, N1807, N1579, N312);
or OR2 (N1963, N1960, N1832);
buf BUF1 (N1964, N1941);
and AND4 (N1965, N1963, N1356, N1057, N1951);
not NOT1 (N1966, N1961);
or OR4 (N1967, N1965, N1738, N1913, N6);
and AND2 (N1968, N1967, N1879);
and AND3 (N1969, N1959, N129, N1804);
nand NAND3 (N1970, N1952, N282, N2);
or OR2 (N1971, N1939, N835);
buf BUF1 (N1972, N1966);
and AND4 (N1973, N1964, N1225, N1533, N716);
or OR2 (N1974, N1969, N1112);
nand NAND4 (N1975, N1970, N400, N726, N991);
nand NAND3 (N1976, N1971, N949, N1359);
not NOT1 (N1977, N1975);
and AND4 (N1978, N1958, N585, N1727, N1645);
or OR2 (N1979, N1977, N1659);
buf BUF1 (N1980, N1956);
not NOT1 (N1981, N1972);
or OR2 (N1982, N1934, N532);
nand NAND4 (N1983, N1974, N710, N480, N1563);
nand NAND4 (N1984, N1962, N373, N1004, N332);
xor XOR2 (N1985, N1984, N19);
not NOT1 (N1986, N1985);
not NOT1 (N1987, N1979);
not NOT1 (N1988, N1973);
xor XOR2 (N1989, N1976, N334);
or OR4 (N1990, N1988, N1370, N396, N552);
xor XOR2 (N1991, N1968, N721);
buf BUF1 (N1992, N1986);
or OR2 (N1993, N1980, N1424);
buf BUF1 (N1994, N1989);
nor NOR3 (N1995, N1991, N1791, N1972);
not NOT1 (N1996, N1983);
buf BUF1 (N1997, N1981);
nor NOR4 (N1998, N1993, N704, N1313, N1526);
buf BUF1 (N1999, N1998);
buf BUF1 (N2000, N1996);
nor NOR2 (N2001, N1992, N918);
nor NOR4 (N2002, N1978, N688, N47, N41);
and AND4 (N2003, N1999, N1546, N1263, N1086);
xor XOR2 (N2004, N1994, N116);
nor NOR4 (N2005, N2004, N918, N849, N1407);
not NOT1 (N2006, N2003);
xor XOR2 (N2007, N2005, N1013);
buf BUF1 (N2008, N2007);
and AND4 (N2009, N1995, N1207, N1964, N176);
and AND4 (N2010, N2008, N1752, N1662, N623);
xor XOR2 (N2011, N2009, N185);
xor XOR2 (N2012, N1987, N141);
buf BUF1 (N2013, N2001);
nor NOR3 (N2014, N2002, N1042, N1171);
nand NAND4 (N2015, N2014, N711, N1987, N730);
not NOT1 (N2016, N2011);
or OR2 (N2017, N1982, N1904);
nand NAND2 (N2018, N2000, N715);
xor XOR2 (N2019, N1990, N21);
not NOT1 (N2020, N1997);
or OR4 (N2021, N2018, N1428, N417, N1587);
buf BUF1 (N2022, N2019);
buf BUF1 (N2023, N2006);
or OR4 (N2024, N2012, N1576, N282, N1088);
not NOT1 (N2025, N2023);
or OR2 (N2026, N2017, N216);
and AND3 (N2027, N2015, N1543, N1950);
nor NOR3 (N2028, N2021, N302, N419);
nand NAND4 (N2029, N2020, N179, N1223, N846);
and AND4 (N2030, N2025, N1989, N513, N2018);
nor NOR4 (N2031, N2010, N1441, N1638, N979);
xor XOR2 (N2032, N2027, N630);
and AND4 (N2033, N2028, N895, N271, N1112);
and AND3 (N2034, N2026, N1579, N1891);
or OR2 (N2035, N2031, N1075);
xor XOR2 (N2036, N2029, N737);
buf BUF1 (N2037, N2034);
and AND3 (N2038, N2013, N425, N230);
buf BUF1 (N2039, N2024);
buf BUF1 (N2040, N2032);
nand NAND4 (N2041, N2038, N1588, N1135, N1561);
and AND2 (N2042, N2039, N127);
or OR2 (N2043, N2040, N2040);
and AND2 (N2044, N2022, N717);
nand NAND4 (N2045, N2030, N1101, N1969, N334);
buf BUF1 (N2046, N2016);
or OR4 (N2047, N2033, N1888, N1765, N2036);
nand NAND4 (N2048, N1358, N1841, N397, N119);
nor NOR2 (N2049, N2043, N117);
nand NAND2 (N2050, N2049, N91);
and AND4 (N2051, N2047, N702, N419, N1083);
or OR3 (N2052, N2037, N1123, N1338);
nand NAND3 (N2053, N2046, N158, N1407);
nand NAND3 (N2054, N2035, N1556, N560);
buf BUF1 (N2055, N2044);
nor NOR2 (N2056, N2042, N817);
nand NAND2 (N2057, N2051, N60);
not NOT1 (N2058, N2045);
nand NAND3 (N2059, N2055, N1845, N1739);
or OR2 (N2060, N2056, N1213);
buf BUF1 (N2061, N2054);
buf BUF1 (N2062, N2053);
xor XOR2 (N2063, N2062, N1182);
not NOT1 (N2064, N2063);
or OR2 (N2065, N2057, N487);
nor NOR3 (N2066, N2058, N1284, N71);
nor NOR4 (N2067, N2064, N661, N720, N84);
not NOT1 (N2068, N2061);
buf BUF1 (N2069, N2060);
and AND2 (N2070, N2059, N1544);
buf BUF1 (N2071, N2041);
xor XOR2 (N2072, N2070, N1466);
buf BUF1 (N2073, N2048);
nand NAND2 (N2074, N2050, N514);
nand NAND2 (N2075, N2071, N1404);
nand NAND2 (N2076, N2068, N1729);
xor XOR2 (N2077, N2072, N1402);
not NOT1 (N2078, N2077);
buf BUF1 (N2079, N2073);
nand NAND3 (N2080, N2069, N803, N846);
xor XOR2 (N2081, N2080, N312);
nor NOR3 (N2082, N2081, N1088, N443);
xor XOR2 (N2083, N2074, N881);
or OR2 (N2084, N2082, N1867);
nand NAND2 (N2085, N2083, N1376);
nand NAND2 (N2086, N2084, N946);
and AND3 (N2087, N2079, N617, N1733);
buf BUF1 (N2088, N2066);
not NOT1 (N2089, N2086);
or OR3 (N2090, N2085, N1827, N216);
nor NOR4 (N2091, N2067, N1749, N1743, N89);
or OR4 (N2092, N2075, N820, N347, N1021);
buf BUF1 (N2093, N2091);
not NOT1 (N2094, N2088);
nand NAND2 (N2095, N2093, N1322);
xor XOR2 (N2096, N2065, N1363);
and AND3 (N2097, N2076, N163, N922);
buf BUF1 (N2098, N2094);
nand NAND4 (N2099, N2096, N1003, N1915, N1679);
nand NAND3 (N2100, N2078, N306, N1020);
nand NAND2 (N2101, N2087, N1182);
nor NOR2 (N2102, N2100, N1436);
not NOT1 (N2103, N2102);
nor NOR3 (N2104, N2089, N641, N88);
xor XOR2 (N2105, N2052, N274);
and AND4 (N2106, N2103, N1281, N921, N1126);
not NOT1 (N2107, N2101);
nand NAND4 (N2108, N2107, N1440, N1736, N1605);
nand NAND2 (N2109, N2108, N1107);
xor XOR2 (N2110, N2109, N1937);
nand NAND2 (N2111, N2098, N933);
nand NAND2 (N2112, N2110, N1110);
not NOT1 (N2113, N2111);
not NOT1 (N2114, N2106);
and AND2 (N2115, N2092, N1524);
xor XOR2 (N2116, N2104, N1455);
buf BUF1 (N2117, N2113);
or OR3 (N2118, N2105, N1258, N1559);
and AND2 (N2119, N2112, N1898);
or OR4 (N2120, N2114, N1579, N2039, N1989);
and AND3 (N2121, N2095, N399, N1450);
nor NOR2 (N2122, N2119, N2034);
nand NAND2 (N2123, N2117, N1485);
nor NOR4 (N2124, N2123, N318, N245, N556);
not NOT1 (N2125, N2099);
nor NOR3 (N2126, N2121, N554, N1917);
buf BUF1 (N2127, N2115);
buf BUF1 (N2128, N2118);
nand NAND4 (N2129, N2090, N1593, N1152, N361);
nand NAND4 (N2130, N2125, N1588, N1903, N544);
and AND2 (N2131, N2122, N1556);
nand NAND4 (N2132, N2130, N1361, N1240, N776);
not NOT1 (N2133, N2126);
nor NOR2 (N2134, N2127, N534);
nand NAND4 (N2135, N2131, N1035, N1930, N1023);
nand NAND4 (N2136, N2120, N1895, N1778, N768);
nand NAND2 (N2137, N2128, N144);
nand NAND4 (N2138, N2136, N2055, N49, N660);
not NOT1 (N2139, N2116);
or OR2 (N2140, N2135, N709);
or OR4 (N2141, N2133, N1259, N1964, N1733);
buf BUF1 (N2142, N2129);
not NOT1 (N2143, N2097);
or OR3 (N2144, N2140, N1095, N1358);
xor XOR2 (N2145, N2124, N617);
or OR3 (N2146, N2144, N184, N649);
buf BUF1 (N2147, N2141);
xor XOR2 (N2148, N2139, N366);
or OR3 (N2149, N2132, N892, N1372);
and AND4 (N2150, N2146, N2005, N149, N1585);
nor NOR3 (N2151, N2150, N762, N540);
nand NAND4 (N2152, N2138, N1420, N219, N940);
xor XOR2 (N2153, N2143, N1038);
nor NOR3 (N2154, N2152, N94, N1417);
buf BUF1 (N2155, N2134);
or OR2 (N2156, N2137, N1985);
not NOT1 (N2157, N2151);
nand NAND3 (N2158, N2154, N1730, N1656);
buf BUF1 (N2159, N2153);
not NOT1 (N2160, N2155);
and AND3 (N2161, N2145, N637, N1163);
xor XOR2 (N2162, N2158, N734);
nand NAND4 (N2163, N2148, N646, N2072, N1739);
nand NAND3 (N2164, N2161, N1764, N1558);
or OR4 (N2165, N2159, N135, N835, N2149);
nor NOR3 (N2166, N951, N1118, N1218);
not NOT1 (N2167, N2157);
and AND4 (N2168, N2167, N103, N1711, N1101);
xor XOR2 (N2169, N2156, N256);
buf BUF1 (N2170, N2147);
nor NOR4 (N2171, N2170, N2025, N1434, N613);
not NOT1 (N2172, N2165);
nand NAND2 (N2173, N2162, N1520);
xor XOR2 (N2174, N2164, N2134);
nand NAND2 (N2175, N2142, N1172);
or OR4 (N2176, N2173, N1451, N1501, N284);
xor XOR2 (N2177, N2160, N1309);
xor XOR2 (N2178, N2169, N1377);
or OR3 (N2179, N2174, N806, N1013);
and AND4 (N2180, N2168, N442, N1716, N224);
nor NOR3 (N2181, N2175, N985, N777);
nor NOR4 (N2182, N2181, N786, N217, N301);
and AND2 (N2183, N2177, N1625);
or OR3 (N2184, N2178, N1444, N2121);
buf BUF1 (N2185, N2179);
not NOT1 (N2186, N2171);
nor NOR4 (N2187, N2182, N1860, N2022, N580);
nor NOR4 (N2188, N2166, N119, N1562, N1074);
buf BUF1 (N2189, N2186);
and AND2 (N2190, N2188, N1240);
or OR4 (N2191, N2163, N1384, N1762, N836);
xor XOR2 (N2192, N2180, N713);
nor NOR4 (N2193, N2185, N1027, N10, N1191);
or OR4 (N2194, N2190, N208, N853, N1398);
xor XOR2 (N2195, N2187, N355);
xor XOR2 (N2196, N2192, N654);
or OR3 (N2197, N2172, N500, N491);
xor XOR2 (N2198, N2195, N2047);
buf BUF1 (N2199, N2197);
and AND2 (N2200, N2194, N953);
and AND2 (N2201, N2196, N619);
xor XOR2 (N2202, N2198, N929);
and AND3 (N2203, N2189, N1656, N1736);
and AND4 (N2204, N2203, N1101, N2104, N1606);
nand NAND2 (N2205, N2184, N1093);
not NOT1 (N2206, N2191);
nand NAND3 (N2207, N2193, N1325, N769);
or OR3 (N2208, N2199, N357, N128);
nand NAND3 (N2209, N2207, N217, N996);
nor NOR2 (N2210, N2206, N1024);
or OR4 (N2211, N2205, N1459, N1867, N1995);
not NOT1 (N2212, N2210);
or OR3 (N2213, N2209, N1161, N1079);
buf BUF1 (N2214, N2176);
or OR4 (N2215, N2183, N284, N1384, N256);
nor NOR4 (N2216, N2211, N1159, N1218, N2037);
or OR3 (N2217, N2202, N1701, N957);
buf BUF1 (N2218, N2216);
or OR4 (N2219, N2214, N1792, N475, N646);
and AND3 (N2220, N2213, N1543, N709);
not NOT1 (N2221, N2200);
buf BUF1 (N2222, N2215);
buf BUF1 (N2223, N2201);
nor NOR4 (N2224, N2217, N647, N250, N558);
xor XOR2 (N2225, N2218, N2224);
not NOT1 (N2226, N1178);
and AND2 (N2227, N2223, N281);
not NOT1 (N2228, N2212);
nand NAND2 (N2229, N2225, N2120);
xor XOR2 (N2230, N2228, N184);
or OR2 (N2231, N2219, N191);
not NOT1 (N2232, N2231);
or OR3 (N2233, N2230, N856, N354);
or OR4 (N2234, N2204, N428, N1264, N1731);
nor NOR4 (N2235, N2208, N465, N1864, N846);
xor XOR2 (N2236, N2234, N1957);
buf BUF1 (N2237, N2232);
nand NAND4 (N2238, N2235, N2206, N1045, N1314);
or OR4 (N2239, N2237, N1115, N244, N814);
buf BUF1 (N2240, N2239);
or OR3 (N2241, N2220, N1471, N2063);
not NOT1 (N2242, N2238);
and AND4 (N2243, N2236, N1083, N2088, N541);
nor NOR2 (N2244, N2243, N1655);
and AND4 (N2245, N2240, N1783, N1429, N342);
buf BUF1 (N2246, N2229);
or OR2 (N2247, N2233, N1346);
and AND3 (N2248, N2242, N251, N639);
or OR2 (N2249, N2227, N591);
or OR4 (N2250, N2226, N1418, N119, N2040);
not NOT1 (N2251, N2241);
xor XOR2 (N2252, N2245, N1709);
nand NAND2 (N2253, N2244, N592);
or OR2 (N2254, N2250, N654);
nor NOR4 (N2255, N2222, N1095, N1410, N2118);
nor NOR4 (N2256, N2249, N1190, N646, N1001);
nor NOR3 (N2257, N2256, N767, N1985);
buf BUF1 (N2258, N2255);
nor NOR4 (N2259, N2253, N88, N1524, N2106);
buf BUF1 (N2260, N2254);
nand NAND2 (N2261, N2259, N1511);
and AND2 (N2262, N2248, N364);
nand NAND4 (N2263, N2221, N2213, N2088, N1350);
nor NOR2 (N2264, N2247, N1422);
nor NOR2 (N2265, N2246, N1214);
nor NOR4 (N2266, N2263, N1688, N461, N874);
buf BUF1 (N2267, N2251);
xor XOR2 (N2268, N2265, N60);
xor XOR2 (N2269, N2267, N1110);
or OR2 (N2270, N2269, N533);
buf BUF1 (N2271, N2268);
nand NAND2 (N2272, N2261, N551);
nor NOR4 (N2273, N2257, N917, N1381, N1230);
not NOT1 (N2274, N2271);
buf BUF1 (N2275, N2272);
nand NAND3 (N2276, N2275, N626, N1808);
buf BUF1 (N2277, N2270);
or OR3 (N2278, N2260, N152, N1780);
nor NOR3 (N2279, N2278, N1920, N694);
or OR4 (N2280, N2266, N1848, N1537, N1911);
or OR2 (N2281, N2274, N1465);
nand NAND3 (N2282, N2280, N886, N1650);
nor NOR4 (N2283, N2279, N116, N527, N1882);
nand NAND4 (N2284, N2252, N633, N794, N1396);
nor NOR4 (N2285, N2283, N565, N1596, N1761);
and AND2 (N2286, N2258, N2063);
and AND3 (N2287, N2262, N558, N379);
and AND3 (N2288, N2282, N1382, N252);
nor NOR2 (N2289, N2288, N2022);
not NOT1 (N2290, N2286);
nand NAND4 (N2291, N2284, N1551, N184, N163);
and AND2 (N2292, N2273, N1504);
and AND4 (N2293, N2289, N1893, N181, N579);
nor NOR3 (N2294, N2285, N2132, N251);
nor NOR3 (N2295, N2292, N1743, N2173);
or OR4 (N2296, N2287, N269, N2047, N940);
and AND2 (N2297, N2291, N19);
nand NAND3 (N2298, N2276, N2180, N1513);
not NOT1 (N2299, N2296);
xor XOR2 (N2300, N2281, N1368);
nor NOR2 (N2301, N2295, N1171);
buf BUF1 (N2302, N2293);
not NOT1 (N2303, N2301);
or OR2 (N2304, N2297, N584);
nand NAND4 (N2305, N2300, N1936, N809, N981);
not NOT1 (N2306, N2277);
buf BUF1 (N2307, N2294);
buf BUF1 (N2308, N2290);
or OR2 (N2309, N2298, N2183);
or OR4 (N2310, N2304, N1301, N2243, N1180);
nand NAND4 (N2311, N2309, N819, N2078, N2306);
buf BUF1 (N2312, N253);
buf BUF1 (N2313, N2307);
nand NAND2 (N2314, N2311, N1374);
and AND3 (N2315, N2308, N2070, N961);
and AND3 (N2316, N2310, N1670, N1918);
nor NOR4 (N2317, N2302, N332, N131, N1310);
nand NAND3 (N2318, N2303, N90, N741);
and AND2 (N2319, N2317, N1136);
nor NOR4 (N2320, N2312, N421, N84, N200);
nand NAND3 (N2321, N2299, N1051, N1081);
nor NOR3 (N2322, N2319, N1854, N1375);
buf BUF1 (N2323, N2315);
or OR4 (N2324, N2316, N1412, N1074, N407);
xor XOR2 (N2325, N2321, N324);
and AND2 (N2326, N2314, N273);
nor NOR2 (N2327, N2322, N1348);
and AND4 (N2328, N2320, N831, N2119, N1162);
buf BUF1 (N2329, N2325);
or OR4 (N2330, N2264, N898, N643, N1723);
buf BUF1 (N2331, N2313);
and AND2 (N2332, N2305, N509);
nor NOR3 (N2333, N2324, N1103, N408);
buf BUF1 (N2334, N2318);
xor XOR2 (N2335, N2332, N1475);
buf BUF1 (N2336, N2328);
xor XOR2 (N2337, N2323, N2104);
xor XOR2 (N2338, N2331, N743);
or OR4 (N2339, N2335, N240, N427, N179);
not NOT1 (N2340, N2326);
xor XOR2 (N2341, N2334, N1941);
buf BUF1 (N2342, N2333);
and AND4 (N2343, N2330, N569, N2093, N1240);
not NOT1 (N2344, N2329);
buf BUF1 (N2345, N2341);
or OR2 (N2346, N2336, N923);
nand NAND2 (N2347, N2339, N1078);
nand NAND2 (N2348, N2340, N709);
or OR3 (N2349, N2346, N843, N1520);
nand NAND2 (N2350, N2349, N1232);
nand NAND2 (N2351, N2343, N1031);
not NOT1 (N2352, N2344);
nor NOR2 (N2353, N2350, N759);
or OR2 (N2354, N2342, N1068);
not NOT1 (N2355, N2338);
xor XOR2 (N2356, N2345, N289);
or OR2 (N2357, N2353, N1250);
xor XOR2 (N2358, N2352, N546);
or OR3 (N2359, N2354, N662, N827);
not NOT1 (N2360, N2359);
and AND2 (N2361, N2327, N2194);
nor NOR3 (N2362, N2356, N2110, N1196);
and AND3 (N2363, N2362, N552, N1782);
nor NOR4 (N2364, N2347, N1932, N2162, N1543);
nand NAND2 (N2365, N2361, N764);
or OR3 (N2366, N2355, N640, N1174);
nor NOR4 (N2367, N2348, N605, N2115, N1801);
xor XOR2 (N2368, N2358, N941);
and AND2 (N2369, N2364, N2030);
nand NAND4 (N2370, N2367, N2285, N68, N1416);
or OR2 (N2371, N2357, N427);
or OR4 (N2372, N2365, N1831, N1935, N2288);
xor XOR2 (N2373, N2369, N404);
xor XOR2 (N2374, N2337, N11);
and AND4 (N2375, N2368, N1994, N841, N1588);
not NOT1 (N2376, N2372);
and AND4 (N2377, N2366, N1263, N1447, N2374);
or OR2 (N2378, N1433, N438);
or OR3 (N2379, N2373, N282, N189);
not NOT1 (N2380, N2379);
and AND3 (N2381, N2351, N229, N554);
or OR3 (N2382, N2381, N366, N1603);
or OR2 (N2383, N2375, N2012);
not NOT1 (N2384, N2377);
nand NAND4 (N2385, N2363, N1438, N1676, N894);
or OR2 (N2386, N2380, N25);
and AND3 (N2387, N2360, N1326, N1641);
nand NAND3 (N2388, N2387, N2174, N2370);
or OR4 (N2389, N2005, N1340, N1441, N2267);
xor XOR2 (N2390, N2386, N262);
not NOT1 (N2391, N2385);
nand NAND2 (N2392, N2371, N2231);
not NOT1 (N2393, N2388);
xor XOR2 (N2394, N2383, N1432);
not NOT1 (N2395, N2384);
xor XOR2 (N2396, N2378, N2228);
and AND4 (N2397, N2382, N502, N1402, N1769);
and AND4 (N2398, N2392, N633, N843, N1894);
buf BUF1 (N2399, N2394);
or OR4 (N2400, N2376, N971, N1351, N1959);
and AND3 (N2401, N2396, N24, N1963);
buf BUF1 (N2402, N2390);
buf BUF1 (N2403, N2400);
buf BUF1 (N2404, N2389);
xor XOR2 (N2405, N2399, N793);
and AND2 (N2406, N2397, N2374);
nand NAND3 (N2407, N2398, N1178, N54);
xor XOR2 (N2408, N2401, N1460);
nand NAND3 (N2409, N2393, N1456, N1357);
not NOT1 (N2410, N2395);
nor NOR4 (N2411, N2405, N94, N1351, N87);
nor NOR3 (N2412, N2408, N2136, N884);
or OR3 (N2413, N2402, N273, N1223);
not NOT1 (N2414, N2403);
nand NAND3 (N2415, N2412, N387, N1055);
buf BUF1 (N2416, N2404);
not NOT1 (N2417, N2413);
or OR2 (N2418, N2391, N337);
not NOT1 (N2419, N2416);
not NOT1 (N2420, N2406);
nor NOR4 (N2421, N2414, N2406, N1628, N109);
or OR2 (N2422, N2420, N2072);
nor NOR2 (N2423, N2409, N557);
xor XOR2 (N2424, N2407, N982);
nand NAND2 (N2425, N2421, N721);
xor XOR2 (N2426, N2411, N1927);
not NOT1 (N2427, N2417);
nand NAND3 (N2428, N2426, N648, N1313);
or OR3 (N2429, N2424, N557, N451);
buf BUF1 (N2430, N2422);
nor NOR3 (N2431, N2410, N2201, N1201);
buf BUF1 (N2432, N2430);
and AND2 (N2433, N2418, N1517);
not NOT1 (N2434, N2425);
not NOT1 (N2435, N2433);
or OR2 (N2436, N2432, N1183);
nor NOR4 (N2437, N2428, N861, N86, N961);
nand NAND4 (N2438, N2435, N1641, N1578, N271);
nor NOR4 (N2439, N2434, N764, N1817, N562);
xor XOR2 (N2440, N2427, N1341);
xor XOR2 (N2441, N2438, N1511);
not NOT1 (N2442, N2439);
buf BUF1 (N2443, N2436);
xor XOR2 (N2444, N2443, N1583);
not NOT1 (N2445, N2423);
not NOT1 (N2446, N2442);
buf BUF1 (N2447, N2445);
not NOT1 (N2448, N2415);
or OR4 (N2449, N2444, N2398, N1894, N214);
or OR4 (N2450, N2440, N1271, N432, N490);
nor NOR2 (N2451, N2450, N1279);
nor NOR2 (N2452, N2431, N376);
buf BUF1 (N2453, N2447);
or OR2 (N2454, N2437, N300);
or OR2 (N2455, N2419, N632);
or OR3 (N2456, N2448, N1973, N2424);
and AND3 (N2457, N2456, N2351, N1526);
buf BUF1 (N2458, N2446);
and AND4 (N2459, N2458, N2313, N2310, N2404);
nor NOR2 (N2460, N2454, N1903);
not NOT1 (N2461, N2451);
and AND4 (N2462, N2461, N2044, N1390, N1741);
buf BUF1 (N2463, N2460);
nor NOR3 (N2464, N2463, N59, N1745);
and AND4 (N2465, N2453, N2033, N1297, N796);
buf BUF1 (N2466, N2452);
or OR3 (N2467, N2465, N2457, N1654);
and AND3 (N2468, N861, N546, N724);
or OR2 (N2469, N2449, N2005);
not NOT1 (N2470, N2466);
and AND2 (N2471, N2469, N1512);
nor NOR4 (N2472, N2455, N874, N1321, N2252);
nand NAND3 (N2473, N2470, N1880, N1621);
not NOT1 (N2474, N2441);
nand NAND3 (N2475, N2464, N1903, N1164);
and AND2 (N2476, N2462, N171);
buf BUF1 (N2477, N2467);
not NOT1 (N2478, N2475);
nor NOR2 (N2479, N2429, N579);
or OR2 (N2480, N2471, N2477);
xor XOR2 (N2481, N1074, N99);
and AND4 (N2482, N2476, N546, N138, N1302);
buf BUF1 (N2483, N2473);
not NOT1 (N2484, N2468);
nand NAND3 (N2485, N2481, N1794, N180);
not NOT1 (N2486, N2459);
xor XOR2 (N2487, N2485, N734);
and AND4 (N2488, N2483, N1469, N1408, N59);
or OR2 (N2489, N2479, N1010);
nor NOR3 (N2490, N2478, N947, N915);
nand NAND4 (N2491, N2472, N2062, N749, N572);
buf BUF1 (N2492, N2487);
buf BUF1 (N2493, N2482);
xor XOR2 (N2494, N2484, N747);
xor XOR2 (N2495, N2490, N702);
or OR3 (N2496, N2488, N1069, N2302);
xor XOR2 (N2497, N2494, N109);
not NOT1 (N2498, N2493);
and AND2 (N2499, N2497, N2029);
nand NAND2 (N2500, N2498, N321);
buf BUF1 (N2501, N2489);
or OR2 (N2502, N2486, N400);
not NOT1 (N2503, N2501);
not NOT1 (N2504, N2499);
buf BUF1 (N2505, N2474);
and AND3 (N2506, N2492, N1407, N1857);
or OR4 (N2507, N2502, N2031, N1770, N59);
not NOT1 (N2508, N2507);
or OR4 (N2509, N2495, N1170, N837, N1539);
nand NAND4 (N2510, N2496, N2044, N1523, N1519);
not NOT1 (N2511, N2503);
nand NAND4 (N2512, N2510, N386, N104, N2474);
buf BUF1 (N2513, N2508);
or OR3 (N2514, N2491, N190, N1453);
and AND2 (N2515, N2511, N1020);
and AND3 (N2516, N2506, N1389, N879);
xor XOR2 (N2517, N2480, N463);
nand NAND3 (N2518, N2516, N1664, N316);
not NOT1 (N2519, N2515);
buf BUF1 (N2520, N2505);
or OR4 (N2521, N2500, N2163, N1156, N1303);
or OR2 (N2522, N2518, N1633);
or OR3 (N2523, N2514, N2326, N1764);
nor NOR3 (N2524, N2517, N2372, N282);
or OR4 (N2525, N2520, N947, N1998, N1873);
xor XOR2 (N2526, N2522, N1153);
or OR4 (N2527, N2504, N498, N1451, N449);
or OR4 (N2528, N2509, N1438, N650, N973);
buf BUF1 (N2529, N2519);
buf BUF1 (N2530, N2526);
nand NAND3 (N2531, N2524, N878, N2486);
xor XOR2 (N2532, N2528, N857);
not NOT1 (N2533, N2532);
xor XOR2 (N2534, N2531, N51);
or OR2 (N2535, N2527, N2452);
buf BUF1 (N2536, N2530);
nand NAND4 (N2537, N2534, N1357, N1889, N1431);
buf BUF1 (N2538, N2525);
nand NAND2 (N2539, N2513, N1819);
and AND2 (N2540, N2512, N1828);
xor XOR2 (N2541, N2538, N2520);
nor NOR4 (N2542, N2537, N1710, N537, N2048);
buf BUF1 (N2543, N2523);
nand NAND4 (N2544, N2536, N1324, N1989, N1324);
and AND3 (N2545, N2543, N1622, N1761);
xor XOR2 (N2546, N2535, N262);
not NOT1 (N2547, N2540);
xor XOR2 (N2548, N2529, N1385);
and AND3 (N2549, N2542, N2397, N1094);
and AND4 (N2550, N2544, N1182, N1590, N29);
xor XOR2 (N2551, N2546, N818);
nor NOR4 (N2552, N2547, N995, N503, N2228);
xor XOR2 (N2553, N2550, N2088);
xor XOR2 (N2554, N2549, N210);
buf BUF1 (N2555, N2539);
or OR2 (N2556, N2552, N1107);
xor XOR2 (N2557, N2548, N1998);
or OR2 (N2558, N2553, N2424);
buf BUF1 (N2559, N2521);
xor XOR2 (N2560, N2554, N1293);
and AND2 (N2561, N2558, N1754);
not NOT1 (N2562, N2541);
xor XOR2 (N2563, N2561, N2252);
not NOT1 (N2564, N2563);
nor NOR4 (N2565, N2560, N125, N1443, N1644);
not NOT1 (N2566, N2533);
nand NAND3 (N2567, N2557, N1311, N1517);
and AND3 (N2568, N2562, N1260, N1238);
nor NOR2 (N2569, N2551, N1833);
nand NAND4 (N2570, N2565, N1906, N586, N1666);
buf BUF1 (N2571, N2570);
xor XOR2 (N2572, N2555, N1188);
buf BUF1 (N2573, N2571);
buf BUF1 (N2574, N2568);
nor NOR3 (N2575, N2545, N1300, N2187);
not NOT1 (N2576, N2567);
and AND4 (N2577, N2569, N811, N1574, N914);
buf BUF1 (N2578, N2559);
and AND2 (N2579, N2556, N376);
xor XOR2 (N2580, N2575, N375);
not NOT1 (N2581, N2572);
or OR3 (N2582, N2580, N710, N107);
not NOT1 (N2583, N2573);
or OR2 (N2584, N2566, N1626);
and AND4 (N2585, N2577, N1908, N154, N1318);
xor XOR2 (N2586, N2584, N590);
nand NAND2 (N2587, N2564, N1648);
xor XOR2 (N2588, N2582, N354);
xor XOR2 (N2589, N2579, N2521);
and AND4 (N2590, N2576, N180, N1628, N2126);
nand NAND4 (N2591, N2587, N431, N2203, N1583);
and AND2 (N2592, N2581, N1866);
and AND2 (N2593, N2591, N2094);
nand NAND3 (N2594, N2586, N1029, N857);
nor NOR2 (N2595, N2592, N259);
xor XOR2 (N2596, N2595, N851);
nand NAND2 (N2597, N2589, N1214);
xor XOR2 (N2598, N2585, N709);
buf BUF1 (N2599, N2596);
and AND4 (N2600, N2599, N738, N1007, N1276);
buf BUF1 (N2601, N2588);
buf BUF1 (N2602, N2598);
and AND2 (N2603, N2593, N2472);
xor XOR2 (N2604, N2590, N1528);
buf BUF1 (N2605, N2597);
nor NOR2 (N2606, N2578, N602);
not NOT1 (N2607, N2594);
nand NAND2 (N2608, N2600, N1797);
buf BUF1 (N2609, N2603);
nor NOR3 (N2610, N2601, N2137, N97);
xor XOR2 (N2611, N2608, N437);
buf BUF1 (N2612, N2611);
nor NOR2 (N2613, N2574, N2170);
buf BUF1 (N2614, N2607);
xor XOR2 (N2615, N2609, N1197);
nand NAND2 (N2616, N2605, N177);
nand NAND2 (N2617, N2602, N353);
nor NOR2 (N2618, N2617, N1559);
xor XOR2 (N2619, N2583, N2177);
not NOT1 (N2620, N2604);
and AND3 (N2621, N2612, N582, N1044);
nand NAND2 (N2622, N2614, N1488);
or OR4 (N2623, N2615, N740, N1604, N842);
buf BUF1 (N2624, N2606);
xor XOR2 (N2625, N2621, N1971);
nor NOR3 (N2626, N2613, N315, N681);
or OR2 (N2627, N2610, N1651);
nand NAND2 (N2628, N2624, N2378);
not NOT1 (N2629, N2616);
and AND3 (N2630, N2626, N789, N23);
buf BUF1 (N2631, N2630);
or OR3 (N2632, N2623, N1791, N1913);
not NOT1 (N2633, N2632);
xor XOR2 (N2634, N2633, N565);
nor NOR3 (N2635, N2634, N843, N318);
xor XOR2 (N2636, N2625, N1339);
nor NOR4 (N2637, N2627, N1409, N1107, N43);
not NOT1 (N2638, N2619);
or OR3 (N2639, N2631, N1410, N1498);
and AND3 (N2640, N2637, N2225, N2569);
nand NAND4 (N2641, N2618, N28, N2188, N1546);
nand NAND4 (N2642, N2628, N44, N1122, N1692);
and AND2 (N2643, N2640, N2072);
not NOT1 (N2644, N2629);
not NOT1 (N2645, N2638);
buf BUF1 (N2646, N2635);
buf BUF1 (N2647, N2620);
buf BUF1 (N2648, N2644);
and AND3 (N2649, N2622, N630, N429);
xor XOR2 (N2650, N2642, N2464);
buf BUF1 (N2651, N2639);
and AND3 (N2652, N2645, N2115, N306);
not NOT1 (N2653, N2648);
not NOT1 (N2654, N2653);
xor XOR2 (N2655, N2643, N1434);
or OR4 (N2656, N2655, N1548, N678, N2418);
and AND4 (N2657, N2654, N2020, N682, N2380);
nor NOR4 (N2658, N2647, N1331, N1930, N1549);
xor XOR2 (N2659, N2641, N1581);
and AND3 (N2660, N2650, N79, N428);
nand NAND2 (N2661, N2651, N1922);
xor XOR2 (N2662, N2661, N302);
nand NAND4 (N2663, N2659, N188, N1037, N134);
xor XOR2 (N2664, N2658, N1405);
buf BUF1 (N2665, N2662);
nor NOR4 (N2666, N2652, N2256, N2394, N2162);
nand NAND4 (N2667, N2664, N2127, N1859, N143);
and AND4 (N2668, N2649, N1362, N2385, N375);
buf BUF1 (N2669, N2668);
not NOT1 (N2670, N2656);
and AND3 (N2671, N2663, N101, N1961);
not NOT1 (N2672, N2660);
nor NOR2 (N2673, N2646, N1283);
xor XOR2 (N2674, N2671, N1175);
xor XOR2 (N2675, N2665, N2416);
or OR4 (N2676, N2673, N2668, N1750, N362);
buf BUF1 (N2677, N2669);
xor XOR2 (N2678, N2636, N393);
and AND3 (N2679, N2666, N1212, N696);
nor NOR3 (N2680, N2674, N1890, N296);
nor NOR4 (N2681, N2667, N608, N2047, N1783);
xor XOR2 (N2682, N2672, N2555);
xor XOR2 (N2683, N2657, N1331);
buf BUF1 (N2684, N2678);
nor NOR2 (N2685, N2670, N1406);
nand NAND2 (N2686, N2676, N2380);
buf BUF1 (N2687, N2683);
xor XOR2 (N2688, N2685, N801);
nor NOR4 (N2689, N2686, N1169, N2305, N792);
nand NAND3 (N2690, N2689, N1097, N1850);
nor NOR3 (N2691, N2684, N1040, N317);
and AND2 (N2692, N2682, N2505);
or OR4 (N2693, N2692, N75, N1808, N526);
xor XOR2 (N2694, N2687, N989);
nor NOR3 (N2695, N2693, N2554, N64);
and AND2 (N2696, N2690, N2378);
xor XOR2 (N2697, N2679, N852);
nand NAND4 (N2698, N2677, N1374, N2489, N1005);
nor NOR2 (N2699, N2694, N1888);
or OR3 (N2700, N2688, N908, N497);
and AND3 (N2701, N2675, N1707, N469);
or OR4 (N2702, N2698, N1796, N2623, N1583);
xor XOR2 (N2703, N2695, N1403);
not NOT1 (N2704, N2681);
not NOT1 (N2705, N2691);
or OR2 (N2706, N2699, N2627);
buf BUF1 (N2707, N2703);
xor XOR2 (N2708, N2697, N2259);
nor NOR4 (N2709, N2696, N2403, N1512, N883);
and AND2 (N2710, N2705, N2679);
nor NOR3 (N2711, N2704, N275, N2286);
nor NOR3 (N2712, N2700, N1078, N759);
not NOT1 (N2713, N2707);
xor XOR2 (N2714, N2709, N1133);
buf BUF1 (N2715, N2708);
not NOT1 (N2716, N2714);
xor XOR2 (N2717, N2711, N2053);
nand NAND2 (N2718, N2680, N2715);
buf BUF1 (N2719, N2247);
nand NAND4 (N2720, N2718, N1641, N1526, N1975);
buf BUF1 (N2721, N2719);
nand NAND3 (N2722, N2713, N2298, N1031);
nand NAND2 (N2723, N2722, N2385);
and AND3 (N2724, N2706, N2338, N1525);
or OR4 (N2725, N2720, N2614, N1370, N1986);
not NOT1 (N2726, N2725);
or OR4 (N2727, N2717, N1188, N1072, N2598);
and AND3 (N2728, N2710, N2200, N1501);
not NOT1 (N2729, N2726);
xor XOR2 (N2730, N2702, N496);
or OR2 (N2731, N2712, N634);
buf BUF1 (N2732, N2721);
and AND4 (N2733, N2716, N143, N2118, N482);
buf BUF1 (N2734, N2733);
nor NOR2 (N2735, N2732, N1557);
nand NAND2 (N2736, N2731, N2679);
and AND3 (N2737, N2723, N118, N820);
not NOT1 (N2738, N2728);
nor NOR4 (N2739, N2727, N1257, N2157, N2389);
xor XOR2 (N2740, N2724, N1850);
not NOT1 (N2741, N2730);
or OR2 (N2742, N2729, N1168);
nand NAND2 (N2743, N2735, N1754);
nor NOR2 (N2744, N2739, N182);
not NOT1 (N2745, N2740);
and AND3 (N2746, N2736, N784, N1897);
not NOT1 (N2747, N2742);
nand NAND2 (N2748, N2746, N2168);
and AND3 (N2749, N2743, N297, N1010);
nand NAND4 (N2750, N2734, N2384, N486, N2742);
and AND3 (N2751, N2737, N1809, N900);
buf BUF1 (N2752, N2749);
not NOT1 (N2753, N2750);
or OR4 (N2754, N2753, N943, N1229, N2424);
or OR2 (N2755, N2701, N974);
nand NAND4 (N2756, N2738, N391, N869, N1798);
nor NOR4 (N2757, N2754, N2104, N1593, N1937);
buf BUF1 (N2758, N2751);
nor NOR4 (N2759, N2747, N804, N1225, N33);
and AND2 (N2760, N2758, N21);
and AND4 (N2761, N2741, N1323, N2350, N2461);
nor NOR4 (N2762, N2761, N1743, N1121, N50);
buf BUF1 (N2763, N2748);
and AND4 (N2764, N2752, N2651, N889, N1795);
nor NOR4 (N2765, N2759, N1202, N1228, N2060);
nand NAND3 (N2766, N2756, N1389, N1816);
or OR2 (N2767, N2763, N647);
xor XOR2 (N2768, N2755, N2743);
nand NAND4 (N2769, N2767, N93, N2368, N983);
or OR3 (N2770, N2768, N940, N1936);
buf BUF1 (N2771, N2766);
or OR4 (N2772, N2765, N1194, N1961, N2119);
not NOT1 (N2773, N2762);
xor XOR2 (N2774, N2745, N1509);
nand NAND4 (N2775, N2773, N2319, N1165, N789);
and AND3 (N2776, N2775, N2707, N2401);
nor NOR3 (N2777, N2772, N128, N2453);
not NOT1 (N2778, N2771);
buf BUF1 (N2779, N2776);
buf BUF1 (N2780, N2760);
nor NOR3 (N2781, N2777, N1491, N2004);
not NOT1 (N2782, N2764);
nor NOR2 (N2783, N2770, N190);
and AND4 (N2784, N2781, N551, N445, N2482);
and AND2 (N2785, N2782, N1732);
nor NOR4 (N2786, N2780, N1384, N2247, N1762);
nand NAND3 (N2787, N2757, N673, N2320);
xor XOR2 (N2788, N2774, N2173);
buf BUF1 (N2789, N2784);
nor NOR2 (N2790, N2786, N2234);
xor XOR2 (N2791, N2783, N779);
buf BUF1 (N2792, N2769);
nor NOR4 (N2793, N2788, N2760, N2713, N2053);
buf BUF1 (N2794, N2787);
buf BUF1 (N2795, N2789);
nand NAND2 (N2796, N2792, N242);
buf BUF1 (N2797, N2796);
and AND2 (N2798, N2778, N962);
xor XOR2 (N2799, N2793, N2015);
or OR2 (N2800, N2795, N594);
nand NAND4 (N2801, N2744, N969, N450, N1086);
nand NAND2 (N2802, N2794, N1195);
nor NOR4 (N2803, N2802, N342, N1148, N2047);
nand NAND2 (N2804, N2791, N35);
or OR2 (N2805, N2779, N1189);
nor NOR3 (N2806, N2799, N1965, N140);
nor NOR3 (N2807, N2800, N1023, N2751);
or OR3 (N2808, N2790, N452, N1934);
xor XOR2 (N2809, N2804, N460);
nand NAND4 (N2810, N2785, N1101, N1033, N615);
and AND4 (N2811, N2806, N2102, N1589, N2535);
nor NOR3 (N2812, N2807, N2042, N1844);
xor XOR2 (N2813, N2810, N511);
not NOT1 (N2814, N2797);
nand NAND2 (N2815, N2805, N1593);
buf BUF1 (N2816, N2809);
and AND4 (N2817, N2803, N569, N937, N649);
not NOT1 (N2818, N2813);
or OR4 (N2819, N2814, N241, N1575, N2158);
nor NOR3 (N2820, N2815, N1280, N1464);
nand NAND4 (N2821, N2819, N662, N983, N2453);
or OR4 (N2822, N2820, N1639, N1939, N669);
buf BUF1 (N2823, N2801);
or OR2 (N2824, N2818, N727);
nand NAND2 (N2825, N2824, N950);
nor NOR4 (N2826, N2825, N1743, N1723, N1295);
not NOT1 (N2827, N2811);
not NOT1 (N2828, N2821);
or OR3 (N2829, N2798, N2221, N1775);
nor NOR3 (N2830, N2827, N1736, N2130);
xor XOR2 (N2831, N2826, N2509);
nand NAND3 (N2832, N2830, N2085, N1120);
xor XOR2 (N2833, N2831, N2077);
and AND3 (N2834, N2832, N2589, N872);
not NOT1 (N2835, N2828);
or OR4 (N2836, N2808, N2505, N1182, N1115);
nand NAND2 (N2837, N2836, N1483);
nor NOR3 (N2838, N2823, N1043, N523);
nor NOR3 (N2839, N2816, N713, N848);
nand NAND2 (N2840, N2817, N1263);
and AND2 (N2841, N2829, N1614);
not NOT1 (N2842, N2812);
buf BUF1 (N2843, N2834);
buf BUF1 (N2844, N2822);
nand NAND2 (N2845, N2835, N2510);
or OR3 (N2846, N2841, N1495, N1717);
buf BUF1 (N2847, N2843);
or OR2 (N2848, N2840, N488);
and AND2 (N2849, N2847, N1325);
nor NOR4 (N2850, N2845, N442, N2687, N2207);
xor XOR2 (N2851, N2849, N1748);
nand NAND4 (N2852, N2844, N769, N2647, N2286);
or OR4 (N2853, N2839, N1854, N1983, N806);
xor XOR2 (N2854, N2837, N2725);
buf BUF1 (N2855, N2846);
buf BUF1 (N2856, N2852);
xor XOR2 (N2857, N2855, N1298);
xor XOR2 (N2858, N2857, N441);
nand NAND2 (N2859, N2858, N2766);
xor XOR2 (N2860, N2854, N985);
and AND3 (N2861, N2833, N371, N786);
nor NOR3 (N2862, N2860, N1260, N2223);
and AND4 (N2863, N2838, N2355, N2259, N1078);
nor NOR3 (N2864, N2856, N728, N1408);
not NOT1 (N2865, N2842);
and AND3 (N2866, N2863, N1769, N1522);
and AND4 (N2867, N2850, N394, N2385, N2502);
nand NAND2 (N2868, N2864, N2590);
nand NAND2 (N2869, N2851, N2074);
or OR3 (N2870, N2868, N2806, N181);
buf BUF1 (N2871, N2865);
or OR4 (N2872, N2862, N1001, N1412, N1645);
or OR3 (N2873, N2872, N339, N127);
nand NAND2 (N2874, N2873, N2358);
not NOT1 (N2875, N2870);
xor XOR2 (N2876, N2848, N1017);
xor XOR2 (N2877, N2875, N45);
xor XOR2 (N2878, N2869, N2460);
or OR2 (N2879, N2878, N2264);
nor NOR4 (N2880, N2877, N453, N204, N1057);
buf BUF1 (N2881, N2866);
nor NOR3 (N2882, N2876, N51, N224);
or OR2 (N2883, N2882, N1620);
nand NAND2 (N2884, N2853, N2257);
nor NOR3 (N2885, N2867, N1638, N2846);
and AND2 (N2886, N2871, N337);
not NOT1 (N2887, N2885);
nor NOR4 (N2888, N2879, N953, N1362, N2776);
nand NAND3 (N2889, N2883, N211, N2104);
xor XOR2 (N2890, N2889, N1109);
not NOT1 (N2891, N2888);
not NOT1 (N2892, N2880);
buf BUF1 (N2893, N2859);
xor XOR2 (N2894, N2874, N2395);
not NOT1 (N2895, N2861);
not NOT1 (N2896, N2893);
nand NAND3 (N2897, N2887, N1859, N2881);
not NOT1 (N2898, N2273);
and AND2 (N2899, N2891, N1649);
buf BUF1 (N2900, N2894);
not NOT1 (N2901, N2884);
nand NAND4 (N2902, N2890, N1772, N28, N12);
and AND2 (N2903, N2900, N1773);
not NOT1 (N2904, N2895);
not NOT1 (N2905, N2892);
nand NAND2 (N2906, N2902, N117);
xor XOR2 (N2907, N2905, N2421);
nor NOR4 (N2908, N2886, N779, N2008, N1078);
xor XOR2 (N2909, N2896, N1182);
and AND3 (N2910, N2906, N919, N1695);
nand NAND3 (N2911, N2898, N1904, N2582);
not NOT1 (N2912, N2907);
nand NAND3 (N2913, N2908, N2767, N1613);
or OR2 (N2914, N2912, N1494);
not NOT1 (N2915, N2904);
and AND4 (N2916, N2914, N511, N546, N1870);
buf BUF1 (N2917, N2913);
not NOT1 (N2918, N2916);
or OR2 (N2919, N2909, N2412);
or OR4 (N2920, N2915, N308, N139, N866);
buf BUF1 (N2921, N2920);
nor NOR2 (N2922, N2910, N2800);
or OR2 (N2923, N2901, N1178);
xor XOR2 (N2924, N2899, N1337);
xor XOR2 (N2925, N2903, N1244);
xor XOR2 (N2926, N2923, N2801);
or OR2 (N2927, N2918, N390);
and AND2 (N2928, N2922, N1774);
xor XOR2 (N2929, N2924, N2423);
nand NAND2 (N2930, N2925, N1475);
xor XOR2 (N2931, N2917, N2582);
or OR2 (N2932, N2929, N445);
not NOT1 (N2933, N2930);
nor NOR4 (N2934, N2919, N2509, N2022, N2046);
nand NAND3 (N2935, N2926, N2818, N2129);
and AND3 (N2936, N2935, N958, N808);
buf BUF1 (N2937, N2936);
xor XOR2 (N2938, N2934, N335);
not NOT1 (N2939, N2897);
xor XOR2 (N2940, N2921, N167);
xor XOR2 (N2941, N2911, N2575);
nor NOR2 (N2942, N2938, N715);
nand NAND2 (N2943, N2933, N2647);
or OR3 (N2944, N2927, N1258, N68);
nand NAND3 (N2945, N2932, N461, N499);
buf BUF1 (N2946, N2945);
or OR3 (N2947, N2939, N1399, N1466);
or OR4 (N2948, N2937, N589, N2930, N708);
nor NOR2 (N2949, N2941, N46);
not NOT1 (N2950, N2928);
nand NAND4 (N2951, N2931, N2324, N2588, N537);
not NOT1 (N2952, N2943);
nor NOR4 (N2953, N2947, N2186, N2029, N1919);
and AND3 (N2954, N2942, N2766, N588);
nor NOR3 (N2955, N2950, N2208, N119);
or OR3 (N2956, N2948, N512, N1382);
or OR3 (N2957, N2946, N2478, N2001);
nand NAND4 (N2958, N2940, N2308, N2151, N2525);
and AND3 (N2959, N2956, N1967, N1615);
not NOT1 (N2960, N2944);
xor XOR2 (N2961, N2954, N2048);
xor XOR2 (N2962, N2959, N455);
buf BUF1 (N2963, N2962);
not NOT1 (N2964, N2952);
and AND3 (N2965, N2961, N849, N1463);
xor XOR2 (N2966, N2949, N679);
or OR3 (N2967, N2963, N1363, N1739);
nor NOR2 (N2968, N2960, N2832);
or OR3 (N2969, N2967, N338, N2458);
or OR2 (N2970, N2955, N1495);
nor NOR3 (N2971, N2964, N1659, N750);
nand NAND4 (N2972, N2970, N2240, N2068, N2061);
not NOT1 (N2973, N2972);
buf BUF1 (N2974, N2958);
and AND2 (N2975, N2971, N2759);
not NOT1 (N2976, N2951);
buf BUF1 (N2977, N2957);
buf BUF1 (N2978, N2977);
nor NOR3 (N2979, N2978, N2000, N2868);
and AND2 (N2980, N2953, N1541);
not NOT1 (N2981, N2968);
not NOT1 (N2982, N2980);
nor NOR2 (N2983, N2974, N1258);
xor XOR2 (N2984, N2982, N2407);
nand NAND4 (N2985, N2979, N427, N352, N2218);
and AND4 (N2986, N2981, N2410, N499, N945);
nor NOR4 (N2987, N2985, N2138, N1410, N2789);
not NOT1 (N2988, N2966);
nor NOR2 (N2989, N2975, N2155);
and AND4 (N2990, N2984, N18, N1218, N2965);
and AND3 (N2991, N2095, N1736, N64);
nand NAND4 (N2992, N2976, N2447, N1382, N2071);
nand NAND3 (N2993, N2986, N2738, N31);
or OR3 (N2994, N2983, N747, N1016);
and AND4 (N2995, N2994, N1010, N2351, N2528);
buf BUF1 (N2996, N2995);
xor XOR2 (N2997, N2989, N126);
xor XOR2 (N2998, N2992, N2606);
nor NOR3 (N2999, N2987, N383, N324);
nand NAND2 (N3000, N2990, N2234);
and AND4 (N3001, N2999, N1544, N939, N1086);
nor NOR4 (N3002, N2973, N1900, N355, N2515);
or OR3 (N3003, N2988, N1493, N2361);
nor NOR4 (N3004, N2969, N2297, N1670, N1091);
nor NOR2 (N3005, N3001, N2067);
xor XOR2 (N3006, N3002, N2594);
or OR3 (N3007, N2993, N1059, N2638);
or OR4 (N3008, N2991, N2150, N1310, N1501);
not NOT1 (N3009, N3008);
not NOT1 (N3010, N3007);
or OR2 (N3011, N2998, N2467);
and AND4 (N3012, N3010, N2510, N1068, N1574);
buf BUF1 (N3013, N3009);
buf BUF1 (N3014, N3013);
not NOT1 (N3015, N2996);
buf BUF1 (N3016, N3012);
or OR4 (N3017, N3014, N2302, N1087, N424);
buf BUF1 (N3018, N2997);
or OR2 (N3019, N3017, N2052);
xor XOR2 (N3020, N3019, N1322);
not NOT1 (N3021, N3020);
xor XOR2 (N3022, N3015, N1790);
not NOT1 (N3023, N3016);
not NOT1 (N3024, N3005);
xor XOR2 (N3025, N3011, N2438);
xor XOR2 (N3026, N3018, N961);
nand NAND4 (N3027, N3026, N2284, N2356, N2736);
xor XOR2 (N3028, N3000, N12);
buf BUF1 (N3029, N3028);
nand NAND3 (N3030, N3006, N2212, N2093);
buf BUF1 (N3031, N3029);
xor XOR2 (N3032, N3031, N4);
nand NAND4 (N3033, N3030, N175, N1605, N2162);
nand NAND3 (N3034, N3004, N457, N2103);
not NOT1 (N3035, N3032);
buf BUF1 (N3036, N3023);
or OR3 (N3037, N3024, N6, N2951);
and AND3 (N3038, N3033, N571, N1949);
nand NAND2 (N3039, N3037, N954);
xor XOR2 (N3040, N3025, N2414);
nand NAND2 (N3041, N3021, N1903);
and AND2 (N3042, N3038, N810);
and AND4 (N3043, N3039, N2027, N947, N613);
buf BUF1 (N3044, N3003);
nand NAND2 (N3045, N3027, N2132);
xor XOR2 (N3046, N3041, N333);
xor XOR2 (N3047, N3044, N1462);
buf BUF1 (N3048, N3042);
buf BUF1 (N3049, N3046);
nor NOR4 (N3050, N3022, N1260, N835, N1167);
nand NAND3 (N3051, N3048, N1576, N1105);
and AND4 (N3052, N3036, N2739, N1405, N194);
buf BUF1 (N3053, N3050);
and AND2 (N3054, N3045, N1604);
or OR4 (N3055, N3047, N2071, N1585, N1269);
xor XOR2 (N3056, N3054, N1577);
not NOT1 (N3057, N3056);
buf BUF1 (N3058, N3053);
buf BUF1 (N3059, N3040);
nor NOR2 (N3060, N3058, N52);
xor XOR2 (N3061, N3049, N1229);
not NOT1 (N3062, N3052);
nand NAND3 (N3063, N3043, N1034, N756);
or OR4 (N3064, N3062, N196, N2553, N1073);
not NOT1 (N3065, N3057);
xor XOR2 (N3066, N3060, N1958);
nand NAND4 (N3067, N3055, N808, N2882, N2854);
xor XOR2 (N3068, N3035, N1488);
xor XOR2 (N3069, N3068, N1147);
and AND4 (N3070, N3063, N1669, N1090, N1220);
nor NOR2 (N3071, N3034, N2847);
not NOT1 (N3072, N3066);
and AND2 (N3073, N3067, N1569);
and AND4 (N3074, N3064, N1209, N2901, N2114);
nor NOR3 (N3075, N3070, N1582, N844);
nand NAND2 (N3076, N3071, N1213);
and AND3 (N3077, N3061, N504, N2641);
xor XOR2 (N3078, N3075, N2131);
or OR2 (N3079, N3069, N1428);
nand NAND2 (N3080, N3074, N2056);
buf BUF1 (N3081, N3078);
buf BUF1 (N3082, N3080);
nand NAND3 (N3083, N3051, N2856, N1762);
xor XOR2 (N3084, N3076, N1328);
or OR2 (N3085, N3065, N357);
nor NOR4 (N3086, N3083, N2970, N1639, N1076);
xor XOR2 (N3087, N3081, N1241);
nand NAND4 (N3088, N3072, N1081, N2746, N2716);
buf BUF1 (N3089, N3086);
xor XOR2 (N3090, N3089, N122);
xor XOR2 (N3091, N3084, N1522);
or OR4 (N3092, N3085, N2313, N3083, N922);
or OR4 (N3093, N3059, N2183, N21, N1279);
buf BUF1 (N3094, N3092);
nor NOR3 (N3095, N3093, N2052, N2938);
xor XOR2 (N3096, N3095, N506);
or OR4 (N3097, N3077, N943, N1985, N673);
nor NOR4 (N3098, N3091, N214, N2845, N1562);
buf BUF1 (N3099, N3073);
nand NAND3 (N3100, N3090, N1124, N2883);
or OR3 (N3101, N3099, N1675, N1585);
and AND4 (N3102, N3094, N3037, N1993, N3073);
and AND4 (N3103, N3102, N2188, N2949, N1460);
buf BUF1 (N3104, N3079);
nand NAND4 (N3105, N3104, N1852, N690, N2020);
nand NAND3 (N3106, N3088, N2830, N667);
or OR4 (N3107, N3097, N367, N1444, N2594);
and AND4 (N3108, N3103, N2481, N3075, N659);
nand NAND4 (N3109, N3101, N931, N1391, N2339);
buf BUF1 (N3110, N3105);
or OR4 (N3111, N3109, N880, N3079, N822);
not NOT1 (N3112, N3087);
nor NOR3 (N3113, N3096, N1166, N2303);
buf BUF1 (N3114, N3082);
not NOT1 (N3115, N3114);
not NOT1 (N3116, N3110);
nand NAND4 (N3117, N3098, N2639, N3091, N2986);
or OR3 (N3118, N3100, N2176, N2658);
xor XOR2 (N3119, N3116, N135);
buf BUF1 (N3120, N3119);
nor NOR4 (N3121, N3115, N776, N101, N2187);
not NOT1 (N3122, N3120);
xor XOR2 (N3123, N3106, N1815);
and AND4 (N3124, N3118, N2494, N894, N1928);
nand NAND2 (N3125, N3124, N2142);
not NOT1 (N3126, N3117);
buf BUF1 (N3127, N3125);
and AND3 (N3128, N3113, N1175, N2386);
nand NAND2 (N3129, N3112, N1506);
nor NOR3 (N3130, N3121, N1992, N2814);
nand NAND2 (N3131, N3123, N2886);
buf BUF1 (N3132, N3108);
nand NAND2 (N3133, N3111, N2689);
not NOT1 (N3134, N3131);
xor XOR2 (N3135, N3130, N264);
or OR3 (N3136, N3127, N371, N2172);
buf BUF1 (N3137, N3136);
and AND3 (N3138, N3129, N1620, N870);
not NOT1 (N3139, N3132);
xor XOR2 (N3140, N3134, N1802);
xor XOR2 (N3141, N3126, N1220);
nand NAND4 (N3142, N3128, N93, N1225, N2425);
nand NAND4 (N3143, N3107, N2779, N678, N814);
and AND4 (N3144, N3135, N2578, N2080, N3140);
and AND4 (N3145, N2184, N2718, N2010, N91);
not NOT1 (N3146, N3145);
xor XOR2 (N3147, N3143, N1228);
xor XOR2 (N3148, N3137, N2569);
and AND4 (N3149, N3122, N1526, N2871, N1690);
not NOT1 (N3150, N3139);
not NOT1 (N3151, N3138);
nand NAND3 (N3152, N3144, N1042, N3151);
nand NAND2 (N3153, N1537, N1365);
nand NAND2 (N3154, N3150, N951);
not NOT1 (N3155, N3153);
nand NAND2 (N3156, N3142, N2197);
and AND3 (N3157, N3155, N741, N2639);
nor NOR2 (N3158, N3141, N457);
buf BUF1 (N3159, N3148);
or OR3 (N3160, N3154, N2259, N165);
and AND3 (N3161, N3157, N2765, N2419);
not NOT1 (N3162, N3147);
buf BUF1 (N3163, N3133);
buf BUF1 (N3164, N3152);
nor NOR4 (N3165, N3160, N2067, N2379, N1430);
nor NOR3 (N3166, N3161, N2522, N2566);
and AND2 (N3167, N3158, N2852);
or OR3 (N3168, N3164, N890, N2343);
or OR2 (N3169, N3149, N1529);
and AND4 (N3170, N3165, N1121, N1347, N1794);
nand NAND2 (N3171, N3156, N918);
buf BUF1 (N3172, N3169);
nor NOR3 (N3173, N3171, N2420, N1531);
not NOT1 (N3174, N3146);
not NOT1 (N3175, N3174);
nand NAND3 (N3176, N3173, N1112, N1867);
buf BUF1 (N3177, N3167);
xor XOR2 (N3178, N3162, N1043);
not NOT1 (N3179, N3177);
nor NOR4 (N3180, N3176, N32, N328, N929);
and AND4 (N3181, N3159, N135, N2358, N1414);
nand NAND4 (N3182, N3166, N781, N1742, N1893);
or OR3 (N3183, N3180, N1659, N794);
nand NAND2 (N3184, N3178, N511);
not NOT1 (N3185, N3181);
and AND4 (N3186, N3172, N2117, N151, N1184);
and AND3 (N3187, N3175, N1971, N2558);
nand NAND2 (N3188, N3179, N2873);
not NOT1 (N3189, N3185);
nor NOR3 (N3190, N3163, N1005, N95);
nor NOR2 (N3191, N3190, N1724);
nand NAND3 (N3192, N3189, N1569, N1563);
not NOT1 (N3193, N3182);
not NOT1 (N3194, N3183);
xor XOR2 (N3195, N3184, N1017);
and AND4 (N3196, N3170, N1800, N2313, N726);
or OR2 (N3197, N3196, N3148);
and AND2 (N3198, N3187, N1861);
or OR3 (N3199, N3197, N2873, N1342);
or OR3 (N3200, N3186, N1889, N1053);
not NOT1 (N3201, N3191);
xor XOR2 (N3202, N3193, N848);
not NOT1 (N3203, N3202);
or OR3 (N3204, N3199, N2874, N1565);
nand NAND2 (N3205, N3192, N1988);
buf BUF1 (N3206, N3194);
xor XOR2 (N3207, N3168, N1864);
and AND2 (N3208, N3200, N2720);
xor XOR2 (N3209, N3198, N241);
buf BUF1 (N3210, N3207);
nand NAND4 (N3211, N3195, N2085, N3136, N1850);
or OR2 (N3212, N3210, N2724);
and AND3 (N3213, N3204, N2428, N1518);
xor XOR2 (N3214, N3212, N3005);
nand NAND3 (N3215, N3201, N330, N315);
not NOT1 (N3216, N3214);
or OR4 (N3217, N3216, N2038, N2771, N468);
buf BUF1 (N3218, N3211);
nor NOR2 (N3219, N3215, N1731);
not NOT1 (N3220, N3205);
buf BUF1 (N3221, N3206);
buf BUF1 (N3222, N3203);
nor NOR2 (N3223, N3221, N1085);
buf BUF1 (N3224, N3213);
nand NAND2 (N3225, N3220, N1249);
xor XOR2 (N3226, N3223, N1038);
or OR4 (N3227, N3217, N620, N184, N1378);
nor NOR3 (N3228, N3226, N1687, N2384);
not NOT1 (N3229, N3208);
xor XOR2 (N3230, N3228, N2401);
and AND4 (N3231, N3229, N180, N2996, N553);
not NOT1 (N3232, N3227);
nor NOR3 (N3233, N3219, N1382, N964);
or OR2 (N3234, N3209, N861);
nor NOR2 (N3235, N3225, N868);
not NOT1 (N3236, N3222);
nor NOR2 (N3237, N3224, N2537);
nand NAND4 (N3238, N3232, N2240, N59, N2191);
or OR2 (N3239, N3218, N477);
not NOT1 (N3240, N3238);
not NOT1 (N3241, N3235);
or OR2 (N3242, N3241, N1039);
not NOT1 (N3243, N3240);
or OR3 (N3244, N3236, N1444, N2530);
or OR3 (N3245, N3188, N395, N2);
nor NOR2 (N3246, N3234, N1540);
buf BUF1 (N3247, N3233);
nor NOR3 (N3248, N3245, N372, N1188);
and AND4 (N3249, N3246, N2071, N645, N656);
or OR3 (N3250, N3237, N1387, N2610);
nor NOR2 (N3251, N3243, N996);
and AND4 (N3252, N3251, N3014, N1251, N2969);
and AND2 (N3253, N3244, N2845);
xor XOR2 (N3254, N3250, N3246);
buf BUF1 (N3255, N3230);
buf BUF1 (N3256, N3253);
nor NOR2 (N3257, N3242, N2546);
buf BUF1 (N3258, N3231);
xor XOR2 (N3259, N3252, N930);
nand NAND3 (N3260, N3247, N352, N240);
buf BUF1 (N3261, N3249);
nand NAND4 (N3262, N3239, N2822, N1983, N2162);
buf BUF1 (N3263, N3254);
nor NOR3 (N3264, N3259, N2397, N778);
or OR3 (N3265, N3264, N2558, N2973);
and AND3 (N3266, N3265, N1000, N2049);
and AND4 (N3267, N3255, N2048, N2688, N2610);
buf BUF1 (N3268, N3261);
or OR2 (N3269, N3248, N2376);
not NOT1 (N3270, N3256);
not NOT1 (N3271, N3263);
not NOT1 (N3272, N3270);
nor NOR2 (N3273, N3262, N72);
or OR2 (N3274, N3273, N1154);
not NOT1 (N3275, N3266);
nand NAND4 (N3276, N3258, N1359, N2867, N131);
xor XOR2 (N3277, N3268, N2857);
buf BUF1 (N3278, N3274);
buf BUF1 (N3279, N3260);
not NOT1 (N3280, N3269);
nand NAND4 (N3281, N3267, N2031, N533, N21);
not NOT1 (N3282, N3275);
not NOT1 (N3283, N3278);
not NOT1 (N3284, N3272);
buf BUF1 (N3285, N3283);
xor XOR2 (N3286, N3271, N2588);
or OR4 (N3287, N3284, N298, N2811, N455);
and AND3 (N3288, N3286, N2155, N1590);
nand NAND4 (N3289, N3257, N2220, N1190, N2938);
xor XOR2 (N3290, N3288, N75);
not NOT1 (N3291, N3285);
nand NAND3 (N3292, N3281, N2447, N1182);
not NOT1 (N3293, N3292);
buf BUF1 (N3294, N3282);
and AND2 (N3295, N3294, N39);
nand NAND2 (N3296, N3279, N303);
nand NAND2 (N3297, N3277, N2099);
buf BUF1 (N3298, N3295);
xor XOR2 (N3299, N3290, N1274);
nand NAND3 (N3300, N3291, N3140, N2293);
buf BUF1 (N3301, N3298);
nand NAND4 (N3302, N3297, N2788, N2519, N1342);
or OR3 (N3303, N3280, N936, N2235);
buf BUF1 (N3304, N3300);
or OR2 (N3305, N3304, N1981);
nand NAND4 (N3306, N3296, N1251, N122, N2847);
and AND4 (N3307, N3299, N1191, N2136, N1914);
or OR4 (N3308, N3303, N144, N1168, N1363);
nand NAND3 (N3309, N3293, N3249, N1318);
xor XOR2 (N3310, N3307, N420);
xor XOR2 (N3311, N3302, N3215);
xor XOR2 (N3312, N3311, N392);
or OR2 (N3313, N3289, N2453);
xor XOR2 (N3314, N3306, N14);
buf BUF1 (N3315, N3305);
not NOT1 (N3316, N3315);
buf BUF1 (N3317, N3276);
xor XOR2 (N3318, N3312, N2730);
and AND3 (N3319, N3318, N2851, N2584);
and AND2 (N3320, N3310, N845);
buf BUF1 (N3321, N3287);
xor XOR2 (N3322, N3321, N3228);
not NOT1 (N3323, N3319);
nand NAND2 (N3324, N3317, N319);
not NOT1 (N3325, N3313);
xor XOR2 (N3326, N3309, N2865);
xor XOR2 (N3327, N3316, N2108);
nand NAND3 (N3328, N3325, N110, N1675);
xor XOR2 (N3329, N3322, N1962);
and AND3 (N3330, N3327, N1587, N862);
or OR4 (N3331, N3330, N1112, N1191, N1983);
not NOT1 (N3332, N3329);
nand NAND3 (N3333, N3326, N28, N685);
not NOT1 (N3334, N3332);
nor NOR3 (N3335, N3314, N1191, N1532);
or OR4 (N3336, N3333, N2752, N762, N2837);
not NOT1 (N3337, N3308);
not NOT1 (N3338, N3320);
nand NAND4 (N3339, N3331, N1888, N1657, N1426);
buf BUF1 (N3340, N3301);
not NOT1 (N3341, N3334);
xor XOR2 (N3342, N3328, N2484);
and AND2 (N3343, N3338, N2621);
buf BUF1 (N3344, N3342);
buf BUF1 (N3345, N3343);
xor XOR2 (N3346, N3324, N134);
xor XOR2 (N3347, N3345, N2507);
nand NAND4 (N3348, N3336, N2244, N1950, N1026);
and AND4 (N3349, N3335, N1967, N2700, N2320);
and AND3 (N3350, N3348, N1742, N49);
buf BUF1 (N3351, N3350);
or OR4 (N3352, N3351, N1646, N1999, N764);
not NOT1 (N3353, N3344);
nand NAND3 (N3354, N3347, N1670, N706);
and AND4 (N3355, N3337, N1174, N2313, N1432);
or OR2 (N3356, N3346, N679);
nand NAND4 (N3357, N3339, N985, N173, N272);
nor NOR3 (N3358, N3341, N1492, N2945);
not NOT1 (N3359, N3358);
nor NOR3 (N3360, N3353, N1072, N88);
not NOT1 (N3361, N3355);
not NOT1 (N3362, N3359);
nand NAND3 (N3363, N3357, N1823, N3208);
not NOT1 (N3364, N3323);
or OR2 (N3365, N3354, N2175);
and AND4 (N3366, N3340, N909, N190, N1557);
nand NAND4 (N3367, N3361, N1715, N563, N2413);
buf BUF1 (N3368, N3366);
and AND3 (N3369, N3368, N1740, N2998);
not NOT1 (N3370, N3356);
buf BUF1 (N3371, N3363);
buf BUF1 (N3372, N3365);
buf BUF1 (N3373, N3362);
not NOT1 (N3374, N3371);
nand NAND4 (N3375, N3373, N1342, N2707, N177);
nor NOR4 (N3376, N3375, N901, N3345, N121);
or OR2 (N3377, N3367, N2687);
nor NOR4 (N3378, N3377, N2942, N569, N2518);
and AND2 (N3379, N3378, N74);
nand NAND3 (N3380, N3379, N2086, N2687);
nor NOR4 (N3381, N3369, N1920, N2996, N1959);
or OR2 (N3382, N3360, N1460);
nor NOR3 (N3383, N3376, N1611, N1718);
and AND2 (N3384, N3370, N2207);
and AND2 (N3385, N3374, N2832);
nor NOR4 (N3386, N3383, N2512, N735, N826);
or OR4 (N3387, N3381, N1142, N2660, N3230);
not NOT1 (N3388, N3352);
or OR4 (N3389, N3372, N3155, N1755, N2485);
or OR4 (N3390, N3386, N2258, N3153, N1929);
or OR4 (N3391, N3382, N3097, N37, N3209);
and AND4 (N3392, N3380, N2857, N265, N2477);
nor NOR4 (N3393, N3392, N312, N651, N2946);
buf BUF1 (N3394, N3388);
nor NOR4 (N3395, N3384, N2630, N1666, N2063);
and AND3 (N3396, N3385, N2737, N2814);
and AND2 (N3397, N3395, N472);
not NOT1 (N3398, N3393);
nor NOR2 (N3399, N3396, N2788);
not NOT1 (N3400, N3349);
nor NOR4 (N3401, N3398, N3087, N2666, N2914);
xor XOR2 (N3402, N3390, N216);
xor XOR2 (N3403, N3397, N1661);
nand NAND3 (N3404, N3403, N726, N598);
nor NOR4 (N3405, N3404, N395, N1124, N2662);
xor XOR2 (N3406, N3364, N2422);
xor XOR2 (N3407, N3401, N167);
and AND4 (N3408, N3406, N2583, N1647, N1238);
xor XOR2 (N3409, N3391, N909);
not NOT1 (N3410, N3399);
not NOT1 (N3411, N3402);
xor XOR2 (N3412, N3405, N2685);
not NOT1 (N3413, N3410);
nand NAND2 (N3414, N3411, N2519);
nor NOR3 (N3415, N3409, N1968, N2297);
xor XOR2 (N3416, N3400, N905);
not NOT1 (N3417, N3414);
or OR3 (N3418, N3416, N2903, N204);
or OR2 (N3419, N3418, N1692);
nor NOR4 (N3420, N3413, N2796, N687, N2085);
nand NAND2 (N3421, N3412, N1534);
xor XOR2 (N3422, N3408, N2020);
xor XOR2 (N3423, N3419, N2397);
buf BUF1 (N3424, N3407);
and AND4 (N3425, N3423, N1958, N2271, N3077);
not NOT1 (N3426, N3422);
nor NOR4 (N3427, N3394, N116, N1199, N3142);
nand NAND3 (N3428, N3387, N1880, N3347);
and AND3 (N3429, N3428, N1860, N2823);
and AND3 (N3430, N3389, N1228, N1763);
xor XOR2 (N3431, N3415, N1803);
and AND4 (N3432, N3417, N1503, N1690, N2902);
nor NOR2 (N3433, N3425, N2505);
buf BUF1 (N3434, N3427);
buf BUF1 (N3435, N3426);
nand NAND2 (N3436, N3431, N2879);
not NOT1 (N3437, N3429);
and AND2 (N3438, N3424, N68);
or OR4 (N3439, N3433, N1010, N3069, N787);
xor XOR2 (N3440, N3432, N2914);
buf BUF1 (N3441, N3436);
nand NAND4 (N3442, N3437, N2521, N2617, N663);
not NOT1 (N3443, N3438);
nor NOR3 (N3444, N3440, N2139, N2556);
nor NOR4 (N3445, N3421, N1565, N39, N1414);
buf BUF1 (N3446, N3443);
or OR4 (N3447, N3439, N2134, N2146, N890);
buf BUF1 (N3448, N3420);
xor XOR2 (N3449, N3444, N2139);
nor NOR2 (N3450, N3435, N3259);
nand NAND4 (N3451, N3448, N8, N2914, N887);
not NOT1 (N3452, N3449);
xor XOR2 (N3453, N3442, N1314);
not NOT1 (N3454, N3446);
or OR2 (N3455, N3454, N1018);
nor NOR4 (N3456, N3452, N227, N2921, N797);
or OR2 (N3457, N3441, N3222);
nor NOR4 (N3458, N3456, N3084, N2217, N2908);
nor NOR2 (N3459, N3447, N1070);
nand NAND4 (N3460, N3450, N877, N2494, N2805);
and AND3 (N3461, N3453, N1073, N2147);
buf BUF1 (N3462, N3458);
buf BUF1 (N3463, N3457);
nor NOR2 (N3464, N3455, N1271);
or OR4 (N3465, N3462, N979, N2164, N543);
not NOT1 (N3466, N3434);
and AND4 (N3467, N3465, N2928, N3268, N3174);
not NOT1 (N3468, N3461);
nor NOR2 (N3469, N3445, N1723);
and AND4 (N3470, N3467, N1963, N1836, N2686);
nand NAND2 (N3471, N3430, N1454);
nor NOR4 (N3472, N3464, N2825, N2693, N3211);
not NOT1 (N3473, N3472);
xor XOR2 (N3474, N3473, N2373);
nor NOR3 (N3475, N3474, N1685, N2452);
and AND2 (N3476, N3469, N801);
not NOT1 (N3477, N3470);
not NOT1 (N3478, N3476);
nor NOR2 (N3479, N3475, N465);
not NOT1 (N3480, N3466);
and AND4 (N3481, N3463, N3364, N2854, N2289);
nor NOR2 (N3482, N3477, N3430);
or OR2 (N3483, N3459, N1889);
not NOT1 (N3484, N3478);
buf BUF1 (N3485, N3482);
buf BUF1 (N3486, N3481);
xor XOR2 (N3487, N3485, N1318);
buf BUF1 (N3488, N3471);
buf BUF1 (N3489, N3451);
buf BUF1 (N3490, N3489);
and AND4 (N3491, N3480, N3063, N41, N2987);
xor XOR2 (N3492, N3491, N1603);
or OR4 (N3493, N3479, N2838, N1063, N1607);
nor NOR3 (N3494, N3483, N3186, N3155);
nand NAND4 (N3495, N3488, N2285, N746, N2175);
xor XOR2 (N3496, N3492, N672);
not NOT1 (N3497, N3468);
and AND2 (N3498, N3497, N2710);
and AND2 (N3499, N3490, N2843);
or OR3 (N3500, N3493, N524, N2474);
nor NOR2 (N3501, N3495, N2109);
nor NOR3 (N3502, N3487, N162, N1442);
nor NOR3 (N3503, N3501, N979, N1907);
nor NOR3 (N3504, N3486, N1911, N823);
nor NOR3 (N3505, N3460, N426, N1632);
and AND3 (N3506, N3503, N1139, N2696);
buf BUF1 (N3507, N3484);
buf BUF1 (N3508, N3498);
nor NOR2 (N3509, N3496, N1760);
nand NAND3 (N3510, N3506, N2320, N1167);
buf BUF1 (N3511, N3505);
nand NAND4 (N3512, N3511, N1109, N1222, N274);
xor XOR2 (N3513, N3509, N2110);
not NOT1 (N3514, N3508);
or OR4 (N3515, N3514, N3123, N3069, N219);
nor NOR3 (N3516, N3510, N1796, N1874);
xor XOR2 (N3517, N3500, N3095);
buf BUF1 (N3518, N3504);
or OR2 (N3519, N3516, N3065);
buf BUF1 (N3520, N3515);
nand NAND4 (N3521, N3512, N1669, N124, N3267);
or OR2 (N3522, N3502, N3269);
xor XOR2 (N3523, N3518, N1995);
nor NOR2 (N3524, N3521, N745);
and AND3 (N3525, N3507, N3404, N1869);
nor NOR3 (N3526, N3499, N1811, N2824);
nor NOR3 (N3527, N3513, N1321, N2782);
buf BUF1 (N3528, N3522);
or OR3 (N3529, N3519, N1368, N640);
buf BUF1 (N3530, N3526);
and AND2 (N3531, N3528, N1185);
nand NAND2 (N3532, N3520, N1220);
buf BUF1 (N3533, N3530);
nor NOR2 (N3534, N3532, N1595);
or OR2 (N3535, N3533, N2051);
and AND2 (N3536, N3523, N2475);
buf BUF1 (N3537, N3527);
or OR2 (N3538, N3534, N1464);
nor NOR4 (N3539, N3536, N960, N2899, N2607);
or OR2 (N3540, N3525, N168);
nand NAND4 (N3541, N3529, N2595, N2160, N2367);
or OR3 (N3542, N3539, N1643, N1619);
nor NOR2 (N3543, N3537, N2049);
or OR2 (N3544, N3531, N371);
nand NAND4 (N3545, N3494, N1831, N554, N1867);
and AND4 (N3546, N3543, N1788, N2290, N1925);
not NOT1 (N3547, N3517);
nor NOR2 (N3548, N3535, N2772);
not NOT1 (N3549, N3545);
not NOT1 (N3550, N3542);
and AND4 (N3551, N3549, N1979, N2281, N896);
nand NAND2 (N3552, N3547, N381);
or OR2 (N3553, N3550, N1956);
not NOT1 (N3554, N3551);
or OR2 (N3555, N3524, N474);
or OR4 (N3556, N3552, N1235, N1122, N286);
not NOT1 (N3557, N3544);
and AND4 (N3558, N3546, N2889, N713, N784);
or OR4 (N3559, N3557, N3258, N912, N1572);
and AND3 (N3560, N3553, N949, N3179);
buf BUF1 (N3561, N3541);
or OR3 (N3562, N3558, N2866, N1099);
not NOT1 (N3563, N3538);
and AND3 (N3564, N3554, N2823, N1760);
not NOT1 (N3565, N3540);
xor XOR2 (N3566, N3562, N2251);
or OR4 (N3567, N3556, N1188, N3412, N2097);
and AND2 (N3568, N3561, N2774);
and AND4 (N3569, N3555, N675, N1966, N1130);
and AND4 (N3570, N3568, N1939, N631, N2222);
or OR4 (N3571, N3548, N3094, N1726, N366);
nor NOR3 (N3572, N3571, N529, N3046);
nor NOR4 (N3573, N3560, N1782, N1061, N1383);
not NOT1 (N3574, N3565);
buf BUF1 (N3575, N3574);
nand NAND2 (N3576, N3563, N2421);
buf BUF1 (N3577, N3572);
buf BUF1 (N3578, N3569);
or OR3 (N3579, N3578, N261, N946);
nand NAND3 (N3580, N3564, N1987, N1404);
and AND4 (N3581, N3579, N2193, N615, N1617);
not NOT1 (N3582, N3575);
xor XOR2 (N3583, N3573, N22);
and AND3 (N3584, N3567, N3389, N2796);
nor NOR2 (N3585, N3570, N836);
buf BUF1 (N3586, N3580);
not NOT1 (N3587, N3559);
and AND3 (N3588, N3584, N1500, N762);
not NOT1 (N3589, N3577);
buf BUF1 (N3590, N3581);
nand NAND4 (N3591, N3589, N3549, N3221, N279);
buf BUF1 (N3592, N3566);
nor NOR4 (N3593, N3590, N3466, N835, N1974);
not NOT1 (N3594, N3591);
not NOT1 (N3595, N3594);
or OR2 (N3596, N3585, N582);
not NOT1 (N3597, N3596);
and AND4 (N3598, N3597, N1814, N840, N1809);
or OR4 (N3599, N3595, N1761, N916, N666);
xor XOR2 (N3600, N3582, N3020);
buf BUF1 (N3601, N3587);
not NOT1 (N3602, N3599);
buf BUF1 (N3603, N3602);
not NOT1 (N3604, N3588);
or OR4 (N3605, N3604, N1636, N960, N1257);
nor NOR4 (N3606, N3576, N3118, N1471, N3459);
not NOT1 (N3607, N3600);
and AND2 (N3608, N3603, N1246);
nor NOR2 (N3609, N3593, N3202);
nor NOR3 (N3610, N3601, N469, N2595);
not NOT1 (N3611, N3605);
not NOT1 (N3612, N3592);
buf BUF1 (N3613, N3609);
nor NOR2 (N3614, N3586, N2608);
nand NAND4 (N3615, N3612, N3476, N1525, N1649);
buf BUF1 (N3616, N3583);
not NOT1 (N3617, N3598);
xor XOR2 (N3618, N3617, N1560);
not NOT1 (N3619, N3610);
nand NAND2 (N3620, N3606, N338);
nand NAND4 (N3621, N3607, N2354, N735, N2029);
nor NOR3 (N3622, N3616, N1651, N609);
not NOT1 (N3623, N3613);
or OR3 (N3624, N3619, N2035, N2139);
nor NOR3 (N3625, N3614, N1248, N2061);
not NOT1 (N3626, N3625);
xor XOR2 (N3627, N3621, N3296);
not NOT1 (N3628, N3623);
or OR3 (N3629, N3627, N447, N2474);
and AND2 (N3630, N3608, N2038);
or OR4 (N3631, N3611, N1077, N1107, N1775);
and AND2 (N3632, N3615, N2813);
and AND3 (N3633, N3631, N1664, N628);
or OR4 (N3634, N3628, N749, N173, N136);
buf BUF1 (N3635, N3622);
nor NOR3 (N3636, N3632, N1448, N1861);
xor XOR2 (N3637, N3630, N912);
not NOT1 (N3638, N3634);
and AND2 (N3639, N3620, N260);
nand NAND2 (N3640, N3629, N2478);
or OR4 (N3641, N3638, N2476, N3299, N3603);
or OR4 (N3642, N3626, N2098, N1836, N617);
nand NAND3 (N3643, N3636, N1330, N445);
nand NAND2 (N3644, N3624, N595);
nor NOR2 (N3645, N3641, N1330);
not NOT1 (N3646, N3642);
and AND3 (N3647, N3643, N3521, N1063);
not NOT1 (N3648, N3635);
not NOT1 (N3649, N3637);
buf BUF1 (N3650, N3646);
xor XOR2 (N3651, N3640, N635);
xor XOR2 (N3652, N3648, N1848);
xor XOR2 (N3653, N3647, N1209);
nand NAND4 (N3654, N3633, N1497, N956, N1400);
buf BUF1 (N3655, N3650);
nand NAND3 (N3656, N3655, N2233, N2911);
and AND3 (N3657, N3652, N2785, N987);
nor NOR3 (N3658, N3618, N1063, N237);
not NOT1 (N3659, N3651);
not NOT1 (N3660, N3656);
buf BUF1 (N3661, N3654);
and AND3 (N3662, N3660, N2341, N1211);
nor NOR2 (N3663, N3639, N193);
and AND3 (N3664, N3663, N1159, N372);
xor XOR2 (N3665, N3661, N1201);
nor NOR2 (N3666, N3657, N2986);
nand NAND2 (N3667, N3653, N2056);
xor XOR2 (N3668, N3667, N1129);
nand NAND4 (N3669, N3645, N2884, N2270, N3098);
nand NAND3 (N3670, N3669, N1952, N3662);
buf BUF1 (N3671, N665);
and AND2 (N3672, N3649, N2136);
nand NAND2 (N3673, N3668, N2720);
nor NOR4 (N3674, N3670, N2946, N598, N474);
nor NOR3 (N3675, N3665, N1152, N2839);
nand NAND4 (N3676, N3644, N2101, N818, N8);
or OR4 (N3677, N3672, N327, N580, N665);
not NOT1 (N3678, N3671);
and AND2 (N3679, N3674, N328);
and AND4 (N3680, N3678, N1312, N1389, N831);
nand NAND2 (N3681, N3658, N1720);
and AND2 (N3682, N3681, N1069);
not NOT1 (N3683, N3675);
and AND2 (N3684, N3676, N1637);
and AND3 (N3685, N3677, N1092, N1111);
nor NOR2 (N3686, N3679, N2471);
buf BUF1 (N3687, N3682);
nand NAND2 (N3688, N3664, N2655);
nand NAND2 (N3689, N3659, N2759);
buf BUF1 (N3690, N3685);
nand NAND2 (N3691, N3680, N1180);
xor XOR2 (N3692, N3683, N1329);
not NOT1 (N3693, N3684);
or OR3 (N3694, N3692, N534, N1724);
xor XOR2 (N3695, N3693, N1237);
xor XOR2 (N3696, N3691, N1515);
xor XOR2 (N3697, N3689, N1798);
and AND3 (N3698, N3688, N260, N2446);
xor XOR2 (N3699, N3686, N1076);
or OR3 (N3700, N3694, N3249, N714);
buf BUF1 (N3701, N3699);
xor XOR2 (N3702, N3687, N3279);
and AND2 (N3703, N3695, N3526);
and AND2 (N3704, N3697, N221);
nand NAND2 (N3705, N3702, N2008);
not NOT1 (N3706, N3673);
and AND4 (N3707, N3704, N2468, N2937, N1707);
and AND2 (N3708, N3696, N2969);
xor XOR2 (N3709, N3690, N2226);
nand NAND3 (N3710, N3703, N51, N2464);
and AND3 (N3711, N3706, N2450, N825);
nand NAND2 (N3712, N3666, N1656);
buf BUF1 (N3713, N3710);
buf BUF1 (N3714, N3712);
not NOT1 (N3715, N3714);
buf BUF1 (N3716, N3707);
xor XOR2 (N3717, N3715, N1304);
nor NOR2 (N3718, N3713, N2059);
buf BUF1 (N3719, N3711);
nand NAND2 (N3720, N3700, N1949);
and AND2 (N3721, N3716, N2473);
or OR3 (N3722, N3718, N2135, N79);
nor NOR3 (N3723, N3720, N2082, N2926);
nand NAND3 (N3724, N3709, N2458, N3719);
not NOT1 (N3725, N1525);
nor NOR2 (N3726, N3708, N1989);
xor XOR2 (N3727, N3705, N1767);
and AND3 (N3728, N3724, N2395, N2328);
xor XOR2 (N3729, N3723, N1732);
buf BUF1 (N3730, N3725);
not NOT1 (N3731, N3726);
or OR3 (N3732, N3721, N3721, N2274);
and AND3 (N3733, N3729, N3319, N2572);
not NOT1 (N3734, N3730);
not NOT1 (N3735, N3701);
and AND3 (N3736, N3735, N2936, N2246);
and AND3 (N3737, N3733, N3196, N2047);
not NOT1 (N3738, N3728);
and AND2 (N3739, N3738, N2195);
not NOT1 (N3740, N3722);
not NOT1 (N3741, N3734);
nor NOR3 (N3742, N3741, N2059, N3381);
and AND2 (N3743, N3737, N172);
nor NOR2 (N3744, N3739, N2241);
and AND4 (N3745, N3731, N1087, N702, N1471);
not NOT1 (N3746, N3736);
and AND4 (N3747, N3717, N3130, N2252, N350);
or OR4 (N3748, N3732, N612, N1743, N2162);
nor NOR2 (N3749, N3742, N3633);
buf BUF1 (N3750, N3698);
nand NAND2 (N3751, N3727, N3279);
nor NOR4 (N3752, N3744, N1350, N898, N3249);
not NOT1 (N3753, N3743);
nand NAND3 (N3754, N3740, N3352, N2403);
or OR3 (N3755, N3748, N3209, N688);
xor XOR2 (N3756, N3745, N989);
not NOT1 (N3757, N3751);
buf BUF1 (N3758, N3753);
xor XOR2 (N3759, N3752, N2991);
xor XOR2 (N3760, N3757, N2205);
buf BUF1 (N3761, N3747);
xor XOR2 (N3762, N3760, N694);
xor XOR2 (N3763, N3755, N1727);
buf BUF1 (N3764, N3761);
xor XOR2 (N3765, N3758, N2965);
not NOT1 (N3766, N3746);
nor NOR4 (N3767, N3749, N2046, N1203, N1443);
buf BUF1 (N3768, N3754);
buf BUF1 (N3769, N3763);
xor XOR2 (N3770, N3768, N2193);
nor NOR3 (N3771, N3770, N2153, N741);
nor NOR4 (N3772, N3764, N3437, N2692, N507);
or OR4 (N3773, N3771, N3019, N3000, N1531);
or OR4 (N3774, N3772, N938, N1599, N2724);
nor NOR2 (N3775, N3750, N2778);
nand NAND4 (N3776, N3769, N3674, N1088, N2229);
nor NOR2 (N3777, N3773, N2941);
and AND4 (N3778, N3767, N2937, N2984, N2818);
xor XOR2 (N3779, N3778, N1599);
or OR2 (N3780, N3774, N3472);
not NOT1 (N3781, N3780);
not NOT1 (N3782, N3781);
or OR2 (N3783, N3777, N39);
xor XOR2 (N3784, N3756, N1795);
and AND2 (N3785, N3776, N1589);
buf BUF1 (N3786, N3784);
xor XOR2 (N3787, N3765, N12);
or OR4 (N3788, N3775, N2994, N3406, N1707);
buf BUF1 (N3789, N3786);
xor XOR2 (N3790, N3766, N385);
xor XOR2 (N3791, N3785, N1249);
not NOT1 (N3792, N3789);
not NOT1 (N3793, N3779);
or OR4 (N3794, N3782, N988, N3592, N2325);
buf BUF1 (N3795, N3762);
buf BUF1 (N3796, N3788);
or OR3 (N3797, N3795, N274, N655);
nand NAND4 (N3798, N3790, N3318, N2274, N3328);
and AND4 (N3799, N3791, N1356, N1621, N1244);
buf BUF1 (N3800, N3787);
or OR4 (N3801, N3798, N2591, N1613, N2788);
nand NAND2 (N3802, N3792, N3379);
buf BUF1 (N3803, N3783);
and AND2 (N3804, N3794, N998);
xor XOR2 (N3805, N3801, N1389);
buf BUF1 (N3806, N3802);
not NOT1 (N3807, N3799);
not NOT1 (N3808, N3759);
not NOT1 (N3809, N3808);
xor XOR2 (N3810, N3796, N1573);
nor NOR4 (N3811, N3806, N3779, N2740, N3661);
xor XOR2 (N3812, N3803, N3181);
or OR3 (N3813, N3793, N1251, N2348);
nand NAND3 (N3814, N3813, N912, N1613);
nor NOR2 (N3815, N3804, N612);
or OR4 (N3816, N3812, N322, N51, N2637);
xor XOR2 (N3817, N3815, N716);
nor NOR4 (N3818, N3816, N570, N1804, N3150);
or OR3 (N3819, N3814, N177, N464);
xor XOR2 (N3820, N3818, N3187);
and AND3 (N3821, N3807, N1036, N1255);
not NOT1 (N3822, N3811);
nor NOR3 (N3823, N3805, N306, N2587);
buf BUF1 (N3824, N3797);
not NOT1 (N3825, N3809);
nor NOR3 (N3826, N3822, N1503, N1467);
buf BUF1 (N3827, N3810);
nor NOR2 (N3828, N3824, N2735);
or OR4 (N3829, N3817, N2501, N2542, N2693);
xor XOR2 (N3830, N3819, N2754);
nand NAND2 (N3831, N3821, N120);
and AND2 (N3832, N3830, N2764);
or OR4 (N3833, N3820, N3648, N985, N341);
buf BUF1 (N3834, N3825);
nand NAND4 (N3835, N3826, N3055, N1984, N1088);
nor NOR2 (N3836, N3833, N3512);
nor NOR2 (N3837, N3827, N3075);
nor NOR2 (N3838, N3823, N2062);
xor XOR2 (N3839, N3832, N3347);
xor XOR2 (N3840, N3836, N1759);
nor NOR2 (N3841, N3831, N460);
or OR2 (N3842, N3828, N3236);
and AND2 (N3843, N3841, N927);
nand NAND4 (N3844, N3834, N2745, N1981, N1248);
xor XOR2 (N3845, N3838, N2860);
nor NOR3 (N3846, N3800, N414, N3593);
xor XOR2 (N3847, N3846, N2690);
and AND2 (N3848, N3844, N3028);
or OR3 (N3849, N3835, N811, N541);
and AND3 (N3850, N3837, N1627, N2347);
xor XOR2 (N3851, N3849, N2);
xor XOR2 (N3852, N3850, N2203);
xor XOR2 (N3853, N3842, N199);
and AND3 (N3854, N3839, N1381, N3155);
and AND4 (N3855, N3829, N1141, N3342, N611);
xor XOR2 (N3856, N3847, N3044);
buf BUF1 (N3857, N3855);
nand NAND4 (N3858, N3852, N1097, N465, N326);
buf BUF1 (N3859, N3851);
or OR3 (N3860, N3854, N1077, N2433);
nor NOR4 (N3861, N3857, N3091, N2003, N1520);
or OR4 (N3862, N3859, N2964, N674, N1779);
and AND3 (N3863, N3858, N389, N2939);
nor NOR2 (N3864, N3860, N1965);
not NOT1 (N3865, N3863);
xor XOR2 (N3866, N3862, N1642);
nand NAND2 (N3867, N3840, N2528);
not NOT1 (N3868, N3866);
and AND2 (N3869, N3861, N2853);
and AND3 (N3870, N3853, N1371, N784);
not NOT1 (N3871, N3843);
not NOT1 (N3872, N3868);
nand NAND3 (N3873, N3867, N1832, N1988);
buf BUF1 (N3874, N3856);
nor NOR4 (N3875, N3864, N3368, N1068, N3236);
nor NOR4 (N3876, N3874, N2565, N2113, N2011);
nor NOR4 (N3877, N3869, N919, N929, N2661);
not NOT1 (N3878, N3873);
and AND2 (N3879, N3871, N2211);
nor NOR2 (N3880, N3872, N1329);
and AND4 (N3881, N3875, N470, N1897, N3449);
nor NOR3 (N3882, N3876, N2112, N3039);
not NOT1 (N3883, N3877);
or OR2 (N3884, N3883, N3514);
nor NOR3 (N3885, N3884, N683, N1948);
and AND4 (N3886, N3878, N812, N3577, N1823);
and AND2 (N3887, N3881, N1179);
or OR3 (N3888, N3887, N2864, N356);
or OR2 (N3889, N3882, N2682);
buf BUF1 (N3890, N3865);
not NOT1 (N3891, N3888);
xor XOR2 (N3892, N3848, N213);
nand NAND2 (N3893, N3885, N2973);
buf BUF1 (N3894, N3891);
and AND2 (N3895, N3845, N2665);
or OR3 (N3896, N3886, N3049, N3758);
nor NOR2 (N3897, N3893, N721);
nor NOR3 (N3898, N3890, N3077, N559);
or OR2 (N3899, N3892, N1701);
nand NAND2 (N3900, N3879, N2434);
or OR4 (N3901, N3895, N2126, N3394, N3594);
and AND4 (N3902, N3897, N2296, N2749, N1538);
nand NAND3 (N3903, N3899, N1804, N459);
and AND4 (N3904, N3902, N2718, N3751, N698);
and AND2 (N3905, N3904, N711);
or OR3 (N3906, N3901, N1671, N433);
and AND2 (N3907, N3898, N2698);
and AND3 (N3908, N3905, N3152, N3848);
and AND3 (N3909, N3896, N3760, N3358);
not NOT1 (N3910, N3907);
nor NOR2 (N3911, N3880, N1876);
and AND3 (N3912, N3906, N347, N3119);
not NOT1 (N3913, N3908);
buf BUF1 (N3914, N3911);
nor NOR3 (N3915, N3894, N1890, N2608);
buf BUF1 (N3916, N3903);
or OR3 (N3917, N3909, N3582, N426);
not NOT1 (N3918, N3889);
not NOT1 (N3919, N3917);
xor XOR2 (N3920, N3918, N898);
not NOT1 (N3921, N3915);
buf BUF1 (N3922, N3912);
xor XOR2 (N3923, N3919, N1820);
xor XOR2 (N3924, N3910, N1756);
or OR2 (N3925, N3924, N3786);
xor XOR2 (N3926, N3921, N3739);
nand NAND3 (N3927, N3916, N36, N1071);
buf BUF1 (N3928, N3927);
buf BUF1 (N3929, N3920);
and AND4 (N3930, N3925, N1154, N1237, N1063);
nor NOR3 (N3931, N3914, N2719, N1907);
not NOT1 (N3932, N3913);
nand NAND3 (N3933, N3932, N1979, N3698);
nor NOR2 (N3934, N3922, N2716);
xor XOR2 (N3935, N3930, N1139);
or OR3 (N3936, N3929, N413, N2407);
or OR3 (N3937, N3923, N1804, N290);
and AND3 (N3938, N3935, N3443, N661);
buf BUF1 (N3939, N3936);
buf BUF1 (N3940, N3937);
or OR2 (N3941, N3934, N3758);
buf BUF1 (N3942, N3933);
not NOT1 (N3943, N3939);
or OR3 (N3944, N3900, N1447, N316);
nand NAND4 (N3945, N3943, N2268, N1622, N1002);
buf BUF1 (N3946, N3928);
xor XOR2 (N3947, N3938, N1304);
not NOT1 (N3948, N3931);
or OR2 (N3949, N3941, N2768);
and AND3 (N3950, N3945, N2479, N1656);
or OR3 (N3951, N3940, N1287, N2037);
or OR3 (N3952, N3926, N116, N60);
buf BUF1 (N3953, N3947);
or OR2 (N3954, N3952, N1790);
buf BUF1 (N3955, N3870);
nand NAND3 (N3956, N3942, N2132, N541);
nor NOR2 (N3957, N3953, N71);
and AND4 (N3958, N3951, N2604, N3607, N2416);
and AND2 (N3959, N3954, N1957);
nand NAND2 (N3960, N3959, N2963);
or OR3 (N3961, N3944, N3331, N2937);
or OR4 (N3962, N3961, N1662, N2975, N3411);
buf BUF1 (N3963, N3960);
xor XOR2 (N3964, N3949, N2463);
nor NOR3 (N3965, N3946, N987, N3234);
xor XOR2 (N3966, N3957, N2569);
xor XOR2 (N3967, N3966, N1402);
buf BUF1 (N3968, N3948);
not NOT1 (N3969, N3963);
nor NOR2 (N3970, N3950, N390);
xor XOR2 (N3971, N3955, N1643);
nand NAND3 (N3972, N3971, N3776, N3785);
xor XOR2 (N3973, N3968, N1379);
nor NOR4 (N3974, N3964, N1904, N729, N2362);
nand NAND2 (N3975, N3962, N1273);
not NOT1 (N3976, N3958);
xor XOR2 (N3977, N3956, N419);
or OR4 (N3978, N3969, N1235, N3668, N1148);
not NOT1 (N3979, N3975);
buf BUF1 (N3980, N3976);
buf BUF1 (N3981, N3979);
xor XOR2 (N3982, N3972, N507);
not NOT1 (N3983, N3970);
not NOT1 (N3984, N3982);
buf BUF1 (N3985, N3978);
or OR4 (N3986, N3973, N3448, N1827, N787);
nand NAND4 (N3987, N3984, N3662, N2110, N3590);
xor XOR2 (N3988, N3974, N2504);
nand NAND4 (N3989, N3986, N2456, N2870, N921);
nand NAND3 (N3990, N3980, N2889, N3371);
buf BUF1 (N3991, N3983);
and AND2 (N3992, N3977, N1427);
nor NOR3 (N3993, N3987, N774, N3402);
or OR3 (N3994, N3989, N2852, N81);
not NOT1 (N3995, N3988);
or OR3 (N3996, N3994, N2537, N1347);
nor NOR4 (N3997, N3995, N3715, N1499, N2703);
xor XOR2 (N3998, N3997, N3096);
not NOT1 (N3999, N3992);
xor XOR2 (N4000, N3999, N2715);
not NOT1 (N4001, N3967);
and AND4 (N4002, N4001, N1868, N996, N1552);
not NOT1 (N4003, N4002);
or OR3 (N4004, N3996, N3482, N1806);
buf BUF1 (N4005, N3993);
nor NOR2 (N4006, N3985, N114);
xor XOR2 (N4007, N4005, N1975);
nand NAND2 (N4008, N3990, N1914);
nand NAND3 (N4009, N3965, N3864, N220);
nor NOR4 (N4010, N4006, N1003, N2469, N52);
nand NAND2 (N4011, N4009, N1320);
or OR2 (N4012, N4000, N3396);
xor XOR2 (N4013, N4004, N40);
not NOT1 (N4014, N4012);
nor NOR4 (N4015, N3998, N3462, N1567, N3331);
and AND3 (N4016, N3991, N1748, N346);
buf BUF1 (N4017, N3981);
or OR3 (N4018, N4003, N2118, N1474);
buf BUF1 (N4019, N4015);
or OR4 (N4020, N4016, N410, N2567, N1447);
nand NAND2 (N4021, N4018, N3389);
nand NAND3 (N4022, N4019, N2194, N684);
buf BUF1 (N4023, N4010);
nor NOR2 (N4024, N4020, N1951);
nor NOR2 (N4025, N4008, N1121);
or OR2 (N4026, N4025, N253);
or OR2 (N4027, N4024, N763);
xor XOR2 (N4028, N4017, N1577);
xor XOR2 (N4029, N4027, N906);
buf BUF1 (N4030, N4021);
not NOT1 (N4031, N4007);
xor XOR2 (N4032, N4013, N1215);
nor NOR2 (N4033, N4030, N2353);
and AND4 (N4034, N4032, N2929, N2608, N3612);
or OR4 (N4035, N4026, N3478, N2561, N3169);
and AND3 (N4036, N4028, N1070, N2225);
xor XOR2 (N4037, N4033, N2843);
nor NOR4 (N4038, N4014, N3148, N1749, N2984);
nand NAND2 (N4039, N4036, N1379);
not NOT1 (N4040, N4011);
xor XOR2 (N4041, N4037, N1314);
or OR2 (N4042, N4029, N3465);
xor XOR2 (N4043, N4035, N1084);
and AND3 (N4044, N4039, N1008, N2837);
not NOT1 (N4045, N4031);
nand NAND3 (N4046, N4040, N2175, N3217);
and AND2 (N4047, N4038, N1226);
and AND2 (N4048, N4045, N2646);
xor XOR2 (N4049, N4042, N193);
nand NAND4 (N4050, N4034, N1262, N1903, N1325);
nor NOR3 (N4051, N4041, N402, N3018);
nand NAND4 (N4052, N4046, N1545, N2067, N2450);
or OR2 (N4053, N4049, N634);
xor XOR2 (N4054, N4023, N2160);
nor NOR4 (N4055, N4054, N2712, N279, N1567);
and AND2 (N4056, N4047, N3521);
nor NOR4 (N4057, N4051, N3422, N318, N3601);
nand NAND3 (N4058, N4055, N22, N2614);
xor XOR2 (N4059, N4056, N1052);
buf BUF1 (N4060, N4048);
and AND2 (N4061, N4050, N2897);
or OR3 (N4062, N4058, N2929, N3982);
nor NOR3 (N4063, N4053, N1170, N838);
not NOT1 (N4064, N4043);
or OR2 (N4065, N4044, N2762);
nor NOR2 (N4066, N4062, N1854);
or OR2 (N4067, N4057, N1813);
and AND3 (N4068, N4065, N3849, N2285);
nor NOR4 (N4069, N4052, N1066, N3635, N3638);
buf BUF1 (N4070, N4059);
buf BUF1 (N4071, N4068);
or OR3 (N4072, N4070, N1749, N2923);
nor NOR4 (N4073, N4022, N3377, N1420, N787);
nand NAND4 (N4074, N4071, N729, N100, N1083);
buf BUF1 (N4075, N4063);
xor XOR2 (N4076, N4066, N2889);
or OR3 (N4077, N4067, N1989, N1343);
and AND3 (N4078, N4074, N1605, N2703);
or OR3 (N4079, N4061, N2178, N4013);
and AND2 (N4080, N4076, N2378);
nor NOR2 (N4081, N4077, N3613);
or OR2 (N4082, N4075, N684);
buf BUF1 (N4083, N4082);
buf BUF1 (N4084, N4060);
not NOT1 (N4085, N4084);
and AND4 (N4086, N4069, N2963, N1465, N750);
nand NAND4 (N4087, N4064, N47, N2261, N484);
nand NAND3 (N4088, N4080, N172, N639);
buf BUF1 (N4089, N4087);
and AND2 (N4090, N4073, N1141);
or OR3 (N4091, N4083, N604, N1627);
buf BUF1 (N4092, N4089);
nor NOR2 (N4093, N4090, N1806);
xor XOR2 (N4094, N4093, N2999);
not NOT1 (N4095, N4081);
nor NOR3 (N4096, N4095, N2484, N555);
and AND2 (N4097, N4086, N1890);
xor XOR2 (N4098, N4085, N1486);
buf BUF1 (N4099, N4092);
nor NOR2 (N4100, N4096, N368);
and AND2 (N4101, N4094, N506);
not NOT1 (N4102, N4091);
xor XOR2 (N4103, N4102, N2240);
nand NAND2 (N4104, N4099, N242);
nor NOR4 (N4105, N4101, N3044, N3697, N2266);
xor XOR2 (N4106, N4100, N1476);
nor NOR2 (N4107, N4105, N2785);
or OR2 (N4108, N4107, N3103);
or OR2 (N4109, N4079, N1182);
and AND4 (N4110, N4103, N2843, N404, N4007);
nand NAND2 (N4111, N4098, N2684);
buf BUF1 (N4112, N4109);
nor NOR2 (N4113, N4072, N3100);
buf BUF1 (N4114, N4097);
nand NAND3 (N4115, N4078, N1201, N2675);
xor XOR2 (N4116, N4112, N1055);
nand NAND2 (N4117, N4106, N3999);
or OR3 (N4118, N4113, N4115, N1315);
nand NAND2 (N4119, N1847, N2411);
xor XOR2 (N4120, N4110, N4079);
buf BUF1 (N4121, N4088);
and AND2 (N4122, N4118, N1529);
not NOT1 (N4123, N4104);
or OR2 (N4124, N4119, N871);
nor NOR3 (N4125, N4121, N699, N2105);
not NOT1 (N4126, N4125);
not NOT1 (N4127, N4116);
not NOT1 (N4128, N4117);
nand NAND2 (N4129, N4127, N3647);
nand NAND4 (N4130, N4108, N322, N157, N1153);
not NOT1 (N4131, N4124);
nor NOR4 (N4132, N4123, N994, N3646, N2746);
xor XOR2 (N4133, N4122, N2550);
and AND2 (N4134, N4129, N2375);
buf BUF1 (N4135, N4126);
nor NOR3 (N4136, N4114, N877, N660);
and AND2 (N4137, N4132, N2093);
and AND3 (N4138, N4130, N1304, N710);
xor XOR2 (N4139, N4131, N4076);
nor NOR3 (N4140, N4137, N892, N198);
buf BUF1 (N4141, N4135);
nor NOR4 (N4142, N4120, N1443, N2669, N2187);
nand NAND4 (N4143, N4134, N1686, N3708, N3769);
and AND3 (N4144, N4138, N2062, N1782);
nor NOR3 (N4145, N4128, N2960, N2952);
nor NOR4 (N4146, N4140, N2750, N2019, N2770);
and AND3 (N4147, N4146, N743, N1944);
not NOT1 (N4148, N4136);
not NOT1 (N4149, N4142);
xor XOR2 (N4150, N4133, N303);
or OR2 (N4151, N4111, N498);
not NOT1 (N4152, N4141);
or OR4 (N4153, N4148, N4034, N1946, N3799);
buf BUF1 (N4154, N4145);
xor XOR2 (N4155, N4152, N1796);
nand NAND3 (N4156, N4147, N2401, N2956);
xor XOR2 (N4157, N4151, N4086);
nor NOR4 (N4158, N4143, N3061, N945, N1211);
nand NAND4 (N4159, N4158, N344, N639, N820);
buf BUF1 (N4160, N4139);
xor XOR2 (N4161, N4155, N677);
xor XOR2 (N4162, N4150, N3345);
not NOT1 (N4163, N4156);
or OR4 (N4164, N4144, N4090, N3578, N2499);
buf BUF1 (N4165, N4157);
xor XOR2 (N4166, N4162, N1854);
nor NOR3 (N4167, N4166, N3262, N326);
and AND2 (N4168, N4167, N4155);
xor XOR2 (N4169, N4153, N2735);
and AND4 (N4170, N4163, N840, N2703, N3614);
nand NAND4 (N4171, N4168, N1259, N1607, N4160);
and AND4 (N4172, N763, N322, N901, N3308);
nand NAND3 (N4173, N4154, N1985, N1655);
and AND4 (N4174, N4159, N2204, N3563, N3954);
buf BUF1 (N4175, N4172);
and AND2 (N4176, N4165, N1628);
xor XOR2 (N4177, N4170, N113);
not NOT1 (N4178, N4149);
and AND4 (N4179, N4169, N2887, N1494, N577);
not NOT1 (N4180, N4164);
not NOT1 (N4181, N4174);
xor XOR2 (N4182, N4181, N2338);
nand NAND2 (N4183, N4176, N4083);
xor XOR2 (N4184, N4178, N4182);
buf BUF1 (N4185, N2302);
xor XOR2 (N4186, N4177, N4074);
not NOT1 (N4187, N4183);
nor NOR4 (N4188, N4175, N3553, N1711, N580);
and AND3 (N4189, N4179, N675, N2984);
xor XOR2 (N4190, N4184, N574);
xor XOR2 (N4191, N4186, N1587);
and AND2 (N4192, N4188, N3821);
not NOT1 (N4193, N4187);
not NOT1 (N4194, N4192);
and AND4 (N4195, N4173, N3583, N1691, N1788);
nor NOR4 (N4196, N4171, N1442, N1427, N2962);
or OR3 (N4197, N4191, N1384, N1055);
or OR3 (N4198, N4180, N1225, N2926);
or OR3 (N4199, N4189, N2190, N36);
nor NOR2 (N4200, N4185, N2492);
not NOT1 (N4201, N4194);
nand NAND3 (N4202, N4196, N482, N4177);
and AND2 (N4203, N4197, N1856);
and AND3 (N4204, N4202, N1163, N2981);
and AND3 (N4205, N4193, N2381, N4146);
nor NOR3 (N4206, N4161, N2542, N2254);
or OR3 (N4207, N4205, N2724, N4101);
or OR2 (N4208, N4195, N3494);
xor XOR2 (N4209, N4198, N3561);
nor NOR4 (N4210, N4209, N2007, N829, N3220);
nand NAND4 (N4211, N4210, N1722, N3123, N1889);
nand NAND3 (N4212, N4208, N4155, N353);
or OR4 (N4213, N4204, N3489, N3993, N1620);
and AND4 (N4214, N4207, N2545, N3086, N730);
not NOT1 (N4215, N4214);
and AND4 (N4216, N4206, N26, N3539, N1155);
nand NAND3 (N4217, N4201, N2547, N2);
and AND2 (N4218, N4215, N681);
and AND4 (N4219, N4212, N4119, N2444, N913);
or OR3 (N4220, N4200, N2748, N1279);
or OR4 (N4221, N4213, N4122, N846, N2595);
xor XOR2 (N4222, N4211, N3159);
nand NAND4 (N4223, N4221, N3003, N1509, N2264);
not NOT1 (N4224, N4217);
buf BUF1 (N4225, N4218);
xor XOR2 (N4226, N4203, N2938);
buf BUF1 (N4227, N4199);
not NOT1 (N4228, N4222);
and AND4 (N4229, N4225, N181, N1942, N2060);
or OR2 (N4230, N4224, N2737);
nand NAND4 (N4231, N4220, N1825, N2500, N1891);
and AND2 (N4232, N4219, N3930);
buf BUF1 (N4233, N4230);
nor NOR3 (N4234, N4223, N1451, N3632);
xor XOR2 (N4235, N4229, N2619);
and AND4 (N4236, N4232, N3885, N2808, N2380);
buf BUF1 (N4237, N4235);
buf BUF1 (N4238, N4233);
not NOT1 (N4239, N4228);
and AND2 (N4240, N4231, N1730);
nand NAND4 (N4241, N4227, N2741, N15, N3647);
nand NAND2 (N4242, N4190, N789);
nor NOR3 (N4243, N4216, N1732, N1487);
nand NAND3 (N4244, N4240, N3600, N3069);
nor NOR2 (N4245, N4239, N1470);
nand NAND3 (N4246, N4238, N802, N3132);
nor NOR2 (N4247, N4237, N473);
and AND3 (N4248, N4247, N3282, N3878);
buf BUF1 (N4249, N4248);
buf BUF1 (N4250, N4243);
nand NAND3 (N4251, N4250, N3933, N468);
buf BUF1 (N4252, N4245);
nand NAND4 (N4253, N4246, N3771, N2980, N2033);
xor XOR2 (N4254, N4234, N1130);
nor NOR2 (N4255, N4252, N2364);
and AND3 (N4256, N4251, N3561, N265);
nor NOR2 (N4257, N4226, N84);
or OR2 (N4258, N4256, N2637);
nor NOR3 (N4259, N4241, N2539, N2686);
xor XOR2 (N4260, N4242, N922);
or OR2 (N4261, N4259, N1024);
not NOT1 (N4262, N4257);
xor XOR2 (N4263, N4255, N2837);
nand NAND2 (N4264, N4262, N1242);
and AND2 (N4265, N4260, N736);
not NOT1 (N4266, N4264);
nand NAND2 (N4267, N4266, N254);
not NOT1 (N4268, N4244);
or OR2 (N4269, N4265, N281);
nand NAND4 (N4270, N4258, N507, N2126, N1480);
and AND2 (N4271, N4253, N522);
xor XOR2 (N4272, N4254, N1918);
not NOT1 (N4273, N4261);
and AND4 (N4274, N4268, N949, N3396, N54);
nor NOR4 (N4275, N4267, N2287, N2295, N3054);
not NOT1 (N4276, N4269);
buf BUF1 (N4277, N4276);
and AND3 (N4278, N4273, N1004, N3136);
and AND3 (N4279, N4275, N846, N3374);
xor XOR2 (N4280, N4278, N2739);
and AND2 (N4281, N4263, N580);
nand NAND4 (N4282, N4274, N2313, N636, N46);
or OR3 (N4283, N4282, N3024, N1640);
nand NAND3 (N4284, N4271, N1311, N2828);
nor NOR3 (N4285, N4284, N1369, N2591);
not NOT1 (N4286, N4279);
buf BUF1 (N4287, N4283);
or OR4 (N4288, N4272, N4145, N3531, N635);
or OR2 (N4289, N4281, N221);
nor NOR3 (N4290, N4288, N3117, N3557);
not NOT1 (N4291, N4289);
nand NAND2 (N4292, N4236, N2305);
or OR4 (N4293, N4290, N390, N2765, N3719);
nand NAND3 (N4294, N4277, N3736, N2872);
and AND4 (N4295, N4291, N2270, N1220, N92);
not NOT1 (N4296, N4293);
buf BUF1 (N4297, N4292);
not NOT1 (N4298, N4285);
buf BUF1 (N4299, N4286);
not NOT1 (N4300, N4294);
nor NOR3 (N4301, N4297, N3652, N387);
not NOT1 (N4302, N4287);
and AND4 (N4303, N4280, N1432, N3530, N1084);
or OR3 (N4304, N4302, N275, N3369);
and AND3 (N4305, N4298, N1863, N4075);
not NOT1 (N4306, N4295);
not NOT1 (N4307, N4303);
or OR2 (N4308, N4306, N4048);
or OR3 (N4309, N4305, N3145, N2222);
xor XOR2 (N4310, N4249, N2377);
nor NOR4 (N4311, N4301, N1736, N191, N1026);
xor XOR2 (N4312, N4307, N703);
not NOT1 (N4313, N4311);
not NOT1 (N4314, N4270);
xor XOR2 (N4315, N4308, N3695);
and AND2 (N4316, N4300, N803);
nor NOR4 (N4317, N4316, N4243, N283, N3968);
nand NAND2 (N4318, N4313, N249);
buf BUF1 (N4319, N4304);
nor NOR4 (N4320, N4309, N2674, N3367, N786);
not NOT1 (N4321, N4319);
nor NOR4 (N4322, N4310, N2074, N2650, N2667);
xor XOR2 (N4323, N4322, N824);
nor NOR4 (N4324, N4321, N22, N2937, N2255);
buf BUF1 (N4325, N4312);
nand NAND3 (N4326, N4324, N2090, N929);
xor XOR2 (N4327, N4323, N3526);
nand NAND2 (N4328, N4299, N639);
nand NAND2 (N4329, N4317, N1792);
buf BUF1 (N4330, N4325);
not NOT1 (N4331, N4315);
nand NAND2 (N4332, N4296, N392);
xor XOR2 (N4333, N4330, N622);
not NOT1 (N4334, N4318);
nor NOR3 (N4335, N4327, N3860, N3050);
nor NOR2 (N4336, N4320, N3400);
not NOT1 (N4337, N4328);
nand NAND3 (N4338, N4337, N1992, N2762);
xor XOR2 (N4339, N4334, N397);
xor XOR2 (N4340, N4339, N751);
xor XOR2 (N4341, N4333, N2575);
and AND2 (N4342, N4331, N4048);
or OR3 (N4343, N4329, N1517, N2244);
nand NAND3 (N4344, N4343, N4295, N3238);
nor NOR3 (N4345, N4344, N3843, N1485);
nor NOR2 (N4346, N4342, N3361);
or OR3 (N4347, N4314, N2676, N1050);
and AND3 (N4348, N4338, N3914, N846);
and AND3 (N4349, N4340, N4320, N4020);
or OR2 (N4350, N4347, N1285);
nor NOR3 (N4351, N4349, N202, N2226);
nor NOR3 (N4352, N4341, N2028, N2061);
xor XOR2 (N4353, N4326, N3586);
nor NOR2 (N4354, N4336, N1569);
xor XOR2 (N4355, N4352, N3128);
and AND4 (N4356, N4351, N3099, N1079, N2028);
nor NOR2 (N4357, N4345, N4210);
xor XOR2 (N4358, N4332, N1733);
nor NOR3 (N4359, N4358, N2547, N1053);
xor XOR2 (N4360, N4335, N1235);
xor XOR2 (N4361, N4357, N2012);
nor NOR4 (N4362, N4346, N1972, N3142, N2321);
nor NOR3 (N4363, N4360, N1610, N4108);
xor XOR2 (N4364, N4348, N3639);
and AND3 (N4365, N4354, N2486, N3514);
xor XOR2 (N4366, N4363, N2386);
xor XOR2 (N4367, N4365, N3598);
not NOT1 (N4368, N4366);
or OR2 (N4369, N4367, N1647);
xor XOR2 (N4370, N4356, N3002);
and AND2 (N4371, N4355, N3745);
nand NAND4 (N4372, N4359, N1747, N1295, N879);
nor NOR2 (N4373, N4361, N1682);
nand NAND2 (N4374, N4371, N3536);
xor XOR2 (N4375, N4369, N3707);
nor NOR3 (N4376, N4350, N1964, N1359);
nor NOR4 (N4377, N4376, N1270, N1357, N4257);
nor NOR2 (N4378, N4374, N2118);
xor XOR2 (N4379, N4373, N2416);
and AND2 (N4380, N4362, N341);
xor XOR2 (N4381, N4353, N2981);
buf BUF1 (N4382, N4378);
nand NAND4 (N4383, N4364, N4252, N1482, N3648);
xor XOR2 (N4384, N4383, N330);
or OR4 (N4385, N4381, N2491, N3914, N176);
or OR3 (N4386, N4385, N1245, N4200);
and AND2 (N4387, N4375, N2736);
buf BUF1 (N4388, N4384);
nand NAND3 (N4389, N4380, N2558, N3619);
nand NAND4 (N4390, N4370, N1231, N4317, N2708);
nand NAND3 (N4391, N4390, N4308, N1866);
nand NAND4 (N4392, N4386, N1594, N1548, N4095);
or OR3 (N4393, N4379, N3599, N289);
nand NAND4 (N4394, N4382, N436, N1770, N213);
nor NOR3 (N4395, N4392, N1259, N2924);
nor NOR4 (N4396, N4394, N2292, N2424, N2975);
buf BUF1 (N4397, N4389);
and AND4 (N4398, N4377, N1101, N3913, N106);
not NOT1 (N4399, N4391);
xor XOR2 (N4400, N4387, N2019);
nand NAND3 (N4401, N4368, N4022, N1801);
not NOT1 (N4402, N4398);
nor NOR3 (N4403, N4399, N3726, N3142);
or OR2 (N4404, N4400, N1776);
or OR4 (N4405, N4402, N50, N2888, N1103);
nand NAND2 (N4406, N4404, N389);
xor XOR2 (N4407, N4395, N3230);
nor NOR2 (N4408, N4396, N3636);
xor XOR2 (N4409, N4372, N2683);
nor NOR2 (N4410, N4388, N3687);
buf BUF1 (N4411, N4393);
nand NAND2 (N4412, N4401, N1089);
or OR3 (N4413, N4406, N2436, N879);
xor XOR2 (N4414, N4407, N2745);
xor XOR2 (N4415, N4412, N3808);
buf BUF1 (N4416, N4415);
nor NOR4 (N4417, N4397, N108, N16, N731);
or OR4 (N4418, N4408, N1363, N2976, N897);
and AND4 (N4419, N4418, N3781, N3222, N1275);
nor NOR2 (N4420, N4405, N3946);
or OR2 (N4421, N4410, N3893);
nand NAND4 (N4422, N4403, N1435, N1141, N2907);
or OR4 (N4423, N4411, N395, N640, N1479);
nor NOR3 (N4424, N4416, N2816, N155);
xor XOR2 (N4425, N4422, N29);
nand NAND4 (N4426, N4419, N3842, N362, N2407);
buf BUF1 (N4427, N4423);
or OR2 (N4428, N4427, N4120);
or OR4 (N4429, N4420, N2689, N3361, N4416);
not NOT1 (N4430, N4417);
not NOT1 (N4431, N4428);
buf BUF1 (N4432, N4426);
nand NAND2 (N4433, N4413, N3218);
nand NAND3 (N4434, N4421, N2403, N2527);
not NOT1 (N4435, N4425);
not NOT1 (N4436, N4424);
or OR3 (N4437, N4436, N1958, N1853);
and AND4 (N4438, N4430, N139, N2179, N3921);
buf BUF1 (N4439, N4437);
buf BUF1 (N4440, N4439);
or OR2 (N4441, N4429, N2042);
or OR3 (N4442, N4414, N3319, N2378);
and AND2 (N4443, N4442, N4175);
xor XOR2 (N4444, N4433, N2742);
xor XOR2 (N4445, N4438, N440);
buf BUF1 (N4446, N4434);
and AND2 (N4447, N4435, N3341);
not NOT1 (N4448, N4444);
buf BUF1 (N4449, N4445);
nor NOR4 (N4450, N4440, N2303, N4310, N1762);
and AND2 (N4451, N4448, N2526);
not NOT1 (N4452, N4450);
or OR3 (N4453, N4432, N2283, N2761);
nand NAND4 (N4454, N4443, N934, N4099, N1087);
xor XOR2 (N4455, N4451, N3960);
not NOT1 (N4456, N4454);
or OR4 (N4457, N4409, N2657, N1977, N3512);
not NOT1 (N4458, N4441);
nor NOR2 (N4459, N4447, N4352);
xor XOR2 (N4460, N4431, N1436);
xor XOR2 (N4461, N4457, N1439);
xor XOR2 (N4462, N4461, N1894);
nor NOR2 (N4463, N4462, N2304);
nand NAND3 (N4464, N4452, N3553, N4127);
not NOT1 (N4465, N4455);
nor NOR2 (N4466, N4463, N1695);
not NOT1 (N4467, N4449);
nand NAND4 (N4468, N4446, N1398, N1612, N4092);
nand NAND2 (N4469, N4456, N3781);
not NOT1 (N4470, N4453);
nand NAND2 (N4471, N4469, N4269);
or OR2 (N4472, N4471, N2449);
or OR4 (N4473, N4467, N597, N501, N579);
or OR4 (N4474, N4464, N247, N2152, N4137);
nand NAND2 (N4475, N4473, N2922);
or OR4 (N4476, N4470, N4311, N2846, N3521);
nor NOR3 (N4477, N4474, N325, N793);
or OR4 (N4478, N4458, N3648, N3428, N2525);
not NOT1 (N4479, N4477);
nand NAND4 (N4480, N4460, N3127, N582, N2205);
or OR2 (N4481, N4472, N1829);
buf BUF1 (N4482, N4459);
nor NOR3 (N4483, N4481, N2812, N3771);
nor NOR4 (N4484, N4480, N2895, N4358, N1187);
or OR3 (N4485, N4484, N2936, N1681);
and AND4 (N4486, N4466, N4208, N3347, N4299);
nor NOR2 (N4487, N4478, N2840);
or OR2 (N4488, N4487, N4450);
nand NAND3 (N4489, N4465, N1373, N3856);
not NOT1 (N4490, N4479);
nor NOR3 (N4491, N4475, N3998, N1962);
not NOT1 (N4492, N4488);
xor XOR2 (N4493, N4491, N136);
not NOT1 (N4494, N4486);
nand NAND4 (N4495, N4482, N4121, N3142, N468);
and AND2 (N4496, N4468, N1219);
nor NOR3 (N4497, N4489, N1357, N1167);
not NOT1 (N4498, N4476);
xor XOR2 (N4499, N4490, N997);
or OR2 (N4500, N4498, N1986);
nand NAND4 (N4501, N4494, N1538, N738, N4165);
buf BUF1 (N4502, N4497);
nand NAND4 (N4503, N4501, N1790, N1330, N4240);
not NOT1 (N4504, N4499);
or OR2 (N4505, N4496, N389);
or OR2 (N4506, N4502, N3764);
nand NAND3 (N4507, N4503, N2571, N1315);
nand NAND3 (N4508, N4493, N4214, N2083);
and AND3 (N4509, N4500, N4455, N2725);
nor NOR4 (N4510, N4509, N3146, N180, N603);
nand NAND4 (N4511, N4506, N3329, N1922, N1817);
and AND3 (N4512, N4504, N1672, N172);
or OR2 (N4513, N4511, N1712);
buf BUF1 (N4514, N4495);
or OR3 (N4515, N4483, N4449, N3143);
not NOT1 (N4516, N4507);
nor NOR4 (N4517, N4513, N43, N2056, N1252);
buf BUF1 (N4518, N4516);
or OR4 (N4519, N4514, N4412, N4060, N3289);
nand NAND2 (N4520, N4485, N2389);
xor XOR2 (N4521, N4515, N1574);
buf BUF1 (N4522, N4521);
and AND4 (N4523, N4508, N362, N1531, N1568);
xor XOR2 (N4524, N4520, N1390);
nand NAND2 (N4525, N4522, N3502);
or OR2 (N4526, N4505, N941);
or OR2 (N4527, N4519, N245);
nor NOR2 (N4528, N4523, N1469);
buf BUF1 (N4529, N4517);
buf BUF1 (N4530, N4529);
nand NAND3 (N4531, N4524, N3344, N3567);
and AND3 (N4532, N4526, N1184, N743);
buf BUF1 (N4533, N4512);
buf BUF1 (N4534, N4518);
not NOT1 (N4535, N4530);
buf BUF1 (N4536, N4525);
and AND2 (N4537, N4492, N1897);
and AND2 (N4538, N4510, N1669);
not NOT1 (N4539, N4535);
or OR4 (N4540, N4534, N479, N3355, N1652);
or OR2 (N4541, N4533, N3828);
or OR2 (N4542, N4531, N2941);
and AND4 (N4543, N4528, N3592, N4301, N2313);
nor NOR4 (N4544, N4532, N3567, N1159, N269);
not NOT1 (N4545, N4527);
nand NAND3 (N4546, N4537, N2346, N1321);
or OR2 (N4547, N4545, N2058);
not NOT1 (N4548, N4540);
buf BUF1 (N4549, N4542);
buf BUF1 (N4550, N4538);
nor NOR2 (N4551, N4536, N2660);
or OR2 (N4552, N4548, N2493);
and AND3 (N4553, N4541, N1497, N2924);
or OR2 (N4554, N4543, N3574);
and AND4 (N4555, N4552, N1516, N1671, N2036);
or OR2 (N4556, N4549, N2319);
or OR3 (N4557, N4554, N2858, N3676);
nand NAND3 (N4558, N4553, N874, N1264);
xor XOR2 (N4559, N4557, N3679);
buf BUF1 (N4560, N4558);
not NOT1 (N4561, N4550);
nand NAND4 (N4562, N4546, N1935, N1135, N2306);
or OR2 (N4563, N4547, N2443);
and AND2 (N4564, N4562, N4522);
and AND3 (N4565, N4561, N3486, N4144);
xor XOR2 (N4566, N4551, N1683);
not NOT1 (N4567, N4539);
buf BUF1 (N4568, N4559);
buf BUF1 (N4569, N4556);
nor NOR2 (N4570, N4555, N3746);
nor NOR2 (N4571, N4564, N2936);
and AND4 (N4572, N4568, N2441, N905, N1172);
and AND3 (N4573, N4560, N3365, N4553);
nor NOR4 (N4574, N4566, N3924, N260, N3519);
buf BUF1 (N4575, N4573);
or OR3 (N4576, N4569, N57, N799);
buf BUF1 (N4577, N4574);
nand NAND2 (N4578, N4563, N1561);
xor XOR2 (N4579, N4565, N1144);
nor NOR3 (N4580, N4572, N3115, N2056);
buf BUF1 (N4581, N4577);
not NOT1 (N4582, N4571);
not NOT1 (N4583, N4576);
and AND3 (N4584, N4583, N689, N113);
nand NAND3 (N4585, N4578, N4502, N4530);
not NOT1 (N4586, N4567);
and AND4 (N4587, N4581, N1741, N1038, N1215);
or OR3 (N4588, N4585, N4490, N570);
buf BUF1 (N4589, N4586);
not NOT1 (N4590, N4587);
and AND2 (N4591, N4579, N3454);
buf BUF1 (N4592, N4582);
and AND2 (N4593, N4575, N1428);
buf BUF1 (N4594, N4544);
not NOT1 (N4595, N4593);
not NOT1 (N4596, N4591);
nor NOR4 (N4597, N4570, N557, N4233, N3604);
buf BUF1 (N4598, N4580);
not NOT1 (N4599, N4589);
xor XOR2 (N4600, N4584, N171);
nor NOR4 (N4601, N4599, N1320, N3197, N2034);
and AND4 (N4602, N4597, N594, N3110, N3327);
and AND2 (N4603, N4598, N1332);
nand NAND2 (N4604, N4592, N1472);
buf BUF1 (N4605, N4600);
not NOT1 (N4606, N4588);
nand NAND3 (N4607, N4605, N2453, N3004);
buf BUF1 (N4608, N4596);
nand NAND3 (N4609, N4607, N1523, N3884);
nand NAND4 (N4610, N4609, N1305, N4575, N2162);
not NOT1 (N4611, N4608);
not NOT1 (N4612, N4610);
xor XOR2 (N4613, N4590, N1971);
nor NOR2 (N4614, N4611, N1788);
nor NOR3 (N4615, N4604, N4303, N2564);
xor XOR2 (N4616, N4615, N1821);
not NOT1 (N4617, N4603);
not NOT1 (N4618, N4613);
or OR4 (N4619, N4602, N1544, N3448, N2322);
buf BUF1 (N4620, N4594);
xor XOR2 (N4621, N4618, N2859);
xor XOR2 (N4622, N4619, N1761);
not NOT1 (N4623, N4612);
and AND2 (N4624, N4616, N1943);
nor NOR2 (N4625, N4622, N2249);
not NOT1 (N4626, N4625);
xor XOR2 (N4627, N4595, N711);
nand NAND3 (N4628, N4617, N3057, N2230);
and AND2 (N4629, N4614, N2029);
and AND2 (N4630, N4628, N633);
buf BUF1 (N4631, N4630);
and AND3 (N4632, N4629, N3579, N3644);
or OR4 (N4633, N4627, N3666, N2336, N1497);
or OR3 (N4634, N4601, N4565, N2679);
not NOT1 (N4635, N4633);
nor NOR2 (N4636, N4634, N590);
and AND2 (N4637, N4636, N2076);
nand NAND4 (N4638, N4631, N1648, N2362, N628);
nand NAND2 (N4639, N4626, N2252);
xor XOR2 (N4640, N4632, N1023);
not NOT1 (N4641, N4637);
xor XOR2 (N4642, N4623, N2713);
and AND4 (N4643, N4635, N3725, N3388, N241);
nor NOR3 (N4644, N4638, N730, N967);
nor NOR2 (N4645, N4624, N3763);
not NOT1 (N4646, N4620);
or OR2 (N4647, N4621, N3022);
or OR3 (N4648, N4646, N2529, N3345);
nand NAND3 (N4649, N4640, N3216, N20);
or OR4 (N4650, N4606, N3463, N2245, N3058);
buf BUF1 (N4651, N4645);
buf BUF1 (N4652, N4644);
nor NOR2 (N4653, N4652, N15);
xor XOR2 (N4654, N4643, N4330);
not NOT1 (N4655, N4654);
buf BUF1 (N4656, N4648);
xor XOR2 (N4657, N4642, N1770);
buf BUF1 (N4658, N4651);
not NOT1 (N4659, N4656);
or OR3 (N4660, N4647, N2658, N1292);
not NOT1 (N4661, N4649);
nor NOR3 (N4662, N4655, N1218, N28);
nand NAND4 (N4663, N4662, N1901, N2665, N4039);
nand NAND2 (N4664, N4650, N4040);
nand NAND3 (N4665, N4663, N1901, N4454);
not NOT1 (N4666, N4661);
xor XOR2 (N4667, N4641, N2);
xor XOR2 (N4668, N4665, N4599);
or OR4 (N4669, N4658, N4181, N3168, N3383);
nor NOR4 (N4670, N4664, N4199, N3303, N3715);
and AND3 (N4671, N4653, N3179, N1574);
and AND3 (N4672, N4659, N4051, N4434);
and AND3 (N4673, N4671, N1645, N4567);
buf BUF1 (N4674, N4639);
buf BUF1 (N4675, N4674);
xor XOR2 (N4676, N4669, N4001);
nand NAND4 (N4677, N4676, N4448, N1955, N3448);
nor NOR3 (N4678, N4657, N367, N1430);
buf BUF1 (N4679, N4666);
buf BUF1 (N4680, N4660);
xor XOR2 (N4681, N4675, N3136);
not NOT1 (N4682, N4673);
and AND4 (N4683, N4667, N3334, N2391, N391);
nor NOR4 (N4684, N4677, N2223, N194, N880);
nand NAND3 (N4685, N4683, N2897, N845);
nor NOR2 (N4686, N4670, N2784);
or OR4 (N4687, N4668, N3935, N2568, N2087);
not NOT1 (N4688, N4687);
and AND3 (N4689, N4682, N2452, N300);
or OR2 (N4690, N4688, N1426);
or OR2 (N4691, N4685, N4666);
nor NOR3 (N4692, N4686, N3116, N4279);
and AND4 (N4693, N4684, N3037, N4107, N1503);
nor NOR3 (N4694, N4680, N1560, N4684);
buf BUF1 (N4695, N4678);
buf BUF1 (N4696, N4679);
buf BUF1 (N4697, N4693);
nor NOR4 (N4698, N4695, N1565, N4179, N4632);
and AND3 (N4699, N4691, N1719, N3958);
or OR2 (N4700, N4697, N4680);
or OR3 (N4701, N4672, N2603, N894);
xor XOR2 (N4702, N4700, N1603);
and AND2 (N4703, N4689, N1497);
xor XOR2 (N4704, N4702, N2303);
or OR4 (N4705, N4696, N3365, N1542, N3124);
buf BUF1 (N4706, N4690);
and AND3 (N4707, N4706, N3050, N3163);
or OR4 (N4708, N4698, N359, N623, N4421);
not NOT1 (N4709, N4708);
xor XOR2 (N4710, N4701, N4197);
or OR4 (N4711, N4709, N4290, N504, N1925);
not NOT1 (N4712, N4681);
or OR2 (N4713, N4694, N2266);
xor XOR2 (N4714, N4710, N701);
or OR2 (N4715, N4707, N2911);
buf BUF1 (N4716, N4715);
nor NOR4 (N4717, N4703, N2622, N708, N3111);
not NOT1 (N4718, N4699);
nor NOR4 (N4719, N4716, N1549, N498, N2678);
and AND4 (N4720, N4714, N2628, N1321, N3861);
nand NAND4 (N4721, N4692, N2936, N3330, N2166);
and AND2 (N4722, N4705, N4639);
nor NOR2 (N4723, N4717, N1363);
or OR3 (N4724, N4723, N2017, N3018);
and AND2 (N4725, N4713, N4544);
or OR2 (N4726, N4712, N4086);
not NOT1 (N4727, N4725);
nand NAND4 (N4728, N4704, N2716, N3939, N588);
xor XOR2 (N4729, N4721, N1328);
not NOT1 (N4730, N4718);
not NOT1 (N4731, N4727);
xor XOR2 (N4732, N4730, N3596);
or OR2 (N4733, N4728, N3962);
and AND3 (N4734, N4724, N4630, N332);
buf BUF1 (N4735, N4734);
nand NAND3 (N4736, N4735, N3656, N2600);
nor NOR3 (N4737, N4736, N403, N597);
xor XOR2 (N4738, N4711, N3132);
buf BUF1 (N4739, N4732);
xor XOR2 (N4740, N4726, N86);
nand NAND3 (N4741, N4739, N3538, N2148);
buf BUF1 (N4742, N4740);
not NOT1 (N4743, N4719);
nand NAND3 (N4744, N4742, N2053, N2328);
buf BUF1 (N4745, N4737);
not NOT1 (N4746, N4731);
xor XOR2 (N4747, N4744, N35);
nand NAND2 (N4748, N4720, N3828);
xor XOR2 (N4749, N4722, N2630);
nor NOR3 (N4750, N4745, N2029, N1750);
and AND3 (N4751, N4748, N3277, N2845);
nand NAND2 (N4752, N4743, N4571);
buf BUF1 (N4753, N4750);
not NOT1 (N4754, N4738);
and AND2 (N4755, N4754, N2563);
not NOT1 (N4756, N4755);
nor NOR3 (N4757, N4749, N3942, N904);
and AND3 (N4758, N4757, N916, N787);
nand NAND3 (N4759, N4747, N1102, N176);
nor NOR2 (N4760, N4733, N1355);
buf BUF1 (N4761, N4753);
nand NAND4 (N4762, N4741, N4514, N507, N2256);
nand NAND3 (N4763, N4751, N1568, N4214);
nand NAND2 (N4764, N4762, N3002);
xor XOR2 (N4765, N4752, N509);
and AND3 (N4766, N4765, N2315, N4736);
nand NAND2 (N4767, N4729, N2602);
buf BUF1 (N4768, N4767);
not NOT1 (N4769, N4768);
nor NOR4 (N4770, N4756, N3040, N455, N2284);
not NOT1 (N4771, N4769);
nor NOR4 (N4772, N4771, N4122, N4549, N722);
buf BUF1 (N4773, N4764);
buf BUF1 (N4774, N4759);
or OR4 (N4775, N4763, N334, N3698, N1790);
nand NAND2 (N4776, N4760, N1861);
nor NOR4 (N4777, N4772, N1823, N2813, N1186);
nor NOR4 (N4778, N4774, N295, N3876, N3489);
or OR4 (N4779, N4761, N3403, N1399, N1488);
or OR2 (N4780, N4758, N1106);
nand NAND2 (N4781, N4777, N3314);
buf BUF1 (N4782, N4778);
or OR3 (N4783, N4773, N4626, N3744);
and AND2 (N4784, N4781, N4734);
xor XOR2 (N4785, N4775, N3264);
nor NOR3 (N4786, N4785, N1003, N2262);
buf BUF1 (N4787, N4776);
xor XOR2 (N4788, N4746, N3742);
nor NOR2 (N4789, N4788, N2174);
and AND4 (N4790, N4770, N574, N82, N4104);
nand NAND4 (N4791, N4783, N3900, N1106, N4366);
buf BUF1 (N4792, N4789);
not NOT1 (N4793, N4784);
nand NAND2 (N4794, N4792, N796);
nand NAND3 (N4795, N4782, N1853, N1079);
xor XOR2 (N4796, N4793, N1390);
buf BUF1 (N4797, N4794);
buf BUF1 (N4798, N4786);
and AND2 (N4799, N4791, N2653);
or OR4 (N4800, N4787, N876, N3247, N1026);
not NOT1 (N4801, N4790);
xor XOR2 (N4802, N4798, N3543);
buf BUF1 (N4803, N4802);
nand NAND3 (N4804, N4801, N3767, N510);
nor NOR3 (N4805, N4796, N1585, N2118);
buf BUF1 (N4806, N4779);
nor NOR3 (N4807, N4800, N2971, N2543);
nor NOR3 (N4808, N4780, N36, N240);
nand NAND4 (N4809, N4795, N1037, N210, N4786);
buf BUF1 (N4810, N4809);
not NOT1 (N4811, N4807);
xor XOR2 (N4812, N4806, N1954);
nand NAND2 (N4813, N4766, N1769);
buf BUF1 (N4814, N4808);
xor XOR2 (N4815, N4803, N351);
not NOT1 (N4816, N4811);
xor XOR2 (N4817, N4813, N2312);
xor XOR2 (N4818, N4797, N4628);
buf BUF1 (N4819, N4804);
and AND2 (N4820, N4819, N1533);
xor XOR2 (N4821, N4805, N308);
xor XOR2 (N4822, N4814, N1233);
or OR3 (N4823, N4815, N4210, N2960);
or OR3 (N4824, N4823, N3729, N770);
not NOT1 (N4825, N4817);
and AND2 (N4826, N4799, N1155);
xor XOR2 (N4827, N4816, N1057);
nor NOR4 (N4828, N4824, N1382, N1532, N2359);
not NOT1 (N4829, N4825);
buf BUF1 (N4830, N4829);
xor XOR2 (N4831, N4826, N1101);
not NOT1 (N4832, N4821);
buf BUF1 (N4833, N4822);
buf BUF1 (N4834, N4833);
nand NAND4 (N4835, N4818, N2034, N1709, N2354);
nand NAND3 (N4836, N4831, N4648, N3763);
not NOT1 (N4837, N4834);
and AND4 (N4838, N4832, N2301, N3971, N2907);
nor NOR4 (N4839, N4820, N3447, N4481, N442);
buf BUF1 (N4840, N4839);
and AND2 (N4841, N4827, N1115);
not NOT1 (N4842, N4838);
xor XOR2 (N4843, N4840, N1079);
xor XOR2 (N4844, N4836, N1978);
or OR3 (N4845, N4842, N1633, N636);
not NOT1 (N4846, N4843);
buf BUF1 (N4847, N4830);
not NOT1 (N4848, N4828);
nand NAND4 (N4849, N4810, N3405, N4574, N2579);
or OR4 (N4850, N4835, N4700, N1609, N554);
not NOT1 (N4851, N4848);
not NOT1 (N4852, N4841);
not NOT1 (N4853, N4849);
buf BUF1 (N4854, N4844);
xor XOR2 (N4855, N4854, N2525);
not NOT1 (N4856, N4837);
and AND3 (N4857, N4853, N2365, N3728);
nand NAND3 (N4858, N4852, N2597, N2201);
or OR4 (N4859, N4858, N1557, N3122, N2141);
buf BUF1 (N4860, N4845);
nand NAND2 (N4861, N4859, N1949);
buf BUF1 (N4862, N4855);
buf BUF1 (N4863, N4850);
nand NAND4 (N4864, N4863, N1016, N4127, N43);
nor NOR4 (N4865, N4857, N1333, N2100, N1196);
nand NAND3 (N4866, N4861, N2979, N3502);
xor XOR2 (N4867, N4864, N422);
and AND3 (N4868, N4812, N1437, N278);
buf BUF1 (N4869, N4866);
nor NOR2 (N4870, N4846, N476);
buf BUF1 (N4871, N4860);
nand NAND4 (N4872, N4847, N4794, N1913, N423);
xor XOR2 (N4873, N4867, N3904);
and AND2 (N4874, N4856, N4546);
or OR4 (N4875, N4865, N2337, N178, N1458);
nor NOR4 (N4876, N4868, N1709, N3041, N1860);
or OR2 (N4877, N4874, N2296);
nor NOR3 (N4878, N4869, N3593, N3583);
buf BUF1 (N4879, N4875);
nor NOR2 (N4880, N4878, N3673);
xor XOR2 (N4881, N4877, N747);
buf BUF1 (N4882, N4876);
xor XOR2 (N4883, N4880, N1744);
not NOT1 (N4884, N4862);
not NOT1 (N4885, N4851);
or OR2 (N4886, N4873, N1024);
and AND4 (N4887, N4883, N1734, N603, N85);
buf BUF1 (N4888, N4882);
xor XOR2 (N4889, N4879, N3718);
nand NAND3 (N4890, N4872, N1064, N3948);
xor XOR2 (N4891, N4884, N1710);
nor NOR2 (N4892, N4871, N1566);
nor NOR3 (N4893, N4886, N3674, N250);
nor NOR4 (N4894, N4888, N4178, N2929, N1061);
buf BUF1 (N4895, N4894);
nand NAND3 (N4896, N4885, N2764, N3217);
nand NAND3 (N4897, N4893, N336, N3139);
buf BUF1 (N4898, N4887);
and AND2 (N4899, N4881, N4511);
nand NAND2 (N4900, N4892, N3264);
and AND3 (N4901, N4898, N4073, N4205);
nand NAND2 (N4902, N4897, N1388);
xor XOR2 (N4903, N4889, N4782);
buf BUF1 (N4904, N4902);
nor NOR4 (N4905, N4903, N4808, N663, N4417);
nor NOR4 (N4906, N4899, N2151, N713, N4684);
xor XOR2 (N4907, N4896, N3793);
nor NOR3 (N4908, N4890, N3254, N519);
not NOT1 (N4909, N4905);
nor NOR3 (N4910, N4909, N2158, N986);
or OR4 (N4911, N4900, N562, N3009, N2873);
xor XOR2 (N4912, N4911, N4747);
buf BUF1 (N4913, N4908);
or OR4 (N4914, N4910, N580, N1940, N1812);
nor NOR3 (N4915, N4904, N937, N1015);
and AND2 (N4916, N4895, N3444);
nand NAND3 (N4917, N4912, N1395, N297);
xor XOR2 (N4918, N4913, N942);
not NOT1 (N4919, N4917);
nor NOR2 (N4920, N4919, N1735);
and AND2 (N4921, N4915, N4180);
not NOT1 (N4922, N4907);
nor NOR2 (N4923, N4891, N2370);
not NOT1 (N4924, N4923);
nor NOR4 (N4925, N4920, N4212, N253, N1211);
nand NAND2 (N4926, N4906, N828);
xor XOR2 (N4927, N4926, N3877);
xor XOR2 (N4928, N4918, N592);
or OR3 (N4929, N4924, N2463, N622);
nand NAND4 (N4930, N4928, N4358, N3199, N2143);
nand NAND3 (N4931, N4921, N381, N3965);
buf BUF1 (N4932, N4870);
buf BUF1 (N4933, N4914);
xor XOR2 (N4934, N4916, N4122);
not NOT1 (N4935, N4901);
nor NOR3 (N4936, N4930, N4780, N626);
or OR2 (N4937, N4925, N1471);
buf BUF1 (N4938, N4927);
not NOT1 (N4939, N4933);
or OR3 (N4940, N4934, N3407, N2938);
xor XOR2 (N4941, N4935, N3861);
and AND2 (N4942, N4939, N1088);
nor NOR3 (N4943, N4937, N4606, N92);
nand NAND4 (N4944, N4936, N2360, N2154, N1361);
nor NOR3 (N4945, N4944, N2984, N240);
nand NAND3 (N4946, N4931, N128, N2384);
nor NOR4 (N4947, N4942, N2840, N186, N4871);
not NOT1 (N4948, N4929);
or OR2 (N4949, N4922, N812);
not NOT1 (N4950, N4940);
and AND3 (N4951, N4943, N3239, N2565);
buf BUF1 (N4952, N4941);
and AND4 (N4953, N4948, N848, N2512, N450);
nor NOR2 (N4954, N4949, N2392);
and AND2 (N4955, N4953, N2008);
nor NOR2 (N4956, N4947, N2446);
not NOT1 (N4957, N4945);
and AND2 (N4958, N4955, N1746);
or OR4 (N4959, N4957, N4028, N711, N913);
buf BUF1 (N4960, N4946);
buf BUF1 (N4961, N4938);
or OR4 (N4962, N4961, N2621, N1876, N4290);
nand NAND4 (N4963, N4951, N825, N586, N1544);
or OR3 (N4964, N4932, N1285, N2802);
not NOT1 (N4965, N4958);
and AND4 (N4966, N4956, N1344, N3367, N3012);
xor XOR2 (N4967, N4952, N427);
nand NAND4 (N4968, N4959, N2993, N1551, N1633);
buf BUF1 (N4969, N4962);
nand NAND3 (N4970, N4965, N1332, N4952);
or OR3 (N4971, N4954, N3190, N795);
nor NOR2 (N4972, N4967, N2790);
not NOT1 (N4973, N4964);
nor NOR4 (N4974, N4971, N1870, N2822, N2114);
not NOT1 (N4975, N4974);
not NOT1 (N4976, N4966);
and AND4 (N4977, N4969, N666, N3435, N3025);
nor NOR2 (N4978, N4976, N4895);
and AND3 (N4979, N4970, N1880, N4923);
xor XOR2 (N4980, N4960, N1347);
not NOT1 (N4981, N4968);
xor XOR2 (N4982, N4977, N2128);
or OR2 (N4983, N4973, N4636);
or OR3 (N4984, N4950, N3935, N1929);
xor XOR2 (N4985, N4972, N2297);
not NOT1 (N4986, N4980);
and AND4 (N4987, N4985, N3685, N2392, N466);
nand NAND3 (N4988, N4987, N3664, N502);
and AND2 (N4989, N4981, N1068);
buf BUF1 (N4990, N4986);
nor NOR2 (N4991, N4978, N2081);
nor NOR2 (N4992, N4979, N83);
or OR3 (N4993, N4975, N123, N3507);
not NOT1 (N4994, N4963);
and AND2 (N4995, N4993, N146);
or OR3 (N4996, N4992, N1217, N1648);
not NOT1 (N4997, N4988);
or OR4 (N4998, N4982, N4149, N1888, N53);
xor XOR2 (N4999, N4995, N3922);
nor NOR4 (N5000, N4991, N1040, N4875, N2422);
not NOT1 (N5001, N4990);
nand NAND4 (N5002, N4983, N4855, N1438, N2171);
not NOT1 (N5003, N5001);
nand NAND2 (N5004, N4989, N1750);
nor NOR3 (N5005, N4996, N560, N877);
not NOT1 (N5006, N4998);
and AND2 (N5007, N4997, N4160);
xor XOR2 (N5008, N4999, N935);
or OR2 (N5009, N5002, N4129);
nand NAND4 (N5010, N4994, N3130, N2226, N2733);
or OR2 (N5011, N5007, N1586);
or OR3 (N5012, N4984, N4107, N3080);
or OR2 (N5013, N5000, N2376);
and AND2 (N5014, N5004, N2238);
nor NOR3 (N5015, N5003, N2464, N312);
nor NOR2 (N5016, N5005, N2205);
or OR2 (N5017, N5008, N1573);
xor XOR2 (N5018, N5011, N3481);
not NOT1 (N5019, N5017);
nand NAND4 (N5020, N5013, N5011, N1864, N3036);
nand NAND4 (N5021, N5016, N1386, N2558, N4410);
nor NOR3 (N5022, N5006, N3844, N304);
xor XOR2 (N5023, N5010, N4567);
not NOT1 (N5024, N5019);
nand NAND2 (N5025, N5018, N4034);
nand NAND2 (N5026, N5022, N4717);
and AND4 (N5027, N5015, N572, N3613, N3913);
xor XOR2 (N5028, N5026, N3950);
and AND4 (N5029, N5014, N1309, N1825, N2002);
or OR4 (N5030, N5025, N821, N1706, N1339);
xor XOR2 (N5031, N5023, N3626);
or OR4 (N5032, N5020, N65, N3287, N2333);
nand NAND2 (N5033, N5009, N3544);
nor NOR3 (N5034, N5031, N2222, N4261);
and AND4 (N5035, N5029, N1330, N3602, N251);
and AND2 (N5036, N5030, N3027);
nor NOR3 (N5037, N5033, N4300, N956);
nand NAND2 (N5038, N5012, N2553);
buf BUF1 (N5039, N5037);
not NOT1 (N5040, N5027);
and AND2 (N5041, N5024, N4483);
and AND4 (N5042, N5038, N186, N2631, N4289);
nand NAND2 (N5043, N5036, N2977);
and AND4 (N5044, N5039, N2084, N3651, N4286);
nand NAND4 (N5045, N5021, N3166, N4998, N2086);
nor NOR2 (N5046, N5032, N249);
not NOT1 (N5047, N5028);
nor NOR2 (N5048, N5044, N4746);
or OR2 (N5049, N5045, N381);
nand NAND2 (N5050, N5048, N5047);
nand NAND4 (N5051, N3843, N2978, N4157, N3384);
or OR4 (N5052, N5049, N3684, N4155, N2993);
not NOT1 (N5053, N5052);
nand NAND3 (N5054, N5040, N770, N2095);
and AND4 (N5055, N5054, N1632, N5031, N4718);
nor NOR3 (N5056, N5050, N1926, N2049);
xor XOR2 (N5057, N5042, N4587);
not NOT1 (N5058, N5046);
nand NAND2 (N5059, N5034, N2051);
buf BUF1 (N5060, N5053);
and AND2 (N5061, N5041, N700);
xor XOR2 (N5062, N5058, N2093);
buf BUF1 (N5063, N5055);
and AND3 (N5064, N5061, N798, N2542);
buf BUF1 (N5065, N5063);
buf BUF1 (N5066, N5060);
nor NOR3 (N5067, N5056, N3178, N3743);
xor XOR2 (N5068, N5066, N1212);
or OR4 (N5069, N5059, N3055, N4925, N481);
nor NOR4 (N5070, N5062, N4922, N3261, N4479);
not NOT1 (N5071, N5035);
nand NAND2 (N5072, N5071, N3029);
nand NAND3 (N5073, N5051, N1994, N4614);
xor XOR2 (N5074, N5043, N3165);
not NOT1 (N5075, N5069);
nand NAND3 (N5076, N5070, N4641, N2699);
and AND3 (N5077, N5065, N4035, N2486);
xor XOR2 (N5078, N5076, N1333);
buf BUF1 (N5079, N5077);
or OR3 (N5080, N5078, N3027, N1295);
and AND4 (N5081, N5073, N1046, N2701, N4233);
not NOT1 (N5082, N5079);
not NOT1 (N5083, N5081);
buf BUF1 (N5084, N5057);
or OR2 (N5085, N5075, N352);
and AND2 (N5086, N5085, N4676);
nor NOR4 (N5087, N5064, N1863, N2667, N2095);
and AND3 (N5088, N5080, N1797, N1184);
nor NOR2 (N5089, N5086, N1695);
nor NOR2 (N5090, N5088, N3825);
or OR2 (N5091, N5084, N3921);
and AND3 (N5092, N5091, N678, N2515);
nor NOR2 (N5093, N5067, N799);
buf BUF1 (N5094, N5093);
xor XOR2 (N5095, N5082, N1397);
nor NOR3 (N5096, N5089, N1206, N3798);
or OR2 (N5097, N5094, N4299);
buf BUF1 (N5098, N5072);
or OR3 (N5099, N5098, N703, N1294);
or OR2 (N5100, N5095, N781);
or OR3 (N5101, N5099, N1080, N2747);
buf BUF1 (N5102, N5096);
xor XOR2 (N5103, N5087, N3867);
and AND4 (N5104, N5101, N2054, N3666, N2443);
xor XOR2 (N5105, N5097, N4616);
or OR2 (N5106, N5083, N3612);
or OR2 (N5107, N5090, N1998);
not NOT1 (N5108, N5100);
not NOT1 (N5109, N5103);
and AND4 (N5110, N5107, N1623, N3508, N3);
buf BUF1 (N5111, N5074);
not NOT1 (N5112, N5110);
buf BUF1 (N5113, N5104);
not NOT1 (N5114, N5113);
xor XOR2 (N5115, N5102, N3604);
or OR2 (N5116, N5114, N3357);
nor NOR2 (N5117, N5112, N382);
xor XOR2 (N5118, N5109, N1348);
xor XOR2 (N5119, N5108, N3474);
and AND2 (N5120, N5119, N428);
or OR3 (N5121, N5116, N4599, N2475);
or OR4 (N5122, N5111, N4521, N4442, N971);
nor NOR4 (N5123, N5117, N3701, N4264, N5116);
nor NOR2 (N5124, N5120, N959);
buf BUF1 (N5125, N5092);
and AND4 (N5126, N5106, N2975, N3571, N75);
and AND2 (N5127, N5118, N766);
or OR2 (N5128, N5127, N829);
nor NOR4 (N5129, N5124, N1078, N310, N2928);
nand NAND2 (N5130, N5105, N3999);
and AND2 (N5131, N5068, N3886);
buf BUF1 (N5132, N5122);
xor XOR2 (N5133, N5128, N3697);
xor XOR2 (N5134, N5129, N3450);
nand NAND3 (N5135, N5121, N961, N3144);
and AND3 (N5136, N5135, N1951, N3182);
nor NOR2 (N5137, N5131, N616);
buf BUF1 (N5138, N5126);
or OR4 (N5139, N5123, N558, N3335, N3800);
nor NOR4 (N5140, N5134, N1808, N2297, N1871);
nor NOR3 (N5141, N5133, N1128, N4112);
and AND2 (N5142, N5115, N3511);
buf BUF1 (N5143, N5140);
or OR2 (N5144, N5137, N4876);
nand NAND4 (N5145, N5142, N4060, N2152, N3455);
nand NAND4 (N5146, N5132, N4312, N3122, N2957);
nor NOR3 (N5147, N5144, N314, N1121);
or OR4 (N5148, N5139, N700, N1665, N2835);
not NOT1 (N5149, N5147);
or OR3 (N5150, N5130, N5015, N3626);
xor XOR2 (N5151, N5141, N4000);
or OR4 (N5152, N5136, N817, N3094, N4581);
buf BUF1 (N5153, N5138);
or OR2 (N5154, N5143, N2837);
nand NAND2 (N5155, N5154, N1779);
and AND4 (N5156, N5153, N4130, N455, N507);
buf BUF1 (N5157, N5146);
buf BUF1 (N5158, N5145);
nand NAND4 (N5159, N5151, N2551, N239, N3852);
not NOT1 (N5160, N5157);
or OR2 (N5161, N5149, N2002);
and AND4 (N5162, N5158, N4589, N4559, N210);
nand NAND4 (N5163, N5152, N4901, N1173, N3133);
and AND2 (N5164, N5159, N212);
not NOT1 (N5165, N5155);
xor XOR2 (N5166, N5162, N3597);
or OR3 (N5167, N5156, N2267, N4225);
nor NOR3 (N5168, N5163, N3143, N591);
nor NOR2 (N5169, N5161, N4138);
xor XOR2 (N5170, N5168, N4013);
not NOT1 (N5171, N5150);
or OR4 (N5172, N5160, N4660, N5151, N4621);
nand NAND4 (N5173, N5125, N3395, N3421, N4240);
nand NAND3 (N5174, N5171, N4713, N2772);
xor XOR2 (N5175, N5164, N1480);
xor XOR2 (N5176, N5165, N3985);
or OR3 (N5177, N5166, N1563, N5108);
nand NAND4 (N5178, N5175, N5095, N3485, N369);
buf BUF1 (N5179, N5169);
nor NOR4 (N5180, N5178, N1836, N3970, N1995);
and AND4 (N5181, N5148, N248, N4573, N4333);
xor XOR2 (N5182, N5180, N1530);
and AND2 (N5183, N5170, N1435);
nand NAND4 (N5184, N5183, N1728, N3134, N670);
and AND2 (N5185, N5177, N778);
buf BUF1 (N5186, N5167);
and AND3 (N5187, N5176, N4106, N3037);
nand NAND3 (N5188, N5185, N4508, N4572);
buf BUF1 (N5189, N5186);
not NOT1 (N5190, N5189);
xor XOR2 (N5191, N5181, N848);
and AND4 (N5192, N5179, N4705, N4697, N4105);
and AND2 (N5193, N5187, N4226);
xor XOR2 (N5194, N5192, N5132);
xor XOR2 (N5195, N5182, N3245);
and AND4 (N5196, N5194, N2674, N1106, N1773);
xor XOR2 (N5197, N5184, N3265);
or OR3 (N5198, N5174, N1799, N2278);
nor NOR2 (N5199, N5193, N4106);
xor XOR2 (N5200, N5196, N4905);
xor XOR2 (N5201, N5173, N3327);
xor XOR2 (N5202, N5200, N2956);
or OR2 (N5203, N5197, N4307);
xor XOR2 (N5204, N5202, N4870);
or OR4 (N5205, N5199, N1465, N1105, N5034);
buf BUF1 (N5206, N5201);
xor XOR2 (N5207, N5188, N884);
or OR4 (N5208, N5172, N2567, N2083, N3750);
nand NAND4 (N5209, N5191, N964, N2562, N3607);
or OR4 (N5210, N5208, N1871, N4548, N1062);
buf BUF1 (N5211, N5198);
nand NAND4 (N5212, N5195, N3793, N3827, N3855);
and AND4 (N5213, N5207, N2117, N2235, N487);
or OR4 (N5214, N5209, N4527, N4533, N1159);
or OR2 (N5215, N5212, N2580);
xor XOR2 (N5216, N5210, N2285);
and AND4 (N5217, N5190, N194, N3365, N2890);
nand NAND3 (N5218, N5205, N2693, N2604);
nand NAND4 (N5219, N5214, N4649, N1500, N4122);
and AND4 (N5220, N5204, N32, N3563, N3531);
buf BUF1 (N5221, N5218);
nand NAND3 (N5222, N5221, N3062, N2932);
and AND2 (N5223, N5213, N2607);
xor XOR2 (N5224, N5222, N4673);
xor XOR2 (N5225, N5216, N4134);
and AND2 (N5226, N5206, N2874);
or OR4 (N5227, N5223, N2557, N684, N4758);
nand NAND3 (N5228, N5219, N4326, N2686);
buf BUF1 (N5229, N5203);
buf BUF1 (N5230, N5220);
or OR4 (N5231, N5211, N2856, N2849, N54);
nand NAND2 (N5232, N5231, N4053);
nand NAND2 (N5233, N5217, N25);
buf BUF1 (N5234, N5224);
not NOT1 (N5235, N5227);
buf BUF1 (N5236, N5229);
or OR3 (N5237, N5228, N1212, N2194);
or OR3 (N5238, N5236, N4095, N4965);
nor NOR3 (N5239, N5238, N4004, N3770);
nand NAND3 (N5240, N5232, N2487, N2754);
nor NOR4 (N5241, N5215, N1985, N3317, N1792);
buf BUF1 (N5242, N5240);
xor XOR2 (N5243, N5225, N4195);
buf BUF1 (N5244, N5241);
and AND3 (N5245, N5244, N165, N3670);
nand NAND3 (N5246, N5237, N3864, N1622);
xor XOR2 (N5247, N5239, N2945);
or OR2 (N5248, N5234, N2136);
and AND3 (N5249, N5226, N1293, N4008);
or OR2 (N5250, N5248, N4072);
nor NOR2 (N5251, N5247, N3218);
buf BUF1 (N5252, N5230);
or OR3 (N5253, N5246, N2843, N3213);
and AND3 (N5254, N5245, N3621, N5231);
buf BUF1 (N5255, N5250);
and AND2 (N5256, N5249, N4567);
buf BUF1 (N5257, N5256);
or OR4 (N5258, N5255, N4101, N1586, N3774);
nand NAND3 (N5259, N5242, N5156, N1741);
xor XOR2 (N5260, N5235, N1285);
or OR4 (N5261, N5251, N5161, N3122, N279);
or OR2 (N5262, N5257, N4021);
buf BUF1 (N5263, N5252);
nor NOR2 (N5264, N5263, N4899);
or OR3 (N5265, N5253, N3746, N4433);
or OR2 (N5266, N5262, N3000);
or OR4 (N5267, N5258, N305, N545, N2683);
and AND3 (N5268, N5254, N4724, N4242);
nor NOR4 (N5269, N5261, N1085, N1050, N1718);
buf BUF1 (N5270, N5268);
xor XOR2 (N5271, N5233, N115);
nand NAND2 (N5272, N5265, N2869);
or OR2 (N5273, N5259, N614);
buf BUF1 (N5274, N5271);
xor XOR2 (N5275, N5269, N2776);
nor NOR3 (N5276, N5264, N2957, N2576);
nand NAND3 (N5277, N5266, N2729, N1880);
nor NOR3 (N5278, N5260, N3664, N1549);
nor NOR2 (N5279, N5276, N1742);
and AND4 (N5280, N5279, N2821, N2510, N4644);
and AND3 (N5281, N5273, N4765, N4206);
buf BUF1 (N5282, N5270);
nor NOR4 (N5283, N5243, N352, N2262, N3220);
nand NAND4 (N5284, N5267, N3032, N2169, N3774);
or OR3 (N5285, N5282, N74, N1188);
nor NOR3 (N5286, N5278, N193, N3394);
or OR3 (N5287, N5281, N2289, N2139);
buf BUF1 (N5288, N5285);
or OR2 (N5289, N5287, N4503);
nor NOR4 (N5290, N5280, N5182, N1897, N1553);
nor NOR4 (N5291, N5284, N5182, N4475, N1198);
buf BUF1 (N5292, N5289);
not NOT1 (N5293, N5286);
nor NOR3 (N5294, N5291, N3702, N5263);
xor XOR2 (N5295, N5275, N4069);
xor XOR2 (N5296, N5274, N1202);
nor NOR2 (N5297, N5290, N991);
xor XOR2 (N5298, N5297, N356);
and AND2 (N5299, N5296, N3962);
nand NAND3 (N5300, N5294, N2210, N2996);
nand NAND4 (N5301, N5300, N2405, N1442, N3447);
not NOT1 (N5302, N5298);
xor XOR2 (N5303, N5293, N1470);
not NOT1 (N5304, N5292);
nor NOR3 (N5305, N5301, N2464, N4852);
or OR4 (N5306, N5303, N4218, N3771, N193);
nand NAND2 (N5307, N5299, N611);
nand NAND4 (N5308, N5295, N4076, N3304, N93);
not NOT1 (N5309, N5277);
nor NOR2 (N5310, N5304, N4369);
nand NAND3 (N5311, N5306, N75, N1359);
nor NOR3 (N5312, N5305, N1228, N3005);
and AND2 (N5313, N5272, N3887);
nor NOR3 (N5314, N5288, N3049, N4178);
or OR4 (N5315, N5308, N337, N2215, N3826);
nand NAND4 (N5316, N5307, N4027, N3969, N3934);
xor XOR2 (N5317, N5309, N4036);
nand NAND2 (N5318, N5313, N595);
nor NOR2 (N5319, N5315, N717);
not NOT1 (N5320, N5319);
buf BUF1 (N5321, N5317);
nand NAND4 (N5322, N5311, N2207, N4079, N3104);
or OR2 (N5323, N5312, N3118);
buf BUF1 (N5324, N5283);
not NOT1 (N5325, N5302);
xor XOR2 (N5326, N5322, N1500);
not NOT1 (N5327, N5324);
nor NOR2 (N5328, N5310, N3401);
and AND4 (N5329, N5320, N1844, N3600, N2092);
xor XOR2 (N5330, N5325, N4555);
not NOT1 (N5331, N5329);
nand NAND2 (N5332, N5323, N2822);
not NOT1 (N5333, N5314);
nand NAND2 (N5334, N5318, N28);
or OR4 (N5335, N5328, N4832, N4790, N4240);
and AND2 (N5336, N5326, N4061);
and AND2 (N5337, N5321, N3590);
buf BUF1 (N5338, N5336);
nand NAND3 (N5339, N5327, N5008, N2347);
nand NAND4 (N5340, N5316, N4495, N4313, N21);
nand NAND4 (N5341, N5339, N2566, N4420, N3504);
nor NOR2 (N5342, N5333, N2391);
and AND4 (N5343, N5342, N3069, N3465, N1947);
not NOT1 (N5344, N5331);
not NOT1 (N5345, N5330);
not NOT1 (N5346, N5332);
nor NOR3 (N5347, N5345, N4140, N3558);
or OR3 (N5348, N5346, N868, N1699);
and AND2 (N5349, N5340, N5078);
or OR4 (N5350, N5347, N4837, N1785, N3892);
xor XOR2 (N5351, N5337, N2407);
not NOT1 (N5352, N5351);
xor XOR2 (N5353, N5352, N700);
buf BUF1 (N5354, N5338);
and AND4 (N5355, N5335, N4722, N2338, N3337);
nor NOR2 (N5356, N5353, N4609);
nor NOR3 (N5357, N5334, N750, N3303);
nor NOR3 (N5358, N5344, N1534, N1589);
nor NOR4 (N5359, N5343, N437, N320, N962);
buf BUF1 (N5360, N5355);
and AND3 (N5361, N5360, N4672, N18);
buf BUF1 (N5362, N5349);
or OR3 (N5363, N5356, N2687, N2286);
or OR3 (N5364, N5350, N981, N600);
and AND3 (N5365, N5354, N1704, N1340);
xor XOR2 (N5366, N5358, N2959);
nor NOR4 (N5367, N5366, N1153, N2459, N4187);
buf BUF1 (N5368, N5361);
or OR3 (N5369, N5367, N496, N5103);
nand NAND3 (N5370, N5368, N594, N124);
xor XOR2 (N5371, N5363, N404);
or OR2 (N5372, N5348, N4483);
not NOT1 (N5373, N5362);
and AND2 (N5374, N5365, N1927);
not NOT1 (N5375, N5373);
nand NAND2 (N5376, N5371, N1210);
or OR2 (N5377, N5364, N1521);
or OR2 (N5378, N5341, N3869);
nor NOR4 (N5379, N5359, N1191, N4738, N1968);
nor NOR3 (N5380, N5357, N1294, N3404);
or OR4 (N5381, N5376, N3982, N2041, N974);
buf BUF1 (N5382, N5378);
not NOT1 (N5383, N5381);
and AND4 (N5384, N5377, N5314, N3129, N979);
nand NAND4 (N5385, N5379, N3675, N4355, N2321);
nor NOR2 (N5386, N5372, N980);
nor NOR2 (N5387, N5383, N1365);
xor XOR2 (N5388, N5384, N3498);
not NOT1 (N5389, N5370);
and AND2 (N5390, N5375, N3637);
or OR4 (N5391, N5388, N1059, N2485, N4836);
xor XOR2 (N5392, N5389, N322);
not NOT1 (N5393, N5374);
nor NOR2 (N5394, N5382, N1689);
or OR2 (N5395, N5391, N1615);
and AND3 (N5396, N5395, N2157, N3627);
nand NAND3 (N5397, N5392, N3256, N3444);
not NOT1 (N5398, N5390);
buf BUF1 (N5399, N5396);
and AND4 (N5400, N5387, N809, N3651, N1693);
nand NAND4 (N5401, N5399, N319, N4736, N3140);
nand NAND2 (N5402, N5397, N556);
nand NAND4 (N5403, N5401, N3375, N4145, N4430);
or OR4 (N5404, N5393, N5191, N3423, N4451);
xor XOR2 (N5405, N5403, N2575);
or OR2 (N5406, N5405, N4298);
or OR4 (N5407, N5385, N198, N4026, N2146);
xor XOR2 (N5408, N5402, N4383);
xor XOR2 (N5409, N5408, N1283);
nand NAND4 (N5410, N5386, N620, N4991, N1193);
not NOT1 (N5411, N5409);
and AND2 (N5412, N5410, N2719);
buf BUF1 (N5413, N5412);
or OR3 (N5414, N5404, N4792, N4681);
and AND3 (N5415, N5380, N3071, N2942);
xor XOR2 (N5416, N5411, N3753);
buf BUF1 (N5417, N5394);
xor XOR2 (N5418, N5398, N859);
xor XOR2 (N5419, N5413, N2078);
xor XOR2 (N5420, N5400, N4782);
nor NOR2 (N5421, N5420, N897);
xor XOR2 (N5422, N5416, N2201);
or OR4 (N5423, N5419, N2047, N348, N3941);
and AND2 (N5424, N5415, N4519);
and AND3 (N5425, N5424, N5222, N2338);
not NOT1 (N5426, N5406);
and AND2 (N5427, N5369, N135);
not NOT1 (N5428, N5421);
buf BUF1 (N5429, N5422);
buf BUF1 (N5430, N5427);
nand NAND2 (N5431, N5429, N2338);
nand NAND4 (N5432, N5431, N964, N3699, N1710);
xor XOR2 (N5433, N5432, N4482);
nor NOR2 (N5434, N5426, N4349);
nor NOR3 (N5435, N5417, N3214, N37);
nand NAND2 (N5436, N5428, N763);
or OR4 (N5437, N5434, N3510, N408, N4855);
or OR3 (N5438, N5418, N3383, N2146);
buf BUF1 (N5439, N5438);
and AND2 (N5440, N5439, N4580);
nor NOR2 (N5441, N5407, N4722);
xor XOR2 (N5442, N5414, N943);
buf BUF1 (N5443, N5425);
buf BUF1 (N5444, N5442);
not NOT1 (N5445, N5441);
buf BUF1 (N5446, N5437);
nor NOR2 (N5447, N5446, N1701);
buf BUF1 (N5448, N5443);
nor NOR4 (N5449, N5445, N4541, N4968, N3333);
xor XOR2 (N5450, N5440, N3667);
xor XOR2 (N5451, N5447, N4073);
or OR3 (N5452, N5448, N424, N1587);
or OR3 (N5453, N5436, N506, N3046);
nand NAND2 (N5454, N5450, N2412);
or OR2 (N5455, N5453, N3860);
not NOT1 (N5456, N5444);
not NOT1 (N5457, N5433);
not NOT1 (N5458, N5454);
nor NOR3 (N5459, N5455, N2242, N3699);
nand NAND3 (N5460, N5430, N2344, N2843);
not NOT1 (N5461, N5423);
xor XOR2 (N5462, N5452, N5074);
xor XOR2 (N5463, N5461, N520);
buf BUF1 (N5464, N5451);
and AND4 (N5465, N5456, N3863, N2982, N433);
or OR4 (N5466, N5463, N83, N533, N3085);
nor NOR2 (N5467, N5457, N3064);
not NOT1 (N5468, N5464);
nor NOR2 (N5469, N5462, N5029);
xor XOR2 (N5470, N5468, N996);
and AND4 (N5471, N5435, N2702, N3863, N3472);
xor XOR2 (N5472, N5470, N4803);
nand NAND3 (N5473, N5466, N3469, N5463);
xor XOR2 (N5474, N5473, N777);
and AND2 (N5475, N5459, N2460);
and AND4 (N5476, N5467, N517, N2880, N3498);
or OR4 (N5477, N5469, N2794, N2815, N645);
nand NAND4 (N5478, N5476, N1494, N2176, N1754);
nor NOR4 (N5479, N5460, N1909, N2734, N4);
xor XOR2 (N5480, N5477, N2649);
nor NOR2 (N5481, N5475, N4078);
nand NAND3 (N5482, N5449, N3922, N3254);
or OR2 (N5483, N5465, N3259);
xor XOR2 (N5484, N5472, N4445);
nor NOR3 (N5485, N5479, N3436, N1033);
nor NOR2 (N5486, N5474, N3742);
xor XOR2 (N5487, N5458, N3040);
or OR4 (N5488, N5487, N4360, N1054, N4914);
nand NAND3 (N5489, N5486, N1223, N3574);
not NOT1 (N5490, N5471);
nand NAND3 (N5491, N5489, N1492, N4361);
or OR4 (N5492, N5488, N2771, N1555, N5217);
xor XOR2 (N5493, N5484, N1609);
or OR2 (N5494, N5480, N902);
nand NAND2 (N5495, N5490, N2735);
buf BUF1 (N5496, N5492);
and AND2 (N5497, N5491, N1680);
and AND3 (N5498, N5483, N4733, N5228);
xor XOR2 (N5499, N5478, N1238);
not NOT1 (N5500, N5482);
nand NAND4 (N5501, N5494, N207, N26, N4482);
xor XOR2 (N5502, N5485, N2366);
or OR4 (N5503, N5501, N938, N619, N4351);
or OR2 (N5504, N5502, N5269);
xor XOR2 (N5505, N5499, N131);
or OR2 (N5506, N5493, N4849);
and AND3 (N5507, N5495, N3149, N2241);
or OR3 (N5508, N5500, N777, N4987);
nand NAND2 (N5509, N5506, N2986);
nand NAND2 (N5510, N5503, N527);
and AND3 (N5511, N5504, N69, N4392);
xor XOR2 (N5512, N5508, N1308);
xor XOR2 (N5513, N5507, N3850);
and AND3 (N5514, N5498, N1507, N2724);
buf BUF1 (N5515, N5497);
not NOT1 (N5516, N5515);
nand NAND4 (N5517, N5496, N1244, N926, N3741);
nor NOR2 (N5518, N5509, N3556);
buf BUF1 (N5519, N5517);
nand NAND4 (N5520, N5505, N3575, N3254, N1258);
or OR3 (N5521, N5511, N5322, N1079);
not NOT1 (N5522, N5510);
xor XOR2 (N5523, N5481, N3241);
not NOT1 (N5524, N5516);
nand NAND2 (N5525, N5514, N2815);
xor XOR2 (N5526, N5523, N576);
nor NOR3 (N5527, N5524, N4397, N2807);
nor NOR2 (N5528, N5527, N2996);
and AND4 (N5529, N5512, N1939, N273, N5331);
xor XOR2 (N5530, N5522, N1272);
or OR4 (N5531, N5521, N2493, N281, N3223);
not NOT1 (N5532, N5513);
xor XOR2 (N5533, N5531, N5455);
buf BUF1 (N5534, N5518);
or OR2 (N5535, N5525, N4551);
xor XOR2 (N5536, N5532, N3042);
and AND3 (N5537, N5536, N3021, N1613);
xor XOR2 (N5538, N5526, N4180);
xor XOR2 (N5539, N5529, N407);
buf BUF1 (N5540, N5535);
nand NAND3 (N5541, N5528, N113, N3669);
and AND2 (N5542, N5539, N1311);
xor XOR2 (N5543, N5542, N1310);
nor NOR4 (N5544, N5537, N226, N2798, N1682);
xor XOR2 (N5545, N5541, N200);
and AND2 (N5546, N5533, N1334);
buf BUF1 (N5547, N5520);
nor NOR2 (N5548, N5519, N1367);
xor XOR2 (N5549, N5546, N3290);
or OR4 (N5550, N5543, N4919, N3197, N2351);
nand NAND2 (N5551, N5548, N2648);
not NOT1 (N5552, N5549);
or OR4 (N5553, N5550, N2332, N1115, N1407);
or OR2 (N5554, N5552, N2986);
nor NOR4 (N5555, N5551, N4241, N1836, N3647);
nor NOR2 (N5556, N5555, N5105);
xor XOR2 (N5557, N5545, N4361);
nand NAND2 (N5558, N5556, N1649);
not NOT1 (N5559, N5558);
nor NOR4 (N5560, N5553, N5107, N1933, N4702);
nand NAND3 (N5561, N5554, N1044, N4132);
buf BUF1 (N5562, N5561);
or OR2 (N5563, N5547, N1035);
nor NOR4 (N5564, N5560, N758, N2523, N4973);
nand NAND2 (N5565, N5563, N1190);
xor XOR2 (N5566, N5564, N116);
and AND3 (N5567, N5566, N744, N598);
nor NOR4 (N5568, N5540, N1424, N5021, N5532);
nor NOR4 (N5569, N5534, N172, N2113, N461);
not NOT1 (N5570, N5544);
nand NAND4 (N5571, N5557, N2048, N1082, N726);
not NOT1 (N5572, N5570);
and AND4 (N5573, N5569, N2351, N3317, N4373);
nor NOR2 (N5574, N5572, N1354);
nor NOR3 (N5575, N5562, N3326, N39);
xor XOR2 (N5576, N5530, N23);
nand NAND3 (N5577, N5559, N4103, N4997);
nor NOR3 (N5578, N5577, N2825, N4833);
and AND4 (N5579, N5578, N2887, N3329, N159);
xor XOR2 (N5580, N5579, N3282);
not NOT1 (N5581, N5565);
not NOT1 (N5582, N5576);
or OR2 (N5583, N5538, N5399);
and AND2 (N5584, N5573, N2524);
not NOT1 (N5585, N5583);
nor NOR2 (N5586, N5571, N3901);
and AND3 (N5587, N5581, N3300, N962);
buf BUF1 (N5588, N5586);
buf BUF1 (N5589, N5588);
and AND2 (N5590, N5574, N172);
not NOT1 (N5591, N5580);
xor XOR2 (N5592, N5582, N4473);
and AND2 (N5593, N5592, N4979);
or OR4 (N5594, N5589, N1267, N930, N4223);
and AND2 (N5595, N5594, N4529);
nand NAND2 (N5596, N5575, N285);
and AND3 (N5597, N5568, N4018, N1653);
xor XOR2 (N5598, N5590, N130);
and AND4 (N5599, N5585, N5076, N4758, N2028);
nor NOR2 (N5600, N5584, N2345);
xor XOR2 (N5601, N5595, N889);
buf BUF1 (N5602, N5596);
nor NOR4 (N5603, N5597, N5500, N1607, N5329);
and AND2 (N5604, N5567, N1036);
nor NOR2 (N5605, N5591, N2060);
or OR3 (N5606, N5600, N3775, N5577);
or OR4 (N5607, N5604, N1515, N204, N4095);
or OR2 (N5608, N5603, N2127);
buf BUF1 (N5609, N5601);
buf BUF1 (N5610, N5607);
xor XOR2 (N5611, N5606, N3656);
nor NOR3 (N5612, N5602, N625, N4500);
and AND2 (N5613, N5611, N1976);
xor XOR2 (N5614, N5605, N4295);
not NOT1 (N5615, N5612);
nor NOR3 (N5616, N5610, N2845, N4631);
or OR4 (N5617, N5608, N1050, N1200, N587);
buf BUF1 (N5618, N5609);
or OR3 (N5619, N5617, N4698, N4727);
not NOT1 (N5620, N5613);
and AND3 (N5621, N5599, N290, N739);
and AND2 (N5622, N5618, N5080);
and AND4 (N5623, N5598, N248, N2029, N3547);
and AND3 (N5624, N5616, N2844, N1758);
or OR3 (N5625, N5615, N2572, N361);
buf BUF1 (N5626, N5622);
or OR4 (N5627, N5623, N5251, N5189, N3473);
nand NAND2 (N5628, N5619, N3389);
not NOT1 (N5629, N5627);
xor XOR2 (N5630, N5587, N4170);
and AND3 (N5631, N5624, N1575, N3043);
and AND2 (N5632, N5620, N1102);
buf BUF1 (N5633, N5632);
not NOT1 (N5634, N5614);
and AND3 (N5635, N5633, N3799, N2202);
not NOT1 (N5636, N5629);
and AND2 (N5637, N5635, N4577);
xor XOR2 (N5638, N5637, N4520);
not NOT1 (N5639, N5631);
nor NOR4 (N5640, N5625, N4775, N4880, N133);
and AND4 (N5641, N5640, N782, N700, N2074);
not NOT1 (N5642, N5634);
not NOT1 (N5643, N5626);
nor NOR2 (N5644, N5621, N1014);
buf BUF1 (N5645, N5644);
and AND2 (N5646, N5636, N3839);
xor XOR2 (N5647, N5639, N4681);
nor NOR3 (N5648, N5641, N2643, N425);
xor XOR2 (N5649, N5638, N5010);
or OR3 (N5650, N5630, N3209, N5017);
not NOT1 (N5651, N5593);
and AND4 (N5652, N5647, N5583, N3923, N3051);
nor NOR2 (N5653, N5650, N2989);
not NOT1 (N5654, N5646);
and AND2 (N5655, N5648, N3137);
nor NOR3 (N5656, N5652, N5602, N4682);
xor XOR2 (N5657, N5653, N2898);
not NOT1 (N5658, N5655);
and AND3 (N5659, N5643, N3564, N3857);
xor XOR2 (N5660, N5656, N1647);
and AND4 (N5661, N5659, N5633, N3879, N1176);
not NOT1 (N5662, N5628);
and AND4 (N5663, N5651, N3014, N1325, N1474);
nand NAND2 (N5664, N5657, N1055);
and AND3 (N5665, N5658, N3894, N4147);
and AND3 (N5666, N5661, N4194, N2973);
and AND2 (N5667, N5665, N3084);
not NOT1 (N5668, N5645);
not NOT1 (N5669, N5649);
nand NAND3 (N5670, N5669, N2745, N5090);
or OR3 (N5671, N5667, N597, N4740);
not NOT1 (N5672, N5668);
buf BUF1 (N5673, N5672);
xor XOR2 (N5674, N5660, N5595);
xor XOR2 (N5675, N5662, N5637);
and AND4 (N5676, N5664, N4234, N4322, N5529);
and AND4 (N5677, N5673, N3576, N5492, N1093);
and AND4 (N5678, N5677, N1673, N1608, N1729);
not NOT1 (N5679, N5666);
nor NOR2 (N5680, N5671, N260);
not NOT1 (N5681, N5675);
or OR3 (N5682, N5654, N2170, N4368);
nor NOR4 (N5683, N5679, N834, N1241, N1244);
or OR3 (N5684, N5670, N3966, N4093);
buf BUF1 (N5685, N5678);
not NOT1 (N5686, N5682);
buf BUF1 (N5687, N5642);
not NOT1 (N5688, N5687);
buf BUF1 (N5689, N5685);
nand NAND4 (N5690, N5680, N830, N4259, N3577);
xor XOR2 (N5691, N5676, N1443);
or OR4 (N5692, N5683, N4418, N1872, N5184);
and AND4 (N5693, N5692, N390, N4562, N65);
xor XOR2 (N5694, N5663, N420);
xor XOR2 (N5695, N5693, N4213);
or OR3 (N5696, N5688, N2722, N5611);
nand NAND3 (N5697, N5691, N3728, N3813);
or OR2 (N5698, N5694, N3680);
nand NAND3 (N5699, N5684, N743, N5031);
nand NAND3 (N5700, N5695, N1074, N1329);
and AND4 (N5701, N5700, N5292, N2842, N4304);
xor XOR2 (N5702, N5697, N842);
xor XOR2 (N5703, N5690, N1110);
nand NAND2 (N5704, N5681, N1388);
xor XOR2 (N5705, N5702, N2119);
xor XOR2 (N5706, N5686, N1248);
and AND3 (N5707, N5696, N50, N5084);
nand NAND3 (N5708, N5704, N2298, N4578);
and AND4 (N5709, N5703, N4298, N2802, N75);
nand NAND4 (N5710, N5707, N32, N2579, N2673);
nand NAND2 (N5711, N5710, N5213);
nand NAND3 (N5712, N5689, N3060, N3665);
nand NAND2 (N5713, N5674, N5701);
and AND2 (N5714, N5602, N2980);
nand NAND2 (N5715, N5709, N3899);
buf BUF1 (N5716, N5711);
xor XOR2 (N5717, N5698, N58);
nor NOR3 (N5718, N5716, N5703, N911);
and AND2 (N5719, N5705, N5694);
xor XOR2 (N5720, N5718, N5051);
nand NAND4 (N5721, N5699, N2669, N2556, N828);
and AND4 (N5722, N5717, N1105, N885, N2305);
or OR3 (N5723, N5713, N3000, N4518);
or OR4 (N5724, N5714, N751, N2785, N5545);
and AND2 (N5725, N5715, N703);
nand NAND2 (N5726, N5712, N3232);
not NOT1 (N5727, N5708);
or OR4 (N5728, N5726, N4212, N579, N1883);
not NOT1 (N5729, N5723);
and AND4 (N5730, N5721, N272, N3592, N615);
not NOT1 (N5731, N5722);
nor NOR4 (N5732, N5731, N2649, N1013, N2529);
nand NAND3 (N5733, N5720, N581, N2877);
or OR2 (N5734, N5730, N28);
nand NAND2 (N5735, N5725, N361);
xor XOR2 (N5736, N5734, N4582);
buf BUF1 (N5737, N5736);
xor XOR2 (N5738, N5733, N2647);
not NOT1 (N5739, N5727);
nor NOR3 (N5740, N5728, N2387, N3511);
buf BUF1 (N5741, N5729);
not NOT1 (N5742, N5724);
xor XOR2 (N5743, N5706, N654);
not NOT1 (N5744, N5743);
or OR4 (N5745, N5741, N320, N1956, N226);
and AND2 (N5746, N5742, N5086);
xor XOR2 (N5747, N5719, N2532);
buf BUF1 (N5748, N5739);
and AND2 (N5749, N5738, N730);
xor XOR2 (N5750, N5749, N4778);
and AND3 (N5751, N5737, N2751, N3755);
nor NOR4 (N5752, N5745, N4172, N3557, N5587);
or OR3 (N5753, N5746, N4265, N3287);
and AND4 (N5754, N5752, N1167, N3610, N649);
not NOT1 (N5755, N5753);
nand NAND3 (N5756, N5747, N4064, N3599);
not NOT1 (N5757, N5750);
buf BUF1 (N5758, N5744);
xor XOR2 (N5759, N5740, N5182);
and AND4 (N5760, N5755, N5514, N861, N4077);
nor NOR3 (N5761, N5748, N2885, N4548);
nand NAND4 (N5762, N5732, N3216, N3377, N5645);
and AND4 (N5763, N5754, N2569, N3763, N3180);
nor NOR4 (N5764, N5761, N836, N2511, N2708);
and AND2 (N5765, N5757, N1122);
buf BUF1 (N5766, N5762);
nand NAND4 (N5767, N5760, N4466, N5258, N4763);
not NOT1 (N5768, N5766);
or OR2 (N5769, N5756, N3893);
nor NOR4 (N5770, N5735, N308, N3594, N2072);
buf BUF1 (N5771, N5770);
xor XOR2 (N5772, N5764, N1266);
not NOT1 (N5773, N5772);
buf BUF1 (N5774, N5773);
not NOT1 (N5775, N5767);
and AND4 (N5776, N5751, N639, N729, N4795);
xor XOR2 (N5777, N5776, N4927);
nor NOR3 (N5778, N5768, N1036, N5638);
nor NOR3 (N5779, N5774, N3055, N95);
nand NAND3 (N5780, N5771, N1155, N4132);
nand NAND3 (N5781, N5778, N5738, N629);
or OR4 (N5782, N5781, N765, N499, N2714);
nand NAND2 (N5783, N5775, N649);
nor NOR2 (N5784, N5779, N3825);
nor NOR4 (N5785, N5758, N2306, N3763, N4408);
nand NAND2 (N5786, N5780, N2255);
or OR4 (N5787, N5784, N3394, N1223, N4815);
buf BUF1 (N5788, N5769);
nor NOR4 (N5789, N5787, N2342, N136, N3335);
or OR4 (N5790, N5763, N128, N3193, N3793);
or OR3 (N5791, N5788, N764, N3493);
xor XOR2 (N5792, N5789, N3653);
not NOT1 (N5793, N5783);
not NOT1 (N5794, N5777);
not NOT1 (N5795, N5793);
not NOT1 (N5796, N5791);
and AND4 (N5797, N5795, N3349, N886, N827);
not NOT1 (N5798, N5794);
or OR3 (N5799, N5765, N191, N547);
nand NAND2 (N5800, N5796, N4268);
buf BUF1 (N5801, N5800);
nor NOR2 (N5802, N5801, N4020);
buf BUF1 (N5803, N5798);
not NOT1 (N5804, N5790);
or OR2 (N5805, N5759, N2099);
or OR3 (N5806, N5792, N2313, N5330);
nor NOR3 (N5807, N5803, N821, N4448);
not NOT1 (N5808, N5805);
not NOT1 (N5809, N5806);
or OR2 (N5810, N5802, N3698);
nand NAND4 (N5811, N5804, N4373, N4509, N5117);
not NOT1 (N5812, N5807);
and AND4 (N5813, N5810, N3410, N63, N2325);
buf BUF1 (N5814, N5812);
xor XOR2 (N5815, N5813, N5049);
not NOT1 (N5816, N5811);
or OR2 (N5817, N5785, N1463);
xor XOR2 (N5818, N5808, N1470);
not NOT1 (N5819, N5818);
not NOT1 (N5820, N5817);
nor NOR4 (N5821, N5819, N5431, N5445, N4782);
or OR3 (N5822, N5799, N851, N982);
not NOT1 (N5823, N5821);
not NOT1 (N5824, N5822);
and AND4 (N5825, N5823, N795, N2159, N506);
xor XOR2 (N5826, N5786, N5622);
nor NOR3 (N5827, N5816, N5206, N795);
or OR4 (N5828, N5797, N3283, N3790, N1263);
not NOT1 (N5829, N5827);
xor XOR2 (N5830, N5814, N2323);
nor NOR4 (N5831, N5829, N586, N2420, N4768);
buf BUF1 (N5832, N5820);
xor XOR2 (N5833, N5809, N1506);
nand NAND2 (N5834, N5833, N5396);
nand NAND2 (N5835, N5834, N1351);
not NOT1 (N5836, N5828);
or OR2 (N5837, N5830, N2619);
not NOT1 (N5838, N5782);
xor XOR2 (N5839, N5836, N3137);
or OR2 (N5840, N5839, N4484);
nor NOR3 (N5841, N5838, N4137, N5313);
nor NOR3 (N5842, N5826, N31, N4228);
or OR3 (N5843, N5815, N5833, N1377);
nand NAND2 (N5844, N5831, N1511);
not NOT1 (N5845, N5824);
nand NAND2 (N5846, N5845, N4553);
and AND4 (N5847, N5837, N1148, N2025, N1289);
or OR3 (N5848, N5844, N789, N2205);
not NOT1 (N5849, N5842);
nand NAND3 (N5850, N5848, N2873, N2515);
nand NAND4 (N5851, N5847, N3445, N3666, N5207);
nor NOR2 (N5852, N5840, N1534);
nand NAND3 (N5853, N5825, N5282, N2021);
buf BUF1 (N5854, N5835);
xor XOR2 (N5855, N5852, N3699);
not NOT1 (N5856, N5846);
or OR4 (N5857, N5854, N937, N954, N2589);
not NOT1 (N5858, N5855);
buf BUF1 (N5859, N5857);
not NOT1 (N5860, N5832);
nor NOR4 (N5861, N5856, N2496, N1561, N3097);
buf BUF1 (N5862, N5859);
xor XOR2 (N5863, N5849, N4675);
and AND2 (N5864, N5861, N325);
nand NAND2 (N5865, N5858, N3947);
not NOT1 (N5866, N5851);
xor XOR2 (N5867, N5862, N3722);
nand NAND2 (N5868, N5843, N402);
or OR4 (N5869, N5868, N79, N2985, N4690);
buf BUF1 (N5870, N5863);
nor NOR3 (N5871, N5850, N3241, N4805);
not NOT1 (N5872, N5860);
xor XOR2 (N5873, N5871, N3623);
not NOT1 (N5874, N5869);
or OR4 (N5875, N5870, N2595, N4702, N1093);
xor XOR2 (N5876, N5865, N3841);
buf BUF1 (N5877, N5853);
nand NAND2 (N5878, N5872, N3730);
xor XOR2 (N5879, N5876, N180);
buf BUF1 (N5880, N5879);
buf BUF1 (N5881, N5873);
nor NOR2 (N5882, N5881, N2744);
buf BUF1 (N5883, N5882);
not NOT1 (N5884, N5874);
not NOT1 (N5885, N5864);
and AND2 (N5886, N5884, N4716);
xor XOR2 (N5887, N5877, N1302);
and AND2 (N5888, N5887, N3723);
buf BUF1 (N5889, N5878);
nor NOR2 (N5890, N5841, N3398);
or OR2 (N5891, N5867, N62);
nor NOR4 (N5892, N5875, N3544, N1983, N4938);
nand NAND2 (N5893, N5880, N4317);
and AND3 (N5894, N5886, N504, N3062);
or OR3 (N5895, N5890, N3508, N1275);
xor XOR2 (N5896, N5893, N3483);
not NOT1 (N5897, N5896);
nor NOR2 (N5898, N5895, N3492);
buf BUF1 (N5899, N5897);
or OR4 (N5900, N5885, N2544, N3420, N3963);
xor XOR2 (N5901, N5894, N863);
nor NOR4 (N5902, N5883, N4071, N2274, N2806);
buf BUF1 (N5903, N5891);
nand NAND3 (N5904, N5892, N5710, N1427);
not NOT1 (N5905, N5898);
not NOT1 (N5906, N5904);
and AND3 (N5907, N5866, N5397, N1066);
or OR3 (N5908, N5906, N5487, N3682);
or OR2 (N5909, N5903, N4106);
nor NOR4 (N5910, N5889, N5623, N2779, N3389);
not NOT1 (N5911, N5888);
xor XOR2 (N5912, N5908, N197);
or OR2 (N5913, N5900, N877);
nor NOR4 (N5914, N5907, N3596, N5006, N1190);
nand NAND3 (N5915, N5902, N498, N97);
not NOT1 (N5916, N5912);
not NOT1 (N5917, N5905);
nand NAND4 (N5918, N5911, N5368, N2878, N4234);
not NOT1 (N5919, N5913);
and AND4 (N5920, N5915, N2003, N3266, N5239);
nor NOR3 (N5921, N5910, N4042, N4286);
nand NAND2 (N5922, N5917, N5130);
and AND2 (N5923, N5901, N2419);
nand NAND3 (N5924, N5899, N4827, N5434);
and AND2 (N5925, N5921, N3839);
nand NAND3 (N5926, N5923, N2926, N2495);
and AND3 (N5927, N5914, N1132, N2632);
nand NAND2 (N5928, N5924, N1695);
xor XOR2 (N5929, N5909, N3106);
xor XOR2 (N5930, N5928, N104);
buf BUF1 (N5931, N5927);
not NOT1 (N5932, N5916);
nor NOR3 (N5933, N5919, N3818, N571);
buf BUF1 (N5934, N5931);
buf BUF1 (N5935, N5925);
and AND4 (N5936, N5918, N68, N483, N3510);
nor NOR2 (N5937, N5922, N2493);
nor NOR2 (N5938, N5926, N5336);
not NOT1 (N5939, N5937);
nor NOR4 (N5940, N5934, N4096, N2427, N2437);
and AND4 (N5941, N5932, N2502, N2315, N781);
nand NAND2 (N5942, N5929, N2473);
xor XOR2 (N5943, N5936, N1677);
not NOT1 (N5944, N5943);
not NOT1 (N5945, N5930);
nand NAND3 (N5946, N5944, N4167, N4958);
nor NOR3 (N5947, N5942, N1188, N4226);
and AND3 (N5948, N5946, N3422, N4526);
not NOT1 (N5949, N5947);
nand NAND4 (N5950, N5935, N1861, N4530, N4737);
nand NAND4 (N5951, N5948, N3579, N2020, N5259);
buf BUF1 (N5952, N5949);
nand NAND2 (N5953, N5945, N443);
and AND4 (N5954, N5939, N3344, N5792, N3270);
and AND4 (N5955, N5950, N580, N3322, N3160);
buf BUF1 (N5956, N5920);
buf BUF1 (N5957, N5953);
xor XOR2 (N5958, N5940, N3459);
or OR2 (N5959, N5933, N383);
nor NOR2 (N5960, N5941, N2668);
nor NOR3 (N5961, N5938, N3858, N2111);
or OR2 (N5962, N5951, N4007);
not NOT1 (N5963, N5961);
nor NOR4 (N5964, N5962, N2497, N414, N1342);
xor XOR2 (N5965, N5957, N5163);
and AND3 (N5966, N5965, N3231, N938);
and AND2 (N5967, N5954, N5484);
buf BUF1 (N5968, N5966);
nand NAND3 (N5969, N5955, N1753, N5118);
or OR4 (N5970, N5958, N1543, N2170, N2003);
or OR4 (N5971, N5968, N839, N3491, N933);
nor NOR2 (N5972, N5952, N549);
not NOT1 (N5973, N5967);
buf BUF1 (N5974, N5956);
and AND2 (N5975, N5969, N5210);
and AND3 (N5976, N5964, N737, N1499);
xor XOR2 (N5977, N5970, N3340);
or OR3 (N5978, N5971, N5478, N1601);
xor XOR2 (N5979, N5959, N3498);
xor XOR2 (N5980, N5974, N5625);
and AND4 (N5981, N5963, N3078, N429, N2297);
or OR4 (N5982, N5976, N704, N5181, N3643);
not NOT1 (N5983, N5979);
or OR3 (N5984, N5981, N3234, N2728);
and AND2 (N5985, N5975, N3838);
nand NAND3 (N5986, N5984, N4494, N3570);
nand NAND3 (N5987, N5986, N5155, N5104);
and AND2 (N5988, N5980, N2213);
buf BUF1 (N5989, N5977);
buf BUF1 (N5990, N5972);
nand NAND2 (N5991, N5989, N326);
buf BUF1 (N5992, N5991);
and AND3 (N5993, N5973, N1054, N5004);
nand NAND2 (N5994, N5985, N3201);
nand NAND3 (N5995, N5988, N3338, N2952);
nand NAND4 (N5996, N5990, N3884, N2795, N2399);
and AND2 (N5997, N5994, N3736);
buf BUF1 (N5998, N5987);
and AND2 (N5999, N5992, N838);
and AND4 (N6000, N5982, N1793, N4528, N1310);
xor XOR2 (N6001, N5960, N3956);
nor NOR4 (N6002, N5999, N4975, N1300, N4958);
or OR2 (N6003, N6002, N4624);
not NOT1 (N6004, N5993);
and AND3 (N6005, N6001, N347, N901);
buf BUF1 (N6006, N6005);
not NOT1 (N6007, N6004);
nand NAND4 (N6008, N6003, N3172, N1733, N1498);
and AND4 (N6009, N6006, N4336, N736, N3293);
nor NOR3 (N6010, N5978, N2657, N5713);
not NOT1 (N6011, N6008);
and AND2 (N6012, N6010, N5902);
nor NOR3 (N6013, N6009, N1880, N3818);
or OR2 (N6014, N6012, N3987);
nand NAND2 (N6015, N5996, N3027);
nor NOR4 (N6016, N5997, N4067, N2016, N2986);
not NOT1 (N6017, N6007);
nor NOR2 (N6018, N6000, N45);
nor NOR4 (N6019, N6014, N2500, N4015, N2041);
nor NOR2 (N6020, N5983, N2225);
buf BUF1 (N6021, N6018);
xor XOR2 (N6022, N6016, N3678);
and AND3 (N6023, N5995, N1723, N1391);
not NOT1 (N6024, N5998);
buf BUF1 (N6025, N6013);
nor NOR2 (N6026, N6015, N2445);
or OR2 (N6027, N6025, N5476);
buf BUF1 (N6028, N6023);
xor XOR2 (N6029, N6011, N2174);
or OR4 (N6030, N6024, N2119, N642, N5088);
nand NAND2 (N6031, N6020, N1317);
nor NOR4 (N6032, N6022, N2747, N1552, N5341);
nor NOR3 (N6033, N6030, N1263, N2069);
xor XOR2 (N6034, N6033, N3579);
buf BUF1 (N6035, N6028);
buf BUF1 (N6036, N6035);
not NOT1 (N6037, N6029);
and AND3 (N6038, N6027, N811, N2201);
not NOT1 (N6039, N6019);
buf BUF1 (N6040, N6039);
not NOT1 (N6041, N6040);
buf BUF1 (N6042, N6037);
not NOT1 (N6043, N6021);
or OR3 (N6044, N6043, N4994, N5073);
or OR2 (N6045, N6017, N1291);
nor NOR2 (N6046, N6036, N294);
nor NOR3 (N6047, N6031, N3224, N5880);
xor XOR2 (N6048, N6026, N842);
buf BUF1 (N6049, N6041);
nand NAND2 (N6050, N6038, N2270);
not NOT1 (N6051, N6048);
nand NAND4 (N6052, N6042, N1902, N456, N4576);
xor XOR2 (N6053, N6034, N2940);
or OR2 (N6054, N6053, N4273);
nand NAND4 (N6055, N6032, N1489, N4011, N2991);
nand NAND3 (N6056, N6045, N4626, N1854);
not NOT1 (N6057, N6054);
xor XOR2 (N6058, N6044, N4615);
nand NAND4 (N6059, N6047, N5716, N2738, N5252);
or OR4 (N6060, N6056, N2292, N4900, N5550);
or OR4 (N6061, N6051, N5689, N5095, N1183);
not NOT1 (N6062, N6061);
nand NAND3 (N6063, N6052, N5036, N1413);
buf BUF1 (N6064, N6055);
and AND4 (N6065, N6060, N2184, N5060, N5432);
and AND4 (N6066, N6058, N3360, N3113, N3162);
buf BUF1 (N6067, N6064);
nor NOR3 (N6068, N6063, N1523, N5199);
or OR3 (N6069, N6067, N4702, N3967);
nand NAND4 (N6070, N6065, N987, N1838, N2614);
xor XOR2 (N6071, N6069, N1059);
or OR2 (N6072, N6049, N5962);
not NOT1 (N6073, N6070);
buf BUF1 (N6074, N6050);
or OR2 (N6075, N6046, N447);
buf BUF1 (N6076, N6075);
buf BUF1 (N6077, N6059);
xor XOR2 (N6078, N6076, N1997);
buf BUF1 (N6079, N6073);
not NOT1 (N6080, N6071);
not NOT1 (N6081, N6079);
xor XOR2 (N6082, N6072, N3534);
not NOT1 (N6083, N6080);
xor XOR2 (N6084, N6068, N1721);
nand NAND4 (N6085, N6057, N4800, N3137, N1020);
xor XOR2 (N6086, N6066, N4796);
and AND2 (N6087, N6083, N4277);
or OR3 (N6088, N6078, N2273, N932);
xor XOR2 (N6089, N6074, N182);
xor XOR2 (N6090, N6089, N1271);
xor XOR2 (N6091, N6086, N3753);
or OR2 (N6092, N6077, N5678);
or OR4 (N6093, N6084, N5082, N5536, N113);
and AND3 (N6094, N6088, N5962, N2520);
xor XOR2 (N6095, N6093, N1869);
nand NAND4 (N6096, N6062, N6019, N1422, N4571);
xor XOR2 (N6097, N6082, N4590);
buf BUF1 (N6098, N6081);
or OR4 (N6099, N6085, N1879, N1180, N4037);
xor XOR2 (N6100, N6097, N2490);
not NOT1 (N6101, N6087);
buf BUF1 (N6102, N6100);
nor NOR3 (N6103, N6096, N2955, N3977);
nor NOR4 (N6104, N6103, N5171, N1468, N4525);
xor XOR2 (N6105, N6090, N5182);
xor XOR2 (N6106, N6098, N5209);
buf BUF1 (N6107, N6102);
not NOT1 (N6108, N6104);
nor NOR2 (N6109, N6105, N1240);
xor XOR2 (N6110, N6109, N2655);
or OR4 (N6111, N6107, N1350, N2729, N485);
nand NAND3 (N6112, N6106, N3570, N254);
nor NOR2 (N6113, N6099, N903);
or OR3 (N6114, N6101, N1847, N5448);
nor NOR2 (N6115, N6111, N4814);
and AND2 (N6116, N6110, N5156);
nor NOR2 (N6117, N6115, N439);
or OR4 (N6118, N6117, N4130, N4430, N4170);
not NOT1 (N6119, N6114);
not NOT1 (N6120, N6118);
nand NAND3 (N6121, N6091, N1201, N4383);
and AND4 (N6122, N6120, N1095, N4425, N3644);
nor NOR3 (N6123, N6113, N5797, N5101);
or OR3 (N6124, N6122, N5858, N3981);
nor NOR4 (N6125, N6121, N81, N5631, N5105);
xor XOR2 (N6126, N6116, N527);
buf BUF1 (N6127, N6092);
nor NOR2 (N6128, N6124, N2033);
nor NOR3 (N6129, N6128, N1101, N5653);
nor NOR2 (N6130, N6112, N934);
nor NOR4 (N6131, N6130, N3129, N1216, N2074);
and AND2 (N6132, N6095, N4052);
not NOT1 (N6133, N6108);
or OR3 (N6134, N6094, N920, N6003);
or OR3 (N6135, N6123, N3758, N3047);
xor XOR2 (N6136, N6132, N4986);
or OR4 (N6137, N6127, N4025, N2875, N206);
nor NOR2 (N6138, N6137, N445);
and AND2 (N6139, N6133, N692);
nor NOR3 (N6140, N6131, N3309, N2377);
xor XOR2 (N6141, N6136, N1662);
nand NAND4 (N6142, N6140, N2211, N3155, N1695);
nor NOR2 (N6143, N6119, N4795);
nor NOR3 (N6144, N6138, N3625, N4295);
or OR4 (N6145, N6129, N4090, N190, N1287);
nor NOR3 (N6146, N6144, N1071, N5248);
not NOT1 (N6147, N6146);
nor NOR2 (N6148, N6142, N4048);
buf BUF1 (N6149, N6148);
nand NAND4 (N6150, N6149, N4913, N5447, N3151);
nor NOR4 (N6151, N6134, N5452, N3, N4413);
nor NOR3 (N6152, N6143, N4807, N656);
nand NAND2 (N6153, N6147, N3325);
buf BUF1 (N6154, N6125);
or OR2 (N6155, N6151, N269);
not NOT1 (N6156, N6154);
and AND2 (N6157, N6145, N3939);
buf BUF1 (N6158, N6139);
xor XOR2 (N6159, N6135, N3241);
xor XOR2 (N6160, N6156, N2010);
or OR4 (N6161, N6141, N5863, N3573, N2892);
nor NOR4 (N6162, N6155, N5641, N4166, N1228);
not NOT1 (N6163, N6150);
xor XOR2 (N6164, N6160, N5170);
not NOT1 (N6165, N6153);
not NOT1 (N6166, N6163);
and AND4 (N6167, N6165, N3947, N178, N4577);
xor XOR2 (N6168, N6152, N2204);
xor XOR2 (N6169, N6167, N632);
buf BUF1 (N6170, N6159);
not NOT1 (N6171, N6157);
buf BUF1 (N6172, N6166);
nor NOR4 (N6173, N6169, N819, N3497, N503);
and AND4 (N6174, N6161, N2795, N3658, N3419);
nand NAND3 (N6175, N6170, N3932, N3448);
and AND4 (N6176, N6175, N4709, N1238, N3812);
xor XOR2 (N6177, N6162, N704);
nand NAND3 (N6178, N6171, N568, N3595);
buf BUF1 (N6179, N6168);
buf BUF1 (N6180, N6172);
buf BUF1 (N6181, N6179);
nor NOR3 (N6182, N6180, N5292, N4924);
not NOT1 (N6183, N6164);
nand NAND4 (N6184, N6177, N4814, N1919, N1175);
or OR2 (N6185, N6181, N2837);
nor NOR2 (N6186, N6174, N3563);
xor XOR2 (N6187, N6186, N5885);
not NOT1 (N6188, N6126);
and AND2 (N6189, N6176, N965);
nand NAND2 (N6190, N6182, N5107);
or OR2 (N6191, N6187, N80);
not NOT1 (N6192, N6184);
xor XOR2 (N6193, N6189, N1447);
and AND4 (N6194, N6178, N4687, N6025, N2124);
xor XOR2 (N6195, N6193, N3343);
nand NAND2 (N6196, N6183, N1945);
and AND3 (N6197, N6185, N1016, N2945);
nand NAND2 (N6198, N6195, N3642);
not NOT1 (N6199, N6188);
nor NOR4 (N6200, N6198, N4527, N181, N818);
nand NAND4 (N6201, N6200, N148, N6068, N5300);
nand NAND2 (N6202, N6190, N1946);
and AND2 (N6203, N6202, N5573);
and AND3 (N6204, N6197, N1417, N2355);
nor NOR4 (N6205, N6173, N5105, N2669, N3717);
nor NOR4 (N6206, N6203, N4643, N1558, N863);
not NOT1 (N6207, N6158);
and AND3 (N6208, N6204, N632, N1009);
not NOT1 (N6209, N6208);
buf BUF1 (N6210, N6199);
not NOT1 (N6211, N6210);
not NOT1 (N6212, N6207);
buf BUF1 (N6213, N6205);
nor NOR3 (N6214, N6209, N643, N4171);
and AND4 (N6215, N6192, N1976, N5910, N6169);
not NOT1 (N6216, N6191);
xor XOR2 (N6217, N6201, N2488);
not NOT1 (N6218, N6212);
nand NAND4 (N6219, N6196, N5403, N2634, N1260);
not NOT1 (N6220, N6216);
or OR2 (N6221, N6211, N4430);
nand NAND4 (N6222, N6194, N5865, N5866, N4606);
or OR3 (N6223, N6221, N5649, N3591);
xor XOR2 (N6224, N6213, N1288);
nor NOR4 (N6225, N6214, N1957, N1819, N5954);
nand NAND2 (N6226, N6217, N2912);
xor XOR2 (N6227, N6215, N5763);
nand NAND2 (N6228, N6227, N5377);
nor NOR4 (N6229, N6206, N4688, N5965, N920);
nor NOR4 (N6230, N6222, N1415, N3958, N3003);
not NOT1 (N6231, N6229);
xor XOR2 (N6232, N6218, N1617);
or OR4 (N6233, N6230, N1137, N5639, N5994);
buf BUF1 (N6234, N6223);
nand NAND3 (N6235, N6234, N5160, N6061);
not NOT1 (N6236, N6228);
buf BUF1 (N6237, N6219);
xor XOR2 (N6238, N6225, N16);
or OR4 (N6239, N6232, N2662, N980, N470);
not NOT1 (N6240, N6220);
not NOT1 (N6241, N6235);
or OR3 (N6242, N6241, N4365, N2416);
not NOT1 (N6243, N6236);
not NOT1 (N6244, N6233);
nand NAND2 (N6245, N6231, N784);
not NOT1 (N6246, N6240);
xor XOR2 (N6247, N6224, N352);
nor NOR3 (N6248, N6244, N6130, N3408);
and AND3 (N6249, N6238, N2379, N3396);
and AND3 (N6250, N6245, N3707, N2931);
nand NAND2 (N6251, N6226, N4784);
buf BUF1 (N6252, N6250);
and AND4 (N6253, N6252, N3559, N5614, N3734);
nand NAND2 (N6254, N6239, N3317);
not NOT1 (N6255, N6243);
nor NOR2 (N6256, N6246, N1152);
xor XOR2 (N6257, N6247, N4350);
xor XOR2 (N6258, N6242, N5864);
or OR4 (N6259, N6237, N1974, N134, N2530);
nand NAND4 (N6260, N6258, N2759, N739, N5273);
and AND2 (N6261, N6255, N2373);
nand NAND2 (N6262, N6256, N3809);
nand NAND4 (N6263, N6249, N1135, N1386, N3139);
buf BUF1 (N6264, N6251);
nand NAND2 (N6265, N6257, N5390);
nor NOR3 (N6266, N6260, N4878, N4619);
nor NOR4 (N6267, N6248, N5736, N4332, N6145);
xor XOR2 (N6268, N6265, N3508);
xor XOR2 (N6269, N6268, N2333);
nand NAND4 (N6270, N6253, N5239, N2392, N3959);
not NOT1 (N6271, N6269);
xor XOR2 (N6272, N6262, N5307);
nor NOR4 (N6273, N6263, N2565, N1380, N6137);
nor NOR4 (N6274, N6270, N481, N3103, N291);
or OR4 (N6275, N6266, N5621, N5534, N2921);
xor XOR2 (N6276, N6274, N2978);
buf BUF1 (N6277, N6275);
not NOT1 (N6278, N6271);
nor NOR4 (N6279, N6277, N1785, N6127, N99);
nor NOR2 (N6280, N6279, N5075);
buf BUF1 (N6281, N6273);
or OR4 (N6282, N6267, N3141, N2882, N3837);
nand NAND2 (N6283, N6276, N3397);
nor NOR2 (N6284, N6280, N2732);
not NOT1 (N6285, N6284);
and AND3 (N6286, N6259, N4397, N2434);
nand NAND2 (N6287, N6264, N1185);
nand NAND4 (N6288, N6286, N5840, N5523, N901);
and AND3 (N6289, N6285, N1317, N333);
xor XOR2 (N6290, N6278, N1869);
or OR2 (N6291, N6283, N416);
buf BUF1 (N6292, N6290);
or OR4 (N6293, N6287, N3638, N475, N2721);
xor XOR2 (N6294, N6261, N4559);
xor XOR2 (N6295, N6272, N2380);
xor XOR2 (N6296, N6288, N3340);
buf BUF1 (N6297, N6254);
not NOT1 (N6298, N6294);
not NOT1 (N6299, N6293);
and AND4 (N6300, N6281, N3929, N2935, N5740);
nand NAND4 (N6301, N6296, N2637, N4449, N552);
nor NOR2 (N6302, N6289, N2012);
nand NAND4 (N6303, N6282, N5913, N2256, N2196);
not NOT1 (N6304, N6300);
and AND4 (N6305, N6303, N1830, N1288, N4357);
nor NOR3 (N6306, N6302, N6088, N5240);
nor NOR3 (N6307, N6297, N4731, N4410);
xor XOR2 (N6308, N6301, N3390);
and AND2 (N6309, N6298, N3373);
and AND3 (N6310, N6306, N295, N5147);
buf BUF1 (N6311, N6307);
and AND4 (N6312, N6291, N6051, N179, N4774);
nand NAND2 (N6313, N6305, N3178);
nand NAND2 (N6314, N6310, N3903);
nor NOR2 (N6315, N6311, N688);
nand NAND4 (N6316, N6315, N2340, N4206, N5834);
nor NOR3 (N6317, N6295, N1489, N812);
nand NAND3 (N6318, N6313, N2082, N4167);
or OR2 (N6319, N6309, N1322);
not NOT1 (N6320, N6314);
xor XOR2 (N6321, N6316, N5466);
nand NAND4 (N6322, N6318, N943, N1963, N3063);
and AND2 (N6323, N6299, N1571);
xor XOR2 (N6324, N6292, N6253);
not NOT1 (N6325, N6323);
buf BUF1 (N6326, N6321);
nand NAND3 (N6327, N6324, N3434, N1328);
not NOT1 (N6328, N6319);
or OR3 (N6329, N6308, N4923, N613);
and AND4 (N6330, N6327, N5371, N5749, N3340);
not NOT1 (N6331, N6329);
and AND2 (N6332, N6328, N6036);
nor NOR2 (N6333, N6325, N5252);
not NOT1 (N6334, N6304);
xor XOR2 (N6335, N6330, N2882);
nand NAND2 (N6336, N6317, N5710);
buf BUF1 (N6337, N6312);
not NOT1 (N6338, N6333);
nor NOR2 (N6339, N6337, N1935);
nand NAND2 (N6340, N6326, N4725);
nor NOR3 (N6341, N6332, N2219, N5332);
or OR2 (N6342, N6340, N5184);
not NOT1 (N6343, N6335);
or OR3 (N6344, N6334, N5274, N492);
and AND4 (N6345, N6331, N6099, N4446, N76);
or OR4 (N6346, N6341, N4282, N3157, N2946);
buf BUF1 (N6347, N6345);
nand NAND3 (N6348, N6343, N4590, N5143);
not NOT1 (N6349, N6322);
buf BUF1 (N6350, N6339);
nor NOR2 (N6351, N6347, N2840);
buf BUF1 (N6352, N6336);
and AND2 (N6353, N6338, N4184);
nand NAND4 (N6354, N6353, N433, N5401, N4679);
nand NAND3 (N6355, N6352, N726, N1048);
buf BUF1 (N6356, N6342);
or OR3 (N6357, N6350, N2279, N6164);
not NOT1 (N6358, N6348);
xor XOR2 (N6359, N6346, N2981);
xor XOR2 (N6360, N6355, N2604);
buf BUF1 (N6361, N6358);
or OR2 (N6362, N6349, N6344);
xor XOR2 (N6363, N5908, N2120);
nand NAND4 (N6364, N6362, N1406, N75, N5762);
xor XOR2 (N6365, N6361, N5448);
buf BUF1 (N6366, N6359);
or OR4 (N6367, N6360, N1573, N4281, N4163);
xor XOR2 (N6368, N6365, N2035);
nand NAND2 (N6369, N6363, N3120);
buf BUF1 (N6370, N6356);
or OR2 (N6371, N6368, N86);
nor NOR2 (N6372, N6371, N5957);
xor XOR2 (N6373, N6367, N2359);
xor XOR2 (N6374, N6351, N1350);
nor NOR4 (N6375, N6354, N2352, N756, N4649);
xor XOR2 (N6376, N6373, N5474);
nor NOR4 (N6377, N6376, N2522, N3923, N265);
buf BUF1 (N6378, N6357);
or OR4 (N6379, N6370, N1644, N5394, N2114);
not NOT1 (N6380, N6374);
nand NAND2 (N6381, N6366, N2799);
not NOT1 (N6382, N6369);
nor NOR3 (N6383, N6379, N4103, N3845);
or OR4 (N6384, N6375, N6058, N1647, N3918);
buf BUF1 (N6385, N6372);
not NOT1 (N6386, N6380);
nand NAND2 (N6387, N6386, N4762);
nor NOR2 (N6388, N6384, N491);
and AND4 (N6389, N6364, N3064, N4456, N151);
or OR2 (N6390, N6320, N4062);
buf BUF1 (N6391, N6387);
not NOT1 (N6392, N6391);
nand NAND2 (N6393, N6383, N1287);
and AND2 (N6394, N6392, N5762);
and AND3 (N6395, N6377, N556, N2598);
nand NAND4 (N6396, N6395, N6060, N5671, N5979);
and AND3 (N6397, N6378, N2176, N243);
not NOT1 (N6398, N6389);
buf BUF1 (N6399, N6390);
or OR3 (N6400, N6396, N4865, N2518);
nor NOR3 (N6401, N6382, N1197, N5764);
nand NAND3 (N6402, N6385, N1831, N4734);
and AND3 (N6403, N6381, N3711, N5077);
nor NOR3 (N6404, N6398, N5768, N5631);
nor NOR4 (N6405, N6400, N2433, N2419, N705);
xor XOR2 (N6406, N6402, N326);
or OR4 (N6407, N6394, N1750, N3213, N2170);
or OR4 (N6408, N6407, N5247, N2771, N946);
and AND4 (N6409, N6397, N5080, N3200, N3215);
or OR3 (N6410, N6403, N3342, N5898);
or OR2 (N6411, N6406, N569);
buf BUF1 (N6412, N6410);
buf BUF1 (N6413, N6401);
xor XOR2 (N6414, N6388, N2962);
and AND3 (N6415, N6405, N3263, N3837);
not NOT1 (N6416, N6393);
nor NOR3 (N6417, N6412, N3437, N6337);
nand NAND3 (N6418, N6399, N6196, N762);
not NOT1 (N6419, N6417);
xor XOR2 (N6420, N6409, N5020);
nor NOR3 (N6421, N6415, N458, N599);
nor NOR2 (N6422, N6413, N2911);
nor NOR2 (N6423, N6421, N703);
buf BUF1 (N6424, N6418);
buf BUF1 (N6425, N6416);
not NOT1 (N6426, N6414);
xor XOR2 (N6427, N6426, N3190);
nor NOR4 (N6428, N6427, N4226, N4166, N4338);
nand NAND2 (N6429, N6423, N4559);
and AND3 (N6430, N6420, N1580, N4349);
xor XOR2 (N6431, N6429, N1908);
buf BUF1 (N6432, N6422);
xor XOR2 (N6433, N6431, N1739);
buf BUF1 (N6434, N6408);
and AND2 (N6435, N6425, N3483);
buf BUF1 (N6436, N6433);
and AND4 (N6437, N6434, N1344, N1136, N1888);
xor XOR2 (N6438, N6430, N2577);
buf BUF1 (N6439, N6432);
not NOT1 (N6440, N6428);
buf BUF1 (N6441, N6435);
xor XOR2 (N6442, N6436, N5920);
or OR4 (N6443, N6440, N2734, N2871, N2082);
not NOT1 (N6444, N6424);
xor XOR2 (N6445, N6404, N2160);
not NOT1 (N6446, N6439);
or OR3 (N6447, N6444, N631, N4438);
xor XOR2 (N6448, N6445, N2313);
not NOT1 (N6449, N6419);
and AND3 (N6450, N6442, N3010, N6149);
nand NAND4 (N6451, N6450, N1191, N5546, N3491);
and AND3 (N6452, N6448, N5680, N5753);
or OR2 (N6453, N6437, N2959);
buf BUF1 (N6454, N6447);
buf BUF1 (N6455, N6438);
xor XOR2 (N6456, N6446, N1024);
and AND4 (N6457, N6452, N3795, N4778, N3859);
not NOT1 (N6458, N6441);
xor XOR2 (N6459, N6457, N4283);
and AND4 (N6460, N6443, N1079, N806, N4250);
xor XOR2 (N6461, N6453, N1722);
or OR3 (N6462, N6451, N5077, N4577);
not NOT1 (N6463, N6462);
xor XOR2 (N6464, N6459, N2318);
nor NOR4 (N6465, N6456, N1753, N1815, N2418);
nor NOR4 (N6466, N6464, N2259, N13, N4096);
not NOT1 (N6467, N6461);
nor NOR2 (N6468, N6455, N4590);
buf BUF1 (N6469, N6411);
nor NOR4 (N6470, N6460, N1938, N6387, N3567);
buf BUF1 (N6471, N6467);
and AND2 (N6472, N6466, N29);
and AND3 (N6473, N6458, N1385, N3347);
or OR3 (N6474, N6469, N3000, N1495);
nand NAND4 (N6475, N6465, N1687, N2904, N172);
or OR4 (N6476, N6468, N4016, N2246, N4668);
and AND3 (N6477, N6470, N5689, N5550);
not NOT1 (N6478, N6475);
not NOT1 (N6479, N6473);
buf BUF1 (N6480, N6474);
and AND3 (N6481, N6454, N4338, N829);
nor NOR2 (N6482, N6480, N4504);
buf BUF1 (N6483, N6471);
nor NOR3 (N6484, N6478, N5595, N2975);
xor XOR2 (N6485, N6479, N4495);
xor XOR2 (N6486, N6477, N5);
buf BUF1 (N6487, N6463);
buf BUF1 (N6488, N6484);
xor XOR2 (N6489, N6485, N6234);
buf BUF1 (N6490, N6487);
and AND4 (N6491, N6488, N3826, N444, N2531);
or OR2 (N6492, N6490, N851);
not NOT1 (N6493, N6472);
not NOT1 (N6494, N6493);
buf BUF1 (N6495, N6494);
not NOT1 (N6496, N6481);
buf BUF1 (N6497, N6483);
xor XOR2 (N6498, N6486, N4555);
nand NAND4 (N6499, N6489, N2911, N1860, N4919);
or OR3 (N6500, N6496, N805, N5200);
nand NAND2 (N6501, N6482, N5075);
buf BUF1 (N6502, N6497);
xor XOR2 (N6503, N6498, N3453);
nand NAND2 (N6504, N6501, N4529);
buf BUF1 (N6505, N6503);
not NOT1 (N6506, N6449);
nand NAND2 (N6507, N6504, N2660);
not NOT1 (N6508, N6507);
nor NOR2 (N6509, N6502, N4014);
not NOT1 (N6510, N6505);
nor NOR2 (N6511, N6492, N3045);
not NOT1 (N6512, N6500);
xor XOR2 (N6513, N6476, N5466);
or OR3 (N6514, N6510, N6047, N5177);
xor XOR2 (N6515, N6512, N5855);
xor XOR2 (N6516, N6495, N3441);
or OR3 (N6517, N6515, N2388, N5732);
or OR2 (N6518, N6511, N1946);
nand NAND4 (N6519, N6508, N5272, N6472, N4805);
nand NAND4 (N6520, N6506, N1888, N3611, N5566);
xor XOR2 (N6521, N6516, N2997);
not NOT1 (N6522, N6499);
or OR4 (N6523, N6521, N1404, N1944, N459);
buf BUF1 (N6524, N6517);
nor NOR4 (N6525, N6513, N2759, N4897, N320);
nor NOR2 (N6526, N6491, N4519);
xor XOR2 (N6527, N6526, N4093);
xor XOR2 (N6528, N6527, N2698);
not NOT1 (N6529, N6525);
not NOT1 (N6530, N6524);
nor NOR2 (N6531, N6519, N2525);
or OR3 (N6532, N6523, N869, N640);
and AND4 (N6533, N6520, N1856, N3124, N5174);
nand NAND4 (N6534, N6514, N3068, N655, N40);
and AND3 (N6535, N6518, N5578, N5373);
not NOT1 (N6536, N6531);
or OR3 (N6537, N6509, N2865, N3661);
buf BUF1 (N6538, N6533);
not NOT1 (N6539, N6528);
not NOT1 (N6540, N6538);
or OR4 (N6541, N6539, N4461, N865, N1171);
buf BUF1 (N6542, N6540);
or OR3 (N6543, N6537, N6531, N3061);
nor NOR4 (N6544, N6543, N3679, N5064, N1305);
nor NOR2 (N6545, N6532, N663);
nor NOR2 (N6546, N6542, N5787);
nor NOR2 (N6547, N6535, N6365);
and AND2 (N6548, N6536, N1834);
or OR2 (N6549, N6548, N3740);
nand NAND2 (N6550, N6529, N738);
not NOT1 (N6551, N6522);
or OR2 (N6552, N6549, N2655);
or OR2 (N6553, N6547, N6162);
nor NOR4 (N6554, N6541, N1568, N4775, N5523);
nand NAND4 (N6555, N6534, N533, N3961, N5967);
nand NAND3 (N6556, N6554, N5377, N632);
xor XOR2 (N6557, N6545, N1789);
nor NOR4 (N6558, N6557, N5859, N5089, N5756);
nand NAND2 (N6559, N6551, N1064);
xor XOR2 (N6560, N6544, N2969);
and AND2 (N6561, N6553, N2012);
xor XOR2 (N6562, N6560, N5382);
not NOT1 (N6563, N6556);
not NOT1 (N6564, N6559);
or OR3 (N6565, N6562, N2677, N4793);
not NOT1 (N6566, N6555);
nor NOR2 (N6567, N6565, N4324);
or OR4 (N6568, N6566, N3473, N204, N5271);
and AND4 (N6569, N6561, N4948, N4321, N2990);
nand NAND4 (N6570, N6550, N5126, N1116, N2277);
not NOT1 (N6571, N6564);
or OR4 (N6572, N6570, N295, N1031, N1181);
or OR2 (N6573, N6567, N4032);
nand NAND3 (N6574, N6569, N2387, N522);
xor XOR2 (N6575, N6574, N1200);
or OR4 (N6576, N6563, N432, N3821, N4119);
nor NOR4 (N6577, N6552, N6498, N1915, N4154);
buf BUF1 (N6578, N6546);
xor XOR2 (N6579, N6558, N5604);
xor XOR2 (N6580, N6573, N4316);
xor XOR2 (N6581, N6578, N200);
buf BUF1 (N6582, N6530);
nor NOR2 (N6583, N6582, N4383);
nand NAND3 (N6584, N6577, N3494, N3385);
nand NAND3 (N6585, N6568, N49, N1120);
or OR4 (N6586, N6584, N5097, N2770, N2975);
or OR4 (N6587, N6575, N530, N1889, N3185);
buf BUF1 (N6588, N6579);
nor NOR4 (N6589, N6583, N2015, N978, N5494);
or OR4 (N6590, N6585, N1209, N415, N4143);
or OR2 (N6591, N6590, N4802);
and AND2 (N6592, N6587, N5609);
nand NAND4 (N6593, N6589, N26, N5239, N566);
buf BUF1 (N6594, N6576);
or OR3 (N6595, N6581, N3071, N3950);
not NOT1 (N6596, N6571);
buf BUF1 (N6597, N6572);
nor NOR4 (N6598, N6586, N4458, N4288, N4355);
or OR3 (N6599, N6593, N1758, N188);
buf BUF1 (N6600, N6592);
not NOT1 (N6601, N6599);
buf BUF1 (N6602, N6594);
or OR3 (N6603, N6598, N6300, N3471);
and AND4 (N6604, N6602, N5817, N5249, N922);
not NOT1 (N6605, N6597);
and AND4 (N6606, N6605, N822, N3816, N434);
or OR4 (N6607, N6603, N2916, N5392, N6251);
nor NOR4 (N6608, N6607, N4285, N4853, N1549);
nand NAND3 (N6609, N6595, N3017, N6361);
buf BUF1 (N6610, N6596);
nor NOR4 (N6611, N6609, N6336, N2533, N6542);
nor NOR3 (N6612, N6604, N2578, N4860);
and AND4 (N6613, N6591, N6379, N5957, N1367);
nor NOR2 (N6614, N6606, N2019);
or OR2 (N6615, N6613, N1688);
nor NOR4 (N6616, N6588, N5548, N4062, N3381);
or OR4 (N6617, N6608, N2862, N5074, N6380);
or OR4 (N6618, N6600, N1012, N1950, N1553);
xor XOR2 (N6619, N6580, N114);
nor NOR3 (N6620, N6601, N896, N1413);
and AND3 (N6621, N6618, N785, N616);
xor XOR2 (N6622, N6616, N2171);
nand NAND4 (N6623, N6620, N4550, N385, N2715);
and AND2 (N6624, N6614, N2987);
buf BUF1 (N6625, N6617);
nor NOR3 (N6626, N6612, N806, N6580);
and AND3 (N6627, N6621, N5725, N5938);
and AND3 (N6628, N6622, N215, N4722);
xor XOR2 (N6629, N6610, N1830);
xor XOR2 (N6630, N6624, N4284);
or OR4 (N6631, N6623, N1770, N6282, N4118);
not NOT1 (N6632, N6627);
xor XOR2 (N6633, N6629, N6608);
and AND2 (N6634, N6625, N4291);
not NOT1 (N6635, N6633);
buf BUF1 (N6636, N6611);
nand NAND2 (N6637, N6632, N5757);
not NOT1 (N6638, N6615);
buf BUF1 (N6639, N6631);
or OR2 (N6640, N6619, N524);
nor NOR3 (N6641, N6639, N2840, N2256);
and AND4 (N6642, N6635, N5521, N206, N888);
buf BUF1 (N6643, N6641);
nor NOR3 (N6644, N6634, N252, N2071);
nand NAND3 (N6645, N6638, N5002, N340);
xor XOR2 (N6646, N6637, N887);
or OR2 (N6647, N6643, N2285);
not NOT1 (N6648, N6630);
buf BUF1 (N6649, N6648);
buf BUF1 (N6650, N6628);
or OR3 (N6651, N6646, N5037, N6406);
or OR2 (N6652, N6651, N579);
buf BUF1 (N6653, N6649);
nand NAND3 (N6654, N6645, N4362, N4382);
buf BUF1 (N6655, N6652);
buf BUF1 (N6656, N6654);
nor NOR3 (N6657, N6636, N2170, N680);
or OR2 (N6658, N6650, N5601);
and AND4 (N6659, N6642, N2044, N1393, N3069);
xor XOR2 (N6660, N6656, N868);
or OR3 (N6661, N6647, N283, N3046);
nor NOR3 (N6662, N6657, N4975, N460);
buf BUF1 (N6663, N6662);
not NOT1 (N6664, N6644);
buf BUF1 (N6665, N6655);
and AND2 (N6666, N6659, N3844);
or OR2 (N6667, N6663, N848);
not NOT1 (N6668, N6665);
and AND2 (N6669, N6661, N2394);
not NOT1 (N6670, N6669);
not NOT1 (N6671, N6658);
nand NAND2 (N6672, N6671, N1665);
nand NAND4 (N6673, N6672, N3000, N5895, N3504);
buf BUF1 (N6674, N6668);
and AND2 (N6675, N6674, N3834);
and AND3 (N6676, N6670, N2182, N6651);
buf BUF1 (N6677, N6667);
buf BUF1 (N6678, N6675);
or OR4 (N6679, N6677, N2402, N5938, N4883);
not NOT1 (N6680, N6666);
nor NOR4 (N6681, N6679, N4758, N2470, N2917);
nor NOR3 (N6682, N6681, N6105, N3580);
and AND3 (N6683, N6673, N2994, N5920);
nor NOR2 (N6684, N6680, N234);
xor XOR2 (N6685, N6664, N4813);
and AND3 (N6686, N6684, N2434, N729);
nor NOR2 (N6687, N6660, N3067);
nor NOR3 (N6688, N6676, N870, N5139);
buf BUF1 (N6689, N6678);
buf BUF1 (N6690, N6685);
not NOT1 (N6691, N6690);
not NOT1 (N6692, N6683);
nand NAND4 (N6693, N6687, N2308, N6486, N4784);
and AND2 (N6694, N6691, N457);
and AND4 (N6695, N6686, N1914, N2464, N4972);
buf BUF1 (N6696, N6640);
nand NAND4 (N6697, N6693, N2277, N41, N4068);
nand NAND4 (N6698, N6626, N6350, N2878, N3426);
buf BUF1 (N6699, N6698);
buf BUF1 (N6700, N6688);
not NOT1 (N6701, N6696);
nand NAND3 (N6702, N6699, N73, N4340);
buf BUF1 (N6703, N6697);
and AND4 (N6704, N6695, N2460, N4986, N1623);
not NOT1 (N6705, N6692);
buf BUF1 (N6706, N6700);
or OR4 (N6707, N6706, N4522, N2064, N1837);
nor NOR2 (N6708, N6705, N2702);
and AND3 (N6709, N6694, N3539, N767);
buf BUF1 (N6710, N6701);
xor XOR2 (N6711, N6707, N3972);
nor NOR3 (N6712, N6689, N3849, N1133);
nand NAND3 (N6713, N6711, N5907, N4457);
not NOT1 (N6714, N6682);
buf BUF1 (N6715, N6702);
and AND2 (N6716, N6653, N4854);
buf BUF1 (N6717, N6715);
not NOT1 (N6718, N6713);
not NOT1 (N6719, N6718);
not NOT1 (N6720, N6714);
not NOT1 (N6721, N6709);
nor NOR3 (N6722, N6719, N789, N2992);
or OR4 (N6723, N6720, N225, N2455, N518);
or OR2 (N6724, N6710, N452);
or OR3 (N6725, N6722, N5935, N3459);
buf BUF1 (N6726, N6725);
buf BUF1 (N6727, N6724);
nor NOR2 (N6728, N6726, N6613);
xor XOR2 (N6729, N6716, N1782);
nand NAND3 (N6730, N6717, N738, N2324);
not NOT1 (N6731, N6708);
buf BUF1 (N6732, N6703);
not NOT1 (N6733, N6732);
buf BUF1 (N6734, N6704);
nand NAND4 (N6735, N6730, N1652, N2393, N4289);
nor NOR2 (N6736, N6721, N4925);
and AND4 (N6737, N6723, N5694, N4804, N3512);
and AND4 (N6738, N6735, N4175, N3691, N3560);
not NOT1 (N6739, N6712);
not NOT1 (N6740, N6733);
nand NAND3 (N6741, N6739, N4768, N6328);
nand NAND4 (N6742, N6731, N1903, N1166, N1344);
or OR2 (N6743, N6734, N5049);
buf BUF1 (N6744, N6741);
xor XOR2 (N6745, N6744, N1961);
and AND3 (N6746, N6738, N5115, N506);
xor XOR2 (N6747, N6745, N6510);
and AND3 (N6748, N6740, N9, N482);
nand NAND2 (N6749, N6737, N1554);
xor XOR2 (N6750, N6728, N3652);
and AND4 (N6751, N6736, N2802, N2924, N4029);
nand NAND3 (N6752, N6747, N6104, N4639);
nand NAND4 (N6753, N6743, N3649, N5041, N5557);
nor NOR4 (N6754, N6753, N1829, N5048, N5516);
nor NOR3 (N6755, N6751, N4387, N3637);
xor XOR2 (N6756, N6749, N564);
xor XOR2 (N6757, N6748, N4950);
and AND4 (N6758, N6746, N3808, N4905, N1423);
buf BUF1 (N6759, N6727);
not NOT1 (N6760, N6752);
and AND4 (N6761, N6759, N6423, N4920, N6152);
xor XOR2 (N6762, N6750, N1423);
nand NAND4 (N6763, N6761, N6164, N4848, N991);
nand NAND2 (N6764, N6763, N586);
xor XOR2 (N6765, N6762, N410);
nand NAND2 (N6766, N6758, N318);
nand NAND4 (N6767, N6765, N6488, N3757, N6055);
and AND3 (N6768, N6764, N5479, N4707);
and AND3 (N6769, N6742, N3783, N1290);
or OR2 (N6770, N6760, N3254);
and AND2 (N6771, N6729, N1210);
not NOT1 (N6772, N6757);
nor NOR2 (N6773, N6766, N3518);
xor XOR2 (N6774, N6771, N123);
nor NOR3 (N6775, N6772, N22, N6055);
xor XOR2 (N6776, N6756, N2800);
xor XOR2 (N6777, N6768, N3413);
not NOT1 (N6778, N6755);
not NOT1 (N6779, N6778);
or OR3 (N6780, N6775, N2418, N1048);
nand NAND2 (N6781, N6777, N572);
or OR4 (N6782, N6754, N1274, N6014, N1538);
or OR2 (N6783, N6780, N2851);
or OR4 (N6784, N6770, N4351, N650, N4654);
and AND4 (N6785, N6779, N4855, N5631, N2805);
or OR4 (N6786, N6782, N3037, N4865, N2128);
nand NAND2 (N6787, N6767, N2833);
nor NOR2 (N6788, N6769, N5779);
nor NOR2 (N6789, N6776, N3729);
nand NAND3 (N6790, N6781, N6281, N4094);
not NOT1 (N6791, N6787);
not NOT1 (N6792, N6773);
xor XOR2 (N6793, N6785, N3857);
nor NOR3 (N6794, N6788, N5880, N1268);
and AND2 (N6795, N6789, N922);
buf BUF1 (N6796, N6783);
not NOT1 (N6797, N6784);
and AND2 (N6798, N6786, N2929);
or OR4 (N6799, N6791, N3487, N2506, N1862);
or OR4 (N6800, N6798, N3010, N2834, N6225);
and AND4 (N6801, N6797, N1337, N5991, N3612);
not NOT1 (N6802, N6796);
nor NOR3 (N6803, N6774, N2934, N6025);
xor XOR2 (N6804, N6800, N2185);
and AND3 (N6805, N6803, N3600, N1237);
and AND2 (N6806, N6802, N2444);
buf BUF1 (N6807, N6795);
not NOT1 (N6808, N6806);
and AND2 (N6809, N6793, N3230);
not NOT1 (N6810, N6790);
xor XOR2 (N6811, N6809, N781);
or OR3 (N6812, N6808, N4762, N134);
nor NOR4 (N6813, N6805, N3162, N2894, N3766);
or OR3 (N6814, N6804, N906, N2791);
nor NOR4 (N6815, N6812, N2121, N2890, N5508);
buf BUF1 (N6816, N6813);
buf BUF1 (N6817, N6816);
nand NAND2 (N6818, N6817, N2547);
and AND4 (N6819, N6814, N3833, N6668, N3279);
nor NOR4 (N6820, N6799, N5405, N6124, N6144);
or OR3 (N6821, N6819, N2799, N551);
and AND4 (N6822, N6807, N6679, N709, N2348);
buf BUF1 (N6823, N6801);
xor XOR2 (N6824, N6822, N3049);
or OR2 (N6825, N6811, N5703);
not NOT1 (N6826, N6823);
nor NOR3 (N6827, N6820, N3062, N462);
and AND3 (N6828, N6815, N5794, N6404);
nor NOR4 (N6829, N6810, N5468, N4777, N1465);
nor NOR4 (N6830, N6821, N2161, N2841, N5353);
nor NOR2 (N6831, N6792, N1745);
and AND4 (N6832, N6824, N1833, N4909, N4395);
or OR4 (N6833, N6830, N951, N6074, N2965);
buf BUF1 (N6834, N6833);
and AND4 (N6835, N6834, N1974, N426, N4603);
nor NOR3 (N6836, N6832, N3633, N1257);
and AND4 (N6837, N6835, N820, N835, N1466);
not NOT1 (N6838, N6794);
nand NAND2 (N6839, N6829, N4388);
buf BUF1 (N6840, N6818);
nand NAND3 (N6841, N6828, N1816, N4753);
buf BUF1 (N6842, N6836);
nor NOR4 (N6843, N6840, N6358, N2596, N4815);
nor NOR4 (N6844, N6839, N1909, N6789, N5839);
not NOT1 (N6845, N6843);
nor NOR3 (N6846, N6826, N4629, N5854);
nand NAND2 (N6847, N6846, N2859);
nor NOR4 (N6848, N6842, N1917, N2402, N4324);
nand NAND2 (N6849, N6838, N3025);
and AND3 (N6850, N6848, N3015, N4315);
nor NOR2 (N6851, N6845, N4584);
or OR3 (N6852, N6827, N6068, N3142);
or OR2 (N6853, N6841, N3570);
not NOT1 (N6854, N6849);
and AND4 (N6855, N6844, N455, N3447, N546);
nand NAND2 (N6856, N6850, N2356);
nand NAND4 (N6857, N6851, N1881, N1621, N5867);
buf BUF1 (N6858, N6847);
nand NAND2 (N6859, N6858, N5505);
and AND2 (N6860, N6856, N1710);
buf BUF1 (N6861, N6857);
buf BUF1 (N6862, N6855);
not NOT1 (N6863, N6859);
nor NOR2 (N6864, N6852, N5503);
and AND2 (N6865, N6837, N5524);
or OR3 (N6866, N6864, N5047, N1986);
xor XOR2 (N6867, N6865, N5244);
and AND2 (N6868, N6862, N1783);
xor XOR2 (N6869, N6868, N3189);
or OR3 (N6870, N6867, N2270, N1190);
nor NOR3 (N6871, N6870, N2113, N5729);
or OR2 (N6872, N6866, N5344);
and AND3 (N6873, N6825, N658, N5060);
xor XOR2 (N6874, N6869, N6430);
nand NAND3 (N6875, N6853, N5952, N3040);
nor NOR2 (N6876, N6863, N5013);
nand NAND4 (N6877, N6861, N377, N5821, N2141);
and AND2 (N6878, N6877, N712);
buf BUF1 (N6879, N6871);
nor NOR4 (N6880, N6878, N2139, N704, N1248);
nand NAND3 (N6881, N6875, N350, N6114);
or OR3 (N6882, N6880, N6410, N2011);
nor NOR3 (N6883, N6873, N815, N6441);
xor XOR2 (N6884, N6881, N70);
nor NOR3 (N6885, N6854, N2238, N747);
nand NAND4 (N6886, N6885, N2145, N1596, N4151);
nor NOR3 (N6887, N6872, N1628, N4052);
and AND3 (N6888, N6883, N6750, N4918);
nor NOR4 (N6889, N6888, N4585, N5417, N2114);
and AND2 (N6890, N6874, N2140);
and AND4 (N6891, N6876, N530, N4568, N3602);
buf BUF1 (N6892, N6891);
nand NAND3 (N6893, N6879, N6710, N5465);
and AND2 (N6894, N6884, N2989);
buf BUF1 (N6895, N6886);
nand NAND2 (N6896, N6831, N5195);
or OR3 (N6897, N6889, N6345, N2284);
or OR4 (N6898, N6882, N2600, N5991, N5547);
xor XOR2 (N6899, N6892, N5707);
and AND4 (N6900, N6896, N2637, N723, N3044);
or OR3 (N6901, N6898, N1607, N1815);
and AND4 (N6902, N6900, N6507, N1218, N6690);
buf BUF1 (N6903, N6899);
buf BUF1 (N6904, N6887);
nand NAND2 (N6905, N6904, N1799);
nor NOR2 (N6906, N6905, N806);
nor NOR2 (N6907, N6893, N4197);
or OR2 (N6908, N6860, N1555);
xor XOR2 (N6909, N6906, N5038);
or OR4 (N6910, N6895, N6347, N3184, N995);
not NOT1 (N6911, N6901);
or OR4 (N6912, N6909, N3840, N6499, N4707);
nand NAND4 (N6913, N6894, N5263, N1820, N3991);
or OR3 (N6914, N6908, N6205, N3865);
and AND2 (N6915, N6897, N5803);
nand NAND4 (N6916, N6902, N142, N5537, N3690);
xor XOR2 (N6917, N6914, N4978);
not NOT1 (N6918, N6915);
or OR4 (N6919, N6890, N2151, N4480, N1806);
and AND2 (N6920, N6910, N3893);
and AND2 (N6921, N6911, N439);
nor NOR4 (N6922, N6916, N1444, N4806, N2591);
xor XOR2 (N6923, N6921, N749);
or OR2 (N6924, N6903, N501);
nand NAND3 (N6925, N6923, N4971, N4260);
or OR3 (N6926, N6918, N5022, N5821);
not NOT1 (N6927, N6912);
nand NAND4 (N6928, N6922, N4366, N6712, N3726);
nand NAND4 (N6929, N6928, N3011, N3878, N5795);
and AND3 (N6930, N6920, N5486, N5951);
or OR4 (N6931, N6927, N791, N45, N6474);
nor NOR2 (N6932, N6913, N4655);
not NOT1 (N6933, N6917);
and AND2 (N6934, N6932, N411);
nor NOR2 (N6935, N6933, N5407);
and AND3 (N6936, N6907, N2313, N1469);
buf BUF1 (N6937, N6936);
not NOT1 (N6938, N6931);
not NOT1 (N6939, N6935);
not NOT1 (N6940, N6938);
nor NOR2 (N6941, N6934, N1298);
buf BUF1 (N6942, N6926);
xor XOR2 (N6943, N6930, N328);
nand NAND3 (N6944, N6924, N6756, N5270);
xor XOR2 (N6945, N6944, N4702);
nand NAND2 (N6946, N6937, N4438);
nor NOR4 (N6947, N6929, N6773, N5271, N2561);
buf BUF1 (N6948, N6940);
and AND2 (N6949, N6941, N1839);
nor NOR3 (N6950, N6925, N2161, N1768);
buf BUF1 (N6951, N6947);
and AND2 (N6952, N6943, N5487);
not NOT1 (N6953, N6948);
nor NOR2 (N6954, N6952, N3103);
buf BUF1 (N6955, N6953);
or OR2 (N6956, N6919, N6567);
and AND3 (N6957, N6955, N1803, N1162);
not NOT1 (N6958, N6956);
nand NAND2 (N6959, N6939, N1002);
buf BUF1 (N6960, N6949);
buf BUF1 (N6961, N6958);
not NOT1 (N6962, N6951);
nor NOR4 (N6963, N6950, N2044, N6747, N5061);
nor NOR3 (N6964, N6946, N1877, N371);
not NOT1 (N6965, N6942);
not NOT1 (N6966, N6957);
nand NAND4 (N6967, N6964, N4161, N6113, N5822);
and AND4 (N6968, N6945, N5059, N3751, N2191);
xor XOR2 (N6969, N6967, N6579);
and AND3 (N6970, N6965, N1806, N2102);
buf BUF1 (N6971, N6954);
not NOT1 (N6972, N6970);
nor NOR2 (N6973, N6959, N3630);
not NOT1 (N6974, N6972);
buf BUF1 (N6975, N6974);
nand NAND3 (N6976, N6971, N733, N876);
buf BUF1 (N6977, N6973);
buf BUF1 (N6978, N6977);
nand NAND3 (N6979, N6961, N5203, N335);
or OR4 (N6980, N6978, N2247, N4250, N1784);
nand NAND2 (N6981, N6969, N3056);
not NOT1 (N6982, N6968);
buf BUF1 (N6983, N6982);
or OR2 (N6984, N6962, N4234);
or OR4 (N6985, N6984, N898, N3911, N6352);
nor NOR4 (N6986, N6960, N3277, N859, N232);
nor NOR4 (N6987, N6963, N2184, N1013, N1412);
and AND4 (N6988, N6986, N874, N5569, N1809);
nand NAND3 (N6989, N6985, N6656, N296);
and AND4 (N6990, N6976, N1534, N1668, N2076);
not NOT1 (N6991, N6990);
nor NOR4 (N6992, N6980, N1509, N6856, N3041);
or OR2 (N6993, N6981, N6558);
and AND2 (N6994, N6991, N2012);
nor NOR3 (N6995, N6975, N2602, N702);
and AND2 (N6996, N6995, N5887);
nor NOR4 (N6997, N6992, N855, N557, N4635);
buf BUF1 (N6998, N6994);
buf BUF1 (N6999, N6987);
nor NOR4 (N7000, N6979, N6506, N3119, N3492);
buf BUF1 (N7001, N6983);
nand NAND2 (N7002, N6996, N3275);
not NOT1 (N7003, N6997);
nor NOR2 (N7004, N6998, N5562);
and AND3 (N7005, N7003, N6080, N5916);
or OR3 (N7006, N6989, N189, N3085);
xor XOR2 (N7007, N6988, N1241);
and AND4 (N7008, N7005, N2354, N255, N5105);
nor NOR3 (N7009, N7008, N3004, N796);
and AND3 (N7010, N7009, N6521, N5550);
not NOT1 (N7011, N6966);
buf BUF1 (N7012, N7010);
nand NAND3 (N7013, N6993, N4172, N619);
buf BUF1 (N7014, N7013);
not NOT1 (N7015, N7014);
nand NAND4 (N7016, N7006, N6429, N2538, N4869);
and AND3 (N7017, N7001, N302, N1072);
nand NAND4 (N7018, N7011, N5733, N2581, N6063);
buf BUF1 (N7019, N7018);
or OR4 (N7020, N7016, N416, N4984, N1577);
nand NAND3 (N7021, N7017, N3311, N511);
and AND2 (N7022, N7019, N1614);
xor XOR2 (N7023, N7000, N6);
or OR2 (N7024, N7002, N3022);
nand NAND3 (N7025, N7012, N3469, N2373);
xor XOR2 (N7026, N7024, N1266);
and AND2 (N7027, N7021, N1069);
buf BUF1 (N7028, N7025);
xor XOR2 (N7029, N7007, N6417);
not NOT1 (N7030, N7027);
or OR2 (N7031, N7029, N2759);
nand NAND2 (N7032, N7028, N211);
buf BUF1 (N7033, N7032);
buf BUF1 (N7034, N6999);
xor XOR2 (N7035, N7033, N5762);
xor XOR2 (N7036, N7015, N166);
or OR3 (N7037, N7034, N3841, N1180);
and AND2 (N7038, N7023, N6216);
or OR3 (N7039, N7020, N1841, N866);
xor XOR2 (N7040, N7031, N5469);
or OR3 (N7041, N7030, N3415, N6253);
xor XOR2 (N7042, N7039, N571);
xor XOR2 (N7043, N7040, N6395);
buf BUF1 (N7044, N7037);
nand NAND4 (N7045, N7035, N6072, N3719, N2329);
nor NOR3 (N7046, N7038, N964, N2029);
nand NAND4 (N7047, N7036, N6987, N2734, N4193);
nor NOR4 (N7048, N7026, N4331, N3230, N4222);
or OR2 (N7049, N7043, N5999);
and AND4 (N7050, N7044, N632, N2777, N3978);
buf BUF1 (N7051, N7041);
xor XOR2 (N7052, N7051, N3018);
buf BUF1 (N7053, N7022);
xor XOR2 (N7054, N7052, N3728);
xor XOR2 (N7055, N7049, N365);
xor XOR2 (N7056, N7054, N4830);
not NOT1 (N7057, N7004);
and AND4 (N7058, N7055, N4148, N885, N5253);
nand NAND3 (N7059, N7053, N2059, N6720);
nand NAND4 (N7060, N7057, N5278, N1942, N3798);
buf BUF1 (N7061, N7050);
not NOT1 (N7062, N7045);
or OR3 (N7063, N7062, N2578, N5503);
xor XOR2 (N7064, N7061, N1545);
xor XOR2 (N7065, N7042, N3828);
and AND2 (N7066, N7064, N5213);
and AND4 (N7067, N7065, N2204, N2249, N6370);
and AND2 (N7068, N7060, N3388);
nor NOR2 (N7069, N7067, N2452);
xor XOR2 (N7070, N7047, N3105);
buf BUF1 (N7071, N7070);
nor NOR2 (N7072, N7056, N5307);
xor XOR2 (N7073, N7058, N4256);
buf BUF1 (N7074, N7059);
xor XOR2 (N7075, N7073, N421);
or OR2 (N7076, N7071, N3860);
xor XOR2 (N7077, N7048, N5977);
not NOT1 (N7078, N7063);
and AND2 (N7079, N7069, N887);
nand NAND2 (N7080, N7076, N1780);
buf BUF1 (N7081, N7072);
buf BUF1 (N7082, N7078);
and AND4 (N7083, N7046, N2545, N6385, N2001);
not NOT1 (N7084, N7068);
nand NAND3 (N7085, N7079, N2847, N3074);
nand NAND3 (N7086, N7085, N564, N1105);
buf BUF1 (N7087, N7074);
nand NAND2 (N7088, N7075, N6491);
xor XOR2 (N7089, N7084, N3018);
and AND3 (N7090, N7082, N257, N3708);
and AND4 (N7091, N7090, N4451, N3260, N2902);
not NOT1 (N7092, N7088);
nor NOR2 (N7093, N7066, N393);
not NOT1 (N7094, N7091);
buf BUF1 (N7095, N7089);
nand NAND2 (N7096, N7093, N3448);
or OR3 (N7097, N7087, N1502, N6849);
or OR2 (N7098, N7095, N2310);
not NOT1 (N7099, N7083);
xor XOR2 (N7100, N7092, N152);
buf BUF1 (N7101, N7080);
nand NAND3 (N7102, N7100, N6850, N3573);
and AND3 (N7103, N7096, N374, N3977);
buf BUF1 (N7104, N7086);
nor NOR4 (N7105, N7101, N1312, N4699, N4872);
or OR2 (N7106, N7104, N4009);
nand NAND3 (N7107, N7106, N1868, N2475);
nand NAND4 (N7108, N7105, N1031, N1017, N6926);
and AND2 (N7109, N7099, N6628);
nor NOR4 (N7110, N7103, N5064, N6682, N1296);
nand NAND2 (N7111, N7109, N6446);
or OR4 (N7112, N7081, N3823, N7082, N2802);
xor XOR2 (N7113, N7108, N6521);
nor NOR2 (N7114, N7094, N812);
xor XOR2 (N7115, N7102, N6478);
xor XOR2 (N7116, N7112, N130);
nor NOR3 (N7117, N7098, N4053, N2762);
nor NOR4 (N7118, N7115, N1685, N5061, N4203);
nand NAND2 (N7119, N7118, N3913);
and AND2 (N7120, N7077, N182);
or OR4 (N7121, N7120, N5122, N863, N2697);
not NOT1 (N7122, N7113);
xor XOR2 (N7123, N7122, N6071);
nand NAND3 (N7124, N7111, N6489, N6473);
and AND2 (N7125, N7123, N1972);
nor NOR4 (N7126, N7097, N5173, N6787, N715);
nand NAND4 (N7127, N7110, N3417, N4648, N4684);
xor XOR2 (N7128, N7124, N6241);
nand NAND3 (N7129, N7125, N6430, N3483);
buf BUF1 (N7130, N7126);
buf BUF1 (N7131, N7116);
buf BUF1 (N7132, N7129);
and AND2 (N7133, N7128, N2896);
buf BUF1 (N7134, N7127);
nor NOR4 (N7135, N7133, N1191, N2272, N4955);
nand NAND2 (N7136, N7134, N5421);
nand NAND4 (N7137, N7117, N5878, N1250, N1873);
nand NAND4 (N7138, N7136, N2728, N2319, N5124);
not NOT1 (N7139, N7131);
or OR4 (N7140, N7139, N4962, N218, N3392);
or OR3 (N7141, N7138, N1547, N4938);
or OR2 (N7142, N7135, N4583);
not NOT1 (N7143, N7140);
and AND2 (N7144, N7114, N2567);
or OR3 (N7145, N7143, N7122, N4014);
nand NAND3 (N7146, N7141, N5740, N3157);
nand NAND2 (N7147, N7121, N5524);
and AND2 (N7148, N7145, N1894);
and AND4 (N7149, N7132, N5637, N1312, N4391);
nand NAND4 (N7150, N7144, N4651, N5348, N1101);
not NOT1 (N7151, N7107);
or OR2 (N7152, N7119, N5057);
nor NOR2 (N7153, N7152, N118);
xor XOR2 (N7154, N7151, N977);
nor NOR3 (N7155, N7148, N2396, N7006);
and AND3 (N7156, N7137, N5782, N1385);
nor NOR2 (N7157, N7150, N550);
or OR3 (N7158, N7153, N2660, N1563);
or OR4 (N7159, N7156, N1719, N5229, N1731);
nand NAND2 (N7160, N7155, N3826);
xor XOR2 (N7161, N7158, N3993);
nor NOR4 (N7162, N7157, N5354, N3745, N721);
buf BUF1 (N7163, N7130);
and AND4 (N7164, N7159, N6084, N2140, N2084);
and AND2 (N7165, N7163, N5725);
and AND4 (N7166, N7164, N5040, N260, N6597);
and AND3 (N7167, N7149, N300, N857);
buf BUF1 (N7168, N7165);
nor NOR2 (N7169, N7147, N2401);
or OR2 (N7170, N7167, N5623);
and AND4 (N7171, N7162, N2591, N3018, N937);
nor NOR4 (N7172, N7146, N851, N6579, N5253);
and AND2 (N7173, N7168, N3170);
nand NAND2 (N7174, N7173, N2409);
or OR3 (N7175, N7161, N4161, N4942);
and AND4 (N7176, N7154, N1789, N2750, N3994);
or OR4 (N7177, N7175, N5536, N3080, N4611);
nand NAND4 (N7178, N7177, N6498, N1447, N5211);
xor XOR2 (N7179, N7171, N1027);
buf BUF1 (N7180, N7160);
buf BUF1 (N7181, N7172);
buf BUF1 (N7182, N7176);
nand NAND2 (N7183, N7179, N963);
buf BUF1 (N7184, N7142);
or OR3 (N7185, N7174, N4772, N4309);
not NOT1 (N7186, N7169);
or OR3 (N7187, N7186, N208, N4372);
not NOT1 (N7188, N7187);
nor NOR3 (N7189, N7184, N4435, N2194);
and AND3 (N7190, N7188, N713, N6977);
buf BUF1 (N7191, N7189);
or OR4 (N7192, N7183, N2859, N4362, N6717);
xor XOR2 (N7193, N7178, N1635);
nand NAND2 (N7194, N7180, N4659);
buf BUF1 (N7195, N7193);
nor NOR4 (N7196, N7182, N3164, N2325, N4888);
xor XOR2 (N7197, N7196, N312);
not NOT1 (N7198, N7170);
nand NAND4 (N7199, N7195, N1294, N6098, N5360);
nand NAND2 (N7200, N7199, N3485);
and AND4 (N7201, N7191, N775, N1156, N6346);
xor XOR2 (N7202, N7185, N1805);
buf BUF1 (N7203, N7201);
and AND2 (N7204, N7200, N3192);
nand NAND2 (N7205, N7204, N5034);
nor NOR4 (N7206, N7205, N3268, N3506, N1212);
nand NAND3 (N7207, N7198, N1685, N1986);
buf BUF1 (N7208, N7192);
and AND4 (N7209, N7202, N2926, N6027, N6798);
buf BUF1 (N7210, N7166);
xor XOR2 (N7211, N7207, N148);
or OR2 (N7212, N7190, N4996);
and AND2 (N7213, N7208, N3486);
nand NAND2 (N7214, N7209, N5455);
nor NOR4 (N7215, N7212, N1780, N4254, N4808);
nor NOR4 (N7216, N7210, N1772, N2392, N5276);
not NOT1 (N7217, N7194);
or OR3 (N7218, N7217, N860, N5193);
nor NOR3 (N7219, N7218, N5503, N3062);
not NOT1 (N7220, N7206);
and AND2 (N7221, N7213, N4276);
xor XOR2 (N7222, N7215, N3527);
buf BUF1 (N7223, N7211);
nor NOR4 (N7224, N7197, N5629, N3530, N86);
not NOT1 (N7225, N7223);
xor XOR2 (N7226, N7181, N109);
and AND2 (N7227, N7225, N1157);
xor XOR2 (N7228, N7220, N676);
nand NAND3 (N7229, N7227, N107, N715);
nand NAND2 (N7230, N7203, N6901);
or OR2 (N7231, N7230, N782);
and AND4 (N7232, N7221, N6796, N1284, N1870);
xor XOR2 (N7233, N7219, N4131);
nand NAND3 (N7234, N7216, N4413, N4027);
or OR3 (N7235, N7226, N6622, N3855);
nor NOR2 (N7236, N7233, N5619);
or OR2 (N7237, N7232, N4138);
nand NAND4 (N7238, N7231, N4983, N2470, N3311);
and AND4 (N7239, N7224, N1951, N5716, N2111);
nor NOR3 (N7240, N7236, N5586, N6596);
buf BUF1 (N7241, N7239);
xor XOR2 (N7242, N7229, N1241);
not NOT1 (N7243, N7235);
and AND4 (N7244, N7228, N3964, N5182, N2204);
or OR2 (N7245, N7243, N744);
nand NAND4 (N7246, N7238, N6939, N407, N6528);
buf BUF1 (N7247, N7214);
not NOT1 (N7248, N7237);
not NOT1 (N7249, N7222);
nand NAND4 (N7250, N7240, N6061, N5323, N4125);
xor XOR2 (N7251, N7249, N7040);
and AND3 (N7252, N7234, N4053, N1100);
xor XOR2 (N7253, N7245, N3360);
nor NOR3 (N7254, N7244, N6214, N2766);
not NOT1 (N7255, N7250);
buf BUF1 (N7256, N7252);
xor XOR2 (N7257, N7256, N3280);
xor XOR2 (N7258, N7254, N4970);
and AND3 (N7259, N7248, N5703, N3359);
nor NOR3 (N7260, N7242, N2490, N867);
not NOT1 (N7261, N7253);
nor NOR2 (N7262, N7246, N3547);
not NOT1 (N7263, N7251);
or OR3 (N7264, N7259, N6946, N6543);
and AND4 (N7265, N7247, N6770, N2428, N6416);
not NOT1 (N7266, N7257);
and AND3 (N7267, N7263, N3206, N7218);
nand NAND2 (N7268, N7265, N6024);
or OR3 (N7269, N7267, N3532, N6174);
nand NAND3 (N7270, N7262, N644, N6349);
nor NOR4 (N7271, N7255, N4444, N697, N5509);
and AND3 (N7272, N7264, N6599, N5246);
buf BUF1 (N7273, N7269);
not NOT1 (N7274, N7272);
not NOT1 (N7275, N7274);
and AND2 (N7276, N7268, N3468);
buf BUF1 (N7277, N7276);
and AND3 (N7278, N7277, N5013, N5965);
nor NOR2 (N7279, N7271, N3409);
buf BUF1 (N7280, N7241);
not NOT1 (N7281, N7280);
nor NOR4 (N7282, N7258, N817, N1144, N293);
not NOT1 (N7283, N7279);
not NOT1 (N7284, N7281);
and AND4 (N7285, N7275, N4896, N447, N2538);
not NOT1 (N7286, N7270);
buf BUF1 (N7287, N7260);
or OR4 (N7288, N7261, N6945, N1659, N3081);
buf BUF1 (N7289, N7282);
and AND4 (N7290, N7285, N749, N4313, N4956);
not NOT1 (N7291, N7287);
nor NOR2 (N7292, N7283, N6080);
or OR3 (N7293, N7291, N4214, N1318);
not NOT1 (N7294, N7289);
or OR2 (N7295, N7292, N1896);
nor NOR3 (N7296, N7288, N6137, N3840);
or OR4 (N7297, N7296, N601, N95, N3179);
xor XOR2 (N7298, N7294, N3847);
or OR4 (N7299, N7284, N2433, N4186, N3840);
buf BUF1 (N7300, N7293);
and AND3 (N7301, N7299, N5421, N5259);
not NOT1 (N7302, N7273);
xor XOR2 (N7303, N7295, N2910);
or OR2 (N7304, N7303, N1254);
and AND3 (N7305, N7298, N3470, N504);
or OR3 (N7306, N7290, N2957, N3368);
nand NAND4 (N7307, N7300, N3375, N1128, N2732);
or OR3 (N7308, N7304, N3398, N4718);
nor NOR3 (N7309, N7266, N6894, N5496);
nor NOR3 (N7310, N7297, N4431, N1109);
buf BUF1 (N7311, N7310);
nand NAND3 (N7312, N7309, N3157, N309);
buf BUF1 (N7313, N7305);
buf BUF1 (N7314, N7307);
buf BUF1 (N7315, N7314);
not NOT1 (N7316, N7278);
xor XOR2 (N7317, N7301, N3249);
nand NAND2 (N7318, N7286, N5982);
nor NOR3 (N7319, N7313, N2317, N2253);
or OR2 (N7320, N7306, N6200);
or OR3 (N7321, N7316, N5368, N6784);
nand NAND2 (N7322, N7302, N6534);
not NOT1 (N7323, N7322);
nor NOR2 (N7324, N7308, N2396);
xor XOR2 (N7325, N7323, N4938);
not NOT1 (N7326, N7312);
not NOT1 (N7327, N7324);
and AND2 (N7328, N7327, N4917);
xor XOR2 (N7329, N7326, N5772);
or OR3 (N7330, N7311, N489, N6975);
nand NAND2 (N7331, N7319, N3309);
xor XOR2 (N7332, N7315, N5813);
not NOT1 (N7333, N7329);
or OR4 (N7334, N7332, N1613, N6651, N3047);
buf BUF1 (N7335, N7334);
buf BUF1 (N7336, N7330);
nand NAND4 (N7337, N7325, N6638, N2223, N6672);
nor NOR2 (N7338, N7328, N2786);
xor XOR2 (N7339, N7335, N6669);
or OR3 (N7340, N7336, N1568, N4472);
xor XOR2 (N7341, N7317, N3415);
not NOT1 (N7342, N7337);
xor XOR2 (N7343, N7342, N2313);
xor XOR2 (N7344, N7331, N6805);
not NOT1 (N7345, N7318);
or OR3 (N7346, N7341, N7121, N4842);
buf BUF1 (N7347, N7338);
buf BUF1 (N7348, N7339);
nor NOR4 (N7349, N7340, N2774, N1279, N1590);
and AND2 (N7350, N7347, N5946);
nand NAND3 (N7351, N7321, N5554, N6891);
not NOT1 (N7352, N7343);
nand NAND3 (N7353, N7345, N4467, N5158);
not NOT1 (N7354, N7349);
or OR4 (N7355, N7352, N6431, N4538, N6675);
nand NAND3 (N7356, N7354, N1529, N2826);
and AND4 (N7357, N7348, N4666, N3417, N5154);
and AND4 (N7358, N7351, N6242, N5368, N2210);
not NOT1 (N7359, N7353);
nand NAND2 (N7360, N7356, N1369);
or OR2 (N7361, N7360, N6701);
or OR2 (N7362, N7358, N420);
or OR3 (N7363, N7362, N418, N1181);
not NOT1 (N7364, N7357);
buf BUF1 (N7365, N7333);
buf BUF1 (N7366, N7361);
not NOT1 (N7367, N7355);
or OR3 (N7368, N7365, N1063, N3726);
nand NAND3 (N7369, N7363, N7295, N4786);
xor XOR2 (N7370, N7366, N5621);
not NOT1 (N7371, N7346);
nor NOR4 (N7372, N7344, N1320, N604, N5931);
and AND2 (N7373, N7368, N2264);
and AND3 (N7374, N7371, N2157, N5487);
xor XOR2 (N7375, N7350, N2780);
and AND2 (N7376, N7375, N1991);
and AND4 (N7377, N7359, N1745, N329, N2911);
buf BUF1 (N7378, N7370);
xor XOR2 (N7379, N7320, N7067);
xor XOR2 (N7380, N7374, N7357);
nor NOR3 (N7381, N7380, N1340, N1095);
xor XOR2 (N7382, N7376, N5427);
and AND3 (N7383, N7364, N4123, N809);
nor NOR4 (N7384, N7367, N4958, N6571, N1099);
or OR2 (N7385, N7369, N7282);
not NOT1 (N7386, N7381);
buf BUF1 (N7387, N7384);
and AND4 (N7388, N7382, N3497, N2199, N3481);
nor NOR3 (N7389, N7387, N4570, N1991);
and AND3 (N7390, N7386, N6080, N3312);
nand NAND2 (N7391, N7379, N2474);
xor XOR2 (N7392, N7390, N1149);
and AND3 (N7393, N7392, N3912, N228);
xor XOR2 (N7394, N7385, N6155);
and AND3 (N7395, N7393, N1835, N1502);
buf BUF1 (N7396, N7378);
and AND2 (N7397, N7389, N5579);
nand NAND3 (N7398, N7391, N4436, N299);
and AND4 (N7399, N7373, N4802, N2861, N385);
or OR2 (N7400, N7398, N4924);
xor XOR2 (N7401, N7400, N6254);
not NOT1 (N7402, N7399);
not NOT1 (N7403, N7394);
and AND3 (N7404, N7383, N1472, N481);
or OR3 (N7405, N7403, N5649, N5281);
buf BUF1 (N7406, N7396);
buf BUF1 (N7407, N7404);
or OR3 (N7408, N7377, N5603, N1156);
buf BUF1 (N7409, N7402);
buf BUF1 (N7410, N7372);
nand NAND4 (N7411, N7388, N7028, N3656, N6545);
and AND4 (N7412, N7410, N4056, N4507, N2128);
buf BUF1 (N7413, N7412);
not NOT1 (N7414, N7401);
not NOT1 (N7415, N7413);
nor NOR4 (N7416, N7411, N4530, N1550, N3109);
nor NOR2 (N7417, N7407, N4636);
buf BUF1 (N7418, N7406);
xor XOR2 (N7419, N7418, N3690);
not NOT1 (N7420, N7415);
xor XOR2 (N7421, N7416, N6179);
or OR2 (N7422, N7405, N5115);
buf BUF1 (N7423, N7422);
nor NOR2 (N7424, N7414, N5951);
buf BUF1 (N7425, N7424);
nor NOR3 (N7426, N7397, N7312, N98);
nor NOR4 (N7427, N7417, N3816, N6457, N7402);
and AND4 (N7428, N7427, N2301, N7384, N4992);
and AND4 (N7429, N7420, N3147, N383, N2020);
xor XOR2 (N7430, N7408, N758);
xor XOR2 (N7431, N7428, N2356);
nor NOR2 (N7432, N7430, N2778);
and AND3 (N7433, N7426, N3825, N1092);
nor NOR3 (N7434, N7409, N4562, N1881);
xor XOR2 (N7435, N7421, N1613);
xor XOR2 (N7436, N7431, N5184);
and AND2 (N7437, N7429, N3725);
nand NAND4 (N7438, N7434, N4263, N7215, N3714);
nor NOR3 (N7439, N7423, N6177, N5124);
not NOT1 (N7440, N7425);
and AND2 (N7441, N7438, N4030);
or OR3 (N7442, N7435, N6218, N480);
xor XOR2 (N7443, N7433, N3035);
buf BUF1 (N7444, N7441);
nor NOR2 (N7445, N7395, N5255);
buf BUF1 (N7446, N7436);
or OR2 (N7447, N7443, N5433);
nand NAND4 (N7448, N7446, N2056, N2202, N2377);
or OR2 (N7449, N7437, N7233);
nand NAND2 (N7450, N7439, N6035);
and AND3 (N7451, N7419, N30, N3299);
buf BUF1 (N7452, N7440);
xor XOR2 (N7453, N7448, N5060);
not NOT1 (N7454, N7450);
and AND3 (N7455, N7442, N7453, N4555);
and AND2 (N7456, N7131, N1675);
and AND2 (N7457, N7444, N6487);
buf BUF1 (N7458, N7455);
not NOT1 (N7459, N7447);
and AND2 (N7460, N7451, N378);
buf BUF1 (N7461, N7445);
nor NOR3 (N7462, N7458, N5007, N4772);
nand NAND3 (N7463, N7456, N6722, N6308);
and AND2 (N7464, N7449, N6772);
or OR4 (N7465, N7459, N5410, N4337, N6041);
or OR2 (N7466, N7462, N7388);
or OR4 (N7467, N7466, N2143, N4113, N4795);
nand NAND4 (N7468, N7452, N1005, N5699, N1646);
nand NAND2 (N7469, N7461, N2034);
and AND4 (N7470, N7432, N4087, N4885, N2602);
buf BUF1 (N7471, N7464);
buf BUF1 (N7472, N7465);
xor XOR2 (N7473, N7469, N5126);
nand NAND2 (N7474, N7457, N1834);
and AND4 (N7475, N7470, N1781, N5487, N6545);
xor XOR2 (N7476, N7467, N727);
and AND2 (N7477, N7472, N6384);
and AND4 (N7478, N7473, N845, N7126, N2880);
or OR2 (N7479, N7468, N2874);
xor XOR2 (N7480, N7454, N4392);
not NOT1 (N7481, N7477);
nand NAND2 (N7482, N7476, N2946);
or OR4 (N7483, N7481, N1867, N862, N7376);
or OR2 (N7484, N7480, N3241);
or OR3 (N7485, N7471, N1680, N4337);
nand NAND4 (N7486, N7474, N3184, N523, N6042);
nand NAND4 (N7487, N7460, N3754, N4948, N1848);
xor XOR2 (N7488, N7479, N1616);
nor NOR3 (N7489, N7482, N4123, N5882);
xor XOR2 (N7490, N7489, N4168);
and AND2 (N7491, N7490, N3020);
or OR3 (N7492, N7491, N5811, N1707);
xor XOR2 (N7493, N7484, N7425);
xor XOR2 (N7494, N7488, N1948);
nor NOR2 (N7495, N7483, N7487);
xor XOR2 (N7496, N6017, N2474);
not NOT1 (N7497, N7492);
or OR3 (N7498, N7494, N6415, N4666);
or OR3 (N7499, N7495, N136, N5406);
nand NAND4 (N7500, N7497, N3252, N7147, N7176);
nor NOR3 (N7501, N7496, N4612, N6283);
nand NAND3 (N7502, N7501, N7428, N1107);
not NOT1 (N7503, N7500);
buf BUF1 (N7504, N7502);
nor NOR2 (N7505, N7493, N5980);
or OR2 (N7506, N7499, N51);
not NOT1 (N7507, N7475);
or OR4 (N7508, N7506, N7189, N4827, N5378);
or OR2 (N7509, N7508, N63);
not NOT1 (N7510, N7507);
and AND2 (N7511, N7478, N4000);
xor XOR2 (N7512, N7485, N93);
or OR2 (N7513, N7512, N6783);
xor XOR2 (N7514, N7503, N885);
or OR3 (N7515, N7504, N3018, N3983);
nand NAND4 (N7516, N7515, N3301, N6575, N6582);
xor XOR2 (N7517, N7498, N6500);
and AND4 (N7518, N7513, N6373, N837, N844);
xor XOR2 (N7519, N7509, N4673);
nor NOR3 (N7520, N7518, N6474, N7031);
nor NOR2 (N7521, N7510, N2772);
buf BUF1 (N7522, N7517);
or OR4 (N7523, N7486, N407, N7024, N3860);
and AND4 (N7524, N7521, N4835, N6723, N3613);
not NOT1 (N7525, N7524);
nor NOR4 (N7526, N7523, N2711, N6750, N5283);
and AND2 (N7527, N7522, N5306);
xor XOR2 (N7528, N7505, N4149);
or OR4 (N7529, N7528, N6848, N3513, N5091);
or OR3 (N7530, N7516, N1377, N5667);
buf BUF1 (N7531, N7463);
nor NOR3 (N7532, N7530, N5671, N6044);
xor XOR2 (N7533, N7526, N6071);
not NOT1 (N7534, N7511);
xor XOR2 (N7535, N7514, N3004);
buf BUF1 (N7536, N7532);
and AND4 (N7537, N7529, N5159, N877, N6848);
xor XOR2 (N7538, N7533, N3935);
xor XOR2 (N7539, N7536, N1516);
buf BUF1 (N7540, N7539);
and AND2 (N7541, N7537, N1537);
and AND3 (N7542, N7519, N1461, N4664);
not NOT1 (N7543, N7542);
or OR4 (N7544, N7520, N2245, N3429, N5657);
nor NOR2 (N7545, N7540, N3181);
nor NOR3 (N7546, N7525, N7533, N6444);
xor XOR2 (N7547, N7545, N1997);
not NOT1 (N7548, N7534);
xor XOR2 (N7549, N7546, N3807);
xor XOR2 (N7550, N7549, N5919);
buf BUF1 (N7551, N7544);
or OR2 (N7552, N7541, N1217);
nor NOR4 (N7553, N7538, N5438, N2017, N1676);
not NOT1 (N7554, N7552);
xor XOR2 (N7555, N7535, N1067);
or OR4 (N7556, N7548, N1329, N233, N2274);
and AND3 (N7557, N7547, N2907, N6523);
nor NOR3 (N7558, N7553, N6917, N1628);
not NOT1 (N7559, N7557);
nand NAND3 (N7560, N7555, N3593, N3029);
nor NOR4 (N7561, N7543, N2843, N110, N4941);
nor NOR2 (N7562, N7556, N6176);
or OR3 (N7563, N7551, N2046, N4695);
and AND4 (N7564, N7550, N3506, N2093, N4916);
or OR3 (N7565, N7563, N16, N3337);
and AND2 (N7566, N7554, N3464);
buf BUF1 (N7567, N7527);
or OR4 (N7568, N7560, N6901, N6976, N2044);
buf BUF1 (N7569, N7565);
xor XOR2 (N7570, N7566, N3372);
xor XOR2 (N7571, N7562, N5587);
nor NOR3 (N7572, N7571, N3560, N5507);
buf BUF1 (N7573, N7558);
xor XOR2 (N7574, N7573, N501);
not NOT1 (N7575, N7559);
nand NAND4 (N7576, N7575, N1420, N1899, N280);
buf BUF1 (N7577, N7531);
not NOT1 (N7578, N7576);
nand NAND2 (N7579, N7572, N638);
nand NAND4 (N7580, N7564, N6037, N2641, N4744);
or OR4 (N7581, N7580, N4178, N2344, N1069);
not NOT1 (N7582, N7568);
or OR2 (N7583, N7569, N6729);
nor NOR4 (N7584, N7577, N2393, N2383, N904);
nor NOR4 (N7585, N7561, N4719, N4167, N176);
not NOT1 (N7586, N7584);
and AND2 (N7587, N7582, N6070);
not NOT1 (N7588, N7585);
nor NOR4 (N7589, N7581, N1214, N1213, N3946);
and AND4 (N7590, N7588, N1497, N623, N1101);
and AND3 (N7591, N7587, N1152, N7180);
not NOT1 (N7592, N7574);
or OR4 (N7593, N7592, N2965, N4318, N2593);
not NOT1 (N7594, N7570);
buf BUF1 (N7595, N7578);
buf BUF1 (N7596, N7590);
and AND2 (N7597, N7593, N640);
buf BUF1 (N7598, N7579);
or OR3 (N7599, N7567, N4259, N319);
nor NOR4 (N7600, N7595, N5459, N7514, N4655);
nand NAND3 (N7601, N7589, N3323, N3979);
xor XOR2 (N7602, N7599, N3779);
buf BUF1 (N7603, N7583);
nand NAND4 (N7604, N7598, N2963, N1792, N2691);
buf BUF1 (N7605, N7594);
nor NOR4 (N7606, N7605, N2620, N5813, N3872);
or OR2 (N7607, N7601, N2283);
or OR2 (N7608, N7586, N1541);
xor XOR2 (N7609, N7597, N3239);
not NOT1 (N7610, N7606);
nand NAND2 (N7611, N7610, N5208);
buf BUF1 (N7612, N7600);
xor XOR2 (N7613, N7604, N6829);
nor NOR2 (N7614, N7612, N2497);
not NOT1 (N7615, N7609);
not NOT1 (N7616, N7603);
or OR2 (N7617, N7615, N1965);
not NOT1 (N7618, N7616);
nand NAND3 (N7619, N7618, N2858, N4050);
buf BUF1 (N7620, N7614);
not NOT1 (N7621, N7591);
not NOT1 (N7622, N7617);
buf BUF1 (N7623, N7613);
not NOT1 (N7624, N7622);
xor XOR2 (N7625, N7596, N560);
or OR3 (N7626, N7625, N6259, N5242);
nor NOR2 (N7627, N7619, N2311);
not NOT1 (N7628, N7623);
buf BUF1 (N7629, N7611);
or OR4 (N7630, N7628, N825, N5990, N2294);
and AND4 (N7631, N7626, N5198, N11, N5674);
buf BUF1 (N7632, N7608);
or OR2 (N7633, N7630, N1537);
buf BUF1 (N7634, N7629);
buf BUF1 (N7635, N7607);
nor NOR2 (N7636, N7627, N6581);
buf BUF1 (N7637, N7621);
buf BUF1 (N7638, N7636);
and AND2 (N7639, N7632, N5093);
or OR2 (N7640, N7639, N3536);
and AND3 (N7641, N7624, N7129, N3623);
or OR3 (N7642, N7634, N3066, N3138);
and AND4 (N7643, N7641, N1965, N2525, N143);
xor XOR2 (N7644, N7638, N2135);
nand NAND4 (N7645, N7602, N652, N5478, N450);
xor XOR2 (N7646, N7637, N3630);
and AND4 (N7647, N7620, N5604, N5702, N565);
not NOT1 (N7648, N7633);
not NOT1 (N7649, N7647);
nor NOR2 (N7650, N7643, N2612);
or OR2 (N7651, N7631, N2263);
not NOT1 (N7652, N7650);
and AND2 (N7653, N7635, N2832);
buf BUF1 (N7654, N7649);
nand NAND4 (N7655, N7654, N4602, N5359, N5328);
and AND2 (N7656, N7646, N634);
xor XOR2 (N7657, N7652, N4687);
buf BUF1 (N7658, N7644);
and AND2 (N7659, N7645, N4395);
buf BUF1 (N7660, N7657);
nand NAND2 (N7661, N7655, N5894);
or OR3 (N7662, N7651, N3474, N2979);
not NOT1 (N7663, N7656);
and AND4 (N7664, N7648, N6048, N6467, N3898);
nor NOR3 (N7665, N7661, N6025, N7307);
buf BUF1 (N7666, N7662);
not NOT1 (N7667, N7659);
nor NOR2 (N7668, N7653, N5832);
and AND4 (N7669, N7663, N886, N2586, N7536);
nand NAND3 (N7670, N7666, N921, N5140);
not NOT1 (N7671, N7640);
nand NAND2 (N7672, N7667, N7064);
not NOT1 (N7673, N7665);
or OR2 (N7674, N7669, N4560);
or OR4 (N7675, N7658, N332, N3355, N3175);
nand NAND2 (N7676, N7673, N5152);
not NOT1 (N7677, N7675);
and AND2 (N7678, N7671, N3119);
not NOT1 (N7679, N7664);
xor XOR2 (N7680, N7642, N1065);
buf BUF1 (N7681, N7674);
and AND4 (N7682, N7679, N290, N6350, N7665);
nand NAND4 (N7683, N7681, N2698, N4473, N4914);
and AND3 (N7684, N7683, N6909, N6305);
nand NAND2 (N7685, N7680, N4386);
nor NOR2 (N7686, N7670, N234);
or OR2 (N7687, N7686, N439);
nand NAND3 (N7688, N7687, N3108, N537);
nor NOR3 (N7689, N7672, N1738, N1698);
xor XOR2 (N7690, N7689, N5562);
and AND4 (N7691, N7676, N1468, N4123, N1423);
or OR3 (N7692, N7691, N3245, N6682);
nand NAND3 (N7693, N7685, N3445, N2059);
or OR4 (N7694, N7678, N5657, N3918, N2421);
or OR4 (N7695, N7677, N6094, N5837, N3484);
nand NAND2 (N7696, N7690, N3977);
or OR2 (N7697, N7668, N7162);
and AND4 (N7698, N7695, N6255, N987, N2764);
not NOT1 (N7699, N7697);
buf BUF1 (N7700, N7688);
buf BUF1 (N7701, N7699);
nor NOR4 (N7702, N7684, N2850, N4625, N46);
not NOT1 (N7703, N7692);
and AND2 (N7704, N7682, N3118);
or OR3 (N7705, N7694, N5837, N4674);
not NOT1 (N7706, N7693);
nand NAND4 (N7707, N7700, N788, N136, N22);
or OR4 (N7708, N7704, N7159, N6114, N6425);
xor XOR2 (N7709, N7706, N3850);
nor NOR4 (N7710, N7701, N4283, N3723, N4362);
buf BUF1 (N7711, N7696);
xor XOR2 (N7712, N7705, N4753);
nand NAND3 (N7713, N7711, N2753, N4085);
nand NAND4 (N7714, N7713, N7675, N7295, N4041);
or OR2 (N7715, N7660, N1267);
xor XOR2 (N7716, N7710, N4785);
xor XOR2 (N7717, N7709, N1010);
or OR3 (N7718, N7708, N2150, N614);
nor NOR2 (N7719, N7712, N3092);
nand NAND4 (N7720, N7716, N4068, N4992, N5015);
xor XOR2 (N7721, N7702, N4751);
not NOT1 (N7722, N7703);
xor XOR2 (N7723, N7714, N5478);
and AND2 (N7724, N7698, N2653);
xor XOR2 (N7725, N7719, N43);
buf BUF1 (N7726, N7707);
xor XOR2 (N7727, N7723, N173);
xor XOR2 (N7728, N7726, N4354);
and AND4 (N7729, N7721, N2248, N6761, N5525);
nor NOR3 (N7730, N7728, N5600, N1606);
nor NOR4 (N7731, N7718, N3024, N3838, N7052);
xor XOR2 (N7732, N7715, N3203);
nor NOR3 (N7733, N7730, N185, N3659);
not NOT1 (N7734, N7717);
xor XOR2 (N7735, N7725, N4831);
nor NOR3 (N7736, N7729, N5790, N6302);
nor NOR2 (N7737, N7735, N2540);
buf BUF1 (N7738, N7736);
xor XOR2 (N7739, N7722, N1731);
nor NOR3 (N7740, N7739, N7709, N981);
not NOT1 (N7741, N7732);
nand NAND3 (N7742, N7738, N3511, N637);
not NOT1 (N7743, N7733);
nor NOR3 (N7744, N7741, N7296, N830);
nor NOR3 (N7745, N7720, N1056, N6635);
nand NAND3 (N7746, N7743, N2652, N4127);
or OR3 (N7747, N7731, N7401, N4673);
not NOT1 (N7748, N7734);
and AND3 (N7749, N7742, N1104, N6711);
buf BUF1 (N7750, N7744);
and AND3 (N7751, N7747, N7477, N2460);
buf BUF1 (N7752, N7727);
and AND2 (N7753, N7745, N5578);
and AND2 (N7754, N7752, N1635);
not NOT1 (N7755, N7751);
not NOT1 (N7756, N7746);
or OR3 (N7757, N7755, N7463, N2496);
not NOT1 (N7758, N7756);
nor NOR3 (N7759, N7724, N6265, N7701);
and AND2 (N7760, N7754, N5734);
xor XOR2 (N7761, N7760, N7082);
buf BUF1 (N7762, N7740);
nand NAND4 (N7763, N7748, N2368, N3608, N3388);
nand NAND2 (N7764, N7750, N6073);
buf BUF1 (N7765, N7757);
nor NOR3 (N7766, N7762, N232, N6942);
nor NOR2 (N7767, N7765, N6822);
nor NOR3 (N7768, N7759, N897, N720);
not NOT1 (N7769, N7768);
or OR4 (N7770, N7753, N7316, N7570, N3878);
xor XOR2 (N7771, N7749, N1771);
buf BUF1 (N7772, N7763);
xor XOR2 (N7773, N7771, N2834);
xor XOR2 (N7774, N7761, N6195);
buf BUF1 (N7775, N7772);
nand NAND2 (N7776, N7764, N2365);
buf BUF1 (N7777, N7774);
or OR2 (N7778, N7776, N3305);
and AND2 (N7779, N7777, N427);
nor NOR2 (N7780, N7778, N2193);
not NOT1 (N7781, N7769);
or OR3 (N7782, N7779, N2110, N2951);
or OR3 (N7783, N7758, N6580, N7762);
and AND4 (N7784, N7781, N6258, N7020, N2692);
or OR2 (N7785, N7783, N4504);
and AND3 (N7786, N7775, N2587, N2265);
and AND2 (N7787, N7767, N1229);
nor NOR3 (N7788, N7787, N6012, N4621);
not NOT1 (N7789, N7782);
and AND3 (N7790, N7785, N1746, N7449);
or OR2 (N7791, N7789, N3240);
not NOT1 (N7792, N7786);
or OR4 (N7793, N7792, N7558, N7673, N3848);
nand NAND2 (N7794, N7770, N1606);
xor XOR2 (N7795, N7794, N1745);
buf BUF1 (N7796, N7795);
or OR2 (N7797, N7773, N3725);
nor NOR2 (N7798, N7788, N5146);
and AND2 (N7799, N7797, N5908);
nand NAND2 (N7800, N7793, N2910);
xor XOR2 (N7801, N7737, N270);
buf BUF1 (N7802, N7784);
xor XOR2 (N7803, N7791, N409);
and AND4 (N7804, N7798, N3075, N3684, N3034);
xor XOR2 (N7805, N7802, N7628);
nor NOR3 (N7806, N7796, N728, N4622);
or OR3 (N7807, N7805, N3783, N1530);
or OR4 (N7808, N7806, N2198, N258, N2525);
not NOT1 (N7809, N7790);
and AND3 (N7810, N7807, N5856, N2634);
nand NAND4 (N7811, N7801, N2038, N1209, N7785);
buf BUF1 (N7812, N7811);
xor XOR2 (N7813, N7810, N6527);
or OR2 (N7814, N7812, N4353);
and AND2 (N7815, N7814, N399);
or OR4 (N7816, N7803, N6182, N177, N5100);
buf BUF1 (N7817, N7809);
and AND2 (N7818, N7808, N1033);
not NOT1 (N7819, N7817);
not NOT1 (N7820, N7819);
nor NOR2 (N7821, N7780, N3578);
not NOT1 (N7822, N7818);
or OR4 (N7823, N7799, N679, N7385, N5498);
buf BUF1 (N7824, N7800);
and AND4 (N7825, N7766, N1480, N6595, N4915);
not NOT1 (N7826, N7822);
xor XOR2 (N7827, N7815, N442);
buf BUF1 (N7828, N7816);
not NOT1 (N7829, N7813);
nand NAND4 (N7830, N7827, N7706, N4230, N5743);
buf BUF1 (N7831, N7823);
nor NOR4 (N7832, N7824, N56, N1335, N6433);
xor XOR2 (N7833, N7804, N1020);
xor XOR2 (N7834, N7820, N6618);
nand NAND3 (N7835, N7831, N6487, N5008);
xor XOR2 (N7836, N7833, N3810);
nor NOR3 (N7837, N7828, N7095, N3340);
xor XOR2 (N7838, N7821, N4626);
not NOT1 (N7839, N7829);
nor NOR3 (N7840, N7830, N927, N2135);
not NOT1 (N7841, N7832);
buf BUF1 (N7842, N7826);
xor XOR2 (N7843, N7825, N564);
or OR3 (N7844, N7834, N3912, N2812);
not NOT1 (N7845, N7842);
nand NAND2 (N7846, N7840, N7013);
not NOT1 (N7847, N7844);
not NOT1 (N7848, N7837);
not NOT1 (N7849, N7838);
nand NAND3 (N7850, N7841, N1069, N7209);
nor NOR4 (N7851, N7848, N1700, N2132, N723);
xor XOR2 (N7852, N7849, N659);
not NOT1 (N7853, N7835);
not NOT1 (N7854, N7852);
or OR4 (N7855, N7836, N2463, N4801, N3857);
or OR2 (N7856, N7851, N171);
and AND4 (N7857, N7853, N6895, N3467, N6013);
not NOT1 (N7858, N7855);
not NOT1 (N7859, N7854);
and AND2 (N7860, N7857, N836);
and AND3 (N7861, N7845, N1500, N835);
not NOT1 (N7862, N7847);
nor NOR2 (N7863, N7861, N3056);
and AND3 (N7864, N7856, N2844, N3608);
xor XOR2 (N7865, N7863, N3409);
nand NAND2 (N7866, N7839, N7396);
not NOT1 (N7867, N7858);
and AND3 (N7868, N7859, N7259, N7211);
or OR4 (N7869, N7867, N6979, N3710, N2507);
buf BUF1 (N7870, N7869);
nor NOR4 (N7871, N7870, N6360, N5095, N7196);
nor NOR4 (N7872, N7850, N658, N6581, N6169);
nor NOR4 (N7873, N7843, N134, N2648, N6049);
nand NAND4 (N7874, N7873, N7233, N4779, N6992);
nand NAND3 (N7875, N7865, N64, N6731);
buf BUF1 (N7876, N7868);
buf BUF1 (N7877, N7875);
or OR3 (N7878, N7862, N866, N204);
or OR2 (N7879, N7874, N5303);
nand NAND3 (N7880, N7876, N5408, N1994);
not NOT1 (N7881, N7879);
xor XOR2 (N7882, N7881, N5347);
not NOT1 (N7883, N7880);
xor XOR2 (N7884, N7864, N1028);
or OR4 (N7885, N7884, N2886, N727, N3943);
not NOT1 (N7886, N7883);
nor NOR3 (N7887, N7886, N2702, N5638);
and AND3 (N7888, N7882, N5782, N4628);
nor NOR4 (N7889, N7878, N7711, N7340, N3276);
or OR2 (N7890, N7889, N2041);
buf BUF1 (N7891, N7846);
xor XOR2 (N7892, N7866, N214);
and AND2 (N7893, N7872, N1621);
and AND4 (N7894, N7877, N6081, N7682, N6766);
nand NAND3 (N7895, N7893, N3220, N4039);
nand NAND4 (N7896, N7871, N5967, N2685, N1788);
not NOT1 (N7897, N7860);
nor NOR3 (N7898, N7892, N5022, N4774);
buf BUF1 (N7899, N7891);
nor NOR3 (N7900, N7885, N453, N7655);
or OR4 (N7901, N7888, N7702, N34, N5763);
not NOT1 (N7902, N7887);
and AND4 (N7903, N7890, N2681, N4932, N4858);
buf BUF1 (N7904, N7901);
or OR3 (N7905, N7904, N5532, N5749);
buf BUF1 (N7906, N7898);
buf BUF1 (N7907, N7896);
nor NOR2 (N7908, N7900, N6982);
not NOT1 (N7909, N7906);
xor XOR2 (N7910, N7903, N7230);
xor XOR2 (N7911, N7897, N3424);
or OR4 (N7912, N7905, N4247, N7165, N6402);
xor XOR2 (N7913, N7907, N1067);
not NOT1 (N7914, N7894);
nand NAND2 (N7915, N7913, N5071);
xor XOR2 (N7916, N7899, N2703);
buf BUF1 (N7917, N7916);
xor XOR2 (N7918, N7912, N1191);
or OR3 (N7919, N7914, N827, N2566);
nor NOR3 (N7920, N7895, N5670, N2887);
or OR2 (N7921, N7911, N2707);
buf BUF1 (N7922, N7908);
and AND3 (N7923, N7920, N6817, N3671);
or OR4 (N7924, N7921, N5725, N4560, N289);
nand NAND2 (N7925, N7918, N572);
not NOT1 (N7926, N7922);
nand NAND3 (N7927, N7926, N7716, N735);
nor NOR2 (N7928, N7910, N6566);
nand NAND4 (N7929, N7924, N1073, N2231, N4478);
and AND2 (N7930, N7902, N1879);
xor XOR2 (N7931, N7927, N7882);
xor XOR2 (N7932, N7909, N2335);
nand NAND4 (N7933, N7932, N3908, N7150, N2381);
xor XOR2 (N7934, N7925, N1147);
buf BUF1 (N7935, N7919);
xor XOR2 (N7936, N7930, N5735);
or OR4 (N7937, N7935, N1421, N6902, N261);
or OR4 (N7938, N7929, N2345, N4546, N7261);
not NOT1 (N7939, N7917);
and AND4 (N7940, N7938, N6685, N1201, N5537);
nor NOR2 (N7941, N7937, N5942);
xor XOR2 (N7942, N7933, N7107);
or OR2 (N7943, N7941, N2960);
buf BUF1 (N7944, N7928);
nor NOR2 (N7945, N7934, N3439);
nand NAND2 (N7946, N7936, N237);
or OR4 (N7947, N7931, N4200, N5634, N7235);
xor XOR2 (N7948, N7940, N3246);
xor XOR2 (N7949, N7942, N2700);
nor NOR3 (N7950, N7948, N7937, N3521);
and AND4 (N7951, N7950, N2231, N3725, N4577);
nor NOR4 (N7952, N7949, N3455, N6559, N7209);
or OR3 (N7953, N7946, N2858, N7113);
buf BUF1 (N7954, N7945);
nand NAND3 (N7955, N7953, N5145, N6523);
or OR2 (N7956, N7923, N1376);
not NOT1 (N7957, N7955);
buf BUF1 (N7958, N7944);
and AND3 (N7959, N7947, N287, N7513);
buf BUF1 (N7960, N7954);
or OR2 (N7961, N7958, N3679);
buf BUF1 (N7962, N7956);
buf BUF1 (N7963, N7959);
or OR3 (N7964, N7915, N6120, N7517);
not NOT1 (N7965, N7939);
and AND4 (N7966, N7951, N1164, N3922, N1158);
not NOT1 (N7967, N7952);
nor NOR4 (N7968, N7962, N7723, N3922, N3612);
not NOT1 (N7969, N7966);
not NOT1 (N7970, N7968);
buf BUF1 (N7971, N7969);
xor XOR2 (N7972, N7970, N2246);
and AND2 (N7973, N7957, N4463);
buf BUF1 (N7974, N7971);
xor XOR2 (N7975, N7961, N6750);
or OR3 (N7976, N7973, N3641, N6364);
or OR3 (N7977, N7963, N3474, N5041);
nor NOR4 (N7978, N7967, N4296, N3755, N4506);
xor XOR2 (N7979, N7964, N5764);
not NOT1 (N7980, N7960);
buf BUF1 (N7981, N7943);
buf BUF1 (N7982, N7976);
and AND3 (N7983, N7977, N1894, N7806);
nand NAND2 (N7984, N7983, N7192);
not NOT1 (N7985, N7972);
nand NAND3 (N7986, N7975, N7722, N5413);
or OR4 (N7987, N7979, N5917, N1340, N4245);
xor XOR2 (N7988, N7986, N5494);
nand NAND4 (N7989, N7984, N4483, N6843, N3316);
or OR4 (N7990, N7980, N6998, N1279, N7297);
not NOT1 (N7991, N7989);
buf BUF1 (N7992, N7982);
and AND4 (N7993, N7991, N4332, N2288, N1642);
buf BUF1 (N7994, N7974);
buf BUF1 (N7995, N7993);
xor XOR2 (N7996, N7985, N3970);
or OR2 (N7997, N7965, N7507);
xor XOR2 (N7998, N7990, N7388);
nand NAND4 (N7999, N7981, N7896, N4000, N5787);
buf BUF1 (N8000, N7992);
and AND2 (N8001, N7994, N4851);
and AND3 (N8002, N8000, N6465, N2019);
nor NOR4 (N8003, N7995, N443, N7692, N4747);
buf BUF1 (N8004, N8003);
and AND4 (N8005, N7996, N4809, N1595, N4050);
nor NOR4 (N8006, N8001, N2402, N6128, N200);
or OR4 (N8007, N7999, N3625, N5580, N3491);
nor NOR3 (N8008, N7997, N1049, N3879);
nor NOR4 (N8009, N7987, N1465, N6552, N398);
nor NOR2 (N8010, N8005, N6389);
nand NAND2 (N8011, N8006, N7018);
not NOT1 (N8012, N8002);
nor NOR3 (N8013, N8004, N139, N3737);
not NOT1 (N8014, N7978);
not NOT1 (N8015, N8012);
buf BUF1 (N8016, N8015);
buf BUF1 (N8017, N8013);
not NOT1 (N8018, N7998);
and AND4 (N8019, N8017, N5330, N7410, N7055);
nand NAND2 (N8020, N8008, N4835);
not NOT1 (N8021, N8016);
not NOT1 (N8022, N8009);
and AND3 (N8023, N8011, N2710, N4696);
buf BUF1 (N8024, N8019);
nor NOR3 (N8025, N8007, N914, N7116);
buf BUF1 (N8026, N7988);
not NOT1 (N8027, N8020);
buf BUF1 (N8028, N8026);
buf BUF1 (N8029, N8014);
nand NAND3 (N8030, N8029, N6050, N1219);
nand NAND4 (N8031, N8028, N1712, N3413, N1160);
or OR4 (N8032, N8023, N6950, N5975, N565);
not NOT1 (N8033, N8010);
buf BUF1 (N8034, N8030);
xor XOR2 (N8035, N8031, N6821);
nand NAND3 (N8036, N8021, N428, N7526);
nand NAND3 (N8037, N8025, N6452, N6299);
nand NAND3 (N8038, N8035, N6014, N2713);
nand NAND4 (N8039, N8037, N2495, N428, N1770);
and AND4 (N8040, N8024, N5125, N7303, N457);
nand NAND2 (N8041, N8036, N7356);
or OR3 (N8042, N8038, N1438, N3436);
not NOT1 (N8043, N8040);
xor XOR2 (N8044, N8022, N6902);
and AND4 (N8045, N8044, N3504, N7061, N2258);
and AND2 (N8046, N8045, N6657);
nor NOR4 (N8047, N8039, N1239, N5342, N6057);
nor NOR3 (N8048, N8034, N1120, N3580);
nand NAND4 (N8049, N8042, N6142, N809, N5661);
or OR4 (N8050, N8046, N7438, N7396, N323);
nor NOR4 (N8051, N8047, N2794, N5289, N7732);
xor XOR2 (N8052, N8051, N5116);
nand NAND2 (N8053, N8049, N4466);
not NOT1 (N8054, N8043);
buf BUF1 (N8055, N8027);
xor XOR2 (N8056, N8052, N2830);
not NOT1 (N8057, N8054);
buf BUF1 (N8058, N8050);
and AND2 (N8059, N8048, N7732);
buf BUF1 (N8060, N8053);
and AND4 (N8061, N8058, N6743, N8005, N3768);
buf BUF1 (N8062, N8033);
not NOT1 (N8063, N8041);
not NOT1 (N8064, N8056);
and AND3 (N8065, N8057, N575, N7165);
and AND2 (N8066, N8060, N4709);
not NOT1 (N8067, N8059);
buf BUF1 (N8068, N8032);
not NOT1 (N8069, N8018);
nor NOR4 (N8070, N8066, N532, N1415, N5498);
xor XOR2 (N8071, N8067, N6485);
and AND4 (N8072, N8071, N5857, N1123, N6245);
or OR3 (N8073, N8064, N3008, N6764);
not NOT1 (N8074, N8055);
buf BUF1 (N8075, N8061);
buf BUF1 (N8076, N8065);
not NOT1 (N8077, N8062);
not NOT1 (N8078, N8070);
xor XOR2 (N8079, N8069, N1378);
buf BUF1 (N8080, N8076);
or OR2 (N8081, N8075, N4632);
or OR4 (N8082, N8063, N6329, N7372, N6784);
nand NAND3 (N8083, N8079, N6026, N1033);
xor XOR2 (N8084, N8068, N7112);
not NOT1 (N8085, N8084);
or OR2 (N8086, N8074, N7676);
or OR2 (N8087, N8086, N1064);
or OR3 (N8088, N8078, N7741, N4497);
or OR3 (N8089, N8081, N7484, N4370);
or OR4 (N8090, N8080, N2443, N7233, N7439);
and AND3 (N8091, N8072, N2744, N2777);
or OR3 (N8092, N8082, N4740, N6972);
buf BUF1 (N8093, N8090);
xor XOR2 (N8094, N8093, N4769);
and AND3 (N8095, N8088, N6961, N330);
or OR4 (N8096, N8094, N5738, N278, N661);
nor NOR2 (N8097, N8095, N488);
not NOT1 (N8098, N8077);
not NOT1 (N8099, N8085);
nor NOR4 (N8100, N8098, N3078, N2996, N6624);
xor XOR2 (N8101, N8096, N4054);
nand NAND2 (N8102, N8073, N4470);
and AND2 (N8103, N8087, N3458);
and AND2 (N8104, N8091, N5332);
nand NAND2 (N8105, N8100, N7932);
or OR2 (N8106, N8104, N3526);
buf BUF1 (N8107, N8103);
nand NAND4 (N8108, N8107, N7634, N950, N5471);
buf BUF1 (N8109, N8089);
not NOT1 (N8110, N8106);
xor XOR2 (N8111, N8099, N2106);
xor XOR2 (N8112, N8109, N3133);
not NOT1 (N8113, N8112);
nand NAND3 (N8114, N8113, N7191, N6090);
nand NAND4 (N8115, N8101, N7146, N4010, N7550);
nor NOR2 (N8116, N8115, N746);
nand NAND3 (N8117, N8116, N6606, N3622);
nor NOR4 (N8118, N8102, N1956, N6140, N6948);
xor XOR2 (N8119, N8114, N5481);
not NOT1 (N8120, N8105);
and AND4 (N8121, N8097, N3795, N4750, N7829);
nand NAND3 (N8122, N8092, N4738, N1014);
or OR2 (N8123, N8122, N7759);
and AND3 (N8124, N8108, N3403, N2363);
nand NAND4 (N8125, N8121, N3106, N4790, N4339);
not NOT1 (N8126, N8120);
or OR3 (N8127, N8118, N3585, N6127);
or OR4 (N8128, N8083, N1822, N4925, N1051);
not NOT1 (N8129, N8111);
or OR3 (N8130, N8127, N1835, N5941);
nand NAND4 (N8131, N8129, N3203, N2036, N6194);
xor XOR2 (N8132, N8124, N4811);
buf BUF1 (N8133, N8119);
not NOT1 (N8134, N8128);
nor NOR3 (N8135, N8126, N7178, N1904);
buf BUF1 (N8136, N8132);
and AND3 (N8137, N8123, N8086, N5169);
nor NOR3 (N8138, N8134, N4077, N6145);
buf BUF1 (N8139, N8117);
not NOT1 (N8140, N8110);
nand NAND2 (N8141, N8139, N4102);
and AND4 (N8142, N8138, N5690, N1609, N4253);
buf BUF1 (N8143, N8140);
not NOT1 (N8144, N8143);
nand NAND4 (N8145, N8133, N4668, N3687, N5970);
nand NAND2 (N8146, N8142, N2796);
or OR3 (N8147, N8131, N44, N6196);
not NOT1 (N8148, N8141);
xor XOR2 (N8149, N8145, N8115);
nand NAND2 (N8150, N8147, N2038);
not NOT1 (N8151, N8149);
buf BUF1 (N8152, N8125);
or OR4 (N8153, N8144, N3883, N7800, N9);
and AND4 (N8154, N8130, N3135, N2640, N7554);
nand NAND2 (N8155, N8152, N6658);
buf BUF1 (N8156, N8154);
xor XOR2 (N8157, N8155, N3585);
or OR2 (N8158, N8136, N499);
buf BUF1 (N8159, N8151);
or OR3 (N8160, N8157, N6336, N4385);
nor NOR4 (N8161, N8146, N3357, N4851, N6427);
or OR4 (N8162, N8156, N7604, N6537, N3754);
xor XOR2 (N8163, N8150, N6231);
or OR3 (N8164, N8137, N2972, N8052);
buf BUF1 (N8165, N8158);
nor NOR4 (N8166, N8135, N6913, N7449, N2059);
nor NOR2 (N8167, N8160, N6157);
or OR2 (N8168, N8167, N2262);
not NOT1 (N8169, N8163);
not NOT1 (N8170, N8161);
buf BUF1 (N8171, N8169);
xor XOR2 (N8172, N8159, N3692);
buf BUF1 (N8173, N8168);
and AND2 (N8174, N8162, N3463);
nand NAND3 (N8175, N8166, N7208, N5519);
nor NOR2 (N8176, N8164, N149);
not NOT1 (N8177, N8165);
not NOT1 (N8178, N8173);
nand NAND2 (N8179, N8153, N3771);
and AND2 (N8180, N8178, N6773);
buf BUF1 (N8181, N8172);
xor XOR2 (N8182, N8179, N815);
nor NOR2 (N8183, N8181, N6901);
not NOT1 (N8184, N8171);
nand NAND3 (N8185, N8183, N6685, N3954);
nand NAND4 (N8186, N8177, N4649, N5033, N2912);
nand NAND2 (N8187, N8176, N1909);
xor XOR2 (N8188, N8185, N6958);
buf BUF1 (N8189, N8182);
not NOT1 (N8190, N8170);
nand NAND3 (N8191, N8175, N7612, N1674);
or OR2 (N8192, N8189, N3675);
and AND2 (N8193, N8191, N3432);
xor XOR2 (N8194, N8187, N4785);
and AND2 (N8195, N8194, N1750);
xor XOR2 (N8196, N8192, N5843);
xor XOR2 (N8197, N8186, N519);
or OR3 (N8198, N8188, N3047, N1207);
not NOT1 (N8199, N8196);
not NOT1 (N8200, N8198);
not NOT1 (N8201, N8197);
buf BUF1 (N8202, N8199);
and AND3 (N8203, N8200, N4771, N1417);
nor NOR3 (N8204, N8174, N76, N1503);
or OR4 (N8205, N8202, N5116, N6165, N7425);
or OR4 (N8206, N8180, N8049, N2130, N5641);
or OR4 (N8207, N8190, N2779, N3356, N5942);
buf BUF1 (N8208, N8204);
or OR3 (N8209, N8184, N7652, N6809);
or OR3 (N8210, N8193, N326, N4047);
and AND2 (N8211, N8203, N2277);
nor NOR2 (N8212, N8210, N1902);
or OR3 (N8213, N8212, N581, N7905);
xor XOR2 (N8214, N8206, N2136);
nand NAND4 (N8215, N8201, N5185, N1437, N792);
and AND3 (N8216, N8205, N7790, N4010);
xor XOR2 (N8217, N8211, N2878);
nand NAND4 (N8218, N8215, N4570, N1096, N4998);
xor XOR2 (N8219, N8148, N3096);
not NOT1 (N8220, N8209);
and AND3 (N8221, N8213, N4009, N1542);
buf BUF1 (N8222, N8207);
nand NAND2 (N8223, N8221, N3500);
buf BUF1 (N8224, N8217);
or OR4 (N8225, N8208, N1617, N6811, N810);
not NOT1 (N8226, N8214);
nor NOR3 (N8227, N8195, N568, N6915);
nor NOR2 (N8228, N8218, N6237);
and AND4 (N8229, N8223, N859, N6651, N8066);
and AND3 (N8230, N8219, N7892, N5210);
xor XOR2 (N8231, N8226, N1575);
nor NOR2 (N8232, N8229, N1644);
not NOT1 (N8233, N8224);
or OR4 (N8234, N8231, N4144, N5741, N5713);
buf BUF1 (N8235, N8225);
xor XOR2 (N8236, N8233, N2130);
not NOT1 (N8237, N8235);
nand NAND4 (N8238, N8222, N5251, N6233, N1394);
not NOT1 (N8239, N8216);
nor NOR4 (N8240, N8236, N5473, N4231, N3882);
nor NOR4 (N8241, N8239, N4894, N2600, N5646);
nor NOR2 (N8242, N8227, N5792);
buf BUF1 (N8243, N8238);
nand NAND2 (N8244, N8243, N6765);
xor XOR2 (N8245, N8244, N3057);
xor XOR2 (N8246, N8234, N593);
not NOT1 (N8247, N8230);
nand NAND4 (N8248, N8245, N8208, N4475, N2466);
and AND3 (N8249, N8220, N2053, N1656);
not NOT1 (N8250, N8246);
or OR3 (N8251, N8242, N7012, N1343);
nor NOR4 (N8252, N8251, N1706, N8020, N1039);
xor XOR2 (N8253, N8240, N7210);
xor XOR2 (N8254, N8249, N3475);
not NOT1 (N8255, N8252);
or OR2 (N8256, N8248, N787);
nand NAND3 (N8257, N8228, N2446, N782);
buf BUF1 (N8258, N8250);
and AND2 (N8259, N8253, N7123);
nor NOR2 (N8260, N8232, N2777);
buf BUF1 (N8261, N8258);
buf BUF1 (N8262, N8237);
nor NOR3 (N8263, N8261, N3980, N7273);
or OR4 (N8264, N8256, N1940, N227, N5956);
and AND3 (N8265, N8255, N6487, N7815);
buf BUF1 (N8266, N8265);
nand NAND4 (N8267, N8266, N7789, N306, N5416);
not NOT1 (N8268, N8263);
xor XOR2 (N8269, N8267, N5040);
or OR2 (N8270, N8268, N7404);
nor NOR4 (N8271, N8264, N3925, N4502, N3455);
or OR2 (N8272, N8270, N5845);
nor NOR3 (N8273, N8260, N5942, N7507);
xor XOR2 (N8274, N8254, N3582);
nor NOR2 (N8275, N8271, N6230);
buf BUF1 (N8276, N8273);
nand NAND3 (N8277, N8257, N7672, N1721);
buf BUF1 (N8278, N8247);
not NOT1 (N8279, N8276);
or OR3 (N8280, N8269, N3668, N1209);
xor XOR2 (N8281, N8262, N8108);
or OR3 (N8282, N8279, N176, N5919);
nor NOR4 (N8283, N8278, N7914, N6732, N2891);
xor XOR2 (N8284, N8241, N5353);
and AND2 (N8285, N8282, N3259);
not NOT1 (N8286, N8272);
and AND2 (N8287, N8275, N4726);
or OR2 (N8288, N8274, N4498);
buf BUF1 (N8289, N8281);
buf BUF1 (N8290, N8283);
not NOT1 (N8291, N8259);
buf BUF1 (N8292, N8287);
or OR2 (N8293, N8290, N6374);
nor NOR2 (N8294, N8293, N6995);
nand NAND3 (N8295, N8285, N7519, N8083);
nand NAND3 (N8296, N8291, N1192, N1013);
not NOT1 (N8297, N8284);
nor NOR2 (N8298, N8280, N8265);
nand NAND3 (N8299, N8298, N6646, N5018);
nand NAND4 (N8300, N8286, N7664, N8202, N5726);
xor XOR2 (N8301, N8296, N858);
and AND3 (N8302, N8295, N7439, N551);
or OR2 (N8303, N8294, N1026);
xor XOR2 (N8304, N8297, N264);
buf BUF1 (N8305, N8299);
xor XOR2 (N8306, N8305, N581);
or OR3 (N8307, N8302, N2850, N1644);
not NOT1 (N8308, N8303);
not NOT1 (N8309, N8300);
xor XOR2 (N8310, N8307, N142);
nor NOR4 (N8311, N8301, N3933, N3475, N7738);
not NOT1 (N8312, N8309);
xor XOR2 (N8313, N8312, N1294);
nor NOR4 (N8314, N8289, N2515, N3206, N5436);
buf BUF1 (N8315, N8304);
nand NAND4 (N8316, N8277, N6404, N7481, N1705);
xor XOR2 (N8317, N8314, N5526);
and AND4 (N8318, N8315, N4897, N3082, N1606);
not NOT1 (N8319, N8308);
or OR2 (N8320, N8313, N3072);
nor NOR4 (N8321, N8288, N3446, N8001, N7325);
not NOT1 (N8322, N8320);
xor XOR2 (N8323, N8318, N509);
buf BUF1 (N8324, N8292);
and AND2 (N8325, N8319, N6015);
and AND4 (N8326, N8311, N7230, N4265, N4735);
nand NAND2 (N8327, N8323, N6023);
xor XOR2 (N8328, N8310, N2027);
buf BUF1 (N8329, N8327);
xor XOR2 (N8330, N8325, N4665);
not NOT1 (N8331, N8321);
not NOT1 (N8332, N8324);
nand NAND3 (N8333, N8328, N7841, N6978);
not NOT1 (N8334, N8329);
buf BUF1 (N8335, N8317);
or OR3 (N8336, N8316, N5778, N5349);
and AND3 (N8337, N8336, N1549, N6770);
and AND4 (N8338, N8326, N7705, N5317, N5214);
and AND2 (N8339, N8334, N2670);
nor NOR2 (N8340, N8335, N6915);
nor NOR3 (N8341, N8332, N76, N6098);
xor XOR2 (N8342, N8306, N6845);
or OR2 (N8343, N8331, N4641);
nand NAND3 (N8344, N8330, N3089, N6925);
or OR2 (N8345, N8339, N2265);
not NOT1 (N8346, N8340);
or OR4 (N8347, N8344, N6145, N8066, N4435);
xor XOR2 (N8348, N8342, N5730);
or OR2 (N8349, N8346, N4282);
and AND4 (N8350, N8341, N6919, N6990, N5094);
nor NOR2 (N8351, N8343, N280);
xor XOR2 (N8352, N8337, N2862);
buf BUF1 (N8353, N8322);
nand NAND3 (N8354, N8349, N2262, N7641);
and AND2 (N8355, N8347, N8112);
not NOT1 (N8356, N8351);
or OR2 (N8357, N8352, N504);
xor XOR2 (N8358, N8348, N7914);
nor NOR2 (N8359, N8338, N3002);
nor NOR3 (N8360, N8353, N4428, N4507);
buf BUF1 (N8361, N8357);
or OR3 (N8362, N8359, N4532, N2203);
and AND2 (N8363, N8356, N5384);
xor XOR2 (N8364, N8358, N6364);
and AND2 (N8365, N8361, N6486);
or OR2 (N8366, N8345, N8256);
nand NAND2 (N8367, N8360, N4597);
nor NOR4 (N8368, N8367, N2406, N3659, N2376);
not NOT1 (N8369, N8355);
and AND4 (N8370, N8362, N7907, N3366, N6618);
nor NOR4 (N8371, N8364, N7342, N5938, N3820);
not NOT1 (N8372, N8368);
xor XOR2 (N8373, N8366, N3478);
and AND4 (N8374, N8363, N7616, N4048, N6221);
not NOT1 (N8375, N8333);
buf BUF1 (N8376, N8369);
buf BUF1 (N8377, N8354);
not NOT1 (N8378, N8370);
or OR4 (N8379, N8378, N4478, N4220, N6520);
buf BUF1 (N8380, N8371);
xor XOR2 (N8381, N8380, N4918);
nor NOR2 (N8382, N8375, N2200);
nand NAND4 (N8383, N8377, N7907, N3992, N4164);
or OR3 (N8384, N8382, N5987, N3296);
nor NOR3 (N8385, N8376, N1049, N8021);
nand NAND3 (N8386, N8384, N3722, N5920);
buf BUF1 (N8387, N8383);
xor XOR2 (N8388, N8373, N775);
buf BUF1 (N8389, N8374);
nor NOR4 (N8390, N8350, N422, N6551, N7192);
xor XOR2 (N8391, N8387, N3704);
nor NOR3 (N8392, N8388, N5770, N1411);
or OR4 (N8393, N8379, N1053, N6971, N734);
nor NOR3 (N8394, N8381, N5218, N6036);
not NOT1 (N8395, N8393);
or OR3 (N8396, N8391, N2727, N3025);
or OR3 (N8397, N8385, N478, N2596);
nand NAND3 (N8398, N8390, N286, N4452);
not NOT1 (N8399, N8398);
nor NOR3 (N8400, N8397, N4599, N3438);
and AND4 (N8401, N8400, N283, N6722, N6832);
and AND2 (N8402, N8396, N2121);
not NOT1 (N8403, N8392);
xor XOR2 (N8404, N8402, N1349);
or OR4 (N8405, N8399, N2443, N3256, N4209);
nor NOR3 (N8406, N8401, N6188, N451);
nand NAND4 (N8407, N8395, N6990, N1739, N1574);
and AND4 (N8408, N8404, N191, N5895, N5820);
buf BUF1 (N8409, N8394);
nand NAND3 (N8410, N8407, N1447, N5707);
or OR4 (N8411, N8389, N7923, N7528, N1558);
nor NOR2 (N8412, N8406, N4779);
not NOT1 (N8413, N8411);
nand NAND3 (N8414, N8403, N101, N7953);
xor XOR2 (N8415, N8386, N7555);
nand NAND4 (N8416, N8412, N8127, N4966, N8242);
buf BUF1 (N8417, N8408);
nor NOR3 (N8418, N8417, N2578, N6149);
buf BUF1 (N8419, N8410);
or OR3 (N8420, N8418, N3192, N7658);
buf BUF1 (N8421, N8372);
buf BUF1 (N8422, N8409);
buf BUF1 (N8423, N8415);
and AND4 (N8424, N8416, N6333, N4383, N1515);
nor NOR4 (N8425, N8424, N5796, N1312, N4012);
nor NOR3 (N8426, N8413, N7776, N7877);
nand NAND2 (N8427, N8423, N3142);
nand NAND2 (N8428, N8425, N7982);
or OR3 (N8429, N8422, N277, N6396);
or OR3 (N8430, N8414, N1945, N595);
and AND3 (N8431, N8426, N5855, N3598);
nand NAND4 (N8432, N8420, N4066, N752, N1476);
xor XOR2 (N8433, N8432, N3776);
and AND4 (N8434, N8431, N1290, N463, N2546);
xor XOR2 (N8435, N8430, N6807);
buf BUF1 (N8436, N8365);
nor NOR2 (N8437, N8436, N4523);
nor NOR2 (N8438, N8433, N4427);
nand NAND4 (N8439, N8419, N4456, N1102, N2428);
or OR2 (N8440, N8439, N8360);
not NOT1 (N8441, N8437);
nor NOR3 (N8442, N8438, N6491, N8105);
not NOT1 (N8443, N8405);
and AND4 (N8444, N8427, N7118, N5818, N360);
buf BUF1 (N8445, N8442);
or OR2 (N8446, N8434, N5109);
or OR3 (N8447, N8444, N5209, N6480);
and AND4 (N8448, N8428, N7550, N299, N4209);
and AND4 (N8449, N8440, N5361, N2996, N2753);
not NOT1 (N8450, N8445);
buf BUF1 (N8451, N8450);
or OR2 (N8452, N8448, N4580);
or OR3 (N8453, N8435, N4615, N3223);
nand NAND2 (N8454, N8446, N6629);
xor XOR2 (N8455, N8451, N6110);
xor XOR2 (N8456, N8452, N816);
not NOT1 (N8457, N8456);
nor NOR2 (N8458, N8453, N4710);
nand NAND4 (N8459, N8429, N6950, N864, N6499);
not NOT1 (N8460, N8455);
nand NAND2 (N8461, N8457, N3327);
nand NAND4 (N8462, N8459, N2516, N1816, N3138);
nand NAND4 (N8463, N8458, N3043, N6499, N4442);
nor NOR4 (N8464, N8462, N108, N4329, N7739);
buf BUF1 (N8465, N8460);
not NOT1 (N8466, N8421);
nand NAND4 (N8467, N8465, N7948, N7301, N2352);
buf BUF1 (N8468, N8464);
or OR2 (N8469, N8441, N7922);
nand NAND2 (N8470, N8467, N1766);
buf BUF1 (N8471, N8468);
nand NAND2 (N8472, N8443, N1083);
nand NAND4 (N8473, N8449, N3651, N5354, N3659);
xor XOR2 (N8474, N8461, N2721);
not NOT1 (N8475, N8454);
buf BUF1 (N8476, N8472);
buf BUF1 (N8477, N8476);
buf BUF1 (N8478, N8474);
nand NAND3 (N8479, N8477, N8305, N1613);
nand NAND4 (N8480, N8475, N4464, N8293, N7576);
or OR4 (N8481, N8473, N8051, N1017, N6390);
nand NAND4 (N8482, N8480, N7642, N7198, N624);
and AND3 (N8483, N8478, N6702, N7992);
not NOT1 (N8484, N8463);
xor XOR2 (N8485, N8470, N1960);
xor XOR2 (N8486, N8466, N4072);
xor XOR2 (N8487, N8485, N7602);
nand NAND2 (N8488, N8483, N4906);
nor NOR2 (N8489, N8469, N3840);
nand NAND3 (N8490, N8479, N4526, N1468);
buf BUF1 (N8491, N8487);
not NOT1 (N8492, N8486);
nor NOR4 (N8493, N8488, N7674, N8134, N7126);
or OR4 (N8494, N8491, N5846, N909, N2000);
not NOT1 (N8495, N8489);
nor NOR4 (N8496, N8471, N3415, N7315, N799);
or OR3 (N8497, N8490, N7838, N6541);
xor XOR2 (N8498, N8493, N5338);
buf BUF1 (N8499, N8481);
nand NAND4 (N8500, N8495, N3845, N6471, N5118);
nor NOR3 (N8501, N8484, N1181, N8031);
buf BUF1 (N8502, N8501);
xor XOR2 (N8503, N8498, N6625);
nor NOR4 (N8504, N8503, N3479, N2894, N1389);
or OR3 (N8505, N8494, N4476, N3342);
not NOT1 (N8506, N8499);
or OR4 (N8507, N8506, N3806, N3659, N7188);
nand NAND2 (N8508, N8500, N7079);
and AND3 (N8509, N8507, N1677, N463);
xor XOR2 (N8510, N8497, N4744);
and AND2 (N8511, N8492, N1576);
nor NOR3 (N8512, N8496, N5783, N2933);
not NOT1 (N8513, N8508);
not NOT1 (N8514, N8482);
or OR2 (N8515, N8505, N4750);
and AND3 (N8516, N8512, N1621, N1929);
not NOT1 (N8517, N8511);
or OR3 (N8518, N8515, N6506, N4461);
or OR2 (N8519, N8509, N369);
or OR2 (N8520, N8516, N3508);
or OR3 (N8521, N8519, N364, N1663);
not NOT1 (N8522, N8520);
nand NAND4 (N8523, N8514, N230, N1208, N4811);
or OR4 (N8524, N8518, N2790, N2635, N4350);
nor NOR2 (N8525, N8513, N1733);
buf BUF1 (N8526, N8517);
nor NOR4 (N8527, N8523, N2080, N3587, N3999);
nand NAND3 (N8528, N8447, N6890, N4102);
and AND3 (N8529, N8526, N3386, N7866);
not NOT1 (N8530, N8510);
nand NAND3 (N8531, N8529, N1161, N8003);
nor NOR2 (N8532, N8502, N4720);
nand NAND3 (N8533, N8504, N1604, N2330);
nor NOR4 (N8534, N8532, N5399, N4841, N4955);
xor XOR2 (N8535, N8534, N2484);
and AND4 (N8536, N8522, N1404, N1210, N3144);
buf BUF1 (N8537, N8527);
buf BUF1 (N8538, N8524);
or OR3 (N8539, N8535, N4385, N8454);
not NOT1 (N8540, N8525);
xor XOR2 (N8541, N8538, N135);
nand NAND3 (N8542, N8528, N5939, N2497);
not NOT1 (N8543, N8536);
nand NAND2 (N8544, N8531, N6446);
and AND4 (N8545, N8537, N5270, N7432, N6390);
nand NAND3 (N8546, N8541, N1755, N7046);
xor XOR2 (N8547, N8533, N2774);
xor XOR2 (N8548, N8547, N1309);
and AND4 (N8549, N8543, N1987, N6497, N186);
or OR2 (N8550, N8542, N5230);
buf BUF1 (N8551, N8545);
nand NAND4 (N8552, N8551, N1481, N155, N2052);
and AND4 (N8553, N8530, N5093, N159, N6082);
or OR4 (N8554, N8550, N3372, N1254, N1730);
not NOT1 (N8555, N8553);
xor XOR2 (N8556, N8544, N1367);
not NOT1 (N8557, N8521);
not NOT1 (N8558, N8546);
nand NAND3 (N8559, N8558, N3742, N7639);
nor NOR2 (N8560, N8554, N5061);
xor XOR2 (N8561, N8556, N7205);
or OR2 (N8562, N8539, N511);
or OR3 (N8563, N8549, N6626, N7183);
buf BUF1 (N8564, N8560);
not NOT1 (N8565, N8559);
nand NAND4 (N8566, N8552, N6992, N1170, N94);
nand NAND3 (N8567, N8555, N7212, N3535);
nand NAND2 (N8568, N8548, N916);
not NOT1 (N8569, N8561);
nor NOR3 (N8570, N8567, N2084, N7535);
or OR3 (N8571, N8540, N3050, N3413);
not NOT1 (N8572, N8565);
nand NAND3 (N8573, N8570, N4839, N6351);
or OR4 (N8574, N8566, N21, N1739, N4705);
or OR2 (N8575, N8569, N6096);
or OR3 (N8576, N8574, N7029, N6740);
or OR4 (N8577, N8576, N8125, N3494, N2006);
not NOT1 (N8578, N8568);
buf BUF1 (N8579, N8578);
and AND4 (N8580, N8557, N4726, N2559, N2177);
or OR3 (N8581, N8564, N6637, N5545);
or OR3 (N8582, N8573, N3766, N2052);
and AND4 (N8583, N8575, N2074, N7681, N5509);
buf BUF1 (N8584, N8580);
not NOT1 (N8585, N8562);
xor XOR2 (N8586, N8583, N1172);
or OR3 (N8587, N8571, N8481, N316);
nand NAND4 (N8588, N8585, N143, N6489, N1809);
or OR3 (N8589, N8572, N3864, N669);
or OR2 (N8590, N8588, N1600);
or OR2 (N8591, N8563, N1665);
nand NAND2 (N8592, N8582, N6316);
and AND2 (N8593, N8586, N4181);
nor NOR3 (N8594, N8579, N8137, N8394);
xor XOR2 (N8595, N8584, N1892);
xor XOR2 (N8596, N8593, N2996);
buf BUF1 (N8597, N8581);
and AND4 (N8598, N8590, N1061, N7692, N1957);
xor XOR2 (N8599, N8577, N388);
nand NAND2 (N8600, N8591, N5891);
nor NOR4 (N8601, N8599, N7331, N918, N8191);
nand NAND2 (N8602, N8592, N4062);
or OR4 (N8603, N8601, N2771, N3216, N2695);
nand NAND4 (N8604, N8603, N3931, N220, N5850);
nor NOR4 (N8605, N8602, N2418, N3360, N5266);
or OR2 (N8606, N8596, N6963);
not NOT1 (N8607, N8594);
and AND2 (N8608, N8606, N3395);
buf BUF1 (N8609, N8595);
not NOT1 (N8610, N8589);
xor XOR2 (N8611, N8598, N8302);
nor NOR2 (N8612, N8597, N3810);
xor XOR2 (N8613, N8610, N5659);
nor NOR3 (N8614, N8609, N7915, N3985);
or OR2 (N8615, N8600, N7912);
buf BUF1 (N8616, N8614);
or OR2 (N8617, N8616, N349);
buf BUF1 (N8618, N8607);
nand NAND2 (N8619, N8604, N5548);
xor XOR2 (N8620, N8608, N3525);
and AND2 (N8621, N8617, N991);
buf BUF1 (N8622, N8587);
and AND2 (N8623, N8615, N5325);
not NOT1 (N8624, N8623);
not NOT1 (N8625, N8621);
not NOT1 (N8626, N8605);
or OR4 (N8627, N8611, N2969, N2160, N4067);
and AND2 (N8628, N8626, N3556);
xor XOR2 (N8629, N8627, N174);
xor XOR2 (N8630, N8625, N5937);
or OR4 (N8631, N8629, N1637, N1291, N6488);
buf BUF1 (N8632, N8612);
and AND3 (N8633, N8619, N3666, N7044);
xor XOR2 (N8634, N8628, N6929);
nor NOR4 (N8635, N8622, N5439, N7478, N2149);
xor XOR2 (N8636, N8632, N5188);
buf BUF1 (N8637, N8630);
or OR3 (N8638, N8637, N4470, N3525);
xor XOR2 (N8639, N8618, N3475);
xor XOR2 (N8640, N8624, N2989);
nor NOR2 (N8641, N8631, N3908);
and AND4 (N8642, N8613, N2465, N4178, N5259);
buf BUF1 (N8643, N8640);
buf BUF1 (N8644, N8639);
and AND4 (N8645, N8644, N8314, N35, N1715);
and AND4 (N8646, N8642, N3230, N5430, N7189);
or OR3 (N8647, N8646, N7657, N7116);
or OR2 (N8648, N8634, N483);
nand NAND3 (N8649, N8645, N1061, N8014);
nand NAND3 (N8650, N8620, N6658, N2417);
xor XOR2 (N8651, N8638, N1011);
or OR3 (N8652, N8635, N8413, N5908);
xor XOR2 (N8653, N8648, N1006);
buf BUF1 (N8654, N8647);
xor XOR2 (N8655, N8641, N234);
buf BUF1 (N8656, N8650);
nand NAND3 (N8657, N8654, N31, N8507);
nand NAND2 (N8658, N8651, N145);
nor NOR3 (N8659, N8633, N8227, N7659);
nand NAND2 (N8660, N8655, N3168);
buf BUF1 (N8661, N8652);
buf BUF1 (N8662, N8660);
xor XOR2 (N8663, N8649, N1439);
or OR2 (N8664, N8636, N92);
not NOT1 (N8665, N8643);
buf BUF1 (N8666, N8658);
not NOT1 (N8667, N8656);
and AND4 (N8668, N8665, N6056, N8366, N7622);
xor XOR2 (N8669, N8659, N5504);
or OR2 (N8670, N8666, N4151);
nor NOR2 (N8671, N8670, N4407);
nand NAND4 (N8672, N8663, N3521, N206, N7515);
nand NAND3 (N8673, N8661, N3902, N520);
nand NAND2 (N8674, N8673, N3590);
xor XOR2 (N8675, N8669, N3653);
and AND2 (N8676, N8675, N3101);
not NOT1 (N8677, N8672);
or OR3 (N8678, N8653, N6894, N4893);
not NOT1 (N8679, N8657);
not NOT1 (N8680, N8678);
and AND4 (N8681, N8671, N6143, N1372, N6926);
nand NAND3 (N8682, N8677, N7120, N6650);
buf BUF1 (N8683, N8667);
and AND3 (N8684, N8682, N7974, N6972);
nand NAND2 (N8685, N8676, N120);
or OR4 (N8686, N8664, N5406, N5808, N7116);
nor NOR3 (N8687, N8685, N4046, N4635);
not NOT1 (N8688, N8680);
nor NOR2 (N8689, N8681, N4595);
or OR2 (N8690, N8686, N4327);
nor NOR4 (N8691, N8679, N3264, N3569, N4080);
and AND3 (N8692, N8688, N8308, N4361);
and AND3 (N8693, N8683, N2203, N5475);
or OR2 (N8694, N8690, N3495);
nor NOR2 (N8695, N8668, N3271);
nor NOR4 (N8696, N8692, N983, N7217, N4525);
not NOT1 (N8697, N8696);
buf BUF1 (N8698, N8674);
nor NOR4 (N8699, N8698, N2527, N8412, N2146);
buf BUF1 (N8700, N8697);
buf BUF1 (N8701, N8699);
and AND4 (N8702, N8689, N4217, N4165, N3015);
xor XOR2 (N8703, N8691, N1706);
and AND2 (N8704, N8662, N4758);
xor XOR2 (N8705, N8693, N5554);
or OR4 (N8706, N8695, N6721, N1661, N5923);
and AND3 (N8707, N8701, N5659, N3631);
and AND4 (N8708, N8706, N5904, N1364, N6679);
not NOT1 (N8709, N8702);
buf BUF1 (N8710, N8687);
buf BUF1 (N8711, N8700);
buf BUF1 (N8712, N8708);
buf BUF1 (N8713, N8710);
or OR3 (N8714, N8709, N6210, N4288);
nor NOR3 (N8715, N8703, N3916, N6646);
xor XOR2 (N8716, N8711, N5412);
nand NAND4 (N8717, N8714, N7821, N76, N3727);
buf BUF1 (N8718, N8712);
nand NAND2 (N8719, N8717, N8090);
nor NOR2 (N8720, N8715, N3143);
not NOT1 (N8721, N8719);
nand NAND2 (N8722, N8716, N2388);
xor XOR2 (N8723, N8722, N1853);
nor NOR3 (N8724, N8704, N4463, N8258);
nor NOR2 (N8725, N8707, N4734);
not NOT1 (N8726, N8713);
nand NAND2 (N8727, N8723, N7371);
xor XOR2 (N8728, N8724, N7461);
not NOT1 (N8729, N8727);
or OR4 (N8730, N8729, N7597, N2120, N8632);
buf BUF1 (N8731, N8726);
xor XOR2 (N8732, N8684, N546);
nand NAND2 (N8733, N8718, N8091);
nand NAND2 (N8734, N8732, N3986);
nand NAND4 (N8735, N8728, N3063, N1526, N6142);
and AND3 (N8736, N8730, N8704, N2290);
xor XOR2 (N8737, N8731, N8034);
nor NOR4 (N8738, N8736, N7361, N5443, N8386);
nand NAND4 (N8739, N8733, N5454, N3752, N3953);
xor XOR2 (N8740, N8737, N4989);
xor XOR2 (N8741, N8738, N2663);
and AND4 (N8742, N8694, N6598, N5732, N4305);
nand NAND4 (N8743, N8742, N7074, N8351, N6620);
xor XOR2 (N8744, N8720, N5569);
xor XOR2 (N8745, N8740, N4070);
not NOT1 (N8746, N8739);
nor NOR2 (N8747, N8734, N7401);
xor XOR2 (N8748, N8741, N5915);
not NOT1 (N8749, N8743);
or OR4 (N8750, N8746, N7419, N7148, N7027);
and AND3 (N8751, N8747, N5871, N1516);
nor NOR2 (N8752, N8745, N6079);
and AND3 (N8753, N8725, N4317, N2544);
and AND3 (N8754, N8705, N2118, N1821);
xor XOR2 (N8755, N8749, N3848);
nand NAND4 (N8756, N8748, N7424, N3417, N5102);
nor NOR3 (N8757, N8755, N3984, N4100);
or OR2 (N8758, N8744, N466);
nand NAND2 (N8759, N8750, N6605);
and AND4 (N8760, N8756, N3982, N6655, N7270);
xor XOR2 (N8761, N8753, N4554);
nand NAND4 (N8762, N8758, N1397, N5862, N3795);
nand NAND3 (N8763, N8760, N1277, N7795);
xor XOR2 (N8764, N8761, N3683);
or OR2 (N8765, N8762, N2436);
nand NAND4 (N8766, N8763, N5551, N5670, N7973);
or OR4 (N8767, N8752, N7689, N2487, N3531);
nor NOR2 (N8768, N8764, N1838);
xor XOR2 (N8769, N8767, N8660);
nand NAND2 (N8770, N8721, N3039);
xor XOR2 (N8771, N8770, N8332);
or OR2 (N8772, N8751, N1048);
nor NOR3 (N8773, N8754, N4691, N1171);
buf BUF1 (N8774, N8759);
and AND4 (N8775, N8765, N5806, N599, N2880);
or OR3 (N8776, N8773, N3995, N8724);
xor XOR2 (N8777, N8774, N296);
or OR4 (N8778, N8775, N7252, N5813, N6703);
nand NAND3 (N8779, N8778, N544, N30);
buf BUF1 (N8780, N8771);
or OR4 (N8781, N8768, N3021, N155, N7985);
and AND3 (N8782, N8766, N2121, N2499);
nor NOR3 (N8783, N8735, N5521, N7671);
and AND4 (N8784, N8772, N3939, N3050, N121);
buf BUF1 (N8785, N8779);
not NOT1 (N8786, N8776);
nor NOR4 (N8787, N8781, N1065, N1779, N5740);
buf BUF1 (N8788, N8784);
nor NOR2 (N8789, N8780, N4169);
xor XOR2 (N8790, N8787, N473);
and AND3 (N8791, N8769, N7859, N8060);
buf BUF1 (N8792, N8790);
nor NOR3 (N8793, N8788, N3825, N476);
buf BUF1 (N8794, N8785);
and AND3 (N8795, N8782, N6714, N5856);
xor XOR2 (N8796, N8757, N4452);
nand NAND4 (N8797, N8793, N5261, N6863, N2063);
nand NAND4 (N8798, N8786, N3156, N2565, N5568);
nor NOR3 (N8799, N8777, N8490, N3303);
and AND2 (N8800, N8797, N7169);
buf BUF1 (N8801, N8791);
xor XOR2 (N8802, N8799, N6914);
not NOT1 (N8803, N8796);
not NOT1 (N8804, N8792);
nor NOR3 (N8805, N8803, N6548, N658);
buf BUF1 (N8806, N8794);
nor NOR2 (N8807, N8806, N3329);
not NOT1 (N8808, N8798);
nand NAND4 (N8809, N8783, N2150, N2513, N4084);
nor NOR2 (N8810, N8801, N3435);
not NOT1 (N8811, N8808);
or OR3 (N8812, N8809, N4996, N773);
not NOT1 (N8813, N8795);
xor XOR2 (N8814, N8800, N7092);
not NOT1 (N8815, N8814);
or OR3 (N8816, N8805, N272, N4091);
buf BUF1 (N8817, N8812);
not NOT1 (N8818, N8807);
nor NOR3 (N8819, N8815, N4458, N5407);
nand NAND2 (N8820, N8816, N3152);
nand NAND4 (N8821, N8817, N6165, N4645, N2535);
buf BUF1 (N8822, N8820);
and AND2 (N8823, N8818, N3154);
not NOT1 (N8824, N8810);
xor XOR2 (N8825, N8789, N3112);
or OR4 (N8826, N8811, N2979, N8719, N3723);
buf BUF1 (N8827, N8823);
or OR3 (N8828, N8804, N3854, N4748);
and AND4 (N8829, N8819, N8109, N2221, N4903);
xor XOR2 (N8830, N8826, N1401);
nand NAND4 (N8831, N8825, N3017, N1490, N874);
buf BUF1 (N8832, N8824);
buf BUF1 (N8833, N8813);
not NOT1 (N8834, N8827);
not NOT1 (N8835, N8834);
xor XOR2 (N8836, N8829, N7613);
buf BUF1 (N8837, N8836);
nand NAND2 (N8838, N8833, N7160);
and AND2 (N8839, N8835, N6642);
or OR4 (N8840, N8802, N2119, N468, N3003);
not NOT1 (N8841, N8840);
buf BUF1 (N8842, N8830);
and AND3 (N8843, N8821, N3904, N4692);
not NOT1 (N8844, N8841);
and AND2 (N8845, N8844, N7035);
or OR2 (N8846, N8843, N2931);
not NOT1 (N8847, N8846);
or OR3 (N8848, N8831, N7692, N4731);
buf BUF1 (N8849, N8822);
nor NOR4 (N8850, N8837, N1215, N6409, N3282);
xor XOR2 (N8851, N8838, N76);
or OR2 (N8852, N8832, N848);
nand NAND2 (N8853, N8847, N896);
nor NOR4 (N8854, N8852, N2469, N6100, N8140);
not NOT1 (N8855, N8842);
nor NOR3 (N8856, N8848, N3242, N3345);
buf BUF1 (N8857, N8845);
and AND3 (N8858, N8849, N8843, N4928);
or OR2 (N8859, N8850, N7843);
not NOT1 (N8860, N8853);
not NOT1 (N8861, N8856);
xor XOR2 (N8862, N8851, N2872);
buf BUF1 (N8863, N8861);
and AND4 (N8864, N8863, N4571, N4811, N5101);
nand NAND3 (N8865, N8864, N958, N1095);
xor XOR2 (N8866, N8865, N5938);
nand NAND2 (N8867, N8839, N2280);
nor NOR2 (N8868, N8855, N1591);
and AND2 (N8869, N8866, N5076);
not NOT1 (N8870, N8869);
xor XOR2 (N8871, N8867, N3291);
xor XOR2 (N8872, N8870, N6181);
not NOT1 (N8873, N8854);
or OR4 (N8874, N8862, N3571, N5425, N5303);
and AND4 (N8875, N8871, N1748, N7152, N6393);
not NOT1 (N8876, N8874);
not NOT1 (N8877, N8857);
nand NAND2 (N8878, N8858, N5398);
nand NAND2 (N8879, N8878, N2570);
nor NOR4 (N8880, N8876, N5508, N1872, N3966);
not NOT1 (N8881, N8859);
and AND4 (N8882, N8868, N5938, N5819, N2822);
not NOT1 (N8883, N8860);
or OR4 (N8884, N8881, N3839, N5330, N7037);
and AND4 (N8885, N8873, N2798, N2290, N6388);
not NOT1 (N8886, N8879);
and AND4 (N8887, N8885, N2396, N8236, N6813);
nand NAND3 (N8888, N8887, N4586, N8162);
buf BUF1 (N8889, N8828);
not NOT1 (N8890, N8877);
nand NAND2 (N8891, N8875, N2811);
not NOT1 (N8892, N8888);
and AND2 (N8893, N8872, N6512);
or OR2 (N8894, N8891, N3538);
buf BUF1 (N8895, N8890);
buf BUF1 (N8896, N8894);
and AND4 (N8897, N8889, N2636, N3224, N6099);
and AND3 (N8898, N8892, N5041, N908);
nand NAND3 (N8899, N8898, N5089, N3508);
not NOT1 (N8900, N8884);
not NOT1 (N8901, N8900);
nand NAND2 (N8902, N8886, N2237);
not NOT1 (N8903, N8893);
and AND4 (N8904, N8901, N5687, N2209, N4227);
buf BUF1 (N8905, N8895);
not NOT1 (N8906, N8904);
or OR4 (N8907, N8906, N3865, N2479, N4348);
and AND4 (N8908, N8903, N6225, N752, N6556);
buf BUF1 (N8909, N8897);
xor XOR2 (N8910, N8896, N4260);
nor NOR4 (N8911, N8880, N6856, N5653, N7766);
not NOT1 (N8912, N8882);
buf BUF1 (N8913, N8883);
nor NOR4 (N8914, N8909, N5916, N7894, N8680);
buf BUF1 (N8915, N8905);
and AND2 (N8916, N8915, N6544);
not NOT1 (N8917, N8902);
nand NAND2 (N8918, N8910, N8076);
xor XOR2 (N8919, N8916, N4070);
not NOT1 (N8920, N8899);
and AND4 (N8921, N8913, N1159, N5378, N6135);
nand NAND4 (N8922, N8907, N3246, N8654, N6968);
nand NAND4 (N8923, N8917, N90, N6348, N1065);
and AND2 (N8924, N8922, N3345);
nand NAND2 (N8925, N8919, N7634);
xor XOR2 (N8926, N8920, N6087);
xor XOR2 (N8927, N8924, N8342);
or OR2 (N8928, N8908, N1753);
buf BUF1 (N8929, N8923);
nor NOR2 (N8930, N8911, N1267);
not NOT1 (N8931, N8925);
nor NOR3 (N8932, N8926, N5522, N6674);
nor NOR2 (N8933, N8928, N1575);
and AND2 (N8934, N8914, N5781);
and AND3 (N8935, N8931, N341, N5880);
buf BUF1 (N8936, N8935);
nand NAND3 (N8937, N8927, N7622, N2680);
xor XOR2 (N8938, N8933, N6757);
buf BUF1 (N8939, N8938);
not NOT1 (N8940, N8936);
xor XOR2 (N8941, N8934, N2559);
or OR4 (N8942, N8939, N600, N1266, N6282);
buf BUF1 (N8943, N8918);
not NOT1 (N8944, N8942);
buf BUF1 (N8945, N8932);
nor NOR4 (N8946, N8945, N4440, N970, N7135);
buf BUF1 (N8947, N8921);
nand NAND2 (N8948, N8946, N2276);
nand NAND3 (N8949, N8929, N3042, N8540);
and AND3 (N8950, N8944, N6816, N1135);
not NOT1 (N8951, N8937);
buf BUF1 (N8952, N8940);
nor NOR3 (N8953, N8930, N8347, N6980);
xor XOR2 (N8954, N8953, N7327);
not NOT1 (N8955, N8949);
not NOT1 (N8956, N8951);
buf BUF1 (N8957, N8943);
xor XOR2 (N8958, N8954, N3917);
or OR4 (N8959, N8956, N3016, N5922, N8278);
xor XOR2 (N8960, N8948, N8759);
not NOT1 (N8961, N8941);
or OR2 (N8962, N8947, N7393);
not NOT1 (N8963, N8962);
or OR2 (N8964, N8958, N7301);
or OR4 (N8965, N8964, N4947, N5070, N6650);
buf BUF1 (N8966, N8950);
and AND4 (N8967, N8966, N3404, N3202, N7921);
nor NOR4 (N8968, N8961, N8607, N8430, N5729);
xor XOR2 (N8969, N8968, N6289);
not NOT1 (N8970, N8967);
nand NAND2 (N8971, N8963, N8808);
and AND2 (N8972, N8957, N6208);
nor NOR3 (N8973, N8971, N3426, N6448);
or OR2 (N8974, N8959, N1004);
not NOT1 (N8975, N8965);
nor NOR3 (N8976, N8912, N2410, N8071);
nor NOR3 (N8977, N8970, N8410, N4016);
nand NAND4 (N8978, N8973, N6734, N2221, N6952);
or OR3 (N8979, N8960, N7670, N7787);
xor XOR2 (N8980, N8979, N8171);
and AND3 (N8981, N8974, N1503, N8484);
and AND4 (N8982, N8955, N442, N7067, N279);
buf BUF1 (N8983, N8975);
not NOT1 (N8984, N8980);
buf BUF1 (N8985, N8984);
or OR3 (N8986, N8969, N7194, N4699);
nor NOR4 (N8987, N8985, N2043, N3527, N2307);
nand NAND3 (N8988, N8982, N7145, N7295);
nand NAND4 (N8989, N8981, N8441, N4309, N3131);
and AND4 (N8990, N8986, N6505, N2795, N7029);
not NOT1 (N8991, N8983);
nand NAND2 (N8992, N8991, N8360);
nand NAND3 (N8993, N8987, N3798, N472);
buf BUF1 (N8994, N8976);
not NOT1 (N8995, N8994);
nand NAND3 (N8996, N8993, N4161, N5060);
buf BUF1 (N8997, N8996);
buf BUF1 (N8998, N8972);
nor NOR3 (N8999, N8997, N1951, N7487);
or OR4 (N9000, N8992, N6609, N464, N4422);
not NOT1 (N9001, N8999);
not NOT1 (N9002, N9001);
or OR4 (N9003, N8998, N1050, N7715, N5687);
nor NOR4 (N9004, N8977, N4779, N2220, N4502);
and AND4 (N9005, N9004, N2059, N527, N4979);
or OR4 (N9006, N8978, N3006, N4213, N3912);
nand NAND4 (N9007, N9005, N7013, N8173, N4018);
nand NAND3 (N9008, N9003, N5761, N622);
xor XOR2 (N9009, N8990, N8990);
not NOT1 (N9010, N8988);
nand NAND3 (N9011, N9007, N5653, N4160);
nand NAND2 (N9012, N8989, N4913);
nor NOR2 (N9013, N8995, N4786);
buf BUF1 (N9014, N9002);
or OR2 (N9015, N9012, N4259);
not NOT1 (N9016, N9006);
nand NAND2 (N9017, N9008, N1871);
xor XOR2 (N9018, N9013, N4063);
buf BUF1 (N9019, N9000);
nor NOR2 (N9020, N9010, N1499);
not NOT1 (N9021, N9019);
buf BUF1 (N9022, N9011);
nor NOR4 (N9023, N9020, N7769, N8064, N7882);
xor XOR2 (N9024, N9016, N5172);
or OR2 (N9025, N9017, N8278);
nand NAND4 (N9026, N9022, N653, N4717, N4064);
not NOT1 (N9027, N9009);
not NOT1 (N9028, N9026);
and AND4 (N9029, N9024, N1917, N4649, N2270);
nor NOR3 (N9030, N9028, N6562, N705);
buf BUF1 (N9031, N9025);
nor NOR2 (N9032, N9015, N1283);
not NOT1 (N9033, N9031);
buf BUF1 (N9034, N9018);
and AND2 (N9035, N9033, N2939);
nand NAND2 (N9036, N9030, N3711);
nand NAND3 (N9037, N9023, N7154, N3425);
buf BUF1 (N9038, N9036);
xor XOR2 (N9039, N9021, N8376);
or OR3 (N9040, N9014, N5075, N515);
nor NOR4 (N9041, N9037, N3802, N4832, N7424);
and AND2 (N9042, N9027, N5689);
xor XOR2 (N9043, N9038, N3843);
nor NOR2 (N9044, N9029, N3737);
or OR4 (N9045, N8952, N4389, N2228, N6949);
nand NAND2 (N9046, N9034, N4502);
buf BUF1 (N9047, N9040);
and AND4 (N9048, N9043, N1806, N2818, N8152);
and AND2 (N9049, N9046, N2583);
xor XOR2 (N9050, N9032, N6882);
nand NAND2 (N9051, N9041, N4443);
nand NAND3 (N9052, N9044, N3380, N4456);
or OR2 (N9053, N9051, N7008);
nand NAND4 (N9054, N9035, N438, N4996, N4876);
nor NOR2 (N9055, N9047, N3760);
and AND3 (N9056, N9050, N8822, N7347);
nor NOR4 (N9057, N9053, N864, N7034, N5002);
nand NAND3 (N9058, N9054, N7730, N4362);
buf BUF1 (N9059, N9039);
xor XOR2 (N9060, N9052, N5214);
or OR3 (N9061, N9058, N9043, N8761);
nand NAND2 (N9062, N9060, N7977);
not NOT1 (N9063, N9045);
not NOT1 (N9064, N9055);
and AND2 (N9065, N9062, N7924);
buf BUF1 (N9066, N9061);
or OR3 (N9067, N9048, N3163, N8687);
or OR2 (N9068, N9059, N1961);
xor XOR2 (N9069, N9042, N5005);
and AND2 (N9070, N9067, N8844);
not NOT1 (N9071, N9068);
nor NOR3 (N9072, N9056, N4888, N4278);
nor NOR2 (N9073, N9049, N1069);
and AND4 (N9074, N9065, N8644, N6777, N8370);
nor NOR3 (N9075, N9066, N8386, N3924);
and AND2 (N9076, N9069, N852);
buf BUF1 (N9077, N9076);
not NOT1 (N9078, N9057);
buf BUF1 (N9079, N9070);
nand NAND4 (N9080, N9071, N6146, N6832, N5449);
buf BUF1 (N9081, N9063);
nor NOR4 (N9082, N9064, N5582, N6577, N7819);
nor NOR2 (N9083, N9082, N5536);
or OR4 (N9084, N9073, N5701, N4773, N1440);
or OR3 (N9085, N9080, N3366, N2325);
not NOT1 (N9086, N9083);
and AND4 (N9087, N9075, N3158, N1993, N8342);
or OR4 (N9088, N9081, N8917, N1469, N6492);
or OR2 (N9089, N9087, N8366);
xor XOR2 (N9090, N9077, N2035);
or OR3 (N9091, N9074, N3233, N2435);
or OR3 (N9092, N9084, N1668, N3149);
and AND4 (N9093, N9089, N2310, N1183, N3885);
not NOT1 (N9094, N9079);
buf BUF1 (N9095, N9072);
xor XOR2 (N9096, N9088, N5472);
and AND3 (N9097, N9085, N4981, N6619);
and AND4 (N9098, N9095, N8940, N8376, N502);
nand NAND4 (N9099, N9091, N6611, N5187, N888);
buf BUF1 (N9100, N9094);
xor XOR2 (N9101, N9086, N353);
nand NAND4 (N9102, N9099, N6429, N8333, N4734);
nand NAND3 (N9103, N9090, N1262, N4092);
not NOT1 (N9104, N9100);
nand NAND4 (N9105, N9101, N2980, N7711, N6046);
not NOT1 (N9106, N9097);
nand NAND3 (N9107, N9092, N659, N5537);
nor NOR3 (N9108, N9096, N6476, N5584);
xor XOR2 (N9109, N9106, N961);
or OR2 (N9110, N9103, N2557);
not NOT1 (N9111, N9078);
or OR4 (N9112, N9109, N6756, N2170, N5806);
xor XOR2 (N9113, N9102, N5449);
xor XOR2 (N9114, N9108, N2515);
xor XOR2 (N9115, N9113, N629);
and AND4 (N9116, N9114, N806, N3360, N2475);
nand NAND4 (N9117, N9115, N5972, N209, N1220);
not NOT1 (N9118, N9093);
xor XOR2 (N9119, N9110, N8400);
buf BUF1 (N9120, N9107);
xor XOR2 (N9121, N9105, N2827);
nor NOR4 (N9122, N9118, N6808, N1841, N3622);
nor NOR3 (N9123, N9122, N4625, N7509);
or OR4 (N9124, N9112, N7279, N8202, N3582);
not NOT1 (N9125, N9121);
not NOT1 (N9126, N9125);
nor NOR2 (N9127, N9119, N4714);
and AND3 (N9128, N9120, N1784, N8459);
buf BUF1 (N9129, N9126);
nor NOR4 (N9130, N9127, N760, N6314, N1400);
not NOT1 (N9131, N9098);
nor NOR2 (N9132, N9117, N3098);
nor NOR4 (N9133, N9104, N2931, N4416, N4502);
and AND4 (N9134, N9123, N2801, N2398, N7804);
xor XOR2 (N9135, N9124, N290);
not NOT1 (N9136, N9133);
and AND2 (N9137, N9128, N8976);
or OR2 (N9138, N9131, N6480);
nand NAND2 (N9139, N9116, N3324);
buf BUF1 (N9140, N9129);
and AND3 (N9141, N9136, N4625, N3249);
buf BUF1 (N9142, N9135);
and AND4 (N9143, N9132, N2480, N1127, N2945);
not NOT1 (N9144, N9143);
xor XOR2 (N9145, N9130, N5623);
nor NOR2 (N9146, N9137, N158);
not NOT1 (N9147, N9141);
xor XOR2 (N9148, N9140, N7972);
or OR2 (N9149, N9145, N8474);
nand NAND2 (N9150, N9138, N6333);
or OR4 (N9151, N9146, N4535, N8599, N8037);
nor NOR3 (N9152, N9139, N1844, N6173);
xor XOR2 (N9153, N9111, N1136);
and AND2 (N9154, N9148, N7979);
not NOT1 (N9155, N9147);
and AND2 (N9156, N9144, N3906);
xor XOR2 (N9157, N9134, N6801);
buf BUF1 (N9158, N9156);
or OR3 (N9159, N9151, N8626, N4501);
and AND4 (N9160, N9159, N1713, N1692, N5158);
xor XOR2 (N9161, N9155, N225);
and AND2 (N9162, N9142, N3922);
buf BUF1 (N9163, N9161);
or OR2 (N9164, N9149, N1141);
not NOT1 (N9165, N9158);
nand NAND3 (N9166, N9162, N364, N899);
or OR2 (N9167, N9160, N1596);
xor XOR2 (N9168, N9164, N95);
nand NAND2 (N9169, N9163, N9026);
buf BUF1 (N9170, N9169);
xor XOR2 (N9171, N9170, N6517);
and AND4 (N9172, N9152, N6484, N5714, N6288);
or OR2 (N9173, N9150, N1450);
or OR2 (N9174, N9167, N8575);
buf BUF1 (N9175, N9153);
not NOT1 (N9176, N9171);
or OR3 (N9177, N9154, N509, N9059);
or OR3 (N9178, N9168, N6594, N6189);
nor NOR4 (N9179, N9175, N8369, N7289, N8227);
xor XOR2 (N9180, N9177, N65);
not NOT1 (N9181, N9176);
and AND4 (N9182, N9178, N1776, N6710, N2009);
nand NAND2 (N9183, N9166, N6915);
not NOT1 (N9184, N9181);
xor XOR2 (N9185, N9165, N6573);
buf BUF1 (N9186, N9185);
nor NOR3 (N9187, N9183, N6793, N7061);
nor NOR2 (N9188, N9179, N5414);
nand NAND3 (N9189, N9173, N5397, N4019);
not NOT1 (N9190, N9172);
and AND2 (N9191, N9188, N2986);
nor NOR3 (N9192, N9174, N7046, N1352);
or OR4 (N9193, N9191, N5378, N4604, N1230);
nand NAND2 (N9194, N9157, N3253);
or OR4 (N9195, N9182, N8245, N7509, N4420);
not NOT1 (N9196, N9193);
not NOT1 (N9197, N9190);
buf BUF1 (N9198, N9180);
nand NAND3 (N9199, N9197, N1756, N3415);
and AND4 (N9200, N9199, N3065, N6688, N8349);
nand NAND2 (N9201, N9194, N4480);
nand NAND2 (N9202, N9192, N5515);
buf BUF1 (N9203, N9184);
not NOT1 (N9204, N9202);
nand NAND3 (N9205, N9204, N1441, N4680);
nand NAND3 (N9206, N9195, N26, N5817);
buf BUF1 (N9207, N9198);
xor XOR2 (N9208, N9196, N6328);
and AND2 (N9209, N9189, N5986);
and AND2 (N9210, N9208, N504);
and AND3 (N9211, N9201, N7762, N4299);
or OR2 (N9212, N9187, N7328);
nand NAND4 (N9213, N9209, N3284, N4109, N9160);
buf BUF1 (N9214, N9213);
or OR3 (N9215, N9186, N1149, N3716);
not NOT1 (N9216, N9207);
or OR2 (N9217, N9205, N6488);
and AND4 (N9218, N9215, N248, N2004, N3932);
buf BUF1 (N9219, N9210);
and AND2 (N9220, N9206, N3654);
not NOT1 (N9221, N9220);
and AND2 (N9222, N9219, N3486);
or OR4 (N9223, N9221, N4097, N2277, N6705);
buf BUF1 (N9224, N9216);
not NOT1 (N9225, N9212);
nand NAND3 (N9226, N9203, N2373, N3815);
nor NOR2 (N9227, N9218, N791);
nor NOR2 (N9228, N9214, N8144);
not NOT1 (N9229, N9223);
nor NOR4 (N9230, N9227, N3154, N8104, N71);
or OR2 (N9231, N9225, N1607);
or OR4 (N9232, N9200, N2218, N1257, N5513);
xor XOR2 (N9233, N9230, N2907);
buf BUF1 (N9234, N9211);
nand NAND2 (N9235, N9233, N8956);
or OR4 (N9236, N9231, N1654, N4384, N2817);
not NOT1 (N9237, N9217);
not NOT1 (N9238, N9234);
nor NOR3 (N9239, N9237, N2338, N5399);
not NOT1 (N9240, N9226);
xor XOR2 (N9241, N9239, N807);
nand NAND4 (N9242, N9235, N1995, N183, N1233);
nor NOR4 (N9243, N9228, N3381, N820, N4971);
buf BUF1 (N9244, N9241);
not NOT1 (N9245, N9222);
nand NAND2 (N9246, N9232, N9188);
nand NAND2 (N9247, N9244, N4503);
buf BUF1 (N9248, N9236);
not NOT1 (N9249, N9247);
and AND4 (N9250, N9224, N7478, N8093, N5053);
or OR2 (N9251, N9229, N8203);
buf BUF1 (N9252, N9243);
buf BUF1 (N9253, N9249);
not NOT1 (N9254, N9252);
buf BUF1 (N9255, N9251);
and AND4 (N9256, N9245, N5351, N5858, N4553);
or OR3 (N9257, N9242, N2849, N1354);
nor NOR3 (N9258, N9246, N2935, N2108);
nor NOR4 (N9259, N9258, N7774, N5659, N9005);
buf BUF1 (N9260, N9250);
and AND3 (N9261, N9238, N5296, N8536);
nand NAND3 (N9262, N9261, N5953, N2591);
xor XOR2 (N9263, N9262, N7462);
nor NOR4 (N9264, N9253, N6999, N6823, N7240);
nand NAND4 (N9265, N9259, N387, N3800, N1988);
xor XOR2 (N9266, N9264, N649);
and AND4 (N9267, N9255, N2894, N8863, N8133);
buf BUF1 (N9268, N9267);
not NOT1 (N9269, N9254);
xor XOR2 (N9270, N9263, N7577);
nand NAND3 (N9271, N9265, N2483, N6460);
nor NOR4 (N9272, N9248, N3670, N303, N1628);
and AND4 (N9273, N9260, N8873, N1515, N8322);
nand NAND4 (N9274, N9256, N8857, N5525, N8609);
or OR4 (N9275, N9269, N770, N8713, N2349);
xor XOR2 (N9276, N9275, N3641);
or OR2 (N9277, N9266, N2451);
nor NOR2 (N9278, N9271, N949);
buf BUF1 (N9279, N9274);
and AND3 (N9280, N9257, N2404, N3809);
nor NOR4 (N9281, N9268, N8510, N3030, N4244);
buf BUF1 (N9282, N9281);
not NOT1 (N9283, N9240);
and AND3 (N9284, N9273, N1063, N5789);
or OR3 (N9285, N9277, N1923, N2663);
buf BUF1 (N9286, N9285);
xor XOR2 (N9287, N9282, N1316);
or OR3 (N9288, N9270, N133, N4424);
xor XOR2 (N9289, N9279, N8905);
xor XOR2 (N9290, N9288, N5796);
xor XOR2 (N9291, N9284, N3588);
xor XOR2 (N9292, N9290, N8978);
and AND2 (N9293, N9291, N8609);
xor XOR2 (N9294, N9278, N8353);
xor XOR2 (N9295, N9289, N1758);
or OR2 (N9296, N9283, N9142);
not NOT1 (N9297, N9296);
buf BUF1 (N9298, N9276);
nor NOR3 (N9299, N9294, N3962, N85);
xor XOR2 (N9300, N9280, N3341);
or OR4 (N9301, N9298, N7937, N1325, N1187);
not NOT1 (N9302, N9293);
nand NAND4 (N9303, N9299, N5601, N4180, N1814);
nor NOR2 (N9304, N9301, N6461);
nor NOR4 (N9305, N9292, N4183, N3153, N5777);
not NOT1 (N9306, N9287);
xor XOR2 (N9307, N9272, N1947);
and AND3 (N9308, N9306, N3922, N1053);
not NOT1 (N9309, N9308);
and AND4 (N9310, N9307, N4124, N9112, N3748);
buf BUF1 (N9311, N9304);
buf BUF1 (N9312, N9295);
nor NOR3 (N9313, N9312, N4914, N3714);
not NOT1 (N9314, N9297);
not NOT1 (N9315, N9305);
nand NAND3 (N9316, N9303, N4115, N4656);
or OR4 (N9317, N9313, N3229, N3010, N1366);
nand NAND4 (N9318, N9310, N3434, N291, N9285);
or OR4 (N9319, N9286, N7348, N7814, N2414);
or OR3 (N9320, N9318, N3500, N2832);
and AND3 (N9321, N9311, N1721, N2554);
xor XOR2 (N9322, N9302, N4696);
and AND4 (N9323, N9300, N5723, N6449, N8321);
nand NAND3 (N9324, N9309, N5645, N4284);
nand NAND3 (N9325, N9323, N2171, N9295);
buf BUF1 (N9326, N9319);
nor NOR4 (N9327, N9324, N6271, N7914, N2950);
not NOT1 (N9328, N9322);
nand NAND3 (N9329, N9326, N587, N2076);
not NOT1 (N9330, N9314);
or OR2 (N9331, N9325, N2979);
xor XOR2 (N9332, N9320, N8421);
or OR2 (N9333, N9321, N6886);
or OR3 (N9334, N9332, N6790, N9067);
nand NAND3 (N9335, N9330, N9217, N8914);
xor XOR2 (N9336, N9327, N7852);
xor XOR2 (N9337, N9333, N7750);
nand NAND2 (N9338, N9315, N8362);
not NOT1 (N9339, N9335);
buf BUF1 (N9340, N9329);
buf BUF1 (N9341, N9338);
xor XOR2 (N9342, N9331, N6240);
and AND2 (N9343, N9341, N7929);
buf BUF1 (N9344, N9339);
nor NOR4 (N9345, N9328, N7981, N8875, N2386);
or OR2 (N9346, N9337, N2227);
not NOT1 (N9347, N9345);
xor XOR2 (N9348, N9344, N1547);
not NOT1 (N9349, N9347);
not NOT1 (N9350, N9317);
xor XOR2 (N9351, N9348, N8748);
buf BUF1 (N9352, N9343);
nand NAND4 (N9353, N9349, N5561, N5403, N9342);
nor NOR4 (N9354, N4866, N3930, N8525, N8481);
or OR4 (N9355, N9354, N1458, N9120, N5606);
not NOT1 (N9356, N9316);
nor NOR2 (N9357, N9350, N5825);
xor XOR2 (N9358, N9334, N1179);
xor XOR2 (N9359, N9358, N7483);
nor NOR2 (N9360, N9340, N2235);
nor NOR3 (N9361, N9352, N372, N1153);
not NOT1 (N9362, N9360);
and AND2 (N9363, N9351, N2497);
buf BUF1 (N9364, N9362);
nand NAND4 (N9365, N9361, N1399, N5868, N2040);
xor XOR2 (N9366, N9357, N874);
or OR2 (N9367, N9364, N1115);
and AND4 (N9368, N9336, N1120, N6513, N4934);
buf BUF1 (N9369, N9346);
nand NAND3 (N9370, N9363, N5258, N3598);
buf BUF1 (N9371, N9366);
not NOT1 (N9372, N9359);
nor NOR2 (N9373, N9371, N2197);
nor NOR2 (N9374, N9370, N7498);
nand NAND2 (N9375, N9368, N5219);
not NOT1 (N9376, N9367);
or OR3 (N9377, N9374, N3711, N4828);
or OR4 (N9378, N9356, N8577, N9028, N680);
nand NAND2 (N9379, N9365, N2797);
nand NAND4 (N9380, N9355, N3177, N1814, N356);
buf BUF1 (N9381, N9377);
nand NAND3 (N9382, N9375, N4528, N4002);
buf BUF1 (N9383, N9379);
nand NAND4 (N9384, N9378, N3376, N6312, N1685);
xor XOR2 (N9385, N9372, N5885);
xor XOR2 (N9386, N9373, N5808);
buf BUF1 (N9387, N9380);
or OR3 (N9388, N9369, N8159, N6152);
or OR2 (N9389, N9381, N5794);
and AND2 (N9390, N9386, N244);
buf BUF1 (N9391, N9353);
nand NAND2 (N9392, N9391, N6647);
nor NOR4 (N9393, N9376, N7591, N5238, N998);
nand NAND3 (N9394, N9393, N5567, N8624);
or OR2 (N9395, N9390, N3261);
xor XOR2 (N9396, N9394, N6441);
nand NAND4 (N9397, N9396, N7663, N4693, N235);
or OR3 (N9398, N9388, N4828, N4740);
or OR4 (N9399, N9387, N7266, N4213, N9160);
not NOT1 (N9400, N9383);
buf BUF1 (N9401, N9398);
nor NOR3 (N9402, N9399, N3622, N5662);
nor NOR4 (N9403, N9389, N9351, N8892, N3878);
not NOT1 (N9404, N9402);
not NOT1 (N9405, N9401);
xor XOR2 (N9406, N9397, N7713);
nand NAND3 (N9407, N9395, N3870, N6205);
or OR2 (N9408, N9403, N7778);
nor NOR2 (N9409, N9392, N7093);
buf BUF1 (N9410, N9400);
nor NOR4 (N9411, N9410, N4225, N1712, N8623);
nand NAND4 (N9412, N9411, N2749, N5450, N7838);
not NOT1 (N9413, N9409);
nor NOR4 (N9414, N9384, N2699, N6098, N5854);
buf BUF1 (N9415, N9413);
buf BUF1 (N9416, N9415);
buf BUF1 (N9417, N9412);
and AND4 (N9418, N9414, N822, N1084, N2365);
buf BUF1 (N9419, N9385);
nand NAND4 (N9420, N9419, N6940, N8753, N2629);
nor NOR4 (N9421, N9416, N7941, N896, N5749);
buf BUF1 (N9422, N9418);
or OR3 (N9423, N9417, N8373, N3353);
not NOT1 (N9424, N9407);
not NOT1 (N9425, N9408);
nand NAND4 (N9426, N9404, N5821, N8375, N1778);
and AND4 (N9427, N9406, N3978, N4107, N1945);
or OR3 (N9428, N9427, N3672, N4504);
nor NOR3 (N9429, N9424, N192, N5507);
or OR2 (N9430, N9420, N683);
or OR2 (N9431, N9425, N8747);
nand NAND3 (N9432, N9428, N2937, N5331);
nand NAND3 (N9433, N9432, N2361, N8341);
buf BUF1 (N9434, N9430);
xor XOR2 (N9435, N9429, N644);
or OR4 (N9436, N9382, N1709, N6947, N3524);
nand NAND4 (N9437, N9434, N2110, N7463, N6211);
not NOT1 (N9438, N9421);
and AND2 (N9439, N9435, N156);
xor XOR2 (N9440, N9423, N6997);
xor XOR2 (N9441, N9440, N8041);
buf BUF1 (N9442, N9426);
or OR3 (N9443, N9442, N6241, N8992);
or OR4 (N9444, N9441, N8540, N5076, N5261);
nand NAND4 (N9445, N9443, N6288, N5053, N2201);
or OR3 (N9446, N9437, N719, N119);
buf BUF1 (N9447, N9436);
and AND3 (N9448, N9444, N6973, N2152);
nand NAND4 (N9449, N9431, N63, N5417, N886);
xor XOR2 (N9450, N9433, N4714);
not NOT1 (N9451, N9449);
xor XOR2 (N9452, N9438, N8166);
not NOT1 (N9453, N9405);
xor XOR2 (N9454, N9439, N3427);
xor XOR2 (N9455, N9452, N830);
and AND4 (N9456, N9422, N3056, N2742, N6320);
not NOT1 (N9457, N9455);
buf BUF1 (N9458, N9451);
nand NAND3 (N9459, N9450, N2182, N2885);
buf BUF1 (N9460, N9446);
buf BUF1 (N9461, N9448);
or OR4 (N9462, N9460, N6209, N5940, N3141);
buf BUF1 (N9463, N9447);
and AND4 (N9464, N9453, N1404, N733, N1298);
nor NOR2 (N9465, N9461, N1009);
nor NOR4 (N9466, N9457, N5557, N4129, N3364);
buf BUF1 (N9467, N9445);
nor NOR2 (N9468, N9459, N222);
and AND2 (N9469, N9462, N727);
nand NAND3 (N9470, N9458, N8726, N760);
buf BUF1 (N9471, N9466);
nand NAND2 (N9472, N9465, N6611);
xor XOR2 (N9473, N9454, N2062);
and AND2 (N9474, N9463, N2335);
not NOT1 (N9475, N9471);
xor XOR2 (N9476, N9473, N1330);
and AND3 (N9477, N9456, N1476, N4399);
xor XOR2 (N9478, N9475, N3014);
nand NAND3 (N9479, N9467, N3353, N4181);
nor NOR2 (N9480, N9477, N585);
xor XOR2 (N9481, N9479, N6722);
and AND3 (N9482, N9476, N5930, N4835);
or OR4 (N9483, N9481, N5267, N1249, N6481);
buf BUF1 (N9484, N9482);
nor NOR4 (N9485, N9483, N4031, N7949, N6252);
and AND3 (N9486, N9484, N3713, N8074);
not NOT1 (N9487, N9468);
nand NAND2 (N9488, N9486, N4095);
buf BUF1 (N9489, N9487);
not NOT1 (N9490, N9464);
buf BUF1 (N9491, N9474);
xor XOR2 (N9492, N9469, N326);
not NOT1 (N9493, N9492);
nand NAND2 (N9494, N9489, N32);
nand NAND3 (N9495, N9478, N689, N3079);
nand NAND2 (N9496, N9493, N2735);
xor XOR2 (N9497, N9491, N8801);
nor NOR2 (N9498, N9470, N250);
or OR3 (N9499, N9494, N1287, N3032);
nand NAND4 (N9500, N9485, N3120, N5036, N379);
nor NOR2 (N9501, N9500, N8080);
nor NOR4 (N9502, N9480, N3334, N7418, N8336);
buf BUF1 (N9503, N9498);
nand NAND4 (N9504, N9503, N6029, N8728, N7505);
buf BUF1 (N9505, N9497);
or OR2 (N9506, N9490, N6854);
buf BUF1 (N9507, N9488);
and AND3 (N9508, N9504, N3362, N5199);
nand NAND2 (N9509, N9472, N8581);
buf BUF1 (N9510, N9508);
and AND3 (N9511, N9499, N3301, N3602);
nor NOR2 (N9512, N9505, N2741);
xor XOR2 (N9513, N9511, N9315);
not NOT1 (N9514, N9509);
nor NOR3 (N9515, N9507, N1962, N5525);
buf BUF1 (N9516, N9512);
not NOT1 (N9517, N9510);
not NOT1 (N9518, N9501);
nand NAND2 (N9519, N9513, N2903);
nor NOR3 (N9520, N9519, N713, N8825);
nand NAND4 (N9521, N9502, N2600, N8920, N9264);
not NOT1 (N9522, N9496);
and AND3 (N9523, N9495, N8607, N5084);
buf BUF1 (N9524, N9517);
buf BUF1 (N9525, N9521);
or OR3 (N9526, N9524, N2084, N9296);
nor NOR2 (N9527, N9515, N4790);
not NOT1 (N9528, N9522);
xor XOR2 (N9529, N9506, N1690);
and AND2 (N9530, N9529, N8198);
and AND3 (N9531, N9528, N9022, N8265);
and AND3 (N9532, N9525, N3615, N872);
or OR4 (N9533, N9516, N4624, N3649, N6391);
not NOT1 (N9534, N9523);
nor NOR2 (N9535, N9530, N6293);
nand NAND2 (N9536, N9527, N7152);
not NOT1 (N9537, N9533);
xor XOR2 (N9538, N9514, N4437);
buf BUF1 (N9539, N9518);
nor NOR2 (N9540, N9539, N9212);
nand NAND4 (N9541, N9538, N7566, N5423, N5408);
nor NOR2 (N9542, N9537, N7109);
xor XOR2 (N9543, N9541, N6515);
not NOT1 (N9544, N9535);
not NOT1 (N9545, N9520);
not NOT1 (N9546, N9542);
nand NAND2 (N9547, N9546, N3390);
nand NAND4 (N9548, N9532, N8256, N6095, N9447);
nand NAND3 (N9549, N9540, N7940, N4739);
buf BUF1 (N9550, N9534);
xor XOR2 (N9551, N9531, N6785);
not NOT1 (N9552, N9548);
and AND4 (N9553, N9536, N538, N419, N3095);
nand NAND4 (N9554, N9553, N1707, N16, N5486);
nor NOR4 (N9555, N9526, N2834, N9106, N3858);
nor NOR3 (N9556, N9551, N3407, N4751);
nand NAND2 (N9557, N9555, N9117);
and AND2 (N9558, N9554, N5092);
and AND4 (N9559, N9549, N1032, N2999, N1633);
or OR2 (N9560, N9559, N1235);
and AND2 (N9561, N9545, N8364);
or OR3 (N9562, N9552, N1398, N8521);
not NOT1 (N9563, N9557);
or OR3 (N9564, N9543, N8829, N8796);
nor NOR4 (N9565, N9544, N4427, N2812, N2988);
nand NAND2 (N9566, N9564, N2396);
or OR4 (N9567, N9563, N991, N6554, N3680);
and AND3 (N9568, N9558, N9116, N2088);
xor XOR2 (N9569, N9560, N9510);
nor NOR2 (N9570, N9562, N9032);
not NOT1 (N9571, N9556);
and AND3 (N9572, N9571, N5546, N5213);
nor NOR2 (N9573, N9569, N7293);
nand NAND4 (N9574, N9566, N176, N3568, N1803);
and AND4 (N9575, N9561, N1027, N9199, N1175);
buf BUF1 (N9576, N9573);
or OR4 (N9577, N9575, N2064, N5918, N8760);
xor XOR2 (N9578, N9570, N1554);
nand NAND2 (N9579, N9578, N2492);
nor NOR4 (N9580, N9574, N6537, N7946, N2707);
buf BUF1 (N9581, N9579);
nand NAND4 (N9582, N9550, N5980, N8054, N751);
and AND4 (N9583, N9581, N7555, N5492, N8317);
not NOT1 (N9584, N9567);
nand NAND4 (N9585, N9580, N6485, N5813, N4892);
or OR3 (N9586, N9576, N5899, N8662);
or OR4 (N9587, N9577, N125, N7999, N8344);
buf BUF1 (N9588, N9568);
nand NAND4 (N9589, N9565, N3362, N1070, N7260);
and AND2 (N9590, N9589, N5605);
nor NOR2 (N9591, N9588, N4590);
nor NOR4 (N9592, N9547, N5939, N4047, N6779);
and AND4 (N9593, N9590, N4142, N2426, N3433);
xor XOR2 (N9594, N9582, N7221);
buf BUF1 (N9595, N9584);
nand NAND4 (N9596, N9593, N6709, N7563, N9114);
and AND4 (N9597, N9596, N6014, N5035, N7052);
buf BUF1 (N9598, N9587);
xor XOR2 (N9599, N9597, N1301);
not NOT1 (N9600, N9585);
or OR2 (N9601, N9583, N3559);
not NOT1 (N9602, N9600);
or OR2 (N9603, N9586, N4007);
not NOT1 (N9604, N9602);
xor XOR2 (N9605, N9572, N6166);
or OR4 (N9606, N9595, N9128, N855, N7444);
xor XOR2 (N9607, N9603, N5854);
nor NOR2 (N9608, N9604, N5630);
nor NOR2 (N9609, N9606, N1686);
not NOT1 (N9610, N9608);
not NOT1 (N9611, N9591);
nor NOR2 (N9612, N9607, N7363);
or OR4 (N9613, N9592, N8130, N477, N6764);
not NOT1 (N9614, N9605);
buf BUF1 (N9615, N9611);
and AND4 (N9616, N9613, N3356, N9450, N938);
buf BUF1 (N9617, N9612);
nand NAND3 (N9618, N9610, N6722, N2509);
xor XOR2 (N9619, N9599, N9077);
not NOT1 (N9620, N9615);
buf BUF1 (N9621, N9609);
nand NAND4 (N9622, N9601, N7734, N1518, N7410);
buf BUF1 (N9623, N9616);
buf BUF1 (N9624, N9623);
buf BUF1 (N9625, N9620);
not NOT1 (N9626, N9619);
and AND2 (N9627, N9626, N4387);
nand NAND4 (N9628, N9621, N2093, N3454, N3081);
not NOT1 (N9629, N9617);
not NOT1 (N9630, N9594);
xor XOR2 (N9631, N9624, N7725);
or OR2 (N9632, N9598, N4460);
or OR4 (N9633, N9630, N4485, N2428, N4510);
or OR2 (N9634, N9627, N8861);
not NOT1 (N9635, N9618);
buf BUF1 (N9636, N9635);
nand NAND4 (N9637, N9625, N9162, N4127, N3473);
nor NOR2 (N9638, N9636, N4231);
nor NOR4 (N9639, N9614, N7228, N8993, N2859);
and AND3 (N9640, N9634, N7326, N1216);
xor XOR2 (N9641, N9628, N1524);
and AND2 (N9642, N9633, N5566);
buf BUF1 (N9643, N9642);
not NOT1 (N9644, N9622);
xor XOR2 (N9645, N9631, N1980);
not NOT1 (N9646, N9641);
not NOT1 (N9647, N9645);
nand NAND3 (N9648, N9647, N2758, N893);
xor XOR2 (N9649, N9639, N2760);
nand NAND3 (N9650, N9648, N7429, N4566);
nor NOR2 (N9651, N9629, N1173);
buf BUF1 (N9652, N9643);
not NOT1 (N9653, N9638);
nor NOR3 (N9654, N9632, N1796, N8278);
buf BUF1 (N9655, N9637);
not NOT1 (N9656, N9654);
or OR2 (N9657, N9649, N5814);
not NOT1 (N9658, N9640);
xor XOR2 (N9659, N9653, N5411);
or OR4 (N9660, N9656, N6511, N6628, N8520);
nand NAND2 (N9661, N9660, N9011);
buf BUF1 (N9662, N9659);
buf BUF1 (N9663, N9650);
nand NAND4 (N9664, N9661, N5091, N6000, N5281);
or OR4 (N9665, N9664, N4688, N2225, N36);
nand NAND2 (N9666, N9657, N1069);
or OR3 (N9667, N9651, N3207, N6893);
or OR3 (N9668, N9663, N5404, N3676);
xor XOR2 (N9669, N9666, N4516);
xor XOR2 (N9670, N9667, N1030);
buf BUF1 (N9671, N9658);
xor XOR2 (N9672, N9662, N9037);
or OR3 (N9673, N9646, N6633, N7613);
and AND3 (N9674, N9671, N7546, N3782);
xor XOR2 (N9675, N9670, N7490);
nand NAND2 (N9676, N9655, N5092);
buf BUF1 (N9677, N9675);
not NOT1 (N9678, N9672);
nand NAND2 (N9679, N9668, N2872);
and AND3 (N9680, N9677, N4394, N2782);
or OR2 (N9681, N9652, N1979);
nand NAND2 (N9682, N9681, N9040);
or OR2 (N9683, N9673, N14);
xor XOR2 (N9684, N9683, N6304);
or OR3 (N9685, N9676, N8870, N6486);
or OR4 (N9686, N9669, N3591, N9417, N8232);
not NOT1 (N9687, N9684);
not NOT1 (N9688, N9680);
not NOT1 (N9689, N9678);
xor XOR2 (N9690, N9644, N9554);
buf BUF1 (N9691, N9687);
not NOT1 (N9692, N9688);
not NOT1 (N9693, N9674);
xor XOR2 (N9694, N9689, N4450);
buf BUF1 (N9695, N9692);
and AND2 (N9696, N9695, N7113);
xor XOR2 (N9697, N9686, N2635);
not NOT1 (N9698, N9690);
not NOT1 (N9699, N9682);
and AND4 (N9700, N9685, N2998, N4825, N4656);
nand NAND4 (N9701, N9696, N3881, N180, N8876);
buf BUF1 (N9702, N9691);
not NOT1 (N9703, N9694);
buf BUF1 (N9704, N9697);
nand NAND2 (N9705, N9699, N8974);
not NOT1 (N9706, N9700);
buf BUF1 (N9707, N9706);
or OR4 (N9708, N9702, N2181, N6159, N7720);
or OR4 (N9709, N9705, N651, N6860, N849);
nand NAND3 (N9710, N9703, N5895, N1571);
nand NAND2 (N9711, N9665, N308);
nand NAND3 (N9712, N9711, N1725, N4020);
xor XOR2 (N9713, N9679, N1705);
nand NAND3 (N9714, N9710, N7610, N342);
and AND4 (N9715, N9712, N9711, N801, N1461);
or OR3 (N9716, N9713, N2667, N7548);
not NOT1 (N9717, N9707);
or OR4 (N9718, N9701, N5357, N3233, N7951);
and AND3 (N9719, N9708, N8426, N8495);
and AND4 (N9720, N9717, N7399, N6189, N7701);
or OR4 (N9721, N9698, N2085, N804, N365);
buf BUF1 (N9722, N9720);
nand NAND2 (N9723, N9709, N792);
nor NOR4 (N9724, N9723, N6494, N3933, N6603);
nor NOR4 (N9725, N9722, N5674, N4742, N6747);
nor NOR2 (N9726, N9714, N7857);
not NOT1 (N9727, N9725);
buf BUF1 (N9728, N9718);
and AND4 (N9729, N9726, N9169, N5404, N7304);
nor NOR2 (N9730, N9716, N891);
and AND4 (N9731, N9728, N2632, N5165, N6196);
xor XOR2 (N9732, N9727, N7754);
nand NAND4 (N9733, N9731, N1366, N8140, N5171);
nand NAND3 (N9734, N9719, N8092, N2610);
buf BUF1 (N9735, N9724);
not NOT1 (N9736, N9733);
nor NOR4 (N9737, N9734, N2323, N3543, N1914);
buf BUF1 (N9738, N9704);
and AND3 (N9739, N9737, N6597, N1042);
nand NAND3 (N9740, N9693, N4872, N2833);
xor XOR2 (N9741, N9730, N9085);
buf BUF1 (N9742, N9732);
xor XOR2 (N9743, N9715, N2422);
nand NAND2 (N9744, N9740, N8354);
buf BUF1 (N9745, N9743);
not NOT1 (N9746, N9745);
buf BUF1 (N9747, N9736);
nor NOR3 (N9748, N9739, N5031, N5505);
nor NOR3 (N9749, N9744, N2201, N356);
not NOT1 (N9750, N9738);
nor NOR2 (N9751, N9729, N7796);
not NOT1 (N9752, N9750);
nand NAND4 (N9753, N9747, N7419, N1442, N2208);
not NOT1 (N9754, N9742);
or OR3 (N9755, N9735, N4748, N4518);
or OR4 (N9756, N9741, N6405, N9502, N2418);
and AND3 (N9757, N9754, N2890, N5050);
not NOT1 (N9758, N9749);
not NOT1 (N9759, N9755);
and AND3 (N9760, N9757, N3691, N3418);
not NOT1 (N9761, N9760);
nor NOR2 (N9762, N9759, N8797);
and AND4 (N9763, N9751, N2710, N987, N1947);
not NOT1 (N9764, N9763);
nand NAND4 (N9765, N9758, N119, N7229, N8124);
nand NAND2 (N9766, N9748, N386);
or OR4 (N9767, N9761, N4883, N6830, N8306);
buf BUF1 (N9768, N9766);
or OR4 (N9769, N9764, N4304, N4137, N3969);
or OR3 (N9770, N9769, N8826, N6759);
buf BUF1 (N9771, N9753);
xor XOR2 (N9772, N9762, N204);
not NOT1 (N9773, N9721);
and AND4 (N9774, N9767, N6540, N520, N3909);
buf BUF1 (N9775, N9770);
and AND4 (N9776, N9772, N3490, N5930, N7986);
or OR2 (N9777, N9771, N4795);
nor NOR4 (N9778, N9765, N3738, N3172, N4344);
nor NOR4 (N9779, N9776, N1928, N3700, N8608);
nor NOR4 (N9780, N9768, N1517, N2682, N8322);
and AND4 (N9781, N9780, N5431, N4038, N6700);
nand NAND2 (N9782, N9752, N251);
not NOT1 (N9783, N9774);
nand NAND2 (N9784, N9783, N4977);
not NOT1 (N9785, N9756);
or OR4 (N9786, N9784, N7642, N9584, N5519);
and AND4 (N9787, N9786, N180, N2473, N366);
and AND4 (N9788, N9777, N9070, N4452, N5321);
buf BUF1 (N9789, N9787);
or OR2 (N9790, N9781, N3435);
not NOT1 (N9791, N9785);
and AND4 (N9792, N9779, N4952, N2118, N3890);
xor XOR2 (N9793, N9775, N3443);
xor XOR2 (N9794, N9792, N5278);
buf BUF1 (N9795, N9790);
and AND4 (N9796, N9794, N6822, N3605, N8257);
nand NAND4 (N9797, N9791, N8774, N7351, N3607);
buf BUF1 (N9798, N9795);
nand NAND2 (N9799, N9782, N2626);
not NOT1 (N9800, N9796);
or OR3 (N9801, N9773, N9751, N3102);
or OR2 (N9802, N9778, N8007);
or OR4 (N9803, N9788, N4150, N1714, N1553);
and AND4 (N9804, N9797, N6901, N7031, N8431);
or OR2 (N9805, N9746, N4198);
buf BUF1 (N9806, N9803);
nand NAND2 (N9807, N9802, N3859);
and AND2 (N9808, N9789, N6724);
or OR4 (N9809, N9793, N3369, N3779, N8265);
not NOT1 (N9810, N9808);
and AND3 (N9811, N9807, N5015, N9803);
nor NOR2 (N9812, N9800, N5958);
or OR3 (N9813, N9811, N2173, N4274);
and AND4 (N9814, N9812, N8405, N8079, N6212);
not NOT1 (N9815, N9809);
xor XOR2 (N9816, N9801, N4480);
xor XOR2 (N9817, N9799, N9742);
not NOT1 (N9818, N9805);
xor XOR2 (N9819, N9806, N7300);
nor NOR3 (N9820, N9816, N4449, N1554);
not NOT1 (N9821, N9820);
nand NAND3 (N9822, N9815, N3468, N8612);
nand NAND2 (N9823, N9814, N854);
and AND2 (N9824, N9813, N4445);
xor XOR2 (N9825, N9824, N6612);
nor NOR4 (N9826, N9819, N3948, N8483, N4348);
not NOT1 (N9827, N9818);
xor XOR2 (N9828, N9798, N3779);
nor NOR4 (N9829, N9822, N4562, N586, N1700);
or OR3 (N9830, N9827, N2767, N7213);
nand NAND4 (N9831, N9828, N2067, N683, N4463);
and AND2 (N9832, N9817, N8944);
xor XOR2 (N9833, N9825, N6884);
buf BUF1 (N9834, N9831);
xor XOR2 (N9835, N9823, N2240);
nand NAND4 (N9836, N9835, N383, N7785, N1874);
buf BUF1 (N9837, N9833);
xor XOR2 (N9838, N9830, N7914);
not NOT1 (N9839, N9834);
not NOT1 (N9840, N9837);
xor XOR2 (N9841, N9838, N9437);
xor XOR2 (N9842, N9810, N3459);
xor XOR2 (N9843, N9826, N4677);
nor NOR3 (N9844, N9832, N8279, N3418);
not NOT1 (N9845, N9840);
nand NAND2 (N9846, N9843, N3930);
nand NAND4 (N9847, N9836, N3696, N5984, N1831);
not NOT1 (N9848, N9842);
and AND2 (N9849, N9846, N223);
xor XOR2 (N9850, N9845, N6388);
not NOT1 (N9851, N9841);
nor NOR3 (N9852, N9829, N3566, N4958);
not NOT1 (N9853, N9821);
xor XOR2 (N9854, N9844, N6354);
not NOT1 (N9855, N9849);
nor NOR4 (N9856, N9847, N4256, N9039, N2359);
xor XOR2 (N9857, N9848, N8593);
nor NOR4 (N9858, N9804, N860, N9242, N8871);
or OR2 (N9859, N9858, N7806);
xor XOR2 (N9860, N9857, N7931);
buf BUF1 (N9861, N9851);
not NOT1 (N9862, N9859);
xor XOR2 (N9863, N9839, N2578);
nand NAND4 (N9864, N9854, N3587, N3361, N4623);
not NOT1 (N9865, N9853);
nand NAND2 (N9866, N9861, N2512);
and AND4 (N9867, N9863, N1515, N6689, N7740);
nor NOR3 (N9868, N9865, N4399, N3714);
or OR3 (N9869, N9866, N8701, N4700);
nand NAND2 (N9870, N9856, N9669);
or OR4 (N9871, N9850, N8958, N7922, N8903);
and AND2 (N9872, N9860, N8921);
nand NAND4 (N9873, N9867, N2641, N7408, N2511);
or OR3 (N9874, N9864, N1396, N109);
not NOT1 (N9875, N9868);
xor XOR2 (N9876, N9875, N3515);
nand NAND4 (N9877, N9874, N8827, N4005, N3023);
xor XOR2 (N9878, N9852, N9624);
not NOT1 (N9879, N9862);
or OR3 (N9880, N9870, N4074, N6777);
xor XOR2 (N9881, N9855, N7661);
buf BUF1 (N9882, N9871);
and AND4 (N9883, N9876, N8869, N5121, N4445);
nand NAND3 (N9884, N9881, N3128, N612);
nand NAND3 (N9885, N9879, N6580, N43);
nor NOR2 (N9886, N9884, N7619);
xor XOR2 (N9887, N9886, N5408);
nand NAND3 (N9888, N9873, N3761, N2349);
nor NOR3 (N9889, N9888, N1219, N7866);
or OR4 (N9890, N9885, N8763, N9182, N5197);
and AND3 (N9891, N9877, N1341, N1977);
xor XOR2 (N9892, N9869, N6853);
nand NAND3 (N9893, N9889, N1451, N2864);
or OR2 (N9894, N9891, N4982);
xor XOR2 (N9895, N9882, N261);
nor NOR3 (N9896, N9880, N5730, N2806);
nand NAND3 (N9897, N9878, N5311, N4090);
and AND3 (N9898, N9872, N3172, N6337);
nand NAND4 (N9899, N9887, N1953, N2309, N4018);
and AND3 (N9900, N9890, N2722, N6831);
or OR3 (N9901, N9883, N763, N5503);
nand NAND2 (N9902, N9899, N641);
or OR4 (N9903, N9896, N5553, N4891, N6620);
nor NOR2 (N9904, N9895, N1648);
not NOT1 (N9905, N9897);
and AND4 (N9906, N9900, N2027, N2038, N2657);
and AND3 (N9907, N9898, N6808, N634);
and AND2 (N9908, N9904, N7411);
not NOT1 (N9909, N9892);
and AND3 (N9910, N9893, N7892, N3862);
or OR4 (N9911, N9908, N5463, N5679, N8118);
buf BUF1 (N9912, N9907);
or OR4 (N9913, N9905, N9069, N668, N775);
nor NOR4 (N9914, N9911, N8303, N3403, N4567);
nor NOR2 (N9915, N9901, N3395);
nor NOR4 (N9916, N9894, N7492, N4498, N3535);
or OR4 (N9917, N9909, N443, N6666, N3234);
and AND2 (N9918, N9912, N6620);
and AND3 (N9919, N9913, N1594, N2101);
and AND4 (N9920, N9918, N1355, N7338, N4682);
xor XOR2 (N9921, N9919, N6084);
buf BUF1 (N9922, N9906);
not NOT1 (N9923, N9903);
nor NOR2 (N9924, N9917, N360);
nand NAND4 (N9925, N9921, N832, N4583, N4711);
not NOT1 (N9926, N9920);
or OR2 (N9927, N9925, N7987);
or OR4 (N9928, N9902, N1893, N9464, N101);
and AND2 (N9929, N9915, N8751);
nand NAND3 (N9930, N9916, N191, N522);
and AND4 (N9931, N9928, N9299, N3100, N1738);
or OR2 (N9932, N9926, N6002);
and AND2 (N9933, N9923, N1239);
and AND3 (N9934, N9910, N5594, N7206);
nand NAND3 (N9935, N9934, N231, N964);
nor NOR4 (N9936, N9929, N6162, N7451, N349);
xor XOR2 (N9937, N9914, N4124);
and AND2 (N9938, N9933, N5097);
not NOT1 (N9939, N9922);
nor NOR3 (N9940, N9927, N4080, N2972);
or OR2 (N9941, N9935, N6465);
xor XOR2 (N9942, N9938, N8203);
or OR2 (N9943, N9931, N5857);
and AND3 (N9944, N9924, N1011, N754);
and AND4 (N9945, N9941, N7610, N9639, N3837);
or OR3 (N9946, N9945, N2982, N1805);
not NOT1 (N9947, N9939);
nand NAND2 (N9948, N9936, N1091);
nor NOR3 (N9949, N9946, N375, N8530);
nor NOR2 (N9950, N9942, N6391);
not NOT1 (N9951, N9940);
not NOT1 (N9952, N9949);
xor XOR2 (N9953, N9944, N4898);
or OR4 (N9954, N9937, N1297, N6694, N4983);
nand NAND3 (N9955, N9947, N1126, N9828);
not NOT1 (N9956, N9943);
xor XOR2 (N9957, N9951, N7814);
and AND3 (N9958, N9932, N9608, N9258);
buf BUF1 (N9959, N9956);
nand NAND3 (N9960, N9950, N3373, N8595);
not NOT1 (N9961, N9953);
or OR3 (N9962, N9960, N9399, N8143);
nand NAND3 (N9963, N9959, N4999, N7936);
xor XOR2 (N9964, N9957, N6957);
and AND2 (N9965, N9948, N5816);
and AND3 (N9966, N9962, N8857, N8866);
nor NOR3 (N9967, N9961, N8296, N9326);
buf BUF1 (N9968, N9965);
buf BUF1 (N9969, N9968);
or OR4 (N9970, N9963, N5325, N6364, N1059);
not NOT1 (N9971, N9952);
or OR3 (N9972, N9970, N255, N4068);
or OR3 (N9973, N9930, N7440, N1535);
xor XOR2 (N9974, N9973, N777);
not NOT1 (N9975, N9966);
nand NAND2 (N9976, N9954, N3288);
nor NOR2 (N9977, N9955, N4013);
buf BUF1 (N9978, N9967);
buf BUF1 (N9979, N9974);
not NOT1 (N9980, N9972);
nand NAND4 (N9981, N9977, N8494, N1446, N7810);
nor NOR2 (N9982, N9979, N333);
xor XOR2 (N9983, N9980, N9111);
nor NOR2 (N9984, N9971, N7503);
not NOT1 (N9985, N9964);
and AND4 (N9986, N9982, N8973, N9194, N7496);
nor NOR3 (N9987, N9983, N7486, N7240);
nand NAND3 (N9988, N9978, N1214, N8236);
nor NOR2 (N9989, N9985, N1717);
not NOT1 (N9990, N9958);
nand NAND4 (N9991, N9984, N2624, N989, N5661);
xor XOR2 (N9992, N9981, N2612);
nor NOR2 (N9993, N9975, N5312);
not NOT1 (N9994, N9990);
nor NOR4 (N9995, N9991, N5046, N4020, N4200);
xor XOR2 (N9996, N9976, N7811);
not NOT1 (N9997, N9988);
xor XOR2 (N9998, N9987, N8782);
and AND4 (N9999, N9969, N3601, N1888, N1175);
not NOT1 (N10000, N9999);
not NOT1 (N10001, N9992);
not NOT1 (N10002, N9996);
nor NOR3 (N10003, N9989, N4591, N8784);
xor XOR2 (N10004, N10000, N615);
nand NAND3 (N10005, N9997, N4976, N1571);
buf BUF1 (N10006, N10001);
and AND4 (N10007, N10006, N8424, N7138, N8617);
xor XOR2 (N10008, N10005, N2380);
nand NAND2 (N10009, N10008, N9292);
nand NAND3 (N10010, N10003, N4100, N4914);
xor XOR2 (N10011, N9994, N1405);
not NOT1 (N10012, N10007);
buf BUF1 (N10013, N10009);
buf BUF1 (N10014, N10004);
nand NAND4 (N10015, N9993, N9121, N8465, N7138);
xor XOR2 (N10016, N10013, N9944);
xor XOR2 (N10017, N10012, N6341);
nor NOR4 (N10018, N10015, N2927, N8215, N7679);
buf BUF1 (N10019, N10010);
and AND3 (N10020, N10014, N6620, N1227);
xor XOR2 (N10021, N9986, N924);
buf BUF1 (N10022, N10021);
not NOT1 (N10023, N9995);
nor NOR2 (N10024, N10020, N128);
and AND4 (N10025, N10024, N3777, N829, N6320);
nor NOR4 (N10026, N9998, N4388, N150, N4434);
xor XOR2 (N10027, N10026, N334);
or OR3 (N10028, N10027, N2825, N2661);
xor XOR2 (N10029, N10022, N980);
or OR2 (N10030, N10029, N2655);
or OR4 (N10031, N10028, N1241, N5145, N4045);
not NOT1 (N10032, N10017);
or OR4 (N10033, N10025, N2262, N3153, N2652);
nand NAND4 (N10034, N10011, N7241, N6877, N1594);
or OR2 (N10035, N10031, N951);
not NOT1 (N10036, N10034);
buf BUF1 (N10037, N10023);
or OR2 (N10038, N10016, N2706);
nor NOR2 (N10039, N10035, N409);
buf BUF1 (N10040, N10038);
nand NAND2 (N10041, N10037, N963);
not NOT1 (N10042, N10002);
or OR2 (N10043, N10041, N3355);
not NOT1 (N10044, N10042);
nand NAND4 (N10045, N10018, N9046, N2261, N5655);
or OR4 (N10046, N10030, N6168, N2788, N4239);
nor NOR4 (N10047, N10044, N9900, N7457, N2126);
xor XOR2 (N10048, N10045, N5228);
nor NOR3 (N10049, N10047, N7802, N1074);
nand NAND3 (N10050, N10019, N1866, N9801);
nand NAND4 (N10051, N10039, N5828, N8452, N5391);
xor XOR2 (N10052, N10046, N7659);
buf BUF1 (N10053, N10043);
or OR2 (N10054, N10050, N5350);
nor NOR3 (N10055, N10054, N2823, N853);
xor XOR2 (N10056, N10052, N10030);
not NOT1 (N10057, N10055);
and AND2 (N10058, N10036, N2966);
or OR3 (N10059, N10048, N6505, N7462);
nor NOR2 (N10060, N10053, N8169);
xor XOR2 (N10061, N10056, N6142);
nor NOR2 (N10062, N10061, N1529);
nor NOR2 (N10063, N10062, N6879);
nand NAND3 (N10064, N10063, N4364, N4512);
xor XOR2 (N10065, N10057, N3472);
and AND4 (N10066, N10033, N8957, N5824, N4095);
xor XOR2 (N10067, N10051, N8653);
xor XOR2 (N10068, N10064, N9637);
nand NAND3 (N10069, N10040, N2966, N5321);
buf BUF1 (N10070, N10059);
buf BUF1 (N10071, N10070);
or OR3 (N10072, N10069, N9429, N1554);
not NOT1 (N10073, N10058);
or OR4 (N10074, N10066, N4116, N8609, N59);
and AND4 (N10075, N10065, N1885, N6554, N4155);
and AND3 (N10076, N10073, N3854, N6503);
buf BUF1 (N10077, N10076);
buf BUF1 (N10078, N10072);
not NOT1 (N10079, N10049);
xor XOR2 (N10080, N10071, N4292);
or OR4 (N10081, N10075, N8784, N7933, N4575);
nand NAND2 (N10082, N10077, N8086);
or OR3 (N10083, N10067, N4581, N5277);
buf BUF1 (N10084, N10080);
and AND4 (N10085, N10081, N8587, N3770, N2053);
nor NOR4 (N10086, N10084, N856, N5387, N9134);
not NOT1 (N10087, N10079);
and AND2 (N10088, N10074, N7161);
not NOT1 (N10089, N10088);
or OR3 (N10090, N10083, N1679, N221);
and AND3 (N10091, N10078, N333, N655);
nor NOR4 (N10092, N10060, N2097, N5449, N3730);
not NOT1 (N10093, N10087);
not NOT1 (N10094, N10086);
and AND4 (N10095, N10092, N698, N6034, N9514);
xor XOR2 (N10096, N10068, N2063);
nor NOR3 (N10097, N10096, N6099, N3717);
nand NAND2 (N10098, N10094, N4441);
not NOT1 (N10099, N10093);
xor XOR2 (N10100, N10098, N2198);
nor NOR3 (N10101, N10100, N9944, N6532);
not NOT1 (N10102, N10090);
buf BUF1 (N10103, N10102);
nor NOR3 (N10104, N10082, N3856, N4626);
xor XOR2 (N10105, N10099, N8731);
nor NOR3 (N10106, N10032, N563, N5349);
buf BUF1 (N10107, N10097);
and AND2 (N10108, N10095, N5347);
not NOT1 (N10109, N10106);
nor NOR3 (N10110, N10089, N6321, N6678);
not NOT1 (N10111, N10105);
not NOT1 (N10112, N10104);
nor NOR2 (N10113, N10101, N9233);
or OR2 (N10114, N10113, N5610);
nor NOR4 (N10115, N10109, N5659, N664, N1299);
xor XOR2 (N10116, N10108, N321);
or OR4 (N10117, N10112, N4576, N10104, N7466);
or OR3 (N10118, N10107, N4487, N9110);
not NOT1 (N10119, N10114);
nand NAND3 (N10120, N10119, N8782, N3357);
nand NAND4 (N10121, N10120, N8344, N741, N6060);
nand NAND2 (N10122, N10110, N873);
and AND2 (N10123, N10085, N9212);
nor NOR4 (N10124, N10118, N96, N3391, N5148);
nand NAND2 (N10125, N10117, N3458);
xor XOR2 (N10126, N10121, N1279);
nor NOR3 (N10127, N10111, N2883, N9103);
xor XOR2 (N10128, N10127, N7441);
not NOT1 (N10129, N10128);
or OR4 (N10130, N10091, N5237, N292, N5123);
and AND2 (N10131, N10129, N4194);
xor XOR2 (N10132, N10126, N4964);
and AND4 (N10133, N10132, N9500, N9459, N9669);
or OR3 (N10134, N10131, N937, N4183);
or OR2 (N10135, N10115, N1157);
buf BUF1 (N10136, N10125);
nand NAND4 (N10137, N10122, N3341, N6243, N2289);
nand NAND3 (N10138, N10130, N7224, N8330);
and AND2 (N10139, N10116, N927);
nor NOR4 (N10140, N10133, N10032, N2421, N3450);
xor XOR2 (N10141, N10140, N6002);
nand NAND3 (N10142, N10138, N835, N35);
nor NOR3 (N10143, N10135, N3293, N2624);
nand NAND4 (N10144, N10134, N1672, N9371, N2763);
buf BUF1 (N10145, N10141);
nand NAND2 (N10146, N10144, N2748);
nor NOR2 (N10147, N10123, N5543);
xor XOR2 (N10148, N10139, N6092);
not NOT1 (N10149, N10137);
nor NOR4 (N10150, N10149, N3215, N8502, N8645);
buf BUF1 (N10151, N10124);
not NOT1 (N10152, N10145);
nor NOR4 (N10153, N10136, N337, N2447, N8551);
nand NAND4 (N10154, N10103, N6434, N3272, N6029);
xor XOR2 (N10155, N10152, N4273);
buf BUF1 (N10156, N10143);
buf BUF1 (N10157, N10153);
xor XOR2 (N10158, N10151, N3013);
not NOT1 (N10159, N10154);
xor XOR2 (N10160, N10155, N9182);
xor XOR2 (N10161, N10158, N8265);
and AND3 (N10162, N10148, N7143, N1275);
or OR2 (N10163, N10157, N5648);
xor XOR2 (N10164, N10150, N8921);
or OR2 (N10165, N10162, N6589);
and AND4 (N10166, N10163, N9027, N3184, N4804);
xor XOR2 (N10167, N10165, N3201);
and AND4 (N10168, N10159, N5304, N980, N653);
nor NOR4 (N10169, N10168, N7811, N5216, N3411);
not NOT1 (N10170, N10167);
not NOT1 (N10171, N10160);
buf BUF1 (N10172, N10142);
xor XOR2 (N10173, N10161, N6219);
and AND2 (N10174, N10164, N2859);
xor XOR2 (N10175, N10166, N2373);
and AND2 (N10176, N10146, N2385);
and AND4 (N10177, N10175, N600, N7367, N2465);
buf BUF1 (N10178, N10169);
not NOT1 (N10179, N10177);
buf BUF1 (N10180, N10172);
and AND4 (N10181, N10180, N3824, N5806, N1219);
and AND2 (N10182, N10171, N4344);
nand NAND3 (N10183, N10179, N8453, N1346);
nand NAND4 (N10184, N10173, N8223, N6790, N9640);
nand NAND2 (N10185, N10184, N7415);
or OR2 (N10186, N10185, N1286);
xor XOR2 (N10187, N10170, N7083);
not NOT1 (N10188, N10181);
xor XOR2 (N10189, N10178, N9415);
nand NAND2 (N10190, N10176, N35);
and AND4 (N10191, N10174, N9742, N6948, N9399);
xor XOR2 (N10192, N10182, N6003);
or OR3 (N10193, N10190, N195, N55);
xor XOR2 (N10194, N10187, N6049);
not NOT1 (N10195, N10188);
not NOT1 (N10196, N10193);
or OR3 (N10197, N10189, N5656, N3930);
nor NOR4 (N10198, N10194, N9349, N6887, N97);
xor XOR2 (N10199, N10197, N8180);
not NOT1 (N10200, N10156);
xor XOR2 (N10201, N10200, N4319);
nor NOR3 (N10202, N10198, N6475, N8379);
not NOT1 (N10203, N10192);
xor XOR2 (N10204, N10202, N6296);
nor NOR3 (N10205, N10186, N3104, N3398);
not NOT1 (N10206, N10199);
and AND2 (N10207, N10196, N1178);
or OR3 (N10208, N10183, N8695, N1402);
nor NOR4 (N10209, N10204, N7028, N6526, N4651);
buf BUF1 (N10210, N10191);
nor NOR2 (N10211, N10207, N1796);
or OR2 (N10212, N10147, N9370);
and AND4 (N10213, N10203, N8874, N5988, N2309);
or OR3 (N10214, N10211, N4434, N4523);
buf BUF1 (N10215, N10213);
or OR2 (N10216, N10212, N6692);
xor XOR2 (N10217, N10214, N10043);
xor XOR2 (N10218, N10195, N1500);
nor NOR4 (N10219, N10209, N1926, N3450, N8257);
xor XOR2 (N10220, N10216, N587);
or OR3 (N10221, N10219, N587, N9900);
or OR2 (N10222, N10220, N7999);
xor XOR2 (N10223, N10218, N2999);
not NOT1 (N10224, N10215);
xor XOR2 (N10225, N10224, N1102);
and AND3 (N10226, N10221, N256, N8167);
buf BUF1 (N10227, N10206);
xor XOR2 (N10228, N10223, N5556);
and AND4 (N10229, N10225, N3022, N7632, N2683);
nor NOR4 (N10230, N10222, N1413, N6706, N8816);
not NOT1 (N10231, N10228);
or OR4 (N10232, N10210, N6584, N2816, N4464);
nand NAND2 (N10233, N10229, N9319);
buf BUF1 (N10234, N10230);
buf BUF1 (N10235, N10234);
or OR2 (N10236, N10217, N5458);
and AND2 (N10237, N10201, N8140);
and AND3 (N10238, N10232, N3070, N3975);
buf BUF1 (N10239, N10231);
not NOT1 (N10240, N10205);
xor XOR2 (N10241, N10233, N2592);
nor NOR2 (N10242, N10208, N2276);
or OR2 (N10243, N10227, N850);
nand NAND2 (N10244, N10239, N3076);
or OR3 (N10245, N10226, N2704, N3797);
buf BUF1 (N10246, N10243);
or OR2 (N10247, N10244, N9853);
xor XOR2 (N10248, N10235, N9864);
or OR3 (N10249, N10242, N7217, N4215);
not NOT1 (N10250, N10237);
buf BUF1 (N10251, N10238);
xor XOR2 (N10252, N10247, N1848);
buf BUF1 (N10253, N10245);
xor XOR2 (N10254, N10252, N8852);
and AND2 (N10255, N10236, N7756);
nor NOR3 (N10256, N10255, N4391, N1662);
and AND2 (N10257, N10246, N4830);
or OR3 (N10258, N10253, N3509, N8868);
not NOT1 (N10259, N10254);
nor NOR3 (N10260, N10257, N1941, N1418);
not NOT1 (N10261, N10250);
or OR3 (N10262, N10241, N4838, N2328);
or OR2 (N10263, N10249, N5501);
buf BUF1 (N10264, N10256);
nand NAND2 (N10265, N10261, N8361);
or OR2 (N10266, N10248, N1750);
nand NAND4 (N10267, N10251, N7853, N585, N5639);
nor NOR4 (N10268, N10258, N3032, N9204, N8054);
nand NAND4 (N10269, N10267, N8593, N7753, N5863);
nand NAND3 (N10270, N10265, N6859, N1957);
or OR2 (N10271, N10266, N698);
xor XOR2 (N10272, N10269, N4063);
buf BUF1 (N10273, N10263);
xor XOR2 (N10274, N10268, N7074);
nand NAND4 (N10275, N10271, N5639, N1476, N6867);
nor NOR4 (N10276, N10274, N8334, N7143, N380);
not NOT1 (N10277, N10259);
xor XOR2 (N10278, N10273, N9172);
nor NOR2 (N10279, N10270, N7531);
nor NOR2 (N10280, N10277, N7501);
not NOT1 (N10281, N10272);
nand NAND2 (N10282, N10278, N1405);
not NOT1 (N10283, N10279);
buf BUF1 (N10284, N10283);
or OR2 (N10285, N10280, N2081);
buf BUF1 (N10286, N10275);
and AND2 (N10287, N10284, N1137);
nor NOR2 (N10288, N10286, N715);
buf BUF1 (N10289, N10282);
nor NOR2 (N10290, N10288, N4645);
not NOT1 (N10291, N10281);
buf BUF1 (N10292, N10291);
nor NOR2 (N10293, N10240, N5426);
or OR3 (N10294, N10290, N271, N7720);
nand NAND4 (N10295, N10276, N135, N3850, N887);
buf BUF1 (N10296, N10294);
buf BUF1 (N10297, N10260);
not NOT1 (N10298, N10297);
buf BUF1 (N10299, N10262);
buf BUF1 (N10300, N10292);
or OR2 (N10301, N10285, N4139);
nand NAND3 (N10302, N10299, N6679, N4829);
or OR2 (N10303, N10289, N1434);
and AND4 (N10304, N10302, N9455, N3957, N3569);
or OR4 (N10305, N10287, N9391, N1632, N4112);
or OR2 (N10306, N10296, N825);
xor XOR2 (N10307, N10301, N469);
nand NAND3 (N10308, N10306, N2226, N4078);
or OR3 (N10309, N10293, N2384, N4445);
or OR2 (N10310, N10308, N7264);
nor NOR2 (N10311, N10300, N1710);
nand NAND2 (N10312, N10310, N9692);
nand NAND2 (N10313, N10311, N4244);
or OR4 (N10314, N10307, N9078, N7283, N6653);
buf BUF1 (N10315, N10312);
xor XOR2 (N10316, N10303, N6134);
not NOT1 (N10317, N10316);
xor XOR2 (N10318, N10313, N4897);
or OR2 (N10319, N10264, N5432);
not NOT1 (N10320, N10314);
and AND4 (N10321, N10309, N8378, N2532, N6385);
nand NAND2 (N10322, N10318, N7291);
xor XOR2 (N10323, N10320, N305);
nand NAND2 (N10324, N10319, N4988);
buf BUF1 (N10325, N10295);
buf BUF1 (N10326, N10304);
and AND4 (N10327, N10305, N5837, N83, N6571);
and AND2 (N10328, N10322, N1934);
nor NOR2 (N10329, N10324, N8730);
nor NOR3 (N10330, N10321, N9125, N4560);
xor XOR2 (N10331, N10327, N4154);
not NOT1 (N10332, N10331);
or OR3 (N10333, N10330, N7684, N9289);
nor NOR3 (N10334, N10333, N8635, N2356);
not NOT1 (N10335, N10298);
or OR2 (N10336, N10334, N4314);
and AND4 (N10337, N10326, N9781, N4628, N4024);
or OR3 (N10338, N10336, N4614, N2495);
buf BUF1 (N10339, N10335);
xor XOR2 (N10340, N10315, N9412);
nand NAND4 (N10341, N10328, N7555, N6222, N9824);
nand NAND3 (N10342, N10337, N2941, N3760);
and AND2 (N10343, N10329, N944);
or OR2 (N10344, N10338, N6996);
or OR4 (N10345, N10325, N9514, N6032, N5397);
nor NOR3 (N10346, N10332, N9852, N3536);
and AND4 (N10347, N10341, N3536, N8763, N9466);
xor XOR2 (N10348, N10346, N8422);
nor NOR2 (N10349, N10344, N10205);
not NOT1 (N10350, N10342);
nor NOR4 (N10351, N10343, N9381, N6639, N3660);
buf BUF1 (N10352, N10350);
nand NAND2 (N10353, N10317, N155);
xor XOR2 (N10354, N10345, N8372);
nor NOR4 (N10355, N10348, N8003, N8828, N4154);
not NOT1 (N10356, N10355);
nand NAND4 (N10357, N10354, N8457, N5338, N2436);
xor XOR2 (N10358, N10351, N8089);
nor NOR4 (N10359, N10339, N2986, N2143, N2504);
or OR4 (N10360, N10352, N1124, N6890, N4786);
xor XOR2 (N10361, N10323, N9700);
nor NOR4 (N10362, N10359, N2480, N5149, N334);
and AND4 (N10363, N10347, N7632, N3126, N2799);
not NOT1 (N10364, N10358);
xor XOR2 (N10365, N10357, N8162);
not NOT1 (N10366, N10363);
xor XOR2 (N10367, N10353, N8635);
nand NAND2 (N10368, N10367, N4714);
not NOT1 (N10369, N10340);
nor NOR3 (N10370, N10366, N9202, N5480);
and AND4 (N10371, N10361, N1998, N7586, N2158);
xor XOR2 (N10372, N10360, N6059);
buf BUF1 (N10373, N10370);
not NOT1 (N10374, N10362);
nor NOR3 (N10375, N10365, N7771, N9519);
or OR4 (N10376, N10374, N1559, N5657, N4058);
not NOT1 (N10377, N10369);
nand NAND3 (N10378, N10364, N9070, N6126);
not NOT1 (N10379, N10378);
xor XOR2 (N10380, N10372, N6803);
and AND3 (N10381, N10349, N4677, N10316);
and AND4 (N10382, N10377, N2409, N7503, N7448);
not NOT1 (N10383, N10379);
nor NOR4 (N10384, N10375, N8480, N8044, N5332);
xor XOR2 (N10385, N10380, N144);
and AND4 (N10386, N10371, N10183, N10258, N6390);
nor NOR4 (N10387, N10356, N1897, N1428, N4833);
nand NAND3 (N10388, N10384, N9683, N152);
nor NOR2 (N10389, N10381, N8223);
xor XOR2 (N10390, N10386, N8556);
and AND3 (N10391, N10383, N7888, N900);
or OR4 (N10392, N10385, N7514, N3077, N1731);
buf BUF1 (N10393, N10391);
and AND4 (N10394, N10387, N4862, N9570, N371);
xor XOR2 (N10395, N10382, N6072);
buf BUF1 (N10396, N10390);
nor NOR2 (N10397, N10392, N5677);
or OR4 (N10398, N10368, N6584, N6602, N2646);
or OR3 (N10399, N10396, N5861, N5440);
nand NAND4 (N10400, N10394, N4705, N1563, N8074);
nand NAND2 (N10401, N10389, N8558);
nor NOR3 (N10402, N10400, N6604, N8559);
buf BUF1 (N10403, N10373);
xor XOR2 (N10404, N10388, N2057);
not NOT1 (N10405, N10393);
not NOT1 (N10406, N10404);
buf BUF1 (N10407, N10376);
not NOT1 (N10408, N10405);
nand NAND4 (N10409, N10401, N4766, N5996, N1525);
or OR3 (N10410, N10397, N3778, N5459);
buf BUF1 (N10411, N10408);
not NOT1 (N10412, N10406);
nor NOR4 (N10413, N10410, N9594, N9465, N1214);
not NOT1 (N10414, N10409);
not NOT1 (N10415, N10413);
and AND2 (N10416, N10415, N8755);
or OR2 (N10417, N10395, N7600);
buf BUF1 (N10418, N10407);
buf BUF1 (N10419, N10399);
or OR4 (N10420, N10414, N4086, N57, N3200);
not NOT1 (N10421, N10412);
buf BUF1 (N10422, N10421);
not NOT1 (N10423, N10398);
nor NOR3 (N10424, N10411, N1059, N152);
nand NAND4 (N10425, N10402, N1410, N4674, N5485);
or OR3 (N10426, N10417, N7758, N8953);
not NOT1 (N10427, N10419);
nor NOR2 (N10428, N10424, N5761);
nor NOR3 (N10429, N10403, N3103, N4616);
xor XOR2 (N10430, N10420, N9784);
and AND3 (N10431, N10422, N6919, N7207);
xor XOR2 (N10432, N10429, N6121);
xor XOR2 (N10433, N10416, N1256);
nor NOR2 (N10434, N10430, N3934);
xor XOR2 (N10435, N10428, N5151);
or OR3 (N10436, N10427, N2287, N917);
not NOT1 (N10437, N10425);
not NOT1 (N10438, N10431);
buf BUF1 (N10439, N10438);
xor XOR2 (N10440, N10436, N8901);
nor NOR3 (N10441, N10433, N9302, N6160);
not NOT1 (N10442, N10437);
nand NAND2 (N10443, N10434, N9426);
xor XOR2 (N10444, N10423, N6017);
xor XOR2 (N10445, N10443, N2790);
buf BUF1 (N10446, N10445);
and AND2 (N10447, N10440, N3683);
buf BUF1 (N10448, N10442);
xor XOR2 (N10449, N10426, N2609);
not NOT1 (N10450, N10435);
and AND4 (N10451, N10449, N9989, N6263, N2083);
or OR2 (N10452, N10444, N696);
nor NOR4 (N10453, N10450, N6626, N9757, N5028);
or OR3 (N10454, N10446, N1744, N5197);
or OR4 (N10455, N10454, N5976, N1204, N671);
nor NOR4 (N10456, N10439, N4060, N2237, N1069);
and AND4 (N10457, N10451, N4313, N4470, N3934);
xor XOR2 (N10458, N10447, N2982);
buf BUF1 (N10459, N10452);
and AND3 (N10460, N10456, N9358, N2315);
buf BUF1 (N10461, N10455);
nor NOR3 (N10462, N10448, N2621, N683);
buf BUF1 (N10463, N10462);
not NOT1 (N10464, N10432);
nand NAND4 (N10465, N10461, N3006, N7354, N3384);
buf BUF1 (N10466, N10459);
nand NAND4 (N10467, N10464, N919, N5872, N2035);
and AND3 (N10468, N10457, N8568, N5445);
buf BUF1 (N10469, N10460);
nor NOR4 (N10470, N10453, N5301, N8773, N4086);
not NOT1 (N10471, N10458);
buf BUF1 (N10472, N10418);
nand NAND3 (N10473, N10463, N10468, N7224);
and AND4 (N10474, N9588, N7266, N8895, N10024);
nor NOR4 (N10475, N10472, N9060, N2686, N10252);
nand NAND2 (N10476, N10465, N4215);
xor XOR2 (N10477, N10470, N9542);
buf BUF1 (N10478, N10476);
buf BUF1 (N10479, N10469);
and AND3 (N10480, N10478, N3054, N4066);
and AND2 (N10481, N10479, N6673);
nor NOR3 (N10482, N10466, N5243, N7513);
and AND2 (N10483, N10441, N2069);
nand NAND4 (N10484, N10483, N4121, N6401, N3781);
buf BUF1 (N10485, N10467);
nor NOR4 (N10486, N10485, N5016, N3694, N5560);
not NOT1 (N10487, N10486);
nor NOR2 (N10488, N10482, N7352);
or OR3 (N10489, N10480, N1685, N2269);
and AND2 (N10490, N10487, N9587);
xor XOR2 (N10491, N10488, N499);
xor XOR2 (N10492, N10481, N10140);
xor XOR2 (N10493, N10489, N8336);
or OR2 (N10494, N10492, N977);
nand NAND3 (N10495, N10474, N10249, N6800);
xor XOR2 (N10496, N10484, N6504);
nor NOR3 (N10497, N10490, N9034, N3029);
buf BUF1 (N10498, N10491);
xor XOR2 (N10499, N10493, N17);
and AND4 (N10500, N10471, N7229, N2116, N4820);
or OR4 (N10501, N10496, N1201, N10199, N6557);
nor NOR2 (N10502, N10497, N5405);
xor XOR2 (N10503, N10500, N8356);
or OR2 (N10504, N10499, N3952);
xor XOR2 (N10505, N10477, N3715);
not NOT1 (N10506, N10494);
xor XOR2 (N10507, N10506, N6981);
nor NOR4 (N10508, N10501, N10159, N2510, N3956);
nand NAND4 (N10509, N10504, N620, N7285, N1510);
nand NAND3 (N10510, N10473, N2289, N8264);
xor XOR2 (N10511, N10475, N343);
and AND4 (N10512, N10498, N3542, N8228, N59);
nand NAND4 (N10513, N10510, N9887, N5490, N8817);
nand NAND2 (N10514, N10507, N1588);
and AND4 (N10515, N10511, N6075, N6761, N3060);
and AND2 (N10516, N10509, N6376);
or OR4 (N10517, N10502, N4757, N822, N3862);
nor NOR4 (N10518, N10495, N8075, N8461, N5359);
xor XOR2 (N10519, N10505, N3856);
or OR4 (N10520, N10514, N3601, N803, N6361);
buf BUF1 (N10521, N10515);
and AND2 (N10522, N10517, N8607);
buf BUF1 (N10523, N10520);
and AND3 (N10524, N10503, N10246, N2916);
buf BUF1 (N10525, N10512);
or OR2 (N10526, N10525, N9277);
nor NOR2 (N10527, N10521, N4789);
nand NAND4 (N10528, N10518, N2838, N2114, N4512);
nor NOR4 (N10529, N10522, N1555, N7068, N4254);
and AND4 (N10530, N10513, N6324, N9056, N4202);
or OR4 (N10531, N10527, N7694, N5553, N44);
not NOT1 (N10532, N10528);
not NOT1 (N10533, N10532);
buf BUF1 (N10534, N10508);
or OR4 (N10535, N10529, N3219, N4892, N8194);
or OR2 (N10536, N10531, N968);
nand NAND2 (N10537, N10524, N2114);
xor XOR2 (N10538, N10519, N6525);
buf BUF1 (N10539, N10535);
nand NAND3 (N10540, N10526, N1540, N8218);
nor NOR4 (N10541, N10530, N4969, N1219, N560);
nand NAND3 (N10542, N10538, N4383, N2466);
buf BUF1 (N10543, N10537);
nor NOR3 (N10544, N10543, N9611, N7746);
and AND4 (N10545, N10523, N4395, N10146, N539);
xor XOR2 (N10546, N10540, N8873);
nor NOR4 (N10547, N10534, N6394, N6222, N7769);
and AND2 (N10548, N10546, N1658);
nor NOR2 (N10549, N10536, N2754);
and AND3 (N10550, N10548, N8470, N10433);
and AND3 (N10551, N10533, N9748, N5017);
nor NOR4 (N10552, N10551, N4746, N3796, N3277);
or OR3 (N10553, N10545, N10023, N1064);
and AND2 (N10554, N10544, N5534);
not NOT1 (N10555, N10516);
nor NOR4 (N10556, N10542, N4872, N3971, N4141);
or OR2 (N10557, N10554, N4433);
nand NAND3 (N10558, N10552, N7, N2454);
or OR4 (N10559, N10549, N8387, N8996, N4369);
not NOT1 (N10560, N10553);
xor XOR2 (N10561, N10541, N2792);
not NOT1 (N10562, N10555);
and AND2 (N10563, N10558, N7052);
nand NAND2 (N10564, N10562, N4916);
xor XOR2 (N10565, N10557, N2281);
and AND3 (N10566, N10564, N1147, N724);
not NOT1 (N10567, N10539);
buf BUF1 (N10568, N10563);
not NOT1 (N10569, N10547);
xor XOR2 (N10570, N10560, N9996);
nor NOR4 (N10571, N10566, N10556, N2214, N8134);
nand NAND3 (N10572, N1238, N6898, N5132);
and AND4 (N10573, N10561, N9854, N9019, N7728);
nand NAND4 (N10574, N10569, N9572, N5785, N4864);
xor XOR2 (N10575, N10572, N8059);
not NOT1 (N10576, N10575);
buf BUF1 (N10577, N10573);
or OR2 (N10578, N10571, N6574);
nand NAND2 (N10579, N10578, N8188);
not NOT1 (N10580, N10567);
nand NAND3 (N10581, N10579, N3802, N1470);
nor NOR3 (N10582, N10581, N10383, N7422);
nor NOR3 (N10583, N10568, N10259, N4058);
nor NOR2 (N10584, N10576, N1468);
nor NOR2 (N10585, N10584, N1607);
nor NOR3 (N10586, N10550, N1008, N6393);
nand NAND2 (N10587, N10570, N3091);
buf BUF1 (N10588, N10582);
or OR4 (N10589, N10559, N3866, N554, N8812);
and AND3 (N10590, N10565, N10367, N339);
buf BUF1 (N10591, N10585);
and AND3 (N10592, N10577, N8932, N2549);
or OR3 (N10593, N10587, N9787, N9519);
or OR4 (N10594, N10593, N223, N6363, N5531);
not NOT1 (N10595, N10589);
not NOT1 (N10596, N10583);
nand NAND2 (N10597, N10590, N10043);
xor XOR2 (N10598, N10586, N1081);
nor NOR2 (N10599, N10598, N6335);
and AND4 (N10600, N10595, N2160, N3303, N7907);
xor XOR2 (N10601, N10588, N7776);
buf BUF1 (N10602, N10600);
not NOT1 (N10603, N10599);
or OR3 (N10604, N10591, N9087, N8911);
xor XOR2 (N10605, N10604, N9125);
buf BUF1 (N10606, N10592);
and AND3 (N10607, N10596, N9582, N2673);
nand NAND4 (N10608, N10597, N9062, N10143, N2455);
and AND3 (N10609, N10603, N9791, N10115);
or OR3 (N10610, N10574, N1752, N1127);
not NOT1 (N10611, N10580);
or OR3 (N10612, N10602, N4461, N4249);
xor XOR2 (N10613, N10606, N676);
nand NAND3 (N10614, N10610, N8036, N415);
not NOT1 (N10615, N10611);
nor NOR3 (N10616, N10605, N5914, N1733);
not NOT1 (N10617, N10615);
buf BUF1 (N10618, N10601);
not NOT1 (N10619, N10608);
nor NOR4 (N10620, N10607, N9857, N1336, N6306);
or OR3 (N10621, N10594, N1413, N9627);
buf BUF1 (N10622, N10614);
or OR4 (N10623, N10622, N8394, N2668, N6173);
xor XOR2 (N10624, N10616, N2785);
nand NAND4 (N10625, N10613, N6063, N5471, N2798);
nor NOR3 (N10626, N10620, N7492, N10049);
buf BUF1 (N10627, N10621);
buf BUF1 (N10628, N10624);
and AND4 (N10629, N10609, N3502, N1265, N5533);
nor NOR4 (N10630, N10627, N8899, N2601, N8983);
buf BUF1 (N10631, N10628);
buf BUF1 (N10632, N10612);
not NOT1 (N10633, N10619);
nor NOR4 (N10634, N10632, N8679, N1239, N4431);
xor XOR2 (N10635, N10630, N9617);
or OR3 (N10636, N10617, N7678, N2675);
and AND2 (N10637, N10629, N4398);
nor NOR4 (N10638, N10626, N7473, N2193, N1545);
not NOT1 (N10639, N10637);
and AND3 (N10640, N10638, N9431, N128);
xor XOR2 (N10641, N10639, N6675);
and AND4 (N10642, N10633, N8062, N7555, N8817);
or OR3 (N10643, N10641, N9145, N3392);
nand NAND4 (N10644, N10636, N7249, N80, N9050);
xor XOR2 (N10645, N10634, N4550);
or OR3 (N10646, N10642, N6958, N5168);
nand NAND3 (N10647, N10645, N5231, N9742);
or OR4 (N10648, N10623, N7981, N497, N9801);
not NOT1 (N10649, N10646);
and AND2 (N10650, N10648, N4208);
not NOT1 (N10651, N10650);
buf BUF1 (N10652, N10631);
nor NOR3 (N10653, N10625, N5068, N8489);
nor NOR2 (N10654, N10647, N8666);
buf BUF1 (N10655, N10649);
and AND3 (N10656, N10654, N9756, N521);
not NOT1 (N10657, N10643);
nor NOR3 (N10658, N10644, N8938, N745);
not NOT1 (N10659, N10618);
or OR4 (N10660, N10656, N2394, N5908, N1156);
xor XOR2 (N10661, N10651, N6745);
buf BUF1 (N10662, N10660);
nor NOR2 (N10663, N10661, N6052);
nand NAND4 (N10664, N10662, N4064, N8451, N6184);
nand NAND2 (N10665, N10657, N3368);
not NOT1 (N10666, N10665);
not NOT1 (N10667, N10653);
not NOT1 (N10668, N10664);
buf BUF1 (N10669, N10652);
and AND3 (N10670, N10667, N504, N3850);
nand NAND2 (N10671, N10640, N3792);
xor XOR2 (N10672, N10666, N4843);
and AND4 (N10673, N10671, N7330, N10414, N3379);
and AND4 (N10674, N10672, N5048, N1801, N5986);
or OR2 (N10675, N10663, N1137);
nand NAND4 (N10676, N10669, N3249, N7812, N5042);
nand NAND4 (N10677, N10674, N4336, N314, N2284);
nor NOR2 (N10678, N10675, N8874);
nand NAND2 (N10679, N10655, N9581);
or OR2 (N10680, N10678, N1261);
buf BUF1 (N10681, N10680);
not NOT1 (N10682, N10670);
buf BUF1 (N10683, N10677);
or OR2 (N10684, N10679, N10430);
buf BUF1 (N10685, N10659);
not NOT1 (N10686, N10685);
xor XOR2 (N10687, N10673, N197);
xor XOR2 (N10688, N10681, N4089);
buf BUF1 (N10689, N10676);
or OR4 (N10690, N10688, N3681, N10038, N3043);
xor XOR2 (N10691, N10635, N3651);
xor XOR2 (N10692, N10690, N3356);
xor XOR2 (N10693, N10692, N2382);
nand NAND3 (N10694, N10658, N10091, N8519);
or OR4 (N10695, N10684, N3725, N4919, N7271);
buf BUF1 (N10696, N10682);
and AND4 (N10697, N10689, N10291, N4912, N1081);
xor XOR2 (N10698, N10691, N658);
nor NOR4 (N10699, N10698, N5549, N10308, N9513);
buf BUF1 (N10700, N10697);
not NOT1 (N10701, N10693);
nand NAND3 (N10702, N10699, N3809, N2661);
not NOT1 (N10703, N10695);
nor NOR3 (N10704, N10696, N2602, N3128);
buf BUF1 (N10705, N10702);
and AND2 (N10706, N10694, N7372);
not NOT1 (N10707, N10668);
not NOT1 (N10708, N10705);
nor NOR2 (N10709, N10708, N10437);
nor NOR4 (N10710, N10707, N3957, N5823, N10189);
buf BUF1 (N10711, N10704);
nand NAND2 (N10712, N10710, N3625);
buf BUF1 (N10713, N10700);
or OR3 (N10714, N10706, N9301, N192);
nand NAND4 (N10715, N10711, N1316, N126, N9588);
nand NAND2 (N10716, N10714, N6840);
nor NOR3 (N10717, N10703, N8125, N1751);
buf BUF1 (N10718, N10709);
not NOT1 (N10719, N10701);
or OR4 (N10720, N10719, N814, N9591, N5241);
nor NOR2 (N10721, N10715, N10122);
nor NOR2 (N10722, N10683, N4959);
nor NOR2 (N10723, N10721, N10060);
or OR2 (N10724, N10720, N1369);
nor NOR2 (N10725, N10686, N8777);
and AND4 (N10726, N10712, N747, N2268, N8178);
and AND2 (N10727, N10726, N6610);
nand NAND2 (N10728, N10727, N2174);
nand NAND3 (N10729, N10718, N5854, N8097);
buf BUF1 (N10730, N10728);
or OR2 (N10731, N10716, N1931);
buf BUF1 (N10732, N10713);
nor NOR3 (N10733, N10717, N2909, N2741);
nand NAND2 (N10734, N10731, N5852);
buf BUF1 (N10735, N10723);
and AND3 (N10736, N10735, N5175, N4190);
buf BUF1 (N10737, N10732);
or OR4 (N10738, N10736, N1090, N3738, N5318);
buf BUF1 (N10739, N10722);
and AND3 (N10740, N10730, N796, N8380);
xor XOR2 (N10741, N10738, N2241);
or OR3 (N10742, N10725, N1159, N3140);
not NOT1 (N10743, N10739);
nor NOR3 (N10744, N10742, N1490, N169);
xor XOR2 (N10745, N10743, N5106);
buf BUF1 (N10746, N10724);
nand NAND2 (N10747, N10733, N8831);
xor XOR2 (N10748, N10740, N10159);
and AND2 (N10749, N10746, N8877);
not NOT1 (N10750, N10729);
not NOT1 (N10751, N10745);
not NOT1 (N10752, N10737);
nand NAND2 (N10753, N10687, N1371);
nor NOR2 (N10754, N10749, N2007);
or OR2 (N10755, N10748, N10139);
nor NOR4 (N10756, N10744, N9805, N4263, N217);
and AND2 (N10757, N10755, N2732);
nor NOR2 (N10758, N10741, N9756);
and AND2 (N10759, N10753, N10461);
nand NAND4 (N10760, N10759, N7338, N7488, N10);
nor NOR3 (N10761, N10747, N4998, N8809);
or OR2 (N10762, N10752, N7219);
buf BUF1 (N10763, N10757);
xor XOR2 (N10764, N10763, N3676);
or OR4 (N10765, N10754, N9519, N8095, N10591);
nand NAND2 (N10766, N10734, N10415);
nand NAND4 (N10767, N10758, N4202, N5307, N83);
buf BUF1 (N10768, N10762);
buf BUF1 (N10769, N10765);
nand NAND2 (N10770, N10750, N10750);
and AND3 (N10771, N10769, N332, N5547);
not NOT1 (N10772, N10761);
buf BUF1 (N10773, N10772);
or OR2 (N10774, N10771, N1676);
nor NOR4 (N10775, N10760, N1473, N523, N6090);
xor XOR2 (N10776, N10775, N6133);
and AND2 (N10777, N10770, N5761);
buf BUF1 (N10778, N10764);
not NOT1 (N10779, N10777);
not NOT1 (N10780, N10773);
nand NAND4 (N10781, N10774, N26, N8129, N3766);
xor XOR2 (N10782, N10780, N2017);
not NOT1 (N10783, N10756);
xor XOR2 (N10784, N10767, N8202);
or OR2 (N10785, N10783, N709);
buf BUF1 (N10786, N10766);
or OR2 (N10787, N10768, N4671);
not NOT1 (N10788, N10776);
not NOT1 (N10789, N10751);
nor NOR4 (N10790, N10788, N5567, N5948, N187);
or OR2 (N10791, N10784, N7106);
buf BUF1 (N10792, N10789);
xor XOR2 (N10793, N10785, N9246);
nand NAND2 (N10794, N10791, N4084);
nor NOR4 (N10795, N10787, N5206, N9323, N2231);
and AND4 (N10796, N10779, N10448, N9935, N7259);
xor XOR2 (N10797, N10794, N8284);
and AND4 (N10798, N10786, N4581, N5657, N155);
and AND3 (N10799, N10782, N1839, N5178);
nand NAND2 (N10800, N10781, N8674);
xor XOR2 (N10801, N10799, N3742);
not NOT1 (N10802, N10778);
xor XOR2 (N10803, N10793, N1519);
nand NAND4 (N10804, N10803, N10401, N4383, N3546);
buf BUF1 (N10805, N10796);
or OR3 (N10806, N10800, N496, N10321);
buf BUF1 (N10807, N10804);
or OR4 (N10808, N10806, N5544, N6389, N9931);
xor XOR2 (N10809, N10792, N9626);
buf BUF1 (N10810, N10797);
xor XOR2 (N10811, N10809, N9335);
nor NOR3 (N10812, N10805, N6943, N4401);
xor XOR2 (N10813, N10801, N8291);
nand NAND2 (N10814, N10807, N8112);
or OR3 (N10815, N10814, N6099, N8041);
not NOT1 (N10816, N10795);
and AND2 (N10817, N10802, N9906);
nor NOR4 (N10818, N10810, N8266, N1123, N6686);
xor XOR2 (N10819, N10790, N2422);
xor XOR2 (N10820, N10816, N1057);
buf BUF1 (N10821, N10815);
not NOT1 (N10822, N10808);
not NOT1 (N10823, N10811);
xor XOR2 (N10824, N10820, N3997);
and AND2 (N10825, N10823, N1724);
buf BUF1 (N10826, N10822);
and AND3 (N10827, N10812, N3175, N8326);
nor NOR3 (N10828, N10817, N5124, N6353);
or OR2 (N10829, N10819, N1187);
not NOT1 (N10830, N10798);
or OR4 (N10831, N10826, N4167, N5465, N9956);
xor XOR2 (N10832, N10831, N391);
buf BUF1 (N10833, N10830);
and AND4 (N10834, N10828, N6684, N4845, N8394);
nand NAND2 (N10835, N10834, N2353);
or OR4 (N10836, N10813, N7915, N71, N3681);
not NOT1 (N10837, N10827);
not NOT1 (N10838, N10837);
xor XOR2 (N10839, N10833, N6462);
nor NOR4 (N10840, N10838, N1576, N8907, N3636);
nor NOR4 (N10841, N10821, N8635, N4782, N3535);
nor NOR2 (N10842, N10839, N2889);
and AND2 (N10843, N10825, N913);
not NOT1 (N10844, N10836);
nand NAND4 (N10845, N10841, N4163, N3400, N2511);
nand NAND2 (N10846, N10840, N2250);
not NOT1 (N10847, N10832);
and AND3 (N10848, N10845, N5908, N10643);
buf BUF1 (N10849, N10843);
and AND3 (N10850, N10844, N1170, N3840);
or OR4 (N10851, N10829, N1083, N3540, N10812);
buf BUF1 (N10852, N10846);
nand NAND2 (N10853, N10818, N904);
buf BUF1 (N10854, N10852);
xor XOR2 (N10855, N10854, N6972);
not NOT1 (N10856, N10842);
and AND2 (N10857, N10848, N2474);
and AND3 (N10858, N10855, N10740, N3827);
nor NOR3 (N10859, N10858, N9148, N9791);
not NOT1 (N10860, N10851);
not NOT1 (N10861, N10857);
nor NOR4 (N10862, N10860, N458, N1453, N3389);
or OR2 (N10863, N10850, N6870);
and AND2 (N10864, N10847, N2446);
xor XOR2 (N10865, N10856, N8226);
buf BUF1 (N10866, N10863);
buf BUF1 (N10867, N10862);
nand NAND4 (N10868, N10865, N3154, N7720, N4688);
not NOT1 (N10869, N10861);
buf BUF1 (N10870, N10867);
nand NAND3 (N10871, N10859, N6628, N53);
not NOT1 (N10872, N10824);
xor XOR2 (N10873, N10835, N10796);
buf BUF1 (N10874, N10866);
not NOT1 (N10875, N10870);
nor NOR4 (N10876, N10874, N76, N6561, N5588);
not NOT1 (N10877, N10875);
buf BUF1 (N10878, N10871);
xor XOR2 (N10879, N10868, N3796);
and AND3 (N10880, N10872, N5039, N9553);
nand NAND2 (N10881, N10876, N3762);
or OR4 (N10882, N10869, N3180, N9101, N7207);
nand NAND3 (N10883, N10853, N7389, N9648);
xor XOR2 (N10884, N10873, N7076);
not NOT1 (N10885, N10881);
or OR2 (N10886, N10879, N8099);
xor XOR2 (N10887, N10884, N265);
buf BUF1 (N10888, N10849);
nand NAND2 (N10889, N10864, N5735);
xor XOR2 (N10890, N10885, N3536);
buf BUF1 (N10891, N10888);
and AND2 (N10892, N10889, N550);
xor XOR2 (N10893, N10891, N6724);
nand NAND2 (N10894, N10893, N6498);
and AND2 (N10895, N10878, N10763);
buf BUF1 (N10896, N10886);
not NOT1 (N10897, N10880);
nand NAND2 (N10898, N10897, N8494);
buf BUF1 (N10899, N10890);
buf BUF1 (N10900, N10892);
nor NOR3 (N10901, N10895, N4366, N8547);
nand NAND3 (N10902, N10898, N7178, N2941);
and AND2 (N10903, N10882, N9448);
and AND4 (N10904, N10901, N1452, N632, N158);
and AND3 (N10905, N10900, N2555, N10256);
xor XOR2 (N10906, N10896, N9130);
buf BUF1 (N10907, N10904);
buf BUF1 (N10908, N10907);
and AND3 (N10909, N10908, N1010, N10068);
nor NOR4 (N10910, N10909, N3115, N8509, N8265);
nand NAND3 (N10911, N10910, N2690, N10806);
xor XOR2 (N10912, N10877, N10573);
buf BUF1 (N10913, N10903);
nand NAND2 (N10914, N10906, N1028);
or OR3 (N10915, N10883, N3898, N8818);
not NOT1 (N10916, N10913);
not NOT1 (N10917, N10902);
and AND4 (N10918, N10899, N3956, N1272, N4712);
buf BUF1 (N10919, N10905);
buf BUF1 (N10920, N10915);
or OR4 (N10921, N10916, N7145, N8457, N7923);
nor NOR3 (N10922, N10917, N10209, N3548);
and AND3 (N10923, N10887, N9740, N8288);
buf BUF1 (N10924, N10920);
xor XOR2 (N10925, N10912, N602);
not NOT1 (N10926, N10911);
or OR2 (N10927, N10921, N5148);
xor XOR2 (N10928, N10924, N9172);
xor XOR2 (N10929, N10918, N10801);
xor XOR2 (N10930, N10926, N6740);
buf BUF1 (N10931, N10925);
or OR3 (N10932, N10931, N2320, N7999);
nand NAND4 (N10933, N10919, N325, N6949, N41);
not NOT1 (N10934, N10928);
not NOT1 (N10935, N10927);
buf BUF1 (N10936, N10933);
buf BUF1 (N10937, N10932);
buf BUF1 (N10938, N10936);
and AND2 (N10939, N10922, N3915);
and AND3 (N10940, N10937, N3222, N6958);
nor NOR4 (N10941, N10914, N1215, N8585, N9602);
and AND4 (N10942, N10894, N9916, N7750, N8293);
xor XOR2 (N10943, N10939, N8115);
buf BUF1 (N10944, N10943);
xor XOR2 (N10945, N10935, N3633);
and AND3 (N10946, N10938, N9931, N9244);
xor XOR2 (N10947, N10942, N1843);
and AND3 (N10948, N10940, N10291, N2164);
xor XOR2 (N10949, N10947, N132);
buf BUF1 (N10950, N10946);
or OR2 (N10951, N10941, N6379);
nand NAND2 (N10952, N10929, N1912);
or OR4 (N10953, N10950, N5943, N6282, N1161);
xor XOR2 (N10954, N10952, N2406);
not NOT1 (N10955, N10923);
and AND4 (N10956, N10954, N8225, N4739, N3195);
not NOT1 (N10957, N10930);
and AND2 (N10958, N10944, N9569);
nor NOR4 (N10959, N10951, N1851, N4373, N1359);
buf BUF1 (N10960, N10957);
or OR2 (N10961, N10955, N2621);
nand NAND2 (N10962, N10960, N460);
not NOT1 (N10963, N10958);
or OR4 (N10964, N10956, N2794, N1854, N9023);
not NOT1 (N10965, N10934);
xor XOR2 (N10966, N10962, N4821);
not NOT1 (N10967, N10948);
buf BUF1 (N10968, N10959);
and AND4 (N10969, N10945, N517, N7858, N3172);
or OR4 (N10970, N10967, N10742, N9517, N6660);
nand NAND4 (N10971, N10963, N7823, N2498, N1823);
xor XOR2 (N10972, N10971, N4068);
or OR4 (N10973, N10968, N9872, N5486, N2642);
nor NOR3 (N10974, N10949, N5638, N5067);
buf BUF1 (N10975, N10965);
nor NOR4 (N10976, N10964, N7331, N9781, N9043);
nor NOR2 (N10977, N10969, N2256);
buf BUF1 (N10978, N10977);
or OR4 (N10979, N10972, N309, N10944, N3855);
xor XOR2 (N10980, N10975, N1132);
or OR4 (N10981, N10974, N7656, N3051, N7789);
or OR4 (N10982, N10953, N8118, N3834, N944);
and AND3 (N10983, N10966, N403, N4973);
not NOT1 (N10984, N10973);
not NOT1 (N10985, N10983);
xor XOR2 (N10986, N10961, N3288);
buf BUF1 (N10987, N10982);
nor NOR2 (N10988, N10979, N10764);
and AND4 (N10989, N10978, N6379, N5292, N4509);
not NOT1 (N10990, N10976);
or OR4 (N10991, N10981, N7172, N618, N3777);
and AND2 (N10992, N10980, N1793);
nor NOR3 (N10993, N10970, N1802, N3186);
nand NAND4 (N10994, N10992, N370, N1696, N2976);
nor NOR4 (N10995, N10990, N2823, N8229, N2051);
xor XOR2 (N10996, N10988, N7736);
and AND4 (N10997, N10993, N10575, N9337, N828);
nor NOR2 (N10998, N10994, N3122);
and AND2 (N10999, N10985, N3420);
nor NOR2 (N11000, N10984, N460);
or OR3 (N11001, N10997, N1597, N5288);
or OR2 (N11002, N10998, N5718);
and AND4 (N11003, N10986, N2740, N10769, N10717);
xor XOR2 (N11004, N10991, N10522);
and AND3 (N11005, N10999, N10083, N4422);
nand NAND3 (N11006, N11004, N2320, N4081);
and AND4 (N11007, N11006, N7434, N7756, N8162);
not NOT1 (N11008, N11005);
buf BUF1 (N11009, N11003);
and AND4 (N11010, N10995, N1340, N8728, N1493);
or OR4 (N11011, N11010, N4185, N10057, N234);
nand NAND2 (N11012, N11001, N274);
nor NOR3 (N11013, N11002, N10493, N3818);
buf BUF1 (N11014, N11000);
xor XOR2 (N11015, N11008, N4779);
or OR4 (N11016, N11011, N2232, N9585, N7130);
nor NOR2 (N11017, N10996, N5855);
nand NAND2 (N11018, N11017, N9695);
and AND2 (N11019, N11016, N7461);
xor XOR2 (N11020, N11009, N7124);
not NOT1 (N11021, N11020);
nand NAND2 (N11022, N10989, N8864);
and AND3 (N11023, N11022, N2416, N1690);
or OR4 (N11024, N11007, N2035, N8589, N6652);
or OR4 (N11025, N11018, N3443, N566, N10807);
and AND2 (N11026, N11019, N10659);
xor XOR2 (N11027, N11023, N6786);
xor XOR2 (N11028, N11026, N696);
or OR4 (N11029, N11025, N7541, N9343, N6528);
nand NAND4 (N11030, N11015, N487, N9438, N5224);
nor NOR2 (N11031, N10987, N7283);
and AND4 (N11032, N11027, N5850, N7450, N10761);
buf BUF1 (N11033, N11012);
or OR3 (N11034, N11030, N5868, N7099);
nor NOR2 (N11035, N11013, N3472);
buf BUF1 (N11036, N11028);
or OR4 (N11037, N11014, N8128, N8173, N5338);
not NOT1 (N11038, N11021);
nand NAND3 (N11039, N11033, N7147, N5469);
nor NOR3 (N11040, N11031, N8471, N6628);
or OR4 (N11041, N11039, N2567, N1887, N7709);
xor XOR2 (N11042, N11032, N10685);
nand NAND3 (N11043, N11040, N8730, N9873);
buf BUF1 (N11044, N11029);
xor XOR2 (N11045, N11035, N1024);
nand NAND3 (N11046, N11045, N4083, N388);
buf BUF1 (N11047, N11037);
and AND2 (N11048, N11036, N10139);
xor XOR2 (N11049, N11044, N3248);
nor NOR3 (N11050, N11041, N498, N9573);
nor NOR4 (N11051, N11047, N10547, N1248, N7328);
nand NAND4 (N11052, N11034, N8105, N10772, N7770);
xor XOR2 (N11053, N11051, N1018);
xor XOR2 (N11054, N11043, N1650);
buf BUF1 (N11055, N11050);
and AND2 (N11056, N11054, N2865);
and AND4 (N11057, N11038, N776, N6879, N3771);
or OR3 (N11058, N11053, N4488, N2852);
xor XOR2 (N11059, N11046, N9265);
nand NAND4 (N11060, N11049, N9411, N1182, N2451);
nor NOR2 (N11061, N11060, N3093);
not NOT1 (N11062, N11055);
nor NOR2 (N11063, N11052, N200);
not NOT1 (N11064, N11062);
and AND4 (N11065, N11057, N830, N209, N1133);
and AND3 (N11066, N11063, N9677, N7949);
nand NAND4 (N11067, N11048, N4518, N7541, N2019);
nand NAND3 (N11068, N11042, N6465, N7729);
nand NAND3 (N11069, N11067, N9294, N2344);
nor NOR2 (N11070, N11056, N6617);
or OR2 (N11071, N11024, N3444);
buf BUF1 (N11072, N11065);
nand NAND4 (N11073, N11072, N2000, N9791, N385);
xor XOR2 (N11074, N11058, N2719);
nand NAND4 (N11075, N11061, N8909, N6040, N1868);
nor NOR2 (N11076, N11071, N7121);
nand NAND4 (N11077, N11064, N4958, N53, N2073);
and AND2 (N11078, N11066, N5349);
nand NAND2 (N11079, N11077, N1663);
nor NOR2 (N11080, N11074, N9730);
not NOT1 (N11081, N11073);
nor NOR4 (N11082, N11070, N4641, N10635, N5670);
nand NAND4 (N11083, N11078, N4480, N7037, N7578);
or OR4 (N11084, N11068, N3598, N3245, N7470);
not NOT1 (N11085, N11080);
nand NAND2 (N11086, N11083, N11053);
nor NOR2 (N11087, N11076, N2636);
and AND4 (N11088, N11087, N3572, N4654, N2340);
buf BUF1 (N11089, N11069);
nor NOR3 (N11090, N11059, N9649, N6474);
xor XOR2 (N11091, N11085, N6431);
and AND2 (N11092, N11088, N8244);
not NOT1 (N11093, N11086);
nand NAND2 (N11094, N11090, N4039);
not NOT1 (N11095, N11082);
and AND2 (N11096, N11092, N6078);
buf BUF1 (N11097, N11091);
or OR4 (N11098, N11075, N8982, N2227, N9364);
xor XOR2 (N11099, N11098, N11074);
buf BUF1 (N11100, N11097);
and AND2 (N11101, N11081, N7987);
and AND3 (N11102, N11084, N8608, N6176);
nand NAND3 (N11103, N11101, N2718, N9216);
nand NAND2 (N11104, N11096, N3645);
xor XOR2 (N11105, N11089, N7972);
buf BUF1 (N11106, N11104);
nor NOR2 (N11107, N11093, N4231);
or OR2 (N11108, N11095, N8765);
or OR4 (N11109, N11103, N969, N5550, N281);
xor XOR2 (N11110, N11102, N8260);
buf BUF1 (N11111, N11106);
or OR4 (N11112, N11094, N8612, N8744, N21);
nand NAND2 (N11113, N11079, N4282);
or OR4 (N11114, N11099, N8444, N10871, N3323);
xor XOR2 (N11115, N11100, N10202);
and AND4 (N11116, N11109, N3017, N6038, N7087);
not NOT1 (N11117, N11107);
nand NAND2 (N11118, N11110, N9987);
nor NOR3 (N11119, N11112, N7218, N2907);
xor XOR2 (N11120, N11111, N9183);
and AND2 (N11121, N11115, N5708);
xor XOR2 (N11122, N11120, N3960);
not NOT1 (N11123, N11119);
nor NOR2 (N11124, N11118, N6183);
nand NAND2 (N11125, N11123, N4306);
and AND4 (N11126, N11114, N8636, N511, N9955);
nor NOR3 (N11127, N11124, N2862, N3071);
buf BUF1 (N11128, N11127);
nand NAND4 (N11129, N11126, N6840, N7775, N6672);
nand NAND3 (N11130, N11129, N6826, N7778);
nand NAND2 (N11131, N11125, N3506);
and AND4 (N11132, N11130, N1483, N1714, N2507);
xor XOR2 (N11133, N11131, N5181);
and AND4 (N11134, N11132, N10065, N2463, N8208);
nand NAND2 (N11135, N11122, N1782);
nand NAND4 (N11136, N11135, N9133, N3633, N5788);
or OR4 (N11137, N11113, N7054, N286, N3546);
nand NAND3 (N11138, N11128, N8370, N9732);
xor XOR2 (N11139, N11108, N5403);
buf BUF1 (N11140, N11133);
nand NAND3 (N11141, N11116, N1538, N5425);
nand NAND2 (N11142, N11137, N4706);
and AND2 (N11143, N11142, N9033);
or OR3 (N11144, N11143, N6104, N8714);
buf BUF1 (N11145, N11117);
or OR4 (N11146, N11136, N4063, N10377, N10667);
or OR4 (N11147, N11144, N3820, N3587, N4860);
nor NOR4 (N11148, N11141, N1549, N1333, N4020);
and AND2 (N11149, N11140, N5135);
xor XOR2 (N11150, N11146, N5009);
not NOT1 (N11151, N11134);
buf BUF1 (N11152, N11147);
buf BUF1 (N11153, N11139);
not NOT1 (N11154, N11148);
buf BUF1 (N11155, N11145);
buf BUF1 (N11156, N11138);
xor XOR2 (N11157, N11105, N577);
or OR4 (N11158, N11157, N7136, N4693, N3026);
xor XOR2 (N11159, N11151, N9475);
and AND4 (N11160, N11152, N9735, N10877, N9809);
nand NAND3 (N11161, N11155, N244, N2551);
or OR2 (N11162, N11158, N9069);
and AND3 (N11163, N11159, N5088, N2703);
nor NOR3 (N11164, N11162, N779, N6674);
buf BUF1 (N11165, N11154);
buf BUF1 (N11166, N11153);
nand NAND4 (N11167, N11121, N4606, N9655, N7654);
and AND4 (N11168, N11165, N1721, N3857, N1515);
not NOT1 (N11169, N11160);
not NOT1 (N11170, N11149);
or OR3 (N11171, N11169, N9730, N10747);
not NOT1 (N11172, N11171);
buf BUF1 (N11173, N11161);
nor NOR3 (N11174, N11156, N5853, N10272);
not NOT1 (N11175, N11170);
or OR4 (N11176, N11164, N9701, N4639, N151);
nand NAND3 (N11177, N11176, N9481, N2164);
xor XOR2 (N11178, N11150, N8022);
and AND4 (N11179, N11178, N3849, N4057, N10157);
nor NOR3 (N11180, N11175, N2136, N1376);
and AND4 (N11181, N11172, N3574, N1656, N9823);
not NOT1 (N11182, N11168);
and AND2 (N11183, N11163, N10590);
nand NAND2 (N11184, N11183, N4525);
not NOT1 (N11185, N11182);
buf BUF1 (N11186, N11167);
and AND3 (N11187, N11181, N5468, N2713);
or OR2 (N11188, N11185, N7973);
xor XOR2 (N11189, N11184, N6868);
not NOT1 (N11190, N11174);
nor NOR2 (N11191, N11173, N1746);
not NOT1 (N11192, N11187);
or OR3 (N11193, N11180, N2851, N3475);
and AND4 (N11194, N11179, N3629, N8401, N8159);
and AND3 (N11195, N11188, N2558, N781);
nand NAND4 (N11196, N11194, N10015, N6986, N2556);
not NOT1 (N11197, N11189);
xor XOR2 (N11198, N11195, N5428);
and AND4 (N11199, N11186, N10301, N10728, N4988);
buf BUF1 (N11200, N11198);
xor XOR2 (N11201, N11177, N7579);
xor XOR2 (N11202, N11190, N8629);
nor NOR2 (N11203, N11192, N10961);
nand NAND2 (N11204, N11202, N9675);
nor NOR4 (N11205, N11166, N739, N9610, N2396);
or OR4 (N11206, N11196, N1129, N9422, N580);
buf BUF1 (N11207, N11197);
and AND3 (N11208, N11204, N6972, N1620);
xor XOR2 (N11209, N11203, N2895);
buf BUF1 (N11210, N11208);
not NOT1 (N11211, N11201);
xor XOR2 (N11212, N11211, N10);
nand NAND4 (N11213, N11212, N2636, N9950, N226);
and AND4 (N11214, N11210, N8196, N8272, N11208);
xor XOR2 (N11215, N11214, N8146);
nand NAND4 (N11216, N11193, N4716, N770, N10439);
and AND3 (N11217, N11200, N9807, N6958);
and AND3 (N11218, N11205, N9014, N7688);
nor NOR3 (N11219, N11216, N1327, N10265);
nand NAND3 (N11220, N11219, N2140, N4194);
not NOT1 (N11221, N11217);
nand NAND3 (N11222, N11221, N7154, N579);
buf BUF1 (N11223, N11220);
not NOT1 (N11224, N11206);
buf BUF1 (N11225, N11224);
xor XOR2 (N11226, N11209, N5802);
and AND3 (N11227, N11207, N11156, N8901);
xor XOR2 (N11228, N11227, N4558);
nor NOR3 (N11229, N11213, N7507, N4324);
and AND2 (N11230, N11222, N7973);
buf BUF1 (N11231, N11215);
and AND4 (N11232, N11199, N793, N6856, N3527);
nand NAND2 (N11233, N11225, N2211);
buf BUF1 (N11234, N11226);
not NOT1 (N11235, N11234);
and AND4 (N11236, N11229, N4812, N6231, N1979);
nor NOR3 (N11237, N11230, N2610, N1041);
and AND4 (N11238, N11232, N1939, N3629, N5270);
nor NOR2 (N11239, N11218, N4978);
or OR2 (N11240, N11231, N8318);
not NOT1 (N11241, N11240);
nor NOR2 (N11242, N11239, N5830);
and AND2 (N11243, N11242, N8193);
not NOT1 (N11244, N11241);
nor NOR4 (N11245, N11228, N2636, N7186, N867);
nor NOR4 (N11246, N11191, N9763, N6867, N4058);
nand NAND2 (N11247, N11244, N5969);
not NOT1 (N11248, N11223);
and AND3 (N11249, N11246, N1448, N5821);
and AND3 (N11250, N11245, N11143, N7941);
nor NOR4 (N11251, N11249, N2573, N854, N10593);
or OR3 (N11252, N11247, N8006, N9639);
or OR4 (N11253, N11248, N2971, N10947, N1414);
buf BUF1 (N11254, N11251);
or OR2 (N11255, N11243, N5635);
buf BUF1 (N11256, N11238);
nand NAND3 (N11257, N11237, N2203, N4031);
buf BUF1 (N11258, N11253);
or OR2 (N11259, N11255, N6413);
not NOT1 (N11260, N11233);
nand NAND3 (N11261, N11257, N7101, N9332);
and AND4 (N11262, N11256, N600, N7278, N4792);
not NOT1 (N11263, N11235);
not NOT1 (N11264, N11254);
not NOT1 (N11265, N11252);
buf BUF1 (N11266, N11265);
buf BUF1 (N11267, N11259);
xor XOR2 (N11268, N11258, N6292);
or OR3 (N11269, N11263, N4311, N6801);
or OR4 (N11270, N11266, N11081, N3298, N6639);
nor NOR4 (N11271, N11262, N7153, N3172, N11115);
nor NOR4 (N11272, N11268, N423, N3366, N10876);
buf BUF1 (N11273, N11264);
buf BUF1 (N11274, N11250);
xor XOR2 (N11275, N11274, N4347);
xor XOR2 (N11276, N11272, N10350);
nor NOR4 (N11277, N11276, N6670, N6958, N1316);
buf BUF1 (N11278, N11236);
nor NOR3 (N11279, N11271, N9641, N2930);
buf BUF1 (N11280, N11260);
xor XOR2 (N11281, N11279, N6403);
and AND3 (N11282, N11281, N9569, N9981);
nor NOR2 (N11283, N11280, N9665);
nand NAND4 (N11284, N11270, N10372, N3254, N7087);
and AND3 (N11285, N11278, N3958, N458);
xor XOR2 (N11286, N11282, N19);
nand NAND2 (N11287, N11286, N7368);
nand NAND2 (N11288, N11283, N10976);
xor XOR2 (N11289, N11273, N4021);
xor XOR2 (N11290, N11287, N858);
buf BUF1 (N11291, N11267);
nor NOR2 (N11292, N11275, N11039);
not NOT1 (N11293, N11291);
nand NAND4 (N11294, N11292, N7746, N6837, N5446);
xor XOR2 (N11295, N11294, N79);
nor NOR4 (N11296, N11289, N6348, N7879, N8789);
and AND2 (N11297, N11290, N7811);
xor XOR2 (N11298, N11285, N2639);
or OR2 (N11299, N11284, N6441);
and AND2 (N11300, N11288, N4435);
nand NAND4 (N11301, N11298, N7487, N4042, N6164);
buf BUF1 (N11302, N11295);
or OR3 (N11303, N11293, N8287, N377);
nor NOR3 (N11304, N11300, N10052, N4861);
nor NOR4 (N11305, N11261, N768, N9030, N7501);
and AND3 (N11306, N11302, N6722, N1768);
or OR3 (N11307, N11301, N8085, N1012);
and AND3 (N11308, N11306, N10492, N10339);
xor XOR2 (N11309, N11299, N11293);
buf BUF1 (N11310, N11277);
nand NAND4 (N11311, N11303, N10107, N5451, N2168);
or OR2 (N11312, N11297, N6983);
xor XOR2 (N11313, N11269, N9346);
or OR2 (N11314, N11296, N9284);
xor XOR2 (N11315, N11308, N9393);
xor XOR2 (N11316, N11313, N6532);
nand NAND4 (N11317, N11310, N10289, N1535, N8110);
nor NOR3 (N11318, N11312, N6368, N6900);
buf BUF1 (N11319, N11305);
buf BUF1 (N11320, N11309);
and AND4 (N11321, N11304, N3921, N2345, N10724);
nand NAND4 (N11322, N11307, N4227, N9986, N2218);
buf BUF1 (N11323, N11317);
xor XOR2 (N11324, N11321, N10638);
not NOT1 (N11325, N11324);
nand NAND4 (N11326, N11311, N8155, N10682, N10210);
not NOT1 (N11327, N11325);
and AND3 (N11328, N11316, N5733, N2538);
and AND4 (N11329, N11326, N5198, N270, N8312);
nand NAND4 (N11330, N11320, N3672, N6433, N5253);
or OR4 (N11331, N11323, N8794, N114, N5527);
not NOT1 (N11332, N11319);
or OR3 (N11333, N11330, N3166, N8782);
nand NAND2 (N11334, N11315, N5768);
not NOT1 (N11335, N11329);
xor XOR2 (N11336, N11328, N5431);
buf BUF1 (N11337, N11335);
buf BUF1 (N11338, N11327);
or OR2 (N11339, N11334, N1315);
xor XOR2 (N11340, N11314, N1342);
and AND3 (N11341, N11318, N4393, N1510);
or OR2 (N11342, N11332, N2477);
and AND2 (N11343, N11337, N11314);
not NOT1 (N11344, N11338);
nor NOR2 (N11345, N11342, N9406);
and AND2 (N11346, N11340, N507);
not NOT1 (N11347, N11339);
nand NAND4 (N11348, N11343, N4932, N6385, N180);
and AND3 (N11349, N11331, N4076, N9317);
xor XOR2 (N11350, N11346, N1560);
nor NOR2 (N11351, N11341, N1176);
nand NAND4 (N11352, N11350, N10254, N10880, N2783);
buf BUF1 (N11353, N11345);
or OR2 (N11354, N11322, N1034);
or OR3 (N11355, N11349, N2778, N6182);
nor NOR2 (N11356, N11352, N2728);
nand NAND3 (N11357, N11344, N4202, N2430);
buf BUF1 (N11358, N11351);
not NOT1 (N11359, N11355);
nor NOR2 (N11360, N11359, N918);
nand NAND2 (N11361, N11360, N6598);
xor XOR2 (N11362, N11361, N8291);
buf BUF1 (N11363, N11336);
buf BUF1 (N11364, N11357);
not NOT1 (N11365, N11358);
or OR3 (N11366, N11347, N4268, N9858);
nor NOR3 (N11367, N11348, N4693, N10491);
not NOT1 (N11368, N11366);
buf BUF1 (N11369, N11363);
or OR2 (N11370, N11353, N2029);
or OR4 (N11371, N11333, N7551, N5390, N6371);
nand NAND2 (N11372, N11362, N11254);
xor XOR2 (N11373, N11369, N5137);
and AND2 (N11374, N11364, N10986);
xor XOR2 (N11375, N11370, N6918);
buf BUF1 (N11376, N11374);
not NOT1 (N11377, N11354);
xor XOR2 (N11378, N11373, N8131);
xor XOR2 (N11379, N11375, N1277);
buf BUF1 (N11380, N11376);
buf BUF1 (N11381, N11380);
xor XOR2 (N11382, N11368, N10477);
or OR2 (N11383, N11377, N3557);
xor XOR2 (N11384, N11367, N9985);
xor XOR2 (N11385, N11365, N8020);
buf BUF1 (N11386, N11381);
not NOT1 (N11387, N11379);
or OR2 (N11388, N11372, N11283);
nor NOR4 (N11389, N11383, N10459, N2281, N7183);
and AND3 (N11390, N11388, N834, N5477);
not NOT1 (N11391, N11386);
buf BUF1 (N11392, N11382);
nand NAND3 (N11393, N11390, N10447, N6003);
nand NAND2 (N11394, N11389, N1310);
nor NOR2 (N11395, N11394, N9903);
nand NAND4 (N11396, N11371, N4105, N7954, N2469);
not NOT1 (N11397, N11391);
or OR4 (N11398, N11393, N1118, N7737, N5386);
nor NOR3 (N11399, N11385, N9148, N1126);
xor XOR2 (N11400, N11396, N3283);
buf BUF1 (N11401, N11400);
nor NOR3 (N11402, N11384, N8210, N638);
xor XOR2 (N11403, N11399, N190);
and AND4 (N11404, N11395, N9238, N9926, N8720);
and AND3 (N11405, N11403, N1103, N9830);
buf BUF1 (N11406, N11397);
xor XOR2 (N11407, N11405, N5064);
and AND4 (N11408, N11356, N10087, N9269, N7518);
nand NAND4 (N11409, N11387, N2019, N8999, N6802);
nand NAND3 (N11410, N11398, N8007, N7488);
nor NOR3 (N11411, N11407, N7196, N9810);
or OR3 (N11412, N11406, N130, N6548);
and AND4 (N11413, N11402, N7761, N9758, N7685);
nand NAND3 (N11414, N11401, N5833, N10963);
and AND4 (N11415, N11378, N7031, N5385, N3755);
or OR4 (N11416, N11414, N4187, N1661, N10152);
buf BUF1 (N11417, N11412);
nand NAND4 (N11418, N11413, N2170, N7376, N1286);
and AND2 (N11419, N11417, N2926);
nand NAND4 (N11420, N11411, N5530, N7715, N388);
buf BUF1 (N11421, N11419);
or OR2 (N11422, N11392, N71);
nor NOR2 (N11423, N11421, N7880);
or OR4 (N11424, N11416, N11209, N9042, N254);
or OR4 (N11425, N11418, N8979, N5912, N7560);
and AND2 (N11426, N11409, N4670);
nand NAND4 (N11427, N11422, N9993, N9511, N7834);
xor XOR2 (N11428, N11410, N3392);
nor NOR2 (N11429, N11408, N4310);
not NOT1 (N11430, N11420);
xor XOR2 (N11431, N11425, N533);
buf BUF1 (N11432, N11426);
not NOT1 (N11433, N11424);
nand NAND3 (N11434, N11432, N3773, N2744);
xor XOR2 (N11435, N11431, N472);
nand NAND3 (N11436, N11427, N10183, N6629);
nor NOR3 (N11437, N11423, N11226, N722);
or OR4 (N11438, N11433, N5732, N3997, N4598);
nand NAND2 (N11439, N11438, N934);
nand NAND2 (N11440, N11429, N1799);
or OR4 (N11441, N11430, N9735, N2126, N10376);
nand NAND3 (N11442, N11441, N2163, N740);
not NOT1 (N11443, N11440);
nor NOR2 (N11444, N11436, N7766);
nor NOR3 (N11445, N11434, N1146, N7560);
xor XOR2 (N11446, N11428, N7719);
and AND4 (N11447, N11443, N4898, N2865, N10849);
and AND2 (N11448, N11435, N5032);
not NOT1 (N11449, N11442);
not NOT1 (N11450, N11439);
nand NAND4 (N11451, N11404, N1605, N7149, N3526);
buf BUF1 (N11452, N11437);
nand NAND2 (N11453, N11446, N9642);
buf BUF1 (N11454, N11444);
xor XOR2 (N11455, N11450, N183);
or OR4 (N11456, N11415, N9593, N4379, N6665);
nor NOR2 (N11457, N11451, N5371);
buf BUF1 (N11458, N11455);
or OR3 (N11459, N11456, N8095, N6138);
buf BUF1 (N11460, N11454);
nor NOR2 (N11461, N11447, N6386);
not NOT1 (N11462, N11452);
nor NOR3 (N11463, N11445, N2413, N5780);
nand NAND2 (N11464, N11461, N6319);
and AND3 (N11465, N11464, N5085, N9929);
nand NAND4 (N11466, N11458, N7810, N5717, N4290);
not NOT1 (N11467, N11457);
and AND2 (N11468, N11448, N8534);
nor NOR2 (N11469, N11467, N11139);
or OR4 (N11470, N11453, N925, N1598, N3184);
or OR2 (N11471, N11468, N3992);
nand NAND2 (N11472, N11462, N10464);
or OR3 (N11473, N11463, N6366, N6069);
xor XOR2 (N11474, N11473, N2032);
buf BUF1 (N11475, N11449);
nor NOR2 (N11476, N11474, N11001);
nor NOR3 (N11477, N11470, N3597, N3519);
xor XOR2 (N11478, N11459, N4894);
nor NOR3 (N11479, N11471, N3892, N3239);
nand NAND2 (N11480, N11472, N271);
and AND2 (N11481, N11479, N7440);
or OR4 (N11482, N11460, N6336, N3702, N802);
nand NAND3 (N11483, N11478, N10487, N8761);
or OR4 (N11484, N11482, N5311, N1421, N6555);
buf BUF1 (N11485, N11481);
not NOT1 (N11486, N11483);
or OR4 (N11487, N11486, N1278, N2257, N8503);
nand NAND3 (N11488, N11465, N7261, N1111);
not NOT1 (N11489, N11475);
or OR4 (N11490, N11477, N8397, N7781, N11113);
xor XOR2 (N11491, N11489, N2914);
xor XOR2 (N11492, N11485, N998);
or OR3 (N11493, N11466, N10042, N9158);
xor XOR2 (N11494, N11487, N1051);
not NOT1 (N11495, N11490);
buf BUF1 (N11496, N11495);
xor XOR2 (N11497, N11491, N10217);
xor XOR2 (N11498, N11488, N10539);
or OR4 (N11499, N11496, N1237, N10872, N2132);
xor XOR2 (N11500, N11480, N11244);
and AND4 (N11501, N11500, N3775, N9489, N2283);
nand NAND3 (N11502, N11494, N10565, N5932);
not NOT1 (N11503, N11476);
buf BUF1 (N11504, N11498);
nor NOR3 (N11505, N11499, N8922, N9651);
and AND4 (N11506, N11502, N1722, N11332, N10136);
nor NOR3 (N11507, N11506, N1329, N8876);
xor XOR2 (N11508, N11497, N4184);
buf BUF1 (N11509, N11501);
nand NAND2 (N11510, N11505, N6781);
nand NAND2 (N11511, N11508, N2823);
nand NAND4 (N11512, N11504, N5290, N7777, N9071);
xor XOR2 (N11513, N11507, N1438);
and AND3 (N11514, N11511, N9860, N1120);
not NOT1 (N11515, N11493);
nor NOR3 (N11516, N11513, N3276, N1330);
and AND2 (N11517, N11516, N8865);
not NOT1 (N11518, N11503);
buf BUF1 (N11519, N11517);
and AND4 (N11520, N11518, N2640, N7229, N7545);
xor XOR2 (N11521, N11484, N5608);
nor NOR2 (N11522, N11492, N1719);
nor NOR2 (N11523, N11509, N9166);
or OR3 (N11524, N11522, N8998, N10732);
or OR3 (N11525, N11512, N6588, N605);
buf BUF1 (N11526, N11523);
or OR4 (N11527, N11525, N9474, N1978, N4937);
or OR3 (N11528, N11515, N1918, N5594);
buf BUF1 (N11529, N11469);
nand NAND4 (N11530, N11527, N1704, N6463, N3909);
nand NAND2 (N11531, N11520, N708);
and AND2 (N11532, N11524, N2735);
nor NOR2 (N11533, N11521, N10145);
nand NAND3 (N11534, N11528, N2210, N3705);
not NOT1 (N11535, N11530);
nor NOR3 (N11536, N11534, N4100, N3660);
xor XOR2 (N11537, N11532, N7763);
not NOT1 (N11538, N11535);
nor NOR4 (N11539, N11529, N941, N5211, N5646);
nand NAND3 (N11540, N11537, N6460, N1712);
not NOT1 (N11541, N11540);
xor XOR2 (N11542, N11539, N7964);
nor NOR2 (N11543, N11519, N7079);
xor XOR2 (N11544, N11538, N2749);
xor XOR2 (N11545, N11533, N3323);
nor NOR2 (N11546, N11531, N3060);
nand NAND4 (N11547, N11543, N5096, N7017, N1598);
not NOT1 (N11548, N11545);
and AND4 (N11549, N11536, N4937, N7572, N10287);
buf BUF1 (N11550, N11544);
or OR4 (N11551, N11514, N7327, N443, N1221);
not NOT1 (N11552, N11547);
xor XOR2 (N11553, N11526, N59);
nand NAND4 (N11554, N11552, N5939, N6684, N9776);
or OR3 (N11555, N11553, N8698, N2657);
nor NOR4 (N11556, N11549, N7085, N1423, N8901);
buf BUF1 (N11557, N11555);
and AND3 (N11558, N11542, N3715, N11437);
nand NAND4 (N11559, N11554, N716, N5867, N6702);
nand NAND3 (N11560, N11551, N10007, N7459);
or OR4 (N11561, N11558, N4151, N10283, N9526);
xor XOR2 (N11562, N11541, N10420);
or OR3 (N11563, N11562, N8790, N4060);
or OR3 (N11564, N11510, N7082, N1870);
nand NAND3 (N11565, N11559, N6482, N10354);
xor XOR2 (N11566, N11561, N589);
nand NAND4 (N11567, N11557, N3238, N1230, N91);
not NOT1 (N11568, N11563);
nand NAND4 (N11569, N11568, N4057, N11430, N2842);
nor NOR3 (N11570, N11550, N776, N3400);
and AND4 (N11571, N11565, N1679, N1650, N11114);
nor NOR3 (N11572, N11567, N11082, N7003);
and AND4 (N11573, N11566, N9531, N2318, N9651);
nand NAND3 (N11574, N11570, N3080, N5760);
and AND2 (N11575, N11571, N7283);
and AND3 (N11576, N11564, N1737, N642);
xor XOR2 (N11577, N11560, N4622);
and AND3 (N11578, N11575, N2676, N92);
nor NOR2 (N11579, N11574, N8608);
or OR2 (N11580, N11578, N11010);
xor XOR2 (N11581, N11572, N7646);
or OR2 (N11582, N11569, N1696);
nor NOR3 (N11583, N11579, N11119, N3815);
buf BUF1 (N11584, N11577);
and AND2 (N11585, N11573, N6194);
xor XOR2 (N11586, N11556, N7251);
or OR2 (N11587, N11548, N6417);
xor XOR2 (N11588, N11576, N10843);
nor NOR3 (N11589, N11583, N6332, N3975);
not NOT1 (N11590, N11580);
xor XOR2 (N11591, N11588, N2966);
buf BUF1 (N11592, N11590);
nor NOR3 (N11593, N11591, N8010, N5664);
xor XOR2 (N11594, N11584, N9342);
or OR4 (N11595, N11594, N7413, N9860, N11086);
or OR4 (N11596, N11592, N9403, N6184, N305);
nand NAND4 (N11597, N11585, N11058, N4462, N5308);
buf BUF1 (N11598, N11582);
nand NAND4 (N11599, N11581, N2344, N9105, N2133);
not NOT1 (N11600, N11599);
xor XOR2 (N11601, N11546, N1403);
nor NOR3 (N11602, N11596, N5715, N2945);
buf BUF1 (N11603, N11598);
nand NAND2 (N11604, N11602, N8355);
and AND2 (N11605, N11586, N1093);
nand NAND4 (N11606, N11593, N140, N4628, N7988);
xor XOR2 (N11607, N11603, N9286);
nand NAND2 (N11608, N11597, N8533);
or OR3 (N11609, N11606, N9538, N10871);
or OR4 (N11610, N11609, N1783, N5555, N4248);
and AND2 (N11611, N11600, N11491);
buf BUF1 (N11612, N11607);
and AND4 (N11613, N11611, N4392, N4052, N10705);
nor NOR2 (N11614, N11589, N9094);
nand NAND2 (N11615, N11604, N6039);
buf BUF1 (N11616, N11587);
nand NAND3 (N11617, N11616, N4258, N2356);
nor NOR4 (N11618, N11605, N5140, N6881, N317);
or OR2 (N11619, N11613, N8563);
buf BUF1 (N11620, N11617);
xor XOR2 (N11621, N11608, N11035);
and AND2 (N11622, N11620, N8321);
nor NOR2 (N11623, N11619, N4757);
nand NAND4 (N11624, N11621, N8509, N1208, N7522);
xor XOR2 (N11625, N11622, N2795);
nor NOR2 (N11626, N11614, N3431);
and AND3 (N11627, N11612, N6389, N5868);
and AND4 (N11628, N11610, N9424, N5873, N7058);
not NOT1 (N11629, N11623);
xor XOR2 (N11630, N11625, N5877);
nor NOR3 (N11631, N11630, N3134, N6606);
xor XOR2 (N11632, N11629, N117);
not NOT1 (N11633, N11627);
buf BUF1 (N11634, N11633);
or OR3 (N11635, N11632, N1418, N5270);
not NOT1 (N11636, N11634);
or OR2 (N11637, N11631, N8350);
nor NOR4 (N11638, N11626, N2016, N1530, N4738);
buf BUF1 (N11639, N11637);
or OR3 (N11640, N11635, N9527, N2237);
nand NAND2 (N11641, N11615, N7968);
not NOT1 (N11642, N11641);
xor XOR2 (N11643, N11624, N11306);
not NOT1 (N11644, N11618);
nand NAND4 (N11645, N11644, N7037, N5888, N7735);
buf BUF1 (N11646, N11639);
nor NOR4 (N11647, N11636, N5873, N11365, N2334);
buf BUF1 (N11648, N11628);
not NOT1 (N11649, N11646);
buf BUF1 (N11650, N11601);
nand NAND2 (N11651, N11649, N9161);
buf BUF1 (N11652, N11650);
and AND4 (N11653, N11638, N5870, N8140, N7339);
and AND2 (N11654, N11651, N129);
and AND2 (N11655, N11648, N5513);
nor NOR2 (N11656, N11655, N11614);
or OR4 (N11657, N11654, N8634, N385, N10229);
not NOT1 (N11658, N11595);
or OR4 (N11659, N11642, N2238, N5892, N6957);
nor NOR3 (N11660, N11643, N80, N378);
buf BUF1 (N11661, N11660);
nand NAND3 (N11662, N11659, N8333, N4536);
xor XOR2 (N11663, N11653, N10902);
or OR2 (N11664, N11658, N9964);
buf BUF1 (N11665, N11661);
buf BUF1 (N11666, N11657);
or OR3 (N11667, N11647, N1024, N9488);
and AND3 (N11668, N11640, N9699, N7232);
and AND4 (N11669, N11656, N7619, N6680, N3159);
or OR3 (N11670, N11645, N10405, N8210);
nand NAND2 (N11671, N11662, N10707);
nor NOR3 (N11672, N11663, N7656, N798);
buf BUF1 (N11673, N11669);
nand NAND3 (N11674, N11673, N3779, N5094);
xor XOR2 (N11675, N11664, N5465);
xor XOR2 (N11676, N11675, N1826);
not NOT1 (N11677, N11672);
nor NOR3 (N11678, N11676, N545, N10057);
not NOT1 (N11679, N11670);
not NOT1 (N11680, N11666);
buf BUF1 (N11681, N11680);
nor NOR3 (N11682, N11678, N1618, N10465);
xor XOR2 (N11683, N11682, N10134);
buf BUF1 (N11684, N11681);
xor XOR2 (N11685, N11668, N10909);
and AND4 (N11686, N11679, N6777, N5259, N4357);
not NOT1 (N11687, N11684);
nand NAND2 (N11688, N11686, N2210);
not NOT1 (N11689, N11665);
and AND2 (N11690, N11674, N9656);
xor XOR2 (N11691, N11688, N198);
nand NAND2 (N11692, N11683, N10738);
nand NAND4 (N11693, N11690, N9413, N10990, N7569);
nand NAND4 (N11694, N11685, N3883, N6313, N100);
and AND2 (N11695, N11652, N1380);
not NOT1 (N11696, N11692);
buf BUF1 (N11697, N11689);
not NOT1 (N11698, N11693);
nand NAND4 (N11699, N11667, N6351, N1918, N10586);
buf BUF1 (N11700, N11671);
nand NAND2 (N11701, N11696, N9134);
and AND2 (N11702, N11677, N2965);
and AND2 (N11703, N11700, N10269);
or OR3 (N11704, N11694, N8111, N3113);
and AND4 (N11705, N11691, N7254, N10087, N2530);
not NOT1 (N11706, N11704);
xor XOR2 (N11707, N11695, N1862);
not NOT1 (N11708, N11703);
nor NOR2 (N11709, N11701, N8083);
not NOT1 (N11710, N11702);
and AND2 (N11711, N11707, N8891);
not NOT1 (N11712, N11710);
and AND4 (N11713, N11687, N9564, N4990, N2238);
xor XOR2 (N11714, N11698, N6797);
not NOT1 (N11715, N11714);
and AND2 (N11716, N11712, N3060);
xor XOR2 (N11717, N11716, N6535);
not NOT1 (N11718, N11697);
or OR2 (N11719, N11699, N2663);
or OR2 (N11720, N11706, N3099);
nand NAND2 (N11721, N11709, N8057);
or OR3 (N11722, N11720, N10214, N9079);
not NOT1 (N11723, N11718);
or OR2 (N11724, N11711, N11392);
xor XOR2 (N11725, N11715, N11063);
or OR3 (N11726, N11719, N1499, N751);
nand NAND2 (N11727, N11717, N8944);
nor NOR4 (N11728, N11723, N2154, N1166, N237);
nand NAND3 (N11729, N11727, N7543, N2093);
buf BUF1 (N11730, N11729);
nand NAND4 (N11731, N11725, N10715, N8856, N4594);
or OR3 (N11732, N11728, N7763, N3831);
and AND2 (N11733, N11726, N4545);
or OR4 (N11734, N11713, N6874, N8330, N2783);
nand NAND2 (N11735, N11732, N464);
nor NOR3 (N11736, N11722, N10643, N8978);
nor NOR3 (N11737, N11731, N4477, N5203);
nor NOR2 (N11738, N11734, N9776);
and AND4 (N11739, N11724, N4295, N3235, N266);
nand NAND2 (N11740, N11733, N954);
xor XOR2 (N11741, N11737, N3607);
nor NOR2 (N11742, N11739, N5479);
nor NOR2 (N11743, N11705, N5547);
not NOT1 (N11744, N11742);
and AND2 (N11745, N11721, N1255);
buf BUF1 (N11746, N11730);
nand NAND4 (N11747, N11745, N4320, N6000, N10148);
not NOT1 (N11748, N11740);
buf BUF1 (N11749, N11747);
xor XOR2 (N11750, N11738, N9381);
nand NAND3 (N11751, N11708, N2974, N1196);
nand NAND4 (N11752, N11751, N155, N16, N1407);
xor XOR2 (N11753, N11741, N11264);
nand NAND4 (N11754, N11735, N6786, N11331, N7810);
or OR3 (N11755, N11749, N9194, N9492);
xor XOR2 (N11756, N11744, N845);
xor XOR2 (N11757, N11746, N1293);
nand NAND3 (N11758, N11756, N1091, N1009);
not NOT1 (N11759, N11758);
nor NOR4 (N11760, N11748, N7196, N9756, N499);
xor XOR2 (N11761, N11760, N7215);
buf BUF1 (N11762, N11761);
and AND3 (N11763, N11736, N1200, N1933);
buf BUF1 (N11764, N11743);
not NOT1 (N11765, N11764);
and AND3 (N11766, N11754, N5956, N9350);
buf BUF1 (N11767, N11763);
buf BUF1 (N11768, N11767);
or OR3 (N11769, N11753, N5009, N6812);
nand NAND2 (N11770, N11759, N6117);
and AND3 (N11771, N11750, N2464, N11316);
xor XOR2 (N11772, N11770, N4398);
nand NAND4 (N11773, N11768, N8929, N4385, N8966);
buf BUF1 (N11774, N11765);
nor NOR3 (N11775, N11774, N2636, N1967);
buf BUF1 (N11776, N11755);
xor XOR2 (N11777, N11766, N10611);
xor XOR2 (N11778, N11769, N1312);
or OR2 (N11779, N11762, N10117);
or OR4 (N11780, N11752, N1656, N4131, N5902);
and AND4 (N11781, N11780, N8054, N6413, N2721);
buf BUF1 (N11782, N11772);
or OR3 (N11783, N11782, N9273, N30);
buf BUF1 (N11784, N11771);
nand NAND4 (N11785, N11776, N9529, N759, N10770);
xor XOR2 (N11786, N11775, N6562);
not NOT1 (N11787, N11786);
or OR4 (N11788, N11778, N10526, N5004, N10327);
buf BUF1 (N11789, N11788);
nor NOR2 (N11790, N11787, N8615);
and AND3 (N11791, N11781, N3754, N4527);
not NOT1 (N11792, N11777);
nor NOR4 (N11793, N11785, N2493, N4070, N7936);
nand NAND4 (N11794, N11791, N11316, N11132, N6854);
not NOT1 (N11795, N11792);
buf BUF1 (N11796, N11757);
and AND3 (N11797, N11779, N11078, N2899);
not NOT1 (N11798, N11797);
buf BUF1 (N11799, N11798);
buf BUF1 (N11800, N11783);
nor NOR2 (N11801, N11796, N9146);
buf BUF1 (N11802, N11784);
and AND4 (N11803, N11799, N84, N1469, N4541);
or OR3 (N11804, N11803, N1402, N6830);
nor NOR3 (N11805, N11794, N723, N10138);
nand NAND3 (N11806, N11802, N5650, N1800);
not NOT1 (N11807, N11805);
xor XOR2 (N11808, N11790, N1226);
and AND2 (N11809, N11806, N1808);
and AND2 (N11810, N11808, N6445);
not NOT1 (N11811, N11773);
not NOT1 (N11812, N11811);
nor NOR3 (N11813, N11789, N1582, N925);
or OR2 (N11814, N11813, N3247);
not NOT1 (N11815, N11795);
buf BUF1 (N11816, N11793);
buf BUF1 (N11817, N11814);
xor XOR2 (N11818, N11817, N252);
and AND4 (N11819, N11812, N29, N5617, N9005);
nand NAND3 (N11820, N11804, N2266, N8990);
nand NAND3 (N11821, N11801, N3439, N7583);
or OR3 (N11822, N11816, N7454, N6354);
not NOT1 (N11823, N11820);
nor NOR2 (N11824, N11822, N11368);
or OR2 (N11825, N11821, N8486);
buf BUF1 (N11826, N11823);
or OR3 (N11827, N11818, N6527, N7667);
not NOT1 (N11828, N11826);
and AND3 (N11829, N11810, N3302, N11143);
and AND2 (N11830, N11825, N3260);
nor NOR2 (N11831, N11800, N9500);
xor XOR2 (N11832, N11827, N5691);
xor XOR2 (N11833, N11832, N11529);
nor NOR3 (N11834, N11833, N5571, N6201);
or OR2 (N11835, N11807, N1334);
nor NOR2 (N11836, N11824, N6273);
not NOT1 (N11837, N11834);
or OR4 (N11838, N11836, N7024, N8245, N7419);
not NOT1 (N11839, N11819);
nand NAND4 (N11840, N11809, N2312, N1791, N10707);
nor NOR3 (N11841, N11835, N400, N6885);
nand NAND2 (N11842, N11838, N2292);
buf BUF1 (N11843, N11841);
nand NAND2 (N11844, N11829, N376);
and AND3 (N11845, N11839, N8796, N11119);
xor XOR2 (N11846, N11843, N10077);
or OR4 (N11847, N11831, N10791, N5351, N133);
and AND3 (N11848, N11844, N6786, N8662);
buf BUF1 (N11849, N11830);
or OR3 (N11850, N11845, N6759, N1543);
buf BUF1 (N11851, N11848);
buf BUF1 (N11852, N11828);
buf BUF1 (N11853, N11837);
and AND2 (N11854, N11852, N2759);
not NOT1 (N11855, N11842);
buf BUF1 (N11856, N11847);
xor XOR2 (N11857, N11855, N5803);
buf BUF1 (N11858, N11851);
nor NOR4 (N11859, N11857, N11083, N11052, N11409);
buf BUF1 (N11860, N11858);
not NOT1 (N11861, N11846);
and AND2 (N11862, N11840, N10096);
buf BUF1 (N11863, N11856);
nor NOR3 (N11864, N11861, N3452, N7877);
and AND4 (N11865, N11815, N8469, N8258, N6885);
nor NOR3 (N11866, N11864, N9859, N2073);
not NOT1 (N11867, N11862);
nor NOR2 (N11868, N11866, N8909);
not NOT1 (N11869, N11853);
and AND3 (N11870, N11860, N9275, N8070);
nor NOR3 (N11871, N11869, N7070, N6180);
buf BUF1 (N11872, N11850);
nor NOR4 (N11873, N11868, N1325, N10895, N5042);
nor NOR4 (N11874, N11871, N285, N1, N3384);
or OR3 (N11875, N11859, N9192, N5803);
nand NAND2 (N11876, N11874, N9878);
and AND2 (N11877, N11876, N3899);
nor NOR4 (N11878, N11875, N11621, N8186, N84);
buf BUF1 (N11879, N11863);
xor XOR2 (N11880, N11849, N7855);
and AND2 (N11881, N11870, N2700);
xor XOR2 (N11882, N11872, N9184);
not NOT1 (N11883, N11882);
or OR3 (N11884, N11879, N397, N1108);
not NOT1 (N11885, N11881);
nand NAND4 (N11886, N11867, N325, N1516, N6355);
nand NAND2 (N11887, N11885, N8965);
and AND4 (N11888, N11877, N10138, N7079, N7332);
xor XOR2 (N11889, N11878, N11833);
nor NOR4 (N11890, N11873, N11729, N3163, N8597);
nand NAND4 (N11891, N11884, N6697, N2880, N10723);
and AND2 (N11892, N11888, N11756);
nor NOR2 (N11893, N11890, N9127);
or OR4 (N11894, N11880, N8058, N11830, N8164);
or OR2 (N11895, N11893, N1771);
and AND4 (N11896, N11886, N11674, N9457, N2197);
and AND2 (N11897, N11891, N6549);
nor NOR2 (N11898, N11889, N8833);
nor NOR3 (N11899, N11896, N4516, N570);
and AND3 (N11900, N11895, N7115, N6913);
nand NAND3 (N11901, N11898, N6775, N8283);
buf BUF1 (N11902, N11897);
buf BUF1 (N11903, N11883);
or OR2 (N11904, N11894, N206);
not NOT1 (N11905, N11903);
nor NOR3 (N11906, N11901, N11699, N10068);
xor XOR2 (N11907, N11854, N1396);
not NOT1 (N11908, N11902);
nor NOR3 (N11909, N11899, N10611, N10529);
and AND4 (N11910, N11887, N11645, N11447, N11879);
xor XOR2 (N11911, N11905, N7743);
not NOT1 (N11912, N11906);
not NOT1 (N11913, N11907);
xor XOR2 (N11914, N11908, N8594);
nand NAND3 (N11915, N11910, N6468, N3355);
and AND4 (N11916, N11915, N1327, N166, N10457);
xor XOR2 (N11917, N11892, N5821);
nor NOR4 (N11918, N11916, N1841, N5914, N2749);
nand NAND3 (N11919, N11912, N1761, N7930);
not NOT1 (N11920, N11900);
and AND4 (N11921, N11917, N9602, N88, N6995);
xor XOR2 (N11922, N11918, N6609);
buf BUF1 (N11923, N11913);
and AND2 (N11924, N11914, N3658);
xor XOR2 (N11925, N11904, N4782);
and AND4 (N11926, N11920, N518, N8590, N9714);
nand NAND3 (N11927, N11919, N9603, N7384);
nor NOR2 (N11928, N11911, N2224);
and AND4 (N11929, N11928, N2648, N4080, N5801);
xor XOR2 (N11930, N11925, N2615);
and AND3 (N11931, N11923, N9136, N9459);
xor XOR2 (N11932, N11865, N6376);
and AND3 (N11933, N11930, N8999, N10446);
nor NOR2 (N11934, N11932, N8027);
nor NOR2 (N11935, N11922, N4476);
nor NOR2 (N11936, N11926, N7466);
nor NOR3 (N11937, N11936, N9049, N1362);
not NOT1 (N11938, N11934);
buf BUF1 (N11939, N11933);
nand NAND2 (N11940, N11938, N10796);
xor XOR2 (N11941, N11937, N2676);
buf BUF1 (N11942, N11924);
and AND2 (N11943, N11927, N11173);
xor XOR2 (N11944, N11941, N3829);
and AND3 (N11945, N11929, N8128, N10419);
not NOT1 (N11946, N11943);
not NOT1 (N11947, N11921);
xor XOR2 (N11948, N11942, N11123);
nor NOR4 (N11949, N11909, N6946, N4669, N10111);
nand NAND4 (N11950, N11935, N3410, N10243, N5758);
buf BUF1 (N11951, N11945);
xor XOR2 (N11952, N11947, N3042);
nand NAND4 (N11953, N11950, N3566, N1775, N6402);
buf BUF1 (N11954, N11948);
not NOT1 (N11955, N11946);
and AND2 (N11956, N11954, N3817);
xor XOR2 (N11957, N11940, N2160);
not NOT1 (N11958, N11953);
not NOT1 (N11959, N11931);
xor XOR2 (N11960, N11939, N2599);
or OR2 (N11961, N11960, N1797);
buf BUF1 (N11962, N11959);
and AND4 (N11963, N11952, N3218, N4221, N3345);
buf BUF1 (N11964, N11962);
and AND3 (N11965, N11961, N5334, N1901);
or OR2 (N11966, N11957, N8776);
buf BUF1 (N11967, N11963);
buf BUF1 (N11968, N11958);
buf BUF1 (N11969, N11955);
nor NOR2 (N11970, N11956, N10959);
xor XOR2 (N11971, N11944, N7798);
not NOT1 (N11972, N11968);
buf BUF1 (N11973, N11970);
not NOT1 (N11974, N11964);
buf BUF1 (N11975, N11972);
and AND2 (N11976, N11967, N5677);
not NOT1 (N11977, N11971);
and AND4 (N11978, N11969, N10878, N2510, N6196);
or OR3 (N11979, N11966, N5712, N8335);
xor XOR2 (N11980, N11973, N11340);
and AND2 (N11981, N11965, N207);
nor NOR4 (N11982, N11980, N5109, N6327, N9963);
xor XOR2 (N11983, N11981, N8507);
and AND3 (N11984, N11978, N424, N9356);
and AND3 (N11985, N11982, N3378, N10612);
nand NAND4 (N11986, N11977, N8477, N122, N1399);
not NOT1 (N11987, N11984);
nand NAND3 (N11988, N11949, N11054, N4811);
xor XOR2 (N11989, N11975, N9182);
nand NAND4 (N11990, N11989, N1004, N6543, N7978);
not NOT1 (N11991, N11985);
not NOT1 (N11992, N11991);
not NOT1 (N11993, N11987);
xor XOR2 (N11994, N11986, N4448);
nand NAND3 (N11995, N11988, N5658, N6304);
not NOT1 (N11996, N11995);
not NOT1 (N11997, N11992);
not NOT1 (N11998, N11951);
xor XOR2 (N11999, N11974, N8084);
or OR4 (N12000, N11990, N8359, N9061, N3364);
nand NAND3 (N12001, N11997, N10248, N6855);
xor XOR2 (N12002, N11993, N5041);
nor NOR4 (N12003, N11979, N4624, N8069, N3676);
not NOT1 (N12004, N11976);
not NOT1 (N12005, N11994);
nor NOR4 (N12006, N11983, N1661, N4707, N607);
nor NOR2 (N12007, N12004, N9465);
or OR2 (N12008, N12007, N9651);
nor NOR3 (N12009, N12005, N11701, N155);
xor XOR2 (N12010, N12001, N11583);
and AND4 (N12011, N12000, N4846, N5365, N4130);
nor NOR2 (N12012, N12010, N9721);
not NOT1 (N12013, N12009);
or OR2 (N12014, N12012, N6987);
buf BUF1 (N12015, N12002);
nand NAND4 (N12016, N11996, N5613, N12, N9893);
or OR3 (N12017, N11999, N2822, N3573);
nor NOR3 (N12018, N12003, N5411, N2921);
not NOT1 (N12019, N12015);
or OR4 (N12020, N12013, N2972, N11335, N10745);
xor XOR2 (N12021, N12008, N2571);
xor XOR2 (N12022, N12006, N10229);
or OR4 (N12023, N12011, N8511, N7180, N190);
buf BUF1 (N12024, N11998);
and AND2 (N12025, N12020, N2179);
buf BUF1 (N12026, N12014);
nand NAND3 (N12027, N12018, N3667, N10170);
or OR2 (N12028, N12019, N8563);
xor XOR2 (N12029, N12017, N2382);
buf BUF1 (N12030, N12023);
or OR3 (N12031, N12028, N543, N10476);
and AND4 (N12032, N12027, N446, N8742, N6043);
buf BUF1 (N12033, N12024);
nand NAND3 (N12034, N12030, N3795, N9393);
xor XOR2 (N12035, N12033, N2484);
and AND2 (N12036, N12031, N3180);
nand NAND2 (N12037, N12032, N7922);
not NOT1 (N12038, N12022);
nand NAND4 (N12039, N12038, N6823, N8905, N845);
not NOT1 (N12040, N12025);
not NOT1 (N12041, N12021);
and AND4 (N12042, N12029, N5105, N3646, N6466);
and AND2 (N12043, N12037, N4557);
xor XOR2 (N12044, N12036, N8065);
nand NAND2 (N12045, N12035, N9126);
nor NOR3 (N12046, N12016, N8022, N4959);
nand NAND4 (N12047, N12044, N4399, N3647, N5870);
buf BUF1 (N12048, N12047);
or OR2 (N12049, N12043, N2735);
and AND4 (N12050, N12040, N5437, N5157, N1223);
xor XOR2 (N12051, N12039, N6045);
not NOT1 (N12052, N12026);
nor NOR4 (N12053, N12051, N8002, N9249, N6910);
xor XOR2 (N12054, N12041, N7562);
and AND2 (N12055, N12034, N8675);
buf BUF1 (N12056, N12049);
and AND2 (N12057, N12056, N3250);
and AND2 (N12058, N12055, N403);
nand NAND2 (N12059, N12054, N419);
nand NAND2 (N12060, N12057, N10869);
not NOT1 (N12061, N12052);
nand NAND2 (N12062, N12053, N7151);
buf BUF1 (N12063, N12045);
nand NAND4 (N12064, N12059, N351, N16, N4670);
and AND3 (N12065, N12063, N8037, N6092);
nand NAND3 (N12066, N12064, N2670, N7034);
and AND2 (N12067, N12058, N8640);
or OR2 (N12068, N12065, N11360);
nand NAND4 (N12069, N12042, N4876, N7052, N8766);
and AND2 (N12070, N12046, N8480);
not NOT1 (N12071, N12060);
buf BUF1 (N12072, N12068);
buf BUF1 (N12073, N12072);
buf BUF1 (N12074, N12048);
nand NAND4 (N12075, N12066, N11920, N5736, N9462);
xor XOR2 (N12076, N12071, N4681);
nand NAND4 (N12077, N12074, N2845, N1370, N837);
and AND3 (N12078, N12070, N436, N3701);
and AND3 (N12079, N12050, N6488, N5865);
nor NOR4 (N12080, N12079, N24, N2756, N6199);
or OR3 (N12081, N12076, N928, N10885);
nor NOR4 (N12082, N12073, N1898, N8674, N337);
nor NOR2 (N12083, N12077, N2340);
xor XOR2 (N12084, N12062, N944);
nand NAND4 (N12085, N12069, N3157, N8992, N7015);
buf BUF1 (N12086, N12085);
or OR2 (N12087, N12067, N3680);
xor XOR2 (N12088, N12083, N3739);
and AND2 (N12089, N12086, N3691);
nor NOR4 (N12090, N12078, N7359, N4210, N3303);
nand NAND3 (N12091, N12081, N4959, N3572);
or OR2 (N12092, N12082, N3546);
xor XOR2 (N12093, N12089, N2213);
xor XOR2 (N12094, N12091, N9249);
xor XOR2 (N12095, N12061, N6940);
or OR2 (N12096, N12084, N11365);
nor NOR4 (N12097, N12080, N6048, N9496, N7265);
not NOT1 (N12098, N12096);
or OR3 (N12099, N12088, N9424, N5323);
or OR3 (N12100, N12075, N6207, N3479);
nand NAND3 (N12101, N12094, N5629, N6773);
nor NOR4 (N12102, N12090, N10867, N5608, N8501);
nor NOR3 (N12103, N12093, N9326, N1392);
not NOT1 (N12104, N12101);
nand NAND2 (N12105, N12092, N8945);
nor NOR3 (N12106, N12087, N11805, N6815);
or OR4 (N12107, N12104, N4856, N3439, N9028);
nand NAND4 (N12108, N12099, N4970, N9409, N4874);
buf BUF1 (N12109, N12097);
nand NAND2 (N12110, N12108, N10323);
buf BUF1 (N12111, N12100);
nor NOR4 (N12112, N12103, N11143, N4895, N9774);
xor XOR2 (N12113, N12106, N11571);
nor NOR2 (N12114, N12105, N9656);
xor XOR2 (N12115, N12111, N2967);
or OR4 (N12116, N12098, N3861, N5749, N2897);
nand NAND4 (N12117, N12113, N11055, N10205, N8021);
xor XOR2 (N12118, N12114, N760);
buf BUF1 (N12119, N12118);
nand NAND2 (N12120, N12095, N1801);
not NOT1 (N12121, N12110);
nor NOR4 (N12122, N12117, N10093, N4084, N5607);
or OR3 (N12123, N12109, N7414, N8388);
or OR4 (N12124, N12121, N7119, N1736, N1750);
xor XOR2 (N12125, N12124, N12015);
not NOT1 (N12126, N12122);
nor NOR2 (N12127, N12119, N3001);
nor NOR2 (N12128, N12125, N5853);
nor NOR2 (N12129, N12128, N8990);
nor NOR4 (N12130, N12123, N6918, N2770, N5047);
buf BUF1 (N12131, N12129);
buf BUF1 (N12132, N12131);
or OR3 (N12133, N12116, N10274, N8171);
nor NOR3 (N12134, N12127, N5365, N10709);
xor XOR2 (N12135, N12130, N4992);
not NOT1 (N12136, N12115);
buf BUF1 (N12137, N12112);
or OR3 (N12138, N12120, N7436, N3563);
and AND2 (N12139, N12107, N1921);
and AND3 (N12140, N12102, N1665, N8822);
and AND2 (N12141, N12134, N3355);
xor XOR2 (N12142, N12139, N8487);
or OR2 (N12143, N12133, N360);
or OR4 (N12144, N12136, N5154, N5663, N1639);
buf BUF1 (N12145, N12135);
and AND4 (N12146, N12132, N9420, N7575, N6719);
and AND3 (N12147, N12143, N4891, N9533);
buf BUF1 (N12148, N12141);
or OR2 (N12149, N12144, N10231);
xor XOR2 (N12150, N12142, N5766);
nor NOR4 (N12151, N12145, N11379, N11492, N920);
xor XOR2 (N12152, N12140, N4607);
nor NOR3 (N12153, N12152, N8917, N3774);
nor NOR4 (N12154, N12146, N1089, N8622, N5757);
nand NAND4 (N12155, N12149, N2096, N12143, N5115);
not NOT1 (N12156, N12147);
nand NAND4 (N12157, N12150, N2281, N8756, N7683);
nor NOR2 (N12158, N12154, N748);
and AND3 (N12159, N12153, N7918, N5638);
buf BUF1 (N12160, N12151);
buf BUF1 (N12161, N12155);
nand NAND2 (N12162, N12161, N3060);
buf BUF1 (N12163, N12157);
and AND3 (N12164, N12126, N1097, N6442);
or OR2 (N12165, N12138, N8742);
nor NOR4 (N12166, N12137, N9420, N3030, N11225);
or OR3 (N12167, N12159, N7731, N280);
and AND2 (N12168, N12164, N6490);
nand NAND3 (N12169, N12165, N7049, N2721);
buf BUF1 (N12170, N12163);
and AND4 (N12171, N12148, N5830, N9125, N2506);
xor XOR2 (N12172, N12168, N8531);
nand NAND4 (N12173, N12171, N4907, N3166, N3575);
or OR4 (N12174, N12172, N8755, N2904, N7400);
not NOT1 (N12175, N12156);
and AND3 (N12176, N12170, N5284, N5154);
xor XOR2 (N12177, N12158, N1690);
or OR3 (N12178, N12169, N2000, N4166);
nand NAND4 (N12179, N12177, N10958, N10163, N11044);
nor NOR2 (N12180, N12178, N6893);
nor NOR4 (N12181, N12162, N6530, N2033, N1942);
nand NAND2 (N12182, N12179, N10910);
or OR3 (N12183, N12180, N734, N5287);
buf BUF1 (N12184, N12183);
and AND4 (N12185, N12182, N7042, N10044, N1030);
buf BUF1 (N12186, N12184);
buf BUF1 (N12187, N12181);
xor XOR2 (N12188, N12185, N4996);
and AND4 (N12189, N12188, N10977, N9024, N9674);
xor XOR2 (N12190, N12167, N6413);
nor NOR3 (N12191, N12166, N11852, N2518);
nand NAND2 (N12192, N12175, N1467);
nor NOR4 (N12193, N12176, N5869, N1154, N11927);
buf BUF1 (N12194, N12192);
or OR3 (N12195, N12174, N8038, N8362);
and AND3 (N12196, N12191, N1593, N7094);
not NOT1 (N12197, N12160);
nor NOR2 (N12198, N12196, N10440);
nand NAND3 (N12199, N12187, N5238, N8700);
nor NOR2 (N12200, N12198, N3535);
and AND4 (N12201, N12195, N2344, N11428, N6791);
nor NOR3 (N12202, N12199, N8731, N2159);
buf BUF1 (N12203, N12189);
buf BUF1 (N12204, N12186);
not NOT1 (N12205, N12190);
not NOT1 (N12206, N12205);
nand NAND4 (N12207, N12193, N9983, N4276, N8251);
or OR4 (N12208, N12207, N10925, N12185, N10239);
nand NAND3 (N12209, N12203, N8281, N2992);
xor XOR2 (N12210, N12200, N8044);
buf BUF1 (N12211, N12204);
nand NAND3 (N12212, N12197, N5003, N4812);
buf BUF1 (N12213, N12209);
not NOT1 (N12214, N12202);
nor NOR3 (N12215, N12173, N5174, N3649);
nand NAND3 (N12216, N12206, N3024, N11779);
nor NOR3 (N12217, N12215, N505, N2913);
nor NOR2 (N12218, N12214, N4444);
not NOT1 (N12219, N12211);
nand NAND4 (N12220, N12217, N8551, N9465, N9809);
nor NOR3 (N12221, N12208, N8954, N2203);
nand NAND3 (N12222, N12210, N7117, N5032);
xor XOR2 (N12223, N12221, N4326);
buf BUF1 (N12224, N12212);
buf BUF1 (N12225, N12194);
and AND2 (N12226, N12213, N11916);
buf BUF1 (N12227, N12222);
nor NOR3 (N12228, N12220, N805, N5583);
xor XOR2 (N12229, N12219, N10406);
nand NAND2 (N12230, N12218, N81);
xor XOR2 (N12231, N12225, N1692);
nor NOR3 (N12232, N12230, N1457, N4901);
nand NAND4 (N12233, N12232, N10138, N8667, N3865);
xor XOR2 (N12234, N12216, N3314);
buf BUF1 (N12235, N12234);
or OR4 (N12236, N12228, N11723, N5827, N10099);
not NOT1 (N12237, N12201);
nand NAND2 (N12238, N12223, N4488);
and AND2 (N12239, N12227, N3744);
buf BUF1 (N12240, N12239);
not NOT1 (N12241, N12224);
xor XOR2 (N12242, N12235, N9864);
xor XOR2 (N12243, N12242, N3611);
nor NOR2 (N12244, N12226, N1952);
xor XOR2 (N12245, N12244, N3891);
and AND3 (N12246, N12241, N6501, N10551);
xor XOR2 (N12247, N12229, N3827);
not NOT1 (N12248, N12236);
xor XOR2 (N12249, N12245, N2507);
or OR4 (N12250, N12246, N3728, N6336, N968);
xor XOR2 (N12251, N12250, N10728);
and AND4 (N12252, N12238, N85, N3589, N2633);
xor XOR2 (N12253, N12252, N9891);
or OR3 (N12254, N12237, N8754, N11902);
xor XOR2 (N12255, N12233, N3777);
nand NAND4 (N12256, N12248, N9522, N963, N5560);
nor NOR3 (N12257, N12256, N10429, N399);
xor XOR2 (N12258, N12251, N11005);
not NOT1 (N12259, N12257);
and AND3 (N12260, N12243, N7637, N9431);
not NOT1 (N12261, N12247);
xor XOR2 (N12262, N12259, N9303);
not NOT1 (N12263, N12240);
buf BUF1 (N12264, N12255);
xor XOR2 (N12265, N12263, N1864);
xor XOR2 (N12266, N12261, N7200);
or OR3 (N12267, N12253, N2273, N3688);
and AND2 (N12268, N12265, N5196);
nand NAND3 (N12269, N12262, N1203, N6542);
and AND2 (N12270, N12267, N6200);
and AND4 (N12271, N12264, N10717, N11411, N272);
nand NAND3 (N12272, N12268, N7287, N5358);
buf BUF1 (N12273, N12231);
buf BUF1 (N12274, N12273);
not NOT1 (N12275, N12258);
not NOT1 (N12276, N12254);
or OR4 (N12277, N12274, N8158, N10375, N2058);
or OR3 (N12278, N12260, N1100, N12034);
not NOT1 (N12279, N12271);
and AND2 (N12280, N12249, N4548);
and AND2 (N12281, N12272, N10662);
and AND3 (N12282, N12275, N541, N7608);
or OR4 (N12283, N12269, N9760, N4177, N8760);
not NOT1 (N12284, N12280);
or OR4 (N12285, N12278, N10031, N6591, N1139);
not NOT1 (N12286, N12284);
or OR3 (N12287, N12270, N10392, N725);
buf BUF1 (N12288, N12266);
nor NOR4 (N12289, N12283, N8344, N2579, N10007);
not NOT1 (N12290, N12279);
nor NOR3 (N12291, N12285, N11885, N8890);
nor NOR4 (N12292, N12289, N6249, N5799, N1081);
nor NOR2 (N12293, N12287, N10147);
or OR2 (N12294, N12277, N268);
nand NAND2 (N12295, N12291, N949);
not NOT1 (N12296, N12293);
nand NAND3 (N12297, N12282, N12099, N11955);
and AND3 (N12298, N12297, N1049, N1026);
nand NAND4 (N12299, N12286, N6262, N8920, N594);
not NOT1 (N12300, N12294);
xor XOR2 (N12301, N12292, N10472);
nand NAND4 (N12302, N12296, N957, N6636, N787);
nor NOR4 (N12303, N12299, N9754, N4413, N7366);
nand NAND3 (N12304, N12300, N8056, N5781);
buf BUF1 (N12305, N12304);
nor NOR3 (N12306, N12302, N2328, N1305);
nor NOR3 (N12307, N12276, N470, N1193);
or OR4 (N12308, N12290, N8098, N5923, N5029);
or OR2 (N12309, N12306, N7281);
nand NAND4 (N12310, N12298, N1318, N563, N10614);
and AND3 (N12311, N12308, N1412, N5149);
or OR4 (N12312, N12310, N1921, N1009, N4616);
or OR2 (N12313, N12311, N4582);
xor XOR2 (N12314, N12295, N6805);
nand NAND2 (N12315, N12309, N696);
nor NOR4 (N12316, N12315, N9712, N4499, N1546);
nand NAND2 (N12317, N12316, N5573);
not NOT1 (N12318, N12314);
not NOT1 (N12319, N12318);
buf BUF1 (N12320, N12288);
and AND3 (N12321, N12320, N2456, N749);
xor XOR2 (N12322, N12303, N3127);
or OR3 (N12323, N12319, N1167, N4548);
and AND3 (N12324, N12313, N8301, N1772);
and AND4 (N12325, N12324, N2083, N6363, N12035);
or OR4 (N12326, N12305, N415, N3428, N7424);
or OR4 (N12327, N12322, N6722, N10021, N6613);
not NOT1 (N12328, N12323);
or OR3 (N12329, N12321, N3542, N2757);
nor NOR4 (N12330, N12307, N4707, N1349, N11222);
nand NAND4 (N12331, N12325, N11670, N1937, N9863);
buf BUF1 (N12332, N12328);
buf BUF1 (N12333, N12329);
or OR2 (N12334, N12327, N5143);
nand NAND4 (N12335, N12326, N9785, N11998, N7191);
xor XOR2 (N12336, N12281, N9423);
xor XOR2 (N12337, N12336, N11080);
buf BUF1 (N12338, N12333);
nor NOR4 (N12339, N12332, N4133, N413, N9966);
xor XOR2 (N12340, N12337, N4358);
xor XOR2 (N12341, N12334, N2585);
buf BUF1 (N12342, N12301);
or OR4 (N12343, N12312, N2721, N3661, N2296);
buf BUF1 (N12344, N12338);
or OR2 (N12345, N12340, N9601);
not NOT1 (N12346, N12345);
nand NAND4 (N12347, N12344, N10983, N3688, N2323);
nand NAND3 (N12348, N12341, N2403, N2818);
or OR4 (N12349, N12342, N3246, N11389, N8066);
not NOT1 (N12350, N12348);
and AND4 (N12351, N12347, N2370, N3401, N884);
nor NOR4 (N12352, N12335, N4671, N11466, N7992);
or OR2 (N12353, N12346, N6877);
buf BUF1 (N12354, N12352);
not NOT1 (N12355, N12349);
nand NAND3 (N12356, N12343, N6896, N1944);
nor NOR3 (N12357, N12353, N4029, N5249);
nor NOR2 (N12358, N12350, N12134);
not NOT1 (N12359, N12356);
and AND3 (N12360, N12351, N3759, N10352);
and AND3 (N12361, N12355, N474, N6168);
nand NAND3 (N12362, N12331, N1132, N12245);
or OR4 (N12363, N12357, N10521, N6954, N2895);
or OR4 (N12364, N12361, N8293, N7513, N6870);
nand NAND2 (N12365, N12339, N1155);
and AND3 (N12366, N12364, N3374, N5392);
xor XOR2 (N12367, N12365, N3051);
xor XOR2 (N12368, N12362, N6272);
buf BUF1 (N12369, N12317);
buf BUF1 (N12370, N12363);
not NOT1 (N12371, N12358);
nor NOR3 (N12372, N12359, N2018, N3068);
xor XOR2 (N12373, N12366, N8000);
or OR4 (N12374, N12368, N5957, N7843, N7764);
nand NAND2 (N12375, N12367, N6773);
nand NAND3 (N12376, N12330, N4979, N1284);
not NOT1 (N12377, N12369);
xor XOR2 (N12378, N12373, N8677);
buf BUF1 (N12379, N12376);
buf BUF1 (N12380, N12354);
nand NAND2 (N12381, N12370, N716);
xor XOR2 (N12382, N12377, N5469);
nand NAND4 (N12383, N12360, N4880, N4309, N11201);
xor XOR2 (N12384, N12374, N5860);
nor NOR3 (N12385, N12371, N10371, N9012);
not NOT1 (N12386, N12379);
nand NAND4 (N12387, N12380, N3644, N9951, N9710);
or OR2 (N12388, N12383, N3855);
nor NOR4 (N12389, N12378, N1325, N4617, N422);
not NOT1 (N12390, N12385);
nand NAND3 (N12391, N12387, N4990, N11733);
not NOT1 (N12392, N12384);
buf BUF1 (N12393, N12392);
not NOT1 (N12394, N12390);
not NOT1 (N12395, N12393);
xor XOR2 (N12396, N12382, N9091);
xor XOR2 (N12397, N12389, N1299);
xor XOR2 (N12398, N12386, N9335);
xor XOR2 (N12399, N12396, N1612);
nand NAND4 (N12400, N12375, N9331, N8089, N9763);
not NOT1 (N12401, N12397);
xor XOR2 (N12402, N12395, N10094);
nor NOR4 (N12403, N12388, N9889, N4924, N4209);
nand NAND2 (N12404, N12399, N4046);
nor NOR2 (N12405, N12402, N780);
and AND2 (N12406, N12381, N8944);
or OR4 (N12407, N12398, N4867, N3236, N8781);
and AND3 (N12408, N12405, N1437, N6751);
xor XOR2 (N12409, N12403, N9601);
nand NAND2 (N12410, N12391, N10602);
xor XOR2 (N12411, N12406, N11948);
and AND4 (N12412, N12401, N2002, N8707, N1541);
buf BUF1 (N12413, N12410);
not NOT1 (N12414, N12409);
nor NOR2 (N12415, N12400, N838);
xor XOR2 (N12416, N12413, N9067);
buf BUF1 (N12417, N12394);
xor XOR2 (N12418, N12404, N6116);
not NOT1 (N12419, N12407);
xor XOR2 (N12420, N12411, N1965);
xor XOR2 (N12421, N12412, N10781);
not NOT1 (N12422, N12420);
and AND3 (N12423, N12417, N9707, N4264);
buf BUF1 (N12424, N12372);
xor XOR2 (N12425, N12424, N2865);
xor XOR2 (N12426, N12408, N3017);
nand NAND4 (N12427, N12416, N2323, N7885, N2726);
nand NAND2 (N12428, N12427, N8971);
not NOT1 (N12429, N12419);
and AND4 (N12430, N12414, N3018, N6469, N6508);
or OR2 (N12431, N12418, N10992);
buf BUF1 (N12432, N12430);
nand NAND2 (N12433, N12428, N714);
and AND2 (N12434, N12415, N10554);
not NOT1 (N12435, N12432);
not NOT1 (N12436, N12434);
not NOT1 (N12437, N12422);
buf BUF1 (N12438, N12433);
not NOT1 (N12439, N12437);
nand NAND2 (N12440, N12423, N11773);
nor NOR3 (N12441, N12440, N9890, N3803);
and AND3 (N12442, N12436, N2413, N4261);
or OR2 (N12443, N12426, N7697);
and AND3 (N12444, N12441, N8280, N9239);
and AND4 (N12445, N12425, N5782, N8707, N847);
and AND3 (N12446, N12439, N8454, N5915);
and AND2 (N12447, N12443, N8221);
not NOT1 (N12448, N12444);
buf BUF1 (N12449, N12431);
xor XOR2 (N12450, N12442, N1195);
not NOT1 (N12451, N12438);
and AND2 (N12452, N12421, N11441);
not NOT1 (N12453, N12447);
and AND4 (N12454, N12448, N7266, N920, N7304);
not NOT1 (N12455, N12445);
and AND2 (N12456, N12446, N3354);
nor NOR3 (N12457, N12456, N11453, N6467);
buf BUF1 (N12458, N12455);
and AND4 (N12459, N12458, N7490, N2847, N10509);
not NOT1 (N12460, N12451);
xor XOR2 (N12461, N12435, N7144);
nand NAND3 (N12462, N12429, N10876, N5926);
xor XOR2 (N12463, N12454, N7962);
not NOT1 (N12464, N12450);
not NOT1 (N12465, N12461);
buf BUF1 (N12466, N12462);
and AND3 (N12467, N12463, N11239, N4443);
nor NOR3 (N12468, N12452, N9831, N10500);
nor NOR2 (N12469, N12467, N8291);
and AND2 (N12470, N12469, N5296);
nand NAND3 (N12471, N12465, N11872, N2812);
nor NOR3 (N12472, N12470, N5844, N4112);
not NOT1 (N12473, N12471);
nor NOR3 (N12474, N12449, N9423, N1764);
buf BUF1 (N12475, N12460);
not NOT1 (N12476, N12466);
not NOT1 (N12477, N12453);
buf BUF1 (N12478, N12472);
buf BUF1 (N12479, N12475);
nor NOR3 (N12480, N12477, N3275, N10480);
xor XOR2 (N12481, N12479, N4379);
nor NOR4 (N12482, N12474, N5358, N4625, N11040);
buf BUF1 (N12483, N12459);
and AND4 (N12484, N12480, N7188, N10731, N12356);
xor XOR2 (N12485, N12468, N5163);
xor XOR2 (N12486, N12482, N3036);
or OR2 (N12487, N12481, N119);
xor XOR2 (N12488, N12464, N7648);
and AND4 (N12489, N12484, N5681, N11373, N4604);
nor NOR2 (N12490, N12478, N3769);
xor XOR2 (N12491, N12457, N6910);
xor XOR2 (N12492, N12487, N10692);
nand NAND3 (N12493, N12491, N11678, N5465);
buf BUF1 (N12494, N12490);
nand NAND4 (N12495, N12492, N2014, N10039, N424);
buf BUF1 (N12496, N12494);
not NOT1 (N12497, N12493);
not NOT1 (N12498, N12497);
or OR2 (N12499, N12498, N5861);
or OR3 (N12500, N12486, N1233, N1501);
not NOT1 (N12501, N12500);
xor XOR2 (N12502, N12483, N8722);
nand NAND3 (N12503, N12488, N5746, N3007);
buf BUF1 (N12504, N12501);
not NOT1 (N12505, N12473);
buf BUF1 (N12506, N12505);
and AND3 (N12507, N12503, N2847, N7357);
buf BUF1 (N12508, N12495);
and AND4 (N12509, N12485, N9704, N5485, N5695);
and AND3 (N12510, N12509, N1941, N1193);
and AND3 (N12511, N12496, N10051, N7610);
not NOT1 (N12512, N12510);
buf BUF1 (N12513, N12507);
nor NOR2 (N12514, N12504, N9475);
xor XOR2 (N12515, N12514, N7053);
nand NAND2 (N12516, N12499, N7275);
and AND2 (N12517, N12508, N11210);
buf BUF1 (N12518, N12512);
nand NAND3 (N12519, N12518, N963, N8734);
nand NAND3 (N12520, N12476, N11260, N873);
buf BUF1 (N12521, N12520);
nand NAND2 (N12522, N12519, N2915);
not NOT1 (N12523, N12522);
nor NOR3 (N12524, N12506, N7549, N3095);
and AND2 (N12525, N12523, N9418);
or OR3 (N12526, N12515, N5610, N6034);
not NOT1 (N12527, N12526);
nand NAND2 (N12528, N12521, N10708);
and AND2 (N12529, N12513, N663);
nor NOR3 (N12530, N12527, N1530, N12294);
xor XOR2 (N12531, N12489, N9360);
nand NAND2 (N12532, N12528, N1470);
nor NOR4 (N12533, N12525, N10330, N11804, N6498);
not NOT1 (N12534, N12530);
xor XOR2 (N12535, N12531, N3454);
nand NAND2 (N12536, N12534, N6136);
not NOT1 (N12537, N12517);
not NOT1 (N12538, N12537);
or OR3 (N12539, N12535, N9779, N5434);
not NOT1 (N12540, N12529);
or OR2 (N12541, N12502, N4923);
or OR2 (N12542, N12516, N3673);
xor XOR2 (N12543, N12533, N2677);
buf BUF1 (N12544, N12524);
not NOT1 (N12545, N12541);
not NOT1 (N12546, N12536);
not NOT1 (N12547, N12543);
buf BUF1 (N12548, N12545);
xor XOR2 (N12549, N12546, N3507);
or OR3 (N12550, N12540, N4259, N2798);
xor XOR2 (N12551, N12549, N753);
xor XOR2 (N12552, N12538, N9499);
xor XOR2 (N12553, N12550, N3906);
xor XOR2 (N12554, N12547, N7657);
buf BUF1 (N12555, N12551);
nor NOR3 (N12556, N12542, N11589, N8919);
nor NOR3 (N12557, N12539, N8606, N4305);
not NOT1 (N12558, N12532);
and AND2 (N12559, N12555, N4943);
and AND3 (N12560, N12556, N5438, N8587);
not NOT1 (N12561, N12553);
xor XOR2 (N12562, N12559, N11312);
not NOT1 (N12563, N12557);
nor NOR3 (N12564, N12562, N9633, N4015);
xor XOR2 (N12565, N12558, N10024);
nand NAND2 (N12566, N12511, N1416);
xor XOR2 (N12567, N12554, N6661);
or OR4 (N12568, N12567, N761, N3489, N11940);
not NOT1 (N12569, N12568);
nor NOR4 (N12570, N12561, N4937, N11381, N7615);
or OR3 (N12571, N12563, N5239, N12396);
not NOT1 (N12572, N12566);
not NOT1 (N12573, N12564);
buf BUF1 (N12574, N12569);
or OR2 (N12575, N12574, N6780);
xor XOR2 (N12576, N12571, N2353);
or OR2 (N12577, N12575, N7807);
and AND2 (N12578, N12552, N9418);
and AND4 (N12579, N12560, N4879, N6318, N1946);
or OR4 (N12580, N12565, N9320, N2757, N9360);
nor NOR4 (N12581, N12572, N9703, N12536, N6396);
or OR3 (N12582, N12573, N9964, N12335);
buf BUF1 (N12583, N12581);
nand NAND2 (N12584, N12579, N8097);
and AND3 (N12585, N12584, N652, N1448);
xor XOR2 (N12586, N12577, N3982);
nor NOR3 (N12587, N12586, N2944, N7016);
not NOT1 (N12588, N12587);
or OR2 (N12589, N12582, N225);
not NOT1 (N12590, N12548);
buf BUF1 (N12591, N12588);
nand NAND2 (N12592, N12589, N6724);
and AND4 (N12593, N12580, N2809, N4124, N5369);
and AND2 (N12594, N12590, N10866);
or OR2 (N12595, N12594, N2917);
xor XOR2 (N12596, N12576, N5925);
not NOT1 (N12597, N12591);
and AND4 (N12598, N12578, N4254, N2288, N10794);
not NOT1 (N12599, N12544);
nand NAND2 (N12600, N12593, N7421);
not NOT1 (N12601, N12583);
buf BUF1 (N12602, N12595);
xor XOR2 (N12603, N12602, N10834);
or OR3 (N12604, N12603, N11841, N9584);
buf BUF1 (N12605, N12604);
and AND3 (N12606, N12597, N3362, N871);
xor XOR2 (N12607, N12606, N8858);
xor XOR2 (N12608, N12596, N9466);
or OR4 (N12609, N12601, N3446, N11278, N4541);
xor XOR2 (N12610, N12600, N858);
nor NOR4 (N12611, N12608, N1364, N2434, N6870);
xor XOR2 (N12612, N12599, N9381);
not NOT1 (N12613, N12570);
buf BUF1 (N12614, N12610);
or OR2 (N12615, N12585, N2886);
or OR4 (N12616, N12607, N7561, N751, N12239);
not NOT1 (N12617, N12598);
xor XOR2 (N12618, N12613, N8911);
xor XOR2 (N12619, N12611, N5754);
xor XOR2 (N12620, N12605, N11390);
nand NAND2 (N12621, N12615, N3379);
nand NAND4 (N12622, N12614, N11941, N3217, N6005);
or OR2 (N12623, N12592, N10394);
nand NAND4 (N12624, N12616, N8910, N8042, N941);
or OR3 (N12625, N12617, N4831, N354);
and AND2 (N12626, N12625, N9083);
buf BUF1 (N12627, N12612);
or OR4 (N12628, N12623, N4356, N5838, N9359);
not NOT1 (N12629, N12626);
or OR2 (N12630, N12622, N6310);
nand NAND2 (N12631, N12627, N2265);
xor XOR2 (N12632, N12618, N11904);
xor XOR2 (N12633, N12628, N5111);
xor XOR2 (N12634, N12619, N11701);
nand NAND4 (N12635, N12621, N9416, N106, N1175);
or OR3 (N12636, N12620, N5438, N11036);
nor NOR4 (N12637, N12634, N3556, N6198, N7106);
xor XOR2 (N12638, N12631, N9507);
buf BUF1 (N12639, N12609);
and AND4 (N12640, N12637, N11283, N10340, N290);
or OR2 (N12641, N12640, N12234);
or OR3 (N12642, N12638, N11425, N6228);
buf BUF1 (N12643, N12641);
nand NAND2 (N12644, N12642, N8881);
xor XOR2 (N12645, N12636, N8081);
nand NAND2 (N12646, N12644, N11000);
and AND4 (N12647, N12635, N5889, N7826, N7499);
buf BUF1 (N12648, N12646);
xor XOR2 (N12649, N12624, N5275);
not NOT1 (N12650, N12647);
nand NAND4 (N12651, N12648, N234, N6205, N4308);
not NOT1 (N12652, N12643);
buf BUF1 (N12653, N12629);
xor XOR2 (N12654, N12651, N7076);
and AND4 (N12655, N12632, N9848, N8266, N9878);
nor NOR4 (N12656, N12652, N12015, N12030, N5556);
nand NAND3 (N12657, N12654, N2225, N7701);
buf BUF1 (N12658, N12645);
nor NOR3 (N12659, N12639, N6028, N2868);
and AND4 (N12660, N12659, N3931, N8600, N5386);
or OR3 (N12661, N12653, N12068, N993);
buf BUF1 (N12662, N12656);
and AND3 (N12663, N12661, N8706, N866);
nand NAND2 (N12664, N12663, N9105);
xor XOR2 (N12665, N12649, N9331);
or OR3 (N12666, N12665, N10370, N5224);
nor NOR3 (N12667, N12664, N3564, N12516);
nand NAND4 (N12668, N12630, N6149, N3274, N2404);
buf BUF1 (N12669, N12668);
xor XOR2 (N12670, N12666, N3387);
and AND3 (N12671, N12660, N2333, N6575);
nor NOR2 (N12672, N12671, N11461);
and AND4 (N12673, N12662, N5514, N8051, N12320);
nand NAND2 (N12674, N12655, N12245);
xor XOR2 (N12675, N12650, N10829);
or OR2 (N12676, N12674, N4387);
or OR4 (N12677, N12667, N5205, N12206, N11833);
nand NAND3 (N12678, N12633, N12416, N8207);
not NOT1 (N12679, N12677);
not NOT1 (N12680, N12676);
or OR4 (N12681, N12657, N2092, N6999, N3023);
not NOT1 (N12682, N12679);
or OR4 (N12683, N12669, N3080, N10103, N2467);
xor XOR2 (N12684, N12672, N12449);
buf BUF1 (N12685, N12658);
xor XOR2 (N12686, N12681, N4853);
and AND4 (N12687, N12682, N2645, N4755, N7306);
or OR3 (N12688, N12684, N10330, N3545);
nor NOR2 (N12689, N12673, N6593);
not NOT1 (N12690, N12688);
not NOT1 (N12691, N12690);
or OR2 (N12692, N12680, N6858);
nor NOR4 (N12693, N12686, N11391, N10537, N393);
not NOT1 (N12694, N12678);
nor NOR4 (N12695, N12689, N1177, N2847, N9217);
nand NAND4 (N12696, N12693, N8211, N12585, N2699);
buf BUF1 (N12697, N12685);
or OR4 (N12698, N12670, N9127, N12164, N10459);
xor XOR2 (N12699, N12696, N4943);
nand NAND2 (N12700, N12695, N3015);
nand NAND3 (N12701, N12700, N7751, N8638);
not NOT1 (N12702, N12687);
not NOT1 (N12703, N12699);
xor XOR2 (N12704, N12694, N4790);
or OR2 (N12705, N12692, N8129);
or OR4 (N12706, N12702, N2794, N1753, N10808);
buf BUF1 (N12707, N12703);
buf BUF1 (N12708, N12707);
or OR4 (N12709, N12704, N2655, N1074, N5410);
buf BUF1 (N12710, N12697);
or OR2 (N12711, N12683, N10324);
nand NAND2 (N12712, N12705, N5141);
not NOT1 (N12713, N12675);
and AND4 (N12714, N12708, N954, N8046, N787);
nor NOR2 (N12715, N12714, N1957);
nor NOR3 (N12716, N12691, N1799, N12495);
not NOT1 (N12717, N12709);
xor XOR2 (N12718, N12717, N941);
and AND2 (N12719, N12712, N6794);
nand NAND2 (N12720, N12718, N11752);
not NOT1 (N12721, N12715);
nor NOR4 (N12722, N12720, N12344, N12462, N7053);
buf BUF1 (N12723, N12719);
xor XOR2 (N12724, N12701, N11076);
not NOT1 (N12725, N12722);
not NOT1 (N12726, N12710);
xor XOR2 (N12727, N12716, N4313);
nand NAND2 (N12728, N12698, N729);
nor NOR2 (N12729, N12725, N2616);
and AND4 (N12730, N12706, N9809, N9060, N9184);
nand NAND3 (N12731, N12711, N1094, N3877);
buf BUF1 (N12732, N12726);
buf BUF1 (N12733, N12713);
nor NOR2 (N12734, N12730, N8713);
and AND3 (N12735, N12732, N2999, N5595);
nor NOR3 (N12736, N12733, N3355, N5450);
nand NAND3 (N12737, N12727, N11591, N11117);
and AND2 (N12738, N12728, N3064);
xor XOR2 (N12739, N12735, N1773);
nor NOR2 (N12740, N12738, N5409);
not NOT1 (N12741, N12729);
buf BUF1 (N12742, N12723);
nand NAND4 (N12743, N12736, N2364, N5789, N9409);
or OR4 (N12744, N12731, N11289, N2557, N2384);
nor NOR3 (N12745, N12741, N10310, N12661);
or OR2 (N12746, N12734, N7913);
xor XOR2 (N12747, N12724, N12060);
xor XOR2 (N12748, N12742, N1545);
and AND2 (N12749, N12746, N2067);
xor XOR2 (N12750, N12739, N5993);
and AND3 (N12751, N12744, N10494, N7008);
buf BUF1 (N12752, N12749);
or OR4 (N12753, N12747, N11861, N134, N7275);
xor XOR2 (N12754, N12753, N11664);
nor NOR2 (N12755, N12752, N3255);
nand NAND3 (N12756, N12754, N5997, N3869);
nor NOR4 (N12757, N12755, N5567, N3665, N1353);
nor NOR4 (N12758, N12757, N8811, N11227, N6639);
xor XOR2 (N12759, N12737, N9997);
nand NAND3 (N12760, N12745, N194, N2114);
xor XOR2 (N12761, N12740, N8657);
buf BUF1 (N12762, N12743);
not NOT1 (N12763, N12751);
and AND2 (N12764, N12762, N5771);
or OR4 (N12765, N12761, N2227, N7372, N7742);
nand NAND3 (N12766, N12760, N12167, N10635);
nand NAND3 (N12767, N12748, N12183, N1340);
xor XOR2 (N12768, N12756, N9764);
nand NAND2 (N12769, N12763, N12349);
buf BUF1 (N12770, N12750);
nor NOR4 (N12771, N12766, N10567, N11970, N1762);
or OR2 (N12772, N12770, N9302);
or OR2 (N12773, N12772, N11853);
nand NAND4 (N12774, N12764, N4079, N7882, N9880);
or OR3 (N12775, N12758, N9351, N10876);
and AND3 (N12776, N12769, N8003, N1887);
nand NAND4 (N12777, N12773, N1045, N4800, N7131);
nand NAND4 (N12778, N12776, N3802, N401, N393);
nor NOR3 (N12779, N12765, N6334, N2170);
nor NOR3 (N12780, N12779, N2340, N3147);
not NOT1 (N12781, N12774);
not NOT1 (N12782, N12781);
buf BUF1 (N12783, N12780);
xor XOR2 (N12784, N12767, N6662);
or OR3 (N12785, N12721, N3582, N8771);
and AND2 (N12786, N12783, N5557);
and AND2 (N12787, N12785, N11824);
and AND4 (N12788, N12771, N4567, N5943, N6370);
buf BUF1 (N12789, N12775);
buf BUF1 (N12790, N12784);
buf BUF1 (N12791, N12788);
and AND4 (N12792, N12768, N3560, N4625, N6554);
and AND4 (N12793, N12792, N9926, N798, N6816);
and AND4 (N12794, N12778, N5033, N2603, N11288);
nand NAND4 (N12795, N12787, N1587, N9926, N1515);
and AND3 (N12796, N12759, N11008, N5404);
not NOT1 (N12797, N12795);
nand NAND2 (N12798, N12777, N11543);
xor XOR2 (N12799, N12797, N1191);
nand NAND3 (N12800, N12796, N1126, N8374);
nor NOR3 (N12801, N12786, N9044, N12155);
nand NAND3 (N12802, N12782, N3393, N1027);
not NOT1 (N12803, N12790);
not NOT1 (N12804, N12800);
not NOT1 (N12805, N12802);
nand NAND4 (N12806, N12793, N1511, N3109, N10864);
xor XOR2 (N12807, N12804, N1740);
or OR3 (N12808, N12799, N5913, N12019);
and AND4 (N12809, N12794, N7470, N9988, N2242);
nand NAND4 (N12810, N12801, N7807, N12565, N5392);
or OR4 (N12811, N12809, N3918, N4743, N4170);
and AND3 (N12812, N12805, N7195, N5629);
or OR2 (N12813, N12810, N3739);
or OR3 (N12814, N12803, N8899, N608);
buf BUF1 (N12815, N12798);
not NOT1 (N12816, N12806);
nor NOR4 (N12817, N12789, N7031, N2270, N9907);
not NOT1 (N12818, N12816);
nand NAND3 (N12819, N12813, N3893, N7468);
nand NAND3 (N12820, N12819, N10856, N4024);
nand NAND2 (N12821, N12791, N4491);
not NOT1 (N12822, N12818);
buf BUF1 (N12823, N12807);
buf BUF1 (N12824, N12808);
buf BUF1 (N12825, N12814);
buf BUF1 (N12826, N12823);
buf BUF1 (N12827, N12812);
not NOT1 (N12828, N12811);
buf BUF1 (N12829, N12817);
or OR3 (N12830, N12825, N10794, N3863);
nor NOR3 (N12831, N12826, N1129, N3034);
xor XOR2 (N12832, N12831, N6567);
nand NAND3 (N12833, N12821, N8144, N397);
and AND2 (N12834, N12822, N7599);
not NOT1 (N12835, N12834);
buf BUF1 (N12836, N12815);
and AND3 (N12837, N12824, N3994, N3295);
and AND3 (N12838, N12832, N2103, N729);
nor NOR3 (N12839, N12836, N4205, N10445);
nand NAND4 (N12840, N12828, N6087, N863, N9062);
not NOT1 (N12841, N12827);
and AND3 (N12842, N12820, N7909, N1336);
or OR3 (N12843, N12833, N12656, N7184);
nor NOR3 (N12844, N12835, N6930, N2482);
and AND3 (N12845, N12839, N12708, N12026);
xor XOR2 (N12846, N12837, N12669);
xor XOR2 (N12847, N12846, N3555);
nand NAND3 (N12848, N12847, N111, N9943);
xor XOR2 (N12849, N12848, N2923);
and AND4 (N12850, N12845, N4077, N3442, N395);
and AND4 (N12851, N12849, N410, N6766, N9982);
and AND3 (N12852, N12841, N7322, N2290);
nor NOR3 (N12853, N12843, N8068, N1877);
buf BUF1 (N12854, N12830);
nand NAND2 (N12855, N12844, N12000);
or OR2 (N12856, N12842, N5441);
not NOT1 (N12857, N12840);
nand NAND3 (N12858, N12829, N12517, N6182);
and AND4 (N12859, N12857, N2970, N8656, N1117);
and AND2 (N12860, N12838, N8849);
and AND3 (N12861, N12855, N300, N1008);
xor XOR2 (N12862, N12856, N4750);
and AND2 (N12863, N12861, N6777);
nor NOR3 (N12864, N12851, N6829, N9640);
and AND2 (N12865, N12858, N4679);
xor XOR2 (N12866, N12864, N11996);
not NOT1 (N12867, N12850);
xor XOR2 (N12868, N12862, N7781);
or OR4 (N12869, N12860, N8632, N6832, N7662);
not NOT1 (N12870, N12868);
nor NOR3 (N12871, N12866, N10524, N7004);
and AND4 (N12872, N12870, N5948, N7203, N10790);
or OR2 (N12873, N12869, N6192);
and AND4 (N12874, N12867, N4870, N6741, N12859);
xor XOR2 (N12875, N12402, N6290);
and AND3 (N12876, N12853, N7940, N10759);
xor XOR2 (N12877, N12865, N1687);
buf BUF1 (N12878, N12854);
not NOT1 (N12879, N12871);
xor XOR2 (N12880, N12852, N3829);
or OR3 (N12881, N12872, N3821, N3895);
xor XOR2 (N12882, N12879, N9892);
nor NOR3 (N12883, N12881, N9990, N5040);
nor NOR2 (N12884, N12880, N7892);
buf BUF1 (N12885, N12878);
nor NOR3 (N12886, N12863, N477, N5908);
nor NOR4 (N12887, N12876, N10899, N4975, N4026);
buf BUF1 (N12888, N12882);
not NOT1 (N12889, N12875);
nor NOR2 (N12890, N12888, N11588);
xor XOR2 (N12891, N12873, N9694);
or OR4 (N12892, N12887, N8115, N11764, N738);
not NOT1 (N12893, N12883);
nor NOR3 (N12894, N12874, N10241, N612);
not NOT1 (N12895, N12890);
buf BUF1 (N12896, N12885);
nor NOR3 (N12897, N12896, N9637, N5834);
xor XOR2 (N12898, N12894, N6346);
or OR3 (N12899, N12884, N11770, N12561);
and AND3 (N12900, N12897, N12052, N7991);
nand NAND2 (N12901, N12895, N12295);
not NOT1 (N12902, N12886);
and AND4 (N12903, N12877, N2290, N1216, N2561);
buf BUF1 (N12904, N12893);
buf BUF1 (N12905, N12899);
nor NOR2 (N12906, N12889, N5271);
not NOT1 (N12907, N12906);
nand NAND4 (N12908, N12898, N11010, N7267, N9002);
and AND3 (N12909, N12892, N434, N9890);
xor XOR2 (N12910, N12908, N10110);
buf BUF1 (N12911, N12907);
nand NAND3 (N12912, N12909, N4684, N7296);
buf BUF1 (N12913, N12904);
buf BUF1 (N12914, N12903);
not NOT1 (N12915, N12905);
or OR3 (N12916, N12911, N1921, N10005);
or OR4 (N12917, N12914, N3, N1358, N5651);
not NOT1 (N12918, N12917);
not NOT1 (N12919, N12891);
xor XOR2 (N12920, N12902, N10126);
nand NAND3 (N12921, N12901, N10201, N7221);
nand NAND4 (N12922, N12910, N6958, N8173, N4413);
buf BUF1 (N12923, N12913);
nand NAND3 (N12924, N12915, N2287, N9646);
or OR3 (N12925, N12921, N5735, N9623);
nand NAND3 (N12926, N12920, N4787, N9296);
xor XOR2 (N12927, N12919, N10887);
buf BUF1 (N12928, N12916);
and AND2 (N12929, N12927, N9902);
and AND2 (N12930, N12929, N10189);
and AND3 (N12931, N12925, N11298, N445);
nor NOR4 (N12932, N12900, N1374, N3432, N11517);
or OR3 (N12933, N12931, N6375, N12359);
not NOT1 (N12934, N12924);
or OR2 (N12935, N12912, N6206);
and AND4 (N12936, N12935, N7317, N10431, N12223);
and AND3 (N12937, N12930, N5848, N519);
nor NOR4 (N12938, N12933, N12418, N5839, N391);
nor NOR2 (N12939, N12926, N12474);
and AND2 (N12940, N12938, N1925);
nand NAND3 (N12941, N12940, N8497, N1784);
or OR3 (N12942, N12941, N6263, N320);
nand NAND4 (N12943, N12923, N2666, N4253, N1492);
and AND2 (N12944, N12928, N7137);
xor XOR2 (N12945, N12943, N10983);
or OR2 (N12946, N12944, N6965);
and AND3 (N12947, N12922, N5483, N4157);
nand NAND3 (N12948, N12934, N11689, N11193);
xor XOR2 (N12949, N12937, N7997);
not NOT1 (N12950, N12947);
xor XOR2 (N12951, N12950, N8113);
nor NOR3 (N12952, N12949, N10405, N8517);
nor NOR3 (N12953, N12918, N3595, N2274);
xor XOR2 (N12954, N12939, N4354);
or OR2 (N12955, N12942, N10815);
and AND3 (N12956, N12953, N12758, N2943);
buf BUF1 (N12957, N12951);
nor NOR2 (N12958, N12955, N7305);
and AND2 (N12959, N12952, N12342);
and AND2 (N12960, N12958, N1840);
xor XOR2 (N12961, N12960, N2675);
nand NAND2 (N12962, N12936, N8610);
xor XOR2 (N12963, N12961, N5352);
not NOT1 (N12964, N12962);
not NOT1 (N12965, N12954);
nand NAND3 (N12966, N12948, N268, N7423);
nand NAND2 (N12967, N12957, N2295);
or OR2 (N12968, N12946, N8296);
buf BUF1 (N12969, N12968);
and AND2 (N12970, N12966, N9182);
not NOT1 (N12971, N12965);
not NOT1 (N12972, N12945);
or OR3 (N12973, N12959, N12255, N1119);
buf BUF1 (N12974, N12967);
and AND2 (N12975, N12974, N3440);
xor XOR2 (N12976, N12973, N4683);
not NOT1 (N12977, N12932);
nand NAND4 (N12978, N12975, N11139, N6802, N5161);
or OR4 (N12979, N12963, N1530, N3925, N3222);
buf BUF1 (N12980, N12976);
nor NOR3 (N12981, N12956, N12269, N4119);
nor NOR3 (N12982, N12969, N3333, N9209);
buf BUF1 (N12983, N12972);
xor XOR2 (N12984, N12983, N1964);
or OR3 (N12985, N12977, N2307, N3614);
or OR2 (N12986, N12970, N9315);
not NOT1 (N12987, N12980);
nand NAND3 (N12988, N12971, N7951, N994);
nor NOR4 (N12989, N12985, N1798, N1175, N798);
and AND4 (N12990, N12978, N5115, N528, N9886);
or OR2 (N12991, N12989, N9043);
not NOT1 (N12992, N12987);
nand NAND3 (N12993, N12981, N8656, N11858);
nand NAND4 (N12994, N12964, N7942, N658, N9577);
nand NAND4 (N12995, N12982, N2353, N3041, N10505);
not NOT1 (N12996, N12991);
nand NAND2 (N12997, N12995, N4650);
buf BUF1 (N12998, N12996);
buf BUF1 (N12999, N12986);
not NOT1 (N13000, N12999);
xor XOR2 (N13001, N12993, N10316);
buf BUF1 (N13002, N12988);
and AND3 (N13003, N12997, N12157, N10213);
buf BUF1 (N13004, N13002);
nand NAND2 (N13005, N13003, N8695);
or OR4 (N13006, N12998, N11304, N10054, N10221);
buf BUF1 (N13007, N13001);
buf BUF1 (N13008, N12994);
not NOT1 (N13009, N13000);
not NOT1 (N13010, N12992);
nor NOR4 (N13011, N13010, N7068, N2323, N1366);
xor XOR2 (N13012, N13008, N11117);
and AND2 (N13013, N13009, N1536);
not NOT1 (N13014, N13007);
or OR2 (N13015, N12990, N10150);
and AND2 (N13016, N13004, N9674);
buf BUF1 (N13017, N13016);
not NOT1 (N13018, N12984);
buf BUF1 (N13019, N13005);
and AND4 (N13020, N13015, N11714, N10398, N5067);
not NOT1 (N13021, N13014);
xor XOR2 (N13022, N13021, N7927);
buf BUF1 (N13023, N13020);
buf BUF1 (N13024, N13018);
and AND2 (N13025, N13022, N3934);
nor NOR2 (N13026, N13023, N6340);
xor XOR2 (N13027, N13026, N11432);
nor NOR2 (N13028, N13011, N8857);
and AND3 (N13029, N13017, N11628, N1125);
nor NOR3 (N13030, N13024, N8448, N3675);
nand NAND3 (N13031, N13012, N1738, N7168);
nor NOR4 (N13032, N13019, N566, N5089, N5531);
not NOT1 (N13033, N12979);
xor XOR2 (N13034, N13032, N10462);
xor XOR2 (N13035, N13013, N2930);
and AND3 (N13036, N13031, N6396, N1762);
buf BUF1 (N13037, N13034);
buf BUF1 (N13038, N13027);
or OR3 (N13039, N13037, N11941, N134);
nand NAND4 (N13040, N13030, N5938, N2934, N6020);
buf BUF1 (N13041, N13006);
xor XOR2 (N13042, N13028, N1479);
xor XOR2 (N13043, N13025, N9213);
nor NOR3 (N13044, N13043, N8377, N5082);
and AND3 (N13045, N13035, N2524, N4891);
not NOT1 (N13046, N13041);
buf BUF1 (N13047, N13038);
buf BUF1 (N13048, N13029);
not NOT1 (N13049, N13048);
xor XOR2 (N13050, N13040, N1445);
nor NOR4 (N13051, N13044, N10391, N1515, N1733);
nor NOR4 (N13052, N13042, N442, N853, N4058);
buf BUF1 (N13053, N13047);
buf BUF1 (N13054, N13052);
nor NOR4 (N13055, N13054, N8897, N6892, N10653);
and AND4 (N13056, N13046, N8841, N1040, N6463);
not NOT1 (N13057, N13051);
buf BUF1 (N13058, N13053);
buf BUF1 (N13059, N13049);
buf BUF1 (N13060, N13036);
xor XOR2 (N13061, N13060, N8396);
and AND3 (N13062, N13033, N2432, N8715);
buf BUF1 (N13063, N13056);
xor XOR2 (N13064, N13039, N10635);
or OR3 (N13065, N13055, N4843, N11173);
nor NOR4 (N13066, N13063, N10964, N7267, N6667);
and AND2 (N13067, N13057, N1607);
nand NAND2 (N13068, N13050, N8306);
buf BUF1 (N13069, N13067);
nor NOR3 (N13070, N13058, N9413, N7506);
xor XOR2 (N13071, N13045, N8583);
nor NOR2 (N13072, N13059, N10146);
nand NAND4 (N13073, N13064, N499, N993, N1202);
and AND4 (N13074, N13068, N3967, N6624, N207);
or OR3 (N13075, N13065, N8363, N1424);
xor XOR2 (N13076, N13062, N7264);
nor NOR3 (N13077, N13066, N4504, N1551);
nand NAND2 (N13078, N13061, N885);
and AND4 (N13079, N13070, N12324, N6240, N4023);
nor NOR4 (N13080, N13069, N10583, N10766, N394);
buf BUF1 (N13081, N13078);
nor NOR2 (N13082, N13075, N1665);
xor XOR2 (N13083, N13081, N8947);
xor XOR2 (N13084, N13079, N301);
buf BUF1 (N13085, N13084);
nand NAND3 (N13086, N13077, N12432, N2233);
nand NAND2 (N13087, N13073, N4397);
or OR3 (N13088, N13072, N4591, N1589);
and AND2 (N13089, N13082, N4462);
or OR3 (N13090, N13086, N130, N2381);
buf BUF1 (N13091, N13074);
and AND3 (N13092, N13089, N1832, N10057);
nand NAND2 (N13093, N13080, N1651);
and AND2 (N13094, N13090, N7477);
nor NOR4 (N13095, N13091, N1016, N368, N8262);
nor NOR4 (N13096, N13095, N9941, N11108, N5373);
not NOT1 (N13097, N13096);
or OR3 (N13098, N13087, N6923, N2573);
or OR2 (N13099, N13097, N4471);
nand NAND4 (N13100, N13083, N8633, N2303, N6916);
buf BUF1 (N13101, N13085);
and AND4 (N13102, N13071, N7315, N8249, N6952);
not NOT1 (N13103, N13102);
buf BUF1 (N13104, N13088);
nand NAND4 (N13105, N13099, N3887, N9432, N133);
xor XOR2 (N13106, N13103, N12017);
or OR4 (N13107, N13105, N10616, N9842, N10365);
or OR3 (N13108, N13076, N4325, N3993);
nand NAND4 (N13109, N13107, N4983, N10579, N5262);
or OR2 (N13110, N13109, N13044);
buf BUF1 (N13111, N13098);
or OR4 (N13112, N13104, N1346, N3796, N7126);
nand NAND3 (N13113, N13100, N1978, N8732);
nor NOR2 (N13114, N13112, N2403);
not NOT1 (N13115, N13101);
nand NAND3 (N13116, N13115, N9366, N6653);
and AND3 (N13117, N13092, N940, N10245);
xor XOR2 (N13118, N13094, N7456);
buf BUF1 (N13119, N13111);
nand NAND3 (N13120, N13106, N4032, N9711);
buf BUF1 (N13121, N13117);
or OR4 (N13122, N13120, N9501, N1088, N6673);
buf BUF1 (N13123, N13121);
or OR2 (N13124, N13113, N6821);
xor XOR2 (N13125, N13123, N6132);
not NOT1 (N13126, N13124);
or OR2 (N13127, N13110, N3020);
or OR2 (N13128, N13108, N10079);
and AND2 (N13129, N13114, N9790);
and AND4 (N13130, N13118, N11226, N9818, N8734);
xor XOR2 (N13131, N13119, N5100);
xor XOR2 (N13132, N13126, N4404);
and AND2 (N13133, N13093, N9577);
nand NAND4 (N13134, N13116, N3553, N6276, N11006);
nand NAND2 (N13135, N13133, N182);
buf BUF1 (N13136, N13128);
xor XOR2 (N13137, N13134, N2246);
or OR4 (N13138, N13137, N6406, N4688, N5638);
nor NOR4 (N13139, N13136, N9548, N7856, N12302);
not NOT1 (N13140, N13127);
nor NOR4 (N13141, N13130, N8657, N8548, N8481);
buf BUF1 (N13142, N13122);
nor NOR2 (N13143, N13129, N11837);
nand NAND4 (N13144, N13125, N5807, N8267, N11527);
nor NOR4 (N13145, N13131, N8757, N2487, N9834);
or OR4 (N13146, N13138, N1682, N5663, N2396);
or OR4 (N13147, N13132, N3243, N13063, N1915);
buf BUF1 (N13148, N13146);
nand NAND4 (N13149, N13135, N5919, N10317, N6904);
and AND2 (N13150, N13143, N2589);
nor NOR2 (N13151, N13141, N9574);
buf BUF1 (N13152, N13145);
not NOT1 (N13153, N13150);
not NOT1 (N13154, N13147);
xor XOR2 (N13155, N13149, N11152);
not NOT1 (N13156, N13155);
and AND2 (N13157, N13156, N574);
not NOT1 (N13158, N13140);
nand NAND4 (N13159, N13153, N304, N2542, N12622);
or OR2 (N13160, N13144, N12463);
or OR2 (N13161, N13139, N13032);
nor NOR2 (N13162, N13151, N6748);
or OR4 (N13163, N13157, N9494, N11792, N1359);
buf BUF1 (N13164, N13162);
xor XOR2 (N13165, N13161, N747);
and AND4 (N13166, N13160, N3591, N9838, N1349);
not NOT1 (N13167, N13164);
xor XOR2 (N13168, N13163, N11114);
and AND4 (N13169, N13148, N12529, N9705, N1269);
and AND4 (N13170, N13169, N9651, N3548, N11267);
buf BUF1 (N13171, N13152);
and AND2 (N13172, N13170, N4992);
nand NAND3 (N13173, N13154, N6315, N8397);
buf BUF1 (N13174, N13168);
nand NAND4 (N13175, N13159, N7341, N4737, N8334);
or OR3 (N13176, N13172, N11968, N10902);
nand NAND4 (N13177, N13174, N486, N3181, N5625);
buf BUF1 (N13178, N13177);
buf BUF1 (N13179, N13166);
or OR3 (N13180, N13167, N9690, N10408);
and AND4 (N13181, N13175, N624, N9965, N3783);
or OR4 (N13182, N13171, N4201, N2750, N12953);
buf BUF1 (N13183, N13179);
or OR2 (N13184, N13173, N9814);
buf BUF1 (N13185, N13176);
or OR2 (N13186, N13183, N10682);
nand NAND4 (N13187, N13182, N1943, N1709, N3455);
buf BUF1 (N13188, N13185);
and AND2 (N13189, N13180, N3191);
not NOT1 (N13190, N13181);
and AND3 (N13191, N13158, N11155, N10);
xor XOR2 (N13192, N13178, N211);
and AND3 (N13193, N13187, N4588, N704);
and AND3 (N13194, N13165, N1965, N10616);
nand NAND4 (N13195, N13190, N3890, N7223, N4367);
and AND2 (N13196, N13142, N2013);
nand NAND3 (N13197, N13188, N3922, N11532);
and AND2 (N13198, N13192, N11883);
xor XOR2 (N13199, N13186, N1247);
or OR3 (N13200, N13196, N3184, N1540);
nand NAND2 (N13201, N13191, N11283);
xor XOR2 (N13202, N13189, N12090);
buf BUF1 (N13203, N13195);
xor XOR2 (N13204, N13193, N9476);
nand NAND3 (N13205, N13200, N12435, N714);
nand NAND3 (N13206, N13203, N8978, N10074);
nor NOR2 (N13207, N13202, N7052);
or OR4 (N13208, N13197, N1642, N8803, N742);
or OR2 (N13209, N13198, N3612);
nand NAND4 (N13210, N13184, N1368, N11826, N7127);
and AND4 (N13211, N13210, N12070, N12386, N11651);
buf BUF1 (N13212, N13211);
nand NAND3 (N13213, N13206, N11279, N7336);
nand NAND2 (N13214, N13204, N8086);
or OR3 (N13215, N13208, N2443, N6458);
not NOT1 (N13216, N13209);
nand NAND3 (N13217, N13215, N12506, N9128);
xor XOR2 (N13218, N13199, N4777);
nor NOR2 (N13219, N13207, N6356);
and AND3 (N13220, N13214, N6611, N11004);
nand NAND4 (N13221, N13219, N13145, N6176, N5813);
nor NOR2 (N13222, N13217, N8736);
xor XOR2 (N13223, N13218, N353);
and AND2 (N13224, N13221, N10088);
not NOT1 (N13225, N13222);
and AND3 (N13226, N13224, N4976, N1949);
nand NAND3 (N13227, N13213, N1872, N13124);
nand NAND2 (N13228, N13212, N8700);
buf BUF1 (N13229, N13226);
and AND4 (N13230, N13201, N3804, N166, N8417);
and AND4 (N13231, N13230, N10504, N4709, N3124);
or OR4 (N13232, N13229, N9428, N302, N10213);
nand NAND4 (N13233, N13194, N10742, N7109, N6174);
or OR3 (N13234, N13228, N9373, N6352);
xor XOR2 (N13235, N13233, N1323);
nor NOR4 (N13236, N13216, N1320, N3933, N10486);
nand NAND2 (N13237, N13205, N12176);
and AND4 (N13238, N13236, N11100, N7667, N9902);
and AND2 (N13239, N13220, N761);
xor XOR2 (N13240, N13231, N7071);
or OR3 (N13241, N13238, N12113, N8059);
or OR4 (N13242, N13223, N7351, N8764, N3927);
and AND2 (N13243, N13242, N11199);
nand NAND4 (N13244, N13225, N9541, N8648, N3068);
nor NOR4 (N13245, N13234, N7733, N8922, N9834);
xor XOR2 (N13246, N13227, N12306);
buf BUF1 (N13247, N13246);
not NOT1 (N13248, N13237);
not NOT1 (N13249, N13247);
not NOT1 (N13250, N13249);
and AND2 (N13251, N13245, N8409);
or OR3 (N13252, N13235, N4112, N5468);
nor NOR3 (N13253, N13241, N2654, N2394);
not NOT1 (N13254, N13243);
and AND4 (N13255, N13251, N5972, N12622, N8347);
buf BUF1 (N13256, N13253);
xor XOR2 (N13257, N13252, N508);
nor NOR2 (N13258, N13248, N11484);
nor NOR4 (N13259, N13256, N9530, N7551, N1386);
nor NOR3 (N13260, N13240, N5660, N697);
buf BUF1 (N13261, N13255);
or OR2 (N13262, N13239, N4736);
not NOT1 (N13263, N13250);
nand NAND4 (N13264, N13261, N5960, N2396, N4879);
nand NAND3 (N13265, N13259, N11152, N862);
buf BUF1 (N13266, N13258);
or OR2 (N13267, N13232, N11340);
nor NOR4 (N13268, N13265, N1911, N10994, N6008);
or OR4 (N13269, N13262, N8703, N10275, N5623);
or OR3 (N13270, N13254, N5470, N1977);
or OR4 (N13271, N13266, N823, N5491, N12524);
nor NOR4 (N13272, N13263, N11328, N7896, N2870);
nand NAND4 (N13273, N13244, N7479, N5509, N4354);
and AND4 (N13274, N13272, N5334, N449, N6540);
nand NAND3 (N13275, N13264, N12454, N6995);
nand NAND4 (N13276, N13260, N7296, N210, N5887);
nand NAND2 (N13277, N13276, N10144);
and AND3 (N13278, N13267, N4383, N8608);
nor NOR4 (N13279, N13277, N6557, N10513, N6682);
buf BUF1 (N13280, N13273);
xor XOR2 (N13281, N13280, N874);
nand NAND2 (N13282, N13270, N7239);
xor XOR2 (N13283, N13281, N4101);
or OR4 (N13284, N13275, N2920, N12932, N124);
and AND3 (N13285, N13268, N11891, N5441);
and AND3 (N13286, N13284, N1149, N8344);
and AND2 (N13287, N13283, N11327);
not NOT1 (N13288, N13282);
or OR2 (N13289, N13287, N7877);
not NOT1 (N13290, N13289);
xor XOR2 (N13291, N13257, N178);
nand NAND2 (N13292, N13291, N11987);
buf BUF1 (N13293, N13288);
not NOT1 (N13294, N13274);
or OR4 (N13295, N13279, N5803, N3212, N6993);
and AND2 (N13296, N13295, N4272);
and AND3 (N13297, N13269, N12625, N5412);
and AND2 (N13298, N13297, N9649);
or OR3 (N13299, N13293, N8219, N5427);
nand NAND2 (N13300, N13299, N1473);
or OR3 (N13301, N13271, N10834, N6974);
buf BUF1 (N13302, N13300);
nand NAND2 (N13303, N13298, N7383);
or OR4 (N13304, N13292, N4036, N3783, N895);
xor XOR2 (N13305, N13303, N965);
and AND2 (N13306, N13285, N12009);
or OR4 (N13307, N13302, N10295, N3445, N7276);
xor XOR2 (N13308, N13307, N7937);
and AND3 (N13309, N13294, N6534, N11407);
and AND3 (N13310, N13306, N10026, N7316);
xor XOR2 (N13311, N13296, N11897);
xor XOR2 (N13312, N13278, N4824);
nand NAND3 (N13313, N13309, N6793, N3879);
xor XOR2 (N13314, N13310, N2808);
xor XOR2 (N13315, N13305, N11030);
or OR4 (N13316, N13290, N9521, N5898, N8381);
nor NOR4 (N13317, N13313, N7528, N6767, N9683);
buf BUF1 (N13318, N13311);
nor NOR2 (N13319, N13317, N5253);
xor XOR2 (N13320, N13308, N5405);
xor XOR2 (N13321, N13301, N3660);
nor NOR4 (N13322, N13286, N9191, N12438, N12494);
xor XOR2 (N13323, N13304, N11496);
or OR3 (N13324, N13322, N11117, N1947);
or OR2 (N13325, N13323, N2214);
or OR4 (N13326, N13316, N3498, N9941, N7948);
and AND2 (N13327, N13318, N4732);
not NOT1 (N13328, N13314);
and AND3 (N13329, N13321, N4184, N11335);
nor NOR3 (N13330, N13325, N3638, N2266);
buf BUF1 (N13331, N13319);
or OR4 (N13332, N13330, N6119, N1425, N2846);
or OR4 (N13333, N13328, N10706, N8484, N12774);
xor XOR2 (N13334, N13326, N3914);
xor XOR2 (N13335, N13320, N12121);
nor NOR2 (N13336, N13329, N8335);
and AND2 (N13337, N13327, N12326);
not NOT1 (N13338, N13337);
nand NAND3 (N13339, N13315, N5902, N135);
not NOT1 (N13340, N13339);
buf BUF1 (N13341, N13335);
buf BUF1 (N13342, N13312);
not NOT1 (N13343, N13332);
and AND4 (N13344, N13333, N4875, N11936, N6789);
or OR2 (N13345, N13343, N4574);
nand NAND3 (N13346, N13334, N11755, N4489);
buf BUF1 (N13347, N13331);
buf BUF1 (N13348, N13324);
or OR3 (N13349, N13341, N9163, N10133);
xor XOR2 (N13350, N13336, N7745);
buf BUF1 (N13351, N13349);
not NOT1 (N13352, N13338);
xor XOR2 (N13353, N13346, N7060);
or OR4 (N13354, N13342, N2359, N9737, N13142);
buf BUF1 (N13355, N13340);
nor NOR3 (N13356, N13347, N7161, N3237);
or OR3 (N13357, N13356, N9290, N7208);
xor XOR2 (N13358, N13352, N2198);
buf BUF1 (N13359, N13348);
nand NAND2 (N13360, N13353, N12580);
buf BUF1 (N13361, N13354);
nand NAND4 (N13362, N13344, N10733, N11986, N3167);
or OR2 (N13363, N13350, N5729);
nand NAND4 (N13364, N13355, N5560, N6552, N3199);
not NOT1 (N13365, N13357);
and AND4 (N13366, N13363, N3935, N3544, N9627);
nand NAND4 (N13367, N13351, N1643, N12550, N1209);
buf BUF1 (N13368, N13359);
nor NOR3 (N13369, N13360, N11129, N5016);
and AND3 (N13370, N13358, N11670, N10217);
not NOT1 (N13371, N13368);
xor XOR2 (N13372, N13366, N3172);
xor XOR2 (N13373, N13364, N5451);
buf BUF1 (N13374, N13369);
and AND2 (N13375, N13367, N7734);
not NOT1 (N13376, N13361);
or OR3 (N13377, N13371, N2843, N3365);
or OR3 (N13378, N13365, N3793, N248);
xor XOR2 (N13379, N13362, N4765);
or OR2 (N13380, N13374, N1598);
buf BUF1 (N13381, N13376);
xor XOR2 (N13382, N13345, N13082);
not NOT1 (N13383, N13377);
buf BUF1 (N13384, N13382);
or OR2 (N13385, N13375, N9265);
nor NOR3 (N13386, N13370, N683, N3975);
not NOT1 (N13387, N13381);
nor NOR3 (N13388, N13386, N8217, N5322);
buf BUF1 (N13389, N13373);
nand NAND2 (N13390, N13385, N4310);
and AND4 (N13391, N13390, N8300, N9840, N2116);
nor NOR4 (N13392, N13384, N2777, N2656, N7844);
or OR3 (N13393, N13380, N3730, N2992);
or OR3 (N13394, N13372, N9894, N8858);
not NOT1 (N13395, N13379);
xor XOR2 (N13396, N13383, N3856);
nor NOR4 (N13397, N13393, N6651, N8984, N6538);
or OR3 (N13398, N13397, N9233, N429);
or OR3 (N13399, N13398, N12637, N7672);
and AND2 (N13400, N13388, N6159);
nor NOR3 (N13401, N13396, N9701, N445);
not NOT1 (N13402, N13401);
buf BUF1 (N13403, N13399);
and AND3 (N13404, N13392, N9982, N7901);
not NOT1 (N13405, N13395);
nand NAND4 (N13406, N13404, N5696, N523, N11623);
not NOT1 (N13407, N13394);
nand NAND2 (N13408, N13391, N8253);
xor XOR2 (N13409, N13402, N606);
and AND2 (N13410, N13407, N6535);
not NOT1 (N13411, N13400);
and AND4 (N13412, N13387, N5409, N2055, N11235);
nand NAND2 (N13413, N13409, N9017);
buf BUF1 (N13414, N13412);
xor XOR2 (N13415, N13411, N2416);
and AND2 (N13416, N13408, N7990);
not NOT1 (N13417, N13403);
not NOT1 (N13418, N13413);
or OR4 (N13419, N13415, N4647, N3355, N12267);
nand NAND4 (N13420, N13419, N1010, N4500, N813);
xor XOR2 (N13421, N13420, N713);
buf BUF1 (N13422, N13414);
not NOT1 (N13423, N13418);
nor NOR3 (N13424, N13405, N11978, N2956);
and AND3 (N13425, N13417, N13354, N10974);
not NOT1 (N13426, N13425);
or OR3 (N13427, N13416, N762, N11111);
and AND3 (N13428, N13422, N4043, N9626);
and AND2 (N13429, N13410, N11222);
buf BUF1 (N13430, N13427);
and AND2 (N13431, N13423, N9701);
nand NAND2 (N13432, N13429, N7905);
not NOT1 (N13433, N13428);
nand NAND2 (N13434, N13424, N7564);
and AND2 (N13435, N13431, N7435);
nand NAND2 (N13436, N13421, N10050);
nand NAND4 (N13437, N13432, N8998, N3898, N7867);
buf BUF1 (N13438, N13378);
and AND4 (N13439, N13434, N12453, N1892, N2597);
and AND4 (N13440, N13406, N1560, N897, N9722);
not NOT1 (N13441, N13433);
nand NAND2 (N13442, N13435, N11198);
and AND4 (N13443, N13439, N4773, N13032, N10074);
xor XOR2 (N13444, N13430, N4999);
not NOT1 (N13445, N13426);
nor NOR3 (N13446, N13438, N9155, N6165);
xor XOR2 (N13447, N13444, N33);
or OR4 (N13448, N13443, N6190, N421, N399);
not NOT1 (N13449, N13437);
and AND2 (N13450, N13436, N8910);
xor XOR2 (N13451, N13389, N10127);
nor NOR2 (N13452, N13447, N12711);
or OR4 (N13453, N13440, N7957, N54, N2064);
or OR3 (N13454, N13448, N9822, N2012);
buf BUF1 (N13455, N13452);
and AND2 (N13456, N13445, N6438);
xor XOR2 (N13457, N13442, N10809);
buf BUF1 (N13458, N13451);
nand NAND4 (N13459, N13450, N11104, N3464, N3867);
and AND3 (N13460, N13453, N3120, N10705);
and AND2 (N13461, N13458, N11997);
or OR2 (N13462, N13457, N2582);
buf BUF1 (N13463, N13449);
buf BUF1 (N13464, N13461);
not NOT1 (N13465, N13463);
or OR4 (N13466, N13462, N4650, N12491, N10209);
and AND3 (N13467, N13456, N166, N5610);
xor XOR2 (N13468, N13465, N1591);
or OR2 (N13469, N13467, N2325);
buf BUF1 (N13470, N13454);
and AND4 (N13471, N13460, N6288, N13395, N124);
buf BUF1 (N13472, N13455);
not NOT1 (N13473, N13446);
or OR4 (N13474, N13470, N12396, N10589, N12332);
xor XOR2 (N13475, N13464, N4191);
not NOT1 (N13476, N13471);
xor XOR2 (N13477, N13476, N12783);
nor NOR2 (N13478, N13441, N12097);
or OR4 (N13479, N13477, N11289, N12663, N1766);
xor XOR2 (N13480, N13472, N5366);
xor XOR2 (N13481, N13480, N12781);
nor NOR2 (N13482, N13459, N2617);
or OR3 (N13483, N13475, N11765, N11098);
buf BUF1 (N13484, N13468);
not NOT1 (N13485, N13469);
and AND2 (N13486, N13474, N5676);
not NOT1 (N13487, N13479);
nand NAND4 (N13488, N13466, N10120, N1023, N1247);
or OR2 (N13489, N13478, N4369);
nor NOR4 (N13490, N13473, N2933, N3225, N10324);
nor NOR3 (N13491, N13481, N3346, N7549);
nor NOR3 (N13492, N13488, N10555, N12996);
nand NAND4 (N13493, N13482, N5861, N3716, N8094);
nand NAND2 (N13494, N13490, N4282);
buf BUF1 (N13495, N13493);
xor XOR2 (N13496, N13495, N6672);
xor XOR2 (N13497, N13489, N2254);
nand NAND3 (N13498, N13492, N338, N8490);
xor XOR2 (N13499, N13483, N9682);
not NOT1 (N13500, N13491);
nand NAND3 (N13501, N13498, N7328, N5642);
and AND4 (N13502, N13494, N1159, N7663, N9036);
xor XOR2 (N13503, N13485, N6123);
and AND4 (N13504, N13501, N13137, N7813, N11361);
nand NAND2 (N13505, N13500, N8290);
xor XOR2 (N13506, N13499, N12206);
and AND2 (N13507, N13497, N3487);
nand NAND4 (N13508, N13487, N9896, N3501, N7807);
and AND2 (N13509, N13496, N3924);
nand NAND2 (N13510, N13506, N13044);
xor XOR2 (N13511, N13486, N7816);
nor NOR4 (N13512, N13508, N12071, N7682, N4064);
xor XOR2 (N13513, N13504, N6833);
or OR3 (N13514, N13511, N2776, N859);
nand NAND2 (N13515, N13510, N11396);
buf BUF1 (N13516, N13509);
or OR2 (N13517, N13484, N1962);
xor XOR2 (N13518, N13507, N3182);
nand NAND3 (N13519, N13505, N878, N4178);
not NOT1 (N13520, N13519);
and AND3 (N13521, N13512, N9358, N4097);
xor XOR2 (N13522, N13521, N11880);
xor XOR2 (N13523, N13517, N5991);
nand NAND4 (N13524, N13503, N574, N10089, N2986);
not NOT1 (N13525, N13514);
or OR4 (N13526, N13520, N8916, N8534, N3414);
buf BUF1 (N13527, N13513);
nor NOR2 (N13528, N13516, N12929);
xor XOR2 (N13529, N13518, N4801);
buf BUF1 (N13530, N13525);
and AND2 (N13531, N13522, N1978);
nor NOR4 (N13532, N13527, N6887, N1303, N8522);
buf BUF1 (N13533, N13526);
nand NAND3 (N13534, N13524, N4883, N9467);
not NOT1 (N13535, N13531);
not NOT1 (N13536, N13532);
nor NOR2 (N13537, N13534, N11333);
nor NOR4 (N13538, N13515, N7824, N6368, N11034);
nand NAND2 (N13539, N13523, N2618);
buf BUF1 (N13540, N13537);
nand NAND3 (N13541, N13533, N10784, N10002);
or OR3 (N13542, N13538, N1073, N7026);
xor XOR2 (N13543, N13535, N6734);
and AND2 (N13544, N13539, N11354);
nand NAND3 (N13545, N13536, N10702, N4316);
xor XOR2 (N13546, N13502, N5684);
and AND3 (N13547, N13544, N10928, N9909);
not NOT1 (N13548, N13540);
buf BUF1 (N13549, N13529);
nand NAND2 (N13550, N13545, N9436);
buf BUF1 (N13551, N13541);
or OR3 (N13552, N13550, N6281, N2816);
nand NAND4 (N13553, N13528, N7487, N1653, N9107);
nor NOR3 (N13554, N13542, N10070, N1671);
buf BUF1 (N13555, N13554);
or OR3 (N13556, N13543, N3168, N12431);
nand NAND3 (N13557, N13549, N7435, N5781);
nor NOR3 (N13558, N13551, N6214, N4433);
or OR3 (N13559, N13548, N8458, N12358);
nor NOR2 (N13560, N13546, N2092);
buf BUF1 (N13561, N13559);
nand NAND3 (N13562, N13557, N5134, N12753);
or OR4 (N13563, N13547, N7447, N2019, N7363);
nand NAND4 (N13564, N13562, N2738, N6900, N4707);
not NOT1 (N13565, N13552);
nor NOR2 (N13566, N13558, N7884);
nand NAND3 (N13567, N13565, N677, N11211);
or OR3 (N13568, N13530, N7564, N4182);
not NOT1 (N13569, N13564);
or OR4 (N13570, N13556, N2157, N2582, N6495);
nand NAND3 (N13571, N13570, N8341, N1119);
nand NAND4 (N13572, N13563, N2736, N1381, N10464);
or OR4 (N13573, N13553, N4425, N11926, N1330);
or OR4 (N13574, N13571, N12266, N3952, N7722);
nand NAND4 (N13575, N13567, N3866, N11213, N11243);
buf BUF1 (N13576, N13568);
or OR2 (N13577, N13555, N11608);
buf BUF1 (N13578, N13566);
or OR4 (N13579, N13573, N10742, N7558, N1279);
and AND3 (N13580, N13575, N3563, N12216);
and AND3 (N13581, N13572, N10255, N13069);
and AND4 (N13582, N13569, N6000, N5408, N6186);
buf BUF1 (N13583, N13582);
or OR3 (N13584, N13561, N11470, N13289);
buf BUF1 (N13585, N13580);
and AND2 (N13586, N13577, N2688);
not NOT1 (N13587, N13586);
nor NOR3 (N13588, N13576, N12576, N8995);
or OR4 (N13589, N13587, N7435, N9016, N4146);
xor XOR2 (N13590, N13560, N8359);
nand NAND2 (N13591, N13589, N11590);
and AND2 (N13592, N13585, N2104);
not NOT1 (N13593, N13583);
xor XOR2 (N13594, N13592, N6224);
and AND2 (N13595, N13593, N12841);
nor NOR3 (N13596, N13579, N3475, N423);
xor XOR2 (N13597, N13578, N13581);
nand NAND2 (N13598, N2386, N9864);
nand NAND3 (N13599, N13595, N12136, N5101);
nor NOR4 (N13600, N13597, N1233, N5830, N7270);
or OR2 (N13601, N13598, N7108);
or OR4 (N13602, N13600, N289, N9839, N3584);
and AND4 (N13603, N13591, N1753, N3650, N3893);
nand NAND4 (N13604, N13588, N2585, N8115, N10722);
or OR2 (N13605, N13603, N8869);
or OR2 (N13606, N13599, N12793);
xor XOR2 (N13607, N13590, N8355);
or OR4 (N13608, N13606, N12329, N6043, N542);
and AND2 (N13609, N13594, N11136);
xor XOR2 (N13610, N13602, N7506);
not NOT1 (N13611, N13605);
nor NOR4 (N13612, N13611, N11128, N4019, N6689);
nand NAND2 (N13613, N13596, N2412);
buf BUF1 (N13614, N13604);
or OR2 (N13615, N13609, N8261);
nand NAND2 (N13616, N13614, N3865);
or OR2 (N13617, N13615, N12608);
buf BUF1 (N13618, N13607);
buf BUF1 (N13619, N13616);
nor NOR4 (N13620, N13610, N12336, N6748, N13369);
nor NOR3 (N13621, N13617, N8588, N3558);
not NOT1 (N13622, N13601);
or OR2 (N13623, N13612, N2582);
buf BUF1 (N13624, N13623);
xor XOR2 (N13625, N13622, N9165);
nor NOR2 (N13626, N13621, N3903);
and AND3 (N13627, N13613, N4962, N12024);
not NOT1 (N13628, N13608);
xor XOR2 (N13629, N13618, N9759);
xor XOR2 (N13630, N13629, N4592);
not NOT1 (N13631, N13628);
nor NOR2 (N13632, N13584, N8941);
and AND3 (N13633, N13619, N4673, N7056);
buf BUF1 (N13634, N13632);
not NOT1 (N13635, N13574);
buf BUF1 (N13636, N13630);
not NOT1 (N13637, N13624);
xor XOR2 (N13638, N13620, N10363);
nor NOR4 (N13639, N13625, N8624, N6907, N5813);
and AND4 (N13640, N13634, N8066, N2707, N13014);
buf BUF1 (N13641, N13631);
nor NOR3 (N13642, N13638, N6215, N10904);
nor NOR3 (N13643, N13642, N7664, N7485);
nand NAND4 (N13644, N13635, N10964, N3515, N556);
or OR3 (N13645, N13637, N3730, N8669);
nor NOR2 (N13646, N13643, N6539);
or OR2 (N13647, N13640, N9108);
buf BUF1 (N13648, N13626);
or OR3 (N13649, N13644, N6761, N616);
buf BUF1 (N13650, N13647);
xor XOR2 (N13651, N13641, N2133);
buf BUF1 (N13652, N13648);
and AND4 (N13653, N13636, N11135, N9409, N6382);
buf BUF1 (N13654, N13639);
and AND2 (N13655, N13627, N4450);
xor XOR2 (N13656, N13652, N6391);
and AND3 (N13657, N13650, N44, N4139);
xor XOR2 (N13658, N13654, N10331);
nand NAND4 (N13659, N13649, N9485, N6980, N487);
and AND3 (N13660, N13651, N6601, N11157);
nand NAND3 (N13661, N13655, N6188, N8387);
or OR2 (N13662, N13653, N3094);
not NOT1 (N13663, N13646);
nand NAND4 (N13664, N13656, N175, N7190, N6767);
buf BUF1 (N13665, N13661);
not NOT1 (N13666, N13658);
nand NAND4 (N13667, N13663, N7901, N638, N2410);
and AND4 (N13668, N13659, N1066, N5248, N2995);
nand NAND3 (N13669, N13633, N2339, N8433);
buf BUF1 (N13670, N13662);
nor NOR2 (N13671, N13669, N6060);
xor XOR2 (N13672, N13665, N1975);
xor XOR2 (N13673, N13672, N3719);
or OR2 (N13674, N13664, N9202);
not NOT1 (N13675, N13674);
buf BUF1 (N13676, N13675);
not NOT1 (N13677, N13667);
xor XOR2 (N13678, N13657, N13659);
or OR4 (N13679, N13668, N2051, N7032, N1791);
nor NOR4 (N13680, N13645, N1911, N2166, N11686);
and AND2 (N13681, N13676, N3156);
nor NOR4 (N13682, N13671, N6660, N11790, N6385);
xor XOR2 (N13683, N13666, N9563);
not NOT1 (N13684, N13681);
buf BUF1 (N13685, N13679);
nand NAND4 (N13686, N13677, N11074, N13022, N140);
nand NAND2 (N13687, N13673, N4129);
xor XOR2 (N13688, N13680, N13270);
and AND3 (N13689, N13684, N3856, N1171);
and AND2 (N13690, N13682, N13329);
or OR4 (N13691, N13670, N10278, N11094, N8770);
nor NOR2 (N13692, N13690, N4519);
nand NAND4 (N13693, N13686, N8235, N5975, N10470);
buf BUF1 (N13694, N13688);
buf BUF1 (N13695, N13689);
xor XOR2 (N13696, N13683, N4375);
nor NOR3 (N13697, N13678, N7775, N6443);
buf BUF1 (N13698, N13687);
nand NAND4 (N13699, N13697, N13439, N10781, N5852);
not NOT1 (N13700, N13693);
buf BUF1 (N13701, N13700);
or OR3 (N13702, N13692, N1684, N7983);
xor XOR2 (N13703, N13691, N7161);
and AND2 (N13704, N13701, N10552);
xor XOR2 (N13705, N13704, N2490);
buf BUF1 (N13706, N13698);
and AND4 (N13707, N13702, N7529, N3601, N1188);
nor NOR4 (N13708, N13703, N13416, N7384, N702);
buf BUF1 (N13709, N13660);
nor NOR4 (N13710, N13694, N11706, N8077, N13079);
buf BUF1 (N13711, N13705);
nand NAND2 (N13712, N13685, N8723);
not NOT1 (N13713, N13709);
not NOT1 (N13714, N13696);
or OR2 (N13715, N13708, N2781);
or OR4 (N13716, N13710, N10255, N898, N11096);
nand NAND2 (N13717, N13699, N7639);
not NOT1 (N13718, N13717);
nor NOR2 (N13719, N13713, N7749);
and AND2 (N13720, N13695, N38);
buf BUF1 (N13721, N13716);
and AND4 (N13722, N13720, N12444, N6086, N5741);
and AND4 (N13723, N13714, N1782, N10610, N9357);
and AND3 (N13724, N13707, N5284, N5741);
not NOT1 (N13725, N13723);
xor XOR2 (N13726, N13706, N13062);
not NOT1 (N13727, N13725);
or OR2 (N13728, N13718, N11734);
xor XOR2 (N13729, N13726, N2178);
xor XOR2 (N13730, N13724, N6133);
xor XOR2 (N13731, N13715, N12420);
and AND3 (N13732, N13712, N456, N693);
nor NOR3 (N13733, N13711, N5953, N701);
nand NAND4 (N13734, N13727, N1276, N7830, N9666);
and AND4 (N13735, N13721, N8612, N3669, N7835);
buf BUF1 (N13736, N13734);
buf BUF1 (N13737, N13732);
or OR4 (N13738, N13719, N11478, N7374, N13368);
and AND3 (N13739, N13738, N4978, N6104);
and AND2 (N13740, N13735, N2852);
buf BUF1 (N13741, N13730);
xor XOR2 (N13742, N13729, N2252);
xor XOR2 (N13743, N13728, N1798);
and AND4 (N13744, N13722, N7489, N1486, N9490);
buf BUF1 (N13745, N13740);
nand NAND3 (N13746, N13743, N12729, N10618);
xor XOR2 (N13747, N13744, N9866);
or OR3 (N13748, N13746, N9779, N3472);
buf BUF1 (N13749, N13748);
nand NAND4 (N13750, N13733, N13156, N11969, N2904);
xor XOR2 (N13751, N13747, N1385);
or OR3 (N13752, N13741, N4460, N7958);
or OR3 (N13753, N13751, N5489, N3794);
buf BUF1 (N13754, N13731);
nor NOR2 (N13755, N13737, N970);
not NOT1 (N13756, N13745);
not NOT1 (N13757, N13754);
not NOT1 (N13758, N13753);
nor NOR4 (N13759, N13752, N8579, N3637, N13578);
or OR2 (N13760, N13742, N4818);
nand NAND2 (N13761, N13756, N11432);
not NOT1 (N13762, N13760);
xor XOR2 (N13763, N13739, N12417);
nand NAND3 (N13764, N13762, N7785, N12728);
xor XOR2 (N13765, N13750, N1638);
and AND3 (N13766, N13758, N10210, N12986);
nor NOR3 (N13767, N13755, N6924, N9846);
and AND3 (N13768, N13749, N10042, N11985);
xor XOR2 (N13769, N13757, N8000);
or OR2 (N13770, N13765, N4168);
nor NOR4 (N13771, N13764, N9088, N6991, N11892);
nand NAND3 (N13772, N13766, N8800, N7682);
xor XOR2 (N13773, N13769, N9701);
nor NOR3 (N13774, N13761, N1728, N4688);
buf BUF1 (N13775, N13772);
buf BUF1 (N13776, N13763);
nand NAND2 (N13777, N13774, N12227);
not NOT1 (N13778, N13771);
nand NAND3 (N13779, N13776, N2169, N1783);
buf BUF1 (N13780, N13775);
and AND3 (N13781, N13770, N11035, N12570);
or OR3 (N13782, N13778, N11781, N5583);
and AND2 (N13783, N13781, N2093);
or OR3 (N13784, N13777, N10313, N7324);
not NOT1 (N13785, N13782);
not NOT1 (N13786, N13785);
nand NAND2 (N13787, N13786, N1153);
xor XOR2 (N13788, N13767, N1231);
xor XOR2 (N13789, N13783, N963);
nand NAND2 (N13790, N13784, N5011);
nor NOR3 (N13791, N13779, N9974, N5297);
not NOT1 (N13792, N13759);
or OR2 (N13793, N13787, N13331);
and AND4 (N13794, N13789, N12355, N8258, N7132);
nand NAND3 (N13795, N13780, N7671, N4061);
buf BUF1 (N13796, N13773);
nand NAND3 (N13797, N13795, N10618, N9874);
nand NAND3 (N13798, N13796, N13143, N13562);
or OR2 (N13799, N13797, N8484);
nand NAND2 (N13800, N13791, N2060);
and AND3 (N13801, N13768, N434, N10972);
not NOT1 (N13802, N13736);
and AND2 (N13803, N13799, N6791);
nand NAND2 (N13804, N13801, N658);
not NOT1 (N13805, N13793);
nand NAND4 (N13806, N13790, N1094, N11691, N10331);
nor NOR2 (N13807, N13804, N2358);
and AND2 (N13808, N13807, N7076);
and AND4 (N13809, N13798, N6156, N7857, N4092);
and AND3 (N13810, N13802, N10677, N6776);
and AND3 (N13811, N13794, N13473, N12670);
xor XOR2 (N13812, N13800, N8425);
and AND4 (N13813, N13809, N9606, N12429, N7049);
buf BUF1 (N13814, N13803);
buf BUF1 (N13815, N13805);
or OR3 (N13816, N13814, N946, N4872);
xor XOR2 (N13817, N13811, N10582);
or OR3 (N13818, N13808, N778, N5315);
and AND4 (N13819, N13812, N12232, N12133, N5480);
nand NAND4 (N13820, N13806, N7767, N12996, N3505);
nor NOR2 (N13821, N13816, N8375);
nor NOR4 (N13822, N13810, N1895, N11424, N10972);
and AND3 (N13823, N13821, N11212, N11462);
nand NAND2 (N13824, N13822, N2731);
or OR3 (N13825, N13820, N12238, N11340);
not NOT1 (N13826, N13815);
not NOT1 (N13827, N13823);
nand NAND3 (N13828, N13788, N11438, N2497);
nor NOR4 (N13829, N13827, N12903, N2295, N5039);
not NOT1 (N13830, N13819);
nand NAND2 (N13831, N13825, N1571);
buf BUF1 (N13832, N13828);
or OR2 (N13833, N13824, N3017);
and AND2 (N13834, N13792, N1014);
not NOT1 (N13835, N13830);
nor NOR4 (N13836, N13826, N12376, N8378, N2032);
not NOT1 (N13837, N13818);
or OR3 (N13838, N13817, N2032, N1199);
and AND2 (N13839, N13836, N7500);
and AND4 (N13840, N13831, N2192, N2033, N9369);
buf BUF1 (N13841, N13834);
and AND2 (N13842, N13841, N1786);
buf BUF1 (N13843, N13829);
xor XOR2 (N13844, N13842, N9916);
or OR4 (N13845, N13813, N10825, N7055, N8820);
nor NOR3 (N13846, N13839, N2051, N4117);
not NOT1 (N13847, N13846);
nor NOR2 (N13848, N13835, N9132);
buf BUF1 (N13849, N13833);
not NOT1 (N13850, N13840);
not NOT1 (N13851, N13847);
buf BUF1 (N13852, N13844);
nor NOR4 (N13853, N13852, N9733, N13411, N5300);
nor NOR2 (N13854, N13837, N7481);
and AND3 (N13855, N13849, N3665, N823);
buf BUF1 (N13856, N13838);
buf BUF1 (N13857, N13845);
xor XOR2 (N13858, N13853, N11047);
not NOT1 (N13859, N13832);
nor NOR2 (N13860, N13859, N5462);
buf BUF1 (N13861, N13851);
nor NOR4 (N13862, N13858, N9230, N5908, N12134);
or OR4 (N13863, N13850, N11825, N834, N10029);
buf BUF1 (N13864, N13855);
not NOT1 (N13865, N13860);
or OR3 (N13866, N13843, N3308, N5526);
and AND3 (N13867, N13865, N3321, N1408);
xor XOR2 (N13868, N13866, N7513);
nand NAND3 (N13869, N13867, N12730, N12778);
nor NOR3 (N13870, N13862, N7680, N9211);
and AND2 (N13871, N13869, N8958);
xor XOR2 (N13872, N13861, N3803);
xor XOR2 (N13873, N13848, N150);
buf BUF1 (N13874, N13863);
xor XOR2 (N13875, N13872, N2983);
xor XOR2 (N13876, N13857, N7665);
and AND3 (N13877, N13870, N652, N7898);
not NOT1 (N13878, N13856);
xor XOR2 (N13879, N13864, N10116);
not NOT1 (N13880, N13875);
xor XOR2 (N13881, N13854, N4988);
nor NOR2 (N13882, N13874, N2545);
nand NAND4 (N13883, N13879, N1873, N8946, N5542);
buf BUF1 (N13884, N13880);
nor NOR3 (N13885, N13871, N12288, N5122);
not NOT1 (N13886, N13881);
nor NOR3 (N13887, N13885, N13218, N9255);
or OR3 (N13888, N13884, N5, N4569);
and AND4 (N13889, N13878, N7593, N6392, N5013);
xor XOR2 (N13890, N13888, N471);
not NOT1 (N13891, N13889);
and AND4 (N13892, N13890, N10019, N11252, N7651);
nor NOR4 (N13893, N13868, N3013, N5146, N8465);
nor NOR3 (N13894, N13887, N4695, N597);
nand NAND4 (N13895, N13876, N3728, N10473, N10106);
and AND3 (N13896, N13882, N6491, N7683);
and AND4 (N13897, N13894, N11719, N6533, N13726);
nor NOR3 (N13898, N13895, N8853, N6468);
buf BUF1 (N13899, N13877);
nor NOR4 (N13900, N13899, N1257, N10119, N11222);
buf BUF1 (N13901, N13898);
buf BUF1 (N13902, N13892);
nor NOR4 (N13903, N13902, N6020, N4686, N1108);
not NOT1 (N13904, N13897);
nand NAND4 (N13905, N13893, N5298, N8643, N8979);
not NOT1 (N13906, N13883);
xor XOR2 (N13907, N13886, N9366);
not NOT1 (N13908, N13903);
nand NAND2 (N13909, N13906, N2896);
and AND3 (N13910, N13904, N8987, N7765);
and AND3 (N13911, N13905, N3818, N820);
nand NAND2 (N13912, N13911, N3636);
not NOT1 (N13913, N13908);
xor XOR2 (N13914, N13912, N8145);
buf BUF1 (N13915, N13910);
nor NOR4 (N13916, N13915, N2158, N2679, N8419);
xor XOR2 (N13917, N13900, N2068);
nand NAND4 (N13918, N13891, N1525, N4090, N757);
or OR4 (N13919, N13907, N666, N9934, N10484);
and AND2 (N13920, N13918, N7261);
xor XOR2 (N13921, N13916, N9112);
and AND3 (N13922, N13909, N12254, N1054);
nor NOR2 (N13923, N13896, N1955);
nand NAND3 (N13924, N13873, N7539, N9049);
and AND2 (N13925, N13920, N10372);
and AND2 (N13926, N13924, N547);
or OR4 (N13927, N13926, N7791, N8478, N12625);
nand NAND4 (N13928, N13901, N9648, N7558, N10988);
nand NAND3 (N13929, N13922, N5107, N2919);
xor XOR2 (N13930, N13928, N12504);
and AND4 (N13931, N13930, N591, N4137, N8002);
xor XOR2 (N13932, N13914, N8341);
and AND3 (N13933, N13931, N2309, N10246);
and AND3 (N13934, N13932, N1300, N11094);
xor XOR2 (N13935, N13919, N11149);
buf BUF1 (N13936, N13917);
and AND2 (N13937, N13925, N9267);
nor NOR3 (N13938, N13935, N5086, N4460);
and AND4 (N13939, N13933, N691, N284, N7749);
not NOT1 (N13940, N13921);
and AND2 (N13941, N13937, N12054);
buf BUF1 (N13942, N13913);
nand NAND3 (N13943, N13942, N8897, N3981);
buf BUF1 (N13944, N13938);
or OR3 (N13945, N13929, N6626, N11005);
not NOT1 (N13946, N13941);
not NOT1 (N13947, N13934);
not NOT1 (N13948, N13927);
not NOT1 (N13949, N13939);
nor NOR4 (N13950, N13923, N5785, N8564, N1480);
or OR2 (N13951, N13940, N9281);
nor NOR4 (N13952, N13948, N1426, N5973, N13019);
nand NAND4 (N13953, N13945, N2123, N3595, N10961);
or OR4 (N13954, N13943, N4090, N9, N3132);
xor XOR2 (N13955, N13950, N10681);
not NOT1 (N13956, N13936);
nand NAND3 (N13957, N13952, N4357, N10497);
or OR4 (N13958, N13946, N4539, N2787, N9017);
buf BUF1 (N13959, N13947);
not NOT1 (N13960, N13957);
buf BUF1 (N13961, N13960);
buf BUF1 (N13962, N13958);
nor NOR4 (N13963, N13955, N1552, N906, N2130);
and AND3 (N13964, N13962, N11100, N13108);
nand NAND4 (N13965, N13963, N6178, N499, N7192);
not NOT1 (N13966, N13965);
and AND3 (N13967, N13961, N1382, N2099);
nor NOR3 (N13968, N13967, N717, N818);
buf BUF1 (N13969, N13959);
nor NOR3 (N13970, N13954, N12626, N11286);
and AND2 (N13971, N13970, N6857);
not NOT1 (N13972, N13964);
or OR3 (N13973, N13949, N11654, N4098);
buf BUF1 (N13974, N13973);
buf BUF1 (N13975, N13951);
and AND4 (N13976, N13974, N2483, N10590, N7992);
nor NOR3 (N13977, N13972, N6798, N6489);
nand NAND2 (N13978, N13956, N1066);
or OR3 (N13979, N13977, N3852, N6821);
or OR4 (N13980, N13978, N325, N1056, N8024);
or OR2 (N13981, N13975, N4912);
and AND3 (N13982, N13968, N3402, N13498);
buf BUF1 (N13983, N13953);
xor XOR2 (N13984, N13979, N9981);
xor XOR2 (N13985, N13944, N8864);
xor XOR2 (N13986, N13971, N2856);
nor NOR4 (N13987, N13986, N5077, N12269, N6359);
buf BUF1 (N13988, N13981);
or OR4 (N13989, N13966, N7620, N13276, N5268);
nor NOR3 (N13990, N13980, N5888, N10054);
or OR4 (N13991, N13985, N1552, N5421, N6525);
not NOT1 (N13992, N13982);
nand NAND3 (N13993, N13983, N7938, N1496);
xor XOR2 (N13994, N13987, N6274);
or OR3 (N13995, N13984, N13660, N8865);
buf BUF1 (N13996, N13995);
not NOT1 (N13997, N13988);
nor NOR2 (N13998, N13991, N6337);
and AND2 (N13999, N13993, N1129);
nor NOR2 (N14000, N13997, N13012);
nor NOR3 (N14001, N13969, N3598, N8800);
buf BUF1 (N14002, N14001);
and AND4 (N14003, N13998, N12642, N13751, N2295);
xor XOR2 (N14004, N13992, N204);
nor NOR2 (N14005, N13989, N1476);
not NOT1 (N14006, N14002);
buf BUF1 (N14007, N13996);
not NOT1 (N14008, N14004);
buf BUF1 (N14009, N13976);
not NOT1 (N14010, N14005);
nand NAND2 (N14011, N13999, N6858);
buf BUF1 (N14012, N14007);
nor NOR2 (N14013, N14011, N8092);
buf BUF1 (N14014, N14003);
xor XOR2 (N14015, N13994, N3206);
and AND2 (N14016, N14008, N4112);
buf BUF1 (N14017, N14014);
buf BUF1 (N14018, N14006);
nand NAND4 (N14019, N14012, N2177, N2355, N9236);
buf BUF1 (N14020, N13990);
not NOT1 (N14021, N14018);
buf BUF1 (N14022, N14020);
nor NOR2 (N14023, N14022, N7387);
nor NOR2 (N14024, N14016, N2661);
xor XOR2 (N14025, N14013, N6989);
not NOT1 (N14026, N14023);
not NOT1 (N14027, N14015);
not NOT1 (N14028, N14017);
and AND4 (N14029, N14024, N12697, N1349, N10342);
buf BUF1 (N14030, N14027);
buf BUF1 (N14031, N14021);
buf BUF1 (N14032, N14019);
not NOT1 (N14033, N14000);
nand NAND2 (N14034, N14028, N7656);
and AND2 (N14035, N14010, N9264);
buf BUF1 (N14036, N14029);
buf BUF1 (N14037, N14026);
nand NAND3 (N14038, N14033, N9048, N3429);
and AND4 (N14039, N14034, N10958, N9972, N6016);
xor XOR2 (N14040, N14030, N6395);
buf BUF1 (N14041, N14009);
nor NOR4 (N14042, N14035, N10065, N1916, N1191);
nor NOR3 (N14043, N14040, N2760, N1769);
xor XOR2 (N14044, N14038, N10489);
and AND3 (N14045, N14032, N6807, N4821);
or OR4 (N14046, N14036, N8666, N9628, N5608);
not NOT1 (N14047, N14042);
buf BUF1 (N14048, N14037);
or OR4 (N14049, N14047, N1551, N11283, N5072);
or OR2 (N14050, N14043, N9380);
buf BUF1 (N14051, N14049);
not NOT1 (N14052, N14031);
nand NAND2 (N14053, N14025, N3377);
not NOT1 (N14054, N14053);
buf BUF1 (N14055, N14045);
or OR2 (N14056, N14046, N7680);
or OR3 (N14057, N14050, N10759, N13021);
xor XOR2 (N14058, N14051, N7562);
nor NOR2 (N14059, N14057, N1162);
not NOT1 (N14060, N14054);
xor XOR2 (N14061, N14041, N1744);
buf BUF1 (N14062, N14061);
or OR2 (N14063, N14058, N13169);
nand NAND3 (N14064, N14056, N9709, N9453);
nand NAND4 (N14065, N14062, N8212, N4314, N6427);
nor NOR2 (N14066, N14065, N1617);
and AND2 (N14067, N14052, N7281);
buf BUF1 (N14068, N14066);
xor XOR2 (N14069, N14060, N8782);
nand NAND4 (N14070, N14064, N5726, N5408, N6005);
and AND4 (N14071, N14039, N5690, N640, N3096);
buf BUF1 (N14072, N14063);
not NOT1 (N14073, N14044);
not NOT1 (N14074, N14071);
or OR4 (N14075, N14072, N4788, N2461, N6385);
or OR3 (N14076, N14059, N2855, N13449);
nand NAND4 (N14077, N14070, N12061, N12764, N1438);
nand NAND2 (N14078, N14073, N11204);
not NOT1 (N14079, N14077);
not NOT1 (N14080, N14076);
or OR4 (N14081, N14075, N12385, N9029, N8098);
nand NAND4 (N14082, N14081, N6993, N9152, N884);
nor NOR3 (N14083, N14074, N8726, N10816);
nor NOR2 (N14084, N14083, N9499);
or OR3 (N14085, N14048, N2155, N8035);
nand NAND2 (N14086, N14084, N4514);
or OR3 (N14087, N14086, N3778, N3254);
xor XOR2 (N14088, N14082, N650);
nand NAND3 (N14089, N14085, N1310, N12890);
xor XOR2 (N14090, N14088, N9481);
buf BUF1 (N14091, N14080);
nand NAND3 (N14092, N14091, N7283, N12713);
nand NAND4 (N14093, N14067, N12019, N12291, N2829);
nor NOR2 (N14094, N14055, N9047);
or OR2 (N14095, N14093, N7230);
or OR2 (N14096, N14094, N12668);
and AND3 (N14097, N14092, N5048, N7422);
or OR4 (N14098, N14079, N14028, N8040, N12056);
and AND3 (N14099, N14089, N8238, N3674);
buf BUF1 (N14100, N14096);
buf BUF1 (N14101, N14068);
xor XOR2 (N14102, N14069, N8987);
and AND4 (N14103, N14101, N7385, N11083, N440);
nor NOR2 (N14104, N14095, N4850);
and AND3 (N14105, N14098, N10182, N12210);
nor NOR2 (N14106, N14097, N7749);
nor NOR4 (N14107, N14078, N1074, N6284, N11946);
not NOT1 (N14108, N14100);
or OR4 (N14109, N14108, N9937, N3251, N12569);
nand NAND2 (N14110, N14087, N4137);
nor NOR3 (N14111, N14090, N11243, N10174);
nand NAND3 (N14112, N14110, N4003, N7658);
and AND4 (N14113, N14103, N13447, N10851, N9721);
not NOT1 (N14114, N14107);
nand NAND3 (N14115, N14109, N3326, N42);
xor XOR2 (N14116, N14105, N4897);
and AND3 (N14117, N14111, N8402, N13301);
or OR3 (N14118, N14099, N4438, N11097);
buf BUF1 (N14119, N14113);
xor XOR2 (N14120, N14118, N6343);
or OR3 (N14121, N14117, N2488, N2319);
or OR3 (N14122, N14115, N11959, N415);
xor XOR2 (N14123, N14104, N9990);
nor NOR4 (N14124, N14123, N11779, N11884, N10888);
nand NAND4 (N14125, N14112, N4721, N3493, N754);
not NOT1 (N14126, N14122);
xor XOR2 (N14127, N14124, N2680);
and AND2 (N14128, N14127, N5369);
and AND2 (N14129, N14125, N8425);
and AND4 (N14130, N14119, N6637, N127, N11798);
nor NOR3 (N14131, N14116, N13297, N2464);
buf BUF1 (N14132, N14114);
nor NOR3 (N14133, N14120, N102, N10985);
nand NAND2 (N14134, N14102, N12563);
and AND4 (N14135, N14129, N10914, N9399, N12048);
not NOT1 (N14136, N14128);
nand NAND3 (N14137, N14121, N2246, N7709);
buf BUF1 (N14138, N14130);
and AND2 (N14139, N14133, N287);
nand NAND2 (N14140, N14131, N8826);
xor XOR2 (N14141, N14132, N13099);
nand NAND3 (N14142, N14134, N9596, N5284);
buf BUF1 (N14143, N14138);
and AND3 (N14144, N14140, N11865, N4539);
xor XOR2 (N14145, N14136, N12118);
and AND3 (N14146, N14145, N12096, N11177);
or OR3 (N14147, N14139, N11761, N1496);
buf BUF1 (N14148, N14142);
or OR2 (N14149, N14137, N3783);
and AND3 (N14150, N14126, N13987, N4177);
and AND3 (N14151, N14147, N13823, N1140);
nand NAND4 (N14152, N14146, N697, N408, N8695);
nand NAND4 (N14153, N14144, N5431, N10949, N8084);
or OR4 (N14154, N14141, N10992, N7278, N11148);
nand NAND2 (N14155, N14153, N2628);
and AND2 (N14156, N14152, N1587);
buf BUF1 (N14157, N14155);
and AND3 (N14158, N14150, N4173, N3357);
or OR4 (N14159, N14106, N3863, N9524, N4529);
xor XOR2 (N14160, N14154, N8058);
and AND4 (N14161, N14135, N1866, N9002, N11614);
xor XOR2 (N14162, N14158, N11674);
not NOT1 (N14163, N14149);
or OR2 (N14164, N14159, N5441);
xor XOR2 (N14165, N14162, N2460);
and AND2 (N14166, N14151, N785);
xor XOR2 (N14167, N14164, N12675);
and AND2 (N14168, N14157, N12083);
buf BUF1 (N14169, N14143);
xor XOR2 (N14170, N14166, N5865);
buf BUF1 (N14171, N14148);
buf BUF1 (N14172, N14165);
buf BUF1 (N14173, N14172);
xor XOR2 (N14174, N14161, N3619);
or OR4 (N14175, N14171, N11071, N13678, N2178);
nor NOR4 (N14176, N14174, N4542, N952, N1857);
nand NAND3 (N14177, N14160, N13357, N9748);
nor NOR2 (N14178, N14170, N7962);
nand NAND4 (N14179, N14176, N3172, N8616, N13338);
nand NAND3 (N14180, N14175, N10964, N4377);
xor XOR2 (N14181, N14179, N1721);
not NOT1 (N14182, N14178);
nor NOR2 (N14183, N14173, N4900);
buf BUF1 (N14184, N14169);
not NOT1 (N14185, N14181);
buf BUF1 (N14186, N14182);
nand NAND4 (N14187, N14163, N8359, N13432, N793);
and AND2 (N14188, N14184, N890);
or OR4 (N14189, N14186, N2584, N3080, N12544);
not NOT1 (N14190, N14187);
nor NOR3 (N14191, N14168, N13532, N6589);
and AND4 (N14192, N14167, N7943, N10354, N7635);
not NOT1 (N14193, N14191);
nand NAND3 (N14194, N14156, N4480, N2982);
nand NAND2 (N14195, N14183, N1663);
and AND2 (N14196, N14185, N7384);
not NOT1 (N14197, N14190);
xor XOR2 (N14198, N14189, N2770);
and AND4 (N14199, N14180, N8637, N10743, N13503);
or OR2 (N14200, N14177, N4797);
buf BUF1 (N14201, N14199);
and AND3 (N14202, N14192, N6369, N9613);
xor XOR2 (N14203, N14193, N9536);
nand NAND3 (N14204, N14203, N3682, N10228);
buf BUF1 (N14205, N14200);
buf BUF1 (N14206, N14194);
or OR2 (N14207, N14195, N8475);
or OR2 (N14208, N14205, N6146);
nor NOR2 (N14209, N14196, N11881);
or OR4 (N14210, N14202, N11745, N5158, N5245);
nand NAND3 (N14211, N14197, N4336, N586);
buf BUF1 (N14212, N14211);
xor XOR2 (N14213, N14198, N6100);
xor XOR2 (N14214, N14207, N4091);
or OR3 (N14215, N14212, N1742, N12467);
nand NAND3 (N14216, N14188, N7213, N5362);
buf BUF1 (N14217, N14208);
nand NAND4 (N14218, N14215, N3851, N5344, N9328);
xor XOR2 (N14219, N14209, N1765);
nand NAND2 (N14220, N14201, N1674);
and AND3 (N14221, N14206, N10115, N124);
not NOT1 (N14222, N14214);
and AND4 (N14223, N14221, N7079, N8832, N1479);
xor XOR2 (N14224, N14216, N439);
or OR2 (N14225, N14223, N8637);
nand NAND2 (N14226, N14210, N6384);
nor NOR3 (N14227, N14204, N12617, N6070);
nand NAND4 (N14228, N14224, N8222, N1338, N1621);
nand NAND3 (N14229, N14217, N2074, N12544);
nand NAND4 (N14230, N14213, N8232, N599, N3181);
xor XOR2 (N14231, N14226, N12228);
and AND3 (N14232, N14220, N2979, N5038);
nor NOR4 (N14233, N14227, N10631, N14088, N5647);
and AND2 (N14234, N14232, N10672);
nor NOR2 (N14235, N14229, N10672);
not NOT1 (N14236, N14233);
not NOT1 (N14237, N14235);
nand NAND2 (N14238, N14219, N5920);
nor NOR2 (N14239, N14230, N13228);
not NOT1 (N14240, N14228);
or OR3 (N14241, N14222, N1946, N14057);
buf BUF1 (N14242, N14239);
nand NAND4 (N14243, N14231, N12792, N13425, N11047);
xor XOR2 (N14244, N14241, N12290);
or OR3 (N14245, N14243, N12870, N1633);
xor XOR2 (N14246, N14225, N11649);
nand NAND4 (N14247, N14246, N11605, N5780, N2710);
xor XOR2 (N14248, N14245, N6647);
xor XOR2 (N14249, N14238, N37);
nand NAND2 (N14250, N14237, N898);
not NOT1 (N14251, N14244);
nor NOR4 (N14252, N14236, N11599, N9956, N2883);
not NOT1 (N14253, N14247);
nor NOR2 (N14254, N14252, N7241);
and AND4 (N14255, N14253, N6405, N9943, N3217);
xor XOR2 (N14256, N14234, N4595);
xor XOR2 (N14257, N14255, N7383);
and AND4 (N14258, N14249, N9662, N1382, N5970);
and AND2 (N14259, N14258, N1930);
or OR3 (N14260, N14240, N8499, N8544);
and AND3 (N14261, N14250, N13189, N12857);
buf BUF1 (N14262, N14259);
and AND3 (N14263, N14260, N14175, N9839);
not NOT1 (N14264, N14242);
nor NOR4 (N14265, N14256, N6982, N14107, N902);
and AND3 (N14266, N14248, N2807, N3902);
not NOT1 (N14267, N14263);
not NOT1 (N14268, N14251);
nand NAND4 (N14269, N14261, N10740, N3604, N7972);
or OR2 (N14270, N14265, N11928);
nor NOR2 (N14271, N14267, N13740);
not NOT1 (N14272, N14254);
not NOT1 (N14273, N14272);
buf BUF1 (N14274, N14266);
nand NAND3 (N14275, N14269, N2697, N1547);
xor XOR2 (N14276, N14262, N11262);
or OR2 (N14277, N14218, N13207);
nand NAND3 (N14278, N14276, N4019, N3415);
nand NAND2 (N14279, N14271, N3356);
buf BUF1 (N14280, N14273);
or OR3 (N14281, N14274, N9453, N978);
xor XOR2 (N14282, N14264, N13178);
buf BUF1 (N14283, N14279);
xor XOR2 (N14284, N14282, N2030);
xor XOR2 (N14285, N14283, N3853);
buf BUF1 (N14286, N14268);
xor XOR2 (N14287, N14270, N8123);
xor XOR2 (N14288, N14277, N13093);
not NOT1 (N14289, N14287);
not NOT1 (N14290, N14289);
nor NOR3 (N14291, N14284, N11962, N357);
buf BUF1 (N14292, N14280);
and AND2 (N14293, N14291, N13443);
nor NOR3 (N14294, N14275, N4848, N10919);
buf BUF1 (N14295, N14257);
and AND2 (N14296, N14292, N3132);
nor NOR3 (N14297, N14281, N8041, N891);
buf BUF1 (N14298, N14285);
nand NAND4 (N14299, N14293, N2617, N8650, N10350);
buf BUF1 (N14300, N14299);
xor XOR2 (N14301, N14288, N9786);
xor XOR2 (N14302, N14300, N8374);
not NOT1 (N14303, N14294);
not NOT1 (N14304, N14302);
and AND2 (N14305, N14286, N8828);
and AND2 (N14306, N14303, N3358);
or OR4 (N14307, N14295, N3269, N11235, N8840);
xor XOR2 (N14308, N14301, N11841);
nor NOR2 (N14309, N14296, N78);
and AND2 (N14310, N14305, N4176);
and AND2 (N14311, N14297, N662);
and AND2 (N14312, N14304, N2125);
nand NAND4 (N14313, N14311, N3306, N7178, N10776);
not NOT1 (N14314, N14309);
and AND2 (N14315, N14298, N3764);
nand NAND3 (N14316, N14278, N12213, N9474);
xor XOR2 (N14317, N14290, N7108);
not NOT1 (N14318, N14306);
buf BUF1 (N14319, N14307);
and AND3 (N14320, N14315, N3801, N1991);
xor XOR2 (N14321, N14313, N6857);
nand NAND3 (N14322, N14321, N12286, N13917);
and AND3 (N14323, N14310, N278, N8716);
xor XOR2 (N14324, N14317, N6454);
nand NAND3 (N14325, N14320, N8184, N10854);
or OR4 (N14326, N14319, N13258, N2109, N13493);
nor NOR4 (N14327, N14312, N14263, N1735, N13717);
nand NAND3 (N14328, N14308, N12774, N8613);
nor NOR2 (N14329, N14322, N40);
nand NAND2 (N14330, N14326, N6842);
nand NAND3 (N14331, N14318, N2385, N13048);
nand NAND4 (N14332, N14330, N8871, N5799, N7784);
buf BUF1 (N14333, N14331);
xor XOR2 (N14334, N14323, N7502);
not NOT1 (N14335, N14332);
and AND3 (N14336, N14316, N8531, N11300);
not NOT1 (N14337, N14333);
not NOT1 (N14338, N14325);
nor NOR2 (N14339, N14328, N8790);
not NOT1 (N14340, N14338);
nor NOR3 (N14341, N14329, N345, N2302);
xor XOR2 (N14342, N14327, N5208);
xor XOR2 (N14343, N14342, N5541);
or OR3 (N14344, N14336, N3803, N11350);
nand NAND3 (N14345, N14341, N6762, N9078);
buf BUF1 (N14346, N14344);
and AND2 (N14347, N14345, N4411);
or OR3 (N14348, N14334, N10358, N4716);
xor XOR2 (N14349, N14324, N11511);
buf BUF1 (N14350, N14347);
and AND4 (N14351, N14337, N6927, N10748, N7193);
nor NOR4 (N14352, N14349, N13007, N11746, N4060);
xor XOR2 (N14353, N14350, N1033);
or OR2 (N14354, N14353, N12550);
nor NOR3 (N14355, N14335, N9908, N3372);
or OR3 (N14356, N14343, N285, N12454);
nand NAND4 (N14357, N14340, N260, N341, N11023);
and AND4 (N14358, N14354, N3286, N10174, N4483);
nand NAND2 (N14359, N14348, N9003);
buf BUF1 (N14360, N14314);
or OR2 (N14361, N14356, N11410);
buf BUF1 (N14362, N14360);
buf BUF1 (N14363, N14358);
nand NAND3 (N14364, N14351, N11837, N2829);
xor XOR2 (N14365, N14362, N8219);
not NOT1 (N14366, N14355);
and AND3 (N14367, N14361, N3219, N4368);
not NOT1 (N14368, N14365);
buf BUF1 (N14369, N14346);
not NOT1 (N14370, N14364);
buf BUF1 (N14371, N14370);
nand NAND2 (N14372, N14367, N12783);
nor NOR2 (N14373, N14357, N12944);
not NOT1 (N14374, N14371);
nand NAND4 (N14375, N14366, N9154, N11559, N9428);
nand NAND2 (N14376, N14373, N13304);
nor NOR2 (N14377, N14368, N7642);
nand NAND3 (N14378, N14377, N7073, N2994);
nand NAND4 (N14379, N14374, N9233, N7491, N3909);
nand NAND3 (N14380, N14378, N3429, N2434);
not NOT1 (N14381, N14359);
and AND2 (N14382, N14372, N11967);
nor NOR3 (N14383, N14363, N13587, N1191);
nor NOR4 (N14384, N14376, N13804, N5778, N11563);
not NOT1 (N14385, N14375);
or OR3 (N14386, N14369, N13816, N6654);
or OR2 (N14387, N14383, N13393);
nor NOR3 (N14388, N14385, N3214, N10400);
nand NAND4 (N14389, N14381, N9145, N7250, N886);
or OR4 (N14390, N14382, N13578, N11364, N1027);
nand NAND4 (N14391, N14387, N10346, N323, N6075);
not NOT1 (N14392, N14390);
not NOT1 (N14393, N14391);
not NOT1 (N14394, N14379);
nand NAND4 (N14395, N14386, N4904, N9300, N4599);
nor NOR2 (N14396, N14393, N1097);
nor NOR2 (N14397, N14392, N6200);
nand NAND2 (N14398, N14352, N12218);
nor NOR4 (N14399, N14389, N3201, N7206, N7557);
nor NOR4 (N14400, N14388, N958, N8428, N2866);
xor XOR2 (N14401, N14397, N2938);
or OR3 (N14402, N14380, N4023, N9252);
buf BUF1 (N14403, N14396);
nand NAND4 (N14404, N14401, N13285, N3984, N195);
xor XOR2 (N14405, N14384, N5029);
nand NAND3 (N14406, N14405, N5470, N870);
buf BUF1 (N14407, N14394);
xor XOR2 (N14408, N14407, N9226);
xor XOR2 (N14409, N14400, N13054);
or OR2 (N14410, N14409, N9379);
or OR3 (N14411, N14398, N571, N4585);
not NOT1 (N14412, N14402);
not NOT1 (N14413, N14408);
xor XOR2 (N14414, N14403, N7794);
nand NAND3 (N14415, N14404, N11192, N3426);
or OR2 (N14416, N14415, N211);
not NOT1 (N14417, N14411);
not NOT1 (N14418, N14339);
xor XOR2 (N14419, N14417, N4161);
nand NAND3 (N14420, N14418, N7719, N10717);
not NOT1 (N14421, N14399);
and AND3 (N14422, N14410, N11442, N5281);
not NOT1 (N14423, N14416);
or OR2 (N14424, N14406, N7773);
nand NAND3 (N14425, N14420, N5489, N10627);
buf BUF1 (N14426, N14419);
nor NOR2 (N14427, N14422, N11012);
nor NOR4 (N14428, N14425, N13624, N11222, N8653);
xor XOR2 (N14429, N14426, N4705);
xor XOR2 (N14430, N14413, N7931);
nor NOR3 (N14431, N14395, N4489, N10067);
nor NOR3 (N14432, N14430, N13251, N12419);
xor XOR2 (N14433, N14427, N9486);
nand NAND4 (N14434, N14429, N7849, N9954, N9056);
nor NOR2 (N14435, N14431, N10215);
buf BUF1 (N14436, N14434);
nor NOR3 (N14437, N14424, N8092, N11667);
buf BUF1 (N14438, N14436);
buf BUF1 (N14439, N14437);
xor XOR2 (N14440, N14433, N7505);
buf BUF1 (N14441, N14435);
nor NOR2 (N14442, N14412, N13715);
not NOT1 (N14443, N14414);
or OR3 (N14444, N14439, N3317, N12917);
nor NOR3 (N14445, N14442, N5001, N7038);
nor NOR4 (N14446, N14443, N8244, N4950, N4246);
xor XOR2 (N14447, N14445, N8282);
nor NOR2 (N14448, N14440, N13661);
or OR3 (N14449, N14438, N7950, N1433);
buf BUF1 (N14450, N14447);
nor NOR4 (N14451, N14448, N4581, N7402, N13401);
and AND3 (N14452, N14432, N1135, N10330);
buf BUF1 (N14453, N14423);
buf BUF1 (N14454, N14444);
nand NAND2 (N14455, N14446, N12851);
or OR3 (N14456, N14449, N10110, N10341);
or OR3 (N14457, N14456, N785, N2439);
buf BUF1 (N14458, N14421);
or OR2 (N14459, N14451, N8373);
nand NAND3 (N14460, N14457, N8043, N11300);
buf BUF1 (N14461, N14454);
buf BUF1 (N14462, N14450);
and AND3 (N14463, N14462, N13983, N7476);
xor XOR2 (N14464, N14461, N4548);
or OR2 (N14465, N14464, N4481);
nand NAND4 (N14466, N14465, N3326, N10564, N8400);
buf BUF1 (N14467, N14455);
and AND4 (N14468, N14460, N355, N3502, N10226);
not NOT1 (N14469, N14428);
buf BUF1 (N14470, N14468);
and AND3 (N14471, N14463, N11576, N2671);
buf BUF1 (N14472, N14466);
or OR2 (N14473, N14471, N4689);
nor NOR2 (N14474, N14459, N1569);
buf BUF1 (N14475, N14453);
and AND3 (N14476, N14452, N2090, N4439);
and AND4 (N14477, N14441, N3005, N14384, N5267);
or OR2 (N14478, N14475, N3575);
or OR3 (N14479, N14477, N6073, N3012);
or OR4 (N14480, N14479, N3639, N1124, N11577);
and AND2 (N14481, N14469, N9644);
not NOT1 (N14482, N14472);
buf BUF1 (N14483, N14480);
nor NOR2 (N14484, N14481, N5228);
nand NAND3 (N14485, N14482, N1155, N10823);
and AND2 (N14486, N14474, N9315);
buf BUF1 (N14487, N14458);
xor XOR2 (N14488, N14467, N13609);
and AND2 (N14489, N14483, N5722);
and AND2 (N14490, N14486, N7150);
nor NOR4 (N14491, N14476, N3516, N7679, N13001);
xor XOR2 (N14492, N14487, N228);
nand NAND2 (N14493, N14488, N8425);
buf BUF1 (N14494, N14484);
nor NOR3 (N14495, N14470, N6677, N1256);
not NOT1 (N14496, N14485);
not NOT1 (N14497, N14490);
nand NAND2 (N14498, N14492, N12675);
nand NAND4 (N14499, N14495, N3488, N11384, N210);
nand NAND3 (N14500, N14497, N7024, N2487);
or OR4 (N14501, N14473, N6047, N11366, N2896);
buf BUF1 (N14502, N14496);
nand NAND2 (N14503, N14491, N12808);
and AND3 (N14504, N14500, N4383, N4461);
not NOT1 (N14505, N14504);
xor XOR2 (N14506, N14498, N13842);
or OR4 (N14507, N14505, N14081, N8345, N13373);
nand NAND4 (N14508, N14489, N10858, N6236, N11881);
nor NOR3 (N14509, N14508, N10453, N6223);
xor XOR2 (N14510, N14494, N4400);
and AND3 (N14511, N14478, N12676, N421);
nor NOR3 (N14512, N14506, N1025, N10993);
xor XOR2 (N14513, N14499, N9339);
and AND2 (N14514, N14503, N13279);
buf BUF1 (N14515, N14513);
buf BUF1 (N14516, N14501);
buf BUF1 (N14517, N14510);
nand NAND4 (N14518, N14517, N9852, N10575, N10948);
xor XOR2 (N14519, N14493, N3666);
not NOT1 (N14520, N14507);
buf BUF1 (N14521, N14512);
not NOT1 (N14522, N14514);
buf BUF1 (N14523, N14520);
or OR2 (N14524, N14511, N6821);
not NOT1 (N14525, N14521);
not NOT1 (N14526, N14509);
or OR3 (N14527, N14524, N1565, N4344);
nand NAND3 (N14528, N14526, N3425, N9494);
nor NOR2 (N14529, N14525, N12325);
or OR4 (N14530, N14516, N8529, N9528, N3097);
and AND4 (N14531, N14502, N11216, N1899, N1709);
not NOT1 (N14532, N14523);
nand NAND4 (N14533, N14522, N4723, N5897, N944);
nand NAND4 (N14534, N14529, N7572, N9499, N876);
or OR3 (N14535, N14533, N7424, N3366);
xor XOR2 (N14536, N14534, N1467);
not NOT1 (N14537, N14515);
not NOT1 (N14538, N14530);
or OR4 (N14539, N14538, N9590, N1025, N11231);
or OR2 (N14540, N14531, N3733);
buf BUF1 (N14541, N14532);
or OR4 (N14542, N14535, N10460, N14188, N5112);
or OR2 (N14543, N14540, N6604);
and AND4 (N14544, N14518, N12478, N5412, N5257);
nor NOR4 (N14545, N14528, N3486, N10843, N1540);
buf BUF1 (N14546, N14539);
and AND4 (N14547, N14527, N835, N8640, N13003);
and AND4 (N14548, N14546, N5957, N11156, N2571);
and AND3 (N14549, N14542, N1261, N617);
or OR3 (N14550, N14537, N9295, N2668);
not NOT1 (N14551, N14545);
or OR3 (N14552, N14536, N8768, N2548);
nor NOR4 (N14553, N14543, N12097, N4760, N2963);
xor XOR2 (N14554, N14544, N873);
nor NOR2 (N14555, N14541, N5007);
nand NAND4 (N14556, N14551, N6376, N12501, N2697);
buf BUF1 (N14557, N14555);
buf BUF1 (N14558, N14548);
nand NAND4 (N14559, N14557, N10115, N7673, N11250);
buf BUF1 (N14560, N14559);
and AND2 (N14561, N14549, N13393);
nor NOR3 (N14562, N14552, N7033, N3410);
nor NOR3 (N14563, N14562, N13312, N7176);
and AND4 (N14564, N14553, N6780, N8044, N12682);
or OR3 (N14565, N14550, N5310, N2372);
nand NAND4 (N14566, N14554, N3819, N1064, N7405);
xor XOR2 (N14567, N14563, N10782);
not NOT1 (N14568, N14567);
nor NOR2 (N14569, N14547, N4244);
and AND2 (N14570, N14564, N9796);
and AND3 (N14571, N14519, N10318, N6140);
or OR2 (N14572, N14565, N13528);
nand NAND2 (N14573, N14566, N1365);
and AND4 (N14574, N14569, N1854, N2900, N12248);
not NOT1 (N14575, N14572);
not NOT1 (N14576, N14568);
buf BUF1 (N14577, N14575);
and AND4 (N14578, N14560, N8409, N420, N2794);
buf BUF1 (N14579, N14576);
not NOT1 (N14580, N14573);
nand NAND4 (N14581, N14574, N12469, N6517, N8310);
buf BUF1 (N14582, N14570);
nand NAND4 (N14583, N14558, N13768, N10589, N8018);
not NOT1 (N14584, N14571);
not NOT1 (N14585, N14577);
not NOT1 (N14586, N14582);
and AND4 (N14587, N14580, N5199, N6783, N11966);
not NOT1 (N14588, N14579);
not NOT1 (N14589, N14584);
buf BUF1 (N14590, N14587);
or OR4 (N14591, N14561, N2108, N3950, N11169);
buf BUF1 (N14592, N14578);
not NOT1 (N14593, N14589);
nor NOR4 (N14594, N14581, N7927, N260, N389);
nand NAND3 (N14595, N14590, N11718, N2350);
and AND2 (N14596, N14595, N6755);
xor XOR2 (N14597, N14594, N504);
not NOT1 (N14598, N14586);
nor NOR2 (N14599, N14597, N8963);
and AND3 (N14600, N14592, N6748, N2269);
or OR2 (N14601, N14600, N6538);
nand NAND4 (N14602, N14596, N2017, N3482, N2942);
or OR3 (N14603, N14585, N5475, N4579);
not NOT1 (N14604, N14602);
or OR4 (N14605, N14604, N2390, N3007, N3704);
buf BUF1 (N14606, N14588);
and AND3 (N14607, N14591, N11790, N2728);
xor XOR2 (N14608, N14601, N13918);
and AND3 (N14609, N14608, N4007, N9349);
and AND4 (N14610, N14607, N4384, N11797, N2700);
xor XOR2 (N14611, N14605, N9347);
and AND3 (N14612, N14593, N4307, N13752);
buf BUF1 (N14613, N14599);
xor XOR2 (N14614, N14612, N6439);
not NOT1 (N14615, N14610);
not NOT1 (N14616, N14556);
xor XOR2 (N14617, N14606, N1959);
not NOT1 (N14618, N14603);
or OR2 (N14619, N14583, N6626);
not NOT1 (N14620, N14615);
or OR4 (N14621, N14614, N6115, N365, N7014);
xor XOR2 (N14622, N14619, N6178);
and AND2 (N14623, N14616, N6238);
xor XOR2 (N14624, N14598, N415);
buf BUF1 (N14625, N14623);
and AND3 (N14626, N14624, N4222, N4304);
and AND4 (N14627, N14613, N5573, N121, N2683);
nand NAND2 (N14628, N14622, N14015);
buf BUF1 (N14629, N14626);
not NOT1 (N14630, N14625);
not NOT1 (N14631, N14611);
buf BUF1 (N14632, N14620);
nor NOR2 (N14633, N14627, N6455);
not NOT1 (N14634, N14617);
not NOT1 (N14635, N14629);
xor XOR2 (N14636, N14634, N113);
nand NAND4 (N14637, N14635, N520, N8884, N1883);
or OR4 (N14638, N14618, N5148, N9936, N5932);
nor NOR2 (N14639, N14628, N8894);
or OR4 (N14640, N14637, N2967, N5940, N2422);
nand NAND4 (N14641, N14632, N7040, N2181, N10846);
nand NAND3 (N14642, N14621, N574, N9850);
nand NAND4 (N14643, N14642, N8883, N11361, N13562);
and AND3 (N14644, N14639, N14243, N7000);
or OR4 (N14645, N14638, N10517, N4023, N7859);
nor NOR3 (N14646, N14636, N3126, N13970);
xor XOR2 (N14647, N14646, N12744);
xor XOR2 (N14648, N14630, N4541);
xor XOR2 (N14649, N14633, N13872);
xor XOR2 (N14650, N14609, N5195);
not NOT1 (N14651, N14641);
buf BUF1 (N14652, N14648);
buf BUF1 (N14653, N14644);
nor NOR2 (N14654, N14650, N5710);
or OR4 (N14655, N14645, N3237, N9682, N6218);
or OR2 (N14656, N14651, N12759);
nor NOR2 (N14657, N14640, N5685);
or OR3 (N14658, N14643, N4506, N11818);
and AND3 (N14659, N14654, N1565, N12690);
buf BUF1 (N14660, N14656);
buf BUF1 (N14661, N14631);
not NOT1 (N14662, N14660);
xor XOR2 (N14663, N14653, N2875);
xor XOR2 (N14664, N14657, N10963);
or OR3 (N14665, N14652, N8256, N8071);
not NOT1 (N14666, N14661);
not NOT1 (N14667, N14665);
xor XOR2 (N14668, N14655, N7441);
xor XOR2 (N14669, N14649, N11628);
not NOT1 (N14670, N14647);
and AND3 (N14671, N14669, N7879, N8338);
nand NAND3 (N14672, N14658, N14256, N11511);
buf BUF1 (N14673, N14663);
buf BUF1 (N14674, N14673);
nand NAND3 (N14675, N14659, N14028, N12659);
nor NOR3 (N14676, N14664, N7458, N11289);
buf BUF1 (N14677, N14670);
or OR2 (N14678, N14662, N7179);
or OR2 (N14679, N14667, N7012);
nor NOR4 (N14680, N14672, N11746, N473, N4828);
not NOT1 (N14681, N14676);
nand NAND4 (N14682, N14671, N54, N9635, N201);
not NOT1 (N14683, N14678);
xor XOR2 (N14684, N14666, N6302);
xor XOR2 (N14685, N14677, N12693);
or OR3 (N14686, N14675, N4286, N2427);
and AND2 (N14687, N14682, N7747);
not NOT1 (N14688, N14680);
nand NAND3 (N14689, N14681, N5773, N11535);
and AND2 (N14690, N14684, N4399);
or OR3 (N14691, N14679, N88, N2841);
nor NOR4 (N14692, N14683, N5845, N10652, N5069);
buf BUF1 (N14693, N14687);
nor NOR4 (N14694, N14693, N5830, N9345, N73);
nand NAND4 (N14695, N14692, N11864, N1151, N712);
nand NAND4 (N14696, N14694, N1396, N13213, N1227);
not NOT1 (N14697, N14691);
nor NOR3 (N14698, N14668, N12102, N1302);
nor NOR3 (N14699, N14688, N32, N9048);
not NOT1 (N14700, N14674);
xor XOR2 (N14701, N14696, N8198);
buf BUF1 (N14702, N14695);
xor XOR2 (N14703, N14686, N3204);
or OR4 (N14704, N14685, N7967, N1883, N4257);
buf BUF1 (N14705, N14703);
and AND4 (N14706, N14699, N9693, N91, N11602);
or OR3 (N14707, N14705, N1958, N13674);
and AND3 (N14708, N14707, N9456, N9110);
buf BUF1 (N14709, N14700);
and AND3 (N14710, N14697, N12624, N5706);
nor NOR2 (N14711, N14706, N6524);
nor NOR4 (N14712, N14689, N9335, N1415, N12503);
and AND4 (N14713, N14701, N6814, N11072, N14364);
buf BUF1 (N14714, N14708);
xor XOR2 (N14715, N14690, N4118);
buf BUF1 (N14716, N14713);
and AND2 (N14717, N14710, N9058);
buf BUF1 (N14718, N14704);
nor NOR2 (N14719, N14711, N1301);
buf BUF1 (N14720, N14709);
nor NOR2 (N14721, N14718, N5943);
buf BUF1 (N14722, N14714);
and AND3 (N14723, N14712, N13984, N3789);
xor XOR2 (N14724, N14721, N489);
nor NOR2 (N14725, N14702, N1026);
or OR4 (N14726, N14717, N9445, N8969, N766);
nor NOR3 (N14727, N14698, N12759, N12510);
nor NOR4 (N14728, N14715, N13964, N2811, N2445);
nand NAND2 (N14729, N14726, N7471);
or OR4 (N14730, N14719, N334, N12676, N401);
buf BUF1 (N14731, N14729);
xor XOR2 (N14732, N14725, N7171);
and AND2 (N14733, N14722, N11954);
nor NOR3 (N14734, N14732, N14486, N10989);
nor NOR2 (N14735, N14716, N8932);
nor NOR4 (N14736, N14728, N11636, N13628, N11278);
buf BUF1 (N14737, N14731);
nor NOR2 (N14738, N14737, N14559);
nand NAND2 (N14739, N14723, N5268);
and AND4 (N14740, N14724, N842, N10207, N8604);
buf BUF1 (N14741, N14740);
xor XOR2 (N14742, N14741, N7048);
buf BUF1 (N14743, N14730);
and AND3 (N14744, N14734, N11153, N7831);
xor XOR2 (N14745, N14743, N5178);
buf BUF1 (N14746, N14745);
nand NAND2 (N14747, N14744, N11364);
not NOT1 (N14748, N14727);
buf BUF1 (N14749, N14736);
nor NOR4 (N14750, N14738, N10637, N10835, N9169);
buf BUF1 (N14751, N14749);
and AND3 (N14752, N14733, N5818, N13338);
buf BUF1 (N14753, N14748);
xor XOR2 (N14754, N14746, N7567);
buf BUF1 (N14755, N14747);
buf BUF1 (N14756, N14735);
buf BUF1 (N14757, N14756);
xor XOR2 (N14758, N14757, N5141);
and AND2 (N14759, N14751, N13151);
nor NOR3 (N14760, N14739, N677, N8360);
or OR2 (N14761, N14752, N4253);
and AND3 (N14762, N14754, N12744, N2740);
nand NAND3 (N14763, N14720, N2178, N9887);
nor NOR4 (N14764, N14761, N13104, N3373, N1233);
xor XOR2 (N14765, N14763, N1460);
or OR3 (N14766, N14742, N14042, N6789);
nand NAND2 (N14767, N14758, N14194);
or OR4 (N14768, N14759, N12875, N4155, N12639);
nor NOR4 (N14769, N14765, N10664, N9390, N8751);
nand NAND2 (N14770, N14767, N544);
and AND3 (N14771, N14768, N14304, N12885);
xor XOR2 (N14772, N14762, N11432);
nand NAND2 (N14773, N14771, N13215);
xor XOR2 (N14774, N14769, N10849);
buf BUF1 (N14775, N14773);
nor NOR3 (N14776, N14750, N2597, N6325);
or OR2 (N14777, N14764, N300);
not NOT1 (N14778, N14776);
and AND2 (N14779, N14760, N5524);
xor XOR2 (N14780, N14766, N4246);
or OR2 (N14781, N14775, N13836);
not NOT1 (N14782, N14772);
buf BUF1 (N14783, N14753);
or OR4 (N14784, N14779, N8546, N8391, N4766);
nand NAND3 (N14785, N14783, N13702, N2311);
xor XOR2 (N14786, N14781, N9422);
nor NOR3 (N14787, N14774, N8317, N11075);
buf BUF1 (N14788, N14770);
nand NAND2 (N14789, N14780, N9876);
xor XOR2 (N14790, N14787, N11830);
nand NAND3 (N14791, N14755, N7734, N12523);
nor NOR3 (N14792, N14782, N1675, N1900);
not NOT1 (N14793, N14785);
or OR4 (N14794, N14784, N6751, N3578, N4911);
xor XOR2 (N14795, N14790, N8800);
xor XOR2 (N14796, N14794, N11409);
not NOT1 (N14797, N14777);
and AND4 (N14798, N14796, N10407, N4984, N6930);
nor NOR3 (N14799, N14791, N6577, N6546);
buf BUF1 (N14800, N14792);
not NOT1 (N14801, N14800);
and AND2 (N14802, N14798, N6071);
not NOT1 (N14803, N14788);
nand NAND3 (N14804, N14778, N5727, N4741);
nor NOR3 (N14805, N14789, N14685, N1122);
buf BUF1 (N14806, N14797);
nand NAND3 (N14807, N14806, N8344, N456);
not NOT1 (N14808, N14807);
buf BUF1 (N14809, N14799);
xor XOR2 (N14810, N14795, N5271);
nor NOR3 (N14811, N14802, N13524, N5692);
xor XOR2 (N14812, N14801, N454);
or OR4 (N14813, N14809, N7306, N10595, N7938);
nand NAND2 (N14814, N14811, N10236);
nor NOR4 (N14815, N14812, N8045, N8807, N10503);
xor XOR2 (N14816, N14805, N12275);
not NOT1 (N14817, N14786);
and AND2 (N14818, N14793, N7007);
and AND4 (N14819, N14818, N7129, N2529, N2573);
not NOT1 (N14820, N14816);
and AND4 (N14821, N14808, N6086, N11163, N5370);
buf BUF1 (N14822, N14817);
nand NAND4 (N14823, N14813, N9839, N12735, N4064);
nand NAND4 (N14824, N14804, N12072, N4370, N14136);
nand NAND4 (N14825, N14815, N3270, N9057, N6073);
nor NOR2 (N14826, N14803, N1492);
or OR2 (N14827, N14821, N1547);
nand NAND2 (N14828, N14825, N7378);
or OR3 (N14829, N14820, N12358, N1985);
nor NOR2 (N14830, N14824, N12537);
nand NAND2 (N14831, N14819, N6029);
not NOT1 (N14832, N14826);
xor XOR2 (N14833, N14829, N3528);
not NOT1 (N14834, N14814);
not NOT1 (N14835, N14810);
or OR3 (N14836, N14823, N6685, N13922);
buf BUF1 (N14837, N14836);
or OR3 (N14838, N14828, N6726, N8771);
and AND3 (N14839, N14822, N4797, N7580);
buf BUF1 (N14840, N14838);
nor NOR3 (N14841, N14833, N2153, N14140);
nand NAND2 (N14842, N14830, N6078);
and AND3 (N14843, N14839, N6843, N8797);
xor XOR2 (N14844, N14831, N14469);
or OR3 (N14845, N14827, N945, N13775);
buf BUF1 (N14846, N14835);
nor NOR2 (N14847, N14834, N5777);
xor XOR2 (N14848, N14843, N6629);
buf BUF1 (N14849, N14847);
nor NOR2 (N14850, N14837, N9800);
not NOT1 (N14851, N14832);
nor NOR3 (N14852, N14848, N4511, N13946);
and AND4 (N14853, N14846, N8150, N2526, N6460);
or OR4 (N14854, N14852, N8836, N10793, N4650);
and AND2 (N14855, N14853, N10322);
not NOT1 (N14856, N14844);
nor NOR3 (N14857, N14840, N2277, N3201);
buf BUF1 (N14858, N14854);
nor NOR3 (N14859, N14851, N14139, N8705);
nand NAND2 (N14860, N14858, N9186);
not NOT1 (N14861, N14841);
nor NOR4 (N14862, N14859, N2775, N2548, N6005);
nand NAND2 (N14863, N14857, N7824);
or OR3 (N14864, N14855, N6999, N3303);
nand NAND3 (N14865, N14863, N3, N8615);
or OR4 (N14866, N14845, N451, N1283, N14422);
not NOT1 (N14867, N14850);
nor NOR3 (N14868, N14842, N12212, N5155);
and AND4 (N14869, N14866, N12170, N3506, N1062);
and AND2 (N14870, N14864, N9796);
and AND4 (N14871, N14860, N11611, N13836, N3813);
nand NAND2 (N14872, N14868, N10854);
not NOT1 (N14873, N14861);
or OR4 (N14874, N14865, N9203, N10649, N13421);
or OR3 (N14875, N14871, N13973, N12586);
xor XOR2 (N14876, N14867, N12267);
nand NAND2 (N14877, N14874, N4578);
not NOT1 (N14878, N14873);
and AND2 (N14879, N14877, N8028);
not NOT1 (N14880, N14862);
and AND2 (N14881, N14870, N10797);
xor XOR2 (N14882, N14869, N10137);
and AND2 (N14883, N14880, N2909);
xor XOR2 (N14884, N14879, N4263);
nor NOR4 (N14885, N14884, N9943, N6569, N3928);
or OR4 (N14886, N14878, N7885, N1813, N2359);
not NOT1 (N14887, N14883);
or OR3 (N14888, N14886, N3633, N12857);
nand NAND2 (N14889, N14888, N9034);
not NOT1 (N14890, N14887);
not NOT1 (N14891, N14882);
nand NAND2 (N14892, N14881, N2710);
not NOT1 (N14893, N14856);
nand NAND2 (N14894, N14875, N11888);
xor XOR2 (N14895, N14876, N11115);
or OR4 (N14896, N14893, N10537, N7350, N2164);
or OR2 (N14897, N14872, N2196);
and AND2 (N14898, N14895, N5360);
not NOT1 (N14899, N14898);
and AND3 (N14900, N14892, N4156, N3727);
nand NAND3 (N14901, N14891, N4516, N10656);
or OR2 (N14902, N14894, N1412);
not NOT1 (N14903, N14896);
or OR4 (N14904, N14885, N14644, N9870, N6764);
or OR4 (N14905, N14899, N3373, N2906, N121);
not NOT1 (N14906, N14897);
and AND3 (N14907, N14902, N13999, N13293);
or OR2 (N14908, N14907, N14550);
not NOT1 (N14909, N14890);
nor NOR2 (N14910, N14903, N6587);
buf BUF1 (N14911, N14901);
nor NOR2 (N14912, N14911, N13591);
or OR2 (N14913, N14904, N2058);
xor XOR2 (N14914, N14905, N9215);
xor XOR2 (N14915, N14909, N4909);
xor XOR2 (N14916, N14914, N12795);
buf BUF1 (N14917, N14906);
nor NOR3 (N14918, N14910, N14723, N4117);
xor XOR2 (N14919, N14889, N10876);
and AND4 (N14920, N14913, N12304, N9750, N7529);
or OR2 (N14921, N14916, N3019);
buf BUF1 (N14922, N14849);
nor NOR4 (N14923, N14919, N10478, N4834, N1737);
or OR4 (N14924, N14920, N542, N13283, N8736);
and AND3 (N14925, N14908, N12369, N5844);
xor XOR2 (N14926, N14918, N1984);
nor NOR3 (N14927, N14917, N4902, N6121);
xor XOR2 (N14928, N14926, N12572);
nand NAND2 (N14929, N14928, N7051);
or OR2 (N14930, N14925, N14112);
nand NAND3 (N14931, N14924, N10517, N7141);
nand NAND4 (N14932, N14929, N6314, N6796, N12507);
and AND3 (N14933, N14900, N10016, N5357);
nand NAND2 (N14934, N14923, N3914);
not NOT1 (N14935, N14912);
nor NOR3 (N14936, N14932, N2787, N155);
xor XOR2 (N14937, N14936, N12341);
nor NOR2 (N14938, N14931, N4419);
not NOT1 (N14939, N14930);
nor NOR2 (N14940, N14934, N5657);
and AND4 (N14941, N14927, N6797, N12924, N7376);
nor NOR2 (N14942, N14921, N8087);
nand NAND4 (N14943, N14937, N524, N1885, N2537);
and AND3 (N14944, N14942, N8634, N6838);
or OR2 (N14945, N14915, N12033);
nor NOR4 (N14946, N14938, N11207, N1699, N6589);
buf BUF1 (N14947, N14922);
nand NAND3 (N14948, N14944, N1332, N988);
xor XOR2 (N14949, N14933, N182);
not NOT1 (N14950, N14948);
nand NAND2 (N14951, N14949, N14540);
and AND4 (N14952, N14935, N5093, N6642, N5551);
not NOT1 (N14953, N14941);
buf BUF1 (N14954, N14950);
xor XOR2 (N14955, N14940, N10828);
and AND4 (N14956, N14946, N6480, N5182, N2641);
or OR4 (N14957, N14956, N13539, N11390, N9026);
and AND2 (N14958, N14952, N13301);
buf BUF1 (N14959, N14945);
xor XOR2 (N14960, N14939, N14900);
not NOT1 (N14961, N14958);
or OR2 (N14962, N14955, N7639);
and AND2 (N14963, N14957, N14560);
xor XOR2 (N14964, N14943, N14936);
buf BUF1 (N14965, N14962);
buf BUF1 (N14966, N14951);
buf BUF1 (N14967, N14960);
not NOT1 (N14968, N14954);
not NOT1 (N14969, N14964);
not NOT1 (N14970, N14965);
xor XOR2 (N14971, N14969, N7155);
nor NOR4 (N14972, N14970, N11520, N6078, N4903);
nor NOR4 (N14973, N14963, N7777, N206, N6860);
buf BUF1 (N14974, N14961);
xor XOR2 (N14975, N14973, N933);
not NOT1 (N14976, N14974);
and AND4 (N14977, N14947, N1665, N8266, N3155);
nor NOR2 (N14978, N14971, N7511);
buf BUF1 (N14979, N14976);
or OR4 (N14980, N14979, N5192, N14819, N8725);
nor NOR4 (N14981, N14967, N13886, N8789, N6885);
nand NAND3 (N14982, N14977, N5758, N3274);
nor NOR2 (N14983, N14982, N1569);
nor NOR2 (N14984, N14968, N1597);
nor NOR3 (N14985, N14953, N6468, N10645);
nor NOR3 (N14986, N14981, N2281, N11690);
nand NAND2 (N14987, N14959, N7947);
nand NAND3 (N14988, N14984, N5167, N2619);
nor NOR3 (N14989, N14978, N7220, N7676);
xor XOR2 (N14990, N14988, N12627);
xor XOR2 (N14991, N14983, N13983);
nor NOR4 (N14992, N14991, N8133, N4390, N5007);
nand NAND2 (N14993, N14987, N7913);
buf BUF1 (N14994, N14990);
and AND3 (N14995, N14992, N4919, N277);
not NOT1 (N14996, N14994);
and AND4 (N14997, N14986, N7271, N8293, N9138);
nand NAND2 (N14998, N14985, N10211);
nand NAND3 (N14999, N14966, N4396, N5864);
buf BUF1 (N15000, N14989);
and AND4 (N15001, N14972, N13498, N9111, N4972);
or OR2 (N15002, N14975, N13659);
nand NAND3 (N15003, N15000, N7686, N629);
or OR2 (N15004, N15003, N10536);
or OR4 (N15005, N15001, N7658, N3549, N11582);
buf BUF1 (N15006, N14999);
or OR4 (N15007, N14998, N8683, N3366, N14128);
not NOT1 (N15008, N14995);
buf BUF1 (N15009, N14993);
buf BUF1 (N15010, N14980);
buf BUF1 (N15011, N15009);
and AND2 (N15012, N15008, N6006);
nand NAND2 (N15013, N15010, N13071);
nand NAND2 (N15014, N15006, N7937);
and AND3 (N15015, N15014, N2990, N8729);
nor NOR3 (N15016, N15002, N154, N12702);
or OR2 (N15017, N14997, N10141);
nor NOR2 (N15018, N15011, N1269);
nand NAND2 (N15019, N14996, N453);
buf BUF1 (N15020, N15015);
and AND2 (N15021, N15013, N5732);
or OR3 (N15022, N15020, N8401, N6897);
not NOT1 (N15023, N15021);
not NOT1 (N15024, N15017);
nand NAND3 (N15025, N15023, N2620, N1995);
or OR2 (N15026, N15019, N11418);
xor XOR2 (N15027, N15016, N10260);
nand NAND3 (N15028, N15018, N9969, N12696);
and AND4 (N15029, N15028, N7153, N2111, N8957);
and AND2 (N15030, N15027, N3463);
and AND4 (N15031, N15022, N11387, N8651, N2311);
buf BUF1 (N15032, N15024);
nand NAND4 (N15033, N15026, N8513, N1867, N10476);
buf BUF1 (N15034, N15005);
or OR4 (N15035, N15030, N1048, N4191, N10908);
nor NOR2 (N15036, N15025, N2264);
nor NOR4 (N15037, N15033, N14725, N4476, N9423);
or OR3 (N15038, N15037, N3305, N12114);
xor XOR2 (N15039, N15007, N13635);
xor XOR2 (N15040, N15036, N7708);
nor NOR2 (N15041, N15034, N9149);
nor NOR4 (N15042, N15035, N10088, N12988, N9770);
nor NOR2 (N15043, N15032, N9383);
or OR3 (N15044, N15038, N11185, N8516);
buf BUF1 (N15045, N15012);
buf BUF1 (N15046, N15045);
and AND4 (N15047, N15004, N4041, N7402, N8075);
buf BUF1 (N15048, N15040);
nand NAND4 (N15049, N15047, N8132, N8364, N1994);
not NOT1 (N15050, N15049);
not NOT1 (N15051, N15048);
buf BUF1 (N15052, N15046);
buf BUF1 (N15053, N15031);
xor XOR2 (N15054, N15051, N11096);
nand NAND2 (N15055, N15044, N14159);
and AND2 (N15056, N15050, N6160);
buf BUF1 (N15057, N15052);
xor XOR2 (N15058, N15055, N6745);
nand NAND4 (N15059, N15043, N14158, N14206, N12419);
nor NOR3 (N15060, N15056, N6372, N13345);
and AND2 (N15061, N15057, N10760);
and AND4 (N15062, N15041, N7505, N11640, N14455);
nand NAND4 (N15063, N15039, N13080, N3610, N3560);
or OR2 (N15064, N15058, N684);
nor NOR2 (N15065, N15062, N3814);
nand NAND2 (N15066, N15061, N1758);
nand NAND2 (N15067, N15029, N7705);
or OR3 (N15068, N15063, N8959, N2740);
nor NOR4 (N15069, N15059, N13505, N8772, N9068);
buf BUF1 (N15070, N15068);
or OR2 (N15071, N15053, N5842);
nor NOR3 (N15072, N15070, N833, N5944);
not NOT1 (N15073, N15066);
not NOT1 (N15074, N15067);
not NOT1 (N15075, N15060);
and AND2 (N15076, N15065, N1427);
and AND3 (N15077, N15073, N9691, N9048);
buf BUF1 (N15078, N15074);
nor NOR2 (N15079, N15075, N6340);
xor XOR2 (N15080, N15054, N6298);
xor XOR2 (N15081, N15069, N13536);
not NOT1 (N15082, N15042);
and AND4 (N15083, N15064, N1611, N3848, N13562);
or OR3 (N15084, N15079, N3268, N6507);
nor NOR4 (N15085, N15082, N13215, N7723, N14597);
or OR3 (N15086, N15081, N8527, N135);
xor XOR2 (N15087, N15071, N8819);
not NOT1 (N15088, N15078);
not NOT1 (N15089, N15083);
buf BUF1 (N15090, N15086);
and AND2 (N15091, N15084, N9363);
not NOT1 (N15092, N15077);
and AND3 (N15093, N15090, N8402, N8837);
nand NAND4 (N15094, N15072, N997, N2059, N10345);
nand NAND2 (N15095, N15085, N4856);
xor XOR2 (N15096, N15080, N2302);
not NOT1 (N15097, N15092);
nor NOR3 (N15098, N15087, N7997, N8070);
xor XOR2 (N15099, N15091, N2774);
nand NAND2 (N15100, N15096, N6952);
and AND2 (N15101, N15098, N12364);
nand NAND4 (N15102, N15089, N202, N3428, N8602);
nor NOR4 (N15103, N15076, N5920, N10514, N8287);
nand NAND4 (N15104, N15095, N9473, N7044, N14491);
and AND4 (N15105, N15104, N9993, N11022, N3163);
buf BUF1 (N15106, N15088);
not NOT1 (N15107, N15099);
not NOT1 (N15108, N15105);
nand NAND3 (N15109, N15106, N13986, N13696);
not NOT1 (N15110, N15102);
xor XOR2 (N15111, N15110, N1485);
xor XOR2 (N15112, N15097, N3208);
or OR4 (N15113, N15108, N7300, N14028, N8858);
not NOT1 (N15114, N15100);
or OR4 (N15115, N15109, N998, N402, N3276);
not NOT1 (N15116, N15107);
not NOT1 (N15117, N15113);
or OR2 (N15118, N15114, N1290);
buf BUF1 (N15119, N15103);
and AND3 (N15120, N15119, N11642, N11293);
or OR4 (N15121, N15117, N890, N13666, N9926);
xor XOR2 (N15122, N15121, N2886);
nor NOR3 (N15123, N15112, N10008, N3198);
nor NOR2 (N15124, N15094, N6480);
nand NAND4 (N15125, N15101, N12928, N3223, N2642);
buf BUF1 (N15126, N15123);
or OR3 (N15127, N15122, N4775, N7844);
buf BUF1 (N15128, N15127);
xor XOR2 (N15129, N15126, N6330);
buf BUF1 (N15130, N15129);
not NOT1 (N15131, N15124);
or OR4 (N15132, N15128, N4071, N2454, N10203);
nand NAND2 (N15133, N15132, N6752);
or OR3 (N15134, N15093, N12886, N9374);
xor XOR2 (N15135, N15125, N4164);
xor XOR2 (N15136, N15135, N3217);
and AND4 (N15137, N15130, N12934, N1061, N9329);
nor NOR3 (N15138, N15133, N1682, N11076);
nand NAND4 (N15139, N15131, N525, N9855, N850);
or OR4 (N15140, N15115, N6777, N1978, N11367);
and AND4 (N15141, N15118, N235, N9694, N8534);
buf BUF1 (N15142, N15137);
not NOT1 (N15143, N15140);
xor XOR2 (N15144, N15142, N5027);
or OR2 (N15145, N15134, N11665);
xor XOR2 (N15146, N15139, N12146);
not NOT1 (N15147, N15144);
xor XOR2 (N15148, N15111, N3246);
not NOT1 (N15149, N15138);
and AND4 (N15150, N15143, N15022, N5976, N13366);
not NOT1 (N15151, N15141);
not NOT1 (N15152, N15150);
xor XOR2 (N15153, N15152, N4750);
and AND4 (N15154, N15145, N117, N14990, N13908);
buf BUF1 (N15155, N15147);
xor XOR2 (N15156, N15116, N501);
nand NAND2 (N15157, N15148, N12076);
not NOT1 (N15158, N15153);
not NOT1 (N15159, N15136);
nand NAND2 (N15160, N15158, N12249);
nand NAND3 (N15161, N15159, N1492, N6645);
or OR4 (N15162, N15156, N3971, N6681, N5405);
or OR4 (N15163, N15120, N14903, N4770, N1864);
nor NOR3 (N15164, N15149, N5806, N8679);
and AND4 (N15165, N15154, N4786, N11714, N70);
not NOT1 (N15166, N15160);
nand NAND4 (N15167, N15162, N3592, N12904, N2842);
nor NOR2 (N15168, N15151, N1576);
nand NAND4 (N15169, N15164, N8974, N5256, N11556);
nand NAND4 (N15170, N15157, N3858, N10609, N1822);
nor NOR3 (N15171, N15146, N4665, N12040);
buf BUF1 (N15172, N15169);
not NOT1 (N15173, N15168);
not NOT1 (N15174, N15171);
xor XOR2 (N15175, N15166, N14132);
and AND4 (N15176, N15170, N5111, N10307, N516);
and AND2 (N15177, N15173, N7020);
xor XOR2 (N15178, N15161, N13924);
not NOT1 (N15179, N15155);
or OR4 (N15180, N15175, N9502, N10059, N2811);
nor NOR4 (N15181, N15172, N9606, N2841, N2140);
nor NOR4 (N15182, N15165, N11855, N4073, N12235);
and AND2 (N15183, N15177, N2028);
buf BUF1 (N15184, N15167);
nand NAND4 (N15185, N15180, N9510, N11127, N946);
or OR4 (N15186, N15179, N10366, N3269, N14871);
nor NOR2 (N15187, N15174, N13979);
not NOT1 (N15188, N15178);
and AND2 (N15189, N15187, N1924);
xor XOR2 (N15190, N15181, N6469);
not NOT1 (N15191, N15182);
nor NOR4 (N15192, N15176, N5106, N1186, N1262);
nor NOR3 (N15193, N15192, N203, N14715);
and AND3 (N15194, N15183, N8218, N324);
xor XOR2 (N15195, N15186, N15143);
nor NOR4 (N15196, N15193, N5299, N2515, N2406);
and AND4 (N15197, N15189, N14114, N455, N14026);
or OR2 (N15198, N15190, N12656);
nor NOR4 (N15199, N15184, N5895, N9931, N7904);
and AND2 (N15200, N15188, N1051);
not NOT1 (N15201, N15191);
not NOT1 (N15202, N15185);
buf BUF1 (N15203, N15197);
xor XOR2 (N15204, N15199, N936);
not NOT1 (N15205, N15201);
or OR3 (N15206, N15195, N8058, N8707);
nor NOR3 (N15207, N15203, N13447, N1457);
or OR3 (N15208, N15202, N5366, N2127);
or OR3 (N15209, N15206, N11655, N7848);
buf BUF1 (N15210, N15200);
buf BUF1 (N15211, N15205);
not NOT1 (N15212, N15204);
not NOT1 (N15213, N15208);
xor XOR2 (N15214, N15210, N6617);
buf BUF1 (N15215, N15163);
not NOT1 (N15216, N15207);
or OR4 (N15217, N15216, N10571, N6973, N5499);
not NOT1 (N15218, N15215);
not NOT1 (N15219, N15209);
buf BUF1 (N15220, N15217);
or OR2 (N15221, N15220, N6016);
nor NOR2 (N15222, N15212, N10653);
or OR2 (N15223, N15198, N4542);
xor XOR2 (N15224, N15222, N2617);
nand NAND2 (N15225, N15221, N11050);
and AND4 (N15226, N15225, N2481, N7612, N1304);
buf BUF1 (N15227, N15219);
nor NOR3 (N15228, N15211, N9028, N1939);
nand NAND2 (N15229, N15214, N6378);
not NOT1 (N15230, N15213);
or OR2 (N15231, N15230, N2583);
nor NOR3 (N15232, N15231, N13383, N2403);
nand NAND2 (N15233, N15218, N4856);
xor XOR2 (N15234, N15226, N4960);
nor NOR2 (N15235, N15232, N11845);
or OR2 (N15236, N15223, N5896);
nand NAND4 (N15237, N15229, N13243, N11643, N13075);
buf BUF1 (N15238, N15233);
xor XOR2 (N15239, N15238, N10852);
buf BUF1 (N15240, N15196);
nand NAND2 (N15241, N15227, N12478);
not NOT1 (N15242, N15234);
or OR3 (N15243, N15235, N12725, N4234);
buf BUF1 (N15244, N15236);
or OR3 (N15245, N15244, N1601, N9589);
buf BUF1 (N15246, N15194);
or OR3 (N15247, N15239, N11564, N3674);
xor XOR2 (N15248, N15241, N11753);
nand NAND4 (N15249, N15228, N38, N527, N2759);
nand NAND3 (N15250, N15237, N1660, N9190);
or OR4 (N15251, N15242, N5572, N12075, N3457);
and AND4 (N15252, N15250, N179, N14328, N4259);
or OR3 (N15253, N15247, N8037, N7673);
or OR4 (N15254, N15243, N7959, N12356, N9164);
or OR2 (N15255, N15248, N12795);
nor NOR3 (N15256, N15255, N2294, N11307);
nand NAND3 (N15257, N15254, N7754, N14000);
not NOT1 (N15258, N15245);
nor NOR2 (N15259, N15256, N12069);
buf BUF1 (N15260, N15240);
buf BUF1 (N15261, N15253);
not NOT1 (N15262, N15246);
not NOT1 (N15263, N15224);
nor NOR2 (N15264, N15261, N12589);
nor NOR3 (N15265, N15262, N2523, N438);
nor NOR2 (N15266, N15259, N334);
and AND2 (N15267, N15260, N1950);
buf BUF1 (N15268, N15258);
not NOT1 (N15269, N15268);
nor NOR2 (N15270, N15249, N11284);
not NOT1 (N15271, N15263);
or OR2 (N15272, N15271, N10275);
not NOT1 (N15273, N15266);
and AND3 (N15274, N15265, N5511, N6879);
buf BUF1 (N15275, N15251);
nand NAND4 (N15276, N15267, N5488, N964, N8879);
and AND2 (N15277, N15275, N14180);
or OR2 (N15278, N15273, N3617);
not NOT1 (N15279, N15264);
not NOT1 (N15280, N15272);
and AND2 (N15281, N15274, N6207);
or OR3 (N15282, N15280, N14141, N11262);
nor NOR4 (N15283, N15281, N4976, N10194, N12513);
xor XOR2 (N15284, N15276, N6958);
xor XOR2 (N15285, N15252, N10215);
nand NAND3 (N15286, N15282, N11233, N10571);
not NOT1 (N15287, N15277);
and AND3 (N15288, N15283, N9331, N5437);
nand NAND3 (N15289, N15269, N5234, N4477);
and AND4 (N15290, N15284, N12554, N1860, N12383);
not NOT1 (N15291, N15289);
nand NAND2 (N15292, N15270, N6323);
xor XOR2 (N15293, N15290, N12537);
nor NOR3 (N15294, N15293, N2402, N2717);
not NOT1 (N15295, N15292);
and AND2 (N15296, N15295, N11246);
xor XOR2 (N15297, N15285, N7537);
not NOT1 (N15298, N15279);
nand NAND2 (N15299, N15294, N8095);
buf BUF1 (N15300, N15296);
nor NOR3 (N15301, N15298, N2765, N10545);
nand NAND4 (N15302, N15278, N6823, N12650, N15281);
not NOT1 (N15303, N15301);
nand NAND4 (N15304, N15286, N12656, N12209, N6066);
xor XOR2 (N15305, N15300, N13533);
not NOT1 (N15306, N15291);
or OR4 (N15307, N15305, N8167, N13130, N5309);
or OR4 (N15308, N15303, N3874, N14099, N1568);
or OR3 (N15309, N15299, N804, N8125);
not NOT1 (N15310, N15257);
buf BUF1 (N15311, N15297);
or OR2 (N15312, N15304, N11113);
nand NAND4 (N15313, N15308, N7999, N2704, N2899);
nand NAND3 (N15314, N15312, N14549, N9158);
xor XOR2 (N15315, N15288, N8207);
nor NOR3 (N15316, N15313, N7212, N3751);
buf BUF1 (N15317, N15315);
not NOT1 (N15318, N15311);
or OR4 (N15319, N15316, N9755, N2004, N663);
xor XOR2 (N15320, N15310, N8972);
nor NOR2 (N15321, N15307, N4250);
and AND2 (N15322, N15302, N13691);
xor XOR2 (N15323, N15322, N10082);
buf BUF1 (N15324, N15287);
buf BUF1 (N15325, N15314);
not NOT1 (N15326, N15325);
or OR2 (N15327, N15319, N1307);
or OR4 (N15328, N15318, N2015, N14940, N4983);
or OR3 (N15329, N15321, N2290, N12692);
xor XOR2 (N15330, N15317, N7172);
nand NAND4 (N15331, N15326, N4524, N1755, N4536);
buf BUF1 (N15332, N15329);
and AND2 (N15333, N15328, N14298);
not NOT1 (N15334, N15306);
not NOT1 (N15335, N15309);
or OR4 (N15336, N15324, N7577, N14495, N4844);
buf BUF1 (N15337, N15331);
and AND3 (N15338, N15333, N9344, N1674);
nand NAND2 (N15339, N15337, N8482);
nand NAND3 (N15340, N15336, N3087, N3798);
and AND2 (N15341, N15334, N3838);
buf BUF1 (N15342, N15320);
or OR3 (N15343, N15323, N11197, N7653);
nor NOR2 (N15344, N15338, N14367);
nor NOR4 (N15345, N15330, N7849, N12915, N4862);
buf BUF1 (N15346, N15335);
xor XOR2 (N15347, N15341, N12914);
buf BUF1 (N15348, N15332);
not NOT1 (N15349, N15327);
or OR3 (N15350, N15348, N5615, N14511);
xor XOR2 (N15351, N15346, N11513);
nand NAND2 (N15352, N15351, N447);
nand NAND2 (N15353, N15350, N8248);
and AND3 (N15354, N15342, N2214, N5728);
and AND2 (N15355, N15353, N1938);
nor NOR2 (N15356, N15340, N9106);
or OR4 (N15357, N15356, N11284, N10017, N8371);
nor NOR2 (N15358, N15344, N7121);
nand NAND4 (N15359, N15339, N4751, N10039, N10172);
or OR3 (N15360, N15345, N4472, N14588);
buf BUF1 (N15361, N15360);
nor NOR2 (N15362, N15349, N1649);
not NOT1 (N15363, N15355);
and AND4 (N15364, N15343, N12434, N6346, N1026);
buf BUF1 (N15365, N15361);
not NOT1 (N15366, N15352);
nor NOR4 (N15367, N15363, N15105, N3292, N1917);
nor NOR3 (N15368, N15358, N9147, N12546);
buf BUF1 (N15369, N15366);
xor XOR2 (N15370, N15365, N12371);
or OR3 (N15371, N15369, N2745, N4226);
nand NAND2 (N15372, N15368, N4048);
or OR3 (N15373, N15362, N11369, N1713);
not NOT1 (N15374, N15372);
and AND4 (N15375, N15370, N4008, N10243, N6539);
or OR4 (N15376, N15367, N1030, N10696, N580);
nor NOR2 (N15377, N15375, N4456);
nand NAND2 (N15378, N15374, N3779);
buf BUF1 (N15379, N15347);
nor NOR4 (N15380, N15371, N4623, N3915, N12797);
buf BUF1 (N15381, N15359);
or OR4 (N15382, N15379, N3784, N14539, N5145);
nor NOR4 (N15383, N15354, N5449, N10192, N7319);
or OR4 (N15384, N15377, N2541, N8993, N9031);
nor NOR3 (N15385, N15382, N6555, N10704);
nand NAND4 (N15386, N15376, N5650, N6306, N7874);
buf BUF1 (N15387, N15383);
buf BUF1 (N15388, N15378);
and AND2 (N15389, N15385, N2653);
nand NAND4 (N15390, N15384, N15092, N10917, N8343);
xor XOR2 (N15391, N15387, N8625);
nand NAND3 (N15392, N15357, N14615, N6276);
or OR2 (N15393, N15381, N9856);
xor XOR2 (N15394, N15393, N4110);
not NOT1 (N15395, N15394);
not NOT1 (N15396, N15390);
not NOT1 (N15397, N15392);
nand NAND3 (N15398, N15373, N15252, N3471);
not NOT1 (N15399, N15398);
nor NOR4 (N15400, N15364, N3923, N9630, N6047);
nand NAND2 (N15401, N15395, N10758);
nor NOR4 (N15402, N15391, N1002, N10431, N12797);
or OR2 (N15403, N15397, N3202);
or OR3 (N15404, N15386, N12198, N3153);
nor NOR2 (N15405, N15403, N8039);
xor XOR2 (N15406, N15389, N9524);
buf BUF1 (N15407, N15401);
not NOT1 (N15408, N15406);
nand NAND2 (N15409, N15399, N14416);
nor NOR2 (N15410, N15402, N4459);
buf BUF1 (N15411, N15388);
or OR4 (N15412, N15405, N10112, N566, N8235);
not NOT1 (N15413, N15380);
or OR3 (N15414, N15396, N6728, N8061);
or OR3 (N15415, N15408, N3699, N9481);
not NOT1 (N15416, N15410);
nand NAND3 (N15417, N15415, N9007, N14474);
xor XOR2 (N15418, N15413, N333);
and AND2 (N15419, N15412, N14771);
nor NOR2 (N15420, N15411, N4727);
xor XOR2 (N15421, N15417, N3908);
not NOT1 (N15422, N15421);
nand NAND2 (N15423, N15422, N9802);
buf BUF1 (N15424, N15416);
nor NOR2 (N15425, N15424, N4347);
nand NAND3 (N15426, N15420, N14649, N15165);
and AND3 (N15427, N15400, N12959, N11230);
buf BUF1 (N15428, N15426);
buf BUF1 (N15429, N15414);
nand NAND3 (N15430, N15418, N9121, N6062);
and AND3 (N15431, N15409, N2809, N8302);
or OR4 (N15432, N15431, N12194, N4023, N6620);
nor NOR2 (N15433, N15430, N8369);
xor XOR2 (N15434, N15419, N117);
nor NOR2 (N15435, N15404, N765);
not NOT1 (N15436, N15425);
and AND2 (N15437, N15435, N782);
or OR4 (N15438, N15428, N12404, N7057, N8478);
and AND3 (N15439, N15433, N12710, N8497);
not NOT1 (N15440, N15438);
or OR4 (N15441, N15439, N9422, N10888, N7650);
and AND3 (N15442, N15441, N11701, N11286);
nand NAND4 (N15443, N15434, N13207, N12438, N4952);
nor NOR4 (N15444, N15442, N686, N5393, N10945);
nand NAND4 (N15445, N15443, N12488, N4833, N6193);
or OR4 (N15446, N15432, N13624, N14089, N11971);
nand NAND4 (N15447, N15423, N10682, N8637, N15094);
not NOT1 (N15448, N15437);
or OR2 (N15449, N15440, N7104);
and AND2 (N15450, N15444, N14881);
xor XOR2 (N15451, N15449, N4646);
or OR4 (N15452, N15427, N11080, N4724, N1819);
or OR2 (N15453, N15407, N630);
and AND3 (N15454, N15450, N14081, N13900);
and AND4 (N15455, N15436, N1867, N13623, N4509);
or OR2 (N15456, N15445, N13520);
nor NOR3 (N15457, N15453, N11492, N1310);
xor XOR2 (N15458, N15446, N13029);
xor XOR2 (N15459, N15429, N9369);
or OR4 (N15460, N15452, N13155, N14801, N9968);
and AND2 (N15461, N15459, N12840);
and AND2 (N15462, N15447, N114);
buf BUF1 (N15463, N15460);
buf BUF1 (N15464, N15456);
not NOT1 (N15465, N15462);
xor XOR2 (N15466, N15463, N15234);
nor NOR4 (N15467, N15461, N9069, N12576, N4568);
buf BUF1 (N15468, N15458);
nand NAND2 (N15469, N15455, N6);
or OR2 (N15470, N15466, N5414);
nor NOR4 (N15471, N15451, N14299, N1579, N12374);
nand NAND2 (N15472, N15465, N4958);
or OR2 (N15473, N15467, N6904);
or OR3 (N15474, N15464, N3078, N12917);
nand NAND2 (N15475, N15457, N12415);
nand NAND2 (N15476, N15471, N14854);
not NOT1 (N15477, N15474);
nand NAND3 (N15478, N15472, N14878, N10910);
and AND4 (N15479, N15448, N5246, N15230, N1799);
buf BUF1 (N15480, N15475);
buf BUF1 (N15481, N15470);
buf BUF1 (N15482, N15478);
nor NOR2 (N15483, N15477, N10759);
or OR4 (N15484, N15473, N11269, N11236, N6070);
nor NOR2 (N15485, N15483, N3245);
nor NOR2 (N15486, N15469, N9273);
buf BUF1 (N15487, N15482);
nor NOR4 (N15488, N15485, N2907, N12550, N7881);
not NOT1 (N15489, N15487);
nand NAND4 (N15490, N15484, N10386, N10309, N12289);
xor XOR2 (N15491, N15490, N442);
not NOT1 (N15492, N15468);
xor XOR2 (N15493, N15486, N3513);
or OR2 (N15494, N15481, N9012);
buf BUF1 (N15495, N15480);
and AND4 (N15496, N15479, N5773, N15145, N41);
not NOT1 (N15497, N15489);
buf BUF1 (N15498, N15491);
nand NAND4 (N15499, N15454, N5710, N12806, N15008);
nand NAND3 (N15500, N15493, N6153, N9577);
nand NAND3 (N15501, N15476, N10684, N13611);
buf BUF1 (N15502, N15488);
nor NOR3 (N15503, N15495, N4870, N4422);
or OR2 (N15504, N15500, N6475);
not NOT1 (N15505, N15503);
and AND3 (N15506, N15492, N8581, N12599);
nand NAND2 (N15507, N15504, N11920);
or OR3 (N15508, N15494, N6778, N7145);
xor XOR2 (N15509, N15507, N10023);
or OR2 (N15510, N15499, N14031);
or OR3 (N15511, N15506, N12251, N8359);
or OR2 (N15512, N15496, N6003);
nand NAND4 (N15513, N15501, N3335, N1163, N11824);
not NOT1 (N15514, N15508);
or OR2 (N15515, N15511, N3897);
and AND2 (N15516, N15512, N5158);
or OR3 (N15517, N15514, N4728, N7952);
xor XOR2 (N15518, N15513, N10469);
nand NAND3 (N15519, N15498, N9222, N4395);
and AND4 (N15520, N15518, N11864, N1701, N9047);
or OR4 (N15521, N15516, N9457, N9306, N6466);
or OR4 (N15522, N15519, N7716, N7344, N13635);
buf BUF1 (N15523, N15521);
and AND2 (N15524, N15509, N13959);
and AND2 (N15525, N15497, N1754);
nor NOR4 (N15526, N15523, N12633, N2350, N14127);
nand NAND4 (N15527, N15520, N1350, N12434, N13997);
xor XOR2 (N15528, N15527, N9081);
and AND4 (N15529, N15526, N4794, N15060, N14109);
buf BUF1 (N15530, N15529);
not NOT1 (N15531, N15515);
nor NOR3 (N15532, N15510, N1980, N6708);
nor NOR2 (N15533, N15532, N1406);
and AND3 (N15534, N15525, N6767, N14642);
buf BUF1 (N15535, N15528);
and AND4 (N15536, N15502, N13106, N10352, N5169);
or OR4 (N15537, N15522, N548, N8279, N11192);
buf BUF1 (N15538, N15533);
and AND4 (N15539, N15534, N12118, N2128, N4188);
xor XOR2 (N15540, N15535, N3493);
buf BUF1 (N15541, N15517);
and AND4 (N15542, N15531, N3821, N10279, N14641);
or OR2 (N15543, N15540, N6835);
nor NOR2 (N15544, N15542, N8313);
not NOT1 (N15545, N15543);
nand NAND4 (N15546, N15538, N2524, N11859, N2739);
nand NAND3 (N15547, N15505, N8666, N11654);
not NOT1 (N15548, N15539);
nor NOR3 (N15549, N15536, N4601, N5390);
xor XOR2 (N15550, N15547, N6231);
buf BUF1 (N15551, N15544);
not NOT1 (N15552, N15546);
nor NOR2 (N15553, N15530, N14285);
nand NAND3 (N15554, N15553, N3557, N669);
xor XOR2 (N15555, N15537, N1206);
buf BUF1 (N15556, N15545);
nand NAND3 (N15557, N15524, N9990, N1513);
nor NOR2 (N15558, N15552, N5531);
nand NAND2 (N15559, N15555, N8176);
nor NOR2 (N15560, N15551, N5467);
nor NOR3 (N15561, N15549, N10874, N5399);
and AND4 (N15562, N15554, N2509, N8444, N1632);
or OR4 (N15563, N15557, N12264, N12681, N11881);
nor NOR4 (N15564, N15560, N6925, N13342, N13096);
xor XOR2 (N15565, N15562, N13618);
nand NAND4 (N15566, N15561, N6889, N7026, N7314);
not NOT1 (N15567, N15541);
and AND2 (N15568, N15563, N5222);
or OR2 (N15569, N15567, N4051);
xor XOR2 (N15570, N15559, N2040);
and AND4 (N15571, N15564, N4660, N3569, N10361);
xor XOR2 (N15572, N15550, N8927);
buf BUF1 (N15573, N15548);
not NOT1 (N15574, N15573);
nor NOR2 (N15575, N15572, N8881);
nand NAND3 (N15576, N15566, N10271, N9554);
and AND2 (N15577, N15568, N13185);
not NOT1 (N15578, N15571);
not NOT1 (N15579, N15575);
not NOT1 (N15580, N15577);
buf BUF1 (N15581, N15580);
not NOT1 (N15582, N15581);
or OR3 (N15583, N15565, N10134, N2342);
xor XOR2 (N15584, N15570, N13370);
or OR2 (N15585, N15576, N9206);
or OR2 (N15586, N15584, N13167);
nor NOR2 (N15587, N15578, N6922);
and AND3 (N15588, N15569, N15530, N256);
nor NOR2 (N15589, N15587, N4744);
buf BUF1 (N15590, N15558);
buf BUF1 (N15591, N15588);
and AND2 (N15592, N15579, N13589);
nand NAND3 (N15593, N15556, N6686, N6715);
xor XOR2 (N15594, N15591, N9058);
nand NAND3 (N15595, N15585, N1567, N13258);
xor XOR2 (N15596, N15593, N2094);
and AND3 (N15597, N15590, N12150, N9892);
buf BUF1 (N15598, N15592);
buf BUF1 (N15599, N15598);
nand NAND3 (N15600, N15599, N15457, N14446);
nand NAND3 (N15601, N15597, N2159, N7199);
xor XOR2 (N15602, N15586, N7082);
nand NAND2 (N15603, N15574, N1177);
nor NOR3 (N15604, N15583, N12906, N4720);
buf BUF1 (N15605, N15596);
or OR4 (N15606, N15602, N10248, N1397, N7894);
nor NOR4 (N15607, N15582, N2809, N3, N11471);
not NOT1 (N15608, N15589);
xor XOR2 (N15609, N15608, N12316);
xor XOR2 (N15610, N15607, N3785);
xor XOR2 (N15611, N15606, N8384);
and AND3 (N15612, N15594, N9027, N3611);
not NOT1 (N15613, N15611);
not NOT1 (N15614, N15613);
nor NOR2 (N15615, N15605, N960);
not NOT1 (N15616, N15615);
and AND3 (N15617, N15600, N1313, N10679);
xor XOR2 (N15618, N15617, N14239);
or OR4 (N15619, N15614, N14919, N5854, N2492);
not NOT1 (N15620, N15603);
or OR2 (N15621, N15618, N7034);
nand NAND3 (N15622, N15601, N7886, N5486);
xor XOR2 (N15623, N15620, N121);
or OR2 (N15624, N15612, N12358);
or OR4 (N15625, N15622, N9548, N4727, N638);
or OR4 (N15626, N15625, N7671, N13027, N10422);
and AND2 (N15627, N15619, N794);
not NOT1 (N15628, N15610);
nor NOR2 (N15629, N15621, N10209);
buf BUF1 (N15630, N15616);
buf BUF1 (N15631, N15628);
buf BUF1 (N15632, N15627);
or OR4 (N15633, N15626, N1966, N4936, N12436);
or OR3 (N15634, N15631, N8333, N7428);
or OR2 (N15635, N15624, N14201);
buf BUF1 (N15636, N15595);
nor NOR3 (N15637, N15632, N6174, N7146);
nor NOR2 (N15638, N15623, N8105);
and AND4 (N15639, N15604, N15608, N645, N15571);
nand NAND4 (N15640, N15633, N14979, N4021, N14959);
xor XOR2 (N15641, N15635, N4966);
and AND2 (N15642, N15636, N10767);
nor NOR3 (N15643, N15642, N6565, N239);
buf BUF1 (N15644, N15609);
nand NAND3 (N15645, N15638, N8964, N13189);
nor NOR2 (N15646, N15634, N12539);
buf BUF1 (N15647, N15646);
not NOT1 (N15648, N15639);
nor NOR4 (N15649, N15637, N1515, N2839, N3860);
and AND4 (N15650, N15629, N7095, N8912, N11477);
not NOT1 (N15651, N15650);
or OR2 (N15652, N15645, N6240);
buf BUF1 (N15653, N15649);
or OR2 (N15654, N15641, N11585);
not NOT1 (N15655, N15653);
and AND2 (N15656, N15651, N8297);
and AND2 (N15657, N15656, N1350);
not NOT1 (N15658, N15630);
not NOT1 (N15659, N15655);
and AND3 (N15660, N15647, N7169, N7815);
and AND4 (N15661, N15654, N9427, N1854, N3336);
buf BUF1 (N15662, N15660);
nand NAND4 (N15663, N15648, N10604, N3283, N3836);
nand NAND4 (N15664, N15652, N4700, N9191, N2359);
buf BUF1 (N15665, N15640);
or OR4 (N15666, N15658, N13886, N12084, N583);
buf BUF1 (N15667, N15661);
or OR2 (N15668, N15662, N8126);
and AND4 (N15669, N15657, N14283, N6732, N9077);
nand NAND3 (N15670, N15659, N640, N13984);
xor XOR2 (N15671, N15670, N5307);
xor XOR2 (N15672, N15668, N4214);
nand NAND3 (N15673, N15672, N7691, N10026);
not NOT1 (N15674, N15664);
xor XOR2 (N15675, N15671, N5356);
xor XOR2 (N15676, N15669, N12158);
buf BUF1 (N15677, N15676);
or OR3 (N15678, N15643, N14750, N2145);
nor NOR3 (N15679, N15675, N6522, N15132);
nand NAND3 (N15680, N15666, N5255, N10859);
not NOT1 (N15681, N15680);
or OR3 (N15682, N15674, N3295, N7959);
buf BUF1 (N15683, N15665);
nand NAND2 (N15684, N15667, N5903);
buf BUF1 (N15685, N15678);
or OR2 (N15686, N15679, N683);
xor XOR2 (N15687, N15686, N13743);
nand NAND2 (N15688, N15681, N3770);
nand NAND4 (N15689, N15684, N12622, N5085, N11579);
xor XOR2 (N15690, N15689, N15643);
and AND4 (N15691, N15687, N2525, N10048, N12400);
not NOT1 (N15692, N15685);
nand NAND4 (N15693, N15691, N14232, N10402, N7430);
or OR3 (N15694, N15692, N637, N10849);
and AND4 (N15695, N15694, N645, N3979, N2764);
and AND2 (N15696, N15688, N7851);
buf BUF1 (N15697, N15690);
or OR4 (N15698, N15697, N5666, N551, N840);
nor NOR4 (N15699, N15695, N8835, N7646, N549);
buf BUF1 (N15700, N15698);
and AND3 (N15701, N15693, N6571, N14931);
nor NOR3 (N15702, N15677, N12741, N13764);
buf BUF1 (N15703, N15644);
buf BUF1 (N15704, N15700);
or OR2 (N15705, N15673, N7514);
and AND2 (N15706, N15705, N6795);
or OR2 (N15707, N15701, N5808);
and AND2 (N15708, N15663, N15656);
and AND3 (N15709, N15703, N9746, N470);
xor XOR2 (N15710, N15704, N2651);
nor NOR2 (N15711, N15708, N1474);
xor XOR2 (N15712, N15711, N6152);
buf BUF1 (N15713, N15709);
nor NOR3 (N15714, N15706, N9660, N14257);
or OR3 (N15715, N15714, N1471, N13874);
and AND4 (N15716, N15710, N6548, N13227, N13707);
or OR3 (N15717, N15716, N9159, N12626);
nand NAND2 (N15718, N15712, N2304);
or OR4 (N15719, N15699, N2831, N6458, N1147);
nor NOR2 (N15720, N15718, N10332);
buf BUF1 (N15721, N15719);
nor NOR4 (N15722, N15702, N10460, N14399, N13472);
xor XOR2 (N15723, N15683, N15429);
nand NAND2 (N15724, N15713, N9213);
nor NOR4 (N15725, N15720, N6721, N12363, N2106);
and AND3 (N15726, N15707, N7682, N9374);
nor NOR4 (N15727, N15721, N6513, N7427, N9165);
not NOT1 (N15728, N15682);
or OR3 (N15729, N15726, N1343, N14815);
not NOT1 (N15730, N15724);
xor XOR2 (N15731, N15728, N14075);
nand NAND4 (N15732, N15729, N2011, N306, N6266);
not NOT1 (N15733, N15722);
xor XOR2 (N15734, N15731, N6016);
buf BUF1 (N15735, N15730);
not NOT1 (N15736, N15715);
buf BUF1 (N15737, N15727);
or OR4 (N15738, N15696, N3405, N1668, N5733);
and AND3 (N15739, N15735, N1082, N5681);
or OR4 (N15740, N15732, N2718, N5353, N12627);
nor NOR2 (N15741, N15734, N11851);
and AND4 (N15742, N15740, N2064, N528, N7715);
nor NOR4 (N15743, N15733, N92, N3234, N3446);
xor XOR2 (N15744, N15738, N6633);
nand NAND3 (N15745, N15737, N13299, N10571);
nand NAND4 (N15746, N15739, N10870, N11925, N14432);
or OR4 (N15747, N15717, N8658, N15589, N9293);
and AND2 (N15748, N15741, N9413);
buf BUF1 (N15749, N15725);
nand NAND4 (N15750, N15742, N3556, N13339, N4150);
nor NOR3 (N15751, N15748, N1374, N10644);
xor XOR2 (N15752, N15736, N1329);
not NOT1 (N15753, N15752);
nor NOR4 (N15754, N15747, N12947, N9519, N9471);
nor NOR4 (N15755, N15751, N2739, N8429, N5520);
buf BUF1 (N15756, N15746);
buf BUF1 (N15757, N15755);
buf BUF1 (N15758, N15754);
buf BUF1 (N15759, N15758);
xor XOR2 (N15760, N15749, N7888);
not NOT1 (N15761, N15744);
buf BUF1 (N15762, N15750);
nand NAND2 (N15763, N15743, N9476);
and AND3 (N15764, N15753, N11332, N8643);
nand NAND4 (N15765, N15760, N9037, N6394, N11834);
nor NOR4 (N15766, N15763, N8999, N8966, N4267);
xor XOR2 (N15767, N15766, N5890);
nand NAND3 (N15768, N15757, N4040, N2935);
buf BUF1 (N15769, N15756);
not NOT1 (N15770, N15761);
and AND2 (N15771, N15759, N13752);
not NOT1 (N15772, N15768);
nor NOR2 (N15773, N15769, N3198);
nor NOR3 (N15774, N15772, N3679, N5641);
nand NAND4 (N15775, N15771, N854, N1048, N1460);
buf BUF1 (N15776, N15767);
buf BUF1 (N15777, N15764);
xor XOR2 (N15778, N15776, N2316);
nor NOR4 (N15779, N15762, N14854, N8528, N3302);
buf BUF1 (N15780, N15774);
or OR2 (N15781, N15723, N12702);
or OR2 (N15782, N15780, N3245);
buf BUF1 (N15783, N15779);
not NOT1 (N15784, N15775);
buf BUF1 (N15785, N15770);
nor NOR4 (N15786, N15781, N5478, N6272, N11834);
not NOT1 (N15787, N15778);
and AND3 (N15788, N15782, N13612, N12632);
nor NOR3 (N15789, N15745, N14803, N13471);
nand NAND2 (N15790, N15783, N11961);
nor NOR2 (N15791, N15787, N829);
not NOT1 (N15792, N15788);
or OR2 (N15793, N15789, N3187);
not NOT1 (N15794, N15777);
and AND3 (N15795, N15794, N10535, N12571);
nor NOR2 (N15796, N15786, N12361);
buf BUF1 (N15797, N15796);
not NOT1 (N15798, N15793);
buf BUF1 (N15799, N15784);
not NOT1 (N15800, N15799);
not NOT1 (N15801, N15797);
nor NOR2 (N15802, N15785, N4180);
xor XOR2 (N15803, N15792, N10808);
not NOT1 (N15804, N15798);
or OR2 (N15805, N15800, N15246);
and AND3 (N15806, N15802, N11153, N490);
xor XOR2 (N15807, N15795, N10664);
nor NOR2 (N15808, N15807, N4700);
not NOT1 (N15809, N15806);
and AND3 (N15810, N15790, N10596, N7024);
xor XOR2 (N15811, N15809, N13426);
or OR3 (N15812, N15773, N2305, N14474);
buf BUF1 (N15813, N15812);
nand NAND3 (N15814, N15803, N6122, N8136);
nor NOR2 (N15815, N15808, N13495);
buf BUF1 (N15816, N15791);
not NOT1 (N15817, N15810);
not NOT1 (N15818, N15814);
buf BUF1 (N15819, N15818);
or OR3 (N15820, N15811, N12275, N4476);
buf BUF1 (N15821, N15820);
nor NOR4 (N15822, N15805, N10580, N385, N5757);
and AND2 (N15823, N15804, N15666);
or OR4 (N15824, N15765, N14408, N8965, N5138);
and AND3 (N15825, N15801, N6611, N11830);
xor XOR2 (N15826, N15815, N6781);
nand NAND3 (N15827, N15823, N2792, N184);
xor XOR2 (N15828, N15821, N3945);
and AND4 (N15829, N15819, N13001, N13391, N14353);
and AND2 (N15830, N15829, N14440);
nand NAND2 (N15831, N15817, N10412);
buf BUF1 (N15832, N15825);
and AND3 (N15833, N15832, N15224, N2003);
nor NOR4 (N15834, N15830, N9720, N2310, N15050);
not NOT1 (N15835, N15831);
or OR3 (N15836, N15824, N11885, N13474);
xor XOR2 (N15837, N15816, N12211);
or OR4 (N15838, N15833, N8221, N6791, N5039);
nand NAND4 (N15839, N15838, N10, N6696, N10479);
nor NOR2 (N15840, N15839, N906);
not NOT1 (N15841, N15827);
or OR2 (N15842, N15837, N15588);
or OR2 (N15843, N15826, N2525);
and AND3 (N15844, N15836, N1879, N6818);
nand NAND2 (N15845, N15835, N604);
buf BUF1 (N15846, N15845);
or OR3 (N15847, N15828, N5674, N7875);
xor XOR2 (N15848, N15813, N4409);
and AND2 (N15849, N15834, N12540);
nor NOR2 (N15850, N15822, N9625);
buf BUF1 (N15851, N15846);
or OR2 (N15852, N15847, N6085);
or OR3 (N15853, N15849, N5413, N4779);
and AND4 (N15854, N15848, N6663, N5617, N6343);
nand NAND3 (N15855, N15841, N9851, N10635);
xor XOR2 (N15856, N15855, N2795);
not NOT1 (N15857, N15840);
buf BUF1 (N15858, N15857);
or OR3 (N15859, N15854, N12135, N12113);
nor NOR3 (N15860, N15852, N13549, N9422);
or OR4 (N15861, N15850, N15200, N11359, N6847);
not NOT1 (N15862, N15860);
not NOT1 (N15863, N15843);
or OR3 (N15864, N15851, N824, N11320);
buf BUF1 (N15865, N15862);
xor XOR2 (N15866, N15853, N11285);
and AND3 (N15867, N15865, N2513, N15787);
not NOT1 (N15868, N15856);
nand NAND4 (N15869, N15866, N13049, N10847, N8592);
nand NAND2 (N15870, N15869, N12772);
buf BUF1 (N15871, N15844);
and AND3 (N15872, N15859, N13041, N11716);
not NOT1 (N15873, N15842);
not NOT1 (N15874, N15873);
buf BUF1 (N15875, N15864);
or OR4 (N15876, N15868, N14121, N10115, N4752);
nand NAND2 (N15877, N15875, N14637);
not NOT1 (N15878, N15872);
not NOT1 (N15879, N15874);
nand NAND2 (N15880, N15877, N13387);
not NOT1 (N15881, N15879);
xor XOR2 (N15882, N15881, N14605);
or OR3 (N15883, N15880, N1417, N6646);
nand NAND2 (N15884, N15882, N11390);
nand NAND2 (N15885, N15867, N361);
buf BUF1 (N15886, N15878);
buf BUF1 (N15887, N15883);
nor NOR3 (N15888, N15876, N10004, N5544);
nand NAND2 (N15889, N15888, N3425);
nor NOR2 (N15890, N15871, N7588);
not NOT1 (N15891, N15863);
and AND4 (N15892, N15884, N383, N8883, N14070);
xor XOR2 (N15893, N15885, N14742);
xor XOR2 (N15894, N15889, N14798);
buf BUF1 (N15895, N15891);
nand NAND3 (N15896, N15894, N3991, N9188);
nor NOR4 (N15897, N15858, N835, N10173, N1730);
nor NOR2 (N15898, N15897, N737);
buf BUF1 (N15899, N15896);
buf BUF1 (N15900, N15887);
buf BUF1 (N15901, N15900);
nand NAND2 (N15902, N15861, N15729);
nand NAND3 (N15903, N15895, N4051, N2808);
xor XOR2 (N15904, N15901, N3208);
or OR3 (N15905, N15892, N6358, N12491);
not NOT1 (N15906, N15890);
nand NAND2 (N15907, N15906, N13875);
buf BUF1 (N15908, N15886);
or OR2 (N15909, N15904, N2963);
not NOT1 (N15910, N15898);
nand NAND2 (N15911, N15907, N12122);
buf BUF1 (N15912, N15908);
nor NOR2 (N15913, N15909, N14933);
xor XOR2 (N15914, N15870, N10559);
or OR2 (N15915, N15910, N11016);
and AND4 (N15916, N15905, N15551, N14725, N12245);
not NOT1 (N15917, N15915);
buf BUF1 (N15918, N15902);
nor NOR3 (N15919, N15899, N2733, N8782);
buf BUF1 (N15920, N15911);
nand NAND3 (N15921, N15918, N9853, N1488);
nor NOR2 (N15922, N15914, N5159);
xor XOR2 (N15923, N15921, N4104);
or OR4 (N15924, N15920, N14983, N1201, N13902);
buf BUF1 (N15925, N15913);
and AND4 (N15926, N15923, N4506, N231, N12103);
xor XOR2 (N15927, N15922, N1897);
nor NOR4 (N15928, N15916, N280, N8574, N11469);
buf BUF1 (N15929, N15917);
nor NOR2 (N15930, N15919, N6760);
nor NOR2 (N15931, N15926, N13000);
xor XOR2 (N15932, N15893, N408);
xor XOR2 (N15933, N15925, N14628);
or OR3 (N15934, N15928, N12457, N799);
and AND2 (N15935, N15927, N13653);
nand NAND2 (N15936, N15934, N7665);
and AND3 (N15937, N15936, N2016, N4378);
nand NAND2 (N15938, N15912, N5897);
not NOT1 (N15939, N15938);
or OR4 (N15940, N15935, N13791, N13206, N10158);
or OR4 (N15941, N15903, N4153, N15038, N4049);
nor NOR4 (N15942, N15930, N3307, N11902, N11889);
buf BUF1 (N15943, N15937);
or OR2 (N15944, N15941, N4399);
xor XOR2 (N15945, N15932, N7581);
nor NOR3 (N15946, N15945, N4055, N6378);
not NOT1 (N15947, N15933);
xor XOR2 (N15948, N15929, N12619);
nand NAND4 (N15949, N15931, N14613, N11892, N13570);
buf BUF1 (N15950, N15942);
nand NAND2 (N15951, N15947, N10066);
nand NAND4 (N15952, N15946, N4391, N11071, N14805);
xor XOR2 (N15953, N15940, N4275);
nor NOR4 (N15954, N15950, N3983, N9978, N8207);
xor XOR2 (N15955, N15952, N10344);
not NOT1 (N15956, N15949);
not NOT1 (N15957, N15943);
xor XOR2 (N15958, N15924, N12084);
and AND3 (N15959, N15953, N14124, N11528);
nor NOR4 (N15960, N15958, N12807, N11741, N8226);
buf BUF1 (N15961, N15939);
buf BUF1 (N15962, N15960);
nand NAND2 (N15963, N15944, N2814);
not NOT1 (N15964, N15963);
nand NAND4 (N15965, N15964, N1323, N10336, N2565);
nand NAND2 (N15966, N15955, N5717);
or OR4 (N15967, N15962, N6927, N7210, N14576);
xor XOR2 (N15968, N15965, N3306);
buf BUF1 (N15969, N15967);
xor XOR2 (N15970, N15968, N541);
and AND3 (N15971, N15961, N1531, N7637);
buf BUF1 (N15972, N15957);
nor NOR3 (N15973, N15969, N12600, N5182);
nand NAND4 (N15974, N15956, N14504, N14823, N8965);
nand NAND4 (N15975, N15951, N529, N13278, N9953);
nand NAND4 (N15976, N15954, N2853, N11269, N7334);
or OR4 (N15977, N15974, N14408, N12857, N11959);
xor XOR2 (N15978, N15977, N14775);
nor NOR3 (N15979, N15966, N13533, N3122);
xor XOR2 (N15980, N15979, N12190);
nor NOR3 (N15981, N15972, N6708, N2943);
xor XOR2 (N15982, N15980, N1799);
not NOT1 (N15983, N15948);
not NOT1 (N15984, N15982);
and AND4 (N15985, N15983, N12869, N9437, N8504);
nand NAND3 (N15986, N15959, N14611, N6995);
nand NAND3 (N15987, N15975, N14102, N12657);
buf BUF1 (N15988, N15986);
nand NAND2 (N15989, N15984, N8253);
nand NAND2 (N15990, N15987, N5112);
and AND4 (N15991, N15990, N3723, N8662, N1576);
not NOT1 (N15992, N15985);
not NOT1 (N15993, N15988);
or OR2 (N15994, N15976, N14910);
xor XOR2 (N15995, N15994, N4308);
or OR4 (N15996, N15970, N15017, N2570, N5504);
nor NOR3 (N15997, N15978, N11598, N7320);
not NOT1 (N15998, N15995);
not NOT1 (N15999, N15997);
and AND2 (N16000, N15971, N5887);
xor XOR2 (N16001, N15992, N14344);
xor XOR2 (N16002, N15996, N7229);
nor NOR3 (N16003, N15998, N1765, N13029);
nor NOR3 (N16004, N15973, N6991, N8445);
not NOT1 (N16005, N16001);
xor XOR2 (N16006, N16002, N15323);
not NOT1 (N16007, N15991);
xor XOR2 (N16008, N15993, N13742);
nand NAND4 (N16009, N16000, N12794, N9500, N13017);
nor NOR2 (N16010, N16006, N14005);
buf BUF1 (N16011, N16004);
and AND2 (N16012, N16011, N8344);
buf BUF1 (N16013, N16005);
or OR3 (N16014, N16003, N13225, N1501);
and AND3 (N16015, N15981, N640, N3117);
buf BUF1 (N16016, N16010);
or OR3 (N16017, N16016, N4613, N5073);
not NOT1 (N16018, N16008);
buf BUF1 (N16019, N15999);
or OR2 (N16020, N15989, N5304);
nor NOR2 (N16021, N16012, N8918);
or OR4 (N16022, N16009, N8820, N1112, N15545);
buf BUF1 (N16023, N16013);
not NOT1 (N16024, N16019);
not NOT1 (N16025, N16007);
nand NAND3 (N16026, N16017, N13862, N5181);
or OR3 (N16027, N16025, N15812, N13260);
not NOT1 (N16028, N16015);
or OR2 (N16029, N16027, N15061);
or OR4 (N16030, N16026, N130, N3915, N2381);
nand NAND3 (N16031, N16022, N2920, N1616);
nor NOR2 (N16032, N16024, N1060);
buf BUF1 (N16033, N16028);
nor NOR3 (N16034, N16030, N12813, N8007);
buf BUF1 (N16035, N16014);
nor NOR3 (N16036, N16023, N10571, N6333);
buf BUF1 (N16037, N16031);
or OR3 (N16038, N16032, N4516, N2015);
xor XOR2 (N16039, N16018, N1107);
buf BUF1 (N16040, N16029);
buf BUF1 (N16041, N16020);
and AND4 (N16042, N16039, N15875, N2195, N5573);
nand NAND3 (N16043, N16035, N12501, N12701);
nor NOR2 (N16044, N16034, N12695);
buf BUF1 (N16045, N16040);
nor NOR4 (N16046, N16045, N13045, N5781, N14254);
nor NOR2 (N16047, N16038, N2344);
buf BUF1 (N16048, N16036);
not NOT1 (N16049, N16021);
and AND3 (N16050, N16041, N8333, N10862);
xor XOR2 (N16051, N16037, N4646);
buf BUF1 (N16052, N16033);
nand NAND2 (N16053, N16050, N4739);
or OR3 (N16054, N16044, N6555, N13623);
nor NOR3 (N16055, N16046, N2689, N6497);
not NOT1 (N16056, N16051);
nand NAND2 (N16057, N16047, N822);
and AND4 (N16058, N16056, N4589, N10747, N2531);
nor NOR4 (N16059, N16048, N9180, N10874, N1725);
buf BUF1 (N16060, N16058);
not NOT1 (N16061, N16042);
and AND4 (N16062, N16053, N1231, N1632, N11731);
and AND2 (N16063, N16060, N5422);
and AND4 (N16064, N16062, N8501, N14265, N11334);
nor NOR4 (N16065, N16052, N14733, N5646, N5133);
buf BUF1 (N16066, N16059);
not NOT1 (N16067, N16065);
nor NOR3 (N16068, N16066, N5752, N2479);
nand NAND2 (N16069, N16055, N930);
and AND4 (N16070, N16054, N1445, N3849, N4408);
not NOT1 (N16071, N16068);
not NOT1 (N16072, N16070);
not NOT1 (N16073, N16069);
not NOT1 (N16074, N16063);
not NOT1 (N16075, N16057);
not NOT1 (N16076, N16043);
not NOT1 (N16077, N16074);
or OR4 (N16078, N16076, N15029, N11813, N15659);
not NOT1 (N16079, N16077);
buf BUF1 (N16080, N16078);
and AND2 (N16081, N16072, N4588);
xor XOR2 (N16082, N16073, N6952);
xor XOR2 (N16083, N16067, N6911);
or OR4 (N16084, N16079, N7955, N13181, N2966);
nand NAND2 (N16085, N16061, N6676);
not NOT1 (N16086, N16071);
and AND4 (N16087, N16080, N1551, N7838, N14327);
nor NOR2 (N16088, N16085, N13650);
not NOT1 (N16089, N16088);
not NOT1 (N16090, N16084);
nand NAND2 (N16091, N16064, N4890);
or OR3 (N16092, N16083, N5595, N11481);
nand NAND4 (N16093, N16081, N14673, N11346, N4019);
or OR3 (N16094, N16093, N1028, N4891);
nand NAND3 (N16095, N16089, N7754, N15654);
and AND2 (N16096, N16086, N12428);
nand NAND4 (N16097, N16082, N7421, N3657, N8983);
or OR2 (N16098, N16095, N4127);
not NOT1 (N16099, N16098);
buf BUF1 (N16100, N16090);
buf BUF1 (N16101, N16099);
buf BUF1 (N16102, N16096);
xor XOR2 (N16103, N16091, N14295);
buf BUF1 (N16104, N16103);
buf BUF1 (N16105, N16075);
nand NAND2 (N16106, N16101, N9930);
buf BUF1 (N16107, N16094);
not NOT1 (N16108, N16104);
nor NOR4 (N16109, N16097, N13140, N14818, N12587);
or OR3 (N16110, N16102, N3123, N10879);
nor NOR4 (N16111, N16100, N12758, N613, N11719);
and AND4 (N16112, N16111, N6085, N5779, N9458);
nand NAND4 (N16113, N16110, N14862, N4843, N12894);
xor XOR2 (N16114, N16106, N4320);
buf BUF1 (N16115, N16087);
or OR4 (N16116, N16113, N4624, N3667, N779);
and AND2 (N16117, N16116, N11689);
buf BUF1 (N16118, N16107);
xor XOR2 (N16119, N16109, N974);
nand NAND2 (N16120, N16049, N5710);
not NOT1 (N16121, N16112);
not NOT1 (N16122, N16108);
buf BUF1 (N16123, N16117);
xor XOR2 (N16124, N16120, N920);
and AND4 (N16125, N16122, N13019, N5424, N12040);
or OR3 (N16126, N16124, N14269, N13193);
or OR3 (N16127, N16121, N3466, N12246);
or OR2 (N16128, N16115, N11141);
nor NOR2 (N16129, N16092, N10283);
not NOT1 (N16130, N16127);
nor NOR3 (N16131, N16105, N3853, N8237);
nand NAND2 (N16132, N16129, N13142);
nor NOR2 (N16133, N16119, N1648);
and AND3 (N16134, N16118, N6117, N2007);
buf BUF1 (N16135, N16114);
buf BUF1 (N16136, N16134);
and AND4 (N16137, N16136, N16026, N6044, N158);
and AND3 (N16138, N16125, N2664, N10105);
xor XOR2 (N16139, N16137, N3319);
nand NAND2 (N16140, N16135, N14680);
xor XOR2 (N16141, N16130, N14928);
not NOT1 (N16142, N16141);
buf BUF1 (N16143, N16126);
xor XOR2 (N16144, N16131, N9498);
and AND4 (N16145, N16142, N13897, N14703, N4524);
not NOT1 (N16146, N16145);
nor NOR2 (N16147, N16139, N14815);
xor XOR2 (N16148, N16128, N9392);
xor XOR2 (N16149, N16143, N3413);
not NOT1 (N16150, N16140);
not NOT1 (N16151, N16149);
nor NOR4 (N16152, N16147, N15204, N13848, N13320);
not NOT1 (N16153, N16150);
nor NOR4 (N16154, N16132, N1890, N1658, N2498);
buf BUF1 (N16155, N16152);
or OR3 (N16156, N16151, N4038, N3195);
buf BUF1 (N16157, N16144);
nand NAND3 (N16158, N16154, N5979, N10329);
buf BUF1 (N16159, N16138);
or OR2 (N16160, N16157, N7500);
or OR4 (N16161, N16156, N4, N10690, N2925);
or OR4 (N16162, N16148, N10268, N3416, N7261);
and AND2 (N16163, N16158, N11751);
nand NAND3 (N16164, N16155, N11498, N11766);
xor XOR2 (N16165, N16133, N2906);
and AND4 (N16166, N16159, N723, N14121, N4349);
nor NOR2 (N16167, N16164, N12410);
xor XOR2 (N16168, N16160, N10248);
xor XOR2 (N16169, N16168, N6032);
nor NOR2 (N16170, N16162, N9933);
or OR2 (N16171, N16167, N1304);
or OR3 (N16172, N16163, N10578, N2072);
xor XOR2 (N16173, N16153, N2653);
nor NOR4 (N16174, N16146, N3200, N9957, N4788);
xor XOR2 (N16175, N16171, N8054);
nand NAND3 (N16176, N16174, N9520, N11227);
not NOT1 (N16177, N16123);
not NOT1 (N16178, N16166);
nor NOR4 (N16179, N16175, N5717, N14724, N10344);
nor NOR2 (N16180, N16170, N7164);
buf BUF1 (N16181, N16179);
buf BUF1 (N16182, N16180);
not NOT1 (N16183, N16181);
buf BUF1 (N16184, N16177);
and AND2 (N16185, N16176, N1061);
nand NAND4 (N16186, N16161, N12832, N15291, N11719);
nand NAND2 (N16187, N16165, N2862);
buf BUF1 (N16188, N16183);
or OR3 (N16189, N16188, N11347, N11518);
not NOT1 (N16190, N16169);
not NOT1 (N16191, N16189);
or OR3 (N16192, N16173, N13337, N9251);
and AND2 (N16193, N16172, N5578);
not NOT1 (N16194, N16187);
xor XOR2 (N16195, N16182, N11368);
xor XOR2 (N16196, N16191, N8587);
or OR3 (N16197, N16193, N4597, N9254);
not NOT1 (N16198, N16196);
nand NAND3 (N16199, N16186, N13077, N5243);
or OR3 (N16200, N16197, N5862, N14840);
buf BUF1 (N16201, N16199);
nor NOR4 (N16202, N16178, N11929, N15062, N1593);
nor NOR4 (N16203, N16184, N15003, N6546, N8569);
xor XOR2 (N16204, N16202, N7183);
and AND2 (N16205, N16198, N1165);
and AND4 (N16206, N16200, N2719, N10042, N5284);
nand NAND4 (N16207, N16203, N7704, N10668, N15883);
not NOT1 (N16208, N16207);
not NOT1 (N16209, N16194);
nand NAND3 (N16210, N16195, N7845, N4842);
buf BUF1 (N16211, N16209);
not NOT1 (N16212, N16190);
or OR4 (N16213, N16206, N13825, N9698, N12155);
xor XOR2 (N16214, N16208, N12864);
or OR2 (N16215, N16210, N8288);
nand NAND4 (N16216, N16211, N5509, N13307, N12451);
not NOT1 (N16217, N16212);
xor XOR2 (N16218, N16204, N14888);
or OR2 (N16219, N16213, N2584);
not NOT1 (N16220, N16215);
or OR2 (N16221, N16217, N15591);
and AND2 (N16222, N16216, N9850);
nand NAND3 (N16223, N16205, N15055, N725);
and AND4 (N16224, N16218, N5637, N12718, N1225);
or OR2 (N16225, N16214, N4353);
not NOT1 (N16226, N16221);
buf BUF1 (N16227, N16222);
nor NOR4 (N16228, N16220, N87, N9827, N6418);
and AND4 (N16229, N16192, N5824, N13889, N16121);
nor NOR4 (N16230, N16228, N2135, N6980, N10748);
or OR4 (N16231, N16201, N5026, N1129, N14930);
or OR4 (N16232, N16226, N15408, N1327, N1669);
not NOT1 (N16233, N16231);
and AND3 (N16234, N16232, N551, N10849);
buf BUF1 (N16235, N16219);
xor XOR2 (N16236, N16223, N7796);
nor NOR2 (N16237, N16233, N11595);
not NOT1 (N16238, N16185);
not NOT1 (N16239, N16236);
and AND3 (N16240, N16234, N4715, N12672);
xor XOR2 (N16241, N16224, N12511);
xor XOR2 (N16242, N16240, N217);
nor NOR3 (N16243, N16225, N4631, N7593);
and AND3 (N16244, N16238, N7383, N7414);
not NOT1 (N16245, N16239);
xor XOR2 (N16246, N16242, N2777);
nor NOR4 (N16247, N16237, N8076, N1775, N15742);
not NOT1 (N16248, N16230);
buf BUF1 (N16249, N16241);
and AND2 (N16250, N16244, N2735);
nand NAND2 (N16251, N16227, N7135);
and AND4 (N16252, N16247, N14091, N2994, N464);
nand NAND3 (N16253, N16229, N8603, N3163);
nand NAND4 (N16254, N16248, N10645, N14925, N7683);
xor XOR2 (N16255, N16252, N1899);
nand NAND2 (N16256, N16253, N9528);
not NOT1 (N16257, N16243);
and AND2 (N16258, N16245, N11019);
not NOT1 (N16259, N16246);
and AND2 (N16260, N16254, N11844);
or OR2 (N16261, N16255, N14620);
nor NOR4 (N16262, N16256, N4995, N14430, N603);
or OR4 (N16263, N16258, N213, N1696, N15764);
not NOT1 (N16264, N16259);
nand NAND2 (N16265, N16235, N5336);
and AND2 (N16266, N16263, N12892);
nand NAND2 (N16267, N16260, N22);
not NOT1 (N16268, N16251);
or OR2 (N16269, N16264, N33);
buf BUF1 (N16270, N16268);
not NOT1 (N16271, N16249);
xor XOR2 (N16272, N16265, N7144);
and AND3 (N16273, N16270, N8606, N9498);
and AND2 (N16274, N16261, N1941);
not NOT1 (N16275, N16262);
nor NOR2 (N16276, N16272, N11188);
buf BUF1 (N16277, N16273);
and AND3 (N16278, N16267, N2799, N2063);
not NOT1 (N16279, N16257);
nor NOR3 (N16280, N16278, N6298, N5047);
buf BUF1 (N16281, N16280);
xor XOR2 (N16282, N16274, N16022);
nor NOR2 (N16283, N16276, N13128);
nor NOR2 (N16284, N16271, N14218);
buf BUF1 (N16285, N16275);
and AND2 (N16286, N16269, N10255);
or OR4 (N16287, N16266, N3727, N6771, N13320);
nand NAND3 (N16288, N16283, N3499, N15781);
xor XOR2 (N16289, N16277, N5689);
xor XOR2 (N16290, N16285, N1228);
not NOT1 (N16291, N16281);
and AND2 (N16292, N16279, N10717);
and AND2 (N16293, N16289, N548);
xor XOR2 (N16294, N16292, N3605);
nor NOR2 (N16295, N16293, N8127);
xor XOR2 (N16296, N16286, N3004);
xor XOR2 (N16297, N16282, N15403);
nor NOR4 (N16298, N16284, N12705, N13489, N4016);
nor NOR2 (N16299, N16295, N8240);
nand NAND2 (N16300, N16294, N5872);
or OR3 (N16301, N16288, N8192, N3739);
not NOT1 (N16302, N16300);
nand NAND3 (N16303, N16287, N6318, N6085);
buf BUF1 (N16304, N16301);
and AND3 (N16305, N16302, N4316, N8796);
and AND4 (N16306, N16304, N2139, N4178, N12259);
not NOT1 (N16307, N16298);
not NOT1 (N16308, N16290);
buf BUF1 (N16309, N16303);
or OR2 (N16310, N16291, N11479);
and AND2 (N16311, N16299, N8611);
xor XOR2 (N16312, N16250, N1746);
nand NAND4 (N16313, N16308, N15849, N13417, N9101);
xor XOR2 (N16314, N16297, N4599);
xor XOR2 (N16315, N16307, N8965);
xor XOR2 (N16316, N16314, N6683);
nand NAND4 (N16317, N16313, N10554, N15203, N15963);
nor NOR2 (N16318, N16311, N4048);
xor XOR2 (N16319, N16318, N14747);
not NOT1 (N16320, N16319);
buf BUF1 (N16321, N16309);
buf BUF1 (N16322, N16316);
nor NOR3 (N16323, N16320, N10081, N13019);
or OR2 (N16324, N16305, N10138);
or OR2 (N16325, N16322, N9923);
and AND2 (N16326, N16324, N1131);
xor XOR2 (N16327, N16323, N10729);
nand NAND3 (N16328, N16315, N10621, N2610);
and AND3 (N16329, N16296, N2299, N4737);
or OR4 (N16330, N16328, N14679, N12151, N12310);
not NOT1 (N16331, N16321);
buf BUF1 (N16332, N16306);
or OR3 (N16333, N16329, N13740, N5089);
buf BUF1 (N16334, N16310);
and AND2 (N16335, N16333, N4100);
buf BUF1 (N16336, N16326);
or OR3 (N16337, N16334, N11815, N5315);
and AND3 (N16338, N16332, N8517, N7889);
nand NAND3 (N16339, N16331, N14253, N6454);
nor NOR4 (N16340, N16312, N6762, N14657, N2228);
buf BUF1 (N16341, N16327);
and AND2 (N16342, N16336, N7940);
buf BUF1 (N16343, N16340);
nand NAND3 (N16344, N16337, N4412, N15917);
or OR3 (N16345, N16330, N8323, N4166);
xor XOR2 (N16346, N16325, N10053);
nor NOR3 (N16347, N16335, N9772, N15544);
not NOT1 (N16348, N16347);
and AND4 (N16349, N16344, N808, N3188, N8273);
not NOT1 (N16350, N16346);
nand NAND3 (N16351, N16338, N11498, N8259);
and AND2 (N16352, N16345, N3090);
and AND4 (N16353, N16352, N8714, N15125, N7373);
nand NAND4 (N16354, N16353, N11589, N6610, N14428);
or OR2 (N16355, N16349, N9039);
nor NOR2 (N16356, N16339, N9221);
not NOT1 (N16357, N16342);
nand NAND3 (N16358, N16355, N6393, N15215);
buf BUF1 (N16359, N16354);
not NOT1 (N16360, N16356);
not NOT1 (N16361, N16360);
or OR2 (N16362, N16350, N3196);
or OR2 (N16363, N16348, N15334);
buf BUF1 (N16364, N16317);
xor XOR2 (N16365, N16364, N3035);
not NOT1 (N16366, N16351);
xor XOR2 (N16367, N16365, N10732);
or OR2 (N16368, N16361, N7077);
not NOT1 (N16369, N16359);
nand NAND2 (N16370, N16362, N13727);
or OR2 (N16371, N16368, N1585);
nand NAND3 (N16372, N16357, N14906, N10554);
and AND3 (N16373, N16343, N14580, N7028);
xor XOR2 (N16374, N16363, N13487);
or OR2 (N16375, N16371, N15306);
or OR4 (N16376, N16373, N11158, N11013, N5086);
not NOT1 (N16377, N16366);
and AND2 (N16378, N16358, N15446);
and AND4 (N16379, N16367, N2771, N13486, N9413);
or OR3 (N16380, N16370, N10122, N6650);
or OR4 (N16381, N16380, N12325, N5771, N6780);
or OR4 (N16382, N16381, N4885, N523, N13502);
xor XOR2 (N16383, N16372, N8763);
or OR3 (N16384, N16376, N5940, N14496);
nand NAND3 (N16385, N16377, N3109, N8672);
and AND4 (N16386, N16378, N396, N12477, N1993);
not NOT1 (N16387, N16369);
nand NAND3 (N16388, N16375, N1597, N5347);
or OR3 (N16389, N16379, N2797, N2061);
xor XOR2 (N16390, N16388, N9665);
not NOT1 (N16391, N16385);
and AND3 (N16392, N16384, N7759, N14719);
buf BUF1 (N16393, N16383);
buf BUF1 (N16394, N16391);
xor XOR2 (N16395, N16341, N3571);
nand NAND3 (N16396, N16389, N16077, N13621);
nand NAND3 (N16397, N16392, N10485, N3869);
or OR3 (N16398, N16390, N6536, N878);
or OR4 (N16399, N16397, N2395, N1592, N9251);
buf BUF1 (N16400, N16382);
xor XOR2 (N16401, N16400, N5029);
nand NAND4 (N16402, N16374, N9802, N16370, N10891);
or OR2 (N16403, N16399, N6244);
not NOT1 (N16404, N16401);
nor NOR2 (N16405, N16404, N6155);
or OR2 (N16406, N16394, N9829);
buf BUF1 (N16407, N16387);
buf BUF1 (N16408, N16405);
not NOT1 (N16409, N16398);
nand NAND3 (N16410, N16403, N4392, N8297);
not NOT1 (N16411, N16386);
xor XOR2 (N16412, N16409, N12925);
or OR3 (N16413, N16393, N2159, N10377);
nor NOR2 (N16414, N16413, N6460);
xor XOR2 (N16415, N16412, N16061);
or OR2 (N16416, N16414, N8496);
xor XOR2 (N16417, N16415, N10558);
buf BUF1 (N16418, N16417);
and AND3 (N16419, N16408, N9946, N14843);
not NOT1 (N16420, N16406);
and AND2 (N16421, N16410, N5180);
xor XOR2 (N16422, N16418, N768);
and AND3 (N16423, N16422, N16092, N12873);
xor XOR2 (N16424, N16416, N7090);
nor NOR4 (N16425, N16411, N11638, N8104, N5035);
or OR4 (N16426, N16419, N4032, N16423, N14900);
nand NAND3 (N16427, N9061, N5660, N2310);
nor NOR2 (N16428, N16424, N3384);
and AND3 (N16429, N16428, N4980, N4942);
and AND2 (N16430, N16420, N11771);
nor NOR3 (N16431, N16426, N13848, N3332);
not NOT1 (N16432, N16425);
buf BUF1 (N16433, N16407);
and AND3 (N16434, N16402, N6880, N7989);
nor NOR2 (N16435, N16431, N3939);
nor NOR4 (N16436, N16432, N2882, N14908, N11378);
not NOT1 (N16437, N16395);
or OR2 (N16438, N16433, N2338);
not NOT1 (N16439, N16434);
xor XOR2 (N16440, N16430, N1690);
and AND2 (N16441, N16440, N8439);
nand NAND4 (N16442, N16421, N6253, N3090, N10447);
nor NOR2 (N16443, N16429, N11684);
xor XOR2 (N16444, N16441, N6229);
nand NAND3 (N16445, N16439, N8148, N14414);
and AND4 (N16446, N16427, N3394, N14669, N2812);
nand NAND3 (N16447, N16446, N11125, N4689);
xor XOR2 (N16448, N16444, N2945);
or OR3 (N16449, N16445, N569, N1491);
nor NOR2 (N16450, N16435, N12899);
xor XOR2 (N16451, N16449, N13420);
xor XOR2 (N16452, N16436, N10759);
buf BUF1 (N16453, N16448);
nor NOR3 (N16454, N16450, N4747, N12894);
and AND2 (N16455, N16438, N4067);
not NOT1 (N16456, N16443);
xor XOR2 (N16457, N16456, N13946);
not NOT1 (N16458, N16447);
xor XOR2 (N16459, N16451, N9528);
nand NAND4 (N16460, N16457, N3161, N11519, N2375);
and AND2 (N16461, N16458, N3005);
nor NOR2 (N16462, N16396, N16294);
nand NAND3 (N16463, N16442, N15681, N6355);
xor XOR2 (N16464, N16463, N10757);
buf BUF1 (N16465, N16460);
or OR2 (N16466, N16455, N940);
nand NAND2 (N16467, N16452, N13484);
or OR4 (N16468, N16459, N5138, N937, N7482);
not NOT1 (N16469, N16464);
buf BUF1 (N16470, N16465);
nand NAND3 (N16471, N16437, N16174, N6421);
nand NAND2 (N16472, N16453, N12459);
xor XOR2 (N16473, N16462, N15559);
or OR4 (N16474, N16469, N14797, N12579, N16068);
xor XOR2 (N16475, N16471, N7092);
not NOT1 (N16476, N16470);
not NOT1 (N16477, N16474);
or OR2 (N16478, N16475, N8751);
nor NOR4 (N16479, N16467, N7263, N2407, N9703);
nor NOR3 (N16480, N16479, N7061, N16272);
and AND3 (N16481, N16478, N8268, N16366);
xor XOR2 (N16482, N16477, N9007);
buf BUF1 (N16483, N16461);
nand NAND4 (N16484, N16466, N12915, N13069, N7961);
and AND4 (N16485, N16482, N6993, N16018, N8804);
or OR2 (N16486, N16481, N6093);
or OR2 (N16487, N16472, N1249);
not NOT1 (N16488, N16486);
not NOT1 (N16489, N16476);
or OR2 (N16490, N16454, N2848);
xor XOR2 (N16491, N16487, N11692);
nor NOR3 (N16492, N16489, N6668, N407);
xor XOR2 (N16493, N16488, N6881);
nor NOR2 (N16494, N16491, N10305);
nand NAND4 (N16495, N16485, N15740, N10205, N11976);
and AND4 (N16496, N16490, N4349, N868, N6621);
nor NOR4 (N16497, N16494, N2184, N622, N11080);
not NOT1 (N16498, N16497);
xor XOR2 (N16499, N16495, N7783);
xor XOR2 (N16500, N16498, N13697);
buf BUF1 (N16501, N16492);
nand NAND3 (N16502, N16500, N9320, N15272);
xor XOR2 (N16503, N16499, N4597);
buf BUF1 (N16504, N16496);
nor NOR2 (N16505, N16503, N15067);
and AND3 (N16506, N16484, N5920, N7137);
or OR2 (N16507, N16493, N6536);
nand NAND2 (N16508, N16473, N15233);
and AND4 (N16509, N16504, N4895, N11399, N7832);
buf BUF1 (N16510, N16468);
nand NAND2 (N16511, N16483, N12982);
nand NAND2 (N16512, N16506, N3023);
xor XOR2 (N16513, N16505, N6651);
and AND3 (N16514, N16511, N2489, N12326);
and AND4 (N16515, N16512, N9505, N6193, N14786);
not NOT1 (N16516, N16507);
or OR3 (N16517, N16513, N13891, N5388);
or OR4 (N16518, N16509, N10725, N10966, N3573);
or OR3 (N16519, N16515, N14155, N450);
and AND2 (N16520, N16508, N2173);
nand NAND3 (N16521, N16516, N10549, N12129);
xor XOR2 (N16522, N16502, N5652);
buf BUF1 (N16523, N16519);
buf BUF1 (N16524, N16522);
or OR4 (N16525, N16514, N13340, N13479, N9252);
or OR4 (N16526, N16480, N13716, N10943, N4643);
buf BUF1 (N16527, N16525);
not NOT1 (N16528, N16521);
nor NOR3 (N16529, N16518, N8999, N11762);
not NOT1 (N16530, N16520);
nor NOR4 (N16531, N16501, N3797, N9238, N1336);
nand NAND2 (N16532, N16527, N15024);
nor NOR4 (N16533, N16531, N1652, N13908, N11104);
not NOT1 (N16534, N16533);
and AND4 (N16535, N16528, N15254, N15132, N8213);
nor NOR2 (N16536, N16524, N8576);
buf BUF1 (N16537, N16517);
and AND4 (N16538, N16530, N11001, N10762, N4277);
buf BUF1 (N16539, N16523);
and AND2 (N16540, N16532, N9615);
not NOT1 (N16541, N16534);
nand NAND3 (N16542, N16539, N8370, N4478);
or OR3 (N16543, N16529, N14653, N12650);
and AND4 (N16544, N16540, N13375, N4636, N6003);
or OR4 (N16545, N16544, N5977, N9145, N7861);
xor XOR2 (N16546, N16541, N2338);
and AND4 (N16547, N16510, N12305, N684, N10471);
buf BUF1 (N16548, N16535);
nor NOR4 (N16549, N16538, N8128, N8550, N4702);
or OR3 (N16550, N16547, N11685, N8011);
nand NAND4 (N16551, N16545, N728, N12097, N15269);
not NOT1 (N16552, N16543);
and AND3 (N16553, N16537, N15412, N10313);
xor XOR2 (N16554, N16546, N1516);
not NOT1 (N16555, N16536);
nor NOR4 (N16556, N16548, N15718, N4282, N13512);
xor XOR2 (N16557, N16542, N7154);
not NOT1 (N16558, N16556);
nor NOR3 (N16559, N16557, N6125, N12581);
nand NAND2 (N16560, N16558, N5536);
not NOT1 (N16561, N16559);
nor NOR4 (N16562, N16554, N11558, N2865, N11100);
nand NAND4 (N16563, N16526, N2125, N8275, N3434);
nor NOR2 (N16564, N16555, N2590);
buf BUF1 (N16565, N16564);
not NOT1 (N16566, N16551);
xor XOR2 (N16567, N16562, N1954);
or OR3 (N16568, N16550, N7124, N2617);
nor NOR4 (N16569, N16549, N12999, N12957, N4071);
not NOT1 (N16570, N16569);
nor NOR3 (N16571, N16552, N6907, N8838);
nand NAND3 (N16572, N16568, N3213, N11148);
xor XOR2 (N16573, N16565, N674);
and AND2 (N16574, N16566, N10458);
nand NAND4 (N16575, N16567, N15832, N3813, N2308);
nand NAND2 (N16576, N16572, N8926);
buf BUF1 (N16577, N16574);
or OR2 (N16578, N16573, N11193);
not NOT1 (N16579, N16578);
not NOT1 (N16580, N16560);
xor XOR2 (N16581, N16571, N12227);
buf BUF1 (N16582, N16576);
nor NOR4 (N16583, N16561, N10169, N7068, N13930);
nand NAND3 (N16584, N16580, N15038, N7647);
or OR4 (N16585, N16581, N8508, N12881, N7828);
buf BUF1 (N16586, N16582);
xor XOR2 (N16587, N16579, N1897);
nor NOR3 (N16588, N16563, N1481, N5566);
nor NOR3 (N16589, N16585, N7333, N11175);
nand NAND2 (N16590, N16587, N13725);
or OR2 (N16591, N16584, N13515);
xor XOR2 (N16592, N16591, N9098);
not NOT1 (N16593, N16570);
not NOT1 (N16594, N16575);
and AND2 (N16595, N16592, N4404);
buf BUF1 (N16596, N16593);
xor XOR2 (N16597, N16589, N5688);
nand NAND4 (N16598, N16586, N10529, N7756, N12311);
nor NOR4 (N16599, N16598, N607, N13747, N16104);
nor NOR3 (N16600, N16596, N12287, N10744);
not NOT1 (N16601, N16588);
nand NAND3 (N16602, N16597, N14320, N3736);
nor NOR4 (N16603, N16595, N10813, N6293, N1577);
and AND4 (N16604, N16590, N13252, N13983, N4068);
or OR4 (N16605, N16594, N7215, N15521, N4108);
xor XOR2 (N16606, N16583, N172);
nand NAND2 (N16607, N16553, N8565);
or OR2 (N16608, N16606, N2988);
not NOT1 (N16609, N16607);
or OR3 (N16610, N16609, N9359, N5490);
xor XOR2 (N16611, N16577, N2534);
and AND4 (N16612, N16601, N5348, N6356, N8658);
not NOT1 (N16613, N16608);
and AND2 (N16614, N16610, N8184);
nor NOR2 (N16615, N16612, N10595);
and AND4 (N16616, N16602, N4720, N12786, N8559);
or OR2 (N16617, N16611, N5593);
xor XOR2 (N16618, N16599, N15315);
xor XOR2 (N16619, N16605, N9664);
nand NAND4 (N16620, N16600, N9296, N7616, N1826);
and AND2 (N16621, N16619, N16394);
buf BUF1 (N16622, N16616);
buf BUF1 (N16623, N16613);
xor XOR2 (N16624, N16620, N16322);
xor XOR2 (N16625, N16618, N8690);
and AND4 (N16626, N16622, N4297, N9677, N14908);
xor XOR2 (N16627, N16604, N2295);
or OR2 (N16628, N16617, N14483);
xor XOR2 (N16629, N16614, N5518);
nand NAND3 (N16630, N16624, N451, N1904);
and AND2 (N16631, N16623, N7799);
not NOT1 (N16632, N16621);
and AND3 (N16633, N16615, N13495, N12012);
or OR4 (N16634, N16632, N8163, N3850, N14239);
and AND2 (N16635, N16629, N3055);
not NOT1 (N16636, N16631);
and AND4 (N16637, N16634, N16535, N3828, N4502);
buf BUF1 (N16638, N16625);
nor NOR2 (N16639, N16636, N15937);
nand NAND2 (N16640, N16628, N14268);
xor XOR2 (N16641, N16639, N12401);
not NOT1 (N16642, N16627);
not NOT1 (N16643, N16642);
nand NAND2 (N16644, N16626, N11208);
or OR4 (N16645, N16603, N7632, N11655, N15733);
nor NOR2 (N16646, N16644, N10201);
not NOT1 (N16647, N16633);
or OR2 (N16648, N16640, N9078);
not NOT1 (N16649, N16647);
or OR2 (N16650, N16641, N11900);
or OR4 (N16651, N16635, N4841, N122, N11330);
nand NAND2 (N16652, N16638, N14420);
not NOT1 (N16653, N16630);
nand NAND3 (N16654, N16649, N3846, N6846);
xor XOR2 (N16655, N16643, N2870);
nand NAND2 (N16656, N16648, N15196);
xor XOR2 (N16657, N16651, N10224);
not NOT1 (N16658, N16656);
nand NAND2 (N16659, N16637, N7012);
and AND4 (N16660, N16653, N10808, N6202, N7794);
nor NOR2 (N16661, N16655, N3086);
not NOT1 (N16662, N16660);
not NOT1 (N16663, N16659);
nand NAND2 (N16664, N16658, N8637);
nor NOR3 (N16665, N16662, N8909, N14280);
nor NOR4 (N16666, N16646, N10459, N1132, N10955);
xor XOR2 (N16667, N16663, N7657);
nand NAND3 (N16668, N16652, N3228, N7847);
and AND4 (N16669, N16645, N16093, N11689, N1640);
nor NOR2 (N16670, N16654, N7150);
buf BUF1 (N16671, N16670);
not NOT1 (N16672, N16657);
not NOT1 (N16673, N16672);
and AND4 (N16674, N16661, N5146, N11122, N15860);
buf BUF1 (N16675, N16668);
xor XOR2 (N16676, N16671, N718);
buf BUF1 (N16677, N16667);
not NOT1 (N16678, N16676);
or OR2 (N16679, N16666, N3591);
or OR4 (N16680, N16679, N4744, N9358, N14863);
not NOT1 (N16681, N16678);
xor XOR2 (N16682, N16669, N1873);
not NOT1 (N16683, N16665);
nor NOR3 (N16684, N16677, N14647, N10942);
nor NOR2 (N16685, N16650, N2737);
buf BUF1 (N16686, N16680);
not NOT1 (N16687, N16674);
nor NOR3 (N16688, N16687, N14052, N16163);
and AND3 (N16689, N16683, N13982, N1064);
or OR3 (N16690, N16685, N9011, N15067);
nor NOR2 (N16691, N16684, N10588);
nand NAND3 (N16692, N16690, N522, N13187);
buf BUF1 (N16693, N16673);
or OR4 (N16694, N16689, N15756, N671, N15446);
or OR2 (N16695, N16688, N13414);
nor NOR3 (N16696, N16686, N4472, N4218);
nor NOR2 (N16697, N16675, N2373);
buf BUF1 (N16698, N16696);
xor XOR2 (N16699, N16694, N2117);
xor XOR2 (N16700, N16681, N12143);
buf BUF1 (N16701, N16700);
nand NAND3 (N16702, N16691, N808, N4851);
buf BUF1 (N16703, N16664);
nand NAND4 (N16704, N16693, N7928, N16357, N10888);
nand NAND2 (N16705, N16695, N3189);
and AND3 (N16706, N16699, N13063, N13822);
nand NAND3 (N16707, N16697, N6538, N456);
buf BUF1 (N16708, N16692);
xor XOR2 (N16709, N16704, N5676);
or OR4 (N16710, N16707, N12285, N12809, N9509);
and AND3 (N16711, N16705, N14581, N8261);
not NOT1 (N16712, N16708);
or OR2 (N16713, N16698, N12550);
nand NAND3 (N16714, N16711, N1560, N3319);
nand NAND2 (N16715, N16709, N9116);
nand NAND2 (N16716, N16701, N2256);
nand NAND3 (N16717, N16703, N5875, N2238);
and AND3 (N16718, N16713, N14241, N269);
not NOT1 (N16719, N16710);
not NOT1 (N16720, N16706);
nor NOR3 (N16721, N16682, N8007, N408);
buf BUF1 (N16722, N16720);
and AND3 (N16723, N16715, N12952, N13877);
or OR3 (N16724, N16716, N5884, N12286);
xor XOR2 (N16725, N16712, N14241);
nor NOR4 (N16726, N16719, N13412, N15568, N10824);
or OR4 (N16727, N16726, N6375, N16209, N11957);
not NOT1 (N16728, N16702);
and AND3 (N16729, N16718, N12740, N14883);
not NOT1 (N16730, N16727);
nor NOR4 (N16731, N16724, N15720, N16263, N13746);
nand NAND3 (N16732, N16730, N12, N15841);
or OR3 (N16733, N16725, N14318, N6479);
not NOT1 (N16734, N16717);
or OR4 (N16735, N16721, N5653, N2948, N10351);
or OR4 (N16736, N16734, N15070, N15105, N7067);
xor XOR2 (N16737, N16733, N16048);
xor XOR2 (N16738, N16731, N13207);
not NOT1 (N16739, N16737);
and AND3 (N16740, N16728, N1620, N16643);
nor NOR3 (N16741, N16729, N14871, N13293);
not NOT1 (N16742, N16739);
buf BUF1 (N16743, N16723);
and AND2 (N16744, N16742, N13492);
buf BUF1 (N16745, N16714);
or OR2 (N16746, N16732, N4105);
nand NAND3 (N16747, N16744, N3507, N7137);
not NOT1 (N16748, N16735);
or OR3 (N16749, N16746, N5425, N14658);
and AND3 (N16750, N16736, N7771, N10419);
not NOT1 (N16751, N16749);
and AND3 (N16752, N16741, N8472, N2726);
nand NAND3 (N16753, N16738, N16074, N2043);
nor NOR4 (N16754, N16751, N13377, N7701, N7993);
or OR4 (N16755, N16752, N15994, N10711, N9145);
and AND4 (N16756, N16755, N4830, N15510, N12823);
nand NAND4 (N16757, N16745, N2100, N11987, N11977);
and AND4 (N16758, N16753, N12352, N13753, N7312);
nor NOR3 (N16759, N16754, N13974, N6983);
nor NOR3 (N16760, N16722, N7461, N12043);
buf BUF1 (N16761, N16748);
buf BUF1 (N16762, N16743);
buf BUF1 (N16763, N16757);
or OR3 (N16764, N16756, N4238, N68);
not NOT1 (N16765, N16763);
or OR3 (N16766, N16758, N7281, N5459);
nor NOR2 (N16767, N16766, N6195);
nor NOR4 (N16768, N16747, N8840, N7142, N13052);
nor NOR4 (N16769, N16760, N14643, N14568, N4692);
buf BUF1 (N16770, N16740);
and AND2 (N16771, N16761, N16611);
and AND3 (N16772, N16771, N16758, N1973);
not NOT1 (N16773, N16764);
or OR2 (N16774, N16773, N5408);
buf BUF1 (N16775, N16769);
buf BUF1 (N16776, N16759);
and AND4 (N16777, N16775, N13797, N8906, N11240);
nor NOR2 (N16778, N16750, N11862);
nand NAND3 (N16779, N16770, N16414, N7717);
not NOT1 (N16780, N16772);
xor XOR2 (N16781, N16768, N15368);
and AND2 (N16782, N16781, N14671);
xor XOR2 (N16783, N16762, N11666);
not NOT1 (N16784, N16783);
not NOT1 (N16785, N16782);
or OR2 (N16786, N16765, N15018);
nand NAND4 (N16787, N16784, N14573, N8553, N11364);
xor XOR2 (N16788, N16777, N3806);
xor XOR2 (N16789, N16776, N8071);
nor NOR4 (N16790, N16774, N3181, N10507, N10199);
and AND2 (N16791, N16785, N15301);
xor XOR2 (N16792, N16779, N9945);
xor XOR2 (N16793, N16786, N644);
xor XOR2 (N16794, N16790, N2865);
buf BUF1 (N16795, N16788);
not NOT1 (N16796, N16792);
xor XOR2 (N16797, N16778, N4176);
buf BUF1 (N16798, N16793);
not NOT1 (N16799, N16767);
nand NAND4 (N16800, N16799, N889, N14148, N8350);
and AND3 (N16801, N16798, N12558, N11024);
or OR3 (N16802, N16797, N11308, N9704);
or OR2 (N16803, N16801, N5610);
nor NOR3 (N16804, N16796, N7144, N14820);
nor NOR3 (N16805, N16780, N12598, N10528);
and AND2 (N16806, N16804, N4176);
xor XOR2 (N16807, N16806, N692);
not NOT1 (N16808, N16794);
nor NOR2 (N16809, N16789, N13761);
not NOT1 (N16810, N16809);
or OR2 (N16811, N16805, N13202);
not NOT1 (N16812, N16811);
not NOT1 (N16813, N16808);
xor XOR2 (N16814, N16802, N323);
not NOT1 (N16815, N16810);
or OR2 (N16816, N16815, N3333);
nor NOR3 (N16817, N16803, N2711, N10686);
nand NAND2 (N16818, N16814, N332);
nand NAND2 (N16819, N16800, N6330);
or OR3 (N16820, N16818, N2601, N9981);
buf BUF1 (N16821, N16787);
nand NAND3 (N16822, N16819, N10690, N683);
or OR4 (N16823, N16820, N4173, N358, N923);
nor NOR4 (N16824, N16817, N3776, N929, N7015);
xor XOR2 (N16825, N16807, N5314);
nor NOR4 (N16826, N16823, N7495, N11921, N2600);
nand NAND3 (N16827, N16812, N3947, N14486);
not NOT1 (N16828, N16821);
or OR2 (N16829, N16828, N9064);
and AND3 (N16830, N16816, N8360, N11381);
xor XOR2 (N16831, N16829, N6336);
xor XOR2 (N16832, N16826, N6856);
xor XOR2 (N16833, N16822, N7300);
or OR4 (N16834, N16824, N13440, N3913, N13149);
buf BUF1 (N16835, N16832);
nor NOR2 (N16836, N16830, N7185);
nand NAND3 (N16837, N16795, N15304, N13512);
nor NOR2 (N16838, N16831, N4529);
and AND3 (N16839, N16825, N5890, N11048);
buf BUF1 (N16840, N16833);
nand NAND3 (N16841, N16827, N8767, N14036);
nand NAND4 (N16842, N16834, N13655, N7126, N9508);
xor XOR2 (N16843, N16836, N14245);
nand NAND4 (N16844, N16791, N14615, N1995, N1470);
and AND3 (N16845, N16840, N16009, N2209);
or OR2 (N16846, N16845, N6753);
and AND4 (N16847, N16839, N15632, N10645, N7918);
xor XOR2 (N16848, N16844, N16709);
and AND4 (N16849, N16841, N4065, N11196, N7008);
or OR3 (N16850, N16843, N176, N4299);
not NOT1 (N16851, N16850);
nand NAND4 (N16852, N16813, N3986, N9164, N12036);
nand NAND4 (N16853, N16846, N14685, N8449, N7112);
not NOT1 (N16854, N16838);
xor XOR2 (N16855, N16837, N9449);
and AND3 (N16856, N16853, N15337, N11053);
nor NOR4 (N16857, N16852, N2241, N101, N6906);
buf BUF1 (N16858, N16851);
nor NOR3 (N16859, N16849, N7752, N6797);
not NOT1 (N16860, N16858);
nand NAND4 (N16861, N16855, N3500, N11677, N8769);
xor XOR2 (N16862, N16848, N10931);
xor XOR2 (N16863, N16835, N813);
and AND4 (N16864, N16854, N15477, N2134, N4048);
not NOT1 (N16865, N16861);
nor NOR3 (N16866, N16857, N5595, N6705);
nand NAND3 (N16867, N16860, N8663, N2697);
nor NOR3 (N16868, N16862, N12072, N9734);
not NOT1 (N16869, N16867);
or OR2 (N16870, N16842, N1948);
not NOT1 (N16871, N16847);
buf BUF1 (N16872, N16869);
nand NAND4 (N16873, N16863, N6455, N3724, N12149);
or OR4 (N16874, N16864, N2129, N16267, N8840);
xor XOR2 (N16875, N16856, N14971);
and AND3 (N16876, N16865, N2636, N5324);
and AND4 (N16877, N16866, N11021, N15455, N7485);
nand NAND3 (N16878, N16877, N5158, N14894);
buf BUF1 (N16879, N16878);
buf BUF1 (N16880, N16876);
nand NAND3 (N16881, N16879, N1181, N8343);
buf BUF1 (N16882, N16881);
nand NAND3 (N16883, N16870, N13976, N992);
buf BUF1 (N16884, N16882);
or OR2 (N16885, N16875, N6127);
nor NOR4 (N16886, N16874, N4884, N13122, N14615);
or OR3 (N16887, N16871, N2498, N4027);
nor NOR3 (N16888, N16859, N6071, N1297);
or OR2 (N16889, N16883, N7884);
and AND4 (N16890, N16868, N9494, N9524, N2078);
or OR2 (N16891, N16884, N16202);
buf BUF1 (N16892, N16888);
xor XOR2 (N16893, N16873, N4923);
nand NAND4 (N16894, N16890, N1336, N9410, N5775);
nand NAND3 (N16895, N16872, N14370, N6147);
nor NOR3 (N16896, N16889, N5462, N725);
or OR3 (N16897, N16894, N7146, N1767);
xor XOR2 (N16898, N16880, N3000);
not NOT1 (N16899, N16896);
nor NOR4 (N16900, N16898, N3144, N13136, N3402);
nor NOR3 (N16901, N16891, N796, N9077);
and AND2 (N16902, N16900, N3860);
xor XOR2 (N16903, N16897, N1814);
and AND3 (N16904, N16902, N10906, N2929);
buf BUF1 (N16905, N16895);
and AND2 (N16906, N16903, N10567);
not NOT1 (N16907, N16893);
nand NAND3 (N16908, N16899, N14442, N3681);
nor NOR4 (N16909, N16885, N2949, N8208, N6690);
not NOT1 (N16910, N16909);
or OR4 (N16911, N16905, N14638, N2342, N7544);
or OR2 (N16912, N16886, N5600);
not NOT1 (N16913, N16911);
or OR4 (N16914, N16887, N42, N8030, N11204);
not NOT1 (N16915, N16901);
xor XOR2 (N16916, N16892, N5302);
or OR2 (N16917, N16904, N13579);
buf BUF1 (N16918, N16914);
buf BUF1 (N16919, N16915);
xor XOR2 (N16920, N16907, N14596);
xor XOR2 (N16921, N16913, N2833);
or OR3 (N16922, N16920, N6884, N14942);
and AND4 (N16923, N16918, N12040, N11628, N15632);
xor XOR2 (N16924, N16908, N9038);
not NOT1 (N16925, N16906);
nand NAND3 (N16926, N16922, N14603, N8457);
nor NOR4 (N16927, N16919, N15242, N527, N12117);
nand NAND4 (N16928, N16923, N4937, N4523, N16260);
not NOT1 (N16929, N16924);
not NOT1 (N16930, N16916);
nand NAND2 (N16931, N16921, N15452);
and AND2 (N16932, N16928, N9660);
and AND4 (N16933, N16930, N14539, N15998, N5700);
not NOT1 (N16934, N16925);
not NOT1 (N16935, N16917);
and AND4 (N16936, N16912, N6344, N16458, N3006);
buf BUF1 (N16937, N16910);
or OR3 (N16938, N16935, N5530, N5917);
nand NAND2 (N16939, N16934, N13280);
and AND4 (N16940, N16936, N7753, N5764, N13008);
nand NAND2 (N16941, N16926, N12116);
or OR3 (N16942, N16932, N3813, N3253);
nand NAND3 (N16943, N16931, N12138, N4823);
nand NAND4 (N16944, N16941, N5522, N2268, N12445);
and AND3 (N16945, N16938, N9564, N10679);
nor NOR3 (N16946, N16943, N12675, N795);
nor NOR4 (N16947, N16937, N209, N12385, N501);
nand NAND2 (N16948, N16942, N4009);
nand NAND2 (N16949, N16940, N2709);
or OR3 (N16950, N16945, N486, N11348);
or OR4 (N16951, N16933, N13076, N13003, N6467);
not NOT1 (N16952, N16944);
and AND2 (N16953, N16948, N11779);
buf BUF1 (N16954, N16950);
buf BUF1 (N16955, N16952);
nand NAND3 (N16956, N16954, N5766, N6891);
or OR4 (N16957, N16927, N16797, N9590, N10840);
xor XOR2 (N16958, N16929, N5251);
nor NOR3 (N16959, N16958, N10827, N8353);
or OR3 (N16960, N16955, N1087, N11228);
not NOT1 (N16961, N16960);
or OR2 (N16962, N16956, N15251);
nor NOR2 (N16963, N16949, N876);
or OR2 (N16964, N16939, N2195);
and AND2 (N16965, N16946, N6705);
xor XOR2 (N16966, N16947, N4836);
buf BUF1 (N16967, N16966);
nand NAND4 (N16968, N16964, N16814, N11104, N14601);
not NOT1 (N16969, N16965);
buf BUF1 (N16970, N16961);
and AND4 (N16971, N16968, N6000, N8370, N13788);
buf BUF1 (N16972, N16957);
not NOT1 (N16973, N16971);
or OR4 (N16974, N16970, N5802, N1693, N2347);
buf BUF1 (N16975, N16967);
not NOT1 (N16976, N16962);
nor NOR3 (N16977, N16951, N10927, N696);
and AND4 (N16978, N16976, N75, N5237, N599);
xor XOR2 (N16979, N16973, N2112);
nor NOR3 (N16980, N16978, N4771, N5687);
nand NAND2 (N16981, N16977, N16532);
and AND2 (N16982, N16981, N15787);
xor XOR2 (N16983, N16959, N918);
nand NAND3 (N16984, N16974, N3590, N7928);
not NOT1 (N16985, N16969);
nor NOR3 (N16986, N16979, N2370, N4243);
nor NOR4 (N16987, N16986, N12539, N2056, N7419);
and AND2 (N16988, N16980, N11057);
nor NOR2 (N16989, N16985, N2422);
and AND3 (N16990, N16989, N3324, N1267);
or OR2 (N16991, N16975, N15768);
xor XOR2 (N16992, N16982, N10458);
nand NAND3 (N16993, N16983, N13502, N7477);
nand NAND4 (N16994, N16972, N11459, N1191, N473);
and AND2 (N16995, N16994, N13702);
and AND2 (N16996, N16988, N3711);
nor NOR4 (N16997, N16991, N12357, N11464, N1363);
not NOT1 (N16998, N16993);
not NOT1 (N16999, N16992);
xor XOR2 (N17000, N16999, N5255);
not NOT1 (N17001, N16987);
not NOT1 (N17002, N16984);
xor XOR2 (N17003, N16995, N5902);
or OR4 (N17004, N17002, N15872, N12535, N13557);
and AND3 (N17005, N17004, N625, N8065);
buf BUF1 (N17006, N17005);
nand NAND3 (N17007, N17000, N11794, N2923);
nor NOR3 (N17008, N16998, N14519, N15990);
buf BUF1 (N17009, N17008);
and AND3 (N17010, N17006, N5330, N7443);
not NOT1 (N17011, N16963);
nor NOR4 (N17012, N16990, N4259, N1651, N10161);
xor XOR2 (N17013, N17012, N15175);
nor NOR2 (N17014, N17013, N3579);
not NOT1 (N17015, N16953);
nor NOR2 (N17016, N17014, N10856);
not NOT1 (N17017, N16997);
nand NAND4 (N17018, N17015, N6722, N4871, N782);
and AND3 (N17019, N17011, N7398, N1678);
nor NOR2 (N17020, N17018, N8723);
not NOT1 (N17021, N17007);
nor NOR2 (N17022, N17019, N5584);
or OR3 (N17023, N16996, N13267, N7087);
buf BUF1 (N17024, N17016);
nor NOR4 (N17025, N17010, N11361, N4266, N9670);
xor XOR2 (N17026, N17022, N2676);
and AND4 (N17027, N17017, N6395, N4684, N8442);
nand NAND4 (N17028, N17024, N9188, N7227, N15981);
xor XOR2 (N17029, N17025, N15860);
xor XOR2 (N17030, N17026, N15831);
nor NOR3 (N17031, N17009, N4705, N13553);
buf BUF1 (N17032, N17023);
buf BUF1 (N17033, N17032);
or OR3 (N17034, N17030, N4850, N9354);
nor NOR4 (N17035, N17020, N9364, N4127, N562);
buf BUF1 (N17036, N17034);
buf BUF1 (N17037, N17021);
nand NAND4 (N17038, N17035, N16856, N8588, N14253);
nand NAND2 (N17039, N17037, N16273);
and AND4 (N17040, N17033, N3279, N254, N6887);
nand NAND2 (N17041, N17040, N730);
xor XOR2 (N17042, N17036, N6360);
nand NAND2 (N17043, N17029, N162);
not NOT1 (N17044, N17041);
not NOT1 (N17045, N17042);
buf BUF1 (N17046, N17028);
nand NAND4 (N17047, N17003, N7574, N13413, N1936);
and AND3 (N17048, N17038, N9491, N9689);
or OR4 (N17049, N17046, N9418, N1608, N15589);
nor NOR2 (N17050, N17044, N10239);
not NOT1 (N17051, N17049);
nand NAND3 (N17052, N17039, N9751, N123);
not NOT1 (N17053, N17001);
nor NOR4 (N17054, N17051, N4800, N17037, N13023);
nand NAND4 (N17055, N17054, N2248, N9177, N13438);
nor NOR2 (N17056, N17048, N7022);
xor XOR2 (N17057, N17053, N12138);
nand NAND2 (N17058, N17045, N15333);
xor XOR2 (N17059, N17056, N2265);
or OR4 (N17060, N17027, N5115, N1414, N7233);
xor XOR2 (N17061, N17057, N7918);
and AND2 (N17062, N17058, N2989);
or OR4 (N17063, N17060, N3344, N9966, N15228);
nor NOR2 (N17064, N17031, N8663);
nand NAND2 (N17065, N17052, N8766);
not NOT1 (N17066, N17064);
nor NOR3 (N17067, N17065, N4081, N14807);
xor XOR2 (N17068, N17055, N13748);
not NOT1 (N17069, N17068);
not NOT1 (N17070, N17050);
xor XOR2 (N17071, N17067, N1169);
and AND3 (N17072, N17043, N7072, N2426);
xor XOR2 (N17073, N17059, N6899);
nand NAND3 (N17074, N17062, N2367, N11929);
and AND3 (N17075, N17066, N10355, N1856);
nand NAND2 (N17076, N17071, N9761);
nand NAND4 (N17077, N17069, N3781, N13502, N3488);
nand NAND2 (N17078, N17063, N7881);
not NOT1 (N17079, N17047);
or OR4 (N17080, N17075, N8150, N10961, N12629);
nand NAND2 (N17081, N17078, N10191);
buf BUF1 (N17082, N17073);
nor NOR3 (N17083, N17079, N2491, N15154);
xor XOR2 (N17084, N17080, N7138);
and AND2 (N17085, N17074, N16858);
buf BUF1 (N17086, N17083);
nor NOR3 (N17087, N17072, N3715, N2480);
nor NOR2 (N17088, N17061, N3671);
buf BUF1 (N17089, N17081);
nor NOR2 (N17090, N17076, N13673);
not NOT1 (N17091, N17086);
and AND4 (N17092, N17084, N16514, N6254, N13089);
or OR4 (N17093, N17077, N13356, N9874, N7335);
and AND2 (N17094, N17085, N15062);
not NOT1 (N17095, N17092);
nor NOR4 (N17096, N17090, N14471, N13701, N9);
not NOT1 (N17097, N17082);
xor XOR2 (N17098, N17093, N11984);
xor XOR2 (N17099, N17087, N7705);
xor XOR2 (N17100, N17095, N6074);
buf BUF1 (N17101, N17096);
nor NOR3 (N17102, N17070, N11310, N4877);
or OR2 (N17103, N17088, N11427);
nand NAND3 (N17104, N17091, N16580, N13380);
nor NOR2 (N17105, N17102, N7442);
and AND2 (N17106, N17094, N13914);
xor XOR2 (N17107, N17100, N8647);
buf BUF1 (N17108, N17104);
buf BUF1 (N17109, N17101);
not NOT1 (N17110, N17107);
and AND4 (N17111, N17108, N3882, N1571, N5066);
xor XOR2 (N17112, N17109, N10971);
xor XOR2 (N17113, N17112, N7505);
nand NAND3 (N17114, N17089, N10777, N13861);
not NOT1 (N17115, N17111);
buf BUF1 (N17116, N17114);
or OR2 (N17117, N17116, N8385);
not NOT1 (N17118, N17113);
and AND3 (N17119, N17099, N8281, N7860);
xor XOR2 (N17120, N17117, N5765);
or OR4 (N17121, N17105, N8740, N3240, N11492);
not NOT1 (N17122, N17118);
or OR2 (N17123, N17110, N10868);
nor NOR4 (N17124, N17097, N16356, N13262, N1117);
nand NAND4 (N17125, N17122, N10613, N16659, N13425);
xor XOR2 (N17126, N17098, N10337);
buf BUF1 (N17127, N17124);
nand NAND2 (N17128, N17120, N17020);
xor XOR2 (N17129, N17121, N9678);
nor NOR4 (N17130, N17129, N11854, N7648, N12563);
not NOT1 (N17131, N17125);
xor XOR2 (N17132, N17103, N2545);
or OR2 (N17133, N17131, N17026);
not NOT1 (N17134, N17127);
nor NOR3 (N17135, N17115, N14401, N12535);
buf BUF1 (N17136, N17123);
xor XOR2 (N17137, N17128, N1068);
or OR2 (N17138, N17134, N38);
nor NOR4 (N17139, N17130, N10009, N10809, N16199);
nor NOR2 (N17140, N17132, N7748);
not NOT1 (N17141, N17135);
nor NOR3 (N17142, N17136, N14525, N12392);
not NOT1 (N17143, N17140);
xor XOR2 (N17144, N17141, N7421);
buf BUF1 (N17145, N17139);
and AND4 (N17146, N17126, N15979, N8717, N14292);
xor XOR2 (N17147, N17119, N15554);
xor XOR2 (N17148, N17142, N11907);
or OR3 (N17149, N17143, N8753, N6270);
buf BUF1 (N17150, N17147);
nand NAND2 (N17151, N17138, N4831);
not NOT1 (N17152, N17106);
or OR2 (N17153, N17148, N10162);
not NOT1 (N17154, N17152);
not NOT1 (N17155, N17145);
xor XOR2 (N17156, N17155, N6089);
or OR4 (N17157, N17133, N4022, N1305, N4318);
buf BUF1 (N17158, N17151);
nand NAND3 (N17159, N17137, N580, N16132);
nor NOR3 (N17160, N17144, N5165, N2997);
xor XOR2 (N17161, N17146, N871);
and AND2 (N17162, N17153, N8228);
and AND2 (N17163, N17159, N6746);
and AND4 (N17164, N17161, N760, N15140, N493);
nor NOR2 (N17165, N17160, N12127);
xor XOR2 (N17166, N17165, N13422);
nor NOR4 (N17167, N17154, N8055, N6214, N3374);
not NOT1 (N17168, N17157);
not NOT1 (N17169, N17167);
not NOT1 (N17170, N17149);
nor NOR4 (N17171, N17164, N9744, N2109, N7925);
xor XOR2 (N17172, N17168, N13252);
nor NOR3 (N17173, N17162, N13928, N12900);
or OR2 (N17174, N17150, N7731);
xor XOR2 (N17175, N17172, N6969);
or OR4 (N17176, N17169, N3786, N2401, N8542);
nor NOR3 (N17177, N17158, N9090, N3714);
not NOT1 (N17178, N17177);
xor XOR2 (N17179, N17174, N13079);
and AND2 (N17180, N17179, N16026);
not NOT1 (N17181, N17156);
nor NOR4 (N17182, N17170, N13211, N15493, N15356);
or OR4 (N17183, N17166, N11434, N9362, N12425);
or OR4 (N17184, N17180, N10071, N15041, N15672);
xor XOR2 (N17185, N17163, N5888);
or OR2 (N17186, N17182, N6310);
or OR3 (N17187, N17181, N6032, N16110);
or OR2 (N17188, N17171, N15860);
nor NOR3 (N17189, N17186, N11985, N10666);
and AND4 (N17190, N17184, N12823, N4029, N7798);
xor XOR2 (N17191, N17188, N8643);
and AND2 (N17192, N17187, N4939);
and AND3 (N17193, N17176, N16410, N15584);
or OR2 (N17194, N17175, N7873);
nor NOR2 (N17195, N17189, N1026);
xor XOR2 (N17196, N17190, N1808);
buf BUF1 (N17197, N17173);
nand NAND2 (N17198, N17185, N16820);
nand NAND2 (N17199, N17193, N14482);
buf BUF1 (N17200, N17192);
not NOT1 (N17201, N17197);
buf BUF1 (N17202, N17196);
nor NOR3 (N17203, N17194, N14226, N12391);
buf BUF1 (N17204, N17202);
nor NOR2 (N17205, N17183, N12302);
buf BUF1 (N17206, N17203);
xor XOR2 (N17207, N17205, N2459);
or OR2 (N17208, N17204, N5038);
buf BUF1 (N17209, N17200);
buf BUF1 (N17210, N17198);
buf BUF1 (N17211, N17210);
xor XOR2 (N17212, N17195, N549);
buf BUF1 (N17213, N17207);
buf BUF1 (N17214, N17199);
nand NAND3 (N17215, N17213, N11303, N7528);
xor XOR2 (N17216, N17212, N5700);
nand NAND2 (N17217, N17206, N6952);
not NOT1 (N17218, N17215);
nor NOR3 (N17219, N17218, N13359, N14152);
not NOT1 (N17220, N17201);
nor NOR3 (N17221, N17209, N9023, N12175);
not NOT1 (N17222, N17178);
buf BUF1 (N17223, N17214);
buf BUF1 (N17224, N17216);
nor NOR2 (N17225, N17222, N12031);
and AND3 (N17226, N17219, N5866, N2240);
nor NOR2 (N17227, N17217, N16100);
or OR3 (N17228, N17225, N14792, N3332);
nor NOR3 (N17229, N17223, N4373, N6222);
buf BUF1 (N17230, N17221);
not NOT1 (N17231, N17208);
buf BUF1 (N17232, N17227);
not NOT1 (N17233, N17230);
or OR3 (N17234, N17231, N16201, N8709);
nand NAND4 (N17235, N17224, N14744, N435, N6192);
nor NOR2 (N17236, N17235, N15432);
or OR3 (N17237, N17228, N8760, N10118);
or OR4 (N17238, N17233, N5453, N14260, N5487);
buf BUF1 (N17239, N17220);
buf BUF1 (N17240, N17191);
xor XOR2 (N17241, N17239, N3052);
nand NAND2 (N17242, N17236, N16169);
nor NOR2 (N17243, N17241, N2683);
nand NAND2 (N17244, N17211, N8433);
nor NOR4 (N17245, N17234, N14085, N12676, N3145);
and AND3 (N17246, N17229, N6858, N6612);
buf BUF1 (N17247, N17243);
not NOT1 (N17248, N17232);
and AND3 (N17249, N17226, N12839, N9512);
xor XOR2 (N17250, N17249, N5885);
nand NAND2 (N17251, N17238, N2909);
nor NOR4 (N17252, N17246, N7344, N15995, N4984);
not NOT1 (N17253, N17240);
nand NAND2 (N17254, N17252, N407);
buf BUF1 (N17255, N17244);
nand NAND3 (N17256, N17255, N4671, N15380);
or OR4 (N17257, N17237, N12669, N3078, N14777);
and AND4 (N17258, N17257, N6627, N17086, N1174);
or OR3 (N17259, N17247, N2170, N15453);
or OR3 (N17260, N17242, N10342, N11677);
xor XOR2 (N17261, N17259, N4163);
nand NAND4 (N17262, N17245, N8004, N11384, N16266);
nand NAND4 (N17263, N17262, N4810, N8939, N14648);
buf BUF1 (N17264, N17261);
or OR2 (N17265, N17264, N6461);
or OR3 (N17266, N17251, N9722, N12051);
or OR3 (N17267, N17248, N5954, N1173);
nand NAND3 (N17268, N17260, N13631, N11114);
nor NOR3 (N17269, N17258, N16211, N16589);
and AND2 (N17270, N17265, N14661);
nand NAND2 (N17271, N17253, N3036);
not NOT1 (N17272, N17256);
not NOT1 (N17273, N17254);
not NOT1 (N17274, N17271);
nand NAND4 (N17275, N17266, N9503, N11842, N7558);
xor XOR2 (N17276, N17275, N11055);
not NOT1 (N17277, N17273);
nand NAND4 (N17278, N17272, N14573, N8640, N6929);
and AND2 (N17279, N17270, N1917);
or OR3 (N17280, N17250, N13057, N13704);
or OR3 (N17281, N17279, N13227, N12459);
xor XOR2 (N17282, N17278, N16344);
or OR2 (N17283, N17282, N17075);
or OR3 (N17284, N17283, N10845, N14823);
nand NAND3 (N17285, N17267, N7035, N15395);
and AND3 (N17286, N17281, N4834, N14504);
nand NAND2 (N17287, N17284, N10743);
xor XOR2 (N17288, N17269, N15342);
or OR3 (N17289, N17288, N8252, N12822);
not NOT1 (N17290, N17285);
not NOT1 (N17291, N17274);
nand NAND3 (N17292, N17287, N14172, N7537);
xor XOR2 (N17293, N17286, N5054);
not NOT1 (N17294, N17292);
buf BUF1 (N17295, N17277);
not NOT1 (N17296, N17290);
xor XOR2 (N17297, N17294, N14802);
nor NOR3 (N17298, N17289, N15155, N318);
nor NOR4 (N17299, N17298, N1392, N7559, N10686);
buf BUF1 (N17300, N17293);
and AND4 (N17301, N17299, N8468, N12500, N10334);
xor XOR2 (N17302, N17268, N10874);
buf BUF1 (N17303, N17295);
xor XOR2 (N17304, N17303, N2673);
buf BUF1 (N17305, N17280);
buf BUF1 (N17306, N17263);
xor XOR2 (N17307, N17300, N13463);
xor XOR2 (N17308, N17297, N6134);
nor NOR2 (N17309, N17301, N597);
and AND3 (N17310, N17306, N13266, N4051);
and AND3 (N17311, N17309, N4373, N7171);
xor XOR2 (N17312, N17311, N601);
not NOT1 (N17313, N17291);
and AND4 (N17314, N17276, N5485, N13969, N9996);
nor NOR4 (N17315, N17310, N7371, N6010, N708);
not NOT1 (N17316, N17313);
nor NOR3 (N17317, N17304, N7531, N16930);
nor NOR3 (N17318, N17296, N1306, N2101);
xor XOR2 (N17319, N17308, N12258);
xor XOR2 (N17320, N17317, N17020);
or OR2 (N17321, N17315, N2396);
and AND3 (N17322, N17302, N8387, N5284);
nand NAND4 (N17323, N17314, N3831, N14021, N11782);
buf BUF1 (N17324, N17305);
nor NOR4 (N17325, N17316, N16646, N5401, N13660);
xor XOR2 (N17326, N17325, N9450);
and AND3 (N17327, N17322, N2164, N177);
and AND2 (N17328, N17327, N16924);
nand NAND3 (N17329, N17312, N2711, N11919);
not NOT1 (N17330, N17328);
or OR4 (N17331, N17330, N16766, N13280, N16996);
not NOT1 (N17332, N17324);
nor NOR2 (N17333, N17321, N3314);
nand NAND3 (N17334, N17307, N1168, N15058);
buf BUF1 (N17335, N17334);
and AND4 (N17336, N17320, N6993, N1941, N14464);
nand NAND3 (N17337, N17335, N9664, N14846);
xor XOR2 (N17338, N17318, N1980);
xor XOR2 (N17339, N17332, N9398);
and AND3 (N17340, N17326, N14189, N7741);
and AND3 (N17341, N17323, N17233, N3887);
nor NOR4 (N17342, N17331, N8828, N4271, N7620);
nand NAND3 (N17343, N17337, N13293, N15904);
not NOT1 (N17344, N17341);
buf BUF1 (N17345, N17340);
not NOT1 (N17346, N17344);
and AND3 (N17347, N17346, N2047, N7395);
not NOT1 (N17348, N17345);
or OR3 (N17349, N17319, N7758, N2802);
or OR2 (N17350, N17347, N6776);
nor NOR4 (N17351, N17336, N6934, N9777, N1741);
nor NOR3 (N17352, N17342, N154, N7747);
xor XOR2 (N17353, N17338, N11972);
buf BUF1 (N17354, N17333);
xor XOR2 (N17355, N17343, N3314);
nor NOR3 (N17356, N17354, N1807, N716);
not NOT1 (N17357, N17355);
and AND2 (N17358, N17352, N15485);
or OR2 (N17359, N17351, N5837);
not NOT1 (N17360, N17357);
not NOT1 (N17361, N17339);
nand NAND2 (N17362, N17348, N17266);
and AND4 (N17363, N17360, N5521, N6545, N14899);
nor NOR2 (N17364, N17361, N7743);
and AND3 (N17365, N17362, N15063, N1667);
or OR4 (N17366, N17359, N14682, N12018, N15997);
xor XOR2 (N17367, N17366, N62);
and AND2 (N17368, N17353, N4795);
nand NAND4 (N17369, N17350, N14416, N8269, N3834);
or OR2 (N17370, N17358, N6402);
buf BUF1 (N17371, N17329);
nand NAND4 (N17372, N17367, N13603, N5608, N12960);
buf BUF1 (N17373, N17371);
and AND3 (N17374, N17370, N14567, N10892);
or OR3 (N17375, N17368, N15358, N7229);
and AND3 (N17376, N17375, N6543, N9474);
and AND3 (N17377, N17373, N10879, N5616);
buf BUF1 (N17378, N17376);
not NOT1 (N17379, N17377);
and AND3 (N17380, N17372, N14341, N6912);
buf BUF1 (N17381, N17365);
buf BUF1 (N17382, N17349);
nor NOR3 (N17383, N17374, N12348, N16862);
xor XOR2 (N17384, N17381, N3092);
nand NAND2 (N17385, N17363, N1614);
or OR2 (N17386, N17385, N8299);
nor NOR2 (N17387, N17384, N1747);
xor XOR2 (N17388, N17386, N7831);
buf BUF1 (N17389, N17380);
nand NAND3 (N17390, N17388, N8988, N8450);
xor XOR2 (N17391, N17382, N8240);
buf BUF1 (N17392, N17364);
nand NAND3 (N17393, N17390, N14702, N12784);
xor XOR2 (N17394, N17356, N11572);
or OR3 (N17395, N17379, N15437, N18);
buf BUF1 (N17396, N17392);
buf BUF1 (N17397, N17395);
buf BUF1 (N17398, N17396);
buf BUF1 (N17399, N17378);
buf BUF1 (N17400, N17399);
or OR3 (N17401, N17383, N10097, N437);
or OR3 (N17402, N17391, N6753, N5640);
nor NOR4 (N17403, N17402, N16693, N10503, N3224);
not NOT1 (N17404, N17393);
not NOT1 (N17405, N17398);
buf BUF1 (N17406, N17401);
buf BUF1 (N17407, N17405);
buf BUF1 (N17408, N17407);
xor XOR2 (N17409, N17404, N176);
nand NAND4 (N17410, N17409, N9142, N9593, N7145);
buf BUF1 (N17411, N17400);
xor XOR2 (N17412, N17410, N1980);
xor XOR2 (N17413, N17408, N10364);
buf BUF1 (N17414, N17412);
nand NAND2 (N17415, N17369, N489);
nand NAND2 (N17416, N17387, N15668);
and AND3 (N17417, N17406, N5644, N16428);
xor XOR2 (N17418, N17411, N13186);
nand NAND3 (N17419, N17389, N10204, N13260);
nor NOR3 (N17420, N17416, N3524, N6193);
or OR2 (N17421, N17415, N16000);
buf BUF1 (N17422, N17419);
or OR2 (N17423, N17417, N9749);
or OR4 (N17424, N17418, N8717, N15624, N7721);
or OR4 (N17425, N17421, N3228, N1071, N15065);
not NOT1 (N17426, N17420);
not NOT1 (N17427, N17414);
nand NAND2 (N17428, N17427, N14906);
not NOT1 (N17429, N17428);
or OR2 (N17430, N17403, N1886);
buf BUF1 (N17431, N17413);
or OR2 (N17432, N17425, N2941);
nor NOR4 (N17433, N17430, N4778, N16492, N14227);
nor NOR2 (N17434, N17429, N16290);
xor XOR2 (N17435, N17424, N9022);
buf BUF1 (N17436, N17433);
or OR4 (N17437, N17434, N12331, N3569, N199);
nor NOR2 (N17438, N17397, N10834);
not NOT1 (N17439, N17438);
buf BUF1 (N17440, N17423);
xor XOR2 (N17441, N17394, N7132);
buf BUF1 (N17442, N17439);
xor XOR2 (N17443, N17422, N14781);
or OR4 (N17444, N17440, N7727, N9089, N12895);
nand NAND2 (N17445, N17432, N4108);
nand NAND2 (N17446, N17436, N11007);
buf BUF1 (N17447, N17443);
or OR2 (N17448, N17444, N15033);
or OR2 (N17449, N17442, N9099);
xor XOR2 (N17450, N17446, N13762);
nor NOR4 (N17451, N17437, N13239, N1340, N1444);
nor NOR3 (N17452, N17450, N12639, N11016);
buf BUF1 (N17453, N17426);
and AND4 (N17454, N17448, N6895, N11422, N14506);
or OR2 (N17455, N17453, N14424);
buf BUF1 (N17456, N17435);
nor NOR4 (N17457, N17452, N16733, N2357, N3239);
and AND3 (N17458, N17451, N1248, N2750);
xor XOR2 (N17459, N17447, N3524);
buf BUF1 (N17460, N17445);
and AND2 (N17461, N17431, N2068);
xor XOR2 (N17462, N17449, N1736);
buf BUF1 (N17463, N17441);
or OR3 (N17464, N17458, N6790, N151);
nor NOR2 (N17465, N17462, N6776);
nand NAND2 (N17466, N17464, N13375);
xor XOR2 (N17467, N17465, N17320);
buf BUF1 (N17468, N17466);
xor XOR2 (N17469, N17454, N4221);
nor NOR4 (N17470, N17459, N1686, N9933, N14688);
not NOT1 (N17471, N17467);
buf BUF1 (N17472, N17469);
and AND3 (N17473, N17455, N1786, N10608);
buf BUF1 (N17474, N17463);
nand NAND2 (N17475, N17461, N1760);
buf BUF1 (N17476, N17470);
or OR4 (N17477, N17474, N15383, N17354, N3819);
nand NAND4 (N17478, N17460, N9839, N8773, N4146);
xor XOR2 (N17479, N17457, N2513);
xor XOR2 (N17480, N17468, N11415);
nand NAND4 (N17481, N17471, N12804, N17278, N7156);
xor XOR2 (N17482, N17477, N3001);
xor XOR2 (N17483, N17481, N9810);
buf BUF1 (N17484, N17478);
buf BUF1 (N17485, N17473);
or OR3 (N17486, N17476, N9859, N2930);
buf BUF1 (N17487, N17472);
or OR3 (N17488, N17484, N15888, N1561);
buf BUF1 (N17489, N17488);
buf BUF1 (N17490, N17487);
or OR3 (N17491, N17479, N17434, N14299);
or OR4 (N17492, N17490, N16356, N13015, N16115);
nand NAND2 (N17493, N17480, N8010);
xor XOR2 (N17494, N17486, N23);
nand NAND4 (N17495, N17493, N8123, N8475, N7875);
xor XOR2 (N17496, N17494, N3167);
or OR3 (N17497, N17456, N17438, N11792);
and AND3 (N17498, N17485, N13883, N14149);
or OR2 (N17499, N17492, N16412);
nand NAND3 (N17500, N17499, N5613, N2394);
or OR3 (N17501, N17491, N4456, N14968);
nand NAND4 (N17502, N17498, N4474, N5569, N3843);
xor XOR2 (N17503, N17501, N4778);
buf BUF1 (N17504, N17483);
nand NAND3 (N17505, N17500, N7279, N5326);
and AND4 (N17506, N17489, N9937, N8278, N15987);
not NOT1 (N17507, N17495);
xor XOR2 (N17508, N17504, N10484);
or OR2 (N17509, N17497, N7366);
xor XOR2 (N17510, N17508, N7101);
or OR4 (N17511, N17475, N2850, N4268, N1791);
nand NAND3 (N17512, N17511, N3150, N13675);
nor NOR2 (N17513, N17482, N2083);
xor XOR2 (N17514, N17513, N14941);
and AND3 (N17515, N17506, N4356, N10966);
nor NOR3 (N17516, N17503, N9524, N4468);
buf BUF1 (N17517, N17507);
not NOT1 (N17518, N17510);
and AND3 (N17519, N17516, N10560, N213);
or OR4 (N17520, N17502, N4451, N5544, N15483);
nand NAND4 (N17521, N17514, N16463, N12651, N1767);
or OR3 (N17522, N17521, N8391, N14891);
or OR3 (N17523, N17522, N16746, N3216);
xor XOR2 (N17524, N17505, N5881);
nand NAND2 (N17525, N17512, N800);
nor NOR4 (N17526, N17496, N13245, N8071, N3812);
nand NAND3 (N17527, N17526, N4058, N10234);
and AND3 (N17528, N17525, N3703, N6842);
nor NOR2 (N17529, N17523, N5421);
xor XOR2 (N17530, N17529, N15067);
xor XOR2 (N17531, N17517, N6426);
buf BUF1 (N17532, N17519);
or OR2 (N17533, N17528, N17403);
buf BUF1 (N17534, N17530);
nor NOR4 (N17535, N17532, N9207, N7853, N6187);
nand NAND2 (N17536, N17534, N11758);
buf BUF1 (N17537, N17527);
buf BUF1 (N17538, N17531);
or OR2 (N17539, N17509, N5046);
xor XOR2 (N17540, N17539, N10361);
nand NAND3 (N17541, N17535, N4895, N1523);
xor XOR2 (N17542, N17540, N11720);
or OR3 (N17543, N17524, N17311, N1455);
and AND3 (N17544, N17533, N13324, N1338);
or OR3 (N17545, N17537, N14372, N1183);
or OR4 (N17546, N17515, N13736, N10302, N5960);
xor XOR2 (N17547, N17546, N15982);
or OR2 (N17548, N17520, N17060);
or OR2 (N17549, N17541, N13448);
buf BUF1 (N17550, N17538);
buf BUF1 (N17551, N17550);
and AND3 (N17552, N17518, N7099, N14788);
xor XOR2 (N17553, N17543, N7002);
or OR3 (N17554, N17553, N3969, N6574);
xor XOR2 (N17555, N17536, N4514);
nand NAND4 (N17556, N17552, N7265, N11920, N8813);
nand NAND4 (N17557, N17555, N9954, N13565, N7456);
nor NOR2 (N17558, N17557, N15019);
buf BUF1 (N17559, N17558);
nor NOR4 (N17560, N17551, N835, N3593, N13908);
xor XOR2 (N17561, N17547, N6553);
nand NAND2 (N17562, N17554, N7777);
or OR3 (N17563, N17549, N5754, N10203);
buf BUF1 (N17564, N17559);
nand NAND4 (N17565, N17564, N7461, N12569, N6676);
nor NOR4 (N17566, N17544, N14625, N11886, N11215);
xor XOR2 (N17567, N17560, N16837);
or OR4 (N17568, N17561, N13347, N3077, N1192);
nor NOR2 (N17569, N17556, N13152);
xor XOR2 (N17570, N17565, N5104);
nor NOR2 (N17571, N17568, N11101);
xor XOR2 (N17572, N17542, N10566);
buf BUF1 (N17573, N17562);
and AND4 (N17574, N17569, N14417, N12870, N12272);
not NOT1 (N17575, N17545);
not NOT1 (N17576, N17548);
not NOT1 (N17577, N17573);
buf BUF1 (N17578, N17571);
and AND2 (N17579, N17574, N17302);
nor NOR2 (N17580, N17579, N4285);
or OR4 (N17581, N17576, N2459, N11841, N17212);
and AND3 (N17582, N17575, N13746, N6967);
or OR2 (N17583, N17572, N5663);
buf BUF1 (N17584, N17578);
buf BUF1 (N17585, N17577);
buf BUF1 (N17586, N17566);
or OR4 (N17587, N17586, N6632, N7270, N17161);
buf BUF1 (N17588, N17587);
nand NAND3 (N17589, N17580, N11494, N12122);
nand NAND3 (N17590, N17582, N8978, N13112);
nor NOR3 (N17591, N17563, N16055, N5269);
not NOT1 (N17592, N17590);
and AND4 (N17593, N17585, N17550, N2719, N2390);
nor NOR4 (N17594, N17588, N6629, N11439, N795);
and AND3 (N17595, N17593, N16737, N905);
or OR3 (N17596, N17581, N1526, N13678);
not NOT1 (N17597, N17589);
xor XOR2 (N17598, N17597, N4732);
nand NAND4 (N17599, N17598, N9003, N2409, N8956);
nor NOR4 (N17600, N17599, N17173, N833, N12470);
not NOT1 (N17601, N17596);
not NOT1 (N17602, N17567);
xor XOR2 (N17603, N17570, N1312);
buf BUF1 (N17604, N17583);
buf BUF1 (N17605, N17604);
or OR4 (N17606, N17600, N11812, N7882, N14327);
buf BUF1 (N17607, N17591);
nand NAND4 (N17608, N17602, N8067, N17454, N10027);
nand NAND3 (N17609, N17608, N10019, N17059);
and AND4 (N17610, N17601, N16101, N13586, N8086);
nand NAND4 (N17611, N17592, N2580, N5520, N3197);
or OR3 (N17612, N17611, N15713, N8499);
or OR3 (N17613, N17603, N3641, N11207);
and AND4 (N17614, N17612, N3204, N13460, N5638);
xor XOR2 (N17615, N17584, N13401);
and AND3 (N17616, N17615, N3611, N8901);
nand NAND2 (N17617, N17616, N13205);
or OR2 (N17618, N17606, N6088);
or OR4 (N17619, N17594, N3276, N14973, N2977);
not NOT1 (N17620, N17614);
nor NOR2 (N17621, N17605, N14385);
buf BUF1 (N17622, N17607);
not NOT1 (N17623, N17595);
buf BUF1 (N17624, N17621);
or OR4 (N17625, N17624, N10499, N13381, N11270);
buf BUF1 (N17626, N17625);
not NOT1 (N17627, N17620);
buf BUF1 (N17628, N17617);
buf BUF1 (N17629, N17623);
nor NOR2 (N17630, N17629, N2337);
or OR3 (N17631, N17628, N10801, N12920);
nand NAND3 (N17632, N17618, N1678, N3325);
or OR2 (N17633, N17622, N8628);
buf BUF1 (N17634, N17626);
or OR3 (N17635, N17613, N8266, N7551);
xor XOR2 (N17636, N17632, N3801);
buf BUF1 (N17637, N17633);
or OR2 (N17638, N17619, N6814);
nand NAND4 (N17639, N17637, N16177, N8476, N11279);
not NOT1 (N17640, N17639);
nor NOR2 (N17641, N17627, N17287);
or OR3 (N17642, N17634, N11301, N2750);
xor XOR2 (N17643, N17635, N15390);
or OR2 (N17644, N17642, N5636);
nor NOR2 (N17645, N17636, N16046);
and AND3 (N17646, N17609, N623, N16381);
nor NOR2 (N17647, N17610, N16578);
nor NOR3 (N17648, N17640, N12453, N13792);
nand NAND3 (N17649, N17643, N12208, N16849);
xor XOR2 (N17650, N17645, N15506);
nor NOR3 (N17651, N17647, N7713, N3635);
and AND3 (N17652, N17646, N7502, N11164);
nor NOR2 (N17653, N17641, N17362);
nor NOR3 (N17654, N17638, N4999, N9987);
buf BUF1 (N17655, N17649);
not NOT1 (N17656, N17648);
or OR3 (N17657, N17631, N12329, N3227);
or OR4 (N17658, N17654, N9606, N308, N10245);
buf BUF1 (N17659, N17656);
xor XOR2 (N17660, N17658, N10645);
xor XOR2 (N17661, N17653, N4431);
not NOT1 (N17662, N17660);
buf BUF1 (N17663, N17657);
not NOT1 (N17664, N17630);
nand NAND2 (N17665, N17655, N14175);
and AND2 (N17666, N17665, N2987);
xor XOR2 (N17667, N17644, N2478);
nand NAND2 (N17668, N17659, N2728);
nor NOR3 (N17669, N17650, N10851, N7804);
buf BUF1 (N17670, N17663);
buf BUF1 (N17671, N17667);
and AND4 (N17672, N17669, N978, N3711, N13017);
and AND3 (N17673, N17670, N14732, N4114);
buf BUF1 (N17674, N17666);
or OR2 (N17675, N17668, N14216);
xor XOR2 (N17676, N17671, N2686);
buf BUF1 (N17677, N17672);
nor NOR2 (N17678, N17661, N5552);
xor XOR2 (N17679, N17678, N73);
buf BUF1 (N17680, N17675);
and AND3 (N17681, N17662, N8055, N14097);
not NOT1 (N17682, N17681);
nand NAND3 (N17683, N17664, N15487, N13731);
xor XOR2 (N17684, N17683, N13339);
nor NOR2 (N17685, N17684, N11494);
buf BUF1 (N17686, N17682);
and AND2 (N17687, N17677, N172);
nor NOR2 (N17688, N17673, N4182);
or OR2 (N17689, N17674, N9031);
buf BUF1 (N17690, N17687);
and AND2 (N17691, N17690, N4903);
buf BUF1 (N17692, N17688);
xor XOR2 (N17693, N17652, N4518);
not NOT1 (N17694, N17686);
or OR3 (N17695, N17689, N14812, N15018);
xor XOR2 (N17696, N17694, N2123);
and AND4 (N17697, N17685, N16209, N4783, N6487);
and AND2 (N17698, N17697, N12913);
or OR3 (N17699, N17680, N8687, N10575);
buf BUF1 (N17700, N17676);
not NOT1 (N17701, N17693);
buf BUF1 (N17702, N17701);
xor XOR2 (N17703, N17696, N17090);
nor NOR4 (N17704, N17702, N1586, N1637, N8969);
and AND3 (N17705, N17698, N14187, N3789);
buf BUF1 (N17706, N17699);
buf BUF1 (N17707, N17679);
buf BUF1 (N17708, N17707);
buf BUF1 (N17709, N17692);
or OR3 (N17710, N17709, N10532, N15676);
not NOT1 (N17711, N17706);
or OR2 (N17712, N17708, N11041);
or OR4 (N17713, N17691, N6521, N4865, N14033);
not NOT1 (N17714, N17711);
or OR4 (N17715, N17695, N15599, N6995, N4435);
or OR2 (N17716, N17704, N10825);
and AND4 (N17717, N17710, N806, N12302, N13569);
buf BUF1 (N17718, N17705);
and AND2 (N17719, N17717, N9818);
nor NOR3 (N17720, N17712, N8982, N1136);
not NOT1 (N17721, N17716);
nand NAND4 (N17722, N17718, N1278, N942, N14844);
not NOT1 (N17723, N17700);
and AND2 (N17724, N17715, N5552);
or OR2 (N17725, N17720, N16300);
nand NAND3 (N17726, N17723, N7673, N6580);
not NOT1 (N17727, N17713);
nand NAND2 (N17728, N17724, N12950);
buf BUF1 (N17729, N17725);
and AND4 (N17730, N17719, N16817, N15336, N8928);
or OR4 (N17731, N17728, N6829, N7748, N9692);
and AND4 (N17732, N17731, N1375, N14806, N1111);
buf BUF1 (N17733, N17732);
nand NAND4 (N17734, N17733, N16219, N5356, N14809);
and AND3 (N17735, N17703, N7158, N15194);
and AND2 (N17736, N17721, N6829);
xor XOR2 (N17737, N17736, N5202);
or OR2 (N17738, N17714, N3614);
not NOT1 (N17739, N17735);
or OR3 (N17740, N17734, N1095, N1226);
nand NAND4 (N17741, N17726, N5812, N6854, N3933);
nand NAND3 (N17742, N17737, N13087, N9440);
or OR4 (N17743, N17727, N10128, N9780, N3077);
nand NAND4 (N17744, N17739, N5190, N4507, N4504);
not NOT1 (N17745, N17738);
and AND4 (N17746, N17729, N12092, N8247, N10775);
xor XOR2 (N17747, N17741, N8986);
or OR3 (N17748, N17744, N6566, N4512);
nand NAND2 (N17749, N17743, N15518);
buf BUF1 (N17750, N17747);
buf BUF1 (N17751, N17651);
xor XOR2 (N17752, N17742, N13159);
nand NAND2 (N17753, N17748, N130);
buf BUF1 (N17754, N17740);
nand NAND3 (N17755, N17730, N16344, N4322);
nand NAND2 (N17756, N17746, N7280);
or OR2 (N17757, N17752, N16411);
xor XOR2 (N17758, N17754, N5459);
nor NOR3 (N17759, N17751, N16131, N12057);
nor NOR3 (N17760, N17749, N8003, N3529);
not NOT1 (N17761, N17750);
buf BUF1 (N17762, N17758);
nand NAND4 (N17763, N17755, N14594, N3634, N944);
buf BUF1 (N17764, N17759);
buf BUF1 (N17765, N17756);
and AND3 (N17766, N17760, N2030, N15916);
buf BUF1 (N17767, N17753);
or OR4 (N17768, N17722, N15508, N11169, N12919);
nor NOR4 (N17769, N17768, N14809, N12480, N9033);
nand NAND2 (N17770, N17769, N7146);
nor NOR3 (N17771, N17757, N10214, N7159);
and AND3 (N17772, N17765, N10143, N16003);
nor NOR4 (N17773, N17745, N9410, N5396, N915);
buf BUF1 (N17774, N17770);
nand NAND4 (N17775, N17766, N17144, N8693, N11406);
nand NAND4 (N17776, N17774, N5821, N10072, N15951);
buf BUF1 (N17777, N17771);
xor XOR2 (N17778, N17775, N1459);
not NOT1 (N17779, N17761);
not NOT1 (N17780, N17773);
buf BUF1 (N17781, N17776);
buf BUF1 (N17782, N17764);
not NOT1 (N17783, N17779);
or OR2 (N17784, N17782, N10780);
buf BUF1 (N17785, N17763);
buf BUF1 (N17786, N17785);
buf BUF1 (N17787, N17762);
not NOT1 (N17788, N17767);
and AND3 (N17789, N17788, N12259, N10493);
buf BUF1 (N17790, N17783);
not NOT1 (N17791, N17784);
xor XOR2 (N17792, N17789, N12638);
buf BUF1 (N17793, N17790);
or OR3 (N17794, N17792, N11645, N8673);
buf BUF1 (N17795, N17781);
or OR3 (N17796, N17793, N4998, N11545);
xor XOR2 (N17797, N17786, N6199);
nand NAND4 (N17798, N17794, N16613, N12485, N17265);
nand NAND3 (N17799, N17777, N13149, N6423);
buf BUF1 (N17800, N17791);
or OR3 (N17801, N17780, N11857, N6137);
nor NOR4 (N17802, N17795, N2520, N10266, N16172);
not NOT1 (N17803, N17797);
or OR4 (N17804, N17803, N12550, N8960, N15676);
buf BUF1 (N17805, N17804);
nand NAND2 (N17806, N17778, N5798);
nand NAND3 (N17807, N17806, N5567, N730);
nor NOR3 (N17808, N17802, N7834, N3040);
buf BUF1 (N17809, N17787);
or OR4 (N17810, N17808, N15821, N4765, N9285);
or OR3 (N17811, N17772, N8414, N4614);
xor XOR2 (N17812, N17805, N1774);
buf BUF1 (N17813, N17810);
and AND3 (N17814, N17799, N11985, N10988);
buf BUF1 (N17815, N17812);
and AND3 (N17816, N17809, N11707, N15634);
not NOT1 (N17817, N17815);
nand NAND4 (N17818, N17811, N17332, N6201, N1008);
not NOT1 (N17819, N17817);
not NOT1 (N17820, N17816);
buf BUF1 (N17821, N17820);
buf BUF1 (N17822, N17800);
nand NAND2 (N17823, N17801, N8481);
nand NAND2 (N17824, N17807, N16288);
xor XOR2 (N17825, N17819, N16850);
buf BUF1 (N17826, N17796);
and AND3 (N17827, N17798, N8610, N2281);
or OR3 (N17828, N17814, N14129, N5071);
buf BUF1 (N17829, N17828);
buf BUF1 (N17830, N17826);
not NOT1 (N17831, N17829);
xor XOR2 (N17832, N17813, N17051);
or OR3 (N17833, N17825, N10374, N11638);
nor NOR4 (N17834, N17821, N10155, N17792, N1501);
or OR3 (N17835, N17834, N11744, N5272);
or OR3 (N17836, N17830, N9031, N17630);
buf BUF1 (N17837, N17818);
nor NOR2 (N17838, N17831, N2930);
xor XOR2 (N17839, N17837, N6826);
nor NOR3 (N17840, N17838, N6202, N15494);
nor NOR4 (N17841, N17823, N7384, N13305, N5325);
and AND2 (N17842, N17822, N14316);
xor XOR2 (N17843, N17842, N3819);
nor NOR2 (N17844, N17839, N14342);
or OR3 (N17845, N17832, N1301, N8118);
and AND4 (N17846, N17840, N6262, N15055, N11083);
and AND3 (N17847, N17835, N12470, N6453);
xor XOR2 (N17848, N17827, N1090);
or OR3 (N17849, N17845, N3986, N11910);
and AND4 (N17850, N17836, N337, N10130, N16007);
and AND2 (N17851, N17849, N6453);
buf BUF1 (N17852, N17841);
or OR4 (N17853, N17844, N7210, N1493, N823);
xor XOR2 (N17854, N17824, N9050);
and AND3 (N17855, N17846, N15122, N15536);
nor NOR2 (N17856, N17851, N6996);
or OR2 (N17857, N17854, N3309);
xor XOR2 (N17858, N17833, N15549);
xor XOR2 (N17859, N17847, N7040);
nor NOR2 (N17860, N17852, N5346);
nor NOR3 (N17861, N17850, N8980, N16361);
nand NAND2 (N17862, N17853, N3172);
buf BUF1 (N17863, N17857);
buf BUF1 (N17864, N17861);
nand NAND4 (N17865, N17859, N3083, N338, N7186);
nor NOR4 (N17866, N17864, N2436, N13024, N2398);
not NOT1 (N17867, N17863);
nor NOR2 (N17868, N17860, N9798);
nand NAND2 (N17869, N17856, N13700);
xor XOR2 (N17870, N17843, N8084);
or OR2 (N17871, N17868, N6160);
xor XOR2 (N17872, N17848, N14840);
and AND2 (N17873, N17862, N16539);
not NOT1 (N17874, N17865);
and AND2 (N17875, N17871, N2844);
not NOT1 (N17876, N17873);
nor NOR3 (N17877, N17866, N15373, N7805);
and AND2 (N17878, N17872, N13734);
and AND3 (N17879, N17855, N9204, N9727);
nand NAND3 (N17880, N17878, N7004, N3836);
nor NOR4 (N17881, N17879, N7051, N12679, N5980);
buf BUF1 (N17882, N17867);
nor NOR2 (N17883, N17881, N12750);
and AND3 (N17884, N17882, N8197, N17463);
or OR2 (N17885, N17880, N10453);
not NOT1 (N17886, N17877);
xor XOR2 (N17887, N17884, N14231);
xor XOR2 (N17888, N17870, N5738);
or OR4 (N17889, N17858, N14606, N3662, N6646);
not NOT1 (N17890, N17875);
nor NOR2 (N17891, N17887, N17192);
buf BUF1 (N17892, N17891);
buf BUF1 (N17893, N17885);
or OR2 (N17894, N17888, N3152);
and AND2 (N17895, N17889, N9189);
and AND4 (N17896, N17894, N11320, N9961, N5825);
nor NOR3 (N17897, N17893, N901, N10248);
nand NAND2 (N17898, N17883, N9174);
not NOT1 (N17899, N17874);
and AND3 (N17900, N17895, N16507, N4378);
buf BUF1 (N17901, N17892);
xor XOR2 (N17902, N17901, N7419);
nand NAND4 (N17903, N17869, N14755, N16829, N12952);
and AND2 (N17904, N17899, N16502);
nand NAND3 (N17905, N17876, N17425, N3380);
xor XOR2 (N17906, N17890, N11120);
not NOT1 (N17907, N17898);
nor NOR4 (N17908, N17900, N3477, N375, N6588);
not NOT1 (N17909, N17904);
nor NOR3 (N17910, N17897, N11553, N4892);
not NOT1 (N17911, N17909);
nand NAND4 (N17912, N17908, N9726, N16564, N6719);
or OR2 (N17913, N17896, N14547);
buf BUF1 (N17914, N17907);
and AND4 (N17915, N17906, N4662, N14709, N4898);
buf BUF1 (N17916, N17915);
not NOT1 (N17917, N17913);
buf BUF1 (N17918, N17905);
and AND3 (N17919, N17903, N11906, N13893);
or OR2 (N17920, N17902, N4712);
or OR2 (N17921, N17919, N914);
nand NAND3 (N17922, N17886, N11696, N10706);
not NOT1 (N17923, N17911);
nand NAND2 (N17924, N17922, N8249);
not NOT1 (N17925, N17923);
not NOT1 (N17926, N17924);
nand NAND2 (N17927, N17920, N14586);
buf BUF1 (N17928, N17918);
nor NOR2 (N17929, N17928, N6920);
or OR3 (N17930, N17910, N10469, N14501);
nand NAND4 (N17931, N17916, N16109, N5020, N13663);
xor XOR2 (N17932, N17926, N9654);
buf BUF1 (N17933, N17925);
xor XOR2 (N17934, N17921, N3385);
nand NAND3 (N17935, N17930, N12909, N17271);
nor NOR3 (N17936, N17927, N616, N3591);
nor NOR2 (N17937, N17917, N8522);
nand NAND3 (N17938, N17929, N457, N12131);
buf BUF1 (N17939, N17934);
not NOT1 (N17940, N17912);
and AND3 (N17941, N17940, N11545, N8428);
nor NOR2 (N17942, N17931, N14929);
xor XOR2 (N17943, N17939, N12858);
and AND3 (N17944, N17941, N4020, N7652);
not NOT1 (N17945, N17937);
or OR4 (N17946, N17943, N12582, N7941, N4997);
nor NOR4 (N17947, N17914, N2403, N10976, N4131);
nand NAND3 (N17948, N17936, N9992, N9169);
nand NAND4 (N17949, N17933, N5612, N16660, N6360);
buf BUF1 (N17950, N17944);
buf BUF1 (N17951, N17945);
or OR4 (N17952, N17946, N3324, N14756, N11222);
and AND2 (N17953, N17952, N11737);
and AND3 (N17954, N17949, N11113, N10978);
and AND3 (N17955, N17935, N12794, N9488);
nand NAND2 (N17956, N17938, N3648);
nand NAND3 (N17957, N17932, N970, N3230);
nor NOR4 (N17958, N17951, N3334, N5930, N366);
xor XOR2 (N17959, N17955, N17920);
not NOT1 (N17960, N17942);
or OR4 (N17961, N17954, N1009, N8040, N1686);
not NOT1 (N17962, N17959);
and AND2 (N17963, N17948, N9543);
and AND3 (N17964, N17957, N17110, N3049);
nor NOR2 (N17965, N17960, N14732);
nand NAND3 (N17966, N17950, N12082, N6041);
nor NOR4 (N17967, N17964, N16578, N12774, N15076);
nand NAND2 (N17968, N17966, N10855);
not NOT1 (N17969, N17953);
not NOT1 (N17970, N17962);
nor NOR2 (N17971, N17956, N17437);
xor XOR2 (N17972, N17969, N2035);
xor XOR2 (N17973, N17965, N1884);
not NOT1 (N17974, N17970);
or OR2 (N17975, N17974, N5149);
not NOT1 (N17976, N17967);
xor XOR2 (N17977, N17972, N212);
or OR3 (N17978, N17973, N14209, N16663);
or OR4 (N17979, N17968, N6427, N8791, N14365);
nand NAND3 (N17980, N17979, N10376, N3936);
buf BUF1 (N17981, N17977);
nor NOR2 (N17982, N17947, N7973);
nand NAND2 (N17983, N17980, N2294);
or OR2 (N17984, N17961, N13033);
nand NAND2 (N17985, N17963, N1356);
xor XOR2 (N17986, N17978, N13903);
or OR3 (N17987, N17976, N1021, N11229);
not NOT1 (N17988, N17971);
nor NOR3 (N17989, N17986, N6971, N1724);
xor XOR2 (N17990, N17981, N17086);
and AND2 (N17991, N17982, N13159);
xor XOR2 (N17992, N17984, N17089);
nand NAND4 (N17993, N17975, N3846, N11058, N16117);
nand NAND3 (N17994, N17987, N16453, N16459);
nand NAND3 (N17995, N17988, N667, N3495);
buf BUF1 (N17996, N17993);
buf BUF1 (N17997, N17995);
nand NAND3 (N17998, N17994, N294, N14365);
buf BUF1 (N17999, N17992);
nor NOR4 (N18000, N17958, N548, N7370, N6319);
and AND4 (N18001, N17999, N2161, N2573, N12620);
buf BUF1 (N18002, N17989);
xor XOR2 (N18003, N17990, N9706);
or OR3 (N18004, N17997, N14417, N16564);
or OR2 (N18005, N18001, N1031);
and AND4 (N18006, N18000, N9698, N9203, N13499);
nand NAND4 (N18007, N18003, N9481, N7348, N1251);
nand NAND4 (N18008, N17991, N6930, N1909, N4423);
xor XOR2 (N18009, N18002, N17812);
or OR4 (N18010, N17998, N2569, N2112, N4373);
and AND2 (N18011, N17983, N1173);
and AND2 (N18012, N17985, N382);
xor XOR2 (N18013, N18006, N2860);
nand NAND3 (N18014, N17996, N6049, N16999);
and AND2 (N18015, N18014, N1600);
nor NOR4 (N18016, N18004, N16047, N10457, N7849);
nor NOR3 (N18017, N18011, N6760, N4133);
xor XOR2 (N18018, N18013, N4492);
buf BUF1 (N18019, N18017);
nand NAND4 (N18020, N18010, N12340, N1290, N15870);
nor NOR2 (N18021, N18012, N9995);
or OR3 (N18022, N18021, N4901, N5051);
nand NAND2 (N18023, N18005, N7695);
nor NOR2 (N18024, N18007, N4591);
and AND2 (N18025, N18024, N1245);
buf BUF1 (N18026, N18015);
not NOT1 (N18027, N18026);
nor NOR3 (N18028, N18008, N6786, N17467);
xor XOR2 (N18029, N18009, N13865);
nor NOR2 (N18030, N18029, N4878);
or OR2 (N18031, N18028, N10344);
or OR2 (N18032, N18025, N13850);
or OR2 (N18033, N18032, N11518);
not NOT1 (N18034, N18023);
or OR4 (N18035, N18020, N8136, N13016, N9762);
nor NOR2 (N18036, N18018, N3386);
nor NOR4 (N18037, N18030, N10236, N16010, N2602);
nor NOR2 (N18038, N18016, N8785);
nand NAND3 (N18039, N18019, N17385, N5547);
or OR4 (N18040, N18035, N5438, N2174, N16173);
nor NOR3 (N18041, N18034, N8319, N10768);
xor XOR2 (N18042, N18033, N3946);
and AND4 (N18043, N18042, N780, N14014, N3546);
buf BUF1 (N18044, N18043);
nand NAND4 (N18045, N18038, N1593, N2392, N4055);
and AND3 (N18046, N18036, N1983, N5502);
nand NAND4 (N18047, N18031, N1727, N9986, N955);
buf BUF1 (N18048, N18044);
xor XOR2 (N18049, N18045, N3334);
xor XOR2 (N18050, N18048, N15401);
nand NAND3 (N18051, N18040, N11539, N10198);
not NOT1 (N18052, N18022);
nor NOR3 (N18053, N18047, N5068, N7867);
xor XOR2 (N18054, N18041, N16891);
nand NAND3 (N18055, N18039, N15475, N7174);
and AND3 (N18056, N18037, N7349, N2184);
or OR4 (N18057, N18054, N6002, N15957, N5815);
nand NAND2 (N18058, N18053, N2000);
buf BUF1 (N18059, N18055);
xor XOR2 (N18060, N18051, N12265);
nand NAND3 (N18061, N18060, N8314, N1595);
not NOT1 (N18062, N18057);
xor XOR2 (N18063, N18059, N4678);
xor XOR2 (N18064, N18063, N13600);
and AND4 (N18065, N18056, N6364, N1947, N11385);
nand NAND4 (N18066, N18046, N12760, N2969, N3411);
nor NOR2 (N18067, N18062, N11890);
or OR2 (N18068, N18064, N7985);
or OR2 (N18069, N18065, N4468);
nor NOR4 (N18070, N18069, N4595, N15093, N17468);
and AND3 (N18071, N18066, N16743, N5153);
and AND4 (N18072, N18071, N11301, N2633, N15231);
nor NOR2 (N18073, N18072, N13752);
nand NAND2 (N18074, N18073, N17895);
or OR4 (N18075, N18049, N1736, N10410, N13309);
not NOT1 (N18076, N18075);
or OR3 (N18077, N18067, N1773, N8811);
buf BUF1 (N18078, N18068);
nor NOR3 (N18079, N18070, N1045, N7243);
xor XOR2 (N18080, N18076, N16783);
buf BUF1 (N18081, N18058);
not NOT1 (N18082, N18050);
and AND2 (N18083, N18078, N412);
not NOT1 (N18084, N18080);
not NOT1 (N18085, N18052);
nor NOR3 (N18086, N18061, N16062, N13456);
not NOT1 (N18087, N18082);
and AND4 (N18088, N18085, N7665, N16148, N13053);
buf BUF1 (N18089, N18086);
or OR3 (N18090, N18027, N14669, N16442);
buf BUF1 (N18091, N18084);
buf BUF1 (N18092, N18081);
xor XOR2 (N18093, N18079, N1252);
not NOT1 (N18094, N18087);
nor NOR3 (N18095, N18091, N17558, N5523);
buf BUF1 (N18096, N18094);
not NOT1 (N18097, N18074);
nor NOR3 (N18098, N18083, N14721, N5754);
buf BUF1 (N18099, N18097);
buf BUF1 (N18100, N18095);
buf BUF1 (N18101, N18100);
and AND3 (N18102, N18092, N17715, N9995);
xor XOR2 (N18103, N18098, N12574);
xor XOR2 (N18104, N18088, N11953);
xor XOR2 (N18105, N18101, N11282);
nand NAND4 (N18106, N18099, N4490, N16374, N1147);
not NOT1 (N18107, N18104);
nand NAND2 (N18108, N18105, N16159);
not NOT1 (N18109, N18106);
nor NOR2 (N18110, N18077, N9050);
nor NOR3 (N18111, N18102, N2760, N8335);
and AND2 (N18112, N18111, N7598);
and AND3 (N18113, N18093, N11724, N2066);
buf BUF1 (N18114, N18103);
xor XOR2 (N18115, N18112, N12885);
nand NAND2 (N18116, N18113, N14645);
nor NOR3 (N18117, N18096, N10832, N1274);
and AND4 (N18118, N18116, N9981, N3902, N9427);
nand NAND2 (N18119, N18108, N4701);
buf BUF1 (N18120, N18119);
not NOT1 (N18121, N18107);
not NOT1 (N18122, N18121);
xor XOR2 (N18123, N18117, N3035);
or OR2 (N18124, N18120, N4475);
and AND2 (N18125, N18114, N12707);
or OR3 (N18126, N18123, N15189, N15101);
nor NOR4 (N18127, N18089, N5965, N12560, N8385);
buf BUF1 (N18128, N18118);
nor NOR3 (N18129, N18115, N5070, N9961);
xor XOR2 (N18130, N18122, N14428);
buf BUF1 (N18131, N18110);
or OR2 (N18132, N18129, N8681);
buf BUF1 (N18133, N18131);
or OR2 (N18134, N18132, N1823);
and AND2 (N18135, N18090, N21);
buf BUF1 (N18136, N18133);
and AND3 (N18137, N18127, N3849, N11102);
not NOT1 (N18138, N18109);
not NOT1 (N18139, N18130);
not NOT1 (N18140, N18138);
and AND2 (N18141, N18134, N7608);
xor XOR2 (N18142, N18135, N133);
nand NAND2 (N18143, N18124, N8897);
not NOT1 (N18144, N18140);
not NOT1 (N18145, N18126);
nor NOR2 (N18146, N18141, N17133);
nand NAND3 (N18147, N18145, N779, N13355);
nand NAND2 (N18148, N18128, N1401);
xor XOR2 (N18149, N18136, N9212);
or OR2 (N18150, N18149, N15770);
not NOT1 (N18151, N18144);
not NOT1 (N18152, N18150);
xor XOR2 (N18153, N18146, N7889);
and AND4 (N18154, N18143, N13215, N9547, N17682);
nand NAND4 (N18155, N18151, N11668, N8154, N10716);
not NOT1 (N18156, N18125);
xor XOR2 (N18157, N18137, N15379);
not NOT1 (N18158, N18148);
nand NAND3 (N18159, N18158, N15299, N4094);
or OR3 (N18160, N18156, N4135, N12457);
or OR2 (N18161, N18155, N8056);
buf BUF1 (N18162, N18160);
buf BUF1 (N18163, N18147);
nand NAND2 (N18164, N18163, N12350);
nand NAND4 (N18165, N18161, N4615, N3814, N2708);
or OR4 (N18166, N18157, N546, N7717, N5573);
nand NAND2 (N18167, N18164, N14155);
not NOT1 (N18168, N18167);
or OR2 (N18169, N18153, N16811);
xor XOR2 (N18170, N18162, N9766);
nor NOR4 (N18171, N18139, N15115, N12792, N10283);
xor XOR2 (N18172, N18168, N16666);
buf BUF1 (N18173, N18142);
nor NOR2 (N18174, N18170, N1222);
or OR3 (N18175, N18173, N10943, N3189);
buf BUF1 (N18176, N18169);
nand NAND2 (N18177, N18171, N10440);
not NOT1 (N18178, N18166);
nor NOR3 (N18179, N18176, N7600, N7888);
or OR3 (N18180, N18174, N10034, N3854);
or OR4 (N18181, N18178, N13911, N1053, N2747);
not NOT1 (N18182, N18175);
or OR4 (N18183, N18154, N1878, N1645, N3129);
not NOT1 (N18184, N18177);
xor XOR2 (N18185, N18182, N17153);
or OR4 (N18186, N18184, N7729, N8314, N360);
or OR4 (N18187, N18179, N13896, N7200, N14457);
not NOT1 (N18188, N18159);
or OR4 (N18189, N18188, N4434, N10884, N3177);
nand NAND2 (N18190, N18186, N1192);
and AND2 (N18191, N18165, N6398);
or OR2 (N18192, N18185, N2130);
buf BUF1 (N18193, N18181);
not NOT1 (N18194, N18152);
not NOT1 (N18195, N18187);
or OR2 (N18196, N18183, N11213);
nand NAND3 (N18197, N18193, N15288, N13342);
nand NAND4 (N18198, N18196, N2873, N1991, N4443);
and AND2 (N18199, N18198, N7738);
nand NAND3 (N18200, N18190, N11293, N18089);
nand NAND3 (N18201, N18192, N8044, N7467);
not NOT1 (N18202, N18189);
buf BUF1 (N18203, N18194);
xor XOR2 (N18204, N18191, N15375);
nand NAND3 (N18205, N18203, N17571, N3711);
and AND3 (N18206, N18199, N9377, N10667);
nor NOR4 (N18207, N18195, N6272, N13799, N16226);
not NOT1 (N18208, N18204);
or OR3 (N18209, N18172, N859, N18149);
and AND2 (N18210, N18209, N609);
buf BUF1 (N18211, N18202);
xor XOR2 (N18212, N18201, N3967);
xor XOR2 (N18213, N18208, N4243);
and AND2 (N18214, N18207, N4808);
or OR4 (N18215, N18197, N881, N957, N5513);
and AND2 (N18216, N18210, N10017);
nor NOR2 (N18217, N18206, N17625);
nor NOR2 (N18218, N18216, N11400);
nand NAND4 (N18219, N18211, N3584, N4612, N9424);
and AND4 (N18220, N18205, N5498, N7126, N6815);
buf BUF1 (N18221, N18200);
nand NAND3 (N18222, N18180, N1011, N279);
buf BUF1 (N18223, N18214);
not NOT1 (N18224, N18222);
nand NAND2 (N18225, N18212, N13941);
not NOT1 (N18226, N18225);
nor NOR3 (N18227, N18213, N15000, N14977);
or OR2 (N18228, N18221, N17092);
and AND2 (N18229, N18218, N245);
xor XOR2 (N18230, N18226, N8808);
not NOT1 (N18231, N18219);
not NOT1 (N18232, N18231);
or OR2 (N18233, N18232, N1632);
buf BUF1 (N18234, N18220);
or OR4 (N18235, N18229, N17759, N4945, N9594);
nand NAND4 (N18236, N18224, N11741, N7045, N16453);
nor NOR2 (N18237, N18217, N5757);
or OR4 (N18238, N18223, N10230, N553, N10539);
or OR4 (N18239, N18227, N1558, N17275, N17860);
and AND3 (N18240, N18215, N6294, N3000);
nand NAND2 (N18241, N18235, N11693);
xor XOR2 (N18242, N18233, N14937);
nor NOR4 (N18243, N18240, N17064, N13933, N5942);
nand NAND2 (N18244, N18237, N11277);
not NOT1 (N18245, N18244);
nand NAND2 (N18246, N18238, N1627);
and AND4 (N18247, N18242, N1798, N16485, N4993);
nand NAND3 (N18248, N18230, N12966, N4697);
buf BUF1 (N18249, N18245);
or OR2 (N18250, N18239, N16564);
nor NOR3 (N18251, N18247, N13868, N4205);
not NOT1 (N18252, N18249);
xor XOR2 (N18253, N18251, N7962);
buf BUF1 (N18254, N18246);
nand NAND3 (N18255, N18243, N11175, N16198);
and AND3 (N18256, N18241, N3533, N11312);
nor NOR2 (N18257, N18253, N7475);
or OR2 (N18258, N18256, N6830);
and AND4 (N18259, N18255, N14279, N5832, N17907);
not NOT1 (N18260, N18236);
nor NOR4 (N18261, N18228, N13905, N3679, N7552);
xor XOR2 (N18262, N18250, N11265);
or OR2 (N18263, N18262, N13246);
nor NOR4 (N18264, N18263, N16749, N16070, N4988);
buf BUF1 (N18265, N18252);
and AND4 (N18266, N18260, N2637, N5654, N4932);
nand NAND2 (N18267, N18264, N3795);
nor NOR2 (N18268, N18265, N2637);
xor XOR2 (N18269, N18267, N15951);
or OR4 (N18270, N18268, N5737, N17301, N9823);
and AND2 (N18271, N18248, N9660);
nor NOR3 (N18272, N18261, N10416, N7739);
and AND3 (N18273, N18257, N12792, N17005);
or OR3 (N18274, N18273, N313, N516);
not NOT1 (N18275, N18269);
nand NAND4 (N18276, N18254, N8777, N14058, N3050);
xor XOR2 (N18277, N18271, N9437);
or OR2 (N18278, N18266, N7007);
nor NOR4 (N18279, N18277, N5420, N3428, N9977);
xor XOR2 (N18280, N18272, N10798);
nor NOR3 (N18281, N18280, N10173, N1519);
not NOT1 (N18282, N18270);
or OR3 (N18283, N18278, N17557, N7391);
buf BUF1 (N18284, N18274);
nor NOR3 (N18285, N18258, N5062, N8306);
or OR3 (N18286, N18282, N5858, N18163);
nor NOR2 (N18287, N18281, N1670);
xor XOR2 (N18288, N18285, N5905);
nor NOR3 (N18289, N18259, N2028, N4865);
xor XOR2 (N18290, N18283, N12220);
and AND3 (N18291, N18279, N7109, N13485);
not NOT1 (N18292, N18284);
xor XOR2 (N18293, N18289, N7660);
nand NAND3 (N18294, N18288, N2325, N14932);
nor NOR3 (N18295, N18276, N12779, N9005);
not NOT1 (N18296, N18287);
xor XOR2 (N18297, N18275, N17615);
nor NOR3 (N18298, N18290, N4076, N1181);
not NOT1 (N18299, N18293);
nor NOR4 (N18300, N18286, N16620, N10244, N17565);
or OR2 (N18301, N18298, N14881);
not NOT1 (N18302, N18301);
not NOT1 (N18303, N18302);
nor NOR2 (N18304, N18295, N15037);
xor XOR2 (N18305, N18304, N17316);
nor NOR3 (N18306, N18297, N6876, N11848);
nor NOR3 (N18307, N18234, N10086, N13377);
buf BUF1 (N18308, N18306);
or OR4 (N18309, N18307, N4497, N1012, N341);
or OR2 (N18310, N18299, N13996);
xor XOR2 (N18311, N18300, N1314);
buf BUF1 (N18312, N18309);
nand NAND4 (N18313, N18310, N17831, N610, N8938);
buf BUF1 (N18314, N18308);
buf BUF1 (N18315, N18294);
buf BUF1 (N18316, N18313);
not NOT1 (N18317, N18303);
not NOT1 (N18318, N18312);
not NOT1 (N18319, N18318);
or OR4 (N18320, N18316, N6013, N10543, N6796);
not NOT1 (N18321, N18320);
or OR4 (N18322, N18305, N8712, N6253, N412);
nand NAND4 (N18323, N18315, N15372, N6353, N7329);
buf BUF1 (N18324, N18319);
buf BUF1 (N18325, N18323);
nand NAND3 (N18326, N18325, N719, N4808);
and AND4 (N18327, N18324, N6729, N2440, N3625);
xor XOR2 (N18328, N18317, N15038);
not NOT1 (N18329, N18328);
buf BUF1 (N18330, N18322);
buf BUF1 (N18331, N18311);
or OR4 (N18332, N18326, N10804, N774, N11461);
nor NOR4 (N18333, N18331, N11148, N1683, N6759);
buf BUF1 (N18334, N18327);
nand NAND3 (N18335, N18314, N16508, N323);
not NOT1 (N18336, N18329);
buf BUF1 (N18337, N18335);
and AND2 (N18338, N18291, N7468);
or OR4 (N18339, N18334, N15214, N16433, N13318);
and AND4 (N18340, N18330, N16432, N7096, N13505);
or OR3 (N18341, N18296, N4806, N8283);
nor NOR2 (N18342, N18338, N7213);
buf BUF1 (N18343, N18321);
buf BUF1 (N18344, N18342);
nor NOR3 (N18345, N18344, N11836, N12585);
nor NOR2 (N18346, N18345, N9247);
and AND2 (N18347, N18336, N12780);
nor NOR4 (N18348, N18333, N10619, N8149, N17138);
nor NOR3 (N18349, N18292, N11708, N14994);
or OR3 (N18350, N18339, N5860, N425);
nand NAND3 (N18351, N18343, N17475, N4776);
not NOT1 (N18352, N18350);
and AND3 (N18353, N18347, N1170, N17099);
buf BUF1 (N18354, N18337);
xor XOR2 (N18355, N18352, N11781);
buf BUF1 (N18356, N18351);
nand NAND2 (N18357, N18332, N12180);
not NOT1 (N18358, N18349);
not NOT1 (N18359, N18348);
and AND2 (N18360, N18356, N16839);
not NOT1 (N18361, N18355);
and AND4 (N18362, N18341, N16694, N5989, N10518);
xor XOR2 (N18363, N18340, N13708);
not NOT1 (N18364, N18363);
nand NAND2 (N18365, N18360, N14511);
nand NAND4 (N18366, N18365, N12449, N17814, N15638);
buf BUF1 (N18367, N18359);
not NOT1 (N18368, N18366);
nand NAND2 (N18369, N18357, N11105);
xor XOR2 (N18370, N18361, N7293);
and AND3 (N18371, N18362, N15756, N1386);
and AND3 (N18372, N18358, N13939, N10959);
nand NAND3 (N18373, N18367, N17343, N6258);
xor XOR2 (N18374, N18372, N16781);
and AND4 (N18375, N18374, N12928, N9289, N18261);
or OR3 (N18376, N18373, N15408, N11419);
or OR4 (N18377, N18371, N14961, N5315, N1760);
nor NOR4 (N18378, N18346, N3103, N11244, N1964);
and AND3 (N18379, N18375, N2891, N10302);
nor NOR4 (N18380, N18376, N174, N10946, N16472);
not NOT1 (N18381, N18364);
not NOT1 (N18382, N18380);
not NOT1 (N18383, N18369);
not NOT1 (N18384, N18354);
xor XOR2 (N18385, N18379, N292);
and AND4 (N18386, N18385, N11414, N9589, N6336);
nor NOR2 (N18387, N18382, N9504);
nor NOR4 (N18388, N18383, N4369, N15946, N10668);
xor XOR2 (N18389, N18377, N17207);
and AND2 (N18390, N18370, N4678);
not NOT1 (N18391, N18384);
not NOT1 (N18392, N18386);
or OR3 (N18393, N18388, N9105, N17725);
nand NAND2 (N18394, N18389, N2990);
nand NAND2 (N18395, N18391, N8384);
nor NOR2 (N18396, N18395, N12610);
or OR4 (N18397, N18353, N10365, N16258, N1412);
xor XOR2 (N18398, N18393, N2471);
or OR4 (N18399, N18387, N2204, N4836, N16563);
or OR2 (N18400, N18392, N16464);
not NOT1 (N18401, N18394);
not NOT1 (N18402, N18401);
xor XOR2 (N18403, N18399, N9574);
nor NOR2 (N18404, N18381, N5438);
not NOT1 (N18405, N18390);
or OR3 (N18406, N18398, N6778, N3411);
buf BUF1 (N18407, N18396);
and AND4 (N18408, N18378, N10424, N794, N4980);
not NOT1 (N18409, N18402);
not NOT1 (N18410, N18409);
xor XOR2 (N18411, N18397, N17223);
nor NOR3 (N18412, N18410, N2528, N15086);
not NOT1 (N18413, N18403);
xor XOR2 (N18414, N18406, N11426);
buf BUF1 (N18415, N18408);
nand NAND4 (N18416, N18407, N7712, N9502, N6286);
and AND2 (N18417, N18368, N7289);
and AND3 (N18418, N18411, N223, N18338);
xor XOR2 (N18419, N18418, N9770);
buf BUF1 (N18420, N18415);
xor XOR2 (N18421, N18419, N10980);
xor XOR2 (N18422, N18405, N4883);
not NOT1 (N18423, N18420);
nor NOR3 (N18424, N18417, N6953, N18285);
xor XOR2 (N18425, N18414, N2685);
nor NOR4 (N18426, N18416, N15502, N1938, N5223);
and AND4 (N18427, N18413, N3567, N7603, N3762);
or OR2 (N18428, N18404, N14041);
or OR3 (N18429, N18412, N10994, N15243);
not NOT1 (N18430, N18421);
or OR2 (N18431, N18426, N12435);
buf BUF1 (N18432, N18431);
buf BUF1 (N18433, N18430);
nor NOR4 (N18434, N18432, N13669, N4628, N9392);
nor NOR3 (N18435, N18434, N14827, N11243);
nand NAND4 (N18436, N18435, N9750, N11047, N11124);
and AND3 (N18437, N18429, N1794, N9312);
buf BUF1 (N18438, N18428);
not NOT1 (N18439, N18436);
or OR4 (N18440, N18423, N10102, N1580, N6668);
xor XOR2 (N18441, N18425, N3860);
and AND2 (N18442, N18422, N6263);
buf BUF1 (N18443, N18433);
xor XOR2 (N18444, N18440, N1028);
not NOT1 (N18445, N18427);
not NOT1 (N18446, N18439);
xor XOR2 (N18447, N18444, N14225);
buf BUF1 (N18448, N18424);
buf BUF1 (N18449, N18443);
nand NAND2 (N18450, N18442, N10664);
not NOT1 (N18451, N18445);
and AND3 (N18452, N18449, N11890, N2037);
nor NOR2 (N18453, N18441, N7641);
xor XOR2 (N18454, N18447, N15516);
not NOT1 (N18455, N18446);
not NOT1 (N18456, N18450);
and AND4 (N18457, N18453, N11824, N4493, N12967);
or OR3 (N18458, N18457, N11758, N11147);
and AND4 (N18459, N18451, N13694, N14768, N18107);
buf BUF1 (N18460, N18458);
buf BUF1 (N18461, N18438);
or OR4 (N18462, N18400, N10982, N5837, N17137);
nand NAND2 (N18463, N18448, N1925);
or OR3 (N18464, N18452, N5903, N6032);
and AND3 (N18465, N18462, N4787, N4715);
or OR2 (N18466, N18463, N12551);
xor XOR2 (N18467, N18466, N13922);
nand NAND3 (N18468, N18460, N16637, N14154);
or OR3 (N18469, N18467, N4475, N18004);
nand NAND2 (N18470, N18454, N3189);
buf BUF1 (N18471, N18456);
xor XOR2 (N18472, N18469, N9182);
buf BUF1 (N18473, N18455);
buf BUF1 (N18474, N18472);
or OR4 (N18475, N18470, N6151, N13048, N16474);
and AND2 (N18476, N18473, N4697);
xor XOR2 (N18477, N18459, N4371);
nand NAND3 (N18478, N18477, N9901, N17440);
buf BUF1 (N18479, N18464);
and AND2 (N18480, N18461, N3919);
nand NAND2 (N18481, N18437, N5917);
not NOT1 (N18482, N18468);
and AND2 (N18483, N18471, N14441);
xor XOR2 (N18484, N18480, N1611);
nor NOR2 (N18485, N18475, N14676);
nand NAND4 (N18486, N18476, N8647, N1442, N13608);
nand NAND2 (N18487, N18465, N5584);
nand NAND2 (N18488, N18484, N10973);
xor XOR2 (N18489, N18482, N5812);
nor NOR3 (N18490, N18486, N11021, N17429);
not NOT1 (N18491, N18488);
buf BUF1 (N18492, N18491);
or OR3 (N18493, N18487, N9107, N9992);
not NOT1 (N18494, N18493);
buf BUF1 (N18495, N18474);
xor XOR2 (N18496, N18489, N12804);
or OR3 (N18497, N18494, N4520, N10114);
nand NAND2 (N18498, N18485, N8544);
and AND4 (N18499, N18498, N15330, N4697, N5600);
or OR4 (N18500, N18490, N13104, N9180, N5579);
nor NOR4 (N18501, N18496, N14258, N2862, N8628);
buf BUF1 (N18502, N18499);
xor XOR2 (N18503, N18483, N18235);
and AND2 (N18504, N18481, N3592);
xor XOR2 (N18505, N18478, N11366);
and AND2 (N18506, N18495, N14114);
xor XOR2 (N18507, N18479, N11655);
and AND4 (N18508, N18497, N5545, N12795, N1164);
nand NAND2 (N18509, N18504, N967);
not NOT1 (N18510, N18509);
buf BUF1 (N18511, N18503);
not NOT1 (N18512, N18506);
nand NAND3 (N18513, N18501, N4506, N5901);
not NOT1 (N18514, N18492);
xor XOR2 (N18515, N18508, N968);
xor XOR2 (N18516, N18511, N15854);
and AND2 (N18517, N18514, N2554);
nand NAND4 (N18518, N18516, N5141, N11992, N5397);
and AND2 (N18519, N18507, N8584);
nor NOR2 (N18520, N18512, N16998);
nor NOR2 (N18521, N18500, N3871);
not NOT1 (N18522, N18517);
not NOT1 (N18523, N18519);
nor NOR3 (N18524, N18510, N10633, N3623);
nor NOR4 (N18525, N18523, N1647, N8178, N15005);
buf BUF1 (N18526, N18513);
xor XOR2 (N18527, N18505, N3294);
and AND2 (N18528, N18524, N17658);
not NOT1 (N18529, N18515);
nor NOR4 (N18530, N18528, N11269, N4440, N15564);
or OR4 (N18531, N18526, N17949, N14640, N18185);
nor NOR4 (N18532, N18525, N18114, N17222, N57);
nand NAND4 (N18533, N18527, N6845, N15104, N18375);
xor XOR2 (N18534, N18531, N11278);
or OR3 (N18535, N18520, N17243, N15459);
xor XOR2 (N18536, N18534, N17976);
nor NOR2 (N18537, N18535, N15502);
buf BUF1 (N18538, N18530);
nor NOR2 (N18539, N18502, N6504);
xor XOR2 (N18540, N18538, N3549);
buf BUF1 (N18541, N18532);
and AND2 (N18542, N18536, N17485);
xor XOR2 (N18543, N18522, N6985);
xor XOR2 (N18544, N18540, N8869);
not NOT1 (N18545, N18533);
nor NOR3 (N18546, N18529, N15768, N8291);
xor XOR2 (N18547, N18537, N5791);
or OR2 (N18548, N18539, N17513);
nor NOR3 (N18549, N18544, N13329, N5392);
or OR2 (N18550, N18547, N16910);
nor NOR4 (N18551, N18541, N18459, N5297, N18332);
not NOT1 (N18552, N18549);
buf BUF1 (N18553, N18545);
and AND4 (N18554, N18551, N12112, N990, N5070);
and AND4 (N18555, N18548, N7166, N3364, N11613);
not NOT1 (N18556, N18553);
buf BUF1 (N18557, N18550);
buf BUF1 (N18558, N18557);
not NOT1 (N18559, N18546);
xor XOR2 (N18560, N18552, N5993);
xor XOR2 (N18561, N18542, N13157);
and AND3 (N18562, N18554, N5960, N12347);
buf BUF1 (N18563, N18556);
nor NOR4 (N18564, N18555, N3501, N16597, N985);
not NOT1 (N18565, N18521);
xor XOR2 (N18566, N18562, N6258);
not NOT1 (N18567, N18560);
buf BUF1 (N18568, N18566);
buf BUF1 (N18569, N18558);
or OR4 (N18570, N18564, N16079, N9623, N18088);
xor XOR2 (N18571, N18569, N13494);
and AND2 (N18572, N18568, N2608);
buf BUF1 (N18573, N18543);
nand NAND2 (N18574, N18518, N1503);
nor NOR2 (N18575, N18563, N7305);
and AND2 (N18576, N18573, N15296);
and AND3 (N18577, N18574, N7152, N13397);
nand NAND2 (N18578, N18576, N16849);
nand NAND2 (N18579, N18570, N1948);
xor XOR2 (N18580, N18571, N12037);
and AND2 (N18581, N18575, N3142);
xor XOR2 (N18582, N18580, N16523);
xor XOR2 (N18583, N18579, N17981);
nor NOR3 (N18584, N18583, N13145, N3866);
not NOT1 (N18585, N18578);
nor NOR3 (N18586, N18584, N11460, N9437);
nand NAND4 (N18587, N18577, N7419, N2762, N7578);
and AND2 (N18588, N18581, N12248);
nand NAND4 (N18589, N18572, N8211, N15325, N11271);
nand NAND2 (N18590, N18559, N9478);
nand NAND2 (N18591, N18582, N8042);
and AND2 (N18592, N18567, N11489);
buf BUF1 (N18593, N18587);
xor XOR2 (N18594, N18565, N17628);
xor XOR2 (N18595, N18589, N826);
buf BUF1 (N18596, N18586);
buf BUF1 (N18597, N18590);
xor XOR2 (N18598, N18597, N12673);
xor XOR2 (N18599, N18592, N8997);
or OR3 (N18600, N18599, N11893, N5746);
or OR4 (N18601, N18561, N6518, N15270, N8776);
xor XOR2 (N18602, N18598, N1038);
xor XOR2 (N18603, N18594, N6687);
or OR4 (N18604, N18591, N2532, N17303, N7886);
and AND2 (N18605, N18600, N17735);
not NOT1 (N18606, N18593);
nand NAND2 (N18607, N18604, N7446);
buf BUF1 (N18608, N18603);
nand NAND4 (N18609, N18595, N12614, N8206, N993);
nand NAND2 (N18610, N18608, N2517);
not NOT1 (N18611, N18602);
not NOT1 (N18612, N18606);
and AND3 (N18613, N18596, N14034, N9621);
buf BUF1 (N18614, N18585);
buf BUF1 (N18615, N18612);
xor XOR2 (N18616, N18611, N10420);
buf BUF1 (N18617, N18610);
nor NOR4 (N18618, N18614, N13257, N13348, N7143);
xor XOR2 (N18619, N18605, N1540);
buf BUF1 (N18620, N18617);
and AND3 (N18621, N18619, N10569, N13177);
buf BUF1 (N18622, N18613);
and AND2 (N18623, N18609, N7410);
and AND4 (N18624, N18618, N16575, N12831, N9667);
or OR3 (N18625, N18616, N8281, N11764);
xor XOR2 (N18626, N18622, N11328);
not NOT1 (N18627, N18615);
nand NAND3 (N18628, N18621, N5254, N12165);
xor XOR2 (N18629, N18624, N11900);
xor XOR2 (N18630, N18601, N11444);
and AND3 (N18631, N18607, N2923, N4700);
or OR3 (N18632, N18628, N8642, N14838);
xor XOR2 (N18633, N18623, N4032);
not NOT1 (N18634, N18629);
and AND2 (N18635, N18634, N6106);
and AND4 (N18636, N18626, N4540, N14542, N18110);
buf BUF1 (N18637, N18588);
or OR4 (N18638, N18630, N8387, N11958, N8220);
not NOT1 (N18639, N18638);
and AND2 (N18640, N18636, N668);
nor NOR2 (N18641, N18625, N2663);
and AND3 (N18642, N18639, N13651, N10202);
and AND4 (N18643, N18631, N7936, N2059, N5334);
not NOT1 (N18644, N18635);
buf BUF1 (N18645, N18643);
xor XOR2 (N18646, N18637, N3328);
buf BUF1 (N18647, N18627);
and AND3 (N18648, N18642, N16657, N14452);
nand NAND3 (N18649, N18647, N15062, N8158);
nand NAND2 (N18650, N18620, N585);
and AND2 (N18651, N18650, N8336);
buf BUF1 (N18652, N18633);
xor XOR2 (N18653, N18646, N8053);
xor XOR2 (N18654, N18651, N1225);
nor NOR3 (N18655, N18645, N8089, N18005);
not NOT1 (N18656, N18648);
nand NAND2 (N18657, N18644, N6493);
or OR4 (N18658, N18649, N1121, N1862, N2526);
and AND2 (N18659, N18653, N363);
not NOT1 (N18660, N18657);
nand NAND2 (N18661, N18641, N2065);
nor NOR4 (N18662, N18655, N3349, N3066, N5695);
or OR2 (N18663, N18652, N14124);
and AND4 (N18664, N18654, N7422, N8155, N17015);
or OR2 (N18665, N18658, N15070);
xor XOR2 (N18666, N18663, N18321);
xor XOR2 (N18667, N18664, N3811);
nor NOR4 (N18668, N18640, N13075, N15234, N6875);
xor XOR2 (N18669, N18660, N1703);
buf BUF1 (N18670, N18666);
nor NOR3 (N18671, N18656, N6798, N18498);
not NOT1 (N18672, N18661);
or OR3 (N18673, N18669, N6956, N16723);
nand NAND3 (N18674, N18671, N5070, N6994);
not NOT1 (N18675, N18668);
nand NAND3 (N18676, N18667, N8639, N2342);
or OR3 (N18677, N18670, N17010, N6977);
buf BUF1 (N18678, N18665);
not NOT1 (N18679, N18672);
or OR3 (N18680, N18677, N6476, N10688);
or OR2 (N18681, N18675, N12951);
buf BUF1 (N18682, N18681);
not NOT1 (N18683, N18678);
nor NOR2 (N18684, N18674, N13129);
not NOT1 (N18685, N18673);
and AND3 (N18686, N18682, N1750, N6694);
and AND4 (N18687, N18683, N470, N15162, N7090);
not NOT1 (N18688, N18686);
buf BUF1 (N18689, N18676);
or OR2 (N18690, N18659, N16288);
not NOT1 (N18691, N18662);
nand NAND4 (N18692, N18679, N5877, N16252, N4292);
buf BUF1 (N18693, N18692);
or OR2 (N18694, N18688, N17858);
buf BUF1 (N18695, N18694);
or OR3 (N18696, N18685, N7917, N4793);
nand NAND2 (N18697, N18687, N13629);
and AND2 (N18698, N18689, N2217);
not NOT1 (N18699, N18695);
xor XOR2 (N18700, N18699, N4556);
and AND4 (N18701, N18691, N14505, N5627, N12300);
not NOT1 (N18702, N18693);
buf BUF1 (N18703, N18698);
buf BUF1 (N18704, N18700);
and AND4 (N18705, N18680, N17789, N1591, N8174);
or OR3 (N18706, N18697, N6944, N207);
nor NOR4 (N18707, N18701, N3641, N12194, N3596);
not NOT1 (N18708, N18703);
xor XOR2 (N18709, N18704, N5368);
xor XOR2 (N18710, N18690, N6394);
nor NOR4 (N18711, N18710, N6582, N2023, N10016);
buf BUF1 (N18712, N18709);
nand NAND2 (N18713, N18696, N8477);
buf BUF1 (N18714, N18712);
buf BUF1 (N18715, N18713);
or OR2 (N18716, N18711, N14179);
buf BUF1 (N18717, N18705);
and AND3 (N18718, N18716, N3010, N4163);
or OR4 (N18719, N18714, N16596, N5046, N4243);
nor NOR4 (N18720, N18708, N18492, N5848, N13350);
xor XOR2 (N18721, N18684, N13843);
xor XOR2 (N18722, N18632, N5906);
nor NOR3 (N18723, N18718, N5759, N8737);
not NOT1 (N18724, N18707);
and AND4 (N18725, N18724, N4449, N15569, N13557);
nand NAND3 (N18726, N18721, N4772, N7428);
nor NOR4 (N18727, N18715, N8462, N12511, N15762);
or OR4 (N18728, N18717, N7561, N17124, N8873);
not NOT1 (N18729, N18726);
nor NOR2 (N18730, N18728, N18584);
xor XOR2 (N18731, N18730, N11877);
not NOT1 (N18732, N18722);
not NOT1 (N18733, N18729);
xor XOR2 (N18734, N18706, N1562);
and AND3 (N18735, N18720, N4532, N17322);
or OR2 (N18736, N18702, N11457);
and AND3 (N18737, N18734, N14611, N3981);
nor NOR2 (N18738, N18735, N18664);
nand NAND2 (N18739, N18737, N6411);
not NOT1 (N18740, N18719);
xor XOR2 (N18741, N18732, N5414);
buf BUF1 (N18742, N18733);
or OR4 (N18743, N18727, N17450, N11819, N8525);
nor NOR4 (N18744, N18738, N14187, N11633, N2654);
or OR2 (N18745, N18731, N10046);
or OR4 (N18746, N18744, N10034, N15370, N13623);
buf BUF1 (N18747, N18736);
and AND3 (N18748, N18743, N14838, N9959);
or OR4 (N18749, N18741, N8744, N10546, N14601);
not NOT1 (N18750, N18725);
or OR3 (N18751, N18739, N13665, N12881);
nand NAND2 (N18752, N18750, N2575);
and AND2 (N18753, N18723, N11258);
and AND4 (N18754, N18749, N10598, N17356, N9353);
not NOT1 (N18755, N18747);
buf BUF1 (N18756, N18748);
or OR3 (N18757, N18754, N5244, N5090);
buf BUF1 (N18758, N18755);
or OR4 (N18759, N18753, N11616, N11530, N2375);
nor NOR4 (N18760, N18740, N1695, N12703, N14185);
xor XOR2 (N18761, N18751, N7906);
xor XOR2 (N18762, N18746, N193);
and AND3 (N18763, N18757, N1527, N15964);
xor XOR2 (N18764, N18759, N14310);
or OR2 (N18765, N18763, N4559);
xor XOR2 (N18766, N18756, N2059);
not NOT1 (N18767, N18761);
not NOT1 (N18768, N18762);
not NOT1 (N18769, N18764);
xor XOR2 (N18770, N18766, N6625);
or OR4 (N18771, N18760, N2021, N12135, N15663);
buf BUF1 (N18772, N18742);
nand NAND2 (N18773, N18745, N1695);
or OR3 (N18774, N18758, N11928, N17560);
nand NAND3 (N18775, N18769, N15448, N15842);
xor XOR2 (N18776, N18752, N12425);
buf BUF1 (N18777, N18767);
xor XOR2 (N18778, N18775, N196);
nand NAND2 (N18779, N18765, N8802);
and AND2 (N18780, N18776, N10773);
buf BUF1 (N18781, N18772);
xor XOR2 (N18782, N18770, N4382);
buf BUF1 (N18783, N18780);
buf BUF1 (N18784, N18777);
buf BUF1 (N18785, N18774);
xor XOR2 (N18786, N18782, N9130);
not NOT1 (N18787, N18786);
or OR4 (N18788, N18771, N8149, N4010, N5286);
xor XOR2 (N18789, N18788, N11019);
buf BUF1 (N18790, N18787);
or OR3 (N18791, N18783, N1122, N11167);
not NOT1 (N18792, N18791);
not NOT1 (N18793, N18778);
nor NOR4 (N18794, N18789, N14726, N3649, N6874);
xor XOR2 (N18795, N18768, N7811);
not NOT1 (N18796, N18779);
and AND4 (N18797, N18793, N7457, N16458, N9964);
xor XOR2 (N18798, N18773, N15596);
or OR2 (N18799, N18795, N4012);
and AND2 (N18800, N18797, N559);
buf BUF1 (N18801, N18799);
buf BUF1 (N18802, N18781);
and AND4 (N18803, N18792, N3764, N16331, N6286);
nand NAND4 (N18804, N18803, N13512, N18117, N13419);
buf BUF1 (N18805, N18785);
buf BUF1 (N18806, N18801);
nand NAND3 (N18807, N18784, N18394, N7301);
and AND3 (N18808, N18805, N16050, N1066);
xor XOR2 (N18809, N18798, N12968);
and AND2 (N18810, N18796, N15860);
nor NOR4 (N18811, N18804, N6113, N9739, N1951);
and AND3 (N18812, N18810, N15300, N11415);
nand NAND2 (N18813, N18808, N10913);
buf BUF1 (N18814, N18794);
and AND2 (N18815, N18802, N10809);
xor XOR2 (N18816, N18814, N18239);
buf BUF1 (N18817, N18811);
nand NAND4 (N18818, N18812, N116, N11965, N10012);
xor XOR2 (N18819, N18806, N4483);
xor XOR2 (N18820, N18809, N13878);
not NOT1 (N18821, N18820);
and AND4 (N18822, N18813, N10236, N11007, N2356);
xor XOR2 (N18823, N18790, N3937);
buf BUF1 (N18824, N18800);
buf BUF1 (N18825, N18817);
buf BUF1 (N18826, N18815);
xor XOR2 (N18827, N18807, N9057);
and AND3 (N18828, N18823, N3668, N9822);
xor XOR2 (N18829, N18826, N10366);
xor XOR2 (N18830, N18824, N651);
buf BUF1 (N18831, N18819);
nand NAND4 (N18832, N18827, N8324, N5048, N8297);
xor XOR2 (N18833, N18825, N12829);
or OR3 (N18834, N18832, N12713, N13000);
not NOT1 (N18835, N18821);
not NOT1 (N18836, N18833);
and AND4 (N18837, N18829, N2910, N7558, N10567);
and AND2 (N18838, N18837, N16019);
nand NAND2 (N18839, N18816, N6187);
and AND4 (N18840, N18835, N5369, N3166, N17966);
nand NAND3 (N18841, N18838, N11517, N5392);
nand NAND4 (N18842, N18818, N6223, N8832, N1863);
xor XOR2 (N18843, N18822, N4362);
not NOT1 (N18844, N18841);
or OR2 (N18845, N18836, N7321);
or OR3 (N18846, N18828, N8097, N8060);
buf BUF1 (N18847, N18831);
and AND2 (N18848, N18845, N9126);
nand NAND4 (N18849, N18834, N15162, N5655, N8040);
nor NOR4 (N18850, N18844, N12220, N1718, N7303);
nor NOR4 (N18851, N18850, N13165, N1518, N2280);
xor XOR2 (N18852, N18842, N4631);
xor XOR2 (N18853, N18852, N15725);
nand NAND2 (N18854, N18843, N15179);
and AND3 (N18855, N18849, N5518, N14171);
nand NAND3 (N18856, N18840, N7817, N3002);
nor NOR4 (N18857, N18847, N18423, N1077, N14581);
nor NOR2 (N18858, N18839, N17781);
not NOT1 (N18859, N18851);
or OR4 (N18860, N18848, N11835, N13405, N12321);
nand NAND2 (N18861, N18859, N8095);
buf BUF1 (N18862, N18855);
not NOT1 (N18863, N18853);
not NOT1 (N18864, N18863);
buf BUF1 (N18865, N18864);
xor XOR2 (N18866, N18862, N1043);
or OR4 (N18867, N18856, N10973, N16809, N113);
and AND3 (N18868, N18861, N10278, N13901);
nor NOR4 (N18869, N18858, N12437, N18137, N17323);
and AND4 (N18870, N18867, N2113, N4650, N16062);
nand NAND3 (N18871, N18830, N2118, N6794);
xor XOR2 (N18872, N18866, N2492);
xor XOR2 (N18873, N18860, N1711);
and AND2 (N18874, N18865, N18826);
and AND3 (N18875, N18874, N2389, N7976);
and AND3 (N18876, N18873, N957, N3091);
nand NAND4 (N18877, N18869, N2364, N13908, N10037);
xor XOR2 (N18878, N18876, N6794);
not NOT1 (N18879, N18846);
not NOT1 (N18880, N18872);
nor NOR2 (N18881, N18870, N2775);
xor XOR2 (N18882, N18871, N747);
xor XOR2 (N18883, N18875, N10803);
xor XOR2 (N18884, N18868, N12268);
xor XOR2 (N18885, N18883, N13757);
nor NOR3 (N18886, N18884, N4440, N6729);
xor XOR2 (N18887, N18881, N14663);
buf BUF1 (N18888, N18877);
or OR4 (N18889, N18854, N18447, N17566, N1965);
nand NAND4 (N18890, N18879, N2739, N5922, N10464);
buf BUF1 (N18891, N18889);
and AND4 (N18892, N18886, N10583, N752, N12437);
xor XOR2 (N18893, N18857, N12731);
nand NAND2 (N18894, N18892, N18335);
xor XOR2 (N18895, N18890, N13911);
nor NOR2 (N18896, N18888, N18429);
nor NOR2 (N18897, N18885, N5389);
or OR2 (N18898, N18895, N6831);
xor XOR2 (N18899, N18898, N3376);
xor XOR2 (N18900, N18880, N3107);
or OR3 (N18901, N18882, N6210, N16924);
nand NAND3 (N18902, N18896, N9472, N11127);
buf BUF1 (N18903, N18899);
and AND4 (N18904, N18902, N5552, N4436, N10260);
nor NOR2 (N18905, N18903, N4793);
xor XOR2 (N18906, N18904, N11398);
nor NOR3 (N18907, N18900, N17468, N560);
and AND4 (N18908, N18894, N13428, N18307, N2331);
nor NOR3 (N18909, N18905, N14458, N16877);
xor XOR2 (N18910, N18906, N16068);
or OR4 (N18911, N18910, N18083, N4432, N3612);
not NOT1 (N18912, N18908);
xor XOR2 (N18913, N18891, N8384);
not NOT1 (N18914, N18909);
not NOT1 (N18915, N18912);
xor XOR2 (N18916, N18914, N7484);
xor XOR2 (N18917, N18911, N10720);
and AND3 (N18918, N18901, N3783, N8482);
and AND4 (N18919, N18907, N8834, N13415, N1958);
and AND4 (N18920, N18918, N15587, N10751, N4173);
xor XOR2 (N18921, N18916, N1913);
nand NAND3 (N18922, N18921, N11320, N15920);
not NOT1 (N18923, N18917);
buf BUF1 (N18924, N18878);
or OR4 (N18925, N18893, N1924, N16107, N5754);
or OR4 (N18926, N18887, N16221, N7898, N6308);
buf BUF1 (N18927, N18924);
buf BUF1 (N18928, N18913);
xor XOR2 (N18929, N18915, N5912);
buf BUF1 (N18930, N18928);
xor XOR2 (N18931, N18926, N9145);
nand NAND2 (N18932, N18927, N15553);
or OR3 (N18933, N18931, N5800, N7703);
nor NOR4 (N18934, N18930, N16291, N9864, N1912);
and AND3 (N18935, N18934, N7759, N10357);
and AND4 (N18936, N18929, N7751, N850, N4777);
xor XOR2 (N18937, N18920, N14061);
or OR3 (N18938, N18933, N13949, N4727);
and AND2 (N18939, N18938, N5231);
or OR3 (N18940, N18935, N15444, N13537);
xor XOR2 (N18941, N18939, N8856);
nor NOR3 (N18942, N18937, N13397, N15075);
nor NOR3 (N18943, N18923, N9081, N11569);
xor XOR2 (N18944, N18925, N2815);
or OR3 (N18945, N18919, N16952, N1112);
nor NOR2 (N18946, N18940, N17309);
nor NOR4 (N18947, N18941, N18200, N7805, N13807);
not NOT1 (N18948, N18897);
buf BUF1 (N18949, N18942);
xor XOR2 (N18950, N18922, N5133);
or OR2 (N18951, N18945, N7031);
not NOT1 (N18952, N18943);
xor XOR2 (N18953, N18949, N16775);
buf BUF1 (N18954, N18932);
not NOT1 (N18955, N18947);
nand NAND3 (N18956, N18953, N14033, N8274);
xor XOR2 (N18957, N18944, N7949);
not NOT1 (N18958, N18955);
buf BUF1 (N18959, N18952);
not NOT1 (N18960, N18954);
nand NAND3 (N18961, N18950, N987, N7689);
and AND2 (N18962, N18961, N2055);
xor XOR2 (N18963, N18951, N6630);
not NOT1 (N18964, N18958);
xor XOR2 (N18965, N18948, N16430);
xor XOR2 (N18966, N18959, N2471);
xor XOR2 (N18967, N18936, N7515);
or OR3 (N18968, N18963, N6795, N2131);
buf BUF1 (N18969, N18966);
nor NOR4 (N18970, N18967, N1939, N7285, N10638);
nor NOR4 (N18971, N18956, N17536, N12406, N16427);
xor XOR2 (N18972, N18946, N7167);
xor XOR2 (N18973, N18971, N12867);
nand NAND4 (N18974, N18968, N12119, N16141, N13461);
nand NAND2 (N18975, N18970, N7543);
nor NOR4 (N18976, N18957, N1816, N5121, N1351);
or OR4 (N18977, N18973, N7185, N1752, N9852);
buf BUF1 (N18978, N18976);
buf BUF1 (N18979, N18974);
nand NAND3 (N18980, N18979, N14470, N8391);
buf BUF1 (N18981, N18975);
buf BUF1 (N18982, N18964);
and AND3 (N18983, N18962, N16198, N14793);
nand NAND2 (N18984, N18980, N2090);
nand NAND4 (N18985, N18978, N6649, N10065, N6311);
not NOT1 (N18986, N18981);
and AND4 (N18987, N18972, N14018, N11536, N7057);
nor NOR4 (N18988, N18977, N1428, N7283, N18533);
buf BUF1 (N18989, N18969);
or OR4 (N18990, N18984, N224, N3685, N12138);
nor NOR2 (N18991, N18990, N8755);
or OR3 (N18992, N18965, N456, N2021);
buf BUF1 (N18993, N18983);
nand NAND4 (N18994, N18987, N7748, N8344, N1439);
xor XOR2 (N18995, N18989, N13928);
and AND4 (N18996, N18992, N394, N14877, N11546);
buf BUF1 (N18997, N18985);
buf BUF1 (N18998, N18991);
nand NAND2 (N18999, N18998, N5518);
not NOT1 (N19000, N18999);
buf BUF1 (N19001, N18997);
or OR3 (N19002, N19000, N18827, N2959);
and AND4 (N19003, N19002, N13476, N15802, N1754);
and AND3 (N19004, N18986, N3749, N12660);
not NOT1 (N19005, N18995);
and AND3 (N19006, N19003, N9893, N13680);
nor NOR3 (N19007, N19001, N13884, N427);
and AND2 (N19008, N18988, N8319);
or OR4 (N19009, N18960, N14785, N14366, N3160);
buf BUF1 (N19010, N18982);
nand NAND3 (N19011, N19007, N12047, N17643);
nor NOR4 (N19012, N19010, N7192, N8452, N18928);
not NOT1 (N19013, N18993);
xor XOR2 (N19014, N19012, N14757);
buf BUF1 (N19015, N19011);
xor XOR2 (N19016, N19008, N15999);
buf BUF1 (N19017, N19015);
buf BUF1 (N19018, N19016);
not NOT1 (N19019, N19017);
and AND2 (N19020, N18996, N13427);
and AND4 (N19021, N19014, N9307, N13627, N4312);
and AND3 (N19022, N19006, N9621, N2381);
xor XOR2 (N19023, N19013, N11577);
and AND2 (N19024, N18994, N15696);
buf BUF1 (N19025, N19022);
not NOT1 (N19026, N19005);
nor NOR4 (N19027, N19020, N1929, N3588, N4171);
nand NAND3 (N19028, N19018, N12657, N1869);
xor XOR2 (N19029, N19004, N14964);
nand NAND2 (N19030, N19021, N10918);
buf BUF1 (N19031, N19030);
buf BUF1 (N19032, N19025);
xor XOR2 (N19033, N19024, N12878);
not NOT1 (N19034, N19029);
xor XOR2 (N19035, N19027, N4711);
xor XOR2 (N19036, N19035, N4282);
buf BUF1 (N19037, N19023);
and AND4 (N19038, N19019, N3771, N14708, N6671);
buf BUF1 (N19039, N19032);
or OR4 (N19040, N19031, N3200, N6451, N15077);
and AND4 (N19041, N19033, N1145, N12944, N11878);
nor NOR3 (N19042, N19037, N8505, N4288);
nand NAND4 (N19043, N19009, N12538, N11799, N9274);
nor NOR3 (N19044, N19042, N3259, N4174);
nand NAND2 (N19045, N19036, N5319);
buf BUF1 (N19046, N19039);
nor NOR4 (N19047, N19044, N10969, N11450, N11011);
nand NAND4 (N19048, N19034, N5612, N18812, N12117);
and AND3 (N19049, N19040, N11026, N6917);
buf BUF1 (N19050, N19049);
buf BUF1 (N19051, N19038);
nand NAND2 (N19052, N19046, N1208);
not NOT1 (N19053, N19050);
buf BUF1 (N19054, N19041);
nor NOR3 (N19055, N19026, N17649, N16384);
buf BUF1 (N19056, N19028);
buf BUF1 (N19057, N19048);
and AND4 (N19058, N19051, N4512, N14781, N5475);
and AND2 (N19059, N19053, N13823);
nand NAND3 (N19060, N19047, N9543, N8764);
nand NAND2 (N19061, N19058, N16567);
buf BUF1 (N19062, N19043);
nand NAND4 (N19063, N19045, N1232, N446, N7489);
nor NOR2 (N19064, N19056, N17985);
not NOT1 (N19065, N19064);
xor XOR2 (N19066, N19059, N10586);
buf BUF1 (N19067, N19060);
xor XOR2 (N19068, N19065, N9300);
nand NAND3 (N19069, N19067, N7259, N13424);
and AND3 (N19070, N19069, N2517, N3693);
buf BUF1 (N19071, N19054);
nand NAND4 (N19072, N19057, N1974, N15980, N13685);
and AND3 (N19073, N19061, N2778, N18709);
nor NOR2 (N19074, N19072, N7072);
buf BUF1 (N19075, N19074);
not NOT1 (N19076, N19075);
not NOT1 (N19077, N19062);
or OR4 (N19078, N19076, N1053, N10790, N1425);
and AND4 (N19079, N19078, N13542, N12938, N12896);
and AND2 (N19080, N19079, N13221);
and AND2 (N19081, N19071, N16351);
or OR3 (N19082, N19077, N13627, N1828);
not NOT1 (N19083, N19073);
nor NOR4 (N19084, N19082, N18712, N262, N1221);
nand NAND4 (N19085, N19052, N11184, N7420, N7226);
buf BUF1 (N19086, N19055);
nand NAND3 (N19087, N19063, N10021, N9491);
nor NOR2 (N19088, N19081, N12962);
xor XOR2 (N19089, N19066, N15467);
xor XOR2 (N19090, N19088, N4928);
buf BUF1 (N19091, N19084);
xor XOR2 (N19092, N19087, N13361);
and AND2 (N19093, N19080, N15349);
not NOT1 (N19094, N19092);
xor XOR2 (N19095, N19070, N14482);
buf BUF1 (N19096, N19090);
not NOT1 (N19097, N19096);
nand NAND2 (N19098, N19093, N6851);
nor NOR3 (N19099, N19095, N1552, N10450);
buf BUF1 (N19100, N19097);
nor NOR4 (N19101, N19086, N3238, N2550, N17078);
nand NAND3 (N19102, N19085, N8915, N16008);
not NOT1 (N19103, N19102);
buf BUF1 (N19104, N19083);
not NOT1 (N19105, N19101);
xor XOR2 (N19106, N19098, N18743);
or OR4 (N19107, N19068, N8835, N17951, N3727);
buf BUF1 (N19108, N19091);
and AND2 (N19109, N19108, N4649);
not NOT1 (N19110, N19103);
not NOT1 (N19111, N19107);
nand NAND3 (N19112, N19089, N1187, N728);
and AND3 (N19113, N19109, N18605, N16223);
or OR4 (N19114, N19104, N18781, N17581, N16081);
and AND3 (N19115, N19112, N4564, N18796);
and AND2 (N19116, N19099, N9819);
nor NOR2 (N19117, N19105, N4957);
buf BUF1 (N19118, N19110);
xor XOR2 (N19119, N19113, N12954);
or OR2 (N19120, N19117, N11374);
and AND4 (N19121, N19100, N17739, N7372, N8058);
and AND3 (N19122, N19106, N13441, N18715);
xor XOR2 (N19123, N19111, N3329);
not NOT1 (N19124, N19121);
buf BUF1 (N19125, N19120);
or OR4 (N19126, N19118, N113, N16547, N14582);
nor NOR4 (N19127, N19115, N10838, N7073, N14972);
nor NOR4 (N19128, N19126, N11047, N18627, N14890);
xor XOR2 (N19129, N19124, N4406);
xor XOR2 (N19130, N19128, N3784);
buf BUF1 (N19131, N19130);
not NOT1 (N19132, N19119);
nand NAND4 (N19133, N19127, N15417, N10900, N4933);
xor XOR2 (N19134, N19131, N17410);
not NOT1 (N19135, N19133);
or OR3 (N19136, N19114, N5547, N5136);
nand NAND4 (N19137, N19094, N14835, N16244, N6659);
nor NOR2 (N19138, N19122, N11245);
nor NOR3 (N19139, N19116, N2424, N3608);
not NOT1 (N19140, N19137);
and AND3 (N19141, N19134, N10518, N18267);
not NOT1 (N19142, N19138);
xor XOR2 (N19143, N19129, N11785);
or OR4 (N19144, N19125, N9055, N16431, N9085);
nor NOR4 (N19145, N19123, N2299, N8047, N4458);
or OR4 (N19146, N19141, N14917, N8546, N17608);
xor XOR2 (N19147, N19139, N16715);
nor NOR3 (N19148, N19136, N2371, N14561);
not NOT1 (N19149, N19140);
xor XOR2 (N19150, N19132, N8348);
or OR4 (N19151, N19144, N321, N2008, N6525);
xor XOR2 (N19152, N19142, N14065);
nand NAND4 (N19153, N19150, N12457, N7307, N8648);
xor XOR2 (N19154, N19152, N7806);
not NOT1 (N19155, N19154);
and AND3 (N19156, N19147, N18078, N9304);
nand NAND2 (N19157, N19145, N7088);
not NOT1 (N19158, N19143);
xor XOR2 (N19159, N19135, N14040);
and AND2 (N19160, N19159, N18241);
or OR3 (N19161, N19149, N267, N11508);
xor XOR2 (N19162, N19158, N5979);
nor NOR4 (N19163, N19160, N12049, N8538, N18019);
buf BUF1 (N19164, N19162);
nor NOR3 (N19165, N19151, N4572, N6970);
or OR2 (N19166, N19163, N18177);
buf BUF1 (N19167, N19161);
buf BUF1 (N19168, N19167);
or OR2 (N19169, N19146, N8227);
and AND3 (N19170, N19155, N7914, N10872);
xor XOR2 (N19171, N19156, N13089);
and AND2 (N19172, N19166, N17952);
nand NAND3 (N19173, N19170, N16319, N12932);
buf BUF1 (N19174, N19165);
not NOT1 (N19175, N19157);
not NOT1 (N19176, N19171);
xor XOR2 (N19177, N19176, N1063);
or OR4 (N19178, N19177, N11592, N3233, N3023);
xor XOR2 (N19179, N19174, N17792);
not NOT1 (N19180, N19173);
nor NOR4 (N19181, N19180, N5715, N11200, N18666);
buf BUF1 (N19182, N19169);
not NOT1 (N19183, N19175);
and AND4 (N19184, N19172, N17154, N4875, N7185);
nand NAND2 (N19185, N19168, N7460);
or OR4 (N19186, N19164, N18838, N4903, N10009);
and AND2 (N19187, N19148, N9434);
not NOT1 (N19188, N19181);
xor XOR2 (N19189, N19187, N14918);
nor NOR3 (N19190, N19184, N7332, N988);
buf BUF1 (N19191, N19189);
xor XOR2 (N19192, N19183, N11441);
buf BUF1 (N19193, N19179);
or OR2 (N19194, N19185, N17177);
nor NOR4 (N19195, N19188, N8013, N15395, N4922);
not NOT1 (N19196, N19195);
nand NAND4 (N19197, N19192, N15972, N15942, N13797);
xor XOR2 (N19198, N19196, N16656);
and AND2 (N19199, N19182, N12539);
nor NOR2 (N19200, N19191, N1484);
or OR3 (N19201, N19200, N19151, N3366);
not NOT1 (N19202, N19194);
nand NAND2 (N19203, N19178, N9280);
nand NAND2 (N19204, N19193, N13246);
and AND2 (N19205, N19201, N631);
nand NAND4 (N19206, N19197, N13224, N11399, N3763);
and AND3 (N19207, N19186, N17218, N3804);
or OR3 (N19208, N19205, N12699, N11621);
buf BUF1 (N19209, N19198);
nand NAND2 (N19210, N19207, N7662);
and AND3 (N19211, N19190, N6670, N1471);
not NOT1 (N19212, N19210);
xor XOR2 (N19213, N19212, N19105);
and AND2 (N19214, N19206, N518);
and AND4 (N19215, N19204, N13340, N6793, N2054);
or OR4 (N19216, N19209, N17774, N2976, N12932);
and AND2 (N19217, N19215, N6193);
not NOT1 (N19218, N19202);
nor NOR3 (N19219, N19203, N14545, N13216);
nand NAND3 (N19220, N19214, N4893, N5336);
nand NAND3 (N19221, N19208, N16470, N2870);
nand NAND4 (N19222, N19199, N18146, N17883, N2162);
nand NAND2 (N19223, N19153, N9807);
xor XOR2 (N19224, N19223, N12780);
nor NOR3 (N19225, N19221, N3098, N4445);
nand NAND4 (N19226, N19217, N15886, N1934, N13521);
or OR4 (N19227, N19225, N11200, N11142, N386);
xor XOR2 (N19228, N19227, N238);
buf BUF1 (N19229, N19219);
and AND2 (N19230, N19213, N16933);
and AND2 (N19231, N19226, N9133);
not NOT1 (N19232, N19228);
buf BUF1 (N19233, N19224);
xor XOR2 (N19234, N19231, N8782);
nor NOR2 (N19235, N19222, N14708);
not NOT1 (N19236, N19220);
nor NOR4 (N19237, N19211, N2491, N16982, N13990);
not NOT1 (N19238, N19237);
or OR2 (N19239, N19238, N5647);
nor NOR3 (N19240, N19216, N8793, N10206);
and AND2 (N19241, N19235, N17596);
nor NOR4 (N19242, N19239, N14415, N9652, N489);
buf BUF1 (N19243, N19218);
buf BUF1 (N19244, N19233);
nand NAND3 (N19245, N19240, N9077, N17986);
nand NAND2 (N19246, N19234, N17342);
xor XOR2 (N19247, N19241, N6802);
nor NOR3 (N19248, N19247, N10760, N16779);
nor NOR3 (N19249, N19232, N5332, N16007);
xor XOR2 (N19250, N19236, N4630);
or OR3 (N19251, N19248, N3961, N15116);
or OR4 (N19252, N19243, N10123, N8668, N13887);
nand NAND2 (N19253, N19242, N4694);
nand NAND2 (N19254, N19253, N13219);
or OR4 (N19255, N19250, N11708, N4979, N13139);
not NOT1 (N19256, N19255);
and AND4 (N19257, N19244, N2271, N4152, N5035);
not NOT1 (N19258, N19251);
nand NAND4 (N19259, N19229, N16184, N11316, N1236);
buf BUF1 (N19260, N19259);
buf BUF1 (N19261, N19246);
nand NAND2 (N19262, N19230, N3758);
or OR2 (N19263, N19260, N12022);
buf BUF1 (N19264, N19245);
xor XOR2 (N19265, N19261, N14432);
buf BUF1 (N19266, N19254);
xor XOR2 (N19267, N19262, N19153);
buf BUF1 (N19268, N19258);
buf BUF1 (N19269, N19266);
and AND2 (N19270, N19264, N8901);
nand NAND4 (N19271, N19269, N4652, N12966, N1924);
xor XOR2 (N19272, N19256, N2649);
buf BUF1 (N19273, N19270);
not NOT1 (N19274, N19267);
or OR4 (N19275, N19273, N13704, N19117, N3085);
not NOT1 (N19276, N19268);
or OR4 (N19277, N19276, N1056, N8316, N5988);
xor XOR2 (N19278, N19277, N8393);
xor XOR2 (N19279, N19278, N8511);
or OR2 (N19280, N19272, N7623);
or OR2 (N19281, N19274, N16002);
buf BUF1 (N19282, N19265);
buf BUF1 (N19283, N19257);
nor NOR3 (N19284, N19252, N9022, N9213);
not NOT1 (N19285, N19263);
buf BUF1 (N19286, N19249);
not NOT1 (N19287, N19271);
nand NAND3 (N19288, N19283, N3074, N10032);
not NOT1 (N19289, N19281);
and AND3 (N19290, N19275, N8643, N13015);
xor XOR2 (N19291, N19286, N2336);
and AND3 (N19292, N19280, N4657, N17013);
or OR2 (N19293, N19282, N4879);
nand NAND3 (N19294, N19279, N11948, N11146);
nor NOR3 (N19295, N19285, N5131, N13250);
and AND3 (N19296, N19290, N5465, N2778);
or OR3 (N19297, N19293, N4154, N2349);
and AND3 (N19298, N19287, N2011, N17283);
and AND4 (N19299, N19298, N13620, N19249, N17125);
or OR3 (N19300, N19292, N15810, N13347);
nor NOR2 (N19301, N19294, N1299);
not NOT1 (N19302, N19291);
buf BUF1 (N19303, N19302);
buf BUF1 (N19304, N19284);
not NOT1 (N19305, N19303);
buf BUF1 (N19306, N19305);
nor NOR3 (N19307, N19297, N18121, N4926);
not NOT1 (N19308, N19306);
nor NOR3 (N19309, N19295, N7854, N17200);
not NOT1 (N19310, N19296);
buf BUF1 (N19311, N19288);
nor NOR3 (N19312, N19310, N7628, N10049);
or OR2 (N19313, N19301, N3713);
nand NAND2 (N19314, N19289, N6682);
or OR4 (N19315, N19311, N12631, N7416, N8611);
and AND3 (N19316, N19304, N16118, N15163);
nor NOR3 (N19317, N19315, N15046, N15283);
or OR4 (N19318, N19299, N9765, N2060, N2304);
not NOT1 (N19319, N19313);
buf BUF1 (N19320, N19319);
nor NOR4 (N19321, N19318, N3599, N14125, N4099);
nand NAND3 (N19322, N19307, N8525, N14849);
buf BUF1 (N19323, N19317);
buf BUF1 (N19324, N19312);
or OR4 (N19325, N19309, N14413, N3254, N11555);
nand NAND4 (N19326, N19325, N1625, N10211, N1729);
or OR3 (N19327, N19324, N5956, N10067);
buf BUF1 (N19328, N19327);
not NOT1 (N19329, N19321);
nand NAND4 (N19330, N19326, N2130, N3870, N15738);
and AND2 (N19331, N19330, N16076);
nand NAND2 (N19332, N19314, N9616);
not NOT1 (N19333, N19316);
or OR2 (N19334, N19308, N18602);
buf BUF1 (N19335, N19323);
nor NOR2 (N19336, N19300, N19088);
buf BUF1 (N19337, N19336);
and AND3 (N19338, N19331, N13667, N8742);
not NOT1 (N19339, N19322);
or OR3 (N19340, N19329, N16794, N1069);
and AND3 (N19341, N19333, N14049, N15517);
nor NOR2 (N19342, N19335, N18699);
xor XOR2 (N19343, N19328, N6920);
and AND3 (N19344, N19339, N3290, N13569);
and AND4 (N19345, N19343, N11300, N19272, N3730);
xor XOR2 (N19346, N19337, N12513);
and AND2 (N19347, N19344, N18838);
nor NOR4 (N19348, N19341, N18414, N11687, N24);
nand NAND2 (N19349, N19348, N714);
nor NOR4 (N19350, N19346, N3532, N5061, N437);
nand NAND2 (N19351, N19332, N19210);
xor XOR2 (N19352, N19345, N10505);
not NOT1 (N19353, N19350);
nand NAND3 (N19354, N19334, N7967, N5943);
buf BUF1 (N19355, N19351);
and AND4 (N19356, N19320, N5595, N4285, N15253);
nor NOR3 (N19357, N19349, N3758, N19113);
buf BUF1 (N19358, N19354);
nand NAND4 (N19359, N19342, N261, N18113, N12016);
xor XOR2 (N19360, N19358, N17042);
or OR3 (N19361, N19352, N5915, N7868);
xor XOR2 (N19362, N19360, N1448);
nor NOR4 (N19363, N19338, N4992, N8743, N5705);
nor NOR4 (N19364, N19362, N18970, N12835, N18177);
or OR3 (N19365, N19363, N4630, N13942);
buf BUF1 (N19366, N19347);
not NOT1 (N19367, N19357);
or OR2 (N19368, N19365, N5879);
buf BUF1 (N19369, N19367);
nand NAND2 (N19370, N19364, N15397);
nand NAND3 (N19371, N19356, N1123, N18444);
xor XOR2 (N19372, N19355, N18959);
buf BUF1 (N19373, N19369);
not NOT1 (N19374, N19340);
nor NOR4 (N19375, N19361, N17675, N4325, N8992);
nor NOR4 (N19376, N19374, N11897, N2254, N8573);
not NOT1 (N19377, N19368);
buf BUF1 (N19378, N19377);
not NOT1 (N19379, N19353);
and AND4 (N19380, N19359, N8889, N11495, N2350);
buf BUF1 (N19381, N19373);
and AND2 (N19382, N19378, N5987);
buf BUF1 (N19383, N19371);
not NOT1 (N19384, N19382);
buf BUF1 (N19385, N19376);
xor XOR2 (N19386, N19370, N1083);
or OR2 (N19387, N19372, N10287);
nor NOR4 (N19388, N19385, N3090, N10086, N18277);
not NOT1 (N19389, N19387);
nor NOR3 (N19390, N19379, N16967, N16904);
nor NOR3 (N19391, N19384, N3131, N4242);
and AND2 (N19392, N19381, N9774);
and AND2 (N19393, N19391, N9867);
nor NOR3 (N19394, N19393, N13282, N10681);
and AND4 (N19395, N19380, N9688, N2607, N4299);
nor NOR4 (N19396, N19388, N11708, N17467, N13937);
xor XOR2 (N19397, N19396, N11352);
or OR4 (N19398, N19375, N3265, N848, N12069);
and AND4 (N19399, N19398, N1059, N10773, N5002);
buf BUF1 (N19400, N19392);
nand NAND4 (N19401, N19390, N404, N4762, N4482);
buf BUF1 (N19402, N19389);
or OR3 (N19403, N19366, N17994, N17760);
not NOT1 (N19404, N19395);
nor NOR3 (N19405, N19394, N18489, N15793);
or OR2 (N19406, N19401, N3287);
nor NOR3 (N19407, N19400, N3116, N5253);
nor NOR3 (N19408, N19405, N886, N1631);
xor XOR2 (N19409, N19404, N11562);
not NOT1 (N19410, N19408);
or OR2 (N19411, N19406, N5124);
and AND3 (N19412, N19383, N6410, N16160);
buf BUF1 (N19413, N19407);
or OR3 (N19414, N19409, N12531, N17674);
xor XOR2 (N19415, N19403, N13766);
and AND2 (N19416, N19414, N17595);
nor NOR4 (N19417, N19410, N14117, N1785, N15287);
not NOT1 (N19418, N19416);
xor XOR2 (N19419, N19402, N19128);
xor XOR2 (N19420, N19415, N11495);
xor XOR2 (N19421, N19413, N5482);
nand NAND3 (N19422, N19399, N6400, N6060);
xor XOR2 (N19423, N19412, N18357);
nor NOR3 (N19424, N19422, N9256, N16876);
buf BUF1 (N19425, N19417);
not NOT1 (N19426, N19420);
buf BUF1 (N19427, N19423);
xor XOR2 (N19428, N19426, N1947);
nand NAND2 (N19429, N19428, N19012);
buf BUF1 (N19430, N19397);
nand NAND4 (N19431, N19421, N15887, N13022, N7481);
not NOT1 (N19432, N19425);
and AND2 (N19433, N19427, N9272);
xor XOR2 (N19434, N19419, N7935);
not NOT1 (N19435, N19429);
nor NOR3 (N19436, N19433, N15624, N10919);
nor NOR3 (N19437, N19424, N16152, N2885);
xor XOR2 (N19438, N19431, N12252);
not NOT1 (N19439, N19430);
buf BUF1 (N19440, N19434);
nand NAND3 (N19441, N19435, N16742, N11187);
and AND3 (N19442, N19436, N14074, N326);
or OR3 (N19443, N19437, N14171, N7813);
nand NAND4 (N19444, N19439, N12179, N13991, N6667);
nand NAND3 (N19445, N19418, N12849, N841);
xor XOR2 (N19446, N19444, N7274);
nand NAND2 (N19447, N19432, N2421);
nand NAND4 (N19448, N19445, N264, N5113, N12665);
and AND4 (N19449, N19442, N18141, N5075, N5278);
nand NAND4 (N19450, N19446, N9680, N8723, N12287);
or OR2 (N19451, N19440, N8715);
or OR2 (N19452, N19451, N15188);
buf BUF1 (N19453, N19448);
not NOT1 (N19454, N19438);
and AND3 (N19455, N19447, N640, N8567);
nor NOR2 (N19456, N19450, N3456);
nor NOR4 (N19457, N19449, N13511, N16894, N5279);
not NOT1 (N19458, N19457);
not NOT1 (N19459, N19441);
xor XOR2 (N19460, N19386, N1702);
and AND3 (N19461, N19411, N5019, N12259);
nand NAND3 (N19462, N19460, N9817, N10829);
buf BUF1 (N19463, N19454);
buf BUF1 (N19464, N19455);
nand NAND2 (N19465, N19453, N15468);
nor NOR2 (N19466, N19452, N4462);
nand NAND4 (N19467, N19465, N18831, N4348, N13933);
buf BUF1 (N19468, N19456);
buf BUF1 (N19469, N19443);
nor NOR2 (N19470, N19462, N3278);
or OR2 (N19471, N19467, N16938);
nor NOR2 (N19472, N19459, N19140);
xor XOR2 (N19473, N19463, N17893);
and AND4 (N19474, N19472, N4741, N9511, N15305);
and AND3 (N19475, N19473, N13676, N14818);
nand NAND4 (N19476, N19468, N7137, N16980, N10242);
and AND2 (N19477, N19476, N14578);
buf BUF1 (N19478, N19470);
and AND3 (N19479, N19469, N11730, N3994);
buf BUF1 (N19480, N19478);
or OR3 (N19481, N19458, N19320, N14649);
or OR4 (N19482, N19474, N14281, N1195, N2456);
and AND4 (N19483, N19477, N5151, N1482, N6700);
xor XOR2 (N19484, N19466, N15528);
nand NAND3 (N19485, N19461, N13627, N17802);
xor XOR2 (N19486, N19481, N3868);
not NOT1 (N19487, N19484);
not NOT1 (N19488, N19486);
not NOT1 (N19489, N19475);
nand NAND3 (N19490, N19471, N16738, N6386);
nand NAND4 (N19491, N19485, N14501, N15938, N6493);
or OR4 (N19492, N19464, N14473, N15222, N14210);
or OR4 (N19493, N19491, N10754, N18495, N8435);
xor XOR2 (N19494, N19487, N8913);
xor XOR2 (N19495, N19482, N2515);
xor XOR2 (N19496, N19495, N17427);
or OR2 (N19497, N19494, N3345);
or OR2 (N19498, N19483, N13852);
buf BUF1 (N19499, N19493);
not NOT1 (N19500, N19479);
buf BUF1 (N19501, N19480);
and AND4 (N19502, N19501, N6212, N17472, N9976);
not NOT1 (N19503, N19500);
and AND3 (N19504, N19498, N3044, N8875);
buf BUF1 (N19505, N19490);
or OR4 (N19506, N19488, N13229, N2244, N19156);
not NOT1 (N19507, N19503);
and AND4 (N19508, N19496, N7061, N13213, N14635);
nor NOR3 (N19509, N19508, N7046, N622);
and AND3 (N19510, N19499, N2075, N6779);
xor XOR2 (N19511, N19510, N5203);
nor NOR3 (N19512, N19506, N19444, N11248);
nand NAND4 (N19513, N19509, N5046, N6264, N3998);
xor XOR2 (N19514, N19507, N9294);
xor XOR2 (N19515, N19513, N16445);
nor NOR3 (N19516, N19502, N30, N5769);
nand NAND4 (N19517, N19512, N6471, N16539, N2177);
not NOT1 (N19518, N19511);
and AND2 (N19519, N19517, N1758);
nor NOR4 (N19520, N19505, N3671, N18251, N2205);
and AND2 (N19521, N19516, N6943);
xor XOR2 (N19522, N19489, N14736);
or OR3 (N19523, N19518, N8074, N8212);
buf BUF1 (N19524, N19492);
nor NOR3 (N19525, N19524, N6442, N4795);
and AND3 (N19526, N19522, N14349, N18578);
nor NOR3 (N19527, N19520, N12024, N7840);
nor NOR2 (N19528, N19521, N7239);
buf BUF1 (N19529, N19527);
nor NOR4 (N19530, N19523, N14423, N7744, N7284);
buf BUF1 (N19531, N19529);
nand NAND4 (N19532, N19504, N2514, N16716, N1426);
or OR2 (N19533, N19497, N8053);
buf BUF1 (N19534, N19531);
nor NOR4 (N19535, N19519, N9648, N7281, N8300);
nor NOR3 (N19536, N19515, N669, N787);
nor NOR2 (N19537, N19533, N1777);
and AND3 (N19538, N19514, N15399, N2932);
not NOT1 (N19539, N19534);
xor XOR2 (N19540, N19530, N10483);
or OR2 (N19541, N19538, N9232);
and AND3 (N19542, N19532, N12539, N9598);
not NOT1 (N19543, N19540);
nor NOR3 (N19544, N19528, N14943, N6461);
nand NAND2 (N19545, N19535, N17544);
xor XOR2 (N19546, N19543, N4364);
xor XOR2 (N19547, N19546, N8485);
nand NAND3 (N19548, N19526, N17804, N571);
buf BUF1 (N19549, N19548);
buf BUF1 (N19550, N19539);
not NOT1 (N19551, N19525);
buf BUF1 (N19552, N19545);
and AND4 (N19553, N19541, N18998, N1227, N10805);
nor NOR3 (N19554, N19550, N14412, N13696);
and AND4 (N19555, N19552, N4388, N3070, N4047);
not NOT1 (N19556, N19537);
not NOT1 (N19557, N19554);
buf BUF1 (N19558, N19553);
nand NAND3 (N19559, N19558, N16148, N13998);
buf BUF1 (N19560, N19557);
xor XOR2 (N19561, N19547, N9265);
and AND3 (N19562, N19549, N17220, N11304);
nand NAND2 (N19563, N19542, N16733);
nand NAND2 (N19564, N19536, N8707);
xor XOR2 (N19565, N19556, N9226);
not NOT1 (N19566, N19555);
not NOT1 (N19567, N19559);
or OR2 (N19568, N19560, N1230);
and AND4 (N19569, N19544, N13690, N11505, N4074);
or OR3 (N19570, N19563, N7070, N12950);
xor XOR2 (N19571, N19564, N1332);
nand NAND4 (N19572, N19570, N3618, N9424, N12961);
not NOT1 (N19573, N19562);
xor XOR2 (N19574, N19572, N4891);
nor NOR2 (N19575, N19551, N5393);
xor XOR2 (N19576, N19575, N6695);
buf BUF1 (N19577, N19565);
xor XOR2 (N19578, N19574, N2716);
and AND4 (N19579, N19561, N12034, N6501, N10996);
or OR4 (N19580, N19569, N1546, N6679, N4410);
buf BUF1 (N19581, N19577);
and AND4 (N19582, N19576, N3946, N6939, N13413);
nor NOR4 (N19583, N19580, N6091, N1161, N2079);
or OR3 (N19584, N19578, N15750, N19288);
xor XOR2 (N19585, N19584, N942);
nand NAND3 (N19586, N19582, N410, N10407);
or OR2 (N19587, N19583, N6865);
not NOT1 (N19588, N19566);
and AND2 (N19589, N19581, N17367);
nor NOR4 (N19590, N19589, N18479, N9387, N8250);
nor NOR3 (N19591, N19590, N7076, N13644);
and AND3 (N19592, N19573, N10024, N14046);
or OR4 (N19593, N19579, N13937, N4563, N11044);
xor XOR2 (N19594, N19571, N17413);
and AND2 (N19595, N19592, N9586);
or OR2 (N19596, N19568, N1073);
and AND3 (N19597, N19593, N19299, N13747);
nand NAND4 (N19598, N19591, N6351, N5955, N9275);
nand NAND4 (N19599, N19596, N3751, N18231, N9823);
and AND2 (N19600, N19587, N18576);
buf BUF1 (N19601, N19594);
xor XOR2 (N19602, N19567, N7821);
xor XOR2 (N19603, N19595, N14491);
nor NOR2 (N19604, N19597, N7625);
xor XOR2 (N19605, N19585, N14677);
nor NOR4 (N19606, N19588, N1562, N1467, N12426);
or OR3 (N19607, N19603, N17117, N18630);
buf BUF1 (N19608, N19598);
not NOT1 (N19609, N19604);
or OR2 (N19610, N19608, N13588);
nor NOR3 (N19611, N19610, N9821, N14267);
nand NAND2 (N19612, N19611, N2569);
and AND2 (N19613, N19607, N14396);
or OR2 (N19614, N19613, N6740);
not NOT1 (N19615, N19602);
or OR2 (N19616, N19614, N12439);
nand NAND3 (N19617, N19615, N11575, N561);
or OR3 (N19618, N19606, N11952, N15846);
nor NOR4 (N19619, N19612, N18696, N8044, N7596);
xor XOR2 (N19620, N19609, N7218);
nand NAND3 (N19621, N19586, N12783, N14179);
nor NOR4 (N19622, N19599, N17268, N15908, N11331);
nor NOR4 (N19623, N19620, N1815, N1502, N9162);
and AND4 (N19624, N19621, N9868, N8024, N17059);
or OR3 (N19625, N19624, N7509, N19473);
and AND2 (N19626, N19619, N11972);
nor NOR3 (N19627, N19626, N9354, N1921);
not NOT1 (N19628, N19600);
buf BUF1 (N19629, N19623);
nor NOR3 (N19630, N19629, N8107, N16646);
nand NAND4 (N19631, N19630, N13953, N17946, N11619);
or OR2 (N19632, N19622, N16846);
and AND4 (N19633, N19616, N14781, N12304, N18682);
not NOT1 (N19634, N19628);
xor XOR2 (N19635, N19632, N3313);
buf BUF1 (N19636, N19617);
or OR3 (N19637, N19635, N13572, N8398);
or OR2 (N19638, N19636, N6185);
nor NOR4 (N19639, N19618, N5618, N5391, N1047);
xor XOR2 (N19640, N19627, N1134);
or OR4 (N19641, N19638, N12920, N16070, N5052);
xor XOR2 (N19642, N19625, N19455);
nand NAND3 (N19643, N19605, N17447, N3543);
nor NOR4 (N19644, N19641, N18918, N16638, N14363);
buf BUF1 (N19645, N19639);
nand NAND3 (N19646, N19631, N1075, N4664);
nand NAND2 (N19647, N19634, N2547);
buf BUF1 (N19648, N19643);
buf BUF1 (N19649, N19644);
nand NAND4 (N19650, N19601, N8865, N5247, N6158);
not NOT1 (N19651, N19633);
xor XOR2 (N19652, N19640, N6155);
xor XOR2 (N19653, N19647, N16843);
nor NOR2 (N19654, N19646, N19299);
buf BUF1 (N19655, N19650);
not NOT1 (N19656, N19652);
nand NAND3 (N19657, N19642, N5445, N15089);
nor NOR2 (N19658, N19656, N10859);
nand NAND2 (N19659, N19657, N8284);
buf BUF1 (N19660, N19658);
buf BUF1 (N19661, N19654);
or OR3 (N19662, N19651, N2179, N7294);
nor NOR2 (N19663, N19662, N9655);
and AND4 (N19664, N19637, N8824, N1186, N15160);
xor XOR2 (N19665, N19661, N6165);
nand NAND3 (N19666, N19648, N9444, N12199);
and AND3 (N19667, N19655, N8837, N2453);
or OR4 (N19668, N19664, N4148, N6535, N92);
buf BUF1 (N19669, N19668);
or OR2 (N19670, N19665, N1373);
nor NOR4 (N19671, N19667, N1982, N5908, N1523);
or OR4 (N19672, N19645, N17657, N11995, N11196);
and AND3 (N19673, N19672, N15385, N1069);
not NOT1 (N19674, N19666);
or OR4 (N19675, N19669, N13536, N2471, N9339);
or OR2 (N19676, N19659, N7664);
nor NOR3 (N19677, N19675, N7575, N16739);
not NOT1 (N19678, N19670);
or OR2 (N19679, N19660, N7146);
and AND3 (N19680, N19677, N1744, N19018);
buf BUF1 (N19681, N19663);
not NOT1 (N19682, N19674);
or OR3 (N19683, N19671, N17071, N667);
nand NAND3 (N19684, N19653, N10084, N15728);
nand NAND2 (N19685, N19679, N8877);
not NOT1 (N19686, N19685);
buf BUF1 (N19687, N19682);
or OR2 (N19688, N19678, N17033);
or OR3 (N19689, N19688, N3303, N958);
or OR2 (N19690, N19683, N3938);
buf BUF1 (N19691, N19676);
and AND4 (N19692, N19686, N13306, N9361, N6127);
and AND4 (N19693, N19690, N14814, N792, N17937);
or OR3 (N19694, N19681, N9825, N18683);
nand NAND4 (N19695, N19689, N4402, N13312, N9519);
or OR4 (N19696, N19687, N3434, N15850, N16946);
buf BUF1 (N19697, N19695);
xor XOR2 (N19698, N19673, N4807);
or OR3 (N19699, N19697, N13355, N11557);
nand NAND4 (N19700, N19699, N6197, N691, N18595);
nand NAND4 (N19701, N19649, N12368, N524, N6997);
and AND3 (N19702, N19694, N18748, N16705);
buf BUF1 (N19703, N19680);
xor XOR2 (N19704, N19692, N15578);
nor NOR4 (N19705, N19698, N4022, N3059, N15469);
and AND3 (N19706, N19704, N16591, N4868);
nor NOR3 (N19707, N19706, N2249, N15181);
nand NAND3 (N19708, N19705, N374, N9377);
and AND3 (N19709, N19684, N8389, N1199);
or OR2 (N19710, N19691, N3287);
xor XOR2 (N19711, N19701, N8867);
or OR4 (N19712, N19710, N10957, N10967, N15359);
xor XOR2 (N19713, N19693, N5184);
and AND4 (N19714, N19696, N5569, N502, N2384);
xor XOR2 (N19715, N19714, N10748);
not NOT1 (N19716, N19709);
nand NAND4 (N19717, N19708, N14669, N19364, N4767);
not NOT1 (N19718, N19713);
buf BUF1 (N19719, N19702);
buf BUF1 (N19720, N19715);
xor XOR2 (N19721, N19718, N14787);
not NOT1 (N19722, N19720);
xor XOR2 (N19723, N19707, N12780);
nor NOR4 (N19724, N19700, N6651, N19149, N9268);
not NOT1 (N19725, N19716);
and AND4 (N19726, N19721, N16182, N17502, N10483);
or OR3 (N19727, N19726, N630, N3113);
nand NAND4 (N19728, N19719, N7597, N14180, N10513);
buf BUF1 (N19729, N19724);
nor NOR2 (N19730, N19728, N3499);
or OR4 (N19731, N19703, N16693, N6019, N6508);
and AND4 (N19732, N19711, N11709, N1780, N458);
and AND2 (N19733, N19729, N6701);
and AND4 (N19734, N19712, N9797, N14113, N8048);
nand NAND4 (N19735, N19731, N1274, N13951, N1502);
and AND3 (N19736, N19723, N8975, N15543);
not NOT1 (N19737, N19722);
buf BUF1 (N19738, N19725);
xor XOR2 (N19739, N19735, N3183);
not NOT1 (N19740, N19738);
buf BUF1 (N19741, N19736);
and AND2 (N19742, N19740, N4844);
xor XOR2 (N19743, N19741, N12031);
not NOT1 (N19744, N19743);
or OR4 (N19745, N19742, N11926, N1677, N7196);
or OR3 (N19746, N19739, N12300, N9299);
or OR3 (N19747, N19730, N18655, N7446);
nor NOR3 (N19748, N19734, N19156, N3454);
or OR4 (N19749, N19727, N3005, N664, N8978);
or OR3 (N19750, N19737, N14802, N5430);
and AND2 (N19751, N19748, N11238);
xor XOR2 (N19752, N19746, N13345);
xor XOR2 (N19753, N19752, N7189);
not NOT1 (N19754, N19751);
or OR3 (N19755, N19732, N6259, N8577);
nor NOR3 (N19756, N19747, N7929, N17694);
not NOT1 (N19757, N19753);
or OR4 (N19758, N19749, N8703, N17603, N16175);
nand NAND3 (N19759, N19745, N5393, N9522);
and AND2 (N19760, N19757, N3462);
not NOT1 (N19761, N19733);
not NOT1 (N19762, N19759);
nor NOR2 (N19763, N19758, N15185);
nor NOR4 (N19764, N19756, N9093, N6695, N17080);
nor NOR2 (N19765, N19761, N12013);
nand NAND2 (N19766, N19744, N17952);
buf BUF1 (N19767, N19766);
nand NAND3 (N19768, N19754, N10974, N13404);
or OR3 (N19769, N19760, N18928, N13781);
not NOT1 (N19770, N19767);
nor NOR4 (N19771, N19763, N18278, N16483, N3205);
nand NAND2 (N19772, N19770, N12576);
and AND2 (N19773, N19769, N17709);
buf BUF1 (N19774, N19762);
not NOT1 (N19775, N19768);
nand NAND3 (N19776, N19773, N4592, N10041);
nand NAND2 (N19777, N19765, N2947);
xor XOR2 (N19778, N19771, N6633);
or OR3 (N19779, N19717, N10932, N4548);
nor NOR4 (N19780, N19755, N2355, N16736, N8416);
nand NAND3 (N19781, N19764, N6160, N6297);
xor XOR2 (N19782, N19776, N5385);
xor XOR2 (N19783, N19778, N6349);
and AND4 (N19784, N19750, N8161, N10303, N15858);
xor XOR2 (N19785, N19772, N1371);
xor XOR2 (N19786, N19779, N3253);
not NOT1 (N19787, N19782);
nor NOR3 (N19788, N19780, N8449, N15514);
and AND4 (N19789, N19784, N9971, N16237, N7365);
or OR3 (N19790, N19789, N10039, N17309);
or OR4 (N19791, N19790, N19175, N9904, N5008);
or OR4 (N19792, N19781, N8642, N14951, N7603);
nor NOR3 (N19793, N19775, N17429, N16039);
xor XOR2 (N19794, N19783, N15770);
nor NOR3 (N19795, N19793, N1764, N6104);
xor XOR2 (N19796, N19786, N17607);
nand NAND4 (N19797, N19791, N18967, N9935, N3854);
and AND4 (N19798, N19794, N10354, N7027, N766);
nand NAND4 (N19799, N19777, N18732, N1392, N17163);
or OR4 (N19800, N19774, N7373, N9564, N18669);
xor XOR2 (N19801, N19796, N15598);
not NOT1 (N19802, N19787);
or OR3 (N19803, N19802, N1598, N5299);
and AND3 (N19804, N19800, N13144, N1440);
or OR2 (N19805, N19795, N13301);
xor XOR2 (N19806, N19797, N9364);
or OR3 (N19807, N19785, N6180, N3021);
not NOT1 (N19808, N19807);
buf BUF1 (N19809, N19808);
and AND3 (N19810, N19792, N3800, N13660);
nor NOR4 (N19811, N19788, N10029, N6041, N860);
xor XOR2 (N19812, N19805, N3235);
and AND3 (N19813, N19811, N10992, N6084);
nand NAND3 (N19814, N19806, N1869, N6825);
or OR4 (N19815, N19804, N7604, N9971, N16010);
buf BUF1 (N19816, N19798);
buf BUF1 (N19817, N19799);
buf BUF1 (N19818, N19814);
xor XOR2 (N19819, N19815, N17569);
or OR2 (N19820, N19803, N16634);
and AND3 (N19821, N19817, N17496, N3713);
not NOT1 (N19822, N19809);
or OR2 (N19823, N19822, N6283);
nand NAND4 (N19824, N19810, N18680, N8361, N5166);
and AND3 (N19825, N19823, N2944, N486);
nand NAND4 (N19826, N19825, N3461, N9691, N10194);
xor XOR2 (N19827, N19816, N17094);
and AND4 (N19828, N19818, N2385, N2114, N12042);
buf BUF1 (N19829, N19813);
xor XOR2 (N19830, N19827, N7048);
buf BUF1 (N19831, N19824);
xor XOR2 (N19832, N19830, N14810);
nor NOR4 (N19833, N19829, N15725, N3937, N1749);
nand NAND4 (N19834, N19819, N7939, N11665, N17909);
or OR3 (N19835, N19833, N3935, N9548);
xor XOR2 (N19836, N19820, N15665);
or OR4 (N19837, N19831, N3118, N19110, N13035);
nor NOR2 (N19838, N19832, N9130);
not NOT1 (N19839, N19821);
xor XOR2 (N19840, N19828, N6660);
nand NAND2 (N19841, N19840, N1885);
buf BUF1 (N19842, N19837);
nor NOR4 (N19843, N19838, N14434, N19341, N11025);
nor NOR4 (N19844, N19826, N13556, N5734, N8221);
or OR3 (N19845, N19801, N19091, N18308);
nor NOR4 (N19846, N19842, N3168, N17356, N14697);
and AND4 (N19847, N19841, N2371, N2213, N1781);
nor NOR3 (N19848, N19847, N19524, N8452);
nand NAND3 (N19849, N19812, N15498, N9779);
nand NAND4 (N19850, N19849, N2912, N15543, N13743);
xor XOR2 (N19851, N19846, N16939);
nand NAND4 (N19852, N19850, N17085, N15542, N17815);
buf BUF1 (N19853, N19852);
nor NOR2 (N19854, N19843, N3015);
nand NAND3 (N19855, N19834, N4919, N2765);
nand NAND3 (N19856, N19845, N13486, N16613);
and AND3 (N19857, N19856, N15552, N5071);
xor XOR2 (N19858, N19853, N18040);
and AND2 (N19859, N19858, N13002);
or OR2 (N19860, N19844, N3145);
not NOT1 (N19861, N19839);
buf BUF1 (N19862, N19859);
or OR3 (N19863, N19855, N9862, N14553);
or OR2 (N19864, N19851, N8942);
buf BUF1 (N19865, N19857);
not NOT1 (N19866, N19862);
buf BUF1 (N19867, N19863);
and AND4 (N19868, N19864, N5467, N18407, N11376);
nor NOR4 (N19869, N19865, N6494, N5445, N9538);
nor NOR4 (N19870, N19867, N13609, N2504, N8501);
not NOT1 (N19871, N19861);
buf BUF1 (N19872, N19848);
nand NAND4 (N19873, N19836, N9991, N18907, N180);
nor NOR3 (N19874, N19866, N16394, N14224);
nand NAND4 (N19875, N19873, N5445, N8742, N2039);
and AND3 (N19876, N19835, N3524, N15030);
nand NAND2 (N19877, N19854, N4255);
buf BUF1 (N19878, N19876);
nand NAND4 (N19879, N19860, N16235, N9355, N8167);
buf BUF1 (N19880, N19872);
not NOT1 (N19881, N19874);
or OR3 (N19882, N19881, N1317, N1438);
not NOT1 (N19883, N19878);
nand NAND3 (N19884, N19869, N7995, N9087);
not NOT1 (N19885, N19884);
xor XOR2 (N19886, N19880, N6191);
nor NOR2 (N19887, N19886, N2231);
nand NAND3 (N19888, N19887, N19605, N1550);
xor XOR2 (N19889, N19871, N11215);
xor XOR2 (N19890, N19888, N11378);
xor XOR2 (N19891, N19889, N17694);
nand NAND4 (N19892, N19877, N16415, N7260, N7425);
buf BUF1 (N19893, N19868);
nor NOR2 (N19894, N19891, N18225);
xor XOR2 (N19895, N19892, N6508);
nor NOR2 (N19896, N19883, N858);
nor NOR3 (N19897, N19896, N19894, N2964);
or OR3 (N19898, N6285, N13847, N12604);
nand NAND2 (N19899, N19885, N721);
buf BUF1 (N19900, N19895);
not NOT1 (N19901, N19899);
nand NAND4 (N19902, N19898, N17756, N16602, N13736);
buf BUF1 (N19903, N19897);
nand NAND4 (N19904, N19882, N15133, N14985, N1714);
not NOT1 (N19905, N19890);
and AND4 (N19906, N19900, N4488, N598, N17069);
not NOT1 (N19907, N19905);
nand NAND4 (N19908, N19902, N6765, N8356, N13850);
or OR2 (N19909, N19903, N17913);
nand NAND4 (N19910, N19870, N2380, N14197, N9964);
and AND4 (N19911, N19910, N11796, N7670, N5119);
xor XOR2 (N19912, N19901, N16609);
not NOT1 (N19913, N19909);
and AND2 (N19914, N19904, N18190);
and AND2 (N19915, N19908, N4741);
not NOT1 (N19916, N19912);
or OR4 (N19917, N19911, N4414, N7060, N13559);
and AND2 (N19918, N19875, N5234);
nor NOR4 (N19919, N19918, N3041, N18791, N12786);
not NOT1 (N19920, N19916);
buf BUF1 (N19921, N19920);
buf BUF1 (N19922, N19906);
nand NAND4 (N19923, N19917, N17335, N7947, N5998);
nor NOR3 (N19924, N19907, N13837, N167);
not NOT1 (N19925, N19914);
or OR3 (N19926, N19924, N5399, N233);
buf BUF1 (N19927, N19925);
buf BUF1 (N19928, N19923);
nor NOR4 (N19929, N19922, N6150, N17098, N9380);
and AND4 (N19930, N19927, N5495, N1356, N8742);
not NOT1 (N19931, N19921);
xor XOR2 (N19932, N19926, N1389);
not NOT1 (N19933, N19929);
nor NOR3 (N19934, N19915, N6078, N5234);
nor NOR2 (N19935, N19930, N18118);
nand NAND4 (N19936, N19928, N14940, N10141, N15138);
and AND4 (N19937, N19893, N9522, N14480, N14359);
and AND2 (N19938, N19934, N4925);
buf BUF1 (N19939, N19936);
nand NAND2 (N19940, N19879, N17159);
and AND3 (N19941, N19933, N5208, N19465);
not NOT1 (N19942, N19935);
not NOT1 (N19943, N19931);
not NOT1 (N19944, N19919);
xor XOR2 (N19945, N19944, N7793);
xor XOR2 (N19946, N19943, N13802);
nor NOR2 (N19947, N19946, N3003);
or OR2 (N19948, N19942, N13821);
and AND2 (N19949, N19938, N11881);
or OR2 (N19950, N19940, N3208);
not NOT1 (N19951, N19945);
nand NAND4 (N19952, N19950, N16955, N13903, N2703);
xor XOR2 (N19953, N19947, N6275);
not NOT1 (N19954, N19939);
and AND2 (N19955, N19954, N1326);
buf BUF1 (N19956, N19932);
xor XOR2 (N19957, N19956, N6166);
and AND3 (N19958, N19948, N5433, N17705);
and AND4 (N19959, N19941, N16019, N1358, N8982);
nor NOR4 (N19960, N19955, N19704, N16625, N19655);
xor XOR2 (N19961, N19958, N16537);
nor NOR3 (N19962, N19951, N2350, N2641);
xor XOR2 (N19963, N19952, N7909);
nand NAND4 (N19964, N19953, N17538, N18021, N13505);
and AND3 (N19965, N19961, N13114, N17);
nor NOR3 (N19966, N19962, N14478, N8065);
and AND4 (N19967, N19966, N3505, N7784, N13635);
not NOT1 (N19968, N19960);
not NOT1 (N19969, N19913);
buf BUF1 (N19970, N19965);
and AND4 (N19971, N19959, N3242, N7102, N146);
nand NAND4 (N19972, N19937, N3476, N9095, N9221);
xor XOR2 (N19973, N19970, N19067);
xor XOR2 (N19974, N19971, N9630);
not NOT1 (N19975, N19964);
not NOT1 (N19976, N19968);
or OR3 (N19977, N19963, N3617, N2016);
not NOT1 (N19978, N19969);
not NOT1 (N19979, N19949);
nand NAND2 (N19980, N19975, N18748);
buf BUF1 (N19981, N19957);
or OR2 (N19982, N19967, N2653);
xor XOR2 (N19983, N19981, N2913);
or OR2 (N19984, N19977, N8186);
nand NAND3 (N19985, N19976, N12190, N13317);
or OR2 (N19986, N19983, N238);
or OR3 (N19987, N19973, N5530, N13096);
not NOT1 (N19988, N19979);
xor XOR2 (N19989, N19986, N7734);
buf BUF1 (N19990, N19982);
buf BUF1 (N19991, N19972);
xor XOR2 (N19992, N19984, N12561);
or OR3 (N19993, N19974, N13776, N12879);
nor NOR4 (N19994, N19989, N19701, N6732, N9363);
nor NOR2 (N19995, N19994, N11786);
xor XOR2 (N19996, N19990, N1787);
xor XOR2 (N19997, N19987, N7135);
nand NAND2 (N19998, N19980, N17447);
not NOT1 (N19999, N19997);
nor NOR4 (N20000, N19995, N8655, N8735, N4409);
and AND3 (N20001, N19985, N15732, N5065);
and AND2 (N20002, N19996, N7002);
not NOT1 (N20003, N19978);
or OR4 (N20004, N19991, N9075, N13090, N4536);
and AND3 (N20005, N20002, N3977, N13941);
buf BUF1 (N20006, N19992);
or OR3 (N20007, N19998, N14210, N264);
not NOT1 (N20008, N20004);
and AND2 (N20009, N20008, N12451);
nand NAND2 (N20010, N20009, N9826);
nand NAND2 (N20011, N19993, N11754);
nor NOR4 (N20012, N20007, N18532, N5199, N11355);
nor NOR4 (N20013, N20011, N11778, N12114, N7754);
and AND2 (N20014, N20013, N449);
buf BUF1 (N20015, N20006);
xor XOR2 (N20016, N20001, N3094);
nor NOR4 (N20017, N20000, N15314, N1974, N11606);
not NOT1 (N20018, N20015);
buf BUF1 (N20019, N19999);
buf BUF1 (N20020, N20003);
buf BUF1 (N20021, N20018);
nor NOR2 (N20022, N19988, N17836);
xor XOR2 (N20023, N20005, N11759);
xor XOR2 (N20024, N20023, N7227);
nor NOR3 (N20025, N20021, N7987, N10699);
xor XOR2 (N20026, N20014, N17765);
or OR4 (N20027, N20020, N6615, N7585, N19230);
xor XOR2 (N20028, N20012, N17405);
xor XOR2 (N20029, N20010, N7392);
or OR2 (N20030, N20024, N2875);
nor NOR2 (N20031, N20019, N6623);
nor NOR4 (N20032, N20027, N14961, N14998, N662);
nor NOR4 (N20033, N20028, N7329, N13510, N10009);
nor NOR3 (N20034, N20029, N4820, N7361);
buf BUF1 (N20035, N20017);
xor XOR2 (N20036, N20035, N17986);
or OR2 (N20037, N20033, N789);
buf BUF1 (N20038, N20025);
and AND4 (N20039, N20034, N7232, N220, N15413);
xor XOR2 (N20040, N20036, N19712);
nand NAND3 (N20041, N20022, N12501, N19463);
nand NAND3 (N20042, N20032, N13811, N5096);
not NOT1 (N20043, N20030);
not NOT1 (N20044, N20037);
nand NAND4 (N20045, N20040, N17200, N363, N760);
xor XOR2 (N20046, N20042, N16212);
nor NOR3 (N20047, N20044, N15237, N3353);
and AND4 (N20048, N20041, N16296, N19416, N12118);
and AND2 (N20049, N20026, N13310);
nand NAND4 (N20050, N20045, N3982, N12514, N12805);
nor NOR2 (N20051, N20039, N13085);
xor XOR2 (N20052, N20043, N14455);
xor XOR2 (N20053, N20031, N16086);
nor NOR4 (N20054, N20046, N5049, N10435, N17272);
or OR3 (N20055, N20053, N8071, N9327);
buf BUF1 (N20056, N20038);
and AND3 (N20057, N20051, N264, N13160);
or OR3 (N20058, N20055, N1350, N7629);
or OR4 (N20059, N20054, N7121, N7559, N18003);
and AND3 (N20060, N20052, N719, N6042);
nand NAND3 (N20061, N20057, N16783, N18004);
not NOT1 (N20062, N20061);
not NOT1 (N20063, N20062);
and AND2 (N20064, N20047, N5323);
nor NOR2 (N20065, N20048, N2314);
and AND4 (N20066, N20016, N16255, N2448, N18975);
nand NAND2 (N20067, N20065, N15557);
nand NAND2 (N20068, N20066, N15344);
buf BUF1 (N20069, N20064);
nand NAND4 (N20070, N20056, N11050, N16332, N14292);
not NOT1 (N20071, N20049);
buf BUF1 (N20072, N20060);
or OR3 (N20073, N20069, N19074, N10441);
or OR4 (N20074, N20070, N8163, N191, N14747);
buf BUF1 (N20075, N20068);
xor XOR2 (N20076, N20050, N13120);
or OR3 (N20077, N20072, N4849, N9170);
nor NOR3 (N20078, N20059, N1371, N15394);
not NOT1 (N20079, N20058);
nand NAND2 (N20080, N20067, N19067);
buf BUF1 (N20081, N20080);
buf BUF1 (N20082, N20074);
xor XOR2 (N20083, N20077, N7726);
or OR2 (N20084, N20071, N2101);
not NOT1 (N20085, N20078);
buf BUF1 (N20086, N20084);
not NOT1 (N20087, N20076);
or OR4 (N20088, N20083, N13049, N11499, N3128);
nor NOR4 (N20089, N20073, N20021, N6840, N9565);
nand NAND3 (N20090, N20085, N19621, N11910);
xor XOR2 (N20091, N20086, N8312);
and AND2 (N20092, N20081, N7177);
and AND3 (N20093, N20079, N14324, N17289);
xor XOR2 (N20094, N20087, N11904);
nand NAND3 (N20095, N20092, N15219, N16033);
nand NAND2 (N20096, N20089, N1385);
or OR4 (N20097, N20095, N19911, N10946, N5571);
nor NOR4 (N20098, N20091, N18595, N11064, N9682);
not NOT1 (N20099, N20098);
nor NOR4 (N20100, N20097, N4079, N15109, N10997);
or OR3 (N20101, N20063, N19421, N19872);
xor XOR2 (N20102, N20101, N3239);
xor XOR2 (N20103, N20090, N6723);
buf BUF1 (N20104, N20082);
buf BUF1 (N20105, N20094);
or OR2 (N20106, N20102, N225);
buf BUF1 (N20107, N20105);
buf BUF1 (N20108, N20075);
or OR3 (N20109, N20104, N3647, N13156);
xor XOR2 (N20110, N20088, N10320);
and AND4 (N20111, N20109, N1720, N9800, N2295);
or OR2 (N20112, N20100, N8320);
nor NOR2 (N20113, N20103, N6887);
xor XOR2 (N20114, N20106, N17187);
nor NOR4 (N20115, N20108, N6627, N12030, N9468);
nor NOR4 (N20116, N20107, N4582, N669, N2631);
nand NAND4 (N20117, N20096, N11712, N13755, N13498);
or OR3 (N20118, N20099, N11049, N9169);
or OR2 (N20119, N20113, N2005);
not NOT1 (N20120, N20116);
nand NAND2 (N20121, N20117, N17464);
buf BUF1 (N20122, N20093);
xor XOR2 (N20123, N20110, N19847);
not NOT1 (N20124, N20122);
buf BUF1 (N20125, N20120);
xor XOR2 (N20126, N20121, N11990);
not NOT1 (N20127, N20119);
or OR4 (N20128, N20127, N14502, N4538, N9778);
buf BUF1 (N20129, N20114);
xor XOR2 (N20130, N20128, N2696);
and AND4 (N20131, N20112, N13525, N9591, N14072);
xor XOR2 (N20132, N20129, N18818);
buf BUF1 (N20133, N20123);
xor XOR2 (N20134, N20131, N10625);
nor NOR2 (N20135, N20124, N5844);
and AND3 (N20136, N20132, N5815, N15430);
nor NOR3 (N20137, N20133, N16532, N19417);
nand NAND2 (N20138, N20115, N9634);
or OR2 (N20139, N20126, N4972);
not NOT1 (N20140, N20134);
nand NAND2 (N20141, N20130, N15934);
not NOT1 (N20142, N20139);
buf BUF1 (N20143, N20111);
and AND2 (N20144, N20136, N12516);
and AND3 (N20145, N20135, N11139, N11408);
nor NOR4 (N20146, N20143, N14213, N14331, N298);
not NOT1 (N20147, N20144);
and AND3 (N20148, N20138, N8124, N8155);
xor XOR2 (N20149, N20137, N3073);
buf BUF1 (N20150, N20118);
and AND4 (N20151, N20149, N15158, N9116, N18499);
buf BUF1 (N20152, N20146);
and AND3 (N20153, N20140, N13988, N16040);
not NOT1 (N20154, N20153);
or OR3 (N20155, N20151, N10909, N15845);
xor XOR2 (N20156, N20142, N12515);
xor XOR2 (N20157, N20150, N7255);
buf BUF1 (N20158, N20145);
xor XOR2 (N20159, N20158, N285);
not NOT1 (N20160, N20147);
xor XOR2 (N20161, N20159, N16056);
and AND2 (N20162, N20154, N8337);
buf BUF1 (N20163, N20161);
or OR3 (N20164, N20125, N15165, N18573);
and AND2 (N20165, N20157, N15353);
buf BUF1 (N20166, N20141);
and AND4 (N20167, N20148, N11480, N9003, N16705);
buf BUF1 (N20168, N20160);
or OR3 (N20169, N20163, N8193, N17355);
buf BUF1 (N20170, N20165);
nand NAND2 (N20171, N20170, N17024);
nor NOR2 (N20172, N20156, N8767);
buf BUF1 (N20173, N20162);
not NOT1 (N20174, N20171);
nand NAND4 (N20175, N20155, N4019, N7982, N17698);
and AND4 (N20176, N20169, N9073, N8611, N5161);
buf BUF1 (N20177, N20164);
buf BUF1 (N20178, N20177);
or OR2 (N20179, N20166, N18976);
nand NAND4 (N20180, N20167, N3045, N7198, N5582);
or OR2 (N20181, N20174, N2973);
or OR3 (N20182, N20172, N10889, N10283);
nand NAND4 (N20183, N20176, N14488, N7198, N19734);
or OR4 (N20184, N20178, N17853, N3119, N4332);
or OR4 (N20185, N20180, N10992, N259, N2816);
buf BUF1 (N20186, N20182);
nor NOR4 (N20187, N20179, N17983, N3786, N2765);
and AND3 (N20188, N20168, N10301, N15836);
nand NAND3 (N20189, N20185, N6730, N15997);
and AND3 (N20190, N20189, N2370, N17078);
or OR4 (N20191, N20173, N206, N11903, N5976);
xor XOR2 (N20192, N20183, N2970);
or OR2 (N20193, N20175, N19882);
nor NOR4 (N20194, N20193, N8379, N132, N1136);
and AND4 (N20195, N20192, N19925, N19172, N7524);
or OR3 (N20196, N20194, N14679, N1349);
buf BUF1 (N20197, N20186);
nor NOR3 (N20198, N20152, N3321, N3036);
not NOT1 (N20199, N20188);
xor XOR2 (N20200, N20196, N14833);
or OR3 (N20201, N20191, N4708, N3960);
and AND4 (N20202, N20184, N19501, N12219, N1004);
and AND4 (N20203, N20199, N353, N4140, N6217);
or OR2 (N20204, N20190, N19576);
buf BUF1 (N20205, N20197);
and AND4 (N20206, N20204, N18702, N4667, N16120);
nor NOR4 (N20207, N20203, N18073, N19228, N14566);
or OR4 (N20208, N20207, N14356, N3562, N5299);
or OR2 (N20209, N20208, N4964);
or OR2 (N20210, N20201, N15434);
nand NAND2 (N20211, N20181, N3841);
nand NAND4 (N20212, N20202, N16897, N11224, N4640);
not NOT1 (N20213, N20195);
nand NAND2 (N20214, N20209, N5345);
or OR2 (N20215, N20213, N12758);
not NOT1 (N20216, N20214);
or OR2 (N20217, N20215, N8783);
or OR3 (N20218, N20198, N7765, N2828);
xor XOR2 (N20219, N20200, N9600);
buf BUF1 (N20220, N20211);
not NOT1 (N20221, N20187);
nand NAND2 (N20222, N20218, N12974);
or OR2 (N20223, N20205, N12073);
xor XOR2 (N20224, N20221, N16517);
nand NAND3 (N20225, N20222, N9867, N5582);
nor NOR2 (N20226, N20224, N7604);
nor NOR3 (N20227, N20223, N16230, N11406);
nand NAND2 (N20228, N20217, N8868);
or OR3 (N20229, N20225, N3539, N18742);
nand NAND3 (N20230, N20226, N9541, N7042);
and AND3 (N20231, N20212, N1666, N16790);
buf BUF1 (N20232, N20206);
and AND2 (N20233, N20231, N13791);
or OR2 (N20234, N20227, N14081);
or OR4 (N20235, N20232, N7313, N8496, N8583);
xor XOR2 (N20236, N20235, N15395);
nor NOR4 (N20237, N20229, N10678, N15842, N11960);
not NOT1 (N20238, N20210);
not NOT1 (N20239, N20220);
xor XOR2 (N20240, N20236, N14407);
nand NAND4 (N20241, N20233, N10541, N17988, N7748);
buf BUF1 (N20242, N20240);
buf BUF1 (N20243, N20230);
nor NOR4 (N20244, N20237, N2530, N19898, N14825);
not NOT1 (N20245, N20228);
buf BUF1 (N20246, N20243);
buf BUF1 (N20247, N20244);
or OR2 (N20248, N20241, N16903);
buf BUF1 (N20249, N20246);
buf BUF1 (N20250, N20249);
or OR2 (N20251, N20248, N5029);
xor XOR2 (N20252, N20216, N18163);
nor NOR2 (N20253, N20247, N7539);
buf BUF1 (N20254, N20242);
xor XOR2 (N20255, N20250, N17648);
and AND4 (N20256, N20245, N6353, N7623, N5740);
nor NOR2 (N20257, N20256, N3333);
nor NOR4 (N20258, N20254, N7786, N5635, N16832);
nor NOR4 (N20259, N20253, N9655, N17495, N747);
not NOT1 (N20260, N20257);
nor NOR3 (N20261, N20255, N11643, N4550);
not NOT1 (N20262, N20252);
xor XOR2 (N20263, N20262, N6995);
and AND4 (N20264, N20239, N11430, N16870, N15310);
buf BUF1 (N20265, N20263);
xor XOR2 (N20266, N20251, N7322);
nor NOR3 (N20267, N20238, N20262, N17558);
or OR3 (N20268, N20267, N771, N18985);
buf BUF1 (N20269, N20266);
not NOT1 (N20270, N20258);
nor NOR4 (N20271, N20234, N6648, N19211, N11576);
xor XOR2 (N20272, N20265, N10350);
and AND2 (N20273, N20260, N2690);
nor NOR4 (N20274, N20219, N12600, N15116, N20051);
nand NAND2 (N20275, N20269, N19825);
not NOT1 (N20276, N20268);
buf BUF1 (N20277, N20275);
nand NAND3 (N20278, N20274, N2075, N17533);
nor NOR4 (N20279, N20270, N20101, N7039, N17637);
not NOT1 (N20280, N20264);
or OR4 (N20281, N20271, N17957, N4815, N2673);
nor NOR3 (N20282, N20273, N12275, N9962);
and AND3 (N20283, N20279, N11518, N5097);
not NOT1 (N20284, N20283);
buf BUF1 (N20285, N20277);
buf BUF1 (N20286, N20284);
buf BUF1 (N20287, N20259);
nor NOR3 (N20288, N20278, N17419, N7519);
and AND3 (N20289, N20276, N16653, N13416);
buf BUF1 (N20290, N20261);
not NOT1 (N20291, N20290);
buf BUF1 (N20292, N20281);
xor XOR2 (N20293, N20291, N10294);
xor XOR2 (N20294, N20286, N18750);
or OR2 (N20295, N20292, N2224);
not NOT1 (N20296, N20272);
not NOT1 (N20297, N20294);
or OR3 (N20298, N20293, N7856, N13317);
xor XOR2 (N20299, N20289, N20038);
or OR4 (N20300, N20280, N17834, N10212, N15093);
nand NAND2 (N20301, N20285, N7353);
and AND2 (N20302, N20288, N10822);
nand NAND2 (N20303, N20296, N10361);
not NOT1 (N20304, N20297);
buf BUF1 (N20305, N20287);
nor NOR4 (N20306, N20303, N16597, N17363, N7880);
buf BUF1 (N20307, N20300);
and AND2 (N20308, N20307, N12371);
nor NOR3 (N20309, N20298, N10223, N12374);
and AND4 (N20310, N20299, N14674, N3018, N10544);
xor XOR2 (N20311, N20282, N15728);
buf BUF1 (N20312, N20295);
buf BUF1 (N20313, N20304);
not NOT1 (N20314, N20305);
xor XOR2 (N20315, N20302, N9059);
nor NOR2 (N20316, N20309, N15257);
nor NOR3 (N20317, N20301, N3139, N2006);
buf BUF1 (N20318, N20317);
xor XOR2 (N20319, N20316, N7248);
nand NAND2 (N20320, N20311, N13307);
and AND4 (N20321, N20318, N11515, N5659, N1777);
not NOT1 (N20322, N20312);
or OR3 (N20323, N20313, N15488, N16016);
and AND4 (N20324, N20322, N7453, N3459, N18072);
not NOT1 (N20325, N20324);
nand NAND4 (N20326, N20323, N3542, N5072, N13364);
and AND3 (N20327, N20306, N15665, N11769);
xor XOR2 (N20328, N20308, N1845);
not NOT1 (N20329, N20328);
not NOT1 (N20330, N20321);
and AND4 (N20331, N20330, N12971, N2510, N333);
or OR2 (N20332, N20310, N14425);
nand NAND3 (N20333, N20329, N1548, N17570);
or OR2 (N20334, N20333, N7446);
nor NOR2 (N20335, N20315, N17553);
not NOT1 (N20336, N20332);
nand NAND3 (N20337, N20334, N359, N15295);
buf BUF1 (N20338, N20320);
or OR4 (N20339, N20319, N19150, N11681, N11767);
nand NAND2 (N20340, N20331, N18267);
not NOT1 (N20341, N20340);
and AND2 (N20342, N20339, N12275);
buf BUF1 (N20343, N20341);
xor XOR2 (N20344, N20314, N9795);
and AND4 (N20345, N20344, N15417, N15661, N5532);
and AND3 (N20346, N20326, N7081, N13685);
buf BUF1 (N20347, N20345);
nand NAND3 (N20348, N20335, N3992, N18477);
nor NOR3 (N20349, N20325, N1452, N4451);
not NOT1 (N20350, N20342);
and AND2 (N20351, N20338, N6333);
or OR3 (N20352, N20347, N1600, N13100);
buf BUF1 (N20353, N20336);
and AND3 (N20354, N20343, N5874, N1440);
buf BUF1 (N20355, N20351);
not NOT1 (N20356, N20353);
buf BUF1 (N20357, N20354);
buf BUF1 (N20358, N20350);
not NOT1 (N20359, N20346);
not NOT1 (N20360, N20356);
xor XOR2 (N20361, N20327, N16980);
xor XOR2 (N20362, N20359, N11496);
xor XOR2 (N20363, N20357, N4623);
xor XOR2 (N20364, N20348, N19251);
and AND3 (N20365, N20362, N3624, N4161);
nand NAND2 (N20366, N20360, N102);
buf BUF1 (N20367, N20337);
nand NAND4 (N20368, N20364, N15872, N2778, N940);
buf BUF1 (N20369, N20352);
buf BUF1 (N20370, N20365);
and AND3 (N20371, N20361, N15145, N6602);
nand NAND2 (N20372, N20363, N705);
xor XOR2 (N20373, N20355, N13240);
buf BUF1 (N20374, N20367);
nor NOR2 (N20375, N20370, N3230);
not NOT1 (N20376, N20349);
and AND3 (N20377, N20375, N9315, N11243);
buf BUF1 (N20378, N20376);
nand NAND2 (N20379, N20373, N1562);
xor XOR2 (N20380, N20366, N1360);
buf BUF1 (N20381, N20369);
nor NOR2 (N20382, N20377, N19631);
not NOT1 (N20383, N20379);
or OR2 (N20384, N20368, N3332);
or OR2 (N20385, N20372, N13650);
and AND4 (N20386, N20380, N9164, N7620, N2983);
buf BUF1 (N20387, N20382);
buf BUF1 (N20388, N20378);
buf BUF1 (N20389, N20381);
buf BUF1 (N20390, N20374);
nand NAND3 (N20391, N20389, N6049, N3251);
or OR2 (N20392, N20358, N4719);
nor NOR3 (N20393, N20387, N20318, N5148);
not NOT1 (N20394, N20383);
not NOT1 (N20395, N20386);
nor NOR3 (N20396, N20385, N9554, N8607);
xor XOR2 (N20397, N20395, N10310);
and AND3 (N20398, N20388, N16001, N9493);
not NOT1 (N20399, N20371);
nor NOR2 (N20400, N20390, N15390);
xor XOR2 (N20401, N20397, N262);
nand NAND4 (N20402, N20394, N11584, N2499, N18085);
or OR2 (N20403, N20384, N3666);
nand NAND2 (N20404, N20398, N8704);
xor XOR2 (N20405, N20402, N12374);
xor XOR2 (N20406, N20403, N2058);
not NOT1 (N20407, N20391);
nand NAND2 (N20408, N20404, N19107);
xor XOR2 (N20409, N20396, N5929);
and AND2 (N20410, N20409, N3416);
xor XOR2 (N20411, N20401, N8105);
nor NOR4 (N20412, N20410, N12762, N8394, N3369);
nand NAND4 (N20413, N20411, N2110, N20038, N15451);
nand NAND2 (N20414, N20406, N8967);
and AND3 (N20415, N20393, N7116, N10734);
buf BUF1 (N20416, N20414);
xor XOR2 (N20417, N20412, N5865);
and AND2 (N20418, N20415, N15150);
nand NAND3 (N20419, N20407, N8080, N16014);
nand NAND3 (N20420, N20417, N19372, N16373);
or OR2 (N20421, N20405, N17212);
not NOT1 (N20422, N20418);
buf BUF1 (N20423, N20416);
not NOT1 (N20424, N20422);
buf BUF1 (N20425, N20408);
or OR4 (N20426, N20400, N827, N3721, N2084);
nand NAND4 (N20427, N20413, N9252, N5614, N1861);
or OR3 (N20428, N20399, N13640, N14517);
not NOT1 (N20429, N20427);
or OR2 (N20430, N20424, N17458);
xor XOR2 (N20431, N20420, N2545);
and AND3 (N20432, N20431, N216, N307);
not NOT1 (N20433, N20426);
xor XOR2 (N20434, N20392, N16940);
or OR2 (N20435, N20430, N2494);
and AND2 (N20436, N20435, N1836);
or OR2 (N20437, N20419, N1512);
not NOT1 (N20438, N20428);
xor XOR2 (N20439, N20421, N6420);
nor NOR4 (N20440, N20425, N7872, N17168, N19215);
nand NAND4 (N20441, N20436, N5251, N6115, N19644);
and AND4 (N20442, N20441, N8369, N4498, N3713);
buf BUF1 (N20443, N20433);
not NOT1 (N20444, N20429);
nor NOR4 (N20445, N20434, N16362, N5008, N14623);
not NOT1 (N20446, N20443);
not NOT1 (N20447, N20446);
not NOT1 (N20448, N20423);
nor NOR4 (N20449, N20448, N4827, N7150, N13433);
and AND3 (N20450, N20442, N15480, N9769);
nand NAND2 (N20451, N20440, N7089);
xor XOR2 (N20452, N20445, N7023);
nor NOR3 (N20453, N20437, N9997, N5231);
not NOT1 (N20454, N20438);
not NOT1 (N20455, N20444);
or OR2 (N20456, N20452, N9704);
nor NOR3 (N20457, N20455, N9885, N6206);
nor NOR3 (N20458, N20432, N14771, N11713);
or OR2 (N20459, N20454, N2656);
not NOT1 (N20460, N20447);
nor NOR2 (N20461, N20456, N8426);
not NOT1 (N20462, N20451);
and AND3 (N20463, N20439, N11798, N2625);
xor XOR2 (N20464, N20461, N14337);
not NOT1 (N20465, N20453);
nand NAND2 (N20466, N20457, N14106);
buf BUF1 (N20467, N20462);
buf BUF1 (N20468, N20465);
not NOT1 (N20469, N20468);
buf BUF1 (N20470, N20450);
buf BUF1 (N20471, N20458);
and AND3 (N20472, N20463, N15108, N19080);
nand NAND4 (N20473, N20459, N11804, N15218, N18146);
or OR2 (N20474, N20472, N17981);
nor NOR4 (N20475, N20474, N16486, N15546, N6187);
and AND3 (N20476, N20475, N19554, N16093);
or OR4 (N20477, N20464, N12990, N10123, N1149);
not NOT1 (N20478, N20470);
and AND4 (N20479, N20477, N5885, N17147, N13048);
or OR2 (N20480, N20469, N19209);
xor XOR2 (N20481, N20473, N19504);
buf BUF1 (N20482, N20480);
nor NOR2 (N20483, N20476, N14943);
xor XOR2 (N20484, N20481, N13773);
nor NOR2 (N20485, N20466, N4998);
or OR4 (N20486, N20449, N4579, N19200, N8106);
buf BUF1 (N20487, N20471);
xor XOR2 (N20488, N20467, N20139);
xor XOR2 (N20489, N20483, N804);
or OR2 (N20490, N20489, N17815);
nand NAND3 (N20491, N20482, N16580, N8256);
xor XOR2 (N20492, N20487, N16142);
or OR2 (N20493, N20478, N9691);
and AND3 (N20494, N20490, N4646, N1256);
buf BUF1 (N20495, N20488);
nor NOR3 (N20496, N20493, N19142, N19425);
xor XOR2 (N20497, N20460, N7174);
buf BUF1 (N20498, N20486);
and AND3 (N20499, N20496, N19464, N5049);
nor NOR3 (N20500, N20495, N8045, N11589);
and AND4 (N20501, N20492, N4807, N20018, N1663);
nand NAND2 (N20502, N20491, N6410);
nand NAND2 (N20503, N20485, N5088);
xor XOR2 (N20504, N20503, N16704);
or OR2 (N20505, N20499, N10212);
buf BUF1 (N20506, N20494);
nand NAND3 (N20507, N20501, N6107, N13635);
nor NOR4 (N20508, N20479, N4178, N14423, N5852);
or OR3 (N20509, N20506, N20233, N13518);
not NOT1 (N20510, N20509);
nand NAND2 (N20511, N20510, N13843);
nand NAND2 (N20512, N20511, N798);
buf BUF1 (N20513, N20508);
and AND3 (N20514, N20497, N1888, N18879);
or OR4 (N20515, N20502, N6037, N5237, N17002);
nor NOR2 (N20516, N20514, N4366);
nand NAND4 (N20517, N20498, N4063, N20202, N5672);
buf BUF1 (N20518, N20512);
nor NOR3 (N20519, N20505, N6297, N3298);
xor XOR2 (N20520, N20507, N3424);
buf BUF1 (N20521, N20519);
xor XOR2 (N20522, N20518, N3439);
not NOT1 (N20523, N20500);
or OR3 (N20524, N20517, N560, N18569);
nor NOR2 (N20525, N20521, N6893);
and AND4 (N20526, N20523, N9773, N1452, N8333);
xor XOR2 (N20527, N20484, N2820);
xor XOR2 (N20528, N20522, N14187);
buf BUF1 (N20529, N20527);
nor NOR4 (N20530, N20528, N9564, N13064, N18418);
not NOT1 (N20531, N20524);
nand NAND4 (N20532, N20504, N10986, N728, N4745);
xor XOR2 (N20533, N20529, N13129);
xor XOR2 (N20534, N20526, N10600);
and AND2 (N20535, N20513, N15519);
xor XOR2 (N20536, N20516, N15180);
nand NAND3 (N20537, N20535, N7239, N8181);
nand NAND3 (N20538, N20533, N9814, N16537);
not NOT1 (N20539, N20515);
or OR3 (N20540, N20530, N13013, N2701);
buf BUF1 (N20541, N20538);
buf BUF1 (N20542, N20532);
not NOT1 (N20543, N20542);
or OR4 (N20544, N20540, N19785, N5859, N5532);
xor XOR2 (N20545, N20531, N11007);
nor NOR2 (N20546, N20536, N383);
buf BUF1 (N20547, N20534);
or OR4 (N20548, N20541, N8082, N19416, N94);
buf BUF1 (N20549, N20520);
or OR4 (N20550, N20546, N1662, N15491, N19017);
nor NOR2 (N20551, N20547, N14119);
nor NOR4 (N20552, N20551, N16949, N10908, N5023);
nand NAND2 (N20553, N20548, N10438);
nor NOR3 (N20554, N20543, N857, N1779);
and AND2 (N20555, N20525, N13473);
nor NOR2 (N20556, N20553, N6133);
nand NAND4 (N20557, N20552, N1767, N10590, N16016);
and AND4 (N20558, N20539, N2150, N5777, N11760);
not NOT1 (N20559, N20545);
not NOT1 (N20560, N20556);
buf BUF1 (N20561, N20557);
nor NOR4 (N20562, N20550, N20084, N10484, N9502);
nor NOR3 (N20563, N20554, N4646, N16227);
nand NAND3 (N20564, N20555, N19905, N1386);
nand NAND2 (N20565, N20563, N10725);
buf BUF1 (N20566, N20560);
and AND2 (N20567, N20562, N9605);
or OR3 (N20568, N20544, N15262, N7015);
buf BUF1 (N20569, N20561);
buf BUF1 (N20570, N20569);
nand NAND3 (N20571, N20565, N8831, N4507);
or OR3 (N20572, N20566, N8847, N12338);
nand NAND3 (N20573, N20549, N19889, N4644);
not NOT1 (N20574, N20564);
nor NOR4 (N20575, N20570, N7535, N3318, N467);
xor XOR2 (N20576, N20559, N9673);
and AND2 (N20577, N20568, N15564);
nand NAND2 (N20578, N20576, N196);
xor XOR2 (N20579, N20558, N18395);
not NOT1 (N20580, N20571);
nor NOR2 (N20581, N20579, N19470);
xor XOR2 (N20582, N20577, N4139);
nor NOR3 (N20583, N20578, N16667, N13218);
buf BUF1 (N20584, N20581);
nor NOR4 (N20585, N20584, N1704, N6512, N8746);
or OR4 (N20586, N20582, N10267, N8982, N5940);
or OR2 (N20587, N20574, N10873);
buf BUF1 (N20588, N20587);
buf BUF1 (N20589, N20588);
buf BUF1 (N20590, N20589);
nor NOR4 (N20591, N20573, N13007, N6015, N17305);
xor XOR2 (N20592, N20537, N6118);
xor XOR2 (N20593, N20585, N17049);
nor NOR3 (N20594, N20591, N12010, N18561);
not NOT1 (N20595, N20592);
xor XOR2 (N20596, N20594, N19614);
nand NAND2 (N20597, N20586, N3479);
and AND4 (N20598, N20596, N10567, N13800, N13786);
buf BUF1 (N20599, N20598);
not NOT1 (N20600, N20567);
nor NOR2 (N20601, N20599, N13584);
buf BUF1 (N20602, N20583);
nor NOR3 (N20603, N20590, N3382, N248);
nand NAND3 (N20604, N20575, N13421, N15993);
not NOT1 (N20605, N20595);
xor XOR2 (N20606, N20604, N6324);
not NOT1 (N20607, N20605);
or OR4 (N20608, N20603, N13478, N2229, N17832);
nand NAND4 (N20609, N20580, N6135, N5312, N17026);
or OR4 (N20610, N20601, N4724, N4281, N2842);
xor XOR2 (N20611, N20609, N3602);
buf BUF1 (N20612, N20572);
xor XOR2 (N20613, N20612, N17673);
nand NAND2 (N20614, N20602, N10511);
buf BUF1 (N20615, N20600);
xor XOR2 (N20616, N20615, N17161);
or OR3 (N20617, N20610, N2027, N17251);
nand NAND4 (N20618, N20614, N19384, N18868, N16694);
buf BUF1 (N20619, N20613);
not NOT1 (N20620, N20597);
not NOT1 (N20621, N20593);
xor XOR2 (N20622, N20607, N12296);
xor XOR2 (N20623, N20616, N2822);
buf BUF1 (N20624, N20622);
nor NOR2 (N20625, N20620, N9518);
or OR2 (N20626, N20608, N18919);
not NOT1 (N20627, N20623);
not NOT1 (N20628, N20624);
not NOT1 (N20629, N20628);
and AND3 (N20630, N20618, N18908, N8244);
and AND3 (N20631, N20619, N18063, N20255);
or OR3 (N20632, N20627, N7845, N2945);
buf BUF1 (N20633, N20625);
or OR3 (N20634, N20633, N16446, N17845);
xor XOR2 (N20635, N20606, N832);
nor NOR2 (N20636, N20631, N12044);
xor XOR2 (N20637, N20626, N17296);
or OR4 (N20638, N20617, N1710, N9714, N10434);
nand NAND4 (N20639, N20638, N3753, N11252, N19448);
and AND4 (N20640, N20630, N16893, N17552, N2922);
nor NOR4 (N20641, N20621, N4264, N2032, N5042);
or OR3 (N20642, N20611, N18148, N1415);
xor XOR2 (N20643, N20637, N13271);
not NOT1 (N20644, N20632);
xor XOR2 (N20645, N20635, N20431);
xor XOR2 (N20646, N20644, N19948);
xor XOR2 (N20647, N20629, N2618);
nand NAND4 (N20648, N20646, N5016, N5075, N91);
not NOT1 (N20649, N20634);
nor NOR2 (N20650, N20648, N384);
nand NAND4 (N20651, N20641, N7411, N6207, N5549);
not NOT1 (N20652, N20645);
and AND3 (N20653, N20643, N7551, N17203);
nor NOR2 (N20654, N20653, N13973);
nor NOR2 (N20655, N20642, N12781);
nor NOR2 (N20656, N20654, N13076);
not NOT1 (N20657, N20636);
and AND2 (N20658, N20656, N14377);
buf BUF1 (N20659, N20649);
nand NAND2 (N20660, N20655, N285);
buf BUF1 (N20661, N20647);
not NOT1 (N20662, N20650);
nand NAND4 (N20663, N20662, N6578, N15841, N4869);
xor XOR2 (N20664, N20652, N19012);
xor XOR2 (N20665, N20657, N14026);
and AND2 (N20666, N20663, N5817);
and AND4 (N20667, N20666, N17487, N7197, N20100);
xor XOR2 (N20668, N20658, N8227);
or OR4 (N20669, N20665, N2313, N14390, N4457);
buf BUF1 (N20670, N20664);
not NOT1 (N20671, N20668);
nor NOR4 (N20672, N20639, N18710, N17781, N11811);
or OR3 (N20673, N20661, N13801, N11700);
xor XOR2 (N20674, N20659, N20214);
nand NAND2 (N20675, N20669, N5829);
xor XOR2 (N20676, N20675, N7777);
nor NOR3 (N20677, N20674, N10445, N12721);
xor XOR2 (N20678, N20676, N10412);
not NOT1 (N20679, N20670);
and AND2 (N20680, N20651, N1251);
and AND2 (N20681, N20677, N9879);
xor XOR2 (N20682, N20678, N8746);
xor XOR2 (N20683, N20660, N19439);
buf BUF1 (N20684, N20681);
xor XOR2 (N20685, N20684, N652);
or OR3 (N20686, N20640, N3461, N14892);
and AND2 (N20687, N20673, N19891);
buf BUF1 (N20688, N20679);
xor XOR2 (N20689, N20667, N13988);
not NOT1 (N20690, N20689);
xor XOR2 (N20691, N20690, N552);
xor XOR2 (N20692, N20691, N7109);
and AND3 (N20693, N20692, N2127, N18750);
buf BUF1 (N20694, N20685);
and AND2 (N20695, N20672, N4106);
and AND3 (N20696, N20687, N19996, N14605);
xor XOR2 (N20697, N20694, N17081);
xor XOR2 (N20698, N20695, N2253);
not NOT1 (N20699, N20682);
nor NOR3 (N20700, N20683, N15726, N1601);
nand NAND3 (N20701, N20688, N9963, N15796);
buf BUF1 (N20702, N20700);
not NOT1 (N20703, N20686);
nor NOR2 (N20704, N20702, N20639);
xor XOR2 (N20705, N20704, N34);
not NOT1 (N20706, N20680);
and AND3 (N20707, N20696, N7776, N8689);
buf BUF1 (N20708, N20697);
nand NAND4 (N20709, N20701, N5746, N1579, N9546);
nand NAND2 (N20710, N20703, N1431);
not NOT1 (N20711, N20709);
nand NAND4 (N20712, N20705, N7170, N2833, N11107);
not NOT1 (N20713, N20710);
nand NAND2 (N20714, N20711, N6060);
nor NOR2 (N20715, N20712, N7303);
buf BUF1 (N20716, N20698);
nand NAND3 (N20717, N20707, N17232, N15928);
or OR4 (N20718, N20713, N3236, N13798, N12008);
xor XOR2 (N20719, N20715, N6066);
and AND3 (N20720, N20671, N3202, N7242);
xor XOR2 (N20721, N20717, N8397);
and AND4 (N20722, N20699, N19124, N8612, N4776);
and AND3 (N20723, N20718, N10997, N2364);
xor XOR2 (N20724, N20716, N17578);
buf BUF1 (N20725, N20720);
nand NAND2 (N20726, N20714, N5197);
and AND2 (N20727, N20693, N6639);
and AND2 (N20728, N20721, N20619);
and AND2 (N20729, N20719, N15165);
nor NOR2 (N20730, N20727, N13737);
xor XOR2 (N20731, N20728, N13601);
xor XOR2 (N20732, N20708, N20380);
and AND4 (N20733, N20726, N1883, N1216, N14922);
or OR3 (N20734, N20732, N5807, N16679);
and AND2 (N20735, N20725, N19815);
buf BUF1 (N20736, N20724);
nor NOR2 (N20737, N20729, N20331);
or OR2 (N20738, N20734, N15389);
nand NAND2 (N20739, N20733, N4955);
not NOT1 (N20740, N20738);
buf BUF1 (N20741, N20722);
and AND4 (N20742, N20735, N19071, N5975, N3104);
nor NOR4 (N20743, N20742, N8689, N18127, N1520);
or OR3 (N20744, N20706, N15737, N8341);
nor NOR4 (N20745, N20737, N4398, N13611, N3395);
or OR2 (N20746, N20741, N2694);
or OR2 (N20747, N20731, N15498);
nand NAND4 (N20748, N20739, N1615, N5335, N10334);
or OR4 (N20749, N20745, N7384, N900, N16178);
or OR2 (N20750, N20740, N8171);
or OR4 (N20751, N20748, N10605, N1810, N17780);
not NOT1 (N20752, N20736);
or OR3 (N20753, N20750, N19381, N16609);
nand NAND2 (N20754, N20751, N3477);
nor NOR3 (N20755, N20723, N3768, N5893);
not NOT1 (N20756, N20754);
nor NOR2 (N20757, N20746, N8686);
or OR3 (N20758, N20747, N9032, N2857);
not NOT1 (N20759, N20756);
buf BUF1 (N20760, N20749);
and AND3 (N20761, N20757, N14947, N9822);
buf BUF1 (N20762, N20760);
and AND3 (N20763, N20730, N8946, N850);
or OR4 (N20764, N20758, N5479, N10500, N6371);
or OR4 (N20765, N20744, N11919, N2619, N15144);
buf BUF1 (N20766, N20753);
xor XOR2 (N20767, N20765, N15070);
or OR4 (N20768, N20762, N9337, N6578, N531);
nand NAND2 (N20769, N20755, N15905);
xor XOR2 (N20770, N20763, N10376);
or OR2 (N20771, N20743, N9851);
nand NAND2 (N20772, N20764, N18041);
xor XOR2 (N20773, N20766, N10094);
xor XOR2 (N20774, N20770, N11590);
buf BUF1 (N20775, N20761);
buf BUF1 (N20776, N20769);
or OR4 (N20777, N20767, N2715, N6033, N1594);
and AND2 (N20778, N20775, N18418);
not NOT1 (N20779, N20771);
not NOT1 (N20780, N20752);
nand NAND4 (N20781, N20772, N18646, N15972, N12256);
nor NOR3 (N20782, N20768, N19091, N12675);
not NOT1 (N20783, N20781);
xor XOR2 (N20784, N20780, N7407);
xor XOR2 (N20785, N20778, N8848);
nand NAND2 (N20786, N20785, N8646);
buf BUF1 (N20787, N20776);
nor NOR2 (N20788, N20779, N17812);
not NOT1 (N20789, N20759);
not NOT1 (N20790, N20789);
nor NOR3 (N20791, N20786, N16434, N20240);
nand NAND4 (N20792, N20783, N19069, N6270, N5760);
nand NAND3 (N20793, N20774, N12920, N17337);
nor NOR3 (N20794, N20784, N7614, N15560);
xor XOR2 (N20795, N20788, N3760);
not NOT1 (N20796, N20782);
nand NAND4 (N20797, N20791, N3534, N16992, N15839);
or OR4 (N20798, N20792, N8387, N5905, N4419);
xor XOR2 (N20799, N20794, N14831);
xor XOR2 (N20800, N20787, N5228);
nand NAND4 (N20801, N20796, N6949, N7319, N3245);
buf BUF1 (N20802, N20795);
and AND2 (N20803, N20799, N20141);
xor XOR2 (N20804, N20802, N11969);
or OR2 (N20805, N20801, N13128);
buf BUF1 (N20806, N20790);
or OR2 (N20807, N20800, N13590);
or OR2 (N20808, N20793, N19754);
and AND3 (N20809, N20808, N2033, N9099);
not NOT1 (N20810, N20798);
and AND4 (N20811, N20797, N20723, N12056, N5914);
or OR4 (N20812, N20809, N18554, N11343, N8723);
nor NOR3 (N20813, N20807, N15062, N11565);
buf BUF1 (N20814, N20812);
or OR3 (N20815, N20810, N11329, N7122);
xor XOR2 (N20816, N20773, N15305);
buf BUF1 (N20817, N20805);
and AND2 (N20818, N20811, N8223);
or OR4 (N20819, N20817, N14096, N13147, N17134);
buf BUF1 (N20820, N20818);
nor NOR3 (N20821, N20806, N17031, N19070);
xor XOR2 (N20822, N20814, N15581);
xor XOR2 (N20823, N20804, N406);
nand NAND2 (N20824, N20822, N5706);
nor NOR2 (N20825, N20815, N6336);
nor NOR2 (N20826, N20821, N4466);
and AND2 (N20827, N20819, N20003);
nand NAND4 (N20828, N20826, N9710, N9582, N8727);
nand NAND4 (N20829, N20803, N1343, N14733, N10554);
nand NAND4 (N20830, N20777, N11534, N7339, N18998);
nand NAND2 (N20831, N20824, N529);
nor NOR2 (N20832, N20830, N19237);
and AND4 (N20833, N20820, N8135, N4910, N19981);
nand NAND4 (N20834, N20813, N7371, N3705, N16986);
nor NOR3 (N20835, N20828, N7381, N7575);
xor XOR2 (N20836, N20825, N15267);
and AND4 (N20837, N20836, N8635, N10188, N6073);
nor NOR4 (N20838, N20832, N5073, N1059, N13332);
nor NOR3 (N20839, N20838, N1944, N17031);
xor XOR2 (N20840, N20827, N20078);
buf BUF1 (N20841, N20837);
or OR2 (N20842, N20833, N11303);
or OR2 (N20843, N20816, N19673);
xor XOR2 (N20844, N20843, N16846);
buf BUF1 (N20845, N20823);
not NOT1 (N20846, N20841);
xor XOR2 (N20847, N20839, N4052);
nand NAND4 (N20848, N20845, N12245, N8003, N13147);
not NOT1 (N20849, N20844);
xor XOR2 (N20850, N20848, N13685);
or OR2 (N20851, N20831, N15414);
and AND2 (N20852, N20840, N8938);
nor NOR3 (N20853, N20852, N19627, N10222);
nor NOR3 (N20854, N20849, N15558, N5410);
and AND2 (N20855, N20853, N987);
nor NOR3 (N20856, N20851, N5044, N12461);
xor XOR2 (N20857, N20842, N23);
nand NAND4 (N20858, N20834, N19558, N14802, N12413);
xor XOR2 (N20859, N20856, N15152);
nand NAND4 (N20860, N20829, N12982, N2343, N1315);
nor NOR3 (N20861, N20854, N16312, N10519);
xor XOR2 (N20862, N20860, N12063);
xor XOR2 (N20863, N20859, N18059);
xor XOR2 (N20864, N20835, N9906);
or OR2 (N20865, N20861, N8745);
and AND4 (N20866, N20862, N5814, N3429, N4765);
or OR3 (N20867, N20863, N7995, N2967);
nor NOR2 (N20868, N20864, N2028);
buf BUF1 (N20869, N20868);
buf BUF1 (N20870, N20846);
and AND3 (N20871, N20858, N17299, N9777);
xor XOR2 (N20872, N20865, N13176);
and AND4 (N20873, N20847, N8377, N455, N15524);
nand NAND3 (N20874, N20857, N16793, N2258);
or OR2 (N20875, N20866, N13795);
or OR3 (N20876, N20855, N10361, N11379);
or OR4 (N20877, N20867, N14389, N3620, N5686);
or OR2 (N20878, N20872, N10866);
not NOT1 (N20879, N20871);
or OR3 (N20880, N20850, N1399, N7869);
and AND2 (N20881, N20875, N16460);
nor NOR4 (N20882, N20878, N1951, N11656, N5513);
nor NOR2 (N20883, N20880, N5186);
nor NOR2 (N20884, N20879, N1488);
xor XOR2 (N20885, N20874, N1249);
xor XOR2 (N20886, N20876, N2956);
nor NOR4 (N20887, N20877, N17251, N3623, N16637);
or OR3 (N20888, N20870, N1308, N19276);
nand NAND3 (N20889, N20869, N5169, N758);
nor NOR3 (N20890, N20881, N8964, N8256);
not NOT1 (N20891, N20886);
buf BUF1 (N20892, N20882);
xor XOR2 (N20893, N20889, N18448);
nor NOR3 (N20894, N20885, N5804, N3047);
buf BUF1 (N20895, N20884);
buf BUF1 (N20896, N20892);
nor NOR4 (N20897, N20887, N16290, N9280, N17555);
and AND4 (N20898, N20891, N12752, N8426, N2576);
nor NOR3 (N20899, N20895, N13296, N14855);
and AND2 (N20900, N20893, N5952);
nand NAND4 (N20901, N20894, N12312, N1572, N12908);
nand NAND4 (N20902, N20890, N6302, N1531, N7831);
nand NAND3 (N20903, N20900, N19616, N19627);
and AND3 (N20904, N20897, N7269, N17446);
buf BUF1 (N20905, N20896);
and AND4 (N20906, N20883, N2136, N15008, N2027);
nor NOR4 (N20907, N20901, N5684, N8681, N8212);
or OR3 (N20908, N20906, N14131, N15237);
or OR3 (N20909, N20908, N18469, N8169);
xor XOR2 (N20910, N20909, N15438);
nand NAND3 (N20911, N20873, N11128, N952);
not NOT1 (N20912, N20904);
buf BUF1 (N20913, N20898);
xor XOR2 (N20914, N20907, N13296);
nor NOR3 (N20915, N20899, N19222, N18088);
not NOT1 (N20916, N20905);
nor NOR2 (N20917, N20915, N5185);
xor XOR2 (N20918, N20912, N4717);
not NOT1 (N20919, N20888);
and AND2 (N20920, N20916, N18723);
and AND3 (N20921, N20918, N9779, N4748);
not NOT1 (N20922, N20910);
not NOT1 (N20923, N20919);
nand NAND3 (N20924, N20914, N6531, N20601);
or OR3 (N20925, N20911, N15258, N10793);
nor NOR4 (N20926, N20913, N1838, N11159, N19920);
nand NAND2 (N20927, N20923, N10571);
or OR2 (N20928, N20902, N11788);
nor NOR2 (N20929, N20920, N17145);
not NOT1 (N20930, N20917);
not NOT1 (N20931, N20921);
nor NOR4 (N20932, N20931, N8700, N10768, N11557);
not NOT1 (N20933, N20922);
and AND3 (N20934, N20903, N2669, N16085);
buf BUF1 (N20935, N20924);
xor XOR2 (N20936, N20930, N14666);
not NOT1 (N20937, N20934);
nand NAND2 (N20938, N20936, N18092);
not NOT1 (N20939, N20928);
or OR4 (N20940, N20939, N5799, N17012, N13507);
xor XOR2 (N20941, N20937, N894);
or OR2 (N20942, N20941, N5144);
nand NAND4 (N20943, N20938, N17836, N1966, N17848);
nand NAND2 (N20944, N20940, N8927);
xor XOR2 (N20945, N20933, N15022);
nor NOR4 (N20946, N20944, N8078, N9271, N17508);
and AND3 (N20947, N20942, N8428, N11421);
nor NOR2 (N20948, N20946, N5792);
and AND2 (N20949, N20926, N6022);
not NOT1 (N20950, N20935);
or OR4 (N20951, N20925, N5469, N1894, N14801);
nor NOR3 (N20952, N20950, N6402, N7453);
and AND2 (N20953, N20951, N7795);
not NOT1 (N20954, N20947);
buf BUF1 (N20955, N20954);
nand NAND3 (N20956, N20927, N11780, N16005);
and AND3 (N20957, N20945, N10572, N15543);
and AND2 (N20958, N20943, N19624);
not NOT1 (N20959, N20958);
nor NOR2 (N20960, N20949, N16028);
and AND4 (N20961, N20955, N11285, N9656, N8657);
or OR2 (N20962, N20932, N15203);
xor XOR2 (N20963, N20962, N4879);
nand NAND3 (N20964, N20953, N9246, N9187);
not NOT1 (N20965, N20948);
buf BUF1 (N20966, N20957);
nand NAND4 (N20967, N20963, N673, N6274, N15352);
nor NOR3 (N20968, N20966, N1002, N15006);
not NOT1 (N20969, N20956);
or OR4 (N20970, N20967, N10226, N19160, N3799);
nor NOR4 (N20971, N20960, N9260, N5451, N11382);
or OR2 (N20972, N20952, N8138);
xor XOR2 (N20973, N20971, N11147);
not NOT1 (N20974, N20964);
nand NAND2 (N20975, N20974, N1492);
and AND3 (N20976, N20961, N3214, N18876);
or OR2 (N20977, N20965, N3491);
nor NOR4 (N20978, N20977, N756, N17065, N18061);
xor XOR2 (N20979, N20969, N9669);
nand NAND3 (N20980, N20975, N13421, N20794);
buf BUF1 (N20981, N20973);
nand NAND2 (N20982, N20929, N3659);
or OR3 (N20983, N20970, N18844, N15889);
nor NOR3 (N20984, N20972, N20823, N9367);
not NOT1 (N20985, N20978);
and AND3 (N20986, N20979, N8752, N19343);
and AND3 (N20987, N20985, N18864, N8152);
nand NAND2 (N20988, N20982, N19897);
or OR3 (N20989, N20981, N20977, N1254);
or OR2 (N20990, N20959, N20418);
or OR4 (N20991, N20983, N10884, N10812, N1465);
nand NAND4 (N20992, N20987, N2767, N82, N1961);
nand NAND2 (N20993, N20984, N13282);
nand NAND4 (N20994, N20991, N4165, N17953, N7597);
not NOT1 (N20995, N20988);
buf BUF1 (N20996, N20980);
nor NOR2 (N20997, N20995, N17957);
nand NAND2 (N20998, N20994, N3791);
xor XOR2 (N20999, N20976, N15796);
or OR2 (N21000, N20992, N3883);
xor XOR2 (N21001, N20997, N1654);
xor XOR2 (N21002, N20998, N19730);
nand NAND4 (N21003, N20996, N3853, N18930, N17632);
nand NAND2 (N21004, N21003, N15597);
and AND2 (N21005, N21004, N15612);
or OR3 (N21006, N20968, N18813, N8854);
and AND4 (N21007, N21006, N12085, N10589, N13925);
xor XOR2 (N21008, N21007, N17216);
nor NOR3 (N21009, N21002, N1712, N17809);
or OR2 (N21010, N20986, N17653);
nand NAND2 (N21011, N20990, N11940);
xor XOR2 (N21012, N21010, N12354);
not NOT1 (N21013, N21008);
not NOT1 (N21014, N20989);
nand NAND4 (N21015, N21000, N16458, N15403, N1926);
not NOT1 (N21016, N21013);
not NOT1 (N21017, N21009);
xor XOR2 (N21018, N21001, N6303);
nand NAND4 (N21019, N20993, N5021, N1035, N1492);
buf BUF1 (N21020, N21017);
and AND2 (N21021, N21016, N13167);
nor NOR3 (N21022, N21018, N11073, N13807);
or OR4 (N21023, N20999, N3508, N19383, N12726);
not NOT1 (N21024, N21020);
xor XOR2 (N21025, N21024, N15526);
nor NOR3 (N21026, N21022, N17574, N17415);
nand NAND3 (N21027, N21021, N4944, N10382);
and AND2 (N21028, N21019, N4829);
not NOT1 (N21029, N21015);
xor XOR2 (N21030, N21028, N11626);
buf BUF1 (N21031, N21023);
or OR4 (N21032, N21027, N20580, N122, N14467);
or OR2 (N21033, N21030, N20092);
and AND2 (N21034, N21005, N5184);
and AND2 (N21035, N21032, N18644);
buf BUF1 (N21036, N21014);
and AND3 (N21037, N21025, N7917, N14391);
or OR2 (N21038, N21011, N2132);
xor XOR2 (N21039, N21031, N20103);
nand NAND4 (N21040, N21036, N5335, N19194, N19178);
or OR2 (N21041, N21038, N229);
buf BUF1 (N21042, N21033);
and AND4 (N21043, N21035, N16935, N1588, N2400);
nor NOR2 (N21044, N21043, N14931);
and AND2 (N21045, N21039, N7003);
not NOT1 (N21046, N21044);
nor NOR4 (N21047, N21041, N12353, N18721, N18947);
xor XOR2 (N21048, N21034, N8497);
and AND4 (N21049, N21037, N10913, N336, N867);
or OR4 (N21050, N21040, N17679, N10675, N4172);
not NOT1 (N21051, N21050);
not NOT1 (N21052, N21049);
nand NAND3 (N21053, N21051, N6947, N17117);
and AND3 (N21054, N21045, N4325, N19437);
and AND2 (N21055, N21047, N2061);
xor XOR2 (N21056, N21054, N2489);
not NOT1 (N21057, N21029);
or OR2 (N21058, N21057, N20630);
nand NAND2 (N21059, N21052, N16040);
buf BUF1 (N21060, N21048);
xor XOR2 (N21061, N21026, N16949);
and AND3 (N21062, N21042, N18932, N4437);
nand NAND4 (N21063, N21012, N7336, N14676, N8715);
nand NAND2 (N21064, N21055, N16220);
and AND3 (N21065, N21064, N14619, N19015);
buf BUF1 (N21066, N21065);
and AND3 (N21067, N21056, N13895, N9181);
nand NAND4 (N21068, N21046, N15276, N11935, N13717);
nor NOR2 (N21069, N21058, N9551);
or OR2 (N21070, N21059, N7094);
not NOT1 (N21071, N21070);
or OR3 (N21072, N21063, N8172, N17761);
xor XOR2 (N21073, N21053, N3996);
xor XOR2 (N21074, N21062, N19274);
buf BUF1 (N21075, N21069);
buf BUF1 (N21076, N21060);
xor XOR2 (N21077, N21075, N4804);
nand NAND3 (N21078, N21074, N7575, N11314);
nand NAND4 (N21079, N21078, N20185, N20365, N16176);
not NOT1 (N21080, N21071);
and AND4 (N21081, N21073, N3779, N5862, N4044);
not NOT1 (N21082, N21066);
and AND4 (N21083, N21079, N4109, N11438, N13981);
xor XOR2 (N21084, N21068, N6759);
nor NOR3 (N21085, N21083, N20074, N1712);
or OR2 (N21086, N21085, N13791);
not NOT1 (N21087, N21072);
nand NAND3 (N21088, N21061, N1426, N4125);
or OR3 (N21089, N21081, N13187, N3328);
nand NAND4 (N21090, N21082, N5468, N13683, N3223);
nand NAND2 (N21091, N21067, N13412);
xor XOR2 (N21092, N21088, N12572);
xor XOR2 (N21093, N21087, N4972);
nand NAND3 (N21094, N21086, N9159, N20766);
or OR2 (N21095, N21090, N6288);
or OR2 (N21096, N21089, N6684);
buf BUF1 (N21097, N21095);
or OR3 (N21098, N21077, N187, N17734);
and AND2 (N21099, N21094, N10814);
nor NOR4 (N21100, N21080, N20944, N490, N6044);
and AND3 (N21101, N21100, N2357, N11799);
and AND2 (N21102, N21084, N13045);
nor NOR3 (N21103, N21096, N3155, N11503);
nand NAND3 (N21104, N21076, N6593, N9779);
buf BUF1 (N21105, N21097);
and AND2 (N21106, N21101, N14526);
or OR2 (N21107, N21104, N6531);
and AND2 (N21108, N21105, N4899);
buf BUF1 (N21109, N21092);
xor XOR2 (N21110, N21098, N14380);
and AND3 (N21111, N21102, N20518, N3356);
or OR3 (N21112, N21109, N8240, N2523);
nor NOR2 (N21113, N21091, N20273);
or OR2 (N21114, N21106, N300);
buf BUF1 (N21115, N21108);
xor XOR2 (N21116, N21113, N9489);
nand NAND2 (N21117, N21115, N13867);
nand NAND3 (N21118, N21110, N3058, N18873);
and AND4 (N21119, N21107, N14995, N18204, N12948);
nor NOR4 (N21120, N21117, N15016, N19843, N6705);
buf BUF1 (N21121, N21103);
or OR3 (N21122, N21093, N669, N8778);
nor NOR3 (N21123, N21112, N10278, N5921);
buf BUF1 (N21124, N21120);
or OR4 (N21125, N21114, N17593, N10348, N13589);
xor XOR2 (N21126, N21116, N2201);
xor XOR2 (N21127, N21119, N18020);
nand NAND2 (N21128, N21111, N3650);
buf BUF1 (N21129, N21128);
not NOT1 (N21130, N21122);
nand NAND2 (N21131, N21099, N19550);
or OR4 (N21132, N21118, N12664, N6942, N11561);
xor XOR2 (N21133, N21127, N7469);
xor XOR2 (N21134, N21131, N15144);
or OR2 (N21135, N21130, N19799);
and AND2 (N21136, N21123, N13325);
not NOT1 (N21137, N21124);
and AND4 (N21138, N21135, N16488, N20757, N13875);
or OR3 (N21139, N21133, N20612, N20980);
or OR3 (N21140, N21121, N3764, N16415);
nor NOR2 (N21141, N21137, N9739);
buf BUF1 (N21142, N21141);
nor NOR3 (N21143, N21129, N8548, N8556);
not NOT1 (N21144, N21142);
or OR2 (N21145, N21126, N18527);
or OR3 (N21146, N21125, N17443, N10458);
and AND2 (N21147, N21144, N3057);
not NOT1 (N21148, N21139);
or OR4 (N21149, N21134, N8490, N5306, N20003);
or OR4 (N21150, N21147, N10897, N9721, N19722);
nor NOR4 (N21151, N21145, N4844, N10291, N2657);
xor XOR2 (N21152, N21151, N1107);
not NOT1 (N21153, N21149);
nor NOR4 (N21154, N21140, N10248, N2680, N16350);
or OR2 (N21155, N21146, N3637);
nand NAND2 (N21156, N21136, N13883);
or OR3 (N21157, N21150, N861, N12320);
nand NAND3 (N21158, N21152, N20347, N16141);
xor XOR2 (N21159, N21153, N7987);
and AND2 (N21160, N21132, N11915);
and AND3 (N21161, N21143, N9408, N14953);
or OR2 (N21162, N21158, N1031);
xor XOR2 (N21163, N21138, N615);
and AND2 (N21164, N21160, N16526);
xor XOR2 (N21165, N21164, N4060);
nor NOR3 (N21166, N21162, N6087, N18729);
nor NOR2 (N21167, N21156, N7184);
nand NAND2 (N21168, N21165, N20644);
nand NAND2 (N21169, N21155, N15445);
or OR2 (N21170, N21166, N2205);
buf BUF1 (N21171, N21161);
buf BUF1 (N21172, N21169);
xor XOR2 (N21173, N21148, N5285);
nor NOR3 (N21174, N21170, N17346, N17796);
nand NAND3 (N21175, N21168, N14824, N11453);
buf BUF1 (N21176, N21173);
and AND4 (N21177, N21167, N6036, N7266, N5691);
nor NOR3 (N21178, N21174, N5240, N1753);
and AND2 (N21179, N21171, N4992);
nand NAND2 (N21180, N21154, N19856);
xor XOR2 (N21181, N21172, N9776);
buf BUF1 (N21182, N21177);
xor XOR2 (N21183, N21178, N7556);
xor XOR2 (N21184, N21163, N10053);
and AND2 (N21185, N21180, N51);
nor NOR4 (N21186, N21183, N18167, N11768, N6252);
and AND4 (N21187, N21185, N13410, N8959, N2261);
buf BUF1 (N21188, N21184);
xor XOR2 (N21189, N21157, N8938);
and AND4 (N21190, N21179, N13292, N1870, N8226);
or OR4 (N21191, N21181, N6680, N11469, N7616);
nand NAND2 (N21192, N21182, N1265);
not NOT1 (N21193, N21192);
xor XOR2 (N21194, N21187, N18781);
not NOT1 (N21195, N21188);
and AND4 (N21196, N21175, N13400, N18594, N12593);
not NOT1 (N21197, N21186);
nand NAND2 (N21198, N21189, N11245);
xor XOR2 (N21199, N21190, N19316);
xor XOR2 (N21200, N21176, N6269);
buf BUF1 (N21201, N21200);
xor XOR2 (N21202, N21199, N6765);
and AND2 (N21203, N21194, N11525);
xor XOR2 (N21204, N21195, N17526);
not NOT1 (N21205, N21196);
buf BUF1 (N21206, N21204);
and AND4 (N21207, N21205, N18662, N7788, N5349);
or OR3 (N21208, N21159, N374, N19634);
nand NAND4 (N21209, N21201, N2963, N4665, N1850);
and AND4 (N21210, N21202, N14868, N9005, N20011);
xor XOR2 (N21211, N21191, N4798);
buf BUF1 (N21212, N21211);
nor NOR3 (N21213, N21203, N15722, N17033);
nand NAND4 (N21214, N21193, N3604, N18605, N17530);
xor XOR2 (N21215, N21206, N10701);
buf BUF1 (N21216, N21208);
and AND4 (N21217, N21197, N1023, N13509, N18493);
xor XOR2 (N21218, N21215, N5366);
and AND4 (N21219, N21214, N20745, N9422, N17191);
or OR3 (N21220, N21212, N20035, N4168);
xor XOR2 (N21221, N21207, N18640);
and AND4 (N21222, N21209, N12912, N14528, N9748);
nand NAND3 (N21223, N21221, N18896, N15204);
and AND3 (N21224, N21217, N18771, N15008);
not NOT1 (N21225, N21198);
nor NOR3 (N21226, N21223, N7433, N1076);
nor NOR4 (N21227, N21213, N20832, N8671, N20604);
nand NAND4 (N21228, N21216, N8505, N5958, N8652);
buf BUF1 (N21229, N21225);
and AND4 (N21230, N21219, N8306, N5620, N11197);
or OR2 (N21231, N21228, N9691);
xor XOR2 (N21232, N21220, N9521);
or OR4 (N21233, N21232, N7500, N7528, N18580);
nor NOR2 (N21234, N21210, N3647);
and AND2 (N21235, N21231, N12840);
nor NOR2 (N21236, N21229, N17829);
xor XOR2 (N21237, N21227, N732);
or OR3 (N21238, N21237, N19741, N16000);
nand NAND4 (N21239, N21222, N14187, N4532, N3859);
xor XOR2 (N21240, N21235, N13140);
xor XOR2 (N21241, N21240, N5280);
nor NOR2 (N21242, N21236, N2823);
nand NAND4 (N21243, N21241, N5569, N6397, N10574);
nor NOR3 (N21244, N21233, N12432, N13154);
buf BUF1 (N21245, N21230);
and AND4 (N21246, N21218, N12466, N18436, N17054);
not NOT1 (N21247, N21226);
not NOT1 (N21248, N21246);
and AND3 (N21249, N21248, N12868, N4914);
buf BUF1 (N21250, N21244);
buf BUF1 (N21251, N21239);
xor XOR2 (N21252, N21224, N9513);
or OR2 (N21253, N21251, N19413);
xor XOR2 (N21254, N21247, N20410);
nor NOR4 (N21255, N21245, N4446, N2183, N19083);
buf BUF1 (N21256, N21250);
or OR2 (N21257, N21253, N1367);
nand NAND4 (N21258, N21252, N19988, N18521, N7892);
nor NOR2 (N21259, N21255, N13156);
nor NOR3 (N21260, N21234, N12288, N1);
or OR2 (N21261, N21257, N5027);
xor XOR2 (N21262, N21259, N11842);
or OR4 (N21263, N21256, N2788, N19697, N20475);
or OR3 (N21264, N21263, N17018, N11199);
nand NAND3 (N21265, N21243, N10590, N15040);
xor XOR2 (N21266, N21254, N17566);
xor XOR2 (N21267, N21260, N13486);
not NOT1 (N21268, N21238);
nor NOR4 (N21269, N21249, N3973, N10649, N14166);
and AND4 (N21270, N21261, N7506, N21113, N5341);
nor NOR3 (N21271, N21270, N21086, N57);
or OR3 (N21272, N21242, N16291, N14340);
and AND4 (N21273, N21266, N12101, N13894, N3306);
or OR3 (N21274, N21272, N16552, N2782);
buf BUF1 (N21275, N21265);
xor XOR2 (N21276, N21273, N1705);
nor NOR3 (N21277, N21264, N13359, N19975);
or OR2 (N21278, N21262, N4693);
nor NOR4 (N21279, N21277, N13643, N6116, N8711);
not NOT1 (N21280, N21267);
nor NOR2 (N21281, N21276, N1613);
buf BUF1 (N21282, N21269);
buf BUF1 (N21283, N21268);
xor XOR2 (N21284, N21275, N8290);
xor XOR2 (N21285, N21258, N7000);
buf BUF1 (N21286, N21282);
buf BUF1 (N21287, N21279);
not NOT1 (N21288, N21281);
buf BUF1 (N21289, N21274);
nand NAND2 (N21290, N21288, N9652);
nor NOR4 (N21291, N21271, N12322, N18048, N6413);
not NOT1 (N21292, N21289);
or OR3 (N21293, N21286, N20917, N20340);
or OR4 (N21294, N21278, N11586, N1197, N5370);
or OR4 (N21295, N21292, N16237, N6914, N1073);
xor XOR2 (N21296, N21285, N10806);
and AND2 (N21297, N21283, N3680);
xor XOR2 (N21298, N21290, N5626);
xor XOR2 (N21299, N21296, N3892);
nor NOR2 (N21300, N21295, N17695);
xor XOR2 (N21301, N21284, N3593);
or OR3 (N21302, N21294, N21117, N16132);
nor NOR3 (N21303, N21301, N16336, N6553);
nand NAND3 (N21304, N21300, N7596, N15731);
buf BUF1 (N21305, N21280);
not NOT1 (N21306, N21298);
buf BUF1 (N21307, N21297);
and AND3 (N21308, N21305, N2936, N8971);
nand NAND3 (N21309, N21308, N17756, N19030);
or OR3 (N21310, N21303, N1608, N9229);
buf BUF1 (N21311, N21310);
xor XOR2 (N21312, N21306, N16622);
nor NOR2 (N21313, N21287, N7715);
nand NAND2 (N21314, N21302, N3491);
nand NAND3 (N21315, N21307, N6783, N5809);
xor XOR2 (N21316, N21314, N10551);
nor NOR2 (N21317, N21311, N989);
buf BUF1 (N21318, N21313);
buf BUF1 (N21319, N21318);
and AND2 (N21320, N21293, N13422);
or OR3 (N21321, N21319, N18221, N7766);
not NOT1 (N21322, N21317);
not NOT1 (N21323, N21291);
buf BUF1 (N21324, N21316);
nor NOR4 (N21325, N21315, N16514, N5782, N13018);
or OR2 (N21326, N21304, N15771);
or OR2 (N21327, N21322, N2586);
buf BUF1 (N21328, N21326);
nand NAND3 (N21329, N21324, N4482, N2092);
nand NAND4 (N21330, N21321, N11538, N1364, N7349);
xor XOR2 (N21331, N21299, N18303);
xor XOR2 (N21332, N21331, N18607);
not NOT1 (N21333, N21329);
nor NOR3 (N21334, N21327, N2127, N19828);
and AND2 (N21335, N21330, N19913);
nand NAND2 (N21336, N21334, N16433);
or OR3 (N21337, N21333, N584, N14401);
buf BUF1 (N21338, N21320);
xor XOR2 (N21339, N21325, N8926);
and AND2 (N21340, N21323, N698);
and AND3 (N21341, N21338, N9812, N20388);
nand NAND4 (N21342, N21332, N14897, N5249, N5289);
buf BUF1 (N21343, N21337);
nand NAND3 (N21344, N21339, N13429, N4233);
or OR3 (N21345, N21344, N1982, N1979);
or OR2 (N21346, N21343, N18788);
buf BUF1 (N21347, N21312);
xor XOR2 (N21348, N21345, N14784);
nand NAND3 (N21349, N21348, N13756, N3727);
or OR3 (N21350, N21342, N16849, N121);
not NOT1 (N21351, N21340);
xor XOR2 (N21352, N21351, N8706);
or OR3 (N21353, N21346, N21248, N11780);
nand NAND3 (N21354, N21336, N11211, N153);
and AND3 (N21355, N21352, N17333, N17771);
not NOT1 (N21356, N21353);
nor NOR4 (N21357, N21347, N11135, N14422, N17642);
not NOT1 (N21358, N21356);
nor NOR2 (N21359, N21335, N10963);
not NOT1 (N21360, N21309);
xor XOR2 (N21361, N21358, N17056);
nor NOR2 (N21362, N21354, N4667);
or OR4 (N21363, N21341, N10542, N20576, N13438);
nand NAND4 (N21364, N21363, N16590, N16243, N13674);
or OR2 (N21365, N21328, N19313);
not NOT1 (N21366, N21364);
or OR2 (N21367, N21366, N5285);
or OR3 (N21368, N21359, N4360, N13221);
and AND3 (N21369, N21368, N14068, N7580);
nand NAND4 (N21370, N21369, N15725, N6650, N20632);
and AND4 (N21371, N21362, N15230, N14755, N6111);
xor XOR2 (N21372, N21370, N7225);
buf BUF1 (N21373, N21360);
nor NOR3 (N21374, N21350, N8036, N16185);
buf BUF1 (N21375, N21357);
xor XOR2 (N21376, N21367, N4500);
buf BUF1 (N21377, N21375);
or OR2 (N21378, N21377, N8415);
and AND4 (N21379, N21373, N2046, N19781, N11169);
nor NOR3 (N21380, N21372, N21082, N21134);
and AND3 (N21381, N21349, N14935, N10995);
and AND4 (N21382, N21378, N5899, N14094, N13456);
and AND2 (N21383, N21374, N16263);
xor XOR2 (N21384, N21365, N17909);
and AND2 (N21385, N21361, N17885);
buf BUF1 (N21386, N21379);
nand NAND3 (N21387, N21384, N6274, N329);
not NOT1 (N21388, N21371);
and AND3 (N21389, N21376, N10050, N6471);
and AND4 (N21390, N21386, N1217, N1424, N18034);
not NOT1 (N21391, N21388);
nand NAND2 (N21392, N21383, N19296);
not NOT1 (N21393, N21391);
nand NAND3 (N21394, N21392, N1329, N1519);
or OR4 (N21395, N21394, N17329, N1409, N18042);
not NOT1 (N21396, N21355);
nand NAND3 (N21397, N21380, N10585, N5572);
and AND3 (N21398, N21397, N14226, N4313);
buf BUF1 (N21399, N21385);
xor XOR2 (N21400, N21395, N16962);
and AND3 (N21401, N21381, N17015, N13177);
and AND3 (N21402, N21396, N12770, N18400);
nand NAND3 (N21403, N21389, N18330, N7180);
nand NAND3 (N21404, N21399, N1395, N2160);
nand NAND3 (N21405, N21401, N7836, N4104);
and AND4 (N21406, N21390, N1671, N19951, N13502);
buf BUF1 (N21407, N21393);
not NOT1 (N21408, N21382);
buf BUF1 (N21409, N21402);
and AND3 (N21410, N21408, N8004, N18969);
nor NOR2 (N21411, N21406, N7308);
buf BUF1 (N21412, N21400);
not NOT1 (N21413, N21398);
nor NOR3 (N21414, N21413, N9939, N12735);
xor XOR2 (N21415, N21404, N17407);
and AND3 (N21416, N21407, N5696, N19366);
or OR4 (N21417, N21416, N4704, N6899, N2473);
xor XOR2 (N21418, N21403, N7216);
xor XOR2 (N21419, N21410, N14642);
nand NAND3 (N21420, N21411, N17332, N5662);
not NOT1 (N21421, N21387);
and AND2 (N21422, N21420, N14491);
not NOT1 (N21423, N21405);
not NOT1 (N21424, N21409);
not NOT1 (N21425, N21418);
or OR4 (N21426, N21415, N3810, N19894, N20710);
nand NAND2 (N21427, N21422, N19912);
xor XOR2 (N21428, N21427, N6492);
or OR3 (N21429, N21421, N19408, N8923);
or OR4 (N21430, N21428, N17027, N12516, N7895);
xor XOR2 (N21431, N21417, N8038);
not NOT1 (N21432, N21425);
or OR3 (N21433, N21431, N6859, N9437);
not NOT1 (N21434, N21432);
xor XOR2 (N21435, N21426, N19958);
or OR4 (N21436, N21435, N17189, N5832, N9944);
and AND3 (N21437, N21414, N12923, N7410);
and AND4 (N21438, N21434, N13063, N16700, N16883);
not NOT1 (N21439, N21436);
nand NAND3 (N21440, N21419, N10995, N20915);
nor NOR2 (N21441, N21424, N12420);
and AND3 (N21442, N21429, N13985, N5981);
or OR3 (N21443, N21440, N18410, N3443);
buf BUF1 (N21444, N21438);
nor NOR4 (N21445, N21439, N19295, N14606, N4344);
xor XOR2 (N21446, N21433, N8071);
nand NAND4 (N21447, N21446, N3270, N10769, N19870);
and AND3 (N21448, N21437, N5850, N8327);
xor XOR2 (N21449, N21443, N1329);
and AND4 (N21450, N21441, N316, N15518, N12960);
xor XOR2 (N21451, N21430, N5475);
not NOT1 (N21452, N21449);
xor XOR2 (N21453, N21444, N16496);
buf BUF1 (N21454, N21423);
nor NOR3 (N21455, N21453, N20098, N19677);
not NOT1 (N21456, N21447);
and AND2 (N21457, N21445, N15634);
nor NOR4 (N21458, N21448, N707, N1545, N14541);
or OR3 (N21459, N21456, N15839, N6493);
not NOT1 (N21460, N21452);
xor XOR2 (N21461, N21460, N17901);
not NOT1 (N21462, N21459);
not NOT1 (N21463, N21458);
buf BUF1 (N21464, N21461);
not NOT1 (N21465, N21463);
buf BUF1 (N21466, N21412);
not NOT1 (N21467, N21454);
nor NOR4 (N21468, N21455, N633, N4874, N341);
nor NOR4 (N21469, N21465, N6738, N3947, N9634);
buf BUF1 (N21470, N21450);
or OR4 (N21471, N21442, N325, N21136, N446);
nand NAND2 (N21472, N21457, N6030);
nand NAND3 (N21473, N21471, N14226, N8699);
buf BUF1 (N21474, N21470);
buf BUF1 (N21475, N21473);
buf BUF1 (N21476, N21451);
nand NAND2 (N21477, N21472, N21009);
not NOT1 (N21478, N21466);
nand NAND2 (N21479, N21467, N5400);
not NOT1 (N21480, N21469);
nor NOR3 (N21481, N21478, N502, N3389);
or OR4 (N21482, N21464, N19643, N15069, N16798);
buf BUF1 (N21483, N21479);
not NOT1 (N21484, N21480);
nand NAND3 (N21485, N21482, N8166, N12245);
nor NOR3 (N21486, N21468, N10734, N1428);
or OR4 (N21487, N21484, N7932, N10004, N12791);
nor NOR4 (N21488, N21477, N15196, N7381, N19970);
xor XOR2 (N21489, N21476, N19341);
and AND2 (N21490, N21481, N2711);
nand NAND2 (N21491, N21486, N13069);
nand NAND2 (N21492, N21490, N1437);
and AND4 (N21493, N21491, N2128, N6271, N10614);
xor XOR2 (N21494, N21485, N18248);
buf BUF1 (N21495, N21474);
or OR2 (N21496, N21462, N17900);
nand NAND4 (N21497, N21495, N946, N14468, N7482);
nor NOR4 (N21498, N21488, N15510, N18873, N16409);
xor XOR2 (N21499, N21493, N5796);
and AND4 (N21500, N21497, N16179, N9207, N4081);
or OR2 (N21501, N21499, N13143);
and AND4 (N21502, N21498, N20685, N14691, N6997);
buf BUF1 (N21503, N21501);
nand NAND2 (N21504, N21502, N6817);
or OR3 (N21505, N21500, N1559, N7112);
buf BUF1 (N21506, N21504);
or OR4 (N21507, N21487, N5306, N5599, N18448);
or OR3 (N21508, N21505, N16826, N13500);
not NOT1 (N21509, N21496);
nand NAND3 (N21510, N21492, N1091, N16964);
xor XOR2 (N21511, N21507, N1660);
nor NOR3 (N21512, N21483, N5605, N12649);
nor NOR4 (N21513, N21506, N526, N2232, N20411);
and AND4 (N21514, N21508, N6033, N17180, N6914);
nand NAND2 (N21515, N21513, N3838);
buf BUF1 (N21516, N21515);
and AND4 (N21517, N21512, N15253, N6390, N17743);
nor NOR4 (N21518, N21511, N8668, N12675, N5163);
xor XOR2 (N21519, N21503, N16783);
not NOT1 (N21520, N21519);
and AND3 (N21521, N21489, N4830, N15211);
xor XOR2 (N21522, N21517, N6358);
buf BUF1 (N21523, N21521);
xor XOR2 (N21524, N21509, N20748);
not NOT1 (N21525, N21475);
xor XOR2 (N21526, N21520, N2583);
xor XOR2 (N21527, N21522, N325);
not NOT1 (N21528, N21525);
nor NOR4 (N21529, N21514, N3208, N5998, N8934);
and AND4 (N21530, N21529, N9710, N4983, N990);
or OR3 (N21531, N21530, N3430, N5174);
nor NOR3 (N21532, N21516, N12511, N10358);
or OR2 (N21533, N21524, N19015);
and AND2 (N21534, N21533, N12533);
nor NOR2 (N21535, N21510, N21168);
buf BUF1 (N21536, N21532);
and AND3 (N21537, N21536, N562, N1426);
buf BUF1 (N21538, N21494);
or OR2 (N21539, N21534, N8271);
or OR3 (N21540, N21539, N8427, N1460);
or OR2 (N21541, N21528, N3864);
and AND4 (N21542, N21518, N15703, N1719, N4978);
nand NAND2 (N21543, N21537, N7717);
not NOT1 (N21544, N21526);
nand NAND2 (N21545, N21542, N18717);
and AND3 (N21546, N21527, N4026, N8871);
nand NAND3 (N21547, N21538, N6669, N1968);
buf BUF1 (N21548, N21547);
buf BUF1 (N21549, N21546);
and AND4 (N21550, N21541, N10496, N19224, N5772);
not NOT1 (N21551, N21540);
or OR3 (N21552, N21535, N17574, N20693);
nor NOR3 (N21553, N21545, N9565, N2014);
xor XOR2 (N21554, N21551, N11939);
and AND2 (N21555, N21543, N19342);
not NOT1 (N21556, N21554);
not NOT1 (N21557, N21552);
not NOT1 (N21558, N21556);
nor NOR4 (N21559, N21544, N15510, N1511, N10707);
buf BUF1 (N21560, N21550);
or OR2 (N21561, N21559, N2044);
or OR2 (N21562, N21560, N14191);
and AND3 (N21563, N21553, N14664, N10184);
or OR3 (N21564, N21561, N12985, N2383);
not NOT1 (N21565, N21564);
nand NAND4 (N21566, N21531, N2774, N566, N7718);
nand NAND4 (N21567, N21563, N11861, N14111, N19056);
nand NAND3 (N21568, N21565, N3187, N443);
nand NAND2 (N21569, N21567, N2294);
nand NAND3 (N21570, N21569, N8229, N3130);
and AND4 (N21571, N21557, N2950, N10307, N19849);
nand NAND2 (N21572, N21568, N13254);
xor XOR2 (N21573, N21555, N1675);
not NOT1 (N21574, N21571);
or OR3 (N21575, N21566, N5291, N14417);
or OR3 (N21576, N21570, N21404, N18699);
or OR3 (N21577, N21548, N9152, N4786);
buf BUF1 (N21578, N21549);
and AND4 (N21579, N21573, N9482, N11145, N38);
buf BUF1 (N21580, N21572);
buf BUF1 (N21581, N21575);
buf BUF1 (N21582, N21579);
xor XOR2 (N21583, N21574, N718);
nand NAND3 (N21584, N21581, N20346, N15924);
xor XOR2 (N21585, N21562, N8757);
nor NOR3 (N21586, N21576, N16796, N5064);
buf BUF1 (N21587, N21523);
not NOT1 (N21588, N21580);
xor XOR2 (N21589, N21578, N13268);
and AND3 (N21590, N21587, N2227, N1964);
and AND3 (N21591, N21577, N7646, N3946);
nor NOR4 (N21592, N21558, N13201, N1345, N16570);
nor NOR2 (N21593, N21585, N16776);
and AND2 (N21594, N21586, N1866);
nor NOR3 (N21595, N21594, N5789, N12957);
nor NOR3 (N21596, N21590, N520, N19245);
nor NOR4 (N21597, N21593, N15544, N11865, N800);
not NOT1 (N21598, N21583);
or OR3 (N21599, N21584, N18958, N17829);
nand NAND2 (N21600, N21599, N5300);
nor NOR4 (N21601, N21595, N5292, N6269, N229);
buf BUF1 (N21602, N21588);
buf BUF1 (N21603, N21597);
nand NAND2 (N21604, N21603, N11176);
not NOT1 (N21605, N21582);
and AND2 (N21606, N21605, N85);
not NOT1 (N21607, N21606);
nor NOR3 (N21608, N21592, N2974, N513);
buf BUF1 (N21609, N21596);
nand NAND2 (N21610, N21600, N9301);
not NOT1 (N21611, N21589);
and AND3 (N21612, N21598, N4088, N18751);
buf BUF1 (N21613, N21591);
nand NAND2 (N21614, N21612, N16955);
and AND4 (N21615, N21609, N16463, N7875, N13352);
nor NOR3 (N21616, N21604, N10758, N13972);
nor NOR2 (N21617, N21601, N7845);
or OR3 (N21618, N21611, N4666, N5188);
not NOT1 (N21619, N21614);
not NOT1 (N21620, N21617);
not NOT1 (N21621, N21616);
or OR2 (N21622, N21618, N5033);
buf BUF1 (N21623, N21622);
or OR3 (N21624, N21621, N10032, N8293);
or OR2 (N21625, N21602, N1478);
and AND4 (N21626, N21625, N6947, N19083, N18167);
or OR2 (N21627, N21623, N3285);
not NOT1 (N21628, N21627);
nand NAND2 (N21629, N21608, N3658);
or OR4 (N21630, N21619, N16283, N18487, N4412);
nor NOR4 (N21631, N21628, N11377, N15423, N4045);
buf BUF1 (N21632, N21626);
nand NAND3 (N21633, N21629, N11085, N19523);
and AND2 (N21634, N21607, N7490);
not NOT1 (N21635, N21630);
not NOT1 (N21636, N21635);
not NOT1 (N21637, N21624);
or OR3 (N21638, N21633, N18279, N8911);
nor NOR2 (N21639, N21636, N10315);
xor XOR2 (N21640, N21615, N11346);
nor NOR2 (N21641, N21632, N15673);
nor NOR2 (N21642, N21637, N1610);
xor XOR2 (N21643, N21642, N16372);
or OR2 (N21644, N21634, N8786);
xor XOR2 (N21645, N21620, N11932);
nand NAND4 (N21646, N21638, N16089, N18034, N6727);
buf BUF1 (N21647, N21631);
xor XOR2 (N21648, N21644, N18030);
nor NOR4 (N21649, N21646, N14171, N3443, N8033);
and AND4 (N21650, N21643, N2367, N7915, N20393);
nand NAND3 (N21651, N21610, N16529, N1441);
xor XOR2 (N21652, N21651, N13704);
buf BUF1 (N21653, N21652);
and AND4 (N21654, N21645, N3860, N3536, N10);
and AND3 (N21655, N21648, N1496, N16851);
buf BUF1 (N21656, N21649);
nor NOR3 (N21657, N21650, N19383, N4580);
not NOT1 (N21658, N21655);
not NOT1 (N21659, N21654);
and AND2 (N21660, N21656, N14817);
nand NAND2 (N21661, N21639, N10568);
buf BUF1 (N21662, N21657);
buf BUF1 (N21663, N21641);
or OR3 (N21664, N21661, N2603, N2475);
and AND2 (N21665, N21613, N20091);
xor XOR2 (N21666, N21653, N18730);
and AND2 (N21667, N21659, N4611);
nor NOR4 (N21668, N21666, N6594, N14229, N12506);
xor XOR2 (N21669, N21658, N9120);
nor NOR3 (N21670, N21668, N12501, N20111);
xor XOR2 (N21671, N21647, N21539);
or OR4 (N21672, N21663, N10696, N6836, N13445);
buf BUF1 (N21673, N21669);
nand NAND3 (N21674, N21671, N20897, N1762);
buf BUF1 (N21675, N21670);
buf BUF1 (N21676, N21673);
and AND3 (N21677, N21672, N5428, N7155);
or OR2 (N21678, N21667, N16491);
not NOT1 (N21679, N21674);
not NOT1 (N21680, N21664);
and AND3 (N21681, N21665, N18699, N4253);
buf BUF1 (N21682, N21640);
buf BUF1 (N21683, N21679);
and AND2 (N21684, N21677, N15537);
nor NOR4 (N21685, N21676, N11402, N388, N4502);
nor NOR4 (N21686, N21682, N9368, N11689, N16843);
or OR3 (N21687, N21681, N10778, N10577);
xor XOR2 (N21688, N21684, N8916);
and AND4 (N21689, N21662, N17676, N8755, N7596);
or OR2 (N21690, N21687, N6795);
buf BUF1 (N21691, N21685);
not NOT1 (N21692, N21680);
and AND4 (N21693, N21689, N9285, N14484, N14323);
and AND2 (N21694, N21678, N968);
and AND4 (N21695, N21690, N6985, N14085, N567);
not NOT1 (N21696, N21688);
not NOT1 (N21697, N21694);
buf BUF1 (N21698, N21683);
xor XOR2 (N21699, N21691, N11251);
or OR2 (N21700, N21660, N285);
and AND2 (N21701, N21696, N13271);
nor NOR3 (N21702, N21697, N15928, N16436);
not NOT1 (N21703, N21700);
nor NOR4 (N21704, N21698, N19012, N8475, N8453);
and AND4 (N21705, N21701, N9890, N2166, N11329);
xor XOR2 (N21706, N21695, N15483);
or OR4 (N21707, N21703, N1658, N13696, N5066);
nand NAND4 (N21708, N21692, N9104, N3412, N20577);
nor NOR4 (N21709, N21702, N4977, N9061, N19146);
nor NOR4 (N21710, N21675, N1854, N12797, N6695);
buf BUF1 (N21711, N21708);
not NOT1 (N21712, N21706);
and AND4 (N21713, N21709, N13454, N14892, N14596);
xor XOR2 (N21714, N21705, N21448);
or OR2 (N21715, N21710, N20400);
xor XOR2 (N21716, N21693, N20457);
buf BUF1 (N21717, N21699);
or OR4 (N21718, N21712, N11805, N10833, N5545);
buf BUF1 (N21719, N21686);
xor XOR2 (N21720, N21711, N1657);
nor NOR3 (N21721, N21717, N4014, N19894);
nor NOR2 (N21722, N21719, N10845);
not NOT1 (N21723, N21715);
or OR2 (N21724, N21723, N2086);
nand NAND2 (N21725, N21716, N19076);
nand NAND4 (N21726, N21720, N12085, N15717, N12183);
and AND4 (N21727, N21718, N4578, N820, N4104);
nor NOR3 (N21728, N21722, N6707, N17260);
or OR2 (N21729, N21721, N16291);
buf BUF1 (N21730, N21725);
not NOT1 (N21731, N21727);
or OR2 (N21732, N21729, N11877);
or OR3 (N21733, N21707, N13737, N5192);
or OR2 (N21734, N21733, N16627);
nand NAND4 (N21735, N21731, N14111, N7358, N12096);
or OR4 (N21736, N21728, N9625, N19236, N9560);
or OR4 (N21737, N21732, N19151, N21611, N14687);
xor XOR2 (N21738, N21735, N10981);
nand NAND4 (N21739, N21738, N1421, N8675, N6413);
nand NAND3 (N21740, N21730, N1616, N4514);
nand NAND3 (N21741, N21740, N2851, N427);
xor XOR2 (N21742, N21726, N3904);
nor NOR3 (N21743, N21741, N16733, N6432);
nand NAND3 (N21744, N21737, N17628, N2293);
nor NOR3 (N21745, N21734, N5788, N7976);
nor NOR3 (N21746, N21742, N20075, N13074);
and AND2 (N21747, N21739, N4250);
nor NOR3 (N21748, N21714, N13842, N13970);
buf BUF1 (N21749, N21747);
buf BUF1 (N21750, N21724);
nand NAND2 (N21751, N21736, N16581);
not NOT1 (N21752, N21743);
nand NAND4 (N21753, N21748, N17207, N20340, N5897);
not NOT1 (N21754, N21750);
buf BUF1 (N21755, N21752);
not NOT1 (N21756, N21749);
or OR4 (N21757, N21751, N16418, N12360, N6276);
nand NAND2 (N21758, N21704, N10966);
buf BUF1 (N21759, N21745);
xor XOR2 (N21760, N21754, N14012);
nand NAND2 (N21761, N21744, N10678);
nor NOR2 (N21762, N21753, N15334);
or OR4 (N21763, N21755, N259, N14284, N20159);
or OR4 (N21764, N21760, N932, N14213, N2233);
or OR4 (N21765, N21758, N8431, N14075, N14813);
xor XOR2 (N21766, N21764, N11431);
nand NAND4 (N21767, N21759, N10404, N9446, N2085);
xor XOR2 (N21768, N21767, N1110);
or OR3 (N21769, N21746, N9003, N14599);
buf BUF1 (N21770, N21763);
nor NOR4 (N21771, N21762, N12515, N9397, N6405);
or OR3 (N21772, N21771, N832, N17685);
nor NOR4 (N21773, N21770, N5051, N6316, N8133);
xor XOR2 (N21774, N21713, N20632);
nor NOR4 (N21775, N21769, N12634, N6734, N1498);
not NOT1 (N21776, N21772);
xor XOR2 (N21777, N21775, N15583);
nand NAND4 (N21778, N21756, N16001, N2081, N12687);
nand NAND2 (N21779, N21774, N982);
or OR2 (N21780, N21757, N7223);
xor XOR2 (N21781, N21779, N4902);
not NOT1 (N21782, N21777);
nor NOR2 (N21783, N21766, N5750);
buf BUF1 (N21784, N21780);
and AND3 (N21785, N21768, N21123, N11574);
nand NAND3 (N21786, N21761, N11237, N3322);
xor XOR2 (N21787, N21782, N17277);
buf BUF1 (N21788, N21778);
and AND4 (N21789, N21781, N10705, N21117, N5622);
nor NOR3 (N21790, N21788, N15134, N14105);
buf BUF1 (N21791, N21773);
nand NAND2 (N21792, N21785, N14691);
xor XOR2 (N21793, N21787, N17749);
nor NOR3 (N21794, N21786, N11315, N8994);
or OR4 (N21795, N21793, N12727, N21604, N9548);
xor XOR2 (N21796, N21792, N4855);
buf BUF1 (N21797, N21784);
not NOT1 (N21798, N21794);
xor XOR2 (N21799, N21789, N6649);
and AND3 (N21800, N21765, N12272, N4827);
and AND3 (N21801, N21799, N17868, N13486);
not NOT1 (N21802, N21800);
or OR3 (N21803, N21801, N449, N19607);
and AND3 (N21804, N21802, N16084, N19309);
nor NOR4 (N21805, N21798, N7977, N5543, N13727);
and AND3 (N21806, N21791, N13279, N10303);
buf BUF1 (N21807, N21805);
nand NAND2 (N21808, N21776, N17774);
nor NOR4 (N21809, N21806, N15998, N11098, N2783);
xor XOR2 (N21810, N21796, N5144);
nor NOR4 (N21811, N21783, N3915, N16370, N9788);
buf BUF1 (N21812, N21810);
nand NAND2 (N21813, N21804, N18155);
buf BUF1 (N21814, N21812);
or OR3 (N21815, N21803, N6230, N17988);
or OR2 (N21816, N21808, N3588);
and AND2 (N21817, N21790, N4620);
not NOT1 (N21818, N21814);
not NOT1 (N21819, N21813);
and AND3 (N21820, N21811, N1548, N18071);
and AND3 (N21821, N21807, N17, N630);
xor XOR2 (N21822, N21818, N841);
nor NOR4 (N21823, N21809, N20900, N4065, N9427);
buf BUF1 (N21824, N21821);
buf BUF1 (N21825, N21815);
buf BUF1 (N21826, N21797);
or OR2 (N21827, N21817, N21723);
or OR3 (N21828, N21795, N12813, N10307);
nor NOR2 (N21829, N21826, N18749);
not NOT1 (N21830, N21820);
buf BUF1 (N21831, N21830);
nor NOR3 (N21832, N21816, N18282, N13622);
buf BUF1 (N21833, N21829);
xor XOR2 (N21834, N21819, N2489);
and AND2 (N21835, N21834, N12771);
and AND3 (N21836, N21828, N12836, N6843);
nand NAND2 (N21837, N21832, N18750);
not NOT1 (N21838, N21831);
nand NAND4 (N21839, N21827, N14504, N3884, N8546);
or OR2 (N21840, N21833, N5660);
nand NAND3 (N21841, N21838, N12507, N9711);
nand NAND2 (N21842, N21824, N21517);
xor XOR2 (N21843, N21839, N226);
nand NAND4 (N21844, N21843, N16088, N11682, N6938);
not NOT1 (N21845, N21837);
or OR4 (N21846, N21841, N2174, N5329, N17807);
xor XOR2 (N21847, N21845, N5628);
xor XOR2 (N21848, N21842, N10385);
buf BUF1 (N21849, N21844);
nand NAND4 (N21850, N21847, N21426, N3638, N6323);
xor XOR2 (N21851, N21850, N1598);
xor XOR2 (N21852, N21846, N10445);
and AND3 (N21853, N21852, N18600, N8700);
not NOT1 (N21854, N21840);
or OR2 (N21855, N21823, N6443);
and AND4 (N21856, N21835, N15833, N18091, N7693);
buf BUF1 (N21857, N21853);
nor NOR2 (N21858, N21857, N5793);
buf BUF1 (N21859, N21836);
buf BUF1 (N21860, N21822);
nor NOR4 (N21861, N21851, N5476, N9244, N8316);
and AND4 (N21862, N21861, N3063, N20974, N16398);
xor XOR2 (N21863, N21858, N1002);
and AND3 (N21864, N21848, N1084, N14460);
or OR3 (N21865, N21860, N17725, N1243);
xor XOR2 (N21866, N21855, N16652);
not NOT1 (N21867, N21825);
nor NOR2 (N21868, N21867, N9608);
nand NAND3 (N21869, N21862, N13622, N12746);
xor XOR2 (N21870, N21866, N4329);
nand NAND3 (N21871, N21859, N3436, N5510);
nand NAND4 (N21872, N21849, N15517, N21697, N4317);
nor NOR4 (N21873, N21856, N7708, N20710, N12578);
xor XOR2 (N21874, N21870, N4509);
or OR3 (N21875, N21871, N15958, N7335);
nor NOR3 (N21876, N21854, N16589, N18039);
and AND3 (N21877, N21868, N4497, N13404);
nor NOR3 (N21878, N21865, N14977, N16786);
nand NAND3 (N21879, N21869, N11740, N17926);
nor NOR3 (N21880, N21864, N8200, N1084);
or OR2 (N21881, N21879, N17827);
not NOT1 (N21882, N21875);
nor NOR4 (N21883, N21882, N15871, N11053, N7366);
buf BUF1 (N21884, N21863);
nor NOR2 (N21885, N21876, N19887);
nor NOR3 (N21886, N21874, N6295, N13984);
buf BUF1 (N21887, N21881);
or OR3 (N21888, N21884, N7133, N15498);
buf BUF1 (N21889, N21877);
nand NAND3 (N21890, N21873, N4928, N19774);
nand NAND4 (N21891, N21883, N17827, N12421, N6128);
buf BUF1 (N21892, N21886);
buf BUF1 (N21893, N21887);
xor XOR2 (N21894, N21889, N15180);
not NOT1 (N21895, N21892);
and AND4 (N21896, N21890, N17966, N6358, N13323);
and AND3 (N21897, N21891, N3943, N14002);
nor NOR3 (N21898, N21894, N699, N12380);
and AND2 (N21899, N21872, N11460);
nor NOR4 (N21900, N21878, N4823, N885, N6971);
nand NAND4 (N21901, N21880, N17875, N17646, N3632);
and AND4 (N21902, N21898, N3707, N17866, N2612);
xor XOR2 (N21903, N21901, N14187);
nand NAND2 (N21904, N21895, N16898);
or OR2 (N21905, N21893, N1741);
nor NOR2 (N21906, N21902, N3346);
xor XOR2 (N21907, N21904, N19279);
xor XOR2 (N21908, N21906, N13304);
nor NOR2 (N21909, N21903, N1081);
and AND2 (N21910, N21907, N10268);
xor XOR2 (N21911, N21888, N16416);
and AND2 (N21912, N21896, N1481);
buf BUF1 (N21913, N21897);
nand NAND4 (N21914, N21911, N3027, N2216, N17266);
xor XOR2 (N21915, N21900, N11653);
or OR2 (N21916, N21913, N12658);
nor NOR2 (N21917, N21909, N12094);
and AND4 (N21918, N21899, N15259, N16008, N2502);
nand NAND4 (N21919, N21905, N11301, N13085, N2487);
buf BUF1 (N21920, N21917);
or OR2 (N21921, N21908, N769);
nand NAND3 (N21922, N21915, N13260, N10824);
xor XOR2 (N21923, N21885, N9775);
or OR2 (N21924, N21910, N3126);
xor XOR2 (N21925, N21918, N18666);
not NOT1 (N21926, N21922);
or OR4 (N21927, N21920, N5928, N9837, N18380);
nand NAND3 (N21928, N21926, N15424, N2572);
nand NAND3 (N21929, N21927, N5378, N12070);
buf BUF1 (N21930, N21929);
and AND3 (N21931, N21930, N21718, N21823);
buf BUF1 (N21932, N21931);
nand NAND3 (N21933, N21914, N12182, N17060);
buf BUF1 (N21934, N21912);
nor NOR4 (N21935, N21933, N5406, N15532, N5683);
buf BUF1 (N21936, N21934);
xor XOR2 (N21937, N21925, N20245);
xor XOR2 (N21938, N21916, N12351);
nand NAND3 (N21939, N21938, N15675, N5192);
xor XOR2 (N21940, N21936, N6661);
buf BUF1 (N21941, N21935);
buf BUF1 (N21942, N21921);
or OR3 (N21943, N21924, N2667, N2892);
not NOT1 (N21944, N21937);
nand NAND2 (N21945, N21923, N2306);
not NOT1 (N21946, N21944);
nor NOR3 (N21947, N21946, N14377, N7904);
and AND3 (N21948, N21942, N19545, N7226);
nand NAND4 (N21949, N21932, N20950, N16528, N9266);
and AND2 (N21950, N21919, N6396);
not NOT1 (N21951, N21950);
nor NOR2 (N21952, N21945, N8321);
not NOT1 (N21953, N21940);
or OR4 (N21954, N21947, N8464, N15213, N19020);
nand NAND4 (N21955, N21948, N13232, N14557, N18168);
not NOT1 (N21956, N21953);
nor NOR4 (N21957, N21949, N11662, N711, N21592);
and AND4 (N21958, N21956, N12338, N13228, N18114);
not NOT1 (N21959, N21957);
xor XOR2 (N21960, N21941, N21178);
nand NAND4 (N21961, N21952, N15541, N4330, N18123);
xor XOR2 (N21962, N21961, N4534);
nor NOR2 (N21963, N21962, N11502);
nor NOR2 (N21964, N21958, N14048);
nor NOR3 (N21965, N21964, N487, N6066);
nor NOR3 (N21966, N21965, N6365, N6293);
buf BUF1 (N21967, N21928);
or OR4 (N21968, N21959, N15591, N12791, N8386);
nand NAND3 (N21969, N21963, N4823, N15995);
buf BUF1 (N21970, N21968);
or OR3 (N21971, N21969, N15745, N4966);
or OR3 (N21972, N21939, N9366, N6926);
buf BUF1 (N21973, N21972);
not NOT1 (N21974, N21943);
not NOT1 (N21975, N21974);
xor XOR2 (N21976, N21960, N19356);
or OR4 (N21977, N21967, N13731, N9722, N11802);
nand NAND2 (N21978, N21951, N1098);
and AND2 (N21979, N21975, N1589);
and AND2 (N21980, N21971, N10736);
nor NOR4 (N21981, N21977, N11021, N17102, N1979);
and AND3 (N21982, N21979, N20823, N11600);
not NOT1 (N21983, N21973);
buf BUF1 (N21984, N21981);
nand NAND2 (N21985, N21982, N267);
and AND4 (N21986, N21966, N5833, N6955, N7092);
xor XOR2 (N21987, N21983, N16581);
buf BUF1 (N21988, N21984);
nand NAND2 (N21989, N21985, N9749);
nand NAND3 (N21990, N21986, N18033, N14009);
and AND4 (N21991, N21988, N14017, N3084, N6228);
or OR3 (N21992, N21954, N18735, N4574);
nor NOR2 (N21993, N21970, N12541);
nand NAND4 (N21994, N21978, N7601, N15805, N234);
buf BUF1 (N21995, N21992);
nand NAND4 (N21996, N21976, N10091, N10081, N11861);
xor XOR2 (N21997, N21990, N122);
nand NAND3 (N21998, N21989, N17242, N11529);
and AND3 (N21999, N21987, N13151, N15503);
nor NOR4 (N22000, N21998, N21910, N20309, N16735);
nand NAND3 (N22001, N22000, N6583, N564);
xor XOR2 (N22002, N21999, N21771);
nor NOR4 (N22003, N21955, N14250, N8462, N14923);
nand NAND4 (N22004, N21993, N8024, N3094, N19171);
xor XOR2 (N22005, N22002, N2112);
and AND3 (N22006, N21997, N10593, N16117);
and AND2 (N22007, N21980, N16977);
nor NOR4 (N22008, N21994, N12808, N17667, N8442);
and AND3 (N22009, N22004, N13289, N10958);
or OR3 (N22010, N21996, N3595, N16384);
nand NAND3 (N22011, N22005, N15773, N6855);
nor NOR3 (N22012, N22006, N314, N1074);
or OR3 (N22013, N22007, N21407, N21402);
and AND2 (N22014, N22008, N9588);
nor NOR4 (N22015, N22003, N4731, N3167, N3378);
buf BUF1 (N22016, N22010);
buf BUF1 (N22017, N22012);
and AND4 (N22018, N21991, N9377, N6337, N25);
nor NOR2 (N22019, N22013, N3209);
buf BUF1 (N22020, N22015);
xor XOR2 (N22021, N22019, N4300);
not NOT1 (N22022, N22014);
or OR4 (N22023, N22009, N9833, N16543, N14130);
nand NAND3 (N22024, N22018, N4561, N5263);
not NOT1 (N22025, N22011);
or OR2 (N22026, N22017, N7156);
or OR4 (N22027, N22021, N15136, N11007, N21174);
not NOT1 (N22028, N22023);
and AND2 (N22029, N22027, N8454);
not NOT1 (N22030, N22025);
and AND3 (N22031, N22028, N19869, N6246);
nor NOR4 (N22032, N22016, N20097, N20103, N11676);
nand NAND4 (N22033, N22022, N332, N21299, N12092);
or OR2 (N22034, N22033, N10293);
and AND4 (N22035, N22029, N8570, N15023, N15841);
nand NAND3 (N22036, N22001, N5905, N14670);
nor NOR4 (N22037, N22026, N19102, N3051, N21466);
nand NAND2 (N22038, N22037, N15120);
and AND3 (N22039, N22035, N13722, N9369);
or OR4 (N22040, N22036, N4702, N6273, N3438);
or OR3 (N22041, N22040, N15017, N14264);
not NOT1 (N22042, N21995);
buf BUF1 (N22043, N22020);
xor XOR2 (N22044, N22039, N5202);
nor NOR4 (N22045, N22041, N16143, N18786, N21438);
nor NOR3 (N22046, N22030, N13992, N15937);
not NOT1 (N22047, N22034);
buf BUF1 (N22048, N22046);
and AND3 (N22049, N22032, N158, N429);
and AND3 (N22050, N22031, N5056, N15269);
nand NAND4 (N22051, N22038, N15008, N1122, N2295);
and AND4 (N22052, N22051, N10003, N1537, N6247);
buf BUF1 (N22053, N22042);
buf BUF1 (N22054, N22052);
and AND3 (N22055, N22047, N13091, N7599);
not NOT1 (N22056, N22044);
or OR2 (N22057, N22043, N20031);
nor NOR3 (N22058, N22053, N14356, N15037);
buf BUF1 (N22059, N22055);
buf BUF1 (N22060, N22050);
or OR3 (N22061, N22060, N13617, N11715);
not NOT1 (N22062, N22048);
not NOT1 (N22063, N22057);
nand NAND2 (N22064, N22061, N1413);
and AND2 (N22065, N22056, N8315);
not NOT1 (N22066, N22045);
or OR4 (N22067, N22062, N5829, N14519, N12732);
xor XOR2 (N22068, N22024, N15164);
nor NOR4 (N22069, N22058, N9508, N17070, N796);
and AND2 (N22070, N22067, N2385);
nor NOR3 (N22071, N22049, N21794, N11945);
nand NAND4 (N22072, N22063, N19075, N8787, N7342);
nand NAND3 (N22073, N22072, N6554, N16220);
or OR2 (N22074, N22059, N1509);
nor NOR3 (N22075, N22071, N16105, N1755);
nor NOR2 (N22076, N22073, N20253);
nor NOR2 (N22077, N22054, N17266);
or OR2 (N22078, N22064, N15774);
nor NOR2 (N22079, N22065, N20699);
and AND4 (N22080, N22076, N1098, N4578, N3798);
and AND2 (N22081, N22066, N7209);
buf BUF1 (N22082, N22079);
not NOT1 (N22083, N22074);
xor XOR2 (N22084, N22082, N17925);
not NOT1 (N22085, N22081);
nor NOR3 (N22086, N22084, N11863, N10552);
or OR4 (N22087, N22069, N7104, N7931, N4116);
or OR3 (N22088, N22085, N4, N11940);
xor XOR2 (N22089, N22086, N5576);
buf BUF1 (N22090, N22070);
buf BUF1 (N22091, N22080);
nor NOR2 (N22092, N22078, N15752);
not NOT1 (N22093, N22077);
buf BUF1 (N22094, N22090);
xor XOR2 (N22095, N22092, N13399);
nand NAND2 (N22096, N22094, N1498);
not NOT1 (N22097, N22088);
or OR2 (N22098, N22068, N12980);
xor XOR2 (N22099, N22075, N11959);
nand NAND3 (N22100, N22089, N4129, N1885);
or OR2 (N22101, N22095, N7652);
not NOT1 (N22102, N22101);
xor XOR2 (N22103, N22099, N20773);
xor XOR2 (N22104, N22096, N9397);
nand NAND4 (N22105, N22093, N8737, N6387, N5924);
and AND4 (N22106, N22100, N15472, N4368, N12614);
not NOT1 (N22107, N22105);
or OR4 (N22108, N22104, N5358, N6502, N14825);
xor XOR2 (N22109, N22106, N6462);
buf BUF1 (N22110, N22103);
not NOT1 (N22111, N22108);
and AND2 (N22112, N22109, N18459);
nand NAND4 (N22113, N22111, N9747, N11089, N21334);
or OR4 (N22114, N22112, N21595, N17743, N2455);
xor XOR2 (N22115, N22113, N10505);
xor XOR2 (N22116, N22102, N5910);
or OR3 (N22117, N22107, N3202, N590);
nor NOR3 (N22118, N22097, N13419, N9769);
or OR4 (N22119, N22114, N20404, N7588, N20664);
and AND4 (N22120, N22083, N7472, N13802, N12796);
nor NOR4 (N22121, N22115, N18094, N19258, N30);
and AND3 (N22122, N22118, N20325, N15903);
xor XOR2 (N22123, N22110, N5597);
buf BUF1 (N22124, N22121);
nand NAND4 (N22125, N22123, N21586, N20809, N14920);
and AND3 (N22126, N22124, N17871, N6950);
and AND2 (N22127, N22091, N16916);
buf BUF1 (N22128, N22117);
xor XOR2 (N22129, N22087, N16230);
and AND4 (N22130, N22128, N2763, N12359, N10006);
or OR3 (N22131, N22126, N16712, N11296);
xor XOR2 (N22132, N22127, N19760);
nor NOR3 (N22133, N22119, N10508, N18858);
and AND3 (N22134, N22116, N8436, N16370);
xor XOR2 (N22135, N22130, N14759);
xor XOR2 (N22136, N22132, N2799);
and AND3 (N22137, N22122, N15701, N8614);
not NOT1 (N22138, N22137);
or OR2 (N22139, N22136, N3166);
not NOT1 (N22140, N22120);
or OR4 (N22141, N22135, N1198, N8766, N12821);
buf BUF1 (N22142, N22140);
xor XOR2 (N22143, N22131, N2339);
or OR4 (N22144, N22138, N16899, N13440, N4617);
not NOT1 (N22145, N22142);
or OR3 (N22146, N22145, N5272, N909);
xor XOR2 (N22147, N22098, N6072);
not NOT1 (N22148, N22141);
buf BUF1 (N22149, N22144);
not NOT1 (N22150, N22149);
buf BUF1 (N22151, N22133);
buf BUF1 (N22152, N22143);
nand NAND2 (N22153, N22150, N16412);
nand NAND4 (N22154, N22146, N12612, N9555, N21305);
or OR3 (N22155, N22129, N16153, N13818);
not NOT1 (N22156, N22153);
nand NAND4 (N22157, N22156, N16358, N1771, N14705);
xor XOR2 (N22158, N22151, N20921);
buf BUF1 (N22159, N22158);
nor NOR2 (N22160, N22134, N6766);
or OR2 (N22161, N22125, N13506);
not NOT1 (N22162, N22154);
buf BUF1 (N22163, N22159);
xor XOR2 (N22164, N22139, N15149);
not NOT1 (N22165, N22160);
buf BUF1 (N22166, N22157);
nand NAND4 (N22167, N22155, N10653, N8046, N5098);
nand NAND2 (N22168, N22152, N19778);
xor XOR2 (N22169, N22168, N4704);
nand NAND2 (N22170, N22162, N13449);
nand NAND3 (N22171, N22167, N20718, N15539);
buf BUF1 (N22172, N22161);
not NOT1 (N22173, N22147);
buf BUF1 (N22174, N22166);
and AND4 (N22175, N22164, N7650, N14881, N5696);
buf BUF1 (N22176, N22165);
nand NAND4 (N22177, N22172, N4605, N21178, N11798);
not NOT1 (N22178, N22173);
not NOT1 (N22179, N22170);
buf BUF1 (N22180, N22171);
not NOT1 (N22181, N22178);
nand NAND2 (N22182, N22163, N7084);
not NOT1 (N22183, N22180);
not NOT1 (N22184, N22181);
xor XOR2 (N22185, N22184, N18640);
buf BUF1 (N22186, N22169);
and AND4 (N22187, N22177, N7298, N9165, N6430);
nand NAND4 (N22188, N22187, N21441, N13603, N15043);
not NOT1 (N22189, N22179);
nor NOR2 (N22190, N22188, N5111);
buf BUF1 (N22191, N22174);
nand NAND3 (N22192, N22183, N1100, N10789);
and AND4 (N22193, N22176, N11638, N10695, N16698);
buf BUF1 (N22194, N22193);
not NOT1 (N22195, N22175);
xor XOR2 (N22196, N22189, N9618);
buf BUF1 (N22197, N22185);
xor XOR2 (N22198, N22148, N3620);
and AND4 (N22199, N22182, N14195, N20078, N18898);
buf BUF1 (N22200, N22191);
buf BUF1 (N22201, N22192);
nor NOR4 (N22202, N22197, N4509, N14575, N12973);
not NOT1 (N22203, N22195);
not NOT1 (N22204, N22201);
and AND4 (N22205, N22194, N10357, N11008, N10193);
buf BUF1 (N22206, N22198);
buf BUF1 (N22207, N22202);
xor XOR2 (N22208, N22196, N19439);
or OR3 (N22209, N22204, N17811, N16504);
and AND2 (N22210, N22207, N3377);
xor XOR2 (N22211, N22190, N1896);
nand NAND3 (N22212, N22203, N14842, N18701);
nand NAND2 (N22213, N22211, N2246);
or OR3 (N22214, N22206, N20081, N8731);
xor XOR2 (N22215, N22186, N13953);
buf BUF1 (N22216, N22214);
buf BUF1 (N22217, N22212);
nor NOR3 (N22218, N22210, N16055, N20234);
nor NOR2 (N22219, N22200, N15946);
not NOT1 (N22220, N22217);
and AND4 (N22221, N22218, N6764, N2068, N17637);
buf BUF1 (N22222, N22215);
xor XOR2 (N22223, N22209, N6586);
or OR3 (N22224, N22221, N20218, N6515);
nor NOR2 (N22225, N22220, N21855);
nor NOR4 (N22226, N22213, N16521, N15499, N5609);
and AND2 (N22227, N22205, N17781);
nor NOR4 (N22228, N22199, N13734, N6070, N3744);
nor NOR2 (N22229, N22227, N11859);
nand NAND2 (N22230, N22208, N11472);
nor NOR2 (N22231, N22224, N2408);
nor NOR3 (N22232, N22219, N7384, N19442);
xor XOR2 (N22233, N22226, N1658);
nor NOR3 (N22234, N22233, N22211, N16640);
buf BUF1 (N22235, N22234);
nand NAND4 (N22236, N22222, N3366, N4638, N6897);
not NOT1 (N22237, N22228);
nor NOR4 (N22238, N22216, N12248, N6912, N4535);
buf BUF1 (N22239, N22231);
xor XOR2 (N22240, N22236, N13351);
nand NAND3 (N22241, N22235, N22222, N16893);
or OR2 (N22242, N22223, N16727);
not NOT1 (N22243, N22239);
nor NOR3 (N22244, N22240, N17173, N9280);
and AND2 (N22245, N22238, N5568);
xor XOR2 (N22246, N22225, N4892);
or OR3 (N22247, N22244, N1131, N2659);
not NOT1 (N22248, N22229);
nor NOR3 (N22249, N22242, N21181, N16141);
or OR2 (N22250, N22237, N10812);
buf BUF1 (N22251, N22241);
not NOT1 (N22252, N22249);
and AND3 (N22253, N22247, N15003, N19986);
or OR3 (N22254, N22246, N18119, N2675);
buf BUF1 (N22255, N22245);
buf BUF1 (N22256, N22250);
or OR3 (N22257, N22248, N2549, N6883);
buf BUF1 (N22258, N22256);
buf BUF1 (N22259, N22252);
or OR4 (N22260, N22254, N15844, N12713, N3465);
nand NAND4 (N22261, N22260, N12872, N21577, N19424);
nor NOR3 (N22262, N22251, N20251, N5822);
buf BUF1 (N22263, N22232);
nor NOR4 (N22264, N22259, N14252, N17035, N17659);
or OR3 (N22265, N22255, N5008, N11399);
or OR4 (N22266, N22243, N9293, N2518, N19042);
or OR3 (N22267, N22230, N8022, N8789);
nor NOR4 (N22268, N22253, N16474, N3182, N5050);
nand NAND4 (N22269, N22265, N12005, N3461, N20496);
buf BUF1 (N22270, N22269);
nand NAND2 (N22271, N22270, N12193);
and AND3 (N22272, N22257, N7444, N14790);
and AND2 (N22273, N22262, N21510);
nor NOR3 (N22274, N22264, N386, N992);
xor XOR2 (N22275, N22274, N20837);
and AND3 (N22276, N22275, N4303, N16307);
nor NOR2 (N22277, N22273, N21329);
buf BUF1 (N22278, N22261);
xor XOR2 (N22279, N22267, N11340);
xor XOR2 (N22280, N22263, N20504);
xor XOR2 (N22281, N22278, N5711);
not NOT1 (N22282, N22266);
not NOT1 (N22283, N22271);
nor NOR2 (N22284, N22268, N13683);
and AND3 (N22285, N22282, N8503, N13143);
and AND2 (N22286, N22285, N828);
or OR4 (N22287, N22276, N21726, N18775, N13560);
or OR4 (N22288, N22280, N3279, N263, N10579);
nand NAND3 (N22289, N22277, N10214, N11593);
not NOT1 (N22290, N22281);
xor XOR2 (N22291, N22284, N7706);
xor XOR2 (N22292, N22286, N4927);
not NOT1 (N22293, N22289);
and AND2 (N22294, N22290, N7262);
or OR3 (N22295, N22291, N6720, N17792);
buf BUF1 (N22296, N22293);
nand NAND2 (N22297, N22295, N10616);
xor XOR2 (N22298, N22287, N5937);
nand NAND3 (N22299, N22258, N8192, N9413);
or OR2 (N22300, N22288, N11577);
nor NOR4 (N22301, N22297, N20139, N8732, N8965);
not NOT1 (N22302, N22294);
and AND3 (N22303, N22298, N6648, N5990);
nand NAND2 (N22304, N22283, N646);
and AND3 (N22305, N22304, N8632, N3868);
xor XOR2 (N22306, N22303, N21899);
xor XOR2 (N22307, N22299, N19158);
and AND4 (N22308, N22279, N9607, N1963, N10250);
nand NAND2 (N22309, N22306, N11431);
or OR4 (N22310, N22302, N19596, N10968, N9206);
and AND2 (N22311, N22307, N3728);
and AND3 (N22312, N22292, N1636, N11871);
or OR4 (N22313, N22296, N14225, N3517, N3895);
or OR4 (N22314, N22305, N6953, N4675, N5930);
not NOT1 (N22315, N22272);
or OR3 (N22316, N22312, N2237, N5331);
and AND4 (N22317, N22311, N2448, N4565, N15053);
and AND3 (N22318, N22308, N18996, N15105);
nor NOR2 (N22319, N22315, N20733);
buf BUF1 (N22320, N22300);
and AND4 (N22321, N22319, N16518, N16945, N19136);
nand NAND4 (N22322, N22313, N3266, N13671, N319);
nand NAND2 (N22323, N22321, N19900);
buf BUF1 (N22324, N22310);
xor XOR2 (N22325, N22301, N1596);
nand NAND4 (N22326, N22317, N19238, N9357, N10932);
not NOT1 (N22327, N22320);
nand NAND2 (N22328, N22326, N5555);
nor NOR2 (N22329, N22314, N4246);
nor NOR2 (N22330, N22316, N14996);
or OR3 (N22331, N22324, N7102, N11100);
xor XOR2 (N22332, N22318, N1318);
or OR2 (N22333, N22322, N11520);
xor XOR2 (N22334, N22332, N9230);
xor XOR2 (N22335, N22334, N21865);
and AND2 (N22336, N22328, N11357);
nand NAND2 (N22337, N22330, N9603);
and AND2 (N22338, N22309, N2598);
nand NAND4 (N22339, N22329, N138, N11328, N21359);
xor XOR2 (N22340, N22336, N5607);
nand NAND3 (N22341, N22323, N8113, N3545);
nand NAND3 (N22342, N22339, N22259, N12016);
or OR4 (N22343, N22340, N2151, N2007, N7379);
nor NOR3 (N22344, N22343, N170, N16613);
or OR3 (N22345, N22333, N6284, N20814);
buf BUF1 (N22346, N22331);
nor NOR2 (N22347, N22335, N2070);
and AND2 (N22348, N22342, N5577);
not NOT1 (N22349, N22337);
nor NOR3 (N22350, N22341, N12798, N22007);
nor NOR4 (N22351, N22325, N16659, N14731, N18315);
xor XOR2 (N22352, N22344, N8289);
xor XOR2 (N22353, N22346, N21127);
nand NAND2 (N22354, N22350, N19268);
or OR2 (N22355, N22338, N18662);
not NOT1 (N22356, N22354);
or OR2 (N22357, N22352, N6216);
not NOT1 (N22358, N22349);
buf BUF1 (N22359, N22327);
xor XOR2 (N22360, N22359, N8141);
nor NOR4 (N22361, N22360, N16136, N18095, N3245);
and AND3 (N22362, N22361, N20335, N21022);
buf BUF1 (N22363, N22347);
xor XOR2 (N22364, N22351, N10339);
xor XOR2 (N22365, N22358, N20232);
buf BUF1 (N22366, N22355);
not NOT1 (N22367, N22356);
xor XOR2 (N22368, N22363, N12938);
not NOT1 (N22369, N22348);
and AND3 (N22370, N22345, N4379, N19405);
nand NAND2 (N22371, N22357, N16043);
nor NOR2 (N22372, N22366, N15578);
or OR4 (N22373, N22372, N21806, N21223, N17508);
buf BUF1 (N22374, N22367);
nor NOR4 (N22375, N22362, N20918, N4803, N1779);
and AND2 (N22376, N22375, N3973);
nor NOR2 (N22377, N22369, N6371);
or OR4 (N22378, N22377, N15579, N10059, N6698);
or OR2 (N22379, N22378, N20212);
nor NOR4 (N22380, N22379, N20311, N21099, N9331);
xor XOR2 (N22381, N22370, N17211);
and AND2 (N22382, N22380, N11116);
nor NOR3 (N22383, N22368, N10308, N13574);
buf BUF1 (N22384, N22365);
nor NOR3 (N22385, N22384, N8229, N21654);
xor XOR2 (N22386, N22373, N9217);
buf BUF1 (N22387, N22382);
and AND3 (N22388, N22376, N14949, N7816);
buf BUF1 (N22389, N22385);
nand NAND2 (N22390, N22374, N16273);
nand NAND4 (N22391, N22387, N21663, N20754, N12123);
not NOT1 (N22392, N22371);
xor XOR2 (N22393, N22390, N291);
not NOT1 (N22394, N22353);
nor NOR3 (N22395, N22386, N10526, N12578);
and AND4 (N22396, N22383, N2001, N20201, N12143);
and AND2 (N22397, N22391, N842);
not NOT1 (N22398, N22392);
and AND3 (N22399, N22364, N2098, N15786);
or OR2 (N22400, N22381, N18633);
and AND4 (N22401, N22397, N15804, N11100, N22279);
nand NAND4 (N22402, N22394, N7671, N15024, N11682);
and AND3 (N22403, N22389, N430, N20891);
or OR4 (N22404, N22388, N10104, N22124, N14136);
nand NAND2 (N22405, N22395, N16060);
not NOT1 (N22406, N22405);
and AND3 (N22407, N22398, N8639, N11729);
not NOT1 (N22408, N22402);
nor NOR4 (N22409, N22400, N8143, N3024, N3937);
xor XOR2 (N22410, N22406, N11927);
nor NOR4 (N22411, N22408, N19207, N18644, N11246);
buf BUF1 (N22412, N22403);
xor XOR2 (N22413, N22404, N15172);
buf BUF1 (N22414, N22393);
or OR4 (N22415, N22407, N16905, N20243, N14311);
nor NOR2 (N22416, N22396, N12517);
nand NAND3 (N22417, N22414, N16709, N9627);
or OR4 (N22418, N22413, N1958, N295, N584);
nand NAND2 (N22419, N22409, N19241);
and AND3 (N22420, N22418, N18263, N16662);
buf BUF1 (N22421, N22417);
or OR2 (N22422, N22411, N10165);
nand NAND4 (N22423, N22419, N16112, N6571, N16887);
xor XOR2 (N22424, N22415, N16832);
and AND3 (N22425, N22410, N4751, N5888);
not NOT1 (N22426, N22423);
xor XOR2 (N22427, N22412, N12194);
nor NOR3 (N22428, N22422, N6026, N10077);
not NOT1 (N22429, N22421);
nand NAND4 (N22430, N22429, N8793, N2410, N18952);
and AND4 (N22431, N22420, N12629, N22178, N18053);
and AND4 (N22432, N22416, N20852, N10922, N14652);
or OR2 (N22433, N22426, N13222);
not NOT1 (N22434, N22430);
xor XOR2 (N22435, N22401, N843);
nor NOR2 (N22436, N22399, N14205);
not NOT1 (N22437, N22433);
or OR3 (N22438, N22431, N3330, N5484);
not NOT1 (N22439, N22428);
not NOT1 (N22440, N22437);
or OR2 (N22441, N22425, N17342);
not NOT1 (N22442, N22434);
nand NAND2 (N22443, N22424, N11324);
not NOT1 (N22444, N22432);
or OR3 (N22445, N22435, N17382, N18780);
buf BUF1 (N22446, N22427);
xor XOR2 (N22447, N22446, N7088);
and AND3 (N22448, N22443, N14300, N8929);
and AND3 (N22449, N22439, N21142, N1940);
not NOT1 (N22450, N22438);
and AND3 (N22451, N22436, N6044, N17853);
buf BUF1 (N22452, N22447);
nand NAND2 (N22453, N22441, N11384);
nand NAND2 (N22454, N22440, N9958);
buf BUF1 (N22455, N22451);
nand NAND4 (N22456, N22442, N14746, N16609, N3850);
buf BUF1 (N22457, N22454);
buf BUF1 (N22458, N22444);
buf BUF1 (N22459, N22450);
and AND3 (N22460, N22456, N13246, N7590);
and AND4 (N22461, N22453, N15717, N15145, N17141);
nor NOR3 (N22462, N22448, N14274, N17846);
nand NAND4 (N22463, N22461, N279, N21024, N4059);
nor NOR4 (N22464, N22458, N6830, N12294, N8769);
nand NAND4 (N22465, N22455, N19024, N11917, N20208);
nand NAND2 (N22466, N22452, N9438);
xor XOR2 (N22467, N22464, N21144);
and AND4 (N22468, N22459, N5455, N11841, N9606);
buf BUF1 (N22469, N22462);
buf BUF1 (N22470, N22465);
and AND2 (N22471, N22468, N14060);
or OR3 (N22472, N22449, N4703, N3831);
not NOT1 (N22473, N22470);
and AND2 (N22474, N22463, N9301);
xor XOR2 (N22475, N22467, N17825);
buf BUF1 (N22476, N22445);
nor NOR2 (N22477, N22471, N121);
buf BUF1 (N22478, N22475);
not NOT1 (N22479, N22472);
nor NOR4 (N22480, N22478, N18091, N3078, N1911);
and AND3 (N22481, N22457, N20345, N2043);
nand NAND3 (N22482, N22460, N12571, N21447);
nand NAND3 (N22483, N22481, N14870, N22378);
and AND2 (N22484, N22479, N20193);
and AND4 (N22485, N22469, N2205, N8, N15399);
or OR2 (N22486, N22477, N4133);
not NOT1 (N22487, N22466);
nand NAND2 (N22488, N22480, N10284);
xor XOR2 (N22489, N22476, N8504);
or OR2 (N22490, N22489, N6546);
nand NAND3 (N22491, N22484, N19291, N787);
xor XOR2 (N22492, N22487, N16960);
xor XOR2 (N22493, N22482, N15209);
xor XOR2 (N22494, N22493, N19243);
not NOT1 (N22495, N22492);
nor NOR4 (N22496, N22485, N10583, N9571, N11928);
buf BUF1 (N22497, N22494);
or OR2 (N22498, N22486, N5039);
or OR4 (N22499, N22473, N12134, N16528, N11495);
not NOT1 (N22500, N22474);
nor NOR4 (N22501, N22496, N5445, N21199, N11788);
buf BUF1 (N22502, N22483);
buf BUF1 (N22503, N22495);
not NOT1 (N22504, N22500);
or OR4 (N22505, N22499, N15468, N15511, N10167);
and AND3 (N22506, N22503, N4524, N19164);
nor NOR3 (N22507, N22502, N4380, N6188);
xor XOR2 (N22508, N22498, N20265);
or OR3 (N22509, N22497, N15608, N17708);
or OR4 (N22510, N22488, N22377, N6921, N7579);
buf BUF1 (N22511, N22491);
not NOT1 (N22512, N22501);
buf BUF1 (N22513, N22507);
nand NAND3 (N22514, N22513, N15825, N22035);
nor NOR3 (N22515, N22511, N17825, N8891);
not NOT1 (N22516, N22509);
nor NOR2 (N22517, N22490, N19480);
not NOT1 (N22518, N22516);
nand NAND2 (N22519, N22508, N13289);
and AND2 (N22520, N22505, N1131);
not NOT1 (N22521, N22514);
or OR2 (N22522, N22518, N14171);
nor NOR3 (N22523, N22517, N11182, N18736);
and AND3 (N22524, N22510, N20300, N6158);
buf BUF1 (N22525, N22522);
or OR3 (N22526, N22524, N10471, N9105);
not NOT1 (N22527, N22520);
not NOT1 (N22528, N22506);
xor XOR2 (N22529, N22527, N10121);
nand NAND2 (N22530, N22512, N19442);
nor NOR2 (N22531, N22530, N14344);
not NOT1 (N22532, N22531);
not NOT1 (N22533, N22526);
and AND3 (N22534, N22525, N21295, N4912);
and AND4 (N22535, N22521, N20763, N18735, N416);
nor NOR4 (N22536, N22528, N305, N15512, N1728);
not NOT1 (N22537, N22534);
or OR4 (N22538, N22504, N2232, N16489, N16255);
and AND4 (N22539, N22537, N14455, N17616, N10194);
or OR4 (N22540, N22523, N14288, N21823, N9452);
buf BUF1 (N22541, N22519);
buf BUF1 (N22542, N22539);
and AND3 (N22543, N22542, N14473, N6928);
buf BUF1 (N22544, N22535);
buf BUF1 (N22545, N22515);
nand NAND3 (N22546, N22532, N6244, N20983);
and AND3 (N22547, N22536, N19115, N10259);
nor NOR4 (N22548, N22545, N14179, N16250, N19034);
nand NAND2 (N22549, N22541, N22441);
and AND2 (N22550, N22544, N12932);
not NOT1 (N22551, N22547);
xor XOR2 (N22552, N22543, N21954);
xor XOR2 (N22553, N22551, N20739);
xor XOR2 (N22554, N22540, N1727);
nand NAND2 (N22555, N22554, N16009);
xor XOR2 (N22556, N22546, N1218);
not NOT1 (N22557, N22552);
or OR4 (N22558, N22557, N6766, N8829, N16961);
nand NAND4 (N22559, N22533, N16342, N1889, N21303);
xor XOR2 (N22560, N22553, N6075);
nor NOR3 (N22561, N22550, N15752, N4284);
nand NAND4 (N22562, N22549, N20521, N5818, N18458);
nor NOR3 (N22563, N22562, N22059, N22468);
not NOT1 (N22564, N22558);
buf BUF1 (N22565, N22559);
nand NAND4 (N22566, N22555, N17440, N19728, N4435);
and AND2 (N22567, N22563, N960);
buf BUF1 (N22568, N22567);
nor NOR4 (N22569, N22560, N20129, N8388, N5469);
and AND3 (N22570, N22564, N14569, N19356);
nand NAND2 (N22571, N22561, N20916);
nor NOR2 (N22572, N22566, N19737);
not NOT1 (N22573, N22565);
nor NOR3 (N22574, N22569, N5115, N21811);
not NOT1 (N22575, N22573);
buf BUF1 (N22576, N22548);
or OR3 (N22577, N22568, N13713, N4602);
not NOT1 (N22578, N22529);
xor XOR2 (N22579, N22556, N6456);
not NOT1 (N22580, N22570);
buf BUF1 (N22581, N22572);
buf BUF1 (N22582, N22579);
xor XOR2 (N22583, N22578, N10616);
buf BUF1 (N22584, N22583);
or OR3 (N22585, N22538, N1193, N22523);
nand NAND4 (N22586, N22577, N18895, N11365, N490);
xor XOR2 (N22587, N22586, N6790);
not NOT1 (N22588, N22580);
xor XOR2 (N22589, N22582, N13431);
or OR2 (N22590, N22584, N14201);
buf BUF1 (N22591, N22587);
nand NAND4 (N22592, N22571, N5625, N12324, N15135);
xor XOR2 (N22593, N22589, N15009);
nor NOR2 (N22594, N22590, N4105);
and AND2 (N22595, N22581, N16468);
nand NAND2 (N22596, N22592, N20529);
xor XOR2 (N22597, N22596, N11842);
buf BUF1 (N22598, N22594);
and AND2 (N22599, N22585, N17667);
nand NAND2 (N22600, N22574, N17170);
xor XOR2 (N22601, N22591, N19089);
not NOT1 (N22602, N22576);
nor NOR3 (N22603, N22593, N5995, N15585);
nand NAND2 (N22604, N22575, N13946);
not NOT1 (N22605, N22598);
nand NAND2 (N22606, N22604, N17814);
nand NAND2 (N22607, N22605, N5132);
and AND3 (N22608, N22603, N7580, N6272);
not NOT1 (N22609, N22588);
buf BUF1 (N22610, N22597);
nand NAND3 (N22611, N22601, N2963, N5385);
nor NOR2 (N22612, N22602, N10826);
not NOT1 (N22613, N22606);
or OR2 (N22614, N22609, N641);
not NOT1 (N22615, N22607);
buf BUF1 (N22616, N22613);
xor XOR2 (N22617, N22615, N19382);
xor XOR2 (N22618, N22616, N917);
and AND3 (N22619, N22608, N7617, N17016);
or OR2 (N22620, N22612, N12758);
not NOT1 (N22621, N22599);
and AND3 (N22622, N22614, N9168, N7509);
or OR4 (N22623, N22621, N11009, N11837, N14662);
buf BUF1 (N22624, N22611);
not NOT1 (N22625, N22622);
buf BUF1 (N22626, N22619);
or OR4 (N22627, N22600, N16600, N4523, N3979);
nand NAND3 (N22628, N22625, N798, N19156);
not NOT1 (N22629, N22595);
xor XOR2 (N22630, N22623, N16791);
and AND3 (N22631, N22626, N1985, N8071);
xor XOR2 (N22632, N22627, N206);
buf BUF1 (N22633, N22630);
nor NOR4 (N22634, N22632, N12878, N9976, N16239);
nand NAND2 (N22635, N22629, N10601);
not NOT1 (N22636, N22620);
nand NAND3 (N22637, N22634, N14844, N5530);
xor XOR2 (N22638, N22635, N22199);
nor NOR4 (N22639, N22624, N2183, N1598, N6020);
buf BUF1 (N22640, N22628);
not NOT1 (N22641, N22638);
not NOT1 (N22642, N22641);
and AND2 (N22643, N22617, N6365);
xor XOR2 (N22644, N22640, N12420);
nor NOR2 (N22645, N22644, N6269);
xor XOR2 (N22646, N22610, N5226);
buf BUF1 (N22647, N22643);
or OR3 (N22648, N22631, N7122, N22298);
and AND2 (N22649, N22647, N14544);
nand NAND3 (N22650, N22639, N19977, N6156);
not NOT1 (N22651, N22618);
not NOT1 (N22652, N22645);
nor NOR4 (N22653, N22633, N21364, N7536, N1838);
nand NAND4 (N22654, N22646, N324, N20881, N5887);
xor XOR2 (N22655, N22649, N7562);
or OR4 (N22656, N22655, N9726, N1607, N10505);
nor NOR3 (N22657, N22653, N22395, N22248);
buf BUF1 (N22658, N22648);
nand NAND3 (N22659, N22658, N17600, N9556);
nor NOR4 (N22660, N22637, N7622, N1851, N532);
buf BUF1 (N22661, N22659);
buf BUF1 (N22662, N22642);
and AND2 (N22663, N22661, N4784);
xor XOR2 (N22664, N22660, N10991);
buf BUF1 (N22665, N22652);
nand NAND3 (N22666, N22664, N18138, N136);
nand NAND2 (N22667, N22665, N7360);
or OR2 (N22668, N22667, N22493);
nand NAND3 (N22669, N22650, N19650, N3083);
nand NAND2 (N22670, N22636, N469);
buf BUF1 (N22671, N22662);
xor XOR2 (N22672, N22666, N22383);
and AND2 (N22673, N22654, N21566);
or OR2 (N22674, N22672, N9374);
or OR4 (N22675, N22657, N22140, N12515, N19488);
nor NOR3 (N22676, N22673, N18796, N6364);
and AND4 (N22677, N22668, N2714, N22516, N3086);
xor XOR2 (N22678, N22674, N15830);
buf BUF1 (N22679, N22678);
not NOT1 (N22680, N22669);
not NOT1 (N22681, N22651);
or OR3 (N22682, N22676, N22095, N7970);
nor NOR3 (N22683, N22680, N9376, N20420);
nor NOR3 (N22684, N22682, N9884, N16250);
nor NOR4 (N22685, N22675, N20777, N20843, N12217);
or OR3 (N22686, N22670, N9643, N20839);
xor XOR2 (N22687, N22685, N15769);
nand NAND2 (N22688, N22671, N8871);
and AND3 (N22689, N22679, N13883, N2064);
nand NAND2 (N22690, N22663, N15428);
buf BUF1 (N22691, N22690);
nor NOR3 (N22692, N22656, N18428, N10748);
or OR3 (N22693, N22681, N18910, N6041);
and AND2 (N22694, N22693, N12714);
nor NOR2 (N22695, N22686, N22437);
not NOT1 (N22696, N22688);
or OR4 (N22697, N22677, N3353, N16665, N4421);
or OR3 (N22698, N22697, N15345, N1647);
nor NOR3 (N22699, N22692, N1018, N5088);
nand NAND4 (N22700, N22698, N14887, N21442, N13772);
nand NAND3 (N22701, N22691, N18632, N16748);
or OR3 (N22702, N22687, N14168, N20329);
buf BUF1 (N22703, N22695);
and AND2 (N22704, N22683, N8212);
not NOT1 (N22705, N22694);
and AND3 (N22706, N22696, N20896, N9163);
and AND3 (N22707, N22704, N6584, N17850);
buf BUF1 (N22708, N22702);
nor NOR4 (N22709, N22684, N6566, N22604, N10428);
or OR4 (N22710, N22708, N9023, N8533, N17619);
buf BUF1 (N22711, N22700);
and AND4 (N22712, N22689, N11896, N16088, N1749);
or OR2 (N22713, N22701, N3641);
nor NOR4 (N22714, N22712, N12062, N9866, N11009);
nand NAND3 (N22715, N22714, N12657, N8274);
nand NAND4 (N22716, N22703, N21969, N3964, N21952);
or OR4 (N22717, N22716, N13078, N3925, N13205);
or OR3 (N22718, N22711, N15910, N5928);
nand NAND2 (N22719, N22718, N21322);
nand NAND2 (N22720, N22715, N6067);
and AND4 (N22721, N22720, N19876, N5799, N13567);
or OR3 (N22722, N22706, N21303, N542);
or OR2 (N22723, N22721, N6308);
buf BUF1 (N22724, N22710);
buf BUF1 (N22725, N22724);
nor NOR3 (N22726, N22709, N5051, N2908);
nor NOR4 (N22727, N22726, N5422, N12539, N22470);
or OR3 (N22728, N22699, N9866, N8073);
xor XOR2 (N22729, N22725, N20500);
buf BUF1 (N22730, N22722);
not NOT1 (N22731, N22728);
nand NAND3 (N22732, N22717, N258, N18272);
xor XOR2 (N22733, N22713, N9564);
not NOT1 (N22734, N22732);
and AND3 (N22735, N22707, N6139, N8354);
nand NAND4 (N22736, N22723, N8131, N19385, N7657);
nand NAND3 (N22737, N22731, N3317, N8249);
or OR2 (N22738, N22727, N14132);
nor NOR2 (N22739, N22736, N11477);
nand NAND2 (N22740, N22705, N6630);
xor XOR2 (N22741, N22733, N3564);
not NOT1 (N22742, N22738);
buf BUF1 (N22743, N22735);
buf BUF1 (N22744, N22730);
xor XOR2 (N22745, N22744, N5417);
xor XOR2 (N22746, N22743, N7550);
xor XOR2 (N22747, N22742, N10632);
nand NAND3 (N22748, N22739, N755, N15524);
not NOT1 (N22749, N22746);
xor XOR2 (N22750, N22740, N9666);
xor XOR2 (N22751, N22719, N21409);
and AND2 (N22752, N22747, N20855);
nor NOR2 (N22753, N22737, N18914);
buf BUF1 (N22754, N22750);
nand NAND3 (N22755, N22729, N10473, N7618);
nor NOR3 (N22756, N22749, N4778, N962);
nor NOR4 (N22757, N22753, N21886, N22747, N5852);
and AND3 (N22758, N22752, N12585, N19694);
nand NAND3 (N22759, N22757, N10870, N22336);
and AND4 (N22760, N22755, N10500, N12450, N8821);
and AND2 (N22761, N22754, N1984);
and AND4 (N22762, N22741, N2673, N18248, N20053);
or OR3 (N22763, N22758, N9609, N7690);
xor XOR2 (N22764, N22759, N9546);
xor XOR2 (N22765, N22756, N15749);
buf BUF1 (N22766, N22748);
not NOT1 (N22767, N22763);
nand NAND3 (N22768, N22767, N11916, N16111);
or OR4 (N22769, N22768, N12231, N13174, N14868);
not NOT1 (N22770, N22734);
nand NAND4 (N22771, N22770, N176, N955, N12532);
nor NOR3 (N22772, N22764, N11710, N6467);
and AND4 (N22773, N22751, N12121, N17739, N15421);
nand NAND3 (N22774, N22769, N8032, N16387);
nor NOR4 (N22775, N22766, N444, N11110, N7874);
nor NOR4 (N22776, N22762, N19038, N19169, N14696);
nor NOR2 (N22777, N22771, N18800);
not NOT1 (N22778, N22745);
or OR4 (N22779, N22778, N20434, N3398, N6538);
nand NAND2 (N22780, N22776, N13718);
buf BUF1 (N22781, N22761);
nor NOR2 (N22782, N22775, N7348);
or OR2 (N22783, N22760, N14859);
nand NAND2 (N22784, N22777, N14358);
nor NOR3 (N22785, N22774, N13942, N18809);
or OR3 (N22786, N22772, N2168, N18037);
xor XOR2 (N22787, N22781, N19883);
nand NAND4 (N22788, N22779, N1234, N12088, N12378);
nor NOR3 (N22789, N22786, N2002, N5061);
or OR2 (N22790, N22787, N4714);
not NOT1 (N22791, N22782);
buf BUF1 (N22792, N22788);
nor NOR3 (N22793, N22792, N2519, N18720);
xor XOR2 (N22794, N22773, N15436);
xor XOR2 (N22795, N22794, N9025);
xor XOR2 (N22796, N22765, N4027);
nor NOR3 (N22797, N22793, N18254, N13868);
or OR2 (N22798, N22797, N6386);
or OR3 (N22799, N22798, N19638, N8218);
xor XOR2 (N22800, N22783, N8732);
nor NOR2 (N22801, N22790, N2440);
buf BUF1 (N22802, N22791);
nor NOR2 (N22803, N22802, N20367);
not NOT1 (N22804, N22803);
buf BUF1 (N22805, N22796);
nor NOR2 (N22806, N22801, N16436);
or OR4 (N22807, N22805, N22242, N8815, N2377);
nor NOR2 (N22808, N22806, N2011);
xor XOR2 (N22809, N22807, N13026);
or OR4 (N22810, N22800, N12253, N5637, N16037);
not NOT1 (N22811, N22799);
xor XOR2 (N22812, N22808, N5545);
buf BUF1 (N22813, N22804);
buf BUF1 (N22814, N22795);
buf BUF1 (N22815, N22812);
xor XOR2 (N22816, N22813, N7935);
or OR3 (N22817, N22814, N3243, N8112);
and AND4 (N22818, N22789, N19331, N20313, N11584);
or OR4 (N22819, N22785, N20649, N13047, N806);
xor XOR2 (N22820, N22818, N15434);
nand NAND3 (N22821, N22816, N21603, N10745);
buf BUF1 (N22822, N22815);
and AND2 (N22823, N22820, N20099);
xor XOR2 (N22824, N22819, N9314);
nand NAND2 (N22825, N22821, N10237);
buf BUF1 (N22826, N22809);
nand NAND2 (N22827, N22780, N1894);
nor NOR3 (N22828, N22825, N6214, N5052);
not NOT1 (N22829, N22817);
and AND4 (N22830, N22822, N17013, N15652, N18822);
nor NOR2 (N22831, N22810, N17424);
and AND3 (N22832, N22824, N3345, N9391);
nor NOR4 (N22833, N22784, N13692, N15485, N7567);
nand NAND4 (N22834, N22827, N3216, N18584, N16734);
xor XOR2 (N22835, N22811, N10398);
buf BUF1 (N22836, N22834);
and AND3 (N22837, N22836, N4643, N22122);
nand NAND4 (N22838, N22829, N1988, N18225, N16561);
nor NOR3 (N22839, N22835, N2494, N20713);
and AND2 (N22840, N22832, N22289);
xor XOR2 (N22841, N22831, N4270);
nand NAND3 (N22842, N22828, N17449, N3589);
nor NOR3 (N22843, N22826, N12141, N21914);
buf BUF1 (N22844, N22838);
not NOT1 (N22845, N22841);
and AND2 (N22846, N22840, N3207);
and AND3 (N22847, N22845, N11018, N14795);
buf BUF1 (N22848, N22842);
buf BUF1 (N22849, N22837);
not NOT1 (N22850, N22839);
nor NOR3 (N22851, N22848, N10037, N668);
buf BUF1 (N22852, N22851);
or OR3 (N22853, N22823, N4009, N3633);
and AND4 (N22854, N22833, N8893, N1256, N10042);
nor NOR4 (N22855, N22849, N21512, N2744, N9631);
nand NAND4 (N22856, N22843, N16395, N3067, N20203);
and AND2 (N22857, N22856, N14808);
xor XOR2 (N22858, N22857, N14667);
nand NAND4 (N22859, N22830, N21557, N21189, N4766);
nand NAND2 (N22860, N22853, N22709);
nor NOR3 (N22861, N22860, N5109, N1107);
nor NOR3 (N22862, N22847, N577, N22810);
and AND4 (N22863, N22862, N20084, N391, N21828);
or OR4 (N22864, N22858, N295, N14761, N15292);
buf BUF1 (N22865, N22859);
nand NAND3 (N22866, N22861, N642, N708);
nor NOR2 (N22867, N22865, N13089);
nor NOR4 (N22868, N22864, N1526, N14064, N8710);
and AND3 (N22869, N22846, N944, N2117);
buf BUF1 (N22870, N22869);
not NOT1 (N22871, N22844);
nor NOR2 (N22872, N22868, N22684);
and AND2 (N22873, N22855, N1832);
xor XOR2 (N22874, N22866, N4540);
xor XOR2 (N22875, N22863, N4404);
nand NAND3 (N22876, N22852, N6017, N1132);
buf BUF1 (N22877, N22876);
nor NOR3 (N22878, N22874, N15331, N21283);
buf BUF1 (N22879, N22871);
buf BUF1 (N22880, N22870);
and AND2 (N22881, N22878, N9258);
or OR3 (N22882, N22873, N20080, N14562);
nand NAND3 (N22883, N22872, N16612, N11790);
nand NAND3 (N22884, N22875, N3205, N16617);
or OR4 (N22885, N22877, N12841, N1836, N2659);
buf BUF1 (N22886, N22881);
buf BUF1 (N22887, N22879);
buf BUF1 (N22888, N22886);
xor XOR2 (N22889, N22883, N9935);
or OR4 (N22890, N22882, N20834, N6361, N21323);
nor NOR2 (N22891, N22867, N15691);
or OR4 (N22892, N22850, N5395, N21482, N7501);
buf BUF1 (N22893, N22880);
or OR4 (N22894, N22885, N5105, N6631, N13797);
and AND2 (N22895, N22888, N1899);
or OR4 (N22896, N22887, N6813, N22235, N393);
nor NOR3 (N22897, N22895, N18397, N14265);
not NOT1 (N22898, N22891);
buf BUF1 (N22899, N22896);
nand NAND3 (N22900, N22898, N859, N123);
nand NAND3 (N22901, N22900, N4464, N8567);
and AND2 (N22902, N22897, N20606);
not NOT1 (N22903, N22893);
nor NOR4 (N22904, N22902, N10657, N6998, N21860);
xor XOR2 (N22905, N22884, N11921);
buf BUF1 (N22906, N22892);
xor XOR2 (N22907, N22904, N5650);
or OR3 (N22908, N22899, N17318, N1678);
buf BUF1 (N22909, N22903);
nor NOR2 (N22910, N22854, N14500);
nand NAND4 (N22911, N22905, N2742, N10326, N19105);
not NOT1 (N22912, N22910);
xor XOR2 (N22913, N22906, N4971);
xor XOR2 (N22914, N22894, N7532);
and AND2 (N22915, N22908, N22198);
nor NOR3 (N22916, N22901, N1051, N10266);
not NOT1 (N22917, N22907);
and AND2 (N22918, N22911, N19546);
and AND4 (N22919, N22914, N9480, N6528, N8780);
nor NOR2 (N22920, N22916, N9824);
nand NAND3 (N22921, N22920, N21055, N5996);
or OR4 (N22922, N22919, N4361, N3902, N9887);
nor NOR4 (N22923, N22922, N8582, N758, N12185);
xor XOR2 (N22924, N22921, N13831);
not NOT1 (N22925, N22924);
and AND4 (N22926, N22909, N553, N4841, N9124);
or OR4 (N22927, N22890, N17803, N10766, N10424);
nor NOR3 (N22928, N22917, N1241, N11855);
or OR3 (N22929, N22923, N13529, N1373);
or OR3 (N22930, N22913, N18636, N3540);
not NOT1 (N22931, N22889);
or OR2 (N22932, N22927, N15155);
nor NOR3 (N22933, N22915, N395, N22539);
xor XOR2 (N22934, N22931, N13534);
nor NOR4 (N22935, N22929, N2299, N4815, N13697);
xor XOR2 (N22936, N22930, N15749);
or OR4 (N22937, N22934, N8657, N6397, N21577);
xor XOR2 (N22938, N22928, N10058);
xor XOR2 (N22939, N22926, N1975);
buf BUF1 (N22940, N22937);
nand NAND3 (N22941, N22918, N22118, N12860);
xor XOR2 (N22942, N22935, N7890);
xor XOR2 (N22943, N22936, N20311);
and AND3 (N22944, N22940, N17798, N11959);
xor XOR2 (N22945, N22938, N11870);
nand NAND4 (N22946, N22941, N1133, N1865, N11101);
xor XOR2 (N22947, N22942, N16429);
not NOT1 (N22948, N22943);
and AND2 (N22949, N22932, N3598);
and AND3 (N22950, N22949, N9466, N12766);
and AND4 (N22951, N22947, N14896, N17111, N1745);
or OR3 (N22952, N22948, N7645, N17140);
not NOT1 (N22953, N22925);
and AND3 (N22954, N22951, N5489, N21078);
or OR2 (N22955, N22912, N20943);
xor XOR2 (N22956, N22945, N10090);
not NOT1 (N22957, N22952);
buf BUF1 (N22958, N22933);
xor XOR2 (N22959, N22957, N8610);
buf BUF1 (N22960, N22954);
nor NOR2 (N22961, N22953, N7686);
nor NOR3 (N22962, N22959, N9366, N19511);
or OR2 (N22963, N22958, N16238);
buf BUF1 (N22964, N22944);
not NOT1 (N22965, N22962);
or OR3 (N22966, N22956, N21998, N20664);
and AND3 (N22967, N22963, N7584, N1284);
buf BUF1 (N22968, N22946);
or OR2 (N22969, N22950, N15297);
buf BUF1 (N22970, N22969);
buf BUF1 (N22971, N22968);
and AND2 (N22972, N22965, N8573);
buf BUF1 (N22973, N22961);
nor NOR4 (N22974, N22967, N180, N19950, N4810);
and AND4 (N22975, N22966, N913, N18416, N2948);
buf BUF1 (N22976, N22974);
nand NAND3 (N22977, N22975, N15143, N3546);
nand NAND3 (N22978, N22977, N5652, N5044);
or OR3 (N22979, N22972, N265, N3370);
or OR4 (N22980, N22960, N19224, N8030, N22031);
nand NAND2 (N22981, N22976, N14825);
nand NAND4 (N22982, N22978, N10177, N9643, N9382);
buf BUF1 (N22983, N22982);
nand NAND3 (N22984, N22955, N850, N6140);
nand NAND4 (N22985, N22983, N20017, N1902, N9295);
or OR4 (N22986, N22964, N10942, N19061, N19891);
buf BUF1 (N22987, N22980);
nand NAND3 (N22988, N22971, N4419, N12944);
buf BUF1 (N22989, N22979);
and AND3 (N22990, N22988, N18010, N16943);
not NOT1 (N22991, N22986);
xor XOR2 (N22992, N22985, N22452);
nor NOR3 (N22993, N22989, N19300, N9123);
buf BUF1 (N22994, N22987);
or OR4 (N22995, N22939, N1553, N11159, N14259);
or OR4 (N22996, N22973, N15235, N8817, N13030);
nand NAND2 (N22997, N22981, N11907);
xor XOR2 (N22998, N22997, N200);
nand NAND4 (N22999, N22994, N2829, N4805, N21865);
and AND4 (N23000, N22995, N17997, N14306, N18901);
and AND2 (N23001, N22984, N11377);
not NOT1 (N23002, N22990);
and AND4 (N23003, N22993, N416, N12429, N322);
xor XOR2 (N23004, N22998, N10397);
xor XOR2 (N23005, N22970, N10070);
nand NAND2 (N23006, N22999, N538);
nand NAND3 (N23007, N22992, N19461, N20340);
buf BUF1 (N23008, N23000);
buf BUF1 (N23009, N22996);
and AND4 (N23010, N23007, N17709, N12879, N10724);
buf BUF1 (N23011, N23008);
and AND3 (N23012, N23004, N19774, N22433);
nand NAND3 (N23013, N22991, N14769, N8774);
nor NOR2 (N23014, N23003, N12848);
xor XOR2 (N23015, N23014, N19598);
buf BUF1 (N23016, N23013);
or OR2 (N23017, N23006, N15947);
or OR3 (N23018, N23010, N14187, N15962);
not NOT1 (N23019, N23015);
nor NOR4 (N23020, N23005, N5168, N18336, N20390);
or OR3 (N23021, N23012, N11351, N10523);
nor NOR4 (N23022, N23019, N7554, N22357, N6547);
not NOT1 (N23023, N23009);
nand NAND2 (N23024, N23018, N7260);
nor NOR2 (N23025, N23001, N13160);
nand NAND3 (N23026, N23017, N8661, N14972);
not NOT1 (N23027, N23023);
not NOT1 (N23028, N23024);
nor NOR2 (N23029, N23016, N9187);
or OR4 (N23030, N23025, N16260, N17855, N17282);
nor NOR3 (N23031, N23030, N15638, N9810);
nor NOR3 (N23032, N23027, N21969, N9606);
nand NAND3 (N23033, N23029, N10669, N14553);
nor NOR3 (N23034, N23031, N10765, N11368);
and AND3 (N23035, N23028, N19251, N10283);
and AND2 (N23036, N23035, N12814);
nor NOR3 (N23037, N23022, N11661, N21450);
not NOT1 (N23038, N23021);
buf BUF1 (N23039, N23034);
xor XOR2 (N23040, N23033, N12349);
nor NOR2 (N23041, N23039, N387);
and AND3 (N23042, N23020, N17593, N12209);
nand NAND4 (N23043, N23041, N16410, N8389, N19053);
buf BUF1 (N23044, N23026);
and AND3 (N23045, N23043, N21288, N11431);
and AND3 (N23046, N23032, N8107, N18457);
not NOT1 (N23047, N23038);
nand NAND4 (N23048, N23037, N17408, N17840, N10633);
buf BUF1 (N23049, N23045);
nand NAND3 (N23050, N23040, N8053, N18395);
or OR3 (N23051, N23047, N2566, N19308);
or OR4 (N23052, N23042, N16273, N22531, N20093);
xor XOR2 (N23053, N23049, N9348);
nand NAND4 (N23054, N23053, N15070, N22368, N22096);
and AND3 (N23055, N23052, N14480, N22058);
or OR3 (N23056, N23048, N16604, N16527);
nor NOR3 (N23057, N23055, N20683, N19603);
xor XOR2 (N23058, N23051, N3857);
not NOT1 (N23059, N23050);
not NOT1 (N23060, N23059);
not NOT1 (N23061, N23046);
buf BUF1 (N23062, N23054);
nor NOR4 (N23063, N23036, N7279, N12434, N14557);
nand NAND2 (N23064, N23056, N21993);
not NOT1 (N23065, N23057);
not NOT1 (N23066, N23064);
nor NOR4 (N23067, N23065, N3072, N22899, N14155);
not NOT1 (N23068, N23058);
xor XOR2 (N23069, N23066, N6008);
and AND4 (N23070, N23063, N7579, N10352, N18280);
not NOT1 (N23071, N23062);
or OR2 (N23072, N23068, N1106);
nand NAND3 (N23073, N23061, N22801, N14815);
buf BUF1 (N23074, N23002);
nor NOR2 (N23075, N23071, N17275);
nor NOR3 (N23076, N23070, N3474, N3631);
buf BUF1 (N23077, N23011);
buf BUF1 (N23078, N23076);
nor NOR3 (N23079, N23077, N11952, N22628);
and AND3 (N23080, N23067, N18527, N9097);
not NOT1 (N23081, N23078);
not NOT1 (N23082, N23075);
not NOT1 (N23083, N23073);
nor NOR2 (N23084, N23079, N2069);
not NOT1 (N23085, N23082);
or OR4 (N23086, N23081, N2106, N15399, N15724);
xor XOR2 (N23087, N23060, N20384);
xor XOR2 (N23088, N23087, N9127);
nor NOR3 (N23089, N23072, N5922, N8926);
buf BUF1 (N23090, N23083);
buf BUF1 (N23091, N23090);
and AND3 (N23092, N23084, N7656, N15676);
and AND2 (N23093, N23086, N1180);
and AND4 (N23094, N23089, N11289, N5008, N21240);
xor XOR2 (N23095, N23093, N5845);
and AND3 (N23096, N23094, N18268, N4258);
buf BUF1 (N23097, N23092);
nand NAND4 (N23098, N23088, N6874, N18290, N19163);
nor NOR3 (N23099, N23097, N18652, N4941);
xor XOR2 (N23100, N23080, N14315);
and AND2 (N23101, N23096, N22727);
not NOT1 (N23102, N23085);
not NOT1 (N23103, N23074);
nor NOR3 (N23104, N23100, N1287, N674);
not NOT1 (N23105, N23101);
buf BUF1 (N23106, N23105);
nand NAND4 (N23107, N23104, N10569, N4164, N7643);
and AND3 (N23108, N23091, N443, N15343);
or OR4 (N23109, N23044, N17291, N13005, N16925);
nor NOR2 (N23110, N23108, N21797);
nor NOR4 (N23111, N23110, N12951, N4208, N2387);
nor NOR4 (N23112, N23111, N4171, N2432, N11269);
not NOT1 (N23113, N23112);
and AND4 (N23114, N23109, N9604, N9929, N20316);
not NOT1 (N23115, N23106);
xor XOR2 (N23116, N23102, N2000);
not NOT1 (N23117, N23113);
buf BUF1 (N23118, N23103);
or OR2 (N23119, N23098, N19896);
and AND2 (N23120, N23095, N1116);
or OR2 (N23121, N23117, N21851);
xor XOR2 (N23122, N23119, N20053);
xor XOR2 (N23123, N23118, N13912);
xor XOR2 (N23124, N23116, N7488);
nand NAND4 (N23125, N23115, N5139, N13660, N6823);
not NOT1 (N23126, N23069);
buf BUF1 (N23127, N23114);
and AND4 (N23128, N23123, N6613, N14727, N4574);
buf BUF1 (N23129, N23099);
not NOT1 (N23130, N23122);
nor NOR3 (N23131, N23129, N19981, N2898);
nor NOR4 (N23132, N23131, N7647, N16914, N258);
and AND2 (N23133, N23124, N6814);
nand NAND2 (N23134, N23126, N20706);
nand NAND2 (N23135, N23127, N19620);
buf BUF1 (N23136, N23134);
or OR2 (N23137, N23132, N15663);
buf BUF1 (N23138, N23137);
xor XOR2 (N23139, N23120, N13909);
not NOT1 (N23140, N23138);
or OR2 (N23141, N23107, N4877);
not NOT1 (N23142, N23133);
nand NAND3 (N23143, N23130, N497, N18202);
buf BUF1 (N23144, N23136);
xor XOR2 (N23145, N23139, N2146);
nor NOR3 (N23146, N23128, N2160, N12555);
nand NAND2 (N23147, N23143, N16508);
nor NOR2 (N23148, N23146, N1662);
or OR2 (N23149, N23145, N13205);
xor XOR2 (N23150, N23144, N7720);
buf BUF1 (N23151, N23135);
xor XOR2 (N23152, N23151, N5388);
buf BUF1 (N23153, N23140);
nand NAND2 (N23154, N23153, N20009);
buf BUF1 (N23155, N23141);
buf BUF1 (N23156, N23154);
buf BUF1 (N23157, N23147);
not NOT1 (N23158, N23150);
nor NOR4 (N23159, N23157, N17508, N21368, N8499);
nor NOR2 (N23160, N23155, N20712);
xor XOR2 (N23161, N23159, N8834);
nor NOR2 (N23162, N23152, N12164);
nand NAND4 (N23163, N23161, N12303, N1779, N7856);
nand NAND3 (N23164, N23125, N1915, N8457);
not NOT1 (N23165, N23149);
not NOT1 (N23166, N23156);
and AND3 (N23167, N23166, N2176, N13557);
nor NOR2 (N23168, N23165, N18853);
buf BUF1 (N23169, N23121);
or OR3 (N23170, N23164, N16009, N21374);
not NOT1 (N23171, N23169);
xor XOR2 (N23172, N23142, N16787);
buf BUF1 (N23173, N23171);
nand NAND4 (N23174, N23158, N10161, N13837, N11736);
nand NAND3 (N23175, N23162, N17381, N20743);
xor XOR2 (N23176, N23167, N5946);
nand NAND3 (N23177, N23170, N20360, N13992);
xor XOR2 (N23178, N23173, N14162);
nor NOR3 (N23179, N23168, N7410, N22373);
nor NOR3 (N23180, N23174, N6551, N7929);
or OR3 (N23181, N23179, N22473, N2724);
or OR4 (N23182, N23176, N14212, N8707, N8489);
buf BUF1 (N23183, N23175);
xor XOR2 (N23184, N23163, N19065);
xor XOR2 (N23185, N23180, N10433);
buf BUF1 (N23186, N23183);
buf BUF1 (N23187, N23178);
and AND2 (N23188, N23181, N22802);
xor XOR2 (N23189, N23172, N12618);
nor NOR4 (N23190, N23186, N11543, N5879, N4551);
and AND3 (N23191, N23184, N23139, N17618);
nand NAND4 (N23192, N23182, N18397, N13477, N22009);
buf BUF1 (N23193, N23177);
or OR2 (N23194, N23193, N12800);
nor NOR4 (N23195, N23192, N9279, N7324, N6535);
buf BUF1 (N23196, N23189);
or OR3 (N23197, N23160, N15378, N4719);
and AND3 (N23198, N23187, N8113, N12172);
and AND3 (N23199, N23190, N15827, N19342);
nand NAND4 (N23200, N23198, N22311, N3258, N20531);
nor NOR2 (N23201, N23191, N10448);
and AND3 (N23202, N23200, N268, N9102);
or OR4 (N23203, N23188, N21491, N1889, N22340);
and AND3 (N23204, N23202, N18870, N13627);
buf BUF1 (N23205, N23148);
buf BUF1 (N23206, N23199);
and AND4 (N23207, N23185, N2313, N1886, N18887);
and AND2 (N23208, N23206, N20221);
nand NAND3 (N23209, N23197, N18106, N3333);
buf BUF1 (N23210, N23208);
or OR3 (N23211, N23207, N4643, N17867);
or OR2 (N23212, N23196, N17697);
nand NAND2 (N23213, N23201, N20406);
xor XOR2 (N23214, N23213, N13945);
and AND3 (N23215, N23214, N9958, N17982);
not NOT1 (N23216, N23212);
xor XOR2 (N23217, N23210, N21592);
xor XOR2 (N23218, N23194, N12010);
and AND4 (N23219, N23204, N3216, N7195, N7198);
xor XOR2 (N23220, N23215, N4192);
buf BUF1 (N23221, N23218);
not NOT1 (N23222, N23219);
xor XOR2 (N23223, N23217, N8531);
xor XOR2 (N23224, N23220, N14833);
nand NAND3 (N23225, N23209, N21567, N17869);
not NOT1 (N23226, N23216);
nand NAND3 (N23227, N23203, N10180, N7605);
nand NAND3 (N23228, N23195, N4219, N11157);
or OR2 (N23229, N23226, N14155);
buf BUF1 (N23230, N23225);
and AND4 (N23231, N23222, N8173, N10540, N7160);
xor XOR2 (N23232, N23231, N11746);
xor XOR2 (N23233, N23205, N22768);
nand NAND3 (N23234, N23211, N21142, N8154);
or OR2 (N23235, N23221, N16511);
not NOT1 (N23236, N23230);
xor XOR2 (N23237, N23232, N14550);
nor NOR3 (N23238, N23233, N13831, N16404);
not NOT1 (N23239, N23238);
xor XOR2 (N23240, N23228, N13723);
xor XOR2 (N23241, N23227, N7239);
xor XOR2 (N23242, N23237, N11786);
nor NOR3 (N23243, N23242, N11789, N16550);
nor NOR3 (N23244, N23243, N19876, N15394);
and AND3 (N23245, N23224, N4368, N11899);
not NOT1 (N23246, N23240);
and AND4 (N23247, N23246, N6342, N18596, N10794);
and AND2 (N23248, N23239, N16390);
nand NAND2 (N23249, N23244, N21771);
nand NAND3 (N23250, N23236, N7901, N1118);
nand NAND4 (N23251, N23235, N3131, N16312, N17053);
nor NOR2 (N23252, N23229, N1274);
xor XOR2 (N23253, N23234, N14457);
buf BUF1 (N23254, N23252);
xor XOR2 (N23255, N23251, N9906);
buf BUF1 (N23256, N23250);
not NOT1 (N23257, N23247);
nand NAND4 (N23258, N23223, N21627, N13758, N4307);
buf BUF1 (N23259, N23245);
and AND4 (N23260, N23241, N11778, N10557, N3143);
xor XOR2 (N23261, N23255, N20624);
not NOT1 (N23262, N23261);
or OR3 (N23263, N23254, N1902, N9982);
nor NOR2 (N23264, N23257, N22912);
and AND2 (N23265, N23264, N17699);
xor XOR2 (N23266, N23262, N7681);
xor XOR2 (N23267, N23265, N13155);
or OR4 (N23268, N23263, N13459, N7116, N11420);
not NOT1 (N23269, N23267);
nand NAND2 (N23270, N23249, N21711);
nor NOR3 (N23271, N23256, N4943, N13418);
buf BUF1 (N23272, N23266);
not NOT1 (N23273, N23258);
nor NOR4 (N23274, N23260, N6502, N20453, N22226);
and AND3 (N23275, N23268, N20700, N19540);
nand NAND2 (N23276, N23274, N21833);
and AND2 (N23277, N23272, N21984);
not NOT1 (N23278, N23275);
and AND4 (N23279, N23248, N7503, N21118, N8146);
nand NAND2 (N23280, N23259, N23044);
buf BUF1 (N23281, N23270);
nand NAND3 (N23282, N23281, N14664, N21944);
nor NOR4 (N23283, N23271, N6309, N5049, N2477);
nor NOR2 (N23284, N23277, N12700);
or OR4 (N23285, N23276, N15232, N23041, N14639);
xor XOR2 (N23286, N23282, N1862);
buf BUF1 (N23287, N23273);
nand NAND4 (N23288, N23286, N1716, N10511, N1827);
nor NOR3 (N23289, N23283, N12318, N22513);
buf BUF1 (N23290, N23278);
not NOT1 (N23291, N23287);
or OR2 (N23292, N23280, N19627);
nand NAND2 (N23293, N23284, N9972);
and AND2 (N23294, N23288, N2880);
xor XOR2 (N23295, N23279, N22689);
xor XOR2 (N23296, N23290, N5753);
or OR3 (N23297, N23293, N3002, N16097);
nand NAND2 (N23298, N23294, N3844);
or OR4 (N23299, N23269, N4222, N7120, N1599);
nand NAND3 (N23300, N23295, N16785, N699);
not NOT1 (N23301, N23285);
and AND4 (N23302, N23298, N16026, N5023, N8671);
buf BUF1 (N23303, N23301);
or OR2 (N23304, N23253, N19402);
xor XOR2 (N23305, N23291, N3739);
xor XOR2 (N23306, N23297, N11180);
buf BUF1 (N23307, N23300);
nor NOR4 (N23308, N23296, N21435, N15665, N3939);
nor NOR3 (N23309, N23306, N13916, N22850);
xor XOR2 (N23310, N23299, N3918);
nor NOR4 (N23311, N23289, N21580, N14881, N13069);
or OR3 (N23312, N23302, N8334, N4784);
xor XOR2 (N23313, N23307, N7486);
not NOT1 (N23314, N23303);
or OR3 (N23315, N23312, N13798, N3122);
xor XOR2 (N23316, N23311, N19130);
and AND3 (N23317, N23315, N9198, N17829);
or OR2 (N23318, N23304, N1287);
nand NAND4 (N23319, N23309, N10281, N6150, N4801);
nand NAND4 (N23320, N23318, N7528, N22020, N14231);
nand NAND2 (N23321, N23305, N5955);
not NOT1 (N23322, N23314);
or OR4 (N23323, N23319, N11458, N14569, N12290);
nor NOR3 (N23324, N23322, N17665, N7310);
buf BUF1 (N23325, N23292);
nand NAND2 (N23326, N23321, N14991);
buf BUF1 (N23327, N23326);
xor XOR2 (N23328, N23323, N18639);
buf BUF1 (N23329, N23327);
xor XOR2 (N23330, N23320, N14439);
buf BUF1 (N23331, N23330);
nor NOR4 (N23332, N23325, N10242, N17227, N7737);
buf BUF1 (N23333, N23329);
and AND2 (N23334, N23331, N12166);
nand NAND2 (N23335, N23333, N388);
nor NOR3 (N23336, N23332, N1932, N16131);
nand NAND3 (N23337, N23316, N12882, N11613);
not NOT1 (N23338, N23324);
not NOT1 (N23339, N23335);
nor NOR4 (N23340, N23310, N5982, N19546, N2211);
nand NAND4 (N23341, N23338, N13392, N9200, N8318);
nand NAND3 (N23342, N23336, N9927, N138);
buf BUF1 (N23343, N23341);
nand NAND2 (N23344, N23317, N17690);
or OR4 (N23345, N23340, N10887, N15017, N10517);
and AND4 (N23346, N23344, N18491, N17394, N5423);
and AND2 (N23347, N23339, N9647);
or OR3 (N23348, N23347, N21757, N13950);
nor NOR2 (N23349, N23346, N12215);
not NOT1 (N23350, N23343);
xor XOR2 (N23351, N23349, N9842);
not NOT1 (N23352, N23350);
or OR2 (N23353, N23313, N12427);
nand NAND2 (N23354, N23342, N14444);
not NOT1 (N23355, N23348);
xor XOR2 (N23356, N23345, N1113);
or OR4 (N23357, N23356, N11688, N22039, N16414);
nor NOR4 (N23358, N23308, N10065, N23124, N22747);
or OR4 (N23359, N23355, N18321, N19089, N6554);
nor NOR4 (N23360, N23351, N9708, N22146, N7309);
and AND3 (N23361, N23359, N2523, N15911);
nand NAND3 (N23362, N23352, N7157, N14401);
nand NAND3 (N23363, N23354, N6735, N818);
buf BUF1 (N23364, N23362);
xor XOR2 (N23365, N23353, N9859);
not NOT1 (N23366, N23365);
or OR2 (N23367, N23328, N256);
and AND3 (N23368, N23334, N12949, N12236);
or OR2 (N23369, N23363, N23066);
xor XOR2 (N23370, N23366, N22464);
xor XOR2 (N23371, N23357, N15444);
buf BUF1 (N23372, N23360);
and AND3 (N23373, N23372, N5578, N6586);
nor NOR2 (N23374, N23358, N508);
nor NOR4 (N23375, N23337, N16909, N21491, N12716);
and AND3 (N23376, N23368, N17383, N1944);
nor NOR4 (N23377, N23374, N1514, N2730, N13754);
xor XOR2 (N23378, N23377, N15567);
xor XOR2 (N23379, N23361, N397);
nand NAND2 (N23380, N23369, N5499);
and AND2 (N23381, N23380, N4925);
or OR4 (N23382, N23375, N22492, N4892, N5437);
xor XOR2 (N23383, N23364, N4067);
not NOT1 (N23384, N23371);
nor NOR3 (N23385, N23384, N5251, N5346);
nor NOR2 (N23386, N23370, N2375);
nor NOR3 (N23387, N23367, N19168, N19383);
and AND2 (N23388, N23376, N8139);
not NOT1 (N23389, N23382);
and AND4 (N23390, N23379, N8420, N13726, N21794);
not NOT1 (N23391, N23383);
buf BUF1 (N23392, N23389);
buf BUF1 (N23393, N23373);
not NOT1 (N23394, N23393);
buf BUF1 (N23395, N23388);
nand NAND2 (N23396, N23387, N19566);
or OR2 (N23397, N23386, N19737);
buf BUF1 (N23398, N23390);
nand NAND4 (N23399, N23395, N20881, N17241, N15268);
nor NOR2 (N23400, N23381, N5218);
and AND3 (N23401, N23378, N11503, N21170);
nor NOR3 (N23402, N23398, N12803, N11166);
nand NAND2 (N23403, N23401, N4860);
buf BUF1 (N23404, N23394);
and AND4 (N23405, N23391, N6084, N18995, N9280);
xor XOR2 (N23406, N23402, N19063);
and AND3 (N23407, N23396, N9153, N19413);
not NOT1 (N23408, N23399);
and AND2 (N23409, N23404, N21397);
not NOT1 (N23410, N23392);
not NOT1 (N23411, N23400);
not NOT1 (N23412, N23409);
nor NOR2 (N23413, N23385, N418);
nand NAND4 (N23414, N23411, N12161, N17088, N17899);
xor XOR2 (N23415, N23410, N13562);
nor NOR3 (N23416, N23403, N10365, N12300);
nor NOR2 (N23417, N23415, N8970);
nand NAND3 (N23418, N23416, N10206, N13301);
xor XOR2 (N23419, N23414, N14874);
or OR3 (N23420, N23413, N23278, N17157);
not NOT1 (N23421, N23408);
nor NOR2 (N23422, N23418, N8769);
nor NOR2 (N23423, N23406, N272);
nor NOR2 (N23424, N23412, N2982);
nor NOR4 (N23425, N23422, N8635, N21194, N2667);
or OR2 (N23426, N23425, N5960);
and AND4 (N23427, N23417, N296, N8523, N7598);
and AND3 (N23428, N23407, N21029, N22783);
and AND3 (N23429, N23423, N18316, N15112);
nor NOR4 (N23430, N23419, N22324, N15932, N3684);
xor XOR2 (N23431, N23426, N17715);
or OR2 (N23432, N23427, N12382);
buf BUF1 (N23433, N23432);
nor NOR4 (N23434, N23420, N20270, N2387, N8883);
and AND3 (N23435, N23434, N1518, N20687);
nand NAND3 (N23436, N23430, N19922, N14935);
nor NOR4 (N23437, N23433, N1902, N19716, N12082);
xor XOR2 (N23438, N23435, N17219);
buf BUF1 (N23439, N23436);
nor NOR4 (N23440, N23405, N6129, N4232, N22766);
and AND2 (N23441, N23421, N22249);
xor XOR2 (N23442, N23428, N19075);
not NOT1 (N23443, N23442);
buf BUF1 (N23444, N23397);
and AND4 (N23445, N23443, N16502, N19593, N10987);
and AND2 (N23446, N23440, N450);
or OR3 (N23447, N23439, N14631, N1120);
nor NOR4 (N23448, N23438, N12068, N2995, N21603);
nor NOR2 (N23449, N23445, N13877);
xor XOR2 (N23450, N23437, N7797);
nand NAND3 (N23451, N23441, N8726, N6665);
or OR4 (N23452, N23429, N11959, N15795, N22437);
nor NOR4 (N23453, N23448, N465, N682, N1653);
not NOT1 (N23454, N23446);
xor XOR2 (N23455, N23450, N3460);
nand NAND4 (N23456, N23453, N11112, N13361, N1017);
nor NOR3 (N23457, N23424, N15799, N10323);
buf BUF1 (N23458, N23444);
buf BUF1 (N23459, N23431);
nor NOR2 (N23460, N23457, N20232);
nand NAND4 (N23461, N23455, N6916, N8847, N10144);
nand NAND2 (N23462, N23458, N9908);
nand NAND4 (N23463, N23456, N8110, N5493, N2005);
nand NAND2 (N23464, N23460, N12967);
and AND4 (N23465, N23461, N9197, N3847, N18290);
buf BUF1 (N23466, N23451);
and AND2 (N23467, N23464, N803);
or OR4 (N23468, N23454, N4148, N17046, N21209);
nor NOR4 (N23469, N23465, N12759, N21444, N11432);
xor XOR2 (N23470, N23468, N22452);
nor NOR2 (N23471, N23449, N280);
and AND3 (N23472, N23466, N15379, N12422);
nand NAND4 (N23473, N23452, N7162, N5467, N17228);
and AND4 (N23474, N23472, N19606, N5995, N6572);
nand NAND3 (N23475, N23471, N21943, N19115);
nor NOR3 (N23476, N23467, N4602, N3165);
xor XOR2 (N23477, N23469, N2903);
and AND2 (N23478, N23447, N5708);
nand NAND2 (N23479, N23474, N18701);
or OR2 (N23480, N23473, N17411);
nand NAND2 (N23481, N23480, N6435);
and AND2 (N23482, N23475, N6751);
xor XOR2 (N23483, N23482, N20251);
buf BUF1 (N23484, N23481);
nor NOR4 (N23485, N23462, N20233, N5923, N7418);
nand NAND4 (N23486, N23463, N21780, N20911, N21864);
xor XOR2 (N23487, N23477, N22089);
buf BUF1 (N23488, N23486);
nor NOR3 (N23489, N23479, N7339, N12126);
xor XOR2 (N23490, N23489, N18004);
or OR2 (N23491, N23478, N21987);
or OR4 (N23492, N23483, N848, N12254, N23412);
nand NAND2 (N23493, N23470, N6166);
buf BUF1 (N23494, N23487);
or OR3 (N23495, N23485, N19616, N14029);
xor XOR2 (N23496, N23476, N15242);
and AND2 (N23497, N23494, N18208);
buf BUF1 (N23498, N23493);
xor XOR2 (N23499, N23495, N7897);
or OR2 (N23500, N23497, N14309);
or OR4 (N23501, N23498, N9804, N6264, N11344);
xor XOR2 (N23502, N23492, N8978);
and AND4 (N23503, N23500, N9360, N5771, N7946);
nor NOR2 (N23504, N23491, N15814);
not NOT1 (N23505, N23490);
xor XOR2 (N23506, N23499, N2403);
not NOT1 (N23507, N23503);
not NOT1 (N23508, N23507);
and AND3 (N23509, N23488, N9282, N2110);
nand NAND2 (N23510, N23459, N6627);
and AND4 (N23511, N23501, N4733, N16214, N21011);
and AND4 (N23512, N23504, N11386, N21504, N14094);
not NOT1 (N23513, N23511);
xor XOR2 (N23514, N23508, N3577);
xor XOR2 (N23515, N23509, N5504);
nor NOR4 (N23516, N23505, N21390, N18808, N16603);
buf BUF1 (N23517, N23513);
or OR2 (N23518, N23512, N2699);
nand NAND2 (N23519, N23484, N16995);
nand NAND2 (N23520, N23510, N10614);
and AND4 (N23521, N23516, N13170, N11631, N1215);
buf BUF1 (N23522, N23496);
nor NOR2 (N23523, N23506, N1842);
buf BUF1 (N23524, N23520);
nand NAND4 (N23525, N23517, N15930, N5919, N15935);
nor NOR4 (N23526, N23502, N21883, N19767, N2322);
and AND2 (N23527, N23526, N13990);
xor XOR2 (N23528, N23523, N12949);
not NOT1 (N23529, N23521);
or OR3 (N23530, N23515, N13784, N600);
nand NAND2 (N23531, N23524, N5747);
xor XOR2 (N23532, N23525, N2989);
and AND4 (N23533, N23518, N6830, N23222, N12110);
buf BUF1 (N23534, N23527);
nor NOR2 (N23535, N23522, N4490);
not NOT1 (N23536, N23528);
buf BUF1 (N23537, N23519);
not NOT1 (N23538, N23534);
nor NOR3 (N23539, N23538, N14427, N23017);
nor NOR2 (N23540, N23529, N11249);
nand NAND4 (N23541, N23536, N6997, N19533, N1685);
and AND2 (N23542, N23532, N2955);
nor NOR4 (N23543, N23530, N22003, N11617, N11967);
buf BUF1 (N23544, N23543);
or OR3 (N23545, N23540, N19650, N11360);
nand NAND3 (N23546, N23545, N6107, N20423);
nor NOR3 (N23547, N23539, N17406, N14779);
xor XOR2 (N23548, N23544, N1880);
or OR3 (N23549, N23541, N12602, N1629);
nor NOR2 (N23550, N23535, N14166);
xor XOR2 (N23551, N23548, N20517);
xor XOR2 (N23552, N23537, N7191);
nand NAND3 (N23553, N23550, N8299, N16918);
or OR3 (N23554, N23549, N16735, N20978);
and AND3 (N23555, N23542, N22204, N511);
nand NAND4 (N23556, N23555, N18141, N5287, N7858);
nand NAND2 (N23557, N23554, N10495);
or OR2 (N23558, N23546, N17653);
nor NOR2 (N23559, N23557, N6428);
and AND4 (N23560, N23553, N17572, N11345, N9989);
xor XOR2 (N23561, N23552, N20059);
xor XOR2 (N23562, N23531, N20167);
and AND4 (N23563, N23562, N19280, N6976, N1860);
buf BUF1 (N23564, N23561);
not NOT1 (N23565, N23560);
nand NAND3 (N23566, N23558, N5867, N20826);
not NOT1 (N23567, N23533);
xor XOR2 (N23568, N23564, N12165);
or OR3 (N23569, N23547, N4993, N4602);
not NOT1 (N23570, N23565);
xor XOR2 (N23571, N23559, N363);
nor NOR2 (N23572, N23570, N20596);
buf BUF1 (N23573, N23571);
xor XOR2 (N23574, N23573, N2090);
not NOT1 (N23575, N23566);
xor XOR2 (N23576, N23514, N890);
nand NAND2 (N23577, N23569, N11235);
nor NOR3 (N23578, N23567, N3858, N8967);
nor NOR2 (N23579, N23575, N1843);
buf BUF1 (N23580, N23578);
nand NAND4 (N23581, N23572, N17065, N5981, N22913);
and AND3 (N23582, N23574, N13488, N1935);
nand NAND3 (N23583, N23563, N4244, N6636);
and AND2 (N23584, N23576, N7991);
nand NAND2 (N23585, N23583, N18523);
nor NOR3 (N23586, N23585, N8570, N9813);
buf BUF1 (N23587, N23580);
nand NAND2 (N23588, N23581, N7858);
nor NOR4 (N23589, N23556, N4460, N12875, N1805);
not NOT1 (N23590, N23587);
nor NOR4 (N23591, N23589, N19884, N10523, N15546);
not NOT1 (N23592, N23590);
nand NAND4 (N23593, N23582, N10961, N13057, N21689);
and AND3 (N23594, N23588, N15438, N16442);
xor XOR2 (N23595, N23594, N590);
nand NAND3 (N23596, N23579, N16253, N13272);
and AND2 (N23597, N23551, N13835);
buf BUF1 (N23598, N23568);
and AND2 (N23599, N23577, N14725);
or OR4 (N23600, N23593, N999, N12729, N15496);
xor XOR2 (N23601, N23595, N23077);
nor NOR4 (N23602, N23586, N17040, N21713, N14692);
nor NOR3 (N23603, N23597, N701, N11450);
or OR3 (N23604, N23598, N15287, N14570);
not NOT1 (N23605, N23584);
buf BUF1 (N23606, N23605);
and AND4 (N23607, N23596, N12158, N11091, N22675);
xor XOR2 (N23608, N23600, N642);
xor XOR2 (N23609, N23607, N21464);
nand NAND2 (N23610, N23606, N6632);
nand NAND2 (N23611, N23601, N2094);
buf BUF1 (N23612, N23608);
not NOT1 (N23613, N23591);
not NOT1 (N23614, N23612);
nand NAND2 (N23615, N23592, N16710);
not NOT1 (N23616, N23610);
not NOT1 (N23617, N23599);
and AND4 (N23618, N23603, N19690, N631, N11145);
nor NOR2 (N23619, N23617, N19113);
xor XOR2 (N23620, N23602, N7324);
nor NOR2 (N23621, N23619, N96);
xor XOR2 (N23622, N23609, N8492);
not NOT1 (N23623, N23604);
nor NOR3 (N23624, N23618, N9615, N1578);
buf BUF1 (N23625, N23622);
or OR4 (N23626, N23620, N920, N10205, N2860);
xor XOR2 (N23627, N23625, N17772);
buf BUF1 (N23628, N23621);
xor XOR2 (N23629, N23628, N18487);
and AND4 (N23630, N23624, N10192, N6489, N3859);
or OR4 (N23631, N23613, N15007, N14781, N14322);
nor NOR4 (N23632, N23611, N20169, N5385, N4703);
xor XOR2 (N23633, N23616, N2476);
not NOT1 (N23634, N23614);
or OR4 (N23635, N23623, N3520, N6280, N8254);
buf BUF1 (N23636, N23634);
and AND2 (N23637, N23632, N6216);
xor XOR2 (N23638, N23636, N4363);
or OR3 (N23639, N23635, N23323, N1310);
nor NOR3 (N23640, N23639, N7523, N13498);
xor XOR2 (N23641, N23631, N15646);
and AND4 (N23642, N23630, N14108, N10889, N5692);
nand NAND2 (N23643, N23641, N1903);
not NOT1 (N23644, N23640);
xor XOR2 (N23645, N23642, N11828);
xor XOR2 (N23646, N23637, N3466);
buf BUF1 (N23647, N23633);
nor NOR3 (N23648, N23638, N6670, N5686);
nor NOR4 (N23649, N23615, N656, N21418, N9235);
or OR2 (N23650, N23649, N4716);
and AND3 (N23651, N23643, N4667, N10142);
buf BUF1 (N23652, N23645);
not NOT1 (N23653, N23644);
not NOT1 (N23654, N23653);
xor XOR2 (N23655, N23650, N16875);
or OR2 (N23656, N23627, N10669);
xor XOR2 (N23657, N23652, N19032);
nand NAND2 (N23658, N23654, N13937);
or OR3 (N23659, N23646, N4219, N3650);
not NOT1 (N23660, N23629);
nand NAND4 (N23661, N23651, N9792, N370, N18068);
and AND2 (N23662, N23647, N716);
buf BUF1 (N23663, N23656);
nor NOR3 (N23664, N23658, N16024, N4970);
buf BUF1 (N23665, N23659);
buf BUF1 (N23666, N23662);
xor XOR2 (N23667, N23657, N3298);
not NOT1 (N23668, N23661);
and AND2 (N23669, N23648, N11357);
xor XOR2 (N23670, N23665, N30);
and AND3 (N23671, N23666, N18549, N15600);
not NOT1 (N23672, N23670);
nand NAND2 (N23673, N23660, N12241);
xor XOR2 (N23674, N23672, N2602);
nand NAND3 (N23675, N23673, N22165, N10337);
nand NAND3 (N23676, N23669, N5394, N20629);
nand NAND3 (N23677, N23668, N20573, N18462);
or OR2 (N23678, N23676, N3382);
and AND2 (N23679, N23667, N23248);
nand NAND2 (N23680, N23674, N2056);
buf BUF1 (N23681, N23671);
buf BUF1 (N23682, N23663);
xor XOR2 (N23683, N23682, N3036);
and AND2 (N23684, N23678, N20665);
not NOT1 (N23685, N23680);
not NOT1 (N23686, N23681);
nand NAND3 (N23687, N23675, N20743, N13775);
not NOT1 (N23688, N23677);
not NOT1 (N23689, N23687);
buf BUF1 (N23690, N23688);
xor XOR2 (N23691, N23664, N15308);
or OR2 (N23692, N23691, N13003);
and AND2 (N23693, N23690, N23401);
or OR4 (N23694, N23686, N23547, N1648, N9997);
buf BUF1 (N23695, N23679);
or OR2 (N23696, N23689, N11084);
or OR4 (N23697, N23655, N21113, N20697, N5434);
or OR4 (N23698, N23697, N10855, N21353, N8509);
nor NOR3 (N23699, N23698, N1109, N16661);
and AND4 (N23700, N23683, N13026, N22548, N18649);
nand NAND3 (N23701, N23626, N14634, N153);
and AND2 (N23702, N23684, N3821);
buf BUF1 (N23703, N23693);
nor NOR2 (N23704, N23695, N5815);
nand NAND4 (N23705, N23703, N13871, N2981, N16478);
not NOT1 (N23706, N23702);
not NOT1 (N23707, N23705);
nor NOR3 (N23708, N23694, N16284, N18716);
xor XOR2 (N23709, N23692, N15167);
and AND4 (N23710, N23701, N3045, N13131, N16913);
nand NAND3 (N23711, N23704, N21779, N21932);
and AND3 (N23712, N23708, N11009, N18067);
buf BUF1 (N23713, N23685);
buf BUF1 (N23714, N23699);
xor XOR2 (N23715, N23700, N21817);
and AND2 (N23716, N23696, N1312);
nor NOR3 (N23717, N23706, N5140, N5327);
and AND3 (N23718, N23711, N6088, N12326);
not NOT1 (N23719, N23717);
not NOT1 (N23720, N23712);
nand NAND2 (N23721, N23719, N4696);
and AND4 (N23722, N23713, N3049, N3182, N19818);
and AND3 (N23723, N23718, N4324, N3264);
xor XOR2 (N23724, N23721, N16213);
xor XOR2 (N23725, N23723, N5280);
and AND3 (N23726, N23710, N22087, N12715);
not NOT1 (N23727, N23725);
or OR2 (N23728, N23707, N5263);
nor NOR2 (N23729, N23727, N9444);
nor NOR3 (N23730, N23726, N5088, N1573);
buf BUF1 (N23731, N23722);
and AND4 (N23732, N23730, N21942, N22086, N23009);
nand NAND2 (N23733, N23729, N2289);
nor NOR2 (N23734, N23716, N17396);
xor XOR2 (N23735, N23731, N3442);
and AND3 (N23736, N23720, N19476, N6329);
nand NAND2 (N23737, N23735, N17504);
and AND2 (N23738, N23734, N11213);
xor XOR2 (N23739, N23724, N12527);
buf BUF1 (N23740, N23714);
not NOT1 (N23741, N23732);
not NOT1 (N23742, N23715);
nor NOR2 (N23743, N23739, N2311);
nor NOR3 (N23744, N23733, N23220, N2839);
nor NOR3 (N23745, N23740, N11813, N18863);
xor XOR2 (N23746, N23745, N1081);
nor NOR2 (N23747, N23743, N17016);
xor XOR2 (N23748, N23737, N5178);
xor XOR2 (N23749, N23736, N19625);
nor NOR4 (N23750, N23741, N2166, N13484, N19307);
nand NAND3 (N23751, N23709, N12026, N2594);
buf BUF1 (N23752, N23728);
nor NOR4 (N23753, N23747, N16093, N19224, N3734);
buf BUF1 (N23754, N23750);
or OR3 (N23755, N23744, N7550, N19728);
nor NOR3 (N23756, N23751, N11998, N3632);
buf BUF1 (N23757, N23754);
buf BUF1 (N23758, N23749);
not NOT1 (N23759, N23757);
or OR3 (N23760, N23753, N9772, N12443);
or OR4 (N23761, N23755, N9658, N18161, N16886);
and AND4 (N23762, N23746, N19185, N8705, N9365);
and AND4 (N23763, N23759, N8134, N6735, N15098);
not NOT1 (N23764, N23760);
xor XOR2 (N23765, N23748, N2521);
not NOT1 (N23766, N23752);
or OR4 (N23767, N23765, N8007, N2191, N7362);
and AND3 (N23768, N23763, N16689, N23616);
and AND4 (N23769, N23766, N19926, N9882, N17536);
buf BUF1 (N23770, N23738);
nand NAND2 (N23771, N23767, N11200);
nor NOR3 (N23772, N23771, N9759, N2385);
nand NAND2 (N23773, N23758, N5042);
or OR4 (N23774, N23762, N20165, N17878, N7445);
not NOT1 (N23775, N23772);
nor NOR4 (N23776, N23742, N226, N9081, N6477);
or OR4 (N23777, N23768, N20963, N11357, N13036);
or OR3 (N23778, N23769, N10584, N1236);
and AND3 (N23779, N23776, N6481, N21598);
buf BUF1 (N23780, N23774);
xor XOR2 (N23781, N23778, N1443);
and AND4 (N23782, N23777, N14217, N16849, N2396);
buf BUF1 (N23783, N23761);
buf BUF1 (N23784, N23779);
buf BUF1 (N23785, N23781);
buf BUF1 (N23786, N23784);
not NOT1 (N23787, N23756);
xor XOR2 (N23788, N23785, N20601);
buf BUF1 (N23789, N23770);
buf BUF1 (N23790, N23782);
not NOT1 (N23791, N23764);
buf BUF1 (N23792, N23780);
nor NOR2 (N23793, N23787, N2980);
not NOT1 (N23794, N23791);
or OR3 (N23795, N23793, N21729, N831);
not NOT1 (N23796, N23790);
or OR3 (N23797, N23773, N20722, N21487);
xor XOR2 (N23798, N23792, N15986);
not NOT1 (N23799, N23798);
buf BUF1 (N23800, N23794);
buf BUF1 (N23801, N23789);
nor NOR2 (N23802, N23799, N5260);
not NOT1 (N23803, N23783);
nand NAND2 (N23804, N23797, N9119);
nor NOR3 (N23805, N23802, N3194, N16377);
nor NOR4 (N23806, N23796, N5520, N3626, N1640);
or OR4 (N23807, N23801, N6902, N7251, N10411);
or OR4 (N23808, N23786, N10293, N9622, N5716);
nor NOR4 (N23809, N23806, N4965, N19087, N21184);
and AND3 (N23810, N23809, N11462, N18265);
nor NOR2 (N23811, N23805, N10625);
nand NAND2 (N23812, N23788, N18718);
nand NAND3 (N23813, N23804, N17885, N9656);
nand NAND2 (N23814, N23807, N17522);
nor NOR2 (N23815, N23775, N3954);
nor NOR3 (N23816, N23812, N17346, N7934);
not NOT1 (N23817, N23795);
buf BUF1 (N23818, N23811);
or OR3 (N23819, N23803, N20720, N1709);
not NOT1 (N23820, N23815);
or OR2 (N23821, N23814, N341);
or OR2 (N23822, N23821, N7643);
nand NAND3 (N23823, N23822, N8401, N1791);
nand NAND3 (N23824, N23818, N4820, N6939);
buf BUF1 (N23825, N23813);
buf BUF1 (N23826, N23800);
nand NAND2 (N23827, N23817, N10046);
and AND4 (N23828, N23808, N14277, N3799, N1953);
xor XOR2 (N23829, N23828, N14923);
nor NOR4 (N23830, N23826, N11535, N847, N19099);
not NOT1 (N23831, N23829);
buf BUF1 (N23832, N23823);
and AND4 (N23833, N23830, N946, N7698, N22318);
and AND4 (N23834, N23810, N15289, N16277, N9583);
and AND2 (N23835, N23834, N4485);
buf BUF1 (N23836, N23833);
nor NOR2 (N23837, N23825, N23144);
nand NAND4 (N23838, N23824, N6010, N16080, N21537);
nor NOR2 (N23839, N23820, N5090);
and AND3 (N23840, N23831, N15731, N23);
and AND4 (N23841, N23832, N5651, N14977, N17691);
nor NOR4 (N23842, N23827, N2390, N18242, N11191);
or OR4 (N23843, N23842, N11969, N2101, N19269);
or OR2 (N23844, N23816, N12587);
and AND3 (N23845, N23819, N9343, N18790);
buf BUF1 (N23846, N23836);
xor XOR2 (N23847, N23845, N428);
xor XOR2 (N23848, N23843, N3956);
not NOT1 (N23849, N23837);
and AND4 (N23850, N23846, N19039, N6866, N7556);
nand NAND3 (N23851, N23847, N21818, N7387);
nor NOR2 (N23852, N23841, N21319);
and AND2 (N23853, N23839, N12091);
xor XOR2 (N23854, N23850, N8008);
nor NOR4 (N23855, N23840, N22999, N12704, N10585);
or OR4 (N23856, N23854, N11730, N22772, N14751);
and AND3 (N23857, N23844, N1383, N15544);
nand NAND2 (N23858, N23853, N22230);
xor XOR2 (N23859, N23855, N15473);
xor XOR2 (N23860, N23835, N23688);
xor XOR2 (N23861, N23857, N1377);
nand NAND2 (N23862, N23860, N10273);
not NOT1 (N23863, N23838);
and AND2 (N23864, N23859, N19584);
or OR3 (N23865, N23863, N6654, N4328);
xor XOR2 (N23866, N23851, N19605);
nor NOR4 (N23867, N23862, N18154, N2782, N21245);
nor NOR4 (N23868, N23858, N13566, N8560, N14207);
buf BUF1 (N23869, N23867);
not NOT1 (N23870, N23849);
buf BUF1 (N23871, N23852);
nand NAND4 (N23872, N23871, N12342, N22735, N21778);
and AND2 (N23873, N23861, N21800);
buf BUF1 (N23874, N23865);
and AND2 (N23875, N23873, N4870);
nand NAND4 (N23876, N23864, N12829, N12791, N2440);
nor NOR2 (N23877, N23869, N11614);
nor NOR2 (N23878, N23848, N19940);
and AND2 (N23879, N23877, N11116);
or OR4 (N23880, N23856, N5982, N16646, N17780);
not NOT1 (N23881, N23879);
nand NAND3 (N23882, N23868, N14048, N12556);
xor XOR2 (N23883, N23874, N3188);
and AND2 (N23884, N23875, N8433);
not NOT1 (N23885, N23870);
and AND4 (N23886, N23880, N6620, N18600, N17387);
buf BUF1 (N23887, N23884);
and AND4 (N23888, N23866, N17727, N18371, N9306);
nand NAND2 (N23889, N23885, N11631);
and AND4 (N23890, N23889, N1769, N10604, N20156);
buf BUF1 (N23891, N23876);
buf BUF1 (N23892, N23891);
and AND3 (N23893, N23881, N22793, N2608);
not NOT1 (N23894, N23893);
xor XOR2 (N23895, N23886, N18408);
nand NAND4 (N23896, N23872, N10414, N18299, N16453);
buf BUF1 (N23897, N23890);
or OR3 (N23898, N23882, N2281, N11315);
xor XOR2 (N23899, N23883, N13204);
buf BUF1 (N23900, N23888);
not NOT1 (N23901, N23892);
nor NOR3 (N23902, N23894, N8880, N19222);
or OR2 (N23903, N23896, N18383);
buf BUF1 (N23904, N23903);
nor NOR4 (N23905, N23898, N11668, N11779, N4020);
or OR3 (N23906, N23899, N17742, N6370);
nand NAND2 (N23907, N23878, N4226);
nor NOR2 (N23908, N23904, N11724);
or OR4 (N23909, N23900, N22045, N23057, N17517);
or OR2 (N23910, N23908, N17973);
nand NAND4 (N23911, N23895, N13811, N3758, N7776);
or OR2 (N23912, N23902, N15649);
buf BUF1 (N23913, N23911);
or OR3 (N23914, N23897, N11644, N20130);
xor XOR2 (N23915, N23906, N15815);
buf BUF1 (N23916, N23905);
buf BUF1 (N23917, N23912);
xor XOR2 (N23918, N23916, N16886);
and AND3 (N23919, N23901, N8986, N18062);
buf BUF1 (N23920, N23914);
not NOT1 (N23921, N23907);
buf BUF1 (N23922, N23921);
buf BUF1 (N23923, N23918);
nor NOR4 (N23924, N23923, N22282, N10241, N19003);
nand NAND4 (N23925, N23913, N1079, N8366, N18649);
not NOT1 (N23926, N23915);
buf BUF1 (N23927, N23924);
buf BUF1 (N23928, N23922);
buf BUF1 (N23929, N23928);
and AND4 (N23930, N23927, N15567, N16841, N18155);
nand NAND3 (N23931, N23926, N9079, N19954);
not NOT1 (N23932, N23930);
not NOT1 (N23933, N23919);
buf BUF1 (N23934, N23887);
and AND3 (N23935, N23931, N22695, N8809);
nor NOR2 (N23936, N23909, N1459);
nor NOR3 (N23937, N23936, N13151, N1119);
not NOT1 (N23938, N23920);
nor NOR3 (N23939, N23932, N5440, N13980);
nand NAND2 (N23940, N23935, N19876);
or OR2 (N23941, N23939, N18227);
and AND3 (N23942, N23917, N23198, N19960);
buf BUF1 (N23943, N23938);
or OR2 (N23944, N23925, N21532);
xor XOR2 (N23945, N23941, N22974);
nor NOR3 (N23946, N23944, N2026, N658);
nor NOR3 (N23947, N23910, N23876, N9043);
buf BUF1 (N23948, N23933);
not NOT1 (N23949, N23945);
xor XOR2 (N23950, N23943, N21157);
buf BUF1 (N23951, N23942);
not NOT1 (N23952, N23949);
nor NOR2 (N23953, N23951, N8566);
not NOT1 (N23954, N23929);
or OR4 (N23955, N23948, N5748, N12049, N3987);
or OR4 (N23956, N23955, N6645, N14607, N19063);
and AND3 (N23957, N23946, N12390, N23786);
nor NOR3 (N23958, N23952, N17749, N17718);
nor NOR3 (N23959, N23940, N2113, N15782);
nor NOR3 (N23960, N23937, N18875, N9932);
xor XOR2 (N23961, N23950, N11677);
and AND4 (N23962, N23959, N21617, N8407, N10179);
not NOT1 (N23963, N23954);
and AND4 (N23964, N23956, N7710, N437, N20603);
xor XOR2 (N23965, N23953, N19709);
not NOT1 (N23966, N23958);
xor XOR2 (N23967, N23962, N11909);
xor XOR2 (N23968, N23965, N21337);
nand NAND2 (N23969, N23963, N4537);
and AND2 (N23970, N23947, N13756);
xor XOR2 (N23971, N23967, N3427);
xor XOR2 (N23972, N23966, N14768);
and AND4 (N23973, N23960, N16614, N17029, N6277);
not NOT1 (N23974, N23934);
not NOT1 (N23975, N23974);
xor XOR2 (N23976, N23970, N8429);
nand NAND4 (N23977, N23976, N15523, N22220, N10638);
nor NOR2 (N23978, N23972, N1814);
and AND2 (N23979, N23964, N19976);
nor NOR4 (N23980, N23957, N19828, N3177, N706);
and AND2 (N23981, N23980, N11473);
or OR4 (N23982, N23981, N22755, N20441, N9229);
or OR3 (N23983, N23968, N15850, N13046);
or OR2 (N23984, N23977, N9762);
xor XOR2 (N23985, N23983, N10004);
nand NAND4 (N23986, N23979, N438, N16784, N3553);
buf BUF1 (N23987, N23971);
not NOT1 (N23988, N23986);
xor XOR2 (N23989, N23975, N21737);
nand NAND2 (N23990, N23988, N7337);
and AND2 (N23991, N23973, N8485);
and AND2 (N23992, N23987, N2765);
xor XOR2 (N23993, N23990, N15668);
nand NAND2 (N23994, N23982, N20499);
not NOT1 (N23995, N23985);
nor NOR3 (N23996, N23989, N8981, N14210);
xor XOR2 (N23997, N23992, N7721);
not NOT1 (N23998, N23984);
and AND3 (N23999, N23961, N11395, N22790);
nand NAND3 (N24000, N23995, N23385, N6120);
nand NAND3 (N24001, N23999, N22711, N7274);
nand NAND2 (N24002, N23997, N11360);
xor XOR2 (N24003, N24001, N15283);
and AND2 (N24004, N23991, N17189);
nand NAND4 (N24005, N24000, N19546, N16757, N10564);
buf BUF1 (N24006, N24005);
nand NAND3 (N24007, N23998, N12113, N21811);
not NOT1 (N24008, N23994);
nand NAND3 (N24009, N23996, N835, N19522);
nand NAND2 (N24010, N24009, N748);
buf BUF1 (N24011, N24007);
buf BUF1 (N24012, N24002);
xor XOR2 (N24013, N24006, N9596);
nor NOR3 (N24014, N24003, N21819, N17513);
xor XOR2 (N24015, N24004, N1134);
nor NOR2 (N24016, N24010, N6490);
buf BUF1 (N24017, N23978);
xor XOR2 (N24018, N24013, N15069);
not NOT1 (N24019, N23969);
or OR2 (N24020, N23993, N262);
not NOT1 (N24021, N24016);
nand NAND2 (N24022, N24017, N1259);
nand NAND3 (N24023, N24021, N19863, N12759);
and AND2 (N24024, N24018, N3113);
xor XOR2 (N24025, N24008, N7297);
or OR3 (N24026, N24024, N11139, N11956);
xor XOR2 (N24027, N24011, N19128);
nor NOR3 (N24028, N24015, N10126, N23547);
not NOT1 (N24029, N24023);
nand NAND3 (N24030, N24020, N1774, N14159);
or OR4 (N24031, N24022, N48, N3814, N10567);
nor NOR4 (N24032, N24019, N16940, N4234, N15829);
nor NOR2 (N24033, N24014, N16806);
and AND2 (N24034, N24032, N12948);
xor XOR2 (N24035, N24034, N950);
nor NOR4 (N24036, N24028, N2956, N11885, N23748);
not NOT1 (N24037, N24025);
or OR4 (N24038, N24033, N849, N8815, N17341);
buf BUF1 (N24039, N24031);
buf BUF1 (N24040, N24039);
nand NAND2 (N24041, N24035, N23239);
nand NAND3 (N24042, N24038, N12127, N4913);
nand NAND2 (N24043, N24036, N7954);
or OR4 (N24044, N24026, N13746, N18684, N19887);
xor XOR2 (N24045, N24042, N12965);
xor XOR2 (N24046, N24041, N4069);
xor XOR2 (N24047, N24043, N3393);
or OR3 (N24048, N24037, N17902, N17009);
nor NOR4 (N24049, N24045, N16167, N10448, N20052);
or OR2 (N24050, N24044, N14698);
and AND4 (N24051, N24012, N19268, N19249, N17424);
or OR3 (N24052, N24049, N13504, N4556);
not NOT1 (N24053, N24048);
not NOT1 (N24054, N24027);
and AND2 (N24055, N24029, N5896);
xor XOR2 (N24056, N24040, N315);
or OR2 (N24057, N24046, N11286);
nor NOR4 (N24058, N24053, N7688, N17206, N110);
xor XOR2 (N24059, N24055, N1475);
and AND2 (N24060, N24050, N6343);
or OR3 (N24061, N24052, N18239, N7080);
or OR2 (N24062, N24060, N145);
not NOT1 (N24063, N24058);
or OR3 (N24064, N24061, N6418, N16318);
not NOT1 (N24065, N24063);
not NOT1 (N24066, N24047);
or OR3 (N24067, N24054, N10423, N13720);
buf BUF1 (N24068, N24051);
not NOT1 (N24069, N24067);
and AND4 (N24070, N24069, N12673, N10550, N7091);
or OR2 (N24071, N24068, N1037);
nor NOR3 (N24072, N24030, N10663, N12771);
or OR4 (N24073, N24066, N4393, N10917, N5476);
and AND3 (N24074, N24065, N20023, N22879);
nand NAND2 (N24075, N24056, N22142);
nor NOR4 (N24076, N24071, N11464, N2244, N9671);
or OR2 (N24077, N24070, N2395);
and AND3 (N24078, N24075, N22852, N21926);
or OR4 (N24079, N24062, N9685, N8115, N20702);
and AND2 (N24080, N24059, N2412);
and AND2 (N24081, N24078, N17131);
xor XOR2 (N24082, N24080, N16673);
nand NAND3 (N24083, N24082, N18776, N3506);
xor XOR2 (N24084, N24081, N5657);
buf BUF1 (N24085, N24057);
buf BUF1 (N24086, N24073);
xor XOR2 (N24087, N24083, N17528);
nand NAND4 (N24088, N24072, N5779, N2395, N10767);
xor XOR2 (N24089, N24085, N3182);
and AND3 (N24090, N24074, N12788, N16943);
xor XOR2 (N24091, N24089, N10828);
nand NAND3 (N24092, N24079, N11235, N13001);
not NOT1 (N24093, N24077);
nor NOR4 (N24094, N24088, N20851, N2071, N16741);
buf BUF1 (N24095, N24084);
xor XOR2 (N24096, N24086, N6629);
or OR2 (N24097, N24094, N18959);
nor NOR4 (N24098, N24087, N21766, N19643, N6971);
or OR2 (N24099, N24092, N665);
nand NAND3 (N24100, N24093, N17024, N4453);
not NOT1 (N24101, N24090);
and AND4 (N24102, N24100, N9314, N3390, N19684);
not NOT1 (N24103, N24099);
and AND2 (N24104, N24101, N18811);
and AND2 (N24105, N24076, N16050);
nor NOR3 (N24106, N24103, N12783, N1313);
nor NOR3 (N24107, N24102, N10373, N17177);
and AND2 (N24108, N24107, N22200);
nand NAND3 (N24109, N24106, N10208, N6686);
xor XOR2 (N24110, N24109, N2707);
xor XOR2 (N24111, N24098, N13604);
not NOT1 (N24112, N24105);
not NOT1 (N24113, N24112);
or OR2 (N24114, N24096, N1627);
nand NAND2 (N24115, N24064, N21153);
not NOT1 (N24116, N24114);
and AND4 (N24117, N24113, N4170, N7185, N12235);
and AND4 (N24118, N24104, N4305, N17963, N5067);
or OR3 (N24119, N24091, N117, N10924);
nand NAND2 (N24120, N24118, N3196);
and AND2 (N24121, N24111, N6336);
buf BUF1 (N24122, N24121);
or OR3 (N24123, N24110, N10585, N11147);
xor XOR2 (N24124, N24120, N6906);
or OR2 (N24125, N24117, N11986);
nor NOR3 (N24126, N24108, N18774, N22168);
nor NOR2 (N24127, N24115, N14665);
xor XOR2 (N24128, N24126, N6364);
xor XOR2 (N24129, N24123, N13144);
nor NOR2 (N24130, N24097, N877);
not NOT1 (N24131, N24124);
buf BUF1 (N24132, N24129);
nand NAND2 (N24133, N24132, N16174);
buf BUF1 (N24134, N24133);
not NOT1 (N24135, N24128);
not NOT1 (N24136, N24125);
nand NAND3 (N24137, N24119, N20896, N5679);
and AND4 (N24138, N24131, N5189, N10897, N18043);
buf BUF1 (N24139, N24134);
nand NAND3 (N24140, N24137, N10314, N21999);
not NOT1 (N24141, N24139);
nand NAND4 (N24142, N24140, N14221, N5913, N9860);
xor XOR2 (N24143, N24141, N11772);
nor NOR2 (N24144, N24135, N7318);
not NOT1 (N24145, N24116);
and AND4 (N24146, N24136, N15682, N22343, N385);
or OR4 (N24147, N24144, N1771, N9300, N19177);
nor NOR4 (N24148, N24142, N6413, N14480, N11692);
nand NAND4 (N24149, N24127, N16010, N1093, N4635);
nand NAND3 (N24150, N24145, N21325, N10628);
buf BUF1 (N24151, N24122);
nor NOR2 (N24152, N24130, N5437);
xor XOR2 (N24153, N24095, N23233);
nor NOR2 (N24154, N24138, N5585);
nor NOR4 (N24155, N24153, N21936, N22728, N243);
and AND4 (N24156, N24152, N6525, N6826, N17983);
nor NOR3 (N24157, N24156, N9992, N4177);
not NOT1 (N24158, N24146);
nor NOR4 (N24159, N24155, N3609, N7724, N15837);
nor NOR4 (N24160, N24148, N8752, N8838, N6265);
nand NAND2 (N24161, N24154, N13768);
not NOT1 (N24162, N24147);
nor NOR3 (N24163, N24150, N17971, N5425);
nand NAND2 (N24164, N24163, N8858);
and AND4 (N24165, N24143, N9559, N16998, N10539);
not NOT1 (N24166, N24157);
nand NAND4 (N24167, N24158, N22510, N15572, N12763);
buf BUF1 (N24168, N24161);
and AND3 (N24169, N24167, N16158, N22672);
buf BUF1 (N24170, N24169);
and AND4 (N24171, N24162, N2664, N8349, N20664);
nand NAND3 (N24172, N24159, N12381, N19886);
nand NAND4 (N24173, N24170, N2054, N2027, N20457);
nand NAND2 (N24174, N24173, N5451);
buf BUF1 (N24175, N24171);
nor NOR3 (N24176, N24160, N13876, N12500);
nor NOR2 (N24177, N24176, N14942);
nand NAND3 (N24178, N24149, N20982, N4923);
nor NOR2 (N24179, N24151, N7410);
not NOT1 (N24180, N24175);
and AND3 (N24181, N24164, N1954, N5060);
and AND4 (N24182, N24174, N20051, N4097, N1252);
nand NAND4 (N24183, N24177, N18415, N19405, N20174);
and AND4 (N24184, N24179, N5071, N9694, N15845);
xor XOR2 (N24185, N24182, N2444);
xor XOR2 (N24186, N24172, N16205);
xor XOR2 (N24187, N24178, N11735);
buf BUF1 (N24188, N24184);
nand NAND2 (N24189, N24181, N23758);
nor NOR3 (N24190, N24180, N398, N11897);
not NOT1 (N24191, N24185);
nor NOR4 (N24192, N24189, N3464, N22742, N12591);
and AND3 (N24193, N24186, N1328, N4351);
or OR3 (N24194, N24183, N8559, N19064);
or OR2 (N24195, N24166, N8484);
nor NOR3 (N24196, N24191, N9340, N4406);
not NOT1 (N24197, N24193);
and AND3 (N24198, N24196, N18180, N4792);
nor NOR2 (N24199, N24197, N354);
nor NOR2 (N24200, N24190, N9639);
or OR4 (N24201, N24168, N11782, N17084, N2862);
buf BUF1 (N24202, N24200);
xor XOR2 (N24203, N24192, N16545);
or OR4 (N24204, N24188, N21254, N7140, N23318);
xor XOR2 (N24205, N24201, N18593);
and AND2 (N24206, N24203, N7661);
nand NAND4 (N24207, N24204, N8855, N15442, N21625);
buf BUF1 (N24208, N24202);
and AND3 (N24209, N24165, N2126, N10600);
or OR2 (N24210, N24198, N7452);
buf BUF1 (N24211, N24209);
nor NOR2 (N24212, N24195, N19431);
nand NAND3 (N24213, N24208, N24011, N23809);
buf BUF1 (N24214, N24187);
or OR4 (N24215, N24205, N22184, N18732, N6981);
buf BUF1 (N24216, N24212);
or OR2 (N24217, N24206, N21244);
nand NAND2 (N24218, N24213, N20412);
or OR2 (N24219, N24210, N13534);
nand NAND3 (N24220, N24207, N1981, N3930);
and AND3 (N24221, N24199, N8147, N12838);
or OR4 (N24222, N24211, N2029, N20295, N8589);
nor NOR3 (N24223, N24220, N3176, N17938);
nor NOR3 (N24224, N24194, N14259, N9348);
not NOT1 (N24225, N24217);
buf BUF1 (N24226, N24216);
and AND2 (N24227, N24218, N6894);
or OR3 (N24228, N24227, N16905, N19158);
or OR3 (N24229, N24219, N16755, N320);
xor XOR2 (N24230, N24225, N5471);
nor NOR4 (N24231, N24226, N1771, N6448, N22002);
xor XOR2 (N24232, N24221, N16723);
nand NAND4 (N24233, N24222, N18021, N1022, N20540);
buf BUF1 (N24234, N24228);
or OR3 (N24235, N24233, N15144, N9673);
not NOT1 (N24236, N24234);
or OR4 (N24237, N24231, N23770, N1603, N20904);
and AND4 (N24238, N24229, N4292, N7960, N17405);
nor NOR3 (N24239, N24232, N21712, N23147);
xor XOR2 (N24240, N24224, N5755);
nand NAND2 (N24241, N24239, N17333);
xor XOR2 (N24242, N24240, N14421);
not NOT1 (N24243, N24236);
xor XOR2 (N24244, N24243, N12737);
nand NAND4 (N24245, N24214, N6094, N6747, N911);
nor NOR4 (N24246, N24245, N16653, N16574, N16691);
buf BUF1 (N24247, N24235);
and AND3 (N24248, N24246, N18452, N23878);
nand NAND4 (N24249, N24241, N24247, N13278, N10216);
not NOT1 (N24250, N4476);
and AND3 (N24251, N24242, N8066, N1084);
nand NAND2 (N24252, N24249, N19943);
and AND4 (N24253, N24230, N16687, N4239, N23095);
nor NOR3 (N24254, N24244, N4829, N13103);
nand NAND2 (N24255, N24253, N21353);
buf BUF1 (N24256, N24237);
or OR3 (N24257, N24256, N10783, N19521);
buf BUF1 (N24258, N24257);
not NOT1 (N24259, N24248);
xor XOR2 (N24260, N24255, N6790);
not NOT1 (N24261, N24238);
xor XOR2 (N24262, N24252, N18821);
or OR3 (N24263, N24254, N11285, N6207);
or OR4 (N24264, N24251, N14508, N2106, N10325);
nand NAND2 (N24265, N24264, N19407);
and AND4 (N24266, N24263, N21549, N4519, N17014);
nor NOR2 (N24267, N24223, N6980);
xor XOR2 (N24268, N24262, N10407);
nand NAND2 (N24269, N24265, N3216);
or OR3 (N24270, N24260, N13378, N18140);
or OR3 (N24271, N24215, N18084, N8866);
xor XOR2 (N24272, N24269, N15259);
not NOT1 (N24273, N24271);
nand NAND3 (N24274, N24259, N6938, N19101);
xor XOR2 (N24275, N24268, N572);
nand NAND3 (N24276, N24261, N14831, N2341);
nand NAND2 (N24277, N24270, N15345);
nand NAND4 (N24278, N24273, N8315, N8798, N22566);
nand NAND2 (N24279, N24277, N7033);
or OR3 (N24280, N24275, N11955, N14405);
xor XOR2 (N24281, N24272, N3023);
nor NOR3 (N24282, N24267, N215, N6995);
nand NAND3 (N24283, N24274, N14672, N17646);
or OR2 (N24284, N24279, N3890);
buf BUF1 (N24285, N24284);
or OR2 (N24286, N24278, N9264);
buf BUF1 (N24287, N24286);
nand NAND2 (N24288, N24282, N2544);
and AND4 (N24289, N24283, N20607, N16886, N8806);
nor NOR4 (N24290, N24285, N20910, N6250, N8589);
buf BUF1 (N24291, N24289);
nor NOR3 (N24292, N24281, N19765, N363);
nor NOR2 (N24293, N24266, N9367);
xor XOR2 (N24294, N24276, N10570);
or OR3 (N24295, N24294, N21629, N15722);
buf BUF1 (N24296, N24287);
nand NAND3 (N24297, N24291, N2327, N7088);
xor XOR2 (N24298, N24292, N17157);
or OR4 (N24299, N24298, N9208, N5251, N11458);
not NOT1 (N24300, N24297);
or OR4 (N24301, N24295, N22180, N15798, N9460);
nor NOR4 (N24302, N24290, N7134, N6287, N22759);
nor NOR2 (N24303, N24300, N13182);
nor NOR3 (N24304, N24301, N261, N8584);
nand NAND4 (N24305, N24293, N23765, N137, N3159);
nor NOR2 (N24306, N24303, N22708);
nand NAND2 (N24307, N24306, N4673);
buf BUF1 (N24308, N24307);
xor XOR2 (N24309, N24258, N10556);
and AND2 (N24310, N24304, N3441);
or OR3 (N24311, N24309, N5490, N19412);
xor XOR2 (N24312, N24311, N22864);
and AND4 (N24313, N24288, N18555, N12268, N14101);
not NOT1 (N24314, N24313);
nand NAND4 (N24315, N24296, N14195, N15084, N18776);
buf BUF1 (N24316, N24312);
not NOT1 (N24317, N24280);
or OR2 (N24318, N24299, N7476);
and AND4 (N24319, N24302, N24121, N19699, N14758);
nand NAND3 (N24320, N24308, N23004, N10394);
nor NOR2 (N24321, N24317, N15975);
and AND4 (N24322, N24321, N21569, N21281, N17273);
or OR4 (N24323, N24319, N1392, N4541, N9014);
buf BUF1 (N24324, N24305);
nand NAND4 (N24325, N24315, N11629, N6912, N14151);
nand NAND2 (N24326, N24316, N13487);
nand NAND4 (N24327, N24320, N16068, N11544, N3322);
nand NAND4 (N24328, N24318, N1932, N18350, N1416);
nand NAND2 (N24329, N24327, N9129);
nor NOR2 (N24330, N24325, N1679);
nand NAND4 (N24331, N24324, N2228, N10113, N20817);
nand NAND3 (N24332, N24328, N5619, N14586);
buf BUF1 (N24333, N24310);
nand NAND3 (N24334, N24331, N18782, N16828);
xor XOR2 (N24335, N24333, N12573);
xor XOR2 (N24336, N24330, N9649);
and AND2 (N24337, N24322, N19792);
buf BUF1 (N24338, N24337);
xor XOR2 (N24339, N24338, N9904);
buf BUF1 (N24340, N24326);
buf BUF1 (N24341, N24329);
buf BUF1 (N24342, N24332);
xor XOR2 (N24343, N24339, N14993);
nor NOR3 (N24344, N24335, N5350, N11560);
xor XOR2 (N24345, N24340, N8463);
not NOT1 (N24346, N24334);
buf BUF1 (N24347, N24344);
or OR4 (N24348, N24345, N8605, N9051, N15169);
not NOT1 (N24349, N24342);
not NOT1 (N24350, N24347);
nand NAND2 (N24351, N24343, N3622);
or OR4 (N24352, N24314, N3262, N4475, N13965);
nand NAND2 (N24353, N24350, N12413);
xor XOR2 (N24354, N24323, N2239);
buf BUF1 (N24355, N24354);
nand NAND2 (N24356, N24336, N12711);
and AND2 (N24357, N24346, N2532);
and AND4 (N24358, N24356, N7982, N17031, N4695);
xor XOR2 (N24359, N24357, N15200);
and AND3 (N24360, N24353, N15132, N9723);
nand NAND2 (N24361, N24349, N841);
xor XOR2 (N24362, N24361, N13013);
nor NOR3 (N24363, N24359, N15800, N13290);
and AND2 (N24364, N24362, N12608);
not NOT1 (N24365, N24355);
or OR2 (N24366, N24358, N10992);
and AND4 (N24367, N24250, N23037, N21478, N6867);
and AND3 (N24368, N24348, N11578, N665);
nand NAND4 (N24369, N24367, N6531, N13046, N13553);
buf BUF1 (N24370, N24368);
and AND4 (N24371, N24360, N2938, N22794, N10280);
or OR2 (N24372, N24370, N12075);
nor NOR3 (N24373, N24352, N11533, N1614);
or OR4 (N24374, N24373, N4072, N2491, N4023);
not NOT1 (N24375, N24372);
nand NAND3 (N24376, N24369, N10615, N14621);
xor XOR2 (N24377, N24376, N8404);
xor XOR2 (N24378, N24341, N18100);
buf BUF1 (N24379, N24375);
not NOT1 (N24380, N24377);
nor NOR3 (N24381, N24366, N14361, N17962);
buf BUF1 (N24382, N24371);
or OR3 (N24383, N24364, N12548, N9996);
xor XOR2 (N24384, N24363, N13956);
buf BUF1 (N24385, N24351);
and AND4 (N24386, N24378, N9173, N16650, N10975);
xor XOR2 (N24387, N24384, N17158);
and AND4 (N24388, N24381, N105, N17341, N12464);
nand NAND4 (N24389, N24380, N13109, N13682, N20650);
nand NAND2 (N24390, N24388, N15814);
buf BUF1 (N24391, N24365);
xor XOR2 (N24392, N24391, N1954);
buf BUF1 (N24393, N24379);
nor NOR3 (N24394, N24383, N22316, N22833);
nand NAND3 (N24395, N24393, N9801, N8863);
buf BUF1 (N24396, N24386);
buf BUF1 (N24397, N24392);
nor NOR3 (N24398, N24387, N16461, N21402);
or OR4 (N24399, N24398, N17123, N7917, N19229);
not NOT1 (N24400, N24385);
nor NOR3 (N24401, N24394, N13708, N3210);
buf BUF1 (N24402, N24401);
buf BUF1 (N24403, N24395);
not NOT1 (N24404, N24399);
nor NOR2 (N24405, N24382, N8495);
nor NOR4 (N24406, N24389, N18983, N10486, N8505);
not NOT1 (N24407, N24405);
nand NAND3 (N24408, N24374, N21995, N1883);
buf BUF1 (N24409, N24396);
not NOT1 (N24410, N24407);
nor NOR4 (N24411, N24408, N3986, N23424, N18142);
nand NAND4 (N24412, N24410, N454, N21194, N18880);
buf BUF1 (N24413, N24404);
xor XOR2 (N24414, N24403, N11435);
or OR3 (N24415, N24412, N8131, N13919);
xor XOR2 (N24416, N24400, N19359);
nand NAND2 (N24417, N24409, N5142);
nor NOR4 (N24418, N24413, N19889, N1912, N1951);
nand NAND3 (N24419, N24415, N3737, N546);
nor NOR2 (N24420, N24414, N21268);
nor NOR2 (N24421, N24418, N3582);
buf BUF1 (N24422, N24390);
or OR3 (N24423, N24411, N8007, N21872);
and AND2 (N24424, N24406, N10300);
not NOT1 (N24425, N24417);
nand NAND3 (N24426, N24419, N6808, N12061);
or OR2 (N24427, N24421, N20363);
and AND2 (N24428, N24424, N6898);
buf BUF1 (N24429, N24428);
buf BUF1 (N24430, N24402);
or OR2 (N24431, N24416, N9219);
nand NAND2 (N24432, N24429, N24316);
xor XOR2 (N24433, N24431, N15538);
nor NOR3 (N24434, N24397, N14343, N5288);
not NOT1 (N24435, N24427);
nand NAND2 (N24436, N24432, N20348);
not NOT1 (N24437, N24433);
nand NAND2 (N24438, N24422, N15310);
xor XOR2 (N24439, N24426, N16950);
not NOT1 (N24440, N24437);
nand NAND2 (N24441, N24425, N11724);
and AND3 (N24442, N24439, N11777, N24337);
xor XOR2 (N24443, N24435, N14610);
buf BUF1 (N24444, N24434);
nand NAND4 (N24445, N24423, N17406, N17606, N1002);
xor XOR2 (N24446, N24441, N6212);
xor XOR2 (N24447, N24436, N20679);
or OR4 (N24448, N24420, N2780, N954, N7939);
buf BUF1 (N24449, N24442);
nor NOR2 (N24450, N24449, N5018);
or OR2 (N24451, N24443, N22359);
nand NAND2 (N24452, N24447, N22671);
xor XOR2 (N24453, N24451, N7256);
not NOT1 (N24454, N24445);
and AND2 (N24455, N24450, N3042);
and AND4 (N24456, N24453, N15633, N23978, N7718);
or OR3 (N24457, N24430, N2233, N6049);
xor XOR2 (N24458, N24448, N292);
not NOT1 (N24459, N24457);
xor XOR2 (N24460, N24455, N6688);
and AND3 (N24461, N24456, N11424, N22454);
nor NOR2 (N24462, N24458, N2441);
nand NAND2 (N24463, N24461, N23916);
nand NAND3 (N24464, N24454, N19231, N2214);
buf BUF1 (N24465, N24440);
and AND4 (N24466, N24446, N3655, N14531, N6042);
buf BUF1 (N24467, N24463);
buf BUF1 (N24468, N24462);
xor XOR2 (N24469, N24460, N7758);
nor NOR4 (N24470, N24452, N3493, N14516, N4181);
nor NOR2 (N24471, N24465, N5662);
xor XOR2 (N24472, N24468, N2071);
not NOT1 (N24473, N24464);
xor XOR2 (N24474, N24466, N439);
buf BUF1 (N24475, N24469);
nor NOR2 (N24476, N24467, N19158);
or OR3 (N24477, N24438, N18962, N13805);
xor XOR2 (N24478, N24475, N17233);
xor XOR2 (N24479, N24474, N20977);
or OR3 (N24480, N24479, N14612, N21553);
buf BUF1 (N24481, N24473);
buf BUF1 (N24482, N24470);
nor NOR3 (N24483, N24476, N16407, N6899);
nor NOR2 (N24484, N24480, N19507);
buf BUF1 (N24485, N24481);
or OR2 (N24486, N24484, N11690);
or OR4 (N24487, N24478, N14633, N20342, N14499);
not NOT1 (N24488, N24459);
not NOT1 (N24489, N24487);
nand NAND3 (N24490, N24472, N5131, N6708);
xor XOR2 (N24491, N24485, N2610);
or OR3 (N24492, N24471, N11798, N20731);
or OR3 (N24493, N24486, N15651, N17677);
nand NAND4 (N24494, N24444, N18994, N18468, N23791);
nand NAND2 (N24495, N24483, N21976);
buf BUF1 (N24496, N24491);
not NOT1 (N24497, N24488);
xor XOR2 (N24498, N24489, N690);
xor XOR2 (N24499, N24495, N5312);
or OR4 (N24500, N24497, N8523, N12270, N10443);
or OR4 (N24501, N24499, N5077, N18216, N20165);
and AND2 (N24502, N24494, N18855);
xor XOR2 (N24503, N24501, N5563);
not NOT1 (N24504, N24492);
not NOT1 (N24505, N24504);
buf BUF1 (N24506, N24477);
not NOT1 (N24507, N24506);
and AND3 (N24508, N24503, N1436, N20715);
nand NAND3 (N24509, N24502, N3848, N7990);
or OR3 (N24510, N24490, N8013, N13334);
nor NOR3 (N24511, N24482, N23378, N22067);
nand NAND2 (N24512, N24511, N7396);
xor XOR2 (N24513, N24498, N1314);
and AND2 (N24514, N24505, N23395);
not NOT1 (N24515, N24493);
nor NOR2 (N24516, N24513, N7755);
and AND2 (N24517, N24507, N21792);
and AND3 (N24518, N24512, N23882, N12342);
nor NOR3 (N24519, N24518, N3740, N5467);
buf BUF1 (N24520, N24515);
buf BUF1 (N24521, N24496);
xor XOR2 (N24522, N24519, N1309);
and AND2 (N24523, N24514, N3657);
and AND3 (N24524, N24521, N3480, N3288);
and AND3 (N24525, N24516, N4588, N20916);
or OR4 (N24526, N24500, N16634, N1015, N18363);
or OR2 (N24527, N24525, N2173);
nand NAND2 (N24528, N24524, N19466);
xor XOR2 (N24529, N24509, N16143);
not NOT1 (N24530, N24508);
nand NAND4 (N24531, N24522, N4228, N4768, N3080);
and AND4 (N24532, N24529, N7275, N2793, N13982);
not NOT1 (N24533, N24526);
buf BUF1 (N24534, N24528);
nand NAND3 (N24535, N24517, N12088, N8511);
xor XOR2 (N24536, N24523, N16554);
nor NOR4 (N24537, N24510, N378, N2352, N9053);
xor XOR2 (N24538, N24530, N2214);
xor XOR2 (N24539, N24527, N12152);
buf BUF1 (N24540, N24537);
and AND2 (N24541, N24536, N19621);
or OR2 (N24542, N24541, N17101);
buf BUF1 (N24543, N24539);
nor NOR4 (N24544, N24538, N10838, N15954, N1515);
nor NOR2 (N24545, N24534, N4712);
or OR3 (N24546, N24542, N13052, N13819);
not NOT1 (N24547, N24544);
or OR4 (N24548, N24520, N218, N3523, N7500);
nand NAND3 (N24549, N24540, N2838, N6550);
not NOT1 (N24550, N24545);
and AND4 (N24551, N24546, N14382, N1408, N20821);
buf BUF1 (N24552, N24547);
and AND3 (N24553, N24535, N2836, N17844);
xor XOR2 (N24554, N24551, N9569);
not NOT1 (N24555, N24548);
and AND4 (N24556, N24554, N3724, N13833, N17899);
xor XOR2 (N24557, N24532, N9765);
not NOT1 (N24558, N24531);
xor XOR2 (N24559, N24553, N22259);
nand NAND3 (N24560, N24557, N20123, N7176);
nand NAND2 (N24561, N24558, N943);
or OR3 (N24562, N24556, N15470, N22423);
buf BUF1 (N24563, N24561);
xor XOR2 (N24564, N24559, N22925);
buf BUF1 (N24565, N24543);
buf BUF1 (N24566, N24564);
not NOT1 (N24567, N24562);
or OR2 (N24568, N24533, N1247);
or OR3 (N24569, N24550, N10768, N16957);
or OR4 (N24570, N24568, N5346, N2739, N74);
or OR3 (N24571, N24552, N5863, N7419);
xor XOR2 (N24572, N24566, N3614);
not NOT1 (N24573, N24570);
xor XOR2 (N24574, N24567, N18746);
or OR3 (N24575, N24563, N5990, N6853);
not NOT1 (N24576, N24549);
not NOT1 (N24577, N24565);
not NOT1 (N24578, N24573);
xor XOR2 (N24579, N24555, N3132);
nor NOR2 (N24580, N24571, N19558);
nor NOR4 (N24581, N24579, N2854, N12857, N20689);
buf BUF1 (N24582, N24580);
nand NAND4 (N24583, N24577, N7896, N12725, N9082);
nor NOR4 (N24584, N24575, N20951, N23347, N15816);
nor NOR4 (N24585, N24576, N9724, N23596, N19113);
buf BUF1 (N24586, N24585);
xor XOR2 (N24587, N24584, N5197);
or OR2 (N24588, N24581, N17308);
xor XOR2 (N24589, N24583, N17563);
nor NOR2 (N24590, N24582, N18882);
and AND3 (N24591, N24578, N270, N19028);
buf BUF1 (N24592, N24569);
nand NAND4 (N24593, N24586, N3520, N21923, N17273);
nand NAND3 (N24594, N24592, N5276, N18558);
and AND2 (N24595, N24572, N6119);
nor NOR2 (N24596, N24589, N13474);
buf BUF1 (N24597, N24593);
not NOT1 (N24598, N24597);
xor XOR2 (N24599, N24591, N1264);
or OR4 (N24600, N24574, N9669, N6184, N4851);
nor NOR2 (N24601, N24587, N20505);
nor NOR3 (N24602, N24598, N953, N22127);
nand NAND3 (N24603, N24599, N17107, N20371);
nor NOR4 (N24604, N24603, N20725, N19417, N21992);
and AND2 (N24605, N24601, N22140);
nand NAND3 (N24606, N24560, N12841, N10793);
nand NAND2 (N24607, N24606, N10241);
not NOT1 (N24608, N24588);
nor NOR3 (N24609, N24607, N20439, N17319);
xor XOR2 (N24610, N24608, N5454);
and AND3 (N24611, N24602, N14586, N15654);
xor XOR2 (N24612, N24594, N21422);
nor NOR2 (N24613, N24611, N20144);
nor NOR2 (N24614, N24613, N9252);
buf BUF1 (N24615, N24596);
not NOT1 (N24616, N24614);
buf BUF1 (N24617, N24609);
buf BUF1 (N24618, N24610);
buf BUF1 (N24619, N24600);
nor NOR3 (N24620, N24617, N8909, N7293);
nor NOR2 (N24621, N24618, N12869);
or OR2 (N24622, N24612, N895);
xor XOR2 (N24623, N24604, N18758);
xor XOR2 (N24624, N24590, N3894);
buf BUF1 (N24625, N24622);
nor NOR2 (N24626, N24595, N23260);
and AND2 (N24627, N24620, N9359);
nand NAND3 (N24628, N24619, N13340, N2299);
nand NAND4 (N24629, N24625, N2837, N401, N23605);
xor XOR2 (N24630, N24626, N23171);
not NOT1 (N24631, N24623);
buf BUF1 (N24632, N24615);
nand NAND2 (N24633, N24621, N22387);
xor XOR2 (N24634, N24624, N12387);
nand NAND3 (N24635, N24634, N11847, N18038);
buf BUF1 (N24636, N24631);
or OR3 (N24637, N24630, N17678, N11481);
buf BUF1 (N24638, N24635);
or OR3 (N24639, N24605, N2528, N21106);
nor NOR2 (N24640, N24616, N7059);
nor NOR3 (N24641, N24639, N17794, N12915);
and AND4 (N24642, N24628, N9502, N20983, N177);
or OR4 (N24643, N24633, N924, N11834, N6854);
xor XOR2 (N24644, N24641, N14849);
and AND3 (N24645, N24636, N14907, N16854);
nor NOR4 (N24646, N24642, N13159, N15101, N23286);
nor NOR4 (N24647, N24644, N11566, N17404, N6018);
and AND4 (N24648, N24645, N11756, N17382, N8366);
nand NAND3 (N24649, N24627, N24354, N23555);
and AND2 (N24650, N24646, N5847);
or OR4 (N24651, N24632, N3771, N21588, N22500);
and AND4 (N24652, N24649, N9185, N19036, N18088);
not NOT1 (N24653, N24648);
buf BUF1 (N24654, N24637);
or OR4 (N24655, N24654, N2813, N21556, N18610);
xor XOR2 (N24656, N24643, N3094);
or OR4 (N24657, N24652, N21466, N13917, N14376);
nor NOR4 (N24658, N24651, N16912, N15053, N19068);
not NOT1 (N24659, N24650);
and AND4 (N24660, N24659, N15858, N4219, N8925);
xor XOR2 (N24661, N24660, N14829);
xor XOR2 (N24662, N24656, N344);
nand NAND2 (N24663, N24640, N12357);
not NOT1 (N24664, N24657);
buf BUF1 (N24665, N24663);
buf BUF1 (N24666, N24653);
nor NOR4 (N24667, N24658, N15411, N15417, N19023);
xor XOR2 (N24668, N24665, N20990);
nand NAND4 (N24669, N24647, N8178, N6091, N5571);
buf BUF1 (N24670, N24661);
nand NAND4 (N24671, N24668, N21898, N13039, N12013);
nor NOR3 (N24672, N24662, N12439, N22324);
nor NOR4 (N24673, N24629, N11333, N323, N19810);
or OR3 (N24674, N24669, N5580, N4433);
xor XOR2 (N24675, N24670, N18034);
not NOT1 (N24676, N24675);
nor NOR2 (N24677, N24667, N2023);
xor XOR2 (N24678, N24638, N1971);
not NOT1 (N24679, N24655);
nor NOR2 (N24680, N24679, N10272);
xor XOR2 (N24681, N24673, N13350);
not NOT1 (N24682, N24674);
not NOT1 (N24683, N24681);
buf BUF1 (N24684, N24682);
nand NAND4 (N24685, N24680, N17720, N9723, N19628);
or OR4 (N24686, N24677, N10123, N19489, N23934);
nand NAND3 (N24687, N24676, N845, N8867);
not NOT1 (N24688, N24686);
buf BUF1 (N24689, N24684);
nor NOR3 (N24690, N24664, N23772, N5551);
or OR2 (N24691, N24688, N12232);
xor XOR2 (N24692, N24678, N447);
buf BUF1 (N24693, N24672);
and AND3 (N24694, N24691, N5469, N23052);
nor NOR3 (N24695, N24690, N15628, N13569);
not NOT1 (N24696, N24671);
nand NAND4 (N24697, N24695, N17712, N20769, N10710);
and AND3 (N24698, N24692, N1485, N9668);
or OR2 (N24699, N24666, N20963);
nand NAND2 (N24700, N24689, N18660);
and AND2 (N24701, N24698, N23330);
and AND2 (N24702, N24693, N13691);
buf BUF1 (N24703, N24702);
or OR3 (N24704, N24703, N14393, N21416);
nor NOR3 (N24705, N24696, N14264, N5722);
xor XOR2 (N24706, N24701, N23508);
buf BUF1 (N24707, N24700);
not NOT1 (N24708, N24683);
xor XOR2 (N24709, N24705, N20757);
not NOT1 (N24710, N24687);
xor XOR2 (N24711, N24708, N4420);
and AND4 (N24712, N24704, N3134, N6506, N9701);
nor NOR4 (N24713, N24697, N20013, N9608, N4465);
or OR4 (N24714, N24694, N3611, N1809, N10555);
xor XOR2 (N24715, N24713, N18550);
and AND4 (N24716, N24709, N17444, N3140, N8206);
and AND2 (N24717, N24716, N19235);
buf BUF1 (N24718, N24710);
or OR3 (N24719, N24715, N9560, N7091);
and AND3 (N24720, N24719, N15994, N15838);
xor XOR2 (N24721, N24706, N5429);
nand NAND4 (N24722, N24721, N616, N3597, N13561);
or OR3 (N24723, N24722, N16767, N17094);
nand NAND3 (N24724, N24707, N13946, N9779);
nand NAND3 (N24725, N24714, N11869, N3410);
or OR2 (N24726, N24718, N17544);
buf BUF1 (N24727, N24685);
nand NAND2 (N24728, N24726, N16530);
or OR2 (N24729, N24699, N21359);
and AND4 (N24730, N24725, N22288, N12521, N8031);
or OR4 (N24731, N24723, N14738, N8779, N18116);
nor NOR3 (N24732, N24712, N9062, N3128);
and AND3 (N24733, N24720, N11675, N10791);
nand NAND4 (N24734, N24711, N2437, N22834, N863);
buf BUF1 (N24735, N24734);
xor XOR2 (N24736, N24729, N10920);
nand NAND3 (N24737, N24732, N19019, N19961);
or OR3 (N24738, N24730, N11114, N219);
not NOT1 (N24739, N24728);
buf BUF1 (N24740, N24731);
not NOT1 (N24741, N24727);
buf BUF1 (N24742, N24737);
or OR4 (N24743, N24740, N7121, N633, N1046);
not NOT1 (N24744, N24733);
nand NAND4 (N24745, N24717, N24512, N24226, N20187);
not NOT1 (N24746, N24736);
and AND4 (N24747, N24742, N19020, N5389, N22876);
xor XOR2 (N24748, N24741, N16147);
xor XOR2 (N24749, N24743, N13383);
nor NOR2 (N24750, N24735, N5008);
not NOT1 (N24751, N24724);
nand NAND2 (N24752, N24748, N23960);
and AND4 (N24753, N24745, N4831, N2449, N3379);
xor XOR2 (N24754, N24750, N8005);
and AND2 (N24755, N24739, N6851);
and AND3 (N24756, N24755, N5028, N10495);
not NOT1 (N24757, N24751);
and AND2 (N24758, N24746, N9566);
nor NOR4 (N24759, N24752, N12210, N11862, N22619);
buf BUF1 (N24760, N24759);
and AND3 (N24761, N24744, N21992, N12060);
xor XOR2 (N24762, N24753, N8910);
nor NOR2 (N24763, N24754, N13375);
nand NAND3 (N24764, N24758, N2843, N84);
and AND2 (N24765, N24762, N22141);
and AND4 (N24766, N24749, N180, N22943, N7450);
nand NAND4 (N24767, N24747, N18295, N3910, N4251);
and AND3 (N24768, N24761, N11825, N3363);
nand NAND4 (N24769, N24757, N5796, N17025, N9012);
and AND4 (N24770, N24738, N15308, N5871, N21776);
buf BUF1 (N24771, N24765);
and AND4 (N24772, N24764, N16166, N20334, N20411);
nor NOR2 (N24773, N24769, N12389);
not NOT1 (N24774, N24771);
not NOT1 (N24775, N24756);
buf BUF1 (N24776, N24767);
buf BUF1 (N24777, N24773);
buf BUF1 (N24778, N24770);
nand NAND3 (N24779, N24763, N17049, N21599);
not NOT1 (N24780, N24772);
not NOT1 (N24781, N24780);
nand NAND4 (N24782, N24760, N8337, N4402, N19504);
nand NAND2 (N24783, N24768, N22919);
nor NOR4 (N24784, N24783, N126, N19738, N20722);
or OR2 (N24785, N24776, N18485);
nor NOR4 (N24786, N24785, N12584, N23293, N12906);
and AND2 (N24787, N24774, N6451);
not NOT1 (N24788, N24782);
not NOT1 (N24789, N24781);
or OR3 (N24790, N24766, N2324, N9004);
xor XOR2 (N24791, N24786, N16410);
xor XOR2 (N24792, N24775, N8788);
not NOT1 (N24793, N24788);
buf BUF1 (N24794, N24779);
buf BUF1 (N24795, N24790);
nand NAND2 (N24796, N24777, N19715);
not NOT1 (N24797, N24794);
not NOT1 (N24798, N24791);
buf BUF1 (N24799, N24797);
nor NOR2 (N24800, N24792, N22578);
not NOT1 (N24801, N24796);
buf BUF1 (N24802, N24798);
not NOT1 (N24803, N24784);
buf BUF1 (N24804, N24799);
xor XOR2 (N24805, N24802, N12373);
and AND4 (N24806, N24801, N3387, N11626, N6832);
not NOT1 (N24807, N24803);
and AND2 (N24808, N24789, N20914);
and AND2 (N24809, N24787, N2698);
not NOT1 (N24810, N24795);
xor XOR2 (N24811, N24807, N3694);
xor XOR2 (N24812, N24778, N21620);
nand NAND2 (N24813, N24811, N23906);
and AND3 (N24814, N24800, N72, N24386);
buf BUF1 (N24815, N24806);
nand NAND4 (N24816, N24805, N6671, N1604, N21976);
nor NOR2 (N24817, N24793, N4274);
nor NOR2 (N24818, N24814, N10406);
or OR3 (N24819, N24808, N18042, N8782);
not NOT1 (N24820, N24812);
not NOT1 (N24821, N24813);
xor XOR2 (N24822, N24818, N11307);
xor XOR2 (N24823, N24821, N13688);
buf BUF1 (N24824, N24819);
nor NOR2 (N24825, N24816, N5542);
buf BUF1 (N24826, N24810);
nand NAND2 (N24827, N24824, N16879);
nand NAND2 (N24828, N24823, N5506);
xor XOR2 (N24829, N24820, N20946);
and AND3 (N24830, N24826, N20334, N19294);
xor XOR2 (N24831, N24827, N948);
or OR4 (N24832, N24829, N20969, N15052, N9368);
not NOT1 (N24833, N24817);
buf BUF1 (N24834, N24833);
or OR3 (N24835, N24809, N8104, N2344);
buf BUF1 (N24836, N24825);
or OR2 (N24837, N24834, N6295);
not NOT1 (N24838, N24835);
nand NAND4 (N24839, N24831, N1262, N1635, N4318);
nor NOR3 (N24840, N24828, N23151, N14941);
not NOT1 (N24841, N24840);
and AND3 (N24842, N24841, N3974, N2643);
nand NAND2 (N24843, N24836, N8765);
not NOT1 (N24844, N24837);
xor XOR2 (N24845, N24822, N18960);
or OR4 (N24846, N24842, N23015, N21595, N6280);
nor NOR3 (N24847, N24839, N23514, N22191);
and AND3 (N24848, N24846, N16065, N18890);
xor XOR2 (N24849, N24838, N8696);
not NOT1 (N24850, N24832);
nor NOR4 (N24851, N24848, N4660, N12915, N24297);
and AND4 (N24852, N24849, N8661, N19297, N24659);
and AND2 (N24853, N24850, N8456);
not NOT1 (N24854, N24830);
and AND2 (N24855, N24845, N22600);
or OR2 (N24856, N24815, N766);
nor NOR4 (N24857, N24856, N11508, N8684, N10112);
not NOT1 (N24858, N24847);
buf BUF1 (N24859, N24858);
nand NAND2 (N24860, N24851, N10180);
buf BUF1 (N24861, N24854);
and AND4 (N24862, N24852, N11735, N11983, N20840);
and AND4 (N24863, N24859, N23865, N9585, N22154);
and AND2 (N24864, N24861, N10893);
xor XOR2 (N24865, N24864, N16370);
nand NAND3 (N24866, N24857, N1877, N23228);
xor XOR2 (N24867, N24853, N16237);
buf BUF1 (N24868, N24855);
nor NOR4 (N24869, N24865, N4899, N5372, N2759);
nor NOR2 (N24870, N24862, N3165);
not NOT1 (N24871, N24870);
or OR3 (N24872, N24860, N625, N5039);
or OR4 (N24873, N24843, N17266, N6593, N1604);
xor XOR2 (N24874, N24844, N4969);
nand NAND4 (N24875, N24871, N1281, N6902, N23421);
nand NAND2 (N24876, N24867, N11689);
nor NOR4 (N24877, N24869, N2231, N6826, N15378);
not NOT1 (N24878, N24875);
nor NOR4 (N24879, N24874, N13333, N9371, N10432);
nor NOR4 (N24880, N24879, N15956, N222, N22076);
or OR4 (N24881, N24873, N9564, N18494, N4920);
not NOT1 (N24882, N24866);
and AND4 (N24883, N24872, N4319, N14205, N23439);
xor XOR2 (N24884, N24868, N6121);
or OR3 (N24885, N24804, N9469, N328);
xor XOR2 (N24886, N24863, N17477);
nor NOR3 (N24887, N24880, N245, N20287);
nand NAND4 (N24888, N24886, N1630, N8867, N13294);
nand NAND3 (N24889, N24885, N5970, N462);
and AND2 (N24890, N24889, N10637);
and AND4 (N24891, N24881, N2510, N10497, N16660);
nand NAND3 (N24892, N24887, N2037, N12163);
nand NAND2 (N24893, N24884, N11154);
and AND2 (N24894, N24878, N2523);
not NOT1 (N24895, N24877);
not NOT1 (N24896, N24892);
buf BUF1 (N24897, N24894);
or OR3 (N24898, N24891, N7714, N21921);
xor XOR2 (N24899, N24883, N20127);
or OR3 (N24900, N24896, N12811, N4604);
xor XOR2 (N24901, N24897, N1352);
nand NAND4 (N24902, N24901, N13800, N10221, N560);
and AND4 (N24903, N24882, N11606, N9073, N12528);
and AND2 (N24904, N24893, N10857);
buf BUF1 (N24905, N24902);
xor XOR2 (N24906, N24888, N15672);
buf BUF1 (N24907, N24903);
buf BUF1 (N24908, N24876);
not NOT1 (N24909, N24890);
xor XOR2 (N24910, N24906, N655);
buf BUF1 (N24911, N24907);
or OR2 (N24912, N24904, N19702);
nor NOR4 (N24913, N24910, N6514, N20661, N3478);
or OR4 (N24914, N24912, N6830, N9695, N15701);
buf BUF1 (N24915, N24914);
not NOT1 (N24916, N24909);
xor XOR2 (N24917, N24899, N8781);
or OR4 (N24918, N24898, N15617, N13324, N23726);
xor XOR2 (N24919, N24918, N16446);
and AND4 (N24920, N24911, N19024, N13777, N24408);
xor XOR2 (N24921, N24920, N22348);
xor XOR2 (N24922, N24900, N20191);
or OR4 (N24923, N24922, N4154, N5974, N10167);
nor NOR3 (N24924, N24905, N88, N14561);
buf BUF1 (N24925, N24916);
nor NOR3 (N24926, N24913, N3881, N7390);
and AND4 (N24927, N24924, N692, N5915, N12348);
and AND3 (N24928, N24919, N10017, N15746);
xor XOR2 (N24929, N24917, N19674);
not NOT1 (N24930, N24895);
nand NAND2 (N24931, N24915, N12147);
xor XOR2 (N24932, N24908, N4067);
buf BUF1 (N24933, N24928);
nand NAND3 (N24934, N24927, N18827, N4487);
or OR2 (N24935, N24930, N20148);
xor XOR2 (N24936, N24935, N10376);
nor NOR2 (N24937, N24926, N12180);
nand NAND3 (N24938, N24931, N9046, N19768);
buf BUF1 (N24939, N24923);
not NOT1 (N24940, N24938);
or OR2 (N24941, N24936, N4268);
not NOT1 (N24942, N24939);
or OR4 (N24943, N24934, N572, N14939, N5550);
not NOT1 (N24944, N24941);
xor XOR2 (N24945, N24942, N19113);
or OR2 (N24946, N24921, N14286);
buf BUF1 (N24947, N24943);
not NOT1 (N24948, N24933);
xor XOR2 (N24949, N24945, N7863);
buf BUF1 (N24950, N24937);
buf BUF1 (N24951, N24929);
and AND2 (N24952, N24925, N6654);
nand NAND3 (N24953, N24940, N18806, N4052);
not NOT1 (N24954, N24951);
not NOT1 (N24955, N24949);
nand NAND3 (N24956, N24946, N3696, N15212);
or OR3 (N24957, N24947, N18244, N7501);
nor NOR2 (N24958, N24954, N24602);
not NOT1 (N24959, N24955);
or OR4 (N24960, N24944, N12825, N13391, N24749);
xor XOR2 (N24961, N24948, N4292);
and AND3 (N24962, N24950, N10649, N16945);
or OR4 (N24963, N24958, N7895, N1694, N19033);
xor XOR2 (N24964, N24960, N3155);
or OR4 (N24965, N24957, N17986, N6141, N24556);
not NOT1 (N24966, N24932);
or OR2 (N24967, N24953, N2442);
or OR2 (N24968, N24959, N18671);
and AND2 (N24969, N24964, N20111);
nor NOR2 (N24970, N24962, N4981);
xor XOR2 (N24971, N24966, N12221);
nand NAND4 (N24972, N24965, N2952, N14451, N7786);
xor XOR2 (N24973, N24963, N22207);
nor NOR2 (N24974, N24968, N23208);
or OR4 (N24975, N24956, N16650, N4295, N12688);
not NOT1 (N24976, N24972);
nor NOR4 (N24977, N24976, N24606, N23071, N18186);
nand NAND3 (N24978, N24970, N17149, N15311);
or OR2 (N24979, N24961, N1513);
buf BUF1 (N24980, N24973);
xor XOR2 (N24981, N24979, N9391);
nor NOR2 (N24982, N24969, N12230);
buf BUF1 (N24983, N24975);
and AND2 (N24984, N24977, N1571);
xor XOR2 (N24985, N24967, N23637);
and AND4 (N24986, N24981, N12499, N13253, N15467);
xor XOR2 (N24987, N24978, N16584);
or OR3 (N24988, N24952, N4321, N12117);
or OR4 (N24989, N24985, N13404, N8189, N14706);
and AND3 (N24990, N24983, N13519, N10190);
or OR3 (N24991, N24987, N15788, N13898);
or OR2 (N24992, N24990, N11770);
nand NAND3 (N24993, N24991, N2559, N10422);
not NOT1 (N24994, N24992);
buf BUF1 (N24995, N24989);
nand NAND4 (N24996, N24993, N5112, N7051, N1430);
buf BUF1 (N24997, N24980);
nand NAND2 (N24998, N24982, N12930);
buf BUF1 (N24999, N24994);
nor NOR2 (N25000, N24971, N11710);
or OR3 (N25001, N24998, N13398, N12219);
buf BUF1 (N25002, N24996);
not NOT1 (N25003, N24986);
not NOT1 (N25004, N24974);
xor XOR2 (N25005, N24999, N9953);
nand NAND4 (N25006, N25004, N13542, N19152, N6859);
buf BUF1 (N25007, N24995);
and AND3 (N25008, N24988, N10093, N15699);
buf BUF1 (N25009, N25002);
buf BUF1 (N25010, N25009);
xor XOR2 (N25011, N25006, N9199);
nand NAND4 (N25012, N25003, N9027, N5531, N14161);
buf BUF1 (N25013, N25007);
and AND4 (N25014, N24997, N8209, N10104, N16401);
nand NAND2 (N25015, N25013, N13918);
or OR2 (N25016, N25012, N7711);
and AND2 (N25017, N25014, N14057);
xor XOR2 (N25018, N25011, N6679);
buf BUF1 (N25019, N25010);
nor NOR3 (N25020, N25008, N18093, N10844);
or OR3 (N25021, N25020, N9486, N19074);
buf BUF1 (N25022, N25001);
nand NAND4 (N25023, N25021, N17980, N10806, N7220);
xor XOR2 (N25024, N25019, N22194);
buf BUF1 (N25025, N25022);
not NOT1 (N25026, N24984);
buf BUF1 (N25027, N25000);
buf BUF1 (N25028, N25025);
and AND4 (N25029, N25026, N12731, N15719, N24394);
and AND2 (N25030, N25005, N19024);
not NOT1 (N25031, N25028);
and AND3 (N25032, N25024, N21987, N59);
nor NOR2 (N25033, N25032, N33);
not NOT1 (N25034, N25031);
and AND2 (N25035, N25033, N19888);
nand NAND4 (N25036, N25030, N17381, N20899, N20557);
not NOT1 (N25037, N25034);
xor XOR2 (N25038, N25027, N16866);
and AND2 (N25039, N25036, N6200);
buf BUF1 (N25040, N25035);
xor XOR2 (N25041, N25017, N15779);
xor XOR2 (N25042, N25023, N8410);
buf BUF1 (N25043, N25016);
xor XOR2 (N25044, N25043, N21745);
nor NOR2 (N25045, N25038, N14750);
buf BUF1 (N25046, N25045);
nand NAND4 (N25047, N25015, N19605, N884, N8447);
and AND4 (N25048, N25041, N7591, N19256, N12992);
not NOT1 (N25049, N25018);
xor XOR2 (N25050, N25039, N15906);
buf BUF1 (N25051, N25042);
xor XOR2 (N25052, N25049, N8865);
not NOT1 (N25053, N25048);
or OR2 (N25054, N25053, N13252);
not NOT1 (N25055, N25029);
nor NOR2 (N25056, N25055, N16578);
xor XOR2 (N25057, N25037, N6468);
buf BUF1 (N25058, N25046);
not NOT1 (N25059, N25044);
and AND3 (N25060, N25050, N2556, N6642);
not NOT1 (N25061, N25040);
not NOT1 (N25062, N25061);
xor XOR2 (N25063, N25062, N14968);
not NOT1 (N25064, N25052);
and AND3 (N25065, N25064, N15813, N6854);
or OR2 (N25066, N25047, N22561);
xor XOR2 (N25067, N25058, N24221);
nor NOR3 (N25068, N25067, N11634, N23210);
and AND3 (N25069, N25056, N11523, N14963);
buf BUF1 (N25070, N25066);
nand NAND2 (N25071, N25069, N24112);
xor XOR2 (N25072, N25068, N20376);
buf BUF1 (N25073, N25060);
or OR2 (N25074, N25070, N13217);
not NOT1 (N25075, N25065);
nor NOR2 (N25076, N25072, N23234);
nand NAND2 (N25077, N25075, N6761);
and AND4 (N25078, N25074, N25030, N18961, N11504);
xor XOR2 (N25079, N25057, N19721);
nand NAND3 (N25080, N25073, N17489, N18182);
or OR3 (N25081, N25051, N21615, N22203);
buf BUF1 (N25082, N25063);
and AND4 (N25083, N25079, N19035, N6798, N6341);
nor NOR4 (N25084, N25078, N20980, N5634, N12596);
xor XOR2 (N25085, N25071, N7603);
nor NOR2 (N25086, N25082, N8671);
not NOT1 (N25087, N25086);
xor XOR2 (N25088, N25080, N13450);
and AND3 (N25089, N25088, N21037, N6267);
nor NOR3 (N25090, N25087, N18783, N15505);
nand NAND4 (N25091, N25054, N17059, N19438, N13333);
nand NAND3 (N25092, N25076, N7911, N6822);
buf BUF1 (N25093, N25059);
or OR4 (N25094, N25085, N24936, N22812, N19690);
nor NOR3 (N25095, N25081, N13642, N10405);
nor NOR3 (N25096, N25091, N16585, N6914);
xor XOR2 (N25097, N25090, N13105);
nor NOR4 (N25098, N25084, N12653, N14436, N14590);
buf BUF1 (N25099, N25089);
nand NAND3 (N25100, N25099, N25047, N25041);
nand NAND2 (N25101, N25093, N23412);
not NOT1 (N25102, N25097);
not NOT1 (N25103, N25101);
nor NOR2 (N25104, N25100, N24040);
nand NAND3 (N25105, N25092, N1802, N9764);
buf BUF1 (N25106, N25077);
xor XOR2 (N25107, N25102, N17436);
and AND3 (N25108, N25103, N17113, N4987);
not NOT1 (N25109, N25083);
nor NOR3 (N25110, N25098, N18103, N24567);
xor XOR2 (N25111, N25095, N17749);
not NOT1 (N25112, N25108);
xor XOR2 (N25113, N25106, N13717);
nor NOR4 (N25114, N25107, N2209, N17278, N12260);
nor NOR2 (N25115, N25105, N20052);
or OR4 (N25116, N25094, N22220, N19802, N23974);
not NOT1 (N25117, N25112);
nor NOR2 (N25118, N25109, N1376);
buf BUF1 (N25119, N25114);
xor XOR2 (N25120, N25116, N17809);
xor XOR2 (N25121, N25120, N5229);
buf BUF1 (N25122, N25110);
nand NAND4 (N25123, N25113, N6605, N2766, N14954);
xor XOR2 (N25124, N25117, N12891);
or OR2 (N25125, N25111, N385);
nand NAND4 (N25126, N25125, N12032, N8746, N15501);
nand NAND2 (N25127, N25119, N18377);
buf BUF1 (N25128, N25115);
not NOT1 (N25129, N25122);
xor XOR2 (N25130, N25127, N10986);
not NOT1 (N25131, N25104);
nor NOR3 (N25132, N25130, N12217, N6073);
or OR2 (N25133, N25118, N12588);
or OR2 (N25134, N25124, N4833);
nor NOR4 (N25135, N25126, N11996, N7720, N13835);
xor XOR2 (N25136, N25123, N15506);
nor NOR3 (N25137, N25121, N3158, N12386);
not NOT1 (N25138, N25096);
buf BUF1 (N25139, N25135);
xor XOR2 (N25140, N25136, N3039);
and AND3 (N25141, N25131, N7608, N22623);
nor NOR3 (N25142, N25138, N606, N22298);
or OR4 (N25143, N25133, N1205, N21543, N6279);
buf BUF1 (N25144, N25140);
nor NOR3 (N25145, N25141, N16206, N10919);
nand NAND3 (N25146, N25143, N2712, N9351);
nor NOR4 (N25147, N25146, N6283, N2613, N6022);
nor NOR4 (N25148, N25139, N6643, N15425, N17487);
buf BUF1 (N25149, N25144);
buf BUF1 (N25150, N25128);
nand NAND3 (N25151, N25137, N21745, N11864);
and AND3 (N25152, N25148, N22394, N17708);
and AND4 (N25153, N25145, N10824, N19671, N16146);
xor XOR2 (N25154, N25149, N15576);
not NOT1 (N25155, N25153);
and AND2 (N25156, N25152, N16992);
nand NAND4 (N25157, N25147, N5514, N9743, N23553);
nand NAND4 (N25158, N25129, N10413, N2905, N14502);
nor NOR4 (N25159, N25151, N6376, N7206, N13810);
nor NOR3 (N25160, N25134, N484, N7328);
buf BUF1 (N25161, N25160);
xor XOR2 (N25162, N25150, N431);
nor NOR2 (N25163, N25161, N7519);
nand NAND2 (N25164, N25163, N11087);
nor NOR2 (N25165, N25132, N14562);
and AND3 (N25166, N25159, N9540, N9133);
or OR4 (N25167, N25142, N20084, N1724, N10885);
not NOT1 (N25168, N25154);
not NOT1 (N25169, N25168);
or OR4 (N25170, N25165, N21324, N15352, N20253);
and AND2 (N25171, N25167, N15418);
not NOT1 (N25172, N25155);
or OR3 (N25173, N25156, N3968, N14548);
buf BUF1 (N25174, N25171);
and AND2 (N25175, N25172, N13651);
or OR3 (N25176, N25166, N24214, N18428);
xor XOR2 (N25177, N25169, N8187);
xor XOR2 (N25178, N25175, N20036);
not NOT1 (N25179, N25158);
nor NOR2 (N25180, N25173, N9497);
buf BUF1 (N25181, N25162);
nor NOR3 (N25182, N25177, N17834, N14472);
nor NOR3 (N25183, N25157, N13764, N20344);
buf BUF1 (N25184, N25182);
or OR3 (N25185, N25178, N3771, N23197);
nor NOR2 (N25186, N25180, N16045);
or OR4 (N25187, N25176, N7111, N22745, N5016);
or OR4 (N25188, N25183, N7885, N14368, N24257);
buf BUF1 (N25189, N25174);
nor NOR3 (N25190, N25187, N10065, N14191);
and AND3 (N25191, N25189, N1524, N8279);
xor XOR2 (N25192, N25170, N6364);
nand NAND3 (N25193, N25190, N9105, N21311);
xor XOR2 (N25194, N25164, N22256);
xor XOR2 (N25195, N25179, N24530);
nand NAND4 (N25196, N25194, N8181, N14091, N2724);
xor XOR2 (N25197, N25188, N20348);
nand NAND3 (N25198, N25195, N14952, N16863);
and AND4 (N25199, N25181, N2109, N9866, N9116);
or OR2 (N25200, N25186, N14044);
xor XOR2 (N25201, N25198, N6241);
buf BUF1 (N25202, N25197);
or OR2 (N25203, N25184, N10609);
and AND4 (N25204, N25191, N6686, N20643, N11740);
not NOT1 (N25205, N25192);
nand NAND4 (N25206, N25201, N6682, N16239, N2941);
not NOT1 (N25207, N25203);
buf BUF1 (N25208, N25202);
not NOT1 (N25209, N25193);
buf BUF1 (N25210, N25209);
nand NAND2 (N25211, N25207, N13973);
xor XOR2 (N25212, N25205, N20160);
nand NAND4 (N25213, N25210, N13137, N23296, N10550);
xor XOR2 (N25214, N25213, N7955);
xor XOR2 (N25215, N25199, N14148);
nand NAND4 (N25216, N25214, N1071, N15743, N80);
not NOT1 (N25217, N25200);
or OR3 (N25218, N25215, N4481, N15338);
or OR2 (N25219, N25211, N19954);
not NOT1 (N25220, N25185);
nand NAND2 (N25221, N25212, N21473);
nor NOR3 (N25222, N25221, N14906, N1559);
buf BUF1 (N25223, N25217);
xor XOR2 (N25224, N25220, N7646);
xor XOR2 (N25225, N25216, N13997);
nand NAND2 (N25226, N25222, N17492);
nor NOR4 (N25227, N25219, N24047, N23490, N1899);
or OR2 (N25228, N25206, N20706);
or OR3 (N25229, N25218, N17254, N8850);
nor NOR2 (N25230, N25227, N20508);
and AND2 (N25231, N25228, N10090);
nand NAND4 (N25232, N25223, N10863, N23280, N9940);
nor NOR2 (N25233, N25196, N5640);
nor NOR3 (N25234, N25208, N10465, N21045);
not NOT1 (N25235, N25204);
or OR4 (N25236, N25229, N4761, N11629, N6368);
buf BUF1 (N25237, N25234);
not NOT1 (N25238, N25235);
not NOT1 (N25239, N25231);
xor XOR2 (N25240, N25237, N10356);
buf BUF1 (N25241, N25226);
buf BUF1 (N25242, N25233);
nand NAND2 (N25243, N25225, N13987);
or OR3 (N25244, N25230, N3542, N173);
nor NOR3 (N25245, N25239, N9482, N13698);
xor XOR2 (N25246, N25236, N1207);
xor XOR2 (N25247, N25224, N15361);
and AND2 (N25248, N25232, N18674);
or OR4 (N25249, N25243, N15618, N5647, N71);
nand NAND3 (N25250, N25249, N1374, N4471);
or OR3 (N25251, N25244, N8148, N19240);
and AND3 (N25252, N25247, N25111, N21189);
xor XOR2 (N25253, N25252, N169);
not NOT1 (N25254, N25240);
nor NOR2 (N25255, N25242, N9693);
xor XOR2 (N25256, N25245, N9860);
nor NOR4 (N25257, N25253, N13523, N19519, N17096);
and AND2 (N25258, N25246, N15257);
nand NAND2 (N25259, N25254, N6955);
xor XOR2 (N25260, N25251, N7282);
or OR3 (N25261, N25250, N18069, N24511);
nand NAND4 (N25262, N25248, N436, N22006, N25138);
nand NAND3 (N25263, N25255, N5194, N15474);
and AND3 (N25264, N25259, N18867, N11770);
and AND3 (N25265, N25263, N5313, N8870);
xor XOR2 (N25266, N25265, N17959);
xor XOR2 (N25267, N25266, N8765);
nor NOR3 (N25268, N25264, N15849, N12977);
nor NOR2 (N25269, N25238, N17822);
not NOT1 (N25270, N25262);
nor NOR2 (N25271, N25241, N23604);
nand NAND3 (N25272, N25267, N12589, N23041);
nor NOR2 (N25273, N25268, N23442);
not NOT1 (N25274, N25271);
or OR3 (N25275, N25261, N2661, N13225);
not NOT1 (N25276, N25272);
xor XOR2 (N25277, N25275, N6921);
nand NAND2 (N25278, N25277, N18888);
nand NAND4 (N25279, N25278, N2541, N7856, N13110);
buf BUF1 (N25280, N25256);
nor NOR3 (N25281, N25257, N4319, N4855);
nor NOR3 (N25282, N25274, N18751, N3089);
buf BUF1 (N25283, N25258);
buf BUF1 (N25284, N25270);
and AND3 (N25285, N25276, N18805, N1503);
and AND4 (N25286, N25273, N12352, N22501, N22294);
and AND3 (N25287, N25281, N15478, N24687);
or OR3 (N25288, N25286, N4731, N23750);
or OR4 (N25289, N25283, N11231, N22345, N24969);
not NOT1 (N25290, N25285);
or OR3 (N25291, N25282, N21576, N10353);
nand NAND3 (N25292, N25279, N2705, N12839);
buf BUF1 (N25293, N25287);
nor NOR3 (N25294, N25289, N13446, N2131);
or OR3 (N25295, N25290, N8052, N18148);
nand NAND4 (N25296, N25294, N3873, N15462, N737);
or OR3 (N25297, N25291, N582, N17269);
and AND2 (N25298, N25269, N21626);
nand NAND3 (N25299, N25288, N1259, N11425);
or OR3 (N25300, N25284, N1291, N18880);
not NOT1 (N25301, N25293);
or OR2 (N25302, N25280, N16303);
or OR2 (N25303, N25301, N16924);
nor NOR3 (N25304, N25260, N14353, N7179);
nand NAND3 (N25305, N25296, N9438, N10157);
nand NAND3 (N25306, N25292, N7519, N20792);
buf BUF1 (N25307, N25297);
and AND3 (N25308, N25305, N18066, N17569);
buf BUF1 (N25309, N25295);
xor XOR2 (N25310, N25308, N22186);
and AND2 (N25311, N25307, N18213);
xor XOR2 (N25312, N25300, N14688);
nor NOR2 (N25313, N25306, N7263);
nor NOR2 (N25314, N25309, N132);
xor XOR2 (N25315, N25314, N25015);
nor NOR4 (N25316, N25311, N21702, N8084, N21820);
and AND4 (N25317, N25313, N17975, N18886, N2888);
and AND2 (N25318, N25298, N6639);
not NOT1 (N25319, N25304);
nor NOR2 (N25320, N25319, N11691);
or OR4 (N25321, N25303, N22006, N1415, N8098);
nor NOR3 (N25322, N25312, N24768, N12988);
or OR4 (N25323, N25315, N19985, N24792, N18795);
or OR2 (N25324, N25310, N2536);
or OR2 (N25325, N25324, N24228);
buf BUF1 (N25326, N25322);
not NOT1 (N25327, N25321);
nand NAND2 (N25328, N25316, N1817);
nor NOR2 (N25329, N25317, N17027);
nor NOR3 (N25330, N25299, N12351, N14658);
or OR3 (N25331, N25327, N2170, N20755);
or OR2 (N25332, N25329, N12193);
xor XOR2 (N25333, N25326, N6632);
or OR2 (N25334, N25323, N9218);
nand NAND4 (N25335, N25318, N4369, N21884, N17627);
buf BUF1 (N25336, N25335);
or OR3 (N25337, N25331, N3898, N13278);
buf BUF1 (N25338, N25330);
not NOT1 (N25339, N25328);
xor XOR2 (N25340, N25337, N8900);
nand NAND2 (N25341, N25302, N9525);
buf BUF1 (N25342, N25338);
and AND4 (N25343, N25341, N18340, N4243, N6609);
nand NAND3 (N25344, N25325, N12728, N13799);
nor NOR3 (N25345, N25342, N18350, N19819);
nor NOR4 (N25346, N25334, N11782, N21876, N23277);
not NOT1 (N25347, N25343);
nand NAND4 (N25348, N25332, N6955, N6653, N20694);
xor XOR2 (N25349, N25344, N4091);
nor NOR3 (N25350, N25346, N24135, N9615);
and AND4 (N25351, N25348, N22795, N14101, N6598);
and AND2 (N25352, N25347, N9164);
xor XOR2 (N25353, N25340, N11622);
or OR3 (N25354, N25351, N7785, N21913);
and AND2 (N25355, N25352, N15372);
not NOT1 (N25356, N25339);
or OR4 (N25357, N25333, N11295, N8503, N6301);
xor XOR2 (N25358, N25354, N10711);
buf BUF1 (N25359, N25336);
xor XOR2 (N25360, N25353, N15324);
buf BUF1 (N25361, N25345);
not NOT1 (N25362, N25358);
nand NAND2 (N25363, N25359, N20347);
nor NOR2 (N25364, N25320, N16167);
and AND4 (N25365, N25350, N5779, N2317, N18649);
buf BUF1 (N25366, N25355);
nand NAND4 (N25367, N25365, N4946, N15518, N19908);
xor XOR2 (N25368, N25356, N5755);
and AND3 (N25369, N25357, N4207, N25173);
or OR2 (N25370, N25366, N23202);
nand NAND3 (N25371, N25360, N4113, N20244);
xor XOR2 (N25372, N25364, N18125);
not NOT1 (N25373, N25363);
or OR2 (N25374, N25367, N4594);
nor NOR2 (N25375, N25373, N311);
or OR3 (N25376, N25370, N8039, N1908);
not NOT1 (N25377, N25361);
nor NOR4 (N25378, N25377, N9070, N24817, N23153);
or OR3 (N25379, N25378, N23034, N20513);
xor XOR2 (N25380, N25362, N7581);
nor NOR4 (N25381, N25369, N7769, N10855, N15557);
nor NOR4 (N25382, N25374, N6200, N15373, N14485);
and AND4 (N25383, N25380, N14951, N274, N14594);
buf BUF1 (N25384, N25383);
not NOT1 (N25385, N25379);
nor NOR4 (N25386, N25371, N5304, N1859, N12625);
nand NAND4 (N25387, N25385, N13458, N15073, N19622);
or OR3 (N25388, N25376, N6262, N1451);
nand NAND3 (N25389, N25388, N23471, N1418);
or OR3 (N25390, N25382, N18561, N24966);
xor XOR2 (N25391, N25384, N22359);
or OR3 (N25392, N25381, N23319, N5111);
xor XOR2 (N25393, N25389, N8218);
not NOT1 (N25394, N25391);
nand NAND2 (N25395, N25394, N5056);
xor XOR2 (N25396, N25387, N15038);
nand NAND3 (N25397, N25393, N16, N10161);
nor NOR2 (N25398, N25375, N975);
buf BUF1 (N25399, N25386);
buf BUF1 (N25400, N25397);
nand NAND4 (N25401, N25396, N1702, N14103, N13126);
not NOT1 (N25402, N25398);
nand NAND2 (N25403, N25368, N23874);
xor XOR2 (N25404, N25392, N22063);
not NOT1 (N25405, N25400);
xor XOR2 (N25406, N25403, N19273);
not NOT1 (N25407, N25401);
or OR2 (N25408, N25390, N17781);
and AND4 (N25409, N25349, N20385, N1701, N16770);
or OR3 (N25410, N25405, N23416, N20849);
nand NAND3 (N25411, N25407, N3168, N24587);
xor XOR2 (N25412, N25406, N18448);
or OR4 (N25413, N25372, N14797, N2680, N24460);
and AND3 (N25414, N25409, N15768, N20437);
not NOT1 (N25415, N25399);
or OR2 (N25416, N25408, N21972);
or OR2 (N25417, N25412, N5781);
or OR4 (N25418, N25415, N8281, N15498, N25416);
nand NAND2 (N25419, N22652, N2868);
or OR3 (N25420, N25402, N15056, N3652);
nand NAND2 (N25421, N25411, N7178);
xor XOR2 (N25422, N25410, N4475);
buf BUF1 (N25423, N25413);
buf BUF1 (N25424, N25423);
or OR3 (N25425, N25419, N3255, N3457);
nor NOR4 (N25426, N25425, N385, N5957, N4084);
buf BUF1 (N25427, N25417);
xor XOR2 (N25428, N25414, N7050);
not NOT1 (N25429, N25424);
buf BUF1 (N25430, N25395);
buf BUF1 (N25431, N25418);
not NOT1 (N25432, N25426);
nand NAND3 (N25433, N25431, N5347, N14742);
buf BUF1 (N25434, N25404);
xor XOR2 (N25435, N25422, N1714);
buf BUF1 (N25436, N25430);
buf BUF1 (N25437, N25420);
or OR4 (N25438, N25421, N15256, N994, N10543);
not NOT1 (N25439, N25435);
or OR2 (N25440, N25436, N19489);
not NOT1 (N25441, N25434);
and AND3 (N25442, N25440, N10446, N22376);
buf BUF1 (N25443, N25441);
nor NOR4 (N25444, N25428, N23682, N13378, N8736);
xor XOR2 (N25445, N25438, N23545);
xor XOR2 (N25446, N25427, N24766);
buf BUF1 (N25447, N25439);
not NOT1 (N25448, N25437);
not NOT1 (N25449, N25447);
not NOT1 (N25450, N25445);
not NOT1 (N25451, N25446);
xor XOR2 (N25452, N25433, N19861);
nor NOR4 (N25453, N25450, N10321, N1132, N22596);
buf BUF1 (N25454, N25452);
not NOT1 (N25455, N25429);
and AND4 (N25456, N25455, N980, N11388, N22444);
and AND4 (N25457, N25456, N17006, N15865, N15485);
and AND4 (N25458, N25457, N5626, N20318, N17502);
nor NOR3 (N25459, N25451, N2333, N19882);
xor XOR2 (N25460, N25448, N12312);
not NOT1 (N25461, N25442);
nand NAND3 (N25462, N25443, N19943, N3835);
and AND2 (N25463, N25432, N19246);
not NOT1 (N25464, N25458);
not NOT1 (N25465, N25449);
xor XOR2 (N25466, N25454, N2970);
nor NOR3 (N25467, N25464, N12137, N1645);
or OR3 (N25468, N25453, N10532, N13115);
nor NOR2 (N25469, N25467, N20710);
nor NOR2 (N25470, N25466, N16297);
and AND4 (N25471, N25460, N12103, N23967, N25341);
nor NOR4 (N25472, N25462, N9030, N25147, N7101);
xor XOR2 (N25473, N25471, N16549);
nor NOR4 (N25474, N25461, N16293, N2964, N14524);
xor XOR2 (N25475, N25473, N9682);
buf BUF1 (N25476, N25474);
xor XOR2 (N25477, N25472, N5817);
not NOT1 (N25478, N25465);
and AND2 (N25479, N25478, N9076);
or OR2 (N25480, N25477, N22469);
nor NOR4 (N25481, N25459, N19386, N7325, N13756);
nor NOR4 (N25482, N25479, N18740, N7632, N19940);
or OR4 (N25483, N25481, N21907, N3491, N16529);
not NOT1 (N25484, N25444);
xor XOR2 (N25485, N25463, N13726);
nand NAND4 (N25486, N25483, N5484, N2108, N21288);
nand NAND2 (N25487, N25476, N8809);
nor NOR4 (N25488, N25468, N9543, N10564, N6542);
not NOT1 (N25489, N25470);
buf BUF1 (N25490, N25484);
and AND3 (N25491, N25488, N19577, N23879);
buf BUF1 (N25492, N25475);
nor NOR4 (N25493, N25485, N14573, N18488, N8801);
buf BUF1 (N25494, N25490);
xor XOR2 (N25495, N25482, N25411);
buf BUF1 (N25496, N25489);
nor NOR4 (N25497, N25492, N1659, N18952, N11397);
and AND4 (N25498, N25469, N931, N9882, N8298);
not NOT1 (N25499, N25497);
xor XOR2 (N25500, N25486, N7857);
xor XOR2 (N25501, N25499, N24242);
nand NAND2 (N25502, N25494, N551);
not NOT1 (N25503, N25501);
buf BUF1 (N25504, N25487);
buf BUF1 (N25505, N25493);
and AND3 (N25506, N25480, N22966, N25490);
buf BUF1 (N25507, N25496);
buf BUF1 (N25508, N25491);
not NOT1 (N25509, N25502);
nor NOR3 (N25510, N25509, N8742, N1214);
not NOT1 (N25511, N25498);
and AND2 (N25512, N25510, N17485);
nor NOR3 (N25513, N25503, N23917, N398);
and AND2 (N25514, N25511, N11607);
xor XOR2 (N25515, N25506, N11092);
xor XOR2 (N25516, N25514, N5111);
and AND3 (N25517, N25500, N22710, N14204);
not NOT1 (N25518, N25505);
nand NAND3 (N25519, N25495, N16457, N22872);
nor NOR4 (N25520, N25512, N6767, N1040, N5974);
nand NAND3 (N25521, N25519, N9165, N22084);
nand NAND2 (N25522, N25515, N24870);
and AND2 (N25523, N25516, N5338);
not NOT1 (N25524, N25521);
xor XOR2 (N25525, N25520, N7089);
and AND2 (N25526, N25524, N23334);
nand NAND2 (N25527, N25523, N5377);
and AND4 (N25528, N25508, N5630, N13261, N9098);
nand NAND2 (N25529, N25526, N9053);
xor XOR2 (N25530, N25527, N16327);
xor XOR2 (N25531, N25528, N18556);
nand NAND2 (N25532, N25530, N9019);
xor XOR2 (N25533, N25531, N9100);
or OR4 (N25534, N25533, N15871, N7132, N20606);
nor NOR2 (N25535, N25507, N14159);
and AND3 (N25536, N25532, N4648, N13677);
nand NAND4 (N25537, N25525, N22236, N14465, N1504);
and AND2 (N25538, N25536, N16025);
nor NOR2 (N25539, N25538, N21294);
or OR3 (N25540, N25535, N10897, N12321);
nand NAND2 (N25541, N25518, N8880);
nand NAND3 (N25542, N25513, N12503, N3222);
and AND2 (N25543, N25522, N17308);
not NOT1 (N25544, N25534);
xor XOR2 (N25545, N25529, N10586);
buf BUF1 (N25546, N25543);
buf BUF1 (N25547, N25539);
or OR3 (N25548, N25544, N12861, N3789);
and AND4 (N25549, N25545, N24972, N25006, N7800);
buf BUF1 (N25550, N25547);
and AND2 (N25551, N25504, N10828);
xor XOR2 (N25552, N25546, N1855);
xor XOR2 (N25553, N25548, N22659);
not NOT1 (N25554, N25551);
nor NOR4 (N25555, N25549, N10665, N18766, N13606);
not NOT1 (N25556, N25552);
or OR4 (N25557, N25550, N22692, N9736, N16787);
buf BUF1 (N25558, N25540);
nor NOR2 (N25559, N25558, N7251);
or OR3 (N25560, N25537, N4611, N1003);
nand NAND3 (N25561, N25541, N2426, N18978);
xor XOR2 (N25562, N25555, N5904);
or OR3 (N25563, N25542, N18210, N5140);
and AND2 (N25564, N25517, N12068);
buf BUF1 (N25565, N25553);
not NOT1 (N25566, N25554);
xor XOR2 (N25567, N25562, N2836);
xor XOR2 (N25568, N25565, N15110);
xor XOR2 (N25569, N25560, N3676);
and AND4 (N25570, N25563, N7462, N14429, N16333);
and AND3 (N25571, N25567, N6055, N9696);
nor NOR3 (N25572, N25564, N4833, N13832);
nor NOR2 (N25573, N25556, N8290);
nor NOR2 (N25574, N25566, N12935);
or OR3 (N25575, N25573, N16736, N14641);
and AND4 (N25576, N25569, N7831, N16221, N23943);
or OR3 (N25577, N25576, N20548, N21629);
not NOT1 (N25578, N25572);
xor XOR2 (N25579, N25574, N24311);
xor XOR2 (N25580, N25559, N13120);
not NOT1 (N25581, N25575);
nand NAND4 (N25582, N25561, N8723, N23155, N5796);
xor XOR2 (N25583, N25577, N9949);
not NOT1 (N25584, N25568);
nor NOR3 (N25585, N25584, N15151, N18797);
buf BUF1 (N25586, N25570);
nor NOR2 (N25587, N25578, N24825);
not NOT1 (N25588, N25583);
buf BUF1 (N25589, N25582);
xor XOR2 (N25590, N25581, N7536);
buf BUF1 (N25591, N25580);
or OR4 (N25592, N25589, N6672, N5339, N8472);
nand NAND2 (N25593, N25591, N20462);
nor NOR3 (N25594, N25590, N8911, N2035);
xor XOR2 (N25595, N25579, N19929);
or OR2 (N25596, N25587, N6030);
nor NOR4 (N25597, N25586, N23107, N8040, N5126);
and AND4 (N25598, N25557, N11271, N20246, N20294);
nand NAND3 (N25599, N25598, N4311, N14903);
and AND2 (N25600, N25596, N5182);
buf BUF1 (N25601, N25592);
and AND3 (N25602, N25600, N4242, N20840);
nand NAND4 (N25603, N25601, N21058, N12846, N23702);
xor XOR2 (N25604, N25585, N23286);
xor XOR2 (N25605, N25597, N16389);
xor XOR2 (N25606, N25603, N4646);
nor NOR3 (N25607, N25593, N14816, N24952);
not NOT1 (N25608, N25605);
nor NOR2 (N25609, N25571, N4200);
nand NAND2 (N25610, N25599, N18914);
and AND4 (N25611, N25606, N12520, N3190, N24480);
not NOT1 (N25612, N25588);
not NOT1 (N25613, N25594);
not NOT1 (N25614, N25602);
not NOT1 (N25615, N25610);
and AND3 (N25616, N25609, N17933, N8922);
not NOT1 (N25617, N25612);
not NOT1 (N25618, N25615);
nor NOR2 (N25619, N25614, N14126);
or OR4 (N25620, N25613, N7585, N18467, N16851);
endmodule