// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N3013,N3018,N2996,N2983,N3015,N3008,N3017,N3014,N3002,N3019;

and AND4 (N20, N5, N10, N16, N12);
nand NAND4 (N21, N5, N11, N9, N6);
not NOT1 (N22, N9);
nor NOR2 (N23, N6, N12);
xor XOR2 (N24, N13, N18);
and AND4 (N25, N2, N16, N17, N3);
nor NOR4 (N26, N21, N22, N6, N5);
nand NAND2 (N27, N22, N21);
not NOT1 (N28, N8);
nand NAND2 (N29, N25, N8);
and AND3 (N30, N5, N23, N28);
xor XOR2 (N31, N25, N12);
xor XOR2 (N32, N31, N7);
nor NOR3 (N33, N7, N3, N28);
nor NOR3 (N34, N14, N16, N1);
nor NOR4 (N35, N5, N6, N33, N17);
and AND3 (N36, N17, N19, N21);
buf BUF1 (N37, N32);
nand NAND2 (N38, N26, N24);
xor XOR2 (N39, N35, N36);
xor XOR2 (N40, N11, N18);
xor XOR2 (N41, N6, N30);
not NOT1 (N42, N25);
buf BUF1 (N43, N41);
xor XOR2 (N44, N34, N16);
nand NAND2 (N45, N42, N8);
and AND2 (N46, N29, N32);
not NOT1 (N47, N40);
or OR2 (N48, N27, N27);
xor XOR2 (N49, N37, N41);
nand NAND4 (N50, N39, N1, N33, N38);
or OR3 (N51, N8, N24, N37);
nand NAND3 (N52, N44, N46, N43);
not NOT1 (N53, N7);
buf BUF1 (N54, N13);
nand NAND4 (N55, N54, N25, N36, N46);
xor XOR2 (N56, N53, N50);
and AND4 (N57, N15, N32, N19, N16);
nand NAND3 (N58, N57, N7, N30);
or OR4 (N59, N20, N44, N40, N36);
not NOT1 (N60, N49);
xor XOR2 (N61, N56, N36);
or OR4 (N62, N45, N38, N31, N29);
not NOT1 (N63, N52);
buf BUF1 (N64, N61);
not NOT1 (N65, N62);
nand NAND2 (N66, N58, N34);
and AND3 (N67, N66, N46, N19);
or OR3 (N68, N47, N64, N65);
xor XOR2 (N69, N37, N50);
not NOT1 (N70, N68);
or OR4 (N71, N21, N59, N36, N54);
nand NAND2 (N72, N58, N36);
nor NOR4 (N73, N63, N52, N66, N22);
xor XOR2 (N74, N71, N49);
and AND4 (N75, N70, N25, N70, N7);
and AND2 (N76, N73, N46);
buf BUF1 (N77, N74);
xor XOR2 (N78, N67, N33);
not NOT1 (N79, N69);
and AND3 (N80, N75, N27, N35);
or OR3 (N81, N48, N44, N44);
or OR2 (N82, N72, N27);
or OR3 (N83, N76, N69, N61);
nand NAND2 (N84, N83, N40);
buf BUF1 (N85, N60);
nor NOR2 (N86, N84, N43);
and AND4 (N87, N86, N6, N86, N78);
nor NOR3 (N88, N83, N22, N40);
not NOT1 (N89, N79);
xor XOR2 (N90, N51, N84);
or OR4 (N91, N77, N69, N5, N5);
not NOT1 (N92, N87);
not NOT1 (N93, N88);
nor NOR3 (N94, N92, N67, N86);
nand NAND3 (N95, N94, N2, N92);
and AND2 (N96, N90, N87);
xor XOR2 (N97, N91, N6);
buf BUF1 (N98, N93);
or OR3 (N99, N97, N45, N25);
and AND4 (N100, N99, N1, N23, N53);
nor NOR4 (N101, N100, N8, N46, N15);
nor NOR4 (N102, N82, N35, N20, N64);
nor NOR3 (N103, N102, N32, N97);
buf BUF1 (N104, N89);
and AND3 (N105, N103, N13, N13);
nor NOR3 (N106, N96, N13, N88);
or OR2 (N107, N106, N78);
nand NAND2 (N108, N81, N76);
xor XOR2 (N109, N85, N67);
xor XOR2 (N110, N108, N60);
nand NAND2 (N111, N95, N62);
not NOT1 (N112, N107);
or OR2 (N113, N98, N56);
xor XOR2 (N114, N80, N83);
nand NAND3 (N115, N114, N1, N66);
and AND4 (N116, N115, N27, N113, N109);
nor NOR3 (N117, N70, N57, N6);
buf BUF1 (N118, N24);
or OR4 (N119, N110, N87, N117, N58);
nand NAND2 (N120, N1, N30);
not NOT1 (N121, N104);
and AND4 (N122, N121, N29, N81, N78);
nor NOR4 (N123, N105, N86, N16, N107);
and AND4 (N124, N112, N55, N25, N102);
nand NAND3 (N125, N69, N17, N81);
and AND3 (N126, N101, N8, N58);
nand NAND3 (N127, N123, N26, N72);
not NOT1 (N128, N116);
nand NAND3 (N129, N128, N83, N110);
or OR2 (N130, N118, N8);
nand NAND3 (N131, N111, N105, N35);
buf BUF1 (N132, N131);
nand NAND2 (N133, N122, N64);
or OR3 (N134, N120, N109, N97);
buf BUF1 (N135, N127);
nand NAND3 (N136, N125, N18, N2);
nor NOR2 (N137, N126, N84);
not NOT1 (N138, N124);
nand NAND2 (N139, N133, N61);
not NOT1 (N140, N130);
xor XOR2 (N141, N134, N58);
and AND4 (N142, N129, N67, N106, N117);
or OR2 (N143, N141, N69);
buf BUF1 (N144, N140);
not NOT1 (N145, N132);
not NOT1 (N146, N137);
buf BUF1 (N147, N143);
not NOT1 (N148, N145);
or OR4 (N149, N144, N128, N134, N106);
or OR2 (N150, N135, N130);
buf BUF1 (N151, N136);
or OR4 (N152, N147, N42, N28, N14);
nor NOR3 (N153, N148, N71, N23);
or OR3 (N154, N146, N78, N55);
and AND3 (N155, N150, N106, N92);
not NOT1 (N156, N152);
nand NAND3 (N157, N119, N111, N153);
or OR2 (N158, N1, N35);
xor XOR2 (N159, N151, N66);
xor XOR2 (N160, N157, N84);
buf BUF1 (N161, N156);
nand NAND2 (N162, N138, N156);
nor NOR2 (N163, N162, N67);
not NOT1 (N164, N163);
and AND3 (N165, N142, N70, N8);
nor NOR2 (N166, N161, N155);
buf BUF1 (N167, N78);
and AND4 (N168, N154, N66, N129, N148);
or OR4 (N169, N160, N58, N128, N156);
buf BUF1 (N170, N169);
and AND2 (N171, N170, N90);
or OR3 (N172, N139, N114, N42);
xor XOR2 (N173, N165, N127);
nand NAND4 (N174, N167, N47, N22, N93);
nor NOR3 (N175, N168, N112, N155);
and AND2 (N176, N174, N116);
nor NOR2 (N177, N171, N21);
nand NAND3 (N178, N158, N135, N169);
buf BUF1 (N179, N178);
nor NOR2 (N180, N149, N119);
buf BUF1 (N181, N176);
nor NOR3 (N182, N177, N95, N70);
or OR2 (N183, N173, N130);
and AND4 (N184, N179, N77, N113, N66);
xor XOR2 (N185, N159, N7);
xor XOR2 (N186, N164, N146);
and AND4 (N187, N182, N40, N140, N123);
or OR2 (N188, N172, N130);
nor NOR3 (N189, N181, N77, N63);
buf BUF1 (N190, N189);
buf BUF1 (N191, N166);
xor XOR2 (N192, N187, N50);
xor XOR2 (N193, N186, N81);
not NOT1 (N194, N175);
not NOT1 (N195, N188);
nand NAND4 (N196, N195, N74, N27, N147);
nand NAND3 (N197, N184, N160, N17);
nor NOR2 (N198, N180, N114);
nand NAND2 (N199, N190, N48);
and AND4 (N200, N199, N104, N187, N47);
or OR4 (N201, N185, N37, N155, N34);
not NOT1 (N202, N183);
and AND2 (N203, N192, N64);
and AND2 (N204, N197, N122);
nand NAND4 (N205, N196, N73, N44, N146);
and AND2 (N206, N205, N42);
not NOT1 (N207, N193);
nand NAND2 (N208, N200, N184);
buf BUF1 (N209, N207);
not NOT1 (N210, N206);
nand NAND3 (N211, N208, N104, N82);
nand NAND4 (N212, N211, N93, N179, N55);
or OR3 (N213, N204, N127, N57);
nand NAND3 (N214, N194, N165, N173);
nor NOR2 (N215, N209, N82);
and AND3 (N216, N198, N100, N99);
nor NOR3 (N217, N216, N213, N17);
buf BUF1 (N218, N178);
nor NOR2 (N219, N210, N180);
or OR3 (N220, N218, N197, N143);
xor XOR2 (N221, N202, N208);
not NOT1 (N222, N203);
and AND4 (N223, N201, N91, N95, N94);
and AND2 (N224, N220, N114);
nand NAND4 (N225, N217, N81, N199, N209);
xor XOR2 (N226, N223, N51);
nand NAND4 (N227, N215, N184, N225, N73);
not NOT1 (N228, N116);
nor NOR2 (N229, N226, N65);
buf BUF1 (N230, N214);
or OR2 (N231, N191, N58);
not NOT1 (N232, N219);
and AND3 (N233, N222, N225, N35);
nand NAND4 (N234, N227, N130, N43, N75);
and AND3 (N235, N224, N31, N102);
and AND4 (N236, N221, N137, N231, N26);
not NOT1 (N237, N57);
nand NAND3 (N238, N229, N228, N63);
or OR4 (N239, N9, N231, N49, N233);
and AND2 (N240, N63, N146);
buf BUF1 (N241, N238);
not NOT1 (N242, N239);
xor XOR2 (N243, N212, N33);
nand NAND3 (N244, N242, N188, N118);
buf BUF1 (N245, N230);
buf BUF1 (N246, N232);
nor NOR2 (N247, N243, N14);
nand NAND2 (N248, N244, N85);
and AND3 (N249, N236, N61, N100);
or OR2 (N250, N249, N219);
or OR4 (N251, N234, N215, N241, N135);
nand NAND3 (N252, N105, N90, N99);
buf BUF1 (N253, N237);
xor XOR2 (N254, N235, N104);
buf BUF1 (N255, N240);
or OR2 (N256, N250, N218);
or OR4 (N257, N256, N5, N32, N80);
nand NAND3 (N258, N253, N169, N94);
and AND2 (N259, N251, N147);
xor XOR2 (N260, N248, N29);
buf BUF1 (N261, N254);
or OR3 (N262, N246, N99, N257);
buf BUF1 (N263, N71);
xor XOR2 (N264, N255, N108);
not NOT1 (N265, N245);
nand NAND4 (N266, N265, N265, N195, N216);
or OR3 (N267, N258, N142, N120);
not NOT1 (N268, N266);
not NOT1 (N269, N268);
nor NOR2 (N270, N264, N269);
xor XOR2 (N271, N156, N253);
nor NOR2 (N272, N247, N6);
nand NAND2 (N273, N259, N102);
buf BUF1 (N274, N270);
xor XOR2 (N275, N262, N56);
buf BUF1 (N276, N267);
xor XOR2 (N277, N271, N261);
nand NAND3 (N278, N106, N220, N131);
and AND3 (N279, N276, N136, N225);
or OR3 (N280, N275, N162, N129);
or OR4 (N281, N280, N166, N48, N76);
or OR4 (N282, N279, N47, N164, N37);
nor NOR2 (N283, N263, N9);
xor XOR2 (N284, N283, N121);
or OR3 (N285, N252, N77, N161);
not NOT1 (N286, N282);
nand NAND3 (N287, N284, N116, N24);
and AND2 (N288, N260, N29);
and AND4 (N289, N274, N142, N191, N260);
not NOT1 (N290, N281);
buf BUF1 (N291, N290);
xor XOR2 (N292, N277, N140);
buf BUF1 (N293, N287);
xor XOR2 (N294, N288, N150);
or OR4 (N295, N272, N237, N33, N162);
buf BUF1 (N296, N293);
buf BUF1 (N297, N286);
or OR4 (N298, N295, N249, N76, N115);
nor NOR4 (N299, N289, N206, N41, N186);
not NOT1 (N300, N273);
xor XOR2 (N301, N296, N277);
and AND4 (N302, N299, N107, N73, N267);
buf BUF1 (N303, N297);
not NOT1 (N304, N303);
and AND2 (N305, N294, N285);
and AND2 (N306, N118, N167);
and AND2 (N307, N298, N89);
or OR2 (N308, N306, N155);
nor NOR3 (N309, N305, N267, N11);
buf BUF1 (N310, N309);
and AND4 (N311, N304, N213, N230, N290);
nand NAND2 (N312, N291, N47);
or OR4 (N313, N312, N116, N240, N220);
or OR4 (N314, N292, N179, N202, N35);
nand NAND4 (N315, N278, N169, N211, N198);
buf BUF1 (N316, N300);
xor XOR2 (N317, N315, N121);
xor XOR2 (N318, N311, N38);
xor XOR2 (N319, N307, N163);
and AND3 (N320, N319, N14, N217);
and AND4 (N321, N316, N159, N131, N106);
nand NAND2 (N322, N318, N292);
not NOT1 (N323, N317);
and AND3 (N324, N323, N124, N218);
xor XOR2 (N325, N314, N118);
not NOT1 (N326, N324);
nand NAND4 (N327, N302, N171, N186, N5);
or OR2 (N328, N327, N211);
or OR3 (N329, N308, N33, N161);
nor NOR3 (N330, N325, N288, N12);
and AND3 (N331, N329, N232, N151);
buf BUF1 (N332, N310);
buf BUF1 (N333, N322);
or OR2 (N334, N313, N288);
and AND3 (N335, N321, N178, N17);
buf BUF1 (N336, N334);
and AND2 (N337, N328, N326);
nand NAND4 (N338, N68, N219, N331, N149);
nor NOR3 (N339, N248, N294, N50);
nand NAND4 (N340, N337, N141, N163, N211);
and AND3 (N341, N335, N84, N140);
or OR3 (N342, N330, N27, N313);
nand NAND2 (N343, N340, N145);
nor NOR4 (N344, N343, N269, N73, N73);
not NOT1 (N345, N336);
not NOT1 (N346, N333);
nand NAND2 (N347, N346, N322);
xor XOR2 (N348, N345, N66);
xor XOR2 (N349, N332, N101);
or OR3 (N350, N339, N210, N87);
buf BUF1 (N351, N347);
not NOT1 (N352, N342);
or OR4 (N353, N351, N119, N52, N38);
or OR2 (N354, N341, N190);
buf BUF1 (N355, N301);
and AND3 (N356, N349, N246, N231);
xor XOR2 (N357, N348, N340);
nor NOR2 (N358, N344, N258);
nor NOR3 (N359, N358, N35, N187);
xor XOR2 (N360, N353, N91);
not NOT1 (N361, N357);
or OR2 (N362, N355, N295);
buf BUF1 (N363, N360);
nor NOR2 (N364, N350, N134);
and AND3 (N365, N359, N344, N318);
nor NOR3 (N366, N320, N110, N94);
and AND3 (N367, N354, N44, N67);
and AND3 (N368, N363, N73, N101);
xor XOR2 (N369, N352, N259);
xor XOR2 (N370, N366, N317);
nor NOR4 (N371, N369, N315, N237, N259);
xor XOR2 (N372, N370, N216);
nand NAND3 (N373, N372, N268, N192);
xor XOR2 (N374, N356, N13);
not NOT1 (N375, N367);
buf BUF1 (N376, N361);
or OR3 (N377, N375, N216, N360);
buf BUF1 (N378, N373);
not NOT1 (N379, N377);
or OR2 (N380, N338, N201);
buf BUF1 (N381, N380);
nand NAND2 (N382, N374, N99);
buf BUF1 (N383, N365);
nand NAND4 (N384, N381, N40, N163, N13);
buf BUF1 (N385, N384);
nor NOR3 (N386, N383, N17, N137);
and AND3 (N387, N378, N365, N66);
and AND4 (N388, N379, N186, N344, N57);
buf BUF1 (N389, N368);
nand NAND2 (N390, N387, N234);
not NOT1 (N391, N386);
and AND3 (N392, N376, N97, N350);
nor NOR4 (N393, N371, N136, N213, N317);
buf BUF1 (N394, N392);
not NOT1 (N395, N364);
nor NOR4 (N396, N395, N281, N167, N240);
or OR2 (N397, N362, N259);
and AND2 (N398, N394, N193);
and AND3 (N399, N397, N39, N20);
xor XOR2 (N400, N393, N160);
buf BUF1 (N401, N398);
nand NAND3 (N402, N382, N134, N328);
or OR4 (N403, N402, N145, N34, N24);
buf BUF1 (N404, N400);
buf BUF1 (N405, N391);
and AND4 (N406, N389, N134, N267, N292);
buf BUF1 (N407, N401);
xor XOR2 (N408, N403, N106);
or OR2 (N409, N388, N54);
or OR4 (N410, N385, N188, N92, N90);
not NOT1 (N411, N408);
xor XOR2 (N412, N404, N113);
or OR3 (N413, N396, N229, N348);
nand NAND2 (N414, N409, N115);
xor XOR2 (N415, N412, N289);
or OR4 (N416, N406, N150, N46, N143);
xor XOR2 (N417, N413, N34);
and AND2 (N418, N415, N308);
and AND2 (N419, N417, N17);
buf BUF1 (N420, N416);
xor XOR2 (N421, N390, N98);
or OR4 (N422, N421, N179, N200, N356);
xor XOR2 (N423, N420, N108);
or OR2 (N424, N399, N368);
or OR3 (N425, N414, N423, N274);
or OR2 (N426, N6, N17);
not NOT1 (N427, N422);
and AND2 (N428, N418, N327);
xor XOR2 (N429, N411, N168);
or OR3 (N430, N425, N355, N352);
and AND4 (N431, N424, N416, N377, N358);
xor XOR2 (N432, N426, N38);
not NOT1 (N433, N419);
buf BUF1 (N434, N407);
nor NOR3 (N435, N434, N109, N125);
nor NOR2 (N436, N431, N266);
or OR3 (N437, N405, N353, N28);
and AND2 (N438, N437, N244);
nor NOR2 (N439, N433, N245);
and AND4 (N440, N439, N340, N52, N166);
and AND2 (N441, N428, N251);
buf BUF1 (N442, N441);
nand NAND2 (N443, N410, N9);
xor XOR2 (N444, N435, N152);
nor NOR4 (N445, N443, N306, N266, N148);
xor XOR2 (N446, N442, N170);
nor NOR4 (N447, N440, N181, N29, N311);
not NOT1 (N448, N446);
or OR3 (N449, N448, N409, N264);
nand NAND4 (N450, N445, N127, N21, N332);
not NOT1 (N451, N438);
nand NAND2 (N452, N427, N288);
buf BUF1 (N453, N450);
and AND2 (N454, N447, N246);
or OR3 (N455, N430, N159, N218);
buf BUF1 (N456, N451);
not NOT1 (N457, N449);
and AND2 (N458, N452, N142);
buf BUF1 (N459, N454);
nor NOR4 (N460, N459, N6, N52, N378);
or OR4 (N461, N436, N235, N233, N97);
or OR3 (N462, N453, N206, N60);
buf BUF1 (N463, N458);
xor XOR2 (N464, N463, N297);
buf BUF1 (N465, N460);
not NOT1 (N466, N464);
or OR4 (N467, N456, N449, N452, N255);
or OR3 (N468, N429, N331, N383);
buf BUF1 (N469, N457);
buf BUF1 (N470, N469);
and AND2 (N471, N465, N5);
and AND3 (N472, N444, N26, N437);
or OR4 (N473, N461, N70, N402, N452);
not NOT1 (N474, N473);
nor NOR2 (N475, N471, N62);
not NOT1 (N476, N475);
nor NOR2 (N477, N462, N437);
nand NAND2 (N478, N470, N108);
buf BUF1 (N479, N478);
not NOT1 (N480, N455);
and AND3 (N481, N480, N414, N389);
xor XOR2 (N482, N477, N263);
not NOT1 (N483, N472);
or OR2 (N484, N481, N71);
not NOT1 (N485, N474);
nand NAND2 (N486, N479, N74);
not NOT1 (N487, N483);
nand NAND3 (N488, N466, N171, N105);
buf BUF1 (N489, N468);
not NOT1 (N490, N484);
nor NOR4 (N491, N432, N222, N355, N458);
nand NAND2 (N492, N467, N347);
or OR2 (N493, N482, N395);
and AND4 (N494, N488, N397, N353, N293);
xor XOR2 (N495, N490, N118);
xor XOR2 (N496, N476, N355);
xor XOR2 (N497, N491, N243);
or OR2 (N498, N497, N417);
nor NOR2 (N499, N486, N8);
and AND3 (N500, N487, N52, N328);
xor XOR2 (N501, N493, N102);
or OR3 (N502, N496, N205, N177);
buf BUF1 (N503, N489);
xor XOR2 (N504, N498, N494);
xor XOR2 (N505, N210, N137);
nand NAND3 (N506, N492, N130, N49);
nand NAND3 (N507, N495, N500, N303);
or OR4 (N508, N92, N93, N366, N232);
xor XOR2 (N509, N503, N207);
or OR2 (N510, N504, N18);
xor XOR2 (N511, N510, N319);
not NOT1 (N512, N501);
xor XOR2 (N513, N512, N292);
or OR4 (N514, N513, N494, N493, N281);
not NOT1 (N515, N507);
or OR3 (N516, N511, N324, N158);
or OR3 (N517, N505, N265, N138);
not NOT1 (N518, N508);
not NOT1 (N519, N516);
nor NOR3 (N520, N514, N293, N386);
buf BUF1 (N521, N506);
not NOT1 (N522, N485);
nand NAND4 (N523, N502, N280, N281, N268);
or OR3 (N524, N522, N266, N404);
buf BUF1 (N525, N519);
and AND3 (N526, N499, N196, N275);
xor XOR2 (N527, N525, N204);
and AND2 (N528, N521, N301);
nor NOR4 (N529, N526, N102, N209, N440);
nor NOR2 (N530, N529, N116);
not NOT1 (N531, N530);
not NOT1 (N532, N524);
nor NOR4 (N533, N520, N298, N391, N489);
not NOT1 (N534, N527);
or OR4 (N535, N533, N227, N393, N176);
buf BUF1 (N536, N515);
and AND3 (N537, N535, N532, N39);
nor NOR3 (N538, N367, N162, N27);
and AND2 (N539, N518, N82);
xor XOR2 (N540, N523, N94);
buf BUF1 (N541, N537);
nor NOR2 (N542, N538, N480);
or OR4 (N543, N531, N480, N247, N48);
nand NAND3 (N544, N539, N427, N77);
xor XOR2 (N545, N517, N255);
not NOT1 (N546, N543);
xor XOR2 (N547, N534, N205);
nand NAND3 (N548, N546, N43, N436);
and AND3 (N549, N548, N373, N417);
and AND3 (N550, N509, N149, N25);
or OR4 (N551, N540, N473, N24, N483);
not NOT1 (N552, N542);
buf BUF1 (N553, N545);
or OR4 (N554, N550, N347, N80, N330);
or OR2 (N555, N554, N147);
or OR3 (N556, N544, N266, N185);
or OR2 (N557, N553, N287);
or OR2 (N558, N528, N424);
nor NOR3 (N559, N536, N493, N282);
xor XOR2 (N560, N559, N224);
nand NAND3 (N561, N552, N548, N63);
nand NAND4 (N562, N541, N49, N530, N68);
and AND3 (N563, N562, N166, N279);
not NOT1 (N564, N556);
not NOT1 (N565, N555);
buf BUF1 (N566, N557);
or OR2 (N567, N549, N340);
or OR4 (N568, N565, N497, N58, N141);
nand NAND2 (N569, N566, N510);
nand NAND4 (N570, N558, N163, N196, N273);
xor XOR2 (N571, N568, N413);
nor NOR2 (N572, N571, N174);
buf BUF1 (N573, N551);
nand NAND4 (N574, N561, N45, N410, N267);
and AND3 (N575, N564, N94, N497);
and AND2 (N576, N570, N137);
buf BUF1 (N577, N563);
nand NAND4 (N578, N567, N187, N104, N409);
and AND3 (N579, N577, N66, N219);
or OR2 (N580, N579, N530);
not NOT1 (N581, N547);
nand NAND3 (N582, N569, N19, N30);
nor NOR3 (N583, N575, N141, N541);
buf BUF1 (N584, N574);
not NOT1 (N585, N572);
nor NOR4 (N586, N578, N290, N418, N293);
xor XOR2 (N587, N582, N339);
not NOT1 (N588, N583);
xor XOR2 (N589, N581, N100);
nor NOR3 (N590, N585, N551, N489);
nor NOR4 (N591, N580, N142, N582, N97);
and AND2 (N592, N560, N422);
nor NOR3 (N593, N587, N313, N390);
buf BUF1 (N594, N591);
nor NOR4 (N595, N589, N13, N405, N267);
or OR2 (N596, N584, N569);
not NOT1 (N597, N595);
and AND2 (N598, N573, N491);
not NOT1 (N599, N586);
or OR4 (N600, N590, N397, N407, N10);
not NOT1 (N601, N594);
xor XOR2 (N602, N598, N407);
or OR4 (N603, N599, N32, N88, N417);
buf BUF1 (N604, N600);
not NOT1 (N605, N576);
buf BUF1 (N606, N602);
nand NAND4 (N607, N593, N416, N466, N234);
nand NAND2 (N608, N592, N450);
buf BUF1 (N609, N606);
and AND4 (N610, N597, N565, N569, N563);
xor XOR2 (N611, N596, N286);
xor XOR2 (N612, N605, N549);
and AND2 (N613, N603, N370);
and AND2 (N614, N612, N202);
and AND3 (N615, N614, N356, N168);
nor NOR3 (N616, N601, N50, N8);
xor XOR2 (N617, N607, N298);
and AND4 (N618, N616, N420, N6, N508);
and AND4 (N619, N604, N603, N408, N23);
xor XOR2 (N620, N588, N264);
buf BUF1 (N621, N615);
buf BUF1 (N622, N609);
nand NAND3 (N623, N611, N359, N528);
nor NOR2 (N624, N621, N162);
not NOT1 (N625, N622);
or OR2 (N626, N613, N244);
buf BUF1 (N627, N608);
xor XOR2 (N628, N626, N102);
and AND2 (N629, N610, N325);
nor NOR2 (N630, N629, N373);
nor NOR2 (N631, N620, N3);
buf BUF1 (N632, N630);
or OR4 (N633, N628, N172, N424, N123);
nand NAND4 (N634, N633, N314, N477, N205);
xor XOR2 (N635, N634, N376);
or OR4 (N636, N617, N575, N570, N581);
nand NAND2 (N637, N625, N86);
buf BUF1 (N638, N627);
nor NOR3 (N639, N623, N630, N385);
nor NOR3 (N640, N636, N302, N377);
nor NOR4 (N641, N618, N620, N456, N117);
nand NAND3 (N642, N641, N73, N248);
not NOT1 (N643, N640);
not NOT1 (N644, N631);
nand NAND4 (N645, N643, N591, N108, N38);
and AND2 (N646, N639, N313);
xor XOR2 (N647, N638, N588);
and AND2 (N648, N637, N48);
and AND2 (N649, N647, N117);
nand NAND2 (N650, N635, N323);
or OR4 (N651, N632, N278, N578, N101);
and AND2 (N652, N651, N584);
not NOT1 (N653, N619);
not NOT1 (N654, N642);
and AND4 (N655, N644, N455, N200, N417);
not NOT1 (N656, N653);
buf BUF1 (N657, N652);
or OR4 (N658, N649, N580, N268, N442);
buf BUF1 (N659, N654);
nor NOR2 (N660, N657, N576);
and AND2 (N661, N655, N608);
xor XOR2 (N662, N660, N635);
nand NAND4 (N663, N646, N52, N31, N613);
or OR3 (N664, N645, N476, N593);
buf BUF1 (N665, N662);
xor XOR2 (N666, N624, N124);
not NOT1 (N667, N658);
buf BUF1 (N668, N661);
xor XOR2 (N669, N656, N381);
and AND3 (N670, N667, N600, N659);
nor NOR2 (N671, N208, N407);
nor NOR3 (N672, N665, N160, N568);
not NOT1 (N673, N669);
buf BUF1 (N674, N671);
nand NAND3 (N675, N650, N368, N308);
xor XOR2 (N676, N670, N582);
nand NAND2 (N677, N674, N653);
buf BUF1 (N678, N663);
nand NAND3 (N679, N677, N585, N200);
nand NAND3 (N680, N664, N117, N309);
buf BUF1 (N681, N668);
nor NOR2 (N682, N680, N281);
nand NAND4 (N683, N678, N669, N295, N651);
and AND3 (N684, N679, N163, N18);
buf BUF1 (N685, N673);
nor NOR4 (N686, N684, N16, N504, N427);
nor NOR2 (N687, N681, N340);
and AND3 (N688, N648, N602, N35);
not NOT1 (N689, N685);
nand NAND3 (N690, N688, N545, N90);
buf BUF1 (N691, N686);
not NOT1 (N692, N675);
nor NOR4 (N693, N666, N381, N661, N674);
nor NOR4 (N694, N693, N320, N665, N658);
nor NOR3 (N695, N694, N302, N276);
buf BUF1 (N696, N683);
buf BUF1 (N697, N687);
nor NOR2 (N698, N691, N516);
or OR4 (N699, N689, N363, N294, N486);
nand NAND4 (N700, N698, N558, N88, N424);
and AND3 (N701, N695, N499, N171);
xor XOR2 (N702, N697, N337);
not NOT1 (N703, N700);
nor NOR3 (N704, N701, N149, N530);
not NOT1 (N705, N676);
not NOT1 (N706, N702);
or OR3 (N707, N703, N151, N411);
buf BUF1 (N708, N682);
buf BUF1 (N709, N708);
not NOT1 (N710, N699);
xor XOR2 (N711, N709, N699);
nand NAND3 (N712, N696, N608, N387);
nor NOR3 (N713, N710, N191, N262);
nand NAND3 (N714, N704, N463, N10);
or OR2 (N715, N711, N423);
nor NOR3 (N716, N713, N673, N311);
nand NAND3 (N717, N714, N65, N60);
or OR3 (N718, N690, N107, N436);
or OR3 (N719, N707, N493, N602);
nand NAND3 (N720, N718, N325, N509);
buf BUF1 (N721, N706);
xor XOR2 (N722, N716, N203);
or OR2 (N723, N672, N620);
nand NAND4 (N724, N712, N363, N505, N278);
and AND4 (N725, N722, N89, N265, N548);
nor NOR4 (N726, N724, N51, N124, N442);
or OR3 (N727, N725, N397, N125);
or OR4 (N728, N692, N505, N258, N179);
nand NAND4 (N729, N728, N153, N558, N140);
and AND3 (N730, N717, N342, N692);
xor XOR2 (N731, N721, N245);
nor NOR2 (N732, N726, N179);
buf BUF1 (N733, N719);
or OR3 (N734, N733, N620, N451);
nand NAND4 (N735, N727, N480, N294, N300);
or OR3 (N736, N730, N358, N360);
buf BUF1 (N737, N731);
buf BUF1 (N738, N715);
nand NAND2 (N739, N723, N192);
buf BUF1 (N740, N738);
or OR4 (N741, N737, N592, N369, N690);
xor XOR2 (N742, N705, N118);
buf BUF1 (N743, N740);
nor NOR2 (N744, N735, N283);
nor NOR4 (N745, N742, N46, N458, N91);
nor NOR2 (N746, N734, N77);
xor XOR2 (N747, N739, N329);
xor XOR2 (N748, N746, N468);
nor NOR2 (N749, N729, N446);
buf BUF1 (N750, N732);
buf BUF1 (N751, N748);
and AND4 (N752, N741, N47, N711, N133);
xor XOR2 (N753, N751, N652);
nand NAND2 (N754, N750, N179);
xor XOR2 (N755, N749, N508);
or OR4 (N756, N754, N742, N615, N688);
xor XOR2 (N757, N745, N695);
not NOT1 (N758, N720);
buf BUF1 (N759, N752);
nor NOR2 (N760, N743, N339);
not NOT1 (N761, N760);
and AND4 (N762, N753, N322, N550, N146);
nand NAND4 (N763, N755, N47, N459, N370);
buf BUF1 (N764, N744);
nand NAND3 (N765, N736, N468, N412);
and AND3 (N766, N756, N112, N587);
nor NOR2 (N767, N762, N636);
nand NAND3 (N768, N757, N494, N341);
buf BUF1 (N769, N747);
or OR3 (N770, N763, N739, N682);
and AND2 (N771, N766, N757);
not NOT1 (N772, N769);
nor NOR2 (N773, N761, N233);
buf BUF1 (N774, N759);
not NOT1 (N775, N767);
nor NOR4 (N776, N772, N737, N241, N114);
and AND2 (N777, N775, N509);
and AND2 (N778, N776, N536);
nand NAND4 (N779, N764, N103, N61, N185);
xor XOR2 (N780, N758, N717);
and AND3 (N781, N774, N207, N482);
nand NAND4 (N782, N771, N427, N203, N489);
and AND4 (N783, N765, N1, N216, N63);
nor NOR4 (N784, N778, N643, N39, N288);
buf BUF1 (N785, N773);
or OR4 (N786, N781, N188, N157, N688);
not NOT1 (N787, N782);
xor XOR2 (N788, N768, N121);
not NOT1 (N789, N770);
nand NAND2 (N790, N783, N169);
not NOT1 (N791, N787);
not NOT1 (N792, N790);
xor XOR2 (N793, N780, N203);
xor XOR2 (N794, N786, N767);
and AND3 (N795, N785, N72, N575);
and AND4 (N796, N789, N260, N88, N736);
and AND4 (N797, N777, N789, N262, N417);
not NOT1 (N798, N794);
nor NOR3 (N799, N788, N229, N25);
nor NOR2 (N800, N792, N329);
xor XOR2 (N801, N798, N217);
nor NOR3 (N802, N784, N330, N406);
buf BUF1 (N803, N801);
or OR3 (N804, N797, N521, N495);
buf BUF1 (N805, N779);
and AND2 (N806, N802, N187);
nor NOR3 (N807, N799, N114, N42);
xor XOR2 (N808, N803, N727);
nand NAND3 (N809, N796, N8, N46);
or OR3 (N810, N807, N802, N103);
or OR4 (N811, N804, N603, N278, N104);
and AND4 (N812, N809, N533, N208, N286);
buf BUF1 (N813, N811);
and AND3 (N814, N805, N26, N316);
nand NAND4 (N815, N791, N297, N298, N154);
nor NOR3 (N816, N793, N365, N670);
xor XOR2 (N817, N815, N277);
not NOT1 (N818, N806);
xor XOR2 (N819, N817, N170);
not NOT1 (N820, N816);
nor NOR3 (N821, N800, N780, N748);
xor XOR2 (N822, N818, N559);
buf BUF1 (N823, N821);
nand NAND2 (N824, N808, N278);
xor XOR2 (N825, N810, N743);
or OR3 (N826, N795, N368, N141);
and AND2 (N827, N814, N174);
or OR4 (N828, N824, N621, N815, N404);
nand NAND2 (N829, N825, N470);
nor NOR2 (N830, N826, N379);
buf BUF1 (N831, N829);
or OR2 (N832, N823, N772);
buf BUF1 (N833, N812);
nor NOR3 (N834, N822, N462, N38);
not NOT1 (N835, N820);
nand NAND4 (N836, N830, N727, N592, N370);
nor NOR4 (N837, N828, N316, N270, N815);
nand NAND4 (N838, N833, N392, N718, N510);
nand NAND4 (N839, N819, N4, N481, N589);
and AND4 (N840, N831, N459, N240, N24);
nor NOR2 (N841, N827, N100);
not NOT1 (N842, N835);
not NOT1 (N843, N836);
not NOT1 (N844, N838);
or OR2 (N845, N841, N273);
nand NAND2 (N846, N844, N392);
buf BUF1 (N847, N839);
buf BUF1 (N848, N845);
not NOT1 (N849, N832);
xor XOR2 (N850, N847, N157);
not NOT1 (N851, N848);
nor NOR4 (N852, N849, N566, N350, N840);
xor XOR2 (N853, N57, N193);
nor NOR4 (N854, N834, N183, N415, N121);
xor XOR2 (N855, N854, N663);
nor NOR2 (N856, N813, N600);
buf BUF1 (N857, N851);
nand NAND3 (N858, N852, N512, N659);
not NOT1 (N859, N842);
not NOT1 (N860, N858);
buf BUF1 (N861, N859);
nand NAND2 (N862, N853, N271);
or OR4 (N863, N860, N126, N537, N485);
and AND2 (N864, N846, N751);
nand NAND4 (N865, N855, N203, N114, N640);
nand NAND4 (N866, N863, N813, N531, N541);
nand NAND2 (N867, N837, N443);
not NOT1 (N868, N856);
not NOT1 (N869, N861);
nand NAND4 (N870, N866, N457, N748, N603);
and AND3 (N871, N864, N714, N109);
nor NOR3 (N872, N862, N292, N7);
buf BUF1 (N873, N872);
xor XOR2 (N874, N867, N401);
xor XOR2 (N875, N843, N691);
not NOT1 (N876, N874);
buf BUF1 (N877, N870);
nor NOR2 (N878, N873, N52);
buf BUF1 (N879, N871);
xor XOR2 (N880, N878, N222);
not NOT1 (N881, N879);
not NOT1 (N882, N880);
or OR4 (N883, N857, N786, N537, N420);
not NOT1 (N884, N875);
nor NOR2 (N885, N882, N673);
buf BUF1 (N886, N884);
and AND4 (N887, N886, N325, N232, N195);
xor XOR2 (N888, N868, N274);
xor XOR2 (N889, N881, N366);
and AND2 (N890, N889, N228);
nor NOR2 (N891, N890, N487);
and AND4 (N892, N850, N268, N486, N626);
or OR2 (N893, N891, N519);
and AND3 (N894, N893, N302, N772);
buf BUF1 (N895, N885);
buf BUF1 (N896, N894);
nand NAND2 (N897, N876, N696);
xor XOR2 (N898, N897, N60);
buf BUF1 (N899, N898);
nand NAND4 (N900, N892, N250, N787, N39);
nor NOR3 (N901, N888, N699, N83);
nand NAND4 (N902, N887, N329, N879, N514);
nand NAND4 (N903, N902, N524, N596, N274);
xor XOR2 (N904, N896, N852);
and AND3 (N905, N877, N144, N782);
or OR3 (N906, N901, N104, N44);
not NOT1 (N907, N906);
or OR2 (N908, N869, N41);
xor XOR2 (N909, N907, N161);
nor NOR4 (N910, N903, N270, N389, N115);
not NOT1 (N911, N865);
buf BUF1 (N912, N905);
and AND2 (N913, N900, N371);
nor NOR2 (N914, N908, N274);
xor XOR2 (N915, N911, N183);
or OR2 (N916, N909, N868);
nand NAND3 (N917, N914, N505, N591);
not NOT1 (N918, N904);
buf BUF1 (N919, N918);
or OR3 (N920, N910, N171, N139);
or OR4 (N921, N917, N250, N162, N761);
nand NAND4 (N922, N912, N888, N263, N63);
nand NAND4 (N923, N919, N61, N641, N813);
xor XOR2 (N924, N920, N20);
or OR2 (N925, N915, N275);
nand NAND4 (N926, N921, N450, N165, N607);
nand NAND3 (N927, N895, N551, N883);
or OR3 (N928, N12, N326, N546);
xor XOR2 (N929, N924, N698);
nand NAND3 (N930, N927, N564, N121);
nor NOR3 (N931, N928, N364, N533);
xor XOR2 (N932, N931, N294);
and AND4 (N933, N923, N714, N791, N475);
buf BUF1 (N934, N899);
buf BUF1 (N935, N930);
xor XOR2 (N936, N935, N519);
not NOT1 (N937, N933);
not NOT1 (N938, N926);
xor XOR2 (N939, N922, N420);
not NOT1 (N940, N938);
or OR3 (N941, N934, N627, N473);
or OR3 (N942, N936, N498, N683);
xor XOR2 (N943, N913, N676);
and AND2 (N944, N925, N76);
nor NOR3 (N945, N939, N111, N148);
xor XOR2 (N946, N941, N767);
nand NAND2 (N947, N945, N904);
and AND2 (N948, N932, N78);
not NOT1 (N949, N942);
buf BUF1 (N950, N940);
buf BUF1 (N951, N916);
nor NOR4 (N952, N937, N770, N71, N778);
nand NAND4 (N953, N943, N197, N942, N464);
and AND4 (N954, N950, N949, N792, N416);
xor XOR2 (N955, N949, N167);
nand NAND4 (N956, N948, N286, N544, N188);
or OR4 (N957, N947, N626, N284, N906);
not NOT1 (N958, N946);
nor NOR4 (N959, N956, N320, N636, N743);
or OR4 (N960, N951, N72, N610, N40);
or OR2 (N961, N957, N67);
nand NAND3 (N962, N961, N492, N277);
xor XOR2 (N963, N962, N545);
nor NOR3 (N964, N954, N603, N434);
or OR4 (N965, N963, N164, N676, N251);
nand NAND3 (N966, N960, N816, N444);
nand NAND2 (N967, N965, N679);
or OR3 (N968, N967, N663, N373);
nor NOR3 (N969, N968, N624, N515);
xor XOR2 (N970, N969, N767);
not NOT1 (N971, N966);
or OR4 (N972, N964, N624, N707, N421);
not NOT1 (N973, N929);
or OR4 (N974, N973, N686, N179, N891);
or OR3 (N975, N974, N523, N481);
xor XOR2 (N976, N955, N733);
and AND4 (N977, N975, N603, N33, N400);
nor NOR4 (N978, N976, N527, N528, N480);
xor XOR2 (N979, N952, N415);
nand NAND2 (N980, N958, N951);
or OR2 (N981, N944, N578);
nand NAND3 (N982, N980, N624, N762);
and AND4 (N983, N978, N324, N428, N402);
and AND3 (N984, N971, N140, N294);
not NOT1 (N985, N983);
nor NOR4 (N986, N981, N281, N399, N536);
not NOT1 (N987, N982);
buf BUF1 (N988, N970);
and AND4 (N989, N986, N746, N384, N181);
and AND4 (N990, N987, N495, N414, N975);
xor XOR2 (N991, N989, N729);
xor XOR2 (N992, N990, N189);
xor XOR2 (N993, N992, N609);
and AND2 (N994, N979, N748);
and AND3 (N995, N988, N2, N806);
or OR4 (N996, N953, N57, N284, N914);
not NOT1 (N997, N985);
not NOT1 (N998, N959);
nor NOR4 (N999, N997, N356, N107, N549);
or OR3 (N1000, N995, N144, N61);
and AND3 (N1001, N991, N8, N641);
xor XOR2 (N1002, N972, N407);
nand NAND3 (N1003, N999, N55, N915);
nand NAND2 (N1004, N984, N423);
nor NOR2 (N1005, N977, N237);
nor NOR3 (N1006, N998, N40, N451);
nor NOR2 (N1007, N1005, N682);
buf BUF1 (N1008, N1002);
and AND3 (N1009, N996, N394, N269);
xor XOR2 (N1010, N1009, N421);
xor XOR2 (N1011, N1000, N995);
not NOT1 (N1012, N1001);
nand NAND2 (N1013, N1006, N101);
not NOT1 (N1014, N1010);
buf BUF1 (N1015, N1013);
not NOT1 (N1016, N1014);
buf BUF1 (N1017, N1015);
buf BUF1 (N1018, N1016);
nand NAND4 (N1019, N1004, N874, N609, N56);
not NOT1 (N1020, N1007);
not NOT1 (N1021, N1011);
nor NOR3 (N1022, N1019, N1001, N738);
and AND3 (N1023, N1012, N579, N127);
xor XOR2 (N1024, N1017, N892);
nand NAND2 (N1025, N1018, N936);
xor XOR2 (N1026, N1021, N430);
or OR3 (N1027, N1023, N204, N218);
xor XOR2 (N1028, N1025, N598);
xor XOR2 (N1029, N1022, N175);
not NOT1 (N1030, N1029);
or OR3 (N1031, N993, N38, N831);
buf BUF1 (N1032, N1031);
not NOT1 (N1033, N1024);
or OR3 (N1034, N994, N437, N718);
nor NOR4 (N1035, N1026, N791, N1024, N95);
nand NAND4 (N1036, N1003, N412, N228, N756);
nor NOR2 (N1037, N1035, N320);
buf BUF1 (N1038, N1032);
and AND3 (N1039, N1034, N963, N185);
not NOT1 (N1040, N1008);
and AND3 (N1041, N1020, N283, N235);
not NOT1 (N1042, N1033);
nor NOR3 (N1043, N1039, N742, N535);
xor XOR2 (N1044, N1038, N564);
not NOT1 (N1045, N1028);
nor NOR3 (N1046, N1045, N636, N282);
and AND2 (N1047, N1040, N333);
not NOT1 (N1048, N1042);
not NOT1 (N1049, N1027);
buf BUF1 (N1050, N1046);
and AND2 (N1051, N1036, N175);
and AND4 (N1052, N1041, N154, N77, N945);
nor NOR2 (N1053, N1049, N658);
not NOT1 (N1054, N1044);
nand NAND3 (N1055, N1053, N165, N412);
or OR3 (N1056, N1054, N735, N968);
xor XOR2 (N1057, N1047, N480);
not NOT1 (N1058, N1052);
buf BUF1 (N1059, N1055);
nor NOR2 (N1060, N1037, N474);
and AND3 (N1061, N1050, N953, N141);
buf BUF1 (N1062, N1060);
or OR3 (N1063, N1043, N226, N674);
nand NAND4 (N1064, N1063, N300, N839, N363);
not NOT1 (N1065, N1058);
xor XOR2 (N1066, N1057, N845);
or OR2 (N1067, N1064, N1039);
not NOT1 (N1068, N1030);
nor NOR4 (N1069, N1048, N558, N1059, N204);
nand NAND3 (N1070, N167, N335, N266);
nand NAND4 (N1071, N1056, N564, N560, N847);
buf BUF1 (N1072, N1061);
nand NAND2 (N1073, N1066, N534);
nand NAND2 (N1074, N1067, N849);
or OR3 (N1075, N1072, N1018, N83);
xor XOR2 (N1076, N1071, N814);
nand NAND2 (N1077, N1073, N254);
buf BUF1 (N1078, N1069);
or OR4 (N1079, N1076, N624, N667, N438);
nand NAND3 (N1080, N1079, N692, N1055);
and AND3 (N1081, N1078, N147, N66);
nand NAND3 (N1082, N1062, N197, N1071);
nand NAND2 (N1083, N1070, N416);
and AND4 (N1084, N1074, N267, N1007, N624);
buf BUF1 (N1085, N1081);
xor XOR2 (N1086, N1084, N694);
and AND3 (N1087, N1082, N270, N370);
nor NOR2 (N1088, N1075, N206);
nand NAND4 (N1089, N1086, N336, N875, N231);
nand NAND2 (N1090, N1068, N459);
buf BUF1 (N1091, N1051);
buf BUF1 (N1092, N1090);
and AND3 (N1093, N1080, N1073, N923);
not NOT1 (N1094, N1088);
xor XOR2 (N1095, N1094, N154);
and AND2 (N1096, N1083, N163);
nand NAND3 (N1097, N1089, N539, N389);
nor NOR4 (N1098, N1087, N521, N1076, N468);
and AND2 (N1099, N1091, N290);
or OR2 (N1100, N1097, N132);
buf BUF1 (N1101, N1099);
or OR3 (N1102, N1095, N314, N370);
and AND3 (N1103, N1065, N578, N748);
nand NAND2 (N1104, N1101, N289);
and AND3 (N1105, N1093, N974, N193);
not NOT1 (N1106, N1103);
and AND3 (N1107, N1106, N894, N683);
buf BUF1 (N1108, N1092);
nor NOR4 (N1109, N1102, N1021, N1045, N193);
not NOT1 (N1110, N1096);
and AND2 (N1111, N1104, N652);
buf BUF1 (N1112, N1110);
nor NOR2 (N1113, N1107, N840);
xor XOR2 (N1114, N1077, N371);
or OR2 (N1115, N1098, N295);
nand NAND3 (N1116, N1113, N1016, N483);
nor NOR4 (N1117, N1100, N128, N458, N567);
or OR3 (N1118, N1111, N11, N764);
nand NAND3 (N1119, N1116, N412, N393);
not NOT1 (N1120, N1109);
buf BUF1 (N1121, N1117);
nor NOR3 (N1122, N1108, N969, N508);
nor NOR3 (N1123, N1122, N544, N358);
not NOT1 (N1124, N1105);
buf BUF1 (N1125, N1121);
or OR2 (N1126, N1119, N891);
nand NAND2 (N1127, N1126, N486);
nor NOR3 (N1128, N1114, N960, N191);
not NOT1 (N1129, N1128);
buf BUF1 (N1130, N1125);
nand NAND2 (N1131, N1115, N700);
xor XOR2 (N1132, N1118, N519);
buf BUF1 (N1133, N1130);
and AND3 (N1134, N1112, N790, N682);
or OR2 (N1135, N1131, N742);
or OR4 (N1136, N1134, N606, N338, N443);
nor NOR3 (N1137, N1136, N385, N663);
buf BUF1 (N1138, N1132);
nor NOR2 (N1139, N1127, N456);
and AND3 (N1140, N1124, N42, N1075);
buf BUF1 (N1141, N1120);
nor NOR2 (N1142, N1085, N86);
nor NOR4 (N1143, N1133, N1045, N148, N376);
xor XOR2 (N1144, N1140, N127);
or OR3 (N1145, N1123, N501, N222);
not NOT1 (N1146, N1139);
buf BUF1 (N1147, N1137);
nor NOR4 (N1148, N1144, N735, N725, N548);
buf BUF1 (N1149, N1147);
xor XOR2 (N1150, N1148, N1139);
buf BUF1 (N1151, N1150);
buf BUF1 (N1152, N1145);
and AND4 (N1153, N1146, N832, N331, N677);
or OR4 (N1154, N1152, N847, N336, N995);
or OR4 (N1155, N1154, N529, N253, N1028);
buf BUF1 (N1156, N1138);
not NOT1 (N1157, N1155);
not NOT1 (N1158, N1135);
or OR3 (N1159, N1129, N112, N421);
xor XOR2 (N1160, N1158, N577);
nand NAND2 (N1161, N1160, N1015);
nor NOR2 (N1162, N1153, N497);
buf BUF1 (N1163, N1151);
or OR3 (N1164, N1156, N1154, N1107);
or OR3 (N1165, N1143, N66, N561);
or OR4 (N1166, N1164, N315, N627, N1128);
nor NOR4 (N1167, N1166, N19, N1096, N397);
nand NAND4 (N1168, N1167, N846, N36, N628);
buf BUF1 (N1169, N1161);
not NOT1 (N1170, N1149);
or OR4 (N1171, N1163, N224, N350, N553);
or OR2 (N1172, N1171, N125);
buf BUF1 (N1173, N1157);
not NOT1 (N1174, N1168);
and AND2 (N1175, N1170, N253);
buf BUF1 (N1176, N1162);
nand NAND4 (N1177, N1173, N203, N205, N2);
nor NOR3 (N1178, N1165, N113, N1120);
and AND2 (N1179, N1176, N539);
buf BUF1 (N1180, N1142);
not NOT1 (N1181, N1178);
nand NAND3 (N1182, N1175, N691, N790);
not NOT1 (N1183, N1181);
xor XOR2 (N1184, N1174, N544);
xor XOR2 (N1185, N1177, N458);
buf BUF1 (N1186, N1183);
and AND4 (N1187, N1169, N440, N535, N331);
nand NAND3 (N1188, N1186, N1133, N126);
and AND2 (N1189, N1187, N978);
and AND3 (N1190, N1159, N780, N149);
nand NAND2 (N1191, N1182, N573);
buf BUF1 (N1192, N1141);
and AND2 (N1193, N1189, N162);
buf BUF1 (N1194, N1192);
and AND2 (N1195, N1179, N464);
or OR3 (N1196, N1180, N558, N1051);
xor XOR2 (N1197, N1184, N1008);
xor XOR2 (N1198, N1190, N779);
buf BUF1 (N1199, N1193);
not NOT1 (N1200, N1188);
not NOT1 (N1201, N1185);
and AND4 (N1202, N1198, N558, N114, N911);
buf BUF1 (N1203, N1200);
or OR2 (N1204, N1197, N89);
nor NOR3 (N1205, N1203, N75, N860);
nand NAND2 (N1206, N1202, N226);
xor XOR2 (N1207, N1196, N1132);
buf BUF1 (N1208, N1195);
nor NOR4 (N1209, N1206, N878, N559, N231);
nor NOR2 (N1210, N1208, N773);
buf BUF1 (N1211, N1194);
not NOT1 (N1212, N1207);
nand NAND2 (N1213, N1210, N1024);
nor NOR2 (N1214, N1204, N698);
and AND4 (N1215, N1213, N413, N1103, N402);
not NOT1 (N1216, N1172);
xor XOR2 (N1217, N1211, N655);
xor XOR2 (N1218, N1217, N152);
and AND3 (N1219, N1201, N222, N515);
and AND3 (N1220, N1216, N713, N740);
not NOT1 (N1221, N1215);
or OR2 (N1222, N1205, N963);
buf BUF1 (N1223, N1212);
and AND3 (N1224, N1209, N560, N406);
nor NOR4 (N1225, N1191, N839, N928, N1192);
buf BUF1 (N1226, N1223);
not NOT1 (N1227, N1221);
not NOT1 (N1228, N1227);
and AND3 (N1229, N1219, N490, N550);
buf BUF1 (N1230, N1228);
and AND2 (N1231, N1220, N1034);
xor XOR2 (N1232, N1230, N677);
or OR3 (N1233, N1199, N48, N293);
buf BUF1 (N1234, N1214);
xor XOR2 (N1235, N1234, N685);
or OR2 (N1236, N1222, N722);
nor NOR3 (N1237, N1225, N401, N859);
or OR4 (N1238, N1229, N1223, N1012, N616);
and AND3 (N1239, N1232, N728, N763);
xor XOR2 (N1240, N1218, N201);
buf BUF1 (N1241, N1236);
nor NOR2 (N1242, N1224, N1034);
buf BUF1 (N1243, N1231);
nor NOR4 (N1244, N1235, N491, N1016, N753);
or OR3 (N1245, N1239, N777, N1242);
nand NAND4 (N1246, N53, N579, N204, N675);
buf BUF1 (N1247, N1245);
not NOT1 (N1248, N1238);
or OR3 (N1249, N1240, N712, N993);
or OR4 (N1250, N1237, N31, N971, N1015);
and AND3 (N1251, N1241, N795, N1015);
nand NAND4 (N1252, N1247, N232, N1167, N991);
nand NAND2 (N1253, N1250, N674);
nand NAND3 (N1254, N1249, N858, N1250);
nand NAND3 (N1255, N1226, N1096, N827);
buf BUF1 (N1256, N1255);
buf BUF1 (N1257, N1246);
xor XOR2 (N1258, N1244, N41);
not NOT1 (N1259, N1257);
xor XOR2 (N1260, N1254, N97);
nand NAND4 (N1261, N1258, N662, N860, N1174);
not NOT1 (N1262, N1260);
and AND4 (N1263, N1256, N404, N774, N183);
nand NAND2 (N1264, N1243, N761);
or OR3 (N1265, N1264, N336, N810);
xor XOR2 (N1266, N1261, N192);
and AND4 (N1267, N1262, N883, N434, N753);
xor XOR2 (N1268, N1251, N1261);
nor NOR4 (N1269, N1268, N1248, N415, N632);
buf BUF1 (N1270, N673);
not NOT1 (N1271, N1269);
and AND2 (N1272, N1267, N1200);
nor NOR4 (N1273, N1263, N1243, N444, N946);
buf BUF1 (N1274, N1265);
buf BUF1 (N1275, N1259);
and AND3 (N1276, N1275, N143, N570);
or OR3 (N1277, N1271, N974, N1102);
nor NOR3 (N1278, N1252, N854, N1136);
or OR3 (N1279, N1272, N260, N1240);
nand NAND4 (N1280, N1277, N1006, N400, N905);
or OR2 (N1281, N1273, N1110);
xor XOR2 (N1282, N1279, N534);
xor XOR2 (N1283, N1282, N406);
nand NAND2 (N1284, N1253, N200);
nor NOR3 (N1285, N1283, N1148, N996);
and AND4 (N1286, N1270, N1181, N161, N154);
not NOT1 (N1287, N1276);
buf BUF1 (N1288, N1287);
or OR2 (N1289, N1274, N1005);
nand NAND4 (N1290, N1233, N24, N1005, N601);
nor NOR3 (N1291, N1290, N1108, N1087);
and AND4 (N1292, N1286, N785, N393, N204);
nor NOR3 (N1293, N1291, N123, N27);
xor XOR2 (N1294, N1293, N174);
buf BUF1 (N1295, N1280);
or OR4 (N1296, N1281, N152, N537, N399);
not NOT1 (N1297, N1296);
nor NOR2 (N1298, N1288, N246);
or OR4 (N1299, N1297, N412, N1297, N1127);
xor XOR2 (N1300, N1285, N505);
buf BUF1 (N1301, N1295);
nand NAND2 (N1302, N1298, N589);
or OR4 (N1303, N1299, N950, N542, N788);
not NOT1 (N1304, N1284);
nand NAND4 (N1305, N1294, N545, N1281, N397);
xor XOR2 (N1306, N1300, N1207);
and AND2 (N1307, N1303, N950);
nor NOR2 (N1308, N1289, N960);
or OR3 (N1309, N1308, N748, N331);
or OR4 (N1310, N1302, N198, N690, N224);
and AND4 (N1311, N1301, N704, N351, N138);
nor NOR4 (N1312, N1292, N827, N428, N1000);
xor XOR2 (N1313, N1305, N274);
nor NOR3 (N1314, N1313, N371, N1005);
nand NAND4 (N1315, N1312, N81, N180, N780);
and AND4 (N1316, N1307, N739, N1040, N297);
nand NAND4 (N1317, N1316, N758, N334, N529);
nor NOR2 (N1318, N1311, N657);
or OR3 (N1319, N1310, N268, N557);
nand NAND2 (N1320, N1319, N50);
nand NAND3 (N1321, N1317, N551, N1235);
not NOT1 (N1322, N1278);
buf BUF1 (N1323, N1304);
buf BUF1 (N1324, N1318);
and AND2 (N1325, N1322, N109);
not NOT1 (N1326, N1315);
nor NOR2 (N1327, N1323, N1285);
nand NAND4 (N1328, N1327, N1271, N104, N1205);
nand NAND2 (N1329, N1314, N1264);
or OR3 (N1330, N1328, N511, N1311);
buf BUF1 (N1331, N1320);
xor XOR2 (N1332, N1309, N349);
nand NAND2 (N1333, N1330, N1067);
nand NAND4 (N1334, N1332, N718, N1317, N914);
or OR4 (N1335, N1329, N6, N847, N1124);
nor NOR4 (N1336, N1326, N199, N904, N402);
not NOT1 (N1337, N1331);
buf BUF1 (N1338, N1266);
and AND3 (N1339, N1325, N761, N385);
xor XOR2 (N1340, N1321, N505);
buf BUF1 (N1341, N1306);
not NOT1 (N1342, N1339);
and AND3 (N1343, N1336, N567, N377);
nand NAND3 (N1344, N1334, N694, N377);
and AND3 (N1345, N1342, N1244, N656);
xor XOR2 (N1346, N1324, N346);
not NOT1 (N1347, N1340);
not NOT1 (N1348, N1338);
xor XOR2 (N1349, N1347, N1303);
or OR2 (N1350, N1343, N1214);
and AND2 (N1351, N1333, N250);
nor NOR3 (N1352, N1341, N549, N574);
not NOT1 (N1353, N1337);
nand NAND3 (N1354, N1345, N708, N315);
or OR3 (N1355, N1354, N4, N897);
nor NOR2 (N1356, N1351, N1235);
xor XOR2 (N1357, N1346, N604);
or OR4 (N1358, N1350, N1012, N1171, N600);
buf BUF1 (N1359, N1357);
not NOT1 (N1360, N1359);
not NOT1 (N1361, N1358);
and AND3 (N1362, N1335, N790, N1242);
not NOT1 (N1363, N1352);
and AND2 (N1364, N1344, N841);
and AND4 (N1365, N1363, N82, N730, N1250);
xor XOR2 (N1366, N1362, N1352);
nor NOR2 (N1367, N1361, N205);
buf BUF1 (N1368, N1353);
buf BUF1 (N1369, N1356);
not NOT1 (N1370, N1367);
or OR3 (N1371, N1369, N1030, N541);
or OR2 (N1372, N1348, N387);
buf BUF1 (N1373, N1366);
not NOT1 (N1374, N1368);
nor NOR3 (N1375, N1373, N856, N128);
buf BUF1 (N1376, N1349);
and AND2 (N1377, N1374, N363);
xor XOR2 (N1378, N1360, N1322);
nand NAND4 (N1379, N1370, N267, N606, N1290);
buf BUF1 (N1380, N1379);
xor XOR2 (N1381, N1372, N224);
or OR2 (N1382, N1377, N958);
not NOT1 (N1383, N1376);
nor NOR2 (N1384, N1371, N671);
and AND4 (N1385, N1365, N1223, N273, N1028);
or OR4 (N1386, N1382, N508, N27, N554);
not NOT1 (N1387, N1355);
nor NOR2 (N1388, N1381, N618);
not NOT1 (N1389, N1364);
or OR4 (N1390, N1389, N1161, N341, N224);
or OR4 (N1391, N1386, N1014, N281, N587);
nor NOR3 (N1392, N1385, N190, N536);
and AND2 (N1393, N1391, N1264);
xor XOR2 (N1394, N1380, N151);
nand NAND2 (N1395, N1387, N1252);
xor XOR2 (N1396, N1388, N183);
xor XOR2 (N1397, N1394, N1116);
nand NAND4 (N1398, N1378, N66, N499, N1187);
not NOT1 (N1399, N1397);
not NOT1 (N1400, N1392);
and AND4 (N1401, N1383, N38, N636, N1148);
buf BUF1 (N1402, N1393);
not NOT1 (N1403, N1398);
and AND3 (N1404, N1375, N899, N143);
and AND4 (N1405, N1396, N48, N259, N420);
nor NOR2 (N1406, N1395, N625);
and AND3 (N1407, N1404, N734, N876);
and AND2 (N1408, N1405, N430);
nor NOR3 (N1409, N1399, N1171, N94);
not NOT1 (N1410, N1384);
nor NOR3 (N1411, N1407, N317, N983);
nor NOR2 (N1412, N1410, N479);
buf BUF1 (N1413, N1400);
not NOT1 (N1414, N1411);
nor NOR4 (N1415, N1413, N1290, N941, N534);
xor XOR2 (N1416, N1409, N97);
nand NAND4 (N1417, N1406, N1003, N70, N1069);
and AND3 (N1418, N1403, N1107, N912);
xor XOR2 (N1419, N1414, N900);
nor NOR3 (N1420, N1417, N360, N981);
buf BUF1 (N1421, N1402);
nor NOR4 (N1422, N1412, N173, N786, N621);
or OR2 (N1423, N1401, N399);
nand NAND2 (N1424, N1415, N168);
nor NOR4 (N1425, N1422, N700, N644, N448);
or OR2 (N1426, N1418, N563);
buf BUF1 (N1427, N1390);
and AND4 (N1428, N1426, N1301, N286, N563);
nand NAND3 (N1429, N1427, N17, N832);
or OR4 (N1430, N1424, N276, N893, N1296);
and AND3 (N1431, N1408, N958, N531);
nand NAND2 (N1432, N1425, N918);
nor NOR3 (N1433, N1431, N508, N1157);
xor XOR2 (N1434, N1432, N1264);
nor NOR2 (N1435, N1434, N1267);
not NOT1 (N1436, N1435);
or OR4 (N1437, N1429, N877, N1139, N1212);
and AND2 (N1438, N1419, N1062);
xor XOR2 (N1439, N1423, N505);
nor NOR3 (N1440, N1416, N919, N171);
nor NOR3 (N1441, N1437, N82, N20);
xor XOR2 (N1442, N1436, N649);
xor XOR2 (N1443, N1439, N37);
xor XOR2 (N1444, N1443, N1073);
xor XOR2 (N1445, N1430, N188);
xor XOR2 (N1446, N1442, N159);
or OR3 (N1447, N1445, N178, N50);
buf BUF1 (N1448, N1441);
xor XOR2 (N1449, N1421, N1246);
or OR2 (N1450, N1444, N754);
buf BUF1 (N1451, N1420);
not NOT1 (N1452, N1450);
buf BUF1 (N1453, N1446);
buf BUF1 (N1454, N1440);
xor XOR2 (N1455, N1428, N1333);
nand NAND3 (N1456, N1447, N45, N694);
or OR4 (N1457, N1433, N179, N298, N406);
xor XOR2 (N1458, N1456, N338);
buf BUF1 (N1459, N1452);
not NOT1 (N1460, N1458);
nand NAND2 (N1461, N1448, N904);
or OR2 (N1462, N1461, N26);
xor XOR2 (N1463, N1455, N328);
not NOT1 (N1464, N1463);
xor XOR2 (N1465, N1457, N1462);
xor XOR2 (N1466, N857, N1462);
or OR4 (N1467, N1454, N92, N612, N1132);
nand NAND2 (N1468, N1451, N975);
nor NOR2 (N1469, N1460, N916);
xor XOR2 (N1470, N1465, N927);
not NOT1 (N1471, N1467);
nor NOR4 (N1472, N1471, N918, N1304, N1358);
nor NOR4 (N1473, N1468, N1425, N489, N1016);
nor NOR3 (N1474, N1472, N832, N510);
nand NAND4 (N1475, N1469, N1351, N432, N82);
and AND3 (N1476, N1438, N950, N318);
not NOT1 (N1477, N1464);
xor XOR2 (N1478, N1466, N1009);
nand NAND4 (N1479, N1449, N425, N589, N1221);
xor XOR2 (N1480, N1476, N387);
nand NAND4 (N1481, N1478, N882, N268, N517);
nand NAND3 (N1482, N1480, N45, N1307);
or OR4 (N1483, N1459, N611, N104, N560);
nand NAND3 (N1484, N1479, N600, N614);
or OR2 (N1485, N1477, N209);
xor XOR2 (N1486, N1484, N691);
not NOT1 (N1487, N1474);
or OR3 (N1488, N1473, N987, N1121);
not NOT1 (N1489, N1487);
buf BUF1 (N1490, N1486);
and AND2 (N1491, N1470, N1057);
not NOT1 (N1492, N1482);
not NOT1 (N1493, N1489);
or OR3 (N1494, N1483, N1455, N990);
and AND4 (N1495, N1494, N1220, N108, N3);
nand NAND3 (N1496, N1492, N7, N589);
nand NAND3 (N1497, N1485, N994, N67);
xor XOR2 (N1498, N1496, N1041);
xor XOR2 (N1499, N1488, N307);
or OR3 (N1500, N1498, N392, N485);
and AND4 (N1501, N1490, N1182, N890, N314);
nor NOR3 (N1502, N1475, N1065, N928);
or OR2 (N1503, N1499, N141);
nor NOR3 (N1504, N1502, N258, N1079);
or OR2 (N1505, N1500, N383);
nor NOR2 (N1506, N1501, N1412);
buf BUF1 (N1507, N1453);
not NOT1 (N1508, N1505);
buf BUF1 (N1509, N1497);
nor NOR2 (N1510, N1507, N1209);
xor XOR2 (N1511, N1493, N203);
xor XOR2 (N1512, N1509, N24);
and AND3 (N1513, N1503, N209, N493);
not NOT1 (N1514, N1508);
not NOT1 (N1515, N1514);
or OR2 (N1516, N1513, N1116);
not NOT1 (N1517, N1504);
not NOT1 (N1518, N1511);
xor XOR2 (N1519, N1510, N1309);
xor XOR2 (N1520, N1518, N392);
nor NOR4 (N1521, N1516, N1446, N998, N35);
nand NAND3 (N1522, N1495, N132, N1508);
buf BUF1 (N1523, N1515);
and AND3 (N1524, N1517, N487, N1173);
not NOT1 (N1525, N1521);
not NOT1 (N1526, N1519);
buf BUF1 (N1527, N1491);
nor NOR3 (N1528, N1523, N730, N6);
nor NOR2 (N1529, N1522, N438);
and AND2 (N1530, N1526, N927);
or OR3 (N1531, N1506, N1015, N1128);
and AND4 (N1532, N1525, N1029, N613, N111);
nor NOR2 (N1533, N1530, N428);
xor XOR2 (N1534, N1533, N260);
not NOT1 (N1535, N1524);
or OR4 (N1536, N1534, N302, N861, N1293);
buf BUF1 (N1537, N1536);
not NOT1 (N1538, N1520);
nand NAND2 (N1539, N1537, N57);
and AND4 (N1540, N1528, N772, N1323, N253);
not NOT1 (N1541, N1539);
or OR3 (N1542, N1529, N815, N186);
not NOT1 (N1543, N1538);
and AND4 (N1544, N1535, N754, N397, N1058);
not NOT1 (N1545, N1481);
not NOT1 (N1546, N1543);
or OR3 (N1547, N1512, N829, N450);
or OR4 (N1548, N1547, N1240, N200, N1184);
nand NAND2 (N1549, N1544, N1174);
xor XOR2 (N1550, N1546, N521);
or OR3 (N1551, N1550, N1537, N1483);
or OR4 (N1552, N1527, N1435, N361, N547);
xor XOR2 (N1553, N1545, N746);
or OR2 (N1554, N1553, N395);
nor NOR2 (N1555, N1552, N976);
nor NOR4 (N1556, N1532, N582, N992, N1273);
buf BUF1 (N1557, N1555);
xor XOR2 (N1558, N1541, N1278);
xor XOR2 (N1559, N1531, N1222);
or OR4 (N1560, N1542, N1095, N627, N782);
xor XOR2 (N1561, N1559, N1063);
and AND2 (N1562, N1548, N888);
nor NOR4 (N1563, N1554, N872, N38, N1501);
not NOT1 (N1564, N1563);
buf BUF1 (N1565, N1551);
xor XOR2 (N1566, N1561, N465);
nor NOR4 (N1567, N1557, N261, N1566, N311);
buf BUF1 (N1568, N594);
xor XOR2 (N1569, N1540, N913);
not NOT1 (N1570, N1556);
buf BUF1 (N1571, N1568);
not NOT1 (N1572, N1571);
nor NOR3 (N1573, N1549, N414, N1237);
or OR2 (N1574, N1567, N288);
nor NOR4 (N1575, N1565, N882, N193, N682);
or OR3 (N1576, N1560, N169, N143);
or OR4 (N1577, N1575, N592, N422, N924);
not NOT1 (N1578, N1576);
nand NAND4 (N1579, N1573, N1315, N1049, N401);
and AND3 (N1580, N1572, N1505, N41);
nor NOR2 (N1581, N1564, N1428);
and AND3 (N1582, N1562, N590, N246);
xor XOR2 (N1583, N1581, N499);
buf BUF1 (N1584, N1579);
buf BUF1 (N1585, N1570);
xor XOR2 (N1586, N1578, N573);
and AND2 (N1587, N1584, N1328);
xor XOR2 (N1588, N1587, N246);
nand NAND2 (N1589, N1582, N279);
or OR3 (N1590, N1585, N928, N851);
not NOT1 (N1591, N1589);
buf BUF1 (N1592, N1558);
nand NAND4 (N1593, N1591, N1370, N189, N642);
buf BUF1 (N1594, N1583);
xor XOR2 (N1595, N1577, N164);
buf BUF1 (N1596, N1569);
or OR3 (N1597, N1595, N1076, N634);
buf BUF1 (N1598, N1580);
not NOT1 (N1599, N1586);
xor XOR2 (N1600, N1596, N414);
xor XOR2 (N1601, N1590, N1366);
and AND4 (N1602, N1593, N1354, N933, N713);
or OR4 (N1603, N1599, N498, N200, N754);
nand NAND3 (N1604, N1594, N1288, N1312);
nand NAND3 (N1605, N1601, N559, N381);
nor NOR3 (N1606, N1592, N897, N518);
xor XOR2 (N1607, N1603, N647);
xor XOR2 (N1608, N1597, N287);
and AND2 (N1609, N1598, N920);
xor XOR2 (N1610, N1588, N1032);
nor NOR3 (N1611, N1610, N681, N1263);
xor XOR2 (N1612, N1605, N836);
nor NOR2 (N1613, N1604, N1158);
nand NAND2 (N1614, N1608, N612);
buf BUF1 (N1615, N1607);
buf BUF1 (N1616, N1611);
and AND4 (N1617, N1602, N339, N1109, N497);
or OR3 (N1618, N1600, N493, N365);
nor NOR3 (N1619, N1612, N115, N1236);
nand NAND3 (N1620, N1619, N718, N90);
nand NAND4 (N1621, N1617, N714, N671, N1548);
not NOT1 (N1622, N1606);
or OR4 (N1623, N1574, N499, N1335, N1184);
buf BUF1 (N1624, N1616);
nor NOR4 (N1625, N1623, N895, N1309, N1511);
nor NOR3 (N1626, N1618, N1526, N1182);
or OR4 (N1627, N1626, N1399, N881, N1441);
or OR3 (N1628, N1614, N533, N537);
nand NAND4 (N1629, N1624, N929, N695, N1069);
xor XOR2 (N1630, N1609, N1504);
or OR4 (N1631, N1621, N1039, N660, N204);
nand NAND2 (N1632, N1630, N930);
buf BUF1 (N1633, N1629);
not NOT1 (N1634, N1631);
nor NOR2 (N1635, N1628, N338);
xor XOR2 (N1636, N1625, N911);
nor NOR4 (N1637, N1620, N4, N1125, N698);
xor XOR2 (N1638, N1636, N1161);
nand NAND2 (N1639, N1637, N985);
xor XOR2 (N1640, N1638, N1549);
and AND2 (N1641, N1615, N478);
and AND2 (N1642, N1640, N1151);
not NOT1 (N1643, N1634);
nand NAND2 (N1644, N1642, N567);
or OR2 (N1645, N1641, N1156);
nor NOR3 (N1646, N1639, N278, N1145);
buf BUF1 (N1647, N1613);
not NOT1 (N1648, N1644);
nor NOR3 (N1649, N1632, N1520, N442);
not NOT1 (N1650, N1645);
or OR4 (N1651, N1650, N286, N1257, N779);
nor NOR3 (N1652, N1627, N1129, N654);
and AND4 (N1653, N1635, N1597, N840, N1537);
or OR2 (N1654, N1622, N1179);
xor XOR2 (N1655, N1648, N168);
nand NAND4 (N1656, N1646, N1378, N1282, N1581);
not NOT1 (N1657, N1652);
or OR3 (N1658, N1653, N200, N298);
nor NOR4 (N1659, N1633, N621, N1201, N1181);
nand NAND4 (N1660, N1656, N785, N877, N1038);
not NOT1 (N1661, N1649);
or OR4 (N1662, N1660, N1495, N13, N366);
nor NOR2 (N1663, N1651, N1373);
nand NAND4 (N1664, N1659, N557, N1239, N1437);
xor XOR2 (N1665, N1664, N962);
or OR2 (N1666, N1663, N1579);
buf BUF1 (N1667, N1662);
nand NAND3 (N1668, N1666, N865, N1538);
xor XOR2 (N1669, N1643, N1249);
nand NAND2 (N1670, N1654, N770);
xor XOR2 (N1671, N1669, N1072);
buf BUF1 (N1672, N1665);
buf BUF1 (N1673, N1670);
and AND3 (N1674, N1661, N1076, N788);
not NOT1 (N1675, N1672);
and AND2 (N1676, N1667, N1367);
not NOT1 (N1677, N1676);
and AND4 (N1678, N1675, N1298, N1085, N1286);
xor XOR2 (N1679, N1671, N1251);
and AND4 (N1680, N1679, N950, N109, N129);
xor XOR2 (N1681, N1680, N1063);
not NOT1 (N1682, N1673);
or OR4 (N1683, N1655, N174, N145, N820);
and AND4 (N1684, N1658, N400, N17, N932);
and AND2 (N1685, N1681, N333);
nor NOR4 (N1686, N1647, N691, N848, N611);
nor NOR3 (N1687, N1668, N1561, N1073);
xor XOR2 (N1688, N1677, N650);
xor XOR2 (N1689, N1674, N112);
not NOT1 (N1690, N1685);
not NOT1 (N1691, N1678);
and AND2 (N1692, N1691, N1264);
buf BUF1 (N1693, N1687);
or OR3 (N1694, N1692, N366, N1617);
buf BUF1 (N1695, N1688);
nor NOR4 (N1696, N1689, N635, N580, N1354);
nand NAND2 (N1697, N1682, N1693);
and AND3 (N1698, N1370, N667, N480);
nand NAND4 (N1699, N1684, N489, N721, N1443);
nor NOR2 (N1700, N1698, N1077);
or OR2 (N1701, N1683, N1453);
nor NOR3 (N1702, N1694, N1198, N1369);
xor XOR2 (N1703, N1697, N803);
and AND2 (N1704, N1695, N1430);
and AND2 (N1705, N1657, N260);
nand NAND4 (N1706, N1704, N33, N1438, N798);
not NOT1 (N1707, N1703);
and AND2 (N1708, N1699, N570);
buf BUF1 (N1709, N1702);
nor NOR4 (N1710, N1705, N1495, N985, N1636);
buf BUF1 (N1711, N1686);
nand NAND3 (N1712, N1711, N550, N514);
buf BUF1 (N1713, N1712);
nor NOR4 (N1714, N1713, N444, N9, N1222);
nand NAND2 (N1715, N1708, N324);
not NOT1 (N1716, N1707);
nand NAND4 (N1717, N1701, N1446, N1127, N210);
buf BUF1 (N1718, N1700);
and AND2 (N1719, N1696, N274);
nor NOR2 (N1720, N1690, N629);
and AND2 (N1721, N1715, N1633);
xor XOR2 (N1722, N1710, N1327);
buf BUF1 (N1723, N1717);
nor NOR2 (N1724, N1719, N631);
xor XOR2 (N1725, N1718, N386);
nand NAND3 (N1726, N1709, N1117, N448);
not NOT1 (N1727, N1720);
not NOT1 (N1728, N1724);
or OR2 (N1729, N1723, N864);
nand NAND4 (N1730, N1729, N40, N931, N301);
nand NAND2 (N1731, N1725, N1600);
or OR2 (N1732, N1714, N473);
nor NOR3 (N1733, N1706, N1281, N298);
or OR3 (N1734, N1721, N1231, N1653);
buf BUF1 (N1735, N1734);
and AND4 (N1736, N1733, N736, N810, N491);
nor NOR2 (N1737, N1730, N1399);
nor NOR3 (N1738, N1716, N590, N213);
xor XOR2 (N1739, N1731, N770);
or OR2 (N1740, N1739, N1292);
not NOT1 (N1741, N1735);
not NOT1 (N1742, N1736);
and AND3 (N1743, N1732, N1560, N228);
nand NAND3 (N1744, N1742, N500, N278);
nor NOR3 (N1745, N1743, N1355, N1729);
not NOT1 (N1746, N1726);
nor NOR4 (N1747, N1740, N754, N299, N1526);
and AND2 (N1748, N1727, N1690);
buf BUF1 (N1749, N1744);
not NOT1 (N1750, N1738);
nand NAND4 (N1751, N1722, N956, N873, N1634);
nand NAND4 (N1752, N1728, N720, N1308, N1146);
or OR4 (N1753, N1741, N1091, N934, N205);
and AND4 (N1754, N1745, N651, N1726, N1567);
and AND2 (N1755, N1737, N1622);
not NOT1 (N1756, N1751);
xor XOR2 (N1757, N1755, N932);
or OR3 (N1758, N1747, N1268, N321);
nand NAND3 (N1759, N1746, N1047, N1511);
nand NAND3 (N1760, N1759, N947, N732);
not NOT1 (N1761, N1760);
and AND4 (N1762, N1754, N1622, N1449, N1565);
nor NOR4 (N1763, N1756, N1194, N753, N1385);
buf BUF1 (N1764, N1750);
or OR4 (N1765, N1752, N1146, N156, N636);
or OR3 (N1766, N1753, N179, N1429);
buf BUF1 (N1767, N1762);
nor NOR4 (N1768, N1764, N1731, N1582, N1062);
and AND3 (N1769, N1748, N1743, N338);
xor XOR2 (N1770, N1768, N116);
or OR3 (N1771, N1758, N1606, N1444);
or OR4 (N1772, N1763, N1198, N394, N1496);
nor NOR3 (N1773, N1767, N841, N566);
nor NOR2 (N1774, N1766, N208);
xor XOR2 (N1775, N1774, N79);
nor NOR3 (N1776, N1769, N754, N1206);
nor NOR2 (N1777, N1765, N882);
and AND4 (N1778, N1761, N125, N468, N107);
nor NOR3 (N1779, N1777, N251, N418);
or OR4 (N1780, N1779, N724, N337, N390);
and AND3 (N1781, N1749, N440, N602);
buf BUF1 (N1782, N1781);
and AND3 (N1783, N1757, N987, N1270);
xor XOR2 (N1784, N1775, N56);
xor XOR2 (N1785, N1776, N708);
and AND3 (N1786, N1773, N1269, N234);
nand NAND4 (N1787, N1780, N928, N1005, N1100);
or OR2 (N1788, N1784, N141);
nand NAND2 (N1789, N1785, N583);
not NOT1 (N1790, N1782);
and AND4 (N1791, N1788, N72, N930, N1255);
nand NAND3 (N1792, N1787, N825, N1513);
or OR3 (N1793, N1792, N436, N1780);
xor XOR2 (N1794, N1786, N915);
nand NAND3 (N1795, N1770, N1321, N915);
xor XOR2 (N1796, N1771, N127);
nand NAND3 (N1797, N1794, N26, N501);
buf BUF1 (N1798, N1795);
or OR3 (N1799, N1789, N1077, N1324);
or OR2 (N1800, N1796, N228);
and AND2 (N1801, N1798, N193);
not NOT1 (N1802, N1801);
or OR3 (N1803, N1791, N257, N1354);
xor XOR2 (N1804, N1800, N339);
xor XOR2 (N1805, N1802, N1040);
nand NAND3 (N1806, N1803, N271, N1725);
not NOT1 (N1807, N1806);
and AND2 (N1808, N1797, N1292);
xor XOR2 (N1809, N1790, N694);
buf BUF1 (N1810, N1809);
nand NAND4 (N1811, N1772, N630, N1613, N1288);
or OR4 (N1812, N1804, N338, N1661, N630);
xor XOR2 (N1813, N1811, N367);
or OR3 (N1814, N1805, N1754, N1422);
and AND3 (N1815, N1814, N1371, N1418);
nor NOR4 (N1816, N1812, N258, N435, N212);
nand NAND2 (N1817, N1813, N1161);
or OR4 (N1818, N1817, N1197, N1145, N1750);
or OR2 (N1819, N1810, N1569);
not NOT1 (N1820, N1815);
or OR3 (N1821, N1818, N1475, N367);
xor XOR2 (N1822, N1821, N317);
nand NAND4 (N1823, N1820, N1065, N1374, N634);
xor XOR2 (N1824, N1778, N552);
buf BUF1 (N1825, N1819);
xor XOR2 (N1826, N1793, N1702);
nor NOR4 (N1827, N1823, N1660, N159, N694);
nor NOR4 (N1828, N1822, N1628, N789, N631);
xor XOR2 (N1829, N1824, N137);
or OR4 (N1830, N1783, N421, N485, N866);
and AND2 (N1831, N1827, N48);
xor XOR2 (N1832, N1799, N151);
buf BUF1 (N1833, N1807);
not NOT1 (N1834, N1831);
or OR2 (N1835, N1830, N420);
not NOT1 (N1836, N1835);
buf BUF1 (N1837, N1808);
xor XOR2 (N1838, N1836, N728);
not NOT1 (N1839, N1825);
xor XOR2 (N1840, N1829, N1472);
or OR4 (N1841, N1834, N1780, N1238, N771);
nor NOR4 (N1842, N1833, N1541, N1538, N970);
xor XOR2 (N1843, N1828, N835);
or OR4 (N1844, N1843, N989, N1274, N1715);
nand NAND3 (N1845, N1838, N1622, N1624);
buf BUF1 (N1846, N1826);
and AND2 (N1847, N1840, N448);
nor NOR2 (N1848, N1847, N692);
or OR2 (N1849, N1816, N1226);
nor NOR2 (N1850, N1841, N357);
buf BUF1 (N1851, N1850);
buf BUF1 (N1852, N1848);
and AND4 (N1853, N1846, N451, N787, N355);
buf BUF1 (N1854, N1852);
buf BUF1 (N1855, N1854);
or OR2 (N1856, N1842, N1464);
nand NAND2 (N1857, N1855, N672);
or OR4 (N1858, N1832, N1258, N944, N574);
nand NAND2 (N1859, N1839, N1351);
nand NAND4 (N1860, N1857, N1444, N310, N1256);
not NOT1 (N1861, N1849);
and AND3 (N1862, N1851, N835, N364);
and AND4 (N1863, N1860, N60, N1436, N1590);
xor XOR2 (N1864, N1837, N1374);
not NOT1 (N1865, N1864);
xor XOR2 (N1866, N1862, N1198);
buf BUF1 (N1867, N1866);
nor NOR3 (N1868, N1861, N898, N1014);
nor NOR3 (N1869, N1845, N552, N551);
xor XOR2 (N1870, N1867, N1587);
xor XOR2 (N1871, N1863, N1364);
xor XOR2 (N1872, N1853, N907);
nand NAND3 (N1873, N1869, N1641, N1586);
and AND2 (N1874, N1872, N1830);
buf BUF1 (N1875, N1873);
nor NOR2 (N1876, N1858, N1083);
buf BUF1 (N1877, N1865);
nor NOR2 (N1878, N1877, N679);
and AND4 (N1879, N1844, N1647, N1415, N1410);
buf BUF1 (N1880, N1871);
and AND3 (N1881, N1856, N635, N1831);
or OR4 (N1882, N1881, N451, N197, N697);
xor XOR2 (N1883, N1875, N39);
buf BUF1 (N1884, N1868);
xor XOR2 (N1885, N1874, N1490);
and AND3 (N1886, N1883, N766, N504);
buf BUF1 (N1887, N1876);
buf BUF1 (N1888, N1880);
or OR2 (N1889, N1859, N30);
and AND4 (N1890, N1889, N784, N299, N1509);
buf BUF1 (N1891, N1879);
nor NOR4 (N1892, N1890, N1512, N1571, N385);
and AND2 (N1893, N1882, N336);
and AND3 (N1894, N1886, N459, N159);
nand NAND2 (N1895, N1888, N5);
and AND3 (N1896, N1891, N321, N127);
or OR4 (N1897, N1885, N565, N133, N1238);
or OR2 (N1898, N1878, N1890);
nand NAND4 (N1899, N1894, N972, N340, N295);
xor XOR2 (N1900, N1892, N1105);
xor XOR2 (N1901, N1887, N525);
buf BUF1 (N1902, N1897);
or OR4 (N1903, N1884, N1448, N1378, N1464);
or OR4 (N1904, N1893, N770, N890, N609);
and AND3 (N1905, N1900, N39, N1081);
buf BUF1 (N1906, N1870);
nand NAND2 (N1907, N1904, N1751);
and AND3 (N1908, N1903, N1714, N1457);
and AND4 (N1909, N1908, N59, N1282, N1831);
buf BUF1 (N1910, N1906);
not NOT1 (N1911, N1909);
buf BUF1 (N1912, N1896);
buf BUF1 (N1913, N1907);
or OR2 (N1914, N1899, N1597);
and AND4 (N1915, N1902, N825, N1046, N1112);
buf BUF1 (N1916, N1901);
xor XOR2 (N1917, N1915, N1546);
and AND3 (N1918, N1914, N1387, N325);
nor NOR2 (N1919, N1911, N1635);
nor NOR3 (N1920, N1916, N926, N1122);
and AND3 (N1921, N1913, N1573, N1674);
and AND3 (N1922, N1895, N238, N1342);
xor XOR2 (N1923, N1921, N122);
or OR2 (N1924, N1917, N891);
nor NOR2 (N1925, N1910, N1785);
nand NAND3 (N1926, N1920, N642, N108);
nand NAND3 (N1927, N1926, N1599, N1905);
or OR3 (N1928, N1021, N1144, N1909);
xor XOR2 (N1929, N1918, N783);
nor NOR4 (N1930, N1924, N1855, N1238, N1262);
buf BUF1 (N1931, N1928);
nor NOR4 (N1932, N1922, N1825, N558, N410);
nand NAND2 (N1933, N1930, N155);
buf BUF1 (N1934, N1898);
not NOT1 (N1935, N1931);
and AND4 (N1936, N1929, N121, N1445, N1191);
xor XOR2 (N1937, N1925, N1747);
or OR2 (N1938, N1919, N1069);
not NOT1 (N1939, N1934);
or OR2 (N1940, N1923, N981);
and AND3 (N1941, N1935, N1055, N196);
nor NOR3 (N1942, N1933, N381, N163);
xor XOR2 (N1943, N1940, N579);
nor NOR2 (N1944, N1932, N1028);
or OR3 (N1945, N1937, N28, N301);
xor XOR2 (N1946, N1912, N1029);
nand NAND2 (N1947, N1936, N1818);
xor XOR2 (N1948, N1947, N316);
not NOT1 (N1949, N1942);
xor XOR2 (N1950, N1948, N603);
nor NOR4 (N1951, N1941, N1397, N1455, N237);
buf BUF1 (N1952, N1945);
not NOT1 (N1953, N1950);
buf BUF1 (N1954, N1944);
xor XOR2 (N1955, N1943, N847);
buf BUF1 (N1956, N1939);
and AND3 (N1957, N1953, N570, N1844);
nand NAND3 (N1958, N1952, N1511, N476);
or OR4 (N1959, N1951, N1225, N1633, N1266);
buf BUF1 (N1960, N1957);
and AND2 (N1961, N1960, N1262);
xor XOR2 (N1962, N1961, N1587);
xor XOR2 (N1963, N1954, N1914);
or OR4 (N1964, N1949, N1683, N611, N507);
nor NOR4 (N1965, N1938, N1051, N1559, N1354);
not NOT1 (N1966, N1959);
buf BUF1 (N1967, N1958);
xor XOR2 (N1968, N1964, N1415);
or OR2 (N1969, N1967, N786);
buf BUF1 (N1970, N1965);
xor XOR2 (N1971, N1963, N1094);
buf BUF1 (N1972, N1966);
xor XOR2 (N1973, N1970, N1529);
or OR3 (N1974, N1968, N1506, N1110);
nand NAND3 (N1975, N1927, N1121, N970);
xor XOR2 (N1976, N1973, N884);
or OR4 (N1977, N1972, N1547, N483, N1933);
buf BUF1 (N1978, N1977);
not NOT1 (N1979, N1974);
or OR2 (N1980, N1956, N1454);
and AND3 (N1981, N1978, N385, N1902);
not NOT1 (N1982, N1979);
not NOT1 (N1983, N1982);
and AND3 (N1984, N1981, N470, N1329);
nor NOR2 (N1985, N1969, N1639);
xor XOR2 (N1986, N1976, N783);
nor NOR4 (N1987, N1962, N1038, N421, N665);
or OR4 (N1988, N1987, N96, N1040, N850);
not NOT1 (N1989, N1971);
nor NOR2 (N1990, N1946, N966);
xor XOR2 (N1991, N1983, N464);
nand NAND4 (N1992, N1975, N111, N873, N1134);
not NOT1 (N1993, N1984);
xor XOR2 (N1994, N1992, N388);
nor NOR2 (N1995, N1990, N379);
or OR3 (N1996, N1985, N1895, N956);
buf BUF1 (N1997, N1986);
xor XOR2 (N1998, N1993, N1965);
or OR3 (N1999, N1995, N101, N966);
or OR2 (N2000, N1991, N1881);
nand NAND3 (N2001, N1998, N1545, N1579);
not NOT1 (N2002, N1988);
buf BUF1 (N2003, N1980);
buf BUF1 (N2004, N2003);
not NOT1 (N2005, N1999);
nor NOR2 (N2006, N2005, N829);
nor NOR2 (N2007, N1997, N1384);
buf BUF1 (N2008, N2006);
not NOT1 (N2009, N2004);
nor NOR3 (N2010, N2009, N1044, N1217);
nand NAND2 (N2011, N1996, N2001);
xor XOR2 (N2012, N1967, N631);
or OR3 (N2013, N2011, N57, N1086);
nand NAND3 (N2014, N2013, N1898, N319);
not NOT1 (N2015, N1994);
or OR3 (N2016, N1989, N1411, N234);
buf BUF1 (N2017, N2012);
not NOT1 (N2018, N2008);
nor NOR3 (N2019, N1955, N742, N136);
or OR4 (N2020, N2014, N1558, N1378, N426);
not NOT1 (N2021, N2016);
nand NAND4 (N2022, N2020, N127, N1394, N367);
or OR2 (N2023, N2022, N818);
xor XOR2 (N2024, N2015, N415);
nand NAND3 (N2025, N2021, N305, N657);
nor NOR4 (N2026, N2007, N612, N1080, N727);
xor XOR2 (N2027, N2025, N784);
nand NAND3 (N2028, N2027, N1644, N393);
nand NAND4 (N2029, N2026, N1884, N1929, N249);
nand NAND4 (N2030, N2024, N283, N470, N815);
xor XOR2 (N2031, N2017, N304);
not NOT1 (N2032, N2028);
nand NAND2 (N2033, N2019, N1316);
xor XOR2 (N2034, N2018, N365);
nor NOR3 (N2035, N2030, N613, N676);
and AND3 (N2036, N2010, N139, N1103);
xor XOR2 (N2037, N2032, N398);
nand NAND4 (N2038, N2036, N947, N1825, N175);
buf BUF1 (N2039, N2029);
or OR3 (N2040, N2031, N108, N2011);
xor XOR2 (N2041, N2040, N216);
nor NOR3 (N2042, N2035, N1937, N685);
buf BUF1 (N2043, N2037);
nand NAND4 (N2044, N2002, N478, N2032, N1607);
or OR3 (N2045, N2039, N1381, N122);
nand NAND3 (N2046, N2042, N1491, N387);
and AND2 (N2047, N2034, N144);
or OR4 (N2048, N2000, N680, N1297, N1908);
nor NOR4 (N2049, N2047, N72, N1542, N1402);
xor XOR2 (N2050, N2023, N1919);
and AND2 (N2051, N2050, N619);
and AND3 (N2052, N2051, N84, N1739);
not NOT1 (N2053, N2043);
and AND2 (N2054, N2052, N145);
buf BUF1 (N2055, N2048);
nor NOR4 (N2056, N2033, N1340, N338, N1222);
nand NAND4 (N2057, N2049, N1839, N512, N745);
and AND2 (N2058, N2055, N180);
and AND2 (N2059, N2057, N611);
and AND3 (N2060, N2045, N1306, N219);
or OR2 (N2061, N2060, N85);
and AND3 (N2062, N2053, N1570, N797);
and AND3 (N2063, N2041, N741, N2052);
or OR3 (N2064, N2056, N858, N2031);
nand NAND4 (N2065, N2064, N1769, N1344, N1553);
not NOT1 (N2066, N2038);
not NOT1 (N2067, N2058);
buf BUF1 (N2068, N2061);
not NOT1 (N2069, N2054);
nor NOR3 (N2070, N2068, N2009, N1555);
and AND3 (N2071, N2066, N1054, N1024);
nor NOR2 (N2072, N2046, N1553);
nor NOR2 (N2073, N2070, N1722);
or OR2 (N2074, N2073, N1386);
nor NOR2 (N2075, N2065, N1877);
xor XOR2 (N2076, N2074, N932);
nor NOR2 (N2077, N2072, N1314);
and AND2 (N2078, N2044, N728);
and AND3 (N2079, N2078, N1986, N1622);
nand NAND3 (N2080, N2077, N462, N1499);
xor XOR2 (N2081, N2069, N1240);
xor XOR2 (N2082, N2063, N746);
buf BUF1 (N2083, N2080);
buf BUF1 (N2084, N2071);
nor NOR2 (N2085, N2062, N661);
nand NAND3 (N2086, N2067, N1455, N1281);
and AND3 (N2087, N2085, N285, N1239);
and AND2 (N2088, N2087, N717);
and AND3 (N2089, N2076, N375, N1350);
nor NOR3 (N2090, N2082, N844, N1913);
not NOT1 (N2091, N2075);
or OR4 (N2092, N2089, N1454, N751, N1093);
and AND3 (N2093, N2083, N208, N1083);
xor XOR2 (N2094, N2090, N1289);
buf BUF1 (N2095, N2059);
nand NAND3 (N2096, N2091, N705, N1165);
or OR4 (N2097, N2084, N1910, N1118, N763);
buf BUF1 (N2098, N2092);
and AND3 (N2099, N2081, N1770, N854);
and AND4 (N2100, N2096, N658, N27, N284);
or OR4 (N2101, N2099, N1993, N1935, N1166);
nand NAND2 (N2102, N2101, N1804);
not NOT1 (N2103, N2093);
or OR3 (N2104, N2097, N1709, N1191);
not NOT1 (N2105, N2103);
or OR2 (N2106, N2095, N603);
or OR3 (N2107, N2086, N211, N1383);
xor XOR2 (N2108, N2104, N1295);
or OR2 (N2109, N2088, N1510);
and AND3 (N2110, N2108, N1198, N303);
buf BUF1 (N2111, N2107);
nor NOR3 (N2112, N2106, N2052, N606);
and AND2 (N2113, N2111, N1215);
or OR2 (N2114, N2079, N1329);
not NOT1 (N2115, N2110);
nor NOR2 (N2116, N2109, N1585);
buf BUF1 (N2117, N2116);
or OR4 (N2118, N2105, N1984, N1180, N1586);
not NOT1 (N2119, N2118);
xor XOR2 (N2120, N2112, N1447);
or OR4 (N2121, N2100, N2104, N359, N646);
nor NOR3 (N2122, N2121, N1613, N80);
not NOT1 (N2123, N2119);
or OR4 (N2124, N2120, N917, N510, N1790);
not NOT1 (N2125, N2113);
or OR3 (N2126, N2125, N304, N527);
nand NAND2 (N2127, N2114, N1186);
nor NOR2 (N2128, N2117, N25);
nor NOR4 (N2129, N2098, N367, N1289, N1571);
nand NAND3 (N2130, N2094, N501, N463);
or OR4 (N2131, N2127, N1402, N740, N269);
nor NOR3 (N2132, N2102, N760, N1945);
not NOT1 (N2133, N2115);
nand NAND4 (N2134, N2124, N293, N649, N2036);
nand NAND2 (N2135, N2128, N289);
nor NOR4 (N2136, N2132, N1679, N1000, N596);
nor NOR4 (N2137, N2135, N768, N710, N1530);
nand NAND4 (N2138, N2122, N255, N718, N1492);
not NOT1 (N2139, N2123);
buf BUF1 (N2140, N2137);
buf BUF1 (N2141, N2136);
buf BUF1 (N2142, N2130);
and AND4 (N2143, N2131, N360, N132, N215);
xor XOR2 (N2144, N2142, N1408);
buf BUF1 (N2145, N2144);
buf BUF1 (N2146, N2129);
not NOT1 (N2147, N2145);
xor XOR2 (N2148, N2133, N525);
buf BUF1 (N2149, N2139);
or OR3 (N2150, N2148, N324, N1265);
nor NOR4 (N2151, N2143, N102, N1160, N767);
buf BUF1 (N2152, N2147);
xor XOR2 (N2153, N2134, N1695);
not NOT1 (N2154, N2138);
xor XOR2 (N2155, N2152, N647);
and AND3 (N2156, N2155, N598, N2027);
or OR2 (N2157, N2146, N418);
nand NAND4 (N2158, N2151, N1887, N594, N1525);
nand NAND3 (N2159, N2157, N989, N1828);
or OR3 (N2160, N2153, N1891, N848);
nor NOR3 (N2161, N2156, N1657, N1919);
buf BUF1 (N2162, N2149);
and AND2 (N2163, N2150, N1963);
nor NOR4 (N2164, N2162, N919, N1877, N1405);
nor NOR3 (N2165, N2126, N770, N763);
not NOT1 (N2166, N2165);
and AND4 (N2167, N2140, N1846, N1312, N1401);
xor XOR2 (N2168, N2161, N954);
xor XOR2 (N2169, N2160, N305);
xor XOR2 (N2170, N2164, N1973);
xor XOR2 (N2171, N2167, N543);
and AND4 (N2172, N2168, N955, N765, N1884);
and AND3 (N2173, N2170, N36, N383);
xor XOR2 (N2174, N2154, N1401);
not NOT1 (N2175, N2172);
and AND3 (N2176, N2141, N1723, N1006);
nand NAND3 (N2177, N2174, N101, N2143);
not NOT1 (N2178, N2173);
xor XOR2 (N2179, N2169, N384);
not NOT1 (N2180, N2158);
nor NOR2 (N2181, N2179, N1489);
buf BUF1 (N2182, N2175);
xor XOR2 (N2183, N2166, N1384);
xor XOR2 (N2184, N2182, N1835);
xor XOR2 (N2185, N2159, N69);
xor XOR2 (N2186, N2181, N505);
not NOT1 (N2187, N2184);
not NOT1 (N2188, N2183);
or OR4 (N2189, N2177, N1301, N664, N1243);
nor NOR2 (N2190, N2178, N1570);
nand NAND4 (N2191, N2180, N1088, N1716, N507);
buf BUF1 (N2192, N2188);
xor XOR2 (N2193, N2185, N1071);
nand NAND2 (N2194, N2192, N78);
buf BUF1 (N2195, N2163);
xor XOR2 (N2196, N2190, N679);
and AND3 (N2197, N2176, N631, N1080);
and AND4 (N2198, N2187, N1166, N1726, N2014);
or OR3 (N2199, N2198, N494, N1035);
xor XOR2 (N2200, N2196, N26);
or OR2 (N2201, N2197, N1729);
or OR4 (N2202, N2201, N2178, N1033, N1913);
xor XOR2 (N2203, N2199, N1465);
xor XOR2 (N2204, N2189, N983);
not NOT1 (N2205, N2171);
nor NOR2 (N2206, N2204, N825);
buf BUF1 (N2207, N2194);
xor XOR2 (N2208, N2203, N1960);
or OR4 (N2209, N2195, N80, N1821, N1600);
xor XOR2 (N2210, N2206, N564);
xor XOR2 (N2211, N2200, N1964);
not NOT1 (N2212, N2191);
nor NOR2 (N2213, N2205, N1730);
nor NOR3 (N2214, N2210, N473, N1815);
nor NOR3 (N2215, N2214, N959, N2102);
xor XOR2 (N2216, N2207, N1532);
nor NOR2 (N2217, N2213, N2040);
nand NAND3 (N2218, N2186, N1813, N132);
nor NOR4 (N2219, N2211, N882, N1345, N860);
buf BUF1 (N2220, N2193);
nand NAND3 (N2221, N2219, N376, N1050);
buf BUF1 (N2222, N2208);
nor NOR4 (N2223, N2209, N61, N228, N188);
and AND2 (N2224, N2202, N1873);
nand NAND3 (N2225, N2222, N1779, N74);
nor NOR3 (N2226, N2225, N405, N269);
xor XOR2 (N2227, N2215, N2167);
buf BUF1 (N2228, N2227);
or OR2 (N2229, N2221, N1561);
or OR2 (N2230, N2216, N1113);
and AND3 (N2231, N2217, N1101, N1648);
xor XOR2 (N2232, N2220, N2147);
nor NOR3 (N2233, N2232, N1971, N1601);
not NOT1 (N2234, N2226);
not NOT1 (N2235, N2233);
and AND4 (N2236, N2218, N993, N1547, N1192);
nor NOR2 (N2237, N2228, N239);
or OR2 (N2238, N2234, N666);
or OR4 (N2239, N2212, N1480, N1011, N1002);
or OR4 (N2240, N2237, N1218, N791, N513);
not NOT1 (N2241, N2236);
not NOT1 (N2242, N2241);
and AND2 (N2243, N2223, N1769);
xor XOR2 (N2244, N2231, N37);
not NOT1 (N2245, N2243);
not NOT1 (N2246, N2244);
or OR2 (N2247, N2224, N2172);
not NOT1 (N2248, N2230);
xor XOR2 (N2249, N2238, N521);
nor NOR2 (N2250, N2245, N432);
nor NOR3 (N2251, N2239, N116, N510);
or OR4 (N2252, N2242, N1713, N812, N1012);
and AND2 (N2253, N2251, N726);
and AND2 (N2254, N2246, N1087);
buf BUF1 (N2255, N2253);
buf BUF1 (N2256, N2252);
nand NAND3 (N2257, N2247, N1741, N99);
or OR3 (N2258, N2229, N466, N1340);
or OR4 (N2259, N2255, N1593, N1235, N782);
or OR3 (N2260, N2240, N635, N642);
and AND4 (N2261, N2248, N1927, N1250, N1570);
not NOT1 (N2262, N2259);
buf BUF1 (N2263, N2250);
xor XOR2 (N2264, N2258, N1187);
nand NAND4 (N2265, N2249, N2027, N1273, N1706);
xor XOR2 (N2266, N2257, N1739);
not NOT1 (N2267, N2265);
or OR3 (N2268, N2254, N22, N820);
buf BUF1 (N2269, N2266);
nor NOR2 (N2270, N2263, N883);
nand NAND2 (N2271, N2261, N2030);
or OR4 (N2272, N2267, N1932, N1367, N883);
nor NOR3 (N2273, N2270, N1582, N494);
and AND2 (N2274, N2269, N1647);
and AND2 (N2275, N2268, N1784);
and AND2 (N2276, N2260, N194);
nand NAND3 (N2277, N2272, N75, N471);
buf BUF1 (N2278, N2273);
nand NAND3 (N2279, N2264, N2087, N1309);
nand NAND2 (N2280, N2262, N329);
and AND2 (N2281, N2256, N2167);
xor XOR2 (N2282, N2281, N547);
buf BUF1 (N2283, N2275);
nor NOR2 (N2284, N2274, N1682);
xor XOR2 (N2285, N2235, N953);
nand NAND2 (N2286, N2284, N948);
buf BUF1 (N2287, N2282);
buf BUF1 (N2288, N2276);
xor XOR2 (N2289, N2278, N1871);
nand NAND2 (N2290, N2271, N796);
xor XOR2 (N2291, N2288, N871);
xor XOR2 (N2292, N2291, N1696);
and AND2 (N2293, N2279, N1900);
nor NOR3 (N2294, N2280, N1624, N1920);
xor XOR2 (N2295, N2293, N2174);
nor NOR2 (N2296, N2289, N302);
nor NOR3 (N2297, N2285, N2246, N1277);
buf BUF1 (N2298, N2295);
and AND3 (N2299, N2292, N1820, N2174);
xor XOR2 (N2300, N2290, N520);
xor XOR2 (N2301, N2283, N1734);
nor NOR2 (N2302, N2286, N1407);
and AND4 (N2303, N2297, N2017, N182, N2045);
nand NAND3 (N2304, N2287, N352, N2136);
nand NAND2 (N2305, N2299, N1374);
and AND3 (N2306, N2302, N1223, N133);
buf BUF1 (N2307, N2305);
nand NAND4 (N2308, N2303, N1853, N775, N1007);
nor NOR2 (N2309, N2306, N313);
xor XOR2 (N2310, N2296, N595);
and AND4 (N2311, N2310, N25, N310, N1333);
nand NAND4 (N2312, N2307, N1924, N2201, N157);
not NOT1 (N2313, N2294);
or OR2 (N2314, N2300, N822);
not NOT1 (N2315, N2304);
nand NAND4 (N2316, N2308, N476, N208, N1167);
xor XOR2 (N2317, N2313, N2017);
and AND4 (N2318, N2315, N2032, N2019, N2135);
xor XOR2 (N2319, N2309, N1682);
nor NOR3 (N2320, N2319, N875, N90);
not NOT1 (N2321, N2298);
or OR2 (N2322, N2321, N2185);
nor NOR2 (N2323, N2301, N136);
xor XOR2 (N2324, N2323, N1402);
xor XOR2 (N2325, N2320, N707);
xor XOR2 (N2326, N2316, N45);
xor XOR2 (N2327, N2277, N1568);
and AND4 (N2328, N2314, N1565, N2143, N2205);
or OR3 (N2329, N2325, N588, N1643);
not NOT1 (N2330, N2312);
nor NOR2 (N2331, N2328, N576);
nor NOR4 (N2332, N2326, N1773, N1596, N520);
buf BUF1 (N2333, N2318);
and AND4 (N2334, N2327, N1642, N714, N27);
and AND3 (N2335, N2330, N873, N533);
nor NOR4 (N2336, N2322, N2094, N1935, N1847);
nor NOR4 (N2337, N2311, N718, N853, N455);
nor NOR4 (N2338, N2324, N1592, N1954, N423);
xor XOR2 (N2339, N2337, N1946);
buf BUF1 (N2340, N2332);
buf BUF1 (N2341, N2333);
nor NOR3 (N2342, N2331, N1269, N519);
and AND3 (N2343, N2338, N269, N83);
xor XOR2 (N2344, N2329, N668);
buf BUF1 (N2345, N2344);
nand NAND2 (N2346, N2343, N659);
or OR4 (N2347, N2346, N1247, N168, N2198);
buf BUF1 (N2348, N2341);
not NOT1 (N2349, N2340);
not NOT1 (N2350, N2317);
nand NAND2 (N2351, N2342, N1732);
buf BUF1 (N2352, N2348);
nor NOR3 (N2353, N2339, N797, N1965);
nor NOR4 (N2354, N2345, N1243, N949, N1348);
or OR4 (N2355, N2335, N239, N921, N2342);
nand NAND4 (N2356, N2351, N955, N553, N1906);
nand NAND2 (N2357, N2356, N807);
and AND4 (N2358, N2354, N2011, N1302, N1178);
nand NAND3 (N2359, N2336, N1353, N652);
or OR4 (N2360, N2359, N54, N1524, N763);
nand NAND4 (N2361, N2355, N894, N350, N2305);
nand NAND2 (N2362, N2357, N1537);
nand NAND3 (N2363, N2353, N1564, N714);
not NOT1 (N2364, N2360);
xor XOR2 (N2365, N2364, N1289);
buf BUF1 (N2366, N2352);
and AND4 (N2367, N2350, N48, N1351, N1869);
or OR3 (N2368, N2362, N216, N486);
and AND3 (N2369, N2366, N1789, N1302);
and AND3 (N2370, N2363, N146, N721);
and AND4 (N2371, N2347, N343, N2327, N2141);
nor NOR3 (N2372, N2334, N710, N1348);
or OR4 (N2373, N2368, N1480, N1281, N1023);
not NOT1 (N2374, N2361);
nand NAND4 (N2375, N2365, N1503, N2015, N1086);
not NOT1 (N2376, N2367);
not NOT1 (N2377, N2358);
and AND4 (N2378, N2371, N557, N283, N1457);
xor XOR2 (N2379, N2378, N753);
not NOT1 (N2380, N2375);
buf BUF1 (N2381, N2349);
nor NOR2 (N2382, N2379, N1528);
xor XOR2 (N2383, N2372, N646);
nor NOR2 (N2384, N2380, N16);
nand NAND2 (N2385, N2369, N288);
and AND2 (N2386, N2385, N1829);
or OR3 (N2387, N2381, N905, N2104);
nor NOR4 (N2388, N2384, N1402, N1572, N625);
and AND3 (N2389, N2383, N1069, N2181);
buf BUF1 (N2390, N2386);
or OR2 (N2391, N2388, N2213);
or OR3 (N2392, N2377, N1202, N248);
or OR3 (N2393, N2387, N475, N450);
and AND3 (N2394, N2389, N1935, N2355);
or OR3 (N2395, N2374, N1486, N702);
and AND4 (N2396, N2373, N2, N1482, N2389);
buf BUF1 (N2397, N2396);
and AND2 (N2398, N2395, N586);
not NOT1 (N2399, N2394);
nand NAND2 (N2400, N2397, N2089);
or OR4 (N2401, N2392, N1983, N1148, N439);
or OR4 (N2402, N2399, N1474, N618, N1215);
or OR3 (N2403, N2398, N1456, N217);
nor NOR4 (N2404, N2402, N1884, N1416, N1103);
or OR4 (N2405, N2382, N1742, N419, N114);
buf BUF1 (N2406, N2393);
buf BUF1 (N2407, N2406);
nand NAND2 (N2408, N2403, N1143);
not NOT1 (N2409, N2401);
not NOT1 (N2410, N2405);
or OR3 (N2411, N2409, N1000, N1301);
not NOT1 (N2412, N2404);
nor NOR2 (N2413, N2390, N1835);
nand NAND4 (N2414, N2376, N1289, N246, N1944);
or OR2 (N2415, N2410, N1756);
nand NAND4 (N2416, N2408, N2385, N361, N1110);
not NOT1 (N2417, N2400);
and AND4 (N2418, N2391, N727, N608, N65);
not NOT1 (N2419, N2417);
not NOT1 (N2420, N2407);
and AND4 (N2421, N2370, N2231, N1642, N702);
nor NOR3 (N2422, N2412, N1162, N2261);
or OR3 (N2423, N2413, N1909, N118);
xor XOR2 (N2424, N2422, N2386);
buf BUF1 (N2425, N2419);
nand NAND4 (N2426, N2421, N2199, N1146, N812);
buf BUF1 (N2427, N2411);
xor XOR2 (N2428, N2416, N2229);
xor XOR2 (N2429, N2414, N238);
not NOT1 (N2430, N2424);
not NOT1 (N2431, N2423);
or OR3 (N2432, N2427, N1037, N1830);
or OR4 (N2433, N2428, N1358, N1679, N239);
buf BUF1 (N2434, N2426);
not NOT1 (N2435, N2415);
buf BUF1 (N2436, N2432);
nor NOR3 (N2437, N2430, N2338, N146);
not NOT1 (N2438, N2436);
buf BUF1 (N2439, N2435);
nand NAND4 (N2440, N2434, N633, N432, N1004);
and AND2 (N2441, N2431, N1670);
not NOT1 (N2442, N2418);
buf BUF1 (N2443, N2420);
nand NAND2 (N2444, N2425, N2204);
nor NOR3 (N2445, N2438, N2137, N711);
not NOT1 (N2446, N2429);
nand NAND4 (N2447, N2441, N983, N267, N298);
nor NOR3 (N2448, N2442, N2275, N418);
buf BUF1 (N2449, N2445);
buf BUF1 (N2450, N2443);
or OR4 (N2451, N2437, N2307, N869, N493);
or OR4 (N2452, N2449, N1792, N315, N974);
xor XOR2 (N2453, N2440, N825);
buf BUF1 (N2454, N2453);
nand NAND4 (N2455, N2448, N59, N232, N1324);
buf BUF1 (N2456, N2450);
or OR2 (N2457, N2455, N546);
and AND4 (N2458, N2446, N1731, N134, N1822);
xor XOR2 (N2459, N2433, N451);
and AND2 (N2460, N2444, N1157);
nand NAND2 (N2461, N2439, N1439);
buf BUF1 (N2462, N2452);
nor NOR3 (N2463, N2458, N1159, N2289);
nand NAND3 (N2464, N2451, N2015, N1503);
buf BUF1 (N2465, N2461);
buf BUF1 (N2466, N2465);
not NOT1 (N2467, N2454);
nand NAND2 (N2468, N2466, N568);
not NOT1 (N2469, N2463);
nand NAND2 (N2470, N2447, N402);
or OR2 (N2471, N2456, N122);
xor XOR2 (N2472, N2460, N2029);
xor XOR2 (N2473, N2464, N1967);
nand NAND4 (N2474, N2459, N1158, N836, N458);
not NOT1 (N2475, N2469);
nand NAND2 (N2476, N2472, N2152);
not NOT1 (N2477, N2476);
xor XOR2 (N2478, N2477, N1049);
buf BUF1 (N2479, N2468);
nor NOR2 (N2480, N2470, N162);
xor XOR2 (N2481, N2474, N607);
buf BUF1 (N2482, N2480);
xor XOR2 (N2483, N2462, N1907);
nand NAND3 (N2484, N2457, N1233, N1821);
buf BUF1 (N2485, N2484);
nor NOR3 (N2486, N2479, N1583, N1615);
or OR4 (N2487, N2482, N2157, N2103, N1268);
nor NOR2 (N2488, N2473, N427);
nor NOR4 (N2489, N2481, N841, N665, N1699);
not NOT1 (N2490, N2467);
not NOT1 (N2491, N2485);
and AND3 (N2492, N2488, N2274, N2298);
nor NOR4 (N2493, N2486, N1265, N841, N942);
buf BUF1 (N2494, N2491);
buf BUF1 (N2495, N2478);
nor NOR4 (N2496, N2483, N2427, N1495, N408);
or OR4 (N2497, N2495, N1188, N1344, N1442);
buf BUF1 (N2498, N2497);
nor NOR4 (N2499, N2496, N660, N1107, N835);
or OR2 (N2500, N2494, N814);
nor NOR2 (N2501, N2489, N87);
xor XOR2 (N2502, N2487, N2256);
buf BUF1 (N2503, N2501);
nor NOR3 (N2504, N2500, N148, N1266);
and AND4 (N2505, N2490, N2489, N1099, N1887);
buf BUF1 (N2506, N2493);
nor NOR4 (N2507, N2504, N2311, N1482, N2441);
xor XOR2 (N2508, N2498, N1280);
buf BUF1 (N2509, N2505);
not NOT1 (N2510, N2503);
not NOT1 (N2511, N2506);
or OR3 (N2512, N2507, N1017, N484);
buf BUF1 (N2513, N2510);
xor XOR2 (N2514, N2492, N1182);
and AND4 (N2515, N2509, N2285, N2461, N341);
nor NOR3 (N2516, N2513, N1267, N2274);
xor XOR2 (N2517, N2516, N424);
or OR4 (N2518, N2471, N253, N314, N1676);
nand NAND4 (N2519, N2518, N253, N2184, N900);
xor XOR2 (N2520, N2508, N1205);
xor XOR2 (N2521, N2499, N134);
or OR2 (N2522, N2517, N1137);
nand NAND3 (N2523, N2511, N1686, N387);
or OR3 (N2524, N2521, N2293, N2112);
or OR2 (N2525, N2502, N537);
nor NOR3 (N2526, N2523, N314, N2373);
nor NOR2 (N2527, N2526, N562);
nand NAND4 (N2528, N2519, N2023, N1923, N2425);
xor XOR2 (N2529, N2522, N1805);
buf BUF1 (N2530, N2524);
or OR3 (N2531, N2525, N2382, N2217);
buf BUF1 (N2532, N2529);
nand NAND2 (N2533, N2520, N1354);
buf BUF1 (N2534, N2515);
or OR3 (N2535, N2534, N749, N1417);
nor NOR2 (N2536, N2535, N1050);
and AND4 (N2537, N2530, N1701, N2484, N1737);
nor NOR3 (N2538, N2528, N1880, N703);
or OR3 (N2539, N2533, N1666, N1309);
and AND2 (N2540, N2532, N1204);
or OR2 (N2541, N2514, N564);
nand NAND3 (N2542, N2538, N1204, N1374);
nand NAND4 (N2543, N2540, N2283, N1255, N1184);
nor NOR4 (N2544, N2527, N941, N1582, N537);
xor XOR2 (N2545, N2537, N609);
not NOT1 (N2546, N2512);
buf BUF1 (N2547, N2541);
or OR3 (N2548, N2547, N1559, N220);
xor XOR2 (N2549, N2539, N1340);
not NOT1 (N2550, N2549);
and AND4 (N2551, N2531, N2048, N712, N2439);
nor NOR2 (N2552, N2546, N1033);
or OR2 (N2553, N2545, N2112);
nand NAND4 (N2554, N2552, N2265, N2395, N104);
and AND3 (N2555, N2553, N328, N2342);
xor XOR2 (N2556, N2475, N237);
not NOT1 (N2557, N2551);
and AND4 (N2558, N2556, N1734, N2327, N1829);
xor XOR2 (N2559, N2542, N206);
xor XOR2 (N2560, N2559, N1245);
xor XOR2 (N2561, N2557, N1845);
buf BUF1 (N2562, N2560);
nor NOR3 (N2563, N2544, N334, N362);
nand NAND4 (N2564, N2558, N230, N810, N1044);
xor XOR2 (N2565, N2563, N1662);
buf BUF1 (N2566, N2554);
and AND2 (N2567, N2555, N2083);
buf BUF1 (N2568, N2564);
buf BUF1 (N2569, N2550);
or OR4 (N2570, N2569, N76, N2067, N1712);
and AND4 (N2571, N2566, N2531, N1485, N2217);
nor NOR4 (N2572, N2561, N2261, N2239, N1341);
or OR3 (N2573, N2570, N1477, N1528);
buf BUF1 (N2574, N2573);
xor XOR2 (N2575, N2562, N57);
not NOT1 (N2576, N2572);
and AND3 (N2577, N2565, N2453, N836);
xor XOR2 (N2578, N2571, N2528);
nor NOR3 (N2579, N2536, N1749, N684);
nand NAND3 (N2580, N2543, N1564, N695);
and AND4 (N2581, N2568, N502, N1992, N2510);
nand NAND2 (N2582, N2578, N1422);
nand NAND3 (N2583, N2580, N842, N1294);
xor XOR2 (N2584, N2548, N1101);
not NOT1 (N2585, N2577);
nand NAND2 (N2586, N2585, N1587);
xor XOR2 (N2587, N2583, N237);
xor XOR2 (N2588, N2582, N1884);
nor NOR2 (N2589, N2581, N1886);
buf BUF1 (N2590, N2575);
or OR2 (N2591, N2574, N726);
buf BUF1 (N2592, N2586);
nor NOR2 (N2593, N2584, N1435);
not NOT1 (N2594, N2590);
xor XOR2 (N2595, N2592, N549);
and AND4 (N2596, N2589, N1189, N1022, N1169);
not NOT1 (N2597, N2596);
xor XOR2 (N2598, N2597, N1494);
nand NAND3 (N2599, N2598, N1263, N986);
buf BUF1 (N2600, N2576);
xor XOR2 (N2601, N2567, N1295);
buf BUF1 (N2602, N2601);
buf BUF1 (N2603, N2602);
nand NAND4 (N2604, N2588, N514, N2528, N645);
nor NOR4 (N2605, N2587, N1761, N1742, N2407);
nand NAND3 (N2606, N2591, N1914, N80);
xor XOR2 (N2607, N2603, N1605);
not NOT1 (N2608, N2606);
nand NAND2 (N2609, N2608, N626);
buf BUF1 (N2610, N2595);
not NOT1 (N2611, N2600);
not NOT1 (N2612, N2607);
nand NAND4 (N2613, N2599, N787, N2338, N1608);
and AND3 (N2614, N2613, N766, N1953);
nand NAND4 (N2615, N2579, N149, N1875, N1304);
xor XOR2 (N2616, N2611, N2352);
xor XOR2 (N2617, N2593, N2434);
xor XOR2 (N2618, N2614, N1268);
or OR4 (N2619, N2594, N2003, N494, N262);
nor NOR3 (N2620, N2617, N1583, N23);
nor NOR3 (N2621, N2615, N1008, N2018);
or OR4 (N2622, N2605, N215, N2546, N1426);
xor XOR2 (N2623, N2612, N1123);
or OR2 (N2624, N2616, N68);
not NOT1 (N2625, N2620);
and AND4 (N2626, N2610, N2078, N164, N1248);
not NOT1 (N2627, N2621);
nor NOR4 (N2628, N2618, N1161, N1870, N1000);
nor NOR3 (N2629, N2625, N1749, N2571);
or OR2 (N2630, N2624, N2220);
not NOT1 (N2631, N2630);
and AND2 (N2632, N2609, N844);
or OR4 (N2633, N2627, N35, N1062, N1085);
not NOT1 (N2634, N2632);
nor NOR2 (N2635, N2622, N1964);
nor NOR2 (N2636, N2633, N1708);
or OR2 (N2637, N2623, N1267);
or OR3 (N2638, N2636, N1382, N926);
not NOT1 (N2639, N2631);
buf BUF1 (N2640, N2626);
or OR4 (N2641, N2629, N1090, N2145, N1922);
not NOT1 (N2642, N2638);
nand NAND4 (N2643, N2635, N228, N612, N731);
and AND4 (N2644, N2639, N934, N1605, N1864);
nor NOR4 (N2645, N2619, N2555, N78, N2195);
xor XOR2 (N2646, N2634, N2577);
xor XOR2 (N2647, N2628, N1338);
nand NAND4 (N2648, N2643, N16, N1379, N933);
buf BUF1 (N2649, N2640);
and AND4 (N2650, N2604, N1422, N2458, N202);
buf BUF1 (N2651, N2646);
or OR4 (N2652, N2650, N2594, N2529, N2356);
buf BUF1 (N2653, N2648);
nand NAND3 (N2654, N2651, N996, N2545);
nor NOR4 (N2655, N2652, N2005, N2367, N810);
nand NAND4 (N2656, N2637, N1847, N1501, N1166);
nand NAND3 (N2657, N2653, N759, N2568);
buf BUF1 (N2658, N2657);
xor XOR2 (N2659, N2641, N1497);
or OR2 (N2660, N2645, N1413);
and AND2 (N2661, N2656, N1575);
not NOT1 (N2662, N2660);
nor NOR4 (N2663, N2659, N49, N850, N748);
or OR3 (N2664, N2662, N1106, N768);
not NOT1 (N2665, N2644);
not NOT1 (N2666, N2661);
not NOT1 (N2667, N2649);
buf BUF1 (N2668, N2663);
buf BUF1 (N2669, N2665);
not NOT1 (N2670, N2666);
or OR2 (N2671, N2670, N674);
not NOT1 (N2672, N2667);
nor NOR2 (N2673, N2669, N817);
nor NOR4 (N2674, N2664, N1297, N1031, N6);
not NOT1 (N2675, N2672);
and AND2 (N2676, N2658, N1842);
not NOT1 (N2677, N2673);
xor XOR2 (N2678, N2654, N2641);
buf BUF1 (N2679, N2668);
not NOT1 (N2680, N2655);
nor NOR2 (N2681, N2675, N1647);
nor NOR2 (N2682, N2681, N2234);
not NOT1 (N2683, N2676);
or OR3 (N2684, N2642, N1302, N9);
nor NOR4 (N2685, N2684, N2065, N701, N1346);
buf BUF1 (N2686, N2685);
xor XOR2 (N2687, N2671, N1869);
not NOT1 (N2688, N2674);
and AND4 (N2689, N2678, N312, N2290, N98);
and AND2 (N2690, N2677, N2086);
nand NAND2 (N2691, N2682, N1813);
nand NAND3 (N2692, N2691, N2518, N1332);
or OR2 (N2693, N2687, N2529);
nand NAND2 (N2694, N2693, N1990);
xor XOR2 (N2695, N2683, N2516);
buf BUF1 (N2696, N2690);
and AND4 (N2697, N2688, N1013, N1905, N437);
and AND3 (N2698, N2696, N726, N2181);
not NOT1 (N2699, N2679);
nand NAND4 (N2700, N2680, N2558, N78, N2310);
buf BUF1 (N2701, N2689);
and AND4 (N2702, N2698, N219, N333, N2488);
buf BUF1 (N2703, N2702);
or OR2 (N2704, N2647, N981);
nand NAND4 (N2705, N2695, N2602, N995, N1812);
nor NOR3 (N2706, N2700, N2012, N1970);
xor XOR2 (N2707, N2686, N1674);
and AND2 (N2708, N2704, N2410);
nor NOR3 (N2709, N2708, N464, N2223);
not NOT1 (N2710, N2707);
nand NAND2 (N2711, N2703, N2045);
xor XOR2 (N2712, N2711, N6);
nand NAND4 (N2713, N2692, N1747, N2068, N284);
not NOT1 (N2714, N2710);
not NOT1 (N2715, N2714);
nor NOR4 (N2716, N2701, N1373, N2050, N2575);
xor XOR2 (N2717, N2715, N1607);
nand NAND2 (N2718, N2716, N2124);
buf BUF1 (N2719, N2699);
and AND3 (N2720, N2717, N313, N134);
nand NAND3 (N2721, N2705, N607, N2583);
nor NOR3 (N2722, N2706, N2510, N848);
buf BUF1 (N2723, N2718);
buf BUF1 (N2724, N2713);
and AND2 (N2725, N2694, N1333);
nand NAND2 (N2726, N2722, N31);
or OR2 (N2727, N2719, N1688);
nand NAND3 (N2728, N2726, N318, N1433);
or OR2 (N2729, N2709, N1265);
buf BUF1 (N2730, N2723);
nand NAND3 (N2731, N2725, N2429, N2445);
not NOT1 (N2732, N2727);
and AND2 (N2733, N2731, N1032);
nor NOR2 (N2734, N2729, N1259);
not NOT1 (N2735, N2721);
and AND2 (N2736, N2732, N1045);
and AND4 (N2737, N2720, N332, N107, N679);
not NOT1 (N2738, N2724);
nor NOR4 (N2739, N2738, N1580, N2539, N2390);
buf BUF1 (N2740, N2733);
xor XOR2 (N2741, N2740, N2056);
buf BUF1 (N2742, N2697);
not NOT1 (N2743, N2728);
buf BUF1 (N2744, N2735);
and AND3 (N2745, N2742, N2110, N1892);
xor XOR2 (N2746, N2745, N29);
and AND3 (N2747, N2737, N595, N1310);
xor XOR2 (N2748, N2743, N1700);
not NOT1 (N2749, N2712);
xor XOR2 (N2750, N2744, N2578);
nor NOR4 (N2751, N2730, N1902, N1164, N1480);
not NOT1 (N2752, N2751);
or OR4 (N2753, N2750, N2071, N490, N584);
or OR4 (N2754, N2748, N1379, N876, N2691);
not NOT1 (N2755, N2747);
nor NOR2 (N2756, N2753, N1363);
buf BUF1 (N2757, N2734);
buf BUF1 (N2758, N2754);
not NOT1 (N2759, N2752);
not NOT1 (N2760, N2739);
buf BUF1 (N2761, N2749);
nand NAND2 (N2762, N2757, N526);
or OR4 (N2763, N2755, N2352, N2663, N675);
buf BUF1 (N2764, N2763);
nor NOR4 (N2765, N2764, N2364, N313, N1057);
xor XOR2 (N2766, N2761, N1579);
or OR3 (N2767, N2736, N583, N785);
nor NOR4 (N2768, N2767, N2290, N2107, N76);
nand NAND2 (N2769, N2746, N1183);
not NOT1 (N2770, N2769);
buf BUF1 (N2771, N2741);
buf BUF1 (N2772, N2759);
nand NAND4 (N2773, N2768, N707, N2351, N1734);
buf BUF1 (N2774, N2771);
and AND3 (N2775, N2772, N564, N1782);
nor NOR3 (N2776, N2773, N968, N2467);
nand NAND2 (N2777, N2775, N1691);
buf BUF1 (N2778, N2774);
buf BUF1 (N2779, N2762);
nor NOR3 (N2780, N2756, N7, N2688);
and AND3 (N2781, N2780, N2589, N178);
not NOT1 (N2782, N2766);
xor XOR2 (N2783, N2770, N331);
nand NAND4 (N2784, N2779, N545, N464, N1764);
buf BUF1 (N2785, N2781);
or OR3 (N2786, N2784, N1162, N1958);
buf BUF1 (N2787, N2782);
xor XOR2 (N2788, N2785, N374);
not NOT1 (N2789, N2760);
nand NAND2 (N2790, N2777, N2128);
and AND2 (N2791, N2776, N54);
and AND4 (N2792, N2783, N1880, N919, N2035);
nor NOR2 (N2793, N2787, N1232);
not NOT1 (N2794, N2765);
and AND2 (N2795, N2794, N2665);
or OR2 (N2796, N2786, N2032);
buf BUF1 (N2797, N2791);
buf BUF1 (N2798, N2788);
xor XOR2 (N2799, N2789, N1501);
nand NAND3 (N2800, N2758, N839, N577);
and AND3 (N2801, N2799, N2138, N2436);
xor XOR2 (N2802, N2797, N2048);
not NOT1 (N2803, N2795);
and AND4 (N2804, N2778, N415, N1662, N535);
or OR3 (N2805, N2796, N2589, N2202);
buf BUF1 (N2806, N2802);
not NOT1 (N2807, N2801);
nor NOR4 (N2808, N2805, N2484, N2266, N2025);
xor XOR2 (N2809, N2803, N2657);
and AND4 (N2810, N2793, N1612, N2772, N160);
nor NOR4 (N2811, N2810, N2776, N318, N2633);
nor NOR4 (N2812, N2807, N1345, N1815, N629);
buf BUF1 (N2813, N2790);
nand NAND2 (N2814, N2813, N1722);
xor XOR2 (N2815, N2809, N1486);
nor NOR3 (N2816, N2798, N2155, N2052);
and AND2 (N2817, N2792, N1768);
nor NOR2 (N2818, N2816, N2523);
not NOT1 (N2819, N2817);
xor XOR2 (N2820, N2818, N1019);
not NOT1 (N2821, N2812);
and AND2 (N2822, N2819, N713);
and AND4 (N2823, N2806, N1560, N2711, N2756);
and AND2 (N2824, N2814, N2079);
nor NOR4 (N2825, N2815, N1221, N1623, N2747);
and AND2 (N2826, N2820, N2738);
xor XOR2 (N2827, N2823, N1847);
buf BUF1 (N2828, N2827);
buf BUF1 (N2829, N2828);
xor XOR2 (N2830, N2811, N728);
nor NOR3 (N2831, N2824, N229, N980);
xor XOR2 (N2832, N2804, N1350);
nor NOR4 (N2833, N2822, N1144, N60, N928);
buf BUF1 (N2834, N2832);
and AND3 (N2835, N2831, N1444, N1848);
buf BUF1 (N2836, N2808);
nand NAND4 (N2837, N2835, N2388, N1041, N2408);
xor XOR2 (N2838, N2800, N1494);
not NOT1 (N2839, N2830);
not NOT1 (N2840, N2826);
and AND3 (N2841, N2829, N1683, N524);
and AND2 (N2842, N2838, N2399);
buf BUF1 (N2843, N2842);
nand NAND4 (N2844, N2825, N2229, N2190, N159);
or OR3 (N2845, N2841, N250, N2802);
or OR4 (N2846, N2821, N2004, N752, N1559);
nor NOR4 (N2847, N2837, N845, N977, N2682);
and AND3 (N2848, N2844, N1550, N1447);
xor XOR2 (N2849, N2833, N1763);
buf BUF1 (N2850, N2848);
buf BUF1 (N2851, N2847);
buf BUF1 (N2852, N2850);
xor XOR2 (N2853, N2843, N1930);
nand NAND2 (N2854, N2836, N1301);
not NOT1 (N2855, N2834);
buf BUF1 (N2856, N2845);
nor NOR2 (N2857, N2839, N1175);
nor NOR4 (N2858, N2853, N656, N2687, N1487);
xor XOR2 (N2859, N2858, N715);
not NOT1 (N2860, N2840);
nand NAND4 (N2861, N2856, N1811, N2485, N931);
nand NAND2 (N2862, N2849, N2449);
and AND4 (N2863, N2859, N1163, N1448, N720);
and AND3 (N2864, N2857, N813, N626);
nor NOR3 (N2865, N2860, N670, N1918);
or OR4 (N2866, N2854, N332, N532, N2181);
nor NOR3 (N2867, N2846, N1368, N821);
xor XOR2 (N2868, N2852, N1088);
not NOT1 (N2869, N2855);
xor XOR2 (N2870, N2864, N2603);
xor XOR2 (N2871, N2851, N1248);
nor NOR2 (N2872, N2861, N517);
buf BUF1 (N2873, N2863);
xor XOR2 (N2874, N2872, N2862);
xor XOR2 (N2875, N37, N1810);
nor NOR2 (N2876, N2865, N1437);
nand NAND2 (N2877, N2876, N1598);
nor NOR2 (N2878, N2870, N1857);
buf BUF1 (N2879, N2871);
and AND3 (N2880, N2866, N1463, N685);
not NOT1 (N2881, N2868);
nor NOR2 (N2882, N2879, N526);
not NOT1 (N2883, N2881);
xor XOR2 (N2884, N2877, N1970);
nand NAND2 (N2885, N2869, N2759);
and AND3 (N2886, N2875, N1216, N1062);
nand NAND3 (N2887, N2874, N2589, N2554);
and AND4 (N2888, N2873, N720, N612, N79);
nand NAND4 (N2889, N2867, N808, N775, N1548);
or OR2 (N2890, N2880, N2776);
nor NOR2 (N2891, N2887, N2520);
not NOT1 (N2892, N2890);
buf BUF1 (N2893, N2884);
xor XOR2 (N2894, N2891, N993);
or OR2 (N2895, N2889, N301);
not NOT1 (N2896, N2886);
buf BUF1 (N2897, N2892);
buf BUF1 (N2898, N2895);
nor NOR3 (N2899, N2898, N2323, N2044);
buf BUF1 (N2900, N2878);
nor NOR2 (N2901, N2885, N377);
and AND4 (N2902, N2882, N770, N1481, N2081);
nand NAND3 (N2903, N2897, N555, N17);
or OR3 (N2904, N2902, N2149, N1151);
nor NOR3 (N2905, N2901, N1177, N2367);
and AND4 (N2906, N2893, N1493, N895, N1206);
nand NAND4 (N2907, N2903, N515, N2613, N94);
not NOT1 (N2908, N2896);
xor XOR2 (N2909, N2883, N435);
and AND3 (N2910, N2900, N849, N1758);
buf BUF1 (N2911, N2908);
nand NAND3 (N2912, N2906, N2449, N1133);
and AND2 (N2913, N2888, N1303);
not NOT1 (N2914, N2907);
not NOT1 (N2915, N2914);
nand NAND3 (N2916, N2894, N704, N810);
nor NOR2 (N2917, N2904, N663);
or OR2 (N2918, N2911, N1226);
or OR2 (N2919, N2909, N105);
not NOT1 (N2920, N2917);
xor XOR2 (N2921, N2913, N1747);
or OR2 (N2922, N2916, N611);
or OR4 (N2923, N2921, N401, N609, N788);
nand NAND2 (N2924, N2920, N108);
buf BUF1 (N2925, N2905);
xor XOR2 (N2926, N2899, N1988);
nor NOR4 (N2927, N2915, N2801, N1544, N1608);
not NOT1 (N2928, N2918);
nand NAND4 (N2929, N2928, N108, N1882, N2408);
nor NOR2 (N2930, N2926, N1289);
xor XOR2 (N2931, N2925, N1572);
or OR4 (N2932, N2910, N958, N1790, N1347);
not NOT1 (N2933, N2931);
buf BUF1 (N2934, N2927);
nor NOR4 (N2935, N2932, N660, N1644, N653);
nor NOR3 (N2936, N2922, N1055, N1429);
and AND2 (N2937, N2912, N738);
xor XOR2 (N2938, N2919, N2926);
and AND2 (N2939, N2937, N2907);
nor NOR3 (N2940, N2924, N1222, N790);
xor XOR2 (N2941, N2935, N1098);
nand NAND4 (N2942, N2936, N212, N2228, N1954);
nor NOR3 (N2943, N2930, N206, N1464);
nor NOR2 (N2944, N2938, N1320);
and AND4 (N2945, N2943, N2560, N1481, N1789);
buf BUF1 (N2946, N2934);
nor NOR3 (N2947, N2945, N2604, N501);
nor NOR4 (N2948, N2941, N2683, N2257, N28);
nor NOR2 (N2949, N2929, N980);
or OR4 (N2950, N2946, N154, N2892, N2239);
not NOT1 (N2951, N2940);
or OR2 (N2952, N2939, N2444);
and AND2 (N2953, N2944, N1872);
not NOT1 (N2954, N2950);
xor XOR2 (N2955, N2923, N1020);
not NOT1 (N2956, N2952);
and AND3 (N2957, N2947, N328, N2758);
or OR4 (N2958, N2956, N2679, N2081, N2164);
not NOT1 (N2959, N2953);
not NOT1 (N2960, N2933);
not NOT1 (N2961, N2959);
and AND3 (N2962, N2960, N697, N428);
and AND4 (N2963, N2957, N1167, N2592, N2534);
and AND3 (N2964, N2948, N1835, N2493);
and AND4 (N2965, N2962, N1947, N2396, N1936);
or OR4 (N2966, N2963, N347, N2142, N2130);
not NOT1 (N2967, N2961);
nand NAND3 (N2968, N2949, N2689, N1503);
not NOT1 (N2969, N2942);
buf BUF1 (N2970, N2967);
nand NAND4 (N2971, N2955, N1880, N2282, N2278);
not NOT1 (N2972, N2969);
and AND3 (N2973, N2970, N295, N570);
not NOT1 (N2974, N2951);
buf BUF1 (N2975, N2968);
and AND2 (N2976, N2971, N804);
and AND3 (N2977, N2965, N1927, N1733);
not NOT1 (N2978, N2954);
nand NAND3 (N2979, N2974, N1017, N50);
not NOT1 (N2980, N2966);
xor XOR2 (N2981, N2958, N2529);
xor XOR2 (N2982, N2977, N1740);
nand NAND3 (N2983, N2979, N2026, N1975);
and AND3 (N2984, N2976, N1573, N1777);
xor XOR2 (N2985, N2981, N88);
nor NOR3 (N2986, N2980, N730, N2362);
or OR3 (N2987, N2986, N2071, N928);
not NOT1 (N2988, N2982);
xor XOR2 (N2989, N2975, N656);
nand NAND4 (N2990, N2989, N733, N925, N1001);
xor XOR2 (N2991, N2985, N1447);
nand NAND4 (N2992, N2973, N1634, N2474, N2194);
or OR2 (N2993, N2964, N1615);
buf BUF1 (N2994, N2993);
or OR3 (N2995, N2994, N788, N343);
nand NAND3 (N2996, N2987, N1063, N2458);
or OR3 (N2997, N2988, N1838, N2484);
not NOT1 (N2998, N2992);
and AND4 (N2999, N2972, N1093, N925, N214);
nand NAND3 (N3000, N2997, N284, N1509);
not NOT1 (N3001, N2978);
and AND3 (N3002, N2995, N1790, N8);
xor XOR2 (N3003, N2999, N112);
nor NOR3 (N3004, N2998, N366, N442);
xor XOR2 (N3005, N2991, N2988);
not NOT1 (N3006, N2990);
or OR3 (N3007, N3003, N2505, N2420);
and AND3 (N3008, N3007, N2791, N1171);
nor NOR4 (N3009, N3006, N2523, N2071, N2324);
nor NOR3 (N3010, N3001, N2698, N1340);
nor NOR2 (N3011, N3010, N1181);
xor XOR2 (N3012, N3011, N1036);
nand NAND3 (N3013, N3004, N1841, N2518);
not NOT1 (N3014, N3000);
xor XOR2 (N3015, N3009, N2243);
xor XOR2 (N3016, N3005, N1663);
nand NAND3 (N3017, N2984, N1686, N1051);
nor NOR2 (N3018, N3012, N1431);
buf BUF1 (N3019, N3016);
endmodule