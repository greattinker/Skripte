// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;

output N4014,N4015,N4017,N4006,N4016,N4003,N3989,N3995,N4008,N4018;

or OR2 (N19, N2, N4);
nand NAND3 (N20, N18, N17, N2);
not NOT1 (N21, N1);
xor XOR2 (N22, N17, N15);
xor XOR2 (N23, N7, N13);
and AND4 (N24, N5, N6, N16, N18);
xor XOR2 (N25, N7, N14);
not NOT1 (N26, N18);
buf BUF1 (N27, N15);
nand NAND3 (N28, N25, N4, N26);
or OR4 (N29, N7, N18, N21, N16);
not NOT1 (N30, N17);
buf BUF1 (N31, N16);
xor XOR2 (N32, N24, N10);
or OR2 (N33, N32, N30);
xor XOR2 (N34, N4, N14);
or OR3 (N35, N27, N19, N8);
nand NAND4 (N36, N11, N3, N30, N34);
not NOT1 (N37, N33);
nand NAND3 (N38, N9, N22, N29);
xor XOR2 (N39, N32, N18);
or OR4 (N40, N2, N2, N3, N19);
not NOT1 (N41, N31);
or OR3 (N42, N39, N18, N39);
xor XOR2 (N43, N40, N15);
nor NOR3 (N44, N20, N14, N29);
nor NOR2 (N45, N43, N28);
buf BUF1 (N46, N11);
xor XOR2 (N47, N46, N43);
and AND2 (N48, N45, N22);
and AND3 (N49, N48, N28, N43);
and AND3 (N50, N42, N23, N18);
nor NOR4 (N51, N12, N12, N20, N5);
nand NAND3 (N52, N49, N10, N13);
nand NAND3 (N53, N44, N42, N18);
or OR4 (N54, N52, N41, N23, N29);
nor NOR3 (N55, N52, N45, N24);
buf BUF1 (N56, N36);
nor NOR3 (N57, N47, N4, N20);
nor NOR4 (N58, N50, N49, N47, N30);
nand NAND4 (N59, N58, N11, N47, N56);
and AND3 (N60, N1, N17, N24);
buf BUF1 (N61, N57);
and AND4 (N62, N53, N5, N55, N26);
not NOT1 (N63, N36);
nand NAND3 (N64, N37, N61, N57);
nand NAND4 (N65, N55, N14, N56, N9);
nor NOR3 (N66, N35, N41, N56);
buf BUF1 (N67, N59);
nor NOR3 (N68, N67, N56, N6);
nand NAND2 (N69, N66, N48);
or OR4 (N70, N63, N16, N13, N42);
not NOT1 (N71, N51);
xor XOR2 (N72, N70, N21);
buf BUF1 (N73, N71);
not NOT1 (N74, N68);
xor XOR2 (N75, N64, N27);
not NOT1 (N76, N60);
nor NOR4 (N77, N76, N64, N26, N54);
or OR2 (N78, N25, N47);
nor NOR2 (N79, N77, N30);
nor NOR4 (N80, N74, N34, N51, N60);
not NOT1 (N81, N79);
nand NAND2 (N82, N69, N14);
nor NOR2 (N83, N65, N4);
or OR3 (N84, N81, N56, N56);
xor XOR2 (N85, N72, N75);
not NOT1 (N86, N42);
not NOT1 (N87, N62);
buf BUF1 (N88, N87);
nor NOR3 (N89, N80, N13, N59);
and AND3 (N90, N78, N9, N16);
buf BUF1 (N91, N89);
nand NAND3 (N92, N83, N10, N89);
or OR4 (N93, N38, N31, N40, N39);
nand NAND3 (N94, N73, N63, N61);
buf BUF1 (N95, N85);
xor XOR2 (N96, N88, N53);
and AND3 (N97, N93, N73, N33);
nor NOR3 (N98, N91, N13, N52);
or OR2 (N99, N95, N36);
xor XOR2 (N100, N94, N10);
xor XOR2 (N101, N82, N22);
and AND4 (N102, N84, N53, N4, N63);
and AND4 (N103, N96, N26, N4, N71);
nor NOR4 (N104, N103, N93, N11, N83);
xor XOR2 (N105, N97, N37);
xor XOR2 (N106, N98, N2);
buf BUF1 (N107, N92);
nand NAND2 (N108, N90, N100);
xor XOR2 (N109, N60, N48);
nand NAND3 (N110, N106, N31, N82);
nor NOR3 (N111, N105, N76, N83);
nor NOR4 (N112, N107, N72, N59, N28);
and AND4 (N113, N112, N33, N42, N88);
not NOT1 (N114, N101);
nand NAND4 (N115, N110, N29, N100, N49);
nor NOR4 (N116, N86, N104, N25, N107);
nand NAND2 (N117, N17, N5);
xor XOR2 (N118, N113, N47);
buf BUF1 (N119, N102);
nor NOR3 (N120, N117, N48, N11);
not NOT1 (N121, N114);
or OR2 (N122, N109, N88);
xor XOR2 (N123, N111, N90);
and AND3 (N124, N123, N68, N30);
and AND4 (N125, N116, N34, N52, N76);
buf BUF1 (N126, N108);
or OR4 (N127, N99, N89, N86, N125);
buf BUF1 (N128, N11);
buf BUF1 (N129, N124);
or OR4 (N130, N120, N120, N64, N128);
buf BUF1 (N131, N94);
and AND2 (N132, N121, N45);
not NOT1 (N133, N115);
not NOT1 (N134, N133);
buf BUF1 (N135, N127);
nand NAND2 (N136, N130, N127);
or OR3 (N137, N119, N71, N78);
or OR2 (N138, N136, N2);
not NOT1 (N139, N132);
nand NAND4 (N140, N138, N116, N3, N22);
and AND2 (N141, N122, N88);
and AND2 (N142, N131, N30);
xor XOR2 (N143, N139, N88);
not NOT1 (N144, N142);
xor XOR2 (N145, N126, N6);
not NOT1 (N146, N143);
not NOT1 (N147, N129);
not NOT1 (N148, N141);
not NOT1 (N149, N148);
xor XOR2 (N150, N134, N84);
buf BUF1 (N151, N145);
nand NAND2 (N152, N144, N3);
xor XOR2 (N153, N118, N140);
nor NOR2 (N154, N56, N6);
nor NOR2 (N155, N147, N62);
buf BUF1 (N156, N151);
xor XOR2 (N157, N149, N77);
nand NAND3 (N158, N156, N112, N153);
and AND3 (N159, N107, N6, N105);
and AND2 (N160, N154, N50);
or OR2 (N161, N135, N122);
xor XOR2 (N162, N146, N117);
and AND3 (N163, N152, N58, N60);
xor XOR2 (N164, N137, N29);
nand NAND3 (N165, N162, N130, N151);
xor XOR2 (N166, N159, N156);
xor XOR2 (N167, N157, N6);
buf BUF1 (N168, N155);
not NOT1 (N169, N161);
or OR3 (N170, N163, N58, N147);
xor XOR2 (N171, N164, N109);
not NOT1 (N172, N168);
nand NAND2 (N173, N150, N58);
or OR2 (N174, N169, N6);
xor XOR2 (N175, N166, N12);
and AND3 (N176, N167, N115, N123);
nor NOR3 (N177, N160, N162, N4);
xor XOR2 (N178, N174, N144);
nor NOR2 (N179, N170, N156);
nand NAND2 (N180, N175, N64);
and AND2 (N181, N173, N115);
buf BUF1 (N182, N176);
not NOT1 (N183, N180);
xor XOR2 (N184, N165, N79);
nor NOR2 (N185, N183, N117);
buf BUF1 (N186, N178);
or OR2 (N187, N181, N27);
nand NAND4 (N188, N158, N154, N88, N171);
nand NAND2 (N189, N29, N163);
nand NAND4 (N190, N179, N50, N27, N158);
and AND4 (N191, N177, N165, N9, N37);
nor NOR3 (N192, N189, N50, N86);
not NOT1 (N193, N172);
xor XOR2 (N194, N192, N105);
buf BUF1 (N195, N185);
and AND2 (N196, N186, N3);
xor XOR2 (N197, N184, N53);
xor XOR2 (N198, N193, N122);
buf BUF1 (N199, N198);
not NOT1 (N200, N197);
nand NAND2 (N201, N191, N127);
and AND3 (N202, N182, N103, N146);
or OR4 (N203, N196, N120, N156, N80);
nand NAND4 (N204, N194, N152, N11, N84);
or OR4 (N205, N203, N78, N90, N47);
or OR4 (N206, N188, N165, N9, N58);
and AND4 (N207, N190, N40, N122, N127);
nor NOR2 (N208, N206, N159);
buf BUF1 (N209, N187);
nand NAND4 (N210, N204, N23, N92, N198);
nor NOR4 (N211, N209, N8, N48, N94);
or OR4 (N212, N199, N173, N104, N110);
nor NOR2 (N213, N210, N117);
nand NAND3 (N214, N207, N16, N25);
nand NAND3 (N215, N208, N11, N155);
and AND4 (N216, N213, N28, N26, N168);
buf BUF1 (N217, N195);
and AND2 (N218, N216, N9);
or OR3 (N219, N218, N67, N41);
buf BUF1 (N220, N217);
or OR3 (N221, N215, N84, N201);
not NOT1 (N222, N131);
xor XOR2 (N223, N200, N120);
buf BUF1 (N224, N222);
nand NAND3 (N225, N212, N215, N111);
not NOT1 (N226, N220);
not NOT1 (N227, N202);
or OR2 (N228, N205, N52);
not NOT1 (N229, N226);
buf BUF1 (N230, N219);
nand NAND2 (N231, N214, N133);
buf BUF1 (N232, N228);
buf BUF1 (N233, N230);
nand NAND3 (N234, N225, N181, N190);
nand NAND3 (N235, N223, N145, N174);
not NOT1 (N236, N232);
buf BUF1 (N237, N229);
not NOT1 (N238, N237);
or OR2 (N239, N235, N3);
not NOT1 (N240, N211);
xor XOR2 (N241, N240, N4);
buf BUF1 (N242, N239);
and AND4 (N243, N238, N233, N32, N223);
or OR4 (N244, N179, N208, N64, N13);
or OR2 (N245, N243, N106);
nand NAND4 (N246, N224, N29, N123, N56);
nor NOR2 (N247, N246, N62);
buf BUF1 (N248, N221);
buf BUF1 (N249, N227);
and AND2 (N250, N247, N200);
nand NAND4 (N251, N244, N17, N164, N45);
nor NOR4 (N252, N231, N54, N232, N172);
buf BUF1 (N253, N245);
and AND3 (N254, N253, N232, N211);
nand NAND4 (N255, N236, N13, N129, N46);
not NOT1 (N256, N241);
xor XOR2 (N257, N242, N61);
not NOT1 (N258, N252);
nor NOR2 (N259, N249, N254);
nor NOR4 (N260, N258, N49, N189, N204);
and AND3 (N261, N146, N137, N85);
nand NAND2 (N262, N250, N217);
not NOT1 (N263, N251);
not NOT1 (N264, N248);
or OR2 (N265, N257, N10);
buf BUF1 (N266, N264);
not NOT1 (N267, N256);
and AND3 (N268, N261, N230, N265);
or OR2 (N269, N69, N141);
xor XOR2 (N270, N263, N229);
buf BUF1 (N271, N260);
or OR4 (N272, N259, N247, N153, N54);
nor NOR4 (N273, N234, N154, N127, N85);
not NOT1 (N274, N267);
nand NAND3 (N275, N271, N196, N132);
not NOT1 (N276, N272);
and AND4 (N277, N270, N30, N127, N73);
not NOT1 (N278, N255);
xor XOR2 (N279, N262, N99);
and AND4 (N280, N269, N79, N160, N133);
and AND2 (N281, N278, N38);
or OR4 (N282, N280, N185, N228, N75);
buf BUF1 (N283, N276);
nand NAND4 (N284, N273, N132, N261, N173);
not NOT1 (N285, N283);
and AND2 (N286, N268, N168);
not NOT1 (N287, N281);
buf BUF1 (N288, N286);
buf BUF1 (N289, N285);
or OR3 (N290, N275, N76, N161);
xor XOR2 (N291, N288, N55);
nor NOR2 (N292, N284, N118);
nor NOR4 (N293, N274, N5, N198, N287);
not NOT1 (N294, N207);
or OR3 (N295, N293, N228, N87);
nand NAND2 (N296, N289, N99);
not NOT1 (N297, N279);
buf BUF1 (N298, N266);
nor NOR4 (N299, N277, N172, N164, N137);
nand NAND4 (N300, N295, N122, N207, N226);
nor NOR2 (N301, N291, N260);
nor NOR4 (N302, N296, N103, N14, N181);
nor NOR2 (N303, N282, N24);
or OR2 (N304, N294, N287);
xor XOR2 (N305, N299, N296);
nand NAND4 (N306, N302, N133, N268, N158);
buf BUF1 (N307, N304);
buf BUF1 (N308, N290);
nand NAND2 (N309, N301, N229);
xor XOR2 (N310, N292, N142);
buf BUF1 (N311, N305);
nor NOR2 (N312, N306, N143);
xor XOR2 (N313, N309, N68);
nand NAND4 (N314, N307, N202, N48, N306);
not NOT1 (N315, N310);
xor XOR2 (N316, N308, N214);
xor XOR2 (N317, N315, N36);
nand NAND3 (N318, N314, N114, N287);
buf BUF1 (N319, N298);
nor NOR4 (N320, N317, N216, N46, N299);
or OR3 (N321, N318, N310, N40);
buf BUF1 (N322, N313);
nor NOR4 (N323, N322, N71, N257, N248);
nand NAND2 (N324, N321, N100);
buf BUF1 (N325, N324);
nand NAND3 (N326, N320, N32, N189);
not NOT1 (N327, N311);
xor XOR2 (N328, N323, N297);
nor NOR3 (N329, N273, N211, N306);
and AND2 (N330, N328, N16);
not NOT1 (N331, N312);
nand NAND4 (N332, N319, N10, N70, N316);
and AND2 (N333, N289, N285);
buf BUF1 (N334, N325);
xor XOR2 (N335, N332, N99);
xor XOR2 (N336, N300, N256);
not NOT1 (N337, N335);
nor NOR2 (N338, N303, N213);
or OR2 (N339, N331, N90);
buf BUF1 (N340, N337);
xor XOR2 (N341, N327, N281);
xor XOR2 (N342, N336, N235);
not NOT1 (N343, N342);
xor XOR2 (N344, N329, N93);
and AND4 (N345, N339, N156, N263, N69);
nand NAND3 (N346, N333, N206, N322);
nor NOR3 (N347, N344, N31, N255);
or OR3 (N348, N347, N118, N279);
nor NOR4 (N349, N334, N204, N250, N48);
nand NAND3 (N350, N346, N215, N271);
nand NAND4 (N351, N350, N101, N305, N100);
or OR4 (N352, N338, N152, N58, N108);
xor XOR2 (N353, N352, N37);
nor NOR3 (N354, N330, N9, N284);
nor NOR2 (N355, N326, N192);
nand NAND3 (N356, N353, N119, N45);
xor XOR2 (N357, N349, N257);
buf BUF1 (N358, N345);
buf BUF1 (N359, N343);
and AND4 (N360, N355, N215, N349, N26);
nand NAND2 (N361, N340, N298);
buf BUF1 (N362, N354);
nand NAND4 (N363, N356, N139, N352, N133);
xor XOR2 (N364, N360, N7);
or OR3 (N365, N348, N214, N33);
nand NAND3 (N366, N357, N148, N26);
nor NOR3 (N367, N365, N9, N215);
not NOT1 (N368, N359);
nor NOR2 (N369, N351, N250);
nor NOR4 (N370, N367, N241, N344, N280);
nor NOR4 (N371, N362, N21, N180, N100);
nor NOR4 (N372, N369, N70, N244, N80);
buf BUF1 (N373, N372);
not NOT1 (N374, N371);
or OR2 (N375, N368, N154);
xor XOR2 (N376, N370, N178);
nand NAND3 (N377, N358, N111, N268);
nand NAND3 (N378, N341, N108, N11);
nand NAND3 (N379, N361, N103, N309);
buf BUF1 (N380, N374);
xor XOR2 (N381, N375, N223);
not NOT1 (N382, N381);
nand NAND3 (N383, N373, N172, N356);
nor NOR4 (N384, N364, N142, N206, N272);
nor NOR3 (N385, N384, N361, N263);
not NOT1 (N386, N379);
xor XOR2 (N387, N376, N182);
nor NOR3 (N388, N386, N40, N315);
nand NAND3 (N389, N366, N33, N252);
nand NAND3 (N390, N385, N149, N353);
buf BUF1 (N391, N377);
xor XOR2 (N392, N389, N352);
nand NAND2 (N393, N391, N33);
and AND3 (N394, N363, N349, N319);
and AND2 (N395, N380, N170);
buf BUF1 (N396, N390);
nand NAND3 (N397, N392, N133, N25);
not NOT1 (N398, N387);
and AND4 (N399, N378, N22, N322, N80);
or OR2 (N400, N396, N310);
and AND4 (N401, N399, N312, N73, N269);
not NOT1 (N402, N398);
xor XOR2 (N403, N393, N352);
and AND2 (N404, N403, N119);
nand NAND2 (N405, N397, N185);
or OR2 (N406, N401, N316);
or OR4 (N407, N395, N57, N44, N181);
not NOT1 (N408, N383);
xor XOR2 (N409, N405, N332);
or OR3 (N410, N400, N164, N146);
nand NAND2 (N411, N407, N315);
buf BUF1 (N412, N409);
not NOT1 (N413, N411);
and AND3 (N414, N413, N247, N214);
or OR3 (N415, N404, N132, N253);
buf BUF1 (N416, N402);
xor XOR2 (N417, N408, N317);
or OR4 (N418, N417, N180, N130, N103);
xor XOR2 (N419, N406, N58);
xor XOR2 (N420, N394, N258);
xor XOR2 (N421, N420, N148);
not NOT1 (N422, N382);
or OR4 (N423, N418, N342, N371, N87);
and AND3 (N424, N414, N86, N100);
or OR2 (N425, N424, N249);
and AND4 (N426, N415, N397, N132, N292);
nand NAND3 (N427, N412, N83, N13);
not NOT1 (N428, N388);
nand NAND4 (N429, N423, N328, N135, N292);
nor NOR4 (N430, N426, N293, N360, N28);
nor NOR3 (N431, N430, N24, N379);
nand NAND3 (N432, N419, N104, N75);
xor XOR2 (N433, N429, N353);
nand NAND3 (N434, N410, N152, N73);
not NOT1 (N435, N433);
nor NOR2 (N436, N432, N228);
nand NAND2 (N437, N427, N49);
nor NOR2 (N438, N436, N153);
buf BUF1 (N439, N416);
and AND4 (N440, N421, N285, N142, N419);
not NOT1 (N441, N435);
nand NAND3 (N442, N434, N122, N198);
xor XOR2 (N443, N428, N386);
nand NAND4 (N444, N431, N66, N335, N274);
and AND2 (N445, N425, N58);
buf BUF1 (N446, N445);
nand NAND4 (N447, N438, N433, N323, N273);
or OR2 (N448, N442, N266);
nor NOR2 (N449, N439, N447);
buf BUF1 (N450, N160);
xor XOR2 (N451, N449, N45);
or OR4 (N452, N450, N139, N426, N106);
buf BUF1 (N453, N422);
nand NAND4 (N454, N452, N96, N26, N291);
buf BUF1 (N455, N448);
not NOT1 (N456, N441);
and AND3 (N457, N440, N399, N34);
not NOT1 (N458, N437);
buf BUF1 (N459, N456);
xor XOR2 (N460, N444, N387);
not NOT1 (N461, N459);
buf BUF1 (N462, N454);
xor XOR2 (N463, N451, N190);
xor XOR2 (N464, N455, N433);
nand NAND2 (N465, N463, N464);
nor NOR3 (N466, N100, N226, N41);
xor XOR2 (N467, N461, N216);
xor XOR2 (N468, N465, N420);
xor XOR2 (N469, N467, N219);
xor XOR2 (N470, N462, N158);
not NOT1 (N471, N460);
nor NOR2 (N472, N470, N248);
nor NOR3 (N473, N471, N313, N304);
or OR3 (N474, N472, N313, N391);
not NOT1 (N475, N468);
not NOT1 (N476, N443);
buf BUF1 (N477, N476);
nand NAND3 (N478, N453, N338, N47);
nand NAND4 (N479, N474, N226, N245, N189);
buf BUF1 (N480, N475);
not NOT1 (N481, N478);
nor NOR3 (N482, N480, N315, N173);
nor NOR3 (N483, N479, N90, N154);
nand NAND2 (N484, N483, N401);
nand NAND3 (N485, N482, N243, N299);
and AND4 (N486, N457, N384, N120, N326);
or OR3 (N487, N477, N271, N312);
not NOT1 (N488, N466);
buf BUF1 (N489, N446);
nand NAND3 (N490, N484, N48, N166);
nand NAND2 (N491, N490, N329);
or OR2 (N492, N486, N125);
not NOT1 (N493, N481);
xor XOR2 (N494, N473, N402);
nand NAND3 (N495, N491, N130, N437);
not NOT1 (N496, N489);
xor XOR2 (N497, N469, N362);
nor NOR2 (N498, N494, N47);
or OR2 (N499, N458, N385);
buf BUF1 (N500, N495);
xor XOR2 (N501, N496, N408);
and AND3 (N502, N500, N321, N144);
and AND2 (N503, N502, N165);
and AND3 (N504, N493, N283, N246);
nor NOR4 (N505, N498, N490, N374, N378);
xor XOR2 (N506, N499, N40);
and AND2 (N507, N485, N249);
nor NOR3 (N508, N506, N115, N53);
and AND2 (N509, N487, N456);
xor XOR2 (N510, N488, N256);
xor XOR2 (N511, N510, N475);
nor NOR2 (N512, N511, N13);
nand NAND2 (N513, N512, N207);
xor XOR2 (N514, N513, N195);
not NOT1 (N515, N508);
and AND3 (N516, N509, N51, N458);
buf BUF1 (N517, N507);
not NOT1 (N518, N504);
or OR2 (N519, N505, N466);
and AND3 (N520, N517, N167, N418);
nor NOR3 (N521, N518, N469, N326);
or OR2 (N522, N497, N459);
xor XOR2 (N523, N522, N306);
nand NAND4 (N524, N503, N176, N89, N475);
or OR2 (N525, N515, N189);
nand NAND2 (N526, N523, N44);
not NOT1 (N527, N492);
nor NOR3 (N528, N514, N251, N419);
nor NOR3 (N529, N516, N506, N156);
not NOT1 (N530, N525);
xor XOR2 (N531, N529, N160);
not NOT1 (N532, N527);
not NOT1 (N533, N524);
nand NAND4 (N534, N526, N76, N134, N518);
nor NOR2 (N535, N534, N479);
not NOT1 (N536, N535);
xor XOR2 (N537, N520, N292);
and AND3 (N538, N528, N265, N18);
or OR4 (N539, N537, N168, N101, N366);
xor XOR2 (N540, N531, N451);
or OR2 (N541, N538, N179);
or OR4 (N542, N532, N19, N364, N338);
or OR3 (N543, N539, N538, N200);
buf BUF1 (N544, N540);
nand NAND4 (N545, N544, N342, N506, N445);
nand NAND4 (N546, N519, N257, N193, N112);
and AND4 (N547, N542, N242, N415, N64);
not NOT1 (N548, N530);
buf BUF1 (N549, N541);
nand NAND3 (N550, N549, N138, N451);
buf BUF1 (N551, N533);
and AND3 (N552, N550, N268, N462);
and AND4 (N553, N551, N420, N546, N135);
buf BUF1 (N554, N379);
buf BUF1 (N555, N552);
nor NOR4 (N556, N548, N315, N409, N326);
xor XOR2 (N557, N554, N438);
nor NOR2 (N558, N553, N271);
and AND2 (N559, N543, N163);
nor NOR3 (N560, N559, N481, N406);
or OR3 (N561, N545, N396, N10);
buf BUF1 (N562, N555);
nor NOR4 (N563, N558, N559, N38, N522);
or OR2 (N564, N547, N466);
and AND4 (N565, N521, N554, N113, N445);
xor XOR2 (N566, N563, N366);
xor XOR2 (N567, N560, N265);
nand NAND3 (N568, N565, N243, N246);
buf BUF1 (N569, N556);
not NOT1 (N570, N561);
nand NAND2 (N571, N567, N446);
nand NAND3 (N572, N568, N82, N345);
nor NOR3 (N573, N566, N522, N442);
not NOT1 (N574, N573);
buf BUF1 (N575, N501);
buf BUF1 (N576, N575);
nand NAND4 (N577, N569, N426, N293, N314);
or OR4 (N578, N557, N258, N84, N84);
or OR3 (N579, N578, N203, N131);
xor XOR2 (N580, N571, N442);
nand NAND4 (N581, N570, N182, N126, N175);
xor XOR2 (N582, N574, N326);
not NOT1 (N583, N579);
xor XOR2 (N584, N536, N56);
or OR4 (N585, N582, N98, N453, N511);
xor XOR2 (N586, N585, N324);
or OR3 (N587, N564, N361, N250);
buf BUF1 (N588, N586);
nor NOR4 (N589, N588, N435, N190, N29);
nand NAND2 (N590, N581, N263);
nand NAND2 (N591, N580, N426);
buf BUF1 (N592, N576);
nor NOR3 (N593, N577, N45, N408);
buf BUF1 (N594, N591);
xor XOR2 (N595, N584, N397);
not NOT1 (N596, N590);
nand NAND4 (N597, N593, N27, N84, N103);
xor XOR2 (N598, N596, N313);
or OR2 (N599, N592, N225);
not NOT1 (N600, N595);
buf BUF1 (N601, N562);
and AND4 (N602, N601, N579, N53, N155);
nand NAND4 (N603, N594, N413, N6, N269);
or OR2 (N604, N600, N353);
and AND4 (N605, N597, N45, N291, N2);
nand NAND3 (N606, N587, N40, N287);
or OR2 (N607, N605, N132);
not NOT1 (N608, N606);
buf BUF1 (N609, N572);
and AND2 (N610, N607, N555);
not NOT1 (N611, N598);
xor XOR2 (N612, N599, N486);
xor XOR2 (N613, N610, N164);
buf BUF1 (N614, N604);
or OR3 (N615, N602, N217, N418);
or OR3 (N616, N614, N92, N234);
nor NOR3 (N617, N603, N284, N89);
nor NOR2 (N618, N611, N332);
or OR3 (N619, N615, N430, N5);
and AND4 (N620, N613, N446, N414, N564);
or OR3 (N621, N589, N355, N583);
or OR2 (N622, N41, N313);
or OR4 (N623, N620, N483, N198, N164);
and AND2 (N624, N609, N70);
nand NAND4 (N625, N618, N7, N461, N175);
not NOT1 (N626, N623);
or OR4 (N627, N622, N38, N455, N308);
nor NOR4 (N628, N619, N447, N429, N104);
nand NAND3 (N629, N627, N384, N109);
or OR4 (N630, N617, N603, N390, N82);
xor XOR2 (N631, N621, N247);
and AND2 (N632, N631, N159);
xor XOR2 (N633, N628, N433);
nand NAND3 (N634, N630, N243, N280);
nor NOR3 (N635, N633, N331, N58);
not NOT1 (N636, N632);
or OR4 (N637, N608, N271, N472, N468);
nor NOR3 (N638, N636, N49, N53);
or OR4 (N639, N626, N243, N310, N513);
xor XOR2 (N640, N634, N82);
not NOT1 (N641, N635);
or OR3 (N642, N616, N541, N295);
not NOT1 (N643, N642);
not NOT1 (N644, N640);
buf BUF1 (N645, N629);
nand NAND2 (N646, N645, N13);
buf BUF1 (N647, N624);
nor NOR4 (N648, N612, N569, N617, N225);
nor NOR2 (N649, N644, N621);
buf BUF1 (N650, N638);
not NOT1 (N651, N647);
nand NAND3 (N652, N649, N525, N281);
or OR4 (N653, N639, N136, N597, N247);
buf BUF1 (N654, N652);
nor NOR2 (N655, N637, N65);
not NOT1 (N656, N625);
buf BUF1 (N657, N653);
xor XOR2 (N658, N650, N197);
xor XOR2 (N659, N641, N110);
xor XOR2 (N660, N651, N189);
not NOT1 (N661, N648);
or OR2 (N662, N661, N333);
xor XOR2 (N663, N659, N431);
nor NOR3 (N664, N646, N422, N81);
nand NAND4 (N665, N657, N57, N571, N445);
or OR3 (N666, N663, N83, N540);
buf BUF1 (N667, N665);
or OR3 (N668, N654, N494, N477);
xor XOR2 (N669, N667, N391);
nor NOR4 (N670, N666, N272, N315, N189);
nand NAND2 (N671, N656, N470);
buf BUF1 (N672, N660);
buf BUF1 (N673, N669);
nand NAND4 (N674, N671, N46, N328, N529);
nor NOR3 (N675, N674, N668, N504);
nor NOR3 (N676, N509, N632, N627);
and AND4 (N677, N670, N510, N508, N151);
xor XOR2 (N678, N673, N356);
buf BUF1 (N679, N676);
and AND4 (N680, N678, N180, N481, N435);
not NOT1 (N681, N643);
and AND2 (N682, N655, N552);
nand NAND2 (N683, N679, N293);
or OR2 (N684, N683, N571);
nand NAND4 (N685, N658, N661, N493, N138);
buf BUF1 (N686, N662);
buf BUF1 (N687, N682);
nor NOR2 (N688, N681, N371);
not NOT1 (N689, N672);
not NOT1 (N690, N675);
xor XOR2 (N691, N686, N420);
nand NAND2 (N692, N664, N25);
and AND4 (N693, N680, N156, N271, N202);
nand NAND3 (N694, N677, N578, N204);
buf BUF1 (N695, N691);
or OR2 (N696, N690, N302);
or OR4 (N697, N693, N528, N303, N246);
nor NOR3 (N698, N687, N541, N546);
or OR4 (N699, N689, N509, N635, N271);
not NOT1 (N700, N694);
nand NAND4 (N701, N692, N554, N264, N653);
not NOT1 (N702, N696);
nand NAND3 (N703, N702, N521, N369);
or OR3 (N704, N699, N339, N563);
not NOT1 (N705, N685);
buf BUF1 (N706, N684);
xor XOR2 (N707, N700, N575);
or OR4 (N708, N704, N691, N13, N299);
not NOT1 (N709, N701);
nand NAND2 (N710, N706, N206);
xor XOR2 (N711, N697, N645);
xor XOR2 (N712, N703, N250);
xor XOR2 (N713, N710, N496);
buf BUF1 (N714, N707);
nor NOR2 (N715, N705, N303);
nand NAND4 (N716, N708, N350, N154, N66);
or OR4 (N717, N688, N656, N504, N360);
buf BUF1 (N718, N714);
not NOT1 (N719, N717);
nor NOR3 (N720, N711, N263, N285);
nand NAND3 (N721, N713, N701, N525);
or OR4 (N722, N715, N483, N573, N585);
or OR4 (N723, N718, N257, N605, N629);
and AND3 (N724, N722, N67, N197);
nor NOR2 (N725, N712, N670);
buf BUF1 (N726, N709);
nor NOR2 (N727, N721, N594);
buf BUF1 (N728, N724);
nand NAND2 (N729, N698, N97);
xor XOR2 (N730, N716, N571);
or OR4 (N731, N725, N479, N177, N269);
and AND3 (N732, N731, N691, N3);
nand NAND4 (N733, N728, N664, N97, N9);
buf BUF1 (N734, N732);
xor XOR2 (N735, N730, N162);
and AND4 (N736, N720, N631, N351, N14);
not NOT1 (N737, N729);
xor XOR2 (N738, N733, N645);
not NOT1 (N739, N695);
or OR4 (N740, N735, N233, N61, N588);
nand NAND2 (N741, N739, N302);
xor XOR2 (N742, N736, N732);
not NOT1 (N743, N719);
or OR4 (N744, N737, N520, N484, N288);
nor NOR2 (N745, N740, N445);
xor XOR2 (N746, N726, N41);
nand NAND2 (N747, N738, N287);
nand NAND4 (N748, N723, N661, N90, N659);
or OR4 (N749, N741, N54, N80, N357);
not NOT1 (N750, N748);
not NOT1 (N751, N745);
xor XOR2 (N752, N742, N382);
buf BUF1 (N753, N749);
nor NOR2 (N754, N751, N154);
xor XOR2 (N755, N747, N592);
buf BUF1 (N756, N753);
buf BUF1 (N757, N727);
nand NAND2 (N758, N754, N540);
buf BUF1 (N759, N758);
and AND3 (N760, N756, N68, N446);
nor NOR4 (N761, N734, N36, N351, N517);
buf BUF1 (N762, N757);
buf BUF1 (N763, N761);
nor NOR2 (N764, N746, N752);
buf BUF1 (N765, N568);
or OR4 (N766, N762, N242, N671, N394);
nor NOR3 (N767, N755, N130, N87);
nor NOR2 (N768, N744, N85);
not NOT1 (N769, N760);
xor XOR2 (N770, N759, N7);
nand NAND3 (N771, N767, N58, N403);
and AND4 (N772, N769, N509, N275, N558);
nor NOR2 (N773, N763, N524);
or OR2 (N774, N772, N172);
not NOT1 (N775, N768);
xor XOR2 (N776, N774, N739);
xor XOR2 (N777, N766, N181);
or OR2 (N778, N773, N586);
or OR2 (N779, N765, N343);
xor XOR2 (N780, N777, N599);
not NOT1 (N781, N764);
nor NOR3 (N782, N780, N570, N313);
xor XOR2 (N783, N775, N657);
nand NAND4 (N784, N750, N327, N58, N727);
nor NOR2 (N785, N743, N114);
xor XOR2 (N786, N779, N440);
and AND2 (N787, N776, N236);
not NOT1 (N788, N782);
not NOT1 (N789, N783);
nor NOR2 (N790, N787, N157);
nor NOR4 (N791, N785, N711, N684, N539);
not NOT1 (N792, N781);
xor XOR2 (N793, N770, N457);
and AND2 (N794, N786, N177);
xor XOR2 (N795, N790, N407);
and AND3 (N796, N791, N757, N637);
or OR2 (N797, N792, N149);
nand NAND2 (N798, N793, N792);
nand NAND4 (N799, N784, N189, N622, N455);
not NOT1 (N800, N795);
nor NOR3 (N801, N796, N305, N87);
or OR3 (N802, N789, N689, N771);
nand NAND4 (N803, N44, N195, N423, N643);
nand NAND3 (N804, N797, N217, N234);
xor XOR2 (N805, N798, N81);
not NOT1 (N806, N778);
not NOT1 (N807, N806);
and AND4 (N808, N801, N151, N721, N778);
nor NOR3 (N809, N807, N523, N127);
not NOT1 (N810, N800);
or OR3 (N811, N803, N47, N611);
xor XOR2 (N812, N805, N625);
or OR4 (N813, N812, N176, N648, N403);
nor NOR2 (N814, N810, N228);
xor XOR2 (N815, N813, N468);
and AND4 (N816, N815, N468, N25, N418);
and AND2 (N817, N809, N290);
buf BUF1 (N818, N788);
nand NAND3 (N819, N802, N622, N659);
or OR4 (N820, N799, N475, N295, N66);
xor XOR2 (N821, N820, N724);
nor NOR4 (N822, N808, N200, N416, N27);
or OR3 (N823, N822, N771, N368);
buf BUF1 (N824, N811);
and AND3 (N825, N821, N606, N500);
buf BUF1 (N826, N818);
nand NAND3 (N827, N826, N597, N65);
or OR2 (N828, N794, N618);
and AND3 (N829, N823, N817, N641);
or OR3 (N830, N734, N33, N211);
buf BUF1 (N831, N816);
and AND4 (N832, N825, N765, N305, N252);
nand NAND3 (N833, N828, N716, N470);
or OR2 (N834, N833, N462);
buf BUF1 (N835, N804);
nor NOR2 (N836, N832, N644);
buf BUF1 (N837, N819);
nand NAND3 (N838, N827, N2, N138);
xor XOR2 (N839, N830, N584);
xor XOR2 (N840, N836, N196);
xor XOR2 (N841, N839, N153);
xor XOR2 (N842, N841, N249);
buf BUF1 (N843, N831);
not NOT1 (N844, N842);
xor XOR2 (N845, N843, N262);
xor XOR2 (N846, N840, N745);
and AND2 (N847, N829, N663);
and AND4 (N848, N844, N486, N646, N460);
or OR3 (N849, N848, N143, N717);
not NOT1 (N850, N835);
not NOT1 (N851, N849);
buf BUF1 (N852, N847);
or OR3 (N853, N851, N626, N2);
buf BUF1 (N854, N837);
xor XOR2 (N855, N854, N140);
and AND3 (N856, N824, N585, N112);
xor XOR2 (N857, N856, N637);
xor XOR2 (N858, N845, N317);
or OR4 (N859, N838, N164, N665, N410);
not NOT1 (N860, N814);
nand NAND3 (N861, N857, N106, N706);
xor XOR2 (N862, N859, N31);
not NOT1 (N863, N853);
nor NOR4 (N864, N858, N581, N728, N81);
nor NOR3 (N865, N852, N17, N824);
xor XOR2 (N866, N846, N763);
xor XOR2 (N867, N865, N410);
nor NOR2 (N868, N834, N707);
buf BUF1 (N869, N867);
and AND4 (N870, N861, N117, N26, N32);
nand NAND3 (N871, N860, N390, N443);
nand NAND4 (N872, N862, N189, N768, N395);
buf BUF1 (N873, N868);
xor XOR2 (N874, N870, N473);
xor XOR2 (N875, N850, N714);
nand NAND2 (N876, N855, N316);
xor XOR2 (N877, N863, N239);
nor NOR2 (N878, N869, N712);
buf BUF1 (N879, N871);
not NOT1 (N880, N874);
nor NOR2 (N881, N877, N81);
not NOT1 (N882, N864);
or OR4 (N883, N881, N309, N590, N571);
and AND4 (N884, N882, N167, N833, N372);
nor NOR4 (N885, N872, N861, N113, N825);
not NOT1 (N886, N885);
or OR4 (N887, N886, N662, N93, N747);
not NOT1 (N888, N883);
or OR2 (N889, N884, N549);
buf BUF1 (N890, N879);
nand NAND2 (N891, N878, N836);
or OR2 (N892, N876, N19);
xor XOR2 (N893, N880, N826);
or OR3 (N894, N891, N52, N685);
nor NOR2 (N895, N888, N363);
nor NOR4 (N896, N892, N348, N369, N32);
nand NAND4 (N897, N890, N5, N705, N322);
or OR4 (N898, N893, N226, N496, N603);
or OR2 (N899, N873, N570);
nand NAND2 (N900, N898, N755);
not NOT1 (N901, N896);
xor XOR2 (N902, N875, N755);
not NOT1 (N903, N895);
xor XOR2 (N904, N887, N169);
or OR3 (N905, N900, N365, N273);
not NOT1 (N906, N903);
xor XOR2 (N907, N894, N42);
buf BUF1 (N908, N905);
xor XOR2 (N909, N897, N170);
not NOT1 (N910, N904);
and AND3 (N911, N908, N465, N885);
nand NAND2 (N912, N889, N500);
nor NOR4 (N913, N902, N840, N511, N238);
or OR4 (N914, N911, N859, N223, N286);
and AND3 (N915, N913, N63, N417);
buf BUF1 (N916, N901);
nand NAND3 (N917, N916, N302, N549);
nor NOR4 (N918, N914, N339, N765, N99);
xor XOR2 (N919, N912, N907);
nor NOR3 (N920, N743, N397, N237);
not NOT1 (N921, N866);
and AND2 (N922, N899, N669);
buf BUF1 (N923, N910);
xor XOR2 (N924, N920, N574);
nor NOR2 (N925, N921, N627);
nor NOR4 (N926, N906, N855, N738, N31);
xor XOR2 (N927, N922, N429);
nand NAND2 (N928, N924, N303);
not NOT1 (N929, N919);
nor NOR4 (N930, N923, N690, N21, N92);
and AND3 (N931, N909, N806, N177);
buf BUF1 (N932, N930);
not NOT1 (N933, N925);
xor XOR2 (N934, N931, N166);
xor XOR2 (N935, N915, N654);
buf BUF1 (N936, N934);
nor NOR4 (N937, N918, N718, N758, N681);
or OR2 (N938, N928, N937);
nor NOR4 (N939, N873, N664, N16, N454);
buf BUF1 (N940, N933);
and AND4 (N941, N935, N793, N309, N122);
not NOT1 (N942, N917);
or OR2 (N943, N939, N233);
buf BUF1 (N944, N926);
nand NAND4 (N945, N932, N748, N912, N205);
xor XOR2 (N946, N944, N152);
or OR2 (N947, N927, N657);
or OR4 (N948, N943, N100, N365, N536);
nand NAND2 (N949, N948, N250);
not NOT1 (N950, N947);
not NOT1 (N951, N941);
and AND4 (N952, N940, N795, N617, N1);
not NOT1 (N953, N929);
nand NAND4 (N954, N945, N800, N361, N859);
not NOT1 (N955, N952);
not NOT1 (N956, N954);
nand NAND4 (N957, N938, N897, N123, N154);
or OR2 (N958, N942, N172);
nor NOR4 (N959, N956, N561, N463, N313);
nand NAND4 (N960, N949, N245, N551, N538);
not NOT1 (N961, N951);
nand NAND2 (N962, N958, N335);
nand NAND3 (N963, N946, N152, N552);
xor XOR2 (N964, N960, N288);
nor NOR3 (N965, N955, N108, N675);
nor NOR4 (N966, N965, N583, N577, N148);
xor XOR2 (N967, N959, N671);
and AND3 (N968, N953, N792, N208);
buf BUF1 (N969, N964);
not NOT1 (N970, N963);
nand NAND2 (N971, N961, N681);
buf BUF1 (N972, N962);
nor NOR3 (N973, N970, N645, N887);
nor NOR2 (N974, N957, N540);
xor XOR2 (N975, N973, N17);
and AND2 (N976, N969, N609);
xor XOR2 (N977, N968, N4);
nor NOR4 (N978, N971, N629, N909, N436);
nor NOR3 (N979, N967, N328, N635);
or OR4 (N980, N966, N913, N941, N72);
not NOT1 (N981, N980);
and AND3 (N982, N975, N237, N407);
nand NAND2 (N983, N978, N569);
not NOT1 (N984, N982);
or OR4 (N985, N977, N967, N923, N964);
xor XOR2 (N986, N983, N317);
not NOT1 (N987, N981);
xor XOR2 (N988, N974, N19);
nand NAND3 (N989, N987, N680, N740);
nor NOR4 (N990, N985, N117, N875, N714);
buf BUF1 (N991, N990);
nand NAND2 (N992, N972, N896);
nand NAND4 (N993, N991, N52, N82, N865);
nor NOR4 (N994, N993, N188, N58, N301);
nand NAND4 (N995, N988, N677, N946, N814);
xor XOR2 (N996, N992, N429);
nor NOR2 (N997, N936, N982);
nand NAND3 (N998, N989, N87, N80);
and AND2 (N999, N950, N167);
or OR3 (N1000, N986, N82, N265);
not NOT1 (N1001, N998);
and AND4 (N1002, N994, N72, N759, N362);
nor NOR3 (N1003, N1001, N550, N671);
and AND2 (N1004, N984, N759);
and AND2 (N1005, N999, N155);
buf BUF1 (N1006, N1002);
buf BUF1 (N1007, N1004);
not NOT1 (N1008, N976);
buf BUF1 (N1009, N1007);
nor NOR2 (N1010, N997, N688);
xor XOR2 (N1011, N996, N123);
xor XOR2 (N1012, N995, N646);
nand NAND4 (N1013, N1006, N617, N898, N621);
or OR2 (N1014, N1003, N137);
buf BUF1 (N1015, N1011);
not NOT1 (N1016, N1008);
xor XOR2 (N1017, N1009, N426);
nor NOR2 (N1018, N1014, N626);
and AND4 (N1019, N979, N33, N926, N649);
nor NOR2 (N1020, N1012, N491);
and AND2 (N1021, N1010, N483);
nor NOR3 (N1022, N1019, N441, N560);
nand NAND2 (N1023, N1000, N743);
not NOT1 (N1024, N1020);
nand NAND2 (N1025, N1015, N176);
nor NOR4 (N1026, N1005, N578, N505, N930);
and AND3 (N1027, N1016, N334, N403);
xor XOR2 (N1028, N1023, N302);
or OR3 (N1029, N1018, N462, N312);
not NOT1 (N1030, N1028);
and AND2 (N1031, N1013, N594);
nand NAND4 (N1032, N1024, N340, N884, N593);
or OR4 (N1033, N1031, N922, N182, N996);
not NOT1 (N1034, N1026);
xor XOR2 (N1035, N1029, N986);
buf BUF1 (N1036, N1021);
not NOT1 (N1037, N1022);
nand NAND4 (N1038, N1027, N626, N195, N243);
not NOT1 (N1039, N1035);
not NOT1 (N1040, N1025);
buf BUF1 (N1041, N1017);
not NOT1 (N1042, N1038);
or OR3 (N1043, N1032, N568, N624);
nand NAND4 (N1044, N1041, N599, N30, N270);
and AND2 (N1045, N1039, N149);
xor XOR2 (N1046, N1036, N764);
or OR4 (N1047, N1033, N491, N16, N625);
nand NAND4 (N1048, N1044, N39, N565, N873);
buf BUF1 (N1049, N1048);
and AND4 (N1050, N1047, N549, N659, N352);
nand NAND4 (N1051, N1043, N960, N195, N647);
not NOT1 (N1052, N1046);
buf BUF1 (N1053, N1040);
or OR3 (N1054, N1034, N352, N949);
nand NAND3 (N1055, N1042, N939, N1042);
nand NAND4 (N1056, N1030, N967, N930, N261);
buf BUF1 (N1057, N1055);
not NOT1 (N1058, N1045);
xor XOR2 (N1059, N1037, N751);
buf BUF1 (N1060, N1054);
buf BUF1 (N1061, N1049);
buf BUF1 (N1062, N1058);
buf BUF1 (N1063, N1057);
buf BUF1 (N1064, N1051);
nand NAND2 (N1065, N1064, N345);
buf BUF1 (N1066, N1060);
nand NAND4 (N1067, N1050, N330, N1062, N246);
buf BUF1 (N1068, N592);
xor XOR2 (N1069, N1063, N297);
buf BUF1 (N1070, N1053);
and AND4 (N1071, N1061, N351, N778, N356);
not NOT1 (N1072, N1065);
xor XOR2 (N1073, N1070, N515);
nor NOR3 (N1074, N1067, N525, N395);
nor NOR3 (N1075, N1074, N535, N809);
and AND4 (N1076, N1066, N298, N444, N1014);
nand NAND3 (N1077, N1073, N1028, N968);
nor NOR2 (N1078, N1075, N800);
not NOT1 (N1079, N1078);
buf BUF1 (N1080, N1072);
not NOT1 (N1081, N1077);
and AND3 (N1082, N1076, N789, N977);
or OR4 (N1083, N1052, N794, N402, N640);
and AND2 (N1084, N1069, N925);
or OR3 (N1085, N1071, N524, N184);
not NOT1 (N1086, N1081);
nand NAND3 (N1087, N1068, N431, N989);
or OR3 (N1088, N1082, N698, N820);
nor NOR2 (N1089, N1087, N430);
or OR2 (N1090, N1085, N1078);
nor NOR4 (N1091, N1079, N332, N1074, N581);
nor NOR4 (N1092, N1084, N60, N1032, N798);
nand NAND3 (N1093, N1088, N25, N947);
buf BUF1 (N1094, N1092);
or OR4 (N1095, N1091, N582, N468, N150);
and AND2 (N1096, N1094, N778);
buf BUF1 (N1097, N1089);
not NOT1 (N1098, N1095);
buf BUF1 (N1099, N1059);
not NOT1 (N1100, N1080);
or OR2 (N1101, N1098, N212);
and AND4 (N1102, N1093, N538, N777, N517);
nand NAND2 (N1103, N1090, N117);
xor XOR2 (N1104, N1099, N305);
or OR4 (N1105, N1086, N507, N2, N490);
not NOT1 (N1106, N1097);
or OR3 (N1107, N1096, N812, N827);
nor NOR3 (N1108, N1100, N426, N654);
or OR4 (N1109, N1107, N1019, N771, N599);
and AND4 (N1110, N1109, N889, N885, N833);
or OR2 (N1111, N1103, N1058);
not NOT1 (N1112, N1111);
xor XOR2 (N1113, N1102, N955);
not NOT1 (N1114, N1104);
or OR2 (N1115, N1105, N127);
xor XOR2 (N1116, N1106, N994);
nor NOR3 (N1117, N1056, N402, N434);
nor NOR2 (N1118, N1115, N14);
and AND4 (N1119, N1116, N641, N714, N246);
not NOT1 (N1120, N1117);
nor NOR3 (N1121, N1118, N1087, N655);
nor NOR2 (N1122, N1113, N1059);
xor XOR2 (N1123, N1119, N378);
buf BUF1 (N1124, N1110);
nand NAND3 (N1125, N1120, N252, N339);
not NOT1 (N1126, N1122);
and AND3 (N1127, N1124, N1086, N463);
xor XOR2 (N1128, N1083, N1059);
and AND3 (N1129, N1121, N62, N400);
and AND2 (N1130, N1125, N679);
and AND2 (N1131, N1108, N181);
or OR3 (N1132, N1131, N890, N868);
and AND3 (N1133, N1128, N867, N388);
nand NAND4 (N1134, N1130, N265, N252, N420);
xor XOR2 (N1135, N1127, N219);
nor NOR2 (N1136, N1126, N282);
or OR3 (N1137, N1129, N497, N584);
buf BUF1 (N1138, N1133);
or OR2 (N1139, N1114, N1028);
nor NOR2 (N1140, N1134, N635);
xor XOR2 (N1141, N1135, N1112);
nor NOR3 (N1142, N115, N220, N143);
nand NAND3 (N1143, N1137, N228, N611);
xor XOR2 (N1144, N1138, N363);
nor NOR4 (N1145, N1144, N364, N325, N995);
nand NAND2 (N1146, N1136, N868);
nand NAND2 (N1147, N1142, N659);
not NOT1 (N1148, N1147);
and AND4 (N1149, N1145, N92, N466, N954);
xor XOR2 (N1150, N1132, N720);
nor NOR2 (N1151, N1141, N1138);
nand NAND3 (N1152, N1148, N15, N45);
nor NOR3 (N1153, N1101, N822, N477);
nand NAND2 (N1154, N1143, N218);
not NOT1 (N1155, N1146);
not NOT1 (N1156, N1150);
nor NOR2 (N1157, N1140, N307);
nor NOR3 (N1158, N1153, N27, N292);
not NOT1 (N1159, N1123);
or OR2 (N1160, N1157, N284);
not NOT1 (N1161, N1156);
nor NOR4 (N1162, N1159, N91, N890, N144);
xor XOR2 (N1163, N1161, N413);
not NOT1 (N1164, N1151);
buf BUF1 (N1165, N1164);
nor NOR3 (N1166, N1165, N792, N236);
xor XOR2 (N1167, N1155, N149);
nand NAND2 (N1168, N1167, N496);
nand NAND3 (N1169, N1154, N224, N1102);
not NOT1 (N1170, N1160);
buf BUF1 (N1171, N1166);
buf BUF1 (N1172, N1149);
and AND2 (N1173, N1152, N705);
not NOT1 (N1174, N1158);
nor NOR4 (N1175, N1172, N775, N956, N1114);
and AND4 (N1176, N1174, N999, N395, N491);
and AND3 (N1177, N1170, N342, N863);
nand NAND3 (N1178, N1177, N151, N858);
buf BUF1 (N1179, N1176);
xor XOR2 (N1180, N1171, N235);
not NOT1 (N1181, N1173);
and AND4 (N1182, N1180, N159, N236, N214);
nand NAND3 (N1183, N1169, N1098, N641);
or OR4 (N1184, N1168, N231, N443, N401);
and AND4 (N1185, N1182, N1080, N992, N71);
buf BUF1 (N1186, N1184);
not NOT1 (N1187, N1175);
buf BUF1 (N1188, N1183);
and AND3 (N1189, N1162, N682, N407);
buf BUF1 (N1190, N1179);
buf BUF1 (N1191, N1178);
or OR4 (N1192, N1185, N873, N444, N946);
buf BUF1 (N1193, N1139);
nand NAND3 (N1194, N1163, N46, N622);
buf BUF1 (N1195, N1192);
nor NOR3 (N1196, N1189, N705, N542);
xor XOR2 (N1197, N1187, N655);
not NOT1 (N1198, N1190);
nor NOR2 (N1199, N1197, N962);
xor XOR2 (N1200, N1193, N1078);
and AND3 (N1201, N1198, N762, N420);
and AND3 (N1202, N1181, N1141, N685);
not NOT1 (N1203, N1186);
and AND2 (N1204, N1202, N1094);
and AND3 (N1205, N1188, N1053, N609);
buf BUF1 (N1206, N1196);
nand NAND2 (N1207, N1200, N1139);
xor XOR2 (N1208, N1191, N457);
xor XOR2 (N1209, N1203, N537);
xor XOR2 (N1210, N1208, N424);
and AND4 (N1211, N1195, N563, N853, N969);
and AND4 (N1212, N1204, N694, N758, N804);
xor XOR2 (N1213, N1207, N677);
not NOT1 (N1214, N1206);
or OR3 (N1215, N1194, N239, N1067);
xor XOR2 (N1216, N1213, N422);
nor NOR2 (N1217, N1199, N156);
nor NOR2 (N1218, N1214, N672);
xor XOR2 (N1219, N1201, N946);
buf BUF1 (N1220, N1210);
nand NAND3 (N1221, N1215, N200, N987);
xor XOR2 (N1222, N1219, N796);
not NOT1 (N1223, N1216);
xor XOR2 (N1224, N1223, N442);
nand NAND2 (N1225, N1211, N135);
not NOT1 (N1226, N1220);
not NOT1 (N1227, N1218);
xor XOR2 (N1228, N1226, N1184);
not NOT1 (N1229, N1222);
nand NAND4 (N1230, N1228, N1024, N1129, N1128);
nand NAND3 (N1231, N1205, N465, N700);
not NOT1 (N1232, N1230);
not NOT1 (N1233, N1221);
or OR2 (N1234, N1217, N945);
or OR3 (N1235, N1232, N1067, N931);
nor NOR2 (N1236, N1233, N583);
xor XOR2 (N1237, N1235, N1200);
xor XOR2 (N1238, N1229, N573);
nor NOR4 (N1239, N1237, N202, N990, N399);
nand NAND2 (N1240, N1231, N986);
nand NAND4 (N1241, N1239, N785, N584, N755);
nand NAND3 (N1242, N1225, N146, N968);
nor NOR4 (N1243, N1242, N1054, N1035, N311);
or OR3 (N1244, N1234, N1073, N163);
nor NOR2 (N1245, N1212, N532);
or OR4 (N1246, N1224, N1152, N746, N530);
not NOT1 (N1247, N1244);
xor XOR2 (N1248, N1240, N495);
nor NOR4 (N1249, N1243, N962, N324, N968);
and AND2 (N1250, N1248, N874);
not NOT1 (N1251, N1245);
nor NOR4 (N1252, N1246, N216, N56, N789);
nor NOR2 (N1253, N1251, N398);
buf BUF1 (N1254, N1238);
and AND3 (N1255, N1227, N415, N669);
not NOT1 (N1256, N1236);
or OR4 (N1257, N1250, N706, N1027, N1015);
xor XOR2 (N1258, N1256, N215);
nand NAND2 (N1259, N1249, N99);
xor XOR2 (N1260, N1258, N426);
or OR4 (N1261, N1255, N1088, N790, N354);
not NOT1 (N1262, N1241);
or OR2 (N1263, N1254, N10);
not NOT1 (N1264, N1259);
nor NOR3 (N1265, N1260, N642, N7);
buf BUF1 (N1266, N1264);
not NOT1 (N1267, N1209);
and AND2 (N1268, N1253, N1060);
and AND4 (N1269, N1252, N1116, N651, N747);
or OR3 (N1270, N1263, N1130, N393);
or OR2 (N1271, N1265, N1214);
nor NOR2 (N1272, N1269, N697);
nor NOR4 (N1273, N1271, N291, N786, N455);
not NOT1 (N1274, N1257);
xor XOR2 (N1275, N1267, N370);
nor NOR3 (N1276, N1261, N531, N199);
and AND3 (N1277, N1273, N931, N462);
nand NAND3 (N1278, N1247, N760, N421);
or OR3 (N1279, N1274, N142, N311);
buf BUF1 (N1280, N1279);
nand NAND4 (N1281, N1278, N279, N345, N401);
or OR4 (N1282, N1275, N1118, N589, N363);
nand NAND3 (N1283, N1270, N1044, N544);
xor XOR2 (N1284, N1272, N71);
or OR4 (N1285, N1268, N933, N562, N974);
nand NAND2 (N1286, N1262, N479);
buf BUF1 (N1287, N1286);
buf BUF1 (N1288, N1284);
xor XOR2 (N1289, N1276, N749);
nor NOR3 (N1290, N1281, N492, N702);
buf BUF1 (N1291, N1290);
and AND3 (N1292, N1287, N744, N1024);
and AND4 (N1293, N1266, N360, N157, N728);
nor NOR4 (N1294, N1288, N220, N933, N60);
not NOT1 (N1295, N1291);
and AND3 (N1296, N1282, N982, N494);
nand NAND2 (N1297, N1285, N603);
buf BUF1 (N1298, N1292);
buf BUF1 (N1299, N1293);
nand NAND4 (N1300, N1280, N697, N1004, N451);
not NOT1 (N1301, N1295);
or OR3 (N1302, N1298, N590, N326);
nor NOR4 (N1303, N1302, N1144, N1038, N580);
and AND4 (N1304, N1301, N92, N511, N613);
or OR3 (N1305, N1304, N911, N1283);
and AND2 (N1306, N238, N926);
and AND2 (N1307, N1297, N24);
and AND3 (N1308, N1277, N636, N233);
nand NAND4 (N1309, N1308, N226, N599, N234);
buf BUF1 (N1310, N1309);
xor XOR2 (N1311, N1300, N1101);
buf BUF1 (N1312, N1306);
xor XOR2 (N1313, N1311, N539);
xor XOR2 (N1314, N1307, N959);
not NOT1 (N1315, N1305);
buf BUF1 (N1316, N1303);
nor NOR4 (N1317, N1313, N244, N1220, N1195);
or OR4 (N1318, N1310, N876, N605, N356);
or OR4 (N1319, N1315, N536, N170, N778);
nor NOR4 (N1320, N1296, N267, N702, N683);
or OR2 (N1321, N1319, N935);
xor XOR2 (N1322, N1294, N225);
xor XOR2 (N1323, N1321, N178);
nor NOR2 (N1324, N1314, N520);
nor NOR2 (N1325, N1323, N1017);
nor NOR3 (N1326, N1312, N913, N5);
xor XOR2 (N1327, N1324, N544);
nand NAND2 (N1328, N1320, N880);
nor NOR2 (N1329, N1299, N150);
not NOT1 (N1330, N1322);
xor XOR2 (N1331, N1328, N242);
nand NAND4 (N1332, N1327, N118, N360, N514);
and AND4 (N1333, N1330, N1317, N520, N974);
buf BUF1 (N1334, N1081);
or OR3 (N1335, N1332, N556, N795);
not NOT1 (N1336, N1316);
and AND4 (N1337, N1325, N1199, N377, N745);
not NOT1 (N1338, N1318);
nor NOR4 (N1339, N1326, N624, N109, N293);
or OR4 (N1340, N1289, N247, N630, N1011);
xor XOR2 (N1341, N1331, N1200);
nor NOR2 (N1342, N1334, N40);
not NOT1 (N1343, N1337);
xor XOR2 (N1344, N1329, N1217);
not NOT1 (N1345, N1344);
not NOT1 (N1346, N1339);
xor XOR2 (N1347, N1342, N1159);
xor XOR2 (N1348, N1338, N866);
xor XOR2 (N1349, N1346, N1259);
xor XOR2 (N1350, N1348, N336);
not NOT1 (N1351, N1343);
nand NAND2 (N1352, N1351, N341);
not NOT1 (N1353, N1340);
and AND3 (N1354, N1349, N1078, N1101);
xor XOR2 (N1355, N1335, N1339);
buf BUF1 (N1356, N1347);
nor NOR4 (N1357, N1352, N915, N538, N255);
buf BUF1 (N1358, N1341);
or OR3 (N1359, N1345, N725, N21);
nand NAND3 (N1360, N1357, N782, N1151);
xor XOR2 (N1361, N1359, N174);
not NOT1 (N1362, N1361);
and AND4 (N1363, N1358, N51, N1269, N1260);
or OR4 (N1364, N1350, N846, N394, N278);
xor XOR2 (N1365, N1356, N115);
buf BUF1 (N1366, N1363);
or OR4 (N1367, N1355, N987, N274, N861);
nand NAND4 (N1368, N1354, N109, N681, N770);
not NOT1 (N1369, N1353);
or OR3 (N1370, N1366, N751, N1306);
and AND2 (N1371, N1360, N966);
not NOT1 (N1372, N1368);
buf BUF1 (N1373, N1369);
xor XOR2 (N1374, N1333, N993);
buf BUF1 (N1375, N1374);
not NOT1 (N1376, N1365);
nand NAND3 (N1377, N1336, N900, N636);
buf BUF1 (N1378, N1362);
buf BUF1 (N1379, N1376);
xor XOR2 (N1380, N1379, N521);
buf BUF1 (N1381, N1377);
or OR3 (N1382, N1367, N615, N762);
and AND4 (N1383, N1373, N96, N617, N1257);
not NOT1 (N1384, N1381);
and AND2 (N1385, N1372, N808);
nor NOR4 (N1386, N1383, N841, N1004, N919);
nand NAND4 (N1387, N1364, N541, N1044, N1091);
not NOT1 (N1388, N1387);
not NOT1 (N1389, N1384);
xor XOR2 (N1390, N1380, N1247);
or OR2 (N1391, N1370, N353);
nand NAND3 (N1392, N1386, N1131, N430);
nand NAND4 (N1393, N1371, N659, N39, N309);
or OR3 (N1394, N1388, N296, N1199);
buf BUF1 (N1395, N1393);
nor NOR3 (N1396, N1392, N1094, N481);
xor XOR2 (N1397, N1394, N569);
nor NOR4 (N1398, N1378, N1317, N673, N328);
buf BUF1 (N1399, N1398);
or OR4 (N1400, N1390, N1314, N65, N686);
nor NOR3 (N1401, N1400, N955, N1000);
nor NOR3 (N1402, N1385, N1056, N757);
nand NAND2 (N1403, N1391, N192);
not NOT1 (N1404, N1401);
xor XOR2 (N1405, N1403, N765);
and AND2 (N1406, N1404, N1247);
xor XOR2 (N1407, N1395, N433);
not NOT1 (N1408, N1375);
or OR3 (N1409, N1406, N55, N1205);
and AND2 (N1410, N1399, N408);
not NOT1 (N1411, N1402);
nand NAND4 (N1412, N1389, N239, N787, N1251);
nor NOR3 (N1413, N1408, N1100, N768);
and AND4 (N1414, N1412, N1292, N1218, N918);
not NOT1 (N1415, N1414);
buf BUF1 (N1416, N1413);
not NOT1 (N1417, N1397);
nand NAND3 (N1418, N1410, N1172, N755);
nand NAND4 (N1419, N1407, N746, N515, N317);
nor NOR4 (N1420, N1419, N1156, N1069, N190);
or OR3 (N1421, N1416, N1278, N1150);
xor XOR2 (N1422, N1418, N655);
nand NAND4 (N1423, N1396, N326, N1263, N5);
nor NOR4 (N1424, N1409, N1186, N699, N626);
or OR4 (N1425, N1423, N346, N126, N507);
nand NAND3 (N1426, N1411, N886, N723);
nand NAND4 (N1427, N1415, N889, N60, N371);
nor NOR2 (N1428, N1427, N549);
nand NAND4 (N1429, N1421, N102, N899, N1035);
nand NAND2 (N1430, N1405, N715);
buf BUF1 (N1431, N1425);
not NOT1 (N1432, N1420);
nor NOR3 (N1433, N1430, N352, N1066);
or OR2 (N1434, N1382, N1067);
and AND3 (N1435, N1434, N115, N42);
nor NOR2 (N1436, N1424, N955);
nand NAND2 (N1437, N1432, N754);
or OR4 (N1438, N1422, N542, N92, N1010);
buf BUF1 (N1439, N1438);
or OR3 (N1440, N1428, N1209, N227);
not NOT1 (N1441, N1431);
or OR3 (N1442, N1429, N1056, N308);
and AND2 (N1443, N1435, N777);
nand NAND3 (N1444, N1443, N360, N1040);
and AND4 (N1445, N1433, N37, N182, N1393);
xor XOR2 (N1446, N1426, N1246);
xor XOR2 (N1447, N1436, N338);
and AND2 (N1448, N1439, N1417);
not NOT1 (N1449, N715);
buf BUF1 (N1450, N1446);
nor NOR4 (N1451, N1450, N842, N1019, N832);
xor XOR2 (N1452, N1444, N78);
xor XOR2 (N1453, N1449, N318);
and AND4 (N1454, N1437, N1335, N1240, N567);
or OR3 (N1455, N1445, N1192, N361);
nor NOR2 (N1456, N1441, N1140);
nor NOR2 (N1457, N1452, N502);
and AND2 (N1458, N1456, N637);
nand NAND2 (N1459, N1454, N1427);
buf BUF1 (N1460, N1447);
buf BUF1 (N1461, N1457);
not NOT1 (N1462, N1442);
nand NAND4 (N1463, N1460, N1192, N1338, N1337);
xor XOR2 (N1464, N1461, N1373);
or OR4 (N1465, N1448, N591, N7, N1387);
buf BUF1 (N1466, N1464);
or OR2 (N1467, N1463, N1068);
not NOT1 (N1468, N1455);
buf BUF1 (N1469, N1465);
xor XOR2 (N1470, N1469, N867);
nand NAND2 (N1471, N1451, N1072);
buf BUF1 (N1472, N1466);
or OR2 (N1473, N1440, N250);
nand NAND4 (N1474, N1458, N434, N785, N794);
not NOT1 (N1475, N1472);
or OR4 (N1476, N1475, N1373, N311, N785);
nor NOR4 (N1477, N1468, N1437, N1433, N664);
buf BUF1 (N1478, N1476);
xor XOR2 (N1479, N1473, N1395);
and AND2 (N1480, N1467, N1104);
and AND3 (N1481, N1470, N1447, N1038);
xor XOR2 (N1482, N1480, N1117);
buf BUF1 (N1483, N1477);
not NOT1 (N1484, N1459);
and AND3 (N1485, N1484, N1445, N1038);
nand NAND2 (N1486, N1453, N593);
nand NAND2 (N1487, N1486, N751);
nand NAND3 (N1488, N1479, N1033, N653);
or OR2 (N1489, N1483, N938);
buf BUF1 (N1490, N1462);
or OR3 (N1491, N1488, N1076, N627);
nand NAND2 (N1492, N1485, N932);
nor NOR3 (N1493, N1478, N596, N556);
nand NAND3 (N1494, N1482, N125, N892);
nand NAND3 (N1495, N1489, N590, N757);
nand NAND3 (N1496, N1492, N128, N892);
nor NOR3 (N1497, N1481, N1471, N414);
nor NOR4 (N1498, N641, N807, N1112, N890);
or OR2 (N1499, N1490, N67);
nor NOR2 (N1500, N1474, N1323);
or OR2 (N1501, N1499, N1280);
buf BUF1 (N1502, N1491);
xor XOR2 (N1503, N1497, N1334);
xor XOR2 (N1504, N1501, N1087);
xor XOR2 (N1505, N1495, N709);
buf BUF1 (N1506, N1502);
xor XOR2 (N1507, N1500, N129);
and AND3 (N1508, N1506, N754, N766);
not NOT1 (N1509, N1494);
nor NOR4 (N1510, N1487, N770, N745, N87);
nand NAND4 (N1511, N1508, N862, N199, N1449);
buf BUF1 (N1512, N1498);
or OR3 (N1513, N1493, N717, N164);
nor NOR4 (N1514, N1505, N1091, N617, N135);
or OR2 (N1515, N1504, N1294);
xor XOR2 (N1516, N1514, N956);
and AND3 (N1517, N1512, N333, N234);
buf BUF1 (N1518, N1496);
not NOT1 (N1519, N1518);
or OR3 (N1520, N1515, N1042, N299);
nor NOR3 (N1521, N1516, N772, N1502);
or OR3 (N1522, N1511, N1316, N1216);
and AND3 (N1523, N1513, N90, N1218);
and AND3 (N1524, N1517, N754, N429);
xor XOR2 (N1525, N1520, N175);
nor NOR4 (N1526, N1503, N428, N1253, N361);
xor XOR2 (N1527, N1523, N39);
not NOT1 (N1528, N1521);
xor XOR2 (N1529, N1507, N1152);
and AND3 (N1530, N1525, N1520, N173);
nand NAND4 (N1531, N1530, N248, N633, N1470);
not NOT1 (N1532, N1528);
and AND4 (N1533, N1524, N1157, N686, N1497);
or OR2 (N1534, N1531, N1433);
xor XOR2 (N1535, N1527, N589);
nor NOR2 (N1536, N1510, N815);
xor XOR2 (N1537, N1535, N205);
buf BUF1 (N1538, N1537);
xor XOR2 (N1539, N1509, N999);
buf BUF1 (N1540, N1534);
xor XOR2 (N1541, N1522, N1538);
buf BUF1 (N1542, N1308);
nor NOR2 (N1543, N1533, N1320);
not NOT1 (N1544, N1540);
nor NOR4 (N1545, N1532, N1409, N855, N647);
nor NOR3 (N1546, N1519, N987, N582);
xor XOR2 (N1547, N1539, N1012);
nand NAND3 (N1548, N1543, N48, N521);
nand NAND4 (N1549, N1546, N854, N1173, N665);
buf BUF1 (N1550, N1526);
and AND2 (N1551, N1542, N1392);
not NOT1 (N1552, N1545);
nor NOR2 (N1553, N1544, N75);
buf BUF1 (N1554, N1529);
nor NOR2 (N1555, N1536, N1217);
or OR2 (N1556, N1551, N1339);
and AND2 (N1557, N1550, N1517);
buf BUF1 (N1558, N1547);
nand NAND3 (N1559, N1558, N56, N1404);
xor XOR2 (N1560, N1541, N1307);
xor XOR2 (N1561, N1549, N1497);
not NOT1 (N1562, N1552);
nor NOR4 (N1563, N1561, N222, N1309, N1206);
not NOT1 (N1564, N1553);
buf BUF1 (N1565, N1555);
or OR3 (N1566, N1565, N528, N978);
nor NOR4 (N1567, N1548, N175, N296, N1400);
not NOT1 (N1568, N1554);
nor NOR2 (N1569, N1563, N656);
or OR4 (N1570, N1567, N934, N109, N899);
nor NOR4 (N1571, N1566, N221, N1380, N684);
xor XOR2 (N1572, N1569, N412);
nand NAND2 (N1573, N1556, N660);
nor NOR2 (N1574, N1568, N1231);
xor XOR2 (N1575, N1564, N1429);
not NOT1 (N1576, N1560);
nor NOR2 (N1577, N1571, N196);
not NOT1 (N1578, N1575);
buf BUF1 (N1579, N1557);
nand NAND3 (N1580, N1570, N202, N1329);
not NOT1 (N1581, N1577);
buf BUF1 (N1582, N1573);
buf BUF1 (N1583, N1581);
xor XOR2 (N1584, N1579, N369);
not NOT1 (N1585, N1578);
or OR3 (N1586, N1580, N461, N1445);
nor NOR2 (N1587, N1585, N676);
buf BUF1 (N1588, N1584);
or OR4 (N1589, N1559, N1003, N387, N229);
buf BUF1 (N1590, N1574);
and AND3 (N1591, N1562, N783, N909);
nand NAND2 (N1592, N1589, N1192);
xor XOR2 (N1593, N1591, N444);
not NOT1 (N1594, N1587);
or OR4 (N1595, N1592, N611, N507, N1170);
xor XOR2 (N1596, N1572, N263);
or OR3 (N1597, N1583, N606, N389);
buf BUF1 (N1598, N1597);
buf BUF1 (N1599, N1596);
xor XOR2 (N1600, N1588, N1273);
nor NOR2 (N1601, N1590, N436);
not NOT1 (N1602, N1576);
not NOT1 (N1603, N1595);
and AND3 (N1604, N1599, N395, N483);
nor NOR4 (N1605, N1593, N1377, N1315, N1067);
buf BUF1 (N1606, N1582);
and AND2 (N1607, N1602, N833);
xor XOR2 (N1608, N1605, N1184);
nand NAND3 (N1609, N1594, N1540, N897);
not NOT1 (N1610, N1604);
and AND4 (N1611, N1603, N1330, N1320, N516);
nand NAND2 (N1612, N1607, N478);
nand NAND3 (N1613, N1612, N571, N1272);
or OR4 (N1614, N1600, N121, N1108, N128);
and AND2 (N1615, N1601, N127);
buf BUF1 (N1616, N1586);
or OR4 (N1617, N1608, N879, N451, N507);
not NOT1 (N1618, N1606);
or OR3 (N1619, N1613, N207, N1100);
buf BUF1 (N1620, N1598);
buf BUF1 (N1621, N1620);
and AND4 (N1622, N1615, N291, N799, N834);
nor NOR3 (N1623, N1621, N225, N1067);
nand NAND4 (N1624, N1623, N1191, N155, N747);
xor XOR2 (N1625, N1614, N1286);
and AND4 (N1626, N1624, N50, N409, N860);
and AND4 (N1627, N1622, N203, N1163, N6);
and AND3 (N1628, N1617, N1245, N177);
buf BUF1 (N1629, N1618);
nand NAND4 (N1630, N1625, N351, N408, N1384);
buf BUF1 (N1631, N1616);
nor NOR3 (N1632, N1626, N1357, N696);
buf BUF1 (N1633, N1619);
xor XOR2 (N1634, N1611, N1402);
nand NAND2 (N1635, N1627, N468);
and AND4 (N1636, N1632, N137, N899, N1230);
xor XOR2 (N1637, N1609, N890);
nand NAND2 (N1638, N1610, N632);
nor NOR4 (N1639, N1637, N1074, N1158, N894);
and AND3 (N1640, N1629, N833, N885);
xor XOR2 (N1641, N1630, N775);
nand NAND2 (N1642, N1639, N968);
or OR2 (N1643, N1642, N933);
nor NOR4 (N1644, N1636, N1274, N1269, N714);
buf BUF1 (N1645, N1631);
buf BUF1 (N1646, N1645);
nand NAND2 (N1647, N1633, N1281);
nand NAND2 (N1648, N1640, N62);
xor XOR2 (N1649, N1648, N730);
xor XOR2 (N1650, N1643, N1598);
nor NOR2 (N1651, N1628, N1132);
not NOT1 (N1652, N1650);
nand NAND4 (N1653, N1647, N371, N818, N410);
or OR4 (N1654, N1641, N108, N217, N312);
nand NAND3 (N1655, N1649, N417, N958);
buf BUF1 (N1656, N1634);
nor NOR4 (N1657, N1651, N973, N1646, N1296);
and AND4 (N1658, N1218, N22, N713, N297);
and AND3 (N1659, N1655, N274, N1460);
buf BUF1 (N1660, N1652);
not NOT1 (N1661, N1656);
buf BUF1 (N1662, N1635);
not NOT1 (N1663, N1654);
nor NOR4 (N1664, N1657, N838, N528, N565);
nand NAND4 (N1665, N1658, N880, N678, N567);
xor XOR2 (N1666, N1660, N1336);
buf BUF1 (N1667, N1663);
and AND2 (N1668, N1661, N145);
buf BUF1 (N1669, N1653);
not NOT1 (N1670, N1666);
nor NOR4 (N1671, N1667, N817, N107, N1405);
nor NOR4 (N1672, N1668, N1128, N1263, N925);
nand NAND4 (N1673, N1672, N557, N436, N203);
buf BUF1 (N1674, N1659);
xor XOR2 (N1675, N1638, N593);
nand NAND2 (N1676, N1644, N1332);
or OR2 (N1677, N1671, N1522);
nand NAND2 (N1678, N1677, N1434);
and AND2 (N1679, N1675, N545);
and AND2 (N1680, N1674, N823);
xor XOR2 (N1681, N1679, N1304);
nor NOR4 (N1682, N1680, N1552, N257, N1124);
xor XOR2 (N1683, N1681, N765);
buf BUF1 (N1684, N1664);
buf BUF1 (N1685, N1684);
nor NOR2 (N1686, N1676, N958);
and AND3 (N1687, N1670, N584, N963);
nor NOR3 (N1688, N1678, N477, N1165);
buf BUF1 (N1689, N1687);
nand NAND3 (N1690, N1689, N1331, N1424);
buf BUF1 (N1691, N1662);
buf BUF1 (N1692, N1673);
xor XOR2 (N1693, N1686, N1663);
nand NAND2 (N1694, N1665, N1001);
buf BUF1 (N1695, N1685);
and AND3 (N1696, N1682, N1462, N997);
not NOT1 (N1697, N1669);
xor XOR2 (N1698, N1694, N1531);
nand NAND2 (N1699, N1688, N936);
or OR4 (N1700, N1696, N1397, N885, N555);
nor NOR3 (N1701, N1699, N545, N1325);
not NOT1 (N1702, N1683);
or OR2 (N1703, N1692, N621);
and AND4 (N1704, N1700, N1086, N1181, N1349);
and AND3 (N1705, N1691, N1369, N1);
nand NAND3 (N1706, N1690, N719, N422);
nand NAND2 (N1707, N1701, N1669);
nor NOR4 (N1708, N1702, N1032, N1284, N1597);
and AND3 (N1709, N1708, N777, N1373);
buf BUF1 (N1710, N1697);
or OR2 (N1711, N1704, N1284);
and AND4 (N1712, N1703, N999, N1270, N237);
nand NAND4 (N1713, N1709, N622, N1570, N1198);
nor NOR2 (N1714, N1710, N238);
nor NOR3 (N1715, N1712, N1351, N1305);
nor NOR2 (N1716, N1715, N1130);
not NOT1 (N1717, N1714);
xor XOR2 (N1718, N1693, N1189);
nand NAND3 (N1719, N1718, N1203, N221);
xor XOR2 (N1720, N1698, N535);
nand NAND3 (N1721, N1706, N567, N268);
or OR4 (N1722, N1695, N815, N389, N483);
not NOT1 (N1723, N1713);
or OR4 (N1724, N1723, N1011, N1154, N1663);
not NOT1 (N1725, N1716);
and AND3 (N1726, N1705, N802, N1003);
xor XOR2 (N1727, N1724, N378);
nand NAND3 (N1728, N1726, N676, N1299);
nor NOR2 (N1729, N1711, N1385);
nand NAND3 (N1730, N1725, N1224, N258);
not NOT1 (N1731, N1717);
or OR3 (N1732, N1728, N246, N802);
nor NOR4 (N1733, N1732, N828, N910, N726);
or OR2 (N1734, N1720, N71);
nor NOR3 (N1735, N1731, N633, N393);
nor NOR2 (N1736, N1730, N1238);
or OR4 (N1737, N1727, N926, N14, N638);
nor NOR2 (N1738, N1722, N1285);
not NOT1 (N1739, N1738);
nand NAND2 (N1740, N1737, N254);
buf BUF1 (N1741, N1736);
buf BUF1 (N1742, N1707);
and AND2 (N1743, N1741, N66);
xor XOR2 (N1744, N1729, N361);
nand NAND3 (N1745, N1735, N796, N249);
not NOT1 (N1746, N1719);
and AND4 (N1747, N1733, N1339, N1014, N1326);
not NOT1 (N1748, N1746);
buf BUF1 (N1749, N1744);
xor XOR2 (N1750, N1748, N608);
and AND2 (N1751, N1734, N414);
xor XOR2 (N1752, N1721, N33);
nand NAND3 (N1753, N1747, N1069, N180);
nor NOR4 (N1754, N1745, N767, N589, N822);
xor XOR2 (N1755, N1750, N1677);
or OR2 (N1756, N1754, N1039);
or OR3 (N1757, N1752, N207, N1394);
or OR2 (N1758, N1740, N387);
buf BUF1 (N1759, N1757);
and AND3 (N1760, N1755, N1111, N956);
nor NOR2 (N1761, N1760, N1343);
buf BUF1 (N1762, N1749);
nor NOR3 (N1763, N1759, N1640, N48);
nor NOR4 (N1764, N1761, N423, N316, N925);
nor NOR2 (N1765, N1743, N1514);
xor XOR2 (N1766, N1762, N1054);
not NOT1 (N1767, N1758);
nand NAND3 (N1768, N1767, N651, N889);
xor XOR2 (N1769, N1763, N622);
not NOT1 (N1770, N1751);
or OR3 (N1771, N1742, N1769, N1020);
not NOT1 (N1772, N1372);
and AND2 (N1773, N1772, N672);
xor XOR2 (N1774, N1770, N1169);
or OR2 (N1775, N1771, N1061);
and AND3 (N1776, N1756, N1107, N1293);
and AND4 (N1777, N1768, N1263, N297, N563);
xor XOR2 (N1778, N1777, N1215);
not NOT1 (N1779, N1739);
or OR2 (N1780, N1764, N8);
not NOT1 (N1781, N1774);
not NOT1 (N1782, N1765);
nor NOR3 (N1783, N1782, N1466, N503);
and AND4 (N1784, N1766, N676, N552, N827);
and AND4 (N1785, N1775, N21, N1529, N1656);
xor XOR2 (N1786, N1781, N231);
not NOT1 (N1787, N1780);
or OR3 (N1788, N1784, N1782, N1015);
not NOT1 (N1789, N1787);
buf BUF1 (N1790, N1779);
buf BUF1 (N1791, N1753);
or OR2 (N1792, N1773, N1347);
or OR2 (N1793, N1790, N1779);
buf BUF1 (N1794, N1786);
buf BUF1 (N1795, N1788);
or OR2 (N1796, N1794, N1399);
not NOT1 (N1797, N1795);
nor NOR2 (N1798, N1778, N212);
not NOT1 (N1799, N1776);
xor XOR2 (N1800, N1798, N1320);
and AND3 (N1801, N1797, N767, N1795);
or OR4 (N1802, N1783, N294, N545, N863);
xor XOR2 (N1803, N1785, N642);
nor NOR2 (N1804, N1802, N1627);
not NOT1 (N1805, N1803);
xor XOR2 (N1806, N1792, N1797);
or OR3 (N1807, N1799, N172, N920);
or OR4 (N1808, N1804, N903, N993, N78);
buf BUF1 (N1809, N1806);
xor XOR2 (N1810, N1789, N1709);
xor XOR2 (N1811, N1805, N598);
or OR3 (N1812, N1807, N29, N679);
xor XOR2 (N1813, N1812, N791);
nor NOR3 (N1814, N1813, N952, N1543);
and AND3 (N1815, N1811, N836, N71);
nor NOR2 (N1816, N1800, N1218);
not NOT1 (N1817, N1814);
xor XOR2 (N1818, N1809, N1807);
xor XOR2 (N1819, N1801, N1422);
and AND3 (N1820, N1815, N1470, N581);
nand NAND2 (N1821, N1817, N335);
buf BUF1 (N1822, N1808);
not NOT1 (N1823, N1822);
or OR2 (N1824, N1791, N1711);
buf BUF1 (N1825, N1819);
xor XOR2 (N1826, N1816, N495);
nor NOR3 (N1827, N1825, N540, N1541);
or OR3 (N1828, N1818, N1758, N1125);
nor NOR2 (N1829, N1826, N1405);
nor NOR4 (N1830, N1828, N133, N437, N1026);
or OR2 (N1831, N1793, N1399);
nor NOR2 (N1832, N1824, N566);
buf BUF1 (N1833, N1829);
buf BUF1 (N1834, N1830);
or OR2 (N1835, N1827, N1644);
nand NAND2 (N1836, N1834, N507);
or OR2 (N1837, N1810, N780);
or OR2 (N1838, N1835, N1629);
and AND3 (N1839, N1837, N1812, N537);
buf BUF1 (N1840, N1838);
nor NOR2 (N1841, N1836, N1749);
or OR4 (N1842, N1823, N1170, N761, N412);
nor NOR3 (N1843, N1841, N1624, N1811);
nand NAND3 (N1844, N1839, N325, N797);
xor XOR2 (N1845, N1833, N1265);
nand NAND3 (N1846, N1796, N1365, N127);
nor NOR3 (N1847, N1842, N1155, N1761);
not NOT1 (N1848, N1845);
or OR2 (N1849, N1843, N1478);
xor XOR2 (N1850, N1848, N1152);
nor NOR2 (N1851, N1850, N1212);
nand NAND3 (N1852, N1847, N81, N1119);
nor NOR4 (N1853, N1840, N1310, N80, N1663);
nor NOR2 (N1854, N1832, N1022);
nand NAND4 (N1855, N1854, N321, N1228, N1591);
xor XOR2 (N1856, N1852, N1141);
nand NAND2 (N1857, N1853, N1806);
buf BUF1 (N1858, N1855);
not NOT1 (N1859, N1856);
not NOT1 (N1860, N1844);
buf BUF1 (N1861, N1821);
not NOT1 (N1862, N1851);
buf BUF1 (N1863, N1860);
not NOT1 (N1864, N1859);
buf BUF1 (N1865, N1831);
or OR2 (N1866, N1864, N1529);
xor XOR2 (N1867, N1866, N1777);
and AND3 (N1868, N1846, N380, N801);
not NOT1 (N1869, N1863);
nor NOR4 (N1870, N1868, N840, N104, N1606);
nor NOR4 (N1871, N1870, N1388, N1128, N135);
nand NAND4 (N1872, N1861, N679, N1327, N430);
and AND2 (N1873, N1858, N1672);
nand NAND3 (N1874, N1857, N112, N561);
nor NOR3 (N1875, N1820, N1372, N1844);
nor NOR3 (N1876, N1862, N707, N178);
nor NOR2 (N1877, N1872, N1391);
buf BUF1 (N1878, N1875);
nand NAND3 (N1879, N1874, N534, N1054);
nor NOR3 (N1880, N1876, N1004, N721);
xor XOR2 (N1881, N1877, N21);
xor XOR2 (N1882, N1849, N243);
or OR2 (N1883, N1873, N1829);
not NOT1 (N1884, N1883);
not NOT1 (N1885, N1881);
xor XOR2 (N1886, N1882, N287);
and AND2 (N1887, N1885, N943);
not NOT1 (N1888, N1865);
or OR3 (N1889, N1887, N1266, N931);
and AND4 (N1890, N1888, N611, N789, N55);
not NOT1 (N1891, N1867);
not NOT1 (N1892, N1886);
nor NOR3 (N1893, N1890, N1652, N1611);
buf BUF1 (N1894, N1891);
nand NAND4 (N1895, N1869, N168, N508, N1007);
and AND4 (N1896, N1884, N321, N26, N16);
or OR3 (N1897, N1892, N1159, N1353);
or OR4 (N1898, N1894, N849, N430, N574);
buf BUF1 (N1899, N1871);
not NOT1 (N1900, N1897);
nand NAND2 (N1901, N1893, N1671);
buf BUF1 (N1902, N1880);
nor NOR3 (N1903, N1878, N844, N146);
not NOT1 (N1904, N1898);
and AND3 (N1905, N1896, N1523, N577);
nor NOR2 (N1906, N1903, N965);
buf BUF1 (N1907, N1889);
xor XOR2 (N1908, N1879, N1859);
xor XOR2 (N1909, N1908, N523);
and AND4 (N1910, N1904, N868, N288, N1873);
or OR2 (N1911, N1910, N1492);
and AND4 (N1912, N1907, N1788, N1840, N911);
buf BUF1 (N1913, N1905);
xor XOR2 (N1914, N1900, N1767);
nor NOR3 (N1915, N1909, N975, N394);
xor XOR2 (N1916, N1914, N390);
buf BUF1 (N1917, N1913);
buf BUF1 (N1918, N1906);
xor XOR2 (N1919, N1912, N1669);
nor NOR3 (N1920, N1895, N1537, N832);
nor NOR3 (N1921, N1899, N1302, N794);
not NOT1 (N1922, N1917);
buf BUF1 (N1923, N1920);
nand NAND3 (N1924, N1923, N1297, N1032);
or OR2 (N1925, N1918, N1214);
buf BUF1 (N1926, N1924);
nor NOR2 (N1927, N1902, N1449);
and AND3 (N1928, N1916, N1196, N75);
nor NOR3 (N1929, N1915, N1495, N142);
and AND2 (N1930, N1928, N1300);
nor NOR2 (N1931, N1919, N765);
not NOT1 (N1932, N1927);
not NOT1 (N1933, N1925);
or OR3 (N1934, N1933, N1854, N120);
buf BUF1 (N1935, N1930);
nor NOR2 (N1936, N1922, N857);
and AND2 (N1937, N1921, N1445);
nand NAND3 (N1938, N1901, N1006, N150);
xor XOR2 (N1939, N1934, N1790);
buf BUF1 (N1940, N1926);
nor NOR2 (N1941, N1935, N1442);
not NOT1 (N1942, N1932);
not NOT1 (N1943, N1931);
nand NAND4 (N1944, N1941, N769, N857, N1425);
xor XOR2 (N1945, N1911, N1280);
not NOT1 (N1946, N1936);
or OR4 (N1947, N1929, N1024, N43, N236);
not NOT1 (N1948, N1944);
nor NOR4 (N1949, N1947, N1798, N645, N1371);
not NOT1 (N1950, N1940);
nor NOR2 (N1951, N1945, N223);
and AND2 (N1952, N1937, N267);
nand NAND2 (N1953, N1939, N1600);
not NOT1 (N1954, N1948);
or OR4 (N1955, N1946, N1429, N1696, N1885);
buf BUF1 (N1956, N1952);
and AND4 (N1957, N1943, N948, N1952, N574);
not NOT1 (N1958, N1942);
nand NAND4 (N1959, N1950, N1016, N26, N1129);
buf BUF1 (N1960, N1959);
buf BUF1 (N1961, N1954);
buf BUF1 (N1962, N1957);
xor XOR2 (N1963, N1953, N53);
xor XOR2 (N1964, N1961, N754);
buf BUF1 (N1965, N1955);
buf BUF1 (N1966, N1951);
not NOT1 (N1967, N1966);
and AND3 (N1968, N1938, N10, N54);
or OR3 (N1969, N1960, N154, N1930);
buf BUF1 (N1970, N1963);
nor NOR3 (N1971, N1968, N603, N1004);
nor NOR4 (N1972, N1971, N151, N29, N500);
nand NAND2 (N1973, N1970, N1510);
nor NOR2 (N1974, N1949, N287);
buf BUF1 (N1975, N1962);
nor NOR2 (N1976, N1972, N1866);
buf BUF1 (N1977, N1958);
buf BUF1 (N1978, N1967);
xor XOR2 (N1979, N1978, N1364);
and AND4 (N1980, N1964, N369, N44, N993);
nand NAND4 (N1981, N1975, N1125, N144, N1471);
nand NAND4 (N1982, N1976, N8, N1959, N1933);
xor XOR2 (N1983, N1982, N1428);
and AND3 (N1984, N1973, N802, N391);
nor NOR4 (N1985, N1981, N1606, N1617, N853);
nand NAND2 (N1986, N1984, N1256);
or OR4 (N1987, N1977, N887, N860, N622);
xor XOR2 (N1988, N1987, N843);
xor XOR2 (N1989, N1965, N1721);
nor NOR4 (N1990, N1983, N1196, N40, N629);
buf BUF1 (N1991, N1974);
xor XOR2 (N1992, N1969, N212);
or OR4 (N1993, N1979, N881, N1422, N1391);
not NOT1 (N1994, N1991);
and AND2 (N1995, N1986, N94);
nor NOR3 (N1996, N1994, N1847, N1974);
xor XOR2 (N1997, N1990, N1780);
nor NOR4 (N1998, N1988, N1699, N1182, N791);
buf BUF1 (N1999, N1993);
xor XOR2 (N2000, N1997, N386);
nand NAND2 (N2001, N1992, N784);
and AND4 (N2002, N1980, N1262, N984, N1832);
buf BUF1 (N2003, N1998);
nand NAND3 (N2004, N1985, N1929, N288);
nand NAND4 (N2005, N2002, N113, N1232, N1476);
or OR3 (N2006, N2005, N1560, N1969);
nand NAND2 (N2007, N2001, N1274);
and AND4 (N2008, N2000, N1992, N1840, N1982);
buf BUF1 (N2009, N2003);
buf BUF1 (N2010, N2004);
not NOT1 (N2011, N2006);
and AND3 (N2012, N1996, N799, N1963);
not NOT1 (N2013, N2010);
xor XOR2 (N2014, N1995, N2013);
and AND3 (N2015, N728, N1824, N1397);
or OR3 (N2016, N1956, N1097, N1570);
buf BUF1 (N2017, N2011);
buf BUF1 (N2018, N2016);
not NOT1 (N2019, N2009);
nand NAND3 (N2020, N1989, N1979, N1366);
nor NOR3 (N2021, N2012, N1818, N1790);
buf BUF1 (N2022, N2018);
nand NAND2 (N2023, N1999, N1233);
nor NOR3 (N2024, N2008, N1474, N1255);
or OR3 (N2025, N2023, N1191, N499);
not NOT1 (N2026, N2024);
buf BUF1 (N2027, N2021);
nand NAND3 (N2028, N2020, N153, N1424);
not NOT1 (N2029, N2015);
buf BUF1 (N2030, N2017);
or OR4 (N2031, N2014, N1329, N724, N1724);
buf BUF1 (N2032, N2029);
or OR3 (N2033, N2031, N1993, N1385);
nand NAND2 (N2034, N2027, N1273);
or OR2 (N2035, N2032, N1142);
and AND2 (N2036, N2028, N638);
xor XOR2 (N2037, N2036, N1132);
or OR4 (N2038, N2022, N1496, N1509, N13);
or OR3 (N2039, N2025, N845, N296);
buf BUF1 (N2040, N2026);
nand NAND4 (N2041, N2030, N511, N591, N401);
not NOT1 (N2042, N2033);
nor NOR2 (N2043, N2040, N623);
nand NAND2 (N2044, N2039, N770);
buf BUF1 (N2045, N2038);
xor XOR2 (N2046, N2044, N1450);
xor XOR2 (N2047, N2045, N149);
not NOT1 (N2048, N2034);
or OR2 (N2049, N2035, N738);
xor XOR2 (N2050, N2019, N1004);
and AND3 (N2051, N2037, N1988, N491);
nor NOR2 (N2052, N2047, N1971);
buf BUF1 (N2053, N2052);
xor XOR2 (N2054, N2050, N1969);
or OR3 (N2055, N2043, N466, N1514);
xor XOR2 (N2056, N2007, N1403);
or OR2 (N2057, N2051, N1534);
xor XOR2 (N2058, N2049, N363);
or OR2 (N2059, N2041, N1762);
xor XOR2 (N2060, N2053, N780);
and AND2 (N2061, N2042, N1917);
or OR4 (N2062, N2059, N1506, N1146, N1558);
buf BUF1 (N2063, N2061);
not NOT1 (N2064, N2048);
nor NOR3 (N2065, N2063, N878, N1866);
and AND2 (N2066, N2064, N1884);
xor XOR2 (N2067, N2055, N101);
buf BUF1 (N2068, N2058);
or OR2 (N2069, N2068, N713);
nand NAND2 (N2070, N2054, N1161);
or OR3 (N2071, N2046, N1639, N950);
and AND3 (N2072, N2066, N782, N461);
and AND3 (N2073, N2062, N1653, N737);
not NOT1 (N2074, N2060);
or OR3 (N2075, N2069, N660, N1046);
not NOT1 (N2076, N2075);
and AND2 (N2077, N2073, N1608);
not NOT1 (N2078, N2077);
not NOT1 (N2079, N2072);
nand NAND3 (N2080, N2079, N1072, N1355);
not NOT1 (N2081, N2067);
xor XOR2 (N2082, N2071, N571);
and AND3 (N2083, N2081, N2031, N1998);
xor XOR2 (N2084, N2080, N840);
nor NOR2 (N2085, N2076, N866);
xor XOR2 (N2086, N2082, N1002);
nor NOR2 (N2087, N2086, N1593);
and AND2 (N2088, N2074, N1012);
nor NOR4 (N2089, N2057, N510, N1064, N1508);
nor NOR3 (N2090, N2070, N867, N2022);
or OR3 (N2091, N2089, N1770, N805);
xor XOR2 (N2092, N2090, N1345);
buf BUF1 (N2093, N2084);
nand NAND4 (N2094, N2083, N1432, N646, N2012);
and AND3 (N2095, N2094, N1072, N489);
or OR4 (N2096, N2056, N628, N1468, N1980);
and AND3 (N2097, N2078, N257, N1646);
and AND3 (N2098, N2088, N1771, N1310);
and AND4 (N2099, N2093, N1458, N1804, N1745);
nand NAND4 (N2100, N2095, N976, N1766, N1765);
xor XOR2 (N2101, N2091, N368);
nor NOR4 (N2102, N2099, N1099, N1370, N2089);
buf BUF1 (N2103, N2100);
xor XOR2 (N2104, N2087, N968);
or OR2 (N2105, N2092, N76);
xor XOR2 (N2106, N2104, N1837);
buf BUF1 (N2107, N2105);
and AND3 (N2108, N2102, N623, N1538);
not NOT1 (N2109, N2101);
xor XOR2 (N2110, N2103, N440);
and AND2 (N2111, N2110, N725);
xor XOR2 (N2112, N2108, N1776);
xor XOR2 (N2113, N2107, N1413);
not NOT1 (N2114, N2085);
xor XOR2 (N2115, N2113, N1602);
nor NOR3 (N2116, N2106, N573, N60);
xor XOR2 (N2117, N2111, N315);
nand NAND4 (N2118, N2097, N1586, N1147, N1182);
not NOT1 (N2119, N2114);
nand NAND3 (N2120, N2096, N1123, N544);
buf BUF1 (N2121, N2109);
and AND2 (N2122, N2098, N615);
and AND3 (N2123, N2120, N501, N1375);
not NOT1 (N2124, N2065);
nor NOR4 (N2125, N2115, N19, N1152, N1767);
or OR3 (N2126, N2119, N1991, N959);
xor XOR2 (N2127, N2125, N481);
nand NAND3 (N2128, N2116, N851, N1695);
and AND4 (N2129, N2127, N1532, N89, N973);
or OR3 (N2130, N2128, N1506, N1800);
and AND2 (N2131, N2122, N789);
not NOT1 (N2132, N2129);
not NOT1 (N2133, N2123);
or OR3 (N2134, N2132, N633, N423);
not NOT1 (N2135, N2134);
nand NAND3 (N2136, N2130, N681, N1101);
or OR3 (N2137, N2126, N747, N90);
xor XOR2 (N2138, N2136, N1690);
buf BUF1 (N2139, N2138);
and AND3 (N2140, N2124, N1628, N865);
nor NOR4 (N2141, N2118, N735, N833, N184);
nor NOR3 (N2142, N2117, N1711, N265);
and AND3 (N2143, N2135, N452, N541);
and AND4 (N2144, N2140, N850, N594, N1112);
xor XOR2 (N2145, N2121, N202);
buf BUF1 (N2146, N2131);
and AND4 (N2147, N2139, N1292, N347, N134);
and AND4 (N2148, N2146, N483, N1677, N1081);
nand NAND3 (N2149, N2143, N391, N1178);
nand NAND3 (N2150, N2144, N1236, N391);
and AND3 (N2151, N2149, N816, N129);
not NOT1 (N2152, N2141);
or OR4 (N2153, N2151, N1771, N908, N640);
or OR4 (N2154, N2142, N2141, N1476, N1663);
and AND4 (N2155, N2148, N59, N1979, N1748);
not NOT1 (N2156, N2147);
not NOT1 (N2157, N2145);
buf BUF1 (N2158, N2133);
nor NOR2 (N2159, N2150, N482);
not NOT1 (N2160, N2112);
or OR2 (N2161, N2156, N1870);
or OR3 (N2162, N2160, N1155, N496);
xor XOR2 (N2163, N2152, N102);
and AND3 (N2164, N2154, N632, N2112);
or OR4 (N2165, N2159, N1535, N998, N672);
and AND4 (N2166, N2165, N1540, N726, N1485);
or OR4 (N2167, N2162, N463, N984, N617);
not NOT1 (N2168, N2158);
buf BUF1 (N2169, N2168);
and AND3 (N2170, N2163, N2074, N1833);
xor XOR2 (N2171, N2166, N1463);
or OR3 (N2172, N2164, N1960, N462);
not NOT1 (N2173, N2153);
buf BUF1 (N2174, N2157);
or OR3 (N2175, N2161, N831, N1319);
buf BUF1 (N2176, N2174);
and AND4 (N2177, N2172, N614, N150, N1454);
buf BUF1 (N2178, N2155);
and AND3 (N2179, N2177, N335, N348);
nor NOR4 (N2180, N2179, N2063, N810, N1854);
or OR2 (N2181, N2175, N2156);
and AND4 (N2182, N2137, N495, N1272, N1169);
or OR3 (N2183, N2181, N459, N1687);
xor XOR2 (N2184, N2180, N1328);
buf BUF1 (N2185, N2176);
and AND2 (N2186, N2169, N91);
not NOT1 (N2187, N2184);
not NOT1 (N2188, N2167);
xor XOR2 (N2189, N2183, N669);
xor XOR2 (N2190, N2185, N467);
or OR2 (N2191, N2178, N230);
nand NAND2 (N2192, N2190, N2127);
nand NAND2 (N2193, N2182, N1023);
nand NAND3 (N2194, N2187, N1049, N2192);
xor XOR2 (N2195, N859, N479);
buf BUF1 (N2196, N2193);
nor NOR3 (N2197, N2188, N1840, N139);
and AND2 (N2198, N2186, N225);
and AND3 (N2199, N2198, N694, N74);
nor NOR2 (N2200, N2189, N727);
and AND4 (N2201, N2194, N1282, N1625, N510);
or OR3 (N2202, N2170, N1217, N1901);
nand NAND4 (N2203, N2191, N441, N1452, N1736);
not NOT1 (N2204, N2195);
not NOT1 (N2205, N2203);
and AND2 (N2206, N2173, N227);
or OR2 (N2207, N2201, N273);
or OR3 (N2208, N2197, N867, N1642);
nand NAND2 (N2209, N2206, N2076);
xor XOR2 (N2210, N2207, N917);
nand NAND3 (N2211, N2171, N1178, N265);
nor NOR4 (N2212, N2204, N2162, N1578, N2101);
nand NAND3 (N2213, N2212, N1497, N1092);
and AND4 (N2214, N2211, N1640, N491, N1285);
nor NOR2 (N2215, N2210, N668);
or OR4 (N2216, N2208, N2075, N1180, N325);
not NOT1 (N2217, N2214);
nand NAND2 (N2218, N2205, N1788);
xor XOR2 (N2219, N2218, N397);
nor NOR4 (N2220, N2209, N835, N441, N631);
not NOT1 (N2221, N2215);
or OR2 (N2222, N2216, N905);
not NOT1 (N2223, N2196);
nand NAND2 (N2224, N2217, N874);
nor NOR2 (N2225, N2220, N708);
nand NAND3 (N2226, N2213, N502, N1490);
nand NAND4 (N2227, N2223, N1613, N1819, N1191);
xor XOR2 (N2228, N2224, N1856);
nor NOR2 (N2229, N2225, N1656);
or OR4 (N2230, N2227, N255, N1263, N952);
and AND3 (N2231, N2230, N864, N734);
xor XOR2 (N2232, N2200, N1789);
or OR2 (N2233, N2228, N935);
or OR2 (N2234, N2233, N60);
buf BUF1 (N2235, N2219);
nand NAND4 (N2236, N2235, N766, N566, N1526);
not NOT1 (N2237, N2229);
nand NAND2 (N2238, N2222, N912);
xor XOR2 (N2239, N2238, N2059);
nor NOR3 (N2240, N2226, N902, N1056);
and AND2 (N2241, N2237, N707);
buf BUF1 (N2242, N2231);
buf BUF1 (N2243, N2221);
not NOT1 (N2244, N2202);
buf BUF1 (N2245, N2241);
or OR3 (N2246, N2199, N1497, N2206);
and AND2 (N2247, N2244, N693);
buf BUF1 (N2248, N2243);
nand NAND3 (N2249, N2234, N1488, N960);
nor NOR3 (N2250, N2245, N1191, N1271);
or OR4 (N2251, N2249, N312, N1510, N1529);
or OR4 (N2252, N2248, N14, N1315, N1130);
and AND3 (N2253, N2250, N1546, N949);
and AND4 (N2254, N2239, N1402, N732, N852);
nor NOR2 (N2255, N2246, N1288);
and AND2 (N2256, N2255, N444);
buf BUF1 (N2257, N2252);
and AND3 (N2258, N2232, N1217, N662);
and AND2 (N2259, N2242, N1476);
nor NOR2 (N2260, N2251, N480);
nand NAND2 (N2261, N2240, N1292);
nor NOR3 (N2262, N2256, N1663, N2002);
and AND2 (N2263, N2257, N2112);
not NOT1 (N2264, N2254);
and AND2 (N2265, N2260, N1781);
nor NOR2 (N2266, N2259, N366);
nor NOR2 (N2267, N2264, N38);
buf BUF1 (N2268, N2247);
nand NAND3 (N2269, N2258, N1378, N1264);
buf BUF1 (N2270, N2265);
nor NOR2 (N2271, N2253, N975);
and AND4 (N2272, N2262, N1006, N527, N1917);
nor NOR4 (N2273, N2270, N1922, N911, N1965);
not NOT1 (N2274, N2269);
xor XOR2 (N2275, N2267, N1435);
or OR2 (N2276, N2236, N1360);
nand NAND2 (N2277, N2273, N1213);
nand NAND4 (N2278, N2274, N2218, N901, N1126);
nand NAND3 (N2279, N2271, N1001, N1609);
nor NOR2 (N2280, N2279, N68);
xor XOR2 (N2281, N2278, N1531);
xor XOR2 (N2282, N2281, N703);
nor NOR4 (N2283, N2276, N876, N2137, N1287);
buf BUF1 (N2284, N2272);
and AND4 (N2285, N2277, N2199, N268, N907);
nor NOR4 (N2286, N2266, N1283, N2077, N1150);
not NOT1 (N2287, N2280);
nor NOR4 (N2288, N2287, N2110, N1140, N481);
and AND3 (N2289, N2284, N2158, N2150);
xor XOR2 (N2290, N2282, N2120);
nand NAND4 (N2291, N2290, N1891, N656, N1630);
xor XOR2 (N2292, N2285, N202);
or OR2 (N2293, N2292, N2095);
xor XOR2 (N2294, N2263, N1639);
and AND4 (N2295, N2268, N400, N1680, N630);
not NOT1 (N2296, N2291);
not NOT1 (N2297, N2288);
buf BUF1 (N2298, N2283);
xor XOR2 (N2299, N2294, N996);
nand NAND3 (N2300, N2261, N93, N1614);
nand NAND4 (N2301, N2299, N1476, N1008, N555);
not NOT1 (N2302, N2275);
and AND3 (N2303, N2293, N1192, N1990);
or OR3 (N2304, N2286, N1421, N211);
or OR2 (N2305, N2297, N1346);
nand NAND4 (N2306, N2300, N1760, N79, N1471);
nor NOR2 (N2307, N2305, N74);
and AND4 (N2308, N2307, N200, N1055, N1309);
not NOT1 (N2309, N2296);
not NOT1 (N2310, N2298);
xor XOR2 (N2311, N2310, N1859);
buf BUF1 (N2312, N2309);
and AND3 (N2313, N2289, N395, N1812);
nand NAND2 (N2314, N2313, N1774);
or OR3 (N2315, N2301, N1901, N1755);
not NOT1 (N2316, N2311);
nor NOR4 (N2317, N2312, N1412, N1727, N1564);
xor XOR2 (N2318, N2314, N1428);
and AND4 (N2319, N2306, N968, N1289, N1998);
xor XOR2 (N2320, N2304, N321);
not NOT1 (N2321, N2295);
or OR4 (N2322, N2303, N1312, N2189, N980);
buf BUF1 (N2323, N2317);
not NOT1 (N2324, N2319);
not NOT1 (N2325, N2308);
not NOT1 (N2326, N2318);
nand NAND2 (N2327, N2315, N225);
buf BUF1 (N2328, N2327);
buf BUF1 (N2329, N2328);
not NOT1 (N2330, N2326);
not NOT1 (N2331, N2330);
and AND4 (N2332, N2325, N2018, N1243, N1868);
nand NAND2 (N2333, N2321, N934);
or OR4 (N2334, N2324, N2320, N1620, N1401);
nor NOR3 (N2335, N1020, N2212, N1568);
not NOT1 (N2336, N2335);
nor NOR4 (N2337, N2316, N1983, N681, N1508);
nand NAND2 (N2338, N2332, N1005);
xor XOR2 (N2339, N2322, N1913);
nand NAND3 (N2340, N2323, N5, N160);
buf BUF1 (N2341, N2334);
or OR3 (N2342, N2340, N904, N1967);
not NOT1 (N2343, N2339);
xor XOR2 (N2344, N2337, N16);
buf BUF1 (N2345, N2336);
or OR3 (N2346, N2338, N2142, N647);
buf BUF1 (N2347, N2331);
not NOT1 (N2348, N2329);
and AND3 (N2349, N2333, N567, N337);
not NOT1 (N2350, N2341);
or OR3 (N2351, N2302, N945, N684);
not NOT1 (N2352, N2342);
nor NOR4 (N2353, N2343, N554, N2118, N221);
or OR3 (N2354, N2351, N815, N33);
or OR4 (N2355, N2354, N490, N1179, N33);
or OR4 (N2356, N2352, N295, N83, N1725);
and AND2 (N2357, N2355, N1870);
and AND2 (N2358, N2348, N1572);
nand NAND3 (N2359, N2357, N493, N1781);
nor NOR4 (N2360, N2350, N1932, N676, N241);
and AND2 (N2361, N2344, N805);
or OR2 (N2362, N2356, N1038);
nand NAND3 (N2363, N2358, N2289, N1254);
not NOT1 (N2364, N2349);
and AND3 (N2365, N2353, N2211, N2273);
buf BUF1 (N2366, N2360);
xor XOR2 (N2367, N2363, N648);
xor XOR2 (N2368, N2347, N1555);
not NOT1 (N2369, N2365);
nor NOR4 (N2370, N2346, N74, N989, N113);
not NOT1 (N2371, N2370);
nor NOR3 (N2372, N2361, N1351, N2280);
buf BUF1 (N2373, N2367);
or OR2 (N2374, N2371, N155);
or OR2 (N2375, N2372, N829);
or OR3 (N2376, N2364, N508, N220);
buf BUF1 (N2377, N2368);
and AND3 (N2378, N2373, N187, N1663);
and AND3 (N2379, N2359, N1674, N2162);
or OR3 (N2380, N2369, N257, N1197);
or OR4 (N2381, N2376, N2194, N978, N1025);
or OR3 (N2382, N2375, N2268, N1849);
xor XOR2 (N2383, N2380, N704);
nor NOR3 (N2384, N2374, N1794, N1817);
not NOT1 (N2385, N2345);
buf BUF1 (N2386, N2379);
nor NOR3 (N2387, N2377, N735, N780);
nor NOR2 (N2388, N2378, N757);
nand NAND2 (N2389, N2366, N521);
or OR2 (N2390, N2381, N566);
and AND3 (N2391, N2387, N689, N1015);
buf BUF1 (N2392, N2383);
xor XOR2 (N2393, N2388, N1205);
buf BUF1 (N2394, N2393);
buf BUF1 (N2395, N2390);
nand NAND2 (N2396, N2382, N619);
or OR2 (N2397, N2389, N137);
nor NOR2 (N2398, N2395, N1635);
not NOT1 (N2399, N2391);
buf BUF1 (N2400, N2396);
nor NOR4 (N2401, N2399, N226, N2398, N943);
xor XOR2 (N2402, N2110, N186);
nand NAND2 (N2403, N2400, N569);
not NOT1 (N2404, N2362);
buf BUF1 (N2405, N2392);
or OR4 (N2406, N2386, N751, N1461, N202);
nand NAND4 (N2407, N2397, N171, N2193, N416);
nor NOR2 (N2408, N2406, N276);
and AND2 (N2409, N2402, N1355);
nor NOR2 (N2410, N2404, N197);
nand NAND3 (N2411, N2407, N1238, N2031);
or OR2 (N2412, N2409, N387);
nand NAND4 (N2413, N2410, N577, N1989, N780);
xor XOR2 (N2414, N2384, N2330);
or OR2 (N2415, N2405, N407);
and AND4 (N2416, N2401, N144, N2240, N1657);
or OR4 (N2417, N2412, N1702, N468, N1347);
nand NAND2 (N2418, N2403, N308);
xor XOR2 (N2419, N2417, N1470);
or OR2 (N2420, N2394, N649);
and AND2 (N2421, N2411, N989);
and AND3 (N2422, N2416, N1732, N967);
xor XOR2 (N2423, N2414, N724);
nor NOR4 (N2424, N2408, N1469, N2422, N1898);
buf BUF1 (N2425, N1884);
or OR3 (N2426, N2425, N841, N2349);
xor XOR2 (N2427, N2413, N1898);
or OR3 (N2428, N2424, N639, N1522);
not NOT1 (N2429, N2418);
and AND2 (N2430, N2385, N690);
buf BUF1 (N2431, N2419);
nand NAND2 (N2432, N2423, N2126);
nand NAND3 (N2433, N2426, N1672, N946);
nand NAND3 (N2434, N2420, N679, N2035);
xor XOR2 (N2435, N2421, N2372);
and AND3 (N2436, N2428, N1187, N2212);
nand NAND4 (N2437, N2435, N772, N1162, N97);
xor XOR2 (N2438, N2431, N1742);
buf BUF1 (N2439, N2437);
nor NOR4 (N2440, N2436, N447, N889, N1798);
xor XOR2 (N2441, N2434, N2160);
not NOT1 (N2442, N2440);
xor XOR2 (N2443, N2430, N210);
not NOT1 (N2444, N2433);
or OR3 (N2445, N2439, N1745, N697);
buf BUF1 (N2446, N2429);
nor NOR2 (N2447, N2441, N1252);
not NOT1 (N2448, N2444);
and AND3 (N2449, N2446, N1758, N1241);
xor XOR2 (N2450, N2449, N1893);
buf BUF1 (N2451, N2438);
xor XOR2 (N2452, N2447, N1484);
buf BUF1 (N2453, N2427);
nor NOR4 (N2454, N2442, N1021, N323, N1599);
nor NOR4 (N2455, N2450, N2066, N214, N1731);
nand NAND2 (N2456, N2415, N2219);
nor NOR3 (N2457, N2453, N240, N925);
nor NOR2 (N2458, N2448, N1378);
xor XOR2 (N2459, N2443, N331);
nor NOR2 (N2460, N2452, N244);
xor XOR2 (N2461, N2460, N2427);
nor NOR2 (N2462, N2458, N819);
not NOT1 (N2463, N2432);
buf BUF1 (N2464, N2445);
not NOT1 (N2465, N2455);
or OR3 (N2466, N2451, N536, N1149);
or OR4 (N2467, N2463, N1234, N1020, N856);
nand NAND4 (N2468, N2464, N2446, N1470, N794);
buf BUF1 (N2469, N2457);
xor XOR2 (N2470, N2465, N1217);
not NOT1 (N2471, N2466);
buf BUF1 (N2472, N2459);
or OR3 (N2473, N2462, N1148, N2382);
nand NAND4 (N2474, N2473, N2053, N1674, N1424);
nand NAND3 (N2475, N2461, N2322, N967);
xor XOR2 (N2476, N2468, N1973);
nor NOR4 (N2477, N2471, N1776, N771, N669);
or OR4 (N2478, N2454, N470, N4, N1323);
buf BUF1 (N2479, N2467);
not NOT1 (N2480, N2470);
or OR4 (N2481, N2479, N2066, N1379, N547);
buf BUF1 (N2482, N2478);
nand NAND4 (N2483, N2456, N294, N1919, N783);
buf BUF1 (N2484, N2475);
and AND3 (N2485, N2469, N2354, N1111);
nand NAND3 (N2486, N2483, N1333, N2434);
and AND2 (N2487, N2476, N2076);
xor XOR2 (N2488, N2474, N498);
xor XOR2 (N2489, N2488, N139);
nor NOR4 (N2490, N2486, N371, N1748, N1493);
buf BUF1 (N2491, N2472);
not NOT1 (N2492, N2480);
and AND3 (N2493, N2482, N1228, N613);
and AND2 (N2494, N2485, N590);
not NOT1 (N2495, N2489);
and AND3 (N2496, N2492, N1460, N590);
buf BUF1 (N2497, N2493);
not NOT1 (N2498, N2494);
not NOT1 (N2499, N2484);
nand NAND3 (N2500, N2491, N1583, N1299);
and AND4 (N2501, N2481, N189, N2271, N2382);
and AND2 (N2502, N2495, N1058);
nand NAND3 (N2503, N2500, N271, N1207);
not NOT1 (N2504, N2496);
xor XOR2 (N2505, N2503, N70);
nand NAND3 (N2506, N2487, N1368, N109);
and AND4 (N2507, N2490, N2298, N1149, N1938);
buf BUF1 (N2508, N2506);
xor XOR2 (N2509, N2477, N2291);
buf BUF1 (N2510, N2507);
and AND4 (N2511, N2504, N2212, N2212, N193);
xor XOR2 (N2512, N2501, N114);
or OR4 (N2513, N2497, N1111, N577, N924);
xor XOR2 (N2514, N2511, N979);
and AND2 (N2515, N2508, N1773);
nor NOR4 (N2516, N2499, N2249, N1840, N264);
nor NOR2 (N2517, N2509, N1887);
buf BUF1 (N2518, N2516);
nand NAND4 (N2519, N2505, N665, N2011, N545);
xor XOR2 (N2520, N2498, N2043);
and AND2 (N2521, N2520, N2249);
and AND4 (N2522, N2517, N1305, N453, N868);
nor NOR2 (N2523, N2513, N406);
and AND4 (N2524, N2514, N2472, N782, N1618);
or OR4 (N2525, N2521, N2388, N403, N1917);
or OR2 (N2526, N2523, N1394);
not NOT1 (N2527, N2519);
not NOT1 (N2528, N2526);
and AND3 (N2529, N2515, N647, N285);
buf BUF1 (N2530, N2529);
and AND3 (N2531, N2502, N398, N2080);
and AND4 (N2532, N2525, N328, N452, N1074);
and AND4 (N2533, N2531, N2060, N2381, N1691);
nand NAND3 (N2534, N2524, N251, N2423);
not NOT1 (N2535, N2512);
and AND2 (N2536, N2532, N181);
nor NOR2 (N2537, N2528, N210);
xor XOR2 (N2538, N2537, N2503);
buf BUF1 (N2539, N2535);
buf BUF1 (N2540, N2510);
nand NAND4 (N2541, N2539, N2268, N758, N1950);
not NOT1 (N2542, N2522);
or OR3 (N2543, N2536, N269, N2355);
nor NOR3 (N2544, N2542, N2210, N338);
not NOT1 (N2545, N2530);
nand NAND2 (N2546, N2540, N1442);
nor NOR2 (N2547, N2534, N2106);
not NOT1 (N2548, N2545);
and AND4 (N2549, N2541, N819, N236, N1711);
buf BUF1 (N2550, N2543);
nor NOR3 (N2551, N2533, N178, N764);
and AND3 (N2552, N2549, N1282, N469);
nand NAND3 (N2553, N2546, N1245, N234);
xor XOR2 (N2554, N2553, N394);
and AND3 (N2555, N2538, N1447, N611);
nor NOR3 (N2556, N2547, N2279, N455);
and AND3 (N2557, N2548, N691, N1528);
nor NOR4 (N2558, N2556, N1132, N1812, N645);
nor NOR4 (N2559, N2527, N2262, N2062, N1862);
buf BUF1 (N2560, N2544);
nor NOR4 (N2561, N2550, N2556, N594, N1577);
or OR4 (N2562, N2554, N1430, N217, N1083);
not NOT1 (N2563, N2559);
nor NOR4 (N2564, N2551, N1547, N260, N2312);
and AND2 (N2565, N2555, N1586);
not NOT1 (N2566, N2560);
or OR4 (N2567, N2565, N2062, N2538, N2379);
buf BUF1 (N2568, N2563);
buf BUF1 (N2569, N2552);
not NOT1 (N2570, N2567);
nor NOR3 (N2571, N2568, N944, N333);
xor XOR2 (N2572, N2564, N1882);
nand NAND2 (N2573, N2561, N785);
or OR3 (N2574, N2562, N2266, N1759);
and AND4 (N2575, N2574, N2226, N2310, N1102);
nor NOR4 (N2576, N2570, N90, N1130, N2053);
not NOT1 (N2577, N2572);
nor NOR4 (N2578, N2518, N554, N969, N706);
and AND4 (N2579, N2575, N1773, N2185, N289);
not NOT1 (N2580, N2558);
nand NAND2 (N2581, N2571, N2514);
and AND4 (N2582, N2566, N1157, N202, N1283);
xor XOR2 (N2583, N2580, N1635);
nand NAND2 (N2584, N2577, N2411);
buf BUF1 (N2585, N2582);
not NOT1 (N2586, N2557);
and AND4 (N2587, N2583, N2494, N715, N1985);
or OR3 (N2588, N2587, N2257, N1648);
not NOT1 (N2589, N2576);
and AND3 (N2590, N2579, N28, N2362);
xor XOR2 (N2591, N2573, N1881);
nor NOR4 (N2592, N2581, N1007, N689, N856);
nand NAND4 (N2593, N2586, N1319, N66, N296);
or OR3 (N2594, N2578, N1382, N666);
buf BUF1 (N2595, N2593);
xor XOR2 (N2596, N2591, N1060);
or OR3 (N2597, N2589, N653, N1095);
nor NOR4 (N2598, N2592, N1581, N2189, N1210);
xor XOR2 (N2599, N2590, N1378);
not NOT1 (N2600, N2597);
xor XOR2 (N2601, N2598, N2402);
and AND3 (N2602, N2599, N265, N2000);
buf BUF1 (N2603, N2600);
nor NOR3 (N2604, N2595, N2157, N2384);
and AND3 (N2605, N2601, N1658, N2272);
not NOT1 (N2606, N2584);
not NOT1 (N2607, N2585);
nor NOR2 (N2608, N2594, N2374);
nor NOR4 (N2609, N2569, N388, N1000, N317);
nor NOR4 (N2610, N2609, N1001, N1215, N57);
nor NOR2 (N2611, N2607, N1689);
nand NAND4 (N2612, N2608, N1115, N1935, N637);
and AND2 (N2613, N2603, N2582);
nand NAND3 (N2614, N2612, N2290, N2471);
xor XOR2 (N2615, N2588, N1094);
or OR4 (N2616, N2602, N1291, N2091, N1043);
buf BUF1 (N2617, N2615);
nand NAND2 (N2618, N2605, N1030);
and AND3 (N2619, N2616, N469, N1912);
buf BUF1 (N2620, N2614);
buf BUF1 (N2621, N2617);
buf BUF1 (N2622, N2620);
xor XOR2 (N2623, N2596, N1849);
xor XOR2 (N2624, N2604, N2332);
buf BUF1 (N2625, N2619);
xor XOR2 (N2626, N2611, N938);
nor NOR2 (N2627, N2621, N588);
nand NAND3 (N2628, N2613, N109, N1551);
not NOT1 (N2629, N2627);
or OR4 (N2630, N2629, N2426, N589, N2218);
nor NOR2 (N2631, N2630, N173);
nor NOR3 (N2632, N2624, N329, N2091);
not NOT1 (N2633, N2623);
and AND3 (N2634, N2632, N493, N1465);
or OR2 (N2635, N2610, N392);
not NOT1 (N2636, N2635);
nand NAND3 (N2637, N2606, N1783, N2133);
and AND3 (N2638, N2625, N2031, N1298);
and AND4 (N2639, N2631, N1703, N1329, N177);
and AND3 (N2640, N2628, N266, N2405);
nand NAND4 (N2641, N2637, N921, N1516, N1384);
xor XOR2 (N2642, N2640, N1735);
and AND4 (N2643, N2622, N1175, N2126, N389);
xor XOR2 (N2644, N2643, N110);
nand NAND3 (N2645, N2633, N993, N807);
nand NAND2 (N2646, N2638, N2642);
not NOT1 (N2647, N441);
nor NOR4 (N2648, N2641, N328, N2449, N2404);
or OR3 (N2649, N2644, N927, N403);
buf BUF1 (N2650, N2646);
or OR3 (N2651, N2645, N2213, N850);
not NOT1 (N2652, N2626);
buf BUF1 (N2653, N2634);
buf BUF1 (N2654, N2648);
not NOT1 (N2655, N2654);
or OR4 (N2656, N2618, N2547, N1876, N1324);
nand NAND4 (N2657, N2649, N788, N2216, N926);
and AND3 (N2658, N2652, N643, N92);
buf BUF1 (N2659, N2650);
or OR2 (N2660, N2636, N1532);
nand NAND4 (N2661, N2657, N1778, N1312, N1768);
buf BUF1 (N2662, N2659);
and AND2 (N2663, N2660, N825);
not NOT1 (N2664, N2663);
or OR3 (N2665, N2655, N426, N2566);
or OR3 (N2666, N2662, N2511, N1895);
buf BUF1 (N2667, N2651);
not NOT1 (N2668, N2658);
and AND2 (N2669, N2653, N756);
xor XOR2 (N2670, N2667, N924);
not NOT1 (N2671, N2670);
xor XOR2 (N2672, N2661, N271);
nor NOR2 (N2673, N2669, N2020);
nand NAND2 (N2674, N2665, N970);
and AND4 (N2675, N2674, N740, N2277, N2660);
and AND2 (N2676, N2668, N2413);
xor XOR2 (N2677, N2639, N2197);
and AND2 (N2678, N2666, N260);
and AND3 (N2679, N2647, N917, N957);
nor NOR2 (N2680, N2664, N893);
xor XOR2 (N2681, N2676, N2635);
and AND2 (N2682, N2677, N1511);
or OR2 (N2683, N2680, N13);
nand NAND3 (N2684, N2673, N1203, N1937);
nand NAND4 (N2685, N2682, N1787, N930, N92);
xor XOR2 (N2686, N2675, N628);
and AND4 (N2687, N2678, N2674, N234, N2648);
and AND4 (N2688, N2656, N2146, N1850, N374);
xor XOR2 (N2689, N2687, N67);
or OR2 (N2690, N2688, N1644);
and AND3 (N2691, N2689, N388, N1432);
buf BUF1 (N2692, N2681);
nand NAND3 (N2693, N2692, N1550, N741);
or OR4 (N2694, N2684, N1732, N1008, N2658);
xor XOR2 (N2695, N2691, N704);
and AND4 (N2696, N2683, N746, N1674, N2464);
nand NAND2 (N2697, N2695, N2502);
xor XOR2 (N2698, N2693, N1721);
and AND4 (N2699, N2686, N1786, N2512, N230);
and AND4 (N2700, N2698, N1275, N1752, N1964);
nor NOR4 (N2701, N2694, N2306, N1058, N2487);
buf BUF1 (N2702, N2679);
not NOT1 (N2703, N2696);
nor NOR2 (N2704, N2690, N1640);
not NOT1 (N2705, N2700);
buf BUF1 (N2706, N2703);
or OR3 (N2707, N2702, N599, N530);
not NOT1 (N2708, N2701);
or OR3 (N2709, N2699, N700, N886);
not NOT1 (N2710, N2707);
not NOT1 (N2711, N2706);
buf BUF1 (N2712, N2711);
nor NOR4 (N2713, N2697, N940, N540, N794);
nor NOR2 (N2714, N2704, N2004);
nor NOR2 (N2715, N2672, N880);
nand NAND4 (N2716, N2685, N2407, N774, N2042);
not NOT1 (N2717, N2713);
nand NAND3 (N2718, N2709, N1318, N2182);
buf BUF1 (N2719, N2714);
nor NOR3 (N2720, N2719, N256, N834);
and AND4 (N2721, N2716, N302, N1104, N1108);
xor XOR2 (N2722, N2718, N1816);
nand NAND3 (N2723, N2722, N1011, N598);
not NOT1 (N2724, N2723);
buf BUF1 (N2725, N2671);
or OR4 (N2726, N2720, N2595, N660, N345);
or OR3 (N2727, N2726, N89, N782);
buf BUF1 (N2728, N2721);
or OR4 (N2729, N2727, N2093, N142, N526);
or OR4 (N2730, N2715, N1689, N2456, N2216);
or OR4 (N2731, N2724, N388, N1726, N2262);
or OR2 (N2732, N2710, N937);
nor NOR3 (N2733, N2732, N1143, N1368);
xor XOR2 (N2734, N2705, N2569);
and AND4 (N2735, N2731, N2193, N1439, N853);
nand NAND3 (N2736, N2725, N876, N1537);
not NOT1 (N2737, N2733);
and AND4 (N2738, N2734, N961, N1947, N1752);
nand NAND4 (N2739, N2738, N1671, N2592, N2309);
buf BUF1 (N2740, N2730);
and AND4 (N2741, N2712, N2041, N638, N1737);
or OR2 (N2742, N2717, N1888);
buf BUF1 (N2743, N2742);
and AND4 (N2744, N2740, N927, N690, N1841);
buf BUF1 (N2745, N2735);
and AND3 (N2746, N2744, N369, N265);
xor XOR2 (N2747, N2729, N1654);
not NOT1 (N2748, N2743);
or OR2 (N2749, N2746, N251);
xor XOR2 (N2750, N2741, N1350);
nor NOR3 (N2751, N2728, N822, N2282);
nor NOR3 (N2752, N2708, N2016, N1014);
nor NOR3 (N2753, N2749, N1923, N2482);
and AND2 (N2754, N2739, N26);
or OR2 (N2755, N2752, N2592);
not NOT1 (N2756, N2737);
and AND3 (N2757, N2756, N2744, N2525);
xor XOR2 (N2758, N2736, N68);
xor XOR2 (N2759, N2748, N1901);
or OR3 (N2760, N2751, N153, N1870);
buf BUF1 (N2761, N2757);
nand NAND3 (N2762, N2750, N108, N689);
and AND4 (N2763, N2755, N2367, N2735, N2140);
nand NAND2 (N2764, N2762, N274);
or OR2 (N2765, N2758, N23);
or OR4 (N2766, N2759, N212, N1909, N93);
nand NAND3 (N2767, N2747, N1027, N2268);
buf BUF1 (N2768, N2753);
buf BUF1 (N2769, N2763);
buf BUF1 (N2770, N2765);
nor NOR2 (N2771, N2760, N865);
nand NAND4 (N2772, N2761, N1554, N1048, N1964);
or OR3 (N2773, N2767, N2544, N2735);
and AND3 (N2774, N2772, N451, N943);
nand NAND3 (N2775, N2745, N1216, N260);
and AND3 (N2776, N2770, N220, N2496);
nand NAND2 (N2777, N2776, N415);
buf BUF1 (N2778, N2775);
and AND3 (N2779, N2766, N2665, N2468);
and AND4 (N2780, N2774, N1050, N2086, N2249);
and AND2 (N2781, N2778, N701);
nor NOR2 (N2782, N2773, N2641);
nor NOR2 (N2783, N2754, N587);
buf BUF1 (N2784, N2777);
buf BUF1 (N2785, N2781);
nor NOR4 (N2786, N2784, N1225, N1390, N1198);
nor NOR3 (N2787, N2785, N848, N24);
or OR2 (N2788, N2786, N392);
xor XOR2 (N2789, N2764, N1221);
buf BUF1 (N2790, N2788);
xor XOR2 (N2791, N2771, N494);
not NOT1 (N2792, N2779);
nor NOR4 (N2793, N2787, N250, N1243, N867);
nand NAND2 (N2794, N2780, N1619);
nor NOR4 (N2795, N2791, N744, N668, N95);
nor NOR4 (N2796, N2790, N2442, N1806, N2339);
buf BUF1 (N2797, N2789);
or OR3 (N2798, N2768, N612, N566);
nand NAND2 (N2799, N2793, N2379);
buf BUF1 (N2800, N2797);
nand NAND2 (N2801, N2794, N1855);
nor NOR4 (N2802, N2798, N2604, N1484, N160);
not NOT1 (N2803, N2769);
xor XOR2 (N2804, N2803, N600);
or OR3 (N2805, N2783, N568, N1185);
buf BUF1 (N2806, N2795);
nor NOR4 (N2807, N2792, N2447, N311, N2545);
buf BUF1 (N2808, N2806);
not NOT1 (N2809, N2805);
nor NOR4 (N2810, N2800, N1161, N647, N508);
and AND4 (N2811, N2810, N1458, N866, N1201);
or OR3 (N2812, N2807, N2216, N253);
buf BUF1 (N2813, N2799);
nand NAND4 (N2814, N2801, N956, N815, N1034);
buf BUF1 (N2815, N2813);
xor XOR2 (N2816, N2811, N44);
and AND2 (N2817, N2782, N67);
or OR3 (N2818, N2817, N1949, N834);
nor NOR4 (N2819, N2818, N2359, N2198, N1531);
nor NOR3 (N2820, N2812, N190, N794);
xor XOR2 (N2821, N2820, N2344);
buf BUF1 (N2822, N2814);
nand NAND3 (N2823, N2816, N2089, N757);
and AND3 (N2824, N2815, N2816, N1193);
nand NAND3 (N2825, N2809, N2442, N1416);
and AND2 (N2826, N2822, N433);
and AND2 (N2827, N2802, N116);
not NOT1 (N2828, N2827);
nor NOR3 (N2829, N2828, N2471, N758);
xor XOR2 (N2830, N2808, N1305);
and AND4 (N2831, N2819, N2426, N311, N2657);
and AND3 (N2832, N2796, N2237, N558);
nor NOR2 (N2833, N2823, N2373);
not NOT1 (N2834, N2821);
xor XOR2 (N2835, N2804, N1401);
nor NOR4 (N2836, N2829, N486, N405, N755);
buf BUF1 (N2837, N2824);
and AND3 (N2838, N2834, N1652, N503);
xor XOR2 (N2839, N2836, N1957);
nor NOR3 (N2840, N2830, N1421, N2677);
not NOT1 (N2841, N2835);
buf BUF1 (N2842, N2832);
not NOT1 (N2843, N2840);
nand NAND4 (N2844, N2831, N1282, N867, N1601);
nor NOR2 (N2845, N2842, N2275);
xor XOR2 (N2846, N2826, N868);
nor NOR2 (N2847, N2846, N2804);
not NOT1 (N2848, N2833);
nand NAND2 (N2849, N2847, N157);
buf BUF1 (N2850, N2839);
or OR4 (N2851, N2843, N2143, N1039, N2803);
not NOT1 (N2852, N2838);
and AND3 (N2853, N2851, N2542, N2390);
nor NOR4 (N2854, N2841, N1464, N1101, N925);
nor NOR2 (N2855, N2850, N1234);
buf BUF1 (N2856, N2853);
xor XOR2 (N2857, N2849, N2568);
nor NOR4 (N2858, N2848, N1858, N536, N2247);
nand NAND4 (N2859, N2857, N80, N1371, N2466);
or OR3 (N2860, N2844, N2152, N16);
and AND2 (N2861, N2860, N2182);
xor XOR2 (N2862, N2856, N2437);
and AND4 (N2863, N2852, N933, N2834, N1197);
not NOT1 (N2864, N2855);
not NOT1 (N2865, N2854);
xor XOR2 (N2866, N2861, N1647);
or OR2 (N2867, N2859, N862);
or OR2 (N2868, N2865, N2756);
and AND2 (N2869, N2867, N1943);
buf BUF1 (N2870, N2825);
nand NAND4 (N2871, N2866, N60, N1832, N262);
and AND4 (N2872, N2869, N1861, N2603, N1050);
nor NOR2 (N2873, N2868, N1635);
xor XOR2 (N2874, N2862, N414);
nor NOR4 (N2875, N2871, N937, N2542, N2436);
xor XOR2 (N2876, N2858, N1094);
or OR3 (N2877, N2874, N540, N397);
nor NOR2 (N2878, N2875, N1807);
not NOT1 (N2879, N2878);
buf BUF1 (N2880, N2877);
and AND2 (N2881, N2873, N112);
and AND3 (N2882, N2876, N371, N115);
xor XOR2 (N2883, N2845, N1821);
xor XOR2 (N2884, N2883, N1735);
nor NOR4 (N2885, N2879, N2780, N1436, N1392);
nor NOR2 (N2886, N2837, N79);
xor XOR2 (N2887, N2886, N1787);
buf BUF1 (N2888, N2885);
nor NOR2 (N2889, N2870, N1225);
buf BUF1 (N2890, N2864);
nand NAND4 (N2891, N2889, N1585, N1446, N1625);
not NOT1 (N2892, N2863);
xor XOR2 (N2893, N2890, N1910);
buf BUF1 (N2894, N2891);
and AND2 (N2895, N2884, N1838);
not NOT1 (N2896, N2888);
nand NAND4 (N2897, N2892, N1372, N1349, N370);
nor NOR4 (N2898, N2895, N2339, N588, N294);
not NOT1 (N2899, N2894);
and AND4 (N2900, N2882, N627, N1413, N597);
or OR4 (N2901, N2887, N1859, N523, N2153);
buf BUF1 (N2902, N2898);
and AND4 (N2903, N2881, N1326, N531, N83);
and AND2 (N2904, N2896, N301);
xor XOR2 (N2905, N2893, N1029);
or OR2 (N2906, N2872, N270);
nand NAND2 (N2907, N2880, N1395);
or OR4 (N2908, N2907, N1734, N2322, N1590);
nor NOR4 (N2909, N2900, N252, N693, N804);
nand NAND3 (N2910, N2902, N1502, N1124);
buf BUF1 (N2911, N2905);
nor NOR2 (N2912, N2897, N2661);
buf BUF1 (N2913, N2908);
not NOT1 (N2914, N2909);
or OR2 (N2915, N2914, N554);
not NOT1 (N2916, N2910);
nor NOR3 (N2917, N2915, N991, N134);
buf BUF1 (N2918, N2916);
nor NOR4 (N2919, N2906, N2459, N1083, N155);
nand NAND4 (N2920, N2901, N2019, N2889, N1670);
xor XOR2 (N2921, N2920, N2824);
xor XOR2 (N2922, N2904, N737);
nand NAND4 (N2923, N2912, N1497, N639, N2644);
or OR4 (N2924, N2919, N1571, N2638, N300);
nand NAND4 (N2925, N2922, N1783, N2409, N2475);
or OR2 (N2926, N2911, N1392);
not NOT1 (N2927, N2925);
buf BUF1 (N2928, N2917);
buf BUF1 (N2929, N2899);
buf BUF1 (N2930, N2927);
not NOT1 (N2931, N2930);
buf BUF1 (N2932, N2926);
nor NOR3 (N2933, N2913, N1597, N2649);
or OR3 (N2934, N2921, N1448, N1001);
or OR3 (N2935, N2918, N379, N2745);
nand NAND3 (N2936, N2903, N2813, N1502);
and AND4 (N2937, N2936, N2050, N762, N646);
buf BUF1 (N2938, N2933);
buf BUF1 (N2939, N2937);
xor XOR2 (N2940, N2932, N2524);
or OR3 (N2941, N2940, N140, N2496);
nand NAND4 (N2942, N2939, N2357, N992, N1981);
nand NAND2 (N2943, N2938, N1766);
nand NAND3 (N2944, N2935, N1139, N2265);
not NOT1 (N2945, N2942);
buf BUF1 (N2946, N2945);
or OR4 (N2947, N2934, N521, N1584, N113);
not NOT1 (N2948, N2928);
nand NAND2 (N2949, N2948, N2353);
and AND3 (N2950, N2943, N880, N2623);
nor NOR2 (N2951, N2944, N558);
or OR4 (N2952, N2923, N987, N736, N1156);
or OR2 (N2953, N2947, N2479);
not NOT1 (N2954, N2941);
or OR3 (N2955, N2950, N1646, N2261);
not NOT1 (N2956, N2952);
and AND3 (N2957, N2924, N923, N2644);
buf BUF1 (N2958, N2953);
nor NOR2 (N2959, N2955, N1506);
xor XOR2 (N2960, N2957, N1018);
or OR4 (N2961, N2959, N2454, N774, N2459);
and AND4 (N2962, N2946, N634, N1085, N324);
nor NOR4 (N2963, N2929, N1263, N1770, N2325);
not NOT1 (N2964, N2949);
nor NOR3 (N2965, N2961, N337, N1724);
and AND3 (N2966, N2951, N2848, N2192);
xor XOR2 (N2967, N2966, N1578);
nand NAND3 (N2968, N2964, N2888, N2090);
buf BUF1 (N2969, N2956);
buf BUF1 (N2970, N2960);
buf BUF1 (N2971, N2968);
xor XOR2 (N2972, N2931, N193);
and AND3 (N2973, N2970, N735, N1143);
and AND4 (N2974, N2958, N1322, N939, N1108);
nand NAND4 (N2975, N2974, N1826, N1772, N1168);
xor XOR2 (N2976, N2965, N2436);
or OR2 (N2977, N2971, N439);
xor XOR2 (N2978, N2969, N877);
nor NOR3 (N2979, N2972, N108, N1063);
and AND4 (N2980, N2967, N1485, N92, N1735);
or OR2 (N2981, N2962, N2107);
nand NAND2 (N2982, N2973, N1955);
nand NAND4 (N2983, N2978, N1677, N2194, N1584);
nor NOR2 (N2984, N2983, N2276);
nand NAND4 (N2985, N2982, N2367, N952, N917);
xor XOR2 (N2986, N2985, N2683);
nor NOR2 (N2987, N2984, N1237);
buf BUF1 (N2988, N2963);
nor NOR2 (N2989, N2976, N1573);
buf BUF1 (N2990, N2987);
and AND2 (N2991, N2980, N2798);
nand NAND3 (N2992, N2954, N624, N1823);
buf BUF1 (N2993, N2975);
nor NOR4 (N2994, N2981, N1007, N2190, N1517);
xor XOR2 (N2995, N2986, N799);
nand NAND2 (N2996, N2977, N1490);
not NOT1 (N2997, N2994);
not NOT1 (N2998, N2991);
nand NAND4 (N2999, N2998, N1941, N1985, N1095);
buf BUF1 (N3000, N2990);
not NOT1 (N3001, N3000);
and AND4 (N3002, N2993, N2418, N241, N76);
or OR2 (N3003, N2988, N1541);
not NOT1 (N3004, N2979);
nor NOR4 (N3005, N2996, N2955, N240, N2524);
and AND4 (N3006, N2989, N2765, N2892, N1120);
or OR4 (N3007, N2997, N708, N557, N910);
xor XOR2 (N3008, N3004, N2944);
nand NAND4 (N3009, N3006, N638, N920, N363);
buf BUF1 (N3010, N3008);
buf BUF1 (N3011, N3007);
or OR3 (N3012, N2992, N493, N2370);
or OR4 (N3013, N2999, N2058, N2838, N2477);
nor NOR3 (N3014, N3003, N1865, N2978);
xor XOR2 (N3015, N3014, N710);
xor XOR2 (N3016, N3011, N2848);
xor XOR2 (N3017, N3016, N2919);
not NOT1 (N3018, N3001);
buf BUF1 (N3019, N3012);
or OR4 (N3020, N3009, N2741, N1909, N2023);
not NOT1 (N3021, N3018);
nor NOR4 (N3022, N3017, N165, N347, N2891);
nand NAND4 (N3023, N3020, N1548, N557, N1807);
xor XOR2 (N3024, N3021, N12);
not NOT1 (N3025, N3024);
nor NOR3 (N3026, N3023, N2782, N1002);
or OR2 (N3027, N3026, N1181);
nor NOR4 (N3028, N3002, N153, N801, N2285);
buf BUF1 (N3029, N3022);
not NOT1 (N3030, N3015);
or OR2 (N3031, N3005, N3018);
or OR2 (N3032, N3028, N892);
and AND3 (N3033, N3031, N1341, N740);
xor XOR2 (N3034, N3029, N1250);
and AND3 (N3035, N3019, N1552, N1467);
xor XOR2 (N3036, N3034, N1259);
buf BUF1 (N3037, N3032);
nor NOR4 (N3038, N3036, N1743, N1336, N292);
or OR4 (N3039, N3013, N1614, N1845, N172);
and AND3 (N3040, N3010, N560, N1257);
nor NOR2 (N3041, N3037, N1842);
and AND2 (N3042, N3030, N2632);
buf BUF1 (N3043, N3039);
and AND2 (N3044, N3027, N1030);
xor XOR2 (N3045, N2995, N1175);
not NOT1 (N3046, N3044);
or OR3 (N3047, N3042, N3, N1804);
buf BUF1 (N3048, N3040);
not NOT1 (N3049, N3033);
nor NOR2 (N3050, N3035, N198);
or OR2 (N3051, N3050, N2526);
xor XOR2 (N3052, N3047, N2229);
and AND2 (N3053, N3043, N1873);
buf BUF1 (N3054, N3051);
nor NOR2 (N3055, N3048, N1228);
or OR2 (N3056, N3049, N245);
not NOT1 (N3057, N3056);
or OR4 (N3058, N3045, N379, N1133, N156);
buf BUF1 (N3059, N3055);
nor NOR3 (N3060, N3046, N2977, N402);
nand NAND2 (N3061, N3053, N1329);
xor XOR2 (N3062, N3057, N1355);
and AND4 (N3063, N3025, N176, N2178, N717);
and AND2 (N3064, N3054, N149);
not NOT1 (N3065, N3063);
nand NAND3 (N3066, N3058, N811, N2852);
not NOT1 (N3067, N3038);
not NOT1 (N3068, N3065);
buf BUF1 (N3069, N3066);
and AND3 (N3070, N3052, N1251, N1144);
buf BUF1 (N3071, N3068);
or OR4 (N3072, N3062, N2237, N732, N95);
nor NOR4 (N3073, N3041, N2187, N2624, N561);
nand NAND2 (N3074, N3071, N2991);
or OR2 (N3075, N3060, N2595);
not NOT1 (N3076, N3075);
buf BUF1 (N3077, N3076);
and AND4 (N3078, N3074, N2595, N1602, N1833);
xor XOR2 (N3079, N3078, N3055);
buf BUF1 (N3080, N3064);
buf BUF1 (N3081, N3069);
buf BUF1 (N3082, N3079);
not NOT1 (N3083, N3061);
and AND4 (N3084, N3080, N1522, N2304, N186);
or OR3 (N3085, N3059, N2171, N1554);
nand NAND2 (N3086, N3067, N1991);
nand NAND2 (N3087, N3077, N2244);
xor XOR2 (N3088, N3086, N2382);
nand NAND3 (N3089, N3088, N2522, N2512);
or OR3 (N3090, N3072, N964, N2662);
xor XOR2 (N3091, N3090, N2368);
not NOT1 (N3092, N3091);
xor XOR2 (N3093, N3073, N1180);
or OR2 (N3094, N3089, N686);
nor NOR4 (N3095, N3085, N1989, N1766, N1723);
or OR2 (N3096, N3081, N979);
or OR4 (N3097, N3096, N1745, N2365, N1425);
xor XOR2 (N3098, N3070, N282);
nand NAND3 (N3099, N3083, N1986, N2573);
and AND2 (N3100, N3094, N2267);
and AND3 (N3101, N3087, N848, N130);
not NOT1 (N3102, N3092);
buf BUF1 (N3103, N3093);
xor XOR2 (N3104, N3095, N1565);
nor NOR2 (N3105, N3103, N1746);
and AND4 (N3106, N3102, N570, N438, N2484);
xor XOR2 (N3107, N3101, N117);
nand NAND4 (N3108, N3099, N1768, N518, N2031);
buf BUF1 (N3109, N3108);
or OR2 (N3110, N3106, N2576);
and AND4 (N3111, N3104, N495, N1917, N1765);
nor NOR4 (N3112, N3111, N2523, N271, N2469);
or OR3 (N3113, N3107, N576, N2388);
buf BUF1 (N3114, N3109);
or OR4 (N3115, N3112, N452, N3083, N1931);
buf BUF1 (N3116, N3105);
buf BUF1 (N3117, N3082);
nand NAND4 (N3118, N3098, N992, N2485, N218);
nor NOR3 (N3119, N3084, N1989, N2867);
or OR3 (N3120, N3114, N534, N1855);
nand NAND3 (N3121, N3110, N2977, N714);
nor NOR2 (N3122, N3100, N656);
or OR2 (N3123, N3122, N1663);
nor NOR4 (N3124, N3117, N1, N2472, N3066);
or OR2 (N3125, N3124, N2391);
or OR2 (N3126, N3113, N388);
xor XOR2 (N3127, N3119, N1957);
nand NAND3 (N3128, N3125, N2064, N2435);
not NOT1 (N3129, N3123);
nand NAND2 (N3130, N3128, N690);
xor XOR2 (N3131, N3120, N2594);
nand NAND4 (N3132, N3097, N2790, N1865, N216);
nor NOR3 (N3133, N3127, N2997, N1020);
and AND4 (N3134, N3118, N565, N103, N1076);
buf BUF1 (N3135, N3134);
nor NOR2 (N3136, N3131, N2283);
xor XOR2 (N3137, N3136, N3066);
not NOT1 (N3138, N3129);
buf BUF1 (N3139, N3135);
or OR4 (N3140, N3126, N2239, N3090, N175);
or OR4 (N3141, N3132, N1993, N2270, N1964);
nor NOR2 (N3142, N3137, N1269);
nand NAND3 (N3143, N3141, N1297, N1060);
buf BUF1 (N3144, N3116);
xor XOR2 (N3145, N3121, N340);
or OR2 (N3146, N3139, N965);
nor NOR3 (N3147, N3138, N262, N2190);
nor NOR4 (N3148, N3145, N1589, N304, N3012);
nand NAND2 (N3149, N3148, N2815);
and AND4 (N3150, N3115, N1833, N2782, N1859);
nand NAND3 (N3151, N3146, N465, N1621);
buf BUF1 (N3152, N3149);
nor NOR2 (N3153, N3130, N727);
nor NOR4 (N3154, N3152, N597, N1725, N950);
nor NOR4 (N3155, N3153, N1944, N2325, N2240);
nor NOR3 (N3156, N3144, N339, N933);
not NOT1 (N3157, N3143);
nor NOR4 (N3158, N3151, N1840, N1529, N1645);
xor XOR2 (N3159, N3158, N1122);
nor NOR3 (N3160, N3150, N2407, N146);
nand NAND2 (N3161, N3147, N1250);
xor XOR2 (N3162, N3160, N215);
xor XOR2 (N3163, N3157, N1735);
and AND3 (N3164, N3163, N191, N2981);
buf BUF1 (N3165, N3155);
buf BUF1 (N3166, N3165);
or OR2 (N3167, N3156, N450);
nand NAND4 (N3168, N3142, N2232, N1930, N904);
buf BUF1 (N3169, N3159);
and AND4 (N3170, N3166, N2320, N1637, N1097);
and AND2 (N3171, N3168, N3129);
and AND4 (N3172, N3171, N242, N1301, N819);
buf BUF1 (N3173, N3170);
not NOT1 (N3174, N3169);
nand NAND3 (N3175, N3162, N1756, N1338);
nand NAND4 (N3176, N3172, N2604, N953, N2888);
or OR4 (N3177, N3175, N2828, N664, N2072);
xor XOR2 (N3178, N3176, N1164);
nand NAND4 (N3179, N3164, N2080, N1647, N348);
xor XOR2 (N3180, N3177, N2162);
and AND3 (N3181, N3178, N3168, N3139);
not NOT1 (N3182, N3133);
or OR3 (N3183, N3154, N2976, N1273);
nand NAND2 (N3184, N3140, N409);
and AND4 (N3185, N3184, N2369, N2375, N990);
nor NOR4 (N3186, N3182, N2826, N2803, N1939);
or OR2 (N3187, N3173, N2446);
xor XOR2 (N3188, N3181, N2929);
nor NOR2 (N3189, N3180, N744);
not NOT1 (N3190, N3167);
nor NOR3 (N3191, N3161, N1223, N3093);
nand NAND3 (N3192, N3188, N2083, N1235);
and AND3 (N3193, N3190, N2761, N156);
xor XOR2 (N3194, N3193, N1249);
nand NAND3 (N3195, N3191, N2326, N2710);
not NOT1 (N3196, N3194);
nor NOR3 (N3197, N3195, N1434, N2456);
and AND2 (N3198, N3192, N1089);
xor XOR2 (N3199, N3186, N1173);
not NOT1 (N3200, N3199);
and AND3 (N3201, N3174, N3008, N1924);
not NOT1 (N3202, N3183);
or OR4 (N3203, N3198, N2206, N584, N1936);
buf BUF1 (N3204, N3189);
not NOT1 (N3205, N3197);
nand NAND4 (N3206, N3179, N2274, N2639, N2831);
xor XOR2 (N3207, N3205, N1728);
buf BUF1 (N3208, N3204);
and AND2 (N3209, N3203, N1302);
buf BUF1 (N3210, N3201);
nand NAND3 (N3211, N3200, N2437, N261);
not NOT1 (N3212, N3185);
nor NOR3 (N3213, N3187, N2027, N1219);
and AND4 (N3214, N3212, N737, N2766, N1569);
not NOT1 (N3215, N3211);
not NOT1 (N3216, N3206);
and AND3 (N3217, N3209, N762, N1065);
buf BUF1 (N3218, N3214);
not NOT1 (N3219, N3216);
xor XOR2 (N3220, N3219, N119);
buf BUF1 (N3221, N3213);
and AND2 (N3222, N3202, N2668);
or OR3 (N3223, N3217, N249, N1476);
or OR2 (N3224, N3222, N2543);
xor XOR2 (N3225, N3224, N772);
not NOT1 (N3226, N3220);
not NOT1 (N3227, N3196);
not NOT1 (N3228, N3226);
not NOT1 (N3229, N3221);
not NOT1 (N3230, N3225);
nor NOR2 (N3231, N3207, N1496);
nor NOR4 (N3232, N3208, N2556, N474, N1753);
buf BUF1 (N3233, N3223);
buf BUF1 (N3234, N3227);
nor NOR2 (N3235, N3233, N2099);
not NOT1 (N3236, N3232);
xor XOR2 (N3237, N3210, N2090);
not NOT1 (N3238, N3230);
nor NOR3 (N3239, N3238, N2984, N1442);
buf BUF1 (N3240, N3234);
nor NOR2 (N3241, N3231, N197);
not NOT1 (N3242, N3241);
nor NOR3 (N3243, N3229, N502, N1718);
or OR2 (N3244, N3235, N1190);
or OR3 (N3245, N3243, N1822, N1965);
xor XOR2 (N3246, N3218, N67);
not NOT1 (N3247, N3242);
nor NOR3 (N3248, N3240, N961, N2851);
nand NAND2 (N3249, N3247, N1351);
nand NAND2 (N3250, N3236, N2052);
or OR2 (N3251, N3215, N1607);
nor NOR4 (N3252, N3244, N761, N1395, N2875);
xor XOR2 (N3253, N3249, N2243);
or OR4 (N3254, N3228, N759, N1521, N1404);
and AND3 (N3255, N3248, N1256, N2009);
buf BUF1 (N3256, N3239);
or OR4 (N3257, N3253, N1014, N3031, N245);
not NOT1 (N3258, N3257);
or OR2 (N3259, N3250, N740);
xor XOR2 (N3260, N3258, N971);
xor XOR2 (N3261, N3254, N2173);
nand NAND2 (N3262, N3237, N111);
not NOT1 (N3263, N3255);
buf BUF1 (N3264, N3245);
xor XOR2 (N3265, N3246, N248);
and AND4 (N3266, N3261, N1011, N2594, N742);
or OR4 (N3267, N3265, N226, N1692, N1023);
buf BUF1 (N3268, N3260);
or OR2 (N3269, N3256, N1469);
or OR2 (N3270, N3269, N3023);
and AND4 (N3271, N3262, N1796, N1927, N3207);
xor XOR2 (N3272, N3259, N828);
buf BUF1 (N3273, N3267);
nand NAND3 (N3274, N3263, N2844, N2407);
buf BUF1 (N3275, N3274);
nand NAND3 (N3276, N3251, N1599, N1749);
nor NOR2 (N3277, N3270, N71);
and AND4 (N3278, N3271, N1917, N574, N560);
xor XOR2 (N3279, N3273, N833);
buf BUF1 (N3280, N3266);
nor NOR4 (N3281, N3280, N2206, N2346, N166);
nor NOR2 (N3282, N3268, N2929);
xor XOR2 (N3283, N3282, N2342);
xor XOR2 (N3284, N3276, N64);
and AND3 (N3285, N3278, N38, N1821);
nand NAND4 (N3286, N3281, N2560, N498, N1067);
and AND4 (N3287, N3277, N1750, N368, N2817);
xor XOR2 (N3288, N3264, N1757);
or OR2 (N3289, N3252, N39);
buf BUF1 (N3290, N3275);
nand NAND4 (N3291, N3289, N3009, N434, N668);
nor NOR2 (N3292, N3284, N1334);
not NOT1 (N3293, N3286);
and AND2 (N3294, N3288, N219);
nand NAND3 (N3295, N3283, N2484, N855);
buf BUF1 (N3296, N3290);
xor XOR2 (N3297, N3272, N2575);
buf BUF1 (N3298, N3279);
xor XOR2 (N3299, N3297, N2203);
and AND4 (N3300, N3294, N1044, N414, N2981);
nand NAND4 (N3301, N3298, N1873, N2994, N758);
not NOT1 (N3302, N3291);
xor XOR2 (N3303, N3300, N505);
not NOT1 (N3304, N3285);
xor XOR2 (N3305, N3292, N2622);
not NOT1 (N3306, N3295);
nand NAND2 (N3307, N3303, N1771);
and AND4 (N3308, N3305, N2491, N2792, N283);
buf BUF1 (N3309, N3293);
not NOT1 (N3310, N3287);
and AND4 (N3311, N3310, N1209, N673, N2399);
and AND3 (N3312, N3304, N1101, N21);
nand NAND4 (N3313, N3312, N1022, N2459, N2788);
not NOT1 (N3314, N3308);
not NOT1 (N3315, N3301);
buf BUF1 (N3316, N3307);
buf BUF1 (N3317, N3299);
and AND2 (N3318, N3317, N1894);
buf BUF1 (N3319, N3311);
and AND2 (N3320, N3315, N1173);
or OR3 (N3321, N3313, N3021, N1787);
and AND3 (N3322, N3302, N1904, N323);
and AND4 (N3323, N3314, N2578, N781, N253);
or OR2 (N3324, N3296, N2475);
not NOT1 (N3325, N3319);
or OR4 (N3326, N3306, N2444, N2419, N1664);
or OR2 (N3327, N3325, N1703);
and AND4 (N3328, N3326, N2684, N1756, N1203);
nor NOR4 (N3329, N3320, N1263, N2242, N523);
buf BUF1 (N3330, N3324);
xor XOR2 (N3331, N3316, N1958);
buf BUF1 (N3332, N3318);
or OR4 (N3333, N3329, N2957, N2473, N2509);
xor XOR2 (N3334, N3330, N1000);
nand NAND4 (N3335, N3334, N1421, N1863, N525);
or OR3 (N3336, N3328, N652, N1334);
not NOT1 (N3337, N3309);
nand NAND4 (N3338, N3335, N2496, N230, N1496);
buf BUF1 (N3339, N3331);
nand NAND4 (N3340, N3333, N1938, N1306, N2862);
nand NAND4 (N3341, N3321, N1923, N531, N1019);
not NOT1 (N3342, N3332);
nor NOR3 (N3343, N3327, N2255, N1388);
nand NAND3 (N3344, N3339, N568, N2223);
not NOT1 (N3345, N3338);
nand NAND2 (N3346, N3344, N2351);
and AND4 (N3347, N3346, N60, N1954, N1541);
not NOT1 (N3348, N3347);
nor NOR2 (N3349, N3323, N247);
or OR2 (N3350, N3345, N1012);
xor XOR2 (N3351, N3337, N1823);
nand NAND3 (N3352, N3349, N133, N855);
nand NAND4 (N3353, N3343, N2783, N2762, N2353);
and AND4 (N3354, N3342, N459, N1766, N751);
nor NOR4 (N3355, N3352, N3234, N66, N927);
buf BUF1 (N3356, N3341);
xor XOR2 (N3357, N3322, N2864);
or OR3 (N3358, N3354, N2645, N42);
nor NOR2 (N3359, N3355, N668);
or OR3 (N3360, N3356, N1283, N2661);
or OR2 (N3361, N3350, N3249);
buf BUF1 (N3362, N3348);
nand NAND4 (N3363, N3351, N184, N1587, N1872);
and AND2 (N3364, N3336, N1044);
not NOT1 (N3365, N3357);
and AND4 (N3366, N3353, N594, N1797, N98);
nor NOR3 (N3367, N3363, N120, N3211);
nand NAND2 (N3368, N3358, N3181);
buf BUF1 (N3369, N3368);
xor XOR2 (N3370, N3365, N1121);
and AND2 (N3371, N3340, N1887);
and AND3 (N3372, N3361, N3280, N2594);
or OR4 (N3373, N3367, N872, N2390, N1312);
and AND4 (N3374, N3373, N3259, N1312, N1196);
or OR2 (N3375, N3366, N416);
xor XOR2 (N3376, N3364, N2223);
nor NOR2 (N3377, N3371, N1718);
or OR3 (N3378, N3362, N1332, N547);
nand NAND3 (N3379, N3370, N798, N422);
not NOT1 (N3380, N3359);
not NOT1 (N3381, N3376);
nand NAND2 (N3382, N3360, N1075);
nor NOR4 (N3383, N3374, N309, N1623, N2643);
nor NOR3 (N3384, N3369, N3070, N1116);
nand NAND4 (N3385, N3375, N3015, N1232, N3361);
xor XOR2 (N3386, N3382, N2419);
or OR3 (N3387, N3377, N2596, N71);
not NOT1 (N3388, N3378);
xor XOR2 (N3389, N3380, N1038);
nand NAND2 (N3390, N3383, N1917);
nand NAND4 (N3391, N3386, N3122, N2931, N1854);
nand NAND2 (N3392, N3390, N365);
or OR4 (N3393, N3384, N1168, N1748, N1983);
xor XOR2 (N3394, N3391, N3150);
or OR3 (N3395, N3372, N2603, N567);
not NOT1 (N3396, N3394);
xor XOR2 (N3397, N3385, N1007);
nor NOR3 (N3398, N3392, N1829, N675);
buf BUF1 (N3399, N3398);
xor XOR2 (N3400, N3396, N2314);
buf BUF1 (N3401, N3397);
xor XOR2 (N3402, N3388, N1276);
buf BUF1 (N3403, N3400);
nor NOR4 (N3404, N3395, N2132, N138, N1602);
xor XOR2 (N3405, N3401, N1157);
nand NAND3 (N3406, N3403, N399, N1291);
nor NOR3 (N3407, N3387, N3009, N537);
nor NOR4 (N3408, N3405, N1198, N432, N1441);
nand NAND2 (N3409, N3404, N2786);
buf BUF1 (N3410, N3389);
nor NOR2 (N3411, N3406, N1804);
not NOT1 (N3412, N3379);
not NOT1 (N3413, N3407);
or OR4 (N3414, N3402, N2629, N21, N1516);
and AND4 (N3415, N3413, N1982, N1403, N1532);
not NOT1 (N3416, N3411);
buf BUF1 (N3417, N3415);
or OR2 (N3418, N3414, N1161);
and AND3 (N3419, N3412, N2306, N706);
xor XOR2 (N3420, N3417, N1359);
nand NAND4 (N3421, N3393, N3154, N786, N2176);
and AND2 (N3422, N3420, N3066);
buf BUF1 (N3423, N3408);
or OR4 (N3424, N3399, N1139, N2197, N2846);
xor XOR2 (N3425, N3410, N2065);
buf BUF1 (N3426, N3419);
nor NOR2 (N3427, N3381, N814);
not NOT1 (N3428, N3418);
not NOT1 (N3429, N3422);
or OR2 (N3430, N3429, N424);
nor NOR4 (N3431, N3424, N1745, N1606, N757);
xor XOR2 (N3432, N3421, N2950);
nor NOR2 (N3433, N3427, N2100);
not NOT1 (N3434, N3428);
or OR4 (N3435, N3423, N1618, N2940, N2440);
and AND2 (N3436, N3434, N1284);
xor XOR2 (N3437, N3436, N1991);
and AND2 (N3438, N3435, N2816);
not NOT1 (N3439, N3409);
xor XOR2 (N3440, N3437, N2159);
not NOT1 (N3441, N3440);
or OR2 (N3442, N3430, N1350);
buf BUF1 (N3443, N3426);
nor NOR3 (N3444, N3433, N748, N2283);
xor XOR2 (N3445, N3439, N1139);
buf BUF1 (N3446, N3442);
nand NAND4 (N3447, N3431, N1973, N2659, N3062);
buf BUF1 (N3448, N3447);
nor NOR2 (N3449, N3416, N2224);
buf BUF1 (N3450, N3449);
or OR4 (N3451, N3432, N2327, N634, N1884);
nor NOR3 (N3452, N3443, N1311, N1952);
xor XOR2 (N3453, N3452, N477);
buf BUF1 (N3454, N3450);
and AND3 (N3455, N3446, N2732, N1700);
and AND4 (N3456, N3451, N21, N3046, N2050);
nand NAND2 (N3457, N3453, N250);
xor XOR2 (N3458, N3457, N1992);
xor XOR2 (N3459, N3444, N2165);
not NOT1 (N3460, N3455);
nor NOR4 (N3461, N3448, N1671, N2655, N2553);
not NOT1 (N3462, N3445);
and AND4 (N3463, N3425, N2270, N1521, N1421);
not NOT1 (N3464, N3462);
or OR3 (N3465, N3464, N1116, N112);
nor NOR3 (N3466, N3456, N2378, N2452);
or OR3 (N3467, N3441, N2124, N786);
buf BUF1 (N3468, N3465);
buf BUF1 (N3469, N3461);
not NOT1 (N3470, N3463);
not NOT1 (N3471, N3438);
not NOT1 (N3472, N3460);
not NOT1 (N3473, N3467);
not NOT1 (N3474, N3459);
or OR4 (N3475, N3469, N3152, N1273, N1620);
and AND3 (N3476, N3466, N1194, N996);
nand NAND2 (N3477, N3475, N977);
not NOT1 (N3478, N3468);
and AND3 (N3479, N3474, N2409, N457);
not NOT1 (N3480, N3472);
not NOT1 (N3481, N3454);
nand NAND4 (N3482, N3477, N2015, N700, N2814);
and AND2 (N3483, N3481, N3014);
and AND4 (N3484, N3458, N227, N2624, N1554);
not NOT1 (N3485, N3479);
or OR2 (N3486, N3483, N2511);
nor NOR3 (N3487, N3480, N123, N613);
xor XOR2 (N3488, N3482, N60);
nor NOR3 (N3489, N3476, N1600, N2350);
not NOT1 (N3490, N3471);
nor NOR2 (N3491, N3485, N889);
or OR2 (N3492, N3487, N2730);
xor XOR2 (N3493, N3489, N1323);
buf BUF1 (N3494, N3488);
buf BUF1 (N3495, N3484);
nor NOR3 (N3496, N3478, N2549, N2313);
or OR2 (N3497, N3486, N1761);
xor XOR2 (N3498, N3473, N1371);
nand NAND3 (N3499, N3492, N2540, N1534);
xor XOR2 (N3500, N3470, N1294);
xor XOR2 (N3501, N3490, N709);
buf BUF1 (N3502, N3496);
nand NAND2 (N3503, N3497, N3350);
not NOT1 (N3504, N3502);
and AND4 (N3505, N3499, N1937, N2320, N2423);
or OR2 (N3506, N3500, N2416);
and AND4 (N3507, N3504, N989, N2019, N407);
nand NAND2 (N3508, N3493, N2027);
and AND4 (N3509, N3491, N637, N141, N1853);
not NOT1 (N3510, N3494);
and AND3 (N3511, N3508, N1844, N3058);
xor XOR2 (N3512, N3510, N1133);
nand NAND2 (N3513, N3507, N2961);
nand NAND4 (N3514, N3509, N1839, N1887, N950);
xor XOR2 (N3515, N3511, N2107);
buf BUF1 (N3516, N3515);
or OR4 (N3517, N3501, N646, N184, N3073);
not NOT1 (N3518, N3516);
nand NAND2 (N3519, N3506, N661);
xor XOR2 (N3520, N3519, N373);
nand NAND4 (N3521, N3503, N3264, N1070, N1159);
xor XOR2 (N3522, N3520, N2255);
nand NAND3 (N3523, N3522, N1396, N105);
nand NAND3 (N3524, N3513, N493, N1101);
nor NOR4 (N3525, N3523, N1970, N1012, N1056);
and AND2 (N3526, N3514, N2681);
xor XOR2 (N3527, N3521, N2649);
or OR2 (N3528, N3526, N1246);
not NOT1 (N3529, N3495);
nand NAND2 (N3530, N3512, N71);
nand NAND3 (N3531, N3498, N2278, N3185);
nand NAND2 (N3532, N3505, N921);
xor XOR2 (N3533, N3524, N794);
nor NOR3 (N3534, N3518, N1567, N867);
nand NAND3 (N3535, N3532, N2628, N462);
xor XOR2 (N3536, N3534, N2253);
xor XOR2 (N3537, N3536, N515);
xor XOR2 (N3538, N3517, N29);
xor XOR2 (N3539, N3533, N116);
not NOT1 (N3540, N3539);
and AND3 (N3541, N3537, N1133, N341);
or OR3 (N3542, N3525, N2472, N1093);
nand NAND4 (N3543, N3530, N24, N3511, N3039);
not NOT1 (N3544, N3542);
xor XOR2 (N3545, N3531, N1653);
xor XOR2 (N3546, N3529, N2329);
xor XOR2 (N3547, N3543, N942);
nor NOR3 (N3548, N3528, N2576, N489);
not NOT1 (N3549, N3527);
xor XOR2 (N3550, N3546, N2543);
nand NAND4 (N3551, N3545, N2290, N1371, N740);
buf BUF1 (N3552, N3538);
buf BUF1 (N3553, N3552);
buf BUF1 (N3554, N3540);
xor XOR2 (N3555, N3550, N357);
buf BUF1 (N3556, N3547);
or OR4 (N3557, N3544, N261, N1248, N2270);
and AND4 (N3558, N3557, N6, N1903, N2028);
nand NAND3 (N3559, N3551, N161, N493);
and AND2 (N3560, N3548, N2291);
xor XOR2 (N3561, N3555, N30);
nor NOR2 (N3562, N3535, N140);
not NOT1 (N3563, N3562);
buf BUF1 (N3564, N3554);
and AND3 (N3565, N3541, N3562, N1546);
not NOT1 (N3566, N3553);
buf BUF1 (N3567, N3558);
and AND2 (N3568, N3564, N990);
nand NAND3 (N3569, N3559, N96, N2287);
nand NAND4 (N3570, N3567, N614, N3253, N1384);
or OR4 (N3571, N3568, N3330, N800, N2645);
xor XOR2 (N3572, N3560, N1615);
not NOT1 (N3573, N3569);
and AND4 (N3574, N3561, N978, N896, N2099);
and AND3 (N3575, N3571, N677, N2150);
xor XOR2 (N3576, N3570, N812);
not NOT1 (N3577, N3563);
nand NAND3 (N3578, N3576, N3067, N87);
buf BUF1 (N3579, N3575);
nor NOR2 (N3580, N3565, N3260);
or OR2 (N3581, N3549, N2605);
and AND4 (N3582, N3578, N2170, N822, N1381);
nor NOR2 (N3583, N3582, N1075);
xor XOR2 (N3584, N3579, N2905);
nor NOR3 (N3585, N3580, N12, N3060);
xor XOR2 (N3586, N3566, N1639);
or OR3 (N3587, N3584, N3014, N1762);
nor NOR2 (N3588, N3587, N1424);
buf BUF1 (N3589, N3577);
and AND3 (N3590, N3556, N2243, N2257);
nor NOR4 (N3591, N3574, N1099, N876, N2591);
xor XOR2 (N3592, N3591, N1635);
nand NAND3 (N3593, N3581, N1323, N110);
nor NOR2 (N3594, N3592, N1911);
and AND3 (N3595, N3594, N1931, N628);
not NOT1 (N3596, N3590);
nand NAND4 (N3597, N3588, N3433, N3012, N2241);
or OR3 (N3598, N3596, N669, N1427);
xor XOR2 (N3599, N3583, N2369);
buf BUF1 (N3600, N3595);
nand NAND4 (N3601, N3600, N1592, N3446, N943);
nand NAND4 (N3602, N3586, N1849, N2195, N284);
and AND3 (N3603, N3598, N976, N1224);
and AND4 (N3604, N3603, N1016, N2638, N2259);
xor XOR2 (N3605, N3597, N2941);
nor NOR4 (N3606, N3604, N2987, N1324, N2339);
and AND2 (N3607, N3585, N3240);
not NOT1 (N3608, N3605);
nor NOR4 (N3609, N3602, N2161, N1590, N670);
nand NAND4 (N3610, N3593, N533, N2930, N176);
buf BUF1 (N3611, N3601);
or OR2 (N3612, N3610, N2614);
nor NOR4 (N3613, N3589, N2986, N1521, N64);
nand NAND3 (N3614, N3607, N374, N3492);
buf BUF1 (N3615, N3613);
or OR3 (N3616, N3609, N2324, N1017);
or OR2 (N3617, N3606, N2112);
xor XOR2 (N3618, N3611, N2491);
buf BUF1 (N3619, N3608);
and AND2 (N3620, N3599, N1918);
not NOT1 (N3621, N3573);
buf BUF1 (N3622, N3621);
not NOT1 (N3623, N3572);
nor NOR2 (N3624, N3614, N363);
not NOT1 (N3625, N3620);
buf BUF1 (N3626, N3619);
and AND3 (N3627, N3617, N3077, N1626);
not NOT1 (N3628, N3622);
not NOT1 (N3629, N3627);
nor NOR3 (N3630, N3626, N507, N50);
not NOT1 (N3631, N3629);
buf BUF1 (N3632, N3630);
nor NOR4 (N3633, N3631, N2686, N2715, N3500);
and AND2 (N3634, N3623, N1706);
and AND3 (N3635, N3628, N1705, N1429);
not NOT1 (N3636, N3634);
not NOT1 (N3637, N3633);
and AND2 (N3638, N3624, N1159);
nor NOR2 (N3639, N3612, N854);
not NOT1 (N3640, N3618);
nand NAND3 (N3641, N3632, N1794, N771);
buf BUF1 (N3642, N3637);
xor XOR2 (N3643, N3616, N2556);
or OR3 (N3644, N3639, N1800, N1305);
nor NOR2 (N3645, N3642, N1128);
nand NAND2 (N3646, N3641, N400);
buf BUF1 (N3647, N3625);
nand NAND4 (N3648, N3615, N911, N998, N527);
nand NAND2 (N3649, N3636, N708);
nor NOR3 (N3650, N3646, N2567, N372);
nand NAND2 (N3651, N3647, N2694);
and AND4 (N3652, N3645, N1233, N796, N2142);
nor NOR3 (N3653, N3650, N2605, N64);
not NOT1 (N3654, N3651);
not NOT1 (N3655, N3649);
nand NAND3 (N3656, N3648, N3536, N294);
buf BUF1 (N3657, N3656);
nor NOR3 (N3658, N3655, N1391, N350);
and AND3 (N3659, N3653, N1056, N3577);
or OR4 (N3660, N3640, N979, N2219, N3395);
not NOT1 (N3661, N3644);
or OR4 (N3662, N3660, N1301, N1905, N2284);
and AND4 (N3663, N3657, N3349, N1759, N1093);
nor NOR3 (N3664, N3661, N2440, N90);
nor NOR4 (N3665, N3663, N3598, N2004, N1871);
nor NOR2 (N3666, N3658, N142);
xor XOR2 (N3667, N3654, N2309);
or OR2 (N3668, N3643, N3612);
or OR3 (N3669, N3662, N1159, N1538);
nor NOR2 (N3670, N3666, N2385);
and AND4 (N3671, N3669, N97, N1523, N2604);
xor XOR2 (N3672, N3665, N1773);
not NOT1 (N3673, N3659);
nor NOR3 (N3674, N3672, N111, N2345);
not NOT1 (N3675, N3652);
buf BUF1 (N3676, N3670);
nand NAND4 (N3677, N3667, N3039, N2932, N3410);
xor XOR2 (N3678, N3677, N719);
xor XOR2 (N3679, N3678, N650);
not NOT1 (N3680, N3675);
buf BUF1 (N3681, N3671);
not NOT1 (N3682, N3673);
buf BUF1 (N3683, N3681);
or OR3 (N3684, N3679, N1774, N2525);
nand NAND2 (N3685, N3683, N3285);
xor XOR2 (N3686, N3638, N1487);
not NOT1 (N3687, N3668);
nor NOR2 (N3688, N3682, N3459);
or OR4 (N3689, N3687, N2219, N2001, N1867);
nor NOR3 (N3690, N3676, N1404, N2236);
and AND4 (N3691, N3690, N2709, N1417, N1180);
not NOT1 (N3692, N3691);
nor NOR3 (N3693, N3664, N1498, N3581);
nor NOR3 (N3694, N3635, N65, N2824);
not NOT1 (N3695, N3686);
nand NAND2 (N3696, N3692, N1239);
and AND3 (N3697, N3674, N557, N1607);
buf BUF1 (N3698, N3697);
nor NOR4 (N3699, N3688, N1843, N3220, N1835);
not NOT1 (N3700, N3685);
buf BUF1 (N3701, N3695);
nand NAND4 (N3702, N3680, N3592, N3591, N3317);
or OR2 (N3703, N3684, N914);
buf BUF1 (N3704, N3694);
buf BUF1 (N3705, N3704);
or OR4 (N3706, N3703, N898, N2987, N1393);
buf BUF1 (N3707, N3696);
xor XOR2 (N3708, N3698, N1466);
xor XOR2 (N3709, N3708, N2829);
nand NAND2 (N3710, N3709, N803);
not NOT1 (N3711, N3705);
not NOT1 (N3712, N3706);
or OR2 (N3713, N3707, N2301);
nor NOR3 (N3714, N3711, N2498, N582);
or OR2 (N3715, N3693, N2738);
or OR3 (N3716, N3700, N1375, N3437);
and AND2 (N3717, N3689, N3164);
nor NOR3 (N3718, N3717, N801, N3131);
and AND3 (N3719, N3715, N428, N2730);
nand NAND2 (N3720, N3702, N1052);
or OR2 (N3721, N3719, N3449);
not NOT1 (N3722, N3710);
nand NAND4 (N3723, N3714, N2259, N601, N3471);
not NOT1 (N3724, N3718);
buf BUF1 (N3725, N3722);
not NOT1 (N3726, N3720);
nor NOR4 (N3727, N3726, N1830, N3337, N891);
buf BUF1 (N3728, N3699);
not NOT1 (N3729, N3721);
nor NOR2 (N3730, N3713, N327);
not NOT1 (N3731, N3723);
buf BUF1 (N3732, N3725);
buf BUF1 (N3733, N3727);
nor NOR3 (N3734, N3701, N2274, N2267);
or OR3 (N3735, N3732, N1078, N521);
nand NAND2 (N3736, N3729, N2346);
not NOT1 (N3737, N3733);
or OR3 (N3738, N3737, N1516, N1931);
not NOT1 (N3739, N3736);
nand NAND4 (N3740, N3724, N492, N650, N939);
nand NAND3 (N3741, N3728, N3563, N590);
nand NAND3 (N3742, N3716, N2834, N1009);
nor NOR4 (N3743, N3735, N97, N3547, N772);
nand NAND2 (N3744, N3730, N568);
not NOT1 (N3745, N3741);
or OR4 (N3746, N3745, N3668, N3407, N2338);
xor XOR2 (N3747, N3739, N717);
nor NOR2 (N3748, N3740, N2477);
buf BUF1 (N3749, N3743);
and AND3 (N3750, N3748, N1739, N2699);
and AND2 (N3751, N3712, N3561);
and AND2 (N3752, N3744, N2200);
nand NAND4 (N3753, N3731, N1333, N2531, N577);
not NOT1 (N3754, N3746);
not NOT1 (N3755, N3752);
buf BUF1 (N3756, N3742);
xor XOR2 (N3757, N3750, N1755);
and AND3 (N3758, N3757, N1938, N211);
nor NOR4 (N3759, N3738, N1072, N1211, N936);
nand NAND2 (N3760, N3747, N664);
or OR3 (N3761, N3755, N574, N2798);
buf BUF1 (N3762, N3754);
buf BUF1 (N3763, N3761);
not NOT1 (N3764, N3753);
or OR3 (N3765, N3749, N3683, N2350);
not NOT1 (N3766, N3760);
xor XOR2 (N3767, N3763, N1267);
xor XOR2 (N3768, N3759, N2402);
buf BUF1 (N3769, N3766);
nor NOR2 (N3770, N3764, N285);
buf BUF1 (N3771, N3767);
or OR4 (N3772, N3734, N318, N1651, N1176);
not NOT1 (N3773, N3765);
nand NAND2 (N3774, N3751, N2731);
or OR2 (N3775, N3773, N1454);
buf BUF1 (N3776, N3762);
buf BUF1 (N3777, N3756);
not NOT1 (N3778, N3771);
nor NOR3 (N3779, N3758, N268, N2665);
and AND2 (N3780, N3778, N2375);
or OR4 (N3781, N3779, N1942, N689, N2068);
buf BUF1 (N3782, N3781);
not NOT1 (N3783, N3782);
or OR3 (N3784, N3769, N804, N2930);
xor XOR2 (N3785, N3770, N1826);
xor XOR2 (N3786, N3776, N2909);
or OR2 (N3787, N3772, N1074);
nor NOR2 (N3788, N3784, N1853);
or OR3 (N3789, N3783, N1747, N1517);
or OR4 (N3790, N3789, N1035, N3168, N2086);
or OR4 (N3791, N3780, N2375, N787, N256);
nand NAND4 (N3792, N3791, N123, N3400, N558);
xor XOR2 (N3793, N3788, N64);
buf BUF1 (N3794, N3775);
nor NOR4 (N3795, N3786, N1412, N2279, N2574);
and AND4 (N3796, N3794, N2624, N1401, N747);
and AND4 (N3797, N3768, N218, N216, N2662);
xor XOR2 (N3798, N3785, N1095);
or OR3 (N3799, N3796, N2826, N3300);
nand NAND4 (N3800, N3792, N1937, N2998, N3114);
xor XOR2 (N3801, N3774, N830);
xor XOR2 (N3802, N3793, N57);
nor NOR2 (N3803, N3798, N1219);
xor XOR2 (N3804, N3787, N1188);
not NOT1 (N3805, N3803);
and AND3 (N3806, N3800, N1491, N3627);
or OR4 (N3807, N3804, N411, N474, N101);
not NOT1 (N3808, N3799);
nor NOR3 (N3809, N3797, N3045, N3114);
buf BUF1 (N3810, N3806);
xor XOR2 (N3811, N3805, N2852);
nand NAND3 (N3812, N3777, N1955, N3287);
or OR2 (N3813, N3801, N746);
and AND3 (N3814, N3809, N3169, N1179);
or OR3 (N3815, N3795, N3727, N3814);
xor XOR2 (N3816, N345, N3259);
nor NOR4 (N3817, N3815, N1689, N3742, N1203);
nor NOR3 (N3818, N3817, N2933, N2776);
nand NAND4 (N3819, N3808, N1119, N3291, N3307);
nor NOR3 (N3820, N3807, N906, N2032);
nor NOR2 (N3821, N3818, N3552);
nand NAND3 (N3822, N3816, N929, N1336);
nor NOR3 (N3823, N3802, N563, N296);
nor NOR4 (N3824, N3811, N2308, N2566, N1694);
and AND2 (N3825, N3824, N1173);
nor NOR2 (N3826, N3790, N1961);
nor NOR2 (N3827, N3825, N3158);
not NOT1 (N3828, N3826);
buf BUF1 (N3829, N3819);
nor NOR4 (N3830, N3829, N1933, N804, N124);
not NOT1 (N3831, N3820);
or OR3 (N3832, N3830, N2660, N1764);
buf BUF1 (N3833, N3828);
nand NAND2 (N3834, N3831, N1532);
nand NAND4 (N3835, N3827, N3063, N1952, N315);
nand NAND2 (N3836, N3832, N437);
xor XOR2 (N3837, N3834, N192);
buf BUF1 (N3838, N3810);
and AND3 (N3839, N3822, N453, N1730);
not NOT1 (N3840, N3835);
nor NOR4 (N3841, N3840, N3810, N3265, N3077);
nand NAND2 (N3842, N3838, N1193);
and AND4 (N3843, N3823, N938, N3553, N2321);
xor XOR2 (N3844, N3836, N1542);
and AND3 (N3845, N3813, N3078, N3629);
or OR2 (N3846, N3841, N555);
and AND4 (N3847, N3833, N295, N617, N1482);
or OR2 (N3848, N3847, N2568);
not NOT1 (N3849, N3848);
not NOT1 (N3850, N3839);
not NOT1 (N3851, N3821);
nor NOR4 (N3852, N3850, N2905, N391, N3801);
xor XOR2 (N3853, N3852, N3567);
buf BUF1 (N3854, N3837);
nand NAND4 (N3855, N3853, N2472, N433, N2294);
xor XOR2 (N3856, N3851, N3310);
xor XOR2 (N3857, N3812, N1930);
nor NOR3 (N3858, N3846, N2085, N3025);
buf BUF1 (N3859, N3844);
not NOT1 (N3860, N3859);
nand NAND4 (N3861, N3858, N2562, N847, N37);
xor XOR2 (N3862, N3856, N3532);
nand NAND3 (N3863, N3854, N2879, N873);
or OR3 (N3864, N3862, N3159, N1590);
nand NAND4 (N3865, N3842, N1549, N2434, N3387);
and AND3 (N3866, N3849, N533, N1548);
buf BUF1 (N3867, N3857);
or OR2 (N3868, N3845, N3582);
or OR4 (N3869, N3867, N2142, N578, N2411);
nor NOR2 (N3870, N3866, N3019);
xor XOR2 (N3871, N3870, N2552);
nor NOR2 (N3872, N3861, N3604);
nand NAND3 (N3873, N3872, N3618, N3072);
nor NOR3 (N3874, N3869, N3470, N1821);
or OR2 (N3875, N3865, N604);
nor NOR3 (N3876, N3860, N1486, N3800);
xor XOR2 (N3877, N3871, N1517);
and AND4 (N3878, N3876, N407, N2115, N1150);
or OR2 (N3879, N3875, N2914);
nor NOR2 (N3880, N3863, N1077);
xor XOR2 (N3881, N3864, N1854);
buf BUF1 (N3882, N3855);
buf BUF1 (N3883, N3881);
and AND4 (N3884, N3879, N996, N1853, N92);
not NOT1 (N3885, N3843);
buf BUF1 (N3886, N3873);
buf BUF1 (N3887, N3886);
or OR3 (N3888, N3880, N1201, N3728);
nand NAND2 (N3889, N3878, N2807);
buf BUF1 (N3890, N3887);
nand NAND4 (N3891, N3889, N160, N336, N993);
xor XOR2 (N3892, N3868, N2406);
nand NAND4 (N3893, N3890, N2368, N3192, N678);
nor NOR4 (N3894, N3877, N457, N790, N552);
nand NAND4 (N3895, N3892, N601, N2425, N1765);
nand NAND4 (N3896, N3893, N3436, N2547, N1603);
nor NOR3 (N3897, N3896, N2097, N1457);
xor XOR2 (N3898, N3891, N2486);
nor NOR3 (N3899, N3897, N396, N1207);
or OR3 (N3900, N3895, N2694, N98);
or OR4 (N3901, N3884, N3081, N3046, N354);
nand NAND2 (N3902, N3898, N2491);
xor XOR2 (N3903, N3874, N396);
buf BUF1 (N3904, N3883);
buf BUF1 (N3905, N3904);
nand NAND4 (N3906, N3900, N3873, N992, N80);
nand NAND4 (N3907, N3888, N2559, N384, N2039);
not NOT1 (N3908, N3906);
nor NOR3 (N3909, N3885, N3844, N618);
and AND4 (N3910, N3894, N289, N1269, N2960);
not NOT1 (N3911, N3907);
nand NAND4 (N3912, N3905, N2639, N3794, N3341);
not NOT1 (N3913, N3882);
xor XOR2 (N3914, N3908, N2275);
or OR2 (N3915, N3909, N1966);
not NOT1 (N3916, N3899);
and AND4 (N3917, N3916, N1505, N1084, N3871);
and AND4 (N3918, N3903, N3681, N157, N2554);
not NOT1 (N3919, N3913);
and AND3 (N3920, N3918, N2293, N1548);
nand NAND2 (N3921, N3919, N2156);
not NOT1 (N3922, N3921);
or OR4 (N3923, N3912, N1653, N3336, N3705);
nand NAND3 (N3924, N3901, N2542, N42);
not NOT1 (N3925, N3902);
not NOT1 (N3926, N3925);
not NOT1 (N3927, N3915);
buf BUF1 (N3928, N3917);
not NOT1 (N3929, N3924);
nor NOR4 (N3930, N3929, N3284, N2828, N416);
nor NOR2 (N3931, N3930, N2131);
not NOT1 (N3932, N3910);
buf BUF1 (N3933, N3911);
not NOT1 (N3934, N3914);
or OR2 (N3935, N3923, N2773);
xor XOR2 (N3936, N3928, N2742);
nand NAND4 (N3937, N3926, N1676, N2099, N1147);
xor XOR2 (N3938, N3927, N3078);
buf BUF1 (N3939, N3922);
nand NAND4 (N3940, N3931, N1691, N1998, N3130);
xor XOR2 (N3941, N3938, N1607);
xor XOR2 (N3942, N3933, N2095);
nand NAND4 (N3943, N3935, N1180, N3289, N198);
buf BUF1 (N3944, N3932);
or OR3 (N3945, N3936, N321, N2936);
xor XOR2 (N3946, N3945, N724);
buf BUF1 (N3947, N3943);
nand NAND3 (N3948, N3934, N2791, N3378);
nand NAND2 (N3949, N3940, N3122);
nor NOR2 (N3950, N3944, N3455);
not NOT1 (N3951, N3920);
or OR3 (N3952, N3942, N1152, N1311);
not NOT1 (N3953, N3950);
not NOT1 (N3954, N3952);
nand NAND2 (N3955, N3953, N231);
or OR3 (N3956, N3955, N2371, N2778);
nand NAND3 (N3957, N3951, N3570, N2208);
not NOT1 (N3958, N3949);
nor NOR3 (N3959, N3958, N2689, N520);
nand NAND2 (N3960, N3957, N3582);
xor XOR2 (N3961, N3941, N3259);
nor NOR2 (N3962, N3956, N2446);
or OR4 (N3963, N3962, N853, N1421, N2257);
and AND3 (N3964, N3963, N1184, N3795);
not NOT1 (N3965, N3946);
nor NOR4 (N3966, N3954, N3774, N1565, N2826);
not NOT1 (N3967, N3966);
buf BUF1 (N3968, N3967);
xor XOR2 (N3969, N3939, N1528);
or OR4 (N3970, N3937, N3407, N1444, N69);
xor XOR2 (N3971, N3969, N1822);
and AND3 (N3972, N3964, N1063, N1825);
and AND2 (N3973, N3965, N2050);
or OR4 (N3974, N3971, N2241, N2788, N2151);
not NOT1 (N3975, N3968);
nand NAND4 (N3976, N3948, N2793, N3336, N2662);
or OR4 (N3977, N3974, N1727, N3481, N3072);
nand NAND4 (N3978, N3970, N481, N712, N680);
and AND2 (N3979, N3947, N757);
nand NAND2 (N3980, N3959, N1993);
nor NOR4 (N3981, N3961, N2726, N3766, N3077);
nand NAND2 (N3982, N3972, N2065);
nand NAND2 (N3983, N3977, N126);
and AND4 (N3984, N3976, N3124, N2325, N2350);
buf BUF1 (N3985, N3983);
buf BUF1 (N3986, N3960);
nor NOR4 (N3987, N3986, N3482, N1418, N101);
nor NOR4 (N3988, N3984, N3647, N608, N361);
buf BUF1 (N3989, N3980);
nor NOR3 (N3990, N3981, N3228, N643);
nor NOR4 (N3991, N3988, N3690, N492, N42);
not NOT1 (N3992, N3985);
nand NAND2 (N3993, N3973, N1328);
nor NOR4 (N3994, N3991, N228, N2022, N3905);
nor NOR4 (N3995, N3992, N293, N2797, N1491);
or OR4 (N3996, N3975, N2415, N2628, N3914);
xor XOR2 (N3997, N3982, N683);
or OR2 (N3998, N3993, N3699);
buf BUF1 (N3999, N3996);
xor XOR2 (N4000, N3987, N2439);
nor NOR4 (N4001, N4000, N122, N2642, N2447);
or OR2 (N4002, N3999, N2495);
not NOT1 (N4003, N3978);
buf BUF1 (N4004, N3990);
buf BUF1 (N4005, N4001);
buf BUF1 (N4006, N3998);
or OR2 (N4007, N3997, N2652);
nor NOR4 (N4008, N4007, N1017, N1633, N1903);
and AND2 (N4009, N4002, N415);
buf BUF1 (N4010, N3994);
xor XOR2 (N4011, N4005, N452);
buf BUF1 (N4012, N4010);
nand NAND2 (N4013, N4011, N3292);
buf BUF1 (N4014, N4012);
nor NOR4 (N4015, N3979, N2461, N2888, N1357);
not NOT1 (N4016, N4004);
xor XOR2 (N4017, N4009, N2105);
buf BUF1 (N4018, N4013);
endmodule