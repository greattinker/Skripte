// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;

output N611,N622,N619,N609,N587,N621,N620,N617,N603,N623;

nand NAND2 (N24, N8, N7);
or OR4 (N25, N3, N22, N16, N10);
or OR3 (N26, N19, N5, N19);
nor NOR3 (N27, N7, N3, N2);
not NOT1 (N28, N6);
nand NAND3 (N29, N13, N21, N15);
or OR2 (N30, N3, N12);
nand NAND3 (N31, N12, N3, N28);
and AND4 (N32, N7, N17, N30, N6);
or OR4 (N33, N25, N5, N4, N14);
xor XOR2 (N34, N30, N33);
nor NOR4 (N35, N29, N32, N20, N3);
xor XOR2 (N36, N10, N9);
not NOT1 (N37, N23);
nor NOR4 (N38, N13, N21, N27, N29);
not NOT1 (N39, N19);
or OR2 (N40, N1, N11);
buf BUF1 (N41, N40);
not NOT1 (N42, N36);
nor NOR4 (N43, N26, N4, N36, N19);
and AND2 (N44, N35, N27);
nor NOR4 (N45, N39, N40, N12, N23);
or OR2 (N46, N44, N39);
not NOT1 (N47, N43);
or OR4 (N48, N41, N25, N45, N42);
not NOT1 (N49, N35);
nor NOR2 (N50, N6, N22);
nand NAND4 (N51, N34, N36, N15, N34);
not NOT1 (N52, N31);
and AND2 (N53, N52, N8);
nor NOR2 (N54, N51, N52);
not NOT1 (N55, N54);
xor XOR2 (N56, N37, N24);
buf BUF1 (N57, N31);
xor XOR2 (N58, N50, N34);
or OR3 (N59, N56, N6, N17);
nor NOR3 (N60, N53, N2, N21);
or OR3 (N61, N48, N23, N48);
and AND4 (N62, N49, N55, N45, N56);
not NOT1 (N63, N24);
xor XOR2 (N64, N59, N43);
buf BUF1 (N65, N47);
and AND2 (N66, N60, N5);
buf BUF1 (N67, N62);
buf BUF1 (N68, N38);
or OR2 (N69, N58, N31);
not NOT1 (N70, N65);
nand NAND2 (N71, N66, N26);
nor NOR2 (N72, N63, N68);
nand NAND2 (N73, N49, N46);
nand NAND4 (N74, N58, N70, N20, N52);
nand NAND4 (N75, N35, N37, N35, N53);
or OR2 (N76, N67, N37);
or OR4 (N77, N57, N2, N17, N71);
or OR2 (N78, N67, N22);
and AND3 (N79, N77, N44, N59);
not NOT1 (N80, N69);
or OR3 (N81, N78, N50, N28);
buf BUF1 (N82, N79);
nand NAND2 (N83, N80, N44);
nand NAND3 (N84, N72, N56, N1);
xor XOR2 (N85, N81, N76);
buf BUF1 (N86, N62);
not NOT1 (N87, N84);
not NOT1 (N88, N82);
or OR4 (N89, N64, N69, N13, N12);
and AND3 (N90, N74, N21, N85);
and AND3 (N91, N71, N15, N47);
not NOT1 (N92, N83);
xor XOR2 (N93, N88, N92);
xor XOR2 (N94, N58, N42);
and AND3 (N95, N75, N57, N9);
not NOT1 (N96, N87);
not NOT1 (N97, N86);
or OR2 (N98, N93, N49);
nand NAND3 (N99, N90, N58, N98);
and AND3 (N100, N4, N61, N89);
not NOT1 (N101, N72);
nor NOR3 (N102, N3, N44, N47);
or OR2 (N103, N73, N59);
buf BUF1 (N104, N95);
nor NOR4 (N105, N103, N55, N49, N19);
xor XOR2 (N106, N100, N38);
not NOT1 (N107, N105);
xor XOR2 (N108, N94, N30);
xor XOR2 (N109, N102, N19);
and AND2 (N110, N104, N74);
and AND3 (N111, N108, N80, N38);
nand NAND2 (N112, N107, N27);
nand NAND2 (N113, N109, N2);
not NOT1 (N114, N112);
nor NOR3 (N115, N101, N112, N29);
xor XOR2 (N116, N113, N31);
or OR2 (N117, N111, N4);
or OR3 (N118, N117, N65, N83);
not NOT1 (N119, N118);
xor XOR2 (N120, N119, N23);
or OR4 (N121, N110, N106, N59, N37);
and AND3 (N122, N97, N12, N85);
and AND4 (N123, N107, N96, N24, N1);
buf BUF1 (N124, N30);
not NOT1 (N125, N115);
nand NAND3 (N126, N123, N99, N52);
and AND3 (N127, N7, N86, N119);
or OR3 (N128, N120, N71, N6);
or OR2 (N129, N126, N13);
nand NAND4 (N130, N129, N84, N87, N86);
xor XOR2 (N131, N116, N37);
or OR3 (N132, N124, N13, N17);
nand NAND4 (N133, N114, N131, N90, N18);
buf BUF1 (N134, N104);
buf BUF1 (N135, N121);
nor NOR4 (N136, N127, N65, N20, N62);
or OR2 (N137, N125, N56);
buf BUF1 (N138, N128);
not NOT1 (N139, N135);
not NOT1 (N140, N130);
xor XOR2 (N141, N91, N95);
nor NOR3 (N142, N122, N16, N71);
nor NOR4 (N143, N137, N23, N98, N32);
buf BUF1 (N144, N133);
not NOT1 (N145, N140);
not NOT1 (N146, N132);
nor NOR2 (N147, N145, N5);
nand NAND4 (N148, N142, N141, N110, N19);
nor NOR2 (N149, N148, N60);
buf BUF1 (N150, N58);
and AND2 (N151, N134, N142);
nor NOR4 (N152, N139, N35, N60, N19);
or OR2 (N153, N143, N1);
nand NAND3 (N154, N151, N103, N132);
nor NOR4 (N155, N154, N148, N71, N106);
and AND2 (N156, N150, N27);
or OR3 (N157, N146, N84, N98);
and AND3 (N158, N157, N48, N48);
and AND3 (N159, N136, N150, N20);
or OR3 (N160, N158, N143, N133);
nor NOR2 (N161, N147, N75);
buf BUF1 (N162, N155);
and AND2 (N163, N153, N84);
and AND3 (N164, N159, N76, N143);
or OR3 (N165, N138, N123, N1);
not NOT1 (N166, N161);
and AND2 (N167, N160, N117);
nor NOR2 (N168, N152, N143);
or OR4 (N169, N166, N4, N68, N27);
nand NAND4 (N170, N167, N68, N99, N61);
and AND2 (N171, N169, N114);
and AND2 (N172, N163, N120);
and AND3 (N173, N172, N124, N93);
buf BUF1 (N174, N156);
and AND2 (N175, N165, N143);
nor NOR2 (N176, N170, N118);
not NOT1 (N177, N164);
xor XOR2 (N178, N144, N27);
nor NOR2 (N179, N175, N88);
not NOT1 (N180, N168);
or OR2 (N181, N171, N38);
or OR3 (N182, N177, N125, N135);
or OR4 (N183, N179, N72, N98, N14);
and AND2 (N184, N162, N177);
nand NAND3 (N185, N174, N62, N128);
or OR4 (N186, N181, N52, N103, N102);
not NOT1 (N187, N185);
xor XOR2 (N188, N180, N169);
and AND3 (N189, N183, N33, N141);
buf BUF1 (N190, N178);
buf BUF1 (N191, N149);
not NOT1 (N192, N189);
and AND2 (N193, N190, N119);
xor XOR2 (N194, N173, N152);
and AND3 (N195, N186, N116, N80);
nor NOR4 (N196, N194, N76, N65, N2);
buf BUF1 (N197, N187);
xor XOR2 (N198, N193, N106);
nand NAND3 (N199, N197, N132, N144);
nor NOR3 (N200, N191, N63, N153);
or OR2 (N201, N198, N11);
xor XOR2 (N202, N196, N7);
nand NAND2 (N203, N188, N126);
nand NAND3 (N204, N199, N117, N62);
xor XOR2 (N205, N176, N140);
buf BUF1 (N206, N205);
nand NAND3 (N207, N202, N72, N130);
and AND3 (N208, N206, N8, N155);
xor XOR2 (N209, N204, N136);
not NOT1 (N210, N195);
xor XOR2 (N211, N184, N62);
or OR2 (N212, N200, N110);
xor XOR2 (N213, N211, N183);
xor XOR2 (N214, N201, N106);
nand NAND4 (N215, N182, N111, N38, N149);
buf BUF1 (N216, N214);
not NOT1 (N217, N203);
buf BUF1 (N218, N217);
or OR4 (N219, N192, N11, N94, N140);
or OR3 (N220, N215, N146, N167);
or OR2 (N221, N216, N160);
not NOT1 (N222, N210);
not NOT1 (N223, N218);
and AND4 (N224, N208, N78, N96, N223);
xor XOR2 (N225, N56, N147);
xor XOR2 (N226, N209, N119);
or OR4 (N227, N220, N92, N147, N2);
buf BUF1 (N228, N221);
buf BUF1 (N229, N207);
nor NOR4 (N230, N225, N39, N44, N221);
or OR2 (N231, N222, N2);
not NOT1 (N232, N213);
not NOT1 (N233, N228);
or OR3 (N234, N224, N15, N104);
or OR4 (N235, N233, N189, N77, N180);
nor NOR4 (N236, N226, N192, N132, N36);
nor NOR4 (N237, N235, N123, N47, N212);
and AND3 (N238, N138, N180, N233);
or OR2 (N239, N236, N216);
xor XOR2 (N240, N237, N206);
or OR2 (N241, N234, N83);
or OR4 (N242, N238, N12, N212, N145);
or OR3 (N243, N230, N95, N50);
nor NOR3 (N244, N242, N178, N201);
xor XOR2 (N245, N219, N244);
nand NAND4 (N246, N210, N76, N202, N239);
not NOT1 (N247, N238);
nor NOR3 (N248, N229, N152, N28);
buf BUF1 (N249, N241);
xor XOR2 (N250, N227, N240);
or OR2 (N251, N110, N173);
nor NOR2 (N252, N250, N183);
nor NOR3 (N253, N252, N14, N6);
and AND3 (N254, N247, N14, N225);
and AND2 (N255, N245, N100);
and AND4 (N256, N249, N219, N49, N85);
and AND2 (N257, N254, N188);
xor XOR2 (N258, N248, N43);
nand NAND4 (N259, N257, N134, N23, N33);
nand NAND2 (N260, N232, N116);
nor NOR4 (N261, N243, N234, N221, N225);
xor XOR2 (N262, N246, N39);
nor NOR2 (N263, N231, N207);
and AND4 (N264, N262, N59, N27, N217);
not NOT1 (N265, N253);
or OR3 (N266, N261, N25, N148);
not NOT1 (N267, N258);
nor NOR4 (N268, N251, N194, N109, N169);
buf BUF1 (N269, N263);
nand NAND2 (N270, N255, N137);
nand NAND2 (N271, N264, N247);
and AND2 (N272, N271, N77);
nand NAND2 (N273, N268, N87);
and AND2 (N274, N269, N17);
nor NOR2 (N275, N273, N55);
and AND3 (N276, N260, N191, N77);
or OR2 (N277, N259, N106);
and AND4 (N278, N270, N103, N90, N11);
or OR2 (N279, N272, N60);
or OR2 (N280, N267, N273);
nor NOR2 (N281, N280, N19);
nor NOR4 (N282, N277, N134, N194, N36);
nand NAND2 (N283, N274, N255);
xor XOR2 (N284, N276, N197);
not NOT1 (N285, N266);
buf BUF1 (N286, N284);
and AND3 (N287, N265, N126, N266);
or OR3 (N288, N285, N198, N7);
buf BUF1 (N289, N286);
and AND4 (N290, N288, N281, N272, N274);
nand NAND3 (N291, N94, N216, N176);
nand NAND4 (N292, N256, N41, N240, N104);
and AND2 (N293, N290, N96);
nand NAND4 (N294, N282, N237, N1, N225);
buf BUF1 (N295, N283);
or OR2 (N296, N278, N138);
or OR2 (N297, N291, N190);
and AND4 (N298, N294, N175, N58, N185);
not NOT1 (N299, N287);
buf BUF1 (N300, N275);
and AND2 (N301, N300, N274);
xor XOR2 (N302, N299, N103);
or OR4 (N303, N295, N187, N72, N279);
and AND3 (N304, N290, N268, N260);
and AND2 (N305, N298, N158);
buf BUF1 (N306, N305);
or OR3 (N307, N306, N272, N233);
nand NAND2 (N308, N292, N60);
or OR3 (N309, N307, N164, N73);
buf BUF1 (N310, N308);
nand NAND2 (N311, N289, N50);
xor XOR2 (N312, N301, N70);
buf BUF1 (N313, N310);
and AND3 (N314, N297, N9, N30);
not NOT1 (N315, N309);
or OR2 (N316, N304, N118);
and AND3 (N317, N314, N38, N3);
buf BUF1 (N318, N303);
nor NOR4 (N319, N293, N159, N212, N49);
not NOT1 (N320, N319);
not NOT1 (N321, N312);
nor NOR4 (N322, N296, N92, N308, N8);
or OR4 (N323, N316, N6, N42, N73);
nor NOR4 (N324, N313, N220, N223, N151);
buf BUF1 (N325, N321);
nand NAND3 (N326, N322, N148, N284);
buf BUF1 (N327, N317);
and AND4 (N328, N323, N156, N28, N325);
or OR3 (N329, N315, N214, N198);
not NOT1 (N330, N267);
nand NAND3 (N331, N318, N42, N228);
buf BUF1 (N332, N331);
xor XOR2 (N333, N329, N222);
and AND3 (N334, N320, N59, N327);
not NOT1 (N335, N213);
buf BUF1 (N336, N333);
and AND4 (N337, N328, N160, N92, N189);
xor XOR2 (N338, N302, N78);
buf BUF1 (N339, N324);
nand NAND2 (N340, N339, N245);
nand NAND4 (N341, N336, N218, N101, N112);
xor XOR2 (N342, N340, N63);
xor XOR2 (N343, N335, N79);
not NOT1 (N344, N341);
buf BUF1 (N345, N334);
nand NAND3 (N346, N343, N19, N190);
xor XOR2 (N347, N344, N294);
buf BUF1 (N348, N346);
and AND3 (N349, N345, N53, N86);
nor NOR2 (N350, N342, N327);
buf BUF1 (N351, N330);
not NOT1 (N352, N347);
nor NOR4 (N353, N350, N348, N330, N169);
nand NAND3 (N354, N179, N62, N92);
nand NAND2 (N355, N351, N342);
xor XOR2 (N356, N355, N61);
nand NAND4 (N357, N354, N68, N90, N337);
xor XOR2 (N358, N173, N280);
and AND3 (N359, N352, N227, N156);
not NOT1 (N360, N326);
xor XOR2 (N361, N356, N316);
nor NOR2 (N362, N332, N138);
not NOT1 (N363, N359);
xor XOR2 (N364, N357, N324);
not NOT1 (N365, N353);
nand NAND2 (N366, N361, N9);
nor NOR4 (N367, N349, N185, N111, N294);
nor NOR3 (N368, N338, N112, N158);
and AND4 (N369, N368, N80, N157, N328);
or OR4 (N370, N360, N17, N40, N184);
buf BUF1 (N371, N311);
buf BUF1 (N372, N366);
nor NOR2 (N373, N370, N189);
nor NOR3 (N374, N362, N276, N34);
or OR2 (N375, N358, N263);
and AND4 (N376, N373, N170, N259, N212);
nor NOR4 (N377, N372, N291, N296, N31);
and AND4 (N378, N364, N341, N167, N260);
buf BUF1 (N379, N377);
not NOT1 (N380, N379);
nand NAND3 (N381, N376, N99, N316);
and AND3 (N382, N381, N207, N7);
and AND4 (N383, N382, N332, N362, N328);
nand NAND3 (N384, N374, N292, N216);
buf BUF1 (N385, N384);
nor NOR4 (N386, N363, N373, N104, N383);
nor NOR2 (N387, N182, N342);
buf BUF1 (N388, N369);
nor NOR4 (N389, N367, N340, N376, N50);
not NOT1 (N390, N387);
buf BUF1 (N391, N385);
buf BUF1 (N392, N378);
or OR4 (N393, N386, N10, N198, N366);
buf BUF1 (N394, N388);
buf BUF1 (N395, N375);
not NOT1 (N396, N371);
not NOT1 (N397, N393);
buf BUF1 (N398, N390);
xor XOR2 (N399, N391, N84);
buf BUF1 (N400, N398);
xor XOR2 (N401, N396, N268);
xor XOR2 (N402, N397, N332);
and AND3 (N403, N401, N201, N47);
buf BUF1 (N404, N400);
and AND2 (N405, N404, N180);
nand NAND3 (N406, N395, N336, N292);
or OR3 (N407, N406, N386, N196);
buf BUF1 (N408, N402);
xor XOR2 (N409, N399, N144);
nand NAND2 (N410, N409, N37);
buf BUF1 (N411, N405);
nor NOR4 (N412, N411, N353, N283, N42);
buf BUF1 (N413, N410);
buf BUF1 (N414, N389);
not NOT1 (N415, N414);
not NOT1 (N416, N394);
buf BUF1 (N417, N408);
buf BUF1 (N418, N415);
nand NAND4 (N419, N380, N361, N344, N356);
and AND3 (N420, N413, N252, N164);
or OR4 (N421, N420, N240, N28, N138);
and AND2 (N422, N419, N421);
nor NOR2 (N423, N394, N78);
nand NAND3 (N424, N416, N162, N375);
xor XOR2 (N425, N418, N180);
buf BUF1 (N426, N403);
buf BUF1 (N427, N423);
buf BUF1 (N428, N365);
or OR2 (N429, N428, N388);
or OR4 (N430, N412, N250, N211, N51);
nand NAND3 (N431, N424, N324, N279);
and AND4 (N432, N429, N424, N143, N225);
buf BUF1 (N433, N422);
buf BUF1 (N434, N430);
xor XOR2 (N435, N434, N167);
not NOT1 (N436, N392);
or OR4 (N437, N425, N7, N399, N32);
buf BUF1 (N438, N435);
not NOT1 (N439, N433);
xor XOR2 (N440, N439, N241);
nor NOR4 (N441, N436, N85, N206, N277);
and AND4 (N442, N407, N355, N126, N231);
buf BUF1 (N443, N427);
nand NAND4 (N444, N438, N161, N74, N185);
buf BUF1 (N445, N441);
and AND2 (N446, N437, N432);
or OR2 (N447, N116, N364);
buf BUF1 (N448, N417);
not NOT1 (N449, N447);
nand NAND3 (N450, N445, N212, N374);
not NOT1 (N451, N448);
nand NAND3 (N452, N451, N217, N209);
nand NAND4 (N453, N446, N230, N341, N139);
or OR4 (N454, N442, N45, N138, N414);
nor NOR4 (N455, N444, N225, N79, N69);
and AND4 (N456, N450, N281, N112, N221);
nor NOR4 (N457, N456, N396, N53, N200);
or OR3 (N458, N457, N402, N273);
nor NOR2 (N459, N443, N420);
nand NAND2 (N460, N459, N31);
and AND3 (N461, N454, N258, N31);
nor NOR3 (N462, N440, N461, N58);
nor NOR3 (N463, N360, N343, N248);
nor NOR4 (N464, N431, N12, N300, N392);
or OR2 (N465, N460, N420);
buf BUF1 (N466, N464);
buf BUF1 (N467, N453);
not NOT1 (N468, N467);
nor NOR2 (N469, N462, N234);
not NOT1 (N470, N465);
buf BUF1 (N471, N455);
and AND4 (N472, N426, N352, N10, N440);
nand NAND2 (N473, N458, N226);
or OR3 (N474, N469, N45, N56);
nor NOR2 (N475, N463, N301);
or OR4 (N476, N470, N419, N326, N340);
not NOT1 (N477, N452);
buf BUF1 (N478, N449);
buf BUF1 (N479, N473);
or OR2 (N480, N472, N51);
not NOT1 (N481, N480);
or OR4 (N482, N468, N6, N47, N10);
nor NOR3 (N483, N479, N369, N34);
buf BUF1 (N484, N481);
buf BUF1 (N485, N478);
nand NAND4 (N486, N475, N302, N176, N110);
or OR3 (N487, N484, N60, N241);
buf BUF1 (N488, N485);
not NOT1 (N489, N471);
buf BUF1 (N490, N482);
xor XOR2 (N491, N477, N432);
buf BUF1 (N492, N488);
nand NAND3 (N493, N486, N192, N342);
nor NOR2 (N494, N483, N158);
or OR2 (N495, N492, N346);
and AND2 (N496, N491, N177);
nand NAND4 (N497, N489, N324, N396, N449);
not NOT1 (N498, N493);
xor XOR2 (N499, N490, N141);
and AND2 (N500, N498, N151);
nor NOR4 (N501, N494, N373, N299, N379);
not NOT1 (N502, N474);
and AND4 (N503, N500, N119, N483, N402);
nand NAND2 (N504, N502, N191);
not NOT1 (N505, N501);
xor XOR2 (N506, N487, N95);
buf BUF1 (N507, N476);
nor NOR3 (N508, N495, N115, N339);
xor XOR2 (N509, N466, N66);
xor XOR2 (N510, N499, N212);
not NOT1 (N511, N503);
nor NOR2 (N512, N511, N220);
or OR2 (N513, N505, N299);
or OR2 (N514, N513, N274);
buf BUF1 (N515, N512);
not NOT1 (N516, N497);
buf BUF1 (N517, N506);
and AND4 (N518, N496, N168, N105, N269);
buf BUF1 (N519, N507);
and AND3 (N520, N516, N122, N137);
xor XOR2 (N521, N510, N366);
and AND2 (N522, N504, N102);
and AND3 (N523, N522, N231, N413);
nand NAND3 (N524, N509, N353, N382);
xor XOR2 (N525, N517, N276);
and AND3 (N526, N525, N497, N18);
or OR4 (N527, N518, N223, N150, N306);
and AND2 (N528, N521, N221);
nor NOR4 (N529, N527, N427, N121, N448);
and AND3 (N530, N524, N261, N183);
buf BUF1 (N531, N530);
not NOT1 (N532, N519);
not NOT1 (N533, N508);
buf BUF1 (N534, N531);
xor XOR2 (N535, N515, N114);
buf BUF1 (N536, N535);
not NOT1 (N537, N532);
not NOT1 (N538, N534);
xor XOR2 (N539, N528, N184);
xor XOR2 (N540, N537, N139);
buf BUF1 (N541, N538);
nor NOR2 (N542, N523, N381);
or OR2 (N543, N514, N496);
and AND2 (N544, N543, N174);
nor NOR2 (N545, N526, N280);
and AND4 (N546, N536, N316, N128, N314);
nor NOR2 (N547, N541, N202);
and AND3 (N548, N529, N350, N544);
not NOT1 (N549, N250);
or OR4 (N550, N547, N1, N146, N93);
nor NOR3 (N551, N542, N470, N400);
nand NAND4 (N552, N550, N128, N464, N191);
and AND4 (N553, N551, N197, N221, N153);
not NOT1 (N554, N553);
nand NAND2 (N555, N549, N81);
nor NOR4 (N556, N548, N92, N267, N245);
not NOT1 (N557, N552);
or OR3 (N558, N545, N337, N109);
xor XOR2 (N559, N554, N178);
nor NOR3 (N560, N546, N288, N161);
nand NAND4 (N561, N556, N403, N328, N388);
or OR3 (N562, N533, N148, N343);
xor XOR2 (N563, N559, N402);
buf BUF1 (N564, N561);
buf BUF1 (N565, N539);
nor NOR3 (N566, N562, N261, N2);
nor NOR3 (N567, N563, N255, N450);
and AND3 (N568, N560, N18, N355);
buf BUF1 (N569, N566);
xor XOR2 (N570, N565, N452);
or OR3 (N571, N570, N380, N130);
xor XOR2 (N572, N571, N516);
nand NAND4 (N573, N569, N434, N113, N199);
xor XOR2 (N574, N540, N125);
and AND4 (N575, N573, N436, N156, N252);
or OR3 (N576, N574, N312, N364);
or OR2 (N577, N555, N55);
buf BUF1 (N578, N557);
xor XOR2 (N579, N567, N290);
and AND3 (N580, N520, N44, N94);
nor NOR3 (N581, N580, N434, N341);
buf BUF1 (N582, N572);
or OR2 (N583, N579, N232);
nand NAND3 (N584, N576, N507, N483);
buf BUF1 (N585, N577);
nor NOR2 (N586, N558, N155);
or OR3 (N587, N578, N303, N538);
or OR3 (N588, N582, N361, N177);
or OR3 (N589, N568, N163, N91);
buf BUF1 (N590, N575);
nor NOR2 (N591, N581, N112);
not NOT1 (N592, N564);
and AND4 (N593, N584, N112, N315, N458);
not NOT1 (N594, N589);
nor NOR2 (N595, N585, N207);
not NOT1 (N596, N592);
not NOT1 (N597, N591);
and AND4 (N598, N588, N548, N56, N34);
buf BUF1 (N599, N590);
not NOT1 (N600, N586);
not NOT1 (N601, N593);
nand NAND4 (N602, N601, N120, N45, N470);
buf BUF1 (N603, N599);
nand NAND4 (N604, N598, N84, N142, N226);
xor XOR2 (N605, N597, N26);
or OR4 (N606, N594, N565, N435, N287);
xor XOR2 (N607, N602, N513);
buf BUF1 (N608, N606);
nor NOR2 (N609, N607, N32);
xor XOR2 (N610, N583, N532);
nand NAND4 (N611, N605, N51, N216, N194);
not NOT1 (N612, N600);
not NOT1 (N613, N596);
and AND4 (N614, N608, N294, N508, N279);
buf BUF1 (N615, N610);
nor NOR3 (N616, N604, N28, N169);
nor NOR2 (N617, N613, N394);
buf BUF1 (N618, N595);
or OR3 (N619, N616, N163, N541);
xor XOR2 (N620, N618, N123);
xor XOR2 (N621, N615, N149);
buf BUF1 (N622, N612);
nor NOR3 (N623, N614, N505, N59);
endmodule