// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10;

output N4007,N4008,N3995,N3990,N4003,N4005,N4009,N3986,N4004,N4010;

not NOT1 (N11, N5);
buf BUF1 (N12, N8);
nand NAND3 (N13, N8, N12, N10);
nor NOR4 (N14, N5, N5, N7, N9);
xor XOR2 (N15, N1, N6);
not NOT1 (N16, N11);
xor XOR2 (N17, N12, N2);
nand NAND3 (N18, N16, N14, N17);
nand NAND4 (N19, N13, N13, N2, N17);
nor NOR4 (N20, N12, N18, N10, N9);
nand NAND2 (N21, N5, N14);
or OR2 (N22, N9, N2);
nand NAND4 (N23, N1, N3, N21, N3);
buf BUF1 (N24, N8);
and AND2 (N25, N11, N9);
and AND4 (N26, N6, N24, N4, N11);
buf BUF1 (N27, N18);
and AND3 (N28, N11, N11, N19);
nor NOR2 (N29, N13, N25);
xor XOR2 (N30, N2, N13);
nor NOR4 (N31, N27, N11, N14, N2);
nor NOR2 (N32, N27, N11);
xor XOR2 (N33, N20, N3);
and AND4 (N34, N33, N33, N30, N21);
xor XOR2 (N35, N34, N19);
or OR2 (N36, N31, N31);
nor NOR4 (N37, N10, N28, N20, N15);
xor XOR2 (N38, N5, N12);
not NOT1 (N39, N1);
nor NOR2 (N40, N26, N28);
and AND4 (N41, N40, N38, N9, N6);
nand NAND2 (N42, N19, N25);
not NOT1 (N43, N41);
nand NAND3 (N44, N29, N11, N31);
buf BUF1 (N45, N43);
buf BUF1 (N46, N44);
nor NOR4 (N47, N45, N46, N43, N8);
and AND2 (N48, N36, N44);
and AND4 (N49, N35, N5, N14, N11);
nor NOR3 (N50, N49, N41, N1);
and AND2 (N51, N37, N42);
and AND3 (N52, N17, N37, N39);
buf BUF1 (N53, N8);
buf BUF1 (N54, N13);
nand NAND3 (N55, N22, N23, N25);
or OR2 (N56, N36, N22);
or OR3 (N57, N55, N54, N17);
and AND3 (N58, N20, N29, N25);
nor NOR2 (N59, N48, N33);
and AND2 (N60, N52, N38);
nor NOR2 (N61, N47, N32);
not NOT1 (N62, N47);
xor XOR2 (N63, N62, N52);
xor XOR2 (N64, N60, N14);
nor NOR4 (N65, N63, N23, N48, N57);
and AND3 (N66, N31, N22, N61);
buf BUF1 (N67, N27);
nor NOR3 (N68, N59, N15, N28);
or OR3 (N69, N64, N26, N10);
nor NOR2 (N70, N65, N16);
or OR4 (N71, N51, N21, N16, N15);
or OR4 (N72, N69, N69, N43, N47);
and AND2 (N73, N53, N56);
xor XOR2 (N74, N35, N48);
nand NAND2 (N75, N72, N72);
or OR2 (N76, N73, N18);
or OR4 (N77, N50, N69, N55, N4);
buf BUF1 (N78, N66);
xor XOR2 (N79, N67, N59);
nand NAND2 (N80, N76, N20);
not NOT1 (N81, N79);
not NOT1 (N82, N78);
and AND4 (N83, N71, N19, N70, N19);
nor NOR3 (N84, N27, N32, N26);
buf BUF1 (N85, N80);
nand NAND4 (N86, N68, N27, N78, N70);
buf BUF1 (N87, N81);
xor XOR2 (N88, N77, N40);
nand NAND4 (N89, N83, N43, N15, N10);
xor XOR2 (N90, N85, N70);
buf BUF1 (N91, N75);
nand NAND2 (N92, N58, N63);
buf BUF1 (N93, N88);
xor XOR2 (N94, N91, N1);
and AND2 (N95, N87, N70);
and AND2 (N96, N89, N22);
nand NAND2 (N97, N92, N71);
buf BUF1 (N98, N84);
xor XOR2 (N99, N96, N86);
not NOT1 (N100, N58);
xor XOR2 (N101, N94, N84);
xor XOR2 (N102, N90, N64);
nor NOR4 (N103, N82, N67, N68, N7);
xor XOR2 (N104, N100, N48);
or OR3 (N105, N74, N66, N76);
nand NAND2 (N106, N95, N25);
or OR3 (N107, N103, N14, N57);
buf BUF1 (N108, N98);
or OR4 (N109, N93, N15, N42, N33);
nor NOR2 (N110, N107, N99);
not NOT1 (N111, N20);
xor XOR2 (N112, N104, N75);
xor XOR2 (N113, N105, N75);
or OR2 (N114, N102, N113);
nand NAND3 (N115, N95, N95, N41);
nor NOR4 (N116, N115, N107, N105, N69);
buf BUF1 (N117, N101);
xor XOR2 (N118, N108, N48);
not NOT1 (N119, N116);
nand NAND4 (N120, N114, N117, N31, N40);
xor XOR2 (N121, N3, N30);
xor XOR2 (N122, N106, N105);
and AND4 (N123, N122, N53, N80, N84);
nand NAND3 (N124, N119, N97, N36);
or OR4 (N125, N104, N65, N119, N109);
nor NOR3 (N126, N23, N9, N19);
xor XOR2 (N127, N110, N108);
buf BUF1 (N128, N112);
nand NAND3 (N129, N120, N27, N74);
and AND4 (N130, N125, N40, N102, N76);
nor NOR2 (N131, N127, N50);
not NOT1 (N132, N126);
xor XOR2 (N133, N124, N113);
buf BUF1 (N134, N131);
nand NAND2 (N135, N130, N90);
buf BUF1 (N136, N123);
not NOT1 (N137, N128);
not NOT1 (N138, N111);
and AND2 (N139, N118, N54);
nand NAND2 (N140, N137, N91);
not NOT1 (N141, N134);
nand NAND4 (N142, N141, N112, N106, N141);
and AND3 (N143, N138, N96, N90);
and AND3 (N144, N139, N69, N115);
buf BUF1 (N145, N140);
nand NAND3 (N146, N145, N3, N114);
not NOT1 (N147, N135);
or OR2 (N148, N133, N34);
and AND3 (N149, N147, N24, N56);
buf BUF1 (N150, N144);
nor NOR3 (N151, N148, N55, N143);
xor XOR2 (N152, N41, N143);
and AND3 (N153, N132, N109, N2);
nand NAND3 (N154, N151, N99, N46);
nor NOR2 (N155, N121, N98);
not NOT1 (N156, N136);
nand NAND4 (N157, N152, N33, N22, N134);
xor XOR2 (N158, N129, N24);
not NOT1 (N159, N154);
nand NAND4 (N160, N146, N143, N25, N76);
xor XOR2 (N161, N155, N103);
not NOT1 (N162, N159);
and AND3 (N163, N160, N116, N53);
xor XOR2 (N164, N149, N75);
not NOT1 (N165, N156);
nand NAND4 (N166, N164, N13, N35, N105);
buf BUF1 (N167, N162);
or OR4 (N168, N161, N165, N122, N95);
not NOT1 (N169, N57);
nand NAND3 (N170, N169, N142, N115);
nor NOR2 (N171, N95, N118);
or OR3 (N172, N171, N90, N36);
xor XOR2 (N173, N168, N113);
nand NAND4 (N174, N166, N143, N172, N29);
and AND3 (N175, N34, N126, N6);
xor XOR2 (N176, N153, N29);
and AND4 (N177, N176, N24, N171, N18);
or OR4 (N178, N163, N171, N172, N7);
or OR3 (N179, N175, N143, N77);
or OR2 (N180, N179, N18);
and AND3 (N181, N167, N87, N81);
buf BUF1 (N182, N180);
or OR4 (N183, N181, N112, N124, N35);
and AND3 (N184, N150, N152, N167);
buf BUF1 (N185, N174);
or OR3 (N186, N185, N170, N32);
xor XOR2 (N187, N159, N65);
and AND4 (N188, N182, N173, N56, N162);
not NOT1 (N189, N70);
or OR2 (N190, N177, N48);
and AND4 (N191, N158, N119, N97, N91);
and AND3 (N192, N187, N21, N91);
nand NAND2 (N193, N178, N170);
buf BUF1 (N194, N188);
buf BUF1 (N195, N189);
buf BUF1 (N196, N191);
nor NOR3 (N197, N186, N164, N189);
nand NAND4 (N198, N196, N137, N61, N16);
xor XOR2 (N199, N190, N161);
not NOT1 (N200, N184);
not NOT1 (N201, N157);
not NOT1 (N202, N199);
or OR4 (N203, N197, N183, N176, N11);
buf BUF1 (N204, N184);
xor XOR2 (N205, N195, N115);
buf BUF1 (N206, N200);
or OR4 (N207, N204, N138, N56, N6);
or OR3 (N208, N203, N182, N131);
xor XOR2 (N209, N194, N22);
not NOT1 (N210, N206);
and AND4 (N211, N205, N157, N174, N175);
nor NOR2 (N212, N201, N98);
nor NOR4 (N213, N207, N181, N2, N60);
not NOT1 (N214, N213);
xor XOR2 (N215, N198, N17);
and AND3 (N216, N215, N4, N15);
xor XOR2 (N217, N209, N58);
or OR4 (N218, N217, N91, N62, N88);
nor NOR3 (N219, N210, N151, N158);
nor NOR4 (N220, N202, N187, N115, N4);
and AND2 (N221, N211, N24);
or OR2 (N222, N212, N92);
buf BUF1 (N223, N193);
and AND4 (N224, N192, N79, N150, N53);
or OR4 (N225, N220, N170, N90, N117);
and AND2 (N226, N222, N63);
not NOT1 (N227, N225);
and AND3 (N228, N221, N48, N188);
nand NAND4 (N229, N224, N173, N9, N153);
xor XOR2 (N230, N216, N64);
nor NOR2 (N231, N226, N94);
buf BUF1 (N232, N214);
xor XOR2 (N233, N223, N182);
or OR2 (N234, N208, N44);
xor XOR2 (N235, N232, N226);
xor XOR2 (N236, N227, N193);
and AND3 (N237, N234, N98, N66);
nor NOR2 (N238, N230, N55);
and AND2 (N239, N219, N24);
or OR3 (N240, N233, N39, N116);
and AND3 (N241, N239, N82, N38);
xor XOR2 (N242, N240, N208);
buf BUF1 (N243, N237);
not NOT1 (N244, N218);
nor NOR2 (N245, N238, N79);
or OR4 (N246, N231, N195, N61, N100);
or OR2 (N247, N228, N1);
or OR2 (N248, N245, N206);
nand NAND4 (N249, N241, N107, N191, N144);
xor XOR2 (N250, N243, N30);
not NOT1 (N251, N235);
nand NAND2 (N252, N246, N97);
or OR2 (N253, N229, N217);
not NOT1 (N254, N253);
not NOT1 (N255, N251);
and AND4 (N256, N247, N212, N177, N145);
nand NAND2 (N257, N236, N66);
nor NOR3 (N258, N249, N173, N106);
buf BUF1 (N259, N256);
nand NAND3 (N260, N259, N45, N178);
or OR3 (N261, N255, N180, N92);
or OR3 (N262, N260, N68, N147);
nor NOR3 (N263, N261, N3, N71);
nand NAND4 (N264, N254, N1, N101, N79);
buf BUF1 (N265, N264);
or OR4 (N266, N263, N179, N167, N196);
buf BUF1 (N267, N242);
xor XOR2 (N268, N244, N215);
not NOT1 (N269, N252);
or OR4 (N270, N268, N2, N9, N8);
nand NAND3 (N271, N267, N91, N228);
buf BUF1 (N272, N266);
or OR3 (N273, N270, N88, N61);
and AND2 (N274, N258, N202);
nor NOR4 (N275, N271, N219, N87, N30);
and AND2 (N276, N273, N54);
not NOT1 (N277, N262);
or OR3 (N278, N274, N197, N219);
or OR2 (N279, N250, N16);
xor XOR2 (N280, N277, N59);
and AND4 (N281, N257, N137, N48, N92);
xor XOR2 (N282, N280, N45);
xor XOR2 (N283, N279, N1);
nand NAND3 (N284, N281, N143, N48);
buf BUF1 (N285, N276);
not NOT1 (N286, N284);
xor XOR2 (N287, N269, N80);
or OR3 (N288, N282, N226, N278);
nand NAND2 (N289, N131, N62);
nor NOR4 (N290, N288, N28, N110, N255);
buf BUF1 (N291, N287);
buf BUF1 (N292, N285);
not NOT1 (N293, N286);
and AND3 (N294, N283, N187, N46);
or OR4 (N295, N265, N11, N190, N132);
nand NAND3 (N296, N272, N20, N228);
nor NOR4 (N297, N293, N157, N249, N62);
nor NOR3 (N298, N292, N88, N219);
buf BUF1 (N299, N275);
and AND3 (N300, N297, N296, N2);
nor NOR3 (N301, N229, N91, N14);
and AND4 (N302, N301, N137, N127, N157);
nor NOR4 (N303, N300, N169, N225, N44);
nor NOR2 (N304, N294, N131);
and AND2 (N305, N248, N97);
nand NAND3 (N306, N291, N193, N183);
xor XOR2 (N307, N295, N7);
and AND3 (N308, N290, N98, N136);
not NOT1 (N309, N299);
and AND2 (N310, N303, N125);
buf BUF1 (N311, N307);
or OR3 (N312, N309, N57, N85);
and AND3 (N313, N304, N245, N293);
not NOT1 (N314, N305);
or OR3 (N315, N312, N221, N266);
nor NOR2 (N316, N306, N88);
and AND3 (N317, N302, N68, N256);
and AND2 (N318, N311, N70);
nor NOR3 (N319, N308, N251, N118);
not NOT1 (N320, N289);
or OR4 (N321, N320, N135, N78, N107);
nor NOR2 (N322, N310, N94);
buf BUF1 (N323, N314);
not NOT1 (N324, N323);
and AND2 (N325, N324, N265);
buf BUF1 (N326, N321);
and AND3 (N327, N316, N15, N140);
xor XOR2 (N328, N317, N309);
nand NAND3 (N329, N319, N91, N35);
buf BUF1 (N330, N313);
or OR2 (N331, N329, N115);
xor XOR2 (N332, N318, N161);
nand NAND3 (N333, N332, N127, N21);
not NOT1 (N334, N327);
xor XOR2 (N335, N334, N45);
or OR3 (N336, N331, N197, N138);
xor XOR2 (N337, N335, N170);
and AND4 (N338, N315, N48, N178, N41);
nor NOR4 (N339, N330, N295, N38, N126);
xor XOR2 (N340, N322, N52);
not NOT1 (N341, N328);
not NOT1 (N342, N337);
nand NAND3 (N343, N339, N207, N234);
or OR3 (N344, N325, N292, N81);
and AND2 (N345, N336, N291);
xor XOR2 (N346, N326, N46);
not NOT1 (N347, N344);
nand NAND2 (N348, N298, N89);
buf BUF1 (N349, N333);
not NOT1 (N350, N348);
not NOT1 (N351, N343);
buf BUF1 (N352, N338);
buf BUF1 (N353, N346);
nand NAND3 (N354, N340, N300, N112);
xor XOR2 (N355, N345, N339);
xor XOR2 (N356, N355, N62);
not NOT1 (N357, N353);
nor NOR3 (N358, N349, N4, N104);
and AND4 (N359, N350, N253, N61, N314);
buf BUF1 (N360, N351);
nand NAND4 (N361, N341, N13, N70, N62);
buf BUF1 (N362, N354);
buf BUF1 (N363, N359);
xor XOR2 (N364, N356, N132);
and AND4 (N365, N347, N261, N134, N224);
nor NOR2 (N366, N365, N256);
not NOT1 (N367, N357);
xor XOR2 (N368, N352, N246);
not NOT1 (N369, N364);
nor NOR4 (N370, N366, N365, N145, N332);
xor XOR2 (N371, N370, N169);
and AND3 (N372, N360, N75, N249);
not NOT1 (N373, N369);
not NOT1 (N374, N371);
or OR4 (N375, N342, N134, N142, N238);
xor XOR2 (N376, N363, N189);
and AND3 (N377, N361, N302, N163);
nor NOR2 (N378, N375, N357);
xor XOR2 (N379, N378, N315);
xor XOR2 (N380, N373, N168);
xor XOR2 (N381, N368, N204);
or OR4 (N382, N374, N236, N381, N93);
buf BUF1 (N383, N373);
xor XOR2 (N384, N376, N148);
nor NOR4 (N385, N384, N203, N324, N176);
and AND4 (N386, N385, N308, N306, N146);
or OR2 (N387, N362, N287);
buf BUF1 (N388, N380);
and AND3 (N389, N388, N57, N186);
not NOT1 (N390, N367);
xor XOR2 (N391, N358, N13);
buf BUF1 (N392, N383);
xor XOR2 (N393, N389, N216);
nand NAND3 (N394, N387, N154, N12);
and AND2 (N395, N390, N167);
or OR2 (N396, N379, N370);
xor XOR2 (N397, N391, N386);
and AND4 (N398, N130, N64, N35, N369);
and AND3 (N399, N382, N360, N224);
or OR3 (N400, N397, N81, N186);
nor NOR2 (N401, N377, N256);
nor NOR2 (N402, N394, N82);
buf BUF1 (N403, N372);
or OR2 (N404, N396, N243);
or OR3 (N405, N395, N122, N123);
buf BUF1 (N406, N398);
xor XOR2 (N407, N405, N1);
or OR2 (N408, N392, N303);
not NOT1 (N409, N403);
not NOT1 (N410, N402);
nor NOR4 (N411, N410, N331, N175, N95);
nand NAND4 (N412, N393, N79, N269, N131);
xor XOR2 (N413, N409, N392);
or OR4 (N414, N411, N59, N212, N111);
xor XOR2 (N415, N400, N143);
or OR2 (N416, N399, N198);
not NOT1 (N417, N401);
or OR4 (N418, N413, N20, N20, N110);
and AND2 (N419, N407, N368);
buf BUF1 (N420, N417);
not NOT1 (N421, N404);
xor XOR2 (N422, N419, N265);
buf BUF1 (N423, N406);
nor NOR2 (N424, N408, N340);
buf BUF1 (N425, N414);
and AND4 (N426, N422, N185, N187, N319);
buf BUF1 (N427, N418);
xor XOR2 (N428, N424, N381);
or OR4 (N429, N420, N17, N421, N26);
and AND4 (N430, N361, N364, N107, N185);
nand NAND4 (N431, N428, N11, N229, N33);
buf BUF1 (N432, N426);
xor XOR2 (N433, N412, N339);
xor XOR2 (N434, N429, N142);
and AND4 (N435, N434, N425, N286, N416);
buf BUF1 (N436, N206);
buf BUF1 (N437, N237);
not NOT1 (N438, N436);
not NOT1 (N439, N431);
buf BUF1 (N440, N435);
nor NOR2 (N441, N430, N94);
buf BUF1 (N442, N440);
nor NOR3 (N443, N441, N322, N442);
nand NAND2 (N444, N331, N148);
nor NOR2 (N445, N423, N412);
buf BUF1 (N446, N439);
or OR2 (N447, N438, N171);
and AND4 (N448, N433, N264, N321, N71);
not NOT1 (N449, N437);
buf BUF1 (N450, N443);
and AND2 (N451, N445, N212);
nand NAND4 (N452, N446, N364, N287, N385);
or OR2 (N453, N451, N299);
nor NOR3 (N454, N415, N317, N268);
nor NOR4 (N455, N450, N255, N288, N177);
xor XOR2 (N456, N432, N364);
or OR3 (N457, N449, N56, N154);
nand NAND3 (N458, N448, N379, N188);
nor NOR3 (N459, N427, N294, N13);
nor NOR2 (N460, N444, N110);
not NOT1 (N461, N459);
xor XOR2 (N462, N457, N277);
buf BUF1 (N463, N456);
or OR2 (N464, N453, N439);
nor NOR2 (N465, N461, N127);
and AND2 (N466, N452, N269);
or OR2 (N467, N447, N279);
buf BUF1 (N468, N466);
not NOT1 (N469, N460);
buf BUF1 (N470, N469);
buf BUF1 (N471, N465);
xor XOR2 (N472, N464, N114);
or OR3 (N473, N454, N101, N85);
and AND3 (N474, N463, N118, N25);
nand NAND4 (N475, N462, N5, N215, N180);
or OR3 (N476, N472, N81, N297);
xor XOR2 (N477, N468, N411);
and AND2 (N478, N455, N449);
buf BUF1 (N479, N458);
nor NOR2 (N480, N470, N8);
not NOT1 (N481, N473);
not NOT1 (N482, N474);
nand NAND3 (N483, N480, N470, N213);
xor XOR2 (N484, N471, N282);
nand NAND2 (N485, N479, N466);
or OR4 (N486, N481, N468, N11, N120);
not NOT1 (N487, N476);
nand NAND4 (N488, N477, N4, N250, N58);
nand NAND4 (N489, N467, N127, N435, N290);
or OR4 (N490, N489, N241, N422, N268);
or OR2 (N491, N484, N321);
and AND2 (N492, N486, N215);
nor NOR3 (N493, N491, N256, N216);
xor XOR2 (N494, N488, N431);
not NOT1 (N495, N494);
nand NAND3 (N496, N490, N231, N345);
and AND4 (N497, N485, N443, N332, N432);
nor NOR4 (N498, N493, N11, N485, N268);
buf BUF1 (N499, N492);
xor XOR2 (N500, N497, N186);
not NOT1 (N501, N483);
and AND3 (N502, N482, N72, N458);
xor XOR2 (N503, N500, N278);
xor XOR2 (N504, N499, N401);
xor XOR2 (N505, N503, N448);
not NOT1 (N506, N502);
buf BUF1 (N507, N504);
buf BUF1 (N508, N478);
buf BUF1 (N509, N505);
nand NAND3 (N510, N507, N377, N216);
nor NOR3 (N511, N475, N104, N476);
nor NOR4 (N512, N511, N269, N454, N467);
or OR2 (N513, N495, N322);
or OR3 (N514, N501, N271, N167);
nor NOR2 (N515, N513, N242);
or OR3 (N516, N498, N392, N513);
not NOT1 (N517, N487);
xor XOR2 (N518, N514, N89);
not NOT1 (N519, N518);
xor XOR2 (N520, N508, N57);
nor NOR3 (N521, N506, N330, N313);
nand NAND2 (N522, N519, N209);
xor XOR2 (N523, N512, N68);
buf BUF1 (N524, N517);
and AND2 (N525, N523, N470);
nand NAND3 (N526, N509, N278, N128);
xor XOR2 (N527, N510, N507);
buf BUF1 (N528, N521);
nor NOR3 (N529, N527, N279, N5);
nor NOR2 (N530, N525, N324);
and AND2 (N531, N516, N76);
nor NOR4 (N532, N530, N66, N73, N178);
buf BUF1 (N533, N515);
not NOT1 (N534, N528);
nand NAND3 (N535, N533, N242, N479);
nor NOR2 (N536, N522, N89);
nand NAND2 (N537, N529, N491);
and AND4 (N538, N537, N408, N371, N41);
nand NAND2 (N539, N496, N50);
or OR2 (N540, N536, N472);
buf BUF1 (N541, N520);
xor XOR2 (N542, N524, N172);
buf BUF1 (N543, N535);
nand NAND2 (N544, N540, N56);
and AND4 (N545, N544, N16, N335, N227);
buf BUF1 (N546, N545);
not NOT1 (N547, N534);
or OR4 (N548, N546, N294, N281, N420);
not NOT1 (N549, N538);
nand NAND2 (N550, N532, N277);
or OR4 (N551, N531, N375, N190, N528);
nand NAND3 (N552, N539, N550, N176);
or OR4 (N553, N520, N451, N264, N505);
and AND4 (N554, N551, N225, N94, N125);
nor NOR4 (N555, N547, N95, N271, N315);
and AND2 (N556, N552, N345);
and AND3 (N557, N541, N81, N70);
not NOT1 (N558, N548);
buf BUF1 (N559, N543);
nand NAND4 (N560, N555, N244, N107, N558);
or OR2 (N561, N322, N381);
buf BUF1 (N562, N553);
and AND3 (N563, N542, N415, N416);
xor XOR2 (N564, N557, N246);
and AND4 (N565, N549, N127, N170, N371);
xor XOR2 (N566, N565, N352);
not NOT1 (N567, N556);
nand NAND4 (N568, N560, N162, N11, N291);
or OR2 (N569, N562, N30);
nor NOR4 (N570, N564, N182, N479, N282);
not NOT1 (N571, N570);
and AND3 (N572, N526, N190, N508);
and AND4 (N573, N572, N326, N509, N501);
or OR4 (N574, N571, N218, N553, N31);
nor NOR2 (N575, N568, N21);
nor NOR3 (N576, N573, N393, N176);
nand NAND4 (N577, N561, N350, N260, N461);
buf BUF1 (N578, N559);
xor XOR2 (N579, N578, N332);
xor XOR2 (N580, N576, N31);
buf BUF1 (N581, N574);
not NOT1 (N582, N566);
nand NAND3 (N583, N582, N243, N87);
xor XOR2 (N584, N583, N144);
nand NAND3 (N585, N577, N532, N440);
not NOT1 (N586, N567);
not NOT1 (N587, N554);
nand NAND4 (N588, N563, N539, N264, N55);
buf BUF1 (N589, N587);
and AND2 (N590, N584, N96);
xor XOR2 (N591, N585, N418);
nor NOR3 (N592, N575, N110, N422);
or OR3 (N593, N569, N132, N307);
nor NOR2 (N594, N588, N550);
buf BUF1 (N595, N592);
and AND3 (N596, N594, N376, N550);
not NOT1 (N597, N591);
and AND4 (N598, N581, N183, N376, N60);
xor XOR2 (N599, N590, N227);
not NOT1 (N600, N599);
nor NOR3 (N601, N597, N146, N121);
and AND4 (N602, N586, N258, N160, N296);
nor NOR4 (N603, N593, N535, N89, N415);
not NOT1 (N604, N603);
nor NOR2 (N605, N598, N595);
and AND4 (N606, N477, N328, N157, N239);
or OR3 (N607, N604, N543, N274);
xor XOR2 (N608, N602, N520);
not NOT1 (N609, N601);
not NOT1 (N610, N600);
xor XOR2 (N611, N589, N255);
buf BUF1 (N612, N606);
nor NOR3 (N613, N607, N206, N611);
or OR2 (N614, N538, N1);
or OR3 (N615, N605, N541, N561);
xor XOR2 (N616, N610, N309);
nand NAND2 (N617, N612, N29);
nand NAND2 (N618, N579, N6);
not NOT1 (N619, N580);
nor NOR2 (N620, N608, N541);
and AND2 (N621, N616, N212);
not NOT1 (N622, N617);
and AND3 (N623, N619, N4, N204);
not NOT1 (N624, N614);
buf BUF1 (N625, N623);
and AND4 (N626, N609, N391, N265, N609);
not NOT1 (N627, N625);
buf BUF1 (N628, N620);
xor XOR2 (N629, N613, N71);
and AND4 (N630, N627, N339, N24, N364);
nand NAND4 (N631, N615, N258, N99, N393);
xor XOR2 (N632, N618, N494);
xor XOR2 (N633, N631, N259);
buf BUF1 (N634, N621);
not NOT1 (N635, N628);
not NOT1 (N636, N622);
xor XOR2 (N637, N632, N418);
buf BUF1 (N638, N629);
not NOT1 (N639, N630);
xor XOR2 (N640, N634, N631);
not NOT1 (N641, N596);
xor XOR2 (N642, N624, N451);
buf BUF1 (N643, N635);
buf BUF1 (N644, N639);
or OR4 (N645, N633, N552, N416, N440);
not NOT1 (N646, N644);
not NOT1 (N647, N643);
xor XOR2 (N648, N637, N207);
nor NOR3 (N649, N646, N169, N521);
nand NAND2 (N650, N647, N587);
or OR2 (N651, N642, N158);
not NOT1 (N652, N641);
and AND4 (N653, N648, N382, N531, N488);
xor XOR2 (N654, N636, N300);
nor NOR2 (N655, N650, N8);
or OR4 (N656, N638, N378, N472, N290);
nor NOR3 (N657, N645, N169, N164);
nand NAND3 (N658, N655, N604, N32);
buf BUF1 (N659, N626);
not NOT1 (N660, N653);
xor XOR2 (N661, N652, N47);
buf BUF1 (N662, N660);
nand NAND2 (N663, N661, N220);
buf BUF1 (N664, N654);
and AND2 (N665, N640, N580);
not NOT1 (N666, N662);
buf BUF1 (N667, N658);
and AND3 (N668, N656, N161, N199);
or OR3 (N669, N664, N215, N208);
xor XOR2 (N670, N665, N531);
nor NOR4 (N671, N659, N518, N338, N74);
or OR3 (N672, N670, N67, N544);
xor XOR2 (N673, N669, N98);
buf BUF1 (N674, N651);
nor NOR4 (N675, N671, N373, N71, N146);
not NOT1 (N676, N649);
or OR4 (N677, N675, N591, N334, N662);
xor XOR2 (N678, N666, N103);
or OR4 (N679, N667, N71, N492, N438);
or OR2 (N680, N674, N88);
nand NAND3 (N681, N680, N529, N40);
buf BUF1 (N682, N673);
nand NAND2 (N683, N663, N96);
buf BUF1 (N684, N683);
not NOT1 (N685, N677);
and AND4 (N686, N657, N551, N372, N292);
not NOT1 (N687, N679);
nand NAND4 (N688, N686, N275, N464, N229);
buf BUF1 (N689, N684);
nor NOR3 (N690, N687, N231, N109);
not NOT1 (N691, N676);
or OR2 (N692, N690, N446);
buf BUF1 (N693, N689);
nor NOR3 (N694, N693, N636, N373);
xor XOR2 (N695, N692, N507);
not NOT1 (N696, N685);
not NOT1 (N697, N696);
buf BUF1 (N698, N668);
nor NOR2 (N699, N691, N9);
and AND2 (N700, N682, N39);
xor XOR2 (N701, N695, N442);
nor NOR2 (N702, N700, N224);
and AND2 (N703, N698, N513);
buf BUF1 (N704, N672);
nand NAND4 (N705, N702, N637, N538, N470);
and AND4 (N706, N699, N337, N278, N156);
and AND3 (N707, N706, N644, N489);
xor XOR2 (N708, N703, N34);
and AND2 (N709, N697, N412);
xor XOR2 (N710, N708, N500);
nand NAND2 (N711, N678, N565);
xor XOR2 (N712, N701, N554);
and AND2 (N713, N694, N296);
buf BUF1 (N714, N712);
or OR2 (N715, N713, N211);
nor NOR4 (N716, N715, N44, N346, N120);
buf BUF1 (N717, N704);
nor NOR4 (N718, N707, N61, N160, N385);
and AND3 (N719, N681, N671, N173);
and AND4 (N720, N714, N341, N350, N293);
not NOT1 (N721, N719);
nor NOR2 (N722, N716, N540);
not NOT1 (N723, N710);
nand NAND3 (N724, N722, N614, N346);
xor XOR2 (N725, N724, N108);
buf BUF1 (N726, N688);
nand NAND4 (N727, N721, N660, N343, N299);
xor XOR2 (N728, N717, N365);
not NOT1 (N729, N720);
xor XOR2 (N730, N723, N133);
buf BUF1 (N731, N729);
xor XOR2 (N732, N725, N604);
nand NAND3 (N733, N711, N27, N202);
nand NAND4 (N734, N718, N572, N355, N682);
and AND4 (N735, N732, N452, N352, N178);
or OR4 (N736, N709, N642, N204, N607);
nand NAND2 (N737, N727, N516);
nand NAND4 (N738, N734, N12, N494, N69);
not NOT1 (N739, N736);
xor XOR2 (N740, N735, N12);
buf BUF1 (N741, N733);
or OR4 (N742, N726, N463, N682, N626);
xor XOR2 (N743, N739, N718);
or OR2 (N744, N730, N34);
or OR2 (N745, N731, N548);
xor XOR2 (N746, N741, N294);
not NOT1 (N747, N746);
nor NOR4 (N748, N705, N261, N8, N597);
nor NOR4 (N749, N744, N600, N737, N2);
or OR4 (N750, N115, N594, N732, N709);
nor NOR4 (N751, N738, N651, N447, N374);
or OR4 (N752, N747, N110, N254, N119);
buf BUF1 (N753, N752);
xor XOR2 (N754, N745, N356);
and AND4 (N755, N751, N629, N727, N278);
nor NOR3 (N756, N750, N593, N754);
xor XOR2 (N757, N171, N220);
nand NAND3 (N758, N748, N303, N505);
not NOT1 (N759, N740);
nand NAND3 (N760, N743, N539, N652);
not NOT1 (N761, N756);
xor XOR2 (N762, N760, N480);
not NOT1 (N763, N753);
buf BUF1 (N764, N728);
not NOT1 (N765, N759);
xor XOR2 (N766, N762, N424);
nand NAND2 (N767, N755, N699);
buf BUF1 (N768, N767);
nand NAND4 (N769, N764, N498, N102, N724);
not NOT1 (N770, N749);
buf BUF1 (N771, N765);
nand NAND3 (N772, N769, N53, N674);
buf BUF1 (N773, N766);
and AND4 (N774, N763, N241, N650, N122);
buf BUF1 (N775, N758);
nand NAND4 (N776, N757, N771, N96, N161);
or OR4 (N777, N316, N376, N291, N439);
nor NOR3 (N778, N768, N319, N5);
nor NOR2 (N779, N761, N733);
and AND2 (N780, N779, N149);
buf BUF1 (N781, N742);
nor NOR4 (N782, N778, N66, N598, N669);
or OR2 (N783, N781, N545);
buf BUF1 (N784, N780);
or OR2 (N785, N773, N256);
and AND3 (N786, N770, N689, N202);
buf BUF1 (N787, N776);
or OR4 (N788, N783, N439, N424, N489);
and AND2 (N789, N786, N561);
buf BUF1 (N790, N788);
buf BUF1 (N791, N775);
not NOT1 (N792, N789);
buf BUF1 (N793, N782);
xor XOR2 (N794, N772, N748);
nand NAND4 (N795, N784, N382, N139, N424);
xor XOR2 (N796, N787, N623);
nand NAND3 (N797, N774, N431, N302);
and AND2 (N798, N785, N315);
and AND3 (N799, N794, N152, N353);
xor XOR2 (N800, N777, N523);
not NOT1 (N801, N792);
and AND3 (N802, N797, N505, N316);
xor XOR2 (N803, N796, N119);
and AND2 (N804, N790, N548);
or OR3 (N805, N795, N632, N520);
nor NOR4 (N806, N805, N338, N610, N111);
or OR3 (N807, N804, N165, N614);
or OR3 (N808, N799, N215, N5);
buf BUF1 (N809, N791);
xor XOR2 (N810, N800, N206);
and AND2 (N811, N802, N716);
nor NOR4 (N812, N793, N589, N207, N124);
nand NAND2 (N813, N798, N552);
nor NOR3 (N814, N813, N224, N203);
or OR3 (N815, N809, N617, N319);
or OR4 (N816, N801, N53, N779, N138);
or OR4 (N817, N810, N473, N130, N678);
nand NAND2 (N818, N806, N725);
xor XOR2 (N819, N803, N776);
or OR2 (N820, N807, N636);
not NOT1 (N821, N814);
and AND4 (N822, N820, N99, N245, N127);
buf BUF1 (N823, N812);
not NOT1 (N824, N817);
and AND2 (N825, N815, N698);
or OR3 (N826, N816, N557, N133);
nor NOR3 (N827, N825, N331, N443);
or OR2 (N828, N819, N575);
not NOT1 (N829, N808);
not NOT1 (N830, N829);
buf BUF1 (N831, N824);
nor NOR2 (N832, N821, N691);
or OR2 (N833, N832, N753);
xor XOR2 (N834, N830, N471);
nor NOR3 (N835, N822, N129, N595);
nand NAND2 (N836, N827, N588);
not NOT1 (N837, N823);
nand NAND2 (N838, N831, N728);
xor XOR2 (N839, N834, N84);
nor NOR2 (N840, N826, N644);
nor NOR2 (N841, N836, N285);
or OR3 (N842, N841, N490, N20);
nor NOR4 (N843, N811, N464, N711, N816);
nand NAND2 (N844, N840, N437);
buf BUF1 (N845, N835);
buf BUF1 (N846, N838);
or OR4 (N847, N846, N318, N295, N259);
or OR2 (N848, N843, N128);
buf BUF1 (N849, N845);
and AND2 (N850, N837, N521);
and AND2 (N851, N850, N721);
nor NOR4 (N852, N848, N176, N594, N621);
not NOT1 (N853, N818);
nor NOR2 (N854, N851, N216);
buf BUF1 (N855, N842);
xor XOR2 (N856, N828, N772);
xor XOR2 (N857, N855, N91);
nor NOR2 (N858, N853, N658);
not NOT1 (N859, N852);
nand NAND2 (N860, N856, N337);
not NOT1 (N861, N847);
and AND2 (N862, N833, N474);
or OR3 (N863, N844, N585, N567);
not NOT1 (N864, N862);
nor NOR2 (N865, N839, N344);
buf BUF1 (N866, N865);
or OR3 (N867, N863, N657, N98);
not NOT1 (N868, N857);
buf BUF1 (N869, N858);
not NOT1 (N870, N861);
not NOT1 (N871, N860);
not NOT1 (N872, N859);
nand NAND3 (N873, N854, N616, N89);
nor NOR2 (N874, N868, N241);
not NOT1 (N875, N873);
nor NOR3 (N876, N870, N51, N119);
xor XOR2 (N877, N871, N742);
nand NAND4 (N878, N875, N145, N126, N676);
buf BUF1 (N879, N866);
or OR2 (N880, N849, N425);
and AND4 (N881, N872, N680, N63, N94);
xor XOR2 (N882, N878, N227);
or OR4 (N883, N864, N763, N618, N664);
buf BUF1 (N884, N879);
xor XOR2 (N885, N877, N720);
buf BUF1 (N886, N885);
buf BUF1 (N887, N867);
nand NAND2 (N888, N884, N119);
nor NOR2 (N889, N876, N599);
not NOT1 (N890, N882);
not NOT1 (N891, N880);
not NOT1 (N892, N888);
nor NOR2 (N893, N883, N783);
xor XOR2 (N894, N893, N586);
nor NOR4 (N895, N869, N415, N209, N152);
or OR2 (N896, N881, N747);
buf BUF1 (N897, N889);
buf BUF1 (N898, N891);
nand NAND2 (N899, N887, N97);
xor XOR2 (N900, N895, N393);
nand NAND3 (N901, N874, N67, N757);
nor NOR2 (N902, N899, N94);
xor XOR2 (N903, N896, N711);
nor NOR2 (N904, N886, N536);
not NOT1 (N905, N904);
nand NAND2 (N906, N901, N122);
or OR2 (N907, N900, N117);
nor NOR2 (N908, N903, N425);
nand NAND3 (N909, N908, N547, N483);
and AND2 (N910, N906, N758);
and AND2 (N911, N897, N537);
xor XOR2 (N912, N892, N330);
or OR2 (N913, N909, N758);
nor NOR2 (N914, N898, N551);
or OR4 (N915, N907, N465, N745, N701);
and AND3 (N916, N894, N665, N240);
and AND4 (N917, N913, N153, N901, N73);
nor NOR4 (N918, N915, N747, N65, N603);
or OR2 (N919, N916, N163);
and AND3 (N920, N919, N737, N72);
not NOT1 (N921, N902);
nor NOR4 (N922, N921, N255, N677, N810);
not NOT1 (N923, N917);
or OR3 (N924, N918, N685, N502);
and AND2 (N925, N923, N322);
or OR3 (N926, N905, N26, N925);
not NOT1 (N927, N768);
xor XOR2 (N928, N922, N231);
not NOT1 (N929, N910);
buf BUF1 (N930, N924);
not NOT1 (N931, N912);
or OR4 (N932, N930, N231, N397, N860);
and AND2 (N933, N920, N73);
or OR3 (N934, N933, N17, N692);
nor NOR3 (N935, N911, N490, N545);
xor XOR2 (N936, N928, N268);
nor NOR3 (N937, N932, N745, N711);
nand NAND2 (N938, N926, N479);
and AND3 (N939, N929, N826, N387);
nor NOR3 (N940, N914, N848, N512);
buf BUF1 (N941, N935);
not NOT1 (N942, N890);
not NOT1 (N943, N936);
nor NOR3 (N944, N939, N875, N535);
or OR2 (N945, N942, N447);
and AND4 (N946, N943, N625, N854, N195);
buf BUF1 (N947, N938);
buf BUF1 (N948, N944);
nor NOR2 (N949, N941, N878);
buf BUF1 (N950, N947);
buf BUF1 (N951, N940);
xor XOR2 (N952, N950, N189);
nand NAND4 (N953, N945, N857, N6, N793);
not NOT1 (N954, N952);
and AND2 (N955, N927, N240);
nor NOR4 (N956, N953, N566, N259, N297);
buf BUF1 (N957, N948);
not NOT1 (N958, N931);
and AND2 (N959, N956, N530);
and AND2 (N960, N959, N844);
buf BUF1 (N961, N949);
buf BUF1 (N962, N957);
not NOT1 (N963, N934);
nor NOR4 (N964, N962, N410, N956, N694);
buf BUF1 (N965, N937);
nand NAND4 (N966, N960, N854, N483, N55);
buf BUF1 (N967, N963);
nand NAND4 (N968, N951, N712, N952, N625);
nand NAND2 (N969, N955, N941);
xor XOR2 (N970, N966, N122);
nor NOR2 (N971, N968, N691);
xor XOR2 (N972, N961, N526);
nor NOR2 (N973, N967, N784);
not NOT1 (N974, N965);
or OR4 (N975, N958, N889, N50, N440);
or OR4 (N976, N972, N635, N839, N730);
and AND3 (N977, N946, N342, N508);
nor NOR2 (N978, N977, N332);
nand NAND4 (N979, N954, N868, N757, N700);
and AND3 (N980, N969, N92, N519);
and AND2 (N981, N974, N746);
nor NOR2 (N982, N976, N348);
xor XOR2 (N983, N964, N121);
or OR2 (N984, N970, N91);
or OR2 (N985, N973, N545);
nand NAND3 (N986, N979, N859, N846);
or OR3 (N987, N980, N638, N704);
and AND3 (N988, N987, N471, N298);
and AND2 (N989, N983, N234);
or OR2 (N990, N971, N568);
buf BUF1 (N991, N988);
not NOT1 (N992, N986);
xor XOR2 (N993, N981, N708);
nand NAND4 (N994, N978, N710, N52, N583);
not NOT1 (N995, N985);
not NOT1 (N996, N993);
not NOT1 (N997, N992);
nor NOR2 (N998, N990, N592);
or OR3 (N999, N995, N425, N169);
buf BUF1 (N1000, N984);
nor NOR3 (N1001, N999, N576, N788);
or OR3 (N1002, N982, N190, N863);
and AND2 (N1003, N998, N361);
and AND4 (N1004, N994, N344, N20, N977);
xor XOR2 (N1005, N975, N672);
nand NAND3 (N1006, N997, N904, N307);
nor NOR2 (N1007, N996, N263);
nand NAND3 (N1008, N1007, N11, N867);
xor XOR2 (N1009, N1006, N543);
nor NOR2 (N1010, N989, N437);
not NOT1 (N1011, N1010);
buf BUF1 (N1012, N1005);
nand NAND3 (N1013, N1009, N593, N8);
and AND3 (N1014, N1002, N86, N430);
and AND2 (N1015, N1012, N483);
nand NAND2 (N1016, N1004, N853);
buf BUF1 (N1017, N1014);
nand NAND2 (N1018, N991, N113);
and AND3 (N1019, N1016, N341, N100);
nor NOR4 (N1020, N1011, N903, N93, N605);
nor NOR4 (N1021, N1017, N175, N606, N872);
not NOT1 (N1022, N1008);
and AND4 (N1023, N1015, N707, N701, N781);
or OR4 (N1024, N1023, N915, N800, N465);
or OR4 (N1025, N1020, N384, N192, N550);
xor XOR2 (N1026, N1022, N347);
buf BUF1 (N1027, N1021);
xor XOR2 (N1028, N1026, N1012);
or OR2 (N1029, N1025, N812);
or OR4 (N1030, N1001, N1000, N730, N1015);
nor NOR2 (N1031, N687, N90);
nor NOR2 (N1032, N1018, N470);
not NOT1 (N1033, N1024);
and AND2 (N1034, N1033, N799);
not NOT1 (N1035, N1029);
not NOT1 (N1036, N1032);
nor NOR3 (N1037, N1019, N96, N720);
or OR2 (N1038, N1037, N61);
nand NAND3 (N1039, N1003, N1009, N1009);
xor XOR2 (N1040, N1038, N762);
and AND2 (N1041, N1040, N306);
nor NOR2 (N1042, N1027, N507);
nor NOR4 (N1043, N1030, N615, N211, N29);
and AND2 (N1044, N1034, N338);
nor NOR2 (N1045, N1041, N464);
buf BUF1 (N1046, N1013);
not NOT1 (N1047, N1035);
and AND2 (N1048, N1031, N91);
and AND3 (N1049, N1028, N267, N931);
not NOT1 (N1050, N1045);
or OR3 (N1051, N1044, N393, N361);
not NOT1 (N1052, N1050);
or OR2 (N1053, N1046, N170);
nor NOR3 (N1054, N1052, N234, N24);
nor NOR4 (N1055, N1049, N845, N554, N998);
and AND3 (N1056, N1051, N649, N193);
and AND3 (N1057, N1056, N204, N280);
xor XOR2 (N1058, N1053, N979);
or OR3 (N1059, N1057, N86, N665);
nor NOR2 (N1060, N1054, N393);
xor XOR2 (N1061, N1039, N94);
buf BUF1 (N1062, N1042);
buf BUF1 (N1063, N1048);
and AND3 (N1064, N1062, N990, N195);
not NOT1 (N1065, N1059);
buf BUF1 (N1066, N1061);
and AND2 (N1067, N1047, N889);
xor XOR2 (N1068, N1065, N64);
buf BUF1 (N1069, N1055);
and AND3 (N1070, N1068, N255, N748);
or OR4 (N1071, N1058, N20, N473, N695);
nor NOR4 (N1072, N1069, N698, N843, N631);
not NOT1 (N1073, N1071);
not NOT1 (N1074, N1073);
xor XOR2 (N1075, N1063, N832);
nor NOR3 (N1076, N1066, N925, N147);
not NOT1 (N1077, N1075);
nor NOR3 (N1078, N1067, N804, N1037);
nor NOR3 (N1079, N1064, N519, N953);
buf BUF1 (N1080, N1079);
or OR2 (N1081, N1060, N394);
nor NOR4 (N1082, N1076, N78, N503, N376);
and AND2 (N1083, N1081, N398);
not NOT1 (N1084, N1070);
not NOT1 (N1085, N1078);
nor NOR2 (N1086, N1036, N350);
not NOT1 (N1087, N1074);
not NOT1 (N1088, N1072);
and AND2 (N1089, N1088, N358);
not NOT1 (N1090, N1089);
nand NAND2 (N1091, N1077, N786);
nand NAND3 (N1092, N1083, N645, N669);
not NOT1 (N1093, N1082);
and AND4 (N1094, N1085, N271, N951, N170);
xor XOR2 (N1095, N1093, N594);
nand NAND2 (N1096, N1084, N16);
buf BUF1 (N1097, N1090);
nor NOR3 (N1098, N1091, N706, N1028);
and AND4 (N1099, N1095, N63, N366, N575);
buf BUF1 (N1100, N1094);
nand NAND4 (N1101, N1096, N316, N918, N52);
or OR2 (N1102, N1101, N978);
xor XOR2 (N1103, N1080, N63);
or OR3 (N1104, N1100, N865, N144);
or OR4 (N1105, N1103, N941, N339, N971);
xor XOR2 (N1106, N1087, N906);
buf BUF1 (N1107, N1104);
nor NOR2 (N1108, N1106, N725);
nor NOR2 (N1109, N1107, N488);
not NOT1 (N1110, N1105);
xor XOR2 (N1111, N1098, N788);
nor NOR4 (N1112, N1108, N53, N742, N92);
xor XOR2 (N1113, N1110, N799);
not NOT1 (N1114, N1092);
buf BUF1 (N1115, N1109);
xor XOR2 (N1116, N1112, N646);
nand NAND3 (N1117, N1099, N431, N476);
nor NOR3 (N1118, N1116, N336, N63);
nor NOR4 (N1119, N1043, N275, N337, N659);
and AND2 (N1120, N1111, N629);
buf BUF1 (N1121, N1117);
buf BUF1 (N1122, N1119);
buf BUF1 (N1123, N1122);
or OR4 (N1124, N1114, N204, N1118, N248);
nor NOR4 (N1125, N190, N688, N331, N276);
nand NAND3 (N1126, N1123, N62, N195);
or OR2 (N1127, N1124, N22);
and AND4 (N1128, N1086, N318, N695, N530);
nand NAND2 (N1129, N1128, N1125);
not NOT1 (N1130, N335);
nand NAND3 (N1131, N1121, N176, N300);
and AND4 (N1132, N1130, N467, N322, N98);
or OR4 (N1133, N1127, N803, N709, N1102);
xor XOR2 (N1134, N155, N186);
or OR3 (N1135, N1132, N819, N691);
nand NAND3 (N1136, N1126, N14, N425);
nor NOR4 (N1137, N1134, N720, N155, N825);
xor XOR2 (N1138, N1129, N676);
buf BUF1 (N1139, N1097);
not NOT1 (N1140, N1137);
nand NAND2 (N1141, N1138, N1015);
and AND3 (N1142, N1135, N212, N680);
xor XOR2 (N1143, N1139, N187);
and AND3 (N1144, N1113, N653, N831);
xor XOR2 (N1145, N1133, N610);
nand NAND3 (N1146, N1140, N1124, N260);
or OR4 (N1147, N1141, N729, N767, N64);
buf BUF1 (N1148, N1145);
or OR2 (N1149, N1131, N813);
xor XOR2 (N1150, N1120, N100);
xor XOR2 (N1151, N1115, N813);
xor XOR2 (N1152, N1142, N578);
not NOT1 (N1153, N1151);
xor XOR2 (N1154, N1143, N761);
or OR3 (N1155, N1144, N572, N293);
not NOT1 (N1156, N1146);
xor XOR2 (N1157, N1150, N335);
and AND4 (N1158, N1149, N651, N776, N558);
nand NAND4 (N1159, N1147, N477, N1131, N601);
and AND4 (N1160, N1136, N197, N455, N620);
buf BUF1 (N1161, N1156);
nor NOR4 (N1162, N1161, N534, N549, N925);
and AND2 (N1163, N1153, N137);
nor NOR4 (N1164, N1160, N987, N751, N170);
and AND2 (N1165, N1158, N1034);
nor NOR3 (N1166, N1164, N971, N1106);
xor XOR2 (N1167, N1162, N827);
buf BUF1 (N1168, N1155);
nor NOR2 (N1169, N1165, N704);
xor XOR2 (N1170, N1167, N1135);
nor NOR2 (N1171, N1168, N768);
nand NAND2 (N1172, N1166, N46);
nand NAND4 (N1173, N1171, N331, N645, N192);
xor XOR2 (N1174, N1157, N835);
or OR3 (N1175, N1174, N292, N489);
buf BUF1 (N1176, N1170);
not NOT1 (N1177, N1173);
nor NOR4 (N1178, N1176, N550, N593, N734);
or OR2 (N1179, N1159, N741);
nand NAND4 (N1180, N1179, N859, N102, N692);
not NOT1 (N1181, N1178);
not NOT1 (N1182, N1181);
nor NOR4 (N1183, N1163, N663, N780, N182);
not NOT1 (N1184, N1148);
xor XOR2 (N1185, N1169, N264);
nand NAND3 (N1186, N1184, N1164, N819);
nor NOR4 (N1187, N1154, N426, N326, N130);
buf BUF1 (N1188, N1185);
nand NAND4 (N1189, N1175, N1079, N1050, N730);
or OR2 (N1190, N1172, N923);
not NOT1 (N1191, N1182);
nor NOR4 (N1192, N1189, N829, N1149, N903);
xor XOR2 (N1193, N1191, N997);
nor NOR4 (N1194, N1192, N380, N1187, N1078);
not NOT1 (N1195, N71);
and AND2 (N1196, N1183, N261);
and AND4 (N1197, N1188, N643, N448, N337);
xor XOR2 (N1198, N1177, N599);
buf BUF1 (N1199, N1198);
buf BUF1 (N1200, N1197);
not NOT1 (N1201, N1195);
nor NOR3 (N1202, N1180, N532, N535);
buf BUF1 (N1203, N1186);
buf BUF1 (N1204, N1152);
and AND4 (N1205, N1193, N736, N144, N718);
or OR3 (N1206, N1200, N996, N1183);
and AND3 (N1207, N1204, N250, N984);
nor NOR2 (N1208, N1199, N414);
nand NAND2 (N1209, N1207, N167);
nand NAND2 (N1210, N1201, N1118);
not NOT1 (N1211, N1196);
nor NOR2 (N1212, N1205, N542);
buf BUF1 (N1213, N1203);
nor NOR4 (N1214, N1206, N34, N802, N312);
and AND4 (N1215, N1194, N764, N452, N1132);
and AND4 (N1216, N1212, N1062, N895, N1143);
nor NOR2 (N1217, N1215, N57);
nand NAND3 (N1218, N1190, N554, N504);
nor NOR4 (N1219, N1218, N496, N410, N593);
or OR2 (N1220, N1209, N1101);
or OR2 (N1221, N1219, N670);
buf BUF1 (N1222, N1220);
nand NAND3 (N1223, N1211, N898, N462);
nand NAND3 (N1224, N1223, N453, N1216);
not NOT1 (N1225, N1022);
buf BUF1 (N1226, N1210);
buf BUF1 (N1227, N1221);
and AND4 (N1228, N1226, N780, N584, N955);
nand NAND2 (N1229, N1214, N882);
not NOT1 (N1230, N1228);
not NOT1 (N1231, N1213);
nand NAND4 (N1232, N1231, N773, N507, N297);
xor XOR2 (N1233, N1202, N1174);
nand NAND2 (N1234, N1217, N716);
xor XOR2 (N1235, N1233, N994);
and AND2 (N1236, N1222, N968);
not NOT1 (N1237, N1230);
or OR4 (N1238, N1229, N92, N711, N1099);
buf BUF1 (N1239, N1232);
nor NOR2 (N1240, N1237, N881);
not NOT1 (N1241, N1238);
or OR3 (N1242, N1239, N167, N910);
nand NAND2 (N1243, N1240, N996);
nor NOR3 (N1244, N1235, N1158, N1228);
nand NAND2 (N1245, N1227, N485);
buf BUF1 (N1246, N1242);
buf BUF1 (N1247, N1225);
or OR4 (N1248, N1224, N895, N582, N772);
nor NOR3 (N1249, N1248, N224, N247);
xor XOR2 (N1250, N1208, N1101);
or OR3 (N1251, N1234, N313, N754);
not NOT1 (N1252, N1250);
buf BUF1 (N1253, N1247);
nor NOR4 (N1254, N1249, N3, N244, N1001);
and AND3 (N1255, N1251, N966, N204);
or OR4 (N1256, N1252, N445, N990, N1251);
nor NOR3 (N1257, N1243, N437, N322);
or OR4 (N1258, N1255, N1105, N807, N178);
xor XOR2 (N1259, N1245, N132);
or OR2 (N1260, N1236, N547);
and AND4 (N1261, N1257, N353, N1208, N577);
and AND4 (N1262, N1260, N1099, N316, N1049);
xor XOR2 (N1263, N1258, N857);
nor NOR3 (N1264, N1241, N1159, N856);
or OR4 (N1265, N1253, N476, N1251, N298);
and AND2 (N1266, N1256, N550);
nor NOR2 (N1267, N1259, N35);
nand NAND3 (N1268, N1266, N750, N423);
and AND2 (N1269, N1246, N529);
and AND4 (N1270, N1262, N293, N267, N2);
nand NAND2 (N1271, N1261, N259);
nand NAND4 (N1272, N1270, N964, N923, N866);
or OR3 (N1273, N1265, N248, N1256);
nor NOR4 (N1274, N1272, N681, N591, N673);
and AND4 (N1275, N1263, N670, N595, N203);
nor NOR4 (N1276, N1244, N580, N947, N446);
xor XOR2 (N1277, N1276, N242);
not NOT1 (N1278, N1268);
not NOT1 (N1279, N1273);
not NOT1 (N1280, N1264);
nor NOR2 (N1281, N1274, N1081);
nor NOR2 (N1282, N1277, N915);
or OR3 (N1283, N1271, N892, N1163);
buf BUF1 (N1284, N1280);
and AND3 (N1285, N1254, N757, N121);
and AND2 (N1286, N1279, N1175);
nor NOR3 (N1287, N1275, N20, N497);
or OR3 (N1288, N1286, N315, N1090);
not NOT1 (N1289, N1278);
not NOT1 (N1290, N1267);
and AND2 (N1291, N1290, N816);
nand NAND2 (N1292, N1281, N190);
buf BUF1 (N1293, N1292);
and AND2 (N1294, N1293, N259);
and AND3 (N1295, N1283, N690, N724);
xor XOR2 (N1296, N1295, N723);
and AND4 (N1297, N1288, N1145, N325, N233);
nand NAND4 (N1298, N1284, N529, N1149, N635);
nor NOR4 (N1299, N1298, N234, N673, N32);
nor NOR2 (N1300, N1287, N908);
buf BUF1 (N1301, N1285);
not NOT1 (N1302, N1301);
not NOT1 (N1303, N1282);
nor NOR4 (N1304, N1269, N1280, N50, N822);
not NOT1 (N1305, N1303);
buf BUF1 (N1306, N1302);
or OR3 (N1307, N1305, N123, N638);
not NOT1 (N1308, N1294);
buf BUF1 (N1309, N1307);
nand NAND4 (N1310, N1299, N1039, N948, N74);
or OR2 (N1311, N1304, N737);
nand NAND2 (N1312, N1291, N406);
nor NOR4 (N1313, N1309, N1181, N184, N445);
not NOT1 (N1314, N1312);
buf BUF1 (N1315, N1306);
and AND2 (N1316, N1315, N966);
nor NOR4 (N1317, N1308, N119, N210, N1022);
nor NOR3 (N1318, N1316, N486, N919);
not NOT1 (N1319, N1297);
and AND3 (N1320, N1311, N129, N436);
and AND2 (N1321, N1320, N543);
nor NOR4 (N1322, N1319, N532, N1010, N253);
and AND4 (N1323, N1318, N293, N1148, N172);
xor XOR2 (N1324, N1322, N812);
buf BUF1 (N1325, N1321);
xor XOR2 (N1326, N1310, N463);
buf BUF1 (N1327, N1289);
and AND2 (N1328, N1300, N801);
or OR4 (N1329, N1323, N85, N1296, N1176);
and AND3 (N1330, N586, N238, N833);
buf BUF1 (N1331, N1328);
or OR3 (N1332, N1327, N3, N283);
nor NOR4 (N1333, N1317, N137, N718, N958);
xor XOR2 (N1334, N1326, N757);
not NOT1 (N1335, N1334);
nand NAND4 (N1336, N1332, N851, N278, N1198);
nor NOR2 (N1337, N1325, N1035);
nand NAND2 (N1338, N1335, N295);
or OR3 (N1339, N1337, N1336, N1252);
or OR4 (N1340, N1071, N106, N504, N1005);
nand NAND2 (N1341, N1314, N299);
buf BUF1 (N1342, N1330);
buf BUF1 (N1343, N1331);
nor NOR4 (N1344, N1313, N792, N1253, N424);
buf BUF1 (N1345, N1324);
not NOT1 (N1346, N1342);
not NOT1 (N1347, N1343);
buf BUF1 (N1348, N1333);
nor NOR3 (N1349, N1341, N74, N160);
not NOT1 (N1350, N1349);
nor NOR4 (N1351, N1345, N525, N435, N302);
and AND3 (N1352, N1348, N962, N969);
xor XOR2 (N1353, N1340, N336);
and AND4 (N1354, N1339, N499, N35, N521);
and AND3 (N1355, N1351, N1069, N1064);
nor NOR2 (N1356, N1353, N688);
xor XOR2 (N1357, N1350, N1123);
not NOT1 (N1358, N1329);
and AND3 (N1359, N1347, N756, N1139);
not NOT1 (N1360, N1352);
nor NOR2 (N1361, N1355, N1088);
nor NOR2 (N1362, N1354, N147);
buf BUF1 (N1363, N1344);
buf BUF1 (N1364, N1363);
xor XOR2 (N1365, N1361, N143);
and AND2 (N1366, N1364, N153);
and AND3 (N1367, N1358, N935, N721);
xor XOR2 (N1368, N1367, N811);
nor NOR4 (N1369, N1346, N91, N707, N1249);
xor XOR2 (N1370, N1360, N292);
nand NAND3 (N1371, N1357, N272, N376);
nand NAND3 (N1372, N1359, N1092, N718);
xor XOR2 (N1373, N1338, N288);
nor NOR2 (N1374, N1373, N215);
xor XOR2 (N1375, N1362, N1350);
not NOT1 (N1376, N1370);
xor XOR2 (N1377, N1376, N24);
not NOT1 (N1378, N1371);
not NOT1 (N1379, N1372);
or OR2 (N1380, N1369, N764);
not NOT1 (N1381, N1379);
xor XOR2 (N1382, N1381, N230);
xor XOR2 (N1383, N1378, N561);
xor XOR2 (N1384, N1356, N1108);
and AND2 (N1385, N1375, N587);
buf BUF1 (N1386, N1374);
xor XOR2 (N1387, N1383, N236);
xor XOR2 (N1388, N1384, N1106);
buf BUF1 (N1389, N1386);
not NOT1 (N1390, N1366);
nand NAND2 (N1391, N1380, N376);
and AND2 (N1392, N1387, N560);
not NOT1 (N1393, N1368);
and AND2 (N1394, N1393, N764);
and AND4 (N1395, N1365, N472, N745, N1116);
buf BUF1 (N1396, N1388);
and AND3 (N1397, N1389, N688, N8);
not NOT1 (N1398, N1382);
and AND4 (N1399, N1392, N1215, N164, N1080);
buf BUF1 (N1400, N1395);
and AND4 (N1401, N1397, N169, N1147, N787);
not NOT1 (N1402, N1390);
or OR3 (N1403, N1402, N695, N373);
xor XOR2 (N1404, N1399, N889);
and AND2 (N1405, N1400, N676);
and AND3 (N1406, N1391, N1401, N803);
nor NOR2 (N1407, N1306, N208);
not NOT1 (N1408, N1406);
and AND2 (N1409, N1385, N962);
buf BUF1 (N1410, N1409);
buf BUF1 (N1411, N1403);
and AND2 (N1412, N1408, N387);
nor NOR3 (N1413, N1407, N559, N155);
and AND2 (N1414, N1411, N237);
buf BUF1 (N1415, N1377);
and AND4 (N1416, N1404, N497, N1179, N699);
or OR4 (N1417, N1416, N354, N719, N878);
and AND2 (N1418, N1394, N485);
xor XOR2 (N1419, N1398, N427);
or OR2 (N1420, N1412, N909);
xor XOR2 (N1421, N1405, N475);
buf BUF1 (N1422, N1420);
or OR2 (N1423, N1417, N551);
and AND2 (N1424, N1414, N661);
nand NAND3 (N1425, N1413, N970, N536);
nand NAND3 (N1426, N1419, N1188, N751);
nand NAND3 (N1427, N1424, N1071, N797);
nor NOR4 (N1428, N1410, N499, N1139, N727);
buf BUF1 (N1429, N1418);
or OR3 (N1430, N1428, N316, N1149);
buf BUF1 (N1431, N1396);
buf BUF1 (N1432, N1430);
nand NAND2 (N1433, N1423, N1156);
xor XOR2 (N1434, N1432, N1192);
buf BUF1 (N1435, N1415);
and AND4 (N1436, N1434, N1118, N910, N659);
and AND4 (N1437, N1426, N94, N875, N704);
nand NAND3 (N1438, N1437, N562, N159);
or OR4 (N1439, N1431, N221, N8, N90);
and AND2 (N1440, N1435, N54);
nand NAND4 (N1441, N1439, N591, N622, N794);
or OR3 (N1442, N1433, N1295, N222);
buf BUF1 (N1443, N1438);
nor NOR3 (N1444, N1422, N646, N840);
buf BUF1 (N1445, N1429);
xor XOR2 (N1446, N1444, N1011);
and AND3 (N1447, N1445, N870, N950);
not NOT1 (N1448, N1421);
nand NAND3 (N1449, N1441, N1413, N726);
xor XOR2 (N1450, N1447, N1341);
nor NOR2 (N1451, N1440, N864);
or OR2 (N1452, N1449, N888);
buf BUF1 (N1453, N1427);
not NOT1 (N1454, N1451);
or OR3 (N1455, N1452, N1413, N529);
xor XOR2 (N1456, N1455, N390);
buf BUF1 (N1457, N1450);
xor XOR2 (N1458, N1454, N175);
xor XOR2 (N1459, N1448, N1058);
nand NAND2 (N1460, N1457, N1432);
not NOT1 (N1461, N1456);
buf BUF1 (N1462, N1458);
not NOT1 (N1463, N1436);
not NOT1 (N1464, N1443);
nand NAND3 (N1465, N1463, N584, N980);
nor NOR3 (N1466, N1446, N629, N198);
and AND3 (N1467, N1453, N598, N1134);
xor XOR2 (N1468, N1459, N846);
nand NAND2 (N1469, N1465, N844);
or OR4 (N1470, N1460, N116, N1062, N598);
and AND4 (N1471, N1469, N500, N1238, N998);
buf BUF1 (N1472, N1425);
buf BUF1 (N1473, N1464);
and AND2 (N1474, N1470, N1420);
or OR4 (N1475, N1462, N336, N296, N801);
nor NOR3 (N1476, N1442, N879, N328);
and AND4 (N1477, N1471, N510, N192, N942);
nor NOR3 (N1478, N1468, N1351, N1443);
and AND3 (N1479, N1476, N1462, N1156);
and AND2 (N1480, N1473, N923);
nor NOR3 (N1481, N1461, N379, N439);
nor NOR4 (N1482, N1474, N1427, N263, N1312);
and AND2 (N1483, N1477, N1150);
and AND2 (N1484, N1467, N1206);
and AND3 (N1485, N1478, N562, N635);
nand NAND2 (N1486, N1472, N674);
nor NOR3 (N1487, N1479, N1167, N338);
and AND4 (N1488, N1482, N580, N703, N670);
nand NAND2 (N1489, N1481, N599);
or OR2 (N1490, N1483, N660);
buf BUF1 (N1491, N1486);
nand NAND2 (N1492, N1487, N833);
nor NOR4 (N1493, N1466, N1406, N313, N426);
or OR3 (N1494, N1484, N701, N1330);
buf BUF1 (N1495, N1490);
buf BUF1 (N1496, N1475);
not NOT1 (N1497, N1480);
nand NAND3 (N1498, N1494, N1073, N233);
xor XOR2 (N1499, N1491, N12);
nor NOR2 (N1500, N1488, N921);
not NOT1 (N1501, N1497);
and AND3 (N1502, N1489, N1115, N785);
or OR4 (N1503, N1502, N27, N1290, N1303);
and AND2 (N1504, N1498, N369);
nor NOR4 (N1505, N1493, N685, N554, N115);
nor NOR2 (N1506, N1503, N1041);
xor XOR2 (N1507, N1501, N1476);
and AND4 (N1508, N1492, N1080, N417, N631);
nor NOR2 (N1509, N1499, N108);
nand NAND3 (N1510, N1509, N386, N629);
nor NOR3 (N1511, N1507, N1242, N475);
and AND3 (N1512, N1500, N1319, N1238);
xor XOR2 (N1513, N1495, N522);
and AND3 (N1514, N1504, N79, N1118);
buf BUF1 (N1515, N1514);
or OR3 (N1516, N1511, N70, N1306);
xor XOR2 (N1517, N1515, N1086);
nor NOR4 (N1518, N1485, N250, N1091, N548);
nand NAND4 (N1519, N1510, N807, N1274, N1068);
buf BUF1 (N1520, N1508);
and AND4 (N1521, N1506, N1389, N372, N395);
xor XOR2 (N1522, N1518, N1349);
not NOT1 (N1523, N1519);
nand NAND4 (N1524, N1505, N1505, N1024, N1244);
buf BUF1 (N1525, N1523);
and AND3 (N1526, N1512, N692, N876);
nand NAND4 (N1527, N1521, N763, N428, N403);
or OR2 (N1528, N1526, N667);
xor XOR2 (N1529, N1520, N646);
not NOT1 (N1530, N1525);
or OR2 (N1531, N1513, N1028);
and AND3 (N1532, N1531, N721, N1472);
or OR2 (N1533, N1528, N1033);
buf BUF1 (N1534, N1533);
not NOT1 (N1535, N1496);
buf BUF1 (N1536, N1530);
nor NOR2 (N1537, N1529, N1376);
or OR3 (N1538, N1527, N358, N350);
xor XOR2 (N1539, N1537, N80);
and AND2 (N1540, N1539, N1208);
xor XOR2 (N1541, N1536, N720);
xor XOR2 (N1542, N1517, N733);
and AND3 (N1543, N1522, N1471, N195);
xor XOR2 (N1544, N1538, N1062);
and AND3 (N1545, N1532, N367, N193);
or OR4 (N1546, N1540, N145, N880, N387);
and AND3 (N1547, N1516, N933, N748);
nand NAND3 (N1548, N1534, N1449, N243);
and AND4 (N1549, N1547, N611, N203, N331);
or OR2 (N1550, N1548, N248);
and AND3 (N1551, N1541, N1172, N809);
buf BUF1 (N1552, N1542);
not NOT1 (N1553, N1544);
and AND3 (N1554, N1553, N1210, N423);
or OR3 (N1555, N1549, N544, N606);
nand NAND3 (N1556, N1555, N122, N763);
nand NAND2 (N1557, N1524, N1148);
not NOT1 (N1558, N1552);
not NOT1 (N1559, N1535);
nand NAND4 (N1560, N1556, N879, N844, N324);
xor XOR2 (N1561, N1560, N1136);
nor NOR4 (N1562, N1558, N950, N1450, N1008);
and AND2 (N1563, N1546, N2);
nand NAND2 (N1564, N1543, N242);
xor XOR2 (N1565, N1559, N955);
buf BUF1 (N1566, N1562);
or OR2 (N1567, N1565, N261);
and AND3 (N1568, N1545, N244, N1011);
not NOT1 (N1569, N1566);
buf BUF1 (N1570, N1567);
not NOT1 (N1571, N1568);
and AND3 (N1572, N1563, N431, N847);
nand NAND2 (N1573, N1572, N317);
not NOT1 (N1574, N1551);
and AND3 (N1575, N1570, N269, N1303);
and AND4 (N1576, N1564, N205, N1031, N135);
not NOT1 (N1577, N1574);
nor NOR3 (N1578, N1573, N1484, N657);
xor XOR2 (N1579, N1569, N1196);
nor NOR2 (N1580, N1561, N1051);
or OR2 (N1581, N1580, N1429);
or OR4 (N1582, N1577, N1026, N160, N987);
or OR2 (N1583, N1575, N1528);
or OR3 (N1584, N1582, N418, N165);
xor XOR2 (N1585, N1584, N740);
buf BUF1 (N1586, N1557);
or OR4 (N1587, N1554, N955, N1399, N1345);
nand NAND4 (N1588, N1571, N1428, N90, N646);
xor XOR2 (N1589, N1581, N934);
and AND2 (N1590, N1576, N913);
nand NAND4 (N1591, N1583, N555, N232, N176);
buf BUF1 (N1592, N1588);
or OR2 (N1593, N1591, N1177);
and AND4 (N1594, N1590, N583, N92, N1023);
nor NOR4 (N1595, N1592, N1575, N659, N1008);
or OR3 (N1596, N1550, N769, N996);
nor NOR3 (N1597, N1585, N1000, N458);
xor XOR2 (N1598, N1579, N1535);
xor XOR2 (N1599, N1578, N84);
nor NOR4 (N1600, N1596, N1145, N247, N167);
nor NOR2 (N1601, N1597, N743);
or OR4 (N1602, N1598, N121, N1015, N1357);
buf BUF1 (N1603, N1600);
nand NAND2 (N1604, N1595, N650);
and AND2 (N1605, N1586, N754);
xor XOR2 (N1606, N1602, N332);
or OR2 (N1607, N1604, N570);
nand NAND4 (N1608, N1593, N1478, N1004, N161);
or OR3 (N1609, N1608, N476, N1587);
nand NAND2 (N1610, N1545, N453);
nor NOR4 (N1611, N1603, N549, N751, N580);
nor NOR2 (N1612, N1589, N1219);
nand NAND2 (N1613, N1594, N821);
nor NOR3 (N1614, N1607, N122, N1006);
and AND4 (N1615, N1599, N587, N778, N1169);
or OR2 (N1616, N1610, N363);
buf BUF1 (N1617, N1613);
nand NAND3 (N1618, N1614, N783, N981);
nand NAND2 (N1619, N1609, N909);
not NOT1 (N1620, N1616);
and AND2 (N1621, N1601, N435);
not NOT1 (N1622, N1615);
xor XOR2 (N1623, N1611, N301);
and AND2 (N1624, N1619, N326);
nand NAND3 (N1625, N1605, N1613, N1220);
buf BUF1 (N1626, N1624);
not NOT1 (N1627, N1620);
or OR4 (N1628, N1606, N454, N965, N1539);
xor XOR2 (N1629, N1618, N1591);
buf BUF1 (N1630, N1625);
xor XOR2 (N1631, N1612, N879);
xor XOR2 (N1632, N1622, N226);
buf BUF1 (N1633, N1631);
nand NAND2 (N1634, N1623, N824);
and AND4 (N1635, N1632, N409, N1312, N1625);
or OR2 (N1636, N1630, N742);
and AND3 (N1637, N1627, N19, N868);
nor NOR2 (N1638, N1635, N591);
not NOT1 (N1639, N1628);
and AND4 (N1640, N1617, N1568, N80, N993);
or OR2 (N1641, N1621, N35);
nor NOR3 (N1642, N1634, N799, N875);
xor XOR2 (N1643, N1638, N1001);
not NOT1 (N1644, N1633);
not NOT1 (N1645, N1640);
and AND3 (N1646, N1642, N1244, N155);
and AND2 (N1647, N1645, N1168);
not NOT1 (N1648, N1644);
or OR4 (N1649, N1639, N1507, N871, N1514);
and AND2 (N1650, N1649, N228);
or OR3 (N1651, N1646, N1174, N403);
or OR2 (N1652, N1647, N1166);
buf BUF1 (N1653, N1651);
nor NOR3 (N1654, N1643, N1354, N361);
xor XOR2 (N1655, N1629, N1515);
nor NOR4 (N1656, N1626, N1331, N946, N1162);
and AND4 (N1657, N1637, N910, N300, N484);
nand NAND3 (N1658, N1653, N1011, N816);
xor XOR2 (N1659, N1657, N955);
not NOT1 (N1660, N1636);
nor NOR2 (N1661, N1660, N1118);
nand NAND4 (N1662, N1654, N1301, N425, N1447);
not NOT1 (N1663, N1658);
nor NOR4 (N1664, N1655, N1040, N653, N1238);
or OR4 (N1665, N1650, N1587, N1609, N841);
nor NOR2 (N1666, N1659, N564);
buf BUF1 (N1667, N1652);
xor XOR2 (N1668, N1656, N1643);
nand NAND4 (N1669, N1641, N1370, N1635, N1342);
xor XOR2 (N1670, N1666, N1227);
or OR2 (N1671, N1661, N363);
and AND4 (N1672, N1665, N1299, N991, N657);
or OR3 (N1673, N1667, N173, N440);
nand NAND2 (N1674, N1664, N1563);
nor NOR3 (N1675, N1671, N944, N1077);
not NOT1 (N1676, N1675);
xor XOR2 (N1677, N1663, N254);
buf BUF1 (N1678, N1662);
buf BUF1 (N1679, N1673);
not NOT1 (N1680, N1676);
buf BUF1 (N1681, N1678);
or OR4 (N1682, N1670, N1577, N578, N188);
or OR4 (N1683, N1669, N368, N1304, N1513);
nand NAND3 (N1684, N1668, N521, N1317);
buf BUF1 (N1685, N1674);
buf BUF1 (N1686, N1681);
or OR3 (N1687, N1679, N383, N1332);
nand NAND4 (N1688, N1686, N1265, N1236, N890);
buf BUF1 (N1689, N1680);
xor XOR2 (N1690, N1685, N1557);
buf BUF1 (N1691, N1672);
not NOT1 (N1692, N1688);
or OR4 (N1693, N1689, N574, N1599, N1141);
and AND2 (N1694, N1691, N4);
nand NAND2 (N1695, N1690, N1192);
not NOT1 (N1696, N1695);
buf BUF1 (N1697, N1692);
not NOT1 (N1698, N1677);
xor XOR2 (N1699, N1682, N1662);
buf BUF1 (N1700, N1687);
or OR2 (N1701, N1696, N730);
not NOT1 (N1702, N1699);
nand NAND4 (N1703, N1700, N921, N1154, N1097);
nand NAND2 (N1704, N1684, N610);
buf BUF1 (N1705, N1704);
or OR2 (N1706, N1702, N292);
or OR3 (N1707, N1706, N1341, N982);
not NOT1 (N1708, N1701);
nor NOR4 (N1709, N1693, N293, N783, N1525);
nand NAND3 (N1710, N1709, N806, N364);
nor NOR4 (N1711, N1710, N870, N1286, N1686);
not NOT1 (N1712, N1707);
nor NOR2 (N1713, N1703, N1053);
or OR2 (N1714, N1683, N827);
buf BUF1 (N1715, N1708);
nor NOR2 (N1716, N1715, N145);
or OR3 (N1717, N1697, N1496, N902);
or OR3 (N1718, N1648, N956, N868);
not NOT1 (N1719, N1716);
not NOT1 (N1720, N1719);
and AND2 (N1721, N1698, N687);
nand NAND3 (N1722, N1714, N1130, N1314);
or OR4 (N1723, N1720, N1420, N797, N727);
nand NAND4 (N1724, N1694, N1515, N1496, N978);
xor XOR2 (N1725, N1717, N156);
or OR3 (N1726, N1725, N1319, N481);
not NOT1 (N1727, N1713);
nand NAND3 (N1728, N1712, N640, N1106);
buf BUF1 (N1729, N1724);
not NOT1 (N1730, N1723);
nand NAND2 (N1731, N1722, N1669);
and AND4 (N1732, N1731, N254, N978, N343);
xor XOR2 (N1733, N1728, N1689);
and AND4 (N1734, N1727, N485, N109, N581);
not NOT1 (N1735, N1733);
and AND4 (N1736, N1711, N200, N1445, N684);
not NOT1 (N1737, N1732);
nor NOR2 (N1738, N1726, N1478);
or OR2 (N1739, N1729, N1194);
or OR4 (N1740, N1730, N112, N1403, N119);
or OR2 (N1741, N1705, N143);
nor NOR4 (N1742, N1735, N62, N1470, N642);
not NOT1 (N1743, N1738);
nand NAND4 (N1744, N1741, N664, N748, N866);
nand NAND4 (N1745, N1737, N1602, N1187, N151);
xor XOR2 (N1746, N1742, N497);
nand NAND3 (N1747, N1736, N1688, N741);
nand NAND3 (N1748, N1721, N1504, N160);
not NOT1 (N1749, N1734);
xor XOR2 (N1750, N1745, N1262);
not NOT1 (N1751, N1740);
nor NOR4 (N1752, N1750, N963, N995, N1181);
buf BUF1 (N1753, N1751);
buf BUF1 (N1754, N1746);
nor NOR4 (N1755, N1739, N1672, N1162, N138);
nor NOR2 (N1756, N1748, N1603);
buf BUF1 (N1757, N1744);
xor XOR2 (N1758, N1756, N105);
nand NAND4 (N1759, N1754, N983, N1519, N625);
xor XOR2 (N1760, N1757, N1476);
nand NAND4 (N1761, N1755, N1422, N842, N723);
and AND2 (N1762, N1743, N594);
not NOT1 (N1763, N1762);
nand NAND3 (N1764, N1761, N1540, N645);
buf BUF1 (N1765, N1718);
nand NAND3 (N1766, N1753, N954, N1351);
not NOT1 (N1767, N1749);
not NOT1 (N1768, N1765);
xor XOR2 (N1769, N1747, N146);
not NOT1 (N1770, N1763);
nand NAND3 (N1771, N1752, N1074, N1177);
nor NOR4 (N1772, N1770, N937, N1115, N573);
nor NOR3 (N1773, N1760, N419, N1723);
nand NAND3 (N1774, N1766, N55, N1373);
or OR3 (N1775, N1769, N930, N738);
xor XOR2 (N1776, N1774, N983);
xor XOR2 (N1777, N1772, N1116);
nand NAND3 (N1778, N1758, N795, N1509);
not NOT1 (N1779, N1768);
and AND2 (N1780, N1767, N552);
and AND4 (N1781, N1775, N1656, N1239, N863);
xor XOR2 (N1782, N1764, N1034);
and AND2 (N1783, N1780, N1377);
xor XOR2 (N1784, N1783, N1122);
and AND4 (N1785, N1779, N214, N1521, N1179);
nor NOR3 (N1786, N1759, N132, N746);
xor XOR2 (N1787, N1781, N1658);
not NOT1 (N1788, N1778);
not NOT1 (N1789, N1788);
nor NOR3 (N1790, N1777, N196, N1381);
not NOT1 (N1791, N1782);
not NOT1 (N1792, N1791);
xor XOR2 (N1793, N1787, N1489);
and AND4 (N1794, N1785, N1524, N245, N1000);
xor XOR2 (N1795, N1773, N19);
and AND4 (N1796, N1792, N1326, N215, N570);
nor NOR3 (N1797, N1793, N41, N115);
or OR3 (N1798, N1796, N555, N656);
xor XOR2 (N1799, N1776, N760);
and AND4 (N1800, N1797, N1322, N567, N1340);
xor XOR2 (N1801, N1795, N1286);
buf BUF1 (N1802, N1771);
buf BUF1 (N1803, N1800);
and AND3 (N1804, N1789, N670, N1345);
nand NAND4 (N1805, N1799, N1115, N519, N641);
and AND4 (N1806, N1790, N426, N1068, N305);
xor XOR2 (N1807, N1784, N308);
buf BUF1 (N1808, N1803);
buf BUF1 (N1809, N1802);
buf BUF1 (N1810, N1807);
nand NAND4 (N1811, N1804, N599, N436, N618);
or OR4 (N1812, N1801, N1310, N780, N923);
nor NOR2 (N1813, N1786, N395);
or OR3 (N1814, N1794, N1468, N866);
nand NAND3 (N1815, N1806, N1702, N987);
buf BUF1 (N1816, N1808);
xor XOR2 (N1817, N1809, N1612);
nand NAND4 (N1818, N1811, N1156, N979, N1670);
and AND3 (N1819, N1810, N394, N1535);
nand NAND3 (N1820, N1816, N642, N268);
or OR3 (N1821, N1805, N790, N107);
xor XOR2 (N1822, N1818, N916);
not NOT1 (N1823, N1819);
not NOT1 (N1824, N1823);
buf BUF1 (N1825, N1824);
or OR4 (N1826, N1817, N214, N1454, N1368);
xor XOR2 (N1827, N1813, N677);
xor XOR2 (N1828, N1826, N1310);
buf BUF1 (N1829, N1821);
or OR2 (N1830, N1829, N1458);
and AND3 (N1831, N1827, N675, N597);
and AND4 (N1832, N1822, N600, N780, N1471);
or OR2 (N1833, N1815, N922);
not NOT1 (N1834, N1831);
not NOT1 (N1835, N1833);
not NOT1 (N1836, N1812);
xor XOR2 (N1837, N1830, N252);
or OR2 (N1838, N1837, N541);
buf BUF1 (N1839, N1814);
nor NOR3 (N1840, N1828, N739, N1145);
not NOT1 (N1841, N1838);
nor NOR3 (N1842, N1839, N1523, N346);
and AND3 (N1843, N1841, N783, N794);
buf BUF1 (N1844, N1834);
xor XOR2 (N1845, N1798, N1383);
and AND3 (N1846, N1840, N1729, N515);
nor NOR3 (N1847, N1844, N156, N36);
nand NAND2 (N1848, N1836, N651);
nand NAND2 (N1849, N1835, N418);
nand NAND2 (N1850, N1832, N1380);
xor XOR2 (N1851, N1820, N1690);
xor XOR2 (N1852, N1847, N940);
not NOT1 (N1853, N1843);
not NOT1 (N1854, N1842);
xor XOR2 (N1855, N1849, N1776);
nand NAND3 (N1856, N1855, N1432, N264);
xor XOR2 (N1857, N1825, N553);
buf BUF1 (N1858, N1846);
buf BUF1 (N1859, N1856);
not NOT1 (N1860, N1845);
xor XOR2 (N1861, N1853, N265);
and AND4 (N1862, N1848, N1323, N1580, N969);
and AND4 (N1863, N1862, N1212, N180, N561);
buf BUF1 (N1864, N1858);
or OR4 (N1865, N1857, N266, N890, N486);
nand NAND4 (N1866, N1865, N1580, N213, N1598);
xor XOR2 (N1867, N1863, N922);
and AND4 (N1868, N1864, N876, N850, N1247);
nor NOR2 (N1869, N1859, N995);
and AND4 (N1870, N1867, N1289, N1443, N563);
nor NOR4 (N1871, N1868, N494, N1037, N734);
and AND2 (N1872, N1860, N851);
and AND2 (N1873, N1871, N1226);
buf BUF1 (N1874, N1850);
buf BUF1 (N1875, N1869);
nand NAND2 (N1876, N1866, N1690);
nor NOR3 (N1877, N1854, N1611, N1771);
buf BUF1 (N1878, N1874);
buf BUF1 (N1879, N1861);
buf BUF1 (N1880, N1872);
or OR2 (N1881, N1873, N224);
and AND4 (N1882, N1870, N214, N1767, N845);
nand NAND4 (N1883, N1880, N496, N1376, N1223);
and AND4 (N1884, N1875, N61, N640, N470);
not NOT1 (N1885, N1851);
and AND2 (N1886, N1882, N1803);
xor XOR2 (N1887, N1884, N88);
or OR3 (N1888, N1886, N1519, N258);
nor NOR2 (N1889, N1878, N1088);
buf BUF1 (N1890, N1887);
or OR4 (N1891, N1885, N1857, N1334, N1832);
nor NOR2 (N1892, N1877, N1735);
buf BUF1 (N1893, N1883);
buf BUF1 (N1894, N1892);
and AND2 (N1895, N1891, N802);
nand NAND4 (N1896, N1888, N1333, N1773, N1755);
xor XOR2 (N1897, N1893, N646);
and AND4 (N1898, N1894, N117, N340, N299);
nand NAND2 (N1899, N1852, N641);
and AND2 (N1900, N1895, N1627);
nor NOR3 (N1901, N1876, N770, N946);
xor XOR2 (N1902, N1890, N1690);
nor NOR4 (N1903, N1897, N1555, N1538, N141);
buf BUF1 (N1904, N1881);
not NOT1 (N1905, N1903);
and AND2 (N1906, N1879, N1586);
and AND2 (N1907, N1901, N1395);
not NOT1 (N1908, N1904);
nor NOR4 (N1909, N1898, N904, N446, N988);
not NOT1 (N1910, N1906);
and AND4 (N1911, N1889, N1705, N1698, N1786);
buf BUF1 (N1912, N1910);
nor NOR4 (N1913, N1896, N559, N855, N1431);
not NOT1 (N1914, N1905);
buf BUF1 (N1915, N1914);
buf BUF1 (N1916, N1900);
buf BUF1 (N1917, N1909);
buf BUF1 (N1918, N1899);
nor NOR2 (N1919, N1912, N1363);
or OR4 (N1920, N1907, N428, N1721, N66);
nand NAND3 (N1921, N1911, N509, N1174);
xor XOR2 (N1922, N1902, N1143);
not NOT1 (N1923, N1922);
nor NOR3 (N1924, N1913, N477, N1063);
or OR2 (N1925, N1916, N1328);
and AND4 (N1926, N1924, N1658, N1387, N321);
and AND4 (N1927, N1921, N1228, N1227, N781);
not NOT1 (N1928, N1919);
not NOT1 (N1929, N1926);
and AND3 (N1930, N1915, N780, N1250);
buf BUF1 (N1931, N1928);
nor NOR3 (N1932, N1931, N408, N671);
and AND4 (N1933, N1917, N3, N1644, N1522);
or OR4 (N1934, N1929, N1701, N795, N543);
nor NOR3 (N1935, N1930, N599, N1149);
nand NAND4 (N1936, N1932, N831, N1104, N373);
or OR3 (N1937, N1923, N873, N652);
nand NAND2 (N1938, N1927, N290);
nor NOR2 (N1939, N1933, N660);
not NOT1 (N1940, N1935);
or OR2 (N1941, N1940, N1725);
xor XOR2 (N1942, N1937, N1029);
buf BUF1 (N1943, N1941);
nor NOR4 (N1944, N1918, N1894, N1170, N136);
xor XOR2 (N1945, N1944, N1224);
or OR4 (N1946, N1925, N1018, N725, N1013);
nor NOR3 (N1947, N1938, N1034, N1548);
and AND4 (N1948, N1934, N1162, N862, N906);
nor NOR2 (N1949, N1936, N392);
and AND3 (N1950, N1943, N893, N1764);
xor XOR2 (N1951, N1950, N538);
not NOT1 (N1952, N1920);
and AND2 (N1953, N1942, N310);
not NOT1 (N1954, N1953);
buf BUF1 (N1955, N1948);
buf BUF1 (N1956, N1939);
not NOT1 (N1957, N1908);
xor XOR2 (N1958, N1956, N1194);
buf BUF1 (N1959, N1952);
buf BUF1 (N1960, N1946);
not NOT1 (N1961, N1949);
nor NOR3 (N1962, N1951, N709, N1278);
or OR3 (N1963, N1945, N1134, N1052);
buf BUF1 (N1964, N1961);
or OR2 (N1965, N1960, N95);
nand NAND4 (N1966, N1947, N1558, N1588, N1255);
nor NOR4 (N1967, N1957, N786, N1495, N101);
nand NAND4 (N1968, N1963, N645, N748, N1556);
buf BUF1 (N1969, N1968);
or OR2 (N1970, N1969, N758);
and AND2 (N1971, N1964, N1165);
buf BUF1 (N1972, N1954);
xor XOR2 (N1973, N1962, N560);
or OR4 (N1974, N1955, N138, N846, N611);
xor XOR2 (N1975, N1959, N988);
nand NAND4 (N1976, N1975, N556, N295, N1779);
and AND3 (N1977, N1970, N267, N1548);
and AND4 (N1978, N1958, N1976, N523, N1606);
not NOT1 (N1979, N948);
buf BUF1 (N1980, N1979);
buf BUF1 (N1981, N1966);
and AND3 (N1982, N1973, N988, N948);
not NOT1 (N1983, N1967);
and AND3 (N1984, N1977, N559, N51);
nand NAND2 (N1985, N1984, N1029);
or OR2 (N1986, N1974, N1175);
xor XOR2 (N1987, N1981, N1478);
buf BUF1 (N1988, N1965);
xor XOR2 (N1989, N1983, N1425);
not NOT1 (N1990, N1972);
nand NAND4 (N1991, N1990, N587, N1227, N442);
and AND3 (N1992, N1978, N1107, N1052);
nor NOR2 (N1993, N1982, N1644);
xor XOR2 (N1994, N1985, N578);
nor NOR2 (N1995, N1987, N1158);
or OR3 (N1996, N1971, N1509, N326);
not NOT1 (N1997, N1994);
and AND3 (N1998, N1989, N1048, N16);
nand NAND4 (N1999, N1991, N319, N212, N1423);
not NOT1 (N2000, N1986);
and AND2 (N2001, N1980, N1867);
or OR3 (N2002, N1992, N637, N105);
not NOT1 (N2003, N1993);
or OR3 (N2004, N2000, N766, N537);
xor XOR2 (N2005, N1996, N378);
not NOT1 (N2006, N1998);
nand NAND2 (N2007, N1997, N752);
not NOT1 (N2008, N1988);
not NOT1 (N2009, N1995);
nor NOR2 (N2010, N2008, N413);
or OR3 (N2011, N2004, N501, N513);
nor NOR4 (N2012, N2007, N1722, N642, N1691);
nand NAND3 (N2013, N2005, N511, N304);
or OR3 (N2014, N2011, N1829, N2010);
buf BUF1 (N2015, N1132);
and AND3 (N2016, N2003, N955, N1881);
nor NOR3 (N2017, N2001, N629, N1706);
xor XOR2 (N2018, N2013, N1794);
xor XOR2 (N2019, N2009, N1459);
nand NAND2 (N2020, N2014, N993);
and AND3 (N2021, N2019, N808, N1886);
nand NAND4 (N2022, N2021, N1934, N790, N135);
and AND3 (N2023, N2017, N1316, N1422);
not NOT1 (N2024, N2023);
nand NAND4 (N2025, N2022, N1887, N326, N656);
or OR2 (N2026, N2025, N1002);
nand NAND2 (N2027, N2002, N1691);
and AND2 (N2028, N2027, N214);
nand NAND2 (N2029, N1999, N43);
and AND2 (N2030, N2006, N2028);
nor NOR2 (N2031, N1777, N473);
nand NAND2 (N2032, N2030, N1789);
nor NOR2 (N2033, N2020, N1240);
xor XOR2 (N2034, N2024, N1531);
or OR4 (N2035, N2018, N1147, N506, N1820);
nand NAND2 (N2036, N2031, N1536);
or OR4 (N2037, N2016, N836, N117, N202);
nor NOR3 (N2038, N2036, N1484, N1939);
not NOT1 (N2039, N2038);
nor NOR2 (N2040, N2034, N1617);
not NOT1 (N2041, N2012);
and AND2 (N2042, N2026, N1993);
or OR2 (N2043, N2042, N291);
xor XOR2 (N2044, N2040, N875);
or OR2 (N2045, N2043, N287);
or OR2 (N2046, N2015, N18);
nor NOR4 (N2047, N2035, N718, N388, N1659);
nand NAND2 (N2048, N2037, N913);
not NOT1 (N2049, N2039);
xor XOR2 (N2050, N2048, N1055);
nand NAND3 (N2051, N2049, N1896, N688);
nor NOR3 (N2052, N2041, N1545, N1754);
and AND2 (N2053, N2045, N2020);
nand NAND4 (N2054, N2044, N750, N1167, N1702);
not NOT1 (N2055, N2047);
or OR3 (N2056, N2055, N94, N1509);
buf BUF1 (N2057, N2046);
nor NOR4 (N2058, N2053, N1282, N706, N1333);
nand NAND4 (N2059, N2050, N1565, N640, N1644);
buf BUF1 (N2060, N2029);
or OR4 (N2061, N2056, N1612, N773, N600);
nand NAND4 (N2062, N2059, N31, N68, N1765);
or OR2 (N2063, N2062, N1419);
or OR3 (N2064, N2033, N481, N1165);
or OR3 (N2065, N2054, N1373, N1543);
and AND3 (N2066, N2058, N1005, N2045);
and AND3 (N2067, N2063, N322, N1264);
or OR3 (N2068, N2052, N320, N81);
nand NAND2 (N2069, N2066, N1866);
or OR4 (N2070, N2065, N1938, N826, N943);
buf BUF1 (N2071, N2051);
buf BUF1 (N2072, N2071);
not NOT1 (N2073, N2032);
nor NOR4 (N2074, N2070, N1404, N1710, N1620);
not NOT1 (N2075, N2073);
not NOT1 (N2076, N2069);
nand NAND3 (N2077, N2068, N634, N170);
nand NAND2 (N2078, N2076, N1479);
xor XOR2 (N2079, N2074, N1257);
and AND3 (N2080, N2057, N1620, N1678);
and AND3 (N2081, N2067, N123, N1679);
nand NAND4 (N2082, N2081, N537, N1734, N414);
or OR4 (N2083, N2072, N1000, N1990, N306);
or OR4 (N2084, N2083, N1532, N1112, N1107);
xor XOR2 (N2085, N2064, N367);
or OR2 (N2086, N2085, N1393);
buf BUF1 (N2087, N2061);
nor NOR4 (N2088, N2079, N1688, N1948, N979);
xor XOR2 (N2089, N2086, N1248);
nand NAND3 (N2090, N2088, N2011, N1978);
buf BUF1 (N2091, N2080);
nor NOR2 (N2092, N2082, N891);
buf BUF1 (N2093, N2091);
and AND2 (N2094, N2087, N353);
and AND3 (N2095, N2092, N1718, N1169);
buf BUF1 (N2096, N2089);
or OR3 (N2097, N2077, N435, N508);
nor NOR4 (N2098, N2094, N15, N1082, N11);
buf BUF1 (N2099, N2098);
or OR4 (N2100, N2084, N240, N94, N603);
and AND3 (N2101, N2060, N694, N1613);
and AND3 (N2102, N2100, N653, N766);
nand NAND4 (N2103, N2101, N1920, N33, N838);
or OR2 (N2104, N2078, N1912);
nand NAND4 (N2105, N2096, N690, N1146, N40);
buf BUF1 (N2106, N2099);
nand NAND4 (N2107, N2075, N221, N863, N237);
not NOT1 (N2108, N2090);
or OR2 (N2109, N2106, N144);
nor NOR2 (N2110, N2093, N365);
nand NAND2 (N2111, N2104, N476);
not NOT1 (N2112, N2108);
and AND4 (N2113, N2095, N539, N621, N1865);
buf BUF1 (N2114, N2102);
and AND4 (N2115, N2103, N1, N1573, N1073);
not NOT1 (N2116, N2097);
xor XOR2 (N2117, N2111, N2086);
buf BUF1 (N2118, N2117);
buf BUF1 (N2119, N2113);
and AND2 (N2120, N2119, N1200);
buf BUF1 (N2121, N2109);
buf BUF1 (N2122, N2110);
and AND4 (N2123, N2120, N103, N698, N1327);
xor XOR2 (N2124, N2121, N1100);
and AND3 (N2125, N2124, N978, N303);
xor XOR2 (N2126, N2118, N630);
buf BUF1 (N2127, N2107);
nor NOR3 (N2128, N2122, N1371, N1726);
or OR3 (N2129, N2105, N480, N265);
and AND3 (N2130, N2129, N430, N2039);
buf BUF1 (N2131, N2125);
xor XOR2 (N2132, N2130, N765);
buf BUF1 (N2133, N2132);
xor XOR2 (N2134, N2116, N1884);
xor XOR2 (N2135, N2128, N1548);
and AND3 (N2136, N2127, N1939, N929);
not NOT1 (N2137, N2136);
nand NAND2 (N2138, N2114, N1333);
or OR2 (N2139, N2112, N1087);
or OR2 (N2140, N2137, N1900);
xor XOR2 (N2141, N2134, N611);
xor XOR2 (N2142, N2126, N1948);
and AND2 (N2143, N2141, N1347);
or OR2 (N2144, N2139, N402);
or OR3 (N2145, N2131, N1090, N1454);
buf BUF1 (N2146, N2138);
xor XOR2 (N2147, N2142, N437);
nand NAND3 (N2148, N2143, N1896, N1527);
or OR2 (N2149, N2144, N382);
nor NOR4 (N2150, N2135, N112, N375, N473);
and AND2 (N2151, N2146, N252);
or OR3 (N2152, N2149, N1554, N1572);
and AND2 (N2153, N2133, N518);
not NOT1 (N2154, N2123);
buf BUF1 (N2155, N2145);
nand NAND3 (N2156, N2151, N729, N2112);
nor NOR2 (N2157, N2154, N1709);
not NOT1 (N2158, N2152);
nor NOR3 (N2159, N2150, N298, N1304);
and AND3 (N2160, N2140, N1934, N1200);
not NOT1 (N2161, N2157);
xor XOR2 (N2162, N2156, N1441);
and AND2 (N2163, N2115, N1012);
and AND2 (N2164, N2155, N1460);
buf BUF1 (N2165, N2158);
not NOT1 (N2166, N2165);
and AND4 (N2167, N2148, N1375, N1395, N1886);
and AND4 (N2168, N2147, N1643, N162, N2094);
not NOT1 (N2169, N2166);
not NOT1 (N2170, N2163);
buf BUF1 (N2171, N2169);
nand NAND3 (N2172, N2168, N1568, N1076);
nor NOR4 (N2173, N2160, N171, N160, N737);
nand NAND2 (N2174, N2171, N1483);
or OR3 (N2175, N2170, N1644, N803);
xor XOR2 (N2176, N2153, N819);
buf BUF1 (N2177, N2174);
or OR3 (N2178, N2175, N202, N302);
nor NOR4 (N2179, N2176, N1749, N891, N1270);
and AND2 (N2180, N2164, N436);
and AND4 (N2181, N2180, N985, N85, N1577);
xor XOR2 (N2182, N2181, N1654);
xor XOR2 (N2183, N2162, N1419);
buf BUF1 (N2184, N2167);
nand NAND2 (N2185, N2159, N1951);
nor NOR4 (N2186, N2173, N510, N1875, N978);
and AND4 (N2187, N2172, N285, N2001, N1039);
nand NAND2 (N2188, N2178, N753);
and AND3 (N2189, N2187, N266, N775);
not NOT1 (N2190, N2188);
and AND3 (N2191, N2161, N515, N1636);
xor XOR2 (N2192, N2179, N1158);
nor NOR2 (N2193, N2184, N1895);
buf BUF1 (N2194, N2193);
or OR2 (N2195, N2185, N528);
and AND4 (N2196, N2182, N637, N468, N1375);
and AND4 (N2197, N2186, N1689, N1262, N1373);
nor NOR2 (N2198, N2191, N111);
nand NAND4 (N2199, N2194, N717, N1239, N1518);
and AND2 (N2200, N2190, N992);
nor NOR2 (N2201, N2192, N1019);
xor XOR2 (N2202, N2195, N1093);
and AND4 (N2203, N2199, N40, N613, N565);
buf BUF1 (N2204, N2197);
xor XOR2 (N2205, N2202, N300);
nand NAND3 (N2206, N2196, N1233, N1611);
xor XOR2 (N2207, N2200, N1281);
and AND4 (N2208, N2205, N1425, N1344, N61);
or OR2 (N2209, N2208, N1096);
buf BUF1 (N2210, N2204);
or OR3 (N2211, N2206, N1506, N2018);
buf BUF1 (N2212, N2211);
xor XOR2 (N2213, N2201, N1669);
nand NAND3 (N2214, N2177, N399, N841);
not NOT1 (N2215, N2209);
xor XOR2 (N2216, N2212, N2081);
buf BUF1 (N2217, N2214);
nor NOR4 (N2218, N2213, N1726, N329, N580);
nand NAND3 (N2219, N2203, N309, N2063);
or OR4 (N2220, N2198, N701, N1398, N1263);
nor NOR3 (N2221, N2217, N220, N2040);
and AND2 (N2222, N2219, N262);
or OR4 (N2223, N2210, N475, N2056, N1988);
or OR2 (N2224, N2207, N139);
xor XOR2 (N2225, N2183, N1541);
nand NAND4 (N2226, N2216, N1661, N1844, N1207);
nor NOR2 (N2227, N2223, N886);
nor NOR4 (N2228, N2220, N942, N307, N2163);
and AND4 (N2229, N2215, N1206, N1114, N1547);
xor XOR2 (N2230, N2228, N294);
and AND3 (N2231, N2226, N1461, N1432);
nand NAND3 (N2232, N2222, N886, N1449);
or OR2 (N2233, N2227, N204);
not NOT1 (N2234, N2231);
not NOT1 (N2235, N2233);
not NOT1 (N2236, N2225);
xor XOR2 (N2237, N2229, N369);
and AND3 (N2238, N2232, N391, N2044);
not NOT1 (N2239, N2189);
nor NOR2 (N2240, N2236, N874);
or OR4 (N2241, N2218, N498, N464, N667);
not NOT1 (N2242, N2240);
xor XOR2 (N2243, N2221, N1863);
or OR2 (N2244, N2234, N1855);
nand NAND4 (N2245, N2243, N1291, N765, N1033);
nand NAND3 (N2246, N2224, N1052, N1517);
nand NAND3 (N2247, N2246, N262, N1306);
nand NAND2 (N2248, N2238, N1843);
or OR3 (N2249, N2241, N339, N2085);
xor XOR2 (N2250, N2235, N1986);
not NOT1 (N2251, N2239);
xor XOR2 (N2252, N2244, N1858);
buf BUF1 (N2253, N2249);
nor NOR4 (N2254, N2245, N1794, N2052, N222);
or OR3 (N2255, N2248, N518, N694);
nand NAND4 (N2256, N2250, N1089, N1288, N1321);
nand NAND3 (N2257, N2256, N925, N971);
buf BUF1 (N2258, N2247);
nand NAND2 (N2259, N2254, N1549);
and AND4 (N2260, N2237, N556, N1491, N39);
nor NOR3 (N2261, N2257, N271, N1822);
buf BUF1 (N2262, N2252);
or OR3 (N2263, N2255, N1137, N75);
nor NOR4 (N2264, N2260, N2096, N1009, N492);
buf BUF1 (N2265, N2261);
or OR4 (N2266, N2265, N677, N1971, N1428);
not NOT1 (N2267, N2259);
not NOT1 (N2268, N2230);
xor XOR2 (N2269, N2263, N264);
nor NOR4 (N2270, N2264, N382, N2110, N984);
xor XOR2 (N2271, N2268, N2011);
xor XOR2 (N2272, N2258, N2045);
nand NAND3 (N2273, N2242, N2127, N614);
xor XOR2 (N2274, N2251, N750);
not NOT1 (N2275, N2274);
xor XOR2 (N2276, N2275, N2071);
nor NOR3 (N2277, N2253, N555, N968);
buf BUF1 (N2278, N2262);
xor XOR2 (N2279, N2269, N1915);
buf BUF1 (N2280, N2279);
and AND4 (N2281, N2273, N491, N1035, N169);
not NOT1 (N2282, N2266);
buf BUF1 (N2283, N2276);
xor XOR2 (N2284, N2271, N1578);
nand NAND4 (N2285, N2278, N17, N429, N304);
xor XOR2 (N2286, N2280, N2073);
and AND3 (N2287, N2286, N1604, N417);
nand NAND3 (N2288, N2270, N613, N1667);
xor XOR2 (N2289, N2277, N336);
nand NAND2 (N2290, N2267, N1779);
or OR2 (N2291, N2281, N1966);
or OR3 (N2292, N2284, N305, N1000);
or OR4 (N2293, N2283, N1118, N1390, N1020);
nor NOR3 (N2294, N2272, N1469, N1196);
or OR3 (N2295, N2294, N1157, N1108);
and AND3 (N2296, N2287, N462, N1595);
or OR2 (N2297, N2285, N2247);
nand NAND3 (N2298, N2297, N1726, N1573);
or OR2 (N2299, N2282, N1145);
nand NAND3 (N2300, N2291, N1735, N1784);
nand NAND2 (N2301, N2298, N1439);
not NOT1 (N2302, N2299);
or OR2 (N2303, N2300, N2095);
xor XOR2 (N2304, N2293, N1506);
nor NOR2 (N2305, N2290, N482);
xor XOR2 (N2306, N2295, N708);
or OR4 (N2307, N2306, N1150, N600, N656);
nand NAND2 (N2308, N2304, N1713);
xor XOR2 (N2309, N2307, N619);
and AND3 (N2310, N2303, N386, N1586);
nand NAND4 (N2311, N2301, N452, N2255, N2113);
nor NOR3 (N2312, N2292, N2295, N254);
nor NOR4 (N2313, N2302, N333, N565, N1659);
or OR2 (N2314, N2305, N2118);
buf BUF1 (N2315, N2314);
not NOT1 (N2316, N2289);
nand NAND2 (N2317, N2311, N1919);
nand NAND2 (N2318, N2310, N2155);
nand NAND2 (N2319, N2313, N91);
not NOT1 (N2320, N2312);
and AND3 (N2321, N2309, N1668, N1429);
xor XOR2 (N2322, N2321, N1164);
or OR3 (N2323, N2319, N1041, N1924);
xor XOR2 (N2324, N2316, N1683);
nor NOR3 (N2325, N2308, N143, N362);
and AND4 (N2326, N2288, N399, N1442, N1427);
buf BUF1 (N2327, N2315);
nor NOR4 (N2328, N2327, N16, N1194, N591);
nor NOR3 (N2329, N2325, N2039, N1516);
or OR2 (N2330, N2329, N1494);
buf BUF1 (N2331, N2322);
nand NAND3 (N2332, N2320, N1803, N266);
nor NOR3 (N2333, N2296, N1543, N1240);
or OR4 (N2334, N2331, N1766, N114, N2281);
xor XOR2 (N2335, N2330, N883);
not NOT1 (N2336, N2332);
and AND2 (N2337, N2328, N813);
not NOT1 (N2338, N2317);
nand NAND4 (N2339, N2334, N1350, N1110, N1477);
xor XOR2 (N2340, N2333, N184);
buf BUF1 (N2341, N2323);
and AND4 (N2342, N2336, N9, N2125, N1183);
not NOT1 (N2343, N2341);
nor NOR3 (N2344, N2326, N834, N1299);
not NOT1 (N2345, N2344);
not NOT1 (N2346, N2345);
and AND4 (N2347, N2346, N630, N601, N117);
nor NOR3 (N2348, N2339, N645, N1064);
not NOT1 (N2349, N2340);
nor NOR4 (N2350, N2347, N1912, N1041, N378);
or OR3 (N2351, N2343, N426, N834);
nand NAND3 (N2352, N2318, N2313, N1485);
xor XOR2 (N2353, N2324, N1569);
xor XOR2 (N2354, N2348, N1875);
and AND3 (N2355, N2349, N49, N451);
and AND2 (N2356, N2342, N26);
nor NOR2 (N2357, N2356, N2003);
buf BUF1 (N2358, N2351);
nand NAND3 (N2359, N2350, N1711, N402);
xor XOR2 (N2360, N2352, N90);
nand NAND4 (N2361, N2353, N2300, N536, N1365);
nor NOR4 (N2362, N2357, N1732, N1565, N1983);
or OR2 (N2363, N2362, N546);
and AND2 (N2364, N2354, N648);
or OR2 (N2365, N2338, N312);
nand NAND3 (N2366, N2358, N1051, N432);
and AND3 (N2367, N2337, N513, N1391);
and AND2 (N2368, N2335, N1807);
nor NOR3 (N2369, N2361, N595, N1320);
and AND2 (N2370, N2364, N21);
and AND4 (N2371, N2366, N401, N1221, N1486);
xor XOR2 (N2372, N2359, N1461);
or OR3 (N2373, N2363, N382, N1980);
buf BUF1 (N2374, N2367);
buf BUF1 (N2375, N2368);
or OR2 (N2376, N2373, N940);
buf BUF1 (N2377, N2355);
or OR2 (N2378, N2371, N582);
buf BUF1 (N2379, N2369);
nor NOR3 (N2380, N2370, N343, N2199);
or OR4 (N2381, N2360, N608, N498, N248);
or OR4 (N2382, N2379, N1600, N785, N768);
or OR3 (N2383, N2365, N2142, N1137);
buf BUF1 (N2384, N2383);
or OR2 (N2385, N2380, N162);
and AND3 (N2386, N2377, N987, N1848);
and AND4 (N2387, N2375, N697, N132, N1354);
buf BUF1 (N2388, N2381);
nand NAND3 (N2389, N2376, N1001, N1777);
nor NOR4 (N2390, N2378, N332, N1427, N551);
not NOT1 (N2391, N2388);
nand NAND3 (N2392, N2385, N336, N391);
or OR4 (N2393, N2389, N1719, N956, N2256);
buf BUF1 (N2394, N2384);
nor NOR2 (N2395, N2386, N1562);
not NOT1 (N2396, N2393);
nand NAND4 (N2397, N2374, N1722, N1164, N996);
nor NOR2 (N2398, N2392, N484);
nor NOR2 (N2399, N2372, N826);
and AND4 (N2400, N2398, N1260, N1228, N1017);
buf BUF1 (N2401, N2396);
buf BUF1 (N2402, N2400);
nand NAND2 (N2403, N2394, N1702);
or OR4 (N2404, N2401, N1584, N73, N1185);
not NOT1 (N2405, N2402);
buf BUF1 (N2406, N2387);
and AND4 (N2407, N2397, N1533, N1293, N975);
nand NAND3 (N2408, N2390, N1931, N2063);
and AND3 (N2409, N2405, N2146, N604);
nor NOR3 (N2410, N2409, N466, N398);
nand NAND2 (N2411, N2382, N2197);
buf BUF1 (N2412, N2391);
and AND4 (N2413, N2399, N2351, N1712, N1468);
and AND4 (N2414, N2412, N1172, N755, N1794);
xor XOR2 (N2415, N2411, N2027);
nor NOR4 (N2416, N2395, N818, N766, N1706);
not NOT1 (N2417, N2410);
and AND3 (N2418, N2413, N1077, N2153);
nand NAND4 (N2419, N2417, N813, N1614, N2370);
not NOT1 (N2420, N2419);
or OR4 (N2421, N2414, N1320, N1049, N119);
nor NOR4 (N2422, N2416, N2129, N575, N613);
or OR2 (N2423, N2408, N754);
nor NOR2 (N2424, N2421, N467);
not NOT1 (N2425, N2420);
and AND3 (N2426, N2425, N1428, N1317);
xor XOR2 (N2427, N2415, N2036);
nor NOR3 (N2428, N2407, N2197, N1558);
not NOT1 (N2429, N2403);
nor NOR4 (N2430, N2404, N1861, N308, N2055);
nand NAND2 (N2431, N2422, N224);
buf BUF1 (N2432, N2406);
and AND2 (N2433, N2430, N2140);
and AND2 (N2434, N2424, N874);
buf BUF1 (N2435, N2427);
nor NOR2 (N2436, N2432, N633);
xor XOR2 (N2437, N2436, N899);
nand NAND3 (N2438, N2423, N296, N2281);
or OR4 (N2439, N2429, N1387, N2123, N1514);
and AND4 (N2440, N2439, N627, N770, N2107);
or OR3 (N2441, N2428, N21, N1112);
not NOT1 (N2442, N2440);
or OR2 (N2443, N2435, N1818);
buf BUF1 (N2444, N2431);
nand NAND2 (N2445, N2434, N794);
or OR3 (N2446, N2441, N1840, N2178);
xor XOR2 (N2447, N2446, N2392);
not NOT1 (N2448, N2447);
buf BUF1 (N2449, N2443);
nand NAND3 (N2450, N2448, N1380, N1120);
not NOT1 (N2451, N2449);
or OR3 (N2452, N2450, N2020, N1090);
or OR3 (N2453, N2433, N1808, N1069);
and AND2 (N2454, N2418, N1166);
not NOT1 (N2455, N2437);
not NOT1 (N2456, N2426);
nand NAND3 (N2457, N2451, N669, N332);
nor NOR4 (N2458, N2444, N1622, N1527, N2117);
or OR3 (N2459, N2453, N1934, N1204);
and AND4 (N2460, N2459, N1211, N2364, N1944);
not NOT1 (N2461, N2456);
not NOT1 (N2462, N2458);
xor XOR2 (N2463, N2438, N977);
buf BUF1 (N2464, N2454);
and AND2 (N2465, N2460, N1332);
nand NAND3 (N2466, N2457, N1938, N2064);
xor XOR2 (N2467, N2455, N269);
xor XOR2 (N2468, N2464, N1117);
and AND3 (N2469, N2452, N1999, N1889);
or OR2 (N2470, N2461, N268);
xor XOR2 (N2471, N2466, N2335);
or OR3 (N2472, N2442, N1788, N1180);
or OR2 (N2473, N2470, N1205);
xor XOR2 (N2474, N2472, N922);
xor XOR2 (N2475, N2463, N1720);
or OR2 (N2476, N2475, N390);
and AND2 (N2477, N2468, N1555);
buf BUF1 (N2478, N2476);
or OR3 (N2479, N2478, N1439, N2186);
nor NOR3 (N2480, N2479, N1697, N1756);
nand NAND3 (N2481, N2471, N1813, N2437);
nand NAND4 (N2482, N2467, N779, N2243, N2345);
nand NAND2 (N2483, N2465, N509);
or OR4 (N2484, N2482, N225, N463, N1788);
or OR2 (N2485, N2469, N2265);
not NOT1 (N2486, N2477);
not NOT1 (N2487, N2473);
and AND4 (N2488, N2481, N429, N519, N2183);
nor NOR4 (N2489, N2480, N2336, N1847, N198);
xor XOR2 (N2490, N2488, N1077);
xor XOR2 (N2491, N2474, N101);
xor XOR2 (N2492, N2485, N2087);
not NOT1 (N2493, N2445);
nor NOR2 (N2494, N2462, N304);
buf BUF1 (N2495, N2487);
nor NOR4 (N2496, N2494, N868, N1372, N1436);
buf BUF1 (N2497, N2484);
xor XOR2 (N2498, N2493, N268);
xor XOR2 (N2499, N2491, N1754);
buf BUF1 (N2500, N2486);
nand NAND3 (N2501, N2489, N1698, N852);
not NOT1 (N2502, N2501);
nand NAND4 (N2503, N2483, N2100, N1865, N2482);
or OR3 (N2504, N2497, N2250, N573);
nor NOR3 (N2505, N2500, N2054, N2112);
nand NAND4 (N2506, N2504, N1426, N1219, N1148);
nor NOR3 (N2507, N2506, N1113, N295);
nand NAND2 (N2508, N2492, N61);
nand NAND3 (N2509, N2502, N1588, N2123);
nor NOR2 (N2510, N2490, N401);
nand NAND2 (N2511, N2507, N1631);
buf BUF1 (N2512, N2495);
xor XOR2 (N2513, N2499, N500);
nor NOR4 (N2514, N2512, N2025, N665, N468);
and AND2 (N2515, N2509, N769);
xor XOR2 (N2516, N2513, N1451);
nand NAND2 (N2517, N2514, N1153);
not NOT1 (N2518, N2505);
or OR3 (N2519, N2503, N275, N2507);
nand NAND4 (N2520, N2498, N578, N747, N1288);
buf BUF1 (N2521, N2496);
or OR4 (N2522, N2517, N61, N93, N2336);
nor NOR4 (N2523, N2522, N264, N2227, N2325);
not NOT1 (N2524, N2519);
or OR4 (N2525, N2518, N2203, N1286, N563);
or OR2 (N2526, N2525, N2076);
or OR4 (N2527, N2521, N212, N467, N2327);
buf BUF1 (N2528, N2516);
buf BUF1 (N2529, N2511);
nand NAND2 (N2530, N2528, N1530);
not NOT1 (N2531, N2524);
nor NOR3 (N2532, N2523, N2338, N1403);
not NOT1 (N2533, N2527);
buf BUF1 (N2534, N2515);
or OR3 (N2535, N2510, N1230, N2364);
or OR2 (N2536, N2520, N1119);
xor XOR2 (N2537, N2526, N1536);
buf BUF1 (N2538, N2536);
not NOT1 (N2539, N2538);
nor NOR4 (N2540, N2537, N728, N2408, N1313);
and AND3 (N2541, N2530, N1911, N2260);
or OR4 (N2542, N2533, N2284, N995, N2194);
not NOT1 (N2543, N2542);
buf BUF1 (N2544, N2529);
or OR2 (N2545, N2531, N220);
xor XOR2 (N2546, N2532, N1546);
or OR2 (N2547, N2539, N927);
or OR4 (N2548, N2508, N1110, N429, N551);
buf BUF1 (N2549, N2543);
or OR2 (N2550, N2540, N403);
xor XOR2 (N2551, N2549, N251);
nor NOR2 (N2552, N2546, N1578);
xor XOR2 (N2553, N2541, N1477);
nand NAND3 (N2554, N2551, N2458, N1438);
buf BUF1 (N2555, N2553);
nor NOR2 (N2556, N2548, N5);
nor NOR3 (N2557, N2534, N267, N2274);
or OR2 (N2558, N2557, N858);
xor XOR2 (N2559, N2535, N1036);
buf BUF1 (N2560, N2552);
nor NOR4 (N2561, N2547, N1488, N2109, N2034);
xor XOR2 (N2562, N2555, N715);
and AND2 (N2563, N2554, N1678);
nand NAND2 (N2564, N2559, N2327);
nor NOR2 (N2565, N2550, N663);
nor NOR2 (N2566, N2560, N1429);
nand NAND3 (N2567, N2558, N1413, N633);
nand NAND3 (N2568, N2545, N163, N567);
or OR4 (N2569, N2566, N2299, N94, N837);
nor NOR4 (N2570, N2568, N2400, N1941, N745);
buf BUF1 (N2571, N2561);
and AND2 (N2572, N2556, N1422);
not NOT1 (N2573, N2572);
or OR2 (N2574, N2563, N1830);
nor NOR4 (N2575, N2564, N2085, N2514, N1926);
nor NOR4 (N2576, N2571, N1259, N1128, N528);
buf BUF1 (N2577, N2576);
not NOT1 (N2578, N2570);
and AND3 (N2579, N2562, N144, N416);
or OR4 (N2580, N2565, N1890, N223, N640);
not NOT1 (N2581, N2577);
xor XOR2 (N2582, N2575, N1044);
xor XOR2 (N2583, N2581, N1003);
not NOT1 (N2584, N2580);
buf BUF1 (N2585, N2582);
or OR4 (N2586, N2569, N780, N1813, N36);
and AND4 (N2587, N2586, N1599, N2530, N677);
nand NAND2 (N2588, N2579, N497);
nor NOR2 (N2589, N2578, N296);
nand NAND4 (N2590, N2589, N900, N152, N935);
or OR3 (N2591, N2544, N2198, N1564);
xor XOR2 (N2592, N2584, N1903);
not NOT1 (N2593, N2583);
or OR4 (N2594, N2574, N1284, N884, N1038);
xor XOR2 (N2595, N2593, N2324);
nor NOR2 (N2596, N2590, N339);
buf BUF1 (N2597, N2596);
nand NAND2 (N2598, N2588, N2225);
nor NOR2 (N2599, N2594, N2588);
not NOT1 (N2600, N2595);
xor XOR2 (N2601, N2599, N1408);
or OR2 (N2602, N2597, N2211);
and AND4 (N2603, N2600, N268, N725, N285);
nand NAND2 (N2604, N2601, N949);
xor XOR2 (N2605, N2598, N1402);
nand NAND2 (N2606, N2602, N1925);
or OR2 (N2607, N2603, N1444);
xor XOR2 (N2608, N2605, N1308);
and AND2 (N2609, N2585, N207);
buf BUF1 (N2610, N2607);
xor XOR2 (N2611, N2606, N2425);
buf BUF1 (N2612, N2610);
nand NAND3 (N2613, N2608, N1973, N1890);
nand NAND4 (N2614, N2611, N480, N132, N2075);
not NOT1 (N2615, N2609);
buf BUF1 (N2616, N2615);
nand NAND3 (N2617, N2591, N386, N669);
nand NAND2 (N2618, N2616, N989);
not NOT1 (N2619, N2567);
nand NAND4 (N2620, N2618, N548, N334, N2043);
or OR4 (N2621, N2592, N574, N608, N1103);
nand NAND3 (N2622, N2573, N2498, N1456);
nor NOR3 (N2623, N2621, N2251, N2133);
or OR2 (N2624, N2604, N1044);
not NOT1 (N2625, N2623);
or OR3 (N2626, N2625, N939, N120);
and AND4 (N2627, N2619, N381, N219, N2225);
buf BUF1 (N2628, N2613);
nand NAND3 (N2629, N2622, N1772, N1445);
nand NAND2 (N2630, N2612, N2250);
nand NAND2 (N2631, N2628, N2106);
xor XOR2 (N2632, N2587, N501);
nand NAND2 (N2633, N2614, N1327);
nor NOR4 (N2634, N2624, N2270, N2061, N1065);
and AND3 (N2635, N2630, N1951, N1365);
nand NAND3 (N2636, N2626, N1730, N291);
buf BUF1 (N2637, N2631);
buf BUF1 (N2638, N2634);
nand NAND2 (N2639, N2633, N2270);
or OR3 (N2640, N2629, N2046, N500);
not NOT1 (N2641, N2635);
nor NOR3 (N2642, N2639, N538, N368);
nand NAND2 (N2643, N2637, N1948);
xor XOR2 (N2644, N2643, N347);
nand NAND2 (N2645, N2640, N69);
nand NAND2 (N2646, N2638, N1183);
nor NOR4 (N2647, N2636, N469, N210, N2007);
and AND2 (N2648, N2647, N1492);
xor XOR2 (N2649, N2641, N953);
nor NOR4 (N2650, N2642, N1324, N1600, N1037);
buf BUF1 (N2651, N2632);
buf BUF1 (N2652, N2627);
nor NOR4 (N2653, N2644, N654, N1071, N247);
and AND3 (N2654, N2645, N1652, N2606);
or OR4 (N2655, N2654, N313, N1969, N765);
and AND4 (N2656, N2648, N485, N2165, N898);
buf BUF1 (N2657, N2617);
nor NOR2 (N2658, N2650, N1918);
or OR4 (N2659, N2652, N572, N1141, N2457);
or OR2 (N2660, N2655, N1983);
nand NAND2 (N2661, N2649, N1310);
not NOT1 (N2662, N2658);
nand NAND4 (N2663, N2660, N882, N658, N1892);
not NOT1 (N2664, N2656);
nor NOR4 (N2665, N2657, N717, N113, N2462);
nand NAND4 (N2666, N2620, N85, N1822, N494);
and AND4 (N2667, N2646, N2612, N2036, N1766);
not NOT1 (N2668, N2653);
not NOT1 (N2669, N2666);
nor NOR4 (N2670, N2651, N1963, N1915, N1943);
buf BUF1 (N2671, N2661);
or OR3 (N2672, N2667, N2502, N625);
and AND4 (N2673, N2672, N1159, N986, N1649);
or OR2 (N2674, N2669, N999);
or OR3 (N2675, N2671, N1935, N2141);
or OR3 (N2676, N2659, N2079, N1306);
or OR4 (N2677, N2676, N152, N514, N825);
nor NOR4 (N2678, N2665, N2609, N1958, N1004);
xor XOR2 (N2679, N2670, N1137);
buf BUF1 (N2680, N2663);
xor XOR2 (N2681, N2679, N2256);
nand NAND3 (N2682, N2674, N1491, N835);
or OR4 (N2683, N2662, N2616, N711, N2125);
and AND2 (N2684, N2682, N1980);
xor XOR2 (N2685, N2683, N2616);
xor XOR2 (N2686, N2681, N491);
not NOT1 (N2687, N2684);
buf BUF1 (N2688, N2668);
and AND3 (N2689, N2687, N169, N1194);
and AND4 (N2690, N2688, N1964, N867, N1273);
nand NAND2 (N2691, N2690, N690);
nor NOR3 (N2692, N2678, N93, N490);
xor XOR2 (N2693, N2677, N700);
buf BUF1 (N2694, N2693);
not NOT1 (N2695, N2680);
nand NAND3 (N2696, N2664, N172, N1393);
and AND2 (N2697, N2694, N900);
buf BUF1 (N2698, N2685);
not NOT1 (N2699, N2696);
xor XOR2 (N2700, N2692, N2035);
buf BUF1 (N2701, N2695);
nand NAND3 (N2702, N2675, N774, N370);
buf BUF1 (N2703, N2702);
or OR3 (N2704, N2701, N2632, N692);
or OR2 (N2705, N2689, N2410);
and AND4 (N2706, N2699, N520, N1341, N1340);
xor XOR2 (N2707, N2673, N2010);
not NOT1 (N2708, N2698);
or OR3 (N2709, N2705, N408, N2305);
nor NOR4 (N2710, N2707, N2209, N1422, N1977);
or OR2 (N2711, N2700, N2485);
nor NOR4 (N2712, N2706, N695, N2086, N1467);
not NOT1 (N2713, N2709);
and AND2 (N2714, N2691, N237);
buf BUF1 (N2715, N2713);
nand NAND4 (N2716, N2715, N1244, N1224, N2470);
and AND3 (N2717, N2710, N351, N251);
buf BUF1 (N2718, N2716);
buf BUF1 (N2719, N2714);
nand NAND3 (N2720, N2717, N1543, N1227);
xor XOR2 (N2721, N2719, N741);
nor NOR4 (N2722, N2721, N2231, N1859, N772);
xor XOR2 (N2723, N2720, N2401);
and AND3 (N2724, N2703, N479, N2320);
xor XOR2 (N2725, N2722, N79);
not NOT1 (N2726, N2708);
and AND2 (N2727, N2723, N1830);
nand NAND4 (N2728, N2725, N1116, N2035, N2303);
or OR3 (N2729, N2724, N1546, N1721);
buf BUF1 (N2730, N2711);
and AND2 (N2731, N2728, N272);
not NOT1 (N2732, N2712);
nor NOR3 (N2733, N2726, N982, N1749);
buf BUF1 (N2734, N2732);
or OR2 (N2735, N2686, N1571);
nor NOR4 (N2736, N2734, N962, N2445, N329);
or OR3 (N2737, N2735, N858, N1819);
nor NOR3 (N2738, N2697, N1457, N1708);
buf BUF1 (N2739, N2727);
nand NAND2 (N2740, N2737, N1763);
nor NOR3 (N2741, N2704, N1663, N1887);
buf BUF1 (N2742, N2731);
and AND2 (N2743, N2730, N822);
nand NAND4 (N2744, N2740, N2680, N84, N2475);
buf BUF1 (N2745, N2739);
or OR4 (N2746, N2733, N2723, N911, N995);
xor XOR2 (N2747, N2746, N1489);
nand NAND4 (N2748, N2747, N466, N2196, N788);
xor XOR2 (N2749, N2718, N795);
or OR3 (N2750, N2729, N492, N1249);
nor NOR4 (N2751, N2743, N896, N1118, N257);
not NOT1 (N2752, N2738);
buf BUF1 (N2753, N2751);
buf BUF1 (N2754, N2752);
and AND4 (N2755, N2741, N2300, N2003, N2058);
xor XOR2 (N2756, N2748, N2627);
buf BUF1 (N2757, N2736);
xor XOR2 (N2758, N2742, N321);
buf BUF1 (N2759, N2754);
buf BUF1 (N2760, N2758);
buf BUF1 (N2761, N2753);
nor NOR4 (N2762, N2761, N1008, N1541, N1337);
not NOT1 (N2763, N2744);
xor XOR2 (N2764, N2759, N1801);
buf BUF1 (N2765, N2764);
nor NOR2 (N2766, N2763, N2597);
and AND3 (N2767, N2750, N2697, N1611);
or OR4 (N2768, N2756, N826, N1466, N2317);
nor NOR3 (N2769, N2766, N1014, N2039);
or OR3 (N2770, N2765, N1486, N994);
and AND3 (N2771, N2769, N1916, N2726);
and AND4 (N2772, N2770, N729, N96, N908);
xor XOR2 (N2773, N2762, N625);
not NOT1 (N2774, N2772);
xor XOR2 (N2775, N2749, N2567);
nand NAND4 (N2776, N2755, N704, N1992, N494);
nand NAND4 (N2777, N2757, N1612, N2436, N760);
not NOT1 (N2778, N2776);
and AND4 (N2779, N2773, N2356, N456, N372);
or OR4 (N2780, N2778, N1909, N2000, N2330);
and AND2 (N2781, N2779, N1778);
nor NOR3 (N2782, N2767, N624, N1030);
and AND2 (N2783, N2774, N2084);
xor XOR2 (N2784, N2760, N451);
nand NAND2 (N2785, N2783, N35);
and AND3 (N2786, N2780, N1693, N2593);
or OR2 (N2787, N2771, N79);
xor XOR2 (N2788, N2782, N1818);
or OR2 (N2789, N2787, N1836);
buf BUF1 (N2790, N2786);
and AND4 (N2791, N2781, N1741, N1618, N1644);
or OR4 (N2792, N2788, N2179, N1515, N479);
xor XOR2 (N2793, N2768, N61);
and AND2 (N2794, N2775, N2538);
nand NAND3 (N2795, N2794, N1288, N545);
buf BUF1 (N2796, N2784);
nor NOR4 (N2797, N2789, N2236, N898, N2128);
not NOT1 (N2798, N2795);
nor NOR3 (N2799, N2798, N2209, N2168);
nand NAND2 (N2800, N2745, N1997);
or OR4 (N2801, N2793, N395, N87, N852);
and AND4 (N2802, N2791, N1929, N1216, N1601);
or OR2 (N2803, N2799, N190);
or OR4 (N2804, N2801, N315, N351, N2659);
buf BUF1 (N2805, N2804);
and AND2 (N2806, N2785, N1285);
and AND3 (N2807, N2802, N1374, N153);
buf BUF1 (N2808, N2797);
or OR2 (N2809, N2792, N806);
or OR2 (N2810, N2809, N413);
and AND4 (N2811, N2777, N54, N1953, N1853);
and AND4 (N2812, N2810, N183, N760, N1856);
nand NAND4 (N2813, N2805, N1182, N2460, N898);
not NOT1 (N2814, N2790);
and AND4 (N2815, N2803, N2126, N2472, N521);
and AND4 (N2816, N2800, N2208, N2144, N1750);
buf BUF1 (N2817, N2796);
xor XOR2 (N2818, N2807, N2772);
and AND4 (N2819, N2814, N2267, N2080, N1979);
nand NAND4 (N2820, N2815, N260, N1512, N511);
xor XOR2 (N2821, N2817, N739);
not NOT1 (N2822, N2808);
xor XOR2 (N2823, N2820, N1668);
not NOT1 (N2824, N2812);
or OR2 (N2825, N2811, N98);
or OR4 (N2826, N2816, N1630, N1160, N2512);
or OR3 (N2827, N2822, N1558, N1646);
buf BUF1 (N2828, N2823);
nor NOR2 (N2829, N2806, N2272);
or OR3 (N2830, N2828, N29, N2455);
xor XOR2 (N2831, N2825, N1092);
nor NOR2 (N2832, N2831, N1320);
not NOT1 (N2833, N2824);
nand NAND3 (N2834, N2813, N595, N2631);
not NOT1 (N2835, N2826);
nor NOR4 (N2836, N2835, N1326, N532, N838);
or OR2 (N2837, N2834, N1188);
nor NOR2 (N2838, N2837, N1494);
nand NAND3 (N2839, N2829, N517, N370);
nand NAND2 (N2840, N2821, N2112);
or OR4 (N2841, N2818, N1431, N254, N2522);
or OR4 (N2842, N2840, N1248, N405, N2663);
buf BUF1 (N2843, N2827);
not NOT1 (N2844, N2832);
xor XOR2 (N2845, N2833, N1498);
not NOT1 (N2846, N2836);
xor XOR2 (N2847, N2844, N1998);
nor NOR3 (N2848, N2846, N959, N784);
buf BUF1 (N2849, N2848);
xor XOR2 (N2850, N2830, N241);
not NOT1 (N2851, N2843);
nor NOR2 (N2852, N2847, N2502);
nand NAND4 (N2853, N2851, N175, N202, N188);
nand NAND4 (N2854, N2819, N1266, N2367, N1601);
or OR2 (N2855, N2838, N1252);
buf BUF1 (N2856, N2845);
xor XOR2 (N2857, N2854, N2028);
or OR2 (N2858, N2841, N240);
nor NOR3 (N2859, N2857, N2576, N1169);
buf BUF1 (N2860, N2839);
or OR2 (N2861, N2858, N1595);
not NOT1 (N2862, N2861);
nand NAND3 (N2863, N2860, N809, N1723);
or OR2 (N2864, N2853, N1497);
not NOT1 (N2865, N2855);
and AND2 (N2866, N2865, N1693);
and AND4 (N2867, N2859, N847, N1560, N1921);
and AND2 (N2868, N2850, N1758);
nand NAND4 (N2869, N2868, N2529, N267, N2111);
and AND2 (N2870, N2862, N1157);
or OR2 (N2871, N2849, N1976);
nor NOR3 (N2872, N2852, N1150, N1188);
xor XOR2 (N2873, N2856, N1704);
buf BUF1 (N2874, N2873);
xor XOR2 (N2875, N2863, N2402);
and AND3 (N2876, N2867, N1971, N633);
not NOT1 (N2877, N2869);
not NOT1 (N2878, N2864);
and AND3 (N2879, N2871, N274, N168);
or OR4 (N2880, N2875, N1688, N612, N279);
xor XOR2 (N2881, N2879, N1052);
and AND3 (N2882, N2880, N1968, N2445);
buf BUF1 (N2883, N2842);
buf BUF1 (N2884, N2882);
xor XOR2 (N2885, N2878, N1355);
and AND4 (N2886, N2881, N749, N2223, N2855);
not NOT1 (N2887, N2874);
buf BUF1 (N2888, N2870);
and AND2 (N2889, N2887, N721);
and AND4 (N2890, N2884, N1395, N2456, N2124);
not NOT1 (N2891, N2866);
nand NAND2 (N2892, N2876, N2078);
and AND2 (N2893, N2886, N175);
nand NAND4 (N2894, N2888, N2743, N420, N369);
nand NAND2 (N2895, N2872, N1995);
nand NAND4 (N2896, N2895, N1088, N1041, N2184);
nor NOR3 (N2897, N2885, N2831, N282);
nand NAND4 (N2898, N2891, N2302, N552, N1182);
nand NAND2 (N2899, N2892, N2095);
nand NAND4 (N2900, N2894, N2128, N2711, N1427);
and AND4 (N2901, N2899, N375, N683, N1945);
xor XOR2 (N2902, N2898, N1966);
xor XOR2 (N2903, N2877, N1556);
nor NOR3 (N2904, N2901, N1242, N388);
not NOT1 (N2905, N2896);
and AND3 (N2906, N2883, N2587, N340);
nand NAND2 (N2907, N2903, N1280);
and AND4 (N2908, N2890, N1309, N2261, N1222);
and AND2 (N2909, N2907, N806);
and AND4 (N2910, N2889, N918, N2426, N2613);
buf BUF1 (N2911, N2904);
or OR2 (N2912, N2905, N271);
buf BUF1 (N2913, N2909);
or OR4 (N2914, N2912, N511, N2516, N1903);
not NOT1 (N2915, N2908);
or OR4 (N2916, N2902, N603, N2483, N2113);
or OR3 (N2917, N2906, N365, N1738);
not NOT1 (N2918, N2897);
or OR3 (N2919, N2893, N1932, N160);
and AND4 (N2920, N2913, N1696, N682, N1701);
and AND3 (N2921, N2916, N1538, N1396);
nand NAND2 (N2922, N2919, N624);
not NOT1 (N2923, N2910);
xor XOR2 (N2924, N2900, N1188);
buf BUF1 (N2925, N2924);
nor NOR4 (N2926, N2914, N2880, N2613, N1679);
not NOT1 (N2927, N2920);
and AND2 (N2928, N2911, N1835);
not NOT1 (N2929, N2928);
not NOT1 (N2930, N2921);
xor XOR2 (N2931, N2927, N703);
nor NOR4 (N2932, N2926, N2125, N2896, N2390);
or OR4 (N2933, N2915, N1644, N1680, N2203);
buf BUF1 (N2934, N2917);
and AND4 (N2935, N2930, N2002, N345, N2171);
nand NAND2 (N2936, N2923, N2164);
nor NOR2 (N2937, N2935, N592);
xor XOR2 (N2938, N2937, N2937);
and AND3 (N2939, N2938, N573, N1108);
not NOT1 (N2940, N2918);
nor NOR2 (N2941, N2936, N2541);
not NOT1 (N2942, N2922);
or OR3 (N2943, N2932, N2333, N645);
nor NOR3 (N2944, N2929, N493, N2195);
xor XOR2 (N2945, N2931, N1826);
and AND4 (N2946, N2940, N222, N37, N1247);
buf BUF1 (N2947, N2945);
not NOT1 (N2948, N2944);
not NOT1 (N2949, N2939);
buf BUF1 (N2950, N2943);
and AND2 (N2951, N2942, N604);
nor NOR2 (N2952, N2948, N2011);
xor XOR2 (N2953, N2933, N2029);
nand NAND3 (N2954, N2947, N1261, N502);
not NOT1 (N2955, N2950);
and AND3 (N2956, N2955, N647, N1031);
and AND2 (N2957, N2949, N2333);
xor XOR2 (N2958, N2953, N448);
nor NOR2 (N2959, N2934, N316);
not NOT1 (N2960, N2959);
or OR4 (N2961, N2956, N1999, N1635, N229);
and AND4 (N2962, N2954, N732, N2189, N1174);
or OR2 (N2963, N2961, N471);
or OR2 (N2964, N2941, N528);
nand NAND2 (N2965, N2952, N1159);
nand NAND2 (N2966, N2963, N986);
xor XOR2 (N2967, N2964, N1611);
buf BUF1 (N2968, N2925);
and AND2 (N2969, N2968, N906);
nand NAND4 (N2970, N2957, N2876, N1252, N42);
nand NAND2 (N2971, N2958, N2853);
buf BUF1 (N2972, N2971);
nand NAND2 (N2973, N2967, N2782);
buf BUF1 (N2974, N2962);
or OR2 (N2975, N2965, N2092);
or OR2 (N2976, N2966, N2958);
and AND4 (N2977, N2970, N2241, N1841, N784);
and AND2 (N2978, N2975, N560);
nor NOR3 (N2979, N2969, N2510, N2231);
nand NAND3 (N2980, N2976, N566, N2851);
buf BUF1 (N2981, N2980);
xor XOR2 (N2982, N2973, N1383);
xor XOR2 (N2983, N2977, N1750);
xor XOR2 (N2984, N2982, N329);
nor NOR3 (N2985, N2951, N462, N2151);
and AND2 (N2986, N2960, N1860);
and AND4 (N2987, N2985, N412, N1405, N908);
nor NOR3 (N2988, N2979, N2175, N88);
xor XOR2 (N2989, N2983, N914);
nand NAND3 (N2990, N2978, N823, N2102);
or OR3 (N2991, N2988, N2807, N1031);
and AND3 (N2992, N2991, N895, N1220);
nand NAND2 (N2993, N2992, N2572);
or OR2 (N2994, N2990, N2489);
nor NOR4 (N2995, N2986, N1834, N1978, N1185);
nor NOR2 (N2996, N2995, N2350);
buf BUF1 (N2997, N2993);
nand NAND3 (N2998, N2989, N1619, N2888);
or OR3 (N2999, N2996, N2042, N1391);
nand NAND2 (N3000, N2998, N1338);
nor NOR2 (N3001, N2999, N1243);
or OR2 (N3002, N2981, N597);
and AND3 (N3003, N2946, N2099, N2853);
nand NAND2 (N3004, N2994, N600);
or OR2 (N3005, N2972, N2501);
nor NOR3 (N3006, N3003, N2344, N1899);
nor NOR4 (N3007, N2974, N466, N2150, N1045);
nor NOR3 (N3008, N2987, N2632, N1008);
buf BUF1 (N3009, N2997);
nand NAND2 (N3010, N3002, N2863);
nor NOR2 (N3011, N3010, N2503);
or OR2 (N3012, N3007, N1985);
and AND4 (N3013, N3008, N1775, N338, N2374);
or OR4 (N3014, N3006, N1199, N365, N1509);
or OR2 (N3015, N3009, N1927);
or OR2 (N3016, N3014, N1410);
not NOT1 (N3017, N3016);
xor XOR2 (N3018, N2984, N678);
xor XOR2 (N3019, N3005, N1898);
and AND4 (N3020, N3013, N2462, N293, N82);
nor NOR2 (N3021, N3012, N2875);
not NOT1 (N3022, N3004);
nand NAND4 (N3023, N3017, N1436, N855, N1658);
nand NAND3 (N3024, N3000, N252, N549);
buf BUF1 (N3025, N3021);
nor NOR4 (N3026, N3001, N2412, N2625, N78);
buf BUF1 (N3027, N3015);
xor XOR2 (N3028, N3027, N1896);
nand NAND3 (N3029, N3011, N443, N193);
and AND3 (N3030, N3019, N2030, N106);
nand NAND3 (N3031, N3023, N1612, N1596);
xor XOR2 (N3032, N3024, N2652);
not NOT1 (N3033, N3029);
buf BUF1 (N3034, N3025);
nor NOR2 (N3035, N3032, N2002);
and AND2 (N3036, N3033, N2422);
or OR2 (N3037, N3030, N551);
nor NOR3 (N3038, N3031, N1804, N349);
and AND4 (N3039, N3037, N2209, N1327, N1558);
nand NAND4 (N3040, N3036, N434, N100, N954);
buf BUF1 (N3041, N3018);
or OR3 (N3042, N3039, N976, N836);
buf BUF1 (N3043, N3034);
and AND3 (N3044, N3043, N2126, N1078);
nand NAND4 (N3045, N3040, N649, N621, N1878);
or OR2 (N3046, N3038, N1489);
nor NOR4 (N3047, N3028, N1551, N944, N1502);
and AND4 (N3048, N3022, N1506, N2204, N2029);
nor NOR4 (N3049, N3042, N3025, N1773, N1280);
and AND2 (N3050, N3046, N1935);
not NOT1 (N3051, N3041);
xor XOR2 (N3052, N3026, N1483);
xor XOR2 (N3053, N3050, N2768);
or OR3 (N3054, N3049, N471, N1216);
or OR4 (N3055, N3051, N913, N2272, N2731);
not NOT1 (N3056, N3048);
not NOT1 (N3057, N3020);
or OR2 (N3058, N3054, N911);
xor XOR2 (N3059, N3056, N1975);
and AND3 (N3060, N3055, N221, N1246);
xor XOR2 (N3061, N3058, N172);
nor NOR4 (N3062, N3053, N178, N697, N740);
nor NOR3 (N3063, N3061, N1146, N2802);
xor XOR2 (N3064, N3045, N151);
or OR3 (N3065, N3064, N2155, N1272);
nand NAND4 (N3066, N3060, N1663, N1452, N1195);
nand NAND3 (N3067, N3059, N1169, N149);
buf BUF1 (N3068, N3052);
nand NAND3 (N3069, N3062, N1978, N1197);
nand NAND4 (N3070, N3057, N1383, N245, N1166);
nand NAND3 (N3071, N3068, N299, N1059);
nor NOR3 (N3072, N3071, N163, N507);
nor NOR2 (N3073, N3070, N1283);
or OR3 (N3074, N3067, N1080, N1004);
nand NAND4 (N3075, N3065, N2326, N964, N2313);
nor NOR3 (N3076, N3073, N2697, N1245);
not NOT1 (N3077, N3076);
or OR3 (N3078, N3047, N2987, N2376);
or OR2 (N3079, N3044, N3067);
or OR2 (N3080, N3069, N18);
or OR4 (N3081, N3075, N1850, N240, N2604);
buf BUF1 (N3082, N3074);
buf BUF1 (N3083, N3082);
or OR2 (N3084, N3066, N686);
nor NOR3 (N3085, N3080, N1635, N2891);
xor XOR2 (N3086, N3063, N2754);
xor XOR2 (N3087, N3078, N2737);
buf BUF1 (N3088, N3079);
and AND2 (N3089, N3087, N1283);
or OR2 (N3090, N3086, N434);
nor NOR3 (N3091, N3077, N238, N1757);
buf BUF1 (N3092, N3083);
buf BUF1 (N3093, N3085);
not NOT1 (N3094, N3090);
or OR3 (N3095, N3091, N659, N2449);
nand NAND2 (N3096, N3088, N64);
buf BUF1 (N3097, N3093);
not NOT1 (N3098, N3096);
or OR2 (N3099, N3094, N1806);
not NOT1 (N3100, N3099);
nand NAND3 (N3101, N3035, N1624, N1185);
xor XOR2 (N3102, N3100, N1135);
nor NOR2 (N3103, N3072, N2187);
nand NAND4 (N3104, N3098, N2585, N1685, N2391);
nand NAND3 (N3105, N3097, N1716, N1464);
not NOT1 (N3106, N3084);
not NOT1 (N3107, N3095);
not NOT1 (N3108, N3107);
buf BUF1 (N3109, N3108);
nand NAND2 (N3110, N3109, N3049);
buf BUF1 (N3111, N3104);
buf BUF1 (N3112, N3105);
nand NAND4 (N3113, N3111, N1094, N1025, N1228);
buf BUF1 (N3114, N3102);
or OR4 (N3115, N3113, N2456, N1076, N294);
or OR3 (N3116, N3101, N754, N1029);
nor NOR4 (N3117, N3112, N1324, N1921, N2934);
buf BUF1 (N3118, N3116);
or OR3 (N3119, N3103, N476, N82);
buf BUF1 (N3120, N3092);
and AND4 (N3121, N3119, N324, N2370, N1805);
nor NOR2 (N3122, N3089, N688);
and AND4 (N3123, N3110, N1014, N1925, N519);
nor NOR2 (N3124, N3114, N2015);
xor XOR2 (N3125, N3106, N1246);
nor NOR4 (N3126, N3081, N2264, N1538, N1031);
nor NOR2 (N3127, N3123, N600);
not NOT1 (N3128, N3126);
nand NAND3 (N3129, N3125, N574, N2772);
nand NAND2 (N3130, N3121, N2468);
or OR3 (N3131, N3118, N217, N1219);
and AND4 (N3132, N3131, N3098, N2448, N269);
nor NOR2 (N3133, N3132, N2810);
or OR3 (N3134, N3117, N1385, N1231);
and AND4 (N3135, N3134, N1186, N1888, N211);
nand NAND4 (N3136, N3130, N750, N1262, N2290);
not NOT1 (N3137, N3115);
or OR2 (N3138, N3136, N2756);
nand NAND4 (N3139, N3120, N2102, N2775, N2024);
or OR3 (N3140, N3127, N2430, N2813);
and AND3 (N3141, N3137, N2675, N713);
nand NAND3 (N3142, N3135, N1660, N237);
or OR3 (N3143, N3122, N2394, N1899);
nor NOR2 (N3144, N3141, N33);
not NOT1 (N3145, N3143);
not NOT1 (N3146, N3144);
nor NOR4 (N3147, N3128, N1947, N1581, N1021);
and AND3 (N3148, N3140, N666, N2363);
buf BUF1 (N3149, N3146);
not NOT1 (N3150, N3133);
nor NOR4 (N3151, N3139, N1492, N2950, N1538);
not NOT1 (N3152, N3151);
or OR2 (N3153, N3148, N2976);
or OR3 (N3154, N3138, N987, N643);
and AND4 (N3155, N3147, N1239, N2906, N798);
xor XOR2 (N3156, N3152, N2067);
xor XOR2 (N3157, N3153, N2217);
or OR2 (N3158, N3124, N2333);
xor XOR2 (N3159, N3158, N680);
nor NOR3 (N3160, N3145, N307, N2210);
not NOT1 (N3161, N3150);
nand NAND3 (N3162, N3142, N1688, N1930);
not NOT1 (N3163, N3161);
or OR2 (N3164, N3162, N2990);
not NOT1 (N3165, N3129);
nand NAND2 (N3166, N3159, N2179);
nand NAND3 (N3167, N3155, N1101, N1471);
not NOT1 (N3168, N3154);
nand NAND3 (N3169, N3157, N93, N2644);
not NOT1 (N3170, N3156);
or OR4 (N3171, N3170, N1963, N653, N2622);
not NOT1 (N3172, N3163);
nor NOR2 (N3173, N3167, N345);
nor NOR2 (N3174, N3166, N602);
nand NAND3 (N3175, N3168, N2110, N2024);
buf BUF1 (N3176, N3149);
or OR2 (N3177, N3169, N124);
nand NAND3 (N3178, N3175, N2150, N1140);
xor XOR2 (N3179, N3165, N65);
nand NAND4 (N3180, N3172, N1122, N1485, N1867);
xor XOR2 (N3181, N3173, N2416);
and AND3 (N3182, N3179, N270, N2681);
not NOT1 (N3183, N3181);
not NOT1 (N3184, N3174);
nor NOR3 (N3185, N3184, N1401, N2241);
nor NOR3 (N3186, N3164, N2346, N2473);
xor XOR2 (N3187, N3171, N2923);
not NOT1 (N3188, N3160);
buf BUF1 (N3189, N3180);
buf BUF1 (N3190, N3182);
nor NOR3 (N3191, N3176, N804, N2480);
nand NAND2 (N3192, N3186, N1168);
not NOT1 (N3193, N3192);
xor XOR2 (N3194, N3183, N2971);
not NOT1 (N3195, N3189);
not NOT1 (N3196, N3177);
or OR3 (N3197, N3193, N2964, N746);
and AND4 (N3198, N3178, N1889, N2569, N1593);
or OR2 (N3199, N3190, N2384);
or OR2 (N3200, N3187, N653);
nor NOR3 (N3201, N3185, N2136, N2263);
not NOT1 (N3202, N3197);
nor NOR4 (N3203, N3200, N2149, N2183, N3030);
buf BUF1 (N3204, N3194);
nand NAND2 (N3205, N3201, N151);
nand NAND4 (N3206, N3205, N1103, N831, N2931);
and AND2 (N3207, N3203, N2222);
or OR4 (N3208, N3199, N747, N2637, N1900);
buf BUF1 (N3209, N3207);
nand NAND3 (N3210, N3209, N2624, N159);
nor NOR4 (N3211, N3208, N1146, N1066, N1505);
nand NAND2 (N3212, N3211, N722);
nor NOR3 (N3213, N3191, N634, N2243);
buf BUF1 (N3214, N3202);
or OR3 (N3215, N3188, N2224, N2285);
nand NAND4 (N3216, N3198, N1179, N1777, N1774);
buf BUF1 (N3217, N3216);
not NOT1 (N3218, N3215);
buf BUF1 (N3219, N3195);
nor NOR3 (N3220, N3196, N1895, N36);
not NOT1 (N3221, N3213);
not NOT1 (N3222, N3218);
or OR2 (N3223, N3219, N989);
not NOT1 (N3224, N3221);
or OR2 (N3225, N3222, N2505);
not NOT1 (N3226, N3210);
xor XOR2 (N3227, N3224, N2533);
or OR3 (N3228, N3214, N1392, N17);
nor NOR3 (N3229, N3226, N639, N1511);
buf BUF1 (N3230, N3206);
or OR3 (N3231, N3229, N2698, N617);
and AND3 (N3232, N3230, N2579, N745);
and AND3 (N3233, N3227, N1975, N3230);
not NOT1 (N3234, N3217);
nor NOR3 (N3235, N3231, N1097, N2902);
xor XOR2 (N3236, N3235, N342);
buf BUF1 (N3237, N3233);
or OR4 (N3238, N3236, N2021, N2844, N1880);
not NOT1 (N3239, N3225);
xor XOR2 (N3240, N3234, N3192);
buf BUF1 (N3241, N3238);
xor XOR2 (N3242, N3204, N1862);
buf BUF1 (N3243, N3232);
xor XOR2 (N3244, N3223, N3006);
not NOT1 (N3245, N3243);
nand NAND2 (N3246, N3212, N3144);
or OR2 (N3247, N3241, N38);
nor NOR3 (N3248, N3246, N2516, N1383);
not NOT1 (N3249, N3242);
nor NOR3 (N3250, N3228, N962, N1061);
nand NAND2 (N3251, N3220, N1705);
and AND2 (N3252, N3251, N1368);
buf BUF1 (N3253, N3237);
xor XOR2 (N3254, N3248, N2537);
nor NOR3 (N3255, N3244, N3004, N1296);
not NOT1 (N3256, N3255);
nor NOR4 (N3257, N3245, N1808, N1825, N439);
or OR2 (N3258, N3253, N1802);
buf BUF1 (N3259, N3254);
buf BUF1 (N3260, N3239);
nor NOR4 (N3261, N3249, N220, N2591, N404);
nor NOR4 (N3262, N3256, N2207, N3169, N2305);
not NOT1 (N3263, N3261);
buf BUF1 (N3264, N3262);
nand NAND4 (N3265, N3263, N727, N486, N2531);
and AND4 (N3266, N3240, N998, N1422, N1766);
nor NOR3 (N3267, N3252, N803, N2819);
nor NOR4 (N3268, N3266, N981, N2615, N1985);
or OR4 (N3269, N3250, N1873, N2917, N1079);
xor XOR2 (N3270, N3265, N211);
not NOT1 (N3271, N3264);
not NOT1 (N3272, N3258);
or OR3 (N3273, N3260, N3176, N2817);
xor XOR2 (N3274, N3269, N374);
or OR2 (N3275, N3257, N2922);
nand NAND4 (N3276, N3268, N2581, N1527, N173);
nor NOR3 (N3277, N3274, N2196, N3084);
nand NAND2 (N3278, N3272, N412);
nor NOR3 (N3279, N3277, N1335, N873);
buf BUF1 (N3280, N3267);
buf BUF1 (N3281, N3259);
not NOT1 (N3282, N3281);
nor NOR3 (N3283, N3271, N3226, N649);
and AND4 (N3284, N3247, N2354, N506, N1501);
nand NAND3 (N3285, N3279, N2579, N1374);
not NOT1 (N3286, N3283);
or OR4 (N3287, N3282, N625, N895, N1436);
nor NOR2 (N3288, N3273, N2719);
not NOT1 (N3289, N3285);
nand NAND3 (N3290, N3270, N931, N1366);
and AND3 (N3291, N3276, N2026, N1592);
not NOT1 (N3292, N3286);
or OR3 (N3293, N3291, N3027, N1330);
not NOT1 (N3294, N3280);
xor XOR2 (N3295, N3290, N2601);
buf BUF1 (N3296, N3288);
nand NAND3 (N3297, N3287, N152, N2432);
not NOT1 (N3298, N3278);
xor XOR2 (N3299, N3297, N1972);
nand NAND3 (N3300, N3298, N1456, N308);
or OR3 (N3301, N3296, N849, N351);
and AND2 (N3302, N3294, N391);
not NOT1 (N3303, N3284);
or OR2 (N3304, N3300, N1881);
xor XOR2 (N3305, N3295, N688);
not NOT1 (N3306, N3302);
not NOT1 (N3307, N3301);
or OR2 (N3308, N3306, N1503);
not NOT1 (N3309, N3292);
nand NAND3 (N3310, N3307, N2976, N2472);
not NOT1 (N3311, N3309);
buf BUF1 (N3312, N3303);
nor NOR4 (N3313, N3308, N756, N2298, N3299);
and AND4 (N3314, N1994, N63, N2988, N3041);
nor NOR3 (N3315, N3313, N1391, N3194);
buf BUF1 (N3316, N3314);
not NOT1 (N3317, N3289);
buf BUF1 (N3318, N3311);
buf BUF1 (N3319, N3275);
buf BUF1 (N3320, N3317);
nor NOR3 (N3321, N3315, N2283, N2614);
xor XOR2 (N3322, N3320, N803);
not NOT1 (N3323, N3319);
nand NAND4 (N3324, N3318, N3312, N470, N2055);
or OR4 (N3325, N1857, N2657, N581, N159);
buf BUF1 (N3326, N3323);
nor NOR4 (N3327, N3305, N3169, N1623, N2369);
nor NOR4 (N3328, N3322, N285, N3177, N2705);
and AND2 (N3329, N3316, N362);
not NOT1 (N3330, N3304);
not NOT1 (N3331, N3327);
not NOT1 (N3332, N3330);
nand NAND4 (N3333, N3324, N911, N627, N2149);
xor XOR2 (N3334, N3332, N2161);
buf BUF1 (N3335, N3325);
xor XOR2 (N3336, N3333, N2077);
buf BUF1 (N3337, N3328);
nand NAND4 (N3338, N3336, N2196, N3231, N2046);
not NOT1 (N3339, N3337);
or OR3 (N3340, N3293, N2275, N1497);
or OR2 (N3341, N3334, N3135);
nor NOR4 (N3342, N3341, N2153, N2520, N604);
nand NAND3 (N3343, N3340, N852, N2178);
not NOT1 (N3344, N3310);
or OR3 (N3345, N3321, N2197, N2571);
or OR2 (N3346, N3345, N1377);
nor NOR2 (N3347, N3331, N601);
nor NOR3 (N3348, N3347, N2098, N2995);
or OR4 (N3349, N3338, N1656, N600, N1293);
and AND3 (N3350, N3344, N2816, N1910);
nand NAND4 (N3351, N3329, N2537, N1688, N508);
not NOT1 (N3352, N3346);
buf BUF1 (N3353, N3335);
nor NOR3 (N3354, N3326, N2504, N1757);
and AND2 (N3355, N3352, N2148);
xor XOR2 (N3356, N3354, N2471);
xor XOR2 (N3357, N3343, N2362);
nor NOR4 (N3358, N3342, N1981, N1023, N1145);
or OR4 (N3359, N3353, N1881, N317, N2237);
nor NOR4 (N3360, N3339, N1576, N1090, N424);
buf BUF1 (N3361, N3359);
nor NOR2 (N3362, N3357, N3173);
and AND3 (N3363, N3355, N3215, N1981);
buf BUF1 (N3364, N3361);
nor NOR3 (N3365, N3363, N3035, N827);
or OR2 (N3366, N3364, N2697);
nand NAND3 (N3367, N3351, N239, N169);
nor NOR3 (N3368, N3362, N3224, N2729);
not NOT1 (N3369, N3367);
xor XOR2 (N3370, N3368, N2476);
not NOT1 (N3371, N3350);
not NOT1 (N3372, N3360);
and AND3 (N3373, N3348, N2452, N2682);
nand NAND2 (N3374, N3370, N2318);
and AND3 (N3375, N3366, N2525, N121);
nor NOR2 (N3376, N3371, N991);
nor NOR4 (N3377, N3376, N1775, N376, N2226);
not NOT1 (N3378, N3356);
and AND3 (N3379, N3374, N932, N1062);
and AND3 (N3380, N3349, N597, N2194);
nor NOR2 (N3381, N3380, N2296);
not NOT1 (N3382, N3377);
xor XOR2 (N3383, N3372, N1900);
xor XOR2 (N3384, N3358, N372);
or OR2 (N3385, N3382, N856);
xor XOR2 (N3386, N3365, N2287);
not NOT1 (N3387, N3373);
xor XOR2 (N3388, N3378, N366);
or OR3 (N3389, N3383, N2700, N2610);
or OR3 (N3390, N3369, N646, N1313);
or OR4 (N3391, N3386, N1395, N1834, N763);
not NOT1 (N3392, N3385);
not NOT1 (N3393, N3391);
and AND2 (N3394, N3392, N2265);
nand NAND2 (N3395, N3387, N774);
and AND3 (N3396, N3389, N2792, N2143);
or OR4 (N3397, N3388, N1261, N1803, N771);
nor NOR2 (N3398, N3396, N1549);
nor NOR2 (N3399, N3395, N1355);
or OR2 (N3400, N3393, N2374);
nand NAND4 (N3401, N3379, N2582, N1761, N1502);
buf BUF1 (N3402, N3390);
and AND3 (N3403, N3384, N3139, N1765);
buf BUF1 (N3404, N3375);
not NOT1 (N3405, N3401);
buf BUF1 (N3406, N3404);
not NOT1 (N3407, N3406);
or OR4 (N3408, N3407, N377, N1815, N1525);
xor XOR2 (N3409, N3398, N2732);
nand NAND4 (N3410, N3403, N2104, N3154, N3239);
nor NOR3 (N3411, N3394, N1908, N799);
buf BUF1 (N3412, N3411);
or OR3 (N3413, N3405, N2053, N2468);
not NOT1 (N3414, N3410);
nand NAND3 (N3415, N3409, N3413, N1750);
xor XOR2 (N3416, N2103, N243);
buf BUF1 (N3417, N3408);
nor NOR2 (N3418, N3416, N493);
or OR4 (N3419, N3402, N2926, N785, N1350);
and AND4 (N3420, N3397, N84, N810, N1684);
or OR2 (N3421, N3399, N1084);
and AND3 (N3422, N3419, N2389, N3102);
nor NOR4 (N3423, N3421, N3027, N2088, N2568);
buf BUF1 (N3424, N3412);
xor XOR2 (N3425, N3400, N1105);
not NOT1 (N3426, N3425);
not NOT1 (N3427, N3423);
or OR4 (N3428, N3427, N3382, N2977, N214);
and AND4 (N3429, N3426, N3394, N934, N1651);
and AND4 (N3430, N3417, N186, N531, N3205);
buf BUF1 (N3431, N3415);
nor NOR2 (N3432, N3431, N2681);
and AND2 (N3433, N3414, N1337);
xor XOR2 (N3434, N3429, N2338);
xor XOR2 (N3435, N3432, N2226);
not NOT1 (N3436, N3424);
nor NOR2 (N3437, N3381, N3180);
nand NAND3 (N3438, N3437, N1976, N3266);
buf BUF1 (N3439, N3420);
nand NAND4 (N3440, N3430, N791, N18, N1543);
or OR4 (N3441, N3436, N973, N2612, N2637);
nor NOR2 (N3442, N3440, N2619);
and AND4 (N3443, N3439, N1658, N2200, N1795);
or OR3 (N3444, N3435, N257, N1647);
nor NOR4 (N3445, N3441, N1853, N642, N2132);
xor XOR2 (N3446, N3422, N1806);
not NOT1 (N3447, N3428);
nor NOR3 (N3448, N3433, N2519, N324);
nor NOR3 (N3449, N3434, N618, N1610);
xor XOR2 (N3450, N3445, N2892);
nand NAND3 (N3451, N3443, N3021, N831);
xor XOR2 (N3452, N3442, N668);
or OR4 (N3453, N3452, N3373, N2964, N1879);
buf BUF1 (N3454, N3449);
nor NOR2 (N3455, N3448, N225);
nor NOR2 (N3456, N3450, N2372);
nand NAND4 (N3457, N3438, N2245, N3316, N2991);
buf BUF1 (N3458, N3451);
nand NAND3 (N3459, N3458, N2331, N3016);
buf BUF1 (N3460, N3454);
nor NOR2 (N3461, N3447, N1923);
xor XOR2 (N3462, N3459, N2216);
nand NAND4 (N3463, N3460, N406, N2143, N1358);
not NOT1 (N3464, N3455);
and AND2 (N3465, N3464, N2152);
or OR2 (N3466, N3456, N136);
nor NOR4 (N3467, N3463, N1471, N2800, N1);
xor XOR2 (N3468, N3466, N2696);
xor XOR2 (N3469, N3467, N1923);
nor NOR4 (N3470, N3469, N2633, N648, N3039);
xor XOR2 (N3471, N3446, N711);
nand NAND3 (N3472, N3453, N1001, N1467);
nor NOR3 (N3473, N3468, N648, N3111);
and AND4 (N3474, N3473, N1985, N1725, N934);
buf BUF1 (N3475, N3461);
nor NOR4 (N3476, N3470, N2922, N2333, N2271);
nor NOR3 (N3477, N3471, N2043, N2881);
or OR4 (N3478, N3474, N1668, N3355, N260);
xor XOR2 (N3479, N3475, N2090);
buf BUF1 (N3480, N3465);
and AND4 (N3481, N3418, N924, N1463, N1493);
or OR2 (N3482, N3472, N1507);
nor NOR4 (N3483, N3477, N1798, N3300, N2884);
or OR3 (N3484, N3483, N1970, N331);
xor XOR2 (N3485, N3444, N368);
buf BUF1 (N3486, N3457);
buf BUF1 (N3487, N3478);
nand NAND3 (N3488, N3485, N1368, N2354);
and AND2 (N3489, N3476, N603);
not NOT1 (N3490, N3487);
nand NAND2 (N3491, N3486, N2920);
not NOT1 (N3492, N3489);
not NOT1 (N3493, N3491);
nor NOR4 (N3494, N3488, N114, N1617, N1799);
nand NAND4 (N3495, N3481, N3199, N2505, N77);
buf BUF1 (N3496, N3462);
or OR2 (N3497, N3492, N1227);
nand NAND2 (N3498, N3490, N3122);
or OR3 (N3499, N3484, N3136, N1275);
nor NOR2 (N3500, N3497, N1581);
buf BUF1 (N3501, N3496);
not NOT1 (N3502, N3479);
nand NAND2 (N3503, N3494, N3000);
nor NOR2 (N3504, N3501, N365);
not NOT1 (N3505, N3495);
nor NOR2 (N3506, N3500, N3211);
and AND4 (N3507, N3482, N1106, N2303, N2218);
nor NOR4 (N3508, N3480, N2275, N628, N1968);
not NOT1 (N3509, N3498);
or OR2 (N3510, N3506, N3327);
buf BUF1 (N3511, N3504);
nand NAND4 (N3512, N3511, N3252, N2036, N2465);
xor XOR2 (N3513, N3505, N1138);
buf BUF1 (N3514, N3512);
xor XOR2 (N3515, N3509, N147);
or OR3 (N3516, N3513, N3232, N187);
not NOT1 (N3517, N3516);
xor XOR2 (N3518, N3510, N2995);
nor NOR4 (N3519, N3518, N2493, N1484, N323);
not NOT1 (N3520, N3493);
nand NAND3 (N3521, N3502, N687, N1300);
nand NAND4 (N3522, N3508, N1652, N551, N1284);
nor NOR4 (N3523, N3499, N907, N2760, N1635);
nor NOR2 (N3524, N3515, N1686);
not NOT1 (N3525, N3522);
and AND4 (N3526, N3523, N86, N31, N973);
buf BUF1 (N3527, N3503);
not NOT1 (N3528, N3519);
xor XOR2 (N3529, N3507, N1398);
nand NAND2 (N3530, N3526, N1925);
buf BUF1 (N3531, N3520);
not NOT1 (N3532, N3521);
nor NOR2 (N3533, N3531, N577);
not NOT1 (N3534, N3514);
xor XOR2 (N3535, N3524, N849);
buf BUF1 (N3536, N3517);
buf BUF1 (N3537, N3527);
and AND3 (N3538, N3529, N2786, N3429);
and AND4 (N3539, N3537, N2374, N1253, N37);
nor NOR3 (N3540, N3528, N1137, N2513);
nor NOR2 (N3541, N3532, N735);
not NOT1 (N3542, N3525);
nor NOR3 (N3543, N3539, N138, N39);
nand NAND4 (N3544, N3530, N3533, N826, N2876);
nand NAND2 (N3545, N1507, N935);
and AND3 (N3546, N3541, N2302, N1760);
nor NOR4 (N3547, N3544, N3482, N1291, N1800);
and AND3 (N3548, N3536, N2728, N2638);
nand NAND2 (N3549, N3542, N686);
or OR4 (N3550, N3534, N505, N1689, N1986);
or OR4 (N3551, N3547, N1257, N3454, N1234);
and AND3 (N3552, N3538, N3401, N3119);
nor NOR4 (N3553, N3549, N619, N1625, N371);
nand NAND2 (N3554, N3551, N2870);
and AND2 (N3555, N3535, N1207);
and AND3 (N3556, N3545, N2290, N2969);
or OR2 (N3557, N3543, N432);
or OR4 (N3558, N3546, N3021, N492, N1915);
or OR2 (N3559, N3548, N1375);
xor XOR2 (N3560, N3556, N1728);
nand NAND2 (N3561, N3557, N64);
nor NOR2 (N3562, N3552, N644);
buf BUF1 (N3563, N3560);
and AND2 (N3564, N3554, N2968);
or OR2 (N3565, N3540, N449);
buf BUF1 (N3566, N3562);
nor NOR4 (N3567, N3555, N1295, N2242, N9);
nand NAND4 (N3568, N3561, N2646, N124, N2357);
not NOT1 (N3569, N3558);
not NOT1 (N3570, N3553);
buf BUF1 (N3571, N3559);
nand NAND4 (N3572, N3563, N670, N3233, N1793);
not NOT1 (N3573, N3564);
xor XOR2 (N3574, N3573, N1648);
and AND4 (N3575, N3567, N2294, N657, N499);
not NOT1 (N3576, N3566);
nor NOR4 (N3577, N3575, N632, N813, N2018);
buf BUF1 (N3578, N3571);
and AND2 (N3579, N3570, N370);
not NOT1 (N3580, N3569);
xor XOR2 (N3581, N3579, N1811);
nand NAND3 (N3582, N3578, N37, N2236);
xor XOR2 (N3583, N3574, N2295);
nor NOR4 (N3584, N3581, N426, N1422, N13);
nand NAND3 (N3585, N3565, N3539, N1824);
nand NAND4 (N3586, N3580, N2405, N1560, N2648);
buf BUF1 (N3587, N3572);
not NOT1 (N3588, N3568);
not NOT1 (N3589, N3588);
not NOT1 (N3590, N3584);
or OR3 (N3591, N3583, N2468, N1223);
and AND3 (N3592, N3582, N2389, N2893);
not NOT1 (N3593, N3589);
nand NAND2 (N3594, N3585, N1106);
nor NOR4 (N3595, N3576, N211, N639, N696);
nor NOR3 (N3596, N3590, N2541, N54);
nor NOR2 (N3597, N3596, N139);
and AND2 (N3598, N3594, N1793);
not NOT1 (N3599, N3591);
and AND4 (N3600, N3593, N929, N3367, N3252);
xor XOR2 (N3601, N3586, N2778);
buf BUF1 (N3602, N3598);
or OR3 (N3603, N3599, N219, N1255);
nand NAND3 (N3604, N3597, N3130, N3495);
nand NAND4 (N3605, N3604, N498, N848, N566);
nand NAND3 (N3606, N3577, N372, N3585);
not NOT1 (N3607, N3601);
not NOT1 (N3608, N3600);
and AND4 (N3609, N3602, N2009, N1437, N2342);
or OR2 (N3610, N3592, N1817);
nand NAND4 (N3611, N3550, N2766, N1455, N1321);
buf BUF1 (N3612, N3608);
and AND3 (N3613, N3610, N990, N3291);
xor XOR2 (N3614, N3609, N3199);
nand NAND3 (N3615, N3614, N1395, N3007);
and AND4 (N3616, N3613, N254, N2817, N2431);
xor XOR2 (N3617, N3607, N1800);
not NOT1 (N3618, N3616);
nor NOR2 (N3619, N3615, N570);
xor XOR2 (N3620, N3605, N530);
xor XOR2 (N3621, N3618, N327);
xor XOR2 (N3622, N3611, N2564);
or OR3 (N3623, N3603, N3619, N1752);
xor XOR2 (N3624, N1273, N3580);
nand NAND3 (N3625, N3595, N3537, N534);
nor NOR2 (N3626, N3623, N2047);
nor NOR3 (N3627, N3622, N2490, N244);
or OR2 (N3628, N3625, N937);
nor NOR3 (N3629, N3624, N306, N2883);
nor NOR2 (N3630, N3587, N3392);
nand NAND2 (N3631, N3612, N221);
xor XOR2 (N3632, N3628, N496);
nand NAND3 (N3633, N3620, N2451, N3529);
or OR4 (N3634, N3621, N161, N1546, N880);
buf BUF1 (N3635, N3633);
nand NAND3 (N3636, N3631, N2582, N916);
not NOT1 (N3637, N3629);
not NOT1 (N3638, N3637);
nand NAND2 (N3639, N3635, N2823);
or OR4 (N3640, N3634, N2117, N466, N371);
or OR3 (N3641, N3630, N827, N2543);
buf BUF1 (N3642, N3627);
xor XOR2 (N3643, N3638, N752);
buf BUF1 (N3644, N3606);
nor NOR2 (N3645, N3643, N491);
nand NAND3 (N3646, N3641, N2646, N2634);
and AND4 (N3647, N3632, N1826, N268, N2090);
nand NAND4 (N3648, N3644, N622, N729, N1763);
buf BUF1 (N3649, N3646);
and AND4 (N3650, N3617, N3091, N2600, N3514);
not NOT1 (N3651, N3648);
and AND4 (N3652, N3651, N892, N3496, N2931);
xor XOR2 (N3653, N3636, N1929);
nor NOR2 (N3654, N3640, N2989);
nor NOR3 (N3655, N3650, N2316, N3067);
or OR2 (N3656, N3645, N2826);
not NOT1 (N3657, N3655);
or OR2 (N3658, N3657, N3425);
nor NOR2 (N3659, N3639, N2582);
xor XOR2 (N3660, N3642, N2036);
nand NAND2 (N3661, N3656, N2561);
buf BUF1 (N3662, N3647);
nand NAND4 (N3663, N3658, N3046, N2418, N658);
not NOT1 (N3664, N3649);
buf BUF1 (N3665, N3652);
buf BUF1 (N3666, N3626);
nand NAND4 (N3667, N3665, N2460, N2030, N1110);
and AND4 (N3668, N3659, N46, N2086, N1917);
nand NAND2 (N3669, N3654, N742);
nor NOR4 (N3670, N3664, N6, N2040, N2082);
buf BUF1 (N3671, N3669);
and AND2 (N3672, N3670, N1716);
not NOT1 (N3673, N3663);
buf BUF1 (N3674, N3667);
nor NOR2 (N3675, N3661, N1609);
nand NAND4 (N3676, N3672, N1461, N3545, N960);
xor XOR2 (N3677, N3653, N683);
not NOT1 (N3678, N3676);
not NOT1 (N3679, N3674);
not NOT1 (N3680, N3678);
nand NAND4 (N3681, N3666, N2577, N337, N2679);
or OR2 (N3682, N3668, N3108);
buf BUF1 (N3683, N3681);
and AND4 (N3684, N3673, N1513, N3572, N913);
nand NAND2 (N3685, N3679, N928);
xor XOR2 (N3686, N3662, N2021);
or OR3 (N3687, N3671, N2683, N575);
or OR3 (N3688, N3684, N2630, N2779);
xor XOR2 (N3689, N3680, N871);
xor XOR2 (N3690, N3683, N1527);
xor XOR2 (N3691, N3690, N2730);
and AND3 (N3692, N3675, N1845, N1383);
or OR2 (N3693, N3688, N3045);
nor NOR3 (N3694, N3677, N639, N3434);
or OR4 (N3695, N3693, N3227, N1331, N77);
nand NAND2 (N3696, N3660, N227);
and AND4 (N3697, N3694, N1433, N2334, N3477);
or OR2 (N3698, N3682, N298);
or OR4 (N3699, N3686, N3473, N3059, N64);
nand NAND2 (N3700, N3696, N2538);
buf BUF1 (N3701, N3698);
nand NAND3 (N3702, N3692, N3614, N2130);
nand NAND2 (N3703, N3699, N1297);
or OR3 (N3704, N3691, N789, N2369);
nor NOR4 (N3705, N3702, N478, N1896, N3099);
and AND2 (N3706, N3703, N3084);
nand NAND3 (N3707, N3695, N1706, N2592);
or OR2 (N3708, N3706, N1219);
and AND3 (N3709, N3707, N2637, N1281);
buf BUF1 (N3710, N3687);
xor XOR2 (N3711, N3710, N334);
not NOT1 (N3712, N3697);
buf BUF1 (N3713, N3708);
buf BUF1 (N3714, N3713);
xor XOR2 (N3715, N3700, N1545);
not NOT1 (N3716, N3704);
nor NOR4 (N3717, N3712, N3020, N465, N1681);
xor XOR2 (N3718, N3685, N920);
buf BUF1 (N3719, N3716);
xor XOR2 (N3720, N3701, N88);
not NOT1 (N3721, N3705);
xor XOR2 (N3722, N3689, N302);
nand NAND3 (N3723, N3722, N2978, N1332);
xor XOR2 (N3724, N3709, N338);
nor NOR2 (N3725, N3717, N1843);
nand NAND3 (N3726, N3711, N3658, N1879);
nand NAND4 (N3727, N3714, N3492, N197, N2199);
buf BUF1 (N3728, N3726);
or OR3 (N3729, N3724, N144, N2884);
buf BUF1 (N3730, N3727);
and AND4 (N3731, N3729, N3642, N3287, N953);
and AND2 (N3732, N3721, N3703);
not NOT1 (N3733, N3720);
nand NAND4 (N3734, N3730, N34, N3472, N1135);
xor XOR2 (N3735, N3733, N3627);
and AND4 (N3736, N3728, N661, N2032, N3516);
and AND3 (N3737, N3732, N1319, N1051);
and AND4 (N3738, N3718, N2638, N765, N2369);
xor XOR2 (N3739, N3725, N1952);
or OR2 (N3740, N3738, N3295);
not NOT1 (N3741, N3740);
nand NAND2 (N3742, N3719, N3582);
and AND3 (N3743, N3735, N2293, N1764);
or OR3 (N3744, N3739, N3158, N72);
buf BUF1 (N3745, N3743);
or OR3 (N3746, N3745, N1938, N2652);
nor NOR2 (N3747, N3746, N2098);
or OR2 (N3748, N3744, N609);
and AND2 (N3749, N3734, N1266);
or OR2 (N3750, N3715, N3621);
nand NAND2 (N3751, N3750, N3262);
not NOT1 (N3752, N3749);
xor XOR2 (N3753, N3752, N2188);
nor NOR4 (N3754, N3753, N2344, N565, N1638);
and AND4 (N3755, N3754, N1796, N2515, N2112);
and AND4 (N3756, N3737, N1956, N833, N1399);
and AND4 (N3757, N3751, N1154, N1210, N292);
buf BUF1 (N3758, N3736);
or OR2 (N3759, N3756, N2655);
buf BUF1 (N3760, N3741);
nand NAND4 (N3761, N3723, N3209, N2370, N69);
not NOT1 (N3762, N3761);
xor XOR2 (N3763, N3758, N3620);
not NOT1 (N3764, N3742);
buf BUF1 (N3765, N3748);
or OR3 (N3766, N3755, N1660, N1713);
nand NAND3 (N3767, N3764, N3122, N2161);
and AND4 (N3768, N3767, N521, N1734, N2344);
nand NAND4 (N3769, N3731, N1772, N92, N2457);
nand NAND2 (N3770, N3768, N3703);
and AND2 (N3771, N3765, N3437);
nor NOR4 (N3772, N3759, N3635, N2068, N2851);
and AND3 (N3773, N3763, N2691, N3256);
nand NAND4 (N3774, N3760, N1106, N1708, N3498);
nand NAND2 (N3775, N3769, N2404);
not NOT1 (N3776, N3773);
nor NOR2 (N3777, N3772, N2405);
nand NAND2 (N3778, N3771, N1323);
or OR4 (N3779, N3777, N2241, N3756, N1751);
or OR3 (N3780, N3779, N1252, N1690);
or OR4 (N3781, N3780, N752, N1714, N638);
or OR3 (N3782, N3778, N3349, N400);
and AND2 (N3783, N3747, N672);
nand NAND2 (N3784, N3781, N3409);
not NOT1 (N3785, N3776);
nand NAND2 (N3786, N3757, N3480);
buf BUF1 (N3787, N3774);
and AND4 (N3788, N3770, N108, N2116, N973);
xor XOR2 (N3789, N3775, N2288);
or OR4 (N3790, N3785, N300, N472, N1599);
and AND3 (N3791, N3786, N2463, N2486);
and AND4 (N3792, N3766, N2626, N3589, N730);
nand NAND4 (N3793, N3783, N948, N1241, N1232);
not NOT1 (N3794, N3791);
or OR4 (N3795, N3787, N3422, N1384, N3549);
not NOT1 (N3796, N3782);
buf BUF1 (N3797, N3790);
nand NAND4 (N3798, N3789, N1245, N2715, N2545);
and AND3 (N3799, N3793, N3616, N3411);
xor XOR2 (N3800, N3796, N1820);
or OR3 (N3801, N3795, N2343, N1009);
and AND4 (N3802, N3762, N3047, N1811, N2244);
nand NAND4 (N3803, N3784, N1859, N1645, N1305);
and AND3 (N3804, N3794, N1508, N547);
not NOT1 (N3805, N3788);
nor NOR4 (N3806, N3792, N3149, N2484, N10);
or OR2 (N3807, N3805, N2237);
nor NOR4 (N3808, N3800, N3497, N46, N538);
not NOT1 (N3809, N3801);
not NOT1 (N3810, N3802);
or OR2 (N3811, N3808, N3057);
nor NOR2 (N3812, N3803, N3523);
buf BUF1 (N3813, N3804);
nand NAND2 (N3814, N3810, N3756);
buf BUF1 (N3815, N3809);
nor NOR3 (N3816, N3797, N1996, N1927);
or OR3 (N3817, N3813, N2118, N1823);
or OR2 (N3818, N3798, N979);
nand NAND4 (N3819, N3816, N2038, N1863, N359);
xor XOR2 (N3820, N3815, N813);
nand NAND3 (N3821, N3817, N875, N2356);
nand NAND4 (N3822, N3811, N71, N380, N378);
not NOT1 (N3823, N3806);
nand NAND4 (N3824, N3820, N2988, N2969, N2949);
and AND3 (N3825, N3812, N553, N2499);
xor XOR2 (N3826, N3821, N2502);
xor XOR2 (N3827, N3818, N1609);
or OR3 (N3828, N3827, N648, N2641);
or OR4 (N3829, N3799, N3475, N3594, N2102);
xor XOR2 (N3830, N3824, N3705);
or OR4 (N3831, N3822, N746, N3643, N2016);
xor XOR2 (N3832, N3814, N522);
buf BUF1 (N3833, N3823);
nand NAND2 (N3834, N3831, N244);
nand NAND3 (N3835, N3832, N3211, N2934);
or OR4 (N3836, N3830, N3091, N2856, N875);
and AND3 (N3837, N3807, N2632, N2102);
or OR4 (N3838, N3829, N1426, N1472, N3362);
or OR3 (N3839, N3828, N1246, N2513);
buf BUF1 (N3840, N3833);
or OR4 (N3841, N3826, N1834, N344, N1802);
xor XOR2 (N3842, N3839, N3053);
not NOT1 (N3843, N3841);
not NOT1 (N3844, N3837);
and AND4 (N3845, N3835, N1112, N65, N1784);
not NOT1 (N3846, N3834);
buf BUF1 (N3847, N3825);
nor NOR3 (N3848, N3844, N1483, N2286);
xor XOR2 (N3849, N3846, N1958);
buf BUF1 (N3850, N3843);
xor XOR2 (N3851, N3849, N3663);
nor NOR4 (N3852, N3819, N1883, N679, N1285);
buf BUF1 (N3853, N3842);
xor XOR2 (N3854, N3852, N3807);
and AND4 (N3855, N3850, N589, N1791, N3618);
nor NOR4 (N3856, N3840, N3689, N3036, N460);
not NOT1 (N3857, N3853);
buf BUF1 (N3858, N3845);
nand NAND2 (N3859, N3858, N783);
xor XOR2 (N3860, N3848, N436);
buf BUF1 (N3861, N3860);
or OR2 (N3862, N3855, N613);
or OR2 (N3863, N3836, N1354);
or OR3 (N3864, N3851, N1076, N1385);
nor NOR4 (N3865, N3856, N2182, N2166, N973);
xor XOR2 (N3866, N3854, N1968);
xor XOR2 (N3867, N3865, N17);
xor XOR2 (N3868, N3863, N2121);
not NOT1 (N3869, N3864);
nand NAND3 (N3870, N3838, N1330, N2726);
buf BUF1 (N3871, N3847);
or OR3 (N3872, N3866, N2827, N1707);
not NOT1 (N3873, N3861);
nor NOR4 (N3874, N3870, N1128, N2651, N3031);
nor NOR3 (N3875, N3869, N2448, N620);
nand NAND4 (N3876, N3867, N3509, N2550, N2277);
xor XOR2 (N3877, N3868, N3507);
nand NAND3 (N3878, N3871, N2578, N1884);
or OR2 (N3879, N3877, N1526);
or OR4 (N3880, N3874, N1885, N3011, N2697);
xor XOR2 (N3881, N3862, N3692);
xor XOR2 (N3882, N3880, N3514);
xor XOR2 (N3883, N3859, N2192);
buf BUF1 (N3884, N3881);
and AND2 (N3885, N3875, N2466);
not NOT1 (N3886, N3879);
or OR2 (N3887, N3885, N1171);
nor NOR2 (N3888, N3883, N257);
buf BUF1 (N3889, N3876);
not NOT1 (N3890, N3889);
buf BUF1 (N3891, N3873);
and AND4 (N3892, N3890, N714, N900, N739);
nand NAND3 (N3893, N3878, N3284, N2661);
not NOT1 (N3894, N3886);
nand NAND4 (N3895, N3887, N208, N2490, N3851);
xor XOR2 (N3896, N3857, N2511);
nand NAND2 (N3897, N3895, N2500);
nand NAND3 (N3898, N3896, N2089, N2339);
xor XOR2 (N3899, N3891, N3179);
xor XOR2 (N3900, N3882, N2770);
and AND2 (N3901, N3899, N1259);
not NOT1 (N3902, N3884);
not NOT1 (N3903, N3902);
buf BUF1 (N3904, N3892);
or OR4 (N3905, N3894, N253, N21, N2564);
and AND2 (N3906, N3905, N2846);
nand NAND2 (N3907, N3898, N3130);
and AND3 (N3908, N3893, N3533, N2189);
xor XOR2 (N3909, N3897, N663);
buf BUF1 (N3910, N3908);
buf BUF1 (N3911, N3903);
nor NOR4 (N3912, N3906, N2603, N1913, N2823);
and AND2 (N3913, N3907, N3657);
not NOT1 (N3914, N3910);
xor XOR2 (N3915, N3901, N1847);
nor NOR3 (N3916, N3909, N1250, N2596);
not NOT1 (N3917, N3911);
buf BUF1 (N3918, N3913);
xor XOR2 (N3919, N3912, N2742);
buf BUF1 (N3920, N3919);
buf BUF1 (N3921, N3916);
nand NAND3 (N3922, N3900, N1069, N1674);
nor NOR3 (N3923, N3920, N2229, N2296);
nor NOR3 (N3924, N3921, N2201, N2689);
not NOT1 (N3925, N3872);
not NOT1 (N3926, N3914);
buf BUF1 (N3927, N3904);
or OR3 (N3928, N3925, N2224, N2143);
buf BUF1 (N3929, N3927);
not NOT1 (N3930, N3922);
not NOT1 (N3931, N3888);
not NOT1 (N3932, N3929);
nand NAND2 (N3933, N3918, N1881);
not NOT1 (N3934, N3932);
not NOT1 (N3935, N3926);
not NOT1 (N3936, N3928);
nand NAND4 (N3937, N3917, N2887, N613, N451);
buf BUF1 (N3938, N3924);
nand NAND2 (N3939, N3923, N2829);
nand NAND4 (N3940, N3939, N2031, N3720, N741);
xor XOR2 (N3941, N3930, N1893);
or OR3 (N3942, N3935, N3745, N517);
nand NAND3 (N3943, N3934, N1015, N493);
buf BUF1 (N3944, N3915);
or OR4 (N3945, N3943, N3852, N2271, N2544);
nand NAND3 (N3946, N3933, N529, N520);
not NOT1 (N3947, N3940);
xor XOR2 (N3948, N3945, N1959);
not NOT1 (N3949, N3938);
nor NOR4 (N3950, N3936, N1220, N2488, N864);
and AND2 (N3951, N3947, N3716);
nor NOR4 (N3952, N3931, N953, N1575, N1490);
nand NAND2 (N3953, N3950, N3667);
xor XOR2 (N3954, N3951, N1277);
nor NOR4 (N3955, N3953, N1284, N794, N192);
not NOT1 (N3956, N3948);
not NOT1 (N3957, N3946);
xor XOR2 (N3958, N3937, N1356);
nor NOR2 (N3959, N3942, N3080);
and AND3 (N3960, N3955, N1113, N3730);
xor XOR2 (N3961, N3960, N999);
not NOT1 (N3962, N3957);
and AND3 (N3963, N3952, N716, N3219);
nand NAND3 (N3964, N3958, N1011, N3563);
nand NAND4 (N3965, N3961, N2997, N1434, N3540);
nor NOR3 (N3966, N3963, N3162, N3152);
or OR2 (N3967, N3964, N1211);
and AND3 (N3968, N3962, N690, N3530);
xor XOR2 (N3969, N3949, N1910);
nor NOR2 (N3970, N3968, N122);
and AND4 (N3971, N3954, N3586, N2937, N659);
buf BUF1 (N3972, N3965);
nand NAND2 (N3973, N3956, N3187);
nor NOR3 (N3974, N3967, N3491, N13);
nand NAND2 (N3975, N3944, N1078);
buf BUF1 (N3976, N3941);
not NOT1 (N3977, N3959);
buf BUF1 (N3978, N3966);
not NOT1 (N3979, N3976);
not NOT1 (N3980, N3974);
nand NAND2 (N3981, N3971, N816);
nand NAND3 (N3982, N3969, N3581, N2684);
or OR2 (N3983, N3972, N616);
not NOT1 (N3984, N3978);
xor XOR2 (N3985, N3984, N3151);
and AND3 (N3986, N3970, N1214, N375);
or OR4 (N3987, N3982, N1793, N2464, N2452);
buf BUF1 (N3988, N3977);
nand NAND2 (N3989, N3981, N2552);
and AND3 (N3990, N3985, N3355, N1);
buf BUF1 (N3991, N3989);
or OR3 (N3992, N3988, N2940, N1415);
buf BUF1 (N3993, N3983);
not NOT1 (N3994, N3975);
nor NOR3 (N3995, N3992, N829, N1049);
nand NAND4 (N3996, N3991, N2772, N1317, N2968);
or OR4 (N3997, N3987, N183, N2777, N1240);
xor XOR2 (N3998, N3980, N468);
not NOT1 (N3999, N3997);
and AND2 (N4000, N3994, N2238);
buf BUF1 (N4001, N3993);
or OR3 (N4002, N3998, N3607, N3344);
buf BUF1 (N4003, N3996);
and AND2 (N4004, N3979, N2526);
nand NAND3 (N4005, N3973, N613, N2189);
xor XOR2 (N4006, N4001, N459);
buf BUF1 (N4007, N4006);
not NOT1 (N4008, N3999);
or OR2 (N4009, N4000, N848);
nand NAND4 (N4010, N4002, N3900, N252, N3902);
endmodule