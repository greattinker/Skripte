// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19;

output N12808,N12801,N12810,N12815,N12816,N12817,N12803,N12812,N12814,N12819;

or OR3 (N20, N10, N10, N15);
buf BUF1 (N21, N2);
xor XOR2 (N22, N10, N7);
buf BUF1 (N23, N20);
nor NOR2 (N24, N16, N15);
nand NAND4 (N25, N4, N15, N5, N3);
xor XOR2 (N26, N20, N5);
and AND2 (N27, N9, N18);
xor XOR2 (N28, N17, N7);
nor NOR3 (N29, N24, N28, N16);
nand NAND3 (N30, N15, N5, N22);
not NOT1 (N31, N30);
or OR3 (N32, N26, N2, N22);
nor NOR2 (N33, N24, N1);
not NOT1 (N34, N12);
nand NAND4 (N35, N23, N24, N25, N22);
not NOT1 (N36, N33);
xor XOR2 (N37, N17, N11);
not NOT1 (N38, N18);
xor XOR2 (N39, N35, N24);
xor XOR2 (N40, N34, N15);
or OR3 (N41, N40, N34, N15);
or OR2 (N42, N37, N35);
nand NAND2 (N43, N31, N31);
xor XOR2 (N44, N43, N30);
xor XOR2 (N45, N32, N42);
buf BUF1 (N46, N5);
and AND4 (N47, N46, N28, N16, N20);
not NOT1 (N48, N29);
xor XOR2 (N49, N47, N13);
nand NAND4 (N50, N49, N26, N5, N7);
xor XOR2 (N51, N45, N31);
nand NAND2 (N52, N48, N29);
or OR2 (N53, N39, N38);
xor XOR2 (N54, N41, N7);
or OR4 (N55, N46, N47, N49, N16);
xor XOR2 (N56, N27, N51);
or OR3 (N57, N45, N17, N39);
buf BUF1 (N58, N56);
or OR2 (N59, N36, N21);
not NOT1 (N60, N13);
nor NOR4 (N61, N50, N19, N33, N26);
not NOT1 (N62, N54);
and AND4 (N63, N52, N26, N29, N38);
or OR4 (N64, N62, N40, N51, N12);
xor XOR2 (N65, N58, N17);
or OR4 (N66, N44, N65, N28, N6);
nand NAND4 (N67, N41, N42, N7, N35);
nor NOR3 (N68, N55, N10, N13);
and AND4 (N69, N63, N54, N8, N2);
and AND4 (N70, N66, N57, N40, N25);
xor XOR2 (N71, N37, N18);
nand NAND3 (N72, N64, N66, N5);
nand NAND2 (N73, N72, N41);
xor XOR2 (N74, N73, N4);
and AND4 (N75, N69, N1, N34, N13);
xor XOR2 (N76, N67, N20);
or OR2 (N77, N60, N41);
buf BUF1 (N78, N74);
not NOT1 (N79, N53);
or OR2 (N80, N79, N41);
buf BUF1 (N81, N75);
buf BUF1 (N82, N68);
not NOT1 (N83, N61);
or OR4 (N84, N71, N29, N16, N32);
not NOT1 (N85, N76);
and AND4 (N86, N80, N57, N12, N42);
nor NOR4 (N87, N85, N25, N37, N18);
or OR3 (N88, N70, N54, N25);
nor NOR3 (N89, N84, N62, N71);
nor NOR3 (N90, N78, N62, N12);
and AND4 (N91, N82, N46, N49, N5);
nand NAND2 (N92, N89, N46);
nor NOR2 (N93, N88, N38);
nor NOR2 (N94, N86, N36);
not NOT1 (N95, N59);
xor XOR2 (N96, N94, N45);
nand NAND2 (N97, N77, N78);
or OR2 (N98, N87, N55);
or OR3 (N99, N97, N31, N21);
xor XOR2 (N100, N93, N47);
buf BUF1 (N101, N83);
and AND3 (N102, N90, N60, N32);
and AND3 (N103, N92, N77, N9);
xor XOR2 (N104, N81, N17);
not NOT1 (N105, N104);
and AND2 (N106, N91, N47);
nand NAND4 (N107, N106, N35, N4, N32);
and AND2 (N108, N107, N7);
nor NOR4 (N109, N98, N86, N77, N19);
nand NAND3 (N110, N109, N87, N12);
and AND4 (N111, N102, N93, N90, N99);
and AND4 (N112, N20, N67, N92, N32);
buf BUF1 (N113, N100);
nand NAND3 (N114, N95, N82, N13);
nand NAND4 (N115, N108, N64, N77, N61);
nand NAND4 (N116, N105, N73, N33, N44);
nand NAND4 (N117, N101, N61, N15, N41);
buf BUF1 (N118, N96);
nand NAND3 (N119, N114, N27, N1);
buf BUF1 (N120, N103);
nor NOR2 (N121, N119, N27);
not NOT1 (N122, N115);
not NOT1 (N123, N121);
or OR2 (N124, N113, N96);
and AND3 (N125, N120, N6, N15);
nor NOR4 (N126, N110, N112, N86, N17);
and AND2 (N127, N49, N104);
nor NOR2 (N128, N111, N63);
nor NOR2 (N129, N123, N123);
buf BUF1 (N130, N117);
nand NAND2 (N131, N118, N38);
buf BUF1 (N132, N126);
nand NAND3 (N133, N127, N69, N112);
and AND4 (N134, N129, N7, N115, N133);
and AND3 (N135, N111, N63, N129);
not NOT1 (N136, N128);
nand NAND4 (N137, N130, N127, N45, N11);
and AND3 (N138, N124, N1, N67);
xor XOR2 (N139, N125, N38);
buf BUF1 (N140, N116);
nand NAND3 (N141, N136, N132, N115);
or OR4 (N142, N49, N99, N100, N81);
not NOT1 (N143, N122);
and AND4 (N144, N131, N94, N60, N47);
not NOT1 (N145, N134);
and AND3 (N146, N141, N45, N9);
not NOT1 (N147, N143);
nand NAND2 (N148, N142, N63);
buf BUF1 (N149, N137);
buf BUF1 (N150, N145);
or OR4 (N151, N146, N142, N105, N44);
not NOT1 (N152, N150);
xor XOR2 (N153, N147, N122);
xor XOR2 (N154, N140, N15);
nor NOR4 (N155, N139, N83, N140, N15);
xor XOR2 (N156, N135, N99);
nand NAND2 (N157, N138, N30);
buf BUF1 (N158, N149);
or OR2 (N159, N152, N117);
nor NOR3 (N160, N151, N35, N155);
and AND4 (N161, N5, N143, N32, N60);
nor NOR3 (N162, N153, N11, N160);
buf BUF1 (N163, N58);
or OR2 (N164, N163, N155);
nand NAND3 (N165, N156, N82, N35);
or OR2 (N166, N162, N37);
and AND2 (N167, N166, N38);
not NOT1 (N168, N158);
nand NAND2 (N169, N154, N50);
nor NOR4 (N170, N144, N105, N94, N160);
nor NOR4 (N171, N148, N53, N37, N116);
not NOT1 (N172, N157);
nand NAND2 (N173, N159, N109);
and AND4 (N174, N170, N97, N121, N169);
or OR3 (N175, N152, N62, N153);
or OR2 (N176, N161, N133);
xor XOR2 (N177, N165, N59);
or OR3 (N178, N175, N64, N81);
buf BUF1 (N179, N178);
xor XOR2 (N180, N172, N71);
not NOT1 (N181, N179);
nand NAND2 (N182, N177, N40);
or OR2 (N183, N182, N7);
and AND3 (N184, N168, N72, N131);
and AND4 (N185, N184, N64, N98, N2);
nand NAND3 (N186, N176, N137, N177);
not NOT1 (N187, N186);
or OR4 (N188, N173, N55, N20, N78);
and AND3 (N189, N164, N111, N25);
nor NOR3 (N190, N180, N149, N59);
buf BUF1 (N191, N190);
buf BUF1 (N192, N187);
or OR3 (N193, N174, N168, N153);
or OR2 (N194, N192, N33);
nand NAND2 (N195, N191, N121);
or OR4 (N196, N189, N102, N59, N167);
and AND4 (N197, N182, N102, N128, N87);
not NOT1 (N198, N188);
or OR4 (N199, N197, N174, N92, N164);
nand NAND3 (N200, N196, N175, N57);
xor XOR2 (N201, N198, N152);
xor XOR2 (N202, N194, N169);
and AND4 (N203, N201, N101, N72, N111);
nor NOR4 (N204, N185, N106, N39, N88);
or OR2 (N205, N193, N113);
and AND3 (N206, N199, N108, N125);
and AND3 (N207, N203, N57, N182);
or OR2 (N208, N181, N176);
nor NOR3 (N209, N207, N119, N59);
buf BUF1 (N210, N205);
buf BUF1 (N211, N206);
or OR2 (N212, N202, N111);
xor XOR2 (N213, N204, N94);
nand NAND2 (N214, N211, N24);
and AND4 (N215, N214, N93, N126, N158);
xor XOR2 (N216, N210, N102);
buf BUF1 (N217, N195);
xor XOR2 (N218, N171, N130);
nor NOR4 (N219, N213, N93, N197, N200);
buf BUF1 (N220, N95);
or OR2 (N221, N217, N147);
not NOT1 (N222, N220);
buf BUF1 (N223, N208);
xor XOR2 (N224, N209, N166);
nand NAND2 (N225, N222, N34);
xor XOR2 (N226, N225, N86);
nor NOR4 (N227, N216, N197, N182, N131);
and AND4 (N228, N226, N203, N128, N185);
buf BUF1 (N229, N183);
buf BUF1 (N230, N219);
xor XOR2 (N231, N229, N6);
and AND3 (N232, N218, N40, N223);
buf BUF1 (N233, N191);
buf BUF1 (N234, N231);
buf BUF1 (N235, N234);
buf BUF1 (N236, N235);
buf BUF1 (N237, N232);
xor XOR2 (N238, N212, N57);
or OR4 (N239, N233, N14, N31, N100);
buf BUF1 (N240, N236);
xor XOR2 (N241, N227, N1);
or OR3 (N242, N221, N107, N127);
nor NOR4 (N243, N215, N26, N174, N132);
xor XOR2 (N244, N237, N237);
and AND3 (N245, N228, N139, N163);
and AND4 (N246, N242, N226, N168, N131);
xor XOR2 (N247, N224, N12);
or OR2 (N248, N238, N157);
or OR4 (N249, N248, N95, N198, N38);
nor NOR3 (N250, N239, N211, N137);
nand NAND4 (N251, N241, N182, N173, N185);
nor NOR4 (N252, N230, N182, N74, N50);
or OR2 (N253, N251, N235);
and AND4 (N254, N252, N190, N196, N25);
not NOT1 (N255, N247);
nor NOR4 (N256, N244, N16, N198, N6);
and AND4 (N257, N254, N180, N168, N200);
xor XOR2 (N258, N245, N185);
nand NAND3 (N259, N256, N257, N115);
buf BUF1 (N260, N82);
xor XOR2 (N261, N243, N11);
not NOT1 (N262, N253);
not NOT1 (N263, N249);
not NOT1 (N264, N258);
not NOT1 (N265, N259);
xor XOR2 (N266, N262, N251);
xor XOR2 (N267, N250, N136);
and AND4 (N268, N265, N213, N35, N262);
not NOT1 (N269, N268);
nor NOR3 (N270, N266, N214, N54);
nor NOR2 (N271, N264, N71);
or OR2 (N272, N255, N249);
or OR4 (N273, N263, N252, N161, N147);
and AND2 (N274, N271, N184);
nand NAND2 (N275, N272, N24);
and AND2 (N276, N261, N108);
buf BUF1 (N277, N260);
xor XOR2 (N278, N270, N172);
nand NAND3 (N279, N275, N38, N136);
buf BUF1 (N280, N240);
nand NAND3 (N281, N274, N223, N112);
buf BUF1 (N282, N269);
nand NAND3 (N283, N273, N39, N236);
and AND2 (N284, N276, N257);
buf BUF1 (N285, N246);
nand NAND2 (N286, N282, N135);
not NOT1 (N287, N283);
xor XOR2 (N288, N287, N103);
buf BUF1 (N289, N279);
or OR3 (N290, N289, N55, N199);
not NOT1 (N291, N277);
buf BUF1 (N292, N286);
nor NOR4 (N293, N284, N141, N44, N132);
not NOT1 (N294, N285);
and AND3 (N295, N267, N202, N53);
nor NOR3 (N296, N293, N226, N107);
buf BUF1 (N297, N281);
or OR2 (N298, N288, N203);
and AND3 (N299, N290, N207, N7);
nor NOR3 (N300, N296, N286, N208);
nor NOR3 (N301, N280, N39, N102);
xor XOR2 (N302, N295, N7);
nor NOR3 (N303, N297, N245, N35);
or OR3 (N304, N278, N87, N80);
nor NOR4 (N305, N298, N298, N275, N225);
or OR4 (N306, N301, N271, N148, N146);
not NOT1 (N307, N291);
and AND4 (N308, N299, N251, N304, N86);
nand NAND4 (N309, N143, N254, N167, N219);
and AND2 (N310, N300, N200);
buf BUF1 (N311, N306);
and AND4 (N312, N302, N101, N265, N109);
buf BUF1 (N313, N311);
nor NOR4 (N314, N313, N28, N267, N201);
and AND2 (N315, N309, N20);
not NOT1 (N316, N307);
nand NAND3 (N317, N314, N221, N50);
nand NAND2 (N318, N312, N144);
xor XOR2 (N319, N305, N237);
nand NAND3 (N320, N317, N225, N118);
and AND4 (N321, N315, N72, N165, N159);
buf BUF1 (N322, N292);
nand NAND4 (N323, N308, N77, N167, N129);
nor NOR3 (N324, N321, N252, N78);
and AND4 (N325, N316, N222, N302, N20);
buf BUF1 (N326, N322);
nor NOR2 (N327, N323, N100);
not NOT1 (N328, N326);
buf BUF1 (N329, N319);
nand NAND3 (N330, N325, N81, N267);
nor NOR3 (N331, N303, N117, N67);
not NOT1 (N332, N330);
nand NAND4 (N333, N324, N24, N71, N24);
nor NOR3 (N334, N327, N223, N23);
not NOT1 (N335, N294);
nand NAND4 (N336, N333, N125, N79, N35);
and AND3 (N337, N328, N255, N11);
and AND4 (N338, N334, N103, N117, N330);
not NOT1 (N339, N329);
not NOT1 (N340, N332);
not NOT1 (N341, N320);
not NOT1 (N342, N339);
and AND2 (N343, N310, N56);
and AND4 (N344, N340, N282, N282, N216);
nand NAND4 (N345, N336, N287, N249, N44);
nand NAND3 (N346, N342, N267, N229);
nor NOR4 (N347, N346, N304, N271, N252);
or OR3 (N348, N345, N277, N45);
and AND3 (N349, N343, N90, N82);
xor XOR2 (N350, N349, N269);
xor XOR2 (N351, N341, N140);
nor NOR2 (N352, N351, N238);
not NOT1 (N353, N331);
xor XOR2 (N354, N347, N191);
nor NOR2 (N355, N350, N201);
not NOT1 (N356, N344);
nor NOR3 (N357, N354, N328, N244);
and AND2 (N358, N356, N181);
nor NOR3 (N359, N348, N56, N331);
or OR4 (N360, N318, N65, N256, N313);
xor XOR2 (N361, N357, N180);
buf BUF1 (N362, N353);
and AND4 (N363, N360, N331, N177, N27);
not NOT1 (N364, N335);
buf BUF1 (N365, N363);
and AND2 (N366, N337, N150);
nand NAND4 (N367, N355, N68, N72, N354);
xor XOR2 (N368, N365, N28);
buf BUF1 (N369, N358);
nor NOR3 (N370, N361, N325, N366);
nor NOR3 (N371, N153, N271, N342);
or OR2 (N372, N359, N70);
nor NOR2 (N373, N338, N99);
nor NOR2 (N374, N373, N260);
and AND2 (N375, N352, N67);
nor NOR2 (N376, N370, N12);
not NOT1 (N377, N376);
nand NAND2 (N378, N367, N339);
buf BUF1 (N379, N375);
not NOT1 (N380, N368);
xor XOR2 (N381, N371, N172);
or OR2 (N382, N364, N304);
xor XOR2 (N383, N377, N178);
not NOT1 (N384, N381);
and AND3 (N385, N384, N137, N304);
xor XOR2 (N386, N369, N131);
buf BUF1 (N387, N362);
nand NAND2 (N388, N383, N321);
not NOT1 (N389, N387);
buf BUF1 (N390, N382);
xor XOR2 (N391, N390, N93);
nand NAND2 (N392, N372, N106);
nand NAND3 (N393, N391, N244, N364);
not NOT1 (N394, N378);
or OR3 (N395, N386, N148, N186);
or OR3 (N396, N394, N186, N79);
not NOT1 (N397, N385);
nand NAND4 (N398, N392, N70, N241, N173);
or OR3 (N399, N393, N85, N22);
not NOT1 (N400, N379);
or OR2 (N401, N395, N176);
not NOT1 (N402, N401);
xor XOR2 (N403, N397, N210);
buf BUF1 (N404, N398);
and AND4 (N405, N380, N371, N103, N281);
not NOT1 (N406, N399);
nand NAND4 (N407, N389, N23, N355, N398);
nor NOR4 (N408, N396, N269, N152, N275);
buf BUF1 (N409, N374);
nor NOR4 (N410, N407, N408, N102, N90);
nor NOR2 (N411, N377, N110);
xor XOR2 (N412, N388, N178);
nand NAND4 (N413, N406, N273, N6, N379);
not NOT1 (N414, N404);
buf BUF1 (N415, N410);
not NOT1 (N416, N413);
and AND2 (N417, N411, N193);
nand NAND2 (N418, N417, N118);
buf BUF1 (N419, N400);
or OR4 (N420, N415, N230, N43, N302);
xor XOR2 (N421, N412, N85);
nand NAND2 (N422, N403, N108);
not NOT1 (N423, N420);
buf BUF1 (N424, N421);
nor NOR3 (N425, N419, N249, N15);
buf BUF1 (N426, N418);
or OR2 (N427, N422, N72);
and AND4 (N428, N427, N32, N410, N72);
xor XOR2 (N429, N428, N396);
not NOT1 (N430, N402);
or OR3 (N431, N409, N157, N376);
nor NOR4 (N432, N429, N94, N418, N150);
nor NOR4 (N433, N424, N387, N85, N351);
and AND3 (N434, N426, N363, N423);
nand NAND2 (N435, N386, N141);
nor NOR2 (N436, N425, N302);
buf BUF1 (N437, N434);
not NOT1 (N438, N430);
and AND2 (N439, N405, N161);
buf BUF1 (N440, N435);
not NOT1 (N441, N414);
buf BUF1 (N442, N440);
buf BUF1 (N443, N442);
xor XOR2 (N444, N441, N284);
not NOT1 (N445, N432);
xor XOR2 (N446, N443, N158);
not NOT1 (N447, N416);
nor NOR3 (N448, N437, N377, N323);
nand NAND3 (N449, N439, N429, N422);
not NOT1 (N450, N444);
nor NOR2 (N451, N446, N118);
xor XOR2 (N452, N451, N109);
and AND2 (N453, N452, N232);
nand NAND2 (N454, N448, N409);
buf BUF1 (N455, N454);
or OR3 (N456, N447, N3, N240);
nor NOR2 (N457, N456, N30);
or OR3 (N458, N438, N322, N145);
xor XOR2 (N459, N450, N272);
nor NOR3 (N460, N445, N436, N5);
and AND2 (N461, N122, N237);
buf BUF1 (N462, N431);
xor XOR2 (N463, N453, N82);
nand NAND3 (N464, N449, N295, N92);
and AND2 (N465, N459, N15);
buf BUF1 (N466, N464);
buf BUF1 (N467, N457);
xor XOR2 (N468, N466, N128);
or OR3 (N469, N467, N89, N395);
not NOT1 (N470, N433);
nand NAND2 (N471, N469, N7);
not NOT1 (N472, N465);
and AND2 (N473, N455, N4);
nor NOR4 (N474, N461, N469, N16, N319);
buf BUF1 (N475, N470);
xor XOR2 (N476, N460, N264);
and AND4 (N477, N471, N182, N230, N144);
nand NAND4 (N478, N468, N109, N181, N194);
and AND3 (N479, N477, N145, N53);
nand NAND3 (N480, N473, N105, N39);
and AND4 (N481, N472, N67, N304, N124);
buf BUF1 (N482, N476);
or OR4 (N483, N474, N280, N252, N41);
buf BUF1 (N484, N480);
buf BUF1 (N485, N479);
buf BUF1 (N486, N485);
nor NOR2 (N487, N462, N427);
not NOT1 (N488, N482);
and AND3 (N489, N463, N249, N327);
and AND2 (N490, N484, N274);
nor NOR4 (N491, N478, N486, N373, N51);
buf BUF1 (N492, N328);
and AND3 (N493, N458, N19, N278);
not NOT1 (N494, N487);
nand NAND3 (N495, N493, N101, N122);
buf BUF1 (N496, N494);
or OR4 (N497, N496, N357, N217, N163);
nor NOR4 (N498, N488, N14, N113, N420);
or OR2 (N499, N475, N183);
or OR3 (N500, N495, N230, N80);
xor XOR2 (N501, N500, N483);
or OR4 (N502, N260, N338, N60, N182);
not NOT1 (N503, N491);
not NOT1 (N504, N481);
xor XOR2 (N505, N490, N99);
nand NAND2 (N506, N492, N271);
or OR4 (N507, N506, N404, N61, N394);
buf BUF1 (N508, N502);
not NOT1 (N509, N497);
buf BUF1 (N510, N504);
nand NAND3 (N511, N501, N450, N269);
buf BUF1 (N512, N507);
and AND3 (N513, N512, N46, N440);
and AND4 (N514, N505, N489, N278, N117);
and AND3 (N515, N89, N110, N67);
not NOT1 (N516, N509);
or OR4 (N517, N516, N131, N142, N302);
buf BUF1 (N518, N513);
nand NAND4 (N519, N515, N13, N177, N104);
and AND3 (N520, N519, N30, N500);
not NOT1 (N521, N508);
buf BUF1 (N522, N511);
nor NOR2 (N523, N510, N66);
or OR4 (N524, N521, N497, N234, N465);
or OR3 (N525, N520, N472, N501);
nand NAND3 (N526, N523, N470, N123);
buf BUF1 (N527, N517);
xor XOR2 (N528, N503, N115);
nor NOR2 (N529, N527, N135);
xor XOR2 (N530, N514, N190);
not NOT1 (N531, N529);
and AND3 (N532, N498, N29, N6);
or OR3 (N533, N532, N312, N90);
or OR2 (N534, N525, N208);
nand NAND3 (N535, N533, N189, N151);
or OR2 (N536, N531, N183);
nand NAND4 (N537, N518, N180, N519, N418);
nor NOR4 (N538, N528, N442, N100, N312);
buf BUF1 (N539, N537);
or OR2 (N540, N524, N135);
or OR3 (N541, N499, N219, N413);
buf BUF1 (N542, N526);
not NOT1 (N543, N540);
not NOT1 (N544, N542);
not NOT1 (N545, N538);
and AND3 (N546, N541, N142, N47);
buf BUF1 (N547, N522);
xor XOR2 (N548, N539, N248);
nor NOR2 (N549, N545, N344);
buf BUF1 (N550, N546);
not NOT1 (N551, N549);
nor NOR2 (N552, N536, N226);
buf BUF1 (N553, N551);
or OR3 (N554, N544, N88, N434);
or OR3 (N555, N548, N525, N398);
or OR4 (N556, N535, N466, N72, N52);
xor XOR2 (N557, N552, N252);
xor XOR2 (N558, N557, N343);
buf BUF1 (N559, N534);
buf BUF1 (N560, N556);
or OR2 (N561, N554, N142);
not NOT1 (N562, N561);
or OR3 (N563, N547, N97, N425);
not NOT1 (N564, N530);
not NOT1 (N565, N563);
not NOT1 (N566, N564);
xor XOR2 (N567, N562, N386);
not NOT1 (N568, N559);
buf BUF1 (N569, N565);
or OR4 (N570, N567, N237, N376, N264);
xor XOR2 (N571, N560, N381);
nor NOR4 (N572, N571, N356, N325, N500);
buf BUF1 (N573, N566);
and AND2 (N574, N558, N516);
and AND4 (N575, N553, N96, N224, N561);
nor NOR2 (N576, N574, N513);
or OR2 (N577, N576, N184);
not NOT1 (N578, N575);
and AND4 (N579, N578, N461, N51, N490);
or OR4 (N580, N573, N487, N552, N82);
nand NAND2 (N581, N570, N270);
buf BUF1 (N582, N550);
and AND4 (N583, N577, N341, N184, N23);
xor XOR2 (N584, N583, N2);
and AND2 (N585, N581, N68);
nand NAND4 (N586, N569, N59, N312, N201);
not NOT1 (N587, N584);
nand NAND4 (N588, N580, N251, N358, N167);
not NOT1 (N589, N555);
nor NOR4 (N590, N543, N96, N301, N378);
not NOT1 (N591, N589);
nand NAND2 (N592, N572, N400);
nor NOR3 (N593, N585, N565, N203);
buf BUF1 (N594, N568);
nand NAND4 (N595, N579, N174, N34, N294);
and AND3 (N596, N586, N439, N274);
not NOT1 (N597, N595);
not NOT1 (N598, N591);
buf BUF1 (N599, N598);
not NOT1 (N600, N588);
not NOT1 (N601, N597);
not NOT1 (N602, N582);
nand NAND2 (N603, N599, N217);
xor XOR2 (N604, N601, N84);
not NOT1 (N605, N593);
nor NOR4 (N606, N592, N561, N573, N163);
or OR2 (N607, N587, N31);
nor NOR2 (N608, N600, N309);
and AND2 (N609, N603, N77);
not NOT1 (N610, N594);
or OR3 (N611, N608, N492, N110);
or OR4 (N612, N609, N310, N186, N568);
xor XOR2 (N613, N612, N261);
buf BUF1 (N614, N596);
not NOT1 (N615, N602);
or OR3 (N616, N607, N332, N253);
and AND2 (N617, N590, N296);
or OR3 (N618, N615, N406, N317);
nor NOR3 (N619, N610, N543, N270);
buf BUF1 (N620, N613);
not NOT1 (N621, N619);
xor XOR2 (N622, N616, N361);
nor NOR4 (N623, N614, N490, N618, N2);
nor NOR3 (N624, N396, N430, N541);
nand NAND3 (N625, N623, N75, N9);
nor NOR2 (N626, N605, N581);
not NOT1 (N627, N606);
and AND3 (N628, N620, N276, N587);
and AND3 (N629, N626, N329, N202);
not NOT1 (N630, N629);
or OR2 (N631, N604, N122);
not NOT1 (N632, N611);
not NOT1 (N633, N617);
buf BUF1 (N634, N627);
nor NOR4 (N635, N631, N302, N173, N528);
not NOT1 (N636, N625);
and AND4 (N637, N635, N157, N307, N356);
not NOT1 (N638, N634);
xor XOR2 (N639, N636, N533);
or OR2 (N640, N633, N366);
xor XOR2 (N641, N621, N111);
or OR3 (N642, N630, N220, N503);
nand NAND4 (N643, N622, N481, N629, N363);
xor XOR2 (N644, N639, N480);
nand NAND3 (N645, N628, N394, N546);
not NOT1 (N646, N645);
nor NOR2 (N647, N624, N155);
nand NAND3 (N648, N638, N61, N100);
and AND4 (N649, N632, N582, N587, N295);
and AND2 (N650, N649, N203);
or OR4 (N651, N646, N558, N119, N438);
buf BUF1 (N652, N643);
nand NAND2 (N653, N640, N66);
xor XOR2 (N654, N648, N179);
nand NAND2 (N655, N652, N576);
xor XOR2 (N656, N647, N356);
not NOT1 (N657, N637);
not NOT1 (N658, N644);
nor NOR3 (N659, N657, N576, N637);
nand NAND3 (N660, N653, N369, N535);
nor NOR4 (N661, N659, N412, N118, N571);
buf BUF1 (N662, N654);
and AND2 (N663, N641, N97);
buf BUF1 (N664, N658);
xor XOR2 (N665, N650, N92);
or OR4 (N666, N651, N266, N228, N533);
not NOT1 (N667, N666);
buf BUF1 (N668, N665);
xor XOR2 (N669, N655, N566);
nand NAND3 (N670, N664, N397, N666);
or OR4 (N671, N663, N258, N383, N558);
not NOT1 (N672, N667);
nand NAND4 (N673, N660, N571, N247, N650);
nand NAND4 (N674, N668, N456, N268, N288);
and AND3 (N675, N672, N320, N395);
buf BUF1 (N676, N656);
and AND2 (N677, N676, N121);
xor XOR2 (N678, N670, N224);
nor NOR2 (N679, N671, N311);
xor XOR2 (N680, N674, N273);
nor NOR3 (N681, N677, N242, N401);
xor XOR2 (N682, N679, N442);
or OR3 (N683, N662, N213, N317);
not NOT1 (N684, N682);
xor XOR2 (N685, N678, N242);
xor XOR2 (N686, N684, N396);
xor XOR2 (N687, N673, N332);
not NOT1 (N688, N686);
or OR2 (N689, N681, N234);
xor XOR2 (N690, N669, N576);
xor XOR2 (N691, N688, N60);
not NOT1 (N692, N687);
not NOT1 (N693, N691);
nand NAND3 (N694, N642, N122, N1);
nand NAND2 (N695, N689, N343);
or OR3 (N696, N694, N301, N202);
nand NAND3 (N697, N692, N404, N501);
nand NAND2 (N698, N695, N33);
xor XOR2 (N699, N661, N132);
xor XOR2 (N700, N693, N620);
nand NAND3 (N701, N690, N313, N620);
not NOT1 (N702, N680);
not NOT1 (N703, N698);
nand NAND4 (N704, N702, N489, N357, N303);
xor XOR2 (N705, N685, N226);
buf BUF1 (N706, N700);
buf BUF1 (N707, N675);
buf BUF1 (N708, N703);
xor XOR2 (N709, N696, N421);
nor NOR2 (N710, N707, N60);
or OR2 (N711, N705, N617);
xor XOR2 (N712, N708, N607);
nor NOR3 (N713, N704, N185, N157);
or OR3 (N714, N710, N327, N271);
buf BUF1 (N715, N697);
and AND3 (N716, N711, N112, N548);
xor XOR2 (N717, N712, N154);
buf BUF1 (N718, N709);
or OR4 (N719, N715, N203, N417, N604);
not NOT1 (N720, N718);
nor NOR4 (N721, N716, N469, N556, N623);
not NOT1 (N722, N701);
or OR3 (N723, N722, N412, N416);
and AND2 (N724, N717, N155);
nor NOR3 (N725, N720, N112, N47);
and AND4 (N726, N723, N104, N49, N141);
and AND2 (N727, N726, N129);
not NOT1 (N728, N714);
or OR2 (N729, N699, N463);
not NOT1 (N730, N728);
nor NOR2 (N731, N729, N469);
nor NOR4 (N732, N731, N466, N222, N240);
xor XOR2 (N733, N713, N709);
not NOT1 (N734, N724);
nor NOR3 (N735, N721, N192, N536);
xor XOR2 (N736, N706, N516);
or OR3 (N737, N732, N487, N710);
or OR2 (N738, N719, N569);
nand NAND3 (N739, N737, N114, N80);
nor NOR4 (N740, N739, N250, N62, N645);
xor XOR2 (N741, N733, N226);
not NOT1 (N742, N727);
nand NAND4 (N743, N740, N293, N492, N23);
nand NAND3 (N744, N738, N523, N681);
or OR4 (N745, N742, N654, N118, N376);
buf BUF1 (N746, N745);
buf BUF1 (N747, N730);
and AND4 (N748, N734, N636, N327, N457);
nand NAND3 (N749, N735, N249, N510);
and AND3 (N750, N746, N464, N199);
nor NOR2 (N751, N744, N530);
nor NOR3 (N752, N743, N674, N699);
nand NAND3 (N753, N736, N187, N199);
not NOT1 (N754, N752);
nor NOR3 (N755, N753, N113, N173);
and AND2 (N756, N754, N310);
not NOT1 (N757, N756);
and AND2 (N758, N683, N571);
not NOT1 (N759, N750);
buf BUF1 (N760, N751);
or OR4 (N761, N725, N427, N427, N248);
not NOT1 (N762, N760);
and AND2 (N763, N747, N178);
or OR3 (N764, N761, N4, N542);
nand NAND3 (N765, N763, N485, N548);
not NOT1 (N766, N749);
or OR2 (N767, N766, N182);
not NOT1 (N768, N758);
nor NOR3 (N769, N757, N176, N128);
not NOT1 (N770, N768);
nand NAND4 (N771, N759, N321, N270, N449);
nor NOR4 (N772, N767, N268, N128, N164);
not NOT1 (N773, N764);
not NOT1 (N774, N755);
buf BUF1 (N775, N772);
not NOT1 (N776, N748);
nand NAND4 (N777, N770, N545, N57, N769);
and AND4 (N778, N324, N183, N593, N251);
or OR3 (N779, N765, N178, N164);
nor NOR2 (N780, N775, N469);
xor XOR2 (N781, N741, N117);
not NOT1 (N782, N777);
not NOT1 (N783, N779);
nand NAND4 (N784, N774, N145, N502, N724);
nand NAND2 (N785, N762, N195);
not NOT1 (N786, N773);
not NOT1 (N787, N782);
or OR3 (N788, N771, N240, N17);
nor NOR3 (N789, N783, N160, N140);
xor XOR2 (N790, N784, N660);
xor XOR2 (N791, N787, N71);
nor NOR3 (N792, N776, N51, N193);
or OR3 (N793, N778, N672, N226);
buf BUF1 (N794, N789);
nand NAND4 (N795, N780, N34, N499, N13);
and AND2 (N796, N795, N199);
xor XOR2 (N797, N790, N554);
not NOT1 (N798, N796);
nand NAND4 (N799, N781, N75, N243, N227);
nor NOR4 (N800, N788, N440, N33, N246);
buf BUF1 (N801, N800);
nand NAND2 (N802, N792, N742);
nor NOR4 (N803, N794, N625, N609, N497);
not NOT1 (N804, N798);
nand NAND2 (N805, N802, N96);
nand NAND2 (N806, N799, N300);
nand NAND2 (N807, N801, N165);
or OR2 (N808, N805, N153);
nand NAND2 (N809, N786, N504);
not NOT1 (N810, N808);
not NOT1 (N811, N810);
nand NAND4 (N812, N803, N475, N694, N143);
not NOT1 (N813, N797);
or OR4 (N814, N811, N733, N685, N312);
nor NOR4 (N815, N793, N610, N411, N69);
nor NOR3 (N816, N806, N734, N23);
not NOT1 (N817, N813);
not NOT1 (N818, N809);
nor NOR3 (N819, N816, N123, N146);
not NOT1 (N820, N817);
xor XOR2 (N821, N814, N67);
buf BUF1 (N822, N791);
and AND4 (N823, N785, N17, N388, N334);
not NOT1 (N824, N822);
buf BUF1 (N825, N819);
nor NOR2 (N826, N804, N48);
nand NAND2 (N827, N815, N332);
not NOT1 (N828, N825);
not NOT1 (N829, N807);
buf BUF1 (N830, N824);
not NOT1 (N831, N818);
xor XOR2 (N832, N812, N294);
and AND2 (N833, N829, N814);
nand NAND2 (N834, N823, N472);
nand NAND4 (N835, N820, N833, N506, N568);
not NOT1 (N836, N402);
nor NOR3 (N837, N830, N811, N168);
nor NOR3 (N838, N837, N573, N778);
or OR2 (N839, N827, N667);
xor XOR2 (N840, N834, N9);
nand NAND4 (N841, N832, N335, N598, N777);
buf BUF1 (N842, N840);
or OR3 (N843, N839, N6, N173);
nand NAND3 (N844, N842, N160, N360);
nor NOR3 (N845, N828, N815, N98);
buf BUF1 (N846, N844);
buf BUF1 (N847, N821);
nor NOR4 (N848, N826, N823, N750, N746);
and AND4 (N849, N841, N579, N546, N179);
or OR2 (N850, N846, N310);
nand NAND2 (N851, N836, N797);
xor XOR2 (N852, N845, N232);
not NOT1 (N853, N847);
xor XOR2 (N854, N843, N228);
not NOT1 (N855, N838);
nand NAND2 (N856, N849, N266);
not NOT1 (N857, N848);
or OR2 (N858, N831, N91);
xor XOR2 (N859, N854, N439);
and AND4 (N860, N856, N600, N687, N686);
not NOT1 (N861, N857);
buf BUF1 (N862, N853);
or OR3 (N863, N835, N314, N40);
buf BUF1 (N864, N855);
buf BUF1 (N865, N860);
and AND4 (N866, N850, N546, N649, N238);
and AND2 (N867, N852, N331);
nor NOR2 (N868, N859, N670);
xor XOR2 (N869, N865, N829);
or OR4 (N870, N861, N531, N545, N533);
nor NOR2 (N871, N868, N831);
buf BUF1 (N872, N858);
xor XOR2 (N873, N867, N34);
nand NAND4 (N874, N866, N520, N363, N77);
and AND3 (N875, N874, N151, N806);
nand NAND4 (N876, N869, N875, N824, N652);
not NOT1 (N877, N196);
or OR4 (N878, N876, N164, N436, N353);
buf BUF1 (N879, N862);
nand NAND2 (N880, N863, N877);
and AND2 (N881, N178, N267);
buf BUF1 (N882, N873);
nor NOR2 (N883, N871, N496);
buf BUF1 (N884, N878);
buf BUF1 (N885, N884);
xor XOR2 (N886, N881, N395);
nor NOR4 (N887, N851, N643, N678, N588);
xor XOR2 (N888, N887, N783);
nor NOR4 (N889, N882, N45, N477, N582);
and AND2 (N890, N886, N520);
not NOT1 (N891, N872);
nand NAND2 (N892, N864, N44);
buf BUF1 (N893, N888);
or OR4 (N894, N892, N761, N358, N531);
and AND4 (N895, N893, N116, N90, N35);
or OR4 (N896, N890, N143, N655, N180);
nand NAND2 (N897, N895, N389);
xor XOR2 (N898, N870, N383);
xor XOR2 (N899, N889, N404);
and AND4 (N900, N883, N34, N797, N729);
nor NOR3 (N901, N880, N499, N63);
xor XOR2 (N902, N891, N185);
nand NAND2 (N903, N894, N292);
xor XOR2 (N904, N901, N121);
and AND3 (N905, N899, N40, N756);
or OR3 (N906, N902, N612, N219);
or OR2 (N907, N904, N33);
nand NAND4 (N908, N907, N635, N269, N40);
not NOT1 (N909, N885);
xor XOR2 (N910, N903, N271);
buf BUF1 (N911, N900);
not NOT1 (N912, N909);
not NOT1 (N913, N910);
and AND2 (N914, N906, N276);
and AND2 (N915, N912, N293);
nor NOR2 (N916, N915, N788);
and AND2 (N917, N897, N241);
nand NAND3 (N918, N917, N115, N714);
or OR3 (N919, N879, N361, N14);
and AND4 (N920, N898, N233, N651, N663);
nor NOR4 (N921, N918, N619, N823, N261);
and AND2 (N922, N914, N268);
buf BUF1 (N923, N921);
xor XOR2 (N924, N916, N379);
and AND4 (N925, N911, N699, N340, N283);
and AND2 (N926, N905, N415);
xor XOR2 (N927, N919, N556);
buf BUF1 (N928, N920);
not NOT1 (N929, N927);
xor XOR2 (N930, N913, N389);
nand NAND4 (N931, N908, N672, N299, N21);
not NOT1 (N932, N931);
buf BUF1 (N933, N896);
nor NOR3 (N934, N925, N765, N760);
or OR4 (N935, N928, N271, N12, N373);
buf BUF1 (N936, N933);
or OR4 (N937, N935, N76, N883, N268);
not NOT1 (N938, N923);
and AND2 (N939, N932, N714);
and AND4 (N940, N934, N204, N442, N197);
or OR3 (N941, N940, N541, N410);
and AND2 (N942, N926, N29);
nor NOR2 (N943, N937, N144);
nor NOR4 (N944, N943, N795, N496, N90);
nand NAND4 (N945, N930, N839, N670, N341);
nand NAND2 (N946, N922, N371);
nor NOR2 (N947, N945, N412);
or OR4 (N948, N936, N367, N842, N222);
or OR3 (N949, N944, N403, N524);
xor XOR2 (N950, N949, N223);
nor NOR4 (N951, N938, N438, N672, N830);
and AND4 (N952, N942, N647, N232, N200);
not NOT1 (N953, N951);
and AND2 (N954, N946, N491);
nor NOR3 (N955, N950, N212, N294);
buf BUF1 (N956, N954);
or OR4 (N957, N955, N654, N164, N882);
nor NOR3 (N958, N941, N533, N945);
and AND2 (N959, N947, N624);
nor NOR4 (N960, N952, N120, N188, N108);
not NOT1 (N961, N924);
nand NAND2 (N962, N929, N235);
xor XOR2 (N963, N960, N513);
buf BUF1 (N964, N957);
buf BUF1 (N965, N964);
xor XOR2 (N966, N963, N514);
buf BUF1 (N967, N939);
not NOT1 (N968, N967);
not NOT1 (N969, N968);
and AND4 (N970, N956, N944, N482, N336);
xor XOR2 (N971, N953, N826);
nor NOR2 (N972, N959, N602);
xor XOR2 (N973, N962, N443);
and AND3 (N974, N970, N231, N264);
nor NOR3 (N975, N973, N852, N683);
or OR2 (N976, N975, N75);
not NOT1 (N977, N948);
xor XOR2 (N978, N971, N285);
nand NAND4 (N979, N965, N940, N382, N682);
and AND2 (N980, N979, N358);
nand NAND3 (N981, N978, N561, N556);
buf BUF1 (N982, N966);
nand NAND3 (N983, N969, N689, N282);
or OR3 (N984, N977, N220, N63);
or OR4 (N985, N984, N223, N342, N229);
nand NAND4 (N986, N985, N919, N676, N413);
buf BUF1 (N987, N974);
buf BUF1 (N988, N961);
and AND4 (N989, N986, N875, N909, N955);
xor XOR2 (N990, N972, N708);
not NOT1 (N991, N981);
nor NOR2 (N992, N983, N270);
and AND4 (N993, N980, N868, N115, N975);
xor XOR2 (N994, N987, N667);
buf BUF1 (N995, N990);
not NOT1 (N996, N995);
and AND3 (N997, N991, N584, N983);
not NOT1 (N998, N958);
not NOT1 (N999, N998);
xor XOR2 (N1000, N988, N174);
xor XOR2 (N1001, N994, N526);
or OR4 (N1002, N1001, N579, N426, N237);
xor XOR2 (N1003, N996, N276);
nand NAND2 (N1004, N1002, N635);
nand NAND2 (N1005, N1004, N57);
nor NOR4 (N1006, N982, N127, N247, N470);
or OR2 (N1007, N976, N314);
nand NAND2 (N1008, N999, N1001);
buf BUF1 (N1009, N992);
buf BUF1 (N1010, N1000);
not NOT1 (N1011, N989);
or OR2 (N1012, N1005, N972);
and AND2 (N1013, N1010, N825);
buf BUF1 (N1014, N1013);
or OR2 (N1015, N1006, N514);
nor NOR4 (N1016, N997, N686, N839, N235);
xor XOR2 (N1017, N1009, N281);
nor NOR4 (N1018, N1003, N256, N427, N518);
buf BUF1 (N1019, N1008);
nor NOR2 (N1020, N1014, N18);
buf BUF1 (N1021, N1018);
not NOT1 (N1022, N993);
buf BUF1 (N1023, N1016);
nand NAND2 (N1024, N1021, N349);
nor NOR4 (N1025, N1011, N398, N309, N721);
nor NOR3 (N1026, N1007, N528, N74);
and AND2 (N1027, N1012, N961);
nand NAND3 (N1028, N1025, N257, N867);
nand NAND2 (N1029, N1019, N366);
and AND2 (N1030, N1027, N47);
or OR4 (N1031, N1028, N709, N932, N195);
xor XOR2 (N1032, N1017, N986);
and AND4 (N1033, N1023, N691, N478, N11);
nor NOR4 (N1034, N1026, N680, N837, N98);
xor XOR2 (N1035, N1024, N509);
or OR4 (N1036, N1029, N90, N878, N745);
xor XOR2 (N1037, N1030, N387);
and AND4 (N1038, N1036, N376, N321, N1028);
and AND4 (N1039, N1037, N900, N618, N12);
not NOT1 (N1040, N1032);
buf BUF1 (N1041, N1038);
xor XOR2 (N1042, N1034, N63);
xor XOR2 (N1043, N1022, N977);
xor XOR2 (N1044, N1040, N638);
nand NAND4 (N1045, N1031, N743, N416, N696);
or OR2 (N1046, N1044, N595);
not NOT1 (N1047, N1035);
not NOT1 (N1048, N1015);
and AND3 (N1049, N1041, N789, N492);
not NOT1 (N1050, N1045);
and AND4 (N1051, N1020, N91, N814, N771);
buf BUF1 (N1052, N1047);
buf BUF1 (N1053, N1033);
and AND3 (N1054, N1048, N161, N269);
xor XOR2 (N1055, N1039, N131);
nor NOR3 (N1056, N1046, N580, N427);
not NOT1 (N1057, N1050);
buf BUF1 (N1058, N1049);
nand NAND4 (N1059, N1054, N502, N12, N184);
not NOT1 (N1060, N1058);
buf BUF1 (N1061, N1052);
nor NOR4 (N1062, N1043, N49, N41, N363);
nand NAND2 (N1063, N1051, N111);
or OR2 (N1064, N1061, N762);
not NOT1 (N1065, N1059);
xor XOR2 (N1066, N1056, N389);
not NOT1 (N1067, N1066);
xor XOR2 (N1068, N1053, N869);
xor XOR2 (N1069, N1057, N385);
xor XOR2 (N1070, N1068, N740);
nor NOR2 (N1071, N1065, N937);
nand NAND3 (N1072, N1070, N33, N178);
not NOT1 (N1073, N1042);
and AND2 (N1074, N1071, N253);
or OR4 (N1075, N1062, N1035, N321, N704);
nand NAND3 (N1076, N1055, N613, N999);
and AND2 (N1077, N1074, N918);
nand NAND3 (N1078, N1063, N937, N104);
not NOT1 (N1079, N1069);
nand NAND3 (N1080, N1079, N379, N170);
and AND2 (N1081, N1075, N1007);
or OR3 (N1082, N1076, N740, N628);
not NOT1 (N1083, N1064);
nor NOR4 (N1084, N1067, N196, N442, N445);
and AND2 (N1085, N1077, N801);
nand NAND2 (N1086, N1072, N230);
xor XOR2 (N1087, N1086, N727);
nand NAND2 (N1088, N1080, N982);
nand NAND2 (N1089, N1060, N347);
or OR2 (N1090, N1081, N962);
xor XOR2 (N1091, N1085, N351);
nor NOR2 (N1092, N1084, N826);
nand NAND2 (N1093, N1087, N971);
nor NOR2 (N1094, N1083, N637);
nor NOR4 (N1095, N1094, N13, N280, N62);
not NOT1 (N1096, N1091);
not NOT1 (N1097, N1082);
not NOT1 (N1098, N1093);
xor XOR2 (N1099, N1095, N286);
nor NOR2 (N1100, N1097, N302);
buf BUF1 (N1101, N1073);
not NOT1 (N1102, N1099);
xor XOR2 (N1103, N1088, N116);
nor NOR2 (N1104, N1103, N737);
nand NAND3 (N1105, N1096, N686, N313);
and AND3 (N1106, N1090, N18, N440);
xor XOR2 (N1107, N1101, N990);
not NOT1 (N1108, N1098);
nor NOR2 (N1109, N1108, N397);
and AND4 (N1110, N1107, N783, N945, N652);
nor NOR3 (N1111, N1106, N752, N820);
xor XOR2 (N1112, N1089, N100);
and AND2 (N1113, N1105, N393);
nand NAND2 (N1114, N1112, N685);
and AND2 (N1115, N1114, N767);
xor XOR2 (N1116, N1115, N634);
nand NAND4 (N1117, N1116, N866, N692, N943);
nand NAND4 (N1118, N1104, N292, N251, N255);
not NOT1 (N1119, N1109);
buf BUF1 (N1120, N1110);
or OR3 (N1121, N1117, N427, N319);
xor XOR2 (N1122, N1119, N531);
nand NAND2 (N1123, N1092, N47);
not NOT1 (N1124, N1078);
not NOT1 (N1125, N1118);
xor XOR2 (N1126, N1113, N953);
not NOT1 (N1127, N1122);
xor XOR2 (N1128, N1121, N144);
xor XOR2 (N1129, N1128, N723);
and AND2 (N1130, N1100, N991);
nor NOR3 (N1131, N1127, N1106, N450);
nand NAND4 (N1132, N1123, N749, N1086, N175);
xor XOR2 (N1133, N1126, N458);
xor XOR2 (N1134, N1120, N348);
buf BUF1 (N1135, N1130);
or OR4 (N1136, N1134, N730, N967, N1012);
xor XOR2 (N1137, N1136, N864);
nor NOR3 (N1138, N1124, N315, N160);
xor XOR2 (N1139, N1129, N698);
nor NOR2 (N1140, N1111, N355);
nand NAND3 (N1141, N1102, N1093, N1018);
nor NOR4 (N1142, N1141, N802, N616, N9);
and AND4 (N1143, N1138, N79, N256, N476);
nand NAND3 (N1144, N1137, N931, N180);
xor XOR2 (N1145, N1132, N426);
and AND2 (N1146, N1139, N265);
buf BUF1 (N1147, N1135);
xor XOR2 (N1148, N1142, N256);
buf BUF1 (N1149, N1140);
and AND2 (N1150, N1131, N55);
buf BUF1 (N1151, N1146);
xor XOR2 (N1152, N1147, N1056);
nor NOR3 (N1153, N1148, N980, N372);
nand NAND2 (N1154, N1143, N1018);
and AND4 (N1155, N1145, N560, N170, N7);
nand NAND4 (N1156, N1152, N123, N573, N874);
not NOT1 (N1157, N1154);
and AND3 (N1158, N1153, N836, N987);
xor XOR2 (N1159, N1144, N464);
buf BUF1 (N1160, N1158);
buf BUF1 (N1161, N1150);
and AND3 (N1162, N1159, N1048, N571);
or OR4 (N1163, N1162, N1004, N1022, N962);
buf BUF1 (N1164, N1160);
not NOT1 (N1165, N1156);
buf BUF1 (N1166, N1155);
nand NAND2 (N1167, N1165, N1117);
or OR3 (N1168, N1149, N438, N693);
not NOT1 (N1169, N1125);
or OR2 (N1170, N1168, N259);
buf BUF1 (N1171, N1151);
and AND2 (N1172, N1170, N704);
buf BUF1 (N1173, N1166);
and AND2 (N1174, N1169, N809);
buf BUF1 (N1175, N1133);
or OR2 (N1176, N1167, N724);
not NOT1 (N1177, N1172);
and AND2 (N1178, N1157, N246);
nor NOR4 (N1179, N1164, N901, N1092, N551);
buf BUF1 (N1180, N1175);
or OR4 (N1181, N1177, N281, N304, N1144);
nand NAND4 (N1182, N1174, N861, N96, N922);
nand NAND3 (N1183, N1180, N1020, N316);
nand NAND3 (N1184, N1171, N279, N909);
not NOT1 (N1185, N1183);
nand NAND3 (N1186, N1182, N997, N316);
nor NOR3 (N1187, N1186, N463, N707);
nand NAND2 (N1188, N1187, N569);
buf BUF1 (N1189, N1176);
xor XOR2 (N1190, N1184, N639);
and AND3 (N1191, N1173, N111, N1133);
not NOT1 (N1192, N1181);
not NOT1 (N1193, N1189);
nor NOR2 (N1194, N1192, N886);
xor XOR2 (N1195, N1178, N104);
xor XOR2 (N1196, N1193, N1011);
nor NOR3 (N1197, N1196, N663, N1120);
nor NOR2 (N1198, N1161, N942);
xor XOR2 (N1199, N1195, N898);
and AND4 (N1200, N1185, N171, N495, N9);
or OR3 (N1201, N1200, N1028, N591);
and AND4 (N1202, N1179, N35, N1178, N553);
buf BUF1 (N1203, N1198);
buf BUF1 (N1204, N1199);
and AND2 (N1205, N1194, N276);
nand NAND4 (N1206, N1205, N1175, N342, N748);
nor NOR4 (N1207, N1197, N1084, N351, N320);
and AND2 (N1208, N1191, N744);
or OR2 (N1209, N1202, N500);
nor NOR4 (N1210, N1209, N474, N452, N1075);
or OR4 (N1211, N1204, N27, N12, N16);
buf BUF1 (N1212, N1210);
nand NAND4 (N1213, N1207, N999, N728, N710);
nand NAND4 (N1214, N1190, N1212, N962, N82);
xor XOR2 (N1215, N556, N1131);
and AND4 (N1216, N1206, N1046, N333, N934);
xor XOR2 (N1217, N1215, N282);
or OR2 (N1218, N1163, N964);
not NOT1 (N1219, N1208);
or OR2 (N1220, N1216, N550);
and AND4 (N1221, N1203, N58, N222, N100);
buf BUF1 (N1222, N1220);
and AND2 (N1223, N1217, N233);
not NOT1 (N1224, N1218);
buf BUF1 (N1225, N1222);
and AND4 (N1226, N1219, N1056, N1191, N407);
nand NAND3 (N1227, N1224, N1031, N124);
and AND2 (N1228, N1188, N557);
nor NOR4 (N1229, N1221, N1000, N930, N839);
or OR2 (N1230, N1223, N387);
xor XOR2 (N1231, N1211, N1168);
nand NAND3 (N1232, N1230, N235, N16);
xor XOR2 (N1233, N1231, N1142);
buf BUF1 (N1234, N1229);
and AND4 (N1235, N1232, N100, N805, N997);
or OR2 (N1236, N1225, N1045);
xor XOR2 (N1237, N1214, N868);
not NOT1 (N1238, N1235);
nand NAND4 (N1239, N1237, N100, N199, N374);
and AND4 (N1240, N1233, N111, N391, N757);
buf BUF1 (N1241, N1201);
not NOT1 (N1242, N1234);
nor NOR4 (N1243, N1228, N768, N705, N13);
nand NAND2 (N1244, N1238, N305);
xor XOR2 (N1245, N1226, N753);
nor NOR3 (N1246, N1227, N660, N962);
nand NAND4 (N1247, N1245, N838, N912, N1034);
xor XOR2 (N1248, N1241, N1095);
buf BUF1 (N1249, N1247);
nor NOR2 (N1250, N1239, N554);
nand NAND2 (N1251, N1242, N1170);
or OR3 (N1252, N1236, N379, N1076);
or OR3 (N1253, N1244, N1009, N227);
xor XOR2 (N1254, N1249, N1109);
buf BUF1 (N1255, N1253);
and AND3 (N1256, N1251, N222, N1042);
not NOT1 (N1257, N1240);
not NOT1 (N1258, N1254);
and AND3 (N1259, N1255, N1084, N444);
nand NAND4 (N1260, N1256, N119, N319, N592);
nand NAND3 (N1261, N1246, N284, N889);
nand NAND2 (N1262, N1257, N380);
nand NAND4 (N1263, N1250, N982, N852, N949);
xor XOR2 (N1264, N1260, N1131);
or OR4 (N1265, N1259, N827, N174, N1091);
nand NAND3 (N1266, N1263, N780, N37);
or OR2 (N1267, N1248, N613);
nor NOR2 (N1268, N1267, N173);
or OR3 (N1269, N1213, N726, N433);
buf BUF1 (N1270, N1268);
buf BUF1 (N1271, N1258);
buf BUF1 (N1272, N1261);
or OR2 (N1273, N1271, N227);
xor XOR2 (N1274, N1270, N725);
xor XOR2 (N1275, N1274, N163);
nor NOR2 (N1276, N1243, N1122);
nand NAND4 (N1277, N1264, N1275, N179, N1181);
buf BUF1 (N1278, N654);
or OR2 (N1279, N1276, N1117);
nand NAND4 (N1280, N1265, N987, N66, N766);
nand NAND2 (N1281, N1280, N786);
xor XOR2 (N1282, N1277, N624);
or OR4 (N1283, N1279, N654, N1191, N822);
nor NOR3 (N1284, N1262, N421, N97);
nor NOR4 (N1285, N1272, N127, N639, N1268);
nor NOR3 (N1286, N1269, N1012, N378);
and AND4 (N1287, N1281, N211, N946, N215);
buf BUF1 (N1288, N1282);
nor NOR4 (N1289, N1288, N1006, N87, N625);
not NOT1 (N1290, N1273);
and AND3 (N1291, N1290, N969, N1092);
not NOT1 (N1292, N1252);
nand NAND3 (N1293, N1266, N20, N989);
nor NOR2 (N1294, N1285, N1136);
nor NOR4 (N1295, N1278, N555, N27, N713);
buf BUF1 (N1296, N1294);
not NOT1 (N1297, N1283);
not NOT1 (N1298, N1292);
and AND4 (N1299, N1297, N1099, N550, N1270);
and AND4 (N1300, N1291, N1002, N328, N992);
nor NOR3 (N1301, N1287, N376, N279);
or OR2 (N1302, N1284, N1264);
xor XOR2 (N1303, N1293, N752);
nand NAND4 (N1304, N1300, N312, N695, N564);
or OR4 (N1305, N1298, N694, N1163, N1060);
nand NAND3 (N1306, N1286, N758, N1052);
nand NAND4 (N1307, N1296, N1190, N810, N491);
buf BUF1 (N1308, N1299);
or OR4 (N1309, N1306, N778, N1186, N910);
nand NAND4 (N1310, N1309, N69, N1243, N1209);
buf BUF1 (N1311, N1303);
nor NOR2 (N1312, N1305, N576);
not NOT1 (N1313, N1301);
buf BUF1 (N1314, N1310);
nand NAND4 (N1315, N1312, N358, N935, N912);
not NOT1 (N1316, N1315);
nand NAND2 (N1317, N1314, N452);
buf BUF1 (N1318, N1307);
not NOT1 (N1319, N1308);
buf BUF1 (N1320, N1318);
buf BUF1 (N1321, N1304);
and AND4 (N1322, N1295, N111, N765, N1103);
not NOT1 (N1323, N1311);
not NOT1 (N1324, N1322);
and AND3 (N1325, N1321, N588, N59);
or OR2 (N1326, N1320, N922);
nand NAND2 (N1327, N1319, N1300);
nor NOR2 (N1328, N1289, N27);
xor XOR2 (N1329, N1328, N457);
xor XOR2 (N1330, N1325, N402);
nor NOR4 (N1331, N1323, N1308, N38, N1064);
nand NAND4 (N1332, N1316, N264, N619, N549);
nand NAND4 (N1333, N1302, N1162, N618, N618);
not NOT1 (N1334, N1317);
nand NAND3 (N1335, N1327, N399, N54);
not NOT1 (N1336, N1329);
and AND4 (N1337, N1332, N745, N794, N936);
buf BUF1 (N1338, N1336);
nor NOR4 (N1339, N1338, N971, N679, N1316);
xor XOR2 (N1340, N1313, N1332);
not NOT1 (N1341, N1333);
xor XOR2 (N1342, N1326, N280);
buf BUF1 (N1343, N1331);
xor XOR2 (N1344, N1334, N936);
buf BUF1 (N1345, N1342);
buf BUF1 (N1346, N1337);
xor XOR2 (N1347, N1346, N976);
xor XOR2 (N1348, N1335, N197);
buf BUF1 (N1349, N1347);
and AND3 (N1350, N1324, N269, N781);
xor XOR2 (N1351, N1350, N779);
nand NAND3 (N1352, N1340, N841, N1317);
nor NOR3 (N1353, N1344, N713, N1250);
and AND2 (N1354, N1330, N41);
xor XOR2 (N1355, N1351, N942);
not NOT1 (N1356, N1341);
buf BUF1 (N1357, N1354);
buf BUF1 (N1358, N1343);
or OR4 (N1359, N1345, N1281, N506, N822);
or OR2 (N1360, N1353, N569);
nor NOR3 (N1361, N1355, N1052, N364);
and AND4 (N1362, N1360, N927, N265, N539);
not NOT1 (N1363, N1362);
or OR4 (N1364, N1358, N248, N907, N1221);
nand NAND3 (N1365, N1348, N1010, N840);
and AND2 (N1366, N1361, N225);
or OR3 (N1367, N1356, N1151, N963);
nor NOR3 (N1368, N1367, N137, N369);
not NOT1 (N1369, N1366);
xor XOR2 (N1370, N1352, N510);
or OR2 (N1371, N1359, N401);
or OR2 (N1372, N1371, N1309);
buf BUF1 (N1373, N1349);
nand NAND3 (N1374, N1357, N858, N44);
xor XOR2 (N1375, N1365, N214);
and AND3 (N1376, N1339, N919, N1098);
xor XOR2 (N1377, N1373, N1165);
buf BUF1 (N1378, N1375);
nand NAND4 (N1379, N1377, N625, N665, N1129);
not NOT1 (N1380, N1363);
and AND4 (N1381, N1378, N239, N991, N224);
not NOT1 (N1382, N1376);
buf BUF1 (N1383, N1380);
or OR4 (N1384, N1372, N1330, N727, N759);
and AND3 (N1385, N1384, N437, N1371);
not NOT1 (N1386, N1369);
or OR2 (N1387, N1382, N1255);
not NOT1 (N1388, N1387);
nand NAND4 (N1389, N1381, N690, N934, N494);
not NOT1 (N1390, N1386);
buf BUF1 (N1391, N1370);
xor XOR2 (N1392, N1368, N1110);
not NOT1 (N1393, N1364);
not NOT1 (N1394, N1389);
buf BUF1 (N1395, N1393);
or OR3 (N1396, N1395, N359, N762);
nor NOR3 (N1397, N1379, N53, N1193);
nand NAND3 (N1398, N1391, N1008, N1135);
xor XOR2 (N1399, N1392, N224);
nor NOR3 (N1400, N1374, N1260, N865);
buf BUF1 (N1401, N1394);
nand NAND2 (N1402, N1388, N1261);
or OR3 (N1403, N1383, N321, N800);
nand NAND3 (N1404, N1400, N1094, N522);
or OR4 (N1405, N1398, N734, N648, N277);
nand NAND2 (N1406, N1402, N621);
nand NAND4 (N1407, N1397, N1308, N1112, N640);
nor NOR2 (N1408, N1407, N284);
and AND2 (N1409, N1408, N636);
or OR4 (N1410, N1409, N1105, N338, N794);
buf BUF1 (N1411, N1396);
xor XOR2 (N1412, N1410, N633);
not NOT1 (N1413, N1385);
nor NOR2 (N1414, N1406, N937);
nor NOR2 (N1415, N1413, N705);
not NOT1 (N1416, N1415);
buf BUF1 (N1417, N1403);
or OR4 (N1418, N1404, N516, N229, N1244);
not NOT1 (N1419, N1417);
buf BUF1 (N1420, N1401);
buf BUF1 (N1421, N1416);
and AND4 (N1422, N1420, N543, N289, N1420);
xor XOR2 (N1423, N1422, N942);
xor XOR2 (N1424, N1399, N1318);
nor NOR4 (N1425, N1411, N190, N1184, N1165);
and AND2 (N1426, N1425, N840);
not NOT1 (N1427, N1421);
or OR2 (N1428, N1412, N581);
nand NAND2 (N1429, N1426, N221);
xor XOR2 (N1430, N1419, N574);
nor NOR4 (N1431, N1424, N1057, N231, N152);
or OR2 (N1432, N1430, N792);
or OR3 (N1433, N1428, N653, N376);
and AND2 (N1434, N1423, N874);
xor XOR2 (N1435, N1432, N792);
nor NOR3 (N1436, N1431, N860, N433);
nor NOR2 (N1437, N1414, N766);
xor XOR2 (N1438, N1435, N1074);
nor NOR4 (N1439, N1437, N1340, N449, N1071);
xor XOR2 (N1440, N1436, N1195);
xor XOR2 (N1441, N1439, N1279);
not NOT1 (N1442, N1440);
and AND4 (N1443, N1442, N926, N986, N1020);
nor NOR2 (N1444, N1434, N1009);
not NOT1 (N1445, N1444);
and AND4 (N1446, N1443, N916, N516, N821);
not NOT1 (N1447, N1445);
xor XOR2 (N1448, N1446, N754);
or OR2 (N1449, N1390, N1044);
or OR2 (N1450, N1441, N508);
and AND4 (N1451, N1418, N1228, N230, N1388);
xor XOR2 (N1452, N1438, N112);
xor XOR2 (N1453, N1449, N25);
nor NOR2 (N1454, N1447, N1400);
and AND4 (N1455, N1405, N117, N194, N340);
and AND2 (N1456, N1451, N466);
or OR3 (N1457, N1454, N1387, N748);
not NOT1 (N1458, N1453);
nand NAND2 (N1459, N1427, N867);
nand NAND3 (N1460, N1459, N530, N1074);
nand NAND4 (N1461, N1460, N1060, N1302, N1151);
not NOT1 (N1462, N1429);
and AND3 (N1463, N1461, N324, N439);
nand NAND2 (N1464, N1463, N647);
xor XOR2 (N1465, N1455, N1189);
or OR4 (N1466, N1465, N866, N253, N454);
xor XOR2 (N1467, N1456, N279);
not NOT1 (N1468, N1450);
nand NAND4 (N1469, N1452, N409, N1162, N1444);
or OR4 (N1470, N1462, N653, N847, N736);
buf BUF1 (N1471, N1469);
nand NAND4 (N1472, N1471, N457, N245, N1039);
buf BUF1 (N1473, N1466);
or OR2 (N1474, N1464, N1083);
nand NAND2 (N1475, N1433, N731);
or OR3 (N1476, N1457, N759, N1155);
xor XOR2 (N1477, N1475, N1054);
and AND4 (N1478, N1448, N23, N1065, N1196);
nand NAND4 (N1479, N1472, N1083, N548, N1276);
nor NOR2 (N1480, N1479, N910);
nand NAND2 (N1481, N1468, N1348);
nor NOR2 (N1482, N1477, N90);
xor XOR2 (N1483, N1473, N217);
nand NAND2 (N1484, N1476, N1330);
not NOT1 (N1485, N1480);
or OR2 (N1486, N1481, N688);
or OR2 (N1487, N1478, N410);
or OR4 (N1488, N1487, N455, N1166, N987);
not NOT1 (N1489, N1470);
or OR2 (N1490, N1467, N546);
nand NAND2 (N1491, N1488, N513);
buf BUF1 (N1492, N1484);
nand NAND4 (N1493, N1492, N305, N835, N240);
and AND2 (N1494, N1491, N1165);
xor XOR2 (N1495, N1493, N692);
and AND2 (N1496, N1490, N172);
xor XOR2 (N1497, N1485, N66);
nor NOR3 (N1498, N1482, N512, N358);
buf BUF1 (N1499, N1486);
nor NOR4 (N1500, N1489, N349, N99, N586);
nand NAND3 (N1501, N1458, N609, N281);
or OR2 (N1502, N1494, N1404);
and AND3 (N1503, N1495, N319, N1031);
buf BUF1 (N1504, N1498);
buf BUF1 (N1505, N1500);
buf BUF1 (N1506, N1497);
nor NOR2 (N1507, N1474, N793);
nand NAND4 (N1508, N1504, N1128, N909, N772);
or OR4 (N1509, N1499, N147, N755, N653);
or OR2 (N1510, N1502, N89);
not NOT1 (N1511, N1508);
nor NOR4 (N1512, N1496, N1131, N1207, N777);
not NOT1 (N1513, N1505);
nor NOR3 (N1514, N1509, N1388, N431);
or OR3 (N1515, N1483, N958, N1156);
nor NOR3 (N1516, N1512, N524, N400);
xor XOR2 (N1517, N1513, N11);
nor NOR2 (N1518, N1507, N996);
buf BUF1 (N1519, N1517);
buf BUF1 (N1520, N1503);
not NOT1 (N1521, N1511);
nand NAND3 (N1522, N1519, N1123, N345);
and AND3 (N1523, N1501, N799, N1229);
xor XOR2 (N1524, N1506, N163);
not NOT1 (N1525, N1518);
nand NAND3 (N1526, N1523, N1143, N1211);
xor XOR2 (N1527, N1525, N806);
nand NAND4 (N1528, N1510, N973, N898, N702);
xor XOR2 (N1529, N1514, N287);
and AND4 (N1530, N1528, N468, N1100, N1364);
buf BUF1 (N1531, N1516);
buf BUF1 (N1532, N1526);
or OR2 (N1533, N1530, N1297);
not NOT1 (N1534, N1529);
not NOT1 (N1535, N1534);
nor NOR3 (N1536, N1522, N117, N548);
not NOT1 (N1537, N1520);
nor NOR4 (N1538, N1515, N74, N850, N413);
xor XOR2 (N1539, N1521, N300);
and AND3 (N1540, N1533, N1480, N838);
buf BUF1 (N1541, N1536);
nor NOR2 (N1542, N1535, N479);
or OR3 (N1543, N1542, N981, N891);
buf BUF1 (N1544, N1532);
nand NAND2 (N1545, N1538, N566);
or OR4 (N1546, N1541, N1033, N112, N798);
nand NAND2 (N1547, N1544, N990);
buf BUF1 (N1548, N1543);
xor XOR2 (N1549, N1547, N84);
nand NAND3 (N1550, N1537, N40, N1512);
xor XOR2 (N1551, N1524, N1293);
or OR3 (N1552, N1546, N131, N119);
xor XOR2 (N1553, N1545, N212);
not NOT1 (N1554, N1552);
and AND4 (N1555, N1548, N1447, N1364, N912);
xor XOR2 (N1556, N1551, N683);
nor NOR3 (N1557, N1553, N1356, N15);
xor XOR2 (N1558, N1549, N1131);
not NOT1 (N1559, N1531);
xor XOR2 (N1560, N1557, N1377);
nor NOR2 (N1561, N1540, N1516);
nand NAND4 (N1562, N1558, N320, N1081, N1061);
buf BUF1 (N1563, N1562);
buf BUF1 (N1564, N1561);
nor NOR3 (N1565, N1539, N180, N1271);
buf BUF1 (N1566, N1559);
nand NAND2 (N1567, N1554, N119);
and AND2 (N1568, N1567, N1353);
and AND4 (N1569, N1566, N16, N1341, N1522);
buf BUF1 (N1570, N1564);
or OR3 (N1571, N1527, N1542, N1379);
and AND2 (N1572, N1563, N727);
or OR3 (N1573, N1556, N126, N1553);
nor NOR4 (N1574, N1570, N324, N1297, N1071);
and AND3 (N1575, N1550, N515, N1223);
nor NOR4 (N1576, N1574, N1479, N1549, N467);
nand NAND4 (N1577, N1573, N600, N1286, N1066);
xor XOR2 (N1578, N1560, N211);
nor NOR4 (N1579, N1571, N463, N575, N1238);
and AND4 (N1580, N1568, N111, N1225, N1307);
or OR3 (N1581, N1580, N32, N947);
not NOT1 (N1582, N1555);
xor XOR2 (N1583, N1565, N755);
nand NAND4 (N1584, N1572, N1053, N967, N1343);
or OR2 (N1585, N1577, N111);
or OR2 (N1586, N1584, N461);
buf BUF1 (N1587, N1583);
or OR3 (N1588, N1569, N1260, N612);
nor NOR4 (N1589, N1579, N307, N810, N24);
not NOT1 (N1590, N1582);
buf BUF1 (N1591, N1587);
xor XOR2 (N1592, N1585, N266);
xor XOR2 (N1593, N1588, N271);
nand NAND4 (N1594, N1586, N1296, N1351, N153);
buf BUF1 (N1595, N1593);
and AND3 (N1596, N1589, N560, N844);
buf BUF1 (N1597, N1592);
buf BUF1 (N1598, N1578);
xor XOR2 (N1599, N1595, N655);
not NOT1 (N1600, N1576);
buf BUF1 (N1601, N1598);
nor NOR4 (N1602, N1597, N51, N704, N1162);
not NOT1 (N1603, N1601);
buf BUF1 (N1604, N1602);
not NOT1 (N1605, N1590);
and AND2 (N1606, N1594, N344);
not NOT1 (N1607, N1581);
and AND2 (N1608, N1604, N1527);
buf BUF1 (N1609, N1606);
and AND4 (N1610, N1607, N429, N586, N1007);
nor NOR3 (N1611, N1591, N59, N419);
and AND2 (N1612, N1609, N68);
or OR3 (N1613, N1611, N1357, N588);
buf BUF1 (N1614, N1603);
buf BUF1 (N1615, N1612);
and AND2 (N1616, N1610, N1566);
not NOT1 (N1617, N1605);
and AND3 (N1618, N1615, N1602, N448);
or OR2 (N1619, N1599, N30);
buf BUF1 (N1620, N1617);
or OR3 (N1621, N1596, N361, N1096);
nand NAND4 (N1622, N1575, N631, N715, N161);
nor NOR2 (N1623, N1618, N94);
xor XOR2 (N1624, N1623, N1462);
or OR3 (N1625, N1613, N407, N378);
nand NAND3 (N1626, N1624, N852, N365);
not NOT1 (N1627, N1620);
not NOT1 (N1628, N1616);
or OR3 (N1629, N1608, N1546, N1206);
buf BUF1 (N1630, N1628);
nor NOR4 (N1631, N1619, N374, N1603, N1348);
or OR3 (N1632, N1621, N1610, N678);
nor NOR4 (N1633, N1625, N1210, N1083, N175);
and AND2 (N1634, N1629, N227);
and AND2 (N1635, N1631, N1138);
buf BUF1 (N1636, N1633);
xor XOR2 (N1637, N1632, N1493);
nor NOR4 (N1638, N1635, N90, N1560, N520);
nor NOR3 (N1639, N1630, N365, N1574);
nor NOR4 (N1640, N1634, N403, N1451, N1322);
xor XOR2 (N1641, N1640, N641);
not NOT1 (N1642, N1638);
nor NOR4 (N1643, N1600, N248, N150, N906);
not NOT1 (N1644, N1627);
nand NAND3 (N1645, N1642, N675, N1146);
and AND4 (N1646, N1644, N1015, N1497, N16);
nand NAND2 (N1647, N1641, N1608);
buf BUF1 (N1648, N1645);
or OR2 (N1649, N1626, N1297);
nor NOR4 (N1650, N1639, N126, N1126, N1499);
nand NAND3 (N1651, N1648, N919, N1585);
and AND3 (N1652, N1636, N1314, N269);
not NOT1 (N1653, N1651);
buf BUF1 (N1654, N1622);
xor XOR2 (N1655, N1647, N127);
nor NOR2 (N1656, N1614, N920);
buf BUF1 (N1657, N1652);
nand NAND3 (N1658, N1654, N19, N806);
or OR4 (N1659, N1653, N340, N1437, N625);
and AND3 (N1660, N1658, N1153, N845);
not NOT1 (N1661, N1637);
not NOT1 (N1662, N1657);
nand NAND2 (N1663, N1655, N1241);
and AND4 (N1664, N1650, N245, N1333, N1052);
nand NAND2 (N1665, N1663, N693);
buf BUF1 (N1666, N1659);
xor XOR2 (N1667, N1666, N1107);
nor NOR3 (N1668, N1665, N444, N586);
nor NOR4 (N1669, N1660, N472, N1183, N685);
not NOT1 (N1670, N1667);
nand NAND2 (N1671, N1643, N1214);
buf BUF1 (N1672, N1670);
nor NOR4 (N1673, N1646, N217, N1262, N365);
buf BUF1 (N1674, N1656);
or OR3 (N1675, N1664, N687, N250);
and AND4 (N1676, N1661, N935, N486, N1664);
and AND3 (N1677, N1671, N794, N152);
nand NAND4 (N1678, N1672, N185, N1659, N617);
xor XOR2 (N1679, N1649, N275);
nor NOR4 (N1680, N1676, N705, N829, N828);
buf BUF1 (N1681, N1674);
xor XOR2 (N1682, N1679, N68);
and AND3 (N1683, N1673, N795, N1398);
buf BUF1 (N1684, N1678);
xor XOR2 (N1685, N1681, N388);
or OR3 (N1686, N1669, N562, N1340);
buf BUF1 (N1687, N1682);
and AND2 (N1688, N1683, N758);
nor NOR4 (N1689, N1668, N1394, N538, N1404);
buf BUF1 (N1690, N1689);
or OR4 (N1691, N1685, N777, N102, N541);
or OR4 (N1692, N1687, N117, N1070, N999);
or OR4 (N1693, N1684, N376, N445, N964);
nor NOR3 (N1694, N1693, N909, N1505);
nand NAND2 (N1695, N1677, N1333);
xor XOR2 (N1696, N1695, N845);
nand NAND3 (N1697, N1675, N183, N199);
not NOT1 (N1698, N1688);
or OR3 (N1699, N1698, N1284, N743);
nor NOR4 (N1700, N1691, N1437, N495, N870);
nor NOR3 (N1701, N1680, N168, N1126);
nor NOR2 (N1702, N1696, N515);
nand NAND2 (N1703, N1697, N1430);
nand NAND3 (N1704, N1701, N1406, N1071);
xor XOR2 (N1705, N1700, N637);
xor XOR2 (N1706, N1699, N80);
or OR2 (N1707, N1704, N124);
not NOT1 (N1708, N1706);
or OR2 (N1709, N1703, N1028);
or OR2 (N1710, N1692, N197);
xor XOR2 (N1711, N1705, N913);
not NOT1 (N1712, N1690);
or OR2 (N1713, N1662, N16);
not NOT1 (N1714, N1709);
or OR3 (N1715, N1712, N462, N507);
not NOT1 (N1716, N1710);
nand NAND3 (N1717, N1707, N655, N939);
nor NOR2 (N1718, N1711, N983);
or OR3 (N1719, N1715, N1354, N504);
nand NAND2 (N1720, N1714, N1013);
buf BUF1 (N1721, N1708);
xor XOR2 (N1722, N1713, N1012);
buf BUF1 (N1723, N1716);
xor XOR2 (N1724, N1721, N1269);
xor XOR2 (N1725, N1723, N1503);
nand NAND4 (N1726, N1717, N22, N145, N239);
nand NAND4 (N1727, N1726, N349, N1617, N1258);
nand NAND4 (N1728, N1686, N755, N1109, N1306);
or OR2 (N1729, N1694, N1234);
nand NAND2 (N1730, N1724, N353);
not NOT1 (N1731, N1728);
nor NOR2 (N1732, N1720, N1303);
not NOT1 (N1733, N1732);
or OR2 (N1734, N1719, N1102);
xor XOR2 (N1735, N1725, N457);
buf BUF1 (N1736, N1729);
and AND2 (N1737, N1722, N1314);
xor XOR2 (N1738, N1736, N331);
nand NAND4 (N1739, N1718, N1709, N1027, N748);
buf BUF1 (N1740, N1735);
not NOT1 (N1741, N1727);
not NOT1 (N1742, N1738);
and AND3 (N1743, N1741, N786, N1501);
and AND4 (N1744, N1739, N696, N847, N107);
nor NOR2 (N1745, N1743, N158);
or OR3 (N1746, N1734, N1156, N945);
buf BUF1 (N1747, N1733);
nor NOR2 (N1748, N1747, N1541);
buf BUF1 (N1749, N1731);
xor XOR2 (N1750, N1744, N589);
buf BUF1 (N1751, N1746);
nor NOR4 (N1752, N1740, N762, N908, N31);
or OR4 (N1753, N1742, N815, N1001, N1133);
nor NOR3 (N1754, N1748, N65, N196);
buf BUF1 (N1755, N1730);
or OR4 (N1756, N1754, N505, N1288, N598);
or OR4 (N1757, N1702, N1729, N631, N1323);
and AND2 (N1758, N1753, N89);
buf BUF1 (N1759, N1745);
or OR3 (N1760, N1755, N223, N327);
not NOT1 (N1761, N1751);
or OR2 (N1762, N1749, N920);
buf BUF1 (N1763, N1737);
buf BUF1 (N1764, N1756);
buf BUF1 (N1765, N1761);
nand NAND4 (N1766, N1764, N1619, N79, N1094);
buf BUF1 (N1767, N1759);
or OR2 (N1768, N1760, N518);
not NOT1 (N1769, N1763);
not NOT1 (N1770, N1768);
buf BUF1 (N1771, N1758);
buf BUF1 (N1772, N1765);
not NOT1 (N1773, N1750);
xor XOR2 (N1774, N1769, N7);
nand NAND3 (N1775, N1767, N412, N1427);
buf BUF1 (N1776, N1752);
xor XOR2 (N1777, N1762, N1685);
nor NOR3 (N1778, N1777, N1275, N1630);
nand NAND2 (N1779, N1776, N253);
and AND4 (N1780, N1771, N818, N1, N1067);
or OR3 (N1781, N1780, N43, N1100);
nand NAND2 (N1782, N1770, N1184);
nand NAND4 (N1783, N1775, N131, N1039, N1635);
and AND2 (N1784, N1774, N290);
or OR3 (N1785, N1773, N183, N231);
nor NOR3 (N1786, N1783, N142, N777);
and AND4 (N1787, N1784, N468, N1036, N150);
and AND4 (N1788, N1766, N261, N827, N1225);
or OR4 (N1789, N1781, N1150, N1516, N479);
or OR3 (N1790, N1786, N1171, N1729);
buf BUF1 (N1791, N1757);
xor XOR2 (N1792, N1782, N1655);
nor NOR4 (N1793, N1785, N1748, N588, N1444);
nor NOR3 (N1794, N1788, N995, N60);
not NOT1 (N1795, N1787);
not NOT1 (N1796, N1792);
and AND3 (N1797, N1791, N341, N1480);
xor XOR2 (N1798, N1794, N920);
or OR2 (N1799, N1790, N1268);
nand NAND2 (N1800, N1789, N1678);
and AND3 (N1801, N1793, N647, N115);
xor XOR2 (N1802, N1778, N121);
buf BUF1 (N1803, N1801);
xor XOR2 (N1804, N1803, N1730);
not NOT1 (N1805, N1799);
not NOT1 (N1806, N1772);
nand NAND4 (N1807, N1804, N324, N1245, N9);
nor NOR2 (N1808, N1806, N1345);
or OR2 (N1809, N1795, N1221);
not NOT1 (N1810, N1807);
buf BUF1 (N1811, N1808);
not NOT1 (N1812, N1805);
nor NOR4 (N1813, N1779, N1092, N366, N492);
xor XOR2 (N1814, N1797, N1162);
and AND2 (N1815, N1800, N1480);
and AND4 (N1816, N1814, N745, N1204, N1247);
buf BUF1 (N1817, N1812);
or OR3 (N1818, N1817, N764, N477);
and AND3 (N1819, N1810, N1720, N423);
and AND2 (N1820, N1809, N652);
nand NAND2 (N1821, N1813, N954);
not NOT1 (N1822, N1815);
not NOT1 (N1823, N1818);
buf BUF1 (N1824, N1798);
buf BUF1 (N1825, N1824);
xor XOR2 (N1826, N1823, N968);
nand NAND2 (N1827, N1796, N887);
not NOT1 (N1828, N1825);
not NOT1 (N1829, N1816);
nor NOR2 (N1830, N1829, N1251);
not NOT1 (N1831, N1820);
nor NOR3 (N1832, N1830, N815, N409);
and AND2 (N1833, N1802, N1301);
or OR2 (N1834, N1819, N760);
nand NAND3 (N1835, N1821, N715, N228);
buf BUF1 (N1836, N1832);
or OR2 (N1837, N1836, N1791);
xor XOR2 (N1838, N1827, N234);
not NOT1 (N1839, N1835);
not NOT1 (N1840, N1826);
and AND3 (N1841, N1828, N1450, N342);
xor XOR2 (N1842, N1831, N1312);
xor XOR2 (N1843, N1841, N71);
and AND3 (N1844, N1837, N1154, N1352);
nand NAND3 (N1845, N1842, N1373, N1154);
buf BUF1 (N1846, N1834);
buf BUF1 (N1847, N1846);
buf BUF1 (N1848, N1847);
nand NAND3 (N1849, N1839, N774, N891);
nor NOR2 (N1850, N1849, N1026);
nor NOR2 (N1851, N1838, N252);
nand NAND2 (N1852, N1845, N1072);
nand NAND3 (N1853, N1848, N769, N109);
and AND4 (N1854, N1811, N231, N760, N1121);
nand NAND3 (N1855, N1833, N884, N1769);
xor XOR2 (N1856, N1850, N1753);
nor NOR4 (N1857, N1840, N381, N1378, N261);
or OR3 (N1858, N1851, N1090, N1424);
nor NOR4 (N1859, N1855, N1258, N179, N606);
xor XOR2 (N1860, N1854, N1063);
or OR3 (N1861, N1857, N89, N318);
and AND2 (N1862, N1858, N216);
buf BUF1 (N1863, N1843);
xor XOR2 (N1864, N1852, N752);
and AND4 (N1865, N1859, N965, N1749, N765);
nand NAND3 (N1866, N1856, N590, N1634);
or OR2 (N1867, N1860, N1584);
not NOT1 (N1868, N1853);
buf BUF1 (N1869, N1863);
and AND3 (N1870, N1868, N888, N1137);
nand NAND4 (N1871, N1869, N1274, N1229, N1183);
nand NAND4 (N1872, N1864, N189, N1848, N941);
not NOT1 (N1873, N1870);
and AND3 (N1874, N1865, N1407, N1655);
nor NOR3 (N1875, N1862, N1164, N799);
xor XOR2 (N1876, N1871, N268);
xor XOR2 (N1877, N1875, N1159);
xor XOR2 (N1878, N1877, N882);
or OR4 (N1879, N1873, N1788, N985, N529);
xor XOR2 (N1880, N1872, N308);
not NOT1 (N1881, N1861);
nand NAND2 (N1882, N1880, N1819);
xor XOR2 (N1883, N1822, N1754);
xor XOR2 (N1884, N1881, N1676);
and AND2 (N1885, N1867, N143);
not NOT1 (N1886, N1884);
not NOT1 (N1887, N1879);
buf BUF1 (N1888, N1886);
or OR4 (N1889, N1866, N694, N1650, N841);
nor NOR3 (N1890, N1885, N1136, N1640);
and AND3 (N1891, N1844, N680, N1801);
nand NAND2 (N1892, N1876, N1858);
not NOT1 (N1893, N1878);
nand NAND4 (N1894, N1887, N601, N241, N553);
buf BUF1 (N1895, N1889);
xor XOR2 (N1896, N1895, N485);
not NOT1 (N1897, N1896);
buf BUF1 (N1898, N1874);
or OR2 (N1899, N1893, N353);
nand NAND2 (N1900, N1883, N467);
or OR3 (N1901, N1897, N1004, N364);
and AND3 (N1902, N1888, N741, N410);
and AND3 (N1903, N1901, N796, N404);
and AND4 (N1904, N1894, N1691, N946, N429);
buf BUF1 (N1905, N1900);
buf BUF1 (N1906, N1903);
or OR3 (N1907, N1899, N1842, N889);
or OR4 (N1908, N1882, N897, N387, N37);
and AND4 (N1909, N1906, N1785, N1543, N687);
or OR3 (N1910, N1890, N1741, N1048);
nand NAND4 (N1911, N1907, N1330, N403, N814);
not NOT1 (N1912, N1905);
not NOT1 (N1913, N1902);
xor XOR2 (N1914, N1908, N1754);
and AND3 (N1915, N1909, N1037, N160);
nor NOR2 (N1916, N1913, N205);
and AND3 (N1917, N1904, N1521, N361);
or OR4 (N1918, N1910, N1586, N1102, N1202);
and AND4 (N1919, N1912, N462, N1822, N644);
and AND3 (N1920, N1892, N345, N691);
buf BUF1 (N1921, N1920);
nor NOR2 (N1922, N1916, N1670);
or OR4 (N1923, N1891, N194, N1718, N1169);
xor XOR2 (N1924, N1919, N1707);
not NOT1 (N1925, N1918);
not NOT1 (N1926, N1921);
buf BUF1 (N1927, N1898);
nand NAND3 (N1928, N1917, N1496, N240);
nand NAND2 (N1929, N1911, N121);
not NOT1 (N1930, N1925);
xor XOR2 (N1931, N1922, N1274);
not NOT1 (N1932, N1929);
nor NOR2 (N1933, N1926, N1218);
xor XOR2 (N1934, N1932, N1619);
xor XOR2 (N1935, N1934, N1122);
buf BUF1 (N1936, N1933);
and AND4 (N1937, N1927, N1894, N335, N1924);
nor NOR2 (N1938, N1782, N245);
nor NOR2 (N1939, N1914, N147);
nand NAND3 (N1940, N1939, N23, N432);
nand NAND2 (N1941, N1930, N5);
or OR3 (N1942, N1938, N310, N1095);
nand NAND3 (N1943, N1923, N115, N983);
nand NAND3 (N1944, N1940, N196, N7);
nand NAND2 (N1945, N1944, N711);
not NOT1 (N1946, N1937);
nor NOR2 (N1947, N1943, N539);
xor XOR2 (N1948, N1942, N1645);
not NOT1 (N1949, N1948);
or OR2 (N1950, N1931, N863);
or OR2 (N1951, N1928, N872);
not NOT1 (N1952, N1949);
not NOT1 (N1953, N1947);
not NOT1 (N1954, N1915);
nand NAND3 (N1955, N1954, N961, N1114);
not NOT1 (N1956, N1950);
and AND4 (N1957, N1946, N1888, N22, N1350);
buf BUF1 (N1958, N1953);
or OR4 (N1959, N1941, N1302, N1680, N1833);
not NOT1 (N1960, N1959);
buf BUF1 (N1961, N1960);
nand NAND3 (N1962, N1956, N401, N727);
nand NAND4 (N1963, N1935, N1422, N532, N767);
buf BUF1 (N1964, N1957);
nor NOR2 (N1965, N1964, N1103);
nor NOR2 (N1966, N1961, N1416);
or OR3 (N1967, N1962, N601, N18);
not NOT1 (N1968, N1967);
not NOT1 (N1969, N1936);
buf BUF1 (N1970, N1963);
and AND2 (N1971, N1969, N1277);
nand NAND3 (N1972, N1965, N339, N202);
or OR2 (N1973, N1971, N1946);
xor XOR2 (N1974, N1966, N98);
not NOT1 (N1975, N1951);
and AND2 (N1976, N1974, N1676);
buf BUF1 (N1977, N1945);
nor NOR4 (N1978, N1952, N285, N1851, N1115);
not NOT1 (N1979, N1968);
and AND3 (N1980, N1972, N699, N773);
and AND3 (N1981, N1977, N376, N1757);
and AND2 (N1982, N1975, N322);
nand NAND4 (N1983, N1955, N1174, N315, N1950);
buf BUF1 (N1984, N1973);
or OR2 (N1985, N1978, N40);
not NOT1 (N1986, N1983);
nand NAND4 (N1987, N1976, N547, N769, N806);
and AND3 (N1988, N1980, N1959, N507);
buf BUF1 (N1989, N1984);
buf BUF1 (N1990, N1982);
nand NAND2 (N1991, N1990, N27);
and AND3 (N1992, N1970, N1241, N221);
nand NAND4 (N1993, N1985, N1755, N1903, N1064);
or OR2 (N1994, N1958, N994);
xor XOR2 (N1995, N1993, N812);
nor NOR4 (N1996, N1995, N1220, N656, N163);
nor NOR4 (N1997, N1981, N1026, N746, N546);
nor NOR4 (N1998, N1997, N1411, N1603, N1606);
not NOT1 (N1999, N1989);
buf BUF1 (N2000, N1991);
or OR4 (N2001, N1987, N1139, N664, N655);
or OR2 (N2002, N2001, N1700);
not NOT1 (N2003, N2000);
not NOT1 (N2004, N1998);
xor XOR2 (N2005, N1979, N1939);
nand NAND4 (N2006, N1986, N1331, N786, N1086);
nand NAND2 (N2007, N2005, N870);
nand NAND2 (N2008, N1988, N449);
nand NAND2 (N2009, N1994, N556);
or OR4 (N2010, N2003, N1057, N1465, N1655);
nor NOR4 (N2011, N2008, N852, N545, N1776);
or OR2 (N2012, N2006, N181);
nor NOR4 (N2013, N2010, N498, N1060, N1598);
or OR4 (N2014, N1992, N409, N1766, N1915);
nor NOR2 (N2015, N1999, N854);
xor XOR2 (N2016, N2014, N1281);
xor XOR2 (N2017, N2002, N99);
not NOT1 (N2018, N2015);
nand NAND4 (N2019, N2017, N990, N936, N1021);
nand NAND3 (N2020, N2011, N536, N643);
buf BUF1 (N2021, N2020);
or OR3 (N2022, N2013, N1327, N1418);
or OR4 (N2023, N2018, N528, N1712, N654);
nand NAND2 (N2024, N2004, N671);
and AND2 (N2025, N2019, N456);
and AND4 (N2026, N1996, N1992, N177, N805);
and AND4 (N2027, N2023, N1020, N932, N905);
not NOT1 (N2028, N2027);
and AND3 (N2029, N2025, N1537, N1997);
and AND2 (N2030, N2024, N1437);
xor XOR2 (N2031, N2022, N1498);
or OR4 (N2032, N2009, N898, N34, N1577);
xor XOR2 (N2033, N2016, N1127);
or OR2 (N2034, N2032, N1478);
or OR4 (N2035, N2029, N265, N77, N523);
and AND2 (N2036, N2028, N150);
xor XOR2 (N2037, N2036, N756);
and AND3 (N2038, N2033, N420, N468);
nor NOR3 (N2039, N2035, N20, N1173);
nor NOR4 (N2040, N2007, N2028, N376, N149);
not NOT1 (N2041, N2038);
buf BUF1 (N2042, N2041);
nor NOR2 (N2043, N2031, N67);
nand NAND2 (N2044, N2042, N217);
buf BUF1 (N2045, N2037);
xor XOR2 (N2046, N2021, N1432);
or OR3 (N2047, N2034, N1648, N368);
or OR2 (N2048, N2043, N1829);
nand NAND2 (N2049, N2047, N1836);
xor XOR2 (N2050, N2049, N598);
nand NAND2 (N2051, N2026, N648);
not NOT1 (N2052, N2048);
buf BUF1 (N2053, N2050);
and AND4 (N2054, N2052, N1093, N249, N163);
nor NOR3 (N2055, N2046, N52, N960);
nand NAND2 (N2056, N2051, N700);
nor NOR2 (N2057, N2056, N400);
and AND3 (N2058, N2054, N528, N1373);
nor NOR4 (N2059, N2012, N609, N1764, N64);
xor XOR2 (N2060, N2053, N630);
nor NOR3 (N2061, N2059, N860, N1275);
nor NOR4 (N2062, N2030, N259, N2000, N1600);
nand NAND3 (N2063, N2057, N696, N903);
not NOT1 (N2064, N2062);
or OR3 (N2065, N2058, N213, N437);
xor XOR2 (N2066, N2064, N1785);
nor NOR4 (N2067, N2063, N65, N1383, N1228);
nand NAND3 (N2068, N2060, N305, N1502);
nand NAND3 (N2069, N2068, N1800, N357);
xor XOR2 (N2070, N2069, N1716);
not NOT1 (N2071, N2039);
and AND2 (N2072, N2065, N743);
and AND4 (N2073, N2044, N617, N1144, N1878);
buf BUF1 (N2074, N2071);
not NOT1 (N2075, N2040);
not NOT1 (N2076, N2066);
xor XOR2 (N2077, N2070, N1508);
xor XOR2 (N2078, N2073, N1971);
nand NAND4 (N2079, N2055, N432, N1682, N754);
not NOT1 (N2080, N2074);
nor NOR3 (N2081, N2061, N455, N269);
nor NOR2 (N2082, N2045, N1888);
and AND4 (N2083, N2082, N1381, N1662, N1658);
buf BUF1 (N2084, N2080);
nand NAND3 (N2085, N2075, N913, N1219);
not NOT1 (N2086, N2085);
buf BUF1 (N2087, N2072);
nand NAND3 (N2088, N2087, N1394, N1604);
nand NAND4 (N2089, N2078, N1751, N1638, N1678);
or OR3 (N2090, N2067, N429, N1005);
buf BUF1 (N2091, N2084);
xor XOR2 (N2092, N2088, N1254);
or OR3 (N2093, N2077, N686, N1200);
buf BUF1 (N2094, N2079);
not NOT1 (N2095, N2094);
nand NAND4 (N2096, N2089, N746, N993, N1203);
buf BUF1 (N2097, N2081);
nand NAND3 (N2098, N2091, N1884, N1185);
and AND4 (N2099, N2076, N1798, N166, N1109);
nor NOR2 (N2100, N2095, N632);
nor NOR4 (N2101, N2092, N709, N889, N29);
buf BUF1 (N2102, N2096);
buf BUF1 (N2103, N2098);
not NOT1 (N2104, N2102);
and AND4 (N2105, N2083, N1270, N901, N1059);
nor NOR2 (N2106, N2099, N243);
xor XOR2 (N2107, N2086, N11);
buf BUF1 (N2108, N2105);
or OR3 (N2109, N2101, N873, N716);
xor XOR2 (N2110, N2097, N580);
not NOT1 (N2111, N2107);
and AND4 (N2112, N2104, N1016, N1366, N1601);
not NOT1 (N2113, N2103);
or OR3 (N2114, N2110, N622, N1715);
nor NOR2 (N2115, N2100, N1109);
buf BUF1 (N2116, N2115);
xor XOR2 (N2117, N2090, N1141);
not NOT1 (N2118, N2111);
nor NOR3 (N2119, N2112, N1733, N1993);
nand NAND2 (N2120, N2118, N1696);
buf BUF1 (N2121, N2114);
and AND2 (N2122, N2093, N1275);
buf BUF1 (N2123, N2116);
nor NOR4 (N2124, N2109, N439, N1501, N1959);
nor NOR3 (N2125, N2113, N1754, N1705);
buf BUF1 (N2126, N2121);
xor XOR2 (N2127, N2123, N2082);
nand NAND2 (N2128, N2126, N1703);
nor NOR3 (N2129, N2124, N1817, N2102);
nor NOR2 (N2130, N2129, N996);
buf BUF1 (N2131, N2125);
nand NAND2 (N2132, N2117, N1754);
nand NAND2 (N2133, N2108, N526);
or OR4 (N2134, N2106, N1001, N1642, N1300);
nand NAND2 (N2135, N2128, N1729);
xor XOR2 (N2136, N2122, N1399);
xor XOR2 (N2137, N2120, N1448);
and AND3 (N2138, N2135, N1668, N1022);
nand NAND2 (N2139, N2134, N1592);
buf BUF1 (N2140, N2127);
or OR3 (N2141, N2132, N270, N1);
nand NAND3 (N2142, N2139, N2076, N2073);
xor XOR2 (N2143, N2138, N664);
xor XOR2 (N2144, N2140, N957);
and AND2 (N2145, N2136, N271);
or OR2 (N2146, N2143, N121);
nor NOR2 (N2147, N2144, N386);
xor XOR2 (N2148, N2130, N1995);
or OR2 (N2149, N2146, N2139);
not NOT1 (N2150, N2141);
xor XOR2 (N2151, N2131, N985);
not NOT1 (N2152, N2133);
nor NOR3 (N2153, N2151, N714, N1202);
and AND4 (N2154, N2149, N227, N2097, N1810);
buf BUF1 (N2155, N2147);
and AND2 (N2156, N2119, N1325);
buf BUF1 (N2157, N2155);
buf BUF1 (N2158, N2156);
or OR4 (N2159, N2153, N516, N1551, N657);
nand NAND3 (N2160, N2159, N1145, N1004);
xor XOR2 (N2161, N2154, N581);
xor XOR2 (N2162, N2160, N543);
not NOT1 (N2163, N2161);
nand NAND2 (N2164, N2142, N2134);
xor XOR2 (N2165, N2145, N1971);
xor XOR2 (N2166, N2157, N152);
buf BUF1 (N2167, N2148);
and AND4 (N2168, N2165, N1695, N2123, N195);
nand NAND2 (N2169, N2167, N996);
and AND2 (N2170, N2158, N1113);
buf BUF1 (N2171, N2170);
nand NAND4 (N2172, N2171, N608, N37, N196);
buf BUF1 (N2173, N2168);
and AND2 (N2174, N2162, N1971);
nor NOR3 (N2175, N2166, N2054, N328);
and AND3 (N2176, N2164, N792, N1510);
nand NAND4 (N2177, N2175, N426, N1683, N149);
xor XOR2 (N2178, N2173, N1022);
buf BUF1 (N2179, N2152);
buf BUF1 (N2180, N2179);
nor NOR2 (N2181, N2176, N1680);
or OR2 (N2182, N2163, N1307);
or OR2 (N2183, N2174, N1793);
not NOT1 (N2184, N2180);
not NOT1 (N2185, N2183);
xor XOR2 (N2186, N2181, N1050);
buf BUF1 (N2187, N2169);
nor NOR3 (N2188, N2184, N928, N2106);
buf BUF1 (N2189, N2177);
or OR3 (N2190, N2188, N942, N2145);
and AND4 (N2191, N2137, N354, N709, N1034);
nand NAND4 (N2192, N2186, N1871, N1207, N2085);
or OR2 (N2193, N2178, N1736);
not NOT1 (N2194, N2190);
or OR4 (N2195, N2182, N484, N737, N431);
nand NAND4 (N2196, N2185, N2112, N671, N929);
nand NAND3 (N2197, N2194, N649, N840);
xor XOR2 (N2198, N2197, N918);
or OR4 (N2199, N2191, N1457, N2047, N1878);
buf BUF1 (N2200, N2198);
nor NOR4 (N2201, N2172, N1646, N908, N1188);
xor XOR2 (N2202, N2195, N2043);
and AND3 (N2203, N2189, N981, N638);
not NOT1 (N2204, N2199);
and AND3 (N2205, N2202, N1346, N1341);
and AND2 (N2206, N2187, N1544);
not NOT1 (N2207, N2204);
xor XOR2 (N2208, N2150, N1985);
xor XOR2 (N2209, N2196, N1517);
buf BUF1 (N2210, N2200);
or OR3 (N2211, N2203, N77, N899);
or OR2 (N2212, N2209, N1799);
nand NAND3 (N2213, N2193, N1704, N1721);
nor NOR2 (N2214, N2211, N944);
nor NOR3 (N2215, N2201, N962, N273);
or OR2 (N2216, N2207, N2007);
nor NOR3 (N2217, N2214, N2159, N1151);
nand NAND4 (N2218, N2210, N1335, N479, N361);
nand NAND2 (N2219, N2208, N1203);
and AND3 (N2220, N2205, N66, N2033);
xor XOR2 (N2221, N2192, N1748);
buf BUF1 (N2222, N2220);
nor NOR2 (N2223, N2218, N1089);
xor XOR2 (N2224, N2222, N701);
nand NAND4 (N2225, N2215, N850, N1763, N1734);
not NOT1 (N2226, N2213);
not NOT1 (N2227, N2221);
nand NAND4 (N2228, N2224, N1439, N1894, N221);
buf BUF1 (N2229, N2206);
and AND4 (N2230, N2225, N30, N135, N2028);
or OR2 (N2231, N2216, N677);
nor NOR3 (N2232, N2217, N59, N749);
nand NAND3 (N2233, N2219, N619, N732);
or OR3 (N2234, N2212, N1843, N1144);
not NOT1 (N2235, N2233);
buf BUF1 (N2236, N2231);
or OR3 (N2237, N2229, N376, N906);
xor XOR2 (N2238, N2223, N737);
nor NOR3 (N2239, N2236, N642, N972);
nor NOR3 (N2240, N2227, N1846, N1055);
or OR3 (N2241, N2232, N1872, N482);
not NOT1 (N2242, N2234);
xor XOR2 (N2243, N2235, N1728);
xor XOR2 (N2244, N2228, N1888);
not NOT1 (N2245, N2244);
and AND3 (N2246, N2238, N2164, N1030);
buf BUF1 (N2247, N2242);
nor NOR3 (N2248, N2246, N609, N2223);
not NOT1 (N2249, N2247);
xor XOR2 (N2250, N2243, N896);
or OR2 (N2251, N2226, N1724);
xor XOR2 (N2252, N2251, N839);
nor NOR2 (N2253, N2240, N91);
buf BUF1 (N2254, N2253);
buf BUF1 (N2255, N2241);
nor NOR2 (N2256, N2255, N1664);
nand NAND2 (N2257, N2239, N1142);
xor XOR2 (N2258, N2245, N2220);
buf BUF1 (N2259, N2230);
xor XOR2 (N2260, N2259, N1602);
xor XOR2 (N2261, N2252, N90);
not NOT1 (N2262, N2254);
or OR2 (N2263, N2261, N1275);
not NOT1 (N2264, N2260);
nor NOR2 (N2265, N2248, N1172);
not NOT1 (N2266, N2257);
nand NAND3 (N2267, N2264, N1347, N2033);
or OR2 (N2268, N2267, N1181);
buf BUF1 (N2269, N2262);
not NOT1 (N2270, N2256);
nor NOR2 (N2271, N2265, N272);
not NOT1 (N2272, N2250);
buf BUF1 (N2273, N2272);
buf BUF1 (N2274, N2270);
or OR4 (N2275, N2258, N1991, N1710, N960);
not NOT1 (N2276, N2268);
xor XOR2 (N2277, N2271, N2006);
nand NAND4 (N2278, N2266, N1175, N1320, N1337);
not NOT1 (N2279, N2269);
nand NAND3 (N2280, N2275, N2247, N2197);
not NOT1 (N2281, N2277);
buf BUF1 (N2282, N2281);
xor XOR2 (N2283, N2279, N1306);
xor XOR2 (N2284, N2263, N646);
or OR2 (N2285, N2278, N1335);
xor XOR2 (N2286, N2273, N504);
not NOT1 (N2287, N2283);
and AND3 (N2288, N2249, N201, N717);
buf BUF1 (N2289, N2284);
buf BUF1 (N2290, N2287);
nand NAND2 (N2291, N2274, N2139);
nand NAND2 (N2292, N2282, N1938);
not NOT1 (N2293, N2288);
nor NOR3 (N2294, N2289, N1878, N1536);
buf BUF1 (N2295, N2285);
not NOT1 (N2296, N2291);
nor NOR3 (N2297, N2292, N775, N601);
and AND3 (N2298, N2294, N1395, N796);
not NOT1 (N2299, N2280);
nor NOR4 (N2300, N2298, N492, N1783, N39);
not NOT1 (N2301, N2299);
and AND2 (N2302, N2296, N920);
nor NOR4 (N2303, N2286, N2290, N1869, N472);
or OR3 (N2304, N266, N1802, N1574);
not NOT1 (N2305, N2301);
nor NOR4 (N2306, N2304, N1277, N832, N1209);
buf BUF1 (N2307, N2300);
not NOT1 (N2308, N2302);
and AND3 (N2309, N2308, N559, N971);
or OR4 (N2310, N2276, N759, N945, N921);
not NOT1 (N2311, N2310);
not NOT1 (N2312, N2295);
and AND2 (N2313, N2303, N842);
xor XOR2 (N2314, N2313, N3);
nand NAND3 (N2315, N2293, N884, N877);
nand NAND2 (N2316, N2237, N2109);
not NOT1 (N2317, N2314);
not NOT1 (N2318, N2312);
nand NAND2 (N2319, N2315, N2157);
xor XOR2 (N2320, N2319, N1053);
nand NAND2 (N2321, N2318, N1349);
xor XOR2 (N2322, N2309, N2223);
buf BUF1 (N2323, N2306);
nand NAND3 (N2324, N2321, N2087, N1513);
buf BUF1 (N2325, N2311);
and AND4 (N2326, N2320, N813, N1674, N14);
and AND4 (N2327, N2297, N2144, N1884, N573);
nor NOR2 (N2328, N2327, N1075);
nor NOR2 (N2329, N2307, N400);
and AND4 (N2330, N2305, N1330, N2228, N1858);
or OR3 (N2331, N2329, N1868, N1214);
nor NOR4 (N2332, N2324, N1068, N1184, N318);
nor NOR2 (N2333, N2331, N1518);
nand NAND2 (N2334, N2332, N311);
nor NOR2 (N2335, N2325, N1785);
and AND4 (N2336, N2334, N2107, N2005, N272);
or OR4 (N2337, N2336, N55, N1740, N1518);
not NOT1 (N2338, N2322);
or OR2 (N2339, N2328, N528);
nor NOR2 (N2340, N2337, N329);
or OR2 (N2341, N2339, N1615);
xor XOR2 (N2342, N2330, N1396);
nand NAND4 (N2343, N2316, N2265, N1821, N2015);
not NOT1 (N2344, N2335);
nor NOR4 (N2345, N2338, N85, N1702, N1052);
or OR4 (N2346, N2317, N1735, N1259, N38);
nand NAND3 (N2347, N2346, N1541, N1933);
buf BUF1 (N2348, N2340);
not NOT1 (N2349, N2348);
buf BUF1 (N2350, N2347);
or OR4 (N2351, N2349, N17, N1076, N467);
or OR3 (N2352, N2333, N1850, N462);
xor XOR2 (N2353, N2345, N2100);
nand NAND2 (N2354, N2352, N550);
not NOT1 (N2355, N2350);
nand NAND2 (N2356, N2343, N1074);
not NOT1 (N2357, N2351);
nor NOR2 (N2358, N2344, N1203);
not NOT1 (N2359, N2341);
not NOT1 (N2360, N2358);
nor NOR3 (N2361, N2356, N1435, N844);
or OR3 (N2362, N2323, N2068, N598);
not NOT1 (N2363, N2359);
xor XOR2 (N2364, N2342, N2332);
not NOT1 (N2365, N2353);
or OR3 (N2366, N2363, N1947, N62);
buf BUF1 (N2367, N2357);
buf BUF1 (N2368, N2355);
buf BUF1 (N2369, N2354);
xor XOR2 (N2370, N2360, N1263);
not NOT1 (N2371, N2364);
nor NOR3 (N2372, N2365, N170, N1290);
nor NOR2 (N2373, N2370, N1098);
buf BUF1 (N2374, N2366);
xor XOR2 (N2375, N2368, N145);
and AND2 (N2376, N2372, N1660);
nand NAND2 (N2377, N2371, N1157);
and AND2 (N2378, N2367, N1882);
nor NOR2 (N2379, N2377, N278);
or OR3 (N2380, N2369, N525, N1389);
or OR2 (N2381, N2373, N1619);
nor NOR3 (N2382, N2326, N1303, N302);
not NOT1 (N2383, N2380);
or OR2 (N2384, N2381, N2318);
buf BUF1 (N2385, N2375);
buf BUF1 (N2386, N2374);
nor NOR4 (N2387, N2361, N69, N1786, N611);
not NOT1 (N2388, N2386);
and AND3 (N2389, N2383, N730, N1039);
not NOT1 (N2390, N2376);
xor XOR2 (N2391, N2387, N1930);
nor NOR2 (N2392, N2388, N964);
nand NAND2 (N2393, N2392, N554);
or OR3 (N2394, N2389, N1715, N49);
nand NAND4 (N2395, N2378, N919, N2246, N38);
not NOT1 (N2396, N2385);
and AND3 (N2397, N2396, N698, N2064);
nand NAND2 (N2398, N2393, N1917);
or OR2 (N2399, N2398, N507);
buf BUF1 (N2400, N2362);
and AND3 (N2401, N2395, N1984, N447);
or OR3 (N2402, N2394, N2005, N1788);
nor NOR4 (N2403, N2402, N996, N1412, N439);
xor XOR2 (N2404, N2391, N1764);
buf BUF1 (N2405, N2403);
nand NAND3 (N2406, N2379, N775, N1093);
not NOT1 (N2407, N2405);
not NOT1 (N2408, N2407);
not NOT1 (N2409, N2406);
not NOT1 (N2410, N2390);
buf BUF1 (N2411, N2409);
xor XOR2 (N2412, N2382, N247);
buf BUF1 (N2413, N2397);
nand NAND2 (N2414, N2410, N1629);
nor NOR2 (N2415, N2412, N2207);
xor XOR2 (N2416, N2411, N2239);
and AND4 (N2417, N2404, N178, N1125, N268);
xor XOR2 (N2418, N2413, N766);
or OR2 (N2419, N2399, N286);
nor NOR2 (N2420, N2384, N278);
xor XOR2 (N2421, N2408, N2375);
nor NOR3 (N2422, N2420, N1774, N1011);
or OR2 (N2423, N2417, N425);
not NOT1 (N2424, N2414);
or OR2 (N2425, N2422, N852);
and AND2 (N2426, N2419, N1044);
and AND4 (N2427, N2425, N1431, N247, N142);
and AND3 (N2428, N2423, N389, N1536);
not NOT1 (N2429, N2400);
xor XOR2 (N2430, N2416, N348);
nand NAND3 (N2431, N2427, N593, N1894);
nand NAND2 (N2432, N2418, N2376);
nand NAND3 (N2433, N2421, N2368, N2266);
nand NAND4 (N2434, N2432, N485, N2073, N807);
and AND4 (N2435, N2426, N34, N2096, N147);
or OR2 (N2436, N2435, N328);
and AND2 (N2437, N2429, N1375);
buf BUF1 (N2438, N2437);
nand NAND2 (N2439, N2431, N1473);
nand NAND3 (N2440, N2434, N1063, N1828);
nand NAND4 (N2441, N2415, N924, N443, N131);
and AND3 (N2442, N2439, N234, N148);
not NOT1 (N2443, N2442);
nand NAND3 (N2444, N2436, N2157, N2161);
or OR3 (N2445, N2441, N534, N1356);
not NOT1 (N2446, N2443);
nor NOR4 (N2447, N2428, N1341, N1388, N53);
buf BUF1 (N2448, N2447);
xor XOR2 (N2449, N2448, N2238);
xor XOR2 (N2450, N2401, N13);
and AND3 (N2451, N2449, N889, N1501);
not NOT1 (N2452, N2451);
xor XOR2 (N2453, N2445, N2305);
or OR4 (N2454, N2452, N1066, N906, N1532);
nor NOR3 (N2455, N2453, N1637, N1933);
or OR4 (N2456, N2450, N1810, N2383, N723);
xor XOR2 (N2457, N2440, N1687);
xor XOR2 (N2458, N2424, N1921);
and AND4 (N2459, N2433, N1574, N1772, N529);
and AND2 (N2460, N2438, N1088);
and AND3 (N2461, N2455, N1698, N28);
buf BUF1 (N2462, N2459);
nand NAND3 (N2463, N2456, N1621, N1337);
xor XOR2 (N2464, N2458, N301);
and AND4 (N2465, N2462, N1691, N219, N345);
or OR3 (N2466, N2463, N613, N2462);
not NOT1 (N2467, N2460);
and AND3 (N2468, N2446, N1036, N687);
xor XOR2 (N2469, N2444, N2183);
and AND4 (N2470, N2465, N2350, N1255, N1116);
or OR4 (N2471, N2467, N1578, N1871, N2302);
nor NOR4 (N2472, N2430, N1059, N1961, N1547);
nand NAND2 (N2473, N2472, N832);
and AND4 (N2474, N2461, N1427, N542, N1525);
buf BUF1 (N2475, N2454);
xor XOR2 (N2476, N2474, N2457);
nand NAND4 (N2477, N2178, N613, N1171, N113);
not NOT1 (N2478, N2476);
and AND3 (N2479, N2469, N1219, N2023);
nand NAND3 (N2480, N2473, N1168, N1715);
and AND2 (N2481, N2466, N2082);
and AND3 (N2482, N2478, N21, N1273);
nor NOR2 (N2483, N2477, N776);
or OR4 (N2484, N2468, N1117, N1952, N1166);
not NOT1 (N2485, N2479);
nand NAND4 (N2486, N2484, N1344, N1374, N208);
and AND3 (N2487, N2480, N1525, N1352);
xor XOR2 (N2488, N2487, N1144);
nor NOR4 (N2489, N2486, N1195, N1401, N209);
or OR4 (N2490, N2475, N209, N643, N2320);
or OR4 (N2491, N2490, N2458, N1210, N1118);
and AND4 (N2492, N2491, N2263, N2452, N843);
buf BUF1 (N2493, N2489);
and AND3 (N2494, N2471, N1988, N2325);
buf BUF1 (N2495, N2493);
nor NOR4 (N2496, N2483, N2369, N2177, N345);
and AND4 (N2497, N2481, N1244, N1529, N1552);
xor XOR2 (N2498, N2495, N1823);
nand NAND4 (N2499, N2498, N2113, N1954, N1356);
or OR3 (N2500, N2488, N1066, N170);
xor XOR2 (N2501, N2499, N1615);
and AND3 (N2502, N2492, N1094, N468);
not NOT1 (N2503, N2501);
not NOT1 (N2504, N2503);
xor XOR2 (N2505, N2464, N840);
xor XOR2 (N2506, N2485, N1407);
buf BUF1 (N2507, N2470);
not NOT1 (N2508, N2504);
nor NOR4 (N2509, N2494, N666, N1102, N12);
buf BUF1 (N2510, N2505);
nand NAND2 (N2511, N2509, N348);
xor XOR2 (N2512, N2500, N506);
and AND3 (N2513, N2497, N1969, N1425);
nor NOR4 (N2514, N2511, N2083, N1065, N1059);
nand NAND4 (N2515, N2508, N1946, N231, N1911);
not NOT1 (N2516, N2502);
and AND2 (N2517, N2507, N715);
buf BUF1 (N2518, N2496);
nand NAND3 (N2519, N2482, N424, N293);
buf BUF1 (N2520, N2506);
nor NOR3 (N2521, N2512, N370, N622);
xor XOR2 (N2522, N2516, N19);
nor NOR3 (N2523, N2515, N1231, N2182);
nand NAND2 (N2524, N2521, N2268);
or OR2 (N2525, N2520, N360);
or OR2 (N2526, N2513, N517);
buf BUF1 (N2527, N2524);
nand NAND3 (N2528, N2514, N1222, N1919);
xor XOR2 (N2529, N2526, N454);
not NOT1 (N2530, N2523);
xor XOR2 (N2531, N2529, N648);
xor XOR2 (N2532, N2517, N1062);
or OR2 (N2533, N2532, N999);
or OR4 (N2534, N2528, N572, N1877, N2085);
buf BUF1 (N2535, N2518);
or OR4 (N2536, N2525, N1375, N1442, N1556);
nand NAND4 (N2537, N2536, N309, N2295, N408);
not NOT1 (N2538, N2530);
xor XOR2 (N2539, N2534, N1394);
not NOT1 (N2540, N2538);
nand NAND2 (N2541, N2510, N1093);
and AND3 (N2542, N2519, N1480, N1496);
not NOT1 (N2543, N2539);
nor NOR3 (N2544, N2531, N1886, N1571);
nand NAND3 (N2545, N2543, N2289, N1147);
not NOT1 (N2546, N2522);
and AND3 (N2547, N2535, N1124, N836);
and AND3 (N2548, N2533, N1218, N55);
nand NAND2 (N2549, N2527, N1230);
nor NOR3 (N2550, N2537, N1693, N2074);
and AND4 (N2551, N2544, N301, N1311, N1319);
xor XOR2 (N2552, N2547, N801);
and AND2 (N2553, N2545, N887);
or OR2 (N2554, N2541, N401);
nand NAND4 (N2555, N2550, N891, N188, N311);
buf BUF1 (N2556, N2552);
nor NOR3 (N2557, N2546, N1732, N880);
nor NOR3 (N2558, N2549, N916, N2115);
and AND3 (N2559, N2548, N841, N1557);
nor NOR3 (N2560, N2540, N2416, N1283);
or OR3 (N2561, N2551, N998, N526);
xor XOR2 (N2562, N2555, N2158);
nor NOR4 (N2563, N2558, N156, N983, N718);
not NOT1 (N2564, N2556);
or OR4 (N2565, N2560, N1168, N2335, N168);
and AND3 (N2566, N2563, N2054, N27);
or OR2 (N2567, N2557, N196);
nand NAND2 (N2568, N2567, N1394);
xor XOR2 (N2569, N2542, N1643);
nor NOR2 (N2570, N2568, N988);
nor NOR2 (N2571, N2569, N1928);
nand NAND3 (N2572, N2559, N2289, N1239);
not NOT1 (N2573, N2565);
buf BUF1 (N2574, N2562);
not NOT1 (N2575, N2564);
and AND2 (N2576, N2561, N984);
buf BUF1 (N2577, N2566);
not NOT1 (N2578, N2573);
buf BUF1 (N2579, N2576);
xor XOR2 (N2580, N2578, N178);
and AND2 (N2581, N2575, N839);
xor XOR2 (N2582, N2574, N1393);
xor XOR2 (N2583, N2572, N122);
or OR3 (N2584, N2582, N2424, N2578);
and AND4 (N2585, N2577, N1980, N1282, N377);
or OR2 (N2586, N2580, N221);
nor NOR4 (N2587, N2584, N2060, N1833, N220);
and AND3 (N2588, N2570, N832, N562);
buf BUF1 (N2589, N2588);
xor XOR2 (N2590, N2589, N2419);
and AND2 (N2591, N2586, N1678);
buf BUF1 (N2592, N2591);
nor NOR2 (N2593, N2579, N455);
xor XOR2 (N2594, N2590, N1089);
nand NAND4 (N2595, N2593, N353, N2259, N1408);
buf BUF1 (N2596, N2554);
not NOT1 (N2597, N2592);
not NOT1 (N2598, N2587);
xor XOR2 (N2599, N2597, N2520);
nor NOR4 (N2600, N2599, N269, N534, N1113);
nor NOR4 (N2601, N2571, N37, N1067, N2330);
nand NAND4 (N2602, N2598, N1751, N1806, N1359);
xor XOR2 (N2603, N2601, N336);
or OR3 (N2604, N2600, N593, N151);
nor NOR4 (N2605, N2596, N353, N1701, N1405);
xor XOR2 (N2606, N2581, N982);
buf BUF1 (N2607, N2583);
nand NAND4 (N2608, N2585, N1221, N1773, N295);
xor XOR2 (N2609, N2607, N1430);
nor NOR4 (N2610, N2553, N2233, N156, N1295);
and AND2 (N2611, N2606, N929);
or OR2 (N2612, N2604, N2028);
and AND4 (N2613, N2609, N511, N2170, N1488);
xor XOR2 (N2614, N2610, N969);
nand NAND3 (N2615, N2603, N1207, N82);
nor NOR3 (N2616, N2611, N1444, N359);
and AND4 (N2617, N2595, N630, N1789, N192);
or OR3 (N2618, N2617, N27, N2043);
not NOT1 (N2619, N2608);
or OR3 (N2620, N2614, N1369, N1869);
buf BUF1 (N2621, N2619);
and AND4 (N2622, N2605, N1045, N912, N2137);
nor NOR3 (N2623, N2594, N2145, N1311);
not NOT1 (N2624, N2616);
not NOT1 (N2625, N2613);
nand NAND2 (N2626, N2615, N1733);
xor XOR2 (N2627, N2623, N2458);
nand NAND4 (N2628, N2621, N1178, N1876, N1782);
not NOT1 (N2629, N2624);
or OR4 (N2630, N2626, N617, N696, N868);
or OR3 (N2631, N2630, N2567, N2161);
not NOT1 (N2632, N2631);
nor NOR2 (N2633, N2622, N645);
xor XOR2 (N2634, N2628, N2226);
or OR2 (N2635, N2629, N519);
or OR3 (N2636, N2634, N1681, N2635);
not NOT1 (N2637, N852);
not NOT1 (N2638, N2627);
nor NOR2 (N2639, N2633, N2581);
xor XOR2 (N2640, N2620, N870);
buf BUF1 (N2641, N2638);
not NOT1 (N2642, N2641);
nand NAND4 (N2643, N2637, N2604, N1705, N2258);
xor XOR2 (N2644, N2639, N2127);
nor NOR4 (N2645, N2644, N110, N1823, N2500);
nand NAND2 (N2646, N2625, N1899);
nor NOR3 (N2647, N2640, N1058, N735);
nand NAND2 (N2648, N2647, N1719);
nand NAND2 (N2649, N2646, N45);
nand NAND2 (N2650, N2645, N1380);
not NOT1 (N2651, N2618);
or OR2 (N2652, N2642, N1849);
nor NOR2 (N2653, N2651, N450);
or OR2 (N2654, N2636, N2327);
xor XOR2 (N2655, N2649, N2591);
and AND4 (N2656, N2652, N2456, N1811, N1425);
not NOT1 (N2657, N2602);
or OR4 (N2658, N2653, N366, N168, N804);
buf BUF1 (N2659, N2655);
xor XOR2 (N2660, N2612, N839);
and AND3 (N2661, N2632, N2558, N1111);
buf BUF1 (N2662, N2660);
nor NOR3 (N2663, N2662, N349, N748);
nor NOR3 (N2664, N2654, N2447, N475);
nor NOR4 (N2665, N2656, N1736, N2433, N2569);
nand NAND4 (N2666, N2661, N1196, N1630, N10);
nor NOR2 (N2667, N2663, N2209);
nand NAND2 (N2668, N2664, N854);
nand NAND3 (N2669, N2650, N178, N2184);
nor NOR2 (N2670, N2643, N705);
and AND4 (N2671, N2667, N306, N1219, N1904);
or OR3 (N2672, N2666, N2558, N478);
xor XOR2 (N2673, N2665, N448);
not NOT1 (N2674, N2669);
buf BUF1 (N2675, N2648);
and AND2 (N2676, N2674, N2614);
not NOT1 (N2677, N2676);
buf BUF1 (N2678, N2675);
not NOT1 (N2679, N2671);
buf BUF1 (N2680, N2672);
nand NAND3 (N2681, N2680, N2023, N657);
nor NOR3 (N2682, N2679, N2502, N2319);
not NOT1 (N2683, N2657);
nand NAND3 (N2684, N2677, N1517, N64);
or OR4 (N2685, N2658, N1786, N1555, N1992);
nor NOR3 (N2686, N2670, N1394, N2088);
nor NOR4 (N2687, N2684, N794, N1643, N1153);
buf BUF1 (N2688, N2687);
nor NOR4 (N2689, N2678, N1183, N43, N51);
not NOT1 (N2690, N2683);
not NOT1 (N2691, N2659);
nor NOR4 (N2692, N2685, N1026, N520, N986);
nor NOR4 (N2693, N2673, N174, N1538, N174);
nand NAND2 (N2694, N2689, N827);
not NOT1 (N2695, N2668);
buf BUF1 (N2696, N2694);
buf BUF1 (N2697, N2682);
xor XOR2 (N2698, N2696, N902);
buf BUF1 (N2699, N2693);
buf BUF1 (N2700, N2688);
nand NAND2 (N2701, N2681, N653);
nand NAND3 (N2702, N2695, N1336, N2177);
not NOT1 (N2703, N2692);
and AND4 (N2704, N2702, N2327, N1015, N2137);
and AND4 (N2705, N2697, N1526, N1441, N774);
nor NOR4 (N2706, N2700, N2616, N592, N1385);
xor XOR2 (N2707, N2686, N157);
xor XOR2 (N2708, N2706, N1053);
buf BUF1 (N2709, N2703);
or OR2 (N2710, N2707, N1474);
not NOT1 (N2711, N2705);
not NOT1 (N2712, N2701);
nand NAND3 (N2713, N2709, N1694, N1871);
or OR3 (N2714, N2708, N1625, N1856);
and AND2 (N2715, N2711, N1200);
not NOT1 (N2716, N2710);
and AND2 (N2717, N2714, N235);
or OR2 (N2718, N2716, N226);
nand NAND2 (N2719, N2691, N1452);
xor XOR2 (N2720, N2699, N2050);
and AND4 (N2721, N2704, N1321, N313, N2586);
not NOT1 (N2722, N2712);
not NOT1 (N2723, N2690);
or OR4 (N2724, N2698, N1770, N453, N1207);
nor NOR3 (N2725, N2713, N1075, N1938);
nand NAND3 (N2726, N2717, N2509, N1042);
nand NAND3 (N2727, N2724, N419, N1210);
and AND3 (N2728, N2719, N620, N237);
or OR3 (N2729, N2715, N2483, N2728);
nor NOR4 (N2730, N168, N1800, N1220, N1901);
nor NOR3 (N2731, N2720, N71, N1194);
not NOT1 (N2732, N2723);
nor NOR2 (N2733, N2727, N2060);
nor NOR3 (N2734, N2729, N1828, N303);
not NOT1 (N2735, N2722);
nor NOR4 (N2736, N2735, N2118, N1574, N2639);
or OR4 (N2737, N2730, N1164, N592, N205);
xor XOR2 (N2738, N2718, N1832);
and AND4 (N2739, N2737, N156, N1325, N1476);
nor NOR4 (N2740, N2721, N2622, N809, N2271);
nand NAND3 (N2741, N2739, N320, N2172);
nor NOR3 (N2742, N2733, N2485, N1359);
nand NAND2 (N2743, N2726, N519);
buf BUF1 (N2744, N2742);
buf BUF1 (N2745, N2731);
xor XOR2 (N2746, N2745, N121);
and AND2 (N2747, N2738, N597);
or OR4 (N2748, N2734, N2378, N713, N1910);
or OR2 (N2749, N2732, N2020);
xor XOR2 (N2750, N2743, N1677);
nand NAND4 (N2751, N2748, N2439, N1236, N1196);
nor NOR2 (N2752, N2749, N2478);
xor XOR2 (N2753, N2746, N2127);
not NOT1 (N2754, N2753);
and AND3 (N2755, N2750, N2381, N1265);
nor NOR4 (N2756, N2751, N2145, N884, N2522);
or OR4 (N2757, N2755, N110, N1362, N1636);
and AND3 (N2758, N2741, N2502, N1205);
or OR4 (N2759, N2740, N2371, N1971, N1906);
and AND4 (N2760, N2757, N2547, N2355, N825);
or OR2 (N2761, N2754, N1731);
buf BUF1 (N2762, N2760);
nand NAND4 (N2763, N2756, N1679, N409, N2352);
not NOT1 (N2764, N2761);
or OR3 (N2765, N2744, N140, N2568);
xor XOR2 (N2766, N2725, N1662);
not NOT1 (N2767, N2766);
xor XOR2 (N2768, N2747, N329);
not NOT1 (N2769, N2758);
nand NAND3 (N2770, N2762, N761, N111);
xor XOR2 (N2771, N2769, N1028);
or OR4 (N2772, N2763, N1799, N821, N945);
buf BUF1 (N2773, N2770);
nand NAND3 (N2774, N2764, N2727, N124);
nor NOR4 (N2775, N2759, N497, N2621, N2101);
buf BUF1 (N2776, N2773);
and AND3 (N2777, N2765, N244, N1258);
buf BUF1 (N2778, N2752);
not NOT1 (N2779, N2736);
xor XOR2 (N2780, N2774, N915);
not NOT1 (N2781, N2780);
nor NOR4 (N2782, N2768, N542, N1352, N1343);
buf BUF1 (N2783, N2781);
xor XOR2 (N2784, N2772, N1150);
nor NOR2 (N2785, N2782, N66);
or OR2 (N2786, N2767, N2732);
nand NAND2 (N2787, N2776, N2533);
and AND2 (N2788, N2785, N492);
or OR3 (N2789, N2787, N2242, N1662);
and AND2 (N2790, N2778, N1696);
or OR2 (N2791, N2786, N2565);
buf BUF1 (N2792, N2777);
buf BUF1 (N2793, N2788);
and AND4 (N2794, N2775, N868, N1247, N1589);
or OR4 (N2795, N2790, N2057, N2355, N706);
nor NOR3 (N2796, N2789, N2525, N1073);
nor NOR2 (N2797, N2795, N1413);
or OR2 (N2798, N2794, N2415);
not NOT1 (N2799, N2796);
xor XOR2 (N2800, N2799, N1135);
not NOT1 (N2801, N2779);
nor NOR2 (N2802, N2801, N856);
not NOT1 (N2803, N2784);
nand NAND4 (N2804, N2792, N279, N1204, N231);
nor NOR2 (N2805, N2804, N1648);
or OR3 (N2806, N2791, N840, N2381);
and AND2 (N2807, N2803, N1789);
and AND2 (N2808, N2797, N987);
xor XOR2 (N2809, N2802, N1834);
nand NAND4 (N2810, N2783, N995, N1166, N54);
buf BUF1 (N2811, N2800);
nand NAND2 (N2812, N2793, N1832);
xor XOR2 (N2813, N2812, N2787);
and AND3 (N2814, N2808, N1876, N387);
nand NAND3 (N2815, N2805, N582, N1642);
and AND4 (N2816, N2813, N1058, N66, N2152);
nor NOR2 (N2817, N2809, N910);
nor NOR3 (N2818, N2798, N2232, N2060);
and AND2 (N2819, N2771, N2122);
xor XOR2 (N2820, N2807, N56);
buf BUF1 (N2821, N2814);
not NOT1 (N2822, N2810);
nand NAND3 (N2823, N2816, N968, N2049);
or OR4 (N2824, N2823, N2405, N794, N2257);
nand NAND4 (N2825, N2820, N1760, N2361, N2565);
xor XOR2 (N2826, N2811, N1162);
nor NOR3 (N2827, N2825, N982, N1299);
or OR4 (N2828, N2817, N1084, N771, N2008);
buf BUF1 (N2829, N2822);
and AND4 (N2830, N2821, N1465, N1100, N1692);
nor NOR3 (N2831, N2830, N2699, N1226);
xor XOR2 (N2832, N2824, N728);
and AND4 (N2833, N2832, N1438, N2376, N2216);
buf BUF1 (N2834, N2829);
not NOT1 (N2835, N2828);
nor NOR3 (N2836, N2819, N358, N504);
not NOT1 (N2837, N2831);
nand NAND3 (N2838, N2836, N2402, N1570);
or OR4 (N2839, N2838, N662, N1532, N468);
xor XOR2 (N2840, N2827, N1388);
buf BUF1 (N2841, N2818);
and AND3 (N2842, N2841, N640, N638);
not NOT1 (N2843, N2837);
xor XOR2 (N2844, N2806, N602);
and AND3 (N2845, N2843, N1787, N2113);
nand NAND3 (N2846, N2844, N2213, N374);
not NOT1 (N2847, N2815);
or OR4 (N2848, N2833, N1573, N1548, N1092);
or OR3 (N2849, N2847, N1884, N358);
not NOT1 (N2850, N2835);
nand NAND2 (N2851, N2850, N290);
xor XOR2 (N2852, N2826, N1810);
nor NOR4 (N2853, N2845, N929, N2300, N359);
or OR4 (N2854, N2834, N247, N2752, N969);
not NOT1 (N2855, N2849);
and AND2 (N2856, N2848, N234);
nor NOR2 (N2857, N2852, N1391);
xor XOR2 (N2858, N2842, N243);
xor XOR2 (N2859, N2851, N2318);
not NOT1 (N2860, N2858);
xor XOR2 (N2861, N2840, N1768);
xor XOR2 (N2862, N2856, N1464);
nand NAND2 (N2863, N2846, N39);
nand NAND4 (N2864, N2853, N2252, N1860, N1961);
nor NOR2 (N2865, N2863, N366);
buf BUF1 (N2866, N2864);
buf BUF1 (N2867, N2855);
xor XOR2 (N2868, N2839, N960);
buf BUF1 (N2869, N2860);
xor XOR2 (N2870, N2867, N1238);
nor NOR4 (N2871, N2859, N1875, N1138, N2412);
and AND2 (N2872, N2861, N2538);
nor NOR4 (N2873, N2857, N2523, N2583, N90);
nor NOR4 (N2874, N2873, N2854, N1722, N1453);
nor NOR3 (N2875, N439, N1335, N1165);
xor XOR2 (N2876, N2865, N460);
nor NOR4 (N2877, N2871, N2150, N2786, N359);
and AND2 (N2878, N2875, N374);
nor NOR4 (N2879, N2869, N1812, N1291, N2767);
and AND2 (N2880, N2862, N2130);
or OR4 (N2881, N2880, N2042, N164, N2744);
and AND2 (N2882, N2876, N983);
and AND3 (N2883, N2882, N1363, N1045);
buf BUF1 (N2884, N2874);
or OR4 (N2885, N2866, N1452, N748, N1700);
not NOT1 (N2886, N2883);
nor NOR4 (N2887, N2884, N929, N1065, N451);
or OR2 (N2888, N2885, N488);
nor NOR4 (N2889, N2868, N487, N123, N2833);
xor XOR2 (N2890, N2887, N2240);
not NOT1 (N2891, N2886);
or OR4 (N2892, N2872, N615, N2626, N1996);
nand NAND3 (N2893, N2870, N1016, N2761);
xor XOR2 (N2894, N2891, N2341);
not NOT1 (N2895, N2879);
not NOT1 (N2896, N2878);
buf BUF1 (N2897, N2894);
nor NOR3 (N2898, N2881, N1467, N1983);
buf BUF1 (N2899, N2898);
xor XOR2 (N2900, N2899, N70);
nor NOR3 (N2901, N2897, N2710, N315);
and AND2 (N2902, N2896, N911);
nor NOR2 (N2903, N2901, N749);
and AND2 (N2904, N2890, N155);
buf BUF1 (N2905, N2893);
nand NAND4 (N2906, N2895, N2877, N523, N1088);
buf BUF1 (N2907, N404);
and AND4 (N2908, N2902, N1873, N2501, N465);
nand NAND3 (N2909, N2889, N844, N1662);
nor NOR3 (N2910, N2904, N2629, N1325);
buf BUF1 (N2911, N2888);
nand NAND2 (N2912, N2900, N2494);
not NOT1 (N2913, N2905);
not NOT1 (N2914, N2910);
buf BUF1 (N2915, N2914);
buf BUF1 (N2916, N2907);
nor NOR2 (N2917, N2916, N2181);
and AND3 (N2918, N2917, N73, N550);
and AND2 (N2919, N2909, N2331);
or OR2 (N2920, N2911, N2611);
buf BUF1 (N2921, N2915);
nand NAND3 (N2922, N2913, N1424, N1609);
nand NAND3 (N2923, N2912, N1713, N251);
or OR2 (N2924, N2908, N631);
and AND3 (N2925, N2920, N1995, N473);
nor NOR4 (N2926, N2906, N711, N734, N765);
xor XOR2 (N2927, N2919, N2214);
nand NAND4 (N2928, N2903, N240, N1890, N219);
or OR3 (N2929, N2923, N2304, N2664);
nand NAND2 (N2930, N2918, N1116);
and AND3 (N2931, N2930, N2574, N2178);
nand NAND2 (N2932, N2892, N1010);
nor NOR2 (N2933, N2928, N2593);
xor XOR2 (N2934, N2933, N2819);
or OR4 (N2935, N2934, N1309, N2846, N574);
buf BUF1 (N2936, N2927);
buf BUF1 (N2937, N2926);
nor NOR4 (N2938, N2929, N120, N2337, N1454);
buf BUF1 (N2939, N2932);
xor XOR2 (N2940, N2921, N364);
or OR4 (N2941, N2931, N2784, N2730, N2526);
nand NAND2 (N2942, N2925, N2593);
xor XOR2 (N2943, N2938, N2587);
nor NOR4 (N2944, N2922, N1333, N813, N784);
and AND3 (N2945, N2944, N322, N563);
or OR3 (N2946, N2924, N742, N1553);
or OR2 (N2947, N2935, N749);
not NOT1 (N2948, N2945);
nand NAND3 (N2949, N2946, N1330, N2703);
nand NAND2 (N2950, N2936, N2858);
and AND4 (N2951, N2949, N1045, N188, N2262);
nor NOR4 (N2952, N2950, N1777, N2226, N2821);
nand NAND2 (N2953, N2939, N105);
buf BUF1 (N2954, N2947);
nand NAND2 (N2955, N2941, N1977);
or OR2 (N2956, N2948, N1274);
not NOT1 (N2957, N2937);
nand NAND2 (N2958, N2953, N245);
nand NAND4 (N2959, N2958, N234, N512, N2737);
not NOT1 (N2960, N2959);
nor NOR4 (N2961, N2943, N1818, N402, N1950);
and AND3 (N2962, N2961, N754, N1541);
nor NOR3 (N2963, N2942, N1678, N10);
nor NOR3 (N2964, N2962, N1263, N960);
nor NOR3 (N2965, N2955, N1966, N1583);
not NOT1 (N2966, N2951);
not NOT1 (N2967, N2956);
not NOT1 (N2968, N2966);
nand NAND2 (N2969, N2952, N589);
nand NAND3 (N2970, N2967, N2060, N2489);
or OR4 (N2971, N2957, N2911, N628, N2780);
nand NAND3 (N2972, N2963, N1518, N1674);
nand NAND2 (N2973, N2970, N1659);
nor NOR3 (N2974, N2969, N713, N2336);
and AND3 (N2975, N2968, N1278, N2874);
or OR4 (N2976, N2960, N667, N2544, N583);
and AND2 (N2977, N2972, N1007);
not NOT1 (N2978, N2940);
or OR3 (N2979, N2973, N1631, N927);
buf BUF1 (N2980, N2965);
and AND2 (N2981, N2977, N2225);
nor NOR3 (N2982, N2974, N2970, N2363);
nor NOR4 (N2983, N2971, N997, N2274, N2312);
nor NOR2 (N2984, N2981, N2611);
nor NOR4 (N2985, N2954, N2014, N1038, N1065);
and AND4 (N2986, N2979, N847, N1709, N1959);
nor NOR3 (N2987, N2980, N2880, N1555);
and AND2 (N2988, N2986, N1358);
not NOT1 (N2989, N2983);
nor NOR2 (N2990, N2976, N2979);
buf BUF1 (N2991, N2988);
nand NAND2 (N2992, N2987, N113);
and AND2 (N2993, N2978, N2158);
xor XOR2 (N2994, N2992, N1581);
nand NAND2 (N2995, N2990, N2879);
buf BUF1 (N2996, N2985);
and AND2 (N2997, N2991, N1339);
and AND3 (N2998, N2984, N1541, N5);
or OR4 (N2999, N2996, N2713, N2654, N2534);
not NOT1 (N3000, N2997);
nand NAND3 (N3001, N2994, N506, N2527);
nor NOR3 (N3002, N2982, N1416, N2048);
buf BUF1 (N3003, N3002);
nor NOR2 (N3004, N2995, N1910);
not NOT1 (N3005, N3001);
nor NOR4 (N3006, N2989, N1561, N619, N2494);
or OR3 (N3007, N3003, N2071, N1781);
or OR4 (N3008, N2999, N2137, N1800, N1010);
or OR2 (N3009, N3007, N1851);
nor NOR2 (N3010, N2998, N2964);
or OR4 (N3011, N2454, N1929, N2550, N1918);
and AND2 (N3012, N3000, N1783);
and AND4 (N3013, N3006, N2261, N278, N2151);
nand NAND3 (N3014, N3005, N1384, N2192);
buf BUF1 (N3015, N3014);
not NOT1 (N3016, N3010);
not NOT1 (N3017, N3016);
nor NOR3 (N3018, N2993, N2469, N435);
nand NAND4 (N3019, N3011, N262, N979, N1589);
xor XOR2 (N3020, N3013, N1345);
xor XOR2 (N3021, N3009, N416);
buf BUF1 (N3022, N3021);
xor XOR2 (N3023, N3022, N2903);
xor XOR2 (N3024, N3017, N2315);
and AND2 (N3025, N3020, N1512);
nor NOR3 (N3026, N3008, N2412, N435);
buf BUF1 (N3027, N2975);
buf BUF1 (N3028, N3012);
nand NAND4 (N3029, N3004, N525, N954, N1547);
nor NOR3 (N3030, N3028, N872, N2575);
or OR4 (N3031, N3025, N2347, N2833, N1444);
or OR3 (N3032, N3019, N2143, N1828);
nor NOR4 (N3033, N3030, N1460, N2208, N192);
nand NAND2 (N3034, N3024, N2503);
or OR4 (N3035, N3029, N254, N674, N1484);
buf BUF1 (N3036, N3034);
buf BUF1 (N3037, N3027);
nor NOR4 (N3038, N3035, N2662, N445, N911);
not NOT1 (N3039, N3031);
nand NAND2 (N3040, N3026, N1123);
or OR4 (N3041, N3033, N2129, N959, N33);
not NOT1 (N3042, N3040);
and AND2 (N3043, N3015, N2265);
and AND4 (N3044, N3041, N1474, N728, N2556);
and AND3 (N3045, N3038, N2047, N15);
or OR2 (N3046, N3043, N1863);
and AND4 (N3047, N3042, N2356, N936, N1528);
or OR2 (N3048, N3037, N798);
nand NAND2 (N3049, N3045, N2959);
xor XOR2 (N3050, N3032, N2498);
or OR2 (N3051, N3048, N845);
buf BUF1 (N3052, N3050);
or OR2 (N3053, N3036, N74);
xor XOR2 (N3054, N3053, N2827);
buf BUF1 (N3055, N3052);
nand NAND2 (N3056, N3023, N1927);
nand NAND3 (N3057, N3055, N2615, N2573);
nand NAND3 (N3058, N3057, N124, N1651);
or OR4 (N3059, N3054, N378, N2122, N737);
buf BUF1 (N3060, N3056);
xor XOR2 (N3061, N3058, N1199);
not NOT1 (N3062, N3047);
nor NOR2 (N3063, N3039, N2051);
xor XOR2 (N3064, N3062, N2599);
not NOT1 (N3065, N3051);
not NOT1 (N3066, N3049);
xor XOR2 (N3067, N3063, N1125);
nor NOR4 (N3068, N3061, N2632, N2510, N1954);
buf BUF1 (N3069, N3067);
or OR4 (N3070, N3046, N2738, N644, N205);
buf BUF1 (N3071, N3068);
xor XOR2 (N3072, N3018, N1477);
not NOT1 (N3073, N3071);
nand NAND2 (N3074, N3070, N1030);
or OR4 (N3075, N3072, N2022, N1185, N2421);
xor XOR2 (N3076, N3060, N2235);
or OR3 (N3077, N3064, N664, N2307);
not NOT1 (N3078, N3066);
xor XOR2 (N3079, N3075, N201);
nor NOR4 (N3080, N3074, N663, N2209, N2449);
not NOT1 (N3081, N3079);
xor XOR2 (N3082, N3081, N2929);
or OR3 (N3083, N3076, N345, N1408);
or OR2 (N3084, N3082, N2621);
not NOT1 (N3085, N3073);
or OR3 (N3086, N3078, N3072, N1813);
and AND2 (N3087, N3044, N584);
nor NOR2 (N3088, N3065, N125);
nor NOR3 (N3089, N3083, N1067, N864);
or OR4 (N3090, N3077, N609, N1389, N1777);
and AND2 (N3091, N3084, N1126);
nor NOR3 (N3092, N3080, N1382, N1188);
not NOT1 (N3093, N3091);
nor NOR4 (N3094, N3086, N273, N2176, N1134);
buf BUF1 (N3095, N3087);
nand NAND4 (N3096, N3059, N2241, N2317, N2448);
or OR2 (N3097, N3089, N2120);
not NOT1 (N3098, N3096);
not NOT1 (N3099, N3098);
xor XOR2 (N3100, N3092, N653);
or OR3 (N3101, N3100, N2730, N2863);
nand NAND3 (N3102, N3095, N1652, N2259);
nand NAND4 (N3103, N3069, N1820, N396, N1339);
xor XOR2 (N3104, N3090, N1654);
buf BUF1 (N3105, N3102);
buf BUF1 (N3106, N3101);
nand NAND2 (N3107, N3106, N2733);
not NOT1 (N3108, N3085);
buf BUF1 (N3109, N3105);
buf BUF1 (N3110, N3103);
nor NOR2 (N3111, N3097, N2375);
nand NAND4 (N3112, N3109, N1175, N3040, N2508);
nor NOR2 (N3113, N3107, N1213);
not NOT1 (N3114, N3088);
xor XOR2 (N3115, N3111, N2913);
nand NAND3 (N3116, N3114, N1203, N440);
nor NOR3 (N3117, N3093, N2333, N2115);
not NOT1 (N3118, N3113);
not NOT1 (N3119, N3094);
or OR2 (N3120, N3117, N3014);
or OR2 (N3121, N3120, N958);
and AND3 (N3122, N3115, N753, N984);
not NOT1 (N3123, N3110);
or OR2 (N3124, N3123, N1729);
buf BUF1 (N3125, N3119);
nor NOR3 (N3126, N3112, N1128, N535);
or OR4 (N3127, N3121, N2156, N283, N1155);
buf BUF1 (N3128, N3124);
buf BUF1 (N3129, N3127);
buf BUF1 (N3130, N3104);
not NOT1 (N3131, N3126);
and AND3 (N3132, N3130, N1184, N1995);
or OR4 (N3133, N3122, N2436, N985, N463);
nand NAND2 (N3134, N3116, N482);
and AND2 (N3135, N3125, N2952);
and AND3 (N3136, N3108, N1999, N2874);
nand NAND2 (N3137, N3135, N1929);
and AND3 (N3138, N3131, N639, N2720);
or OR4 (N3139, N3128, N1549, N2378, N3121);
and AND2 (N3140, N3134, N3093);
nor NOR2 (N3141, N3138, N1822);
not NOT1 (N3142, N3118);
buf BUF1 (N3143, N3141);
nand NAND4 (N3144, N3136, N2884, N2917, N1497);
buf BUF1 (N3145, N3129);
or OR4 (N3146, N3139, N1892, N2013, N2439);
buf BUF1 (N3147, N3137);
and AND3 (N3148, N3145, N1001, N2270);
nor NOR4 (N3149, N3099, N1835, N1543, N1076);
and AND4 (N3150, N3140, N2934, N1469, N2596);
buf BUF1 (N3151, N3144);
nor NOR2 (N3152, N3150, N1826);
xor XOR2 (N3153, N3149, N578);
not NOT1 (N3154, N3151);
buf BUF1 (N3155, N3133);
nand NAND3 (N3156, N3148, N1839, N790);
xor XOR2 (N3157, N3147, N513);
or OR4 (N3158, N3132, N2485, N536, N1119);
or OR4 (N3159, N3155, N2026, N1298, N2153);
or OR3 (N3160, N3146, N1637, N1174);
nand NAND3 (N3161, N3154, N1387, N1068);
or OR2 (N3162, N3157, N2580);
nand NAND2 (N3163, N3159, N1153);
not NOT1 (N3164, N3143);
nand NAND4 (N3165, N3162, N627, N20, N1601);
nand NAND4 (N3166, N3160, N724, N1528, N2452);
nor NOR2 (N3167, N3161, N2041);
buf BUF1 (N3168, N3142);
nor NOR4 (N3169, N3158, N244, N785, N534);
buf BUF1 (N3170, N3166);
and AND2 (N3171, N3168, N2421);
nor NOR2 (N3172, N3171, N386);
nor NOR3 (N3173, N3163, N3119, N3061);
and AND2 (N3174, N3173, N1865);
and AND2 (N3175, N3174, N1273);
nor NOR2 (N3176, N3156, N1992);
not NOT1 (N3177, N3169);
buf BUF1 (N3178, N3176);
or OR4 (N3179, N3170, N198, N181, N502);
and AND3 (N3180, N3178, N1854, N3160);
or OR4 (N3181, N3165, N268, N2444, N2002);
buf BUF1 (N3182, N3180);
xor XOR2 (N3183, N3172, N1781);
and AND4 (N3184, N3181, N924, N2059, N2478);
buf BUF1 (N3185, N3184);
and AND3 (N3186, N3175, N1878, N2349);
buf BUF1 (N3187, N3167);
xor XOR2 (N3188, N3179, N1999);
and AND2 (N3189, N3153, N1226);
nand NAND2 (N3190, N3164, N424);
xor XOR2 (N3191, N3185, N2180);
nor NOR2 (N3192, N3187, N664);
and AND2 (N3193, N3152, N2429);
not NOT1 (N3194, N3189);
nand NAND4 (N3195, N3186, N546, N3066, N1415);
and AND3 (N3196, N3177, N309, N1188);
and AND3 (N3197, N3188, N1864, N2482);
nor NOR2 (N3198, N3183, N281);
xor XOR2 (N3199, N3195, N590);
not NOT1 (N3200, N3196);
and AND3 (N3201, N3192, N745, N1712);
not NOT1 (N3202, N3200);
not NOT1 (N3203, N3191);
or OR4 (N3204, N3193, N2124, N2863, N2827);
xor XOR2 (N3205, N3203, N3144);
buf BUF1 (N3206, N3198);
or OR4 (N3207, N3204, N2562, N1397, N1845);
nor NOR4 (N3208, N3205, N2910, N2761, N914);
buf BUF1 (N3209, N3197);
nand NAND4 (N3210, N3207, N2565, N2715, N1230);
or OR4 (N3211, N3194, N2563, N2850, N89);
nor NOR3 (N3212, N3190, N2126, N1846);
and AND4 (N3213, N3210, N2768, N1267, N2778);
nor NOR3 (N3214, N3211, N467, N880);
or OR3 (N3215, N3214, N1748, N2395);
nor NOR2 (N3216, N3212, N1383);
buf BUF1 (N3217, N3209);
xor XOR2 (N3218, N3206, N1033);
nor NOR4 (N3219, N3215, N92, N2037, N786);
xor XOR2 (N3220, N3213, N2872);
or OR4 (N3221, N3218, N1013, N795, N691);
buf BUF1 (N3222, N3202);
or OR3 (N3223, N3220, N1949, N1813);
buf BUF1 (N3224, N3216);
nor NOR4 (N3225, N3208, N2352, N838, N915);
not NOT1 (N3226, N3224);
nor NOR4 (N3227, N3217, N1026, N1207, N2257);
and AND4 (N3228, N3222, N1797, N111, N652);
nor NOR3 (N3229, N3182, N901, N886);
not NOT1 (N3230, N3225);
nor NOR2 (N3231, N3226, N443);
xor XOR2 (N3232, N3228, N1631);
and AND3 (N3233, N3230, N166, N936);
not NOT1 (N3234, N3219);
nor NOR3 (N3235, N3232, N1255, N3215);
buf BUF1 (N3236, N3227);
not NOT1 (N3237, N3199);
buf BUF1 (N3238, N3223);
xor XOR2 (N3239, N3201, N3175);
not NOT1 (N3240, N3233);
buf BUF1 (N3241, N3240);
nor NOR2 (N3242, N3231, N955);
nand NAND3 (N3243, N3235, N1645, N2994);
and AND3 (N3244, N3236, N1628, N3200);
buf BUF1 (N3245, N3237);
buf BUF1 (N3246, N3244);
nor NOR4 (N3247, N3242, N521, N483, N2578);
nand NAND2 (N3248, N3229, N2229);
nor NOR4 (N3249, N3245, N1749, N252, N1668);
nor NOR3 (N3250, N3239, N426, N1475);
not NOT1 (N3251, N3250);
nor NOR4 (N3252, N3234, N1618, N2135, N157);
and AND2 (N3253, N3249, N189);
nand NAND2 (N3254, N3247, N1355);
and AND2 (N3255, N3253, N1415);
buf BUF1 (N3256, N3241);
nand NAND4 (N3257, N3252, N1529, N1613, N640);
and AND3 (N3258, N3251, N2052, N738);
nand NAND3 (N3259, N3258, N562, N1666);
nand NAND2 (N3260, N3259, N2068);
or OR3 (N3261, N3221, N1205, N331);
or OR2 (N3262, N3248, N513);
or OR3 (N3263, N3238, N1773, N2970);
not NOT1 (N3264, N3254);
or OR3 (N3265, N3261, N597, N583);
and AND2 (N3266, N3256, N2191);
not NOT1 (N3267, N3260);
nor NOR2 (N3268, N3265, N323);
nor NOR3 (N3269, N3262, N22, N3216);
not NOT1 (N3270, N3246);
nand NAND3 (N3271, N3266, N587, N1958);
and AND3 (N3272, N3255, N2013, N1415);
not NOT1 (N3273, N3269);
buf BUF1 (N3274, N3267);
nor NOR3 (N3275, N3268, N2221, N122);
or OR3 (N3276, N3274, N449, N3164);
nand NAND3 (N3277, N3270, N2996, N3255);
and AND3 (N3278, N3277, N1006, N3025);
nand NAND4 (N3279, N3243, N985, N2818, N1957);
buf BUF1 (N3280, N3273);
and AND4 (N3281, N3271, N1805, N2128, N1010);
or OR4 (N3282, N3264, N1440, N1638, N2403);
xor XOR2 (N3283, N3257, N666);
buf BUF1 (N3284, N3275);
xor XOR2 (N3285, N3279, N2878);
not NOT1 (N3286, N3263);
buf BUF1 (N3287, N3284);
nor NOR2 (N3288, N3287, N2398);
buf BUF1 (N3289, N3278);
nand NAND3 (N3290, N3289, N1946, N710);
xor XOR2 (N3291, N3282, N919);
xor XOR2 (N3292, N3276, N321);
not NOT1 (N3293, N3290);
nand NAND3 (N3294, N3288, N1240, N192);
and AND2 (N3295, N3285, N1771);
nand NAND2 (N3296, N3280, N2580);
and AND4 (N3297, N3293, N1991, N758, N2331);
nand NAND3 (N3298, N3294, N1847, N2091);
and AND4 (N3299, N3283, N2188, N2074, N1012);
nand NAND3 (N3300, N3299, N8, N3117);
or OR3 (N3301, N3281, N78, N2026);
or OR3 (N3302, N3292, N1320, N1103);
nor NOR4 (N3303, N3296, N562, N2728, N280);
buf BUF1 (N3304, N3297);
or OR4 (N3305, N3303, N764, N140, N3046);
or OR4 (N3306, N3295, N1830, N455, N1777);
not NOT1 (N3307, N3305);
xor XOR2 (N3308, N3291, N681);
buf BUF1 (N3309, N3304);
nand NAND4 (N3310, N3298, N856, N1614, N36);
not NOT1 (N3311, N3300);
not NOT1 (N3312, N3310);
nor NOR3 (N3313, N3306, N357, N1986);
nor NOR4 (N3314, N3309, N1755, N3104, N93);
buf BUF1 (N3315, N3313);
nor NOR3 (N3316, N3272, N737, N1460);
not NOT1 (N3317, N3314);
nand NAND3 (N3318, N3307, N1441, N2461);
or OR3 (N3319, N3315, N175, N1226);
or OR2 (N3320, N3301, N760);
nor NOR2 (N3321, N3308, N1579);
nand NAND3 (N3322, N3317, N1680, N145);
not NOT1 (N3323, N3302);
nor NOR4 (N3324, N3318, N1320, N2371, N454);
and AND3 (N3325, N3323, N322, N1127);
nand NAND4 (N3326, N3321, N1948, N270, N2045);
nor NOR3 (N3327, N3286, N1007, N3089);
nor NOR3 (N3328, N3311, N786, N1147);
xor XOR2 (N3329, N3326, N208);
buf BUF1 (N3330, N3316);
buf BUF1 (N3331, N3328);
and AND3 (N3332, N3322, N1018, N2004);
nand NAND2 (N3333, N3330, N2289);
nor NOR4 (N3334, N3320, N355, N2259, N2186);
buf BUF1 (N3335, N3332);
or OR4 (N3336, N3327, N1564, N505, N2519);
buf BUF1 (N3337, N3335);
buf BUF1 (N3338, N3333);
not NOT1 (N3339, N3334);
nor NOR2 (N3340, N3319, N2934);
buf BUF1 (N3341, N3331);
and AND4 (N3342, N3325, N2563, N2164, N2218);
or OR3 (N3343, N3342, N2356, N1286);
buf BUF1 (N3344, N3336);
not NOT1 (N3345, N3329);
xor XOR2 (N3346, N3338, N2674);
xor XOR2 (N3347, N3312, N904);
xor XOR2 (N3348, N3339, N2040);
and AND3 (N3349, N3340, N1355, N3202);
nor NOR2 (N3350, N3324, N1873);
buf BUF1 (N3351, N3344);
or OR4 (N3352, N3341, N2262, N1039, N1687);
and AND4 (N3353, N3347, N2448, N2610, N580);
or OR4 (N3354, N3351, N2970, N1409, N1589);
not NOT1 (N3355, N3350);
nor NOR3 (N3356, N3343, N2719, N800);
nand NAND2 (N3357, N3346, N2152);
not NOT1 (N3358, N3355);
and AND3 (N3359, N3358, N2830, N3031);
nand NAND3 (N3360, N3349, N2773, N2657);
nand NAND2 (N3361, N3354, N648);
or OR3 (N3362, N3353, N2689, N2994);
and AND3 (N3363, N3356, N308, N2382);
nand NAND2 (N3364, N3359, N23);
and AND2 (N3365, N3348, N1086);
nor NOR4 (N3366, N3361, N2174, N1091, N3009);
not NOT1 (N3367, N3352);
nor NOR3 (N3368, N3357, N1214, N2303);
not NOT1 (N3369, N3365);
xor XOR2 (N3370, N3362, N299);
nand NAND2 (N3371, N3367, N3197);
nor NOR3 (N3372, N3363, N1722, N1890);
nor NOR4 (N3373, N3370, N2059, N7, N1905);
buf BUF1 (N3374, N3372);
xor XOR2 (N3375, N3364, N772);
and AND4 (N3376, N3374, N2333, N690, N2066);
or OR2 (N3377, N3368, N3255);
or OR4 (N3378, N3345, N223, N1789, N2576);
xor XOR2 (N3379, N3376, N946);
not NOT1 (N3380, N3378);
nand NAND4 (N3381, N3366, N2072, N1697, N1706);
or OR2 (N3382, N3373, N1072);
and AND4 (N3383, N3377, N1315, N1816, N2029);
not NOT1 (N3384, N3382);
not NOT1 (N3385, N3360);
and AND3 (N3386, N3369, N2004, N316);
or OR4 (N3387, N3379, N1148, N586, N1413);
nand NAND3 (N3388, N3337, N187, N629);
nor NOR4 (N3389, N3385, N1676, N1043, N1727);
nand NAND4 (N3390, N3380, N3049, N3094, N761);
nand NAND4 (N3391, N3375, N161, N1556, N984);
buf BUF1 (N3392, N3388);
nand NAND4 (N3393, N3381, N1579, N290, N2848);
nor NOR4 (N3394, N3386, N1995, N2772, N3356);
nand NAND3 (N3395, N3391, N1791, N2561);
xor XOR2 (N3396, N3389, N810);
and AND2 (N3397, N3371, N1403);
nand NAND4 (N3398, N3394, N1391, N2768, N2096);
nor NOR2 (N3399, N3398, N802);
nor NOR3 (N3400, N3399, N444, N714);
nor NOR3 (N3401, N3397, N860, N1246);
buf BUF1 (N3402, N3383);
and AND2 (N3403, N3387, N3201);
and AND4 (N3404, N3401, N2867, N916, N1580);
nor NOR2 (N3405, N3404, N738);
or OR3 (N3406, N3402, N1255, N904);
not NOT1 (N3407, N3393);
xor XOR2 (N3408, N3390, N2796);
nand NAND4 (N3409, N3406, N1826, N3106, N2495);
or OR2 (N3410, N3395, N240);
and AND4 (N3411, N3409, N2082, N2485, N1813);
nand NAND4 (N3412, N3396, N400, N2899, N1942);
buf BUF1 (N3413, N3412);
nand NAND2 (N3414, N3410, N2462);
or OR3 (N3415, N3414, N2661, N773);
nor NOR2 (N3416, N3405, N2825);
or OR4 (N3417, N3400, N3035, N3159, N1119);
buf BUF1 (N3418, N3411);
xor XOR2 (N3419, N3415, N578);
not NOT1 (N3420, N3407);
or OR3 (N3421, N3416, N2826, N3092);
buf BUF1 (N3422, N3403);
not NOT1 (N3423, N3419);
buf BUF1 (N3424, N3413);
xor XOR2 (N3425, N3421, N1133);
nor NOR4 (N3426, N3425, N662, N1328, N574);
nor NOR2 (N3427, N3424, N1510);
nor NOR4 (N3428, N3427, N2006, N196, N998);
or OR2 (N3429, N3417, N2896);
nor NOR4 (N3430, N3408, N1628, N3409, N1817);
xor XOR2 (N3431, N3384, N2323);
or OR4 (N3432, N3430, N2033, N1247, N1415);
not NOT1 (N3433, N3418);
xor XOR2 (N3434, N3428, N143);
buf BUF1 (N3435, N3420);
not NOT1 (N3436, N3392);
nor NOR3 (N3437, N3422, N2027, N646);
nor NOR2 (N3438, N3436, N2570);
nor NOR3 (N3439, N3438, N947, N2250);
or OR2 (N3440, N3423, N2916);
nand NAND3 (N3441, N3439, N3367, N1538);
nand NAND2 (N3442, N3435, N608);
not NOT1 (N3443, N3426);
nor NOR4 (N3444, N3442, N441, N2315, N3390);
nand NAND2 (N3445, N3444, N1412);
or OR4 (N3446, N3440, N1363, N2315, N525);
buf BUF1 (N3447, N3429);
xor XOR2 (N3448, N3443, N2706);
xor XOR2 (N3449, N3434, N2495);
and AND4 (N3450, N3446, N2380, N2010, N2569);
nor NOR2 (N3451, N3447, N2657);
xor XOR2 (N3452, N3431, N1237);
nor NOR3 (N3453, N3433, N1451, N3307);
or OR4 (N3454, N3452, N77, N1069, N1040);
xor XOR2 (N3455, N3453, N35);
nor NOR2 (N3456, N3445, N2193);
or OR2 (N3457, N3454, N3024);
or OR3 (N3458, N3441, N1321, N1280);
xor XOR2 (N3459, N3448, N1174);
nor NOR4 (N3460, N3437, N46, N59, N1273);
nand NAND4 (N3461, N3451, N1471, N999, N1085);
xor XOR2 (N3462, N3461, N2870);
nand NAND3 (N3463, N3457, N455, N2358);
xor XOR2 (N3464, N3455, N2870);
nor NOR2 (N3465, N3462, N1800);
xor XOR2 (N3466, N3460, N2303);
buf BUF1 (N3467, N3450);
buf BUF1 (N3468, N3432);
nor NOR3 (N3469, N3459, N476, N2495);
nor NOR3 (N3470, N3467, N1407, N619);
nand NAND2 (N3471, N3456, N1605);
nor NOR4 (N3472, N3449, N1895, N2142, N2675);
xor XOR2 (N3473, N3472, N2326);
and AND2 (N3474, N3473, N1955);
and AND4 (N3475, N3468, N854, N3226, N2718);
and AND2 (N3476, N3464, N115);
nand NAND2 (N3477, N3475, N826);
and AND3 (N3478, N3463, N1636, N560);
buf BUF1 (N3479, N3474);
or OR4 (N3480, N3469, N820, N2243, N1396);
or OR4 (N3481, N3479, N1893, N2563, N882);
nor NOR2 (N3482, N3480, N2703);
or OR2 (N3483, N3465, N3109);
xor XOR2 (N3484, N3483, N1196);
and AND4 (N3485, N3466, N1665, N286, N3189);
not NOT1 (N3486, N3471);
buf BUF1 (N3487, N3476);
buf BUF1 (N3488, N3478);
and AND4 (N3489, N3481, N138, N3485, N1581);
or OR2 (N3490, N19, N3324);
or OR3 (N3491, N3470, N503, N2157);
and AND4 (N3492, N3486, N3383, N1476, N2508);
xor XOR2 (N3493, N3492, N388);
nor NOR3 (N3494, N3458, N1757, N1913);
or OR2 (N3495, N3477, N362);
not NOT1 (N3496, N3487);
or OR3 (N3497, N3490, N3202, N3465);
and AND3 (N3498, N3489, N3493, N745);
and AND3 (N3499, N1460, N1055, N1976);
and AND4 (N3500, N3482, N2364, N1238, N1615);
nand NAND2 (N3501, N3484, N594);
nor NOR2 (N3502, N3500, N224);
buf BUF1 (N3503, N3501);
nand NAND2 (N3504, N3491, N1150);
xor XOR2 (N3505, N3498, N3215);
or OR4 (N3506, N3505, N2017, N3187, N2736);
not NOT1 (N3507, N3502);
nor NOR3 (N3508, N3507, N105, N1316);
nor NOR4 (N3509, N3495, N2625, N3258, N548);
and AND4 (N3510, N3506, N234, N1230, N3027);
not NOT1 (N3511, N3503);
nor NOR3 (N3512, N3499, N2524, N531);
buf BUF1 (N3513, N3512);
not NOT1 (N3514, N3513);
not NOT1 (N3515, N3496);
and AND2 (N3516, N3514, N3140);
buf BUF1 (N3517, N3497);
or OR2 (N3518, N3515, N1779);
nor NOR2 (N3519, N3494, N898);
nand NAND2 (N3520, N3488, N1354);
nand NAND2 (N3521, N3504, N1097);
and AND3 (N3522, N3518, N2107, N3125);
and AND4 (N3523, N3517, N512, N926, N3192);
or OR4 (N3524, N3523, N3308, N2214, N1901);
nand NAND2 (N3525, N3524, N1944);
buf BUF1 (N3526, N3521);
and AND2 (N3527, N3525, N472);
and AND2 (N3528, N3511, N3355);
and AND2 (N3529, N3527, N996);
and AND3 (N3530, N3529, N2494, N1658);
nor NOR3 (N3531, N3526, N3138, N2930);
nor NOR4 (N3532, N3519, N2878, N1731, N544);
not NOT1 (N3533, N3509);
xor XOR2 (N3534, N3532, N1966);
buf BUF1 (N3535, N3533);
or OR4 (N3536, N3516, N71, N2486, N2961);
buf BUF1 (N3537, N3531);
not NOT1 (N3538, N3530);
nand NAND2 (N3539, N3537, N3044);
or OR4 (N3540, N3534, N2991, N1246, N2244);
and AND2 (N3541, N3508, N752);
nor NOR3 (N3542, N3541, N656, N1268);
nand NAND3 (N3543, N3520, N3081, N1821);
xor XOR2 (N3544, N3538, N2796);
xor XOR2 (N3545, N3528, N2509);
buf BUF1 (N3546, N3540);
or OR2 (N3547, N3539, N60);
nand NAND2 (N3548, N3522, N3417);
not NOT1 (N3549, N3535);
buf BUF1 (N3550, N3536);
and AND2 (N3551, N3544, N399);
buf BUF1 (N3552, N3546);
nor NOR2 (N3553, N3547, N2930);
nand NAND4 (N3554, N3550, N3280, N764, N2030);
or OR2 (N3555, N3543, N3103);
or OR3 (N3556, N3549, N1409, N1398);
buf BUF1 (N3557, N3542);
xor XOR2 (N3558, N3555, N3298);
nor NOR3 (N3559, N3551, N1921, N1655);
xor XOR2 (N3560, N3557, N222);
xor XOR2 (N3561, N3560, N864);
not NOT1 (N3562, N3553);
not NOT1 (N3563, N3548);
xor XOR2 (N3564, N3556, N2037);
nand NAND2 (N3565, N3545, N8);
and AND4 (N3566, N3558, N1211, N1047, N2493);
not NOT1 (N3567, N3552);
buf BUF1 (N3568, N3565);
and AND2 (N3569, N3567, N757);
nor NOR4 (N3570, N3563, N3445, N2926, N1479);
or OR2 (N3571, N3559, N1521);
buf BUF1 (N3572, N3566);
buf BUF1 (N3573, N3564);
buf BUF1 (N3574, N3569);
and AND4 (N3575, N3562, N2082, N2987, N1047);
nor NOR3 (N3576, N3554, N1341, N2151);
not NOT1 (N3577, N3573);
nor NOR3 (N3578, N3561, N533, N2303);
xor XOR2 (N3579, N3510, N19);
buf BUF1 (N3580, N3578);
or OR4 (N3581, N3572, N1034, N223, N1545);
nand NAND3 (N3582, N3580, N497, N2117);
not NOT1 (N3583, N3570);
not NOT1 (N3584, N3579);
and AND3 (N3585, N3576, N906, N2608);
or OR3 (N3586, N3581, N1227, N2437);
buf BUF1 (N3587, N3568);
not NOT1 (N3588, N3585);
not NOT1 (N3589, N3588);
xor XOR2 (N3590, N3584, N2220);
and AND3 (N3591, N3582, N546, N500);
xor XOR2 (N3592, N3590, N2137);
nand NAND4 (N3593, N3589, N1540, N983, N1113);
buf BUF1 (N3594, N3577);
and AND2 (N3595, N3591, N2196);
and AND4 (N3596, N3574, N1807, N2137, N2928);
and AND3 (N3597, N3571, N3397, N261);
nand NAND2 (N3598, N3593, N1476);
and AND4 (N3599, N3596, N1253, N349, N284);
xor XOR2 (N3600, N3592, N2426);
xor XOR2 (N3601, N3586, N1724);
buf BUF1 (N3602, N3583);
buf BUF1 (N3603, N3600);
xor XOR2 (N3604, N3597, N3199);
or OR4 (N3605, N3595, N2040, N2389, N2585);
not NOT1 (N3606, N3603);
xor XOR2 (N3607, N3594, N1259);
nand NAND2 (N3608, N3601, N2513);
and AND2 (N3609, N3602, N847);
and AND3 (N3610, N3607, N1087, N55);
not NOT1 (N3611, N3609);
or OR4 (N3612, N3606, N2725, N256, N1072);
or OR2 (N3613, N3599, N2534);
or OR4 (N3614, N3587, N2481, N1895, N2538);
and AND4 (N3615, N3613, N3517, N1421, N2752);
and AND3 (N3616, N3575, N356, N686);
nor NOR4 (N3617, N3614, N2989, N666, N2203);
or OR4 (N3618, N3611, N2186, N2267, N979);
not NOT1 (N3619, N3616);
buf BUF1 (N3620, N3612);
buf BUF1 (N3621, N3610);
or OR3 (N3622, N3617, N416, N2213);
or OR4 (N3623, N3615, N1593, N806, N497);
buf BUF1 (N3624, N3622);
buf BUF1 (N3625, N3608);
nor NOR3 (N3626, N3604, N1005, N1438);
nand NAND4 (N3627, N3625, N1683, N1820, N3419);
nor NOR2 (N3628, N3618, N207);
nor NOR2 (N3629, N3598, N2517);
not NOT1 (N3630, N3621);
not NOT1 (N3631, N3605);
nand NAND4 (N3632, N3627, N455, N584, N2535);
not NOT1 (N3633, N3628);
nor NOR3 (N3634, N3632, N1896, N848);
and AND3 (N3635, N3626, N3223, N1600);
buf BUF1 (N3636, N3633);
nor NOR3 (N3637, N3629, N458, N1410);
xor XOR2 (N3638, N3637, N1477);
nand NAND3 (N3639, N3619, N2635, N3117);
or OR2 (N3640, N3636, N1505);
or OR2 (N3641, N3631, N2398);
not NOT1 (N3642, N3630);
nand NAND4 (N3643, N3640, N1699, N1434, N1942);
nand NAND2 (N3644, N3623, N2245);
or OR3 (N3645, N3634, N103, N52);
or OR4 (N3646, N3639, N830, N2861, N2139);
nor NOR2 (N3647, N3643, N1565);
not NOT1 (N3648, N3642);
and AND2 (N3649, N3648, N3424);
and AND3 (N3650, N3624, N3051, N2899);
buf BUF1 (N3651, N3650);
or OR2 (N3652, N3644, N2729);
xor XOR2 (N3653, N3638, N1778);
nor NOR3 (N3654, N3653, N887, N719);
or OR2 (N3655, N3647, N2614);
nand NAND3 (N3656, N3654, N1732, N3468);
not NOT1 (N3657, N3646);
or OR4 (N3658, N3620, N441, N1538, N2421);
buf BUF1 (N3659, N3641);
nand NAND3 (N3660, N3659, N2023, N1189);
nor NOR3 (N3661, N3649, N3181, N591);
buf BUF1 (N3662, N3645);
nor NOR2 (N3663, N3655, N2763);
and AND2 (N3664, N3662, N1347);
buf BUF1 (N3665, N3658);
or OR2 (N3666, N3663, N2723);
nand NAND4 (N3667, N3651, N364, N246, N3072);
nor NOR3 (N3668, N3652, N255, N636);
or OR2 (N3669, N3665, N3352);
buf BUF1 (N3670, N3664);
nor NOR4 (N3671, N3660, N1157, N1583, N2962);
and AND3 (N3672, N3656, N541, N3454);
or OR4 (N3673, N3669, N2075, N2815, N35);
and AND4 (N3674, N3661, N1486, N2783, N371);
and AND2 (N3675, N3672, N3453);
xor XOR2 (N3676, N3666, N1898);
xor XOR2 (N3677, N3671, N3574);
not NOT1 (N3678, N3667);
nor NOR2 (N3679, N3657, N33);
xor XOR2 (N3680, N3678, N2234);
buf BUF1 (N3681, N3677);
nand NAND4 (N3682, N3675, N140, N3633, N2798);
nand NAND4 (N3683, N3676, N2048, N3503, N3663);
or OR4 (N3684, N3681, N2627, N3669, N3264);
nand NAND3 (N3685, N3668, N2489, N2258);
and AND3 (N3686, N3679, N2830, N939);
or OR2 (N3687, N3685, N815);
not NOT1 (N3688, N3683);
or OR2 (N3689, N3674, N1112);
nor NOR4 (N3690, N3673, N646, N2829, N2663);
xor XOR2 (N3691, N3670, N2685);
xor XOR2 (N3692, N3691, N3565);
nor NOR2 (N3693, N3689, N2223);
not NOT1 (N3694, N3680);
and AND3 (N3695, N3687, N1382, N2066);
nor NOR4 (N3696, N3692, N2368, N1072, N1858);
or OR3 (N3697, N3635, N863, N1027);
nand NAND4 (N3698, N3693, N1800, N1325, N614);
buf BUF1 (N3699, N3690);
and AND2 (N3700, N3698, N411);
nor NOR4 (N3701, N3700, N2633, N1074, N1961);
buf BUF1 (N3702, N3694);
or OR2 (N3703, N3701, N3610);
nand NAND3 (N3704, N3703, N1219, N2134);
xor XOR2 (N3705, N3704, N2230);
not NOT1 (N3706, N3686);
or OR4 (N3707, N3705, N91, N946, N821);
or OR2 (N3708, N3695, N153);
buf BUF1 (N3709, N3696);
nor NOR3 (N3710, N3708, N1870, N382);
and AND3 (N3711, N3699, N68, N1910);
nand NAND3 (N3712, N3706, N3106, N2396);
nor NOR2 (N3713, N3712, N2829);
buf BUF1 (N3714, N3713);
or OR2 (N3715, N3710, N32);
buf BUF1 (N3716, N3702);
xor XOR2 (N3717, N3714, N3604);
or OR3 (N3718, N3716, N1048, N2023);
nand NAND3 (N3719, N3709, N3528, N800);
nor NOR3 (N3720, N3711, N2113, N581);
not NOT1 (N3721, N3707);
nor NOR4 (N3722, N3688, N154, N3554, N2389);
xor XOR2 (N3723, N3715, N950);
or OR2 (N3724, N3723, N1765);
buf BUF1 (N3725, N3722);
not NOT1 (N3726, N3718);
buf BUF1 (N3727, N3697);
and AND2 (N3728, N3720, N1572);
buf BUF1 (N3729, N3682);
xor XOR2 (N3730, N3725, N83);
nand NAND2 (N3731, N3730, N1834);
buf BUF1 (N3732, N3717);
nor NOR4 (N3733, N3726, N2420, N2731, N1898);
nand NAND3 (N3734, N3684, N2905, N3443);
not NOT1 (N3735, N3731);
not NOT1 (N3736, N3733);
not NOT1 (N3737, N3724);
or OR3 (N3738, N3734, N127, N1096);
nor NOR2 (N3739, N3721, N3569);
and AND2 (N3740, N3737, N2748);
xor XOR2 (N3741, N3729, N852);
nor NOR3 (N3742, N3727, N2182, N1124);
nand NAND3 (N3743, N3732, N322, N1584);
and AND3 (N3744, N3740, N1723, N2843);
not NOT1 (N3745, N3719);
nand NAND3 (N3746, N3741, N765, N1087);
nor NOR4 (N3747, N3736, N2049, N201, N2113);
not NOT1 (N3748, N3745);
not NOT1 (N3749, N3739);
nor NOR4 (N3750, N3738, N2892, N2940, N33);
or OR2 (N3751, N3747, N1352);
or OR2 (N3752, N3749, N2);
or OR2 (N3753, N3751, N1265);
buf BUF1 (N3754, N3753);
or OR2 (N3755, N3744, N2180);
nand NAND2 (N3756, N3752, N965);
xor XOR2 (N3757, N3743, N898);
and AND2 (N3758, N3756, N3153);
nand NAND2 (N3759, N3758, N1942);
xor XOR2 (N3760, N3759, N391);
or OR3 (N3761, N3728, N1089, N3080);
and AND3 (N3762, N3755, N3647, N2626);
or OR3 (N3763, N3748, N1070, N265);
not NOT1 (N3764, N3742);
xor XOR2 (N3765, N3754, N1575);
or OR3 (N3766, N3763, N3697, N2631);
nor NOR4 (N3767, N3762, N1750, N1532, N2751);
buf BUF1 (N3768, N3757);
not NOT1 (N3769, N3767);
or OR4 (N3770, N3760, N3521, N1348, N2938);
nor NOR2 (N3771, N3735, N875);
xor XOR2 (N3772, N3746, N3402);
buf BUF1 (N3773, N3769);
or OR3 (N3774, N3768, N290, N699);
or OR3 (N3775, N3771, N2447, N3586);
nor NOR4 (N3776, N3764, N1914, N1132, N3090);
nand NAND3 (N3777, N3772, N2468, N1486);
nand NAND4 (N3778, N3765, N2917, N48, N607);
buf BUF1 (N3779, N3778);
and AND2 (N3780, N3773, N1782);
xor XOR2 (N3781, N3780, N90);
nor NOR3 (N3782, N3761, N3545, N815);
buf BUF1 (N3783, N3750);
nand NAND4 (N3784, N3782, N2600, N3733, N3497);
nor NOR3 (N3785, N3776, N2192, N1713);
or OR4 (N3786, N3784, N2948, N1608, N395);
nand NAND2 (N3787, N3775, N2008);
not NOT1 (N3788, N3785);
buf BUF1 (N3789, N3766);
or OR4 (N3790, N3787, N1111, N3485, N1564);
xor XOR2 (N3791, N3789, N338);
and AND2 (N3792, N3790, N1629);
not NOT1 (N3793, N3770);
xor XOR2 (N3794, N3791, N1466);
nand NAND4 (N3795, N3794, N2216, N832, N2766);
xor XOR2 (N3796, N3792, N463);
nand NAND4 (N3797, N3786, N1934, N1833, N3633);
xor XOR2 (N3798, N3777, N1574);
nor NOR2 (N3799, N3781, N682);
or OR2 (N3800, N3795, N697);
not NOT1 (N3801, N3774);
nor NOR3 (N3802, N3779, N2912, N2768);
nor NOR2 (N3803, N3798, N1715);
or OR4 (N3804, N3788, N2833, N1656, N3219);
and AND3 (N3805, N3783, N892, N3760);
xor XOR2 (N3806, N3802, N1559);
nor NOR2 (N3807, N3797, N3245);
xor XOR2 (N3808, N3807, N2980);
and AND3 (N3809, N3799, N317, N147);
or OR4 (N3810, N3803, N2972, N2890, N3294);
xor XOR2 (N3811, N3801, N3002);
buf BUF1 (N3812, N3809);
nor NOR3 (N3813, N3793, N3228, N2106);
not NOT1 (N3814, N3800);
and AND3 (N3815, N3814, N1680, N2064);
nor NOR2 (N3816, N3813, N366);
xor XOR2 (N3817, N3811, N2519);
nor NOR2 (N3818, N3805, N2686);
buf BUF1 (N3819, N3804);
not NOT1 (N3820, N3819);
or OR2 (N3821, N3818, N35);
nand NAND4 (N3822, N3816, N3307, N3367, N1642);
buf BUF1 (N3823, N3817);
xor XOR2 (N3824, N3815, N2669);
or OR3 (N3825, N3812, N981, N2306);
buf BUF1 (N3826, N3796);
nand NAND2 (N3827, N3820, N1882);
nor NOR3 (N3828, N3806, N1361, N101);
nor NOR2 (N3829, N3810, N194);
nand NAND2 (N3830, N3826, N1536);
buf BUF1 (N3831, N3821);
buf BUF1 (N3832, N3825);
or OR4 (N3833, N3822, N1188, N2236, N1783);
or OR4 (N3834, N3808, N723, N1314, N1253);
nor NOR2 (N3835, N3832, N412);
not NOT1 (N3836, N3834);
xor XOR2 (N3837, N3824, N49);
and AND2 (N3838, N3836, N3150);
or OR3 (N3839, N3828, N3487, N61);
buf BUF1 (N3840, N3833);
nor NOR2 (N3841, N3827, N2853);
and AND3 (N3842, N3823, N1363, N1943);
xor XOR2 (N3843, N3837, N3373);
or OR4 (N3844, N3843, N2620, N491, N638);
buf BUF1 (N3845, N3844);
nor NOR4 (N3846, N3841, N1793, N753, N55);
not NOT1 (N3847, N3830);
xor XOR2 (N3848, N3847, N238);
xor XOR2 (N3849, N3842, N689);
xor XOR2 (N3850, N3838, N1717);
and AND3 (N3851, N3848, N1255, N1137);
buf BUF1 (N3852, N3839);
not NOT1 (N3853, N3846);
xor XOR2 (N3854, N3849, N2458);
nor NOR2 (N3855, N3854, N2596);
and AND4 (N3856, N3840, N3127, N3005, N290);
nor NOR2 (N3857, N3851, N3184);
xor XOR2 (N3858, N3856, N3026);
xor XOR2 (N3859, N3858, N2559);
and AND2 (N3860, N3850, N1028);
and AND2 (N3861, N3859, N3263);
nand NAND2 (N3862, N3831, N1700);
or OR4 (N3863, N3861, N583, N2867, N3616);
nand NAND3 (N3864, N3852, N618, N758);
nor NOR2 (N3865, N3853, N1496);
not NOT1 (N3866, N3863);
xor XOR2 (N3867, N3835, N380);
and AND3 (N3868, N3867, N2758, N2897);
nand NAND3 (N3869, N3862, N712, N2552);
buf BUF1 (N3870, N3829);
xor XOR2 (N3871, N3870, N1537);
and AND3 (N3872, N3866, N1117, N2311);
or OR3 (N3873, N3868, N2262, N335);
not NOT1 (N3874, N3857);
or OR2 (N3875, N3873, N1938);
or OR4 (N3876, N3860, N3196, N1122, N1295);
nor NOR3 (N3877, N3876, N3341, N2703);
not NOT1 (N3878, N3874);
nand NAND4 (N3879, N3855, N848, N1220, N85);
xor XOR2 (N3880, N3872, N3596);
buf BUF1 (N3881, N3879);
nand NAND2 (N3882, N3845, N3850);
nor NOR2 (N3883, N3882, N1998);
nor NOR4 (N3884, N3869, N32, N3341, N1267);
nor NOR3 (N3885, N3875, N2928, N3758);
nor NOR4 (N3886, N3878, N2031, N3191, N1367);
xor XOR2 (N3887, N3881, N3612);
buf BUF1 (N3888, N3880);
or OR4 (N3889, N3871, N2814, N2273, N1700);
not NOT1 (N3890, N3883);
nand NAND3 (N3891, N3890, N1436, N125);
not NOT1 (N3892, N3888);
xor XOR2 (N3893, N3877, N3454);
nor NOR4 (N3894, N3892, N1655, N2801, N3788);
or OR2 (N3895, N3889, N3519);
xor XOR2 (N3896, N3894, N3797);
nand NAND2 (N3897, N3886, N2103);
buf BUF1 (N3898, N3895);
buf BUF1 (N3899, N3885);
nand NAND4 (N3900, N3898, N2121, N300, N118);
nor NOR4 (N3901, N3884, N2495, N2581, N3159);
xor XOR2 (N3902, N3865, N2878);
nand NAND4 (N3903, N3893, N2114, N3401, N2591);
xor XOR2 (N3904, N3903, N1530);
nand NAND3 (N3905, N3896, N2441, N2616);
and AND3 (N3906, N3905, N2581, N3361);
nor NOR3 (N3907, N3901, N1314, N3278);
or OR3 (N3908, N3907, N666, N407);
nor NOR3 (N3909, N3900, N2015, N3880);
not NOT1 (N3910, N3906);
nor NOR3 (N3911, N3897, N2337, N3277);
not NOT1 (N3912, N3909);
not NOT1 (N3913, N3864);
nand NAND4 (N3914, N3911, N439, N2161, N1094);
xor XOR2 (N3915, N3912, N317);
nor NOR3 (N3916, N3891, N710, N2162);
xor XOR2 (N3917, N3916, N872);
and AND4 (N3918, N3910, N675, N1506, N3467);
buf BUF1 (N3919, N3915);
or OR4 (N3920, N3917, N3840, N3530, N859);
xor XOR2 (N3921, N3899, N804);
or OR4 (N3922, N3918, N3385, N3655, N1963);
buf BUF1 (N3923, N3920);
xor XOR2 (N3924, N3919, N3827);
nand NAND3 (N3925, N3924, N1156, N742);
nor NOR3 (N3926, N3902, N3832, N676);
and AND2 (N3927, N3887, N594);
xor XOR2 (N3928, N3923, N2918);
not NOT1 (N3929, N3921);
not NOT1 (N3930, N3929);
buf BUF1 (N3931, N3927);
nor NOR2 (N3932, N3913, N1284);
xor XOR2 (N3933, N3932, N64);
or OR3 (N3934, N3922, N99, N2387);
xor XOR2 (N3935, N3928, N439);
buf BUF1 (N3936, N3908);
nor NOR2 (N3937, N3914, N2660);
nand NAND2 (N3938, N3935, N2380);
and AND3 (N3939, N3936, N1375, N866);
and AND2 (N3940, N3904, N1352);
not NOT1 (N3941, N3925);
or OR2 (N3942, N3930, N1519);
and AND4 (N3943, N3926, N1590, N2355, N3191);
buf BUF1 (N3944, N3940);
xor XOR2 (N3945, N3943, N2797);
xor XOR2 (N3946, N3939, N3678);
or OR3 (N3947, N3937, N3825, N2863);
nor NOR3 (N3948, N3941, N1750, N735);
xor XOR2 (N3949, N3942, N1925);
and AND3 (N3950, N3938, N3465, N3226);
or OR4 (N3951, N3946, N2334, N1373, N2837);
not NOT1 (N3952, N3951);
not NOT1 (N3953, N3934);
not NOT1 (N3954, N3947);
nand NAND3 (N3955, N3954, N93, N1076);
buf BUF1 (N3956, N3953);
xor XOR2 (N3957, N3950, N2614);
or OR4 (N3958, N3955, N1153, N2802, N3401);
xor XOR2 (N3959, N3931, N1915);
nor NOR2 (N3960, N3945, N1291);
nand NAND4 (N3961, N3957, N3712, N2815, N1766);
nand NAND4 (N3962, N3961, N165, N1765, N2146);
or OR2 (N3963, N3959, N3315);
buf BUF1 (N3964, N3949);
and AND4 (N3965, N3956, N2423, N392, N3541);
or OR2 (N3966, N3948, N2031);
and AND2 (N3967, N3964, N3165);
buf BUF1 (N3968, N3966);
and AND2 (N3969, N3944, N2725);
xor XOR2 (N3970, N3958, N2485);
or OR3 (N3971, N3968, N355, N214);
not NOT1 (N3972, N3963);
or OR2 (N3973, N3933, N233);
and AND3 (N3974, N3952, N2561, N214);
and AND4 (N3975, N3973, N1052, N1765, N1203);
or OR4 (N3976, N3969, N706, N639, N628);
nor NOR4 (N3977, N3974, N3818, N3670, N2711);
nor NOR2 (N3978, N3970, N3251);
nand NAND4 (N3979, N3971, N471, N1955, N3754);
or OR2 (N3980, N3977, N2438);
or OR4 (N3981, N3965, N3900, N2143, N2070);
nand NAND2 (N3982, N3980, N1412);
buf BUF1 (N3983, N3975);
nand NAND2 (N3984, N3981, N3865);
nor NOR3 (N3985, N3983, N1018, N1900);
xor XOR2 (N3986, N3960, N3317);
not NOT1 (N3987, N3967);
buf BUF1 (N3988, N3979);
and AND3 (N3989, N3982, N409, N1338);
xor XOR2 (N3990, N3985, N1539);
or OR3 (N3991, N3976, N285, N2106);
or OR4 (N3992, N3987, N1857, N2890, N3602);
buf BUF1 (N3993, N3990);
buf BUF1 (N3994, N3992);
buf BUF1 (N3995, N3994);
and AND2 (N3996, N3984, N1446);
and AND4 (N3997, N3993, N796, N3834, N1895);
or OR4 (N3998, N3972, N2434, N1221, N3144);
xor XOR2 (N3999, N3991, N796);
buf BUF1 (N4000, N3989);
nor NOR4 (N4001, N3998, N61, N3907, N3894);
xor XOR2 (N4002, N3999, N1789);
or OR3 (N4003, N3962, N2095, N640);
buf BUF1 (N4004, N3978);
or OR4 (N4005, N3997, N1633, N44, N2975);
or OR2 (N4006, N4000, N639);
buf BUF1 (N4007, N4006);
nor NOR3 (N4008, N4004, N1141, N2643);
or OR3 (N4009, N3996, N955, N2824);
and AND3 (N4010, N4003, N167, N2910);
not NOT1 (N4011, N3988);
or OR4 (N4012, N4007, N150, N649, N2210);
buf BUF1 (N4013, N4005);
xor XOR2 (N4014, N3995, N836);
not NOT1 (N4015, N4014);
nand NAND4 (N4016, N4013, N2534, N415, N2678);
buf BUF1 (N4017, N4012);
or OR2 (N4018, N3986, N3250);
nor NOR4 (N4019, N4015, N3791, N182, N3790);
not NOT1 (N4020, N4018);
or OR3 (N4021, N4008, N1583, N2522);
or OR3 (N4022, N4009, N3471, N138);
buf BUF1 (N4023, N4011);
not NOT1 (N4024, N4016);
and AND2 (N4025, N4001, N323);
nor NOR2 (N4026, N4017, N623);
nor NOR3 (N4027, N4021, N1252, N1939);
and AND4 (N4028, N4020, N120, N420, N2469);
or OR2 (N4029, N4023, N2450);
xor XOR2 (N4030, N4026, N3428);
nand NAND4 (N4031, N4002, N1827, N464, N506);
buf BUF1 (N4032, N4022);
and AND3 (N4033, N4019, N3839, N1225);
nand NAND4 (N4034, N4025, N596, N186, N2755);
or OR2 (N4035, N4034, N3880);
nor NOR4 (N4036, N4027, N3821, N1632, N109);
nor NOR3 (N4037, N4028, N2256, N1185);
not NOT1 (N4038, N4030);
or OR3 (N4039, N4032, N4027, N2180);
buf BUF1 (N4040, N4031);
or OR2 (N4041, N4024, N2511);
buf BUF1 (N4042, N4038);
xor XOR2 (N4043, N4042, N2890);
xor XOR2 (N4044, N4037, N1376);
buf BUF1 (N4045, N4029);
nand NAND3 (N4046, N4035, N1524, N1867);
buf BUF1 (N4047, N4045);
nor NOR2 (N4048, N4010, N2512);
not NOT1 (N4049, N4043);
buf BUF1 (N4050, N4040);
xor XOR2 (N4051, N4049, N380);
and AND4 (N4052, N4047, N3639, N1596, N1097);
nor NOR2 (N4053, N4039, N1121);
not NOT1 (N4054, N4052);
and AND4 (N4055, N4053, N3171, N2079, N3463);
nand NAND3 (N4056, N4051, N1734, N1189);
nand NAND3 (N4057, N4041, N3520, N65);
or OR4 (N4058, N4054, N2041, N3967, N2410);
nor NOR4 (N4059, N4058, N1365, N2562, N1912);
or OR3 (N4060, N4056, N2653, N3827);
nor NOR4 (N4061, N4048, N3680, N2601, N2104);
not NOT1 (N4062, N4055);
or OR3 (N4063, N4062, N1923, N2725);
xor XOR2 (N4064, N4050, N1832);
xor XOR2 (N4065, N4061, N4036);
not NOT1 (N4066, N189);
xor XOR2 (N4067, N4059, N2029);
buf BUF1 (N4068, N4033);
or OR3 (N4069, N4065, N1734, N96);
nand NAND3 (N4070, N4066, N3021, N1360);
nand NAND2 (N4071, N4063, N3138);
not NOT1 (N4072, N4069);
buf BUF1 (N4073, N4071);
nand NAND2 (N4074, N4067, N3637);
buf BUF1 (N4075, N4073);
nor NOR2 (N4076, N4070, N3583);
xor XOR2 (N4077, N4068, N1879);
xor XOR2 (N4078, N4074, N436);
nand NAND2 (N4079, N4078, N3970);
and AND2 (N4080, N4077, N2582);
not NOT1 (N4081, N4080);
not NOT1 (N4082, N4060);
not NOT1 (N4083, N4082);
not NOT1 (N4084, N4083);
buf BUF1 (N4085, N4079);
not NOT1 (N4086, N4084);
nor NOR3 (N4087, N4064, N762, N1954);
and AND4 (N4088, N4057, N2028, N1277, N3269);
buf BUF1 (N4089, N4075);
nor NOR4 (N4090, N4076, N1527, N908, N187);
or OR3 (N4091, N4088, N3460, N2199);
not NOT1 (N4092, N4085);
not NOT1 (N4093, N4089);
buf BUF1 (N4094, N4081);
xor XOR2 (N4095, N4091, N835);
nand NAND2 (N4096, N4046, N2189);
nor NOR4 (N4097, N4094, N2189, N3488, N1876);
not NOT1 (N4098, N4092);
xor XOR2 (N4099, N4044, N1613);
buf BUF1 (N4100, N4087);
nand NAND2 (N4101, N4090, N3370);
xor XOR2 (N4102, N4093, N941);
xor XOR2 (N4103, N4098, N703);
not NOT1 (N4104, N4095);
xor XOR2 (N4105, N4072, N3474);
or OR2 (N4106, N4097, N4010);
and AND2 (N4107, N4103, N1008);
and AND3 (N4108, N4099, N2518, N3445);
buf BUF1 (N4109, N4107);
nand NAND4 (N4110, N4096, N2702, N1922, N3354);
or OR2 (N4111, N4109, N3469);
buf BUF1 (N4112, N4110);
nand NAND4 (N4113, N4086, N722, N2133, N4030);
xor XOR2 (N4114, N4102, N117);
buf BUF1 (N4115, N4114);
nand NAND3 (N4116, N4111, N3472, N3826);
or OR2 (N4117, N4101, N451);
nor NOR3 (N4118, N4113, N531, N3160);
nor NOR2 (N4119, N4100, N3249);
buf BUF1 (N4120, N4117);
nand NAND2 (N4121, N4106, N392);
not NOT1 (N4122, N4112);
nor NOR4 (N4123, N4118, N3601, N2961, N98);
nand NAND3 (N4124, N4115, N3865, N3875);
or OR4 (N4125, N4116, N1481, N590, N992);
buf BUF1 (N4126, N4108);
not NOT1 (N4127, N4123);
or OR3 (N4128, N4126, N2867, N3049);
nor NOR3 (N4129, N4105, N1445, N690);
xor XOR2 (N4130, N4125, N3055);
buf BUF1 (N4131, N4120);
nor NOR3 (N4132, N4131, N3505, N2810);
and AND2 (N4133, N4130, N1846);
and AND4 (N4134, N4124, N2599, N438, N3897);
buf BUF1 (N4135, N4128);
buf BUF1 (N4136, N4119);
buf BUF1 (N4137, N4132);
xor XOR2 (N4138, N4136, N2555);
or OR4 (N4139, N4104, N3477, N379, N1331);
buf BUF1 (N4140, N4122);
nor NOR2 (N4141, N4137, N2639);
not NOT1 (N4142, N4134);
buf BUF1 (N4143, N4138);
xor XOR2 (N4144, N4133, N393);
or OR4 (N4145, N4141, N2907, N513, N1845);
and AND3 (N4146, N4129, N3254, N2160);
and AND2 (N4147, N4139, N147);
and AND3 (N4148, N4145, N3742, N995);
nand NAND2 (N4149, N4146, N629);
nand NAND4 (N4150, N4147, N91, N1076, N2163);
buf BUF1 (N4151, N4142);
not NOT1 (N4152, N4135);
buf BUF1 (N4153, N4121);
not NOT1 (N4154, N4140);
nor NOR4 (N4155, N4143, N2466, N2712, N770);
and AND4 (N4156, N4152, N3853, N512, N3584);
buf BUF1 (N4157, N4148);
not NOT1 (N4158, N4144);
and AND4 (N4159, N4150, N10, N598, N1329);
or OR3 (N4160, N4127, N1617, N2033);
buf BUF1 (N4161, N4156);
buf BUF1 (N4162, N4160);
nand NAND2 (N4163, N4157, N3821);
nor NOR4 (N4164, N4155, N1135, N3466, N1735);
nor NOR4 (N4165, N4163, N3826, N2220, N3618);
not NOT1 (N4166, N4149);
nor NOR3 (N4167, N4166, N2512, N1152);
buf BUF1 (N4168, N4153);
or OR3 (N4169, N4158, N2758, N2638);
nor NOR4 (N4170, N4164, N1195, N1943, N2083);
nor NOR3 (N4171, N4159, N2110, N143);
nand NAND3 (N4172, N4162, N1395, N1916);
or OR3 (N4173, N4171, N1779, N3076);
nand NAND2 (N4174, N4173, N1705);
not NOT1 (N4175, N4172);
buf BUF1 (N4176, N4165);
or OR3 (N4177, N4167, N1982, N1867);
buf BUF1 (N4178, N4174);
nor NOR3 (N4179, N4175, N629, N1678);
and AND3 (N4180, N4168, N2770, N3794);
nor NOR3 (N4181, N4169, N3829, N1005);
buf BUF1 (N4182, N4181);
nand NAND3 (N4183, N4179, N2623, N641);
nor NOR2 (N4184, N4178, N3105);
nor NOR4 (N4185, N4180, N1692, N3395, N3336);
xor XOR2 (N4186, N4182, N324);
and AND3 (N4187, N4186, N3548, N1446);
or OR2 (N4188, N4151, N1762);
xor XOR2 (N4189, N4170, N1101);
nand NAND3 (N4190, N4176, N1555, N1496);
or OR3 (N4191, N4154, N3387, N2138);
and AND4 (N4192, N4184, N2851, N2534, N2514);
xor XOR2 (N4193, N4187, N3854);
buf BUF1 (N4194, N4177);
buf BUF1 (N4195, N4161);
buf BUF1 (N4196, N4188);
nor NOR2 (N4197, N4196, N3059);
and AND2 (N4198, N4192, N1069);
nor NOR2 (N4199, N4197, N3203);
not NOT1 (N4200, N4195);
buf BUF1 (N4201, N4190);
buf BUF1 (N4202, N4183);
buf BUF1 (N4203, N4193);
nand NAND3 (N4204, N4191, N882, N3725);
or OR4 (N4205, N4202, N1720, N527, N2791);
nor NOR3 (N4206, N4201, N498, N3383);
xor XOR2 (N4207, N4205, N3292);
not NOT1 (N4208, N4189);
or OR4 (N4209, N4198, N666, N2699, N223);
not NOT1 (N4210, N4208);
nand NAND2 (N4211, N4194, N447);
or OR4 (N4212, N4200, N648, N1280, N1442);
nor NOR2 (N4213, N4211, N2232);
nor NOR3 (N4214, N4204, N2756, N2189);
buf BUF1 (N4215, N4210);
or OR4 (N4216, N4207, N2798, N2221, N3894);
nand NAND3 (N4217, N4206, N1610, N1318);
or OR3 (N4218, N4199, N3541, N3287);
nor NOR2 (N4219, N4216, N1794);
xor XOR2 (N4220, N4213, N4001);
nor NOR4 (N4221, N4219, N1732, N311, N1991);
nand NAND2 (N4222, N4209, N1379);
and AND3 (N4223, N4217, N2157, N2009);
not NOT1 (N4224, N4220);
not NOT1 (N4225, N4203);
xor XOR2 (N4226, N4218, N1356);
or OR4 (N4227, N4185, N251, N3804, N3012);
nand NAND3 (N4228, N4221, N4116, N4207);
nor NOR4 (N4229, N4225, N654, N2250, N477);
or OR3 (N4230, N4223, N3517, N4137);
and AND2 (N4231, N4212, N4133);
not NOT1 (N4232, N4228);
xor XOR2 (N4233, N4231, N441);
nand NAND2 (N4234, N4214, N429);
xor XOR2 (N4235, N4229, N1675);
and AND2 (N4236, N4232, N2320);
buf BUF1 (N4237, N4227);
not NOT1 (N4238, N4230);
not NOT1 (N4239, N4238);
and AND3 (N4240, N4215, N3296, N2874);
buf BUF1 (N4241, N4236);
or OR4 (N4242, N4224, N3173, N1514, N1162);
nor NOR2 (N4243, N4237, N1590);
buf BUF1 (N4244, N4235);
or OR2 (N4245, N4239, N1064);
nand NAND4 (N4246, N4233, N110, N1281, N3975);
buf BUF1 (N4247, N4244);
buf BUF1 (N4248, N4247);
buf BUF1 (N4249, N4242);
nor NOR4 (N4250, N4234, N882, N2850, N202);
not NOT1 (N4251, N4222);
nand NAND4 (N4252, N4249, N1061, N1786, N709);
not NOT1 (N4253, N4243);
not NOT1 (N4254, N4251);
nor NOR3 (N4255, N4248, N1001, N3686);
and AND4 (N4256, N4226, N4141, N3575, N3515);
or OR2 (N4257, N4253, N811);
and AND4 (N4258, N4256, N2646, N3417, N2847);
and AND3 (N4259, N4257, N639, N2786);
not NOT1 (N4260, N4246);
nor NOR3 (N4261, N4240, N1684, N973);
buf BUF1 (N4262, N4261);
nor NOR4 (N4263, N4252, N332, N2864, N2445);
buf BUF1 (N4264, N4263);
not NOT1 (N4265, N4260);
and AND4 (N4266, N4245, N2529, N968, N3234);
and AND4 (N4267, N4262, N431, N2422, N1904);
and AND4 (N4268, N4266, N2779, N2724, N2312);
buf BUF1 (N4269, N4258);
not NOT1 (N4270, N4267);
not NOT1 (N4271, N4264);
or OR2 (N4272, N4269, N2840);
or OR3 (N4273, N4255, N441, N1474);
buf BUF1 (N4274, N4250);
not NOT1 (N4275, N4268);
nand NAND3 (N4276, N4270, N3873, N2672);
not NOT1 (N4277, N4275);
or OR2 (N4278, N4241, N1392);
nand NAND2 (N4279, N4277, N2310);
nand NAND4 (N4280, N4254, N195, N2423, N1699);
nand NAND3 (N4281, N4265, N3322, N1071);
not NOT1 (N4282, N4276);
nand NAND2 (N4283, N4259, N1371);
not NOT1 (N4284, N4278);
nand NAND4 (N4285, N4280, N1686, N2836, N1121);
or OR3 (N4286, N4281, N2768, N1387);
nand NAND4 (N4287, N4286, N472, N253, N2230);
or OR3 (N4288, N4283, N1546, N4230);
not NOT1 (N4289, N4273);
nand NAND4 (N4290, N4288, N3825, N1921, N3275);
and AND3 (N4291, N4285, N895, N3998);
nand NAND4 (N4292, N4287, N3679, N3921, N1446);
buf BUF1 (N4293, N4290);
or OR3 (N4294, N4279, N79, N3663);
not NOT1 (N4295, N4274);
not NOT1 (N4296, N4272);
buf BUF1 (N4297, N4271);
buf BUF1 (N4298, N4292);
nand NAND4 (N4299, N4298, N3686, N467, N1662);
and AND4 (N4300, N4296, N2944, N486, N2009);
nand NAND2 (N4301, N4297, N942);
buf BUF1 (N4302, N4284);
not NOT1 (N4303, N4291);
not NOT1 (N4304, N4282);
or OR4 (N4305, N4301, N323, N3027, N2038);
not NOT1 (N4306, N4289);
buf BUF1 (N4307, N4293);
not NOT1 (N4308, N4294);
or OR2 (N4309, N4295, N1588);
and AND2 (N4310, N4304, N3775);
nand NAND4 (N4311, N4308, N2141, N1288, N920);
nand NAND4 (N4312, N4302, N2819, N2883, N2349);
or OR4 (N4313, N4303, N1112, N2176, N579);
and AND2 (N4314, N4312, N3635);
nor NOR4 (N4315, N4311, N1076, N2234, N2326);
not NOT1 (N4316, N4309);
buf BUF1 (N4317, N4307);
or OR3 (N4318, N4300, N750, N2789);
buf BUF1 (N4319, N4306);
and AND4 (N4320, N4310, N1787, N3822, N2373);
xor XOR2 (N4321, N4315, N2141);
nor NOR3 (N4322, N4299, N1716, N2198);
nor NOR3 (N4323, N4313, N1427, N193);
or OR4 (N4324, N4305, N2581, N2330, N1861);
or OR2 (N4325, N4316, N2325);
nor NOR2 (N4326, N4319, N1435);
xor XOR2 (N4327, N4318, N3713);
buf BUF1 (N4328, N4320);
and AND4 (N4329, N4326, N190, N269, N742);
and AND4 (N4330, N4328, N4246, N15, N297);
buf BUF1 (N4331, N4330);
xor XOR2 (N4332, N4329, N2044);
xor XOR2 (N4333, N4322, N3499);
or OR2 (N4334, N4333, N619);
not NOT1 (N4335, N4323);
not NOT1 (N4336, N4327);
or OR2 (N4337, N4325, N546);
nor NOR4 (N4338, N4314, N98, N341, N24);
nor NOR4 (N4339, N4336, N39, N3777, N1465);
not NOT1 (N4340, N4317);
nand NAND4 (N4341, N4321, N3599, N567, N2083);
xor XOR2 (N4342, N4324, N3630);
or OR4 (N4343, N4334, N2947, N1191, N1400);
or OR3 (N4344, N4332, N408, N1064);
or OR4 (N4345, N4341, N2608, N3687, N1264);
or OR4 (N4346, N4335, N2998, N3919, N3933);
not NOT1 (N4347, N4345);
and AND4 (N4348, N4337, N2810, N1070, N247);
not NOT1 (N4349, N4344);
nor NOR4 (N4350, N4347, N1055, N2871, N3258);
xor XOR2 (N4351, N4346, N2931);
and AND4 (N4352, N4340, N3414, N3178, N3616);
buf BUF1 (N4353, N4348);
buf BUF1 (N4354, N4352);
buf BUF1 (N4355, N4338);
buf BUF1 (N4356, N4350);
buf BUF1 (N4357, N4342);
nand NAND2 (N4358, N4349, N51);
nand NAND2 (N4359, N4339, N3229);
buf BUF1 (N4360, N4359);
not NOT1 (N4361, N4331);
nand NAND2 (N4362, N4357, N2874);
and AND4 (N4363, N4355, N3438, N3242, N1206);
nand NAND2 (N4364, N4361, N3831);
and AND3 (N4365, N4358, N4327, N2372);
and AND2 (N4366, N4351, N2274);
nand NAND3 (N4367, N4354, N4065, N1686);
nand NAND3 (N4368, N4360, N4173, N99);
and AND4 (N4369, N4362, N1713, N2446, N2915);
and AND2 (N4370, N4369, N1538);
or OR3 (N4371, N4365, N4041, N2020);
xor XOR2 (N4372, N4364, N2298);
not NOT1 (N4373, N4366);
or OR2 (N4374, N4371, N1647);
xor XOR2 (N4375, N4353, N4079);
nor NOR3 (N4376, N4363, N2389, N2204);
or OR3 (N4377, N4373, N3470, N819);
and AND4 (N4378, N4375, N2605, N2237, N2851);
nor NOR3 (N4379, N4377, N2446, N732);
buf BUF1 (N4380, N4356);
or OR2 (N4381, N4343, N1434);
not NOT1 (N4382, N4372);
nor NOR3 (N4383, N4368, N679, N2644);
nand NAND4 (N4384, N4383, N2468, N755, N906);
not NOT1 (N4385, N4384);
xor XOR2 (N4386, N4381, N1291);
xor XOR2 (N4387, N4380, N1363);
xor XOR2 (N4388, N4382, N873);
xor XOR2 (N4389, N4379, N2863);
nand NAND4 (N4390, N4367, N2047, N2741, N2264);
xor XOR2 (N4391, N4376, N2823);
xor XOR2 (N4392, N4385, N3498);
not NOT1 (N4393, N4390);
nand NAND3 (N4394, N4370, N922, N3447);
not NOT1 (N4395, N4374);
not NOT1 (N4396, N4386);
or OR4 (N4397, N4392, N2079, N797, N4098);
nand NAND2 (N4398, N4394, N957);
and AND3 (N4399, N4398, N1673, N868);
nand NAND3 (N4400, N4395, N3538, N787);
or OR2 (N4401, N4378, N2608);
or OR4 (N4402, N4391, N821, N1893, N2511);
or OR3 (N4403, N4387, N4390, N1045);
xor XOR2 (N4404, N4389, N965);
xor XOR2 (N4405, N4401, N3333);
nor NOR3 (N4406, N4405, N1454, N26);
buf BUF1 (N4407, N4402);
xor XOR2 (N4408, N4400, N1353);
buf BUF1 (N4409, N4404);
and AND4 (N4410, N4397, N37, N3945, N1955);
nor NOR3 (N4411, N4408, N3460, N1952);
and AND2 (N4412, N4409, N1855);
xor XOR2 (N4413, N4410, N1858);
or OR3 (N4414, N4396, N2841, N539);
nand NAND2 (N4415, N4406, N1990);
buf BUF1 (N4416, N4388);
xor XOR2 (N4417, N4403, N2907);
or OR2 (N4418, N4413, N4088);
nand NAND3 (N4419, N4393, N3160, N3638);
xor XOR2 (N4420, N4417, N3424);
and AND3 (N4421, N4414, N84, N342);
not NOT1 (N4422, N4415);
buf BUF1 (N4423, N4411);
xor XOR2 (N4424, N4420, N2848);
nand NAND2 (N4425, N4418, N2081);
xor XOR2 (N4426, N4399, N572);
or OR2 (N4427, N4423, N86);
not NOT1 (N4428, N4421);
not NOT1 (N4429, N4412);
or OR2 (N4430, N4419, N3022);
or OR4 (N4431, N4424, N2578, N2635, N2521);
not NOT1 (N4432, N4428);
not NOT1 (N4433, N4422);
xor XOR2 (N4434, N4416, N3502);
buf BUF1 (N4435, N4430);
xor XOR2 (N4436, N4432, N1745);
nor NOR2 (N4437, N4433, N347);
or OR2 (N4438, N4429, N3422);
or OR4 (N4439, N4426, N2851, N3653, N1652);
xor XOR2 (N4440, N4431, N1390);
and AND3 (N4441, N4436, N2959, N4426);
and AND3 (N4442, N4407, N1999, N1077);
and AND2 (N4443, N4438, N2354);
not NOT1 (N4444, N4441);
nand NAND4 (N4445, N4439, N4443, N399, N3036);
nor NOR4 (N4446, N1421, N116, N4090, N1900);
xor XOR2 (N4447, N4437, N522);
and AND3 (N4448, N4447, N3923, N2953);
nor NOR4 (N4449, N4444, N2108, N1920, N1133);
or OR4 (N4450, N4440, N3248, N37, N1823);
and AND3 (N4451, N4435, N1766, N2263);
xor XOR2 (N4452, N4449, N3016);
buf BUF1 (N4453, N4452);
nor NOR2 (N4454, N4450, N716);
or OR4 (N4455, N4454, N2359, N947, N3578);
buf BUF1 (N4456, N4442);
buf BUF1 (N4457, N4455);
or OR3 (N4458, N4434, N3452, N2461);
nand NAND4 (N4459, N4458, N3271, N2559, N1231);
xor XOR2 (N4460, N4453, N645);
xor XOR2 (N4461, N4448, N1793);
nand NAND4 (N4462, N4446, N724, N51, N1978);
nor NOR3 (N4463, N4461, N768, N4330);
and AND2 (N4464, N4427, N670);
not NOT1 (N4465, N4460);
not NOT1 (N4466, N4445);
buf BUF1 (N4467, N4463);
xor XOR2 (N4468, N4464, N4147);
nor NOR4 (N4469, N4468, N97, N3255, N4161);
xor XOR2 (N4470, N4425, N1561);
nand NAND4 (N4471, N4466, N435, N1377, N2182);
not NOT1 (N4472, N4457);
nand NAND3 (N4473, N4465, N1873, N156);
not NOT1 (N4474, N4470);
not NOT1 (N4475, N4467);
or OR2 (N4476, N4474, N1306);
and AND2 (N4477, N4469, N3070);
nand NAND2 (N4478, N4456, N594);
buf BUF1 (N4479, N4459);
and AND3 (N4480, N4471, N2910, N1780);
buf BUF1 (N4481, N4477);
buf BUF1 (N4482, N4476);
nand NAND3 (N4483, N4462, N489, N281);
nor NOR3 (N4484, N4475, N2391, N2327);
and AND2 (N4485, N4483, N1890);
nand NAND2 (N4486, N4479, N3727);
not NOT1 (N4487, N4485);
and AND4 (N4488, N4473, N3204, N71, N3650);
or OR3 (N4489, N4478, N4162, N2124);
and AND3 (N4490, N4484, N3697, N2371);
nor NOR3 (N4491, N4489, N102, N1674);
or OR2 (N4492, N4482, N3515);
nor NOR2 (N4493, N4487, N390);
buf BUF1 (N4494, N4472);
xor XOR2 (N4495, N4494, N1836);
nand NAND4 (N4496, N4492, N1189, N2361, N3450);
and AND4 (N4497, N4480, N2869, N4336, N3558);
buf BUF1 (N4498, N4495);
xor XOR2 (N4499, N4491, N4391);
buf BUF1 (N4500, N4497);
or OR4 (N4501, N4486, N1547, N1174, N2036);
or OR2 (N4502, N4481, N85);
and AND3 (N4503, N4496, N3585, N1261);
and AND2 (N4504, N4502, N3630);
buf BUF1 (N4505, N4503);
or OR3 (N4506, N4493, N2838, N3890);
nand NAND2 (N4507, N4498, N2768);
nand NAND3 (N4508, N4501, N1653, N1620);
and AND4 (N4509, N4505, N2399, N4336, N2654);
and AND4 (N4510, N4508, N825, N2120, N2542);
or OR4 (N4511, N4488, N710, N1542, N2966);
nand NAND4 (N4512, N4507, N1451, N334, N1186);
nor NOR3 (N4513, N4500, N1049, N4432);
xor XOR2 (N4514, N4490, N2223);
xor XOR2 (N4515, N4511, N409);
or OR4 (N4516, N4513, N2986, N926, N3260);
not NOT1 (N4517, N4515);
or OR4 (N4518, N4516, N406, N3587, N3012);
xor XOR2 (N4519, N4504, N4025);
and AND3 (N4520, N4517, N1776, N4039);
buf BUF1 (N4521, N4519);
buf BUF1 (N4522, N4510);
nor NOR4 (N4523, N4509, N2924, N2050, N2081);
xor XOR2 (N4524, N4499, N1370);
not NOT1 (N4525, N4514);
buf BUF1 (N4526, N4524);
nor NOR3 (N4527, N4451, N3365, N3687);
not NOT1 (N4528, N4506);
buf BUF1 (N4529, N4523);
not NOT1 (N4530, N4527);
xor XOR2 (N4531, N4521, N2436);
not NOT1 (N4532, N4518);
or OR2 (N4533, N4530, N4097);
not NOT1 (N4534, N4531);
nand NAND4 (N4535, N4522, N893, N4136, N2601);
buf BUF1 (N4536, N4535);
nor NOR3 (N4537, N4532, N524, N3253);
nand NAND4 (N4538, N4525, N153, N3903, N2365);
nand NAND4 (N4539, N4512, N2538, N3862, N3509);
buf BUF1 (N4540, N4539);
nor NOR2 (N4541, N4538, N629);
or OR2 (N4542, N4520, N3);
not NOT1 (N4543, N4533);
not NOT1 (N4544, N4541);
buf BUF1 (N4545, N4528);
not NOT1 (N4546, N4529);
xor XOR2 (N4547, N4537, N53);
not NOT1 (N4548, N4540);
and AND2 (N4549, N4547, N2166);
or OR2 (N4550, N4546, N1039);
buf BUF1 (N4551, N4545);
nor NOR2 (N4552, N4534, N3803);
nor NOR4 (N4553, N4552, N950, N2966, N2936);
buf BUF1 (N4554, N4542);
or OR3 (N4555, N4526, N1406, N1097);
not NOT1 (N4556, N4549);
nand NAND4 (N4557, N4548, N105, N1676, N68);
buf BUF1 (N4558, N4544);
nand NAND3 (N4559, N4543, N767, N1200);
or OR4 (N4560, N4558, N2237, N1514, N1885);
buf BUF1 (N4561, N4556);
not NOT1 (N4562, N4550);
and AND3 (N4563, N4557, N3040, N2557);
and AND2 (N4564, N4536, N2026);
nor NOR4 (N4565, N4555, N1150, N3140, N3864);
nand NAND4 (N4566, N4562, N2298, N619, N1427);
nor NOR4 (N4567, N4551, N4245, N588, N691);
xor XOR2 (N4568, N4564, N4538);
buf BUF1 (N4569, N4568);
not NOT1 (N4570, N4553);
xor XOR2 (N4571, N4565, N3826);
buf BUF1 (N4572, N4571);
xor XOR2 (N4573, N4559, N2238);
xor XOR2 (N4574, N4567, N2114);
and AND3 (N4575, N4563, N3287, N2800);
xor XOR2 (N4576, N4573, N2716);
and AND3 (N4577, N4554, N727, N904);
nor NOR4 (N4578, N4566, N3848, N3563, N1920);
not NOT1 (N4579, N4561);
not NOT1 (N4580, N4570);
nand NAND4 (N4581, N4574, N2390, N2666, N2692);
xor XOR2 (N4582, N4577, N1379);
not NOT1 (N4583, N4576);
nor NOR2 (N4584, N4579, N2988);
not NOT1 (N4585, N4583);
or OR2 (N4586, N4578, N3076);
xor XOR2 (N4587, N4560, N1593);
and AND3 (N4588, N4569, N3898, N503);
buf BUF1 (N4589, N4572);
nor NOR2 (N4590, N4575, N563);
and AND2 (N4591, N4588, N2892);
xor XOR2 (N4592, N4581, N2741);
nand NAND3 (N4593, N4589, N1243, N3681);
nand NAND2 (N4594, N4587, N1990);
or OR2 (N4595, N4591, N177);
nor NOR4 (N4596, N4594, N1436, N2033, N1847);
nand NAND2 (N4597, N4593, N3841);
xor XOR2 (N4598, N4585, N925);
not NOT1 (N4599, N4592);
or OR4 (N4600, N4595, N2877, N1119, N4162);
or OR2 (N4601, N4582, N3759);
nor NOR2 (N4602, N4598, N4412);
nor NOR3 (N4603, N4596, N4317, N349);
xor XOR2 (N4604, N4601, N2191);
xor XOR2 (N4605, N4580, N3292);
not NOT1 (N4606, N4597);
not NOT1 (N4607, N4584);
or OR3 (N4608, N4603, N1880, N3301);
xor XOR2 (N4609, N4606, N1534);
or OR2 (N4610, N4599, N1705);
and AND2 (N4611, N4602, N4353);
nor NOR4 (N4612, N4586, N1717, N2993, N3258);
or OR4 (N4613, N4611, N4459, N2039, N3699);
buf BUF1 (N4614, N4613);
nor NOR3 (N4615, N4600, N3253, N3398);
nor NOR2 (N4616, N4612, N1237);
nor NOR3 (N4617, N4605, N3086, N905);
not NOT1 (N4618, N4604);
and AND2 (N4619, N4618, N4528);
nor NOR3 (N4620, N4610, N611, N2250);
buf BUF1 (N4621, N4609);
buf BUF1 (N4622, N4607);
nor NOR2 (N4623, N4608, N3121);
or OR4 (N4624, N4623, N4331, N3348, N4573);
xor XOR2 (N4625, N4616, N3101);
buf BUF1 (N4626, N4617);
and AND2 (N4627, N4625, N2371);
buf BUF1 (N4628, N4620);
not NOT1 (N4629, N4590);
nand NAND4 (N4630, N4614, N2729, N1651, N297);
xor XOR2 (N4631, N4626, N994);
nand NAND3 (N4632, N4631, N2463, N3590);
not NOT1 (N4633, N4624);
nor NOR4 (N4634, N4622, N2297, N3714, N1611);
nand NAND4 (N4635, N4634, N3531, N545, N3307);
not NOT1 (N4636, N4615);
or OR3 (N4637, N4636, N877, N650);
and AND3 (N4638, N4621, N364, N4359);
buf BUF1 (N4639, N4638);
not NOT1 (N4640, N4629);
buf BUF1 (N4641, N4635);
and AND4 (N4642, N4633, N2221, N1946, N925);
and AND4 (N4643, N4619, N109, N2246, N4384);
buf BUF1 (N4644, N4630);
buf BUF1 (N4645, N4632);
or OR4 (N4646, N4643, N3124, N1331, N2668);
not NOT1 (N4647, N4645);
nor NOR4 (N4648, N4647, N4402, N44, N2853);
or OR2 (N4649, N4640, N2093);
buf BUF1 (N4650, N4642);
or OR2 (N4651, N4646, N287);
and AND2 (N4652, N4627, N2647);
xor XOR2 (N4653, N4641, N4218);
not NOT1 (N4654, N4649);
nand NAND4 (N4655, N4628, N790, N1410, N3042);
nor NOR3 (N4656, N4639, N3753, N2707);
nand NAND3 (N4657, N4656, N2520, N508);
xor XOR2 (N4658, N4637, N3998);
nand NAND2 (N4659, N4650, N909);
buf BUF1 (N4660, N4659);
nand NAND3 (N4661, N4654, N3030, N1997);
nor NOR4 (N4662, N4644, N1529, N4398, N782);
or OR2 (N4663, N4652, N2410);
buf BUF1 (N4664, N4653);
not NOT1 (N4665, N4663);
xor XOR2 (N4666, N4648, N2679);
nand NAND2 (N4667, N4664, N3958);
xor XOR2 (N4668, N4657, N2557);
xor XOR2 (N4669, N4667, N1916);
buf BUF1 (N4670, N4660);
nand NAND4 (N4671, N4655, N3263, N1206, N2820);
nor NOR2 (N4672, N4666, N729);
not NOT1 (N4673, N4672);
or OR4 (N4674, N4658, N932, N2621, N2678);
nor NOR3 (N4675, N4661, N2129, N3156);
nand NAND2 (N4676, N4668, N3021);
and AND3 (N4677, N4675, N1362, N3362);
xor XOR2 (N4678, N4651, N3426);
buf BUF1 (N4679, N4677);
not NOT1 (N4680, N4670);
nor NOR4 (N4681, N4673, N2731, N1331, N2706);
nor NOR3 (N4682, N4681, N3070, N963);
nor NOR2 (N4683, N4665, N3047);
not NOT1 (N4684, N4680);
and AND4 (N4685, N4676, N3849, N4308, N2018);
not NOT1 (N4686, N4682);
or OR3 (N4687, N4662, N1902, N2502);
not NOT1 (N4688, N4671);
and AND3 (N4689, N4685, N1178, N4376);
buf BUF1 (N4690, N4689);
and AND2 (N4691, N4683, N3380);
nor NOR3 (N4692, N4690, N2298, N1698);
nor NOR4 (N4693, N4687, N1432, N237, N554);
buf BUF1 (N4694, N4688);
xor XOR2 (N4695, N4669, N1816);
nor NOR2 (N4696, N4674, N352);
xor XOR2 (N4697, N4693, N473);
xor XOR2 (N4698, N4686, N2400);
nand NAND4 (N4699, N4684, N1950, N2986, N2665);
not NOT1 (N4700, N4697);
buf BUF1 (N4701, N4679);
and AND4 (N4702, N4694, N4592, N3368, N2822);
and AND2 (N4703, N4701, N3323);
nand NAND4 (N4704, N4703, N1869, N1625, N3360);
and AND4 (N4705, N4699, N948, N2233, N2268);
and AND4 (N4706, N4700, N260, N3859, N611);
or OR4 (N4707, N4691, N1731, N777, N2490);
buf BUF1 (N4708, N4705);
nand NAND3 (N4709, N4695, N543, N3892);
xor XOR2 (N4710, N4702, N1970);
not NOT1 (N4711, N4704);
not NOT1 (N4712, N4698);
nand NAND4 (N4713, N4712, N4491, N3771, N2268);
nor NOR2 (N4714, N4692, N1988);
nand NAND4 (N4715, N4707, N4213, N4008, N843);
nor NOR4 (N4716, N4714, N58, N3121, N3542);
xor XOR2 (N4717, N4678, N4561);
not NOT1 (N4718, N4715);
nand NAND2 (N4719, N4713, N3346);
not NOT1 (N4720, N4696);
and AND3 (N4721, N4717, N3423, N2524);
nand NAND4 (N4722, N4716, N1552, N418, N3469);
xor XOR2 (N4723, N4708, N1059);
nor NOR2 (N4724, N4706, N738);
or OR3 (N4725, N4722, N1516, N262);
buf BUF1 (N4726, N4718);
nor NOR4 (N4727, N4726, N4540, N1426, N3891);
nor NOR4 (N4728, N4727, N1627, N154, N3975);
xor XOR2 (N4729, N4719, N3772);
or OR2 (N4730, N4721, N3608);
xor XOR2 (N4731, N4730, N2260);
nand NAND2 (N4732, N4725, N1026);
not NOT1 (N4733, N4723);
xor XOR2 (N4734, N4733, N4243);
buf BUF1 (N4735, N4731);
not NOT1 (N4736, N4729);
not NOT1 (N4737, N4710);
or OR4 (N4738, N4711, N1563, N1327, N2777);
xor XOR2 (N4739, N4724, N269);
nor NOR4 (N4740, N4732, N522, N2647, N778);
nor NOR2 (N4741, N4739, N3424);
not NOT1 (N4742, N4720);
nand NAND2 (N4743, N4740, N307);
and AND4 (N4744, N4742, N1346, N1030, N1141);
and AND2 (N4745, N4709, N1401);
nor NOR2 (N4746, N4744, N194);
not NOT1 (N4747, N4734);
buf BUF1 (N4748, N4728);
not NOT1 (N4749, N4741);
and AND4 (N4750, N4749, N103, N2882, N1969);
nand NAND2 (N4751, N4743, N2200);
nand NAND4 (N4752, N4747, N200, N4011, N2988);
xor XOR2 (N4753, N4750, N3428);
buf BUF1 (N4754, N4753);
not NOT1 (N4755, N4751);
and AND4 (N4756, N4748, N1305, N3861, N4244);
not NOT1 (N4757, N4756);
nand NAND4 (N4758, N4735, N3714, N1949, N1549);
or OR3 (N4759, N4736, N3242, N1010);
nand NAND4 (N4760, N4759, N3581, N3923, N1092);
not NOT1 (N4761, N4738);
or OR4 (N4762, N4754, N4101, N4671, N2473);
nand NAND2 (N4763, N4745, N4327);
buf BUF1 (N4764, N4762);
buf BUF1 (N4765, N4763);
or OR3 (N4766, N4765, N2610, N1937);
xor XOR2 (N4767, N4760, N3632);
not NOT1 (N4768, N4764);
nor NOR3 (N4769, N4768, N1068, N3867);
and AND3 (N4770, N4767, N4170, N4379);
and AND4 (N4771, N4746, N1101, N2002, N1720);
xor XOR2 (N4772, N4771, N4664);
nor NOR4 (N4773, N4737, N3928, N2981, N759);
nor NOR3 (N4774, N4770, N4707, N1407);
not NOT1 (N4775, N4769);
nand NAND2 (N4776, N4773, N4036);
not NOT1 (N4777, N4755);
and AND3 (N4778, N4757, N2065, N3125);
nor NOR2 (N4779, N4761, N3764);
not NOT1 (N4780, N4758);
not NOT1 (N4781, N4775);
nand NAND2 (N4782, N4766, N609);
and AND2 (N4783, N4752, N4497);
nand NAND2 (N4784, N4778, N788);
not NOT1 (N4785, N4781);
and AND2 (N4786, N4784, N489);
nand NAND2 (N4787, N4783, N606);
nor NOR4 (N4788, N4772, N399, N4177, N3176);
buf BUF1 (N4789, N4785);
not NOT1 (N4790, N4776);
xor XOR2 (N4791, N4789, N3776);
xor XOR2 (N4792, N4779, N2928);
or OR4 (N4793, N4786, N1014, N639, N2767);
nand NAND3 (N4794, N4780, N2648, N892);
nand NAND2 (N4795, N4774, N253);
buf BUF1 (N4796, N4795);
and AND3 (N4797, N4790, N2959, N1035);
nor NOR3 (N4798, N4794, N3044, N2185);
and AND2 (N4799, N4797, N978);
or OR4 (N4800, N4798, N639, N4693, N3445);
buf BUF1 (N4801, N4787);
or OR3 (N4802, N4791, N3135, N904);
xor XOR2 (N4803, N4802, N4343);
not NOT1 (N4804, N4801);
xor XOR2 (N4805, N4796, N2755);
and AND2 (N4806, N4782, N135);
and AND2 (N4807, N4777, N1188);
and AND2 (N4808, N4792, N193);
nand NAND3 (N4809, N4793, N1377, N4210);
not NOT1 (N4810, N4805);
not NOT1 (N4811, N4808);
and AND4 (N4812, N4803, N2430, N4272, N4329);
not NOT1 (N4813, N4806);
not NOT1 (N4814, N4800);
buf BUF1 (N4815, N4814);
buf BUF1 (N4816, N4809);
and AND4 (N4817, N4807, N805, N4698, N764);
not NOT1 (N4818, N4817);
nor NOR3 (N4819, N4818, N403, N134);
buf BUF1 (N4820, N4804);
not NOT1 (N4821, N4788);
not NOT1 (N4822, N4810);
buf BUF1 (N4823, N4799);
xor XOR2 (N4824, N4815, N4133);
buf BUF1 (N4825, N4813);
nor NOR3 (N4826, N4819, N939, N314);
xor XOR2 (N4827, N4816, N2098);
buf BUF1 (N4828, N4812);
xor XOR2 (N4829, N4826, N1436);
xor XOR2 (N4830, N4829, N180);
nor NOR4 (N4831, N4824, N4233, N845, N1985);
nand NAND4 (N4832, N4822, N247, N2946, N1796);
or OR4 (N4833, N4832, N3581, N4767, N2405);
nand NAND4 (N4834, N4827, N223, N1401, N3398);
buf BUF1 (N4835, N4833);
xor XOR2 (N4836, N4828, N3442);
buf BUF1 (N4837, N4835);
not NOT1 (N4838, N4831);
or OR3 (N4839, N4837, N221, N4173);
and AND3 (N4840, N4820, N1344, N3431);
nand NAND4 (N4841, N4830, N3791, N793, N1082);
nand NAND2 (N4842, N4840, N4205);
not NOT1 (N4843, N4838);
not NOT1 (N4844, N4821);
buf BUF1 (N4845, N4839);
and AND4 (N4846, N4834, N2709, N2673, N2604);
nor NOR2 (N4847, N4836, N4493);
not NOT1 (N4848, N4846);
and AND3 (N4849, N4843, N1058, N4450);
xor XOR2 (N4850, N4847, N3654);
buf BUF1 (N4851, N4845);
xor XOR2 (N4852, N4841, N3938);
nand NAND2 (N4853, N4850, N1582);
buf BUF1 (N4854, N4853);
xor XOR2 (N4855, N4848, N3330);
buf BUF1 (N4856, N4852);
or OR4 (N4857, N4856, N4635, N1566, N4605);
and AND3 (N4858, N4849, N611, N585);
or OR4 (N4859, N4854, N2231, N4196, N4431);
buf BUF1 (N4860, N4842);
or OR2 (N4861, N4825, N3765);
or OR3 (N4862, N4844, N397, N574);
not NOT1 (N4863, N4855);
nand NAND2 (N4864, N4851, N857);
or OR2 (N4865, N4811, N2149);
nand NAND3 (N4866, N4857, N2361, N2013);
xor XOR2 (N4867, N4864, N1349);
and AND4 (N4868, N4866, N404, N3548, N280);
not NOT1 (N4869, N4862);
or OR4 (N4870, N4869, N1971, N546, N4635);
buf BUF1 (N4871, N4861);
and AND2 (N4872, N4823, N4173);
not NOT1 (N4873, N4871);
xor XOR2 (N4874, N4870, N4209);
nor NOR2 (N4875, N4860, N4001);
or OR3 (N4876, N4868, N4024, N3709);
buf BUF1 (N4877, N4865);
nor NOR4 (N4878, N4872, N3892, N4296, N790);
and AND2 (N4879, N4874, N3566);
buf BUF1 (N4880, N4863);
nor NOR2 (N4881, N4875, N1909);
and AND3 (N4882, N4876, N3206, N4764);
nand NAND4 (N4883, N4877, N321, N3563, N193);
xor XOR2 (N4884, N4882, N725);
xor XOR2 (N4885, N4878, N3482);
xor XOR2 (N4886, N4881, N1329);
or OR2 (N4887, N4886, N3293);
nand NAND2 (N4888, N4884, N1758);
and AND4 (N4889, N4867, N4321, N1006, N1220);
buf BUF1 (N4890, N4873);
buf BUF1 (N4891, N4887);
and AND4 (N4892, N4880, N3499, N4161, N754);
nor NOR4 (N4893, N4888, N447, N696, N4779);
nand NAND2 (N4894, N4885, N783);
and AND4 (N4895, N4883, N3107, N2591, N1066);
nand NAND4 (N4896, N4890, N1627, N4451, N2238);
and AND2 (N4897, N4892, N3927);
xor XOR2 (N4898, N4858, N1738);
buf BUF1 (N4899, N4859);
or OR4 (N4900, N4893, N3002, N4217, N4251);
not NOT1 (N4901, N4879);
and AND2 (N4902, N4889, N2974);
or OR2 (N4903, N4899, N1151);
xor XOR2 (N4904, N4901, N4348);
nand NAND4 (N4905, N4895, N2671, N4207, N2842);
xor XOR2 (N4906, N4904, N1506);
nor NOR4 (N4907, N4894, N446, N728, N3468);
nor NOR3 (N4908, N4903, N2809, N87);
xor XOR2 (N4909, N4905, N4420);
nand NAND3 (N4910, N4897, N4127, N4592);
xor XOR2 (N4911, N4908, N3645);
xor XOR2 (N4912, N4910, N4757);
or OR4 (N4913, N4911, N2694, N4739, N3966);
nand NAND3 (N4914, N4900, N3608, N2323);
nor NOR2 (N4915, N4914, N1542);
or OR4 (N4916, N4898, N4581, N1033, N1156);
not NOT1 (N4917, N4909);
not NOT1 (N4918, N4891);
nand NAND3 (N4919, N4906, N680, N1781);
nand NAND3 (N4920, N4917, N4608, N4838);
not NOT1 (N4921, N4912);
and AND4 (N4922, N4902, N54, N4342, N1254);
nand NAND3 (N4923, N4918, N3180, N2747);
not NOT1 (N4924, N4896);
nor NOR4 (N4925, N4907, N404, N634, N2870);
and AND3 (N4926, N4919, N3459, N3162);
buf BUF1 (N4927, N4925);
or OR2 (N4928, N4920, N171);
and AND2 (N4929, N4923, N410);
nor NOR2 (N4930, N4926, N4494);
nor NOR3 (N4931, N4915, N1615, N4490);
not NOT1 (N4932, N4928);
not NOT1 (N4933, N4929);
xor XOR2 (N4934, N4916, N260);
not NOT1 (N4935, N4924);
nor NOR2 (N4936, N4921, N2289);
nand NAND3 (N4937, N4933, N2238, N193);
xor XOR2 (N4938, N4913, N145);
nor NOR2 (N4939, N4936, N1245);
nand NAND3 (N4940, N4932, N1103, N889);
and AND4 (N4941, N4940, N4446, N1351, N3400);
nand NAND2 (N4942, N4927, N4727);
buf BUF1 (N4943, N4935);
nand NAND2 (N4944, N4934, N1623);
not NOT1 (N4945, N4941);
buf BUF1 (N4946, N4942);
buf BUF1 (N4947, N4938);
xor XOR2 (N4948, N4937, N1779);
or OR4 (N4949, N4931, N3277, N3932, N248);
and AND2 (N4950, N4949, N3931);
xor XOR2 (N4951, N4950, N1995);
xor XOR2 (N4952, N4943, N935);
buf BUF1 (N4953, N4939);
or OR2 (N4954, N4944, N2522);
xor XOR2 (N4955, N4948, N4681);
or OR2 (N4956, N4954, N4602);
buf BUF1 (N4957, N4946);
not NOT1 (N4958, N4947);
and AND3 (N4959, N4951, N3596, N878);
and AND2 (N4960, N4957, N1197);
xor XOR2 (N4961, N4958, N1810);
or OR3 (N4962, N4922, N2467, N356);
buf BUF1 (N4963, N4956);
or OR2 (N4964, N4963, N3259);
or OR3 (N4965, N4955, N720, N1167);
or OR3 (N4966, N4953, N4545, N3451);
not NOT1 (N4967, N4945);
and AND3 (N4968, N4960, N1465, N1279);
xor XOR2 (N4969, N4962, N4874);
nand NAND2 (N4970, N4930, N4548);
and AND3 (N4971, N4967, N4013, N3050);
and AND4 (N4972, N4970, N4558, N4097, N4941);
and AND4 (N4973, N4968, N3531, N3970, N4161);
buf BUF1 (N4974, N4952);
or OR4 (N4975, N4961, N201, N454, N1899);
xor XOR2 (N4976, N4965, N3365);
buf BUF1 (N4977, N4964);
buf BUF1 (N4978, N4977);
not NOT1 (N4979, N4975);
nand NAND3 (N4980, N4972, N4261, N3109);
buf BUF1 (N4981, N4979);
not NOT1 (N4982, N4980);
or OR2 (N4983, N4982, N226);
not NOT1 (N4984, N4973);
not NOT1 (N4985, N4969);
xor XOR2 (N4986, N4983, N4059);
nor NOR2 (N4987, N4974, N4694);
not NOT1 (N4988, N4966);
xor XOR2 (N4989, N4986, N4390);
nor NOR3 (N4990, N4971, N1587, N3226);
buf BUF1 (N4991, N4990);
xor XOR2 (N4992, N4976, N853);
nor NOR3 (N4993, N4989, N3564, N441);
or OR3 (N4994, N4992, N1584, N203);
nor NOR3 (N4995, N4978, N1066, N3004);
nor NOR3 (N4996, N4994, N2050, N505);
nand NAND4 (N4997, N4995, N4515, N929, N80);
xor XOR2 (N4998, N4993, N1520);
nor NOR3 (N4999, N4984, N1864, N141);
nand NAND2 (N5000, N4987, N1576);
and AND3 (N5001, N4998, N1570, N4436);
buf BUF1 (N5002, N4988);
not NOT1 (N5003, N4991);
not NOT1 (N5004, N4985);
xor XOR2 (N5005, N5002, N4833);
not NOT1 (N5006, N5005);
or OR4 (N5007, N5000, N631, N3204, N1511);
nand NAND4 (N5008, N4999, N3797, N977, N3726);
and AND4 (N5009, N5003, N1895, N3613, N2677);
nand NAND2 (N5010, N4959, N4404);
or OR4 (N5011, N5001, N1216, N3852, N2144);
not NOT1 (N5012, N4996);
nor NOR2 (N5013, N5006, N1217);
and AND2 (N5014, N5007, N1271);
and AND4 (N5015, N5012, N2615, N1298, N1822);
buf BUF1 (N5016, N5013);
and AND3 (N5017, N4997, N2006, N3335);
nor NOR3 (N5018, N4981, N2202, N3303);
nand NAND2 (N5019, N5008, N3962);
and AND3 (N5020, N5004, N4628, N4289);
or OR2 (N5021, N5014, N3628);
buf BUF1 (N5022, N5020);
buf BUF1 (N5023, N5019);
not NOT1 (N5024, N5009);
not NOT1 (N5025, N5018);
nand NAND3 (N5026, N5021, N1057, N3043);
nor NOR4 (N5027, N5016, N4239, N2993, N2535);
and AND3 (N5028, N5022, N4433, N1774);
xor XOR2 (N5029, N5017, N947);
not NOT1 (N5030, N5024);
or OR3 (N5031, N5026, N2748, N4879);
buf BUF1 (N5032, N5015);
xor XOR2 (N5033, N5028, N4859);
xor XOR2 (N5034, N5032, N3545);
or OR3 (N5035, N5023, N2163, N4860);
or OR3 (N5036, N5011, N2442, N3778);
nand NAND4 (N5037, N5027, N1685, N1127, N2576);
nor NOR2 (N5038, N5033, N4486);
and AND3 (N5039, N5030, N4011, N2190);
xor XOR2 (N5040, N5034, N2785);
buf BUF1 (N5041, N5035);
not NOT1 (N5042, N5025);
not NOT1 (N5043, N5042);
buf BUF1 (N5044, N5038);
nand NAND2 (N5045, N5029, N3259);
xor XOR2 (N5046, N5045, N180);
nand NAND2 (N5047, N5010, N2737);
xor XOR2 (N5048, N5046, N3970);
xor XOR2 (N5049, N5047, N4555);
nand NAND3 (N5050, N5036, N838, N4124);
not NOT1 (N5051, N5041);
not NOT1 (N5052, N5037);
nor NOR4 (N5053, N5039, N3308, N4842, N4270);
not NOT1 (N5054, N5048);
nand NAND2 (N5055, N5049, N640);
buf BUF1 (N5056, N5050);
not NOT1 (N5057, N5054);
or OR4 (N5058, N5031, N4742, N1535, N3347);
and AND4 (N5059, N5053, N4450, N3253, N4641);
or OR3 (N5060, N5044, N4126, N2350);
xor XOR2 (N5061, N5059, N1106);
xor XOR2 (N5062, N5061, N4982);
and AND3 (N5063, N5052, N1006, N4279);
buf BUF1 (N5064, N5060);
not NOT1 (N5065, N5051);
and AND3 (N5066, N5058, N2006, N3899);
nand NAND3 (N5067, N5040, N2133, N2438);
xor XOR2 (N5068, N5055, N1734);
xor XOR2 (N5069, N5066, N1414);
buf BUF1 (N5070, N5065);
and AND4 (N5071, N5062, N1407, N1142, N4691);
and AND4 (N5072, N5043, N1205, N4365, N882);
not NOT1 (N5073, N5063);
not NOT1 (N5074, N5056);
xor XOR2 (N5075, N5069, N2629);
nor NOR3 (N5076, N5072, N4012, N2936);
buf BUF1 (N5077, N5076);
buf BUF1 (N5078, N5074);
nand NAND3 (N5079, N5070, N3379, N2208);
nand NAND4 (N5080, N5078, N2116, N3622, N1070);
buf BUF1 (N5081, N5077);
and AND2 (N5082, N5080, N4033);
or OR3 (N5083, N5068, N1025, N1071);
or OR3 (N5084, N5073, N4057, N2312);
or OR3 (N5085, N5082, N3223, N1487);
buf BUF1 (N5086, N5081);
or OR3 (N5087, N5084, N3907, N5064);
buf BUF1 (N5088, N4502);
nand NAND3 (N5089, N5067, N2860, N5055);
or OR2 (N5090, N5083, N2778);
nor NOR2 (N5091, N5086, N5000);
not NOT1 (N5092, N5075);
and AND2 (N5093, N5088, N4691);
not NOT1 (N5094, N5093);
xor XOR2 (N5095, N5092, N3257);
not NOT1 (N5096, N5091);
buf BUF1 (N5097, N5079);
nand NAND4 (N5098, N5089, N1147, N3099, N4459);
xor XOR2 (N5099, N5071, N2007);
buf BUF1 (N5100, N5097);
buf BUF1 (N5101, N5099);
and AND3 (N5102, N5087, N4890, N3663);
or OR2 (N5103, N5085, N5096);
not NOT1 (N5104, N3421);
nand NAND2 (N5105, N5104, N2836);
and AND2 (N5106, N5100, N3586);
xor XOR2 (N5107, N5106, N953);
or OR3 (N5108, N5057, N3506, N38);
and AND2 (N5109, N5094, N733);
nand NAND2 (N5110, N5102, N4316);
or OR3 (N5111, N5101, N103, N886);
and AND4 (N5112, N5105, N1444, N2348, N4286);
or OR3 (N5113, N5110, N709, N4447);
or OR3 (N5114, N5113, N369, N886);
not NOT1 (N5115, N5098);
not NOT1 (N5116, N5103);
nor NOR4 (N5117, N5107, N4189, N3077, N274);
nand NAND2 (N5118, N5114, N127);
nand NAND4 (N5119, N5095, N3686, N1084, N1896);
nor NOR3 (N5120, N5109, N1996, N3156);
not NOT1 (N5121, N5116);
or OR4 (N5122, N5120, N3230, N4071, N2709);
nor NOR3 (N5123, N5090, N1013, N4476);
not NOT1 (N5124, N5122);
or OR3 (N5125, N5111, N4118, N4750);
not NOT1 (N5126, N5112);
or OR2 (N5127, N5126, N3854);
buf BUF1 (N5128, N5117);
nor NOR4 (N5129, N5115, N3302, N2265, N1931);
xor XOR2 (N5130, N5119, N1900);
nand NAND2 (N5131, N5125, N459);
buf BUF1 (N5132, N5121);
nor NOR4 (N5133, N5108, N1728, N1394, N5064);
xor XOR2 (N5134, N5131, N3813);
or OR4 (N5135, N5132, N3013, N4238, N3424);
not NOT1 (N5136, N5133);
not NOT1 (N5137, N5130);
nand NAND4 (N5138, N5124, N1135, N2235, N5025);
or OR4 (N5139, N5128, N4737, N4888, N4801);
nor NOR2 (N5140, N5127, N3136);
nor NOR2 (N5141, N5136, N889);
nor NOR4 (N5142, N5139, N5062, N3946, N3058);
nor NOR2 (N5143, N5138, N868);
not NOT1 (N5144, N5140);
nor NOR4 (N5145, N5141, N2620, N1018, N3288);
buf BUF1 (N5146, N5145);
and AND2 (N5147, N5137, N1209);
xor XOR2 (N5148, N5118, N1560);
buf BUF1 (N5149, N5129);
and AND4 (N5150, N5149, N3637, N3251, N2718);
not NOT1 (N5151, N5146);
nor NOR4 (N5152, N5150, N1753, N713, N2403);
buf BUF1 (N5153, N5151);
nor NOR2 (N5154, N5148, N181);
buf BUF1 (N5155, N5123);
nand NAND3 (N5156, N5154, N4989, N3761);
not NOT1 (N5157, N5153);
buf BUF1 (N5158, N5157);
or OR3 (N5159, N5147, N2919, N2533);
or OR3 (N5160, N5142, N1607, N3220);
and AND3 (N5161, N5135, N1850, N4264);
xor XOR2 (N5162, N5155, N1696);
buf BUF1 (N5163, N5160);
buf BUF1 (N5164, N5158);
and AND3 (N5165, N5162, N4210, N1780);
and AND2 (N5166, N5164, N142);
or OR3 (N5167, N5166, N3626, N3568);
or OR2 (N5168, N5144, N4411);
xor XOR2 (N5169, N5156, N4280);
and AND2 (N5170, N5165, N2151);
not NOT1 (N5171, N5167);
and AND2 (N5172, N5171, N2683);
not NOT1 (N5173, N5143);
or OR2 (N5174, N5159, N2147);
or OR2 (N5175, N5134, N1581);
and AND3 (N5176, N5170, N866, N1660);
or OR2 (N5177, N5152, N5004);
xor XOR2 (N5178, N5172, N385);
or OR3 (N5179, N5178, N2294, N3494);
or OR3 (N5180, N5169, N3597, N788);
and AND2 (N5181, N5180, N722);
nor NOR4 (N5182, N5161, N2439, N732, N4289);
buf BUF1 (N5183, N5174);
xor XOR2 (N5184, N5179, N1357);
nand NAND3 (N5185, N5163, N87, N376);
and AND3 (N5186, N5176, N1292, N1457);
or OR4 (N5187, N5168, N4900, N1117, N716);
xor XOR2 (N5188, N5186, N3341);
xor XOR2 (N5189, N5183, N4635);
buf BUF1 (N5190, N5177);
or OR4 (N5191, N5184, N2828, N185, N516);
nor NOR3 (N5192, N5175, N1873, N1162);
nor NOR3 (N5193, N5187, N2089, N2723);
xor XOR2 (N5194, N5182, N1705);
buf BUF1 (N5195, N5190);
nand NAND4 (N5196, N5192, N4093, N3162, N4629);
and AND3 (N5197, N5188, N4337, N1335);
or OR2 (N5198, N5197, N2140);
and AND2 (N5199, N5181, N225);
and AND4 (N5200, N5194, N1552, N4880, N2546);
not NOT1 (N5201, N5198);
or OR2 (N5202, N5200, N2479);
xor XOR2 (N5203, N5202, N1891);
xor XOR2 (N5204, N5199, N1151);
not NOT1 (N5205, N5173);
nand NAND3 (N5206, N5196, N3986, N455);
xor XOR2 (N5207, N5185, N224);
nor NOR3 (N5208, N5207, N3134, N1151);
and AND3 (N5209, N5206, N3139, N4295);
buf BUF1 (N5210, N5205);
or OR3 (N5211, N5210, N315, N2951);
and AND2 (N5212, N5195, N3275);
or OR3 (N5213, N5191, N3917, N3534);
xor XOR2 (N5214, N5213, N3922);
xor XOR2 (N5215, N5204, N1213);
buf BUF1 (N5216, N5201);
buf BUF1 (N5217, N5203);
nor NOR4 (N5218, N5216, N3262, N1225, N210);
xor XOR2 (N5219, N5208, N1343);
nand NAND2 (N5220, N5209, N990);
buf BUF1 (N5221, N5189);
not NOT1 (N5222, N5215);
nand NAND3 (N5223, N5211, N5011, N3271);
nand NAND4 (N5224, N5218, N4245, N2145, N152);
not NOT1 (N5225, N5220);
xor XOR2 (N5226, N5223, N5039);
nor NOR3 (N5227, N5193, N3108, N1146);
buf BUF1 (N5228, N5212);
nand NAND4 (N5229, N5228, N934, N3029, N419);
and AND3 (N5230, N5225, N619, N3779);
nand NAND3 (N5231, N5222, N3358, N5165);
or OR4 (N5232, N5230, N1577, N2791, N4115);
not NOT1 (N5233, N5221);
nand NAND4 (N5234, N5214, N364, N837, N4167);
or OR2 (N5235, N5224, N4307);
nand NAND2 (N5236, N5231, N3778);
xor XOR2 (N5237, N5233, N3405);
buf BUF1 (N5238, N5229);
buf BUF1 (N5239, N5234);
nand NAND4 (N5240, N5236, N1628, N1619, N2627);
or OR2 (N5241, N5238, N4614);
buf BUF1 (N5242, N5239);
not NOT1 (N5243, N5232);
nand NAND4 (N5244, N5227, N2531, N4015, N1866);
or OR2 (N5245, N5240, N63);
nand NAND3 (N5246, N5245, N3956, N187);
and AND2 (N5247, N5242, N787);
and AND3 (N5248, N5235, N1314, N1818);
nor NOR4 (N5249, N5244, N2580, N2135, N2705);
and AND3 (N5250, N5246, N4023, N1745);
nand NAND2 (N5251, N5237, N1783);
xor XOR2 (N5252, N5247, N1677);
buf BUF1 (N5253, N5217);
xor XOR2 (N5254, N5226, N4749);
nand NAND3 (N5255, N5250, N1899, N4252);
nor NOR3 (N5256, N5249, N5145, N3407);
nor NOR3 (N5257, N5256, N1232, N892);
nand NAND3 (N5258, N5251, N2724, N125);
and AND2 (N5259, N5253, N5239);
nor NOR3 (N5260, N5257, N282, N4653);
nand NAND2 (N5261, N5248, N3074);
buf BUF1 (N5262, N5255);
or OR2 (N5263, N5258, N9);
nor NOR2 (N5264, N5259, N4922);
buf BUF1 (N5265, N5264);
buf BUF1 (N5266, N5254);
or OR2 (N5267, N5263, N1202);
or OR4 (N5268, N5260, N3252, N3842, N3794);
xor XOR2 (N5269, N5219, N1026);
buf BUF1 (N5270, N5261);
not NOT1 (N5271, N5269);
not NOT1 (N5272, N5252);
xor XOR2 (N5273, N5267, N4579);
xor XOR2 (N5274, N5241, N29);
and AND4 (N5275, N5270, N4721, N876, N112);
and AND4 (N5276, N5275, N3275, N4965, N4346);
xor XOR2 (N5277, N5262, N4200);
buf BUF1 (N5278, N5272);
xor XOR2 (N5279, N5268, N4007);
buf BUF1 (N5280, N5279);
nor NOR3 (N5281, N5266, N1960, N116);
and AND3 (N5282, N5243, N3530, N5005);
nand NAND3 (N5283, N5276, N2413, N463);
buf BUF1 (N5284, N5277);
nand NAND3 (N5285, N5281, N5150, N1052);
or OR2 (N5286, N5280, N3580);
xor XOR2 (N5287, N5284, N994);
nand NAND4 (N5288, N5278, N2822, N4489, N405);
not NOT1 (N5289, N5273);
and AND2 (N5290, N5271, N5141);
buf BUF1 (N5291, N5283);
nand NAND2 (N5292, N5282, N845);
not NOT1 (N5293, N5292);
buf BUF1 (N5294, N5274);
not NOT1 (N5295, N5265);
not NOT1 (N5296, N5291);
and AND3 (N5297, N5286, N1721, N3080);
nand NAND2 (N5298, N5285, N3952);
nor NOR2 (N5299, N5289, N1915);
nor NOR2 (N5300, N5295, N741);
and AND2 (N5301, N5300, N537);
nand NAND2 (N5302, N5299, N5111);
or OR4 (N5303, N5293, N421, N5062, N5229);
not NOT1 (N5304, N5296);
or OR3 (N5305, N5301, N3855, N3473);
nand NAND2 (N5306, N5298, N2275);
or OR2 (N5307, N5297, N1386);
not NOT1 (N5308, N5304);
or OR3 (N5309, N5290, N218, N1771);
not NOT1 (N5310, N5288);
nor NOR4 (N5311, N5309, N1226, N1039, N1482);
or OR2 (N5312, N5310, N3832);
nand NAND4 (N5313, N5307, N1182, N556, N883);
xor XOR2 (N5314, N5294, N3495);
not NOT1 (N5315, N5314);
buf BUF1 (N5316, N5305);
not NOT1 (N5317, N5308);
xor XOR2 (N5318, N5312, N5288);
nand NAND4 (N5319, N5287, N4056, N2043, N297);
nand NAND3 (N5320, N5319, N1137, N18);
not NOT1 (N5321, N5318);
xor XOR2 (N5322, N5316, N830);
and AND4 (N5323, N5321, N4946, N1061, N25);
xor XOR2 (N5324, N5315, N4355);
nand NAND3 (N5325, N5306, N1556, N231);
not NOT1 (N5326, N5311);
not NOT1 (N5327, N5317);
nand NAND3 (N5328, N5313, N1505, N2895);
and AND2 (N5329, N5327, N1413);
nor NOR4 (N5330, N5320, N63, N5218, N3537);
and AND3 (N5331, N5328, N3986, N4303);
buf BUF1 (N5332, N5302);
nand NAND3 (N5333, N5324, N3472, N4128);
xor XOR2 (N5334, N5323, N4869);
not NOT1 (N5335, N5303);
buf BUF1 (N5336, N5331);
or OR4 (N5337, N5325, N5182, N4995, N674);
not NOT1 (N5338, N5322);
or OR4 (N5339, N5338, N858, N664, N2607);
not NOT1 (N5340, N5326);
not NOT1 (N5341, N5333);
and AND3 (N5342, N5341, N3049, N833);
nor NOR2 (N5343, N5332, N4851);
buf BUF1 (N5344, N5336);
nand NAND4 (N5345, N5339, N3660, N2093, N5066);
buf BUF1 (N5346, N5343);
nor NOR3 (N5347, N5335, N1564, N4703);
or OR4 (N5348, N5330, N3241, N1216, N2257);
or OR2 (N5349, N5337, N4602);
xor XOR2 (N5350, N5342, N2206);
and AND3 (N5351, N5348, N4231, N3766);
nor NOR2 (N5352, N5340, N2559);
nor NOR3 (N5353, N5351, N4975, N4621);
not NOT1 (N5354, N5334);
nand NAND3 (N5355, N5346, N2381, N3645);
buf BUF1 (N5356, N5345);
xor XOR2 (N5357, N5347, N3628);
xor XOR2 (N5358, N5349, N5250);
nor NOR2 (N5359, N5350, N4349);
buf BUF1 (N5360, N5359);
nor NOR3 (N5361, N5352, N1019, N5257);
xor XOR2 (N5362, N5344, N2019);
xor XOR2 (N5363, N5329, N2523);
and AND2 (N5364, N5361, N3946);
nand NAND3 (N5365, N5364, N4380, N2469);
xor XOR2 (N5366, N5353, N1690);
xor XOR2 (N5367, N5356, N1913);
xor XOR2 (N5368, N5365, N3678);
buf BUF1 (N5369, N5358);
nand NAND2 (N5370, N5368, N1426);
nand NAND3 (N5371, N5367, N5179, N544);
not NOT1 (N5372, N5371);
nor NOR2 (N5373, N5357, N4524);
xor XOR2 (N5374, N5372, N4378);
not NOT1 (N5375, N5370);
buf BUF1 (N5376, N5354);
not NOT1 (N5377, N5360);
or OR2 (N5378, N5355, N2100);
and AND3 (N5379, N5362, N4815, N4232);
or OR4 (N5380, N5378, N1851, N1105, N529);
or OR4 (N5381, N5363, N2251, N3294, N1223);
not NOT1 (N5382, N5381);
or OR4 (N5383, N5376, N2408, N3912, N2952);
nand NAND2 (N5384, N5383, N4589);
or OR4 (N5385, N5380, N4197, N2139, N1029);
not NOT1 (N5386, N5382);
buf BUF1 (N5387, N5373);
or OR2 (N5388, N5377, N481);
and AND3 (N5389, N5366, N4481, N2472);
and AND4 (N5390, N5369, N2413, N1374, N921);
and AND2 (N5391, N5375, N2680);
buf BUF1 (N5392, N5386);
xor XOR2 (N5393, N5384, N1103);
xor XOR2 (N5394, N5374, N1684);
nor NOR4 (N5395, N5388, N424, N692, N5307);
and AND2 (N5396, N5385, N1549);
buf BUF1 (N5397, N5390);
not NOT1 (N5398, N5387);
nand NAND2 (N5399, N5394, N2707);
and AND4 (N5400, N5398, N1291, N3937, N2626);
xor XOR2 (N5401, N5400, N4139);
and AND4 (N5402, N5379, N2083, N1899, N2526);
not NOT1 (N5403, N5391);
or OR3 (N5404, N5399, N3360, N1368);
nor NOR4 (N5405, N5392, N3687, N4378, N1071);
nand NAND3 (N5406, N5403, N1401, N3079);
nor NOR2 (N5407, N5401, N1366);
nand NAND2 (N5408, N5407, N1380);
or OR2 (N5409, N5408, N3613);
and AND2 (N5410, N5402, N4250);
nor NOR2 (N5411, N5396, N1123);
xor XOR2 (N5412, N5395, N3796);
or OR2 (N5413, N5397, N2006);
buf BUF1 (N5414, N5406);
or OR3 (N5415, N5411, N5160, N2767);
xor XOR2 (N5416, N5410, N3989);
or OR3 (N5417, N5415, N5374, N610);
nand NAND4 (N5418, N5393, N1030, N3158, N2770);
and AND2 (N5419, N5409, N1813);
xor XOR2 (N5420, N5419, N1911);
or OR2 (N5421, N5418, N12);
nand NAND4 (N5422, N5412, N2707, N3855, N5364);
xor XOR2 (N5423, N5421, N5413);
and AND4 (N5424, N3441, N4012, N4648, N4284);
nand NAND2 (N5425, N5423, N5140);
not NOT1 (N5426, N5414);
and AND2 (N5427, N5425, N4794);
and AND3 (N5428, N5389, N2800, N3485);
nand NAND3 (N5429, N5416, N4738, N4198);
buf BUF1 (N5430, N5404);
nand NAND4 (N5431, N5430, N1934, N2230, N2481);
not NOT1 (N5432, N5428);
not NOT1 (N5433, N5431);
and AND2 (N5434, N5429, N2309);
xor XOR2 (N5435, N5424, N4877);
not NOT1 (N5436, N5405);
and AND2 (N5437, N5436, N682);
xor XOR2 (N5438, N5417, N2168);
and AND2 (N5439, N5438, N1048);
not NOT1 (N5440, N5437);
xor XOR2 (N5441, N5420, N1663);
xor XOR2 (N5442, N5439, N5367);
or OR3 (N5443, N5442, N3283, N6);
not NOT1 (N5444, N5422);
and AND2 (N5445, N5434, N5281);
or OR4 (N5446, N5441, N3117, N2845, N4180);
nand NAND3 (N5447, N5443, N3232, N4061);
buf BUF1 (N5448, N5445);
nor NOR3 (N5449, N5435, N663, N4623);
or OR4 (N5450, N5432, N2816, N3301, N16);
and AND4 (N5451, N5433, N3163, N5243, N2243);
not NOT1 (N5452, N5426);
or OR4 (N5453, N5440, N1564, N5397, N2150);
nor NOR3 (N5454, N5449, N1102, N1282);
and AND2 (N5455, N5447, N2522);
nand NAND3 (N5456, N5444, N1315, N1432);
nand NAND4 (N5457, N5454, N1429, N1507, N3495);
or OR2 (N5458, N5455, N3641);
buf BUF1 (N5459, N5458);
or OR2 (N5460, N5448, N929);
nand NAND4 (N5461, N5427, N203, N4848, N573);
nor NOR3 (N5462, N5452, N5142, N3398);
nand NAND3 (N5463, N5451, N5247, N1444);
buf BUF1 (N5464, N5453);
nand NAND3 (N5465, N5462, N3664, N3549);
nand NAND2 (N5466, N5461, N4029);
xor XOR2 (N5467, N5465, N1412);
and AND2 (N5468, N5467, N3029);
nor NOR3 (N5469, N5464, N655, N4400);
and AND2 (N5470, N5457, N1580);
not NOT1 (N5471, N5463);
nor NOR3 (N5472, N5456, N4188, N3931);
buf BUF1 (N5473, N5472);
xor XOR2 (N5474, N5469, N5461);
or OR4 (N5475, N5466, N4537, N5001, N4894);
and AND2 (N5476, N5460, N4788);
and AND3 (N5477, N5470, N4630, N2205);
xor XOR2 (N5478, N5468, N4005);
and AND2 (N5479, N5477, N3389);
and AND2 (N5480, N5450, N4431);
or OR4 (N5481, N5480, N2012, N5048, N1620);
buf BUF1 (N5482, N5476);
not NOT1 (N5483, N5446);
or OR2 (N5484, N5459, N4178);
buf BUF1 (N5485, N5484);
xor XOR2 (N5486, N5482, N765);
xor XOR2 (N5487, N5486, N2265);
xor XOR2 (N5488, N5481, N1979);
not NOT1 (N5489, N5479);
buf BUF1 (N5490, N5474);
xor XOR2 (N5491, N5490, N617);
or OR4 (N5492, N5473, N5426, N4706, N3918);
nand NAND2 (N5493, N5475, N648);
not NOT1 (N5494, N5492);
nand NAND3 (N5495, N5471, N1348, N3982);
buf BUF1 (N5496, N5489);
xor XOR2 (N5497, N5485, N655);
not NOT1 (N5498, N5495);
or OR3 (N5499, N5493, N685, N257);
and AND2 (N5500, N5487, N2173);
or OR2 (N5501, N5491, N4349);
not NOT1 (N5502, N5499);
not NOT1 (N5503, N5498);
and AND4 (N5504, N5497, N1940, N2864, N2676);
and AND3 (N5505, N5488, N956, N3987);
nor NOR2 (N5506, N5478, N4049);
nor NOR2 (N5507, N5502, N3061);
buf BUF1 (N5508, N5494);
xor XOR2 (N5509, N5483, N5070);
not NOT1 (N5510, N5509);
xor XOR2 (N5511, N5500, N2859);
buf BUF1 (N5512, N5501);
not NOT1 (N5513, N5511);
buf BUF1 (N5514, N5510);
not NOT1 (N5515, N5513);
nor NOR2 (N5516, N5515, N2077);
buf BUF1 (N5517, N5512);
buf BUF1 (N5518, N5508);
xor XOR2 (N5519, N5506, N3426);
not NOT1 (N5520, N5516);
nor NOR4 (N5521, N5514, N2531, N1889, N2846);
xor XOR2 (N5522, N5517, N2276);
xor XOR2 (N5523, N5505, N2230);
nand NAND2 (N5524, N5503, N1805);
buf BUF1 (N5525, N5496);
buf BUF1 (N5526, N5518);
not NOT1 (N5527, N5524);
and AND3 (N5528, N5520, N785, N4074);
not NOT1 (N5529, N5525);
nor NOR3 (N5530, N5523, N5494, N4273);
and AND2 (N5531, N5521, N3210);
nand NAND2 (N5532, N5527, N2275);
not NOT1 (N5533, N5504);
or OR2 (N5534, N5533, N4038);
nand NAND2 (N5535, N5534, N2783);
not NOT1 (N5536, N5526);
not NOT1 (N5537, N5530);
and AND2 (N5538, N5532, N1988);
nand NAND4 (N5539, N5522, N1595, N3672, N2386);
xor XOR2 (N5540, N5529, N2694);
not NOT1 (N5541, N5535);
or OR4 (N5542, N5528, N3767, N2570, N1242);
and AND4 (N5543, N5539, N4248, N767, N2382);
or OR4 (N5544, N5538, N1470, N1883, N2609);
nor NOR3 (N5545, N5540, N788, N1938);
xor XOR2 (N5546, N5543, N4216);
xor XOR2 (N5547, N5546, N667);
or OR4 (N5548, N5542, N1516, N1848, N4462);
and AND4 (N5549, N5519, N3159, N3130, N408);
nor NOR2 (N5550, N5541, N4148);
nor NOR2 (N5551, N5507, N4514);
nor NOR2 (N5552, N5551, N4562);
and AND2 (N5553, N5545, N4623);
nor NOR2 (N5554, N5550, N2511);
or OR3 (N5555, N5537, N5242, N5478);
or OR4 (N5556, N5547, N1075, N230, N3265);
nand NAND4 (N5557, N5552, N2190, N2525, N53);
not NOT1 (N5558, N5556);
nor NOR4 (N5559, N5558, N3950, N2894, N2937);
nand NAND4 (N5560, N5554, N3373, N5324, N1012);
xor XOR2 (N5561, N5555, N1698);
buf BUF1 (N5562, N5553);
or OR4 (N5563, N5557, N57, N2819, N5005);
not NOT1 (N5564, N5561);
nor NOR3 (N5565, N5548, N3187, N3839);
nor NOR2 (N5566, N5560, N2730);
nor NOR4 (N5567, N5564, N2165, N3494, N633);
or OR4 (N5568, N5544, N918, N4603, N527);
and AND4 (N5569, N5567, N2424, N329, N540);
not NOT1 (N5570, N5568);
xor XOR2 (N5571, N5569, N1610);
buf BUF1 (N5572, N5563);
xor XOR2 (N5573, N5531, N775);
not NOT1 (N5574, N5559);
xor XOR2 (N5575, N5571, N1835);
and AND3 (N5576, N5572, N2745, N5212);
or OR4 (N5577, N5575, N975, N3843, N3829);
or OR3 (N5578, N5570, N731, N2445);
nor NOR3 (N5579, N5562, N185, N1579);
and AND3 (N5580, N5576, N4184, N578);
buf BUF1 (N5581, N5577);
nor NOR2 (N5582, N5536, N5431);
nor NOR4 (N5583, N5578, N5553, N5057, N2631);
not NOT1 (N5584, N5549);
or OR4 (N5585, N5566, N3217, N1134, N2150);
nor NOR3 (N5586, N5584, N3957, N5522);
and AND2 (N5587, N5586, N4419);
or OR2 (N5588, N5565, N2275);
or OR3 (N5589, N5581, N839, N1471);
or OR2 (N5590, N5585, N1142);
buf BUF1 (N5591, N5587);
not NOT1 (N5592, N5589);
or OR2 (N5593, N5574, N2707);
and AND3 (N5594, N5573, N1130, N2311);
nor NOR2 (N5595, N5590, N2779);
nand NAND3 (N5596, N5593, N1673, N4198);
or OR3 (N5597, N5579, N4776, N2362);
buf BUF1 (N5598, N5595);
and AND2 (N5599, N5588, N384);
or OR2 (N5600, N5592, N4054);
not NOT1 (N5601, N5600);
xor XOR2 (N5602, N5583, N5482);
nor NOR2 (N5603, N5591, N2742);
nand NAND3 (N5604, N5601, N143, N1955);
or OR4 (N5605, N5599, N1033, N4466, N2776);
nor NOR4 (N5606, N5602, N3497, N1307, N2900);
buf BUF1 (N5607, N5603);
xor XOR2 (N5608, N5580, N295);
or OR4 (N5609, N5582, N5255, N1305, N3396);
xor XOR2 (N5610, N5596, N288);
buf BUF1 (N5611, N5608);
nand NAND2 (N5612, N5609, N4530);
or OR4 (N5613, N5610, N2040, N4208, N1361);
not NOT1 (N5614, N5607);
nor NOR4 (N5615, N5604, N5125, N2545, N3865);
and AND3 (N5616, N5612, N4351, N138);
nand NAND3 (N5617, N5616, N4105, N3114);
nor NOR2 (N5618, N5611, N4390);
and AND2 (N5619, N5594, N367);
not NOT1 (N5620, N5613);
nor NOR2 (N5621, N5605, N2304);
nand NAND2 (N5622, N5598, N2672);
buf BUF1 (N5623, N5614);
nand NAND3 (N5624, N5617, N4344, N1393);
not NOT1 (N5625, N5621);
or OR3 (N5626, N5623, N5462, N1664);
nor NOR3 (N5627, N5619, N1545, N3792);
xor XOR2 (N5628, N5625, N4161);
and AND4 (N5629, N5618, N13, N5327, N1362);
nor NOR2 (N5630, N5629, N2782);
not NOT1 (N5631, N5615);
xor XOR2 (N5632, N5626, N366);
nor NOR4 (N5633, N5631, N4140, N760, N20);
xor XOR2 (N5634, N5630, N1626);
nand NAND2 (N5635, N5624, N222);
or OR2 (N5636, N5606, N837);
and AND3 (N5637, N5620, N1848, N909);
or OR2 (N5638, N5635, N3036);
nand NAND2 (N5639, N5636, N1081);
buf BUF1 (N5640, N5632);
and AND2 (N5641, N5639, N3781);
and AND2 (N5642, N5634, N3792);
buf BUF1 (N5643, N5597);
buf BUF1 (N5644, N5637);
nor NOR2 (N5645, N5641, N4784);
not NOT1 (N5646, N5638);
and AND3 (N5647, N5627, N2104, N4331);
or OR3 (N5648, N5644, N842, N1218);
or OR2 (N5649, N5647, N2764);
and AND3 (N5650, N5645, N5438, N449);
not NOT1 (N5651, N5640);
xor XOR2 (N5652, N5646, N2501);
nand NAND3 (N5653, N5652, N5625, N4298);
buf BUF1 (N5654, N5648);
buf BUF1 (N5655, N5643);
or OR4 (N5656, N5633, N2104, N3694, N5156);
nand NAND4 (N5657, N5654, N2290, N4440, N4038);
or OR3 (N5658, N5656, N4136, N909);
nor NOR4 (N5659, N5657, N4747, N5506, N3513);
not NOT1 (N5660, N5651);
or OR4 (N5661, N5650, N985, N4136, N1383);
xor XOR2 (N5662, N5660, N463);
and AND4 (N5663, N5622, N86, N1903, N2957);
or OR2 (N5664, N5663, N1101);
not NOT1 (N5665, N5662);
nor NOR2 (N5666, N5628, N949);
or OR4 (N5667, N5666, N2874, N2664, N3226);
or OR3 (N5668, N5642, N438, N5434);
not NOT1 (N5669, N5665);
nor NOR2 (N5670, N5649, N311);
and AND2 (N5671, N5659, N4975);
xor XOR2 (N5672, N5670, N1469);
buf BUF1 (N5673, N5653);
buf BUF1 (N5674, N5655);
xor XOR2 (N5675, N5658, N1035);
and AND2 (N5676, N5673, N5010);
nand NAND3 (N5677, N5664, N4389, N5180);
and AND4 (N5678, N5668, N4262, N218, N4996);
or OR2 (N5679, N5676, N1575);
nor NOR4 (N5680, N5677, N1431, N2767, N3005);
nand NAND2 (N5681, N5678, N3495);
or OR3 (N5682, N5667, N2238, N876);
nor NOR3 (N5683, N5674, N4053, N4731);
nand NAND2 (N5684, N5672, N5128);
buf BUF1 (N5685, N5669);
or OR2 (N5686, N5681, N3955);
xor XOR2 (N5687, N5661, N2651);
nor NOR4 (N5688, N5682, N5167, N1660, N2292);
and AND2 (N5689, N5684, N19);
xor XOR2 (N5690, N5686, N2152);
not NOT1 (N5691, N5679);
not NOT1 (N5692, N5683);
not NOT1 (N5693, N5680);
nor NOR4 (N5694, N5690, N69, N170, N1918);
and AND2 (N5695, N5687, N323);
or OR4 (N5696, N5688, N4307, N906, N492);
nor NOR4 (N5697, N5696, N3454, N1668, N3375);
and AND3 (N5698, N5695, N2893, N4924);
or OR2 (N5699, N5671, N4084);
or OR2 (N5700, N5685, N165);
nor NOR4 (N5701, N5693, N1083, N5083, N2378);
and AND3 (N5702, N5700, N4189, N212);
buf BUF1 (N5703, N5691);
xor XOR2 (N5704, N5694, N2681);
nor NOR4 (N5705, N5689, N2734, N5429, N3160);
not NOT1 (N5706, N5675);
buf BUF1 (N5707, N5706);
nor NOR2 (N5708, N5697, N5469);
not NOT1 (N5709, N5707);
nand NAND2 (N5710, N5705, N5632);
or OR2 (N5711, N5701, N4955);
or OR3 (N5712, N5698, N5638, N3091);
and AND3 (N5713, N5710, N4236, N536);
or OR2 (N5714, N5692, N1239);
buf BUF1 (N5715, N5708);
buf BUF1 (N5716, N5704);
and AND2 (N5717, N5715, N1517);
not NOT1 (N5718, N5703);
nor NOR2 (N5719, N5717, N3170);
buf BUF1 (N5720, N5719);
nand NAND2 (N5721, N5712, N4713);
nor NOR2 (N5722, N5702, N244);
nor NOR2 (N5723, N5722, N1740);
not NOT1 (N5724, N5711);
or OR4 (N5725, N5718, N3054, N4314, N5318);
xor XOR2 (N5726, N5723, N4102);
nor NOR3 (N5727, N5716, N2419, N1788);
not NOT1 (N5728, N5720);
nor NOR2 (N5729, N5699, N4820);
xor XOR2 (N5730, N5709, N3188);
not NOT1 (N5731, N5727);
xor XOR2 (N5732, N5726, N173);
not NOT1 (N5733, N5729);
or OR2 (N5734, N5732, N3963);
nor NOR3 (N5735, N5733, N1130, N5586);
xor XOR2 (N5736, N5724, N5482);
xor XOR2 (N5737, N5731, N3434);
not NOT1 (N5738, N5737);
and AND2 (N5739, N5735, N5647);
not NOT1 (N5740, N5730);
not NOT1 (N5741, N5728);
nor NOR3 (N5742, N5738, N1366, N732);
nand NAND2 (N5743, N5739, N2545);
not NOT1 (N5744, N5736);
or OR4 (N5745, N5741, N1032, N109, N4096);
nor NOR3 (N5746, N5714, N2429, N4312);
not NOT1 (N5747, N5734);
nand NAND4 (N5748, N5743, N185, N3474, N4290);
not NOT1 (N5749, N5721);
nor NOR3 (N5750, N5713, N2276, N931);
not NOT1 (N5751, N5748);
buf BUF1 (N5752, N5745);
nand NAND4 (N5753, N5746, N4705, N3532, N1982);
buf BUF1 (N5754, N5753);
nand NAND3 (N5755, N5749, N1131, N4553);
xor XOR2 (N5756, N5740, N3544);
or OR2 (N5757, N5751, N4843);
buf BUF1 (N5758, N5744);
xor XOR2 (N5759, N5747, N1038);
nor NOR2 (N5760, N5750, N343);
not NOT1 (N5761, N5760);
buf BUF1 (N5762, N5756);
or OR4 (N5763, N5761, N5333, N2620, N3619);
buf BUF1 (N5764, N5752);
or OR2 (N5765, N5725, N4735);
not NOT1 (N5766, N5755);
nand NAND3 (N5767, N5754, N4033, N1847);
not NOT1 (N5768, N5763);
and AND2 (N5769, N5768, N5315);
or OR4 (N5770, N5769, N5143, N3400, N5451);
nand NAND4 (N5771, N5766, N5018, N2432, N2110);
nand NAND3 (N5772, N5764, N5757, N3878);
buf BUF1 (N5773, N1476);
not NOT1 (N5774, N5773);
nand NAND4 (N5775, N5765, N980, N4175, N1345);
or OR4 (N5776, N5775, N1895, N3987, N1081);
buf BUF1 (N5777, N5767);
xor XOR2 (N5778, N5771, N4283);
or OR2 (N5779, N5776, N1032);
not NOT1 (N5780, N5762);
or OR4 (N5781, N5774, N4218, N1860, N2053);
nor NOR2 (N5782, N5781, N5281);
buf BUF1 (N5783, N5759);
not NOT1 (N5784, N5782);
and AND2 (N5785, N5758, N382);
not NOT1 (N5786, N5784);
nand NAND4 (N5787, N5772, N4431, N1514, N1382);
xor XOR2 (N5788, N5777, N3560);
xor XOR2 (N5789, N5787, N3810);
nand NAND3 (N5790, N5783, N3297, N2507);
not NOT1 (N5791, N5779);
not NOT1 (N5792, N5785);
buf BUF1 (N5793, N5786);
nand NAND4 (N5794, N5780, N170, N2624, N5631);
and AND4 (N5795, N5791, N2467, N3180, N2608);
nor NOR3 (N5796, N5790, N5012, N1645);
xor XOR2 (N5797, N5789, N2615);
buf BUF1 (N5798, N5770);
nand NAND3 (N5799, N5778, N4012, N1322);
and AND4 (N5800, N5788, N3899, N4194, N4246);
xor XOR2 (N5801, N5742, N4764);
or OR2 (N5802, N5792, N1207);
nor NOR3 (N5803, N5798, N3315, N5457);
or OR2 (N5804, N5801, N172);
not NOT1 (N5805, N5796);
nor NOR4 (N5806, N5805, N5421, N5653, N4045);
xor XOR2 (N5807, N5793, N5113);
nand NAND3 (N5808, N5800, N2948, N697);
nand NAND4 (N5809, N5795, N616, N3772, N3825);
xor XOR2 (N5810, N5802, N719);
nand NAND3 (N5811, N5807, N720, N444);
nor NOR4 (N5812, N5803, N4582, N1198, N4354);
nand NAND3 (N5813, N5794, N4494, N477);
buf BUF1 (N5814, N5799);
nand NAND3 (N5815, N5811, N936, N4769);
xor XOR2 (N5816, N5814, N1416);
or OR2 (N5817, N5813, N3681);
or OR3 (N5818, N5815, N3446, N2179);
buf BUF1 (N5819, N5818);
or OR4 (N5820, N5817, N980, N5445, N1093);
xor XOR2 (N5821, N5810, N3622);
or OR2 (N5822, N5797, N3500);
nor NOR4 (N5823, N5822, N957, N3160, N3587);
not NOT1 (N5824, N5821);
nand NAND2 (N5825, N5809, N4944);
nor NOR4 (N5826, N5824, N4518, N4604, N4386);
nand NAND3 (N5827, N5808, N4051, N186);
or OR4 (N5828, N5820, N5474, N5550, N845);
xor XOR2 (N5829, N5806, N2402);
buf BUF1 (N5830, N5804);
xor XOR2 (N5831, N5823, N169);
nor NOR4 (N5832, N5826, N309, N3534, N3807);
buf BUF1 (N5833, N5829);
not NOT1 (N5834, N5830);
nand NAND2 (N5835, N5831, N5267);
or OR4 (N5836, N5834, N1167, N491, N3002);
not NOT1 (N5837, N5828);
or OR4 (N5838, N5832, N1267, N5351, N1093);
nor NOR2 (N5839, N5833, N3321);
not NOT1 (N5840, N5819);
or OR2 (N5841, N5840, N3431);
and AND3 (N5842, N5835, N1406, N3997);
nand NAND2 (N5843, N5842, N1277);
nor NOR3 (N5844, N5839, N3276, N1602);
buf BUF1 (N5845, N5812);
not NOT1 (N5846, N5827);
and AND2 (N5847, N5844, N63);
xor XOR2 (N5848, N5841, N1461);
nand NAND2 (N5849, N5836, N3170);
and AND4 (N5850, N5825, N4203, N3395, N3285);
and AND3 (N5851, N5846, N5440, N5487);
nand NAND3 (N5852, N5849, N4399, N5030);
nor NOR2 (N5853, N5850, N1290);
xor XOR2 (N5854, N5848, N1123);
xor XOR2 (N5855, N5847, N1585);
nand NAND4 (N5856, N5845, N4891, N579, N4555);
not NOT1 (N5857, N5854);
xor XOR2 (N5858, N5837, N2834);
nor NOR4 (N5859, N5852, N825, N1924, N2121);
or OR2 (N5860, N5851, N3604);
nor NOR3 (N5861, N5855, N4560, N5719);
and AND3 (N5862, N5838, N829, N4492);
not NOT1 (N5863, N5853);
nor NOR2 (N5864, N5861, N483);
nand NAND2 (N5865, N5858, N2178);
buf BUF1 (N5866, N5865);
or OR3 (N5867, N5856, N71, N3026);
nand NAND4 (N5868, N5863, N3968, N152, N5859);
not NOT1 (N5869, N602);
not NOT1 (N5870, N5843);
or OR3 (N5871, N5870, N2955, N5349);
and AND3 (N5872, N5862, N2876, N5325);
nand NAND3 (N5873, N5867, N5004, N1731);
and AND4 (N5874, N5816, N1833, N3647, N2566);
xor XOR2 (N5875, N5860, N4099);
buf BUF1 (N5876, N5874);
not NOT1 (N5877, N5871);
and AND4 (N5878, N5876, N2294, N767, N2282);
or OR3 (N5879, N5868, N2756, N918);
and AND3 (N5880, N5857, N3977, N3987);
nor NOR4 (N5881, N5879, N1684, N3492, N2045);
xor XOR2 (N5882, N5880, N2927);
and AND4 (N5883, N5872, N2522, N5217, N2577);
buf BUF1 (N5884, N5864);
buf BUF1 (N5885, N5884);
buf BUF1 (N5886, N5883);
nand NAND2 (N5887, N5873, N4223);
xor XOR2 (N5888, N5885, N5531);
nor NOR2 (N5889, N5887, N1520);
not NOT1 (N5890, N5866);
or OR2 (N5891, N5882, N3908);
and AND2 (N5892, N5891, N3279);
or OR3 (N5893, N5877, N468, N2763);
not NOT1 (N5894, N5892);
or OR2 (N5895, N5886, N5723);
nand NAND3 (N5896, N5889, N812, N1881);
xor XOR2 (N5897, N5893, N3788);
nor NOR4 (N5898, N5895, N1159, N3918, N4754);
not NOT1 (N5899, N5881);
or OR3 (N5900, N5888, N1406, N1761);
nand NAND4 (N5901, N5896, N4480, N960, N4261);
buf BUF1 (N5902, N5878);
nor NOR4 (N5903, N5869, N2724, N2748, N191);
not NOT1 (N5904, N5900);
or OR3 (N5905, N5903, N234, N3210);
not NOT1 (N5906, N5890);
or OR3 (N5907, N5901, N481, N3418);
not NOT1 (N5908, N5906);
or OR2 (N5909, N5897, N1586);
xor XOR2 (N5910, N5894, N4573);
nor NOR2 (N5911, N5909, N414);
and AND4 (N5912, N5905, N2570, N3847, N4944);
nor NOR4 (N5913, N5907, N2656, N3179, N5895);
not NOT1 (N5914, N5899);
and AND4 (N5915, N5912, N4249, N2531, N1811);
xor XOR2 (N5916, N5875, N2326);
nand NAND2 (N5917, N5916, N5227);
nor NOR2 (N5918, N5908, N4772);
and AND4 (N5919, N5918, N5909, N3936, N2039);
not NOT1 (N5920, N5917);
buf BUF1 (N5921, N5920);
or OR3 (N5922, N5913, N3120, N5146);
nor NOR4 (N5923, N5910, N561, N5209, N4078);
or OR4 (N5924, N5904, N2524, N3074, N167);
nand NAND2 (N5925, N5921, N3429);
nand NAND4 (N5926, N5923, N854, N2951, N1842);
xor XOR2 (N5927, N5902, N4060);
and AND4 (N5928, N5922, N1095, N321, N2618);
buf BUF1 (N5929, N5915);
or OR3 (N5930, N5926, N4125, N1997);
xor XOR2 (N5931, N5925, N3509);
nand NAND2 (N5932, N5919, N2149);
and AND2 (N5933, N5930, N544);
nor NOR2 (N5934, N5911, N2657);
or OR4 (N5935, N5898, N4869, N1, N3405);
or OR3 (N5936, N5929, N1410, N3845);
xor XOR2 (N5937, N5936, N2971);
and AND3 (N5938, N5927, N970, N5689);
not NOT1 (N5939, N5932);
not NOT1 (N5940, N5931);
xor XOR2 (N5941, N5924, N1419);
buf BUF1 (N5942, N5914);
and AND2 (N5943, N5940, N4497);
or OR4 (N5944, N5933, N4654, N266, N1538);
or OR4 (N5945, N5942, N5605, N1103, N952);
xor XOR2 (N5946, N5945, N4328);
nand NAND3 (N5947, N5935, N1738, N663);
and AND3 (N5948, N5941, N1916, N1005);
and AND3 (N5949, N5943, N2900, N3682);
xor XOR2 (N5950, N5934, N454);
not NOT1 (N5951, N5944);
buf BUF1 (N5952, N5949);
or OR4 (N5953, N5928, N929, N3368, N4805);
nor NOR2 (N5954, N5950, N2276);
xor XOR2 (N5955, N5938, N2180);
buf BUF1 (N5956, N5947);
xor XOR2 (N5957, N5952, N5568);
and AND4 (N5958, N5955, N4441, N2690, N5950);
not NOT1 (N5959, N5948);
nor NOR2 (N5960, N5951, N1523);
or OR2 (N5961, N5958, N4255);
xor XOR2 (N5962, N5961, N4815);
xor XOR2 (N5963, N5960, N5053);
nor NOR4 (N5964, N5953, N5652, N1996, N1170);
buf BUF1 (N5965, N5939);
or OR2 (N5966, N5937, N3631);
or OR2 (N5967, N5959, N2476);
and AND2 (N5968, N5967, N2524);
and AND4 (N5969, N5946, N1523, N2458, N2372);
buf BUF1 (N5970, N5966);
nand NAND2 (N5971, N5968, N4956);
nor NOR2 (N5972, N5971, N206);
xor XOR2 (N5973, N5970, N856);
or OR2 (N5974, N5965, N333);
nor NOR3 (N5975, N5974, N2148, N1679);
buf BUF1 (N5976, N5969);
or OR3 (N5977, N5954, N1275, N5585);
not NOT1 (N5978, N5973);
nand NAND4 (N5979, N5957, N1641, N4188, N4235);
nand NAND2 (N5980, N5977, N2764);
not NOT1 (N5981, N5976);
and AND4 (N5982, N5981, N4142, N1524, N3990);
not NOT1 (N5983, N5963);
nor NOR3 (N5984, N5978, N4124, N5136);
or OR4 (N5985, N5980, N535, N5013, N21);
and AND4 (N5986, N5984, N3378, N3800, N1348);
not NOT1 (N5987, N5962);
or OR2 (N5988, N5986, N3370);
nor NOR4 (N5989, N5956, N3793, N467, N2450);
not NOT1 (N5990, N5985);
nor NOR3 (N5991, N5975, N5293, N2581);
and AND2 (N5992, N5990, N1033);
buf BUF1 (N5993, N5972);
and AND3 (N5994, N5993, N4269, N746);
and AND3 (N5995, N5979, N4451, N3022);
buf BUF1 (N5996, N5983);
xor XOR2 (N5997, N5964, N3681);
nor NOR2 (N5998, N5994, N2199);
xor XOR2 (N5999, N5987, N5296);
xor XOR2 (N6000, N5982, N4638);
and AND3 (N6001, N5996, N1974, N1123);
nand NAND2 (N6002, N5995, N2045);
or OR3 (N6003, N5999, N1702, N5992);
and AND4 (N6004, N4643, N2454, N3228, N5514);
not NOT1 (N6005, N5989);
or OR4 (N6006, N5991, N1891, N4425, N2257);
or OR3 (N6007, N5997, N4568, N4782);
not NOT1 (N6008, N5998);
nand NAND3 (N6009, N6002, N3128, N5488);
or OR3 (N6010, N6005, N270, N4348);
or OR4 (N6011, N6009, N4068, N3147, N4277);
and AND4 (N6012, N5988, N5686, N3940, N5436);
buf BUF1 (N6013, N6001);
not NOT1 (N6014, N6010);
nand NAND3 (N6015, N6012, N1163, N2197);
buf BUF1 (N6016, N6003);
nand NAND2 (N6017, N6007, N3067);
nor NOR3 (N6018, N6006, N3188, N2291);
and AND2 (N6019, N6014, N3250);
not NOT1 (N6020, N6013);
not NOT1 (N6021, N6020);
nor NOR2 (N6022, N6017, N5713);
or OR4 (N6023, N6021, N321, N3746, N5222);
or OR2 (N6024, N6018, N2449);
xor XOR2 (N6025, N6016, N3387);
nand NAND4 (N6026, N6022, N5992, N5329, N5932);
nor NOR2 (N6027, N6008, N657);
xor XOR2 (N6028, N6026, N722);
buf BUF1 (N6029, N6011);
nand NAND4 (N6030, N6028, N4982, N4327, N5983);
xor XOR2 (N6031, N6024, N4967);
and AND4 (N6032, N6029, N1656, N5170, N5867);
and AND2 (N6033, N6031, N1003);
buf BUF1 (N6034, N6015);
or OR4 (N6035, N6032, N604, N3672, N5863);
xor XOR2 (N6036, N6023, N2744);
or OR2 (N6037, N6034, N803);
not NOT1 (N6038, N6000);
or OR3 (N6039, N6030, N5515, N2469);
and AND2 (N6040, N6019, N4135);
xor XOR2 (N6041, N6004, N4982);
or OR3 (N6042, N6040, N5095, N1830);
not NOT1 (N6043, N6035);
and AND3 (N6044, N6043, N325, N415);
xor XOR2 (N6045, N6033, N2934);
nand NAND4 (N6046, N6039, N4081, N5760, N1568);
and AND3 (N6047, N6041, N484, N3644);
buf BUF1 (N6048, N6025);
or OR4 (N6049, N6047, N4252, N4129, N2691);
and AND4 (N6050, N6046, N5989, N2914, N1868);
nand NAND3 (N6051, N6038, N2579, N2001);
nand NAND4 (N6052, N6051, N4315, N3554, N1916);
nor NOR4 (N6053, N6027, N2605, N4604, N427);
or OR3 (N6054, N6042, N2627, N4542);
not NOT1 (N6055, N6037);
and AND4 (N6056, N6044, N4099, N2007, N5601);
buf BUF1 (N6057, N6048);
buf BUF1 (N6058, N6054);
buf BUF1 (N6059, N6055);
or OR2 (N6060, N6036, N2783);
nor NOR3 (N6061, N6050, N1791, N3188);
xor XOR2 (N6062, N6059, N2851);
and AND2 (N6063, N6045, N1233);
or OR2 (N6064, N6060, N1135);
buf BUF1 (N6065, N6063);
or OR4 (N6066, N6049, N4280, N4605, N4176);
or OR2 (N6067, N6056, N52);
not NOT1 (N6068, N6066);
or OR2 (N6069, N6061, N734);
or OR2 (N6070, N6067, N3091);
nand NAND2 (N6071, N6069, N1865);
nand NAND4 (N6072, N6057, N4221, N5667, N2397);
nor NOR4 (N6073, N6053, N4693, N4690, N2118);
nand NAND4 (N6074, N6052, N3347, N220, N1577);
not NOT1 (N6075, N6068);
xor XOR2 (N6076, N6074, N5458);
or OR4 (N6077, N6058, N726, N3593, N720);
buf BUF1 (N6078, N6064);
buf BUF1 (N6079, N6077);
not NOT1 (N6080, N6076);
buf BUF1 (N6081, N6070);
not NOT1 (N6082, N6075);
not NOT1 (N6083, N6081);
and AND3 (N6084, N6073, N2756, N5394);
and AND3 (N6085, N6084, N5354, N2044);
and AND2 (N6086, N6082, N2572);
not NOT1 (N6087, N6071);
not NOT1 (N6088, N6079);
not NOT1 (N6089, N6078);
nand NAND4 (N6090, N6087, N5257, N632, N696);
nor NOR4 (N6091, N6088, N2837, N3525, N4603);
buf BUF1 (N6092, N6083);
buf BUF1 (N6093, N6086);
and AND3 (N6094, N6089, N2223, N4395);
or OR4 (N6095, N6072, N5736, N183, N5166);
nand NAND4 (N6096, N6080, N4116, N1888, N3844);
buf BUF1 (N6097, N6095);
buf BUF1 (N6098, N6091);
xor XOR2 (N6099, N6096, N5538);
buf BUF1 (N6100, N6097);
buf BUF1 (N6101, N6098);
nand NAND4 (N6102, N6093, N2384, N4480, N5029);
nand NAND2 (N6103, N6092, N580);
xor XOR2 (N6104, N6062, N5953);
and AND4 (N6105, N6090, N4624, N3458, N2120);
or OR4 (N6106, N6101, N4741, N2410, N2599);
xor XOR2 (N6107, N6104, N5930);
and AND3 (N6108, N6100, N521, N2575);
and AND4 (N6109, N6065, N1570, N2266, N2708);
not NOT1 (N6110, N6099);
nand NAND3 (N6111, N6085, N1467, N3439);
and AND2 (N6112, N6110, N2496);
not NOT1 (N6113, N6108);
nor NOR2 (N6114, N6102, N3508);
buf BUF1 (N6115, N6114);
nor NOR2 (N6116, N6115, N5064);
or OR3 (N6117, N6112, N92, N1834);
not NOT1 (N6118, N6107);
xor XOR2 (N6119, N6106, N5600);
buf BUF1 (N6120, N6109);
xor XOR2 (N6121, N6118, N3578);
nor NOR4 (N6122, N6105, N4026, N2442, N5254);
nand NAND4 (N6123, N6122, N2968, N4586, N4766);
xor XOR2 (N6124, N6121, N865);
nand NAND4 (N6125, N6103, N3919, N954, N2376);
nor NOR4 (N6126, N6119, N3348, N1802, N6092);
nand NAND2 (N6127, N6124, N3777);
not NOT1 (N6128, N6117);
buf BUF1 (N6129, N6127);
or OR4 (N6130, N6123, N4746, N536, N3184);
buf BUF1 (N6131, N6111);
and AND3 (N6132, N6130, N1012, N1673);
nand NAND4 (N6133, N6128, N4067, N142, N3544);
nor NOR3 (N6134, N6131, N3383, N1542);
nor NOR2 (N6135, N6094, N1145);
or OR4 (N6136, N6135, N3281, N4659, N2895);
not NOT1 (N6137, N6129);
xor XOR2 (N6138, N6116, N2620);
xor XOR2 (N6139, N6113, N5261);
xor XOR2 (N6140, N6137, N2651);
or OR3 (N6141, N6136, N23, N635);
xor XOR2 (N6142, N6138, N4525);
xor XOR2 (N6143, N6141, N433);
nor NOR4 (N6144, N6142, N1635, N4448, N5246);
xor XOR2 (N6145, N6132, N1957);
nand NAND2 (N6146, N6126, N1052);
xor XOR2 (N6147, N6143, N5139);
or OR2 (N6148, N6125, N1725);
buf BUF1 (N6149, N6145);
nor NOR4 (N6150, N6133, N4210, N5387, N1486);
or OR3 (N6151, N6149, N5738, N1909);
xor XOR2 (N6152, N6146, N1142);
xor XOR2 (N6153, N6151, N4701);
buf BUF1 (N6154, N6148);
nand NAND3 (N6155, N6150, N548, N5005);
and AND2 (N6156, N6155, N3761);
or OR4 (N6157, N6144, N3252, N4963, N4335);
buf BUF1 (N6158, N6156);
xor XOR2 (N6159, N6120, N3182);
or OR3 (N6160, N6140, N4280, N5450);
and AND4 (N6161, N6158, N2429, N2206, N2693);
and AND2 (N6162, N6147, N4956);
or OR3 (N6163, N6159, N2716, N234);
and AND3 (N6164, N6153, N110, N5936);
nand NAND4 (N6165, N6162, N4444, N5739, N442);
nor NOR2 (N6166, N6161, N2709);
nand NAND4 (N6167, N6165, N639, N1786, N5232);
or OR3 (N6168, N6166, N4106, N4055);
xor XOR2 (N6169, N6152, N3222);
nand NAND2 (N6170, N6168, N4222);
buf BUF1 (N6171, N6164);
not NOT1 (N6172, N6163);
not NOT1 (N6173, N6171);
buf BUF1 (N6174, N6167);
not NOT1 (N6175, N6169);
buf BUF1 (N6176, N6175);
not NOT1 (N6177, N6170);
nand NAND4 (N6178, N6139, N639, N1575, N1508);
nand NAND3 (N6179, N6176, N4029, N2008);
not NOT1 (N6180, N6179);
xor XOR2 (N6181, N6172, N1180);
nand NAND3 (N6182, N6134, N1251, N4888);
buf BUF1 (N6183, N6182);
not NOT1 (N6184, N6178);
or OR2 (N6185, N6157, N3181);
nand NAND4 (N6186, N6177, N5748, N4935, N788);
nand NAND2 (N6187, N6186, N2882);
buf BUF1 (N6188, N6187);
nor NOR2 (N6189, N6174, N3196);
buf BUF1 (N6190, N6185);
or OR2 (N6191, N6184, N540);
xor XOR2 (N6192, N6181, N3534);
nor NOR3 (N6193, N6183, N4797, N2633);
buf BUF1 (N6194, N6191);
nor NOR3 (N6195, N6154, N4871, N1955);
nand NAND3 (N6196, N6194, N5899, N3195);
or OR2 (N6197, N6193, N780);
nand NAND4 (N6198, N6160, N1674, N1901, N2548);
buf BUF1 (N6199, N6173);
xor XOR2 (N6200, N6196, N2527);
nor NOR4 (N6201, N6199, N569, N2926, N3236);
not NOT1 (N6202, N6197);
nor NOR2 (N6203, N6192, N4847);
or OR3 (N6204, N6201, N3018, N3136);
buf BUF1 (N6205, N6190);
or OR4 (N6206, N6198, N5685, N947, N1714);
and AND4 (N6207, N6205, N4137, N4649, N1195);
buf BUF1 (N6208, N6195);
and AND4 (N6209, N6188, N3378, N813, N3507);
not NOT1 (N6210, N6200);
or OR4 (N6211, N6189, N4794, N234, N5726);
nor NOR4 (N6212, N6204, N4829, N1054, N6048);
not NOT1 (N6213, N6207);
buf BUF1 (N6214, N6180);
and AND2 (N6215, N6203, N6130);
or OR4 (N6216, N6211, N1857, N2195, N4176);
xor XOR2 (N6217, N6209, N3462);
or OR2 (N6218, N6202, N3385);
xor XOR2 (N6219, N6215, N1602);
buf BUF1 (N6220, N6219);
not NOT1 (N6221, N6217);
not NOT1 (N6222, N6206);
nor NOR3 (N6223, N6210, N5654, N1271);
nand NAND2 (N6224, N6216, N93);
nor NOR3 (N6225, N6220, N4710, N6016);
buf BUF1 (N6226, N6222);
not NOT1 (N6227, N6224);
or OR4 (N6228, N6213, N4075, N1242, N724);
and AND3 (N6229, N6218, N3001, N4113);
and AND2 (N6230, N6208, N2025);
nor NOR4 (N6231, N6230, N270, N4720, N811);
nor NOR3 (N6232, N6214, N1266, N148);
nor NOR4 (N6233, N6226, N5827, N3613, N5251);
nand NAND2 (N6234, N6223, N718);
nand NAND3 (N6235, N6233, N4306, N3207);
or OR4 (N6236, N6225, N1138, N1221, N2263);
or OR2 (N6237, N6212, N1556);
not NOT1 (N6238, N6235);
nand NAND3 (N6239, N6231, N4501, N3343);
or OR3 (N6240, N6239, N4086, N4416);
nor NOR2 (N6241, N6221, N3975);
and AND3 (N6242, N6234, N1321, N989);
xor XOR2 (N6243, N6238, N1544);
not NOT1 (N6244, N6236);
not NOT1 (N6245, N6241);
buf BUF1 (N6246, N6232);
not NOT1 (N6247, N6227);
and AND2 (N6248, N6243, N2478);
nand NAND2 (N6249, N6229, N716);
buf BUF1 (N6250, N6244);
nor NOR2 (N6251, N6248, N5745);
xor XOR2 (N6252, N6245, N1552);
and AND2 (N6253, N6247, N4205);
or OR4 (N6254, N6253, N4476, N2859, N3238);
not NOT1 (N6255, N6249);
buf BUF1 (N6256, N6228);
or OR4 (N6257, N6237, N1304, N534, N4315);
and AND3 (N6258, N6240, N2602, N5658);
xor XOR2 (N6259, N6251, N1898);
buf BUF1 (N6260, N6242);
xor XOR2 (N6261, N6255, N5905);
xor XOR2 (N6262, N6250, N3286);
or OR4 (N6263, N6256, N5971, N5316, N4091);
xor XOR2 (N6264, N6260, N4939);
or OR2 (N6265, N6257, N3818);
or OR3 (N6266, N6263, N917, N2530);
or OR2 (N6267, N6252, N882);
and AND2 (N6268, N6254, N5069);
xor XOR2 (N6269, N6258, N3646);
xor XOR2 (N6270, N6266, N647);
xor XOR2 (N6271, N6269, N6239);
and AND4 (N6272, N6271, N962, N3550, N1964);
and AND4 (N6273, N6259, N1404, N3163, N5680);
nand NAND4 (N6274, N6261, N5795, N3362, N2777);
or OR2 (N6275, N6264, N839);
buf BUF1 (N6276, N6268);
buf BUF1 (N6277, N6265);
buf BUF1 (N6278, N6272);
xor XOR2 (N6279, N6273, N4249);
xor XOR2 (N6280, N6270, N507);
buf BUF1 (N6281, N6267);
buf BUF1 (N6282, N6280);
nand NAND2 (N6283, N6246, N160);
xor XOR2 (N6284, N6275, N2086);
or OR3 (N6285, N6282, N1525, N3504);
nor NOR4 (N6286, N6262, N1369, N6047, N17);
not NOT1 (N6287, N6274);
nand NAND4 (N6288, N6286, N295, N2629, N4812);
xor XOR2 (N6289, N6278, N4987);
and AND2 (N6290, N6288, N1596);
not NOT1 (N6291, N6290);
or OR2 (N6292, N6284, N648);
or OR3 (N6293, N6285, N4502, N2093);
nand NAND4 (N6294, N6292, N5913, N5021, N451);
and AND3 (N6295, N6281, N6093, N770);
buf BUF1 (N6296, N6293);
xor XOR2 (N6297, N6283, N2338);
buf BUF1 (N6298, N6297);
nand NAND3 (N6299, N6277, N1496, N4149);
buf BUF1 (N6300, N6279);
not NOT1 (N6301, N6300);
or OR2 (N6302, N6276, N4649);
nand NAND2 (N6303, N6287, N2736);
and AND4 (N6304, N6298, N3550, N1787, N768);
and AND3 (N6305, N6291, N6291, N885);
nor NOR4 (N6306, N6296, N4705, N5079, N6253);
nand NAND4 (N6307, N6303, N2178, N4750, N5522);
nor NOR3 (N6308, N6305, N1700, N4849);
nor NOR3 (N6309, N6295, N60, N137);
nand NAND2 (N6310, N6308, N5512);
not NOT1 (N6311, N6304);
buf BUF1 (N6312, N6310);
nor NOR3 (N6313, N6289, N2319, N2050);
xor XOR2 (N6314, N6306, N3332);
and AND3 (N6315, N6294, N708, N2178);
nand NAND3 (N6316, N6299, N4426, N4420);
nor NOR3 (N6317, N6316, N829, N3197);
buf BUF1 (N6318, N6311);
and AND2 (N6319, N6313, N5593);
not NOT1 (N6320, N6301);
and AND4 (N6321, N6317, N6034, N1403, N2250);
not NOT1 (N6322, N6302);
not NOT1 (N6323, N6322);
or OR3 (N6324, N6312, N5630, N4993);
buf BUF1 (N6325, N6318);
or OR4 (N6326, N6324, N3540, N2109, N6289);
and AND2 (N6327, N6325, N633);
xor XOR2 (N6328, N6309, N1213);
buf BUF1 (N6329, N6320);
not NOT1 (N6330, N6314);
not NOT1 (N6331, N6321);
nand NAND3 (N6332, N6329, N134, N3090);
not NOT1 (N6333, N6326);
xor XOR2 (N6334, N6315, N788);
or OR2 (N6335, N6319, N3346);
nand NAND4 (N6336, N6334, N3952, N535, N2993);
and AND3 (N6337, N6332, N2579, N4827);
xor XOR2 (N6338, N6323, N5969);
nor NOR2 (N6339, N6328, N5533);
xor XOR2 (N6340, N6307, N820);
nand NAND2 (N6341, N6333, N3728);
or OR3 (N6342, N6336, N2988, N608);
and AND4 (N6343, N6337, N4495, N1020, N5475);
xor XOR2 (N6344, N6335, N5437);
or OR3 (N6345, N6343, N5586, N925);
xor XOR2 (N6346, N6331, N1402);
buf BUF1 (N6347, N6339);
xor XOR2 (N6348, N6340, N6333);
and AND4 (N6349, N6330, N1153, N2832, N4535);
nand NAND4 (N6350, N6342, N1742, N3659, N2317);
and AND2 (N6351, N6349, N5143);
nor NOR3 (N6352, N6341, N4288, N1328);
not NOT1 (N6353, N6344);
xor XOR2 (N6354, N6345, N2960);
and AND4 (N6355, N6327, N3949, N6235, N2521);
nand NAND4 (N6356, N6352, N2640, N3451, N4602);
and AND3 (N6357, N6353, N2699, N446);
buf BUF1 (N6358, N6354);
nand NAND3 (N6359, N6358, N4308, N5017);
xor XOR2 (N6360, N6355, N5712);
not NOT1 (N6361, N6348);
xor XOR2 (N6362, N6356, N3150);
and AND4 (N6363, N6351, N3877, N4872, N569);
nand NAND2 (N6364, N6338, N1733);
xor XOR2 (N6365, N6346, N1649);
or OR2 (N6366, N6363, N2623);
buf BUF1 (N6367, N6359);
and AND4 (N6368, N6357, N2222, N1722, N2779);
and AND3 (N6369, N6360, N1497, N2277);
not NOT1 (N6370, N6368);
nor NOR4 (N6371, N6350, N4121, N2724, N3754);
not NOT1 (N6372, N6347);
nor NOR3 (N6373, N6366, N3580, N3461);
nand NAND4 (N6374, N6367, N1075, N1443, N1635);
xor XOR2 (N6375, N6370, N1010);
nor NOR4 (N6376, N6361, N4894, N5879, N4226);
nand NAND3 (N6377, N6369, N1861, N5046);
xor XOR2 (N6378, N6377, N4515);
xor XOR2 (N6379, N6373, N3011);
and AND2 (N6380, N6362, N3993);
buf BUF1 (N6381, N6378);
or OR3 (N6382, N6379, N2698, N1417);
nor NOR3 (N6383, N6380, N6380, N6350);
or OR4 (N6384, N6371, N4441, N5866, N4942);
nand NAND2 (N6385, N6364, N5833);
nand NAND4 (N6386, N6385, N736, N194, N3105);
and AND3 (N6387, N6365, N1010, N3330);
xor XOR2 (N6388, N6386, N2415);
nand NAND4 (N6389, N6382, N118, N2188, N4);
xor XOR2 (N6390, N6389, N359);
or OR3 (N6391, N6387, N2039, N2856);
buf BUF1 (N6392, N6374);
not NOT1 (N6393, N6388);
buf BUF1 (N6394, N6376);
buf BUF1 (N6395, N6375);
not NOT1 (N6396, N6381);
not NOT1 (N6397, N6393);
not NOT1 (N6398, N6390);
nor NOR2 (N6399, N6395, N3485);
and AND2 (N6400, N6399, N2914);
xor XOR2 (N6401, N6398, N5043);
nor NOR4 (N6402, N6400, N2559, N2118, N3283);
nor NOR4 (N6403, N6391, N3243, N3486, N3913);
or OR4 (N6404, N6394, N632, N989, N1066);
nor NOR3 (N6405, N6396, N3739, N1808);
or OR3 (N6406, N6384, N3203, N1262);
not NOT1 (N6407, N6397);
not NOT1 (N6408, N6401);
or OR4 (N6409, N6408, N5459, N2881, N5671);
not NOT1 (N6410, N6383);
or OR2 (N6411, N6404, N2251);
not NOT1 (N6412, N6410);
or OR4 (N6413, N6403, N501, N4495, N4893);
nand NAND2 (N6414, N6392, N6354);
buf BUF1 (N6415, N6409);
nor NOR3 (N6416, N6406, N1736, N1311);
xor XOR2 (N6417, N6414, N1926);
nand NAND4 (N6418, N6405, N2056, N4493, N2404);
or OR3 (N6419, N6411, N5734, N3145);
or OR2 (N6420, N6372, N3969);
xor XOR2 (N6421, N6415, N5750);
or OR4 (N6422, N6407, N4059, N6314, N3637);
and AND4 (N6423, N6413, N3697, N4744, N2860);
nor NOR2 (N6424, N6416, N2329);
not NOT1 (N6425, N6424);
buf BUF1 (N6426, N6420);
nand NAND2 (N6427, N6423, N2181);
or OR4 (N6428, N6412, N1795, N2153, N3873);
or OR4 (N6429, N6422, N5277, N6382, N1065);
nor NOR2 (N6430, N6427, N816);
nor NOR3 (N6431, N6430, N5045, N1953);
xor XOR2 (N6432, N6425, N2823);
or OR4 (N6433, N6417, N3890, N2581, N3452);
or OR3 (N6434, N6419, N678, N680);
nand NAND3 (N6435, N6402, N2994, N2993);
not NOT1 (N6436, N6431);
or OR4 (N6437, N6428, N795, N2510, N4709);
buf BUF1 (N6438, N6426);
nand NAND3 (N6439, N6438, N379, N1686);
nor NOR3 (N6440, N6418, N5892, N2275);
and AND3 (N6441, N6439, N5248, N3621);
nor NOR2 (N6442, N6421, N351);
or OR4 (N6443, N6436, N1841, N4534, N3195);
nor NOR2 (N6444, N6441, N3624);
and AND3 (N6445, N6432, N2933, N3069);
xor XOR2 (N6446, N6435, N4065);
nor NOR3 (N6447, N6442, N3018, N3453);
or OR3 (N6448, N6440, N6316, N4333);
xor XOR2 (N6449, N6437, N4460);
not NOT1 (N6450, N6449);
or OR3 (N6451, N6448, N2094, N5230);
or OR3 (N6452, N6433, N1616, N2453);
not NOT1 (N6453, N6451);
buf BUF1 (N6454, N6444);
xor XOR2 (N6455, N6434, N2614);
or OR2 (N6456, N6443, N2441);
buf BUF1 (N6457, N6456);
xor XOR2 (N6458, N6429, N5413);
and AND3 (N6459, N6445, N5040, N6297);
nand NAND3 (N6460, N6459, N5202, N5594);
not NOT1 (N6461, N6460);
or OR2 (N6462, N6453, N6012);
or OR3 (N6463, N6454, N5840, N2206);
not NOT1 (N6464, N6452);
nor NOR3 (N6465, N6450, N5716, N4952);
and AND2 (N6466, N6463, N1222);
nand NAND4 (N6467, N6457, N1042, N3178, N6279);
nand NAND3 (N6468, N6446, N965, N1365);
nand NAND2 (N6469, N6465, N1702);
not NOT1 (N6470, N6467);
nor NOR2 (N6471, N6469, N1289);
buf BUF1 (N6472, N6447);
not NOT1 (N6473, N6471);
nor NOR4 (N6474, N6472, N5102, N1063, N2160);
or OR3 (N6475, N6464, N4351, N3216);
and AND2 (N6476, N6475, N5887);
or OR4 (N6477, N6468, N5240, N6089, N1557);
buf BUF1 (N6478, N6462);
and AND2 (N6479, N6478, N2551);
and AND3 (N6480, N6461, N1879, N4717);
nor NOR3 (N6481, N6474, N2013, N3758);
and AND4 (N6482, N6479, N1931, N1373, N960);
not NOT1 (N6483, N6455);
not NOT1 (N6484, N6458);
or OR3 (N6485, N6466, N132, N3817);
or OR3 (N6486, N6483, N3464, N5483);
xor XOR2 (N6487, N6480, N1285);
nor NOR4 (N6488, N6473, N2239, N386, N6153);
and AND2 (N6489, N6476, N1894);
and AND3 (N6490, N6486, N5369, N4292);
xor XOR2 (N6491, N6489, N3307);
buf BUF1 (N6492, N6477);
nor NOR2 (N6493, N6492, N5305);
and AND2 (N6494, N6485, N615);
nor NOR3 (N6495, N6482, N1551, N5090);
nor NOR4 (N6496, N6484, N3471, N3304, N2737);
not NOT1 (N6497, N6481);
nand NAND2 (N6498, N6495, N1969);
xor XOR2 (N6499, N6488, N2689);
nor NOR3 (N6500, N6491, N4231, N891);
nor NOR4 (N6501, N6470, N27, N1278, N5981);
buf BUF1 (N6502, N6500);
not NOT1 (N6503, N6494);
and AND3 (N6504, N6498, N1473, N3230);
buf BUF1 (N6505, N6504);
buf BUF1 (N6506, N6503);
and AND2 (N6507, N6501, N3718);
buf BUF1 (N6508, N6496);
not NOT1 (N6509, N6507);
buf BUF1 (N6510, N6487);
and AND4 (N6511, N6508, N2566, N4680, N1322);
nor NOR2 (N6512, N6509, N5539);
and AND3 (N6513, N6511, N947, N3642);
nor NOR3 (N6514, N6502, N2936, N4648);
buf BUF1 (N6515, N6505);
buf BUF1 (N6516, N6510);
nor NOR2 (N6517, N6506, N4927);
or OR2 (N6518, N6516, N4942);
xor XOR2 (N6519, N6497, N2219);
or OR3 (N6520, N6515, N6155, N2680);
nand NAND2 (N6521, N6514, N785);
nand NAND3 (N6522, N6499, N4946, N5370);
buf BUF1 (N6523, N6520);
xor XOR2 (N6524, N6493, N442);
nor NOR4 (N6525, N6522, N2167, N4838, N47);
nand NAND3 (N6526, N6490, N1184, N1619);
or OR4 (N6527, N6524, N2880, N2942, N1687);
buf BUF1 (N6528, N6519);
xor XOR2 (N6529, N6517, N3021);
buf BUF1 (N6530, N6512);
buf BUF1 (N6531, N6525);
buf BUF1 (N6532, N6523);
and AND2 (N6533, N6529, N3513);
or OR4 (N6534, N6526, N461, N661, N2560);
nor NOR4 (N6535, N6527, N2419, N5091, N6124);
not NOT1 (N6536, N6513);
xor XOR2 (N6537, N6534, N6389);
buf BUF1 (N6538, N6535);
buf BUF1 (N6539, N6528);
or OR2 (N6540, N6533, N3309);
and AND2 (N6541, N6538, N1602);
and AND3 (N6542, N6540, N145, N5260);
or OR3 (N6543, N6541, N4823, N731);
xor XOR2 (N6544, N6536, N4964);
buf BUF1 (N6545, N6531);
buf BUF1 (N6546, N6545);
xor XOR2 (N6547, N6521, N1274);
nand NAND4 (N6548, N6543, N6345, N3301, N885);
and AND4 (N6549, N6518, N5327, N4218, N152);
not NOT1 (N6550, N6542);
or OR3 (N6551, N6537, N5881, N6341);
and AND3 (N6552, N6549, N401, N3309);
nand NAND4 (N6553, N6547, N2800, N11, N3185);
nand NAND2 (N6554, N6550, N6317);
and AND2 (N6555, N6544, N1749);
and AND4 (N6556, N6552, N4192, N4978, N1325);
and AND2 (N6557, N6556, N6132);
not NOT1 (N6558, N6548);
nand NAND2 (N6559, N6546, N3902);
not NOT1 (N6560, N6530);
buf BUF1 (N6561, N6555);
xor XOR2 (N6562, N6557, N1848);
xor XOR2 (N6563, N6551, N816);
or OR3 (N6564, N6559, N5188, N5774);
and AND4 (N6565, N6561, N5757, N3082, N1572);
xor XOR2 (N6566, N6554, N3698);
nand NAND4 (N6567, N6564, N4974, N1413, N3007);
and AND4 (N6568, N6532, N3571, N4369, N3407);
and AND3 (N6569, N6558, N4721, N5723);
and AND2 (N6570, N6553, N1763);
not NOT1 (N6571, N6569);
buf BUF1 (N6572, N6567);
not NOT1 (N6573, N6572);
nand NAND2 (N6574, N6570, N2485);
or OR2 (N6575, N6562, N910);
and AND4 (N6576, N6575, N6565, N5198, N5361);
and AND3 (N6577, N3419, N5152, N3364);
nand NAND4 (N6578, N6566, N4853, N5422, N1819);
xor XOR2 (N6579, N6573, N5067);
and AND4 (N6580, N6539, N3687, N2740, N558);
or OR3 (N6581, N6571, N3936, N1850);
not NOT1 (N6582, N6579);
and AND4 (N6583, N6574, N5312, N1335, N1971);
nor NOR4 (N6584, N6582, N3658, N1214, N4105);
not NOT1 (N6585, N6568);
not NOT1 (N6586, N6560);
and AND4 (N6587, N6586, N3515, N4100, N5589);
not NOT1 (N6588, N6583);
nor NOR4 (N6589, N6587, N971, N3403, N1659);
xor XOR2 (N6590, N6563, N3498);
buf BUF1 (N6591, N6588);
and AND3 (N6592, N6584, N4540, N5264);
xor XOR2 (N6593, N6580, N5641);
buf BUF1 (N6594, N6581);
not NOT1 (N6595, N6592);
nand NAND4 (N6596, N6576, N4865, N2997, N6049);
xor XOR2 (N6597, N6593, N4739);
nor NOR3 (N6598, N6577, N164, N76);
buf BUF1 (N6599, N6596);
nor NOR4 (N6600, N6590, N4652, N4046, N1335);
xor XOR2 (N6601, N6600, N3675);
nand NAND2 (N6602, N6585, N4899);
not NOT1 (N6603, N6595);
and AND2 (N6604, N6599, N657);
and AND4 (N6605, N6601, N3150, N5845, N2262);
and AND2 (N6606, N6605, N417);
or OR3 (N6607, N6598, N1664, N1526);
buf BUF1 (N6608, N6594);
and AND2 (N6609, N6589, N3269);
xor XOR2 (N6610, N6607, N5208);
not NOT1 (N6611, N6602);
and AND3 (N6612, N6608, N3631, N327);
not NOT1 (N6613, N6591);
nand NAND3 (N6614, N6611, N5742, N677);
nor NOR4 (N6615, N6604, N2082, N1671, N526);
nor NOR4 (N6616, N6603, N1014, N446, N5304);
buf BUF1 (N6617, N6597);
not NOT1 (N6618, N6616);
xor XOR2 (N6619, N6612, N4666);
nor NOR3 (N6620, N6613, N340, N1269);
nor NOR3 (N6621, N6618, N5587, N881);
nor NOR3 (N6622, N6621, N3267, N4002);
and AND2 (N6623, N6617, N1131);
buf BUF1 (N6624, N6606);
buf BUF1 (N6625, N6609);
buf BUF1 (N6626, N6615);
or OR3 (N6627, N6619, N2073, N4363);
nand NAND2 (N6628, N6578, N291);
xor XOR2 (N6629, N6626, N1479);
nand NAND4 (N6630, N6624, N4566, N5308, N208);
and AND3 (N6631, N6629, N3786, N2137);
or OR4 (N6632, N6631, N3051, N5710, N5495);
or OR4 (N6633, N6630, N6386, N1268, N6034);
buf BUF1 (N6634, N6623);
or OR4 (N6635, N6628, N5452, N1418, N3913);
buf BUF1 (N6636, N6632);
nor NOR4 (N6637, N6610, N1551, N2302, N5637);
not NOT1 (N6638, N6633);
buf BUF1 (N6639, N6620);
and AND4 (N6640, N6637, N1338, N440, N3434);
buf BUF1 (N6641, N6627);
xor XOR2 (N6642, N6614, N1613);
and AND4 (N6643, N6625, N4892, N2761, N140);
not NOT1 (N6644, N6622);
nor NOR4 (N6645, N6634, N2039, N4207, N3084);
not NOT1 (N6646, N6640);
nand NAND2 (N6647, N6638, N1079);
nor NOR2 (N6648, N6647, N4062);
nand NAND2 (N6649, N6635, N2211);
and AND2 (N6650, N6648, N327);
nand NAND3 (N6651, N6639, N875, N2451);
xor XOR2 (N6652, N6644, N2115);
or OR4 (N6653, N6652, N2167, N3383, N6453);
nor NOR2 (N6654, N6646, N5622);
buf BUF1 (N6655, N6645);
not NOT1 (N6656, N6649);
or OR2 (N6657, N6654, N917);
nand NAND3 (N6658, N6656, N4464, N3161);
nand NAND4 (N6659, N6658, N5917, N5350, N562);
and AND3 (N6660, N6650, N4900, N5757);
nand NAND2 (N6661, N6659, N2174);
not NOT1 (N6662, N6661);
buf BUF1 (N6663, N6662);
buf BUF1 (N6664, N6636);
not NOT1 (N6665, N6655);
or OR3 (N6666, N6653, N1201, N69);
nand NAND2 (N6667, N6666, N3047);
buf BUF1 (N6668, N6665);
not NOT1 (N6669, N6664);
not NOT1 (N6670, N6643);
nor NOR4 (N6671, N6663, N86, N5385, N5075);
nand NAND2 (N6672, N6642, N720);
buf BUF1 (N6673, N6651);
nand NAND2 (N6674, N6668, N1645);
nand NAND4 (N6675, N6660, N2876, N1013, N3775);
or OR2 (N6676, N6657, N198);
nand NAND3 (N6677, N6676, N4044, N371);
xor XOR2 (N6678, N6672, N3969);
xor XOR2 (N6679, N6674, N2890);
xor XOR2 (N6680, N6667, N249);
nand NAND2 (N6681, N6679, N1647);
buf BUF1 (N6682, N6673);
xor XOR2 (N6683, N6677, N3491);
not NOT1 (N6684, N6671);
nand NAND4 (N6685, N6675, N419, N693, N2354);
nand NAND2 (N6686, N6684, N1191);
not NOT1 (N6687, N6683);
or OR4 (N6688, N6682, N1564, N3411, N5896);
or OR4 (N6689, N6688, N6362, N1366, N1757);
xor XOR2 (N6690, N6687, N5202);
nand NAND2 (N6691, N6670, N174);
nand NAND3 (N6692, N6681, N573, N5953);
nor NOR2 (N6693, N6685, N3012);
and AND4 (N6694, N6692, N822, N3652, N259);
nor NOR2 (N6695, N6686, N1665);
xor XOR2 (N6696, N6641, N1698);
or OR2 (N6697, N6669, N3838);
buf BUF1 (N6698, N6689);
nand NAND2 (N6699, N6693, N902);
nand NAND2 (N6700, N6690, N2936);
or OR2 (N6701, N6695, N561);
and AND2 (N6702, N6691, N3518);
not NOT1 (N6703, N6697);
not NOT1 (N6704, N6703);
xor XOR2 (N6705, N6699, N355);
not NOT1 (N6706, N6702);
or OR4 (N6707, N6706, N6622, N5977, N5534);
and AND2 (N6708, N6701, N6232);
nand NAND2 (N6709, N6698, N3765);
nand NAND3 (N6710, N6678, N6549, N1582);
buf BUF1 (N6711, N6680);
buf BUF1 (N6712, N6709);
nor NOR2 (N6713, N6708, N5696);
buf BUF1 (N6714, N6707);
not NOT1 (N6715, N6710);
or OR3 (N6716, N6696, N2668, N4063);
nand NAND2 (N6717, N6715, N6613);
and AND3 (N6718, N6712, N2766, N2775);
or OR4 (N6719, N6704, N3258, N3784, N5477);
nand NAND3 (N6720, N6700, N6389, N2320);
nor NOR2 (N6721, N6713, N2277);
not NOT1 (N6722, N6711);
nor NOR3 (N6723, N6716, N4726, N2587);
xor XOR2 (N6724, N6722, N1656);
and AND4 (N6725, N6724, N2131, N4490, N6385);
or OR3 (N6726, N6723, N5947, N2256);
nand NAND4 (N6727, N6717, N3337, N4171, N3171);
nand NAND4 (N6728, N6725, N326, N1744, N4540);
not NOT1 (N6729, N6705);
and AND2 (N6730, N6726, N3348);
buf BUF1 (N6731, N6727);
buf BUF1 (N6732, N6728);
buf BUF1 (N6733, N6730);
nand NAND4 (N6734, N6719, N5096, N502, N6184);
nand NAND3 (N6735, N6732, N4918, N5557);
or OR2 (N6736, N6714, N4101);
buf BUF1 (N6737, N6731);
and AND2 (N6738, N6737, N3939);
not NOT1 (N6739, N6736);
buf BUF1 (N6740, N6718);
nand NAND4 (N6741, N6738, N1910, N4766, N1789);
xor XOR2 (N6742, N6735, N4057);
nand NAND3 (N6743, N6721, N2536, N4763);
and AND4 (N6744, N6720, N6555, N6529, N1992);
and AND2 (N6745, N6739, N2568);
and AND2 (N6746, N6729, N1858);
and AND2 (N6747, N6743, N5190);
and AND2 (N6748, N6746, N1407);
or OR2 (N6749, N6741, N6029);
or OR2 (N6750, N6748, N6232);
not NOT1 (N6751, N6734);
or OR3 (N6752, N6749, N2019, N486);
or OR2 (N6753, N6694, N5);
or OR4 (N6754, N6751, N2870, N5687, N5937);
not NOT1 (N6755, N6752);
and AND4 (N6756, N6740, N2377, N5318, N4586);
buf BUF1 (N6757, N6733);
nor NOR3 (N6758, N6742, N4272, N1520);
and AND3 (N6759, N6747, N1689, N3618);
or OR2 (N6760, N6745, N1964);
not NOT1 (N6761, N6754);
nor NOR3 (N6762, N6758, N2802, N442);
xor XOR2 (N6763, N6757, N2054);
and AND2 (N6764, N6756, N2811);
nor NOR4 (N6765, N6763, N2948, N2636, N5934);
or OR4 (N6766, N6760, N535, N3100, N5263);
or OR2 (N6767, N6750, N2756);
buf BUF1 (N6768, N6767);
nand NAND4 (N6769, N6762, N2032, N4652, N5383);
xor XOR2 (N6770, N6769, N3425);
buf BUF1 (N6771, N6761);
nor NOR3 (N6772, N6759, N2671, N214);
nand NAND4 (N6773, N6768, N3716, N4052, N5644);
and AND2 (N6774, N6771, N5950);
and AND4 (N6775, N6755, N3699, N4089, N6536);
nor NOR2 (N6776, N6773, N6409);
not NOT1 (N6777, N6775);
or OR4 (N6778, N6772, N6424, N5798, N1815);
buf BUF1 (N6779, N6766);
not NOT1 (N6780, N6774);
nor NOR2 (N6781, N6764, N440);
buf BUF1 (N6782, N6779);
nand NAND2 (N6783, N6782, N6273);
not NOT1 (N6784, N6780);
not NOT1 (N6785, N6783);
and AND3 (N6786, N6777, N1573, N3040);
buf BUF1 (N6787, N6770);
xor XOR2 (N6788, N6781, N3369);
not NOT1 (N6789, N6776);
nand NAND3 (N6790, N6765, N498, N6282);
not NOT1 (N6791, N6790);
and AND4 (N6792, N6789, N1941, N6546, N3245);
nand NAND4 (N6793, N6791, N6622, N1364, N798);
or OR3 (N6794, N6744, N3492, N788);
xor XOR2 (N6795, N6778, N6415);
nor NOR2 (N6796, N6787, N5642);
buf BUF1 (N6797, N6794);
nand NAND3 (N6798, N6786, N3232, N4075);
buf BUF1 (N6799, N6788);
xor XOR2 (N6800, N6795, N389);
nor NOR4 (N6801, N6797, N3543, N5854, N3834);
or OR3 (N6802, N6784, N4715, N5973);
or OR4 (N6803, N6753, N751, N1774, N4931);
not NOT1 (N6804, N6803);
and AND4 (N6805, N6785, N4164, N5878, N412);
not NOT1 (N6806, N6804);
not NOT1 (N6807, N6800);
and AND3 (N6808, N6799, N5949, N3689);
xor XOR2 (N6809, N6805, N3895);
not NOT1 (N6810, N6802);
and AND2 (N6811, N6810, N6329);
and AND3 (N6812, N6806, N453, N5152);
or OR2 (N6813, N6809, N2109);
xor XOR2 (N6814, N6798, N3552);
xor XOR2 (N6815, N6796, N2328);
or OR4 (N6816, N6801, N5252, N1111, N995);
nand NAND2 (N6817, N6792, N850);
xor XOR2 (N6818, N6813, N1192);
nand NAND3 (N6819, N6811, N4836, N4019);
or OR4 (N6820, N6815, N5810, N4870, N551);
not NOT1 (N6821, N6818);
or OR4 (N6822, N6819, N4064, N1429, N2568);
and AND3 (N6823, N6793, N6201, N3957);
or OR4 (N6824, N6821, N2412, N5048, N945);
or OR3 (N6825, N6817, N5333, N4812);
nand NAND4 (N6826, N6824, N4851, N392, N4536);
nor NOR4 (N6827, N6816, N3093, N5966, N151);
not NOT1 (N6828, N6827);
nor NOR4 (N6829, N6814, N2493, N748, N2429);
or OR2 (N6830, N6826, N4699);
and AND4 (N6831, N6808, N1606, N1203, N6740);
nor NOR2 (N6832, N6828, N4594);
nor NOR4 (N6833, N6822, N1577, N4890, N1710);
or OR2 (N6834, N6812, N5768);
or OR4 (N6835, N6831, N6730, N884, N6355);
not NOT1 (N6836, N6835);
buf BUF1 (N6837, N6807);
nand NAND3 (N6838, N6833, N73, N2181);
nor NOR2 (N6839, N6820, N5634);
not NOT1 (N6840, N6825);
buf BUF1 (N6841, N6839);
or OR4 (N6842, N6836, N4829, N4114, N5629);
xor XOR2 (N6843, N6840, N1292);
nor NOR3 (N6844, N6843, N3589, N5182);
or OR4 (N6845, N6823, N5904, N4909, N1222);
and AND3 (N6846, N6832, N546, N6384);
xor XOR2 (N6847, N6838, N2120);
nand NAND3 (N6848, N6847, N1171, N1716);
nand NAND4 (N6849, N6834, N3477, N3709, N235);
or OR4 (N6850, N6837, N6293, N2303, N3577);
xor XOR2 (N6851, N6829, N290);
buf BUF1 (N6852, N6841);
and AND3 (N6853, N6852, N6438, N144);
xor XOR2 (N6854, N6846, N5610);
nand NAND4 (N6855, N6850, N1818, N3287, N34);
xor XOR2 (N6856, N6845, N939);
or OR3 (N6857, N6853, N1994, N2017);
buf BUF1 (N6858, N6855);
nand NAND4 (N6859, N6851, N2454, N493, N3867);
xor XOR2 (N6860, N6848, N253);
nand NAND2 (N6861, N6844, N6445);
or OR2 (N6862, N6859, N3605);
buf BUF1 (N6863, N6860);
and AND4 (N6864, N6849, N2265, N5867, N1686);
xor XOR2 (N6865, N6854, N6171);
not NOT1 (N6866, N6857);
buf BUF1 (N6867, N6866);
buf BUF1 (N6868, N6861);
xor XOR2 (N6869, N6830, N4742);
buf BUF1 (N6870, N6863);
nand NAND3 (N6871, N6858, N6134, N3355);
not NOT1 (N6872, N6862);
not NOT1 (N6873, N6865);
not NOT1 (N6874, N6867);
nand NAND3 (N6875, N6869, N2048, N6695);
not NOT1 (N6876, N6871);
not NOT1 (N6877, N6876);
or OR4 (N6878, N6874, N4749, N3068, N5763);
nand NAND2 (N6879, N6875, N3999);
or OR2 (N6880, N6842, N1199);
buf BUF1 (N6881, N6872);
nand NAND3 (N6882, N6870, N4019, N1496);
and AND3 (N6883, N6881, N3807, N4281);
nor NOR3 (N6884, N6856, N2421, N1677);
nand NAND3 (N6885, N6878, N1537, N644);
nor NOR4 (N6886, N6864, N936, N1791, N1135);
nand NAND3 (N6887, N6877, N1038, N293);
xor XOR2 (N6888, N6883, N211);
nand NAND2 (N6889, N6868, N1905);
not NOT1 (N6890, N6889);
nor NOR2 (N6891, N6884, N790);
or OR2 (N6892, N6880, N62);
or OR3 (N6893, N6891, N3157, N1156);
buf BUF1 (N6894, N6888);
and AND4 (N6895, N6886, N1863, N5221, N6892);
and AND2 (N6896, N4028, N1264);
nor NOR4 (N6897, N6890, N460, N584, N2302);
xor XOR2 (N6898, N6879, N444);
xor XOR2 (N6899, N6873, N211);
nand NAND4 (N6900, N6885, N3660, N4622, N2941);
xor XOR2 (N6901, N6895, N3176);
nand NAND4 (N6902, N6893, N641, N1722, N3397);
xor XOR2 (N6903, N6894, N623);
xor XOR2 (N6904, N6897, N2203);
and AND4 (N6905, N6904, N6800, N2588, N312);
not NOT1 (N6906, N6896);
nand NAND4 (N6907, N6882, N3748, N1518, N4824);
or OR4 (N6908, N6899, N6127, N100, N1042);
or OR3 (N6909, N6902, N6147, N4548);
nor NOR3 (N6910, N6903, N6097, N6230);
xor XOR2 (N6911, N6910, N1206);
nor NOR3 (N6912, N6900, N4521, N1846);
buf BUF1 (N6913, N6907);
xor XOR2 (N6914, N6912, N2432);
and AND4 (N6915, N6905, N5291, N6052, N6855);
nor NOR2 (N6916, N6915, N2586);
and AND4 (N6917, N6914, N6266, N2183, N6341);
nor NOR3 (N6918, N6906, N3382, N5753);
nand NAND2 (N6919, N6908, N1401);
xor XOR2 (N6920, N6909, N1967);
not NOT1 (N6921, N6913);
xor XOR2 (N6922, N6911, N6617);
and AND4 (N6923, N6921, N1223, N3886, N5614);
nand NAND3 (N6924, N6917, N6706, N5549);
not NOT1 (N6925, N6916);
xor XOR2 (N6926, N6924, N1391);
nor NOR4 (N6927, N6898, N3825, N2533, N3372);
or OR4 (N6928, N6919, N2755, N532, N5118);
nand NAND3 (N6929, N6922, N2293, N4);
not NOT1 (N6930, N6901);
and AND3 (N6931, N6928, N6462, N3308);
nor NOR4 (N6932, N6927, N4778, N2605, N555);
nand NAND4 (N6933, N6920, N3150, N4132, N71);
buf BUF1 (N6934, N6929);
xor XOR2 (N6935, N6934, N1562);
buf BUF1 (N6936, N6931);
xor XOR2 (N6937, N6926, N6678);
buf BUF1 (N6938, N6937);
and AND3 (N6939, N6938, N330, N3460);
not NOT1 (N6940, N6936);
not NOT1 (N6941, N6940);
nand NAND3 (N6942, N6935, N1472, N4926);
xor XOR2 (N6943, N6933, N4164);
not NOT1 (N6944, N6932);
nor NOR4 (N6945, N6942, N1902, N5344, N4608);
or OR3 (N6946, N6945, N6930, N1836);
or OR3 (N6947, N4059, N5341, N4588);
nand NAND2 (N6948, N6939, N6544);
not NOT1 (N6949, N6925);
nor NOR4 (N6950, N6948, N2977, N557, N758);
xor XOR2 (N6951, N6946, N2421);
and AND4 (N6952, N6947, N1923, N6743, N4841);
nor NOR3 (N6953, N6950, N6578, N4921);
and AND4 (N6954, N6943, N6386, N5256, N787);
buf BUF1 (N6955, N6944);
xor XOR2 (N6956, N6923, N1758);
xor XOR2 (N6957, N6953, N4167);
nand NAND3 (N6958, N6949, N1548, N4875);
and AND4 (N6959, N6955, N6716, N1372, N4320);
xor XOR2 (N6960, N6952, N3556);
not NOT1 (N6961, N6957);
xor XOR2 (N6962, N6918, N1071);
and AND2 (N6963, N6961, N4462);
nor NOR3 (N6964, N6958, N1801, N6387);
and AND3 (N6965, N6960, N3672, N1525);
buf BUF1 (N6966, N6964);
buf BUF1 (N6967, N6965);
buf BUF1 (N6968, N6962);
not NOT1 (N6969, N6887);
and AND4 (N6970, N6956, N2932, N3098, N6351);
not NOT1 (N6971, N6959);
nor NOR3 (N6972, N6963, N3164, N5114);
or OR3 (N6973, N6966, N2563, N6612);
or OR2 (N6974, N6941, N6306);
nand NAND4 (N6975, N6973, N2656, N208, N967);
xor XOR2 (N6976, N6974, N4451);
nand NAND3 (N6977, N6975, N5180, N4085);
buf BUF1 (N6978, N6972);
and AND4 (N6979, N6967, N3138, N4284, N6532);
not NOT1 (N6980, N6977);
buf BUF1 (N6981, N6968);
not NOT1 (N6982, N6976);
and AND2 (N6983, N6981, N1050);
and AND2 (N6984, N6982, N4737);
not NOT1 (N6985, N6954);
xor XOR2 (N6986, N6970, N4336);
not NOT1 (N6987, N6951);
nand NAND2 (N6988, N6987, N4091);
xor XOR2 (N6989, N6984, N821);
not NOT1 (N6990, N6983);
buf BUF1 (N6991, N6971);
nand NAND3 (N6992, N6990, N5339, N4628);
xor XOR2 (N6993, N6978, N1450);
or OR3 (N6994, N6969, N3012, N153);
nand NAND4 (N6995, N6988, N6044, N2418, N2940);
nand NAND4 (N6996, N6979, N6577, N4919, N3532);
and AND4 (N6997, N6995, N3360, N4136, N3259);
nand NAND2 (N6998, N6986, N6757);
buf BUF1 (N6999, N6993);
not NOT1 (N7000, N6989);
nor NOR4 (N7001, N6980, N1934, N5982, N3729);
and AND4 (N7002, N6996, N5006, N6902, N3853);
nand NAND4 (N7003, N6985, N1976, N2732, N3208);
nand NAND3 (N7004, N7000, N674, N6940);
not NOT1 (N7005, N6991);
nand NAND4 (N7006, N6992, N6530, N4208, N4797);
not NOT1 (N7007, N6999);
or OR4 (N7008, N7002, N5062, N5953, N3215);
not NOT1 (N7009, N7006);
or OR4 (N7010, N7005, N496, N6078, N3528);
nor NOR4 (N7011, N6997, N1674, N3125, N3226);
not NOT1 (N7012, N7001);
nor NOR4 (N7013, N6998, N1038, N2205, N543);
not NOT1 (N7014, N7009);
and AND3 (N7015, N7010, N4857, N5533);
xor XOR2 (N7016, N7014, N4559);
or OR4 (N7017, N6994, N4642, N2128, N2094);
and AND4 (N7018, N7003, N3122, N5669, N254);
nand NAND2 (N7019, N7018, N493);
or OR4 (N7020, N7004, N3916, N3278, N5697);
nand NAND2 (N7021, N7007, N6497);
not NOT1 (N7022, N7017);
and AND3 (N7023, N7011, N6843, N1180);
nor NOR3 (N7024, N7008, N2881, N4306);
and AND2 (N7025, N7024, N2271);
or OR3 (N7026, N7013, N1454, N3060);
nand NAND4 (N7027, N7020, N2892, N4429, N6141);
or OR4 (N7028, N7023, N1049, N79, N6581);
nor NOR2 (N7029, N7025, N239);
or OR4 (N7030, N7019, N5506, N5664, N5407);
or OR3 (N7031, N7016, N6053, N3017);
xor XOR2 (N7032, N7027, N5987);
not NOT1 (N7033, N7032);
xor XOR2 (N7034, N7026, N2865);
buf BUF1 (N7035, N7029);
or OR2 (N7036, N7028, N4425);
or OR2 (N7037, N7036, N4910);
or OR3 (N7038, N7034, N489, N3181);
xor XOR2 (N7039, N7038, N1768);
nor NOR4 (N7040, N7035, N6110, N2753, N6938);
not NOT1 (N7041, N7033);
or OR3 (N7042, N7015, N6548, N2502);
xor XOR2 (N7043, N7021, N1390);
not NOT1 (N7044, N7022);
buf BUF1 (N7045, N7039);
or OR2 (N7046, N7045, N638);
nor NOR4 (N7047, N7042, N5972, N5637, N1129);
buf BUF1 (N7048, N7040);
not NOT1 (N7049, N7031);
not NOT1 (N7050, N7030);
or OR2 (N7051, N7037, N3865);
not NOT1 (N7052, N7046);
xor XOR2 (N7053, N7052, N5401);
xor XOR2 (N7054, N7049, N2852);
nor NOR3 (N7055, N7051, N6276, N6419);
buf BUF1 (N7056, N7050);
or OR3 (N7057, N7047, N2553, N874);
xor XOR2 (N7058, N7053, N3070);
and AND4 (N7059, N7056, N6099, N5706, N3003);
nor NOR2 (N7060, N7059, N950);
or OR2 (N7061, N7060, N6182);
or OR4 (N7062, N7061, N3997, N5972, N2508);
and AND2 (N7063, N7012, N1483);
not NOT1 (N7064, N7063);
nand NAND3 (N7065, N7058, N1762, N2477);
not NOT1 (N7066, N7062);
buf BUF1 (N7067, N7065);
and AND2 (N7068, N7057, N5750);
not NOT1 (N7069, N7041);
and AND4 (N7070, N7064, N4295, N4051, N3600);
nand NAND2 (N7071, N7068, N5811);
and AND2 (N7072, N7069, N4145);
nor NOR4 (N7073, N7066, N4989, N6607, N1003);
xor XOR2 (N7074, N7070, N3389);
or OR2 (N7075, N7073, N6592);
not NOT1 (N7076, N7055);
not NOT1 (N7077, N7074);
xor XOR2 (N7078, N7071, N2107);
not NOT1 (N7079, N7078);
and AND2 (N7080, N7067, N6587);
nand NAND3 (N7081, N7080, N862, N3607);
buf BUF1 (N7082, N7054);
and AND4 (N7083, N7075, N1685, N4442, N4392);
nor NOR2 (N7084, N7043, N5423);
buf BUF1 (N7085, N7084);
and AND4 (N7086, N7081, N5217, N1577, N1700);
buf BUF1 (N7087, N7085);
or OR3 (N7088, N7082, N5784, N4050);
and AND3 (N7089, N7076, N1727, N2875);
and AND2 (N7090, N7044, N4045);
xor XOR2 (N7091, N7090, N3224);
buf BUF1 (N7092, N7088);
or OR4 (N7093, N7079, N3608, N6499, N5157);
or OR3 (N7094, N7093, N4497, N6814);
not NOT1 (N7095, N7094);
or OR2 (N7096, N7086, N2593);
not NOT1 (N7097, N7096);
nand NAND3 (N7098, N7095, N5047, N468);
not NOT1 (N7099, N7077);
not NOT1 (N7100, N7072);
nor NOR3 (N7101, N7091, N6453, N1943);
xor XOR2 (N7102, N7092, N2945);
buf BUF1 (N7103, N7089);
xor XOR2 (N7104, N7083, N6950);
xor XOR2 (N7105, N7048, N5451);
buf BUF1 (N7106, N7100);
not NOT1 (N7107, N7103);
nor NOR4 (N7108, N7102, N1974, N3368, N6425);
nor NOR4 (N7109, N7101, N1006, N3198, N5972);
buf BUF1 (N7110, N7106);
and AND3 (N7111, N7107, N6533, N2037);
nand NAND4 (N7112, N7098, N3562, N1309, N701);
buf BUF1 (N7113, N7108);
xor XOR2 (N7114, N7099, N1138);
buf BUF1 (N7115, N7110);
not NOT1 (N7116, N7087);
nor NOR4 (N7117, N7112, N4300, N6694, N296);
xor XOR2 (N7118, N7111, N1227);
nor NOR2 (N7119, N7117, N977);
and AND4 (N7120, N7097, N908, N4119, N1470);
or OR4 (N7121, N7104, N2108, N6790, N4977);
not NOT1 (N7122, N7113);
nand NAND3 (N7123, N7105, N5302, N5840);
and AND3 (N7124, N7116, N5469, N7081);
not NOT1 (N7125, N7118);
nand NAND4 (N7126, N7122, N5684, N56, N729);
xor XOR2 (N7127, N7124, N4416);
nor NOR4 (N7128, N7126, N3326, N2572, N1631);
buf BUF1 (N7129, N7128);
buf BUF1 (N7130, N7129);
not NOT1 (N7131, N7114);
xor XOR2 (N7132, N7131, N1665);
buf BUF1 (N7133, N7130);
not NOT1 (N7134, N7133);
or OR2 (N7135, N7119, N1300);
not NOT1 (N7136, N7125);
not NOT1 (N7137, N7127);
nor NOR3 (N7138, N7136, N1938, N4244);
and AND3 (N7139, N7121, N3178, N2501);
and AND2 (N7140, N7132, N6245);
xor XOR2 (N7141, N7137, N75);
not NOT1 (N7142, N7109);
and AND2 (N7143, N7115, N3340);
buf BUF1 (N7144, N7134);
nand NAND3 (N7145, N7138, N5351, N5529);
xor XOR2 (N7146, N7143, N2602);
and AND4 (N7147, N7120, N3683, N3508, N2790);
and AND4 (N7148, N7135, N5519, N3735, N526);
and AND4 (N7149, N7146, N4795, N4061, N6553);
nand NAND3 (N7150, N7149, N2636, N6676);
and AND3 (N7151, N7139, N1096, N6402);
buf BUF1 (N7152, N7140);
xor XOR2 (N7153, N7144, N743);
or OR2 (N7154, N7150, N4025);
nand NAND2 (N7155, N7123, N279);
buf BUF1 (N7156, N7142);
not NOT1 (N7157, N7151);
buf BUF1 (N7158, N7147);
nor NOR2 (N7159, N7152, N906);
nand NAND2 (N7160, N7153, N4573);
nand NAND4 (N7161, N7160, N4401, N256, N6459);
nand NAND2 (N7162, N7161, N5489);
nand NAND4 (N7163, N7141, N3998, N5556, N1279);
not NOT1 (N7164, N7159);
nor NOR2 (N7165, N7154, N4920);
and AND2 (N7166, N7156, N1301);
or OR3 (N7167, N7162, N6573, N6994);
or OR3 (N7168, N7164, N6641, N3932);
or OR4 (N7169, N7163, N6858, N5671, N226);
not NOT1 (N7170, N7167);
buf BUF1 (N7171, N7169);
not NOT1 (N7172, N7155);
or OR2 (N7173, N7157, N6177);
not NOT1 (N7174, N7172);
or OR3 (N7175, N7171, N2243, N448);
nand NAND4 (N7176, N7175, N6677, N533, N2279);
nor NOR3 (N7177, N7148, N1035, N5314);
buf BUF1 (N7178, N7174);
nand NAND3 (N7179, N7168, N2959, N1762);
xor XOR2 (N7180, N7178, N3486);
nor NOR4 (N7181, N7180, N1491, N4337, N6015);
and AND3 (N7182, N7179, N6122, N5966);
nor NOR3 (N7183, N7165, N6577, N6646);
not NOT1 (N7184, N7158);
nor NOR4 (N7185, N7170, N1593, N381, N2961);
and AND3 (N7186, N7184, N6800, N2820);
or OR4 (N7187, N7166, N6640, N2092, N1213);
or OR2 (N7188, N7176, N2577);
buf BUF1 (N7189, N7182);
xor XOR2 (N7190, N7181, N2574);
not NOT1 (N7191, N7145);
and AND2 (N7192, N7185, N2511);
or OR3 (N7193, N7187, N6348, N5258);
buf BUF1 (N7194, N7190);
and AND2 (N7195, N7188, N6387);
nor NOR2 (N7196, N7193, N4979);
nor NOR2 (N7197, N7192, N5983);
not NOT1 (N7198, N7195);
or OR3 (N7199, N7186, N6443, N3147);
not NOT1 (N7200, N7183);
or OR2 (N7201, N7177, N574);
nand NAND3 (N7202, N7197, N2078, N3642);
and AND2 (N7203, N7189, N335);
nand NAND4 (N7204, N7201, N6594, N5817, N6152);
nor NOR3 (N7205, N7191, N3988, N2598);
not NOT1 (N7206, N7200);
buf BUF1 (N7207, N7199);
nand NAND4 (N7208, N7207, N5984, N4734, N7015);
not NOT1 (N7209, N7208);
xor XOR2 (N7210, N7209, N6953);
not NOT1 (N7211, N7202);
buf BUF1 (N7212, N7206);
and AND2 (N7213, N7204, N3009);
not NOT1 (N7214, N7198);
and AND3 (N7215, N7211, N6449, N2327);
and AND2 (N7216, N7173, N5641);
not NOT1 (N7217, N7196);
nand NAND2 (N7218, N7215, N7120);
buf BUF1 (N7219, N7212);
or OR2 (N7220, N7194, N811);
and AND4 (N7221, N7218, N2095, N1044, N5325);
xor XOR2 (N7222, N7216, N707);
nand NAND2 (N7223, N7221, N3569);
or OR4 (N7224, N7214, N3614, N3934, N6415);
not NOT1 (N7225, N7219);
not NOT1 (N7226, N7217);
nand NAND3 (N7227, N7222, N1626, N357);
and AND4 (N7228, N7205, N1044, N348, N687);
xor XOR2 (N7229, N7213, N2505);
or OR4 (N7230, N7225, N557, N4963, N2145);
not NOT1 (N7231, N7227);
nand NAND3 (N7232, N7226, N4106, N2473);
buf BUF1 (N7233, N7231);
or OR3 (N7234, N7233, N3339, N5391);
xor XOR2 (N7235, N7203, N3385);
xor XOR2 (N7236, N7235, N3968);
xor XOR2 (N7237, N7224, N3335);
nand NAND3 (N7238, N7236, N1288, N4118);
not NOT1 (N7239, N7220);
or OR2 (N7240, N7210, N5986);
and AND3 (N7241, N7237, N5679, N6288);
nand NAND3 (N7242, N7232, N5951, N6564);
or OR3 (N7243, N7234, N3164, N3768);
not NOT1 (N7244, N7223);
nand NAND4 (N7245, N7242, N2282, N1954, N6771);
nand NAND4 (N7246, N7229, N2786, N305, N553);
buf BUF1 (N7247, N7228);
buf BUF1 (N7248, N7239);
buf BUF1 (N7249, N7247);
or OR3 (N7250, N7245, N7062, N3986);
and AND2 (N7251, N7241, N2392);
or OR4 (N7252, N7243, N6313, N2169, N322);
or OR2 (N7253, N7251, N5722);
or OR4 (N7254, N7248, N267, N3883, N5432);
and AND4 (N7255, N7230, N7205, N2149, N1794);
nor NOR3 (N7256, N7255, N6901, N5403);
or OR4 (N7257, N7250, N1220, N4692, N2255);
and AND2 (N7258, N7257, N614);
nor NOR2 (N7259, N7244, N750);
and AND4 (N7260, N7256, N5969, N5717, N7035);
not NOT1 (N7261, N7259);
and AND2 (N7262, N7253, N1499);
not NOT1 (N7263, N7254);
nor NOR3 (N7264, N7262, N3702, N4211);
buf BUF1 (N7265, N7246);
not NOT1 (N7266, N7252);
buf BUF1 (N7267, N7261);
and AND2 (N7268, N7249, N6737);
nor NOR2 (N7269, N7264, N4714);
or OR3 (N7270, N7238, N2697, N3205);
nand NAND4 (N7271, N7266, N2075, N3730, N3338);
nand NAND3 (N7272, N7268, N5496, N1886);
xor XOR2 (N7273, N7263, N2319);
not NOT1 (N7274, N7260);
and AND3 (N7275, N7274, N1314, N7124);
nor NOR2 (N7276, N7270, N5023);
xor XOR2 (N7277, N7258, N2099);
and AND3 (N7278, N7269, N3377, N1703);
and AND4 (N7279, N7267, N1621, N300, N1503);
buf BUF1 (N7280, N7240);
nand NAND3 (N7281, N7277, N6313, N2969);
buf BUF1 (N7282, N7273);
buf BUF1 (N7283, N7271);
not NOT1 (N7284, N7275);
not NOT1 (N7285, N7284);
not NOT1 (N7286, N7278);
nor NOR4 (N7287, N7276, N954, N4819, N1454);
nor NOR3 (N7288, N7280, N2325, N558);
or OR3 (N7289, N7272, N1527, N7172);
and AND3 (N7290, N7286, N2376, N6115);
buf BUF1 (N7291, N7285);
or OR2 (N7292, N7291, N6783);
xor XOR2 (N7293, N7288, N6428);
and AND4 (N7294, N7287, N6132, N5377, N5074);
not NOT1 (N7295, N7293);
xor XOR2 (N7296, N7290, N4561);
nor NOR4 (N7297, N7281, N478, N43, N5093);
nand NAND4 (N7298, N7295, N4307, N590, N187);
xor XOR2 (N7299, N7283, N5917);
nor NOR3 (N7300, N7297, N6599, N7173);
xor XOR2 (N7301, N7282, N2179);
nand NAND2 (N7302, N7289, N5748);
xor XOR2 (N7303, N7296, N6203);
xor XOR2 (N7304, N7299, N2153);
xor XOR2 (N7305, N7302, N5058);
buf BUF1 (N7306, N7305);
nor NOR3 (N7307, N7279, N6729, N3575);
not NOT1 (N7308, N7303);
xor XOR2 (N7309, N7308, N6597);
xor XOR2 (N7310, N7304, N2905);
nor NOR2 (N7311, N7300, N1581);
or OR3 (N7312, N7298, N2885, N1427);
buf BUF1 (N7313, N7311);
not NOT1 (N7314, N7306);
xor XOR2 (N7315, N7313, N5476);
xor XOR2 (N7316, N7309, N6559);
not NOT1 (N7317, N7314);
and AND3 (N7318, N7316, N2684, N667);
buf BUF1 (N7319, N7312);
or OR4 (N7320, N7307, N4715, N4508, N2750);
not NOT1 (N7321, N7319);
nand NAND4 (N7322, N7294, N5734, N5598, N2550);
buf BUF1 (N7323, N7322);
not NOT1 (N7324, N7321);
nor NOR2 (N7325, N7315, N1158);
and AND4 (N7326, N7318, N1719, N1791, N4241);
or OR2 (N7327, N7292, N756);
nand NAND3 (N7328, N7317, N5080, N695);
nor NOR4 (N7329, N7301, N1054, N6939, N5394);
and AND3 (N7330, N7325, N2206, N532);
not NOT1 (N7331, N7324);
and AND4 (N7332, N7326, N658, N1092, N693);
buf BUF1 (N7333, N7328);
xor XOR2 (N7334, N7332, N2825);
buf BUF1 (N7335, N7310);
not NOT1 (N7336, N7330);
or OR4 (N7337, N7333, N3104, N5661, N2019);
nor NOR2 (N7338, N7331, N554);
nor NOR4 (N7339, N7336, N966, N4645, N2292);
buf BUF1 (N7340, N7338);
and AND3 (N7341, N7323, N3053, N5124);
or OR4 (N7342, N7340, N5056, N6908, N616);
or OR3 (N7343, N7329, N4199, N3126);
nand NAND3 (N7344, N7339, N2983, N147);
nand NAND4 (N7345, N7334, N2973, N5916, N1060);
or OR3 (N7346, N7344, N6010, N5424);
nor NOR4 (N7347, N7341, N1357, N1714, N6229);
and AND2 (N7348, N7345, N3956);
xor XOR2 (N7349, N7343, N3701);
not NOT1 (N7350, N7342);
nand NAND4 (N7351, N7265, N6771, N3892, N3338);
and AND2 (N7352, N7320, N1103);
xor XOR2 (N7353, N7349, N6963);
or OR3 (N7354, N7337, N5506, N4755);
and AND4 (N7355, N7346, N6885, N965, N75);
not NOT1 (N7356, N7352);
not NOT1 (N7357, N7347);
nand NAND2 (N7358, N7348, N5436);
not NOT1 (N7359, N7353);
buf BUF1 (N7360, N7355);
xor XOR2 (N7361, N7351, N6509);
buf BUF1 (N7362, N7361);
nor NOR2 (N7363, N7358, N1680);
or OR3 (N7364, N7360, N4425, N4585);
and AND3 (N7365, N7327, N443, N173);
or OR2 (N7366, N7354, N3827);
nand NAND4 (N7367, N7357, N4464, N6376, N113);
xor XOR2 (N7368, N7367, N4843);
nor NOR2 (N7369, N7368, N1282);
buf BUF1 (N7370, N7362);
nor NOR4 (N7371, N7335, N6298, N1168, N167);
nor NOR4 (N7372, N7366, N2412, N2412, N1829);
not NOT1 (N7373, N7370);
and AND2 (N7374, N7364, N6488);
and AND4 (N7375, N7374, N6403, N3278, N2823);
and AND3 (N7376, N7350, N1761, N5341);
and AND2 (N7377, N7359, N2995);
nand NAND3 (N7378, N7369, N2369, N3479);
not NOT1 (N7379, N7356);
xor XOR2 (N7380, N7376, N2905);
and AND2 (N7381, N7363, N2);
nor NOR3 (N7382, N7377, N6868, N816);
buf BUF1 (N7383, N7380);
buf BUF1 (N7384, N7382);
and AND2 (N7385, N7384, N5333);
and AND2 (N7386, N7385, N1308);
xor XOR2 (N7387, N7371, N4205);
and AND2 (N7388, N7379, N6468);
or OR2 (N7389, N7375, N2648);
or OR3 (N7390, N7372, N2610, N679);
nand NAND2 (N7391, N7387, N1846);
nand NAND3 (N7392, N7390, N427, N2012);
and AND2 (N7393, N7392, N336);
not NOT1 (N7394, N7388);
nand NAND3 (N7395, N7386, N1625, N3496);
and AND2 (N7396, N7378, N2091);
not NOT1 (N7397, N7373);
buf BUF1 (N7398, N7381);
and AND3 (N7399, N7393, N296, N6787);
nand NAND3 (N7400, N7389, N1230, N3280);
or OR4 (N7401, N7394, N1242, N1362, N1668);
not NOT1 (N7402, N7396);
and AND2 (N7403, N7401, N2358);
nand NAND3 (N7404, N7395, N5507, N3891);
buf BUF1 (N7405, N7403);
nor NOR4 (N7406, N7391, N6050, N2964, N2863);
xor XOR2 (N7407, N7398, N1168);
or OR2 (N7408, N7402, N1908);
buf BUF1 (N7409, N7407);
buf BUF1 (N7410, N7409);
nand NAND2 (N7411, N7399, N3357);
nand NAND4 (N7412, N7411, N270, N3787, N4492);
xor XOR2 (N7413, N7397, N5001);
not NOT1 (N7414, N7404);
or OR4 (N7415, N7412, N1315, N4908, N745);
nand NAND4 (N7416, N7415, N1205, N3757, N4293);
and AND4 (N7417, N7414, N2206, N4252, N4645);
or OR4 (N7418, N7365, N5641, N6587, N2218);
not NOT1 (N7419, N7400);
or OR2 (N7420, N7405, N922);
nor NOR4 (N7421, N7417, N245, N3515, N5961);
not NOT1 (N7422, N7406);
not NOT1 (N7423, N7408);
nor NOR3 (N7424, N7418, N39, N6638);
nor NOR4 (N7425, N7420, N5666, N3888, N6259);
buf BUF1 (N7426, N7423);
buf BUF1 (N7427, N7424);
or OR2 (N7428, N7421, N3758);
xor XOR2 (N7429, N7427, N3918);
nand NAND3 (N7430, N7413, N5261, N1635);
or OR4 (N7431, N7429, N4802, N6894, N5302);
xor XOR2 (N7432, N7419, N4036);
nand NAND3 (N7433, N7422, N6280, N2717);
or OR2 (N7434, N7416, N915);
nor NOR3 (N7435, N7383, N4952, N192);
nand NAND3 (N7436, N7425, N1314, N2160);
and AND3 (N7437, N7426, N6971, N1805);
nor NOR4 (N7438, N7437, N6657, N7213, N4313);
or OR3 (N7439, N7428, N931, N6116);
nor NOR4 (N7440, N7433, N5845, N3087, N2998);
nand NAND4 (N7441, N7410, N7163, N1943, N1517);
not NOT1 (N7442, N7440);
buf BUF1 (N7443, N7432);
and AND4 (N7444, N7439, N339, N491, N6168);
nor NOR4 (N7445, N7435, N1709, N1650, N5546);
nor NOR2 (N7446, N7436, N6094);
buf BUF1 (N7447, N7445);
buf BUF1 (N7448, N7430);
or OR4 (N7449, N7443, N565, N1716, N3008);
nor NOR4 (N7450, N7449, N691, N5588, N1579);
nand NAND3 (N7451, N7447, N6910, N3775);
nand NAND3 (N7452, N7441, N1993, N1786);
not NOT1 (N7453, N7434);
and AND3 (N7454, N7451, N1120, N3682);
or OR4 (N7455, N7446, N4142, N5502, N3492);
not NOT1 (N7456, N7453);
nand NAND3 (N7457, N7431, N5898, N5963);
buf BUF1 (N7458, N7438);
nand NAND3 (N7459, N7454, N1645, N4676);
nand NAND2 (N7460, N7448, N248);
nand NAND4 (N7461, N7460, N5157, N648, N6498);
not NOT1 (N7462, N7459);
not NOT1 (N7463, N7442);
buf BUF1 (N7464, N7458);
nor NOR4 (N7465, N7452, N2837, N6077, N4188);
nor NOR3 (N7466, N7444, N5583, N2093);
nand NAND3 (N7467, N7462, N141, N2930);
nor NOR2 (N7468, N7457, N1906);
nor NOR4 (N7469, N7465, N4428, N2935, N4501);
nand NAND2 (N7470, N7456, N4885);
xor XOR2 (N7471, N7467, N4080);
not NOT1 (N7472, N7469);
buf BUF1 (N7473, N7468);
nor NOR4 (N7474, N7472, N3569, N1663, N3035);
nand NAND3 (N7475, N7470, N5615, N6244);
and AND3 (N7476, N7461, N2928, N1707);
nor NOR4 (N7477, N7476, N6075, N166, N4456);
not NOT1 (N7478, N7450);
and AND2 (N7479, N7473, N700);
nand NAND4 (N7480, N7474, N5553, N503, N5162);
not NOT1 (N7481, N7475);
nor NOR2 (N7482, N7481, N1862);
or OR3 (N7483, N7463, N4866, N6304);
nand NAND3 (N7484, N7480, N2507, N7024);
buf BUF1 (N7485, N7478);
or OR3 (N7486, N7471, N1491, N732);
nand NAND2 (N7487, N7479, N4474);
or OR2 (N7488, N7485, N2910);
not NOT1 (N7489, N7488);
buf BUF1 (N7490, N7482);
buf BUF1 (N7491, N7486);
nor NOR4 (N7492, N7483, N6897, N2873, N7171);
or OR4 (N7493, N7490, N3384, N2871, N2865);
not NOT1 (N7494, N7464);
or OR3 (N7495, N7477, N1775, N4630);
buf BUF1 (N7496, N7493);
buf BUF1 (N7497, N7455);
buf BUF1 (N7498, N7492);
not NOT1 (N7499, N7495);
buf BUF1 (N7500, N7484);
nand NAND3 (N7501, N7500, N2480, N7217);
nand NAND3 (N7502, N7494, N2262, N4584);
nand NAND2 (N7503, N7497, N993);
and AND3 (N7504, N7501, N2510, N5700);
nor NOR3 (N7505, N7489, N5837, N807);
nand NAND4 (N7506, N7487, N167, N706, N1201);
and AND3 (N7507, N7502, N5367, N5002);
and AND2 (N7508, N7491, N4689);
xor XOR2 (N7509, N7496, N5393);
nand NAND2 (N7510, N7508, N6333);
not NOT1 (N7511, N7510);
or OR4 (N7512, N7509, N4943, N6680, N6988);
not NOT1 (N7513, N7507);
and AND2 (N7514, N7504, N4655);
xor XOR2 (N7515, N7514, N6541);
nor NOR3 (N7516, N7498, N1357, N3719);
or OR4 (N7517, N7506, N4005, N3123, N3413);
or OR4 (N7518, N7505, N1109, N1084, N6320);
xor XOR2 (N7519, N7511, N4698);
buf BUF1 (N7520, N7512);
buf BUF1 (N7521, N7516);
and AND3 (N7522, N7519, N912, N6020);
nand NAND4 (N7523, N7517, N2313, N3031, N1715);
and AND4 (N7524, N7523, N5127, N2251, N651);
not NOT1 (N7525, N7520);
nor NOR4 (N7526, N7525, N4436, N3213, N26);
and AND2 (N7527, N7521, N2358);
nand NAND3 (N7528, N7524, N5613, N3291);
nand NAND2 (N7529, N7528, N3941);
not NOT1 (N7530, N7526);
xor XOR2 (N7531, N7466, N2394);
nor NOR4 (N7532, N7529, N6794, N6312, N5956);
not NOT1 (N7533, N7530);
not NOT1 (N7534, N7531);
and AND2 (N7535, N7515, N2586);
and AND3 (N7536, N7513, N2180, N4653);
buf BUF1 (N7537, N7518);
buf BUF1 (N7538, N7527);
buf BUF1 (N7539, N7522);
or OR3 (N7540, N7536, N995, N1657);
not NOT1 (N7541, N7534);
or OR4 (N7542, N7538, N376, N1526, N1740);
buf BUF1 (N7543, N7533);
buf BUF1 (N7544, N7499);
nor NOR2 (N7545, N7537, N4671);
not NOT1 (N7546, N7544);
xor XOR2 (N7547, N7541, N5183);
xor XOR2 (N7548, N7546, N1338);
nand NAND4 (N7549, N7540, N6503, N3610, N6063);
not NOT1 (N7550, N7543);
and AND4 (N7551, N7550, N789, N2983, N2466);
nor NOR2 (N7552, N7548, N4580);
buf BUF1 (N7553, N7549);
not NOT1 (N7554, N7542);
nor NOR3 (N7555, N7547, N5999, N5289);
and AND2 (N7556, N7554, N5856);
not NOT1 (N7557, N7551);
nor NOR4 (N7558, N7535, N4980, N3037, N2816);
and AND4 (N7559, N7558, N6633, N718, N3127);
nand NAND3 (N7560, N7555, N3854, N6957);
and AND2 (N7561, N7553, N821);
and AND2 (N7562, N7539, N5480);
buf BUF1 (N7563, N7557);
and AND2 (N7564, N7559, N5573);
xor XOR2 (N7565, N7503, N5847);
not NOT1 (N7566, N7560);
nor NOR3 (N7567, N7545, N6177, N1106);
buf BUF1 (N7568, N7563);
not NOT1 (N7569, N7562);
nor NOR3 (N7570, N7532, N2582, N6252);
and AND4 (N7571, N7569, N4421, N4832, N427);
nand NAND2 (N7572, N7571, N5367);
nor NOR2 (N7573, N7556, N7034);
nand NAND4 (N7574, N7565, N4259, N2344, N3407);
and AND4 (N7575, N7564, N1190, N1859, N1228);
or OR3 (N7576, N7561, N6199, N1643);
or OR3 (N7577, N7574, N754, N820);
xor XOR2 (N7578, N7566, N504);
xor XOR2 (N7579, N7572, N4383);
nor NOR3 (N7580, N7579, N5334, N153);
or OR4 (N7581, N7575, N6458, N3045, N2410);
and AND4 (N7582, N7581, N575, N3205, N2828);
nand NAND3 (N7583, N7573, N3954, N2712);
nor NOR3 (N7584, N7578, N3982, N1833);
nand NAND3 (N7585, N7577, N4279, N4595);
or OR4 (N7586, N7584, N6309, N4335, N2495);
or OR2 (N7587, N7570, N1560);
and AND3 (N7588, N7580, N7011, N709);
nand NAND3 (N7589, N7568, N5535, N6709);
xor XOR2 (N7590, N7589, N4288);
nor NOR3 (N7591, N7583, N6728, N215);
nor NOR3 (N7592, N7588, N7201, N4328);
buf BUF1 (N7593, N7590);
xor XOR2 (N7594, N7593, N2998);
and AND4 (N7595, N7567, N1707, N266, N5611);
xor XOR2 (N7596, N7591, N7570);
nor NOR4 (N7597, N7596, N4456, N6800, N7527);
and AND4 (N7598, N7595, N7306, N4071, N4066);
nand NAND4 (N7599, N7586, N1124, N5297, N6897);
xor XOR2 (N7600, N7594, N3631);
xor XOR2 (N7601, N7598, N140);
nor NOR3 (N7602, N7599, N7368, N235);
nand NAND3 (N7603, N7601, N7377, N5290);
and AND3 (N7604, N7597, N725, N6530);
not NOT1 (N7605, N7576);
and AND2 (N7606, N7600, N6234);
buf BUF1 (N7607, N7552);
and AND3 (N7608, N7605, N165, N4330);
not NOT1 (N7609, N7602);
nor NOR4 (N7610, N7582, N3488, N6489, N1195);
nand NAND2 (N7611, N7610, N6710);
nand NAND2 (N7612, N7611, N1258);
not NOT1 (N7613, N7607);
xor XOR2 (N7614, N7606, N2655);
not NOT1 (N7615, N7587);
buf BUF1 (N7616, N7585);
buf BUF1 (N7617, N7614);
buf BUF1 (N7618, N7615);
buf BUF1 (N7619, N7617);
nor NOR2 (N7620, N7609, N966);
not NOT1 (N7621, N7592);
not NOT1 (N7622, N7618);
buf BUF1 (N7623, N7622);
or OR2 (N7624, N7603, N4633);
not NOT1 (N7625, N7612);
or OR4 (N7626, N7619, N941, N7039, N7258);
not NOT1 (N7627, N7625);
nor NOR2 (N7628, N7624, N276);
and AND2 (N7629, N7627, N1901);
not NOT1 (N7630, N7628);
nand NAND2 (N7631, N7608, N3660);
and AND3 (N7632, N7620, N6272, N4620);
or OR3 (N7633, N7630, N3880, N3702);
and AND4 (N7634, N7629, N4526, N401, N7510);
nor NOR2 (N7635, N7634, N1967);
nor NOR3 (N7636, N7616, N3714, N1020);
buf BUF1 (N7637, N7604);
nand NAND2 (N7638, N7623, N7044);
nand NAND2 (N7639, N7635, N953);
not NOT1 (N7640, N7613);
buf BUF1 (N7641, N7632);
and AND3 (N7642, N7639, N5747, N688);
nand NAND3 (N7643, N7626, N6460, N5304);
buf BUF1 (N7644, N7633);
nand NAND2 (N7645, N7644, N6287);
nand NAND3 (N7646, N7640, N1275, N6243);
or OR3 (N7647, N7638, N7492, N2856);
or OR2 (N7648, N7641, N7417);
buf BUF1 (N7649, N7647);
not NOT1 (N7650, N7642);
not NOT1 (N7651, N7621);
or OR2 (N7652, N7651, N5195);
nor NOR2 (N7653, N7636, N3874);
buf BUF1 (N7654, N7645);
or OR3 (N7655, N7646, N5579, N4238);
xor XOR2 (N7656, N7643, N2500);
xor XOR2 (N7657, N7656, N7254);
not NOT1 (N7658, N7650);
xor XOR2 (N7659, N7631, N6335);
and AND4 (N7660, N7659, N336, N2153, N7645);
xor XOR2 (N7661, N7652, N5360);
nand NAND4 (N7662, N7637, N3178, N4222, N2946);
and AND4 (N7663, N7653, N4491, N1355, N6733);
and AND4 (N7664, N7657, N3042, N1178, N7556);
buf BUF1 (N7665, N7658);
nor NOR2 (N7666, N7662, N4387);
not NOT1 (N7667, N7663);
xor XOR2 (N7668, N7655, N6794);
not NOT1 (N7669, N7649);
buf BUF1 (N7670, N7669);
nand NAND3 (N7671, N7661, N1648, N1006);
nor NOR3 (N7672, N7654, N3774, N5037);
nand NAND3 (N7673, N7648, N6838, N1267);
nand NAND3 (N7674, N7670, N2661, N1102);
xor XOR2 (N7675, N7666, N5925);
nand NAND3 (N7676, N7660, N7243, N6252);
buf BUF1 (N7677, N7676);
buf BUF1 (N7678, N7674);
not NOT1 (N7679, N7675);
nand NAND3 (N7680, N7664, N2113, N2816);
nor NOR2 (N7681, N7677, N5536);
buf BUF1 (N7682, N7671);
not NOT1 (N7683, N7667);
nand NAND2 (N7684, N7679, N6602);
not NOT1 (N7685, N7684);
buf BUF1 (N7686, N7678);
xor XOR2 (N7687, N7685, N1859);
or OR2 (N7688, N7668, N7167);
not NOT1 (N7689, N7680);
xor XOR2 (N7690, N7681, N675);
nor NOR2 (N7691, N7688, N5735);
buf BUF1 (N7692, N7689);
or OR3 (N7693, N7691, N1830, N2861);
xor XOR2 (N7694, N7693, N7465);
xor XOR2 (N7695, N7690, N4310);
nor NOR2 (N7696, N7665, N2147);
not NOT1 (N7697, N7692);
or OR2 (N7698, N7686, N3551);
xor XOR2 (N7699, N7694, N3738);
buf BUF1 (N7700, N7672);
buf BUF1 (N7701, N7700);
not NOT1 (N7702, N7699);
nor NOR2 (N7703, N7682, N1111);
buf BUF1 (N7704, N7698);
not NOT1 (N7705, N7673);
and AND3 (N7706, N7702, N2693, N5896);
buf BUF1 (N7707, N7706);
buf BUF1 (N7708, N7696);
nand NAND2 (N7709, N7707, N1274);
nor NOR2 (N7710, N7695, N3772);
nand NAND3 (N7711, N7687, N5138, N4920);
xor XOR2 (N7712, N7704, N2042);
xor XOR2 (N7713, N7701, N7261);
xor XOR2 (N7714, N7703, N5805);
nand NAND3 (N7715, N7713, N2880, N174);
nand NAND3 (N7716, N7714, N4193, N3724);
and AND3 (N7717, N7697, N3447, N5177);
nor NOR4 (N7718, N7709, N6996, N4232, N5167);
or OR2 (N7719, N7711, N272);
not NOT1 (N7720, N7712);
and AND3 (N7721, N7708, N2495, N4717);
nor NOR3 (N7722, N7705, N6928, N4441);
xor XOR2 (N7723, N7683, N1886);
and AND3 (N7724, N7710, N6065, N3440);
and AND3 (N7725, N7723, N6401, N519);
xor XOR2 (N7726, N7725, N312);
and AND4 (N7727, N7719, N5992, N4518, N5854);
nor NOR4 (N7728, N7720, N883, N2110, N4769);
and AND2 (N7729, N7722, N3975);
buf BUF1 (N7730, N7718);
xor XOR2 (N7731, N7717, N5984);
nor NOR3 (N7732, N7728, N1222, N2959);
buf BUF1 (N7733, N7729);
nor NOR3 (N7734, N7730, N4322, N1217);
nand NAND4 (N7735, N7716, N2754, N1803, N6137);
not NOT1 (N7736, N7727);
xor XOR2 (N7737, N7734, N3721);
nand NAND4 (N7738, N7721, N1794, N6507, N3989);
nand NAND4 (N7739, N7731, N5775, N7590, N593);
xor XOR2 (N7740, N7738, N7736);
nor NOR2 (N7741, N6115, N3117);
buf BUF1 (N7742, N7726);
nand NAND4 (N7743, N7737, N7535, N1944, N353);
xor XOR2 (N7744, N7743, N2667);
nor NOR3 (N7745, N7733, N390, N789);
not NOT1 (N7746, N7742);
and AND3 (N7747, N7744, N7524, N432);
xor XOR2 (N7748, N7747, N980);
buf BUF1 (N7749, N7732);
buf BUF1 (N7750, N7745);
nand NAND2 (N7751, N7741, N2607);
or OR2 (N7752, N7724, N4379);
and AND2 (N7753, N7748, N1835);
not NOT1 (N7754, N7751);
buf BUF1 (N7755, N7715);
not NOT1 (N7756, N7752);
buf BUF1 (N7757, N7739);
or OR4 (N7758, N7735, N6964, N5267, N4475);
buf BUF1 (N7759, N7757);
xor XOR2 (N7760, N7754, N4236);
or OR3 (N7761, N7740, N7177, N3794);
and AND2 (N7762, N7750, N4341);
buf BUF1 (N7763, N7753);
buf BUF1 (N7764, N7763);
not NOT1 (N7765, N7749);
buf BUF1 (N7766, N7759);
nand NAND4 (N7767, N7758, N3266, N5705, N3185);
not NOT1 (N7768, N7766);
nand NAND3 (N7769, N7764, N3472, N1098);
xor XOR2 (N7770, N7746, N1631);
nor NOR3 (N7771, N7769, N6865, N3626);
not NOT1 (N7772, N7761);
not NOT1 (N7773, N7756);
nor NOR3 (N7774, N7771, N2330, N1223);
and AND3 (N7775, N7774, N4718, N5643);
not NOT1 (N7776, N7770);
nand NAND4 (N7777, N7768, N2850, N4827, N4796);
or OR4 (N7778, N7777, N4460, N2637, N472);
nand NAND4 (N7779, N7762, N7731, N354, N4731);
not NOT1 (N7780, N7776);
buf BUF1 (N7781, N7773);
nor NOR2 (N7782, N7775, N2553);
and AND4 (N7783, N7780, N1511, N6597, N5741);
nand NAND2 (N7784, N7772, N2691);
or OR3 (N7785, N7778, N1757, N2071);
not NOT1 (N7786, N7784);
and AND3 (N7787, N7755, N7667, N212);
and AND3 (N7788, N7765, N3777, N2341);
xor XOR2 (N7789, N7788, N5234);
nor NOR2 (N7790, N7789, N456);
not NOT1 (N7791, N7767);
nand NAND2 (N7792, N7790, N4232);
nand NAND2 (N7793, N7783, N5532);
and AND3 (N7794, N7791, N621, N4118);
or OR2 (N7795, N7792, N5919);
and AND3 (N7796, N7785, N1701, N3324);
nor NOR4 (N7797, N7760, N7217, N12, N5042);
xor XOR2 (N7798, N7794, N258);
buf BUF1 (N7799, N7795);
nor NOR3 (N7800, N7779, N1531, N5670);
not NOT1 (N7801, N7797);
not NOT1 (N7802, N7796);
not NOT1 (N7803, N7798);
nor NOR3 (N7804, N7781, N3259, N6209);
and AND3 (N7805, N7782, N5535, N5859);
nand NAND3 (N7806, N7793, N5139, N2941);
buf BUF1 (N7807, N7799);
xor XOR2 (N7808, N7787, N3173);
nand NAND3 (N7809, N7801, N5735, N1837);
buf BUF1 (N7810, N7804);
and AND2 (N7811, N7808, N3012);
buf BUF1 (N7812, N7811);
xor XOR2 (N7813, N7807, N259);
nand NAND4 (N7814, N7802, N6935, N1218, N5839);
nand NAND2 (N7815, N7803, N5673);
xor XOR2 (N7816, N7809, N2651);
and AND3 (N7817, N7800, N5661, N2845);
and AND4 (N7818, N7786, N1813, N274, N255);
or OR2 (N7819, N7805, N89);
xor XOR2 (N7820, N7810, N1063);
not NOT1 (N7821, N7818);
or OR2 (N7822, N7815, N3936);
or OR4 (N7823, N7814, N1260, N7720, N5484);
not NOT1 (N7824, N7813);
not NOT1 (N7825, N7824);
or OR2 (N7826, N7817, N5161);
not NOT1 (N7827, N7819);
buf BUF1 (N7828, N7816);
xor XOR2 (N7829, N7826, N3927);
or OR4 (N7830, N7806, N6930, N4440, N595);
xor XOR2 (N7831, N7825, N2553);
not NOT1 (N7832, N7828);
buf BUF1 (N7833, N7820);
or OR4 (N7834, N7833, N2845, N3857, N6111);
buf BUF1 (N7835, N7829);
xor XOR2 (N7836, N7827, N4822);
and AND3 (N7837, N7836, N4009, N7244);
or OR3 (N7838, N7832, N7265, N4814);
buf BUF1 (N7839, N7821);
buf BUF1 (N7840, N7812);
not NOT1 (N7841, N7823);
xor XOR2 (N7842, N7831, N6069);
buf BUF1 (N7843, N7840);
buf BUF1 (N7844, N7838);
xor XOR2 (N7845, N7842, N5876);
and AND2 (N7846, N7845, N1717);
xor XOR2 (N7847, N7846, N5145);
or OR3 (N7848, N7830, N419, N5025);
xor XOR2 (N7849, N7847, N6177);
or OR2 (N7850, N7841, N3545);
and AND2 (N7851, N7843, N5690);
xor XOR2 (N7852, N7822, N1366);
nand NAND2 (N7853, N7848, N3971);
buf BUF1 (N7854, N7839);
nand NAND2 (N7855, N7844, N7734);
xor XOR2 (N7856, N7851, N3118);
nor NOR3 (N7857, N7835, N1871, N6923);
and AND2 (N7858, N7855, N1672);
and AND4 (N7859, N7849, N6148, N194, N3487);
nor NOR3 (N7860, N7852, N6844, N6639);
or OR3 (N7861, N7859, N4655, N7653);
and AND3 (N7862, N7837, N3570, N3230);
or OR3 (N7863, N7861, N2332, N2189);
buf BUF1 (N7864, N7856);
nand NAND2 (N7865, N7834, N358);
buf BUF1 (N7866, N7857);
xor XOR2 (N7867, N7865, N7315);
not NOT1 (N7868, N7853);
xor XOR2 (N7869, N7867, N2086);
buf BUF1 (N7870, N7860);
and AND2 (N7871, N7869, N3731);
nor NOR3 (N7872, N7858, N3665, N7812);
buf BUF1 (N7873, N7864);
or OR3 (N7874, N7854, N4813, N5960);
xor XOR2 (N7875, N7870, N63);
not NOT1 (N7876, N7872);
not NOT1 (N7877, N7876);
nor NOR4 (N7878, N7866, N1110, N2067, N1355);
not NOT1 (N7879, N7875);
nand NAND2 (N7880, N7862, N2578);
and AND2 (N7881, N7871, N6307);
not NOT1 (N7882, N7850);
nor NOR3 (N7883, N7868, N2401, N6138);
not NOT1 (N7884, N7879);
xor XOR2 (N7885, N7873, N1123);
xor XOR2 (N7886, N7881, N2094);
buf BUF1 (N7887, N7885);
xor XOR2 (N7888, N7883, N2978);
or OR2 (N7889, N7887, N719);
buf BUF1 (N7890, N7878);
nand NAND4 (N7891, N7889, N681, N2432, N6372);
nor NOR3 (N7892, N7877, N2477, N5586);
buf BUF1 (N7893, N7886);
and AND2 (N7894, N7888, N5129);
xor XOR2 (N7895, N7880, N3091);
not NOT1 (N7896, N7895);
buf BUF1 (N7897, N7896);
buf BUF1 (N7898, N7897);
nor NOR2 (N7899, N7884, N6714);
and AND3 (N7900, N7892, N470, N335);
and AND4 (N7901, N7899, N3503, N2641, N4112);
nand NAND3 (N7902, N7893, N4376, N6951);
nor NOR3 (N7903, N7891, N3325, N1567);
buf BUF1 (N7904, N7882);
nor NOR4 (N7905, N7898, N1455, N3069, N5327);
nor NOR2 (N7906, N7904, N7100);
xor XOR2 (N7907, N7890, N4584);
xor XOR2 (N7908, N7903, N2821);
or OR2 (N7909, N7908, N195);
xor XOR2 (N7910, N7909, N841);
or OR4 (N7911, N7906, N5062, N3417, N6899);
buf BUF1 (N7912, N7902);
nor NOR3 (N7913, N7907, N281, N6106);
nand NAND4 (N7914, N7910, N919, N3049, N5325);
nor NOR3 (N7915, N7905, N6520, N3441);
nand NAND4 (N7916, N7915, N4392, N5265, N1150);
nand NAND2 (N7917, N7874, N144);
xor XOR2 (N7918, N7917, N6455);
or OR3 (N7919, N7912, N958, N6914);
or OR4 (N7920, N7911, N4235, N6539, N3554);
and AND4 (N7921, N7918, N1510, N488, N1729);
nor NOR4 (N7922, N7901, N89, N5837, N5400);
and AND4 (N7923, N7894, N2188, N5936, N6487);
buf BUF1 (N7924, N7921);
nor NOR3 (N7925, N7923, N308, N2909);
and AND3 (N7926, N7900, N6055, N6497);
or OR3 (N7927, N7924, N3154, N7332);
xor XOR2 (N7928, N7913, N7804);
xor XOR2 (N7929, N7922, N4983);
xor XOR2 (N7930, N7925, N415);
not NOT1 (N7931, N7929);
nand NAND4 (N7932, N7931, N77, N503, N2972);
nor NOR3 (N7933, N7927, N988, N4623);
nand NAND3 (N7934, N7928, N1518, N6819);
buf BUF1 (N7935, N7930);
not NOT1 (N7936, N7935);
nor NOR4 (N7937, N7933, N4703, N307, N6598);
or OR4 (N7938, N7926, N2460, N3663, N3979);
not NOT1 (N7939, N7932);
nand NAND3 (N7940, N7934, N3478, N254);
or OR2 (N7941, N7939, N3419);
not NOT1 (N7942, N7940);
and AND4 (N7943, N7920, N94, N7809, N7894);
buf BUF1 (N7944, N7943);
and AND4 (N7945, N7944, N5647, N933, N3289);
not NOT1 (N7946, N7914);
not NOT1 (N7947, N7946);
and AND4 (N7948, N7936, N1804, N4768, N2517);
xor XOR2 (N7949, N7937, N6347);
nor NOR3 (N7950, N7919, N1711, N3935);
buf BUF1 (N7951, N7950);
buf BUF1 (N7952, N7863);
nand NAND2 (N7953, N7916, N476);
nor NOR4 (N7954, N7942, N2307, N3350, N6755);
nand NAND3 (N7955, N7953, N441, N7656);
nand NAND3 (N7956, N7949, N365, N1120);
or OR3 (N7957, N7941, N418, N7659);
or OR3 (N7958, N7957, N5150, N4871);
or OR2 (N7959, N7948, N233);
xor XOR2 (N7960, N7947, N6689);
or OR3 (N7961, N7955, N7365, N2728);
xor XOR2 (N7962, N7959, N4501);
nand NAND2 (N7963, N7938, N3598);
buf BUF1 (N7964, N7963);
nor NOR2 (N7965, N7964, N6493);
buf BUF1 (N7966, N7961);
not NOT1 (N7967, N7951);
and AND3 (N7968, N7962, N5714, N4147);
and AND4 (N7969, N7952, N4657, N3973, N3706);
not NOT1 (N7970, N7960);
and AND4 (N7971, N7945, N1639, N2634, N4491);
nor NOR3 (N7972, N7966, N1822, N2593);
nand NAND3 (N7973, N7956, N2019, N2950);
buf BUF1 (N7974, N7970);
not NOT1 (N7975, N7954);
nor NOR3 (N7976, N7974, N3379, N5575);
or OR2 (N7977, N7972, N2746);
and AND3 (N7978, N7968, N1876, N1405);
not NOT1 (N7979, N7965);
xor XOR2 (N7980, N7967, N1748);
or OR3 (N7981, N7978, N101, N4854);
buf BUF1 (N7982, N7971);
nor NOR4 (N7983, N7981, N3083, N6349, N5753);
or OR2 (N7984, N7975, N4069);
or OR3 (N7985, N7969, N2913, N6496);
nand NAND3 (N7986, N7979, N628, N5859);
and AND3 (N7987, N7983, N6496, N7609);
buf BUF1 (N7988, N7987);
buf BUF1 (N7989, N7982);
or OR4 (N7990, N7976, N4183, N2182, N6147);
or OR3 (N7991, N7990, N504, N6613);
nand NAND4 (N7992, N7985, N5095, N7486, N5490);
or OR3 (N7993, N7977, N3248, N1991);
nand NAND2 (N7994, N7973, N3971);
not NOT1 (N7995, N7988);
not NOT1 (N7996, N7995);
nand NAND2 (N7997, N7980, N6741);
xor XOR2 (N7998, N7996, N2502);
or OR2 (N7999, N7997, N4202);
and AND2 (N8000, N7999, N3169);
not NOT1 (N8001, N7993);
xor XOR2 (N8002, N7958, N262);
not NOT1 (N8003, N7986);
and AND3 (N8004, N8000, N5961, N5948);
xor XOR2 (N8005, N8002, N3732);
nor NOR2 (N8006, N8004, N5528);
xor XOR2 (N8007, N8001, N1201);
buf BUF1 (N8008, N7989);
nor NOR4 (N8009, N7994, N3286, N7354, N4276);
nor NOR2 (N8010, N7984, N187);
not NOT1 (N8011, N8008);
and AND2 (N8012, N7998, N4992);
nor NOR2 (N8013, N8012, N3500);
and AND3 (N8014, N8011, N2612, N2900);
xor XOR2 (N8015, N8003, N938);
buf BUF1 (N8016, N8014);
nor NOR3 (N8017, N8006, N7025, N6336);
buf BUF1 (N8018, N8016);
not NOT1 (N8019, N7992);
nand NAND4 (N8020, N8013, N6263, N7087, N3890);
xor XOR2 (N8021, N8017, N6448);
buf BUF1 (N8022, N8015);
nor NOR2 (N8023, N8021, N4621);
buf BUF1 (N8024, N8005);
nand NAND3 (N8025, N8024, N167, N811);
nand NAND3 (N8026, N8019, N6383, N1805);
not NOT1 (N8027, N8020);
nor NOR2 (N8028, N8007, N7970);
nor NOR4 (N8029, N8018, N4625, N5577, N7448);
not NOT1 (N8030, N8022);
xor XOR2 (N8031, N8009, N878);
xor XOR2 (N8032, N8025, N2045);
and AND2 (N8033, N8031, N5390);
nand NAND2 (N8034, N8010, N1730);
or OR3 (N8035, N8026, N5231, N7099);
or OR3 (N8036, N8034, N1385, N2516);
and AND4 (N8037, N8029, N2087, N2754, N1216);
nor NOR3 (N8038, N8030, N497, N3671);
buf BUF1 (N8039, N8023);
nand NAND3 (N8040, N8036, N2994, N6985);
xor XOR2 (N8041, N8040, N1501);
not NOT1 (N8042, N7991);
nor NOR4 (N8043, N8041, N992, N6583, N7948);
and AND2 (N8044, N8042, N4669);
buf BUF1 (N8045, N8037);
buf BUF1 (N8046, N8039);
buf BUF1 (N8047, N8043);
xor XOR2 (N8048, N8038, N5777);
xor XOR2 (N8049, N8046, N119);
xor XOR2 (N8050, N8035, N6926);
buf BUF1 (N8051, N8033);
nor NOR3 (N8052, N8049, N6648, N6892);
nor NOR2 (N8053, N8027, N3461);
nand NAND2 (N8054, N8050, N2777);
or OR4 (N8055, N8044, N298, N6429, N6281);
buf BUF1 (N8056, N8045);
buf BUF1 (N8057, N8032);
buf BUF1 (N8058, N8055);
xor XOR2 (N8059, N8053, N3657);
and AND3 (N8060, N8051, N6226, N5036);
xor XOR2 (N8061, N8047, N6047);
nand NAND3 (N8062, N8052, N735, N375);
xor XOR2 (N8063, N8056, N5213);
xor XOR2 (N8064, N8060, N5325);
or OR3 (N8065, N8048, N334, N3669);
nor NOR4 (N8066, N8058, N4523, N692, N2041);
nand NAND3 (N8067, N8063, N5880, N1960);
and AND4 (N8068, N8062, N3451, N1203, N5822);
nor NOR2 (N8069, N8067, N1556);
xor XOR2 (N8070, N8069, N4447);
not NOT1 (N8071, N8059);
xor XOR2 (N8072, N8054, N6838);
and AND3 (N8073, N8070, N88, N933);
nand NAND3 (N8074, N8071, N3550, N2042);
or OR2 (N8075, N8064, N3290);
buf BUF1 (N8076, N8028);
and AND3 (N8077, N8061, N2730, N5224);
or OR2 (N8078, N8068, N2629);
buf BUF1 (N8079, N8066);
buf BUF1 (N8080, N8078);
or OR2 (N8081, N8065, N4397);
not NOT1 (N8082, N8075);
or OR3 (N8083, N8074, N1598, N1290);
nand NAND2 (N8084, N8080, N4643);
xor XOR2 (N8085, N8083, N3167);
or OR2 (N8086, N8081, N2885);
or OR4 (N8087, N8084, N1467, N6855, N4943);
or OR2 (N8088, N8057, N3997);
xor XOR2 (N8089, N8085, N7980);
nand NAND2 (N8090, N8087, N4227);
and AND3 (N8091, N8079, N2477, N5325);
nand NAND3 (N8092, N8086, N3254, N4038);
not NOT1 (N8093, N8088);
or OR2 (N8094, N8077, N6092);
not NOT1 (N8095, N8090);
nor NOR3 (N8096, N8091, N751, N6458);
nor NOR3 (N8097, N8096, N6724, N2218);
nor NOR2 (N8098, N8089, N6123);
nor NOR2 (N8099, N8073, N1501);
not NOT1 (N8100, N8092);
not NOT1 (N8101, N8097);
xor XOR2 (N8102, N8082, N5575);
xor XOR2 (N8103, N8094, N4100);
nand NAND4 (N8104, N8099, N443, N5540, N6609);
nand NAND3 (N8105, N8103, N3028, N1280);
nor NOR3 (N8106, N8095, N671, N44);
not NOT1 (N8107, N8072);
xor XOR2 (N8108, N8101, N5815);
xor XOR2 (N8109, N8098, N2080);
nor NOR4 (N8110, N8104, N4855, N4289, N6115);
not NOT1 (N8111, N8107);
nand NAND4 (N8112, N8076, N5026, N7603, N3388);
nor NOR4 (N8113, N8112, N6815, N3920, N1345);
buf BUF1 (N8114, N8093);
nor NOR4 (N8115, N8108, N1347, N2363, N4819);
buf BUF1 (N8116, N8113);
not NOT1 (N8117, N8102);
not NOT1 (N8118, N8105);
or OR3 (N8119, N8115, N1595, N3527);
xor XOR2 (N8120, N8106, N3989);
or OR4 (N8121, N8110, N5365, N8032, N5331);
not NOT1 (N8122, N8121);
buf BUF1 (N8123, N8109);
or OR4 (N8124, N8118, N4844, N750, N1356);
nor NOR4 (N8125, N8111, N3476, N6237, N738);
not NOT1 (N8126, N8116);
or OR3 (N8127, N8120, N4684, N911);
not NOT1 (N8128, N8122);
nor NOR2 (N8129, N8100, N3377);
nand NAND4 (N8130, N8123, N6384, N5963, N6023);
buf BUF1 (N8131, N8130);
xor XOR2 (N8132, N8131, N1687);
nand NAND4 (N8133, N8128, N7370, N2662, N1212);
nor NOR4 (N8134, N8117, N7748, N2905, N1194);
nor NOR4 (N8135, N8129, N4990, N680, N5123);
buf BUF1 (N8136, N8135);
buf BUF1 (N8137, N8133);
nand NAND2 (N8138, N8114, N8065);
not NOT1 (N8139, N8127);
xor XOR2 (N8140, N8132, N1860);
buf BUF1 (N8141, N8125);
nor NOR2 (N8142, N8136, N3132);
xor XOR2 (N8143, N8124, N7794);
xor XOR2 (N8144, N8141, N4708);
xor XOR2 (N8145, N8143, N4644);
not NOT1 (N8146, N8119);
nand NAND4 (N8147, N8145, N5761, N5557, N3840);
not NOT1 (N8148, N8138);
and AND4 (N8149, N8148, N848, N4707, N2243);
or OR4 (N8150, N8146, N6581, N4591, N4656);
nor NOR2 (N8151, N8147, N194);
nand NAND2 (N8152, N8144, N6593);
not NOT1 (N8153, N8152);
not NOT1 (N8154, N8137);
not NOT1 (N8155, N8149);
nand NAND4 (N8156, N8153, N3966, N424, N2329);
nand NAND2 (N8157, N8156, N6951);
not NOT1 (N8158, N8150);
nor NOR4 (N8159, N8158, N1850, N3836, N388);
xor XOR2 (N8160, N8140, N3328);
xor XOR2 (N8161, N8139, N608);
nand NAND4 (N8162, N8155, N2928, N3978, N6739);
not NOT1 (N8163, N8151);
nand NAND3 (N8164, N8163, N3979, N1968);
nand NAND3 (N8165, N8161, N590, N6541);
buf BUF1 (N8166, N8159);
and AND4 (N8167, N8162, N6664, N6946, N2779);
not NOT1 (N8168, N8154);
nor NOR4 (N8169, N8165, N5596, N5008, N6907);
nand NAND2 (N8170, N8134, N7000);
and AND3 (N8171, N8126, N689, N6148);
not NOT1 (N8172, N8160);
buf BUF1 (N8173, N8168);
nor NOR3 (N8174, N8170, N191, N7620);
and AND3 (N8175, N8157, N5705, N2945);
nand NAND2 (N8176, N8172, N3270);
not NOT1 (N8177, N8174);
xor XOR2 (N8178, N8169, N6105);
nor NOR4 (N8179, N8166, N2535, N5382, N2963);
xor XOR2 (N8180, N8142, N5710);
xor XOR2 (N8181, N8171, N1514);
not NOT1 (N8182, N8181);
or OR4 (N8183, N8176, N1520, N6100, N263);
nor NOR4 (N8184, N8178, N1387, N2128, N8145);
buf BUF1 (N8185, N8179);
buf BUF1 (N8186, N8175);
buf BUF1 (N8187, N8173);
or OR3 (N8188, N8183, N2096, N2134);
buf BUF1 (N8189, N8185);
nor NOR3 (N8190, N8184, N2615, N2658);
not NOT1 (N8191, N8180);
buf BUF1 (N8192, N8189);
and AND2 (N8193, N8191, N4406);
or OR3 (N8194, N8193, N5666, N7601);
or OR4 (N8195, N8190, N1383, N3163, N2027);
nor NOR3 (N8196, N8188, N7310, N3914);
and AND3 (N8197, N8194, N1719, N1616);
nor NOR3 (N8198, N8195, N2588, N2238);
not NOT1 (N8199, N8198);
not NOT1 (N8200, N8177);
nor NOR4 (N8201, N8187, N3487, N3299, N2248);
xor XOR2 (N8202, N8197, N5891);
nand NAND4 (N8203, N8196, N31, N5556, N2176);
nand NAND2 (N8204, N8202, N5769);
nor NOR3 (N8205, N8199, N5452, N6252);
or OR3 (N8206, N8205, N5003, N4625);
or OR4 (N8207, N8182, N6134, N6869, N856);
nor NOR2 (N8208, N8206, N5640);
or OR3 (N8209, N8203, N4623, N6841);
nand NAND4 (N8210, N8208, N5521, N7329, N7265);
buf BUF1 (N8211, N8204);
nand NAND4 (N8212, N8200, N4898, N7673, N6594);
not NOT1 (N8213, N8201);
nor NOR2 (N8214, N8212, N800);
not NOT1 (N8215, N8209);
or OR3 (N8216, N8210, N6663, N1200);
xor XOR2 (N8217, N8216, N6765);
or OR2 (N8218, N8164, N7560);
nor NOR2 (N8219, N8218, N4485);
nor NOR2 (N8220, N8211, N6342);
nor NOR2 (N8221, N8213, N4895);
nand NAND4 (N8222, N8215, N7520, N5640, N350);
and AND4 (N8223, N8221, N7118, N5451, N5087);
not NOT1 (N8224, N8167);
buf BUF1 (N8225, N8217);
or OR4 (N8226, N8214, N7238, N6275, N7655);
and AND2 (N8227, N8225, N4228);
and AND2 (N8228, N8220, N7361);
nor NOR2 (N8229, N8228, N1599);
not NOT1 (N8230, N8186);
xor XOR2 (N8231, N8229, N447);
buf BUF1 (N8232, N8223);
not NOT1 (N8233, N8226);
nor NOR2 (N8234, N8207, N3712);
and AND2 (N8235, N8231, N6250);
buf BUF1 (N8236, N8222);
and AND3 (N8237, N8219, N8083, N3095);
xor XOR2 (N8238, N8237, N3000);
buf BUF1 (N8239, N8224);
nand NAND3 (N8240, N8233, N3123, N5271);
not NOT1 (N8241, N8192);
or OR3 (N8242, N8236, N3974, N3138);
not NOT1 (N8243, N8234);
or OR2 (N8244, N8240, N8203);
nand NAND2 (N8245, N8227, N4078);
or OR2 (N8246, N8235, N7885);
nand NAND2 (N8247, N8244, N3007);
buf BUF1 (N8248, N8238);
nor NOR3 (N8249, N8247, N6246, N8069);
or OR4 (N8250, N8232, N4598, N163, N408);
nand NAND3 (N8251, N8249, N2388, N1419);
xor XOR2 (N8252, N8245, N2857);
or OR2 (N8253, N8250, N6491);
nand NAND3 (N8254, N8252, N2930, N6540);
nand NAND4 (N8255, N8243, N7070, N6785, N8163);
or OR2 (N8256, N8230, N5628);
and AND2 (N8257, N8248, N5895);
and AND2 (N8258, N8253, N7498);
buf BUF1 (N8259, N8258);
nand NAND2 (N8260, N8242, N3383);
or OR4 (N8261, N8256, N1846, N6873, N149);
nand NAND4 (N8262, N8257, N6709, N2931, N3702);
and AND2 (N8263, N8251, N7761);
and AND4 (N8264, N8261, N2321, N6828, N3119);
or OR4 (N8265, N8255, N5623, N5923, N5923);
nand NAND2 (N8266, N8259, N8060);
not NOT1 (N8267, N8241);
buf BUF1 (N8268, N8254);
and AND2 (N8269, N8246, N5106);
xor XOR2 (N8270, N8268, N4386);
buf BUF1 (N8271, N8267);
xor XOR2 (N8272, N8239, N5472);
or OR4 (N8273, N8269, N3808, N5957, N4186);
not NOT1 (N8274, N8271);
buf BUF1 (N8275, N8274);
or OR4 (N8276, N8262, N1307, N955, N5559);
and AND2 (N8277, N8270, N3163);
or OR3 (N8278, N8272, N7771, N1017);
buf BUF1 (N8279, N8260);
nor NOR4 (N8280, N8275, N7667, N8008, N6958);
nand NAND3 (N8281, N8273, N3662, N7958);
and AND2 (N8282, N8281, N5725);
buf BUF1 (N8283, N8264);
not NOT1 (N8284, N8276);
and AND3 (N8285, N8263, N2547, N5356);
nand NAND3 (N8286, N8265, N4202, N2244);
nor NOR2 (N8287, N8266, N7508);
nor NOR3 (N8288, N8286, N3542, N6000);
nand NAND4 (N8289, N8285, N1886, N6532, N166);
nand NAND2 (N8290, N8288, N4240);
xor XOR2 (N8291, N8290, N75);
and AND3 (N8292, N8277, N7222, N2764);
buf BUF1 (N8293, N8292);
or OR2 (N8294, N8291, N3287);
xor XOR2 (N8295, N8294, N4185);
or OR4 (N8296, N8279, N5473, N4919, N6921);
buf BUF1 (N8297, N8280);
buf BUF1 (N8298, N8295);
nor NOR4 (N8299, N8283, N4926, N1439, N7953);
nor NOR3 (N8300, N8298, N8004, N1728);
buf BUF1 (N8301, N8299);
and AND2 (N8302, N8282, N2042);
and AND2 (N8303, N8302, N5500);
xor XOR2 (N8304, N8284, N7270);
and AND3 (N8305, N8278, N5898, N1442);
nor NOR4 (N8306, N8297, N7318, N5678, N7450);
nor NOR2 (N8307, N8306, N7464);
xor XOR2 (N8308, N8301, N2792);
buf BUF1 (N8309, N8296);
and AND4 (N8310, N8289, N4000, N7357, N2635);
not NOT1 (N8311, N8287);
nor NOR4 (N8312, N8307, N4250, N7979, N5409);
or OR2 (N8313, N8310, N7544);
and AND2 (N8314, N8313, N8085);
buf BUF1 (N8315, N8305);
nor NOR4 (N8316, N8312, N3246, N1520, N7952);
not NOT1 (N8317, N8303);
and AND2 (N8318, N8309, N33);
xor XOR2 (N8319, N8316, N803);
xor XOR2 (N8320, N8319, N4222);
nor NOR2 (N8321, N8293, N2561);
not NOT1 (N8322, N8311);
and AND3 (N8323, N8320, N266, N3085);
and AND2 (N8324, N8322, N1532);
buf BUF1 (N8325, N8314);
and AND2 (N8326, N8323, N3746);
buf BUF1 (N8327, N8304);
and AND2 (N8328, N8308, N1310);
buf BUF1 (N8329, N8317);
nand NAND2 (N8330, N8326, N5200);
or OR3 (N8331, N8318, N2998, N1054);
not NOT1 (N8332, N8321);
or OR2 (N8333, N8330, N2042);
not NOT1 (N8334, N8328);
not NOT1 (N8335, N8331);
not NOT1 (N8336, N8332);
or OR2 (N8337, N8300, N173);
not NOT1 (N8338, N8327);
and AND2 (N8339, N8337, N2650);
nor NOR3 (N8340, N8336, N1254, N5725);
not NOT1 (N8341, N8325);
nand NAND2 (N8342, N8335, N5855);
or OR4 (N8343, N8339, N6682, N1119, N7347);
and AND3 (N8344, N8315, N7513, N1535);
or OR2 (N8345, N8329, N1432);
not NOT1 (N8346, N8341);
nor NOR3 (N8347, N8345, N2433, N5151);
xor XOR2 (N8348, N8344, N4713);
nor NOR3 (N8349, N8347, N3138, N2103);
nand NAND3 (N8350, N8333, N6975, N6421);
not NOT1 (N8351, N8346);
and AND2 (N8352, N8324, N4604);
buf BUF1 (N8353, N8350);
or OR2 (N8354, N8349, N3615);
xor XOR2 (N8355, N8338, N6871);
xor XOR2 (N8356, N8343, N5239);
nand NAND2 (N8357, N8356, N2188);
nand NAND2 (N8358, N8353, N4042);
not NOT1 (N8359, N8358);
and AND3 (N8360, N8357, N6754, N4066);
nand NAND3 (N8361, N8351, N2950, N2610);
and AND2 (N8362, N8354, N6391);
or OR3 (N8363, N8342, N2433, N402);
buf BUF1 (N8364, N8362);
and AND4 (N8365, N8340, N5028, N7610, N115);
or OR3 (N8366, N8352, N5674, N2404);
and AND4 (N8367, N8364, N3693, N1256, N1317);
or OR4 (N8368, N8359, N4665, N7550, N4406);
or OR4 (N8369, N8360, N4269, N8208, N686);
or OR2 (N8370, N8365, N4743);
buf BUF1 (N8371, N8369);
nor NOR4 (N8372, N8355, N405, N5890, N774);
or OR3 (N8373, N8348, N3017, N2097);
and AND2 (N8374, N8334, N3740);
not NOT1 (N8375, N8367);
and AND3 (N8376, N8370, N6403, N4653);
and AND2 (N8377, N8375, N7201);
not NOT1 (N8378, N8363);
xor XOR2 (N8379, N8376, N2843);
xor XOR2 (N8380, N8378, N4552);
and AND4 (N8381, N8379, N800, N1227, N6117);
or OR4 (N8382, N8377, N3268, N5582, N1999);
or OR2 (N8383, N8372, N6572);
nand NAND2 (N8384, N8374, N3638);
xor XOR2 (N8385, N8371, N4840);
or OR3 (N8386, N8381, N4553, N1092);
or OR2 (N8387, N8385, N336);
not NOT1 (N8388, N8380);
nor NOR2 (N8389, N8368, N7514);
and AND4 (N8390, N8384, N1275, N2718, N7244);
not NOT1 (N8391, N8383);
and AND3 (N8392, N8388, N634, N5973);
and AND3 (N8393, N8361, N4215, N2637);
or OR2 (N8394, N8373, N792);
nand NAND2 (N8395, N8366, N5696);
or OR2 (N8396, N8386, N6192);
xor XOR2 (N8397, N8389, N1956);
or OR2 (N8398, N8396, N4818);
nor NOR4 (N8399, N8393, N4537, N1241, N3120);
buf BUF1 (N8400, N8398);
and AND2 (N8401, N8392, N5313);
and AND3 (N8402, N8397, N7344, N7136);
nand NAND4 (N8403, N8387, N3608, N921, N370);
and AND2 (N8404, N8401, N7889);
buf BUF1 (N8405, N8400);
nand NAND2 (N8406, N8405, N2204);
xor XOR2 (N8407, N8403, N2065);
or OR3 (N8408, N8399, N7733, N721);
xor XOR2 (N8409, N8402, N6384);
or OR3 (N8410, N8409, N6994, N4246);
buf BUF1 (N8411, N8407);
nor NOR3 (N8412, N8410, N6648, N719);
xor XOR2 (N8413, N8391, N6353);
xor XOR2 (N8414, N8412, N8072);
or OR3 (N8415, N8382, N4321, N2331);
not NOT1 (N8416, N8406);
or OR2 (N8417, N8411, N3568);
or OR3 (N8418, N8395, N1036, N4205);
buf BUF1 (N8419, N8394);
not NOT1 (N8420, N8413);
nand NAND3 (N8421, N8414, N587, N1236);
xor XOR2 (N8422, N8420, N887);
not NOT1 (N8423, N8415);
buf BUF1 (N8424, N8390);
xor XOR2 (N8425, N8408, N7281);
xor XOR2 (N8426, N8419, N4477);
xor XOR2 (N8427, N8422, N7316);
nand NAND3 (N8428, N8423, N2487, N7147);
and AND4 (N8429, N8417, N5398, N4527, N1655);
buf BUF1 (N8430, N8424);
nand NAND4 (N8431, N8429, N8054, N2219, N6554);
not NOT1 (N8432, N8427);
or OR3 (N8433, N8430, N3558, N5874);
and AND3 (N8434, N8404, N6424, N5202);
and AND4 (N8435, N8425, N1543, N8154, N2308);
not NOT1 (N8436, N8431);
or OR2 (N8437, N8421, N2210);
xor XOR2 (N8438, N8428, N474);
xor XOR2 (N8439, N8433, N1682);
and AND3 (N8440, N8435, N4482, N523);
not NOT1 (N8441, N8432);
nor NOR4 (N8442, N8439, N2544, N1905, N5922);
xor XOR2 (N8443, N8418, N6455);
and AND3 (N8444, N8436, N4060, N3809);
nand NAND2 (N8445, N8444, N4642);
nor NOR2 (N8446, N8442, N4151);
not NOT1 (N8447, N8426);
nor NOR2 (N8448, N8443, N7705);
nor NOR2 (N8449, N8448, N6508);
xor XOR2 (N8450, N8446, N4736);
not NOT1 (N8451, N8447);
buf BUF1 (N8452, N8441);
nand NAND3 (N8453, N8437, N7811, N7404);
and AND2 (N8454, N8450, N1877);
nand NAND3 (N8455, N8449, N5500, N4164);
or OR2 (N8456, N8434, N5922);
or OR4 (N8457, N8456, N968, N6883, N416);
and AND3 (N8458, N8454, N6578, N2107);
nor NOR4 (N8459, N8453, N1321, N7554, N4294);
and AND2 (N8460, N8452, N108);
buf BUF1 (N8461, N8445);
nand NAND4 (N8462, N8438, N637, N1621, N319);
nor NOR2 (N8463, N8451, N5782);
buf BUF1 (N8464, N8457);
buf BUF1 (N8465, N8459);
or OR2 (N8466, N8462, N6921);
or OR2 (N8467, N8463, N7637);
buf BUF1 (N8468, N8467);
nand NAND3 (N8469, N8458, N1812, N6369);
nand NAND4 (N8470, N8461, N6942, N7632, N1740);
or OR3 (N8471, N8470, N68, N7537);
nor NOR4 (N8472, N8465, N7583, N6537, N5702);
and AND2 (N8473, N8471, N1224);
nor NOR4 (N8474, N8460, N4803, N1447, N2657);
or OR3 (N8475, N8466, N764, N3918);
or OR3 (N8476, N8469, N1364, N8197);
and AND2 (N8477, N8416, N7014);
nor NOR2 (N8478, N8440, N8432);
nand NAND2 (N8479, N8473, N3381);
buf BUF1 (N8480, N8475);
or OR3 (N8481, N8464, N5203, N735);
xor XOR2 (N8482, N8479, N5115);
nor NOR2 (N8483, N8482, N7850);
nor NOR2 (N8484, N8468, N3772);
or OR2 (N8485, N8483, N8462);
and AND3 (N8486, N8472, N5499, N7407);
nor NOR3 (N8487, N8486, N6176, N1234);
nor NOR4 (N8488, N8478, N8274, N3328, N7271);
nor NOR4 (N8489, N8476, N2641, N8078, N476);
xor XOR2 (N8490, N8455, N2094);
not NOT1 (N8491, N8480);
or OR2 (N8492, N8490, N6136);
not NOT1 (N8493, N8484);
buf BUF1 (N8494, N8488);
nand NAND4 (N8495, N8493, N8051, N1807, N8155);
or OR2 (N8496, N8481, N2575);
nand NAND2 (N8497, N8477, N308);
not NOT1 (N8498, N8496);
or OR2 (N8499, N8494, N1798);
not NOT1 (N8500, N8489);
not NOT1 (N8501, N8491);
nor NOR2 (N8502, N8499, N1620);
buf BUF1 (N8503, N8492);
buf BUF1 (N8504, N8503);
xor XOR2 (N8505, N8474, N94);
nand NAND3 (N8506, N8505, N2669, N4021);
or OR2 (N8507, N8497, N5759);
nand NAND2 (N8508, N8500, N2765);
buf BUF1 (N8509, N8498);
nor NOR3 (N8510, N8501, N2902, N5294);
or OR2 (N8511, N8509, N7484);
and AND4 (N8512, N8511, N5531, N6000, N4795);
and AND2 (N8513, N8502, N4086);
buf BUF1 (N8514, N8506);
buf BUF1 (N8515, N8495);
xor XOR2 (N8516, N8487, N7008);
nor NOR4 (N8517, N8507, N3641, N645, N4175);
nor NOR4 (N8518, N8514, N2862, N1318, N5477);
nand NAND2 (N8519, N8516, N2956);
or OR2 (N8520, N8485, N5175);
and AND3 (N8521, N8508, N7426, N4128);
buf BUF1 (N8522, N8520);
and AND3 (N8523, N8515, N7474, N3687);
nor NOR2 (N8524, N8522, N5020);
not NOT1 (N8525, N8524);
nor NOR3 (N8526, N8525, N3292, N279);
or OR4 (N8527, N8517, N6098, N1645, N5980);
buf BUF1 (N8528, N8512);
and AND4 (N8529, N8527, N5564, N953, N7789);
nand NAND4 (N8530, N8519, N3026, N7801, N5866);
or OR2 (N8531, N8504, N4088);
nor NOR4 (N8532, N8523, N2227, N3617, N2732);
nand NAND3 (N8533, N8531, N219, N2982);
or OR3 (N8534, N8533, N2384, N3342);
xor XOR2 (N8535, N8526, N2110);
or OR4 (N8536, N8528, N1543, N8115, N8366);
nand NAND3 (N8537, N8534, N6454, N1760);
not NOT1 (N8538, N8535);
xor XOR2 (N8539, N8521, N8301);
not NOT1 (N8540, N8513);
or OR4 (N8541, N8510, N6027, N686, N8493);
not NOT1 (N8542, N8536);
nor NOR2 (N8543, N8539, N507);
nand NAND4 (N8544, N8529, N2631, N7387, N2073);
nand NAND3 (N8545, N8532, N5430, N4989);
buf BUF1 (N8546, N8530);
and AND2 (N8547, N8542, N2019);
buf BUF1 (N8548, N8543);
xor XOR2 (N8549, N8540, N7519);
nand NAND2 (N8550, N8518, N2620);
buf BUF1 (N8551, N8537);
nand NAND4 (N8552, N8544, N1647, N4930, N6716);
nand NAND3 (N8553, N8541, N220, N355);
and AND2 (N8554, N8547, N137);
nor NOR2 (N8555, N8549, N3342);
or OR4 (N8556, N8538, N1759, N7656, N5958);
nand NAND3 (N8557, N8554, N1824, N4336);
xor XOR2 (N8558, N8551, N1056);
not NOT1 (N8559, N8545);
buf BUF1 (N8560, N8552);
not NOT1 (N8561, N8560);
buf BUF1 (N8562, N8548);
nor NOR2 (N8563, N8562, N7561);
nor NOR3 (N8564, N8558, N7446, N6275);
or OR2 (N8565, N8550, N2303);
nand NAND2 (N8566, N8556, N6706);
not NOT1 (N8567, N8563);
nand NAND4 (N8568, N8555, N366, N8206, N31);
nor NOR3 (N8569, N8561, N428, N1805);
not NOT1 (N8570, N8546);
buf BUF1 (N8571, N8568);
xor XOR2 (N8572, N8559, N1965);
nand NAND4 (N8573, N8569, N7747, N8534, N333);
buf BUF1 (N8574, N8573);
nor NOR3 (N8575, N8570, N7552, N4789);
nand NAND2 (N8576, N8565, N3387);
or OR3 (N8577, N8575, N7900, N5733);
nor NOR4 (N8578, N8577, N7092, N7290, N6302);
xor XOR2 (N8579, N8567, N7767);
buf BUF1 (N8580, N8571);
nor NOR4 (N8581, N8576, N1094, N8262, N2924);
nand NAND3 (N8582, N8564, N227, N6849);
nor NOR4 (N8583, N8580, N577, N7032, N42);
and AND2 (N8584, N8553, N4190);
not NOT1 (N8585, N8579);
or OR4 (N8586, N8581, N4756, N7165, N3749);
and AND2 (N8587, N8566, N3001);
xor XOR2 (N8588, N8583, N1657);
buf BUF1 (N8589, N8578);
buf BUF1 (N8590, N8574);
buf BUF1 (N8591, N8572);
nor NOR3 (N8592, N8590, N7623, N144);
and AND4 (N8593, N8589, N5552, N5312, N5157);
or OR4 (N8594, N8593, N6132, N2883, N3878);
nand NAND3 (N8595, N8586, N4638, N4328);
and AND3 (N8596, N8585, N7355, N5859);
xor XOR2 (N8597, N8557, N5247);
nor NOR2 (N8598, N8594, N7350);
not NOT1 (N8599, N8591);
not NOT1 (N8600, N8599);
or OR2 (N8601, N8598, N396);
buf BUF1 (N8602, N8584);
nor NOR4 (N8603, N8582, N7170, N7924, N3724);
not NOT1 (N8604, N8596);
nand NAND2 (N8605, N8602, N6856);
nor NOR4 (N8606, N8597, N4601, N7054, N235);
nand NAND3 (N8607, N8606, N6190, N1084);
buf BUF1 (N8608, N8595);
buf BUF1 (N8609, N8592);
nand NAND2 (N8610, N8607, N7579);
nand NAND2 (N8611, N8601, N4409);
xor XOR2 (N8612, N8609, N3500);
or OR3 (N8613, N8600, N5427, N8594);
nor NOR2 (N8614, N8611, N2725);
not NOT1 (N8615, N8614);
or OR3 (N8616, N8610, N1969, N604);
buf BUF1 (N8617, N8608);
or OR2 (N8618, N8588, N5493);
not NOT1 (N8619, N8587);
buf BUF1 (N8620, N8619);
not NOT1 (N8621, N8616);
or OR4 (N8622, N8618, N1380, N2801, N4286);
or OR2 (N8623, N8621, N6598);
or OR2 (N8624, N8613, N1009);
or OR3 (N8625, N8620, N5186, N4267);
nor NOR2 (N8626, N8612, N213);
and AND2 (N8627, N8624, N1067);
buf BUF1 (N8628, N8626);
buf BUF1 (N8629, N8627);
nand NAND2 (N8630, N8617, N2634);
nor NOR3 (N8631, N8605, N8422, N5450);
nand NAND4 (N8632, N8630, N7019, N5352, N6835);
nand NAND4 (N8633, N8622, N4, N5755, N2825);
buf BUF1 (N8634, N8604);
not NOT1 (N8635, N8623);
not NOT1 (N8636, N8625);
and AND4 (N8637, N8631, N3886, N5451, N5954);
not NOT1 (N8638, N8629);
not NOT1 (N8639, N8633);
or OR2 (N8640, N8634, N3851);
nand NAND4 (N8641, N8638, N2813, N7307, N5646);
xor XOR2 (N8642, N8603, N2184);
nand NAND4 (N8643, N8637, N3280, N1953, N8580);
or OR4 (N8644, N8636, N3288, N7961, N509);
xor XOR2 (N8645, N8635, N5840);
nand NAND2 (N8646, N8628, N8381);
or OR3 (N8647, N8644, N6423, N5650);
buf BUF1 (N8648, N8646);
and AND4 (N8649, N8615, N237, N2386, N7600);
not NOT1 (N8650, N8643);
or OR4 (N8651, N8649, N435, N2347, N7440);
and AND2 (N8652, N8648, N5320);
xor XOR2 (N8653, N8650, N6454);
and AND2 (N8654, N8651, N4276);
or OR4 (N8655, N8653, N8165, N6900, N7986);
and AND2 (N8656, N8647, N229);
or OR3 (N8657, N8632, N3638, N3648);
nor NOR2 (N8658, N8656, N7289);
or OR3 (N8659, N8642, N6799, N8546);
nand NAND4 (N8660, N8658, N5234, N6464, N5795);
and AND2 (N8661, N8639, N8227);
nor NOR2 (N8662, N8659, N8392);
xor XOR2 (N8663, N8640, N4328);
buf BUF1 (N8664, N8660);
and AND3 (N8665, N8663, N5502, N1289);
and AND3 (N8666, N8641, N4171, N6486);
nor NOR4 (N8667, N8662, N6134, N1617, N5263);
and AND3 (N8668, N8666, N4941, N8155);
nand NAND3 (N8669, N8667, N2637, N3965);
nor NOR2 (N8670, N8664, N530);
and AND4 (N8671, N8665, N932, N3550, N2015);
nor NOR3 (N8672, N8645, N5703, N8262);
or OR3 (N8673, N8668, N7235, N6792);
buf BUF1 (N8674, N8671);
or OR2 (N8675, N8661, N4907);
xor XOR2 (N8676, N8654, N6504);
xor XOR2 (N8677, N8673, N3931);
and AND3 (N8678, N8670, N4156, N1032);
nand NAND2 (N8679, N8669, N48);
not NOT1 (N8680, N8675);
nand NAND2 (N8681, N8652, N2637);
buf BUF1 (N8682, N8657);
or OR3 (N8683, N8681, N2202, N2994);
and AND4 (N8684, N8677, N6180, N8276, N6131);
and AND3 (N8685, N8655, N751, N7042);
buf BUF1 (N8686, N8683);
and AND2 (N8687, N8682, N6133);
nand NAND4 (N8688, N8678, N5286, N1870, N6108);
or OR4 (N8689, N8685, N5055, N3331, N4182);
or OR2 (N8690, N8679, N2551);
not NOT1 (N8691, N8689);
and AND4 (N8692, N8676, N3112, N8430, N386);
nor NOR4 (N8693, N8692, N7828, N1857, N8545);
and AND2 (N8694, N8691, N3707);
not NOT1 (N8695, N8687);
not NOT1 (N8696, N8688);
and AND3 (N8697, N8690, N4139, N5134);
buf BUF1 (N8698, N8696);
and AND3 (N8699, N8698, N6128, N5445);
or OR3 (N8700, N8674, N7220, N6926);
not NOT1 (N8701, N8695);
or OR2 (N8702, N8693, N6521);
or OR3 (N8703, N8697, N3801, N4635);
buf BUF1 (N8704, N8703);
xor XOR2 (N8705, N8686, N8509);
xor XOR2 (N8706, N8699, N5130);
or OR2 (N8707, N8706, N3993);
nand NAND3 (N8708, N8701, N7684, N5142);
not NOT1 (N8709, N8702);
not NOT1 (N8710, N8672);
and AND4 (N8711, N8680, N7715, N3843, N5374);
nand NAND4 (N8712, N8705, N3512, N5651, N7846);
not NOT1 (N8713, N8712);
xor XOR2 (N8714, N8700, N8036);
buf BUF1 (N8715, N8713);
not NOT1 (N8716, N8694);
buf BUF1 (N8717, N8704);
xor XOR2 (N8718, N8684, N2964);
buf BUF1 (N8719, N8711);
or OR2 (N8720, N8709, N1489);
xor XOR2 (N8721, N8716, N326);
or OR2 (N8722, N8720, N3014);
and AND3 (N8723, N8715, N2888, N1066);
xor XOR2 (N8724, N8722, N7703);
nand NAND2 (N8725, N8719, N8124);
and AND2 (N8726, N8707, N4614);
buf BUF1 (N8727, N8717);
or OR3 (N8728, N8726, N917, N3026);
buf BUF1 (N8729, N8724);
not NOT1 (N8730, N8721);
not NOT1 (N8731, N8710);
nand NAND4 (N8732, N8729, N1528, N6086, N5243);
buf BUF1 (N8733, N8725);
or OR4 (N8734, N8727, N5268, N651, N3381);
and AND4 (N8735, N8733, N6741, N3840, N2356);
not NOT1 (N8736, N8735);
not NOT1 (N8737, N8723);
buf BUF1 (N8738, N8708);
buf BUF1 (N8739, N8734);
buf BUF1 (N8740, N8737);
or OR2 (N8741, N8731, N2210);
nor NOR4 (N8742, N8714, N4539, N7751, N4476);
and AND2 (N8743, N8741, N3423);
and AND4 (N8744, N8732, N4027, N5042, N7429);
not NOT1 (N8745, N8728);
xor XOR2 (N8746, N8738, N3117);
or OR2 (N8747, N8742, N2479);
nor NOR3 (N8748, N8743, N4590, N5974);
and AND4 (N8749, N8740, N95, N2256, N152);
nor NOR3 (N8750, N8745, N1972, N118);
nor NOR4 (N8751, N8744, N1329, N503, N985);
xor XOR2 (N8752, N8748, N5373);
not NOT1 (N8753, N8736);
and AND2 (N8754, N8718, N8508);
and AND3 (N8755, N8750, N7271, N5122);
or OR4 (N8756, N8747, N8357, N6599, N2421);
buf BUF1 (N8757, N8754);
not NOT1 (N8758, N8752);
and AND4 (N8759, N8755, N4439, N5572, N1210);
xor XOR2 (N8760, N8749, N2289);
buf BUF1 (N8761, N8758);
or OR3 (N8762, N8746, N1565, N4294);
xor XOR2 (N8763, N8739, N3137);
nand NAND3 (N8764, N8761, N7801, N8572);
not NOT1 (N8765, N8756);
buf BUF1 (N8766, N8764);
nand NAND3 (N8767, N8730, N2876, N5079);
buf BUF1 (N8768, N8762);
and AND4 (N8769, N8759, N6786, N4809, N4174);
nand NAND2 (N8770, N8765, N5782);
and AND4 (N8771, N8751, N2361, N2460, N6726);
or OR4 (N8772, N8770, N265, N990, N5456);
buf BUF1 (N8773, N8766);
and AND2 (N8774, N8753, N4781);
buf BUF1 (N8775, N8763);
buf BUF1 (N8776, N8771);
nand NAND4 (N8777, N8772, N1631, N2728, N7867);
nor NOR3 (N8778, N8775, N5947, N753);
and AND3 (N8779, N8777, N3195, N628);
or OR2 (N8780, N8779, N2831);
nand NAND4 (N8781, N8757, N6240, N2692, N1065);
not NOT1 (N8782, N8774);
xor XOR2 (N8783, N8769, N5530);
buf BUF1 (N8784, N8776);
and AND3 (N8785, N8760, N586, N6210);
or OR2 (N8786, N8785, N3430);
nor NOR3 (N8787, N8781, N6611, N1639);
buf BUF1 (N8788, N8786);
nand NAND3 (N8789, N8768, N8568, N5788);
nor NOR3 (N8790, N8783, N3299, N2715);
xor XOR2 (N8791, N8788, N7904);
not NOT1 (N8792, N8780);
nand NAND2 (N8793, N8778, N5557);
not NOT1 (N8794, N8791);
xor XOR2 (N8795, N8787, N418);
nor NOR2 (N8796, N8795, N2254);
xor XOR2 (N8797, N8767, N7368);
nand NAND3 (N8798, N8789, N752, N3848);
not NOT1 (N8799, N8793);
or OR4 (N8800, N8798, N7750, N8758, N6959);
or OR3 (N8801, N8784, N7234, N1100);
and AND4 (N8802, N8773, N4811, N8590, N1925);
nand NAND2 (N8803, N8797, N8081);
buf BUF1 (N8804, N8803);
not NOT1 (N8805, N8802);
nor NOR4 (N8806, N8801, N1849, N4275, N5155);
xor XOR2 (N8807, N8806, N1852);
or OR2 (N8808, N8805, N1779);
buf BUF1 (N8809, N8799);
buf BUF1 (N8810, N8809);
nor NOR4 (N8811, N8794, N8497, N2439, N2199);
buf BUF1 (N8812, N8792);
buf BUF1 (N8813, N8790);
nand NAND2 (N8814, N8813, N6309);
buf BUF1 (N8815, N8807);
or OR3 (N8816, N8796, N5482, N348);
or OR4 (N8817, N8815, N1706, N4822, N670);
or OR4 (N8818, N8812, N4898, N5215, N1219);
xor XOR2 (N8819, N8817, N637);
buf BUF1 (N8820, N8800);
nand NAND4 (N8821, N8819, N4272, N2507, N7731);
not NOT1 (N8822, N8811);
buf BUF1 (N8823, N8821);
or OR2 (N8824, N8804, N4788);
not NOT1 (N8825, N8814);
xor XOR2 (N8826, N8820, N4602);
or OR4 (N8827, N8782, N3626, N7662, N7222);
xor XOR2 (N8828, N8827, N2687);
nor NOR2 (N8829, N8825, N7324);
not NOT1 (N8830, N8816);
or OR3 (N8831, N8824, N8108, N4866);
nor NOR3 (N8832, N8818, N2928, N1155);
xor XOR2 (N8833, N8832, N3408);
buf BUF1 (N8834, N8828);
and AND4 (N8835, N8829, N610, N2729, N3533);
xor XOR2 (N8836, N8830, N1947);
buf BUF1 (N8837, N8831);
not NOT1 (N8838, N8836);
nand NAND3 (N8839, N8838, N2646, N7696);
buf BUF1 (N8840, N8834);
or OR4 (N8841, N8826, N3108, N3659, N1993);
or OR2 (N8842, N8840, N26);
or OR4 (N8843, N8823, N5734, N3386, N2907);
or OR4 (N8844, N8822, N6316, N3931, N1981);
not NOT1 (N8845, N8843);
or OR2 (N8846, N8841, N3592);
xor XOR2 (N8847, N8837, N4619);
and AND2 (N8848, N8844, N2458);
nor NOR2 (N8849, N8846, N2568);
and AND2 (N8850, N8845, N6676);
nand NAND3 (N8851, N8808, N4288, N7041);
nand NAND4 (N8852, N8850, N4487, N6338, N1880);
nand NAND3 (N8853, N8852, N8737, N6162);
buf BUF1 (N8854, N8847);
nand NAND4 (N8855, N8851, N6264, N4245, N6432);
nand NAND3 (N8856, N8842, N7996, N895);
and AND3 (N8857, N8854, N8764, N8661);
nor NOR2 (N8858, N8810, N936);
or OR4 (N8859, N8835, N5527, N7055, N2682);
nand NAND2 (N8860, N8858, N2838);
not NOT1 (N8861, N8856);
and AND4 (N8862, N8833, N4168, N5667, N5774);
and AND2 (N8863, N8859, N3367);
and AND3 (N8864, N8860, N6534, N8769);
not NOT1 (N8865, N8855);
or OR3 (N8866, N8865, N5613, N3393);
buf BUF1 (N8867, N8857);
nor NOR3 (N8868, N8867, N5471, N7822);
xor XOR2 (N8869, N8853, N1368);
buf BUF1 (N8870, N8849);
and AND2 (N8871, N8861, N1986);
or OR4 (N8872, N8839, N3302, N6333, N7524);
and AND2 (N8873, N8864, N4391);
buf BUF1 (N8874, N8868);
xor XOR2 (N8875, N8863, N2048);
nand NAND2 (N8876, N8862, N8404);
and AND2 (N8877, N8869, N864);
xor XOR2 (N8878, N8875, N731);
and AND4 (N8879, N8871, N7915, N8469, N8282);
or OR2 (N8880, N8879, N4778);
nor NOR3 (N8881, N8878, N1650, N8861);
buf BUF1 (N8882, N8877);
nor NOR4 (N8883, N8881, N7708, N8708, N1771);
xor XOR2 (N8884, N8882, N6235);
xor XOR2 (N8885, N8866, N4830);
buf BUF1 (N8886, N8874);
xor XOR2 (N8887, N8884, N8568);
xor XOR2 (N8888, N8876, N321);
nor NOR4 (N8889, N8887, N5816, N8242, N1517);
nor NOR3 (N8890, N8880, N7225, N1606);
nand NAND3 (N8891, N8870, N2689, N8544);
nor NOR2 (N8892, N8890, N3132);
buf BUF1 (N8893, N8885);
and AND2 (N8894, N8892, N7017);
xor XOR2 (N8895, N8893, N8003);
xor XOR2 (N8896, N8894, N5625);
nand NAND4 (N8897, N8883, N4763, N6762, N1294);
nand NAND4 (N8898, N8848, N64, N1824, N898);
and AND3 (N8899, N8898, N8399, N3530);
or OR2 (N8900, N8886, N8294);
nor NOR3 (N8901, N8900, N5759, N1321);
and AND4 (N8902, N8896, N6088, N8186, N2691);
nor NOR3 (N8903, N8872, N2078, N2248);
nand NAND4 (N8904, N8889, N931, N5793, N1065);
nor NOR4 (N8905, N8895, N5118, N3706, N7911);
buf BUF1 (N8906, N8888);
not NOT1 (N8907, N8873);
nor NOR2 (N8908, N8906, N188);
buf BUF1 (N8909, N8891);
or OR2 (N8910, N8909, N3395);
buf BUF1 (N8911, N8905);
and AND4 (N8912, N8897, N5306, N4122, N1075);
and AND4 (N8913, N8911, N7259, N4892, N3398);
xor XOR2 (N8914, N8901, N4918);
nor NOR2 (N8915, N8902, N8554);
buf BUF1 (N8916, N8912);
not NOT1 (N8917, N8916);
nand NAND2 (N8918, N8907, N1560);
and AND2 (N8919, N8915, N8180);
nor NOR4 (N8920, N8904, N5950, N6, N6963);
or OR3 (N8921, N8910, N5040, N8013);
nor NOR2 (N8922, N8921, N2407);
and AND4 (N8923, N8914, N4342, N4455, N5173);
or OR3 (N8924, N8908, N647, N6580);
not NOT1 (N8925, N8913);
not NOT1 (N8926, N8903);
or OR3 (N8927, N8923, N837, N4305);
xor XOR2 (N8928, N8922, N2200);
or OR3 (N8929, N8917, N8128, N1313);
buf BUF1 (N8930, N8926);
buf BUF1 (N8931, N8899);
buf BUF1 (N8932, N8919);
buf BUF1 (N8933, N8928);
and AND4 (N8934, N8918, N1970, N6003, N4831);
nor NOR3 (N8935, N8927, N8092, N1157);
or OR2 (N8936, N8934, N3088);
nand NAND4 (N8937, N8931, N6764, N1414, N507);
buf BUF1 (N8938, N8929);
nor NOR4 (N8939, N8932, N6929, N1630, N5290);
xor XOR2 (N8940, N8936, N5439);
and AND4 (N8941, N8930, N5710, N2702, N4894);
or OR2 (N8942, N8933, N6864);
xor XOR2 (N8943, N8940, N3210);
buf BUF1 (N8944, N8942);
buf BUF1 (N8945, N8935);
not NOT1 (N8946, N8944);
not NOT1 (N8947, N8924);
not NOT1 (N8948, N8937);
nand NAND3 (N8949, N8941, N3381, N768);
or OR3 (N8950, N8938, N4360, N7932);
nor NOR4 (N8951, N8943, N2583, N532, N6323);
or OR3 (N8952, N8920, N1852, N6037);
nand NAND3 (N8953, N8925, N6174, N3630);
nor NOR2 (N8954, N8948, N2642);
and AND2 (N8955, N8947, N1289);
not NOT1 (N8956, N8950);
buf BUF1 (N8957, N8939);
xor XOR2 (N8958, N8946, N5454);
and AND2 (N8959, N8953, N6844);
nand NAND3 (N8960, N8957, N7239, N4006);
xor XOR2 (N8961, N8954, N8406);
or OR3 (N8962, N8951, N8817, N5138);
nand NAND3 (N8963, N8962, N5063, N3172);
xor XOR2 (N8964, N8956, N450);
nand NAND2 (N8965, N8958, N5514);
buf BUF1 (N8966, N8961);
and AND4 (N8967, N8952, N2886, N8369, N6750);
buf BUF1 (N8968, N8949);
xor XOR2 (N8969, N8968, N612);
or OR2 (N8970, N8963, N7657);
xor XOR2 (N8971, N8959, N1819);
and AND3 (N8972, N8960, N5155, N4012);
nand NAND4 (N8973, N8964, N8210, N5111, N6107);
xor XOR2 (N8974, N8967, N8971);
nor NOR2 (N8975, N894, N3562);
nand NAND3 (N8976, N8970, N2448, N3085);
xor XOR2 (N8977, N8976, N1945);
xor XOR2 (N8978, N8965, N2631);
nor NOR2 (N8979, N8975, N1323);
nand NAND3 (N8980, N8973, N1226, N760);
or OR3 (N8981, N8980, N4514, N6833);
not NOT1 (N8982, N8978);
and AND3 (N8983, N8972, N6424, N4410);
buf BUF1 (N8984, N8979);
nand NAND2 (N8985, N8984, N2372);
xor XOR2 (N8986, N8985, N5017);
nand NAND2 (N8987, N8966, N6648);
buf BUF1 (N8988, N8955);
or OR3 (N8989, N8983, N7458, N3772);
nor NOR2 (N8990, N8974, N6366);
or OR2 (N8991, N8988, N5994);
buf BUF1 (N8992, N8987);
buf BUF1 (N8993, N8945);
xor XOR2 (N8994, N8991, N5822);
or OR4 (N8995, N8989, N5734, N5558, N7323);
or OR4 (N8996, N8994, N5198, N86, N630);
and AND2 (N8997, N8993, N3180);
not NOT1 (N8998, N8981);
and AND2 (N8999, N8977, N5490);
nand NAND4 (N9000, N8998, N7110, N2647, N2019);
not NOT1 (N9001, N8999);
or OR2 (N9002, N8997, N845);
and AND2 (N9003, N8996, N2381);
xor XOR2 (N9004, N8995, N5029);
nor NOR3 (N9005, N9003, N8420, N2193);
buf BUF1 (N9006, N9004);
or OR3 (N9007, N8986, N110, N2276);
not NOT1 (N9008, N9002);
not NOT1 (N9009, N9001);
nor NOR2 (N9010, N8990, N3315);
buf BUF1 (N9011, N9006);
xor XOR2 (N9012, N9000, N4611);
and AND2 (N9013, N8982, N6358);
or OR4 (N9014, N9008, N3517, N2231, N5523);
or OR4 (N9015, N9005, N6333, N914, N6206);
xor XOR2 (N9016, N8992, N8641);
not NOT1 (N9017, N9007);
buf BUF1 (N9018, N9012);
or OR2 (N9019, N9011, N3194);
nand NAND2 (N9020, N9015, N7787);
or OR2 (N9021, N9018, N2085);
and AND4 (N9022, N9016, N5048, N63, N3534);
nor NOR4 (N9023, N9021, N7661, N7637, N6861);
xor XOR2 (N9024, N9017, N2312);
or OR2 (N9025, N9014, N3605);
not NOT1 (N9026, N9025);
and AND2 (N9027, N9026, N5483);
xor XOR2 (N9028, N9023, N457);
or OR2 (N9029, N9027, N2128);
and AND4 (N9030, N9019, N3939, N1498, N1392);
buf BUF1 (N9031, N9022);
not NOT1 (N9032, N9020);
nor NOR3 (N9033, N9032, N8792, N7284);
xor XOR2 (N9034, N9029, N3750);
buf BUF1 (N9035, N9034);
and AND2 (N9036, N9024, N8706);
and AND2 (N9037, N9013, N7741);
nand NAND2 (N9038, N9030, N1150);
xor XOR2 (N9039, N9035, N8140);
not NOT1 (N9040, N9038);
nand NAND4 (N9041, N9031, N879, N5767, N5838);
and AND4 (N9042, N8969, N6748, N1436, N284);
not NOT1 (N9043, N9036);
or OR3 (N9044, N9043, N1174, N1279);
not NOT1 (N9045, N9040);
xor XOR2 (N9046, N9010, N4401);
buf BUF1 (N9047, N9037);
buf BUF1 (N9048, N9047);
xor XOR2 (N9049, N9042, N7112);
and AND2 (N9050, N9033, N251);
xor XOR2 (N9051, N9044, N4611);
nand NAND2 (N9052, N9041, N7848);
nand NAND2 (N9053, N9049, N7016);
nand NAND4 (N9054, N9039, N4480, N6342, N8987);
and AND2 (N9055, N9053, N4299);
or OR3 (N9056, N9028, N389, N3070);
nand NAND4 (N9057, N9054, N448, N3938, N1143);
and AND4 (N9058, N9048, N708, N6692, N7303);
and AND3 (N9059, N9055, N7467, N3420);
nor NOR3 (N9060, N9056, N8388, N8459);
and AND3 (N9061, N9046, N8091, N4509);
xor XOR2 (N9062, N9058, N2689);
not NOT1 (N9063, N9050);
or OR4 (N9064, N9060, N2361, N6873, N1264);
nand NAND2 (N9065, N9045, N1696);
not NOT1 (N9066, N9061);
xor XOR2 (N9067, N9066, N7182);
not NOT1 (N9068, N9059);
buf BUF1 (N9069, N9068);
nand NAND2 (N9070, N9067, N4844);
or OR3 (N9071, N9009, N4640, N421);
not NOT1 (N9072, N9064);
and AND4 (N9073, N9063, N2303, N5990, N2313);
buf BUF1 (N9074, N9057);
nor NOR4 (N9075, N9069, N4614, N3250, N2918);
or OR3 (N9076, N9074, N559, N2981);
nand NAND3 (N9077, N9052, N7923, N247);
or OR3 (N9078, N9051, N297, N236);
xor XOR2 (N9079, N9071, N7906);
xor XOR2 (N9080, N9062, N3444);
xor XOR2 (N9081, N9072, N3423);
nor NOR2 (N9082, N9075, N323);
xor XOR2 (N9083, N9076, N5060);
xor XOR2 (N9084, N9080, N4550);
nand NAND4 (N9085, N9065, N6599, N1014, N7824);
or OR3 (N9086, N9083, N2365, N7085);
or OR2 (N9087, N9086, N8561);
nor NOR3 (N9088, N9079, N5009, N9087);
not NOT1 (N9089, N761);
buf BUF1 (N9090, N9085);
or OR2 (N9091, N9082, N8412);
not NOT1 (N9092, N9077);
and AND2 (N9093, N9073, N8168);
not NOT1 (N9094, N9092);
nor NOR3 (N9095, N9081, N8917, N6347);
xor XOR2 (N9096, N9084, N99);
not NOT1 (N9097, N9094);
buf BUF1 (N9098, N9091);
buf BUF1 (N9099, N9096);
xor XOR2 (N9100, N9098, N5026);
buf BUF1 (N9101, N9070);
xor XOR2 (N9102, N9090, N3321);
and AND2 (N9103, N9099, N7482);
or OR2 (N9104, N9093, N7496);
and AND4 (N9105, N9103, N4354, N3065, N1461);
nor NOR2 (N9106, N9078, N5470);
nand NAND3 (N9107, N9097, N807, N7277);
nand NAND3 (N9108, N9089, N3484, N2919);
xor XOR2 (N9109, N9088, N4964);
not NOT1 (N9110, N9105);
buf BUF1 (N9111, N9107);
nand NAND4 (N9112, N9100, N5224, N6246, N5257);
not NOT1 (N9113, N9112);
nor NOR2 (N9114, N9108, N7499);
xor XOR2 (N9115, N9106, N2562);
nand NAND4 (N9116, N9095, N2413, N4501, N8626);
not NOT1 (N9117, N9102);
not NOT1 (N9118, N9114);
or OR2 (N9119, N9113, N2878);
or OR4 (N9120, N9111, N3023, N2879, N2423);
or OR4 (N9121, N9120, N948, N8033, N1878);
or OR4 (N9122, N9121, N2151, N6012, N6669);
xor XOR2 (N9123, N9101, N5532);
not NOT1 (N9124, N9115);
not NOT1 (N9125, N9123);
xor XOR2 (N9126, N9117, N3066);
not NOT1 (N9127, N9109);
or OR3 (N9128, N9127, N3051, N1331);
xor XOR2 (N9129, N9124, N3367);
or OR4 (N9130, N9125, N925, N7982, N6931);
nand NAND4 (N9131, N9126, N7609, N5199, N7190);
not NOT1 (N9132, N9119);
xor XOR2 (N9133, N9132, N8902);
nor NOR2 (N9134, N9128, N1765);
nand NAND4 (N9135, N9116, N491, N5992, N2783);
nor NOR4 (N9136, N9122, N7178, N2534, N4335);
nor NOR2 (N9137, N9136, N2741);
nand NAND2 (N9138, N9110, N1063);
nand NAND3 (N9139, N9133, N5045, N5085);
xor XOR2 (N9140, N9134, N1127);
or OR3 (N9141, N9118, N8481, N9044);
and AND2 (N9142, N9104, N4746);
nor NOR4 (N9143, N9138, N4451, N3781, N9091);
buf BUF1 (N9144, N9129);
nand NAND2 (N9145, N9144, N7198);
or OR2 (N9146, N9137, N8240);
xor XOR2 (N9147, N9145, N8393);
and AND3 (N9148, N9131, N4977, N5325);
nand NAND4 (N9149, N9147, N2492, N5254, N168);
xor XOR2 (N9150, N9146, N2933);
nand NAND2 (N9151, N9130, N2567);
or OR4 (N9152, N9141, N6394, N5161, N7845);
and AND2 (N9153, N9140, N5697);
nand NAND3 (N9154, N9149, N1790, N577);
not NOT1 (N9155, N9150);
nand NAND4 (N9156, N9155, N462, N5583, N2289);
or OR4 (N9157, N9156, N5248, N1574, N5716);
buf BUF1 (N9158, N9151);
or OR4 (N9159, N9148, N7089, N8652, N499);
and AND3 (N9160, N9154, N7747, N5021);
not NOT1 (N9161, N9143);
and AND3 (N9162, N9157, N3188, N6206);
buf BUF1 (N9163, N9160);
nand NAND3 (N9164, N9152, N1513, N5552);
or OR2 (N9165, N9163, N7947);
xor XOR2 (N9166, N9153, N8164);
buf BUF1 (N9167, N9139);
or OR3 (N9168, N9164, N3787, N133);
nand NAND2 (N9169, N9168, N142);
or OR2 (N9170, N9159, N5409);
nor NOR4 (N9171, N9170, N7986, N3559, N5394);
buf BUF1 (N9172, N9142);
or OR3 (N9173, N9162, N8140, N2273);
nor NOR4 (N9174, N9166, N1843, N5405, N701);
buf BUF1 (N9175, N9165);
or OR4 (N9176, N9174, N3104, N6992, N4597);
xor XOR2 (N9177, N9171, N6437);
or OR2 (N9178, N9177, N7809);
nor NOR2 (N9179, N9167, N7029);
xor XOR2 (N9180, N9161, N2639);
and AND2 (N9181, N9175, N3691);
xor XOR2 (N9182, N9179, N3366);
nand NAND3 (N9183, N9173, N5426, N2163);
nand NAND2 (N9184, N9183, N707);
not NOT1 (N9185, N9169);
and AND3 (N9186, N9178, N6410, N2126);
xor XOR2 (N9187, N9184, N9066);
nor NOR2 (N9188, N9185, N6789);
not NOT1 (N9189, N9182);
and AND2 (N9190, N9188, N1388);
and AND3 (N9191, N9190, N4936, N3462);
xor XOR2 (N9192, N9176, N3533);
not NOT1 (N9193, N9186);
or OR3 (N9194, N9172, N1341, N5929);
buf BUF1 (N9195, N9191);
xor XOR2 (N9196, N9181, N2429);
not NOT1 (N9197, N9135);
and AND2 (N9198, N9187, N1701);
not NOT1 (N9199, N9195);
or OR3 (N9200, N9194, N6299, N9006);
and AND2 (N9201, N9189, N9134);
nor NOR3 (N9202, N9193, N8945, N7091);
nand NAND3 (N9203, N9197, N756, N6271);
buf BUF1 (N9204, N9196);
nand NAND4 (N9205, N9180, N7472, N4458, N5038);
not NOT1 (N9206, N9199);
or OR3 (N9207, N9205, N7642, N2943);
or OR4 (N9208, N9202, N6502, N850, N2236);
and AND3 (N9209, N9203, N8753, N4584);
xor XOR2 (N9210, N9208, N3938);
and AND2 (N9211, N9209, N4594);
nor NOR2 (N9212, N9204, N3380);
not NOT1 (N9213, N9201);
nor NOR3 (N9214, N9192, N3084, N6573);
xor XOR2 (N9215, N9210, N5184);
buf BUF1 (N9216, N9214);
not NOT1 (N9217, N9216);
buf BUF1 (N9218, N9198);
not NOT1 (N9219, N9206);
or OR3 (N9220, N9207, N8799, N9192);
xor XOR2 (N9221, N9158, N7519);
nor NOR4 (N9222, N9218, N45, N1743, N5230);
buf BUF1 (N9223, N9212);
nor NOR4 (N9224, N9222, N90, N6993, N9089);
nor NOR2 (N9225, N9221, N4851);
or OR2 (N9226, N9200, N5657);
xor XOR2 (N9227, N9220, N8514);
and AND4 (N9228, N9211, N1028, N9003, N6943);
and AND2 (N9229, N9213, N5943);
or OR2 (N9230, N9226, N6457);
nand NAND3 (N9231, N9224, N5192, N4464);
nor NOR3 (N9232, N9229, N3202, N668);
nand NAND3 (N9233, N9228, N1164, N3327);
buf BUF1 (N9234, N9225);
xor XOR2 (N9235, N9232, N267);
xor XOR2 (N9236, N9219, N1734);
buf BUF1 (N9237, N9227);
or OR3 (N9238, N9223, N630, N8329);
buf BUF1 (N9239, N9234);
and AND3 (N9240, N9237, N8388, N7586);
nor NOR2 (N9241, N9215, N3665);
buf BUF1 (N9242, N9240);
nor NOR4 (N9243, N9233, N8160, N5120, N5936);
buf BUF1 (N9244, N9217);
buf BUF1 (N9245, N9238);
not NOT1 (N9246, N9239);
buf BUF1 (N9247, N9235);
and AND2 (N9248, N9230, N1570);
xor XOR2 (N9249, N9248, N3050);
buf BUF1 (N9250, N9244);
and AND4 (N9251, N9247, N4011, N4942, N5143);
buf BUF1 (N9252, N9242);
nor NOR2 (N9253, N9249, N2824);
buf BUF1 (N9254, N9241);
xor XOR2 (N9255, N9245, N3257);
xor XOR2 (N9256, N9252, N4104);
buf BUF1 (N9257, N9253);
nand NAND4 (N9258, N9257, N4992, N1406, N2430);
or OR2 (N9259, N9255, N7759);
not NOT1 (N9260, N9250);
and AND4 (N9261, N9259, N1815, N1747, N5077);
not NOT1 (N9262, N9236);
nor NOR3 (N9263, N9254, N7629, N8008);
or OR2 (N9264, N9256, N8315);
nand NAND3 (N9265, N9258, N6367, N6636);
nand NAND2 (N9266, N9261, N8556);
nand NAND4 (N9267, N9251, N6481, N8698, N4792);
buf BUF1 (N9268, N9267);
buf BUF1 (N9269, N9260);
not NOT1 (N9270, N9263);
and AND3 (N9271, N9265, N6198, N1632);
nand NAND3 (N9272, N9270, N9182, N3603);
nor NOR3 (N9273, N9269, N3463, N2013);
xor XOR2 (N9274, N9264, N945);
and AND2 (N9275, N9246, N5340);
or OR2 (N9276, N9272, N5359);
and AND2 (N9277, N9271, N599);
nand NAND3 (N9278, N9277, N1540, N97);
nand NAND3 (N9279, N9231, N5050, N7750);
and AND4 (N9280, N9262, N6972, N4960, N1996);
xor XOR2 (N9281, N9279, N3998);
and AND3 (N9282, N9243, N3419, N5985);
xor XOR2 (N9283, N9281, N6715);
xor XOR2 (N9284, N9283, N8957);
and AND4 (N9285, N9274, N7369, N6891, N4299);
buf BUF1 (N9286, N9275);
xor XOR2 (N9287, N9268, N8339);
and AND4 (N9288, N9278, N1627, N6870, N3808);
nor NOR2 (N9289, N9280, N3391);
and AND2 (N9290, N9273, N8004);
buf BUF1 (N9291, N9266);
or OR2 (N9292, N9288, N5393);
buf BUF1 (N9293, N9282);
nand NAND2 (N9294, N9289, N7472);
nand NAND3 (N9295, N9294, N9179, N6089);
buf BUF1 (N9296, N9284);
or OR4 (N9297, N9292, N4426, N1563, N2168);
nor NOR3 (N9298, N9276, N1515, N2953);
xor XOR2 (N9299, N9285, N7199);
nor NOR3 (N9300, N9287, N6485, N719);
nand NAND3 (N9301, N9299, N5547, N914);
and AND4 (N9302, N9293, N5009, N9295, N6197);
buf BUF1 (N9303, N1642);
nor NOR3 (N9304, N9301, N7591, N2468);
and AND2 (N9305, N9290, N3365);
nand NAND4 (N9306, N9298, N4261, N2400, N5914);
not NOT1 (N9307, N9303);
nand NAND2 (N9308, N9305, N5673);
buf BUF1 (N9309, N9300);
nand NAND4 (N9310, N9291, N808, N3088, N7538);
or OR2 (N9311, N9307, N9022);
and AND2 (N9312, N9302, N5102);
nor NOR2 (N9313, N9306, N8327);
or OR4 (N9314, N9309, N3147, N5269, N8931);
buf BUF1 (N9315, N9311);
buf BUF1 (N9316, N9312);
nor NOR2 (N9317, N9310, N2222);
and AND4 (N9318, N9296, N5980, N7975, N3884);
and AND4 (N9319, N9313, N1808, N587, N7477);
nor NOR3 (N9320, N9314, N215, N1037);
not NOT1 (N9321, N9297);
nor NOR2 (N9322, N9318, N6391);
and AND3 (N9323, N9319, N1706, N6919);
xor XOR2 (N9324, N9322, N3651);
nand NAND2 (N9325, N9320, N8865);
buf BUF1 (N9326, N9304);
xor XOR2 (N9327, N9286, N2964);
nor NOR4 (N9328, N9324, N8788, N159, N649);
buf BUF1 (N9329, N9316);
not NOT1 (N9330, N9321);
and AND2 (N9331, N9329, N6310);
and AND3 (N9332, N9326, N8704, N5596);
and AND4 (N9333, N9331, N442, N6383, N6520);
or OR4 (N9334, N9308, N5210, N1882, N3724);
or OR3 (N9335, N9327, N6835, N6365);
and AND4 (N9336, N9317, N6350, N434, N4386);
nand NAND3 (N9337, N9323, N5011, N8890);
not NOT1 (N9338, N9336);
xor XOR2 (N9339, N9330, N5259);
xor XOR2 (N9340, N9339, N6539);
and AND4 (N9341, N9337, N1640, N3033, N6274);
nor NOR2 (N9342, N9341, N1098);
and AND4 (N9343, N9328, N7642, N6158, N6298);
not NOT1 (N9344, N9342);
nand NAND3 (N9345, N9344, N2307, N7148);
or OR3 (N9346, N9338, N2577, N2656);
nor NOR2 (N9347, N9333, N3593);
not NOT1 (N9348, N9332);
buf BUF1 (N9349, N9347);
and AND4 (N9350, N9325, N1611, N8185, N4825);
not NOT1 (N9351, N9340);
or OR2 (N9352, N9346, N7800);
nor NOR3 (N9353, N9349, N4772, N2488);
nor NOR4 (N9354, N9315, N6797, N2449, N4499);
not NOT1 (N9355, N9334);
nor NOR4 (N9356, N9355, N3201, N348, N5757);
nor NOR4 (N9357, N9335, N4254, N3802, N2072);
nor NOR3 (N9358, N9351, N4227, N2469);
or OR3 (N9359, N9358, N6038, N5438);
nor NOR3 (N9360, N9343, N2091, N6256);
xor XOR2 (N9361, N9357, N2537);
xor XOR2 (N9362, N9350, N4211);
buf BUF1 (N9363, N9352);
not NOT1 (N9364, N9345);
nand NAND4 (N9365, N9356, N4965, N6753, N5772);
or OR2 (N9366, N9354, N1490);
buf BUF1 (N9367, N9365);
buf BUF1 (N9368, N9366);
not NOT1 (N9369, N9367);
nor NOR4 (N9370, N9368, N4770, N7002, N5538);
buf BUF1 (N9371, N9359);
nand NAND2 (N9372, N9371, N5624);
nand NAND4 (N9373, N9353, N3244, N8002, N6399);
not NOT1 (N9374, N9369);
not NOT1 (N9375, N9370);
not NOT1 (N9376, N9373);
and AND4 (N9377, N9363, N3219, N7253, N3260);
or OR2 (N9378, N9364, N2836);
not NOT1 (N9379, N9362);
nand NAND3 (N9380, N9361, N6834, N7766);
not NOT1 (N9381, N9380);
and AND2 (N9382, N9348, N7181);
nor NOR2 (N9383, N9382, N4939);
and AND2 (N9384, N9377, N753);
and AND4 (N9385, N9381, N1791, N67, N8498);
and AND4 (N9386, N9372, N8482, N3546, N3535);
buf BUF1 (N9387, N9374);
or OR2 (N9388, N9386, N3366);
not NOT1 (N9389, N9384);
not NOT1 (N9390, N9379);
nand NAND2 (N9391, N9375, N3933);
xor XOR2 (N9392, N9389, N7702);
and AND2 (N9393, N9390, N808);
nand NAND3 (N9394, N9392, N5396, N7764);
and AND3 (N9395, N9393, N4477, N1759);
nand NAND3 (N9396, N9388, N3566, N2474);
xor XOR2 (N9397, N9383, N1983);
not NOT1 (N9398, N9394);
buf BUF1 (N9399, N9378);
nor NOR2 (N9400, N9396, N7432);
and AND3 (N9401, N9387, N6926, N5212);
not NOT1 (N9402, N9397);
and AND3 (N9403, N9376, N1200, N591);
buf BUF1 (N9404, N9360);
or OR3 (N9405, N9401, N6773, N2357);
nand NAND4 (N9406, N9395, N4704, N1950, N7913);
and AND3 (N9407, N9403, N7686, N8898);
nor NOR3 (N9408, N9398, N1803, N777);
xor XOR2 (N9409, N9391, N2561);
not NOT1 (N9410, N9405);
nor NOR4 (N9411, N9409, N7717, N5360, N1492);
not NOT1 (N9412, N9402);
not NOT1 (N9413, N9411);
xor XOR2 (N9414, N9413, N9027);
and AND4 (N9415, N9385, N2250, N3198, N1748);
and AND2 (N9416, N9407, N1928);
nand NAND2 (N9417, N9414, N3058);
nand NAND3 (N9418, N9412, N1949, N8399);
buf BUF1 (N9419, N9415);
and AND3 (N9420, N9400, N5358, N5417);
or OR4 (N9421, N9404, N8414, N1224, N3147);
or OR3 (N9422, N9416, N2112, N6375);
buf BUF1 (N9423, N9399);
and AND4 (N9424, N9418, N3481, N5710, N2893);
not NOT1 (N9425, N9417);
and AND4 (N9426, N9408, N3011, N5593, N3625);
or OR2 (N9427, N9421, N5810);
buf BUF1 (N9428, N9425);
not NOT1 (N9429, N9423);
not NOT1 (N9430, N9406);
and AND4 (N9431, N9430, N8144, N820, N572);
and AND3 (N9432, N9410, N8734, N2936);
or OR2 (N9433, N9426, N5194);
or OR4 (N9434, N9431, N6328, N5135, N7509);
nor NOR2 (N9435, N9419, N1632);
xor XOR2 (N9436, N9432, N8489);
buf BUF1 (N9437, N9428);
not NOT1 (N9438, N9433);
nor NOR3 (N9439, N9429, N6874, N8327);
or OR3 (N9440, N9420, N392, N4949);
nand NAND3 (N9441, N9439, N1100, N970);
or OR3 (N9442, N9435, N2670, N5108);
and AND4 (N9443, N9424, N4073, N8655, N1710);
nor NOR4 (N9444, N9437, N2875, N4686, N5412);
xor XOR2 (N9445, N9438, N7107);
or OR4 (N9446, N9445, N6715, N3899, N5202);
xor XOR2 (N9447, N9436, N7873);
xor XOR2 (N9448, N9427, N1126);
xor XOR2 (N9449, N9441, N776);
nand NAND4 (N9450, N9447, N3248, N8897, N1045);
nand NAND3 (N9451, N9422, N5527, N3681);
or OR3 (N9452, N9450, N782, N5180);
buf BUF1 (N9453, N9434);
buf BUF1 (N9454, N9440);
buf BUF1 (N9455, N9444);
nor NOR2 (N9456, N9454, N5834);
buf BUF1 (N9457, N9449);
nor NOR2 (N9458, N9448, N3940);
and AND2 (N9459, N9446, N5547);
nor NOR4 (N9460, N9457, N3227, N5913, N1405);
or OR3 (N9461, N9451, N4570, N4377);
xor XOR2 (N9462, N9452, N5865);
and AND2 (N9463, N9455, N8381);
and AND3 (N9464, N9443, N1303, N8169);
and AND2 (N9465, N9461, N7228);
xor XOR2 (N9466, N9462, N4468);
and AND2 (N9467, N9463, N8095);
buf BUF1 (N9468, N9458);
xor XOR2 (N9469, N9464, N39);
and AND4 (N9470, N9460, N7248, N2569, N4226);
not NOT1 (N9471, N9467);
xor XOR2 (N9472, N9456, N5057);
xor XOR2 (N9473, N9472, N7515);
or OR2 (N9474, N9469, N4699);
nor NOR4 (N9475, N9465, N3072, N7804, N1789);
buf BUF1 (N9476, N9470);
or OR2 (N9477, N9473, N4091);
nor NOR4 (N9478, N9471, N1243, N7029, N137);
not NOT1 (N9479, N9474);
nand NAND4 (N9480, N9442, N3724, N8481, N5276);
or OR2 (N9481, N9475, N723);
and AND3 (N9482, N9480, N2950, N761);
nor NOR4 (N9483, N9466, N9115, N3519, N5509);
and AND4 (N9484, N9478, N612, N483, N1095);
nand NAND2 (N9485, N9482, N3638);
xor XOR2 (N9486, N9485, N4087);
or OR3 (N9487, N9476, N8828, N7776);
nor NOR2 (N9488, N9479, N5936);
not NOT1 (N9489, N9484);
or OR2 (N9490, N9486, N5087);
or OR4 (N9491, N9489, N3275, N7097, N3172);
xor XOR2 (N9492, N9459, N6488);
or OR3 (N9493, N9481, N6571, N670);
xor XOR2 (N9494, N9490, N7421);
buf BUF1 (N9495, N9494);
or OR3 (N9496, N9492, N5236, N6276);
and AND4 (N9497, N9487, N3109, N1306, N8295);
nand NAND2 (N9498, N9453, N6138);
or OR2 (N9499, N9497, N3522);
xor XOR2 (N9500, N9496, N762);
xor XOR2 (N9501, N9495, N7476);
or OR3 (N9502, N9498, N9173, N9041);
or OR4 (N9503, N9493, N3266, N1983, N4921);
not NOT1 (N9504, N9499);
and AND3 (N9505, N9477, N2447, N9258);
nand NAND2 (N9506, N9505, N7007);
buf BUF1 (N9507, N9504);
not NOT1 (N9508, N9506);
nand NAND3 (N9509, N9507, N5691, N2982);
nand NAND3 (N9510, N9501, N4556, N1315);
or OR2 (N9511, N9483, N2647);
nand NAND4 (N9512, N9508, N8429, N2974, N1847);
buf BUF1 (N9513, N9503);
not NOT1 (N9514, N9512);
xor XOR2 (N9515, N9511, N8660);
buf BUF1 (N9516, N9488);
or OR3 (N9517, N9500, N7490, N1016);
nor NOR3 (N9518, N9513, N4263, N4491);
buf BUF1 (N9519, N9514);
not NOT1 (N9520, N9519);
buf BUF1 (N9521, N9509);
buf BUF1 (N9522, N9520);
nand NAND2 (N9523, N9522, N7615);
nor NOR2 (N9524, N9515, N2182);
not NOT1 (N9525, N9524);
and AND2 (N9526, N9502, N9276);
and AND3 (N9527, N9491, N8082, N8377);
not NOT1 (N9528, N9525);
nand NAND2 (N9529, N9521, N5338);
nand NAND4 (N9530, N9517, N3076, N759, N1762);
nor NOR2 (N9531, N9510, N2732);
or OR3 (N9532, N9530, N3462, N7657);
or OR4 (N9533, N9468, N9325, N5059, N6782);
nor NOR4 (N9534, N9523, N3947, N5595, N1148);
nor NOR3 (N9535, N9532, N7416, N6796);
and AND2 (N9536, N9528, N3946);
xor XOR2 (N9537, N9533, N6421);
nor NOR2 (N9538, N9529, N6955);
nand NAND3 (N9539, N9537, N5477, N7960);
nor NOR3 (N9540, N9518, N2902, N6304);
nor NOR4 (N9541, N9540, N144, N5120, N5221);
not NOT1 (N9542, N9516);
not NOT1 (N9543, N9539);
and AND3 (N9544, N9538, N2609, N1683);
or OR2 (N9545, N9535, N2609);
nand NAND4 (N9546, N9541, N4943, N7380, N8217);
or OR3 (N9547, N9544, N5372, N7062);
xor XOR2 (N9548, N9534, N1825);
buf BUF1 (N9549, N9545);
or OR4 (N9550, N9542, N1452, N8780, N8458);
xor XOR2 (N9551, N9549, N7484);
or OR3 (N9552, N9546, N911, N7644);
nand NAND2 (N9553, N9552, N2592);
nand NAND2 (N9554, N9526, N8694);
nand NAND2 (N9555, N9551, N6055);
xor XOR2 (N9556, N9547, N9030);
nor NOR3 (N9557, N9556, N4443, N6745);
not NOT1 (N9558, N9527);
not NOT1 (N9559, N9536);
buf BUF1 (N9560, N9554);
or OR3 (N9561, N9543, N701, N8184);
xor XOR2 (N9562, N9561, N3303);
xor XOR2 (N9563, N9559, N5806);
xor XOR2 (N9564, N9553, N1936);
or OR2 (N9565, N9564, N2135);
not NOT1 (N9566, N9555);
nor NOR2 (N9567, N9565, N1596);
or OR4 (N9568, N9548, N8619, N2335, N1369);
buf BUF1 (N9569, N9562);
not NOT1 (N9570, N9531);
and AND4 (N9571, N9560, N4548, N2440, N7968);
or OR2 (N9572, N9550, N3414);
xor XOR2 (N9573, N9558, N6887);
buf BUF1 (N9574, N9567);
not NOT1 (N9575, N9573);
not NOT1 (N9576, N9571);
not NOT1 (N9577, N9563);
and AND2 (N9578, N9570, N4122);
not NOT1 (N9579, N9557);
buf BUF1 (N9580, N9574);
xor XOR2 (N9581, N9572, N4331);
or OR2 (N9582, N9581, N2930);
and AND4 (N9583, N9575, N1988, N576, N6245);
xor XOR2 (N9584, N9580, N7801);
buf BUF1 (N9585, N9584);
nor NOR4 (N9586, N9577, N5708, N1503, N3486);
nand NAND2 (N9587, N9586, N1140);
and AND2 (N9588, N9583, N4892);
nor NOR4 (N9589, N9568, N5002, N3708, N8635);
nor NOR2 (N9590, N9589, N7802);
nor NOR2 (N9591, N9590, N8455);
xor XOR2 (N9592, N9576, N5687);
nor NOR2 (N9593, N9591, N554);
xor XOR2 (N9594, N9592, N8774);
buf BUF1 (N9595, N9588);
not NOT1 (N9596, N9593);
nor NOR2 (N9597, N9585, N512);
nand NAND2 (N9598, N9582, N1911);
and AND4 (N9599, N9597, N836, N8371, N8841);
or OR4 (N9600, N9569, N4187, N9244, N7196);
nor NOR2 (N9601, N9578, N7900);
not NOT1 (N9602, N9601);
nor NOR4 (N9603, N9596, N7142, N8706, N7908);
or OR4 (N9604, N9587, N422, N4692, N946);
nor NOR4 (N9605, N9594, N8470, N3050, N9334);
or OR4 (N9606, N9598, N5930, N8203, N3673);
nand NAND3 (N9607, N9603, N7393, N2722);
xor XOR2 (N9608, N9566, N2537);
nand NAND4 (N9609, N9595, N1476, N8149, N7199);
nand NAND3 (N9610, N9607, N9387, N3451);
and AND3 (N9611, N9608, N2139, N2191);
nor NOR2 (N9612, N9579, N8566);
and AND2 (N9613, N9612, N2816);
and AND2 (N9614, N9600, N2712);
buf BUF1 (N9615, N9599);
buf BUF1 (N9616, N9605);
and AND4 (N9617, N9614, N4233, N9299, N3875);
buf BUF1 (N9618, N9613);
or OR3 (N9619, N9610, N3088, N6900);
nor NOR2 (N9620, N9619, N1124);
or OR2 (N9621, N9616, N6681);
buf BUF1 (N9622, N9606);
not NOT1 (N9623, N9620);
and AND4 (N9624, N9623, N4610, N5613, N3026);
xor XOR2 (N9625, N9615, N3167);
nor NOR3 (N9626, N9621, N8979, N3680);
nand NAND3 (N9627, N9602, N205, N3142);
nand NAND4 (N9628, N9609, N4698, N8014, N1473);
nand NAND2 (N9629, N9611, N3601);
buf BUF1 (N9630, N9604);
nand NAND2 (N9631, N9629, N7529);
buf BUF1 (N9632, N9630);
nor NOR2 (N9633, N9627, N5377);
or OR4 (N9634, N9632, N3950, N3502, N8332);
and AND3 (N9635, N9617, N8838, N9035);
buf BUF1 (N9636, N9618);
nor NOR4 (N9637, N9631, N7011, N2489, N5868);
or OR4 (N9638, N9622, N5835, N9557, N8359);
nor NOR2 (N9639, N9637, N7374);
or OR3 (N9640, N9636, N2102, N6545);
and AND3 (N9641, N9640, N742, N6882);
xor XOR2 (N9642, N9624, N2965);
xor XOR2 (N9643, N9642, N8617);
nor NOR3 (N9644, N9626, N6890, N6049);
or OR2 (N9645, N9633, N4835);
and AND2 (N9646, N9634, N8905);
xor XOR2 (N9647, N9628, N8601);
xor XOR2 (N9648, N9639, N638);
buf BUF1 (N9649, N9643);
or OR4 (N9650, N9649, N3735, N8271, N6983);
xor XOR2 (N9651, N9644, N869);
nand NAND2 (N9652, N9625, N4033);
nand NAND4 (N9653, N9650, N408, N655, N8622);
not NOT1 (N9654, N9648);
buf BUF1 (N9655, N9654);
nand NAND2 (N9656, N9647, N2105);
or OR3 (N9657, N9651, N1300, N2253);
xor XOR2 (N9658, N9646, N5058);
or OR4 (N9659, N9638, N895, N5858, N7753);
not NOT1 (N9660, N9659);
xor XOR2 (N9661, N9655, N2190);
xor XOR2 (N9662, N9653, N8325);
and AND4 (N9663, N9656, N8422, N2561, N5351);
nor NOR2 (N9664, N9658, N7810);
nor NOR3 (N9665, N9660, N1466, N3661);
or OR2 (N9666, N9635, N6076);
not NOT1 (N9667, N9664);
and AND2 (N9668, N9662, N8443);
or OR3 (N9669, N9645, N835, N3244);
and AND4 (N9670, N9652, N4616, N3849, N9522);
nor NOR4 (N9671, N9661, N2205, N2250, N8240);
xor XOR2 (N9672, N9665, N3464);
and AND4 (N9673, N9669, N2862, N3896, N6913);
and AND2 (N9674, N9671, N6498);
buf BUF1 (N9675, N9668);
nand NAND3 (N9676, N9667, N4467, N715);
nor NOR3 (N9677, N9676, N7648, N700);
or OR4 (N9678, N9677, N4591, N905, N4170);
nor NOR3 (N9679, N9672, N2870, N2737);
buf BUF1 (N9680, N9663);
and AND3 (N9681, N9680, N7617, N8095);
not NOT1 (N9682, N9678);
or OR2 (N9683, N9673, N6492);
nor NOR4 (N9684, N9670, N3716, N6188, N513);
buf BUF1 (N9685, N9641);
nor NOR2 (N9686, N9674, N9178);
nand NAND4 (N9687, N9675, N9462, N5233, N1324);
xor XOR2 (N9688, N9657, N224);
nor NOR3 (N9689, N9682, N9413, N2353);
xor XOR2 (N9690, N9688, N180);
nand NAND2 (N9691, N9679, N648);
or OR3 (N9692, N9666, N543, N2414);
and AND2 (N9693, N9686, N2315);
nor NOR3 (N9694, N9690, N7634, N6707);
or OR3 (N9695, N9694, N2773, N7721);
or OR2 (N9696, N9687, N28);
nand NAND3 (N9697, N9693, N5429, N5944);
nor NOR4 (N9698, N9697, N9597, N5435, N3077);
nand NAND2 (N9699, N9683, N2116);
xor XOR2 (N9700, N9695, N1849);
nand NAND3 (N9701, N9700, N4514, N9040);
nand NAND2 (N9702, N9681, N3575);
or OR3 (N9703, N9685, N2398, N4432);
and AND2 (N9704, N9684, N7141);
not NOT1 (N9705, N9701);
not NOT1 (N9706, N9689);
nand NAND2 (N9707, N9705, N3959);
nor NOR4 (N9708, N9696, N2406, N2864, N319);
xor XOR2 (N9709, N9699, N2795);
nand NAND4 (N9710, N9709, N2656, N5172, N5397);
and AND2 (N9711, N9708, N4721);
nor NOR2 (N9712, N9707, N6675);
or OR4 (N9713, N9691, N3400, N1709, N7205);
nor NOR4 (N9714, N9698, N1753, N993, N6141);
nor NOR2 (N9715, N9704, N6413);
nor NOR2 (N9716, N9692, N4159);
and AND2 (N9717, N9711, N7944);
or OR4 (N9718, N9706, N9326, N6206, N3315);
not NOT1 (N9719, N9716);
nor NOR4 (N9720, N9710, N9354, N2581, N484);
not NOT1 (N9721, N9715);
nor NOR3 (N9722, N9719, N7339, N2831);
xor XOR2 (N9723, N9703, N9210);
nand NAND2 (N9724, N9721, N4990);
buf BUF1 (N9725, N9724);
not NOT1 (N9726, N9717);
xor XOR2 (N9727, N9726, N7886);
or OR4 (N9728, N9722, N8678, N2252, N1253);
xor XOR2 (N9729, N9702, N2497);
nor NOR3 (N9730, N9727, N2188, N3372);
nor NOR3 (N9731, N9720, N7620, N6600);
nand NAND2 (N9732, N9714, N8430);
not NOT1 (N9733, N9728);
or OR3 (N9734, N9731, N1328, N2381);
xor XOR2 (N9735, N9712, N7809);
not NOT1 (N9736, N9734);
buf BUF1 (N9737, N9733);
and AND2 (N9738, N9732, N1099);
not NOT1 (N9739, N9737);
buf BUF1 (N9740, N9725);
xor XOR2 (N9741, N9723, N3340);
and AND2 (N9742, N9739, N1206);
nand NAND3 (N9743, N9738, N3956, N2637);
not NOT1 (N9744, N9740);
nand NAND2 (N9745, N9730, N4978);
and AND2 (N9746, N9741, N2050);
nand NAND2 (N9747, N9735, N4599);
not NOT1 (N9748, N9747);
and AND4 (N9749, N9743, N5669, N3846, N4109);
and AND3 (N9750, N9745, N2985, N6474);
or OR4 (N9751, N9748, N1027, N2237, N4784);
xor XOR2 (N9752, N9718, N9305);
or OR4 (N9753, N9744, N1512, N243, N5889);
xor XOR2 (N9754, N9746, N1161);
and AND2 (N9755, N9752, N8841);
xor XOR2 (N9756, N9749, N9197);
nor NOR2 (N9757, N9753, N3764);
not NOT1 (N9758, N9755);
not NOT1 (N9759, N9713);
buf BUF1 (N9760, N9751);
nor NOR4 (N9761, N9736, N5557, N9141, N346);
buf BUF1 (N9762, N9742);
not NOT1 (N9763, N9757);
nand NAND4 (N9764, N9756, N1271, N8575, N2044);
nand NAND2 (N9765, N9729, N5246);
and AND2 (N9766, N9761, N1057);
and AND3 (N9767, N9754, N2102, N7682);
or OR4 (N9768, N9760, N2982, N723, N4785);
nor NOR3 (N9769, N9759, N5863, N4047);
xor XOR2 (N9770, N9768, N5855);
xor XOR2 (N9771, N9750, N8452);
buf BUF1 (N9772, N9765);
or OR3 (N9773, N9772, N4788, N7726);
buf BUF1 (N9774, N9767);
or OR4 (N9775, N9766, N8560, N365, N205);
and AND4 (N9776, N9774, N3862, N5735, N6686);
xor XOR2 (N9777, N9776, N1157);
not NOT1 (N9778, N9762);
not NOT1 (N9779, N9758);
xor XOR2 (N9780, N9764, N3491);
buf BUF1 (N9781, N9773);
nand NAND4 (N9782, N9781, N2665, N3891, N298);
and AND4 (N9783, N9782, N8911, N5176, N3943);
nor NOR2 (N9784, N9769, N7902);
xor XOR2 (N9785, N9771, N7779);
or OR3 (N9786, N9775, N4081, N7864);
nand NAND2 (N9787, N9770, N699);
and AND2 (N9788, N9783, N6446);
nand NAND2 (N9789, N9784, N9124);
nand NAND3 (N9790, N9763, N88, N4681);
xor XOR2 (N9791, N9786, N486);
and AND3 (N9792, N9779, N9206, N8505);
not NOT1 (N9793, N9780);
and AND4 (N9794, N9788, N9037, N7282, N2433);
not NOT1 (N9795, N9794);
xor XOR2 (N9796, N9777, N21);
or OR3 (N9797, N9785, N6008, N2104);
not NOT1 (N9798, N9796);
nor NOR3 (N9799, N9795, N8676, N2094);
and AND4 (N9800, N9798, N1755, N8836, N5414);
buf BUF1 (N9801, N9789);
nand NAND2 (N9802, N9800, N339);
not NOT1 (N9803, N9801);
buf BUF1 (N9804, N9792);
or OR3 (N9805, N9804, N2745, N5810);
nand NAND2 (N9806, N9803, N1512);
or OR2 (N9807, N9793, N2230);
and AND4 (N9808, N9797, N5905, N9450, N1413);
and AND4 (N9809, N9808, N8473, N3291, N3189);
buf BUF1 (N9810, N9805);
not NOT1 (N9811, N9809);
nand NAND2 (N9812, N9791, N5293);
nor NOR2 (N9813, N9811, N2040);
nor NOR4 (N9814, N9807, N5047, N6523, N9767);
and AND2 (N9815, N9802, N6648);
buf BUF1 (N9816, N9810);
xor XOR2 (N9817, N9790, N7166);
not NOT1 (N9818, N9812);
nor NOR4 (N9819, N9817, N9098, N5297, N2188);
buf BUF1 (N9820, N9816);
and AND3 (N9821, N9819, N2773, N4923);
and AND3 (N9822, N9821, N7258, N8887);
nand NAND2 (N9823, N9787, N5589);
and AND4 (N9824, N9814, N9788, N2631, N1032);
xor XOR2 (N9825, N9818, N9397);
nand NAND3 (N9826, N9824, N9609, N3118);
or OR3 (N9827, N9778, N9775, N2518);
nor NOR4 (N9828, N9815, N8255, N3289, N8163);
buf BUF1 (N9829, N9828);
nor NOR4 (N9830, N9799, N1747, N9714, N3093);
and AND3 (N9831, N9806, N8427, N8957);
nand NAND4 (N9832, N9831, N2963, N3895, N4520);
not NOT1 (N9833, N9827);
nand NAND4 (N9834, N9826, N5977, N4447, N368);
buf BUF1 (N9835, N9834);
nor NOR2 (N9836, N9823, N7772);
and AND4 (N9837, N9832, N7709, N7599, N9800);
buf BUF1 (N9838, N9829);
not NOT1 (N9839, N9813);
nor NOR3 (N9840, N9822, N3740, N7739);
not NOT1 (N9841, N9830);
nand NAND3 (N9842, N9835, N4250, N6812);
nand NAND2 (N9843, N9820, N6695);
nor NOR2 (N9844, N9840, N5819);
or OR4 (N9845, N9836, N8478, N3099, N1705);
and AND4 (N9846, N9844, N7744, N2621, N2961);
nand NAND4 (N9847, N9837, N7986, N4544, N5175);
not NOT1 (N9848, N9825);
not NOT1 (N9849, N9848);
nor NOR3 (N9850, N9843, N2494, N4182);
buf BUF1 (N9851, N9849);
or OR2 (N9852, N9838, N534);
or OR3 (N9853, N9850, N2611, N8865);
xor XOR2 (N9854, N9851, N280);
nor NOR2 (N9855, N9846, N1552);
or OR4 (N9856, N9852, N1486, N3554, N6174);
buf BUF1 (N9857, N9853);
not NOT1 (N9858, N9854);
or OR4 (N9859, N9857, N9439, N1327, N8115);
and AND3 (N9860, N9855, N4705, N1771);
or OR4 (N9861, N9841, N7646, N1595, N6414);
buf BUF1 (N9862, N9860);
nor NOR2 (N9863, N9861, N575);
buf BUF1 (N9864, N9856);
nand NAND3 (N9865, N9842, N2821, N6000);
and AND4 (N9866, N9862, N130, N608, N8514);
and AND3 (N9867, N9839, N9403, N7812);
xor XOR2 (N9868, N9859, N8237);
xor XOR2 (N9869, N9867, N7637);
nor NOR2 (N9870, N9869, N3910);
xor XOR2 (N9871, N9865, N4439);
and AND4 (N9872, N9845, N2824, N6552, N966);
and AND2 (N9873, N9833, N9392);
or OR4 (N9874, N9866, N6458, N973, N7258);
xor XOR2 (N9875, N9874, N786);
nor NOR4 (N9876, N9847, N3509, N3384, N9119);
xor XOR2 (N9877, N9871, N9634);
nand NAND2 (N9878, N9875, N7652);
or OR4 (N9879, N9858, N2818, N9624, N695);
not NOT1 (N9880, N9878);
not NOT1 (N9881, N9863);
nand NAND4 (N9882, N9880, N9061, N3124, N7549);
nor NOR4 (N9883, N9870, N7569, N4100, N6055);
xor XOR2 (N9884, N9882, N166);
nor NOR3 (N9885, N9876, N3208, N993);
and AND2 (N9886, N9864, N7506);
xor XOR2 (N9887, N9881, N2960);
or OR4 (N9888, N9883, N6999, N1403, N2265);
nand NAND4 (N9889, N9877, N6349, N6367, N3730);
and AND3 (N9890, N9868, N4776, N7522);
nand NAND4 (N9891, N9888, N7875, N4456, N5252);
and AND3 (N9892, N9891, N2013, N1243);
and AND3 (N9893, N9890, N5193, N6883);
nand NAND3 (N9894, N9887, N7964, N3062);
and AND2 (N9895, N9873, N3141);
buf BUF1 (N9896, N9889);
not NOT1 (N9897, N9885);
nor NOR2 (N9898, N9872, N2508);
buf BUF1 (N9899, N9884);
not NOT1 (N9900, N9899);
or OR3 (N9901, N9895, N5373, N7421);
nand NAND2 (N9902, N9898, N7194);
xor XOR2 (N9903, N9901, N4456);
buf BUF1 (N9904, N9903);
or OR3 (N9905, N9896, N1168, N349);
nor NOR4 (N9906, N9879, N3568, N6773, N1385);
or OR3 (N9907, N9902, N5015, N8443);
not NOT1 (N9908, N9894);
and AND2 (N9909, N9905, N9621);
nor NOR2 (N9910, N9892, N6383);
nor NOR2 (N9911, N9907, N8371);
nand NAND4 (N9912, N9893, N9635, N5591, N781);
nand NAND3 (N9913, N9886, N8571, N3708);
xor XOR2 (N9914, N9900, N4958);
and AND2 (N9915, N9912, N1990);
nand NAND4 (N9916, N9906, N6427, N8943, N1450);
and AND2 (N9917, N9904, N2175);
and AND4 (N9918, N9913, N9786, N2355, N1027);
not NOT1 (N9919, N9916);
and AND3 (N9920, N9897, N5163, N6867);
nand NAND2 (N9921, N9910, N4903);
or OR4 (N9922, N9914, N130, N1730, N6620);
nor NOR4 (N9923, N9909, N9306, N6786, N8559);
nor NOR2 (N9924, N9915, N9501);
not NOT1 (N9925, N9920);
nor NOR2 (N9926, N9911, N2658);
buf BUF1 (N9927, N9917);
nor NOR4 (N9928, N9922, N7723, N9798, N990);
or OR2 (N9929, N9924, N6579);
or OR2 (N9930, N9927, N8123);
xor XOR2 (N9931, N9918, N2478);
nand NAND2 (N9932, N9908, N9910);
buf BUF1 (N9933, N9928);
and AND3 (N9934, N9932, N7602, N9480);
buf BUF1 (N9935, N9919);
buf BUF1 (N9936, N9925);
nor NOR3 (N9937, N9923, N8839, N2698);
xor XOR2 (N9938, N9935, N7652);
or OR4 (N9939, N9936, N6509, N175, N4155);
nand NAND4 (N9940, N9930, N2260, N8916, N7735);
nand NAND3 (N9941, N9938, N290, N4207);
not NOT1 (N9942, N9933);
buf BUF1 (N9943, N9940);
nor NOR2 (N9944, N9931, N4521);
or OR3 (N9945, N9943, N4210, N8443);
or OR2 (N9946, N9942, N6079);
and AND4 (N9947, N9941, N3028, N5930, N3193);
nor NOR3 (N9948, N9921, N3858, N2676);
xor XOR2 (N9949, N9946, N9250);
nand NAND2 (N9950, N9947, N7438);
xor XOR2 (N9951, N9948, N4300);
nor NOR4 (N9952, N9939, N5043, N8630, N7417);
nor NOR3 (N9953, N9937, N3077, N4074);
and AND4 (N9954, N9953, N2499, N1245, N1043);
nand NAND2 (N9955, N9926, N2320);
nand NAND2 (N9956, N9945, N9777);
nor NOR2 (N9957, N9955, N9955);
nor NOR2 (N9958, N9954, N4589);
xor XOR2 (N9959, N9958, N5731);
nor NOR4 (N9960, N9951, N5962, N4386, N4512);
or OR4 (N9961, N9934, N5221, N8899, N1750);
xor XOR2 (N9962, N9956, N6057);
not NOT1 (N9963, N9961);
xor XOR2 (N9964, N9949, N6115);
buf BUF1 (N9965, N9964);
nor NOR4 (N9966, N9962, N9436, N9890, N6116);
nor NOR3 (N9967, N9960, N3395, N2022);
and AND3 (N9968, N9967, N8492, N4380);
xor XOR2 (N9969, N9929, N4323);
not NOT1 (N9970, N9944);
buf BUF1 (N9971, N9963);
nor NOR2 (N9972, N9965, N1017);
not NOT1 (N9973, N9952);
nand NAND2 (N9974, N9950, N8159);
buf BUF1 (N9975, N9970);
buf BUF1 (N9976, N9959);
not NOT1 (N9977, N9972);
and AND2 (N9978, N9969, N2314);
nor NOR4 (N9979, N9957, N3673, N3388, N2623);
nand NAND3 (N9980, N9968, N3000, N186);
not NOT1 (N9981, N9966);
nor NOR2 (N9982, N9981, N9776);
not NOT1 (N9983, N9974);
not NOT1 (N9984, N9977);
and AND2 (N9985, N9973, N5263);
or OR4 (N9986, N9980, N44, N8930, N3496);
not NOT1 (N9987, N9978);
nand NAND3 (N9988, N9985, N6944, N2159);
nor NOR3 (N9989, N9988, N9538, N9320);
xor XOR2 (N9990, N9983, N1504);
nor NOR4 (N9991, N9976, N6546, N6839, N2521);
or OR4 (N9992, N9989, N469, N9055, N5567);
not NOT1 (N9993, N9971);
not NOT1 (N9994, N9992);
nand NAND4 (N9995, N9991, N6508, N3673, N1299);
nor NOR4 (N9996, N9993, N1435, N4551, N3016);
buf BUF1 (N9997, N9987);
or OR4 (N9998, N9984, N1083, N1408, N9888);
xor XOR2 (N9999, N9975, N9681);
buf BUF1 (N10000, N9994);
not NOT1 (N10001, N9986);
and AND3 (N10002, N9982, N6777, N7388);
nand NAND3 (N10003, N10002, N2375, N5153);
buf BUF1 (N10004, N10003);
not NOT1 (N10005, N9990);
nor NOR4 (N10006, N10005, N3565, N667, N6230);
not NOT1 (N10007, N9979);
and AND4 (N10008, N9999, N2328, N5599, N1741);
nand NAND4 (N10009, N10004, N4665, N6421, N9235);
buf BUF1 (N10010, N9998);
or OR2 (N10011, N10007, N1414);
nand NAND4 (N10012, N10009, N3487, N3012, N526);
nand NAND2 (N10013, N10010, N9092);
nand NAND4 (N10014, N10006, N6383, N3373, N645);
and AND3 (N10015, N10014, N6146, N928);
or OR3 (N10016, N9996, N8945, N3612);
nand NAND2 (N10017, N10015, N7638);
not NOT1 (N10018, N10017);
buf BUF1 (N10019, N10016);
not NOT1 (N10020, N10000);
nand NAND4 (N10021, N10008, N7990, N9594, N5854);
xor XOR2 (N10022, N9995, N3333);
xor XOR2 (N10023, N10019, N515);
nand NAND3 (N10024, N10023, N1841, N1477);
and AND3 (N10025, N9997, N7023, N7658);
nand NAND4 (N10026, N10012, N7790, N2543, N9333);
and AND4 (N10027, N10025, N1562, N7826, N6218);
and AND4 (N10028, N10022, N4848, N3749, N428);
xor XOR2 (N10029, N10027, N4573);
or OR4 (N10030, N10029, N576, N4756, N4254);
not NOT1 (N10031, N10028);
and AND2 (N10032, N10001, N5253);
not NOT1 (N10033, N10011);
not NOT1 (N10034, N10024);
and AND3 (N10035, N10020, N2810, N4752);
nor NOR2 (N10036, N10018, N2366);
nor NOR2 (N10037, N10035, N2202);
and AND4 (N10038, N10037, N8155, N639, N3112);
not NOT1 (N10039, N10033);
buf BUF1 (N10040, N10021);
xor XOR2 (N10041, N10036, N7538);
xor XOR2 (N10042, N10039, N1629);
xor XOR2 (N10043, N10038, N4159);
and AND3 (N10044, N10032, N3835, N1843);
nand NAND2 (N10045, N10040, N5196);
nor NOR3 (N10046, N10044, N6607, N4026);
or OR4 (N10047, N10026, N1716, N6057, N6111);
and AND4 (N10048, N10030, N4586, N9403, N3937);
xor XOR2 (N10049, N10013, N630);
nor NOR4 (N10050, N10049, N584, N5051, N4161);
buf BUF1 (N10051, N10043);
nor NOR3 (N10052, N10042, N9710, N4267);
buf BUF1 (N10053, N10048);
and AND2 (N10054, N10046, N4979);
buf BUF1 (N10055, N10031);
xor XOR2 (N10056, N10047, N7507);
nor NOR2 (N10057, N10053, N5407);
nor NOR2 (N10058, N10050, N8230);
buf BUF1 (N10059, N10058);
nand NAND4 (N10060, N10041, N5435, N2860, N5816);
xor XOR2 (N10061, N10051, N3029);
and AND4 (N10062, N10056, N8923, N9035, N9406);
xor XOR2 (N10063, N10052, N3027);
xor XOR2 (N10064, N10061, N2949);
or OR4 (N10065, N10062, N1524, N3298, N8222);
buf BUF1 (N10066, N10060);
and AND3 (N10067, N10034, N9985, N2255);
and AND2 (N10068, N10057, N12);
not NOT1 (N10069, N10045);
not NOT1 (N10070, N10065);
not NOT1 (N10071, N10069);
xor XOR2 (N10072, N10054, N5321);
nor NOR4 (N10073, N10068, N4768, N7032, N9739);
and AND4 (N10074, N10055, N7119, N9763, N5709);
buf BUF1 (N10075, N10073);
not NOT1 (N10076, N10064);
nand NAND4 (N10077, N10059, N9733, N5299, N6779);
or OR2 (N10078, N10070, N1682);
or OR4 (N10079, N10071, N7771, N6559, N5828);
nand NAND2 (N10080, N10077, N6336);
not NOT1 (N10081, N10072);
buf BUF1 (N10082, N10081);
buf BUF1 (N10083, N10066);
nor NOR4 (N10084, N10080, N8224, N7044, N1058);
or OR4 (N10085, N10076, N9696, N5160, N7724);
not NOT1 (N10086, N10063);
not NOT1 (N10087, N10075);
not NOT1 (N10088, N10085);
nor NOR3 (N10089, N10088, N2360, N7173);
xor XOR2 (N10090, N10089, N9608);
nand NAND4 (N10091, N10067, N8487, N174, N4523);
and AND3 (N10092, N10079, N9521, N10078);
and AND2 (N10093, N8822, N4634);
nand NAND3 (N10094, N10084, N4970, N9893);
not NOT1 (N10095, N10093);
buf BUF1 (N10096, N10086);
buf BUF1 (N10097, N10091);
not NOT1 (N10098, N10092);
buf BUF1 (N10099, N10097);
xor XOR2 (N10100, N10096, N650);
not NOT1 (N10101, N10095);
and AND4 (N10102, N10099, N7672, N71, N9253);
not NOT1 (N10103, N10087);
nand NAND3 (N10104, N10083, N5828, N573);
nor NOR4 (N10105, N10094, N5056, N5730, N6387);
nor NOR3 (N10106, N10082, N9757, N1081);
xor XOR2 (N10107, N10103, N4112);
nor NOR4 (N10108, N10100, N9369, N4248, N374);
or OR3 (N10109, N10106, N7224, N3678);
not NOT1 (N10110, N10090);
nor NOR4 (N10111, N10101, N4416, N7443, N8845);
buf BUF1 (N10112, N10102);
or OR2 (N10113, N10105, N914);
and AND4 (N10114, N10111, N4211, N1394, N9022);
and AND4 (N10115, N10109, N4941, N6156, N7462);
nand NAND3 (N10116, N10108, N489, N9537);
buf BUF1 (N10117, N10115);
not NOT1 (N10118, N10074);
xor XOR2 (N10119, N10118, N9211);
nand NAND4 (N10120, N10104, N3670, N8610, N8346);
or OR3 (N10121, N10116, N5987, N5574);
or OR4 (N10122, N10120, N6032, N2063, N7956);
nand NAND3 (N10123, N10114, N3832, N805);
or OR2 (N10124, N10098, N3022);
or OR2 (N10125, N10113, N3849);
and AND2 (N10126, N10107, N3776);
not NOT1 (N10127, N10110);
buf BUF1 (N10128, N10125);
nand NAND2 (N10129, N10124, N5446);
or OR3 (N10130, N10117, N7066, N8432);
buf BUF1 (N10131, N10128);
xor XOR2 (N10132, N10121, N2198);
not NOT1 (N10133, N10130);
or OR3 (N10134, N10133, N59, N9824);
and AND2 (N10135, N10126, N2988);
nor NOR2 (N10136, N10119, N6474);
nor NOR2 (N10137, N10135, N2566);
not NOT1 (N10138, N10127);
not NOT1 (N10139, N10122);
nor NOR3 (N10140, N10132, N3667, N3708);
or OR3 (N10141, N10112, N8998, N9384);
buf BUF1 (N10142, N10123);
nor NOR2 (N10143, N10131, N1355);
buf BUF1 (N10144, N10134);
nand NAND4 (N10145, N10136, N4251, N4733, N6810);
xor XOR2 (N10146, N10141, N81);
nor NOR2 (N10147, N10145, N8684);
or OR2 (N10148, N10144, N8224);
and AND2 (N10149, N10129, N2092);
buf BUF1 (N10150, N10138);
xor XOR2 (N10151, N10149, N208);
and AND2 (N10152, N10139, N1278);
not NOT1 (N10153, N10148);
nand NAND2 (N10154, N10150, N6162);
or OR2 (N10155, N10147, N9439);
xor XOR2 (N10156, N10142, N6640);
buf BUF1 (N10157, N10151);
xor XOR2 (N10158, N10140, N8065);
nor NOR2 (N10159, N10137, N2124);
and AND3 (N10160, N10153, N2717, N5175);
not NOT1 (N10161, N10146);
buf BUF1 (N10162, N10155);
or OR3 (N10163, N10143, N12, N5300);
nor NOR3 (N10164, N10163, N7933, N9798);
not NOT1 (N10165, N10159);
not NOT1 (N10166, N10165);
nor NOR3 (N10167, N10166, N355, N7227);
xor XOR2 (N10168, N10167, N8576);
or OR2 (N10169, N10168, N9876);
and AND4 (N10170, N10156, N3768, N7720, N9648);
not NOT1 (N10171, N10157);
nor NOR2 (N10172, N10170, N10073);
and AND3 (N10173, N10158, N6809, N313);
or OR4 (N10174, N10173, N5517, N1689, N9563);
or OR3 (N10175, N10161, N2720, N459);
not NOT1 (N10176, N10160);
nand NAND2 (N10177, N10175, N4961);
or OR3 (N10178, N10154, N6065, N2954);
and AND4 (N10179, N10177, N1343, N7220, N4103);
xor XOR2 (N10180, N10162, N10164);
buf BUF1 (N10181, N2028);
nor NOR2 (N10182, N10176, N1495);
nand NAND3 (N10183, N10152, N1211, N5582);
buf BUF1 (N10184, N10180);
buf BUF1 (N10185, N10183);
buf BUF1 (N10186, N10172);
xor XOR2 (N10187, N10178, N6548);
and AND3 (N10188, N10187, N2040, N4456);
or OR4 (N10189, N10188, N3277, N8400, N4977);
or OR4 (N10190, N10184, N8398, N2064, N8652);
or OR2 (N10191, N10189, N8454);
not NOT1 (N10192, N10181);
or OR4 (N10193, N10182, N6884, N4111, N7809);
buf BUF1 (N10194, N10186);
nand NAND3 (N10195, N10192, N7122, N69);
nor NOR3 (N10196, N10190, N1868, N1909);
nor NOR3 (N10197, N10196, N2300, N661);
nand NAND2 (N10198, N10169, N2517);
or OR4 (N10199, N10194, N3527, N371, N9778);
nor NOR3 (N10200, N10191, N3310, N1062);
and AND2 (N10201, N10193, N1069);
nand NAND4 (N10202, N10197, N3230, N9086, N7138);
nand NAND3 (N10203, N10199, N7009, N326);
not NOT1 (N10204, N10179);
buf BUF1 (N10205, N10202);
not NOT1 (N10206, N10198);
nor NOR4 (N10207, N10203, N6014, N1421, N5738);
buf BUF1 (N10208, N10185);
buf BUF1 (N10209, N10195);
not NOT1 (N10210, N10209);
not NOT1 (N10211, N10207);
xor XOR2 (N10212, N10174, N1347);
or OR4 (N10213, N10211, N7333, N8686, N685);
buf BUF1 (N10214, N10200);
nor NOR4 (N10215, N10212, N10059, N4427, N10056);
xor XOR2 (N10216, N10208, N3639);
not NOT1 (N10217, N10201);
nand NAND4 (N10218, N10217, N699, N5702, N6173);
nor NOR4 (N10219, N10204, N6019, N864, N8901);
and AND2 (N10220, N10210, N7093);
xor XOR2 (N10221, N10205, N9797);
nand NAND2 (N10222, N10221, N8905);
or OR3 (N10223, N10214, N3960, N468);
not NOT1 (N10224, N10215);
nor NOR3 (N10225, N10206, N5098, N10048);
and AND2 (N10226, N10213, N732);
xor XOR2 (N10227, N10226, N5371);
and AND4 (N10228, N10220, N5736, N1553, N7607);
not NOT1 (N10229, N10171);
buf BUF1 (N10230, N10225);
xor XOR2 (N10231, N10227, N2025);
nor NOR3 (N10232, N10229, N3628, N7523);
not NOT1 (N10233, N10218);
not NOT1 (N10234, N10216);
buf BUF1 (N10235, N10231);
or OR3 (N10236, N10222, N4110, N609);
nor NOR4 (N10237, N10234, N4687, N6425, N9854);
nor NOR3 (N10238, N10228, N232, N3671);
xor XOR2 (N10239, N10223, N4851);
nor NOR2 (N10240, N10237, N7428);
nor NOR4 (N10241, N10236, N8999, N5374, N8161);
or OR2 (N10242, N10239, N2168);
buf BUF1 (N10243, N10242);
xor XOR2 (N10244, N10232, N6112);
nand NAND3 (N10245, N10230, N744, N7457);
xor XOR2 (N10246, N10219, N5103);
not NOT1 (N10247, N10238);
and AND3 (N10248, N10224, N2304, N7249);
xor XOR2 (N10249, N10247, N1337);
and AND2 (N10250, N10249, N1438);
xor XOR2 (N10251, N10233, N6374);
buf BUF1 (N10252, N10246);
nor NOR2 (N10253, N10244, N9626);
xor XOR2 (N10254, N10243, N7686);
xor XOR2 (N10255, N10253, N7243);
xor XOR2 (N10256, N10235, N9335);
nor NOR2 (N10257, N10255, N4483);
not NOT1 (N10258, N10252);
nor NOR3 (N10259, N10240, N9349, N516);
xor XOR2 (N10260, N10248, N4698);
buf BUF1 (N10261, N10245);
or OR2 (N10262, N10261, N3612);
not NOT1 (N10263, N10241);
xor XOR2 (N10264, N10257, N5921);
nand NAND4 (N10265, N10254, N344, N3481, N10263);
nor NOR3 (N10266, N9632, N7823, N5629);
nor NOR3 (N10267, N10264, N5247, N10171);
nor NOR4 (N10268, N10262, N5931, N4184, N10002);
nand NAND2 (N10269, N10260, N6065);
and AND3 (N10270, N10256, N9934, N4014);
and AND2 (N10271, N10267, N4987);
not NOT1 (N10272, N10250);
and AND4 (N10273, N10271, N7817, N8207, N4686);
nor NOR3 (N10274, N10270, N8325, N8385);
buf BUF1 (N10275, N10259);
not NOT1 (N10276, N10265);
nand NAND3 (N10277, N10266, N4838, N6763);
nand NAND4 (N10278, N10275, N5896, N4477, N1248);
or OR4 (N10279, N10276, N3334, N8257, N1981);
nand NAND4 (N10280, N10278, N6980, N21, N8321);
or OR2 (N10281, N10251, N9782);
xor XOR2 (N10282, N10258, N701);
nor NOR3 (N10283, N10268, N2880, N366);
xor XOR2 (N10284, N10280, N5547);
or OR3 (N10285, N10277, N2494, N3859);
or OR4 (N10286, N10272, N6269, N7404, N6530);
or OR3 (N10287, N10279, N4447, N3140);
buf BUF1 (N10288, N10287);
and AND3 (N10289, N10274, N9300, N4765);
or OR3 (N10290, N10284, N4922, N1583);
xor XOR2 (N10291, N10286, N3019);
and AND3 (N10292, N10291, N9823, N1743);
buf BUF1 (N10293, N10288);
nand NAND4 (N10294, N10281, N2809, N1322, N1429);
and AND4 (N10295, N10273, N5355, N2820, N6199);
not NOT1 (N10296, N10295);
nor NOR2 (N10297, N10294, N9716);
or OR4 (N10298, N10285, N8581, N474, N4797);
buf BUF1 (N10299, N10269);
nand NAND4 (N10300, N10297, N1599, N6067, N6008);
and AND4 (N10301, N10282, N10166, N718, N1734);
and AND4 (N10302, N10300, N8760, N9089, N4777);
or OR2 (N10303, N10296, N2840);
not NOT1 (N10304, N10292);
buf BUF1 (N10305, N10298);
not NOT1 (N10306, N10304);
not NOT1 (N10307, N10303);
or OR4 (N10308, N10289, N6141, N796, N1742);
not NOT1 (N10309, N10283);
nand NAND4 (N10310, N10293, N4437, N680, N21);
nor NOR3 (N10311, N10306, N1810, N9263);
or OR3 (N10312, N10302, N9245, N10204);
not NOT1 (N10313, N10305);
buf BUF1 (N10314, N10309);
nand NAND3 (N10315, N10314, N3598, N8272);
or OR4 (N10316, N10315, N9303, N5940, N3334);
buf BUF1 (N10317, N10313);
not NOT1 (N10318, N10311);
nand NAND2 (N10319, N10307, N5020);
nor NOR3 (N10320, N10308, N6674, N4380);
nand NAND2 (N10321, N10301, N4732);
and AND3 (N10322, N10318, N8991, N36);
nor NOR3 (N10323, N10319, N9342, N1010);
nand NAND4 (N10324, N10321, N2519, N829, N3347);
nor NOR4 (N10325, N10324, N8720, N8581, N588);
not NOT1 (N10326, N10299);
and AND3 (N10327, N10323, N862, N2935);
nand NAND4 (N10328, N10326, N4191, N6651, N7741);
nand NAND2 (N10329, N10320, N1023);
or OR4 (N10330, N10329, N4363, N5169, N1335);
nand NAND4 (N10331, N10328, N596, N7265, N3206);
nor NOR2 (N10332, N10317, N1056);
nor NOR3 (N10333, N10312, N3690, N8492);
nand NAND4 (N10334, N10332, N7704, N6659, N1177);
nor NOR3 (N10335, N10290, N3461, N6732);
not NOT1 (N10336, N10316);
buf BUF1 (N10337, N10330);
nand NAND4 (N10338, N10336, N9570, N9913, N8464);
nor NOR2 (N10339, N10333, N4696);
buf BUF1 (N10340, N10322);
buf BUF1 (N10341, N10325);
xor XOR2 (N10342, N10337, N7263);
xor XOR2 (N10343, N10335, N4960);
xor XOR2 (N10344, N10338, N7865);
or OR3 (N10345, N10327, N9573, N1439);
and AND4 (N10346, N10334, N6219, N2733, N4079);
buf BUF1 (N10347, N10344);
not NOT1 (N10348, N10310);
nor NOR2 (N10349, N10346, N3311);
or OR4 (N10350, N10349, N6408, N1582, N417);
nand NAND2 (N10351, N10342, N7727);
or OR4 (N10352, N10348, N6993, N9648, N7593);
and AND4 (N10353, N10341, N5532, N6574, N6940);
buf BUF1 (N10354, N10339);
nand NAND2 (N10355, N10350, N4848);
xor XOR2 (N10356, N10343, N1981);
not NOT1 (N10357, N10355);
and AND3 (N10358, N10357, N4716, N1281);
nand NAND3 (N10359, N10354, N4903, N9045);
buf BUF1 (N10360, N10353);
xor XOR2 (N10361, N10356, N6765);
nor NOR2 (N10362, N10331, N792);
buf BUF1 (N10363, N10361);
nand NAND2 (N10364, N10352, N7289);
not NOT1 (N10365, N10358);
or OR3 (N10366, N10360, N7504, N5036);
or OR3 (N10367, N10364, N2977, N4333);
or OR3 (N10368, N10359, N9702, N1512);
and AND3 (N10369, N10366, N10083, N3669);
nand NAND2 (N10370, N10347, N3003);
nand NAND2 (N10371, N10370, N5610);
nor NOR2 (N10372, N10340, N1608);
buf BUF1 (N10373, N10351);
not NOT1 (N10374, N10367);
and AND4 (N10375, N10372, N3275, N3536, N9782);
nand NAND3 (N10376, N10345, N8698, N2562);
nand NAND3 (N10377, N10376, N5422, N5);
buf BUF1 (N10378, N10375);
buf BUF1 (N10379, N10377);
not NOT1 (N10380, N10371);
nand NAND2 (N10381, N10362, N79);
nor NOR3 (N10382, N10363, N2884, N6577);
not NOT1 (N10383, N10365);
xor XOR2 (N10384, N10382, N9435);
xor XOR2 (N10385, N10369, N9611);
and AND3 (N10386, N10385, N1213, N8360);
nand NAND2 (N10387, N10373, N9873);
not NOT1 (N10388, N10379);
or OR4 (N10389, N10384, N1143, N10121, N1257);
buf BUF1 (N10390, N10380);
nand NAND2 (N10391, N10390, N3881);
or OR4 (N10392, N10374, N6370, N593, N8382);
not NOT1 (N10393, N10391);
buf BUF1 (N10394, N10378);
xor XOR2 (N10395, N10381, N9638);
not NOT1 (N10396, N10368);
xor XOR2 (N10397, N10383, N5377);
and AND3 (N10398, N10387, N7517, N9132);
nand NAND3 (N10399, N10389, N704, N6093);
xor XOR2 (N10400, N10399, N1513);
or OR2 (N10401, N10398, N9891);
not NOT1 (N10402, N10388);
nand NAND3 (N10403, N10396, N3204, N3);
nand NAND4 (N10404, N10386, N6514, N7443, N1541);
xor XOR2 (N10405, N10402, N7934);
nor NOR4 (N10406, N10392, N146, N3589, N7085);
xor XOR2 (N10407, N10403, N2054);
nand NAND3 (N10408, N10405, N8572, N6093);
buf BUF1 (N10409, N10393);
nand NAND3 (N10410, N10394, N3504, N796);
nand NAND3 (N10411, N10409, N3444, N8262);
xor XOR2 (N10412, N10395, N5532);
nor NOR4 (N10413, N10410, N5097, N9775, N6969);
not NOT1 (N10414, N10407);
nor NOR4 (N10415, N10400, N4330, N6639, N2468);
nand NAND3 (N10416, N10411, N4275, N5100);
nor NOR2 (N10417, N10415, N9163);
not NOT1 (N10418, N10401);
nand NAND4 (N10419, N10417, N2943, N2147, N9938);
nor NOR2 (N10420, N10414, N1436);
nor NOR2 (N10421, N10412, N1189);
not NOT1 (N10422, N10406);
and AND3 (N10423, N10413, N3386, N3546);
nor NOR4 (N10424, N10421, N4033, N1242, N4538);
and AND4 (N10425, N10424, N2452, N3833, N5914);
xor XOR2 (N10426, N10425, N5834);
and AND3 (N10427, N10423, N8439, N10102);
nor NOR4 (N10428, N10404, N10274, N8245, N5081);
nor NOR2 (N10429, N10397, N1282);
nand NAND2 (N10430, N10416, N4140);
nand NAND3 (N10431, N10426, N1822, N311);
nor NOR4 (N10432, N10428, N3149, N2806, N2795);
and AND4 (N10433, N10427, N7124, N5040, N2645);
xor XOR2 (N10434, N10431, N6771);
nor NOR4 (N10435, N10418, N4334, N5945, N8081);
xor XOR2 (N10436, N10434, N5132);
and AND3 (N10437, N10408, N5689, N1461);
buf BUF1 (N10438, N10429);
xor XOR2 (N10439, N10437, N4439);
nor NOR2 (N10440, N10422, N6539);
not NOT1 (N10441, N10419);
not NOT1 (N10442, N10435);
nor NOR4 (N10443, N10420, N8540, N7674, N9750);
and AND3 (N10444, N10436, N2634, N8307);
xor XOR2 (N10445, N10430, N4863);
nor NOR2 (N10446, N10444, N4539);
nand NAND4 (N10447, N10442, N10056, N2798, N2305);
or OR3 (N10448, N10443, N3430, N2094);
or OR2 (N10449, N10433, N8823);
and AND4 (N10450, N10440, N3397, N2384, N6432);
or OR2 (N10451, N10448, N9275);
buf BUF1 (N10452, N10438);
nand NAND4 (N10453, N10447, N7458, N3255, N5787);
buf BUF1 (N10454, N10432);
not NOT1 (N10455, N10451);
buf BUF1 (N10456, N10454);
or OR4 (N10457, N10450, N3644, N852, N10445);
xor XOR2 (N10458, N7438, N8062);
nand NAND4 (N10459, N10455, N9862, N4781, N10365);
buf BUF1 (N10460, N10441);
and AND2 (N10461, N10453, N9984);
buf BUF1 (N10462, N10460);
nor NOR2 (N10463, N10458, N7760);
buf BUF1 (N10464, N10452);
not NOT1 (N10465, N10439);
nor NOR3 (N10466, N10462, N6837, N9888);
nand NAND2 (N10467, N10457, N379);
nor NOR4 (N10468, N10467, N853, N3722, N1576);
not NOT1 (N10469, N10456);
nor NOR2 (N10470, N10459, N7398);
xor XOR2 (N10471, N10466, N929);
nand NAND4 (N10472, N10446, N3653, N9739, N3293);
buf BUF1 (N10473, N10461);
and AND3 (N10474, N10463, N8670, N2055);
nor NOR3 (N10475, N10472, N5627, N6600);
nor NOR3 (N10476, N10465, N4539, N859);
and AND3 (N10477, N10449, N4387, N2354);
nor NOR3 (N10478, N10473, N249, N3069);
nand NAND2 (N10479, N10477, N5832);
and AND2 (N10480, N10471, N7912);
buf BUF1 (N10481, N10469);
buf BUF1 (N10482, N10479);
xor XOR2 (N10483, N10470, N1331);
xor XOR2 (N10484, N10464, N8236);
nand NAND2 (N10485, N10481, N3646);
or OR4 (N10486, N10478, N6165, N9950, N7603);
xor XOR2 (N10487, N10468, N3843);
nand NAND2 (N10488, N10486, N7442);
nor NOR2 (N10489, N10480, N2409);
nand NAND4 (N10490, N10489, N3969, N4458, N2027);
not NOT1 (N10491, N10475);
buf BUF1 (N10492, N10488);
nor NOR3 (N10493, N10485, N8610, N5927);
xor XOR2 (N10494, N10491, N1891);
not NOT1 (N10495, N10493);
nor NOR2 (N10496, N10487, N4752);
or OR4 (N10497, N10482, N1436, N2113, N7033);
or OR3 (N10498, N10495, N6289, N1057);
nor NOR4 (N10499, N10494, N6163, N4898, N7552);
or OR4 (N10500, N10476, N10333, N9663, N6542);
nand NAND3 (N10501, N10492, N5505, N9279);
buf BUF1 (N10502, N10490);
nand NAND3 (N10503, N10501, N2371, N4378);
buf BUF1 (N10504, N10496);
xor XOR2 (N10505, N10484, N688);
not NOT1 (N10506, N10502);
nand NAND2 (N10507, N10474, N10030);
xor XOR2 (N10508, N10498, N3640);
buf BUF1 (N10509, N10483);
buf BUF1 (N10510, N10499);
not NOT1 (N10511, N10503);
xor XOR2 (N10512, N10507, N1827);
nor NOR3 (N10513, N10509, N1907, N1569);
nand NAND4 (N10514, N10510, N10023, N8204, N4767);
xor XOR2 (N10515, N10504, N6482);
nand NAND4 (N10516, N10508, N828, N9198, N4624);
not NOT1 (N10517, N10512);
or OR2 (N10518, N10513, N2574);
buf BUF1 (N10519, N10515);
nor NOR2 (N10520, N10516, N9095);
nand NAND3 (N10521, N10511, N3187, N6942);
nand NAND3 (N10522, N10521, N8550, N5380);
or OR2 (N10523, N10517, N8583);
nor NOR4 (N10524, N10518, N3439, N7834, N6136);
nor NOR4 (N10525, N10522, N911, N4554, N2014);
nor NOR2 (N10526, N10505, N3953);
nor NOR2 (N10527, N10526, N1494);
nor NOR3 (N10528, N10506, N7279, N5438);
nand NAND3 (N10529, N10497, N1340, N10206);
nor NOR4 (N10530, N10527, N5571, N4286, N5088);
nor NOR4 (N10531, N10519, N1729, N5289, N4729);
nand NAND2 (N10532, N10530, N6310);
nor NOR4 (N10533, N10531, N3727, N6931, N7445);
or OR2 (N10534, N10525, N3889);
nand NAND4 (N10535, N10514, N1129, N7436, N5479);
xor XOR2 (N10536, N10535, N7964);
not NOT1 (N10537, N10532);
buf BUF1 (N10538, N10534);
and AND3 (N10539, N10537, N2632, N3224);
or OR3 (N10540, N10529, N736, N640);
buf BUF1 (N10541, N10536);
not NOT1 (N10542, N10524);
nand NAND3 (N10543, N10539, N3330, N4937);
nand NAND3 (N10544, N10520, N297, N8384);
not NOT1 (N10545, N10533);
nor NOR2 (N10546, N10545, N2735);
not NOT1 (N10547, N10543);
xor XOR2 (N10548, N10542, N6984);
not NOT1 (N10549, N10548);
xor XOR2 (N10550, N10549, N4096);
nor NOR3 (N10551, N10523, N9438, N7633);
xor XOR2 (N10552, N10547, N8390);
nor NOR4 (N10553, N10546, N3548, N715, N9348);
or OR4 (N10554, N10544, N8265, N1555, N4309);
buf BUF1 (N10555, N10541);
nand NAND4 (N10556, N10500, N7757, N1434, N4575);
xor XOR2 (N10557, N10528, N3317);
xor XOR2 (N10558, N10553, N9365);
buf BUF1 (N10559, N10538);
nor NOR2 (N10560, N10551, N3660);
or OR2 (N10561, N10556, N3006);
not NOT1 (N10562, N10555);
not NOT1 (N10563, N10559);
nor NOR2 (N10564, N10563, N5414);
xor XOR2 (N10565, N10560, N2417);
buf BUF1 (N10566, N10565);
not NOT1 (N10567, N10566);
buf BUF1 (N10568, N10540);
not NOT1 (N10569, N10568);
and AND2 (N10570, N10567, N4322);
or OR3 (N10571, N10550, N2152, N9917);
buf BUF1 (N10572, N10570);
buf BUF1 (N10573, N10562);
buf BUF1 (N10574, N10572);
or OR2 (N10575, N10554, N9412);
buf BUF1 (N10576, N10571);
xor XOR2 (N10577, N10573, N5368);
and AND4 (N10578, N10575, N6232, N6258, N3787);
and AND2 (N10579, N10564, N4761);
and AND4 (N10580, N10557, N10541, N7500, N2265);
buf BUF1 (N10581, N10576);
and AND4 (N10582, N10574, N8834, N9748, N5051);
buf BUF1 (N10583, N10580);
xor XOR2 (N10584, N10561, N6327);
not NOT1 (N10585, N10583);
nor NOR3 (N10586, N10584, N4842, N10580);
not NOT1 (N10587, N10582);
nor NOR3 (N10588, N10577, N4574, N737);
or OR3 (N10589, N10588, N7508, N4345);
or OR2 (N10590, N10558, N2484);
not NOT1 (N10591, N10587);
not NOT1 (N10592, N10586);
not NOT1 (N10593, N10589);
buf BUF1 (N10594, N10579);
and AND4 (N10595, N10552, N1156, N1126, N6758);
xor XOR2 (N10596, N10590, N3425);
buf BUF1 (N10597, N10569);
nand NAND4 (N10598, N10597, N45, N8036, N5350);
not NOT1 (N10599, N10593);
xor XOR2 (N10600, N10592, N8363);
nand NAND4 (N10601, N10598, N5222, N7681, N3849);
xor XOR2 (N10602, N10581, N8303);
nor NOR4 (N10603, N10594, N3434, N5624, N8376);
nand NAND4 (N10604, N10603, N1216, N10441, N1443);
not NOT1 (N10605, N10604);
nand NAND4 (N10606, N10591, N2845, N8463, N1696);
and AND4 (N10607, N10599, N5483, N8632, N3041);
nor NOR2 (N10608, N10607, N5404);
not NOT1 (N10609, N10602);
nor NOR3 (N10610, N10609, N9176, N792);
xor XOR2 (N10611, N10596, N8236);
nand NAND3 (N10612, N10585, N2451, N7183);
not NOT1 (N10613, N10611);
or OR4 (N10614, N10608, N2502, N10540, N6807);
and AND2 (N10615, N10600, N9024);
and AND3 (N10616, N10610, N9725, N1801);
nor NOR3 (N10617, N10601, N3650, N812);
nand NAND2 (N10618, N10605, N5542);
and AND3 (N10619, N10606, N7075, N2225);
not NOT1 (N10620, N10618);
nand NAND2 (N10621, N10619, N4832);
nand NAND2 (N10622, N10621, N7805);
nand NAND3 (N10623, N10615, N2260, N558);
and AND4 (N10624, N10578, N619, N265, N10106);
nor NOR2 (N10625, N10624, N3893);
and AND3 (N10626, N10616, N7957, N9117);
or OR4 (N10627, N10626, N9539, N4712, N10440);
and AND4 (N10628, N10622, N149, N6693, N5883);
xor XOR2 (N10629, N10628, N1796);
xor XOR2 (N10630, N10629, N4586);
xor XOR2 (N10631, N10595, N5941);
not NOT1 (N10632, N10623);
or OR4 (N10633, N10612, N8054, N4621, N6206);
nand NAND4 (N10634, N10620, N7578, N3860, N8781);
xor XOR2 (N10635, N10613, N990);
and AND4 (N10636, N10627, N729, N5806, N7419);
xor XOR2 (N10637, N10614, N7869);
buf BUF1 (N10638, N10617);
not NOT1 (N10639, N10625);
and AND2 (N10640, N10636, N3792);
nand NAND2 (N10641, N10630, N372);
buf BUF1 (N10642, N10638);
and AND3 (N10643, N10641, N10123, N5549);
and AND3 (N10644, N10631, N6125, N974);
buf BUF1 (N10645, N10637);
not NOT1 (N10646, N10645);
not NOT1 (N10647, N10640);
or OR3 (N10648, N10644, N7760, N3332);
buf BUF1 (N10649, N10632);
buf BUF1 (N10650, N10648);
xor XOR2 (N10651, N10650, N7666);
buf BUF1 (N10652, N10633);
or OR4 (N10653, N10642, N7366, N3939, N9385);
nor NOR3 (N10654, N10646, N1192, N6718);
nor NOR2 (N10655, N10639, N4015);
xor XOR2 (N10656, N10649, N9109);
nand NAND2 (N10657, N10655, N3367);
buf BUF1 (N10658, N10647);
not NOT1 (N10659, N10643);
nor NOR2 (N10660, N10653, N8535);
or OR4 (N10661, N10654, N4911, N7253, N9438);
nand NAND4 (N10662, N10634, N920, N5556, N8597);
and AND3 (N10663, N10659, N9370, N2021);
or OR3 (N10664, N10651, N466, N6817);
xor XOR2 (N10665, N10660, N1504);
buf BUF1 (N10666, N10635);
and AND4 (N10667, N10652, N172, N10196, N6424);
not NOT1 (N10668, N10667);
buf BUF1 (N10669, N10665);
or OR2 (N10670, N10656, N8148);
buf BUF1 (N10671, N10669);
xor XOR2 (N10672, N10668, N2565);
nand NAND2 (N10673, N10663, N9423);
or OR2 (N10674, N10661, N10431);
nand NAND4 (N10675, N10662, N6824, N4138, N7673);
xor XOR2 (N10676, N10666, N10215);
nor NOR4 (N10677, N10676, N4479, N4495, N6417);
and AND4 (N10678, N10664, N9106, N2544, N7881);
xor XOR2 (N10679, N10677, N1075);
nor NOR2 (N10680, N10671, N2247);
xor XOR2 (N10681, N10678, N2346);
buf BUF1 (N10682, N10657);
nor NOR4 (N10683, N10673, N8440, N10425, N6987);
or OR2 (N10684, N10679, N10606);
or OR3 (N10685, N10681, N2654, N4655);
not NOT1 (N10686, N10674);
not NOT1 (N10687, N10686);
nor NOR2 (N10688, N10682, N4809);
xor XOR2 (N10689, N10672, N731);
not NOT1 (N10690, N10675);
nand NAND3 (N10691, N10688, N9913, N6072);
and AND4 (N10692, N10685, N2541, N1093, N6754);
xor XOR2 (N10693, N10687, N1013);
xor XOR2 (N10694, N10693, N4909);
or OR3 (N10695, N10680, N4678, N5893);
not NOT1 (N10696, N10683);
nand NAND3 (N10697, N10695, N5539, N4247);
nor NOR4 (N10698, N10658, N10285, N3247, N2372);
nor NOR3 (N10699, N10692, N7411, N2553);
and AND2 (N10700, N10684, N1484);
buf BUF1 (N10701, N10700);
buf BUF1 (N10702, N10694);
buf BUF1 (N10703, N10696);
nand NAND2 (N10704, N10703, N3754);
xor XOR2 (N10705, N10690, N6071);
or OR4 (N10706, N10705, N1018, N9506, N6532);
xor XOR2 (N10707, N10697, N9335);
nor NOR2 (N10708, N10702, N459);
not NOT1 (N10709, N10704);
or OR4 (N10710, N10701, N9839, N8760, N5547);
xor XOR2 (N10711, N10707, N2192);
buf BUF1 (N10712, N10698);
not NOT1 (N10713, N10689);
xor XOR2 (N10714, N10670, N445);
xor XOR2 (N10715, N10712, N8418);
nor NOR2 (N10716, N10715, N3495);
nand NAND2 (N10717, N10709, N8315);
xor XOR2 (N10718, N10717, N8392);
nor NOR3 (N10719, N10714, N3531, N8604);
xor XOR2 (N10720, N10699, N1130);
or OR4 (N10721, N10718, N9485, N4696, N2302);
or OR2 (N10722, N10706, N5862);
and AND2 (N10723, N10721, N10416);
nand NAND3 (N10724, N10722, N3092, N2545);
buf BUF1 (N10725, N10691);
nand NAND2 (N10726, N10711, N4566);
nand NAND4 (N10727, N10723, N1603, N3057, N1998);
nand NAND4 (N10728, N10713, N10077, N6306, N4276);
xor XOR2 (N10729, N10724, N5504);
buf BUF1 (N10730, N10708);
not NOT1 (N10731, N10726);
nand NAND3 (N10732, N10729, N955, N8893);
nor NOR4 (N10733, N10720, N5828, N1085, N10531);
or OR4 (N10734, N10716, N4294, N9230, N1088);
nand NAND2 (N10735, N10728, N9878);
not NOT1 (N10736, N10733);
xor XOR2 (N10737, N10730, N9572);
buf BUF1 (N10738, N10725);
buf BUF1 (N10739, N10737);
and AND4 (N10740, N10731, N1832, N530, N2261);
or OR2 (N10741, N10739, N7126);
nand NAND4 (N10742, N10738, N8956, N4141, N5196);
and AND2 (N10743, N10732, N7917);
and AND2 (N10744, N10740, N3720);
nand NAND3 (N10745, N10734, N9335, N2402);
xor XOR2 (N10746, N10727, N1455);
buf BUF1 (N10747, N10710);
nor NOR2 (N10748, N10743, N10483);
or OR2 (N10749, N10746, N8300);
buf BUF1 (N10750, N10741);
nor NOR2 (N10751, N10736, N4590);
buf BUF1 (N10752, N10719);
and AND3 (N10753, N10751, N804, N1968);
and AND2 (N10754, N10752, N5872);
or OR2 (N10755, N10753, N1360);
or OR3 (N10756, N10742, N8910, N9191);
nand NAND3 (N10757, N10735, N2274, N9066);
nor NOR3 (N10758, N10747, N6850, N6737);
xor XOR2 (N10759, N10755, N8421);
or OR2 (N10760, N10758, N6047);
xor XOR2 (N10761, N10749, N9115);
buf BUF1 (N10762, N10760);
buf BUF1 (N10763, N10744);
nor NOR2 (N10764, N10748, N8854);
nand NAND3 (N10765, N10764, N523, N1629);
nor NOR3 (N10766, N10757, N10589, N9047);
nor NOR3 (N10767, N10766, N10310, N8971);
nor NOR2 (N10768, N10759, N10355);
nor NOR4 (N10769, N10756, N4482, N2637, N10761);
or OR3 (N10770, N7802, N7789, N10146);
nor NOR3 (N10771, N10745, N7001, N2959);
xor XOR2 (N10772, N10769, N3702);
nand NAND3 (N10773, N10770, N10157, N3991);
and AND4 (N10774, N10750, N6229, N2263, N10613);
nor NOR3 (N10775, N10763, N2004, N169);
or OR4 (N10776, N10774, N10174, N5909, N3235);
buf BUF1 (N10777, N10773);
and AND4 (N10778, N10771, N3581, N6387, N10352);
nor NOR2 (N10779, N10765, N8460);
and AND3 (N10780, N10776, N4112, N10089);
or OR3 (N10781, N10775, N5873, N10654);
buf BUF1 (N10782, N10778);
nor NOR2 (N10783, N10767, N2654);
or OR2 (N10784, N10772, N889);
or OR4 (N10785, N10762, N4458, N9227, N10132);
not NOT1 (N10786, N10754);
not NOT1 (N10787, N10781);
not NOT1 (N10788, N10784);
buf BUF1 (N10789, N10788);
buf BUF1 (N10790, N10789);
xor XOR2 (N10791, N10783, N2939);
and AND4 (N10792, N10779, N9262, N3804, N1290);
not NOT1 (N10793, N10786);
buf BUF1 (N10794, N10768);
xor XOR2 (N10795, N10782, N2005);
xor XOR2 (N10796, N10777, N3515);
xor XOR2 (N10797, N10780, N2967);
not NOT1 (N10798, N10793);
nand NAND2 (N10799, N10785, N9565);
or OR2 (N10800, N10799, N10660);
and AND4 (N10801, N10790, N6408, N6809, N4418);
xor XOR2 (N10802, N10796, N3785);
buf BUF1 (N10803, N10792);
not NOT1 (N10804, N10795);
buf BUF1 (N10805, N10802);
nor NOR4 (N10806, N10797, N3640, N9634, N9210);
not NOT1 (N10807, N10794);
nor NOR4 (N10808, N10806, N2459, N3017, N3767);
not NOT1 (N10809, N10791);
or OR3 (N10810, N10808, N4084, N1795);
buf BUF1 (N10811, N10801);
or OR3 (N10812, N10811, N254, N7410);
nor NOR2 (N10813, N10803, N341);
or OR3 (N10814, N10812, N7857, N7088);
buf BUF1 (N10815, N10807);
or OR4 (N10816, N10814, N9828, N2143, N6657);
and AND2 (N10817, N10813, N8316);
xor XOR2 (N10818, N10800, N1764);
buf BUF1 (N10819, N10787);
buf BUF1 (N10820, N10815);
or OR4 (N10821, N10798, N3868, N99, N3446);
not NOT1 (N10822, N10804);
not NOT1 (N10823, N10821);
nor NOR4 (N10824, N10820, N358, N231, N374);
nor NOR4 (N10825, N10818, N10508, N5074, N5250);
nor NOR3 (N10826, N10817, N1072, N7339);
not NOT1 (N10827, N10809);
nand NAND4 (N10828, N10805, N1957, N2529, N2624);
or OR4 (N10829, N10824, N6779, N1111, N1278);
buf BUF1 (N10830, N10827);
nand NAND3 (N10831, N10819, N4714, N2884);
nor NOR2 (N10832, N10826, N3580);
xor XOR2 (N10833, N10822, N1090);
or OR4 (N10834, N10823, N1384, N3532, N2752);
xor XOR2 (N10835, N10816, N9513);
or OR4 (N10836, N10825, N9635, N2416, N969);
or OR2 (N10837, N10830, N6591);
nor NOR4 (N10838, N10829, N502, N6608, N8294);
buf BUF1 (N10839, N10831);
not NOT1 (N10840, N10834);
and AND2 (N10841, N10828, N9711);
nor NOR2 (N10842, N10833, N7909);
and AND3 (N10843, N10810, N6017, N6709);
xor XOR2 (N10844, N10842, N6041);
nand NAND3 (N10845, N10837, N9326, N5430);
and AND2 (N10846, N10843, N1502);
nand NAND3 (N10847, N10844, N2782, N5082);
not NOT1 (N10848, N10846);
not NOT1 (N10849, N10845);
and AND2 (N10850, N10832, N3205);
and AND3 (N10851, N10836, N6939, N131);
or OR2 (N10852, N10851, N5853);
not NOT1 (N10853, N10841);
nand NAND3 (N10854, N10849, N2145, N3382);
nand NAND2 (N10855, N10848, N9769);
buf BUF1 (N10856, N10850);
buf BUF1 (N10857, N10835);
or OR4 (N10858, N10852, N1299, N1414, N10022);
buf BUF1 (N10859, N10856);
buf BUF1 (N10860, N10838);
nand NAND3 (N10861, N10855, N6231, N6496);
nor NOR3 (N10862, N10847, N6881, N8577);
nand NAND2 (N10863, N10853, N7171);
xor XOR2 (N10864, N10839, N676);
buf BUF1 (N10865, N10861);
not NOT1 (N10866, N10859);
not NOT1 (N10867, N10862);
and AND4 (N10868, N10863, N3120, N583, N6804);
and AND3 (N10869, N10867, N3997, N10610);
nor NOR2 (N10870, N10858, N8546);
xor XOR2 (N10871, N10866, N4130);
and AND3 (N10872, N10868, N1855, N4122);
nand NAND2 (N10873, N10865, N7678);
or OR2 (N10874, N10840, N3253);
nor NOR3 (N10875, N10854, N7129, N9858);
nor NOR2 (N10876, N10857, N3393);
nand NAND3 (N10877, N10873, N4981, N5786);
nor NOR3 (N10878, N10860, N10032, N5300);
nand NAND3 (N10879, N10870, N2659, N1549);
xor XOR2 (N10880, N10875, N9335);
xor XOR2 (N10881, N10876, N9559);
not NOT1 (N10882, N10871);
nor NOR4 (N10883, N10880, N8801, N1861, N5444);
nand NAND2 (N10884, N10881, N4436);
nand NAND3 (N10885, N10872, N8313, N9316);
nand NAND3 (N10886, N10883, N10152, N8647);
not NOT1 (N10887, N10886);
nand NAND3 (N10888, N10882, N7854, N8853);
xor XOR2 (N10889, N10869, N6980);
or OR3 (N10890, N10884, N7009, N7384);
xor XOR2 (N10891, N10879, N8780);
not NOT1 (N10892, N10891);
nand NAND3 (N10893, N10874, N9422, N7712);
nand NAND2 (N10894, N10877, N4961);
nand NAND4 (N10895, N10878, N1135, N4802, N1811);
nand NAND3 (N10896, N10885, N2272, N581);
buf BUF1 (N10897, N10894);
not NOT1 (N10898, N10895);
buf BUF1 (N10899, N10888);
and AND2 (N10900, N10898, N7621);
buf BUF1 (N10901, N10889);
buf BUF1 (N10902, N10899);
nor NOR3 (N10903, N10896, N1140, N9850);
or OR3 (N10904, N10897, N9087, N10781);
or OR4 (N10905, N10864, N3173, N6749, N2731);
xor XOR2 (N10906, N10901, N6746);
and AND2 (N10907, N10893, N3704);
and AND4 (N10908, N10904, N3012, N8105, N10756);
not NOT1 (N10909, N10900);
and AND2 (N10910, N10906, N3506);
and AND3 (N10911, N10902, N4909, N9448);
not NOT1 (N10912, N10909);
xor XOR2 (N10913, N10892, N6818);
buf BUF1 (N10914, N10907);
or OR4 (N10915, N10890, N188, N8431, N2264);
xor XOR2 (N10916, N10915, N8958);
xor XOR2 (N10917, N10912, N4981);
and AND4 (N10918, N10913, N5737, N5261, N9251);
and AND2 (N10919, N10903, N9652);
not NOT1 (N10920, N10918);
and AND3 (N10921, N10905, N8807, N2586);
buf BUF1 (N10922, N10919);
buf BUF1 (N10923, N10908);
nand NAND3 (N10924, N10922, N160, N2138);
nor NOR2 (N10925, N10910, N10592);
buf BUF1 (N10926, N10917);
not NOT1 (N10927, N10920);
buf BUF1 (N10928, N10911);
or OR4 (N10929, N10924, N599, N4001, N3168);
not NOT1 (N10930, N10887);
not NOT1 (N10931, N10914);
nand NAND2 (N10932, N10927, N10037);
and AND3 (N10933, N10923, N5179, N2812);
xor XOR2 (N10934, N10926, N6697);
nand NAND2 (N10935, N10929, N8968);
and AND4 (N10936, N10921, N7546, N8491, N291);
xor XOR2 (N10937, N10936, N618);
and AND4 (N10938, N10916, N3239, N1285, N1729);
buf BUF1 (N10939, N10937);
nor NOR2 (N10940, N10935, N2069);
or OR4 (N10941, N10938, N5534, N5732, N1164);
buf BUF1 (N10942, N10928);
nand NAND4 (N10943, N10931, N5523, N7533, N10302);
nor NOR2 (N10944, N10941, N10456);
xor XOR2 (N10945, N10934, N3906);
nor NOR2 (N10946, N10930, N9290);
xor XOR2 (N10947, N10946, N8734);
and AND3 (N10948, N10945, N7684, N4403);
and AND2 (N10949, N10940, N9773);
or OR2 (N10950, N10942, N4121);
not NOT1 (N10951, N10943);
not NOT1 (N10952, N10950);
xor XOR2 (N10953, N10932, N2418);
not NOT1 (N10954, N10925);
buf BUF1 (N10955, N10944);
xor XOR2 (N10956, N10955, N2078);
nand NAND2 (N10957, N10951, N4879);
and AND3 (N10958, N10957, N8751, N4229);
not NOT1 (N10959, N10953);
or OR4 (N10960, N10949, N3117, N8727, N3347);
nor NOR4 (N10961, N10958, N429, N88, N4334);
or OR3 (N10962, N10959, N9470, N1653);
nand NAND2 (N10963, N10962, N9382);
nor NOR3 (N10964, N10939, N9121, N6795);
buf BUF1 (N10965, N10947);
nand NAND3 (N10966, N10961, N6513, N2361);
buf BUF1 (N10967, N10954);
not NOT1 (N10968, N10965);
nand NAND4 (N10969, N10967, N5884, N3606, N8519);
and AND3 (N10970, N10964, N9599, N1612);
or OR2 (N10971, N10956, N457);
nor NOR3 (N10972, N10966, N6095, N7398);
buf BUF1 (N10973, N10971);
buf BUF1 (N10974, N10960);
xor XOR2 (N10975, N10973, N2057);
nor NOR4 (N10976, N10974, N6230, N7813, N9503);
or OR2 (N10977, N10972, N1857);
buf BUF1 (N10978, N10963);
or OR4 (N10979, N10978, N2631, N7411, N3869);
or OR2 (N10980, N10933, N1053);
or OR4 (N10981, N10977, N10808, N8777, N7853);
and AND2 (N10982, N10952, N10104);
not NOT1 (N10983, N10970);
nor NOR2 (N10984, N10980, N7364);
not NOT1 (N10985, N10976);
xor XOR2 (N10986, N10985, N9067);
not NOT1 (N10987, N10975);
or OR2 (N10988, N10948, N4486);
nand NAND3 (N10989, N10986, N2382, N6045);
or OR3 (N10990, N10981, N5554, N7417);
not NOT1 (N10991, N10982);
or OR3 (N10992, N10989, N6752, N8013);
or OR3 (N10993, N10991, N6648, N3479);
buf BUF1 (N10994, N10983);
or OR3 (N10995, N10968, N5751, N7368);
xor XOR2 (N10996, N10993, N8930);
xor XOR2 (N10997, N10990, N357);
and AND4 (N10998, N10994, N1105, N10837, N5571);
buf BUF1 (N10999, N10979);
nand NAND3 (N11000, N10987, N3442, N5928);
nand NAND4 (N11001, N10988, N9623, N8927, N3723);
nor NOR4 (N11002, N11000, N10184, N8607, N810);
and AND4 (N11003, N10996, N8402, N809, N3555);
nor NOR4 (N11004, N10992, N1979, N523, N6909);
nor NOR4 (N11005, N10995, N6500, N5917, N2952);
and AND2 (N11006, N11004, N3549);
and AND4 (N11007, N11001, N10225, N6736, N3068);
xor XOR2 (N11008, N11005, N1479);
xor XOR2 (N11009, N10997, N5685);
nand NAND2 (N11010, N11003, N8101);
or OR2 (N11011, N11006, N7981);
nor NOR2 (N11012, N11011, N10649);
nor NOR2 (N11013, N10999, N7890);
buf BUF1 (N11014, N10969);
xor XOR2 (N11015, N10998, N8944);
nor NOR3 (N11016, N11009, N10014, N5318);
not NOT1 (N11017, N11013);
buf BUF1 (N11018, N11016);
not NOT1 (N11019, N10984);
and AND2 (N11020, N11014, N6932);
or OR2 (N11021, N11017, N1626);
nor NOR2 (N11022, N11020, N10342);
or OR2 (N11023, N11018, N9164);
and AND4 (N11024, N11010, N5170, N1201, N9631);
nand NAND3 (N11025, N11015, N6071, N6952);
nand NAND3 (N11026, N11002, N3918, N3930);
nand NAND2 (N11027, N11022, N5582);
xor XOR2 (N11028, N11021, N2787);
not NOT1 (N11029, N11027);
buf BUF1 (N11030, N11007);
and AND3 (N11031, N11008, N4609, N7588);
xor XOR2 (N11032, N11030, N1972);
nand NAND4 (N11033, N11026, N7175, N7097, N5154);
not NOT1 (N11034, N11028);
or OR4 (N11035, N11032, N6538, N4495, N5896);
or OR4 (N11036, N11019, N3734, N2579, N2707);
nand NAND2 (N11037, N11023, N448);
or OR4 (N11038, N11024, N3222, N10205, N5362);
nor NOR4 (N11039, N11012, N4376, N9148, N2882);
nand NAND4 (N11040, N11035, N10519, N1813, N7442);
xor XOR2 (N11041, N11038, N8363);
not NOT1 (N11042, N11034);
buf BUF1 (N11043, N11036);
not NOT1 (N11044, N11031);
nand NAND4 (N11045, N11043, N13, N4462, N7423);
xor XOR2 (N11046, N11029, N1183);
not NOT1 (N11047, N11041);
xor XOR2 (N11048, N11046, N10869);
nand NAND4 (N11049, N11042, N5038, N452, N3153);
buf BUF1 (N11050, N11039);
buf BUF1 (N11051, N11045);
nand NAND2 (N11052, N11051, N8512);
or OR2 (N11053, N11050, N2839);
buf BUF1 (N11054, N11047);
nand NAND3 (N11055, N11033, N8129, N7274);
buf BUF1 (N11056, N11053);
buf BUF1 (N11057, N11054);
buf BUF1 (N11058, N11057);
buf BUF1 (N11059, N11055);
nor NOR4 (N11060, N11049, N2551, N8414, N169);
and AND4 (N11061, N11058, N4260, N7777, N1617);
xor XOR2 (N11062, N11025, N8810);
nor NOR2 (N11063, N11044, N132);
buf BUF1 (N11064, N11062);
or OR4 (N11065, N11063, N4259, N3230, N8081);
and AND3 (N11066, N11040, N4127, N2157);
not NOT1 (N11067, N11037);
buf BUF1 (N11068, N11061);
nor NOR4 (N11069, N11056, N10330, N8244, N2974);
nand NAND3 (N11070, N11064, N2190, N5224);
xor XOR2 (N11071, N11069, N6742);
and AND3 (N11072, N11071, N5213, N10683);
xor XOR2 (N11073, N11068, N10481);
or OR3 (N11074, N11070, N2894, N3036);
nor NOR4 (N11075, N11060, N8238, N5559, N9873);
and AND2 (N11076, N11066, N6992);
and AND2 (N11077, N11048, N529);
not NOT1 (N11078, N11072);
not NOT1 (N11079, N11075);
not NOT1 (N11080, N11059);
nand NAND4 (N11081, N11065, N1813, N7623, N5298);
nand NAND3 (N11082, N11081, N10821, N7002);
nand NAND2 (N11083, N11080, N10584);
buf BUF1 (N11084, N11077);
buf BUF1 (N11085, N11076);
or OR2 (N11086, N11078, N6216);
and AND4 (N11087, N11084, N3037, N4283, N3286);
buf BUF1 (N11088, N11085);
not NOT1 (N11089, N11087);
nand NAND4 (N11090, N11052, N311, N10629, N536);
nand NAND2 (N11091, N11079, N2943);
or OR2 (N11092, N11082, N5726);
xor XOR2 (N11093, N11074, N1950);
buf BUF1 (N11094, N11083);
buf BUF1 (N11095, N11091);
or OR2 (N11096, N11095, N7438);
nand NAND4 (N11097, N11090, N8192, N10661, N6838);
nand NAND4 (N11098, N11088, N10979, N5076, N5345);
xor XOR2 (N11099, N11092, N9583);
nand NAND2 (N11100, N11093, N5603);
xor XOR2 (N11101, N11094, N8166);
nor NOR2 (N11102, N11073, N6110);
buf BUF1 (N11103, N11102);
or OR3 (N11104, N11089, N1257, N1757);
nor NOR3 (N11105, N11101, N1658, N1515);
nand NAND4 (N11106, N11105, N8222, N8998, N364);
nand NAND2 (N11107, N11100, N1252);
and AND4 (N11108, N11096, N8977, N1303, N2085);
and AND4 (N11109, N11106, N9899, N4604, N7319);
xor XOR2 (N11110, N11108, N7632);
nor NOR2 (N11111, N11107, N5020);
not NOT1 (N11112, N11104);
nor NOR2 (N11113, N11067, N5490);
nor NOR4 (N11114, N11110, N814, N10092, N842);
and AND2 (N11115, N11113, N144);
and AND4 (N11116, N11099, N5598, N2841, N1400);
not NOT1 (N11117, N11111);
nand NAND3 (N11118, N11086, N7593, N9136);
buf BUF1 (N11119, N11116);
nand NAND2 (N11120, N11114, N4257);
nor NOR3 (N11121, N11117, N10930, N4915);
nand NAND4 (N11122, N11109, N494, N8357, N9935);
not NOT1 (N11123, N11103);
and AND2 (N11124, N11121, N4088);
and AND2 (N11125, N11119, N5816);
buf BUF1 (N11126, N11118);
xor XOR2 (N11127, N11125, N6572);
buf BUF1 (N11128, N11115);
nor NOR2 (N11129, N11098, N3243);
not NOT1 (N11130, N11123);
not NOT1 (N11131, N11126);
xor XOR2 (N11132, N11120, N10091);
or OR2 (N11133, N11131, N9267);
or OR3 (N11134, N11133, N9732, N4658);
buf BUF1 (N11135, N11127);
and AND4 (N11136, N11122, N990, N10091, N4238);
buf BUF1 (N11137, N11112);
not NOT1 (N11138, N11124);
nand NAND4 (N11139, N11138, N9756, N8885, N4627);
nor NOR4 (N11140, N11136, N2645, N7513, N6499);
or OR4 (N11141, N11129, N9891, N1757, N11038);
buf BUF1 (N11142, N11130);
not NOT1 (N11143, N11128);
or OR3 (N11144, N11135, N5886, N9241);
or OR4 (N11145, N11097, N5146, N3696, N9995);
xor XOR2 (N11146, N11141, N1381);
not NOT1 (N11147, N11140);
nand NAND2 (N11148, N11134, N2);
and AND3 (N11149, N11139, N7156, N8917);
nand NAND4 (N11150, N11144, N5666, N629, N5042);
not NOT1 (N11151, N11145);
and AND2 (N11152, N11148, N5630);
nand NAND4 (N11153, N11132, N2009, N5704, N8930);
nand NAND3 (N11154, N11142, N6837, N739);
nand NAND2 (N11155, N11152, N11068);
nand NAND3 (N11156, N11146, N7748, N6773);
buf BUF1 (N11157, N11150);
nor NOR3 (N11158, N11151, N853, N52);
or OR3 (N11159, N11149, N269, N3486);
buf BUF1 (N11160, N11137);
buf BUF1 (N11161, N11157);
or OR4 (N11162, N11159, N2211, N1540, N2749);
or OR4 (N11163, N11147, N5514, N1678, N1674);
nor NOR2 (N11164, N11162, N7910);
buf BUF1 (N11165, N11155);
buf BUF1 (N11166, N11164);
or OR4 (N11167, N11161, N909, N415, N2398);
xor XOR2 (N11168, N11158, N4391);
and AND3 (N11169, N11167, N8087, N5686);
buf BUF1 (N11170, N11168);
not NOT1 (N11171, N11154);
and AND4 (N11172, N11156, N3833, N5040, N9928);
nand NAND2 (N11173, N11160, N8535);
buf BUF1 (N11174, N11153);
or OR3 (N11175, N11174, N8583, N1228);
or OR2 (N11176, N11165, N6951);
nand NAND4 (N11177, N11175, N9061, N5781, N1020);
buf BUF1 (N11178, N11170);
nand NAND2 (N11179, N11143, N3616);
buf BUF1 (N11180, N11163);
or OR4 (N11181, N11169, N3925, N6042, N4432);
and AND3 (N11182, N11166, N690, N6624);
and AND4 (N11183, N11182, N1338, N6857, N3298);
nand NAND4 (N11184, N11176, N9764, N872, N139);
xor XOR2 (N11185, N11184, N10501);
nor NOR4 (N11186, N11178, N6041, N8343, N4081);
xor XOR2 (N11187, N11172, N7177);
or OR4 (N11188, N11173, N17, N7977, N766);
not NOT1 (N11189, N11179);
xor XOR2 (N11190, N11171, N5359);
and AND3 (N11191, N11177, N3745, N8041);
not NOT1 (N11192, N11189);
xor XOR2 (N11193, N11192, N587);
nand NAND3 (N11194, N11181, N9543, N6726);
or OR2 (N11195, N11191, N5136);
not NOT1 (N11196, N11187);
nor NOR4 (N11197, N11188, N4908, N8209, N5087);
buf BUF1 (N11198, N11180);
not NOT1 (N11199, N11195);
and AND4 (N11200, N11194, N7869, N5920, N10874);
or OR3 (N11201, N11186, N622, N10974);
not NOT1 (N11202, N11193);
and AND4 (N11203, N11183, N7324, N6470, N7267);
xor XOR2 (N11204, N11185, N7326);
xor XOR2 (N11205, N11201, N10610);
nand NAND2 (N11206, N11199, N10818);
nor NOR4 (N11207, N11202, N8700, N558, N8820);
nand NAND3 (N11208, N11204, N8894, N9930);
or OR2 (N11209, N11207, N2216);
not NOT1 (N11210, N11196);
xor XOR2 (N11211, N11190, N10308);
nor NOR3 (N11212, N11208, N4298, N2664);
nor NOR3 (N11213, N11206, N6206, N8238);
buf BUF1 (N11214, N11211);
nor NOR3 (N11215, N11197, N9838, N2086);
nor NOR2 (N11216, N11210, N7354);
xor XOR2 (N11217, N11216, N1361);
not NOT1 (N11218, N11214);
or OR2 (N11219, N11205, N4166);
nand NAND4 (N11220, N11203, N10433, N1030, N10600);
not NOT1 (N11221, N11219);
buf BUF1 (N11222, N11200);
not NOT1 (N11223, N11213);
nand NAND2 (N11224, N11217, N3364);
or OR2 (N11225, N11215, N1863);
buf BUF1 (N11226, N11221);
or OR3 (N11227, N11226, N4611, N2928);
or OR4 (N11228, N11224, N5272, N493, N4433);
not NOT1 (N11229, N11218);
nand NAND2 (N11230, N11209, N5547);
nand NAND4 (N11231, N11227, N4976, N4999, N3978);
and AND2 (N11232, N11231, N9172);
buf BUF1 (N11233, N11232);
and AND4 (N11234, N11229, N3485, N6155, N7106);
nor NOR3 (N11235, N11230, N2664, N2988);
nor NOR2 (N11236, N11235, N2377);
or OR4 (N11237, N11225, N6095, N1558, N11132);
nor NOR4 (N11238, N11198, N9553, N1276, N4495);
xor XOR2 (N11239, N11212, N4568);
or OR2 (N11240, N11223, N5799);
or OR3 (N11241, N11233, N4018, N4989);
and AND3 (N11242, N11240, N2708, N2145);
and AND4 (N11243, N11239, N3451, N9518, N5646);
and AND2 (N11244, N11220, N4385);
buf BUF1 (N11245, N11242);
xor XOR2 (N11246, N11236, N9171);
or OR4 (N11247, N11222, N135, N3909, N3059);
buf BUF1 (N11248, N11244);
not NOT1 (N11249, N11243);
buf BUF1 (N11250, N11248);
and AND4 (N11251, N11249, N5119, N4840, N5276);
nor NOR2 (N11252, N11237, N6359);
not NOT1 (N11253, N11251);
not NOT1 (N11254, N11253);
and AND3 (N11255, N11252, N3962, N10446);
and AND3 (N11256, N11241, N6588, N5266);
or OR2 (N11257, N11250, N5905);
nand NAND4 (N11258, N11234, N9989, N5512, N1416);
or OR4 (N11259, N11228, N8286, N10564, N1170);
and AND3 (N11260, N11254, N6565, N3825);
and AND2 (N11261, N11259, N6015);
nor NOR3 (N11262, N11246, N3239, N2293);
and AND4 (N11263, N11247, N6820, N8911, N7934);
and AND2 (N11264, N11245, N3110);
and AND4 (N11265, N11255, N4392, N6576, N1281);
not NOT1 (N11266, N11264);
not NOT1 (N11267, N11257);
nand NAND2 (N11268, N11258, N1954);
nor NOR3 (N11269, N11268, N10169, N2359);
or OR3 (N11270, N11260, N2078, N1472);
or OR2 (N11271, N11270, N7630);
and AND2 (N11272, N11271, N2516);
nor NOR4 (N11273, N11272, N811, N3895, N7098);
and AND3 (N11274, N11256, N10468, N2425);
and AND2 (N11275, N11265, N1403);
nor NOR3 (N11276, N11274, N6056, N5804);
nor NOR3 (N11277, N11262, N6086, N1972);
and AND3 (N11278, N11275, N9990, N880);
or OR3 (N11279, N11266, N9476, N5435);
xor XOR2 (N11280, N11278, N3399);
nand NAND3 (N11281, N11261, N9563, N7331);
nor NOR3 (N11282, N11269, N6753, N11138);
and AND2 (N11283, N11277, N6803);
not NOT1 (N11284, N11281);
or OR3 (N11285, N11267, N3841, N10390);
nand NAND4 (N11286, N11285, N1468, N242, N1850);
and AND4 (N11287, N11279, N8370, N7941, N3592);
xor XOR2 (N11288, N11282, N2314);
and AND4 (N11289, N11238, N10910, N3517, N8366);
nor NOR3 (N11290, N11289, N9776, N4876);
buf BUF1 (N11291, N11290);
or OR3 (N11292, N11286, N3872, N8530);
nor NOR4 (N11293, N11291, N8433, N5493, N6891);
or OR3 (N11294, N11276, N2383, N4726);
nor NOR2 (N11295, N11283, N2201);
or OR4 (N11296, N11273, N9609, N9217, N6683);
or OR3 (N11297, N11293, N10652, N10375);
xor XOR2 (N11298, N11294, N3688);
buf BUF1 (N11299, N11297);
xor XOR2 (N11300, N11295, N590);
xor XOR2 (N11301, N11280, N4444);
not NOT1 (N11302, N11284);
xor XOR2 (N11303, N11296, N8206);
or OR2 (N11304, N11300, N4124);
or OR3 (N11305, N11301, N8226, N7430);
nand NAND4 (N11306, N11305, N6895, N9520, N6942);
nor NOR3 (N11307, N11302, N8710, N10892);
xor XOR2 (N11308, N11298, N11016);
buf BUF1 (N11309, N11288);
or OR4 (N11310, N11304, N3274, N4848, N201);
xor XOR2 (N11311, N11307, N1164);
nor NOR3 (N11312, N11299, N2813, N5274);
nor NOR4 (N11313, N11306, N6615, N4110, N8674);
nor NOR3 (N11314, N11287, N2456, N7668);
nor NOR4 (N11315, N11314, N3997, N2154, N4076);
or OR3 (N11316, N11313, N4201, N2069);
xor XOR2 (N11317, N11316, N2278);
or OR3 (N11318, N11292, N10741, N468);
xor XOR2 (N11319, N11312, N810);
or OR2 (N11320, N11315, N1556);
not NOT1 (N11321, N11263);
and AND2 (N11322, N11320, N9282);
nor NOR3 (N11323, N11317, N1730, N5188);
not NOT1 (N11324, N11323);
nand NAND4 (N11325, N11309, N992, N8782, N9970);
xor XOR2 (N11326, N11318, N9387);
nand NAND3 (N11327, N11322, N5603, N931);
or OR4 (N11328, N11325, N9752, N7555, N6147);
and AND2 (N11329, N11319, N2183);
xor XOR2 (N11330, N11310, N2045);
buf BUF1 (N11331, N11311);
xor XOR2 (N11332, N11328, N10701);
and AND4 (N11333, N11308, N10424, N7374, N4963);
and AND3 (N11334, N11331, N8029, N6858);
nand NAND3 (N11335, N11303, N10735, N8744);
nor NOR3 (N11336, N11326, N4973, N4041);
or OR3 (N11337, N11329, N9491, N5960);
xor XOR2 (N11338, N11330, N4564);
xor XOR2 (N11339, N11336, N2654);
or OR3 (N11340, N11327, N7113, N2276);
or OR4 (N11341, N11340, N8173, N4289, N1540);
or OR2 (N11342, N11338, N6671);
not NOT1 (N11343, N11337);
nand NAND3 (N11344, N11324, N7865, N3836);
nand NAND2 (N11345, N11334, N53);
xor XOR2 (N11346, N11342, N491);
nor NOR2 (N11347, N11335, N9172);
nand NAND4 (N11348, N11341, N666, N7897, N6458);
nand NAND2 (N11349, N11345, N7482);
nor NOR2 (N11350, N11349, N3677);
buf BUF1 (N11351, N11339);
or OR3 (N11352, N11348, N8383, N6153);
xor XOR2 (N11353, N11333, N10227);
xor XOR2 (N11354, N11351, N10059);
or OR3 (N11355, N11346, N11251, N1544);
or OR3 (N11356, N11352, N4839, N5476);
nor NOR2 (N11357, N11332, N1651);
not NOT1 (N11358, N11350);
buf BUF1 (N11359, N11357);
nor NOR3 (N11360, N11343, N10104, N7168);
nor NOR2 (N11361, N11321, N7185);
buf BUF1 (N11362, N11360);
nand NAND2 (N11363, N11344, N4583);
buf BUF1 (N11364, N11353);
or OR4 (N11365, N11362, N8988, N2455, N8018);
or OR3 (N11366, N11355, N2618, N6622);
and AND2 (N11367, N11366, N3368);
nor NOR3 (N11368, N11367, N4234, N5729);
nand NAND4 (N11369, N11368, N6002, N463, N4490);
and AND3 (N11370, N11359, N5997, N6170);
or OR2 (N11371, N11370, N5357);
and AND4 (N11372, N11364, N2278, N8302, N7009);
and AND2 (N11373, N11354, N2457);
not NOT1 (N11374, N11361);
nand NAND4 (N11375, N11365, N812, N2906, N3060);
xor XOR2 (N11376, N11373, N7550);
nand NAND4 (N11377, N11376, N800, N7100, N9219);
buf BUF1 (N11378, N11377);
xor XOR2 (N11379, N11372, N5482);
buf BUF1 (N11380, N11371);
not NOT1 (N11381, N11374);
nand NAND3 (N11382, N11356, N604, N5123);
xor XOR2 (N11383, N11378, N2772);
nor NOR4 (N11384, N11347, N5986, N5514, N2446);
xor XOR2 (N11385, N11375, N1191);
buf BUF1 (N11386, N11382);
and AND4 (N11387, N11383, N3393, N5551, N9622);
not NOT1 (N11388, N11385);
nor NOR3 (N11389, N11388, N9432, N2658);
buf BUF1 (N11390, N11381);
or OR2 (N11391, N11358, N4288);
nor NOR2 (N11392, N11379, N394);
nand NAND3 (N11393, N11387, N5808, N6520);
nand NAND4 (N11394, N11363, N5327, N8062, N4353);
buf BUF1 (N11395, N11391);
nand NAND4 (N11396, N11395, N8686, N5303, N1411);
not NOT1 (N11397, N11390);
not NOT1 (N11398, N11384);
buf BUF1 (N11399, N11393);
xor XOR2 (N11400, N11380, N5928);
and AND4 (N11401, N11397, N2136, N6629, N5992);
buf BUF1 (N11402, N11399);
and AND3 (N11403, N11394, N4479, N6206);
xor XOR2 (N11404, N11400, N3082);
buf BUF1 (N11405, N11389);
buf BUF1 (N11406, N11401);
or OR3 (N11407, N11403, N9348, N1373);
not NOT1 (N11408, N11402);
nor NOR2 (N11409, N11405, N203);
xor XOR2 (N11410, N11407, N5700);
nand NAND2 (N11411, N11406, N9035);
nand NAND2 (N11412, N11398, N10757);
and AND4 (N11413, N11408, N6781, N1228, N5059);
or OR2 (N11414, N11409, N705);
or OR2 (N11415, N11411, N3603);
and AND3 (N11416, N11386, N9817, N7778);
nand NAND4 (N11417, N11414, N9528, N10226, N1066);
buf BUF1 (N11418, N11410);
buf BUF1 (N11419, N11392);
buf BUF1 (N11420, N11419);
and AND4 (N11421, N11396, N7082, N4799, N3084);
or OR4 (N11422, N11415, N2999, N8403, N1752);
and AND3 (N11423, N11404, N10908, N2582);
nand NAND4 (N11424, N11418, N4928, N6699, N2843);
and AND2 (N11425, N11417, N3962);
and AND3 (N11426, N11421, N9456, N9141);
not NOT1 (N11427, N11412);
not NOT1 (N11428, N11420);
xor XOR2 (N11429, N11423, N2478);
or OR4 (N11430, N11429, N7576, N7946, N9279);
not NOT1 (N11431, N11416);
or OR2 (N11432, N11413, N6793);
or OR2 (N11433, N11431, N6937);
or OR2 (N11434, N11426, N332);
or OR2 (N11435, N11428, N7086);
xor XOR2 (N11436, N11434, N11111);
not NOT1 (N11437, N11436);
nand NAND4 (N11438, N11433, N1413, N3079, N1403);
not NOT1 (N11439, N11435);
or OR3 (N11440, N11430, N3171, N3104);
buf BUF1 (N11441, N11437);
xor XOR2 (N11442, N11438, N1856);
buf BUF1 (N11443, N11422);
not NOT1 (N11444, N11369);
nor NOR2 (N11445, N11424, N3635);
nor NOR2 (N11446, N11444, N6888);
not NOT1 (N11447, N11440);
not NOT1 (N11448, N11442);
xor XOR2 (N11449, N11443, N2458);
not NOT1 (N11450, N11446);
nand NAND4 (N11451, N11445, N4274, N4707, N7892);
not NOT1 (N11452, N11448);
and AND3 (N11453, N11447, N526, N2101);
xor XOR2 (N11454, N11451, N10773);
and AND2 (N11455, N11454, N9157);
nand NAND2 (N11456, N11450, N5638);
buf BUF1 (N11457, N11456);
nand NAND3 (N11458, N11449, N3795, N2177);
not NOT1 (N11459, N11425);
buf BUF1 (N11460, N11439);
nand NAND4 (N11461, N11458, N5655, N10419, N5471);
and AND4 (N11462, N11461, N6132, N7706, N7640);
and AND2 (N11463, N11462, N4091);
and AND2 (N11464, N11457, N3042);
not NOT1 (N11465, N11459);
not NOT1 (N11466, N11460);
not NOT1 (N11467, N11463);
buf BUF1 (N11468, N11453);
buf BUF1 (N11469, N11452);
buf BUF1 (N11470, N11468);
and AND2 (N11471, N11441, N1631);
nor NOR2 (N11472, N11466, N5563);
nand NAND2 (N11473, N11470, N9284);
buf BUF1 (N11474, N11469);
xor XOR2 (N11475, N11474, N4447);
and AND4 (N11476, N11467, N9256, N10430, N9352);
not NOT1 (N11477, N11465);
buf BUF1 (N11478, N11455);
not NOT1 (N11479, N11472);
nand NAND2 (N11480, N11427, N4853);
xor XOR2 (N11481, N11480, N5405);
xor XOR2 (N11482, N11479, N4786);
nand NAND3 (N11483, N11432, N2648, N6431);
xor XOR2 (N11484, N11473, N5283);
nor NOR3 (N11485, N11481, N5404, N5927);
buf BUF1 (N11486, N11484);
nor NOR2 (N11487, N11476, N9959);
and AND4 (N11488, N11485, N7925, N1791, N2218);
not NOT1 (N11489, N11488);
buf BUF1 (N11490, N11487);
or OR4 (N11491, N11482, N10170, N7502, N3026);
xor XOR2 (N11492, N11483, N5909);
buf BUF1 (N11493, N11464);
xor XOR2 (N11494, N11490, N10098);
or OR2 (N11495, N11489, N7512);
nand NAND4 (N11496, N11475, N6756, N10813, N9222);
nand NAND4 (N11497, N11492, N9048, N1390, N4237);
nand NAND3 (N11498, N11493, N338, N8792);
and AND4 (N11499, N11478, N3637, N105, N7753);
and AND3 (N11500, N11477, N7856, N11281);
buf BUF1 (N11501, N11499);
and AND2 (N11502, N11496, N1504);
buf BUF1 (N11503, N11491);
buf BUF1 (N11504, N11486);
nor NOR4 (N11505, N11494, N8309, N641, N10700);
and AND3 (N11506, N11502, N9936, N7650);
buf BUF1 (N11507, N11498);
buf BUF1 (N11508, N11507);
xor XOR2 (N11509, N11501, N11229);
buf BUF1 (N11510, N11509);
nand NAND4 (N11511, N11471, N2950, N4249, N4800);
xor XOR2 (N11512, N11510, N9484);
nand NAND4 (N11513, N11512, N2747, N936, N9043);
buf BUF1 (N11514, N11500);
xor XOR2 (N11515, N11514, N4413);
nand NAND2 (N11516, N11506, N10615);
xor XOR2 (N11517, N11511, N5240);
nor NOR3 (N11518, N11504, N6867, N9983);
buf BUF1 (N11519, N11508);
not NOT1 (N11520, N11515);
nand NAND2 (N11521, N11497, N8460);
and AND2 (N11522, N11518, N6837);
and AND4 (N11523, N11522, N9339, N9101, N8311);
nand NAND2 (N11524, N11495, N1396);
nand NAND2 (N11525, N11517, N3019);
not NOT1 (N11526, N11505);
nand NAND3 (N11527, N11516, N2413, N1792);
buf BUF1 (N11528, N11520);
buf BUF1 (N11529, N11528);
buf BUF1 (N11530, N11503);
and AND3 (N11531, N11523, N10941, N4086);
and AND4 (N11532, N11525, N6670, N7146, N7578);
nand NAND3 (N11533, N11530, N4618, N2921);
xor XOR2 (N11534, N11527, N10666);
nand NAND4 (N11535, N11526, N1202, N4309, N2719);
buf BUF1 (N11536, N11531);
xor XOR2 (N11537, N11521, N3449);
and AND4 (N11538, N11533, N1174, N6373, N11262);
xor XOR2 (N11539, N11529, N9867);
nor NOR3 (N11540, N11535, N2537, N8089);
and AND3 (N11541, N11532, N9168, N3403);
xor XOR2 (N11542, N11539, N4365);
xor XOR2 (N11543, N11541, N5383);
nor NOR3 (N11544, N11542, N2764, N1328);
buf BUF1 (N11545, N11513);
xor XOR2 (N11546, N11540, N6437);
and AND3 (N11547, N11543, N4973, N10782);
xor XOR2 (N11548, N11536, N1153);
not NOT1 (N11549, N11547);
nand NAND3 (N11550, N11546, N7488, N2736);
buf BUF1 (N11551, N11537);
nor NOR4 (N11552, N11534, N5961, N10914, N10258);
nand NAND4 (N11553, N11552, N4141, N3323, N2338);
nor NOR2 (N11554, N11545, N6065);
not NOT1 (N11555, N11550);
or OR2 (N11556, N11544, N8783);
xor XOR2 (N11557, N11538, N2820);
or OR3 (N11558, N11548, N8638, N6037);
xor XOR2 (N11559, N11549, N8175);
xor XOR2 (N11560, N11556, N2942);
nor NOR2 (N11561, N11557, N9297);
nor NOR4 (N11562, N11561, N9182, N4723, N5193);
nor NOR4 (N11563, N11555, N1976, N61, N8933);
nor NOR3 (N11564, N11554, N214, N3970);
not NOT1 (N11565, N11564);
xor XOR2 (N11566, N11565, N1551);
buf BUF1 (N11567, N11551);
nand NAND2 (N11568, N11560, N502);
nand NAND3 (N11569, N11559, N3677, N7500);
or OR3 (N11570, N11569, N11516, N9753);
nor NOR4 (N11571, N11570, N3116, N502, N10883);
buf BUF1 (N11572, N11567);
buf BUF1 (N11573, N11572);
or OR3 (N11574, N11558, N1146, N8330);
or OR4 (N11575, N11568, N2650, N8080, N7925);
xor XOR2 (N11576, N11574, N2103);
and AND4 (N11577, N11573, N9534, N3591, N4587);
nand NAND4 (N11578, N11553, N1261, N3014, N4416);
nor NOR4 (N11579, N11575, N9396, N10077, N9823);
nand NAND2 (N11580, N11578, N7380);
buf BUF1 (N11581, N11566);
nor NOR2 (N11582, N11571, N5260);
not NOT1 (N11583, N11577);
buf BUF1 (N11584, N11583);
buf BUF1 (N11585, N11576);
and AND4 (N11586, N11524, N9449, N7500, N4258);
nor NOR4 (N11587, N11580, N1876, N6331, N7120);
xor XOR2 (N11588, N11584, N10637);
not NOT1 (N11589, N11563);
and AND2 (N11590, N11562, N10230);
nor NOR3 (N11591, N11586, N5749, N7071);
buf BUF1 (N11592, N11588);
nand NAND2 (N11593, N11592, N269);
or OR4 (N11594, N11590, N2516, N800, N2868);
xor XOR2 (N11595, N11591, N8964);
and AND2 (N11596, N11595, N2123);
xor XOR2 (N11597, N11585, N5310);
buf BUF1 (N11598, N11597);
nand NAND3 (N11599, N11589, N6654, N11339);
buf BUF1 (N11600, N11587);
and AND3 (N11601, N11594, N5367, N6657);
and AND3 (N11602, N11519, N9508, N3837);
xor XOR2 (N11603, N11579, N3343);
and AND4 (N11604, N11598, N4347, N11209, N5287);
nand NAND4 (N11605, N11601, N11567, N2957, N10957);
nand NAND4 (N11606, N11593, N11282, N5452, N9362);
and AND4 (N11607, N11604, N8493, N6206, N900);
and AND4 (N11608, N11600, N10700, N6832, N9599);
or OR4 (N11609, N11605, N11172, N2917, N5585);
not NOT1 (N11610, N11596);
and AND2 (N11611, N11608, N3014);
buf BUF1 (N11612, N11607);
or OR3 (N11613, N11599, N3195, N2188);
xor XOR2 (N11614, N11602, N8408);
and AND3 (N11615, N11611, N7591, N4182);
not NOT1 (N11616, N11610);
or OR4 (N11617, N11612, N10348, N6113, N1507);
nand NAND2 (N11618, N11616, N8154);
and AND3 (N11619, N11581, N7481, N445);
buf BUF1 (N11620, N11618);
and AND4 (N11621, N11606, N2083, N5927, N3126);
buf BUF1 (N11622, N11613);
not NOT1 (N11623, N11621);
and AND3 (N11624, N11620, N8211, N9175);
or OR2 (N11625, N11619, N3938);
buf BUF1 (N11626, N11624);
xor XOR2 (N11627, N11617, N5379);
or OR3 (N11628, N11615, N10838, N10124);
and AND4 (N11629, N11603, N5131, N6670, N5780);
or OR2 (N11630, N11626, N5158);
nand NAND2 (N11631, N11629, N9774);
nor NOR4 (N11632, N11627, N778, N3332, N152);
and AND4 (N11633, N11614, N9924, N9551, N10757);
and AND3 (N11634, N11630, N3994, N10408);
xor XOR2 (N11635, N11632, N7498);
not NOT1 (N11636, N11634);
xor XOR2 (N11637, N11633, N621);
xor XOR2 (N11638, N11637, N9529);
nand NAND4 (N11639, N11625, N6168, N10430, N7676);
nor NOR4 (N11640, N11631, N7941, N5381, N5191);
not NOT1 (N11641, N11628);
or OR4 (N11642, N11635, N10309, N8597, N6333);
nor NOR4 (N11643, N11639, N3242, N1133, N10155);
nor NOR2 (N11644, N11622, N1798);
nor NOR2 (N11645, N11582, N8884);
not NOT1 (N11646, N11645);
xor XOR2 (N11647, N11641, N1111);
buf BUF1 (N11648, N11609);
not NOT1 (N11649, N11644);
or OR2 (N11650, N11647, N525);
and AND4 (N11651, N11642, N10499, N9357, N5578);
buf BUF1 (N11652, N11643);
not NOT1 (N11653, N11648);
not NOT1 (N11654, N11652);
nand NAND2 (N11655, N11640, N7631);
or OR4 (N11656, N11651, N4455, N7380, N5650);
xor XOR2 (N11657, N11649, N11384);
and AND2 (N11658, N11653, N4581);
buf BUF1 (N11659, N11656);
nor NOR2 (N11660, N11646, N5704);
xor XOR2 (N11661, N11623, N1763);
not NOT1 (N11662, N11636);
and AND3 (N11663, N11655, N8631, N10076);
xor XOR2 (N11664, N11658, N10051);
nor NOR2 (N11665, N11657, N628);
xor XOR2 (N11666, N11663, N461);
buf BUF1 (N11667, N11660);
buf BUF1 (N11668, N11659);
or OR2 (N11669, N11668, N6220);
nor NOR3 (N11670, N11662, N4344, N5748);
buf BUF1 (N11671, N11669);
and AND4 (N11672, N11665, N10002, N3874, N2855);
xor XOR2 (N11673, N11664, N4622);
not NOT1 (N11674, N11667);
nor NOR4 (N11675, N11661, N11006, N256, N3104);
and AND3 (N11676, N11675, N4053, N10307);
buf BUF1 (N11677, N11670);
nor NOR3 (N11678, N11674, N4884, N4859);
nor NOR4 (N11679, N11650, N7256, N10485, N866);
buf BUF1 (N11680, N11676);
buf BUF1 (N11681, N11679);
buf BUF1 (N11682, N11671);
or OR4 (N11683, N11673, N8553, N8459, N6016);
nor NOR4 (N11684, N11666, N4662, N10256, N1044);
xor XOR2 (N11685, N11681, N8679);
nand NAND3 (N11686, N11678, N1843, N5059);
nand NAND3 (N11687, N11684, N10327, N2915);
buf BUF1 (N11688, N11682);
xor XOR2 (N11689, N11687, N6786);
xor XOR2 (N11690, N11688, N6082);
not NOT1 (N11691, N11638);
nor NOR3 (N11692, N11685, N4248, N3273);
buf BUF1 (N11693, N11680);
or OR4 (N11694, N11693, N7514, N8208, N10329);
not NOT1 (N11695, N11686);
xor XOR2 (N11696, N11691, N10179);
nor NOR4 (N11697, N11695, N3942, N5892, N7161);
buf BUF1 (N11698, N11690);
buf BUF1 (N11699, N11692);
nor NOR2 (N11700, N11683, N2924);
not NOT1 (N11701, N11694);
xor XOR2 (N11702, N11700, N11206);
or OR3 (N11703, N11698, N10540, N2277);
nand NAND2 (N11704, N11654, N3014);
and AND3 (N11705, N11677, N1338, N6964);
and AND2 (N11706, N11702, N9106);
or OR3 (N11707, N11705, N201, N4810);
nand NAND2 (N11708, N11701, N1604);
not NOT1 (N11709, N11703);
xor XOR2 (N11710, N11697, N11412);
and AND2 (N11711, N11709, N632);
and AND3 (N11712, N11711, N2291, N11274);
nor NOR4 (N11713, N11672, N5455, N1412, N1030);
not NOT1 (N11714, N11704);
and AND3 (N11715, N11713, N10986, N8585);
buf BUF1 (N11716, N11706);
and AND3 (N11717, N11699, N5665, N138);
xor XOR2 (N11718, N11714, N10525);
or OR2 (N11719, N11715, N881);
or OR4 (N11720, N11712, N7298, N1713, N5910);
and AND2 (N11721, N11720, N135);
and AND4 (N11722, N11721, N236, N7020, N8723);
xor XOR2 (N11723, N11689, N1137);
or OR2 (N11724, N11707, N11201);
nor NOR3 (N11725, N11718, N1850, N11480);
nor NOR2 (N11726, N11708, N1568);
and AND4 (N11727, N11710, N3162, N10579, N5776);
xor XOR2 (N11728, N11716, N265);
xor XOR2 (N11729, N11727, N1630);
xor XOR2 (N11730, N11724, N9760);
buf BUF1 (N11731, N11719);
nor NOR4 (N11732, N11717, N10336, N3291, N6961);
buf BUF1 (N11733, N11696);
buf BUF1 (N11734, N11726);
and AND3 (N11735, N11729, N2713, N9682);
and AND3 (N11736, N11732, N4844, N1240);
buf BUF1 (N11737, N11734);
xor XOR2 (N11738, N11737, N3243);
and AND4 (N11739, N11733, N30, N8632, N8627);
xor XOR2 (N11740, N11725, N5500);
and AND2 (N11741, N11738, N4034);
not NOT1 (N11742, N11722);
nor NOR3 (N11743, N11723, N2591, N1295);
not NOT1 (N11744, N11741);
and AND4 (N11745, N11739, N6863, N11681, N11732);
and AND4 (N11746, N11731, N4305, N3241, N526);
nor NOR2 (N11747, N11745, N1547);
nand NAND2 (N11748, N11730, N7482);
xor XOR2 (N11749, N11743, N3606);
nor NOR2 (N11750, N11747, N4432);
nor NOR2 (N11751, N11740, N5015);
xor XOR2 (N11752, N11742, N10775);
xor XOR2 (N11753, N11751, N5159);
nand NAND3 (N11754, N11752, N4619, N7098);
xor XOR2 (N11755, N11749, N6210);
buf BUF1 (N11756, N11750);
nand NAND3 (N11757, N11736, N1442, N549);
or OR3 (N11758, N11755, N10765, N1813);
or OR4 (N11759, N11754, N10194, N4581, N7035);
not NOT1 (N11760, N11728);
nand NAND3 (N11761, N11748, N4643, N10580);
xor XOR2 (N11762, N11757, N8690);
buf BUF1 (N11763, N11753);
nor NOR2 (N11764, N11758, N7539);
or OR3 (N11765, N11756, N8516, N8755);
and AND4 (N11766, N11761, N3275, N7425, N1646);
or OR3 (N11767, N11763, N10903, N6221);
nand NAND2 (N11768, N11746, N9512);
not NOT1 (N11769, N11765);
or OR4 (N11770, N11767, N6066, N1810, N3407);
nand NAND2 (N11771, N11762, N8698);
not NOT1 (N11772, N11771);
xor XOR2 (N11773, N11760, N5952);
nor NOR3 (N11774, N11773, N6139, N3682);
and AND2 (N11775, N11768, N6320);
buf BUF1 (N11776, N11770);
buf BUF1 (N11777, N11744);
or OR3 (N11778, N11775, N3265, N179);
xor XOR2 (N11779, N11772, N1325);
nand NAND3 (N11780, N11764, N896, N5968);
nand NAND2 (N11781, N11777, N1481);
buf BUF1 (N11782, N11769);
or OR2 (N11783, N11782, N4203);
nand NAND4 (N11784, N11781, N8458, N1086, N2260);
not NOT1 (N11785, N11783);
and AND4 (N11786, N11780, N6804, N5201, N3481);
nor NOR2 (N11787, N11774, N2450);
and AND4 (N11788, N11759, N11493, N2969, N1566);
nor NOR4 (N11789, N11776, N9679, N9935, N3343);
or OR4 (N11790, N11766, N10798, N6742, N10540);
xor XOR2 (N11791, N11787, N7705);
or OR2 (N11792, N11790, N3985);
xor XOR2 (N11793, N11789, N10674);
and AND4 (N11794, N11779, N10806, N336, N10447);
not NOT1 (N11795, N11793);
nor NOR4 (N11796, N11794, N2252, N1779, N7035);
not NOT1 (N11797, N11735);
or OR4 (N11798, N11788, N7264, N6060, N11408);
nand NAND4 (N11799, N11797, N11101, N8432, N9915);
nand NAND4 (N11800, N11778, N3096, N3411, N4261);
buf BUF1 (N11801, N11785);
and AND2 (N11802, N11801, N4795);
nand NAND2 (N11803, N11784, N6308);
nand NAND3 (N11804, N11802, N2743, N7100);
or OR4 (N11805, N11799, N6317, N987, N3326);
buf BUF1 (N11806, N11803);
nor NOR3 (N11807, N11804, N7143, N4165);
xor XOR2 (N11808, N11800, N9546);
nand NAND3 (N11809, N11795, N1400, N3027);
and AND4 (N11810, N11805, N9261, N4062, N2915);
and AND2 (N11811, N11792, N9774);
buf BUF1 (N11812, N11791);
buf BUF1 (N11813, N11812);
and AND2 (N11814, N11806, N2993);
buf BUF1 (N11815, N11811);
xor XOR2 (N11816, N11815, N7308);
or OR3 (N11817, N11809, N769, N5635);
not NOT1 (N11818, N11808);
nand NAND2 (N11819, N11786, N4672);
or OR3 (N11820, N11819, N9587, N10212);
nor NOR3 (N11821, N11810, N10967, N1700);
and AND3 (N11822, N11814, N8779, N5987);
and AND4 (N11823, N11820, N2246, N4246, N3157);
nand NAND2 (N11824, N11822, N5271);
and AND4 (N11825, N11821, N10246, N7624, N4990);
nor NOR3 (N11826, N11823, N8074, N8549);
and AND2 (N11827, N11816, N9037);
nor NOR3 (N11828, N11824, N1152, N7308);
nor NOR4 (N11829, N11798, N2957, N6557, N9203);
nor NOR3 (N11830, N11829, N11605, N7697);
or OR4 (N11831, N11817, N8107, N7953, N9919);
buf BUF1 (N11832, N11831);
not NOT1 (N11833, N11818);
not NOT1 (N11834, N11828);
nand NAND2 (N11835, N11826, N2267);
nor NOR4 (N11836, N11825, N571, N11586, N8477);
nor NOR3 (N11837, N11834, N3531, N3888);
nor NOR4 (N11838, N11837, N8813, N10415, N9621);
buf BUF1 (N11839, N11838);
and AND3 (N11840, N11832, N593, N4589);
not NOT1 (N11841, N11833);
and AND4 (N11842, N11839, N530, N10533, N9336);
and AND4 (N11843, N11841, N8670, N7491, N4964);
nand NAND4 (N11844, N11835, N1388, N6716, N1499);
nand NAND2 (N11845, N11842, N7618);
nand NAND2 (N11846, N11827, N838);
or OR3 (N11847, N11796, N7008, N11668);
xor XOR2 (N11848, N11836, N1623);
buf BUF1 (N11849, N11830);
or OR3 (N11850, N11846, N4131, N2392);
xor XOR2 (N11851, N11845, N8386);
buf BUF1 (N11852, N11850);
and AND3 (N11853, N11844, N8921, N11198);
buf BUF1 (N11854, N11843);
or OR2 (N11855, N11849, N7451);
not NOT1 (N11856, N11848);
nand NAND2 (N11857, N11840, N6211);
buf BUF1 (N11858, N11854);
buf BUF1 (N11859, N11858);
or OR3 (N11860, N11856, N10192, N10477);
nand NAND3 (N11861, N11860, N8048, N10298);
nand NAND4 (N11862, N11852, N8106, N9750, N9754);
nor NOR3 (N11863, N11807, N11035, N1026);
nand NAND2 (N11864, N11861, N9482);
not NOT1 (N11865, N11853);
nand NAND3 (N11866, N11851, N9710, N10289);
xor XOR2 (N11867, N11847, N677);
and AND2 (N11868, N11867, N703);
and AND2 (N11869, N11855, N4041);
or OR2 (N11870, N11862, N6625);
not NOT1 (N11871, N11859);
and AND4 (N11872, N11865, N2008, N5867, N6279);
nand NAND2 (N11873, N11813, N4898);
xor XOR2 (N11874, N11863, N7914);
nor NOR3 (N11875, N11866, N10851, N4083);
and AND2 (N11876, N11857, N7718);
buf BUF1 (N11877, N11864);
nand NAND2 (N11878, N11869, N3192);
nand NAND3 (N11879, N11872, N4441, N7626);
or OR3 (N11880, N11879, N10069, N6543);
xor XOR2 (N11881, N11878, N10487);
xor XOR2 (N11882, N11874, N9013);
buf BUF1 (N11883, N11880);
or OR3 (N11884, N11881, N9678, N987);
not NOT1 (N11885, N11868);
xor XOR2 (N11886, N11875, N7637);
and AND4 (N11887, N11884, N9852, N3152, N2811);
and AND3 (N11888, N11887, N6114, N3061);
or OR3 (N11889, N11888, N4270, N8009);
buf BUF1 (N11890, N11882);
or OR2 (N11891, N11885, N8829);
xor XOR2 (N11892, N11870, N10714);
not NOT1 (N11893, N11876);
nand NAND3 (N11894, N11891, N570, N6802);
xor XOR2 (N11895, N11894, N10295);
xor XOR2 (N11896, N11873, N3255);
buf BUF1 (N11897, N11890);
buf BUF1 (N11898, N11895);
nand NAND2 (N11899, N11886, N2521);
buf BUF1 (N11900, N11898);
nand NAND4 (N11901, N11889, N444, N5256, N1917);
not NOT1 (N11902, N11901);
xor XOR2 (N11903, N11899, N11745);
nand NAND3 (N11904, N11900, N9274, N3235);
not NOT1 (N11905, N11897);
and AND3 (N11906, N11905, N5233, N5382);
or OR4 (N11907, N11871, N10503, N7933, N6352);
and AND2 (N11908, N11893, N7849);
xor XOR2 (N11909, N11906, N8725);
and AND3 (N11910, N11903, N6419, N1324);
and AND3 (N11911, N11904, N9128, N8909);
xor XOR2 (N11912, N11910, N1878);
nand NAND3 (N11913, N11911, N631, N6452);
and AND3 (N11914, N11912, N9120, N9901);
nand NAND2 (N11915, N11914, N5560);
buf BUF1 (N11916, N11896);
xor XOR2 (N11917, N11902, N4004);
not NOT1 (N11918, N11908);
or OR2 (N11919, N11916, N699);
buf BUF1 (N11920, N11892);
not NOT1 (N11921, N11917);
or OR3 (N11922, N11877, N11219, N174);
or OR3 (N11923, N11922, N2184, N3786);
not NOT1 (N11924, N11913);
buf BUF1 (N11925, N11919);
xor XOR2 (N11926, N11883, N3775);
nand NAND3 (N11927, N11923, N11181, N8247);
not NOT1 (N11928, N11920);
nand NAND4 (N11929, N11915, N7777, N10487, N9559);
and AND2 (N11930, N11928, N2762);
not NOT1 (N11931, N11907);
and AND2 (N11932, N11909, N1158);
nor NOR4 (N11933, N11925, N5565, N8052, N5398);
nand NAND4 (N11934, N11933, N9891, N1042, N7593);
buf BUF1 (N11935, N11934);
or OR4 (N11936, N11924, N11783, N6919, N5967);
xor XOR2 (N11937, N11929, N9440);
nand NAND4 (N11938, N11932, N11040, N6419, N906);
and AND3 (N11939, N11931, N5608, N2116);
not NOT1 (N11940, N11930);
or OR2 (N11941, N11921, N6493);
buf BUF1 (N11942, N11926);
buf BUF1 (N11943, N11938);
nor NOR3 (N11944, N11927, N914, N6956);
nand NAND2 (N11945, N11940, N11868);
xor XOR2 (N11946, N11937, N8377);
not NOT1 (N11947, N11939);
buf BUF1 (N11948, N11918);
not NOT1 (N11949, N11935);
and AND3 (N11950, N11946, N11493, N779);
nor NOR3 (N11951, N11949, N1860, N4378);
xor XOR2 (N11952, N11943, N8041);
nand NAND3 (N11953, N11942, N269, N5484);
or OR3 (N11954, N11947, N11000, N3553);
buf BUF1 (N11955, N11941);
nand NAND4 (N11956, N11945, N2388, N2986, N9580);
not NOT1 (N11957, N11951);
or OR3 (N11958, N11952, N6411, N4529);
xor XOR2 (N11959, N11955, N6534);
xor XOR2 (N11960, N11959, N6489);
buf BUF1 (N11961, N11954);
buf BUF1 (N11962, N11948);
nand NAND4 (N11963, N11962, N7842, N3791, N1719);
nand NAND2 (N11964, N11950, N8056);
xor XOR2 (N11965, N11957, N9284);
nor NOR4 (N11966, N11963, N9621, N7392, N3950);
or OR4 (N11967, N11936, N7846, N689, N5359);
not NOT1 (N11968, N11958);
xor XOR2 (N11969, N11944, N6918);
or OR3 (N11970, N11966, N9122, N1549);
xor XOR2 (N11971, N11961, N3679);
and AND2 (N11972, N11971, N10850);
and AND3 (N11973, N11969, N392, N9989);
buf BUF1 (N11974, N11970);
xor XOR2 (N11975, N11964, N11231);
and AND4 (N11976, N11965, N11656, N391, N10420);
and AND3 (N11977, N11953, N7319, N8931);
or OR3 (N11978, N11956, N2731, N10748);
or OR3 (N11979, N11967, N11371, N4877);
nor NOR2 (N11980, N11979, N8959);
nor NOR3 (N11981, N11976, N11717, N8871);
not NOT1 (N11982, N11981);
buf BUF1 (N11983, N11977);
buf BUF1 (N11984, N11980);
or OR2 (N11985, N11973, N3433);
nand NAND2 (N11986, N11982, N11199);
not NOT1 (N11987, N11972);
not NOT1 (N11988, N11987);
not NOT1 (N11989, N11960);
buf BUF1 (N11990, N11968);
nor NOR3 (N11991, N11984, N9927, N4292);
xor XOR2 (N11992, N11985, N9036);
and AND3 (N11993, N11988, N5430, N2017);
or OR2 (N11994, N11983, N8171);
and AND3 (N11995, N11990, N9108, N7081);
and AND2 (N11996, N11993, N9299);
nor NOR2 (N11997, N11989, N3188);
buf BUF1 (N11998, N11986);
nor NOR4 (N11999, N11996, N5553, N11750, N6344);
nor NOR3 (N12000, N11997, N11194, N8458);
xor XOR2 (N12001, N11975, N3306);
nand NAND3 (N12002, N11991, N8125, N2999);
and AND4 (N12003, N11992, N7616, N5026, N5794);
and AND3 (N12004, N11974, N9191, N2157);
nor NOR3 (N12005, N11978, N2340, N3996);
buf BUF1 (N12006, N12001);
and AND3 (N12007, N12003, N5840, N4654);
and AND2 (N12008, N12004, N8617);
nand NAND2 (N12009, N12008, N5824);
xor XOR2 (N12010, N11994, N5132);
and AND2 (N12011, N12002, N9982);
not NOT1 (N12012, N12011);
nor NOR4 (N12013, N12005, N5839, N9265, N1701);
and AND3 (N12014, N12013, N9874, N232);
nand NAND2 (N12015, N12006, N884);
or OR3 (N12016, N12000, N9494, N7561);
and AND2 (N12017, N12015, N3381);
not NOT1 (N12018, N11995);
or OR3 (N12019, N12018, N4478, N7746);
xor XOR2 (N12020, N12017, N8588);
and AND4 (N12021, N12009, N11411, N1423, N8767);
xor XOR2 (N12022, N12019, N10288);
nor NOR2 (N12023, N11998, N2314);
not NOT1 (N12024, N12016);
buf BUF1 (N12025, N12023);
nor NOR4 (N12026, N12020, N7241, N6955, N3815);
xor XOR2 (N12027, N12026, N30);
not NOT1 (N12028, N12007);
nand NAND3 (N12029, N12012, N6232, N7124);
nor NOR2 (N12030, N12022, N6185);
or OR3 (N12031, N12027, N1042, N2601);
and AND4 (N12032, N12028, N4920, N8778, N286);
xor XOR2 (N12033, N12031, N1297);
not NOT1 (N12034, N12021);
not NOT1 (N12035, N12025);
xor XOR2 (N12036, N12033, N1938);
or OR4 (N12037, N12024, N7569, N8279, N1016);
not NOT1 (N12038, N12010);
not NOT1 (N12039, N12037);
or OR3 (N12040, N12030, N1352, N3804);
and AND2 (N12041, N12039, N8286);
nand NAND4 (N12042, N12034, N1014, N8883, N8806);
or OR4 (N12043, N11999, N3682, N10414, N4404);
xor XOR2 (N12044, N12036, N10151);
buf BUF1 (N12045, N12041);
nand NAND3 (N12046, N12044, N6355, N4169);
not NOT1 (N12047, N12035);
nand NAND4 (N12048, N12029, N11226, N7501, N2351);
and AND2 (N12049, N12047, N1593);
xor XOR2 (N12050, N12048, N2458);
nor NOR2 (N12051, N12045, N10015);
buf BUF1 (N12052, N12038);
not NOT1 (N12053, N12046);
nor NOR2 (N12054, N12042, N2732);
xor XOR2 (N12055, N12032, N4811);
nor NOR4 (N12056, N12053, N9904, N9188, N7390);
nor NOR2 (N12057, N12040, N10623);
not NOT1 (N12058, N12050);
or OR4 (N12059, N12051, N8262, N5607, N6922);
nand NAND2 (N12060, N12043, N11254);
nor NOR2 (N12061, N12060, N9266);
buf BUF1 (N12062, N12056);
and AND2 (N12063, N12059, N715);
or OR2 (N12064, N12054, N2622);
and AND2 (N12065, N12064, N6434);
not NOT1 (N12066, N12062);
xor XOR2 (N12067, N12052, N5713);
xor XOR2 (N12068, N12066, N8182);
or OR4 (N12069, N12057, N2965, N9128, N1827);
nor NOR3 (N12070, N12063, N2530, N9810);
xor XOR2 (N12071, N12068, N1328);
nand NAND2 (N12072, N12014, N5728);
not NOT1 (N12073, N12061);
nand NAND4 (N12074, N12065, N10658, N1721, N1880);
nand NAND3 (N12075, N12070, N8228, N1453);
not NOT1 (N12076, N12071);
xor XOR2 (N12077, N12075, N3764);
or OR2 (N12078, N12058, N7584);
xor XOR2 (N12079, N12077, N6534);
nand NAND2 (N12080, N12078, N4100);
and AND2 (N12081, N12072, N3873);
nand NAND4 (N12082, N12069, N8555, N10821, N11932);
and AND2 (N12083, N12067, N10200);
or OR2 (N12084, N12082, N775);
not NOT1 (N12085, N12076);
and AND2 (N12086, N12055, N6034);
and AND4 (N12087, N12080, N2390, N3191, N500);
xor XOR2 (N12088, N12073, N9352);
and AND4 (N12089, N12049, N3165, N6282, N6454);
nand NAND3 (N12090, N12074, N6980, N2953);
nor NOR4 (N12091, N12079, N4144, N3245, N8114);
or OR2 (N12092, N12085, N8905);
xor XOR2 (N12093, N12089, N9321);
nor NOR3 (N12094, N12091, N11899, N3850);
and AND4 (N12095, N12092, N11334, N8626, N3555);
buf BUF1 (N12096, N12095);
nor NOR3 (N12097, N12084, N5304, N5930);
xor XOR2 (N12098, N12096, N3277);
not NOT1 (N12099, N12093);
buf BUF1 (N12100, N12088);
and AND2 (N12101, N12094, N11106);
xor XOR2 (N12102, N12087, N3787);
not NOT1 (N12103, N12100);
nor NOR3 (N12104, N12098, N164, N443);
buf BUF1 (N12105, N12104);
not NOT1 (N12106, N12097);
nand NAND4 (N12107, N12081, N6, N6633, N7474);
or OR2 (N12108, N12105, N3172);
xor XOR2 (N12109, N12090, N6226);
nor NOR3 (N12110, N12101, N8593, N1959);
or OR2 (N12111, N12110, N11638);
xor XOR2 (N12112, N12083, N10631);
and AND2 (N12113, N12102, N1258);
xor XOR2 (N12114, N12099, N9522);
or OR2 (N12115, N12108, N11585);
and AND4 (N12116, N12103, N800, N3154, N3955);
or OR3 (N12117, N12109, N6276, N1888);
buf BUF1 (N12118, N12107);
or OR3 (N12119, N12115, N12066, N8165);
xor XOR2 (N12120, N12111, N1632);
nand NAND4 (N12121, N12106, N9203, N9504, N10269);
xor XOR2 (N12122, N12117, N3123);
buf BUF1 (N12123, N12113);
buf BUF1 (N12124, N12120);
xor XOR2 (N12125, N12112, N5081);
nand NAND3 (N12126, N12123, N5147, N9864);
not NOT1 (N12127, N12121);
xor XOR2 (N12128, N12086, N4644);
or OR3 (N12129, N12125, N9851, N10570);
buf BUF1 (N12130, N12126);
nand NAND3 (N12131, N12119, N4726, N6808);
xor XOR2 (N12132, N12116, N3391);
nand NAND3 (N12133, N12118, N2230, N9414);
or OR4 (N12134, N12129, N5740, N6516, N3274);
or OR3 (N12135, N12127, N222, N6245);
xor XOR2 (N12136, N12135, N2912);
nand NAND3 (N12137, N12132, N3160, N1816);
and AND2 (N12138, N12133, N6006);
not NOT1 (N12139, N12114);
or OR4 (N12140, N12124, N9763, N9593, N9924);
xor XOR2 (N12141, N12130, N1470);
nor NOR4 (N12142, N12138, N8008, N4720, N12003);
xor XOR2 (N12143, N12139, N9913);
buf BUF1 (N12144, N12134);
not NOT1 (N12145, N12144);
nor NOR4 (N12146, N12131, N3584, N5863, N2280);
not NOT1 (N12147, N12146);
or OR3 (N12148, N12145, N3242, N1444);
xor XOR2 (N12149, N12142, N5523);
and AND4 (N12150, N12148, N5667, N1692, N85);
nand NAND2 (N12151, N12147, N145);
nor NOR4 (N12152, N12141, N10283, N5197, N11159);
or OR2 (N12153, N12128, N3827);
or OR3 (N12154, N12153, N9288, N11429);
or OR4 (N12155, N12143, N8061, N11616, N5219);
not NOT1 (N12156, N12151);
nand NAND4 (N12157, N12152, N3972, N566, N10385);
nor NOR4 (N12158, N12155, N11298, N10423, N10503);
not NOT1 (N12159, N12136);
nand NAND3 (N12160, N12122, N10970, N164);
xor XOR2 (N12161, N12140, N10060);
or OR4 (N12162, N12137, N137, N6593, N5404);
or OR4 (N12163, N12159, N9403, N8173, N9880);
or OR3 (N12164, N12158, N8975, N3760);
not NOT1 (N12165, N12150);
buf BUF1 (N12166, N12162);
xor XOR2 (N12167, N12154, N1260);
buf BUF1 (N12168, N12156);
xor XOR2 (N12169, N12161, N483);
nor NOR4 (N12170, N12149, N9383, N8840, N479);
nand NAND4 (N12171, N12157, N2409, N11104, N1089);
xor XOR2 (N12172, N12165, N8208);
xor XOR2 (N12173, N12166, N9172);
or OR2 (N12174, N12160, N2876);
not NOT1 (N12175, N12163);
buf BUF1 (N12176, N12172);
nor NOR4 (N12177, N12170, N5272, N6830, N11211);
nor NOR2 (N12178, N12168, N7908);
or OR2 (N12179, N12164, N7538);
buf BUF1 (N12180, N12179);
or OR4 (N12181, N12175, N7917, N9859, N7415);
nor NOR3 (N12182, N12181, N318, N1885);
buf BUF1 (N12183, N12180);
and AND3 (N12184, N12171, N2869, N9494);
and AND3 (N12185, N12182, N3136, N11871);
and AND2 (N12186, N12167, N5062);
or OR2 (N12187, N12169, N8732);
and AND3 (N12188, N12183, N10520, N633);
not NOT1 (N12189, N12188);
or OR2 (N12190, N12173, N10602);
xor XOR2 (N12191, N12187, N3912);
nand NAND3 (N12192, N12174, N10793, N1538);
not NOT1 (N12193, N12176);
buf BUF1 (N12194, N12177);
and AND3 (N12195, N12193, N9151, N6796);
xor XOR2 (N12196, N12190, N5785);
nand NAND3 (N12197, N12196, N9741, N3069);
or OR4 (N12198, N12184, N4892, N7651, N9716);
not NOT1 (N12199, N12185);
nand NAND4 (N12200, N12186, N4828, N3895, N10617);
nor NOR4 (N12201, N12199, N361, N4434, N5918);
nand NAND4 (N12202, N12194, N6605, N5260, N8779);
nor NOR4 (N12203, N12200, N2070, N5950, N678);
and AND3 (N12204, N12202, N5506, N9206);
buf BUF1 (N12205, N12204);
not NOT1 (N12206, N12198);
or OR4 (N12207, N12197, N5210, N6585, N6567);
not NOT1 (N12208, N12203);
not NOT1 (N12209, N12205);
nand NAND3 (N12210, N12209, N9267, N5185);
nor NOR3 (N12211, N12191, N3394, N6466);
or OR3 (N12212, N12195, N8950, N9101);
and AND3 (N12213, N12189, N9336, N11907);
nor NOR4 (N12214, N12213, N9298, N208, N3037);
not NOT1 (N12215, N12212);
and AND4 (N12216, N12206, N2987, N8360, N7404);
nor NOR3 (N12217, N12192, N5021, N8001);
not NOT1 (N12218, N12210);
buf BUF1 (N12219, N12208);
and AND2 (N12220, N12217, N5812);
nor NOR2 (N12221, N12214, N1612);
and AND2 (N12222, N12218, N631);
not NOT1 (N12223, N12216);
nand NAND4 (N12224, N12178, N1537, N10167, N4655);
nand NAND3 (N12225, N12207, N7830, N6102);
nand NAND3 (N12226, N12222, N4693, N5156);
and AND3 (N12227, N12219, N650, N2570);
and AND2 (N12228, N12226, N3490);
xor XOR2 (N12229, N12211, N3631);
not NOT1 (N12230, N12221);
and AND4 (N12231, N12228, N7112, N5828, N10615);
nor NOR2 (N12232, N12230, N479);
or OR3 (N12233, N12223, N10495, N10554);
not NOT1 (N12234, N12225);
nand NAND2 (N12235, N12234, N39);
nor NOR3 (N12236, N12231, N10690, N4171);
and AND2 (N12237, N12201, N5421);
buf BUF1 (N12238, N12233);
or OR4 (N12239, N12229, N9736, N10183, N1271);
xor XOR2 (N12240, N12236, N3949);
not NOT1 (N12241, N12237);
xor XOR2 (N12242, N12220, N7901);
and AND2 (N12243, N12235, N12045);
nand NAND2 (N12244, N12215, N1354);
xor XOR2 (N12245, N12244, N434);
not NOT1 (N12246, N12224);
nand NAND4 (N12247, N12227, N3341, N9481, N6973);
xor XOR2 (N12248, N12239, N10973);
xor XOR2 (N12249, N12240, N8922);
not NOT1 (N12250, N12248);
not NOT1 (N12251, N12250);
or OR4 (N12252, N12251, N5340, N10102, N5085);
nand NAND4 (N12253, N12247, N5623, N4482, N8634);
nor NOR4 (N12254, N12238, N2469, N9676, N5646);
buf BUF1 (N12255, N12242);
nor NOR4 (N12256, N12246, N9574, N5703, N1779);
or OR3 (N12257, N12243, N5188, N5724);
nand NAND4 (N12258, N12249, N2524, N4403, N2529);
not NOT1 (N12259, N12256);
or OR3 (N12260, N12258, N315, N7885);
nand NAND4 (N12261, N12254, N11148, N6831, N11523);
or OR2 (N12262, N12253, N8243);
nand NAND2 (N12263, N12260, N11929);
or OR4 (N12264, N12262, N5083, N7535, N2009);
buf BUF1 (N12265, N12252);
or OR2 (N12266, N12263, N6586);
and AND4 (N12267, N12245, N9511, N4951, N4761);
not NOT1 (N12268, N12265);
nand NAND3 (N12269, N12232, N8092, N563);
not NOT1 (N12270, N12266);
buf BUF1 (N12271, N12270);
nand NAND4 (N12272, N12268, N6775, N5059, N10476);
nand NAND2 (N12273, N12241, N384);
not NOT1 (N12274, N12264);
nand NAND3 (N12275, N12259, N345, N11376);
xor XOR2 (N12276, N12255, N2672);
nor NOR2 (N12277, N12257, N2990);
and AND4 (N12278, N12275, N8837, N2755, N2474);
nor NOR2 (N12279, N12278, N10317);
buf BUF1 (N12280, N12272);
and AND2 (N12281, N12273, N4251);
not NOT1 (N12282, N12279);
and AND3 (N12283, N12277, N8659, N2664);
not NOT1 (N12284, N12281);
not NOT1 (N12285, N12274);
and AND4 (N12286, N12285, N8683, N4536, N11607);
buf BUF1 (N12287, N12280);
and AND4 (N12288, N12267, N1524, N10176, N6128);
or OR2 (N12289, N12276, N6701);
nor NOR3 (N12290, N12286, N4309, N9758);
xor XOR2 (N12291, N12261, N1442);
xor XOR2 (N12292, N12269, N907);
or OR4 (N12293, N12289, N3111, N4460, N11940);
and AND4 (N12294, N12292, N3945, N5433, N6219);
and AND4 (N12295, N12291, N2846, N8705, N9770);
or OR3 (N12296, N12295, N2784, N5999);
and AND2 (N12297, N12290, N11963);
not NOT1 (N12298, N12287);
nor NOR3 (N12299, N12294, N1647, N933);
or OR4 (N12300, N12288, N4604, N7784, N10064);
or OR4 (N12301, N12271, N3762, N2540, N8347);
nor NOR3 (N12302, N12283, N7917, N3018);
buf BUF1 (N12303, N12284);
nor NOR3 (N12304, N12293, N4602, N435);
nand NAND3 (N12305, N12302, N11838, N2516);
xor XOR2 (N12306, N12297, N10022);
nor NOR2 (N12307, N12299, N7633);
or OR3 (N12308, N12296, N9326, N2271);
nand NAND2 (N12309, N12306, N2528);
xor XOR2 (N12310, N12304, N3611);
nor NOR2 (N12311, N12305, N2908);
and AND2 (N12312, N12311, N489);
nor NOR2 (N12313, N12307, N7804);
and AND4 (N12314, N12308, N2449, N10815, N9140);
and AND4 (N12315, N12309, N9544, N7404, N4052);
nor NOR2 (N12316, N12315, N2792);
nand NAND4 (N12317, N12301, N9107, N2320, N9658);
not NOT1 (N12318, N12313);
nor NOR3 (N12319, N12310, N9592, N1350);
buf BUF1 (N12320, N12314);
buf BUF1 (N12321, N12303);
nor NOR2 (N12322, N12312, N11560);
or OR4 (N12323, N12321, N6849, N4616, N2365);
or OR3 (N12324, N12316, N8698, N10192);
xor XOR2 (N12325, N12322, N3371);
and AND4 (N12326, N12298, N11795, N11113, N4716);
xor XOR2 (N12327, N12300, N10698);
nand NAND4 (N12328, N12325, N9075, N11606, N6790);
not NOT1 (N12329, N12317);
and AND2 (N12330, N12328, N4900);
not NOT1 (N12331, N12318);
not NOT1 (N12332, N12326);
xor XOR2 (N12333, N12323, N4988);
not NOT1 (N12334, N12324);
and AND2 (N12335, N12329, N11384);
xor XOR2 (N12336, N12334, N9177);
not NOT1 (N12337, N12332);
xor XOR2 (N12338, N12319, N4825);
xor XOR2 (N12339, N12333, N8601);
not NOT1 (N12340, N12338);
nand NAND2 (N12341, N12337, N3151);
buf BUF1 (N12342, N12331);
buf BUF1 (N12343, N12341);
xor XOR2 (N12344, N12320, N10936);
and AND2 (N12345, N12282, N8909);
buf BUF1 (N12346, N12339);
and AND2 (N12347, N12330, N7277);
buf BUF1 (N12348, N12335);
or OR4 (N12349, N12327, N10532, N6193, N526);
and AND3 (N12350, N12340, N6772, N4951);
and AND2 (N12351, N12342, N8327);
buf BUF1 (N12352, N12343);
nor NOR2 (N12353, N12344, N11429);
not NOT1 (N12354, N12345);
nor NOR3 (N12355, N12350, N7677, N9165);
nand NAND4 (N12356, N12353, N2105, N11569, N995);
nor NOR4 (N12357, N12351, N5067, N10011, N7571);
or OR4 (N12358, N12346, N8782, N7693, N3558);
buf BUF1 (N12359, N12358);
nand NAND4 (N12360, N12359, N102, N10986, N10173);
nand NAND2 (N12361, N12349, N8095);
buf BUF1 (N12362, N12348);
buf BUF1 (N12363, N12347);
and AND2 (N12364, N12362, N10934);
or OR4 (N12365, N12356, N468, N8016, N820);
buf BUF1 (N12366, N12336);
and AND4 (N12367, N12357, N8692, N7192, N6369);
buf BUF1 (N12368, N12367);
not NOT1 (N12369, N12354);
nand NAND4 (N12370, N12360, N5277, N540, N3548);
buf BUF1 (N12371, N12370);
xor XOR2 (N12372, N12364, N3449);
or OR2 (N12373, N12369, N8333);
xor XOR2 (N12374, N12365, N4164);
and AND4 (N12375, N12355, N1536, N7165, N3988);
and AND2 (N12376, N12373, N11497);
buf BUF1 (N12377, N12374);
buf BUF1 (N12378, N12368);
or OR3 (N12379, N12377, N2939, N1262);
nand NAND4 (N12380, N12366, N3001, N2117, N2673);
or OR3 (N12381, N12380, N9715, N9608);
xor XOR2 (N12382, N12352, N5834);
not NOT1 (N12383, N12381);
xor XOR2 (N12384, N12382, N6041);
and AND3 (N12385, N12361, N4850, N2702);
and AND3 (N12386, N12363, N3970, N6141);
or OR3 (N12387, N12384, N9547, N5734);
or OR4 (N12388, N12375, N9512, N6228, N9001);
and AND4 (N12389, N12379, N9547, N5822, N3977);
nor NOR2 (N12390, N12378, N1475);
buf BUF1 (N12391, N12390);
buf BUF1 (N12392, N12391);
not NOT1 (N12393, N12376);
nor NOR3 (N12394, N12392, N875, N5805);
or OR3 (N12395, N12387, N2360, N9955);
xor XOR2 (N12396, N12388, N9173);
xor XOR2 (N12397, N12385, N6707);
and AND3 (N12398, N12395, N783, N11650);
nor NOR2 (N12399, N12372, N9034);
buf BUF1 (N12400, N12386);
nor NOR4 (N12401, N12399, N4189, N4560, N7572);
xor XOR2 (N12402, N12398, N3282);
and AND4 (N12403, N12397, N9172, N9596, N5619);
not NOT1 (N12404, N12371);
not NOT1 (N12405, N12403);
buf BUF1 (N12406, N12383);
nor NOR4 (N12407, N12393, N4308, N4233, N8852);
nor NOR4 (N12408, N12406, N6660, N10445, N3230);
not NOT1 (N12409, N12405);
nor NOR4 (N12410, N12394, N4643, N12313, N8971);
nor NOR4 (N12411, N12400, N10001, N10495, N891);
or OR3 (N12412, N12389, N787, N389);
buf BUF1 (N12413, N12412);
not NOT1 (N12414, N12404);
nand NAND2 (N12415, N12410, N5863);
xor XOR2 (N12416, N12409, N1430);
or OR2 (N12417, N12415, N992);
xor XOR2 (N12418, N12416, N11451);
buf BUF1 (N12419, N12413);
nand NAND2 (N12420, N12407, N10868);
and AND2 (N12421, N12401, N6538);
nor NOR3 (N12422, N12420, N5496, N2803);
and AND4 (N12423, N12408, N6737, N9977, N175);
nand NAND2 (N12424, N12411, N1774);
not NOT1 (N12425, N12421);
nand NAND3 (N12426, N12422, N474, N8760);
nand NAND3 (N12427, N12414, N3031, N8451);
nor NOR3 (N12428, N12427, N2746, N11924);
and AND3 (N12429, N12426, N3770, N8214);
nand NAND2 (N12430, N12396, N5354);
and AND2 (N12431, N12429, N6741);
nand NAND2 (N12432, N12424, N200);
xor XOR2 (N12433, N12432, N9712);
buf BUF1 (N12434, N12431);
xor XOR2 (N12435, N12425, N3939);
nor NOR2 (N12436, N12434, N10268);
xor XOR2 (N12437, N12428, N1156);
nor NOR2 (N12438, N12435, N9628);
nor NOR4 (N12439, N12438, N6433, N943, N11856);
and AND3 (N12440, N12417, N10897, N3803);
nand NAND3 (N12441, N12433, N2186, N8892);
xor XOR2 (N12442, N12418, N7417);
buf BUF1 (N12443, N12437);
and AND4 (N12444, N12440, N3746, N2958, N7061);
or OR2 (N12445, N12444, N4611);
not NOT1 (N12446, N12402);
nand NAND3 (N12447, N12445, N2770, N1410);
buf BUF1 (N12448, N12430);
and AND4 (N12449, N12443, N5599, N10332, N1832);
nand NAND4 (N12450, N12436, N5490, N11950, N3019);
and AND2 (N12451, N12423, N5924);
nand NAND2 (N12452, N12419, N320);
or OR3 (N12453, N12446, N11125, N6329);
nand NAND4 (N12454, N12453, N2466, N1383, N4452);
or OR4 (N12455, N12442, N4144, N3677, N403);
and AND2 (N12456, N12454, N6516);
nor NOR2 (N12457, N12451, N422);
nor NOR2 (N12458, N12439, N3980);
buf BUF1 (N12459, N12449);
not NOT1 (N12460, N12447);
buf BUF1 (N12461, N12452);
nand NAND3 (N12462, N12441, N9935, N8047);
not NOT1 (N12463, N12448);
xor XOR2 (N12464, N12462, N2258);
xor XOR2 (N12465, N12460, N11909);
not NOT1 (N12466, N12459);
nor NOR2 (N12467, N12457, N7386);
nor NOR4 (N12468, N12466, N8884, N8553, N2300);
buf BUF1 (N12469, N12455);
buf BUF1 (N12470, N12456);
not NOT1 (N12471, N12461);
xor XOR2 (N12472, N12469, N8823);
not NOT1 (N12473, N12471);
or OR2 (N12474, N12470, N6716);
nor NOR2 (N12475, N12474, N6086);
xor XOR2 (N12476, N12450, N10833);
xor XOR2 (N12477, N12473, N8436);
nand NAND4 (N12478, N12463, N1790, N3765, N1126);
buf BUF1 (N12479, N12477);
buf BUF1 (N12480, N12472);
and AND2 (N12481, N12467, N9476);
nand NAND3 (N12482, N12475, N2086, N11357);
or OR4 (N12483, N12482, N11505, N8335, N8368);
buf BUF1 (N12484, N12478);
not NOT1 (N12485, N12483);
or OR3 (N12486, N12484, N5023, N4061);
not NOT1 (N12487, N12480);
nor NOR4 (N12488, N12468, N2098, N8386, N726);
not NOT1 (N12489, N12479);
nor NOR2 (N12490, N12489, N3890);
or OR2 (N12491, N12485, N9097);
nand NAND4 (N12492, N12491, N11630, N10575, N830);
nor NOR2 (N12493, N12476, N9554);
nand NAND2 (N12494, N12493, N780);
and AND2 (N12495, N12490, N6123);
nand NAND2 (N12496, N12492, N8710);
nor NOR2 (N12497, N12488, N6605);
buf BUF1 (N12498, N12458);
or OR3 (N12499, N12498, N11390, N9423);
nor NOR3 (N12500, N12496, N5590, N7279);
or OR3 (N12501, N12495, N9451, N7077);
xor XOR2 (N12502, N12487, N378);
not NOT1 (N12503, N12500);
nor NOR4 (N12504, N12465, N6391, N7540, N128);
and AND3 (N12505, N12502, N5582, N11800);
and AND3 (N12506, N12504, N9917, N6467);
not NOT1 (N12507, N12506);
and AND2 (N12508, N12503, N6091);
xor XOR2 (N12509, N12464, N5846);
xor XOR2 (N12510, N12509, N2157);
and AND2 (N12511, N12501, N7498);
nor NOR4 (N12512, N12494, N3204, N4247, N11902);
xor XOR2 (N12513, N12499, N11883);
xor XOR2 (N12514, N12508, N8080);
nor NOR2 (N12515, N12486, N8434);
buf BUF1 (N12516, N12510);
or OR4 (N12517, N12512, N11319, N7562, N9252);
not NOT1 (N12518, N12505);
or OR3 (N12519, N12518, N7842, N2980);
xor XOR2 (N12520, N12513, N9077);
not NOT1 (N12521, N12515);
nor NOR2 (N12522, N12519, N5399);
buf BUF1 (N12523, N12521);
not NOT1 (N12524, N12514);
buf BUF1 (N12525, N12511);
and AND4 (N12526, N12525, N7777, N2356, N5355);
buf BUF1 (N12527, N12526);
nor NOR3 (N12528, N12497, N3882, N8111);
not NOT1 (N12529, N12516);
or OR2 (N12530, N12529, N4169);
buf BUF1 (N12531, N12530);
buf BUF1 (N12532, N12507);
or OR2 (N12533, N12523, N2600);
and AND2 (N12534, N12531, N11060);
xor XOR2 (N12535, N12517, N2428);
not NOT1 (N12536, N12532);
or OR2 (N12537, N12522, N292);
and AND4 (N12538, N12537, N7676, N4703, N1541);
buf BUF1 (N12539, N12520);
nand NAND4 (N12540, N12535, N3684, N1938, N5169);
and AND4 (N12541, N12536, N161, N2229, N12242);
buf BUF1 (N12542, N12533);
or OR4 (N12543, N12538, N2416, N11818, N5580);
or OR4 (N12544, N12539, N4709, N9291, N8190);
not NOT1 (N12545, N12543);
and AND4 (N12546, N12534, N6520, N12181, N6526);
and AND3 (N12547, N12544, N2616, N568);
or OR2 (N12548, N12541, N7606);
and AND4 (N12549, N12524, N2104, N3641, N6383);
nand NAND4 (N12550, N12545, N11248, N1281, N9882);
nand NAND3 (N12551, N12528, N4851, N8485);
buf BUF1 (N12552, N12546);
xor XOR2 (N12553, N12550, N6490);
nor NOR2 (N12554, N12542, N2488);
nor NOR3 (N12555, N12481, N5063, N6361);
or OR2 (N12556, N12553, N10762);
buf BUF1 (N12557, N12548);
nand NAND3 (N12558, N12527, N9638, N4769);
not NOT1 (N12559, N12555);
nand NAND3 (N12560, N12556, N2273, N11167);
nor NOR2 (N12561, N12551, N3433);
and AND4 (N12562, N12557, N3581, N9673, N11308);
not NOT1 (N12563, N12561);
xor XOR2 (N12564, N12547, N6801);
xor XOR2 (N12565, N12552, N5573);
not NOT1 (N12566, N12560);
and AND3 (N12567, N12562, N10659, N3863);
buf BUF1 (N12568, N12566);
or OR2 (N12569, N12565, N8480);
nor NOR4 (N12570, N12564, N3305, N6358, N4127);
xor XOR2 (N12571, N12569, N9632);
or OR2 (N12572, N12571, N4835);
xor XOR2 (N12573, N12567, N9635);
nand NAND4 (N12574, N12559, N8954, N3741, N11601);
and AND2 (N12575, N12549, N8558);
buf BUF1 (N12576, N12575);
and AND4 (N12577, N12572, N6509, N9936, N8797);
xor XOR2 (N12578, N12563, N1090);
xor XOR2 (N12579, N12554, N11962);
buf BUF1 (N12580, N12578);
nand NAND3 (N12581, N12579, N10231, N12080);
xor XOR2 (N12582, N12581, N3940);
buf BUF1 (N12583, N12576);
not NOT1 (N12584, N12583);
nand NAND2 (N12585, N12580, N3660);
not NOT1 (N12586, N12573);
nand NAND4 (N12587, N12558, N1969, N6620, N12399);
and AND4 (N12588, N12570, N8405, N4215, N6104);
nor NOR3 (N12589, N12568, N9523, N3409);
buf BUF1 (N12590, N12589);
buf BUF1 (N12591, N12582);
or OR4 (N12592, N12577, N2755, N91, N5858);
not NOT1 (N12593, N12587);
or OR4 (N12594, N12592, N2574, N2539, N10553);
buf BUF1 (N12595, N12574);
xor XOR2 (N12596, N12588, N3691);
or OR3 (N12597, N12590, N4164, N2460);
or OR3 (N12598, N12593, N9826, N1119);
or OR3 (N12599, N12594, N10220, N7326);
buf BUF1 (N12600, N12585);
nor NOR3 (N12601, N12540, N144, N8787);
xor XOR2 (N12602, N12597, N3582);
not NOT1 (N12603, N12596);
xor XOR2 (N12604, N12601, N190);
nor NOR2 (N12605, N12604, N2457);
nor NOR2 (N12606, N12602, N5494);
and AND4 (N12607, N12591, N10749, N11027, N856);
not NOT1 (N12608, N12600);
not NOT1 (N12609, N12608);
xor XOR2 (N12610, N12609, N2716);
buf BUF1 (N12611, N12584);
xor XOR2 (N12612, N12598, N10793);
not NOT1 (N12613, N12607);
not NOT1 (N12614, N12586);
nor NOR4 (N12615, N12611, N1582, N7322, N11766);
xor XOR2 (N12616, N12610, N4547);
nor NOR4 (N12617, N12595, N10013, N7841, N6528);
nand NAND3 (N12618, N12612, N3050, N7447);
nor NOR3 (N12619, N12599, N4001, N6421);
not NOT1 (N12620, N12619);
not NOT1 (N12621, N12606);
nand NAND2 (N12622, N12618, N2186);
nor NOR4 (N12623, N12615, N4633, N5402, N2893);
nor NOR3 (N12624, N12616, N2297, N10134);
xor XOR2 (N12625, N12621, N8315);
not NOT1 (N12626, N12605);
and AND3 (N12627, N12614, N9665, N967);
xor XOR2 (N12628, N12625, N7806);
nand NAND4 (N12629, N12613, N8951, N9401, N6630);
xor XOR2 (N12630, N12617, N1939);
xor XOR2 (N12631, N12628, N5972);
xor XOR2 (N12632, N12623, N8782);
nor NOR3 (N12633, N12630, N2061, N4659);
nor NOR3 (N12634, N12624, N3479, N2340);
buf BUF1 (N12635, N12632);
and AND3 (N12636, N12603, N8770, N6871);
nand NAND3 (N12637, N12633, N2293, N8837);
and AND2 (N12638, N12627, N2943);
xor XOR2 (N12639, N12626, N8998);
or OR2 (N12640, N12634, N5606);
xor XOR2 (N12641, N12637, N5561);
xor XOR2 (N12642, N12620, N2226);
nand NAND2 (N12643, N12638, N7787);
nand NAND4 (N12644, N12641, N4202, N10846, N10193);
xor XOR2 (N12645, N12631, N11833);
nand NAND2 (N12646, N12639, N6822);
or OR2 (N12647, N12640, N1335);
or OR3 (N12648, N12642, N6201, N1021);
not NOT1 (N12649, N12645);
xor XOR2 (N12650, N12649, N8585);
nand NAND2 (N12651, N12635, N6256);
or OR4 (N12652, N12651, N7103, N4976, N2122);
or OR4 (N12653, N12648, N1643, N498, N11678);
and AND4 (N12654, N12650, N5565, N243, N923);
or OR3 (N12655, N12622, N12283, N11281);
nor NOR4 (N12656, N12654, N3389, N557, N4346);
or OR2 (N12657, N12655, N3228);
or OR4 (N12658, N12653, N8783, N7036, N9906);
and AND2 (N12659, N12652, N7979);
not NOT1 (N12660, N12659);
xor XOR2 (N12661, N12646, N12313);
nand NAND3 (N12662, N12657, N8190, N5307);
nor NOR3 (N12663, N12643, N10526, N4483);
xor XOR2 (N12664, N12662, N10904);
nand NAND2 (N12665, N12663, N9564);
and AND3 (N12666, N12656, N5694, N12513);
and AND2 (N12667, N12636, N2000);
nand NAND3 (N12668, N12666, N11407, N9085);
and AND3 (N12669, N12664, N6407, N9584);
and AND4 (N12670, N12660, N7488, N5077, N1747);
and AND2 (N12671, N12644, N9208);
buf BUF1 (N12672, N12661);
nand NAND3 (N12673, N12629, N12018, N1357);
and AND3 (N12674, N12672, N1513, N8768);
and AND3 (N12675, N12674, N5533, N8242);
and AND3 (N12676, N12668, N11339, N2024);
buf BUF1 (N12677, N12647);
and AND4 (N12678, N12665, N1493, N6137, N11939);
xor XOR2 (N12679, N12670, N4125);
and AND3 (N12680, N12673, N6252, N5078);
buf BUF1 (N12681, N12680);
nor NOR4 (N12682, N12681, N706, N8723, N1263);
buf BUF1 (N12683, N12679);
not NOT1 (N12684, N12682);
xor XOR2 (N12685, N12676, N226);
xor XOR2 (N12686, N12677, N8554);
or OR3 (N12687, N12667, N8021, N11212);
or OR4 (N12688, N12685, N8100, N5921, N11047);
buf BUF1 (N12689, N12684);
not NOT1 (N12690, N12688);
or OR3 (N12691, N12675, N5663, N1913);
nor NOR2 (N12692, N12683, N3926);
and AND2 (N12693, N12689, N1267);
xor XOR2 (N12694, N12691, N3066);
nor NOR4 (N12695, N12671, N9198, N6158, N3628);
or OR3 (N12696, N12658, N5242, N4975);
or OR2 (N12697, N12693, N4742);
nand NAND2 (N12698, N12686, N11249);
buf BUF1 (N12699, N12690);
and AND2 (N12700, N12669, N7411);
nor NOR3 (N12701, N12678, N1334, N5210);
nand NAND4 (N12702, N12694, N11011, N6125, N1721);
nand NAND2 (N12703, N12702, N8956);
nor NOR2 (N12704, N12700, N2106);
and AND3 (N12705, N12704, N8829, N9882);
or OR3 (N12706, N12687, N9013, N3752);
or OR2 (N12707, N12695, N9055);
nand NAND2 (N12708, N12706, N9614);
nor NOR3 (N12709, N12692, N4301, N6276);
xor XOR2 (N12710, N12699, N7508);
not NOT1 (N12711, N12710);
nand NAND4 (N12712, N12703, N9676, N691, N1464);
nand NAND4 (N12713, N12697, N8370, N11239, N3160);
or OR4 (N12714, N12698, N9606, N12581, N12647);
xor XOR2 (N12715, N12711, N9430);
or OR2 (N12716, N12709, N6369);
xor XOR2 (N12717, N12713, N294);
buf BUF1 (N12718, N12705);
nor NOR2 (N12719, N12712, N7600);
and AND2 (N12720, N12715, N7577);
nand NAND4 (N12721, N12717, N1841, N11455, N4176);
or OR3 (N12722, N12720, N783, N1193);
or OR2 (N12723, N12721, N3086);
or OR3 (N12724, N12701, N248, N9402);
or OR2 (N12725, N12707, N3555);
not NOT1 (N12726, N12718);
buf BUF1 (N12727, N12723);
buf BUF1 (N12728, N12726);
and AND2 (N12729, N12724, N4846);
or OR4 (N12730, N12727, N10300, N4057, N4490);
not NOT1 (N12731, N12725);
buf BUF1 (N12732, N12719);
buf BUF1 (N12733, N12716);
not NOT1 (N12734, N12731);
buf BUF1 (N12735, N12696);
nand NAND4 (N12736, N12734, N3584, N2525, N2323);
nand NAND4 (N12737, N12736, N4476, N6998, N2974);
nand NAND3 (N12738, N12737, N6487, N42);
nor NOR4 (N12739, N12728, N3000, N5414, N11964);
buf BUF1 (N12740, N12735);
xor XOR2 (N12741, N12730, N6887);
nand NAND3 (N12742, N12738, N9138, N5623);
xor XOR2 (N12743, N12714, N8143);
nand NAND4 (N12744, N12743, N9571, N3809, N1282);
xor XOR2 (N12745, N12708, N7560);
xor XOR2 (N12746, N12729, N9921);
or OR2 (N12747, N12741, N8374);
not NOT1 (N12748, N12733);
buf BUF1 (N12749, N12744);
buf BUF1 (N12750, N12745);
and AND2 (N12751, N12732, N9268);
nand NAND4 (N12752, N12746, N8776, N12068, N3505);
nand NAND2 (N12753, N12739, N5132);
and AND2 (N12754, N12748, N6653);
and AND2 (N12755, N12754, N6644);
nor NOR3 (N12756, N12753, N9607, N8475);
and AND3 (N12757, N12749, N5912, N5445);
and AND4 (N12758, N12742, N10206, N8750, N6282);
xor XOR2 (N12759, N12756, N7159);
buf BUF1 (N12760, N12758);
or OR2 (N12761, N12752, N4300);
nand NAND3 (N12762, N12747, N6001, N6629);
buf BUF1 (N12763, N12762);
nor NOR3 (N12764, N12755, N4082, N4660);
or OR4 (N12765, N12763, N6602, N3057, N9962);
nor NOR3 (N12766, N12722, N5418, N5594);
or OR4 (N12767, N12759, N4103, N11120, N2145);
nand NAND3 (N12768, N12760, N6496, N10046);
and AND3 (N12769, N12761, N6978, N5291);
and AND2 (N12770, N12765, N7918);
nand NAND4 (N12771, N12768, N870, N1928, N10769);
or OR4 (N12772, N12740, N11595, N5978, N2140);
xor XOR2 (N12773, N12751, N4135);
nand NAND3 (N12774, N12750, N7485, N4668);
nand NAND3 (N12775, N12764, N10947, N753);
nand NAND3 (N12776, N12766, N1393, N2563);
and AND2 (N12777, N12776, N1177);
or OR3 (N12778, N12757, N8276, N4029);
or OR4 (N12779, N12773, N6189, N12243, N1016);
nor NOR2 (N12780, N12775, N6945);
nor NOR3 (N12781, N12779, N12145, N7201);
nand NAND4 (N12782, N12771, N9162, N4444, N1290);
xor XOR2 (N12783, N12767, N10814);
buf BUF1 (N12784, N12774);
xor XOR2 (N12785, N12780, N8733);
not NOT1 (N12786, N12782);
buf BUF1 (N12787, N12770);
buf BUF1 (N12788, N12778);
not NOT1 (N12789, N12783);
nand NAND4 (N12790, N12785, N8393, N6410, N2153);
buf BUF1 (N12791, N12786);
or OR3 (N12792, N12790, N12006, N5041);
or OR4 (N12793, N12777, N10993, N801, N3644);
nor NOR4 (N12794, N12784, N5990, N3361, N7555);
not NOT1 (N12795, N12794);
xor XOR2 (N12796, N12788, N623);
nor NOR2 (N12797, N12789, N4289);
buf BUF1 (N12798, N12781);
nand NAND4 (N12799, N12795, N1579, N296, N2333);
nand NAND3 (N12800, N12769, N7317, N5930);
not NOT1 (N12801, N12793);
xor XOR2 (N12802, N12797, N12022);
and AND3 (N12803, N12800, N9735, N8575);
buf BUF1 (N12804, N12787);
or OR3 (N12805, N12796, N353, N2525);
buf BUF1 (N12806, N12799);
nand NAND4 (N12807, N12772, N5456, N7516, N9082);
nand NAND2 (N12808, N12807, N3704);
or OR4 (N12809, N12806, N4658, N9499, N234);
or OR3 (N12810, N12798, N10234, N4853);
or OR3 (N12811, N12804, N6462, N4271);
not NOT1 (N12812, N12802);
not NOT1 (N12813, N12791);
and AND4 (N12814, N12792, N4201, N1321, N11248);
nand NAND3 (N12815, N12811, N3221, N10806);
xor XOR2 (N12816, N12813, N3704);
and AND2 (N12817, N12805, N3361);
not NOT1 (N12818, N12809);
nor NOR3 (N12819, N12818, N3834, N4867);
endmodule