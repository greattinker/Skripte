// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N1009,N1001,N1011,N1019,N1005,N1013,N1015,N1017,N998,N1020;

xor XOR2 (N21, N11, N19);
and AND3 (N22, N9, N12, N9);
nand NAND4 (N23, N10, N20, N3, N3);
nand NAND2 (N24, N11, N18);
and AND2 (N25, N16, N1);
not NOT1 (N26, N3);
not NOT1 (N27, N16);
nor NOR2 (N28, N25, N23);
buf BUF1 (N29, N18);
nor NOR2 (N30, N22, N9);
xor XOR2 (N31, N12, N16);
buf BUF1 (N32, N20);
nand NAND4 (N33, N15, N21, N21, N24);
not NOT1 (N34, N19);
nand NAND4 (N35, N31, N16, N9, N12);
nor NOR3 (N36, N15, N32, N30);
buf BUF1 (N37, N11);
nand NAND3 (N38, N21, N9, N6);
buf BUF1 (N39, N37);
buf BUF1 (N40, N39);
not NOT1 (N41, N35);
nand NAND4 (N42, N27, N3, N25, N30);
xor XOR2 (N43, N41, N37);
nand NAND3 (N44, N28, N10, N29);
and AND4 (N45, N6, N16, N37, N25);
or OR3 (N46, N34, N34, N2);
xor XOR2 (N47, N26, N46);
or OR4 (N48, N25, N44, N35, N2);
and AND4 (N49, N40, N1, N14, N2);
buf BUF1 (N50, N24);
not NOT1 (N51, N43);
xor XOR2 (N52, N33, N18);
xor XOR2 (N53, N49, N14);
nand NAND2 (N54, N51, N40);
xor XOR2 (N55, N52, N11);
and AND2 (N56, N47, N11);
buf BUF1 (N57, N56);
nand NAND3 (N58, N54, N12, N37);
nand NAND2 (N59, N45, N33);
nor NOR4 (N60, N48, N31, N58, N34);
or OR4 (N61, N53, N1, N25, N7);
or OR2 (N62, N22, N15);
buf BUF1 (N63, N62);
buf BUF1 (N64, N59);
not NOT1 (N65, N42);
buf BUF1 (N66, N65);
not NOT1 (N67, N36);
not NOT1 (N68, N67);
nand NAND2 (N69, N60, N28);
not NOT1 (N70, N38);
or OR4 (N71, N69, N47, N56, N67);
nand NAND4 (N72, N66, N26, N69, N64);
not NOT1 (N73, N49);
not NOT1 (N74, N70);
buf BUF1 (N75, N63);
or OR3 (N76, N74, N5, N53);
or OR4 (N77, N73, N12, N2, N46);
nor NOR4 (N78, N68, N26, N71, N41);
xor XOR2 (N79, N40, N11);
not NOT1 (N80, N76);
buf BUF1 (N81, N78);
not NOT1 (N82, N75);
buf BUF1 (N83, N81);
not NOT1 (N84, N80);
buf BUF1 (N85, N50);
or OR2 (N86, N57, N28);
or OR3 (N87, N86, N37, N51);
or OR4 (N88, N84, N80, N80, N63);
xor XOR2 (N89, N82, N69);
and AND2 (N90, N55, N40);
nor NOR3 (N91, N79, N65, N89);
xor XOR2 (N92, N46, N8);
nand NAND2 (N93, N77, N39);
xor XOR2 (N94, N88, N93);
nand NAND3 (N95, N22, N39, N20);
nor NOR2 (N96, N85, N33);
not NOT1 (N97, N90);
nor NOR3 (N98, N61, N11, N91);
xor XOR2 (N99, N24, N36);
buf BUF1 (N100, N94);
nand NAND2 (N101, N97, N84);
not NOT1 (N102, N100);
nand NAND4 (N103, N102, N24, N56, N78);
not NOT1 (N104, N95);
or OR4 (N105, N103, N65, N65, N101);
not NOT1 (N106, N64);
xor XOR2 (N107, N92, N105);
and AND4 (N108, N22, N46, N79, N16);
xor XOR2 (N109, N106, N81);
buf BUF1 (N110, N109);
not NOT1 (N111, N107);
and AND4 (N112, N110, N52, N90, N79);
not NOT1 (N113, N98);
nor NOR3 (N114, N108, N79, N56);
and AND4 (N115, N111, N9, N62, N83);
xor XOR2 (N116, N49, N13);
xor XOR2 (N117, N112, N81);
or OR4 (N118, N99, N65, N57, N26);
nor NOR4 (N119, N113, N116, N49, N13);
xor XOR2 (N120, N105, N82);
and AND2 (N121, N72, N25);
xor XOR2 (N122, N120, N79);
and AND2 (N123, N87, N88);
and AND4 (N124, N119, N95, N61, N31);
xor XOR2 (N125, N122, N78);
or OR4 (N126, N114, N107, N121, N11);
nor NOR2 (N127, N124, N126);
nor NOR2 (N128, N79, N34);
buf BUF1 (N129, N113);
nand NAND4 (N130, N117, N32, N127, N14);
xor XOR2 (N131, N44, N35);
buf BUF1 (N132, N128);
buf BUF1 (N133, N115);
nand NAND3 (N134, N133, N7, N31);
xor XOR2 (N135, N96, N100);
nor NOR4 (N136, N118, N105, N130, N67);
not NOT1 (N137, N49);
and AND4 (N138, N125, N86, N15, N109);
or OR3 (N139, N131, N45, N65);
buf BUF1 (N140, N139);
xor XOR2 (N141, N140, N55);
nor NOR4 (N142, N135, N58, N106, N31);
nor NOR4 (N143, N141, N113, N73, N112);
and AND3 (N144, N129, N143, N35);
xor XOR2 (N145, N51, N115);
not NOT1 (N146, N144);
nor NOR2 (N147, N142, N12);
buf BUF1 (N148, N104);
or OR3 (N149, N148, N30, N13);
not NOT1 (N150, N123);
nor NOR2 (N151, N137, N61);
buf BUF1 (N152, N150);
not NOT1 (N153, N138);
not NOT1 (N154, N136);
or OR4 (N155, N152, N108, N21, N74);
and AND3 (N156, N154, N8, N53);
buf BUF1 (N157, N146);
nor NOR3 (N158, N151, N143, N51);
buf BUF1 (N159, N156);
nand NAND3 (N160, N145, N73, N47);
not NOT1 (N161, N155);
buf BUF1 (N162, N159);
nand NAND2 (N163, N132, N84);
nand NAND3 (N164, N149, N52, N29);
not NOT1 (N165, N157);
and AND2 (N166, N162, N148);
and AND2 (N167, N165, N56);
buf BUF1 (N168, N166);
buf BUF1 (N169, N168);
nor NOR4 (N170, N158, N35, N62, N86);
or OR3 (N171, N167, N95, N67);
and AND4 (N172, N170, N89, N34, N29);
nand NAND2 (N173, N171, N159);
and AND3 (N174, N173, N81, N120);
not NOT1 (N175, N160);
xor XOR2 (N176, N172, N14);
xor XOR2 (N177, N164, N48);
not NOT1 (N178, N177);
nand NAND3 (N179, N147, N77, N48);
nor NOR4 (N180, N179, N174, N138, N76);
xor XOR2 (N181, N178, N15);
not NOT1 (N182, N171);
buf BUF1 (N183, N181);
xor XOR2 (N184, N169, N46);
not NOT1 (N185, N183);
nand NAND4 (N186, N185, N30, N43, N102);
or OR2 (N187, N176, N80);
not NOT1 (N188, N180);
buf BUF1 (N189, N134);
buf BUF1 (N190, N188);
not NOT1 (N191, N190);
xor XOR2 (N192, N191, N183);
xor XOR2 (N193, N189, N71);
nand NAND2 (N194, N153, N147);
buf BUF1 (N195, N193);
or OR3 (N196, N186, N6, N193);
buf BUF1 (N197, N182);
nor NOR3 (N198, N192, N184, N100);
buf BUF1 (N199, N133);
nand NAND2 (N200, N196, N77);
buf BUF1 (N201, N194);
or OR2 (N202, N197, N156);
and AND4 (N203, N199, N60, N116, N196);
and AND3 (N204, N198, N10, N193);
nor NOR2 (N205, N163, N68);
and AND4 (N206, N203, N129, N167, N42);
nand NAND4 (N207, N204, N61, N196, N35);
or OR3 (N208, N202, N59, N63);
buf BUF1 (N209, N205);
not NOT1 (N210, N208);
xor XOR2 (N211, N200, N199);
xor XOR2 (N212, N209, N106);
not NOT1 (N213, N175);
nor NOR3 (N214, N212, N12, N34);
xor XOR2 (N215, N206, N114);
buf BUF1 (N216, N201);
or OR2 (N217, N207, N95);
and AND4 (N218, N214, N140, N98, N6);
nor NOR4 (N219, N215, N15, N82, N168);
nand NAND4 (N220, N187, N152, N115, N53);
buf BUF1 (N221, N219);
nor NOR4 (N222, N216, N170, N15, N188);
nand NAND2 (N223, N211, N5);
nor NOR2 (N224, N195, N140);
and AND2 (N225, N213, N21);
nand NAND3 (N226, N210, N204, N3);
xor XOR2 (N227, N220, N58);
xor XOR2 (N228, N217, N108);
xor XOR2 (N229, N228, N210);
nand NAND4 (N230, N222, N47, N48, N52);
xor XOR2 (N231, N227, N186);
xor XOR2 (N232, N221, N47);
xor XOR2 (N233, N230, N25);
xor XOR2 (N234, N218, N20);
and AND3 (N235, N226, N16, N36);
nor NOR3 (N236, N232, N179, N115);
nand NAND2 (N237, N231, N66);
and AND2 (N238, N236, N196);
xor XOR2 (N239, N224, N187);
or OR3 (N240, N225, N199, N77);
or OR2 (N241, N229, N178);
xor XOR2 (N242, N233, N231);
nand NAND4 (N243, N237, N222, N75, N220);
buf BUF1 (N244, N161);
nor NOR2 (N245, N244, N181);
nand NAND3 (N246, N238, N101, N119);
and AND4 (N247, N240, N37, N47, N203);
or OR3 (N248, N245, N11, N28);
buf BUF1 (N249, N223);
or OR4 (N250, N235, N181, N101, N78);
xor XOR2 (N251, N248, N47);
nand NAND4 (N252, N239, N26, N241, N85);
not NOT1 (N253, N171);
xor XOR2 (N254, N252, N209);
and AND4 (N255, N254, N14, N90, N195);
buf BUF1 (N256, N243);
and AND4 (N257, N250, N32, N20, N138);
and AND3 (N258, N255, N48, N83);
nand NAND4 (N259, N246, N68, N133, N28);
or OR4 (N260, N234, N222, N70, N233);
not NOT1 (N261, N258);
buf BUF1 (N262, N249);
xor XOR2 (N263, N260, N7);
and AND3 (N264, N259, N95, N85);
or OR3 (N265, N257, N29, N16);
or OR3 (N266, N265, N87, N220);
nor NOR2 (N267, N264, N88);
xor XOR2 (N268, N261, N98);
or OR3 (N269, N268, N2, N19);
xor XOR2 (N270, N262, N174);
nor NOR4 (N271, N266, N9, N234, N204);
nand NAND2 (N272, N271, N177);
and AND4 (N273, N272, N241, N90, N80);
xor XOR2 (N274, N267, N253);
nor NOR3 (N275, N218, N70, N121);
and AND3 (N276, N269, N77, N81);
nand NAND3 (N277, N242, N266, N63);
not NOT1 (N278, N251);
not NOT1 (N279, N273);
buf BUF1 (N280, N277);
not NOT1 (N281, N280);
xor XOR2 (N282, N256, N17);
buf BUF1 (N283, N270);
nand NAND4 (N284, N274, N116, N176, N194);
buf BUF1 (N285, N278);
nor NOR2 (N286, N284, N80);
xor XOR2 (N287, N263, N199);
xor XOR2 (N288, N276, N270);
nand NAND4 (N289, N283, N21, N193, N176);
nor NOR3 (N290, N285, N53, N21);
not NOT1 (N291, N289);
and AND4 (N292, N275, N270, N2, N21);
xor XOR2 (N293, N291, N153);
or OR4 (N294, N286, N86, N157, N278);
nor NOR4 (N295, N293, N230, N250, N20);
not NOT1 (N296, N292);
xor XOR2 (N297, N247, N188);
buf BUF1 (N298, N295);
not NOT1 (N299, N297);
nor NOR4 (N300, N296, N62, N104, N229);
xor XOR2 (N301, N287, N175);
not NOT1 (N302, N294);
nand NAND2 (N303, N298, N183);
and AND4 (N304, N303, N287, N56, N133);
nand NAND4 (N305, N300, N263, N12, N119);
or OR4 (N306, N304, N263, N101, N177);
xor XOR2 (N307, N281, N245);
nor NOR4 (N308, N279, N149, N188, N232);
nor NOR3 (N309, N288, N239, N77);
and AND2 (N310, N302, N117);
xor XOR2 (N311, N308, N62);
or OR3 (N312, N299, N304, N220);
nand NAND3 (N313, N282, N220, N192);
nor NOR2 (N314, N312, N275);
not NOT1 (N315, N310);
nand NAND3 (N316, N307, N26, N154);
buf BUF1 (N317, N311);
xor XOR2 (N318, N305, N172);
not NOT1 (N319, N317);
buf BUF1 (N320, N316);
and AND3 (N321, N290, N235, N220);
or OR4 (N322, N314, N246, N164, N267);
nor NOR2 (N323, N318, N235);
and AND2 (N324, N322, N119);
or OR4 (N325, N306, N290, N279, N83);
nand NAND4 (N326, N309, N186, N278, N136);
nor NOR4 (N327, N321, N222, N121, N43);
nand NAND4 (N328, N326, N294, N171, N69);
or OR2 (N329, N313, N195);
buf BUF1 (N330, N319);
nand NAND4 (N331, N324, N192, N184, N259);
nor NOR4 (N332, N323, N89, N30, N171);
nor NOR2 (N333, N329, N293);
buf BUF1 (N334, N333);
nor NOR3 (N335, N332, N160, N136);
nand NAND3 (N336, N331, N320, N245);
buf BUF1 (N337, N251);
or OR3 (N338, N301, N13, N265);
nand NAND3 (N339, N328, N86, N268);
nor NOR2 (N340, N315, N26);
and AND3 (N341, N330, N281, N141);
buf BUF1 (N342, N325);
buf BUF1 (N343, N340);
xor XOR2 (N344, N341, N137);
or OR2 (N345, N334, N192);
and AND4 (N346, N339, N20, N138, N104);
nand NAND2 (N347, N336, N277);
nor NOR2 (N348, N342, N192);
nor NOR2 (N349, N344, N89);
not NOT1 (N350, N338);
not NOT1 (N351, N347);
and AND4 (N352, N350, N49, N328, N293);
xor XOR2 (N353, N345, N84);
buf BUF1 (N354, N348);
and AND2 (N355, N327, N84);
xor XOR2 (N356, N354, N329);
xor XOR2 (N357, N356, N81);
xor XOR2 (N358, N352, N90);
or OR3 (N359, N343, N48, N350);
and AND2 (N360, N358, N350);
buf BUF1 (N361, N337);
not NOT1 (N362, N349);
nand NAND3 (N363, N361, N155, N98);
nor NOR3 (N364, N357, N287, N259);
xor XOR2 (N365, N359, N132);
nor NOR3 (N366, N363, N99, N283);
buf BUF1 (N367, N346);
nor NOR3 (N368, N351, N11, N277);
or OR3 (N369, N335, N42, N356);
or OR3 (N370, N364, N13, N260);
xor XOR2 (N371, N353, N124);
not NOT1 (N372, N355);
or OR4 (N373, N372, N69, N354, N57);
nor NOR3 (N374, N371, N78, N179);
or OR4 (N375, N374, N226, N159, N231);
buf BUF1 (N376, N360);
nand NAND3 (N377, N375, N277, N91);
xor XOR2 (N378, N362, N187);
or OR3 (N379, N370, N140, N164);
nor NOR4 (N380, N378, N43, N278, N276);
buf BUF1 (N381, N379);
and AND4 (N382, N366, N308, N349, N120);
nand NAND3 (N383, N369, N378, N348);
nor NOR2 (N384, N377, N319);
nor NOR2 (N385, N382, N120);
not NOT1 (N386, N383);
xor XOR2 (N387, N367, N10);
xor XOR2 (N388, N368, N44);
xor XOR2 (N389, N386, N122);
nand NAND2 (N390, N373, N100);
nor NOR2 (N391, N384, N5);
xor XOR2 (N392, N389, N180);
buf BUF1 (N393, N365);
nor NOR3 (N394, N387, N196, N95);
and AND3 (N395, N376, N242, N36);
buf BUF1 (N396, N388);
nand NAND2 (N397, N395, N248);
nor NOR4 (N398, N396, N124, N318, N55);
nor NOR2 (N399, N381, N271);
and AND2 (N400, N393, N183);
or OR4 (N401, N398, N361, N221, N314);
nor NOR4 (N402, N397, N68, N304, N9);
and AND4 (N403, N394, N145, N144, N61);
xor XOR2 (N404, N380, N151);
nor NOR3 (N405, N390, N120, N189);
nor NOR3 (N406, N405, N281, N124);
nor NOR3 (N407, N402, N344, N153);
and AND4 (N408, N400, N353, N74, N168);
xor XOR2 (N409, N399, N226);
nand NAND2 (N410, N407, N99);
and AND4 (N411, N391, N200, N92, N196);
not NOT1 (N412, N409);
nand NAND4 (N413, N385, N2, N103, N284);
buf BUF1 (N414, N406);
xor XOR2 (N415, N410, N273);
nand NAND2 (N416, N403, N229);
xor XOR2 (N417, N392, N251);
nand NAND4 (N418, N404, N135, N63, N131);
buf BUF1 (N419, N418);
nand NAND4 (N420, N411, N383, N356, N263);
buf BUF1 (N421, N414);
or OR4 (N422, N412, N362, N32, N101);
nor NOR4 (N423, N421, N228, N107, N163);
or OR3 (N424, N423, N391, N157);
not NOT1 (N425, N422);
not NOT1 (N426, N417);
and AND3 (N427, N401, N307, N73);
nand NAND2 (N428, N425, N145);
xor XOR2 (N429, N420, N391);
or OR2 (N430, N424, N97);
buf BUF1 (N431, N408);
not NOT1 (N432, N415);
buf BUF1 (N433, N429);
not NOT1 (N434, N432);
nor NOR3 (N435, N416, N220, N291);
not NOT1 (N436, N426);
nand NAND4 (N437, N413, N436, N186, N227);
buf BUF1 (N438, N374);
xor XOR2 (N439, N430, N367);
nor NOR4 (N440, N439, N245, N370, N322);
buf BUF1 (N441, N435);
buf BUF1 (N442, N433);
not NOT1 (N443, N440);
xor XOR2 (N444, N443, N50);
not NOT1 (N445, N431);
and AND2 (N446, N444, N324);
nor NOR4 (N447, N441, N400, N213, N210);
or OR4 (N448, N442, N318, N14, N37);
and AND2 (N449, N427, N175);
nor NOR4 (N450, N437, N345, N43, N173);
nor NOR3 (N451, N434, N8, N322);
xor XOR2 (N452, N451, N242);
nand NAND3 (N453, N447, N306, N222);
or OR4 (N454, N438, N349, N413, N273);
nor NOR3 (N455, N454, N296, N177);
nand NAND4 (N456, N455, N132, N326, N84);
and AND4 (N457, N445, N339, N392, N138);
and AND3 (N458, N452, N296, N135);
nand NAND4 (N459, N450, N118, N258, N399);
nand NAND3 (N460, N457, N410, N436);
nor NOR3 (N461, N453, N32, N442);
not NOT1 (N462, N448);
not NOT1 (N463, N459);
buf BUF1 (N464, N460);
not NOT1 (N465, N419);
buf BUF1 (N466, N464);
buf BUF1 (N467, N461);
nand NAND3 (N468, N456, N221, N347);
and AND4 (N469, N466, N267, N437, N398);
nor NOR3 (N470, N458, N310, N461);
xor XOR2 (N471, N462, N118);
or OR4 (N472, N428, N337, N227, N400);
xor XOR2 (N473, N469, N327);
or OR3 (N474, N467, N252, N176);
buf BUF1 (N475, N446);
or OR2 (N476, N468, N237);
not NOT1 (N477, N474);
nand NAND2 (N478, N475, N283);
xor XOR2 (N479, N463, N125);
nand NAND4 (N480, N470, N190, N113, N13);
or OR3 (N481, N465, N338, N135);
and AND2 (N482, N481, N224);
nor NOR2 (N483, N449, N293);
xor XOR2 (N484, N478, N46);
not NOT1 (N485, N484);
xor XOR2 (N486, N485, N57);
or OR4 (N487, N483, N298, N460, N45);
nor NOR4 (N488, N471, N62, N211, N251);
nor NOR2 (N489, N480, N389);
xor XOR2 (N490, N479, N449);
and AND2 (N491, N482, N133);
nor NOR4 (N492, N472, N383, N159, N121);
xor XOR2 (N493, N490, N148);
or OR4 (N494, N489, N72, N123, N150);
not NOT1 (N495, N494);
not NOT1 (N496, N476);
not NOT1 (N497, N477);
xor XOR2 (N498, N491, N380);
buf BUF1 (N499, N495);
and AND3 (N500, N492, N170, N101);
not NOT1 (N501, N493);
not NOT1 (N502, N498);
not NOT1 (N503, N473);
and AND4 (N504, N497, N137, N361, N239);
not NOT1 (N505, N504);
buf BUF1 (N506, N496);
and AND2 (N507, N506, N459);
not NOT1 (N508, N501);
not NOT1 (N509, N500);
or OR2 (N510, N486, N141);
nor NOR4 (N511, N509, N228, N506, N461);
or OR2 (N512, N499, N356);
nand NAND3 (N513, N507, N418, N368);
or OR4 (N514, N505, N130, N369, N245);
buf BUF1 (N515, N513);
buf BUF1 (N516, N502);
xor XOR2 (N517, N512, N57);
not NOT1 (N518, N487);
nor NOR3 (N519, N518, N151, N506);
not NOT1 (N520, N508);
and AND4 (N521, N517, N252, N45, N349);
not NOT1 (N522, N514);
not NOT1 (N523, N516);
or OR2 (N524, N511, N304);
xor XOR2 (N525, N519, N25);
xor XOR2 (N526, N510, N99);
and AND4 (N527, N526, N123, N420, N415);
xor XOR2 (N528, N503, N250);
or OR2 (N529, N515, N175);
or OR4 (N530, N521, N124, N29, N492);
not NOT1 (N531, N522);
not NOT1 (N532, N520);
nor NOR3 (N533, N530, N469, N113);
nand NAND4 (N534, N533, N358, N429, N128);
xor XOR2 (N535, N524, N113);
nor NOR3 (N536, N528, N200, N473);
and AND4 (N537, N488, N10, N509, N500);
not NOT1 (N538, N535);
not NOT1 (N539, N537);
xor XOR2 (N540, N531, N55);
not NOT1 (N541, N538);
nand NAND2 (N542, N527, N281);
not NOT1 (N543, N525);
not NOT1 (N544, N523);
or OR4 (N545, N536, N298, N242, N42);
not NOT1 (N546, N540);
nand NAND2 (N547, N542, N444);
nand NAND3 (N548, N529, N59, N318);
nor NOR4 (N549, N543, N336, N39, N32);
nor NOR3 (N550, N544, N312, N500);
nand NAND2 (N551, N550, N465);
not NOT1 (N552, N547);
xor XOR2 (N553, N549, N548);
and AND2 (N554, N291, N46);
not NOT1 (N555, N554);
or OR2 (N556, N539, N304);
buf BUF1 (N557, N555);
or OR4 (N558, N541, N160, N227, N68);
or OR2 (N559, N545, N119);
not NOT1 (N560, N551);
or OR2 (N561, N552, N275);
and AND2 (N562, N553, N424);
not NOT1 (N563, N532);
buf BUF1 (N564, N534);
and AND4 (N565, N546, N121, N405, N241);
and AND3 (N566, N556, N521, N480);
xor XOR2 (N567, N565, N498);
xor XOR2 (N568, N562, N281);
and AND3 (N569, N558, N522, N223);
nand NAND2 (N570, N560, N322);
and AND3 (N571, N566, N366, N217);
nor NOR3 (N572, N557, N451, N428);
nor NOR2 (N573, N572, N70);
xor XOR2 (N574, N571, N202);
or OR4 (N575, N564, N379, N385, N150);
xor XOR2 (N576, N561, N562);
or OR3 (N577, N576, N469, N38);
buf BUF1 (N578, N563);
nand NAND2 (N579, N578, N336);
nor NOR3 (N580, N568, N20, N302);
nand NAND2 (N581, N580, N406);
nand NAND4 (N582, N559, N365, N226, N547);
nand NAND4 (N583, N577, N484, N67, N334);
nor NOR2 (N584, N570, N185);
and AND2 (N585, N579, N533);
or OR4 (N586, N573, N221, N447, N440);
and AND4 (N587, N582, N135, N219, N88);
nand NAND4 (N588, N581, N582, N460, N527);
not NOT1 (N589, N588);
and AND4 (N590, N575, N270, N424, N302);
not NOT1 (N591, N586);
not NOT1 (N592, N590);
buf BUF1 (N593, N585);
xor XOR2 (N594, N584, N102);
and AND3 (N595, N593, N179, N253);
nand NAND3 (N596, N569, N559, N53);
nor NOR2 (N597, N591, N86);
nand NAND2 (N598, N594, N84);
buf BUF1 (N599, N592);
or OR3 (N600, N587, N260, N32);
and AND3 (N601, N596, N141, N291);
and AND4 (N602, N583, N571, N227, N495);
or OR4 (N603, N574, N549, N323, N118);
xor XOR2 (N604, N595, N516);
and AND3 (N605, N604, N283, N513);
not NOT1 (N606, N600);
or OR4 (N607, N603, N372, N126, N494);
not NOT1 (N608, N605);
nor NOR4 (N609, N598, N233, N7, N591);
xor XOR2 (N610, N602, N131);
nor NOR2 (N611, N589, N179);
or OR2 (N612, N607, N337);
buf BUF1 (N613, N610);
not NOT1 (N614, N606);
buf BUF1 (N615, N613);
and AND2 (N616, N608, N160);
nand NAND4 (N617, N567, N359, N230, N604);
not NOT1 (N618, N597);
not NOT1 (N619, N616);
or OR3 (N620, N611, N65, N264);
or OR2 (N621, N618, N619);
nor NOR2 (N622, N433, N481);
buf BUF1 (N623, N617);
not NOT1 (N624, N623);
not NOT1 (N625, N621);
xor XOR2 (N626, N615, N424);
and AND3 (N627, N609, N482, N507);
nor NOR2 (N628, N601, N419);
not NOT1 (N629, N626);
nand NAND4 (N630, N614, N314, N380, N326);
or OR3 (N631, N599, N77, N91);
buf BUF1 (N632, N629);
nor NOR4 (N633, N612, N10, N446, N6);
not NOT1 (N634, N624);
or OR2 (N635, N627, N467);
and AND4 (N636, N630, N120, N282, N119);
and AND4 (N637, N631, N302, N46, N350);
not NOT1 (N638, N628);
or OR3 (N639, N636, N209, N168);
nand NAND4 (N640, N632, N416, N169, N551);
and AND4 (N641, N638, N633, N268, N391);
and AND3 (N642, N614, N513, N408);
and AND2 (N643, N642, N205);
or OR4 (N644, N635, N392, N374, N370);
or OR4 (N645, N639, N266, N614, N345);
not NOT1 (N646, N622);
buf BUF1 (N647, N641);
not NOT1 (N648, N620);
nand NAND4 (N649, N643, N244, N331, N354);
xor XOR2 (N650, N644, N196);
or OR3 (N651, N646, N15, N605);
or OR2 (N652, N650, N530);
xor XOR2 (N653, N651, N213);
not NOT1 (N654, N645);
nand NAND2 (N655, N634, N55);
nor NOR2 (N656, N649, N335);
or OR3 (N657, N656, N180, N355);
or OR3 (N658, N647, N235, N572);
nor NOR3 (N659, N648, N151, N268);
or OR4 (N660, N654, N395, N289, N341);
and AND2 (N661, N657, N445);
buf BUF1 (N662, N640);
and AND2 (N663, N653, N63);
nand NAND3 (N664, N637, N610, N274);
not NOT1 (N665, N625);
nand NAND3 (N666, N665, N456, N277);
or OR4 (N667, N663, N1, N6, N291);
nor NOR3 (N668, N667, N566, N176);
not NOT1 (N669, N661);
buf BUF1 (N670, N666);
nand NAND4 (N671, N659, N361, N643, N279);
and AND3 (N672, N660, N570, N75);
nand NAND3 (N673, N658, N161, N228);
nand NAND4 (N674, N652, N378, N611, N473);
nor NOR3 (N675, N674, N282, N340);
xor XOR2 (N676, N675, N420);
xor XOR2 (N677, N672, N469);
buf BUF1 (N678, N655);
and AND3 (N679, N676, N455, N268);
and AND4 (N680, N671, N142, N94, N336);
xor XOR2 (N681, N670, N544);
not NOT1 (N682, N679);
not NOT1 (N683, N662);
and AND2 (N684, N664, N26);
or OR4 (N685, N684, N254, N664, N193);
not NOT1 (N686, N673);
and AND4 (N687, N669, N135, N272, N25);
and AND2 (N688, N680, N149);
buf BUF1 (N689, N681);
xor XOR2 (N690, N668, N456);
nand NAND2 (N691, N683, N475);
nor NOR2 (N692, N687, N544);
nand NAND4 (N693, N689, N340, N30, N572);
or OR3 (N694, N677, N499, N359);
or OR2 (N695, N693, N325);
nor NOR4 (N696, N688, N494, N590, N409);
not NOT1 (N697, N690);
xor XOR2 (N698, N691, N322);
buf BUF1 (N699, N697);
or OR2 (N700, N699, N315);
or OR3 (N701, N694, N570, N549);
nand NAND3 (N702, N678, N662, N514);
or OR4 (N703, N701, N631, N307, N348);
nor NOR4 (N704, N703, N92, N232, N8);
not NOT1 (N705, N692);
or OR3 (N706, N696, N544, N69);
and AND2 (N707, N686, N463);
not NOT1 (N708, N706);
not NOT1 (N709, N698);
xor XOR2 (N710, N700, N654);
and AND2 (N711, N709, N597);
buf BUF1 (N712, N711);
not NOT1 (N713, N682);
xor XOR2 (N714, N712, N380);
nand NAND2 (N715, N710, N479);
and AND4 (N716, N713, N47, N674, N587);
or OR3 (N717, N685, N608, N160);
xor XOR2 (N718, N702, N187);
nor NOR2 (N719, N715, N609);
nor NOR2 (N720, N708, N642);
or OR2 (N721, N717, N201);
xor XOR2 (N722, N714, N231);
nor NOR4 (N723, N722, N684, N663, N582);
nor NOR4 (N724, N718, N365, N221, N216);
and AND2 (N725, N695, N231);
nand NAND3 (N726, N721, N578, N665);
buf BUF1 (N727, N723);
and AND2 (N728, N716, N258);
and AND4 (N729, N707, N466, N307, N148);
buf BUF1 (N730, N726);
nand NAND4 (N731, N724, N335, N426, N412);
and AND2 (N732, N729, N605);
nor NOR2 (N733, N728, N375);
not NOT1 (N734, N727);
or OR2 (N735, N725, N487);
nand NAND2 (N736, N731, N91);
and AND2 (N737, N730, N729);
nor NOR4 (N738, N737, N209, N236, N376);
xor XOR2 (N739, N719, N650);
or OR3 (N740, N734, N493, N432);
not NOT1 (N741, N720);
nand NAND2 (N742, N738, N310);
buf BUF1 (N743, N733);
or OR3 (N744, N742, N451, N681);
xor XOR2 (N745, N739, N300);
not NOT1 (N746, N736);
not NOT1 (N747, N705);
or OR3 (N748, N744, N309, N177);
or OR3 (N749, N741, N287, N653);
or OR2 (N750, N704, N134);
or OR3 (N751, N745, N198, N209);
nand NAND2 (N752, N748, N694);
and AND3 (N753, N747, N136, N438);
or OR2 (N754, N740, N376);
xor XOR2 (N755, N751, N622);
buf BUF1 (N756, N746);
and AND4 (N757, N735, N419, N48, N165);
xor XOR2 (N758, N756, N157);
xor XOR2 (N759, N749, N450);
xor XOR2 (N760, N753, N72);
nand NAND4 (N761, N750, N592, N579, N60);
xor XOR2 (N762, N760, N617);
or OR3 (N763, N754, N273, N478);
or OR3 (N764, N743, N270, N727);
nand NAND2 (N765, N761, N136);
not NOT1 (N766, N765);
nor NOR3 (N767, N759, N576, N256);
xor XOR2 (N768, N752, N273);
nor NOR3 (N769, N764, N35, N12);
nand NAND3 (N770, N767, N311, N94);
or OR3 (N771, N732, N146, N389);
and AND2 (N772, N758, N768);
buf BUF1 (N773, N41);
nor NOR3 (N774, N769, N422, N505);
and AND4 (N775, N755, N367, N494, N101);
nand NAND2 (N776, N772, N553);
nand NAND4 (N777, N773, N415, N157, N650);
or OR4 (N778, N770, N338, N364, N524);
nor NOR2 (N779, N771, N635);
xor XOR2 (N780, N776, N421);
or OR2 (N781, N775, N775);
nor NOR3 (N782, N779, N219, N302);
xor XOR2 (N783, N782, N134);
buf BUF1 (N784, N777);
and AND3 (N785, N783, N272, N772);
buf BUF1 (N786, N766);
nand NAND2 (N787, N781, N322);
and AND4 (N788, N763, N600, N733, N52);
or OR2 (N789, N785, N144);
buf BUF1 (N790, N774);
not NOT1 (N791, N762);
not NOT1 (N792, N791);
and AND2 (N793, N789, N514);
not NOT1 (N794, N788);
xor XOR2 (N795, N778, N318);
and AND4 (N796, N790, N117, N654, N38);
nand NAND2 (N797, N787, N624);
or OR2 (N798, N792, N367);
and AND4 (N799, N757, N751, N599, N326);
xor XOR2 (N800, N780, N55);
buf BUF1 (N801, N784);
nor NOR2 (N802, N794, N268);
not NOT1 (N803, N800);
nand NAND2 (N804, N796, N413);
nor NOR3 (N805, N801, N45, N597);
xor XOR2 (N806, N795, N2);
or OR3 (N807, N799, N284, N695);
xor XOR2 (N808, N805, N236);
and AND4 (N809, N802, N33, N687, N575);
not NOT1 (N810, N809);
not NOT1 (N811, N806);
and AND3 (N812, N810, N363, N680);
nand NAND3 (N813, N804, N83, N717);
or OR2 (N814, N811, N243);
or OR2 (N815, N812, N291);
and AND3 (N816, N808, N762, N230);
nor NOR3 (N817, N814, N725, N65);
xor XOR2 (N818, N803, N311);
and AND4 (N819, N813, N281, N236, N641);
xor XOR2 (N820, N798, N382);
buf BUF1 (N821, N807);
nand NAND2 (N822, N797, N490);
xor XOR2 (N823, N816, N737);
xor XOR2 (N824, N820, N102);
xor XOR2 (N825, N823, N417);
nor NOR3 (N826, N821, N169, N460);
nor NOR3 (N827, N793, N543, N15);
nor NOR2 (N828, N786, N505);
not NOT1 (N829, N822);
nor NOR3 (N830, N818, N390, N829);
and AND4 (N831, N52, N735, N711, N798);
and AND3 (N832, N819, N105, N474);
buf BUF1 (N833, N830);
nor NOR4 (N834, N824, N360, N117, N617);
not NOT1 (N835, N825);
not NOT1 (N836, N815);
and AND2 (N837, N817, N609);
nand NAND3 (N838, N835, N85, N324);
and AND3 (N839, N837, N801, N282);
buf BUF1 (N840, N827);
buf BUF1 (N841, N839);
not NOT1 (N842, N826);
nand NAND3 (N843, N841, N322, N631);
not NOT1 (N844, N828);
nor NOR2 (N845, N831, N696);
xor XOR2 (N846, N843, N444);
xor XOR2 (N847, N846, N566);
nand NAND4 (N848, N833, N211, N83, N418);
buf BUF1 (N849, N848);
buf BUF1 (N850, N847);
xor XOR2 (N851, N850, N509);
nand NAND4 (N852, N834, N497, N669, N603);
not NOT1 (N853, N845);
nor NOR2 (N854, N832, N335);
and AND3 (N855, N852, N37, N533);
or OR3 (N856, N838, N853, N58);
xor XOR2 (N857, N569, N831);
not NOT1 (N858, N856);
not NOT1 (N859, N854);
nand NAND3 (N860, N844, N54, N513);
or OR3 (N861, N840, N539, N610);
buf BUF1 (N862, N860);
nand NAND4 (N863, N857, N33, N200, N499);
xor XOR2 (N864, N861, N571);
and AND4 (N865, N849, N734, N194, N668);
not NOT1 (N866, N858);
or OR2 (N867, N855, N586);
xor XOR2 (N868, N862, N592);
or OR3 (N869, N836, N638, N235);
or OR4 (N870, N866, N140, N146, N268);
nand NAND2 (N871, N870, N611);
not NOT1 (N872, N867);
buf BUF1 (N873, N842);
or OR2 (N874, N872, N690);
nor NOR3 (N875, N859, N669, N814);
or OR3 (N876, N863, N615, N487);
xor XOR2 (N877, N875, N138);
and AND3 (N878, N851, N436, N692);
xor XOR2 (N879, N873, N221);
buf BUF1 (N880, N864);
or OR3 (N881, N877, N244, N79);
xor XOR2 (N882, N865, N695);
or OR4 (N883, N868, N106, N465, N65);
buf BUF1 (N884, N879);
nand NAND4 (N885, N876, N805, N766, N119);
nor NOR3 (N886, N871, N161, N431);
nor NOR3 (N887, N883, N354, N44);
nand NAND3 (N888, N874, N834, N481);
buf BUF1 (N889, N882);
xor XOR2 (N890, N884, N777);
buf BUF1 (N891, N887);
buf BUF1 (N892, N881);
nand NAND2 (N893, N878, N149);
nand NAND2 (N894, N888, N349);
nand NAND3 (N895, N886, N132, N207);
or OR3 (N896, N885, N632, N199);
buf BUF1 (N897, N895);
buf BUF1 (N898, N894);
nand NAND2 (N899, N898, N468);
and AND2 (N900, N891, N792);
buf BUF1 (N901, N890);
xor XOR2 (N902, N900, N223);
and AND3 (N903, N892, N153, N545);
xor XOR2 (N904, N897, N249);
nor NOR3 (N905, N889, N787, N585);
nand NAND3 (N906, N893, N232, N148);
or OR3 (N907, N906, N744, N457);
nor NOR3 (N908, N903, N349, N591);
nand NAND3 (N909, N905, N562, N25);
and AND2 (N910, N902, N326);
nor NOR2 (N911, N910, N86);
or OR3 (N912, N901, N378, N629);
xor XOR2 (N913, N904, N683);
not NOT1 (N914, N908);
or OR3 (N915, N896, N132, N818);
nor NOR2 (N916, N899, N835);
nand NAND3 (N917, N911, N309, N912);
and AND3 (N918, N9, N625, N427);
nand NAND2 (N919, N869, N845);
nand NAND2 (N920, N919, N37);
not NOT1 (N921, N917);
nand NAND4 (N922, N915, N606, N74, N83);
nor NOR2 (N923, N916, N716);
and AND2 (N924, N921, N477);
nor NOR4 (N925, N918, N70, N657, N766);
nor NOR4 (N926, N920, N531, N665, N402);
not NOT1 (N927, N913);
xor XOR2 (N928, N914, N844);
xor XOR2 (N929, N923, N452);
and AND4 (N930, N924, N716, N69, N340);
xor XOR2 (N931, N926, N6);
or OR4 (N932, N928, N549, N712, N71);
buf BUF1 (N933, N929);
xor XOR2 (N934, N927, N10);
buf BUF1 (N935, N922);
nand NAND2 (N936, N933, N486);
nor NOR3 (N937, N935, N842, N105);
nor NOR3 (N938, N880, N913, N223);
and AND3 (N939, N937, N541, N901);
nor NOR2 (N940, N936, N430);
nand NAND4 (N941, N940, N717, N311, N469);
buf BUF1 (N942, N938);
xor XOR2 (N943, N907, N167);
nand NAND4 (N944, N941, N667, N349, N300);
and AND2 (N945, N943, N141);
nand NAND4 (N946, N931, N381, N934, N681);
or OR2 (N947, N618, N654);
not NOT1 (N948, N932);
or OR2 (N949, N925, N603);
buf BUF1 (N950, N949);
or OR2 (N951, N946, N279);
buf BUF1 (N952, N947);
and AND3 (N953, N942, N726, N492);
and AND4 (N954, N909, N178, N34, N203);
or OR3 (N955, N945, N939, N106);
and AND4 (N956, N557, N371, N205, N122);
not NOT1 (N957, N956);
not NOT1 (N958, N954);
or OR3 (N959, N950, N611, N857);
or OR4 (N960, N948, N815, N423, N311);
nor NOR2 (N961, N952, N700);
not NOT1 (N962, N959);
not NOT1 (N963, N944);
nor NOR2 (N964, N957, N811);
not NOT1 (N965, N963);
xor XOR2 (N966, N965, N615);
and AND2 (N967, N960, N363);
not NOT1 (N968, N930);
xor XOR2 (N969, N964, N335);
or OR4 (N970, N968, N831, N870, N665);
xor XOR2 (N971, N966, N173);
buf BUF1 (N972, N969);
nand NAND4 (N973, N962, N88, N13, N200);
nand NAND3 (N974, N970, N232, N832);
buf BUF1 (N975, N967);
not NOT1 (N976, N971);
buf BUF1 (N977, N976);
buf BUF1 (N978, N973);
buf BUF1 (N979, N972);
and AND3 (N980, N975, N693, N876);
nor NOR4 (N981, N979, N372, N28, N1);
not NOT1 (N982, N951);
buf BUF1 (N983, N977);
nor NOR2 (N984, N961, N476);
buf BUF1 (N985, N958);
and AND2 (N986, N978, N64);
nor NOR4 (N987, N955, N936, N708, N571);
buf BUF1 (N988, N985);
buf BUF1 (N989, N980);
nor NOR3 (N990, N974, N822, N425);
xor XOR2 (N991, N981, N749);
or OR3 (N992, N991, N174, N531);
nor NOR2 (N993, N992, N31);
or OR3 (N994, N953, N31, N897);
not NOT1 (N995, N993);
buf BUF1 (N996, N984);
and AND2 (N997, N996, N810);
nor NOR3 (N998, N997, N818, N345);
nor NOR3 (N999, N990, N323, N266);
not NOT1 (N1000, N988);
and AND3 (N1001, N982, N475, N489);
buf BUF1 (N1002, N995);
buf BUF1 (N1003, N983);
not NOT1 (N1004, N1000);
buf BUF1 (N1005, N986);
nor NOR3 (N1006, N987, N363, N66);
or OR2 (N1007, N989, N760);
nand NAND3 (N1008, N994, N382, N797);
nand NAND2 (N1009, N1007, N497);
or OR3 (N1010, N1003, N61, N631);
nor NOR2 (N1011, N1006, N852);
buf BUF1 (N1012, N1004);
buf BUF1 (N1013, N999);
xor XOR2 (N1014, N1008, N18);
or OR4 (N1015, N1014, N404, N468, N162);
and AND2 (N1016, N1010, N710);
nand NAND4 (N1017, N1002, N893, N74, N711);
nor NOR4 (N1018, N1012, N894, N809, N918);
and AND4 (N1019, N1016, N465, N605, N928);
buf BUF1 (N1020, N1018);
endmodule