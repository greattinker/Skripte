// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17;

output N115,N116,N111,N102,N106,N114,N108,N89,N109,N117;

not NOT1 (N18, N7);
or OR2 (N19, N10, N10);
xor XOR2 (N20, N3, N19);
and AND3 (N21, N5, N4, N8);
buf BUF1 (N22, N20);
xor XOR2 (N23, N15, N8);
nand NAND3 (N24, N5, N14, N21);
xor XOR2 (N25, N4, N18);
and AND2 (N26, N22, N21);
and AND4 (N27, N22, N17, N15, N26);
and AND3 (N28, N7, N7, N18);
and AND2 (N29, N20, N16);
buf BUF1 (N30, N6);
buf BUF1 (N31, N17);
nand NAND4 (N32, N27, N14, N31, N14);
nand NAND4 (N33, N3, N14, N17, N16);
and AND4 (N34, N15, N30, N16, N20);
nor NOR4 (N35, N20, N3, N6, N10);
nand NAND2 (N36, N35, N33);
not NOT1 (N37, N31);
xor XOR2 (N38, N20, N23);
and AND2 (N39, N38, N16);
and AND3 (N40, N27, N39, N5);
and AND4 (N41, N12, N20, N26, N29);
and AND4 (N42, N32, N34, N31, N31);
nor NOR2 (N43, N11, N24);
and AND4 (N44, N8, N29, N37, N10);
nor NOR2 (N45, N32, N31);
nand NAND4 (N46, N42, N32, N44, N38);
nand NAND3 (N47, N35, N19, N13);
not NOT1 (N48, N37);
xor XOR2 (N49, N48, N38);
or OR4 (N50, N46, N1, N41, N2);
xor XOR2 (N51, N13, N18);
buf BUF1 (N52, N50);
nand NAND2 (N53, N47, N50);
buf BUF1 (N54, N43);
nor NOR4 (N55, N28, N16, N11, N40);
xor XOR2 (N56, N43, N38);
buf BUF1 (N57, N45);
or OR4 (N58, N54, N31, N20, N32);
or OR3 (N59, N58, N41, N14);
or OR3 (N60, N56, N5, N6);
not NOT1 (N61, N49);
or OR3 (N62, N55, N59, N10);
or OR2 (N63, N1, N21);
nor NOR2 (N64, N53, N29);
nand NAND4 (N65, N36, N13, N12, N16);
not NOT1 (N66, N25);
nor NOR3 (N67, N57, N53, N5);
and AND4 (N68, N51, N15, N55, N12);
nand NAND2 (N69, N64, N29);
or OR3 (N70, N66, N19, N17);
not NOT1 (N71, N61);
or OR2 (N72, N68, N68);
and AND2 (N73, N67, N49);
or OR3 (N74, N60, N55, N62);
not NOT1 (N75, N40);
nor NOR3 (N76, N75, N42, N45);
nor NOR4 (N77, N74, N9, N73, N53);
not NOT1 (N78, N37);
xor XOR2 (N79, N70, N40);
or OR2 (N80, N72, N6);
or OR2 (N81, N69, N26);
or OR4 (N82, N80, N40, N34, N36);
or OR4 (N83, N77, N51, N11, N25);
and AND3 (N84, N83, N30, N15);
or OR2 (N85, N78, N65);
not NOT1 (N86, N4);
buf BUF1 (N87, N82);
or OR3 (N88, N81, N62, N27);
and AND4 (N89, N88, N60, N50, N71);
xor XOR2 (N90, N41, N49);
not NOT1 (N91, N85);
not NOT1 (N92, N79);
not NOT1 (N93, N86);
and AND2 (N94, N76, N50);
not NOT1 (N95, N94);
nand NAND3 (N96, N90, N28, N35);
or OR3 (N97, N96, N80, N18);
nor NOR4 (N98, N92, N82, N28, N21);
nor NOR2 (N99, N95, N81);
and AND3 (N100, N97, N31, N33);
xor XOR2 (N101, N63, N51);
nand NAND4 (N102, N91, N86, N44, N59);
buf BUF1 (N103, N52);
xor XOR2 (N104, N84, N33);
and AND3 (N105, N98, N68, N7);
nor NOR2 (N106, N101, N75);
xor XOR2 (N107, N100, N41);
not NOT1 (N108, N93);
xor XOR2 (N109, N107, N92);
not NOT1 (N110, N87);
or OR4 (N111, N105, N27, N52, N32);
and AND4 (N112, N103, N107, N84, N44);
not NOT1 (N113, N110);
xor XOR2 (N114, N104, N62);
and AND2 (N115, N113, N98);
not NOT1 (N116, N99);
and AND4 (N117, N112, N47, N60, N72);
endmodule