// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;

output N4019,N4014,N4012,N4017,N4005,N4007,N4018,N4013,N4016,N4020;

nor NOR2 (N21, N5, N15);
not NOT1 (N22, N21);
and AND2 (N23, N12, N2);
nand NAND3 (N24, N8, N16, N9);
and AND3 (N25, N9, N17, N14);
or OR3 (N26, N14, N25, N12);
nand NAND3 (N27, N14, N10, N25);
nand NAND2 (N28, N5, N10);
or OR3 (N29, N19, N11, N27);
xor XOR2 (N30, N7, N29);
buf BUF1 (N31, N3);
or OR2 (N32, N11, N1);
not NOT1 (N33, N6);
not NOT1 (N34, N33);
nor NOR4 (N35, N15, N8, N19, N21);
xor XOR2 (N36, N28, N22);
or OR4 (N37, N4, N33, N31, N19);
or OR4 (N38, N11, N13, N8, N17);
nand NAND4 (N39, N32, N21, N7, N9);
xor XOR2 (N40, N35, N18);
nand NAND4 (N41, N40, N10, N33, N25);
and AND4 (N42, N36, N2, N23, N17);
nor NOR4 (N43, N13, N32, N33, N6);
not NOT1 (N44, N43);
not NOT1 (N45, N26);
nand NAND4 (N46, N24, N2, N24, N20);
xor XOR2 (N47, N46, N2);
or OR2 (N48, N45, N43);
and AND3 (N49, N34, N26, N29);
and AND3 (N50, N39, N19, N44);
buf BUF1 (N51, N33);
nor NOR3 (N52, N30, N34, N22);
nand NAND4 (N53, N37, N10, N48, N52);
nand NAND3 (N54, N31, N44, N3);
or OR2 (N55, N27, N47);
and AND2 (N56, N18, N23);
buf BUF1 (N57, N53);
or OR4 (N58, N50, N30, N49, N26);
not NOT1 (N59, N45);
nor NOR3 (N60, N38, N6, N21);
nor NOR3 (N61, N56, N42, N57);
nand NAND2 (N62, N53, N37);
or OR3 (N63, N58, N6, N32);
not NOT1 (N64, N30);
buf BUF1 (N65, N59);
xor XOR2 (N66, N63, N17);
buf BUF1 (N67, N41);
buf BUF1 (N68, N67);
and AND2 (N69, N54, N32);
xor XOR2 (N70, N60, N9);
or OR3 (N71, N69, N43, N26);
not NOT1 (N72, N61);
nor NOR2 (N73, N64, N70);
buf BUF1 (N74, N71);
buf BUF1 (N75, N30);
and AND3 (N76, N74, N30, N17);
nand NAND4 (N77, N65, N12, N14, N55);
buf BUF1 (N78, N3);
nor NOR4 (N79, N77, N20, N64, N3);
buf BUF1 (N80, N78);
not NOT1 (N81, N62);
or OR4 (N82, N80, N46, N39, N52);
xor XOR2 (N83, N76, N13);
nor NOR2 (N84, N81, N11);
nand NAND4 (N85, N84, N84, N58, N35);
not NOT1 (N86, N68);
not NOT1 (N87, N75);
not NOT1 (N88, N73);
and AND3 (N89, N88, N57, N16);
nor NOR4 (N90, N82, N10, N55, N20);
not NOT1 (N91, N85);
not NOT1 (N92, N86);
and AND2 (N93, N72, N15);
or OR3 (N94, N93, N37, N64);
xor XOR2 (N95, N94, N46);
xor XOR2 (N96, N90, N86);
or OR4 (N97, N96, N89, N5, N7);
not NOT1 (N98, N25);
or OR4 (N99, N51, N72, N86, N17);
or OR4 (N100, N87, N37, N55, N76);
or OR2 (N101, N66, N69);
xor XOR2 (N102, N95, N70);
or OR4 (N103, N98, N39, N15, N69);
or OR2 (N104, N103, N63);
nor NOR3 (N105, N99, N53, N63);
nor NOR4 (N106, N102, N69, N75, N71);
not NOT1 (N107, N101);
buf BUF1 (N108, N79);
not NOT1 (N109, N97);
or OR4 (N110, N92, N21, N50, N24);
nand NAND2 (N111, N105, N41);
xor XOR2 (N112, N107, N53);
buf BUF1 (N113, N100);
not NOT1 (N114, N109);
and AND3 (N115, N110, N18, N21);
and AND3 (N116, N108, N17, N106);
not NOT1 (N117, N9);
buf BUF1 (N118, N83);
nor NOR4 (N119, N104, N64, N47, N90);
buf BUF1 (N120, N115);
xor XOR2 (N121, N117, N44);
or OR2 (N122, N114, N31);
xor XOR2 (N123, N121, N121);
buf BUF1 (N124, N119);
xor XOR2 (N125, N118, N110);
and AND3 (N126, N123, N19, N2);
not NOT1 (N127, N120);
nor NOR3 (N128, N126, N43, N69);
nor NOR3 (N129, N116, N90, N48);
buf BUF1 (N130, N113);
xor XOR2 (N131, N128, N129);
xor XOR2 (N132, N31, N116);
buf BUF1 (N133, N130);
nor NOR4 (N134, N111, N107, N118, N100);
nor NOR2 (N135, N133, N58);
nor NOR3 (N136, N131, N6, N55);
nand NAND2 (N137, N125, N4);
nor NOR2 (N138, N137, N17);
not NOT1 (N139, N124);
nand NAND2 (N140, N112, N36);
not NOT1 (N141, N138);
and AND2 (N142, N135, N29);
nand NAND3 (N143, N136, N132, N63);
xor XOR2 (N144, N58, N110);
and AND4 (N145, N91, N55, N60, N75);
not NOT1 (N146, N143);
xor XOR2 (N147, N134, N28);
xor XOR2 (N148, N127, N83);
not NOT1 (N149, N144);
nor NOR2 (N150, N147, N39);
nand NAND2 (N151, N122, N26);
or OR2 (N152, N150, N131);
and AND3 (N153, N141, N49, N99);
xor XOR2 (N154, N152, N32);
not NOT1 (N155, N140);
nor NOR3 (N156, N139, N125, N89);
not NOT1 (N157, N142);
or OR2 (N158, N157, N104);
not NOT1 (N159, N151);
buf BUF1 (N160, N153);
xor XOR2 (N161, N155, N144);
xor XOR2 (N162, N158, N10);
nor NOR2 (N163, N160, N107);
nor NOR3 (N164, N148, N134, N3);
and AND2 (N165, N163, N115);
nor NOR4 (N166, N149, N69, N162, N51);
buf BUF1 (N167, N61);
not NOT1 (N168, N145);
xor XOR2 (N169, N146, N167);
xor XOR2 (N170, N87, N33);
xor XOR2 (N171, N165, N155);
and AND4 (N172, N169, N149, N83, N41);
buf BUF1 (N173, N166);
nor NOR4 (N174, N164, N74, N131, N114);
and AND3 (N175, N170, N114, N153);
or OR4 (N176, N168, N93, N142, N21);
nor NOR4 (N177, N174, N31, N166, N119);
and AND3 (N178, N177, N19, N77);
or OR2 (N179, N178, N102);
nand NAND2 (N180, N159, N131);
xor XOR2 (N181, N175, N29);
nor NOR3 (N182, N179, N131, N129);
nand NAND3 (N183, N182, N153, N12);
not NOT1 (N184, N154);
or OR2 (N185, N171, N34);
or OR4 (N186, N183, N152, N171, N134);
xor XOR2 (N187, N176, N178);
nor NOR4 (N188, N184, N30, N103, N101);
and AND3 (N189, N180, N44, N108);
not NOT1 (N190, N181);
buf BUF1 (N191, N188);
nor NOR3 (N192, N156, N3, N129);
buf BUF1 (N193, N191);
buf BUF1 (N194, N189);
and AND2 (N195, N173, N104);
xor XOR2 (N196, N161, N144);
buf BUF1 (N197, N196);
nand NAND4 (N198, N187, N164, N146, N76);
nand NAND4 (N199, N190, N3, N25, N134);
not NOT1 (N200, N198);
nor NOR2 (N201, N195, N44);
xor XOR2 (N202, N194, N190);
or OR2 (N203, N186, N5);
and AND2 (N204, N200, N8);
and AND4 (N205, N193, N134, N4, N92);
not NOT1 (N206, N203);
or OR3 (N207, N201, N188, N65);
nand NAND2 (N208, N202, N154);
or OR3 (N209, N205, N72, N66);
not NOT1 (N210, N197);
xor XOR2 (N211, N208, N161);
not NOT1 (N212, N172);
nor NOR3 (N213, N209, N88, N121);
and AND3 (N214, N204, N190, N30);
not NOT1 (N215, N199);
not NOT1 (N216, N206);
buf BUF1 (N217, N210);
nor NOR4 (N218, N207, N152, N39, N98);
buf BUF1 (N219, N215);
nand NAND3 (N220, N185, N32, N28);
not NOT1 (N221, N213);
or OR2 (N222, N212, N211);
buf BUF1 (N223, N110);
xor XOR2 (N224, N219, N1);
or OR2 (N225, N214, N221);
and AND4 (N226, N67, N1, N157, N163);
nand NAND3 (N227, N226, N201, N204);
not NOT1 (N228, N220);
nand NAND4 (N229, N192, N3, N115, N18);
xor XOR2 (N230, N228, N131);
xor XOR2 (N231, N225, N188);
and AND4 (N232, N216, N66, N191, N227);
nor NOR2 (N233, N11, N226);
and AND2 (N234, N229, N24);
or OR3 (N235, N234, N178, N111);
xor XOR2 (N236, N224, N41);
not NOT1 (N237, N231);
not NOT1 (N238, N217);
and AND4 (N239, N232, N102, N206, N184);
nand NAND2 (N240, N233, N122);
buf BUF1 (N241, N236);
or OR2 (N242, N223, N40);
xor XOR2 (N243, N238, N177);
xor XOR2 (N244, N239, N1);
or OR3 (N245, N242, N180, N172);
and AND2 (N246, N240, N138);
buf BUF1 (N247, N218);
nand NAND3 (N248, N241, N131, N74);
nand NAND2 (N249, N237, N238);
buf BUF1 (N250, N246);
nor NOR2 (N251, N222, N110);
nand NAND3 (N252, N243, N169, N201);
not NOT1 (N253, N248);
nand NAND2 (N254, N249, N92);
nand NAND3 (N255, N230, N239, N52);
and AND2 (N256, N247, N75);
buf BUF1 (N257, N245);
or OR2 (N258, N253, N94);
and AND4 (N259, N250, N23, N77, N251);
or OR2 (N260, N57, N228);
and AND3 (N261, N260, N104, N222);
and AND4 (N262, N235, N12, N256, N175);
not NOT1 (N263, N208);
buf BUF1 (N264, N254);
nor NOR3 (N265, N259, N192, N240);
nor NOR2 (N266, N252, N123);
nor NOR2 (N267, N263, N147);
not NOT1 (N268, N255);
and AND4 (N269, N262, N124, N12, N162);
buf BUF1 (N270, N257);
nand NAND2 (N271, N244, N95);
or OR2 (N272, N270, N30);
nand NAND2 (N273, N266, N256);
or OR2 (N274, N269, N85);
not NOT1 (N275, N268);
xor XOR2 (N276, N275, N36);
xor XOR2 (N277, N271, N106);
buf BUF1 (N278, N277);
nor NOR2 (N279, N274, N151);
buf BUF1 (N280, N273);
nand NAND4 (N281, N280, N50, N218, N38);
and AND2 (N282, N272, N12);
and AND4 (N283, N267, N212, N2, N276);
nor NOR2 (N284, N86, N238);
buf BUF1 (N285, N264);
and AND4 (N286, N258, N137, N253, N187);
xor XOR2 (N287, N284, N262);
buf BUF1 (N288, N261);
buf BUF1 (N289, N285);
buf BUF1 (N290, N281);
nor NOR4 (N291, N282, N216, N143, N283);
or OR2 (N292, N236, N110);
and AND2 (N293, N290, N231);
nand NAND2 (N294, N292, N254);
nor NOR2 (N295, N286, N22);
nand NAND3 (N296, N265, N28, N144);
buf BUF1 (N297, N278);
buf BUF1 (N298, N291);
buf BUF1 (N299, N289);
or OR4 (N300, N295, N179, N6, N287);
nor NOR4 (N301, N75, N85, N267, N295);
buf BUF1 (N302, N300);
not NOT1 (N303, N279);
nor NOR4 (N304, N296, N118, N50, N268);
nor NOR2 (N305, N294, N25);
nand NAND4 (N306, N298, N126, N262, N173);
or OR3 (N307, N297, N246, N145);
and AND2 (N308, N293, N1);
or OR4 (N309, N302, N260, N262, N161);
nand NAND4 (N310, N307, N231, N19, N105);
or OR3 (N311, N304, N193, N95);
nand NAND3 (N312, N288, N5, N243);
not NOT1 (N313, N305);
and AND3 (N314, N309, N112, N245);
xor XOR2 (N315, N306, N259);
not NOT1 (N316, N311);
not NOT1 (N317, N312);
not NOT1 (N318, N315);
nand NAND4 (N319, N308, N251, N227, N177);
or OR4 (N320, N301, N198, N294, N289);
and AND3 (N321, N318, N43, N5);
and AND3 (N322, N321, N266, N311);
buf BUF1 (N323, N320);
nor NOR3 (N324, N322, N113, N41);
xor XOR2 (N325, N314, N71);
xor XOR2 (N326, N299, N300);
nand NAND3 (N327, N324, N233, N201);
or OR4 (N328, N317, N273, N299, N42);
nor NOR4 (N329, N326, N59, N14, N152);
not NOT1 (N330, N313);
nand NAND3 (N331, N310, N248, N316);
xor XOR2 (N332, N156, N2);
or OR4 (N333, N303, N76, N208, N285);
and AND3 (N334, N333, N153, N92);
buf BUF1 (N335, N332);
xor XOR2 (N336, N331, N172);
nor NOR2 (N337, N328, N78);
or OR2 (N338, N323, N298);
xor XOR2 (N339, N335, N294);
nand NAND2 (N340, N334, N34);
and AND4 (N341, N339, N88, N261, N144);
buf BUF1 (N342, N325);
xor XOR2 (N343, N342, N293);
not NOT1 (N344, N341);
nor NOR2 (N345, N340, N107);
or OR3 (N346, N329, N202, N109);
not NOT1 (N347, N346);
nor NOR3 (N348, N327, N245, N198);
and AND4 (N349, N348, N76, N289, N260);
nor NOR4 (N350, N319, N155, N180, N343);
not NOT1 (N351, N3);
nand NAND4 (N352, N330, N24, N215, N1);
xor XOR2 (N353, N347, N185);
nor NOR2 (N354, N349, N32);
xor XOR2 (N355, N336, N309);
not NOT1 (N356, N355);
or OR2 (N357, N345, N19);
not NOT1 (N358, N357);
xor XOR2 (N359, N354, N152);
not NOT1 (N360, N359);
not NOT1 (N361, N352);
or OR2 (N362, N356, N3);
nand NAND4 (N363, N358, N123, N332, N32);
and AND2 (N364, N351, N44);
or OR3 (N365, N350, N88, N225);
buf BUF1 (N366, N363);
nor NOR4 (N367, N362, N281, N264, N300);
xor XOR2 (N368, N366, N310);
or OR3 (N369, N337, N311, N329);
and AND2 (N370, N365, N79);
and AND4 (N371, N361, N198, N346, N203);
or OR2 (N372, N353, N38);
nand NAND3 (N373, N344, N229, N39);
nand NAND3 (N374, N370, N350, N39);
nand NAND2 (N375, N373, N263);
not NOT1 (N376, N372);
nor NOR3 (N377, N338, N69, N81);
buf BUF1 (N378, N374);
or OR3 (N379, N364, N258, N198);
xor XOR2 (N380, N378, N364);
not NOT1 (N381, N368);
or OR3 (N382, N376, N328, N328);
not NOT1 (N383, N369);
or OR3 (N384, N383, N307, N5);
nand NAND4 (N385, N367, N167, N12, N173);
or OR3 (N386, N360, N291, N33);
and AND4 (N387, N375, N314, N308, N360);
nand NAND4 (N388, N384, N305, N18, N2);
nand NAND4 (N389, N386, N327, N164, N363);
nor NOR3 (N390, N387, N157, N213);
buf BUF1 (N391, N382);
xor XOR2 (N392, N385, N97);
and AND4 (N393, N379, N314, N362, N388);
buf BUF1 (N394, N332);
xor XOR2 (N395, N389, N363);
xor XOR2 (N396, N394, N168);
nand NAND4 (N397, N393, N115, N312, N89);
xor XOR2 (N398, N395, N257);
and AND2 (N399, N391, N112);
not NOT1 (N400, N392);
not NOT1 (N401, N397);
nor NOR2 (N402, N399, N11);
nor NOR4 (N403, N396, N107, N351, N114);
or OR2 (N404, N380, N237);
nand NAND2 (N405, N404, N99);
or OR2 (N406, N400, N397);
or OR3 (N407, N402, N18, N369);
buf BUF1 (N408, N398);
nand NAND4 (N409, N371, N202, N246, N201);
nor NOR3 (N410, N377, N264, N311);
xor XOR2 (N411, N401, N301);
nor NOR4 (N412, N408, N364, N247, N312);
xor XOR2 (N413, N390, N63);
not NOT1 (N414, N403);
xor XOR2 (N415, N381, N413);
not NOT1 (N416, N352);
xor XOR2 (N417, N409, N249);
nor NOR2 (N418, N405, N377);
and AND2 (N419, N415, N11);
buf BUF1 (N420, N412);
or OR4 (N421, N416, N4, N386, N351);
nand NAND4 (N422, N410, N147, N219, N411);
buf BUF1 (N423, N360);
or OR3 (N424, N406, N331, N382);
xor XOR2 (N425, N421, N158);
xor XOR2 (N426, N407, N335);
and AND3 (N427, N420, N371, N63);
not NOT1 (N428, N423);
buf BUF1 (N429, N428);
xor XOR2 (N430, N414, N286);
or OR2 (N431, N418, N196);
not NOT1 (N432, N417);
buf BUF1 (N433, N419);
buf BUF1 (N434, N426);
xor XOR2 (N435, N433, N48);
nor NOR2 (N436, N427, N10);
nand NAND4 (N437, N429, N289, N370, N276);
nand NAND4 (N438, N422, N146, N291, N78);
or OR3 (N439, N432, N298, N390);
buf BUF1 (N440, N425);
buf BUF1 (N441, N437);
xor XOR2 (N442, N431, N336);
buf BUF1 (N443, N436);
nor NOR4 (N444, N439, N383, N2, N80);
not NOT1 (N445, N434);
nand NAND4 (N446, N435, N108, N400, N219);
and AND4 (N447, N441, N163, N265, N394);
nor NOR2 (N448, N446, N172);
xor XOR2 (N449, N438, N37);
not NOT1 (N450, N449);
not NOT1 (N451, N430);
nand NAND3 (N452, N451, N74, N172);
and AND4 (N453, N445, N237, N424, N375);
not NOT1 (N454, N63);
buf BUF1 (N455, N444);
nand NAND2 (N456, N450, N206);
nor NOR4 (N457, N454, N82, N101, N69);
nor NOR4 (N458, N456, N93, N261, N365);
not NOT1 (N459, N455);
nor NOR2 (N460, N442, N450);
and AND2 (N461, N452, N298);
and AND2 (N462, N440, N95);
or OR2 (N463, N447, N226);
buf BUF1 (N464, N448);
or OR2 (N465, N462, N251);
and AND4 (N466, N464, N236, N139, N123);
nand NAND2 (N467, N443, N104);
xor XOR2 (N468, N466, N22);
nand NAND4 (N469, N467, N44, N215, N165);
and AND2 (N470, N460, N349);
xor XOR2 (N471, N459, N423);
xor XOR2 (N472, N453, N177);
nand NAND3 (N473, N468, N126, N350);
buf BUF1 (N474, N469);
nand NAND3 (N475, N474, N279, N391);
nand NAND2 (N476, N470, N131);
nor NOR4 (N477, N465, N405, N92, N460);
or OR2 (N478, N476, N471);
nor NOR4 (N479, N424, N429, N351, N228);
or OR2 (N480, N472, N227);
or OR4 (N481, N477, N406, N182, N59);
nand NAND4 (N482, N473, N401, N203, N340);
nand NAND3 (N483, N482, N22, N22);
or OR4 (N484, N475, N222, N444, N435);
or OR3 (N485, N483, N272, N48);
buf BUF1 (N486, N480);
or OR2 (N487, N484, N258);
not NOT1 (N488, N458);
or OR4 (N489, N457, N221, N195, N456);
buf BUF1 (N490, N485);
not NOT1 (N491, N490);
nor NOR4 (N492, N491, N379, N293, N174);
not NOT1 (N493, N463);
or OR2 (N494, N486, N146);
not NOT1 (N495, N461);
buf BUF1 (N496, N479);
nand NAND2 (N497, N492, N358);
not NOT1 (N498, N494);
not NOT1 (N499, N493);
or OR4 (N500, N498, N151, N263, N295);
xor XOR2 (N501, N500, N139);
not NOT1 (N502, N489);
nand NAND4 (N503, N478, N400, N247, N399);
and AND2 (N504, N499, N363);
buf BUF1 (N505, N487);
xor XOR2 (N506, N496, N292);
buf BUF1 (N507, N505);
not NOT1 (N508, N503);
not NOT1 (N509, N506);
and AND2 (N510, N509, N493);
buf BUF1 (N511, N501);
or OR4 (N512, N510, N395, N407, N42);
xor XOR2 (N513, N488, N67);
buf BUF1 (N514, N504);
and AND3 (N515, N513, N290, N498);
nand NAND3 (N516, N495, N345, N49);
or OR4 (N517, N515, N223, N114, N456);
nand NAND4 (N518, N516, N160, N428, N271);
nor NOR2 (N519, N518, N481);
xor XOR2 (N520, N491, N489);
buf BUF1 (N521, N511);
or OR3 (N522, N517, N426, N272);
nor NOR2 (N523, N512, N454);
or OR4 (N524, N502, N22, N252, N248);
xor XOR2 (N525, N508, N137);
or OR2 (N526, N523, N262);
xor XOR2 (N527, N524, N105);
nand NAND2 (N528, N497, N137);
not NOT1 (N529, N522);
xor XOR2 (N530, N527, N309);
buf BUF1 (N531, N528);
nor NOR3 (N532, N525, N264, N139);
and AND2 (N533, N519, N361);
xor XOR2 (N534, N526, N212);
buf BUF1 (N535, N533);
xor XOR2 (N536, N531, N449);
buf BUF1 (N537, N520);
or OR2 (N538, N537, N368);
xor XOR2 (N539, N532, N411);
not NOT1 (N540, N514);
buf BUF1 (N541, N529);
and AND2 (N542, N541, N484);
nand NAND3 (N543, N535, N412, N454);
or OR4 (N544, N534, N29, N322, N123);
or OR3 (N545, N536, N410, N132);
or OR4 (N546, N538, N40, N54, N350);
nor NOR2 (N547, N530, N251);
buf BUF1 (N548, N545);
nand NAND2 (N549, N548, N519);
xor XOR2 (N550, N539, N25);
and AND2 (N551, N521, N47);
and AND4 (N552, N542, N37, N519, N454);
nor NOR3 (N553, N552, N166, N463);
buf BUF1 (N554, N547);
nor NOR4 (N555, N549, N40, N305, N400);
or OR2 (N556, N551, N187);
nor NOR3 (N557, N556, N120, N11);
nor NOR2 (N558, N555, N429);
nor NOR2 (N559, N550, N61);
not NOT1 (N560, N507);
nor NOR4 (N561, N544, N427, N526, N388);
nand NAND4 (N562, N557, N383, N92, N64);
xor XOR2 (N563, N561, N471);
buf BUF1 (N564, N546);
nand NAND3 (N565, N560, N200, N451);
xor XOR2 (N566, N540, N547);
buf BUF1 (N567, N558);
buf BUF1 (N568, N564);
nor NOR4 (N569, N565, N316, N381, N88);
not NOT1 (N570, N563);
not NOT1 (N571, N559);
buf BUF1 (N572, N553);
buf BUF1 (N573, N543);
buf BUF1 (N574, N554);
and AND4 (N575, N568, N199, N86, N394);
nand NAND4 (N576, N562, N35, N61, N58);
and AND3 (N577, N576, N351, N149);
not NOT1 (N578, N567);
nor NOR4 (N579, N573, N302, N391, N433);
nor NOR3 (N580, N566, N452, N441);
nor NOR3 (N581, N577, N350, N34);
nand NAND2 (N582, N579, N468);
buf BUF1 (N583, N572);
buf BUF1 (N584, N578);
buf BUF1 (N585, N581);
nand NAND2 (N586, N570, N294);
and AND4 (N587, N575, N313, N218, N78);
nand NAND2 (N588, N583, N545);
nor NOR3 (N589, N580, N480, N279);
xor XOR2 (N590, N571, N327);
nor NOR2 (N591, N588, N461);
or OR4 (N592, N569, N560, N556, N440);
nor NOR4 (N593, N585, N66, N300, N585);
and AND4 (N594, N593, N329, N28, N262);
not NOT1 (N595, N591);
nand NAND2 (N596, N589, N10);
nand NAND2 (N597, N586, N428);
or OR3 (N598, N592, N518, N469);
nand NAND4 (N599, N587, N310, N46, N444);
buf BUF1 (N600, N582);
and AND3 (N601, N584, N240, N145);
xor XOR2 (N602, N597, N62);
nand NAND2 (N603, N601, N415);
and AND2 (N604, N590, N101);
buf BUF1 (N605, N595);
not NOT1 (N606, N602);
xor XOR2 (N607, N606, N238);
nand NAND4 (N608, N604, N150, N115, N541);
nand NAND4 (N609, N599, N234, N191, N497);
nand NAND3 (N610, N608, N384, N157);
buf BUF1 (N611, N574);
buf BUF1 (N612, N598);
nor NOR4 (N613, N611, N523, N578, N70);
not NOT1 (N614, N605);
not NOT1 (N615, N607);
and AND4 (N616, N613, N403, N568, N12);
not NOT1 (N617, N603);
or OR3 (N618, N617, N513, N558);
buf BUF1 (N619, N594);
nand NAND2 (N620, N614, N264);
or OR2 (N621, N615, N54);
not NOT1 (N622, N610);
xor XOR2 (N623, N620, N22);
or OR3 (N624, N619, N310, N373);
or OR4 (N625, N609, N444, N263, N156);
not NOT1 (N626, N623);
nand NAND3 (N627, N596, N358, N282);
nor NOR2 (N628, N622, N60);
xor XOR2 (N629, N624, N539);
buf BUF1 (N630, N618);
or OR4 (N631, N630, N9, N241, N102);
xor XOR2 (N632, N626, N224);
xor XOR2 (N633, N629, N517);
nor NOR3 (N634, N625, N553, N596);
or OR2 (N635, N621, N73);
xor XOR2 (N636, N633, N239);
nand NAND2 (N637, N616, N138);
xor XOR2 (N638, N635, N255);
buf BUF1 (N639, N638);
and AND4 (N640, N637, N88, N192, N638);
nand NAND3 (N641, N632, N545, N56);
or OR3 (N642, N628, N25, N493);
nand NAND4 (N643, N641, N104, N221, N126);
nor NOR3 (N644, N631, N510, N614);
xor XOR2 (N645, N643, N138);
or OR4 (N646, N600, N184, N594, N156);
buf BUF1 (N647, N634);
or OR4 (N648, N627, N259, N501, N430);
nor NOR4 (N649, N636, N544, N356, N483);
and AND4 (N650, N640, N373, N364, N220);
nand NAND2 (N651, N639, N172);
xor XOR2 (N652, N651, N624);
and AND2 (N653, N647, N342);
nor NOR4 (N654, N648, N319, N620, N173);
buf BUF1 (N655, N644);
buf BUF1 (N656, N655);
not NOT1 (N657, N653);
not NOT1 (N658, N642);
buf BUF1 (N659, N654);
and AND4 (N660, N612, N431, N603, N79);
nor NOR2 (N661, N649, N613);
xor XOR2 (N662, N645, N324);
nor NOR4 (N663, N656, N265, N259, N418);
or OR2 (N664, N661, N354);
xor XOR2 (N665, N659, N503);
xor XOR2 (N666, N646, N3);
buf BUF1 (N667, N663);
buf BUF1 (N668, N652);
nor NOR2 (N669, N664, N370);
not NOT1 (N670, N665);
buf BUF1 (N671, N668);
not NOT1 (N672, N670);
not NOT1 (N673, N666);
and AND3 (N674, N657, N514, N491);
nand NAND3 (N675, N667, N608, N209);
xor XOR2 (N676, N660, N301);
and AND2 (N677, N658, N468);
and AND3 (N678, N673, N34, N201);
and AND3 (N679, N650, N451, N479);
and AND3 (N680, N669, N386, N70);
and AND2 (N681, N672, N646);
nor NOR4 (N682, N675, N37, N262, N623);
xor XOR2 (N683, N679, N490);
not NOT1 (N684, N678);
xor XOR2 (N685, N676, N414);
xor XOR2 (N686, N680, N407);
nand NAND2 (N687, N677, N595);
and AND3 (N688, N662, N376, N201);
nand NAND3 (N689, N684, N247, N342);
nand NAND3 (N690, N687, N368, N258);
nor NOR2 (N691, N686, N455);
xor XOR2 (N692, N682, N412);
nor NOR3 (N693, N690, N239, N327);
nand NAND3 (N694, N681, N26, N416);
buf BUF1 (N695, N692);
nor NOR2 (N696, N691, N143);
or OR2 (N697, N695, N440);
nor NOR4 (N698, N674, N418, N254, N600);
and AND4 (N699, N696, N301, N627, N343);
buf BUF1 (N700, N688);
buf BUF1 (N701, N685);
nor NOR4 (N702, N697, N329, N380, N606);
buf BUF1 (N703, N701);
not NOT1 (N704, N700);
buf BUF1 (N705, N702);
or OR2 (N706, N689, N62);
and AND3 (N707, N699, N668, N298);
nand NAND2 (N708, N706, N141);
or OR3 (N709, N704, N230, N411);
nand NAND3 (N710, N671, N697, N384);
nand NAND2 (N711, N709, N608);
buf BUF1 (N712, N710);
nand NAND4 (N713, N708, N32, N571, N437);
not NOT1 (N714, N711);
not NOT1 (N715, N713);
nor NOR3 (N716, N694, N551, N429);
not NOT1 (N717, N693);
nand NAND2 (N718, N683, N232);
xor XOR2 (N719, N715, N13);
and AND4 (N720, N703, N661, N240, N410);
xor XOR2 (N721, N719, N536);
not NOT1 (N722, N716);
xor XOR2 (N723, N720, N148);
or OR2 (N724, N698, N298);
or OR2 (N725, N707, N142);
buf BUF1 (N726, N725);
not NOT1 (N727, N726);
not NOT1 (N728, N718);
nor NOR2 (N729, N717, N386);
and AND2 (N730, N712, N283);
buf BUF1 (N731, N723);
nor NOR3 (N732, N722, N347, N135);
not NOT1 (N733, N727);
and AND2 (N734, N729, N667);
nor NOR3 (N735, N732, N7, N723);
not NOT1 (N736, N731);
xor XOR2 (N737, N735, N95);
xor XOR2 (N738, N705, N39);
buf BUF1 (N739, N734);
and AND3 (N740, N733, N308, N568);
nor NOR2 (N741, N724, N416);
nand NAND4 (N742, N741, N400, N52, N468);
nand NAND2 (N743, N714, N454);
or OR2 (N744, N728, N496);
nor NOR3 (N745, N740, N340, N661);
nor NOR3 (N746, N730, N627, N603);
xor XOR2 (N747, N746, N602);
buf BUF1 (N748, N743);
or OR3 (N749, N737, N615, N579);
nor NOR3 (N750, N739, N432, N699);
nand NAND4 (N751, N749, N656, N586, N630);
nor NOR2 (N752, N750, N4);
not NOT1 (N753, N747);
and AND4 (N754, N721, N729, N445, N416);
or OR3 (N755, N753, N557, N261);
and AND2 (N756, N751, N293);
nand NAND2 (N757, N744, N551);
and AND2 (N758, N754, N229);
or OR3 (N759, N752, N112, N508);
xor XOR2 (N760, N759, N739);
not NOT1 (N761, N745);
not NOT1 (N762, N755);
buf BUF1 (N763, N760);
and AND3 (N764, N756, N626, N540);
or OR4 (N765, N758, N274, N505, N226);
nor NOR2 (N766, N765, N18);
and AND3 (N767, N757, N285, N6);
not NOT1 (N768, N764);
nor NOR2 (N769, N767, N363);
xor XOR2 (N770, N768, N654);
xor XOR2 (N771, N770, N723);
or OR2 (N772, N742, N632);
nor NOR3 (N773, N771, N205, N641);
nand NAND4 (N774, N761, N334, N750, N105);
or OR4 (N775, N769, N705, N765, N161);
not NOT1 (N776, N773);
or OR2 (N777, N776, N705);
and AND2 (N778, N762, N766);
nor NOR4 (N779, N54, N226, N635, N612);
not NOT1 (N780, N736);
nor NOR3 (N781, N779, N670, N440);
or OR4 (N782, N781, N711, N705, N552);
buf BUF1 (N783, N738);
xor XOR2 (N784, N782, N65);
buf BUF1 (N785, N784);
buf BUF1 (N786, N772);
or OR4 (N787, N763, N396, N706, N638);
nor NOR2 (N788, N783, N172);
xor XOR2 (N789, N785, N702);
or OR2 (N790, N786, N220);
not NOT1 (N791, N780);
and AND2 (N792, N775, N124);
nor NOR2 (N793, N748, N221);
nor NOR2 (N794, N791, N581);
nand NAND3 (N795, N774, N702, N90);
xor XOR2 (N796, N795, N588);
or OR2 (N797, N789, N495);
nand NAND4 (N798, N778, N113, N416, N648);
nand NAND3 (N799, N798, N659, N472);
not NOT1 (N800, N797);
xor XOR2 (N801, N794, N737);
nor NOR3 (N802, N800, N497, N281);
buf BUF1 (N803, N793);
and AND4 (N804, N799, N564, N93, N193);
buf BUF1 (N805, N804);
buf BUF1 (N806, N790);
and AND2 (N807, N806, N674);
and AND4 (N808, N788, N802, N289, N46);
or OR3 (N809, N408, N733, N677);
xor XOR2 (N810, N803, N369);
buf BUF1 (N811, N808);
nor NOR4 (N812, N807, N637, N290, N721);
nor NOR3 (N813, N777, N132, N21);
or OR2 (N814, N792, N260);
or OR2 (N815, N810, N714);
nor NOR2 (N816, N812, N586);
xor XOR2 (N817, N814, N552);
and AND2 (N818, N811, N414);
buf BUF1 (N819, N818);
or OR4 (N820, N813, N157, N686, N781);
nor NOR2 (N821, N801, N541);
or OR4 (N822, N796, N140, N197, N667);
xor XOR2 (N823, N822, N776);
buf BUF1 (N824, N787);
and AND4 (N825, N816, N381, N580, N469);
xor XOR2 (N826, N823, N736);
not NOT1 (N827, N805);
not NOT1 (N828, N819);
buf BUF1 (N829, N824);
nand NAND3 (N830, N829, N649, N778);
not NOT1 (N831, N821);
nor NOR3 (N832, N817, N333, N183);
and AND3 (N833, N815, N279, N172);
xor XOR2 (N834, N820, N32);
buf BUF1 (N835, N827);
xor XOR2 (N836, N830, N221);
not NOT1 (N837, N825);
or OR4 (N838, N834, N799, N278, N821);
or OR4 (N839, N831, N610, N98, N427);
not NOT1 (N840, N835);
xor XOR2 (N841, N833, N264);
or OR4 (N842, N832, N114, N370, N532);
nor NOR3 (N843, N836, N24, N453);
nor NOR3 (N844, N840, N32, N175);
buf BUF1 (N845, N839);
nand NAND3 (N846, N844, N77, N352);
buf BUF1 (N847, N828);
buf BUF1 (N848, N837);
and AND4 (N849, N826, N818, N525, N49);
nand NAND2 (N850, N849, N766);
buf BUF1 (N851, N843);
xor XOR2 (N852, N809, N612);
nand NAND3 (N853, N850, N286, N368);
nand NAND3 (N854, N846, N268, N616);
not NOT1 (N855, N852);
nand NAND4 (N856, N847, N363, N412, N534);
nand NAND4 (N857, N848, N782, N526, N669);
nor NOR2 (N858, N838, N246);
and AND4 (N859, N855, N560, N446, N667);
xor XOR2 (N860, N859, N463);
buf BUF1 (N861, N842);
nor NOR4 (N862, N861, N80, N313, N852);
or OR3 (N863, N854, N375, N461);
nor NOR4 (N864, N853, N461, N358, N209);
and AND3 (N865, N858, N351, N619);
or OR4 (N866, N862, N436, N180, N54);
nand NAND4 (N867, N865, N820, N851, N543);
xor XOR2 (N868, N128, N635);
not NOT1 (N869, N841);
xor XOR2 (N870, N857, N288);
buf BUF1 (N871, N868);
or OR2 (N872, N845, N436);
nor NOR2 (N873, N872, N691);
nor NOR2 (N874, N873, N73);
nor NOR2 (N875, N874, N237);
or OR2 (N876, N866, N669);
nor NOR2 (N877, N860, N551);
nand NAND4 (N878, N869, N316, N171, N527);
nor NOR4 (N879, N877, N548, N71, N364);
nor NOR2 (N880, N876, N148);
not NOT1 (N881, N871);
or OR3 (N882, N870, N432, N423);
and AND4 (N883, N878, N182, N207, N38);
nor NOR2 (N884, N879, N658);
not NOT1 (N885, N882);
nor NOR2 (N886, N881, N13);
nor NOR2 (N887, N867, N833);
and AND4 (N888, N886, N802, N856, N325);
and AND4 (N889, N452, N330, N22, N432);
or OR4 (N890, N889, N311, N761, N158);
nand NAND4 (N891, N885, N116, N857, N697);
not NOT1 (N892, N887);
and AND3 (N893, N884, N759, N687);
xor XOR2 (N894, N875, N669);
buf BUF1 (N895, N863);
xor XOR2 (N896, N864, N388);
nor NOR2 (N897, N896, N839);
xor XOR2 (N898, N893, N646);
or OR4 (N899, N892, N474, N196, N271);
xor XOR2 (N900, N883, N557);
nand NAND2 (N901, N897, N653);
or OR2 (N902, N894, N872);
not NOT1 (N903, N890);
nor NOR2 (N904, N899, N491);
nand NAND4 (N905, N903, N761, N747, N449);
buf BUF1 (N906, N901);
buf BUF1 (N907, N905);
and AND3 (N908, N902, N290, N600);
nand NAND3 (N909, N900, N509, N742);
or OR2 (N910, N906, N672);
nand NAND2 (N911, N904, N400);
or OR4 (N912, N911, N592, N794, N639);
not NOT1 (N913, N888);
nand NAND2 (N914, N898, N736);
or OR2 (N915, N910, N838);
and AND3 (N916, N891, N762, N604);
or OR4 (N917, N916, N830, N675, N583);
not NOT1 (N918, N895);
xor XOR2 (N919, N908, N237);
or OR2 (N920, N907, N236);
nor NOR3 (N921, N913, N38, N787);
xor XOR2 (N922, N915, N617);
buf BUF1 (N923, N920);
not NOT1 (N924, N909);
xor XOR2 (N925, N924, N720);
and AND2 (N926, N921, N836);
or OR2 (N927, N926, N799);
and AND3 (N928, N925, N18, N89);
nand NAND4 (N929, N880, N339, N67, N529);
buf BUF1 (N930, N928);
and AND2 (N931, N927, N464);
buf BUF1 (N932, N930);
buf BUF1 (N933, N923);
or OR4 (N934, N919, N288, N845, N921);
not NOT1 (N935, N929);
or OR4 (N936, N934, N262, N200, N242);
and AND2 (N937, N935, N262);
not NOT1 (N938, N932);
nand NAND2 (N939, N922, N89);
and AND3 (N940, N918, N420, N726);
buf BUF1 (N941, N938);
and AND4 (N942, N936, N698, N183, N462);
nor NOR4 (N943, N937, N688, N213, N181);
not NOT1 (N944, N912);
buf BUF1 (N945, N917);
not NOT1 (N946, N941);
and AND2 (N947, N939, N242);
xor XOR2 (N948, N931, N172);
or OR3 (N949, N947, N902, N389);
xor XOR2 (N950, N945, N443);
nand NAND4 (N951, N914, N646, N853, N518);
xor XOR2 (N952, N951, N789);
or OR4 (N953, N949, N111, N830, N860);
nor NOR2 (N954, N950, N43);
xor XOR2 (N955, N953, N380);
xor XOR2 (N956, N943, N64);
nor NOR3 (N957, N952, N804, N846);
not NOT1 (N958, N957);
and AND3 (N959, N954, N552, N635);
or OR2 (N960, N959, N337);
or OR4 (N961, N944, N87, N477, N620);
nor NOR4 (N962, N960, N956, N316, N565);
nand NAND4 (N963, N357, N57, N512, N225);
buf BUF1 (N964, N940);
not NOT1 (N965, N942);
xor XOR2 (N966, N933, N362);
and AND3 (N967, N961, N659, N184);
or OR2 (N968, N966, N822);
xor XOR2 (N969, N963, N50);
not NOT1 (N970, N955);
nor NOR2 (N971, N968, N737);
and AND2 (N972, N964, N73);
or OR4 (N973, N967, N56, N948, N436);
not NOT1 (N974, N828);
buf BUF1 (N975, N974);
xor XOR2 (N976, N946, N861);
nor NOR3 (N977, N958, N591, N740);
not NOT1 (N978, N971);
or OR2 (N979, N975, N327);
xor XOR2 (N980, N978, N588);
or OR4 (N981, N980, N205, N504, N393);
nand NAND2 (N982, N969, N785);
nor NOR2 (N983, N972, N416);
and AND2 (N984, N965, N690);
nor NOR3 (N985, N984, N496, N776);
or OR4 (N986, N979, N629, N887, N261);
buf BUF1 (N987, N977);
and AND3 (N988, N970, N220, N543);
or OR4 (N989, N982, N177, N793, N538);
xor XOR2 (N990, N976, N703);
and AND2 (N991, N973, N370);
nor NOR3 (N992, N985, N190, N450);
buf BUF1 (N993, N983);
xor XOR2 (N994, N993, N487);
buf BUF1 (N995, N988);
nand NAND4 (N996, N986, N151, N651, N686);
buf BUF1 (N997, N994);
nand NAND4 (N998, N991, N217, N17, N979);
nand NAND2 (N999, N997, N982);
and AND2 (N1000, N992, N713);
buf BUF1 (N1001, N998);
buf BUF1 (N1002, N962);
nor NOR2 (N1003, N981, N237);
nor NOR2 (N1004, N989, N692);
nand NAND3 (N1005, N996, N159, N756);
buf BUF1 (N1006, N1002);
nor NOR2 (N1007, N990, N420);
or OR4 (N1008, N1003, N290, N215, N120);
not NOT1 (N1009, N999);
not NOT1 (N1010, N1007);
and AND3 (N1011, N1008, N80, N148);
not NOT1 (N1012, N995);
nor NOR3 (N1013, N1005, N645, N637);
and AND3 (N1014, N1004, N554, N465);
nor NOR3 (N1015, N1012, N717, N549);
nand NAND4 (N1016, N1011, N266, N966, N625);
nand NAND4 (N1017, N1009, N251, N345, N963);
and AND4 (N1018, N1016, N991, N3, N596);
and AND3 (N1019, N1018, N208, N504);
xor XOR2 (N1020, N1013, N609);
and AND4 (N1021, N1019, N228, N409, N72);
nand NAND3 (N1022, N1017, N182, N644);
not NOT1 (N1023, N1020);
nand NAND3 (N1024, N1006, N387, N659);
nand NAND2 (N1025, N1022, N469);
buf BUF1 (N1026, N1014);
xor XOR2 (N1027, N1010, N240);
nor NOR4 (N1028, N1001, N340, N564, N389);
buf BUF1 (N1029, N1025);
and AND4 (N1030, N1000, N941, N32, N15);
not NOT1 (N1031, N1021);
xor XOR2 (N1032, N1024, N78);
or OR3 (N1033, N1027, N860, N687);
buf BUF1 (N1034, N1026);
not NOT1 (N1035, N1029);
and AND3 (N1036, N1023, N571, N951);
or OR3 (N1037, N1036, N841, N693);
nor NOR4 (N1038, N1037, N592, N586, N424);
buf BUF1 (N1039, N1035);
nand NAND2 (N1040, N987, N128);
xor XOR2 (N1041, N1015, N352);
not NOT1 (N1042, N1030);
nand NAND2 (N1043, N1041, N826);
nor NOR4 (N1044, N1028, N136, N245, N49);
and AND3 (N1045, N1042, N394, N651);
and AND4 (N1046, N1045, N580, N719, N744);
buf BUF1 (N1047, N1039);
xor XOR2 (N1048, N1033, N678);
buf BUF1 (N1049, N1038);
or OR3 (N1050, N1043, N465, N450);
not NOT1 (N1051, N1048);
and AND2 (N1052, N1040, N576);
and AND2 (N1053, N1046, N737);
xor XOR2 (N1054, N1031, N206);
buf BUF1 (N1055, N1054);
nand NAND3 (N1056, N1032, N72, N667);
xor XOR2 (N1057, N1051, N194);
nand NAND4 (N1058, N1056, N788, N73, N721);
not NOT1 (N1059, N1044);
xor XOR2 (N1060, N1034, N576);
or OR2 (N1061, N1058, N598);
buf BUF1 (N1062, N1059);
and AND3 (N1063, N1060, N874, N8);
buf BUF1 (N1064, N1061);
or OR4 (N1065, N1062, N687, N838, N992);
not NOT1 (N1066, N1064);
xor XOR2 (N1067, N1049, N190);
or OR3 (N1068, N1052, N1056, N248);
nor NOR4 (N1069, N1050, N238, N28, N502);
nor NOR4 (N1070, N1068, N728, N341, N34);
buf BUF1 (N1071, N1063);
or OR4 (N1072, N1053, N910, N453, N731);
buf BUF1 (N1073, N1072);
buf BUF1 (N1074, N1066);
buf BUF1 (N1075, N1073);
or OR4 (N1076, N1069, N216, N880, N271);
nor NOR4 (N1077, N1075, N8, N806, N249);
buf BUF1 (N1078, N1077);
not NOT1 (N1079, N1065);
and AND4 (N1080, N1057, N151, N547, N302);
or OR3 (N1081, N1047, N551, N998);
xor XOR2 (N1082, N1079, N215);
and AND4 (N1083, N1070, N182, N239, N1076);
xor XOR2 (N1084, N830, N759);
or OR4 (N1085, N1080, N202, N720, N340);
nor NOR4 (N1086, N1078, N549, N381, N752);
not NOT1 (N1087, N1071);
nor NOR2 (N1088, N1074, N766);
and AND4 (N1089, N1084, N946, N210, N680);
or OR2 (N1090, N1085, N1057);
nor NOR3 (N1091, N1067, N929, N76);
nor NOR4 (N1092, N1055, N1037, N474, N467);
xor XOR2 (N1093, N1090, N971);
nand NAND2 (N1094, N1088, N837);
and AND2 (N1095, N1092, N722);
xor XOR2 (N1096, N1095, N1073);
not NOT1 (N1097, N1082);
xor XOR2 (N1098, N1083, N101);
xor XOR2 (N1099, N1098, N86);
nand NAND3 (N1100, N1096, N993, N407);
nor NOR2 (N1101, N1086, N907);
or OR2 (N1102, N1097, N832);
and AND4 (N1103, N1081, N998, N392, N625);
nor NOR3 (N1104, N1102, N221, N291);
and AND2 (N1105, N1093, N932);
not NOT1 (N1106, N1105);
nor NOR3 (N1107, N1087, N699, N406);
not NOT1 (N1108, N1089);
buf BUF1 (N1109, N1106);
and AND2 (N1110, N1107, N772);
nand NAND4 (N1111, N1104, N553, N570, N950);
or OR2 (N1112, N1091, N84);
nand NAND2 (N1113, N1111, N1079);
and AND2 (N1114, N1110, N634);
buf BUF1 (N1115, N1109);
or OR2 (N1116, N1115, N106);
or OR3 (N1117, N1116, N885, N777);
and AND2 (N1118, N1094, N201);
xor XOR2 (N1119, N1118, N299);
or OR2 (N1120, N1113, N130);
nor NOR2 (N1121, N1119, N194);
buf BUF1 (N1122, N1117);
or OR3 (N1123, N1112, N929, N547);
buf BUF1 (N1124, N1099);
xor XOR2 (N1125, N1103, N200);
nor NOR2 (N1126, N1100, N533);
buf BUF1 (N1127, N1101);
buf BUF1 (N1128, N1127);
xor XOR2 (N1129, N1123, N558);
xor XOR2 (N1130, N1129, N703);
and AND3 (N1131, N1120, N193, N588);
buf BUF1 (N1132, N1131);
not NOT1 (N1133, N1125);
buf BUF1 (N1134, N1122);
xor XOR2 (N1135, N1114, N271);
nand NAND2 (N1136, N1121, N251);
nor NOR2 (N1137, N1135, N812);
nand NAND2 (N1138, N1130, N1105);
nor NOR3 (N1139, N1137, N1101, N1012);
nand NAND4 (N1140, N1124, N264, N1018, N642);
nor NOR4 (N1141, N1138, N724, N415, N72);
or OR2 (N1142, N1108, N505);
and AND4 (N1143, N1128, N433, N721, N48);
nand NAND3 (N1144, N1132, N963, N1008);
nor NOR3 (N1145, N1143, N255, N287);
or OR3 (N1146, N1141, N353, N308);
buf BUF1 (N1147, N1146);
nor NOR3 (N1148, N1133, N457, N953);
xor XOR2 (N1149, N1139, N682);
nor NOR2 (N1150, N1148, N674);
and AND3 (N1151, N1136, N366, N146);
nor NOR3 (N1152, N1140, N473, N768);
or OR3 (N1153, N1150, N347, N1033);
nor NOR2 (N1154, N1152, N135);
nand NAND3 (N1155, N1154, N1071, N1028);
or OR3 (N1156, N1151, N387, N922);
xor XOR2 (N1157, N1144, N487);
nand NAND4 (N1158, N1145, N271, N727, N1134);
or OR2 (N1159, N317, N372);
xor XOR2 (N1160, N1157, N754);
nor NOR4 (N1161, N1159, N1048, N121, N1118);
nor NOR3 (N1162, N1147, N260, N182);
not NOT1 (N1163, N1142);
nor NOR2 (N1164, N1155, N404);
nor NOR4 (N1165, N1164, N1013, N569, N567);
and AND2 (N1166, N1126, N1160);
or OR4 (N1167, N290, N1104, N86, N652);
nand NAND2 (N1168, N1153, N167);
not NOT1 (N1169, N1163);
buf BUF1 (N1170, N1169);
or OR4 (N1171, N1166, N548, N975, N8);
xor XOR2 (N1172, N1170, N509);
nand NAND3 (N1173, N1165, N786, N860);
nand NAND2 (N1174, N1167, N144);
and AND4 (N1175, N1174, N805, N142, N590);
and AND4 (N1176, N1172, N696, N131, N1052);
nor NOR4 (N1177, N1176, N198, N683, N103);
not NOT1 (N1178, N1177);
buf BUF1 (N1179, N1149);
and AND3 (N1180, N1171, N1120, N578);
buf BUF1 (N1181, N1175);
and AND3 (N1182, N1180, N84, N350);
or OR4 (N1183, N1179, N521, N914, N1054);
xor XOR2 (N1184, N1158, N893);
or OR3 (N1185, N1184, N477, N486);
nor NOR2 (N1186, N1173, N489);
buf BUF1 (N1187, N1178);
xor XOR2 (N1188, N1156, N1099);
or OR3 (N1189, N1187, N260, N514);
nand NAND4 (N1190, N1168, N1093, N534, N157);
nand NAND2 (N1191, N1189, N62);
nand NAND4 (N1192, N1161, N539, N510, N569);
xor XOR2 (N1193, N1185, N406);
nor NOR2 (N1194, N1188, N424);
nand NAND3 (N1195, N1183, N1103, N938);
nand NAND3 (N1196, N1191, N298, N137);
nor NOR4 (N1197, N1194, N151, N1021, N1100);
buf BUF1 (N1198, N1197);
nor NOR4 (N1199, N1181, N304, N456, N95);
nand NAND4 (N1200, N1182, N205, N1138, N1188);
and AND3 (N1201, N1186, N934, N322);
and AND4 (N1202, N1200, N40, N23, N1009);
nor NOR3 (N1203, N1196, N403, N522);
buf BUF1 (N1204, N1203);
nor NOR4 (N1205, N1190, N281, N898, N1119);
and AND2 (N1206, N1199, N54);
nor NOR4 (N1207, N1198, N716, N191, N946);
buf BUF1 (N1208, N1205);
nand NAND2 (N1209, N1206, N118);
and AND2 (N1210, N1192, N978);
or OR2 (N1211, N1162, N541);
not NOT1 (N1212, N1193);
xor XOR2 (N1213, N1207, N1017);
nor NOR4 (N1214, N1210, N368, N624, N1116);
nor NOR3 (N1215, N1201, N347, N430);
nand NAND4 (N1216, N1215, N269, N376, N645);
and AND3 (N1217, N1213, N979, N678);
nor NOR2 (N1218, N1214, N1032);
nand NAND2 (N1219, N1195, N1161);
buf BUF1 (N1220, N1202);
not NOT1 (N1221, N1204);
xor XOR2 (N1222, N1221, N415);
xor XOR2 (N1223, N1219, N21);
and AND2 (N1224, N1212, N857);
nand NAND3 (N1225, N1217, N121, N874);
not NOT1 (N1226, N1222);
not NOT1 (N1227, N1225);
nor NOR2 (N1228, N1218, N371);
nand NAND2 (N1229, N1216, N530);
and AND2 (N1230, N1227, N869);
or OR3 (N1231, N1223, N81, N1029);
xor XOR2 (N1232, N1229, N1078);
not NOT1 (N1233, N1230);
or OR4 (N1234, N1211, N67, N875, N86);
and AND4 (N1235, N1233, N169, N865, N667);
nand NAND2 (N1236, N1208, N1111);
nand NAND2 (N1237, N1220, N463);
and AND2 (N1238, N1234, N729);
or OR3 (N1239, N1232, N77, N722);
and AND4 (N1240, N1238, N180, N756, N101);
and AND3 (N1241, N1240, N856, N85);
xor XOR2 (N1242, N1209, N617);
xor XOR2 (N1243, N1226, N565);
buf BUF1 (N1244, N1242);
or OR3 (N1245, N1239, N939, N1146);
and AND4 (N1246, N1243, N842, N339, N213);
nor NOR4 (N1247, N1228, N761, N215, N520);
xor XOR2 (N1248, N1237, N552);
not NOT1 (N1249, N1235);
nor NOR3 (N1250, N1247, N621, N160);
xor XOR2 (N1251, N1236, N656);
or OR4 (N1252, N1246, N1086, N676, N865);
not NOT1 (N1253, N1249);
or OR4 (N1254, N1253, N172, N85, N877);
nor NOR3 (N1255, N1248, N232, N1225);
buf BUF1 (N1256, N1250);
or OR3 (N1257, N1241, N297, N1071);
not NOT1 (N1258, N1255);
xor XOR2 (N1259, N1251, N167);
buf BUF1 (N1260, N1224);
and AND4 (N1261, N1254, N391, N1163, N644);
not NOT1 (N1262, N1244);
xor XOR2 (N1263, N1252, N678);
or OR3 (N1264, N1231, N158, N721);
and AND2 (N1265, N1264, N552);
not NOT1 (N1266, N1259);
nand NAND2 (N1267, N1262, N49);
buf BUF1 (N1268, N1263);
buf BUF1 (N1269, N1265);
and AND2 (N1270, N1258, N1163);
xor XOR2 (N1271, N1267, N253);
or OR2 (N1272, N1268, N1210);
nand NAND2 (N1273, N1245, N643);
and AND3 (N1274, N1260, N1271, N827);
or OR2 (N1275, N549, N350);
nor NOR3 (N1276, N1266, N313, N1222);
or OR4 (N1277, N1276, N708, N563, N304);
or OR4 (N1278, N1261, N401, N1262, N448);
or OR2 (N1279, N1269, N347);
nor NOR3 (N1280, N1279, N1181, N433);
nand NAND3 (N1281, N1274, N486, N1070);
nor NOR2 (N1282, N1270, N718);
nand NAND3 (N1283, N1280, N238, N41);
xor XOR2 (N1284, N1277, N649);
not NOT1 (N1285, N1284);
or OR2 (N1286, N1273, N1067);
buf BUF1 (N1287, N1283);
or OR2 (N1288, N1278, N803);
or OR4 (N1289, N1285, N601, N229, N286);
nand NAND3 (N1290, N1257, N379, N97);
nor NOR3 (N1291, N1289, N145, N9);
xor XOR2 (N1292, N1275, N318);
nand NAND2 (N1293, N1292, N1003);
nor NOR3 (N1294, N1281, N1238, N36);
and AND3 (N1295, N1290, N1054, N623);
not NOT1 (N1296, N1286);
not NOT1 (N1297, N1295);
nor NOR2 (N1298, N1256, N454);
xor XOR2 (N1299, N1291, N896);
not NOT1 (N1300, N1297);
or OR4 (N1301, N1298, N153, N752, N1094);
buf BUF1 (N1302, N1294);
or OR3 (N1303, N1293, N903, N374);
or OR2 (N1304, N1272, N319);
not NOT1 (N1305, N1288);
nor NOR4 (N1306, N1303, N792, N1191, N636);
nor NOR3 (N1307, N1306, N147, N221);
nor NOR3 (N1308, N1287, N1193, N1203);
nor NOR4 (N1309, N1308, N514, N614, N1268);
not NOT1 (N1310, N1304);
or OR3 (N1311, N1305, N412, N1290);
nand NAND3 (N1312, N1299, N1248, N381);
nor NOR2 (N1313, N1302, N1232);
and AND4 (N1314, N1310, N337, N1129, N706);
and AND3 (N1315, N1313, N95, N70);
nand NAND3 (N1316, N1312, N789, N848);
nand NAND3 (N1317, N1307, N99, N831);
xor XOR2 (N1318, N1315, N1212);
buf BUF1 (N1319, N1316);
buf BUF1 (N1320, N1296);
nand NAND2 (N1321, N1309, N874);
and AND3 (N1322, N1301, N164, N358);
not NOT1 (N1323, N1321);
or OR2 (N1324, N1318, N547);
or OR4 (N1325, N1282, N568, N690, N1062);
not NOT1 (N1326, N1320);
nand NAND2 (N1327, N1311, N253);
xor XOR2 (N1328, N1325, N1196);
buf BUF1 (N1329, N1326);
and AND4 (N1330, N1328, N991, N642, N685);
nand NAND3 (N1331, N1327, N707, N1195);
xor XOR2 (N1332, N1300, N1135);
nor NOR4 (N1333, N1322, N15, N403, N596);
or OR2 (N1334, N1324, N91);
xor XOR2 (N1335, N1332, N1007);
xor XOR2 (N1336, N1314, N1030);
nand NAND3 (N1337, N1334, N1225, N1043);
nand NAND3 (N1338, N1331, N1164, N628);
or OR2 (N1339, N1329, N421);
or OR3 (N1340, N1333, N160, N772);
xor XOR2 (N1341, N1338, N776);
not NOT1 (N1342, N1336);
nor NOR2 (N1343, N1337, N1337);
and AND2 (N1344, N1339, N246);
nor NOR4 (N1345, N1340, N375, N974, N748);
buf BUF1 (N1346, N1343);
nand NAND3 (N1347, N1319, N419, N520);
nor NOR4 (N1348, N1335, N1060, N1007, N822);
buf BUF1 (N1349, N1347);
or OR4 (N1350, N1342, N895, N397, N633);
buf BUF1 (N1351, N1346);
nand NAND3 (N1352, N1344, N8, N526);
buf BUF1 (N1353, N1323);
nand NAND4 (N1354, N1317, N1338, N746, N170);
xor XOR2 (N1355, N1354, N1214);
not NOT1 (N1356, N1351);
and AND4 (N1357, N1348, N939, N508, N587);
nand NAND2 (N1358, N1353, N744);
or OR2 (N1359, N1330, N755);
nor NOR4 (N1360, N1356, N939, N1141, N529);
and AND3 (N1361, N1359, N259, N160);
nor NOR4 (N1362, N1345, N1061, N543, N954);
xor XOR2 (N1363, N1349, N22);
or OR2 (N1364, N1358, N68);
nor NOR2 (N1365, N1355, N157);
buf BUF1 (N1366, N1361);
or OR3 (N1367, N1350, N99, N516);
nor NOR3 (N1368, N1364, N388, N237);
and AND2 (N1369, N1360, N1293);
and AND4 (N1370, N1365, N1176, N793, N397);
xor XOR2 (N1371, N1357, N630);
xor XOR2 (N1372, N1368, N1322);
nor NOR4 (N1373, N1366, N577, N364, N352);
and AND3 (N1374, N1370, N1319, N251);
or OR4 (N1375, N1352, N222, N774, N1369);
buf BUF1 (N1376, N339);
and AND2 (N1377, N1375, N1329);
buf BUF1 (N1378, N1373);
not NOT1 (N1379, N1341);
xor XOR2 (N1380, N1378, N283);
xor XOR2 (N1381, N1371, N588);
xor XOR2 (N1382, N1374, N1329);
nor NOR4 (N1383, N1379, N164, N759, N688);
nand NAND3 (N1384, N1372, N798, N625);
and AND4 (N1385, N1383, N920, N86, N1167);
not NOT1 (N1386, N1367);
not NOT1 (N1387, N1363);
buf BUF1 (N1388, N1377);
or OR3 (N1389, N1387, N1027, N1053);
and AND2 (N1390, N1386, N1073);
not NOT1 (N1391, N1390);
xor XOR2 (N1392, N1389, N381);
not NOT1 (N1393, N1391);
buf BUF1 (N1394, N1392);
not NOT1 (N1395, N1382);
nand NAND3 (N1396, N1376, N117, N7);
xor XOR2 (N1397, N1394, N276);
not NOT1 (N1398, N1381);
xor XOR2 (N1399, N1380, N533);
nor NOR3 (N1400, N1385, N79, N294);
and AND3 (N1401, N1400, N802, N179);
not NOT1 (N1402, N1362);
nand NAND2 (N1403, N1393, N1349);
and AND2 (N1404, N1397, N981);
and AND3 (N1405, N1399, N426, N1099);
buf BUF1 (N1406, N1401);
or OR3 (N1407, N1395, N289, N927);
not NOT1 (N1408, N1396);
and AND4 (N1409, N1407, N1248, N1207, N1239);
or OR2 (N1410, N1406, N620);
nor NOR4 (N1411, N1408, N955, N1058, N676);
not NOT1 (N1412, N1398);
or OR2 (N1413, N1412, N1288);
or OR2 (N1414, N1402, N564);
buf BUF1 (N1415, N1403);
buf BUF1 (N1416, N1410);
buf BUF1 (N1417, N1414);
nor NOR2 (N1418, N1415, N1211);
nor NOR3 (N1419, N1416, N226, N1103);
not NOT1 (N1420, N1409);
xor XOR2 (N1421, N1388, N1188);
nand NAND4 (N1422, N1384, N1197, N1063, N997);
or OR3 (N1423, N1411, N524, N104);
and AND4 (N1424, N1413, N1028, N467, N1205);
xor XOR2 (N1425, N1420, N699);
nor NOR4 (N1426, N1417, N1001, N1093, N1339);
nand NAND2 (N1427, N1404, N1286);
or OR4 (N1428, N1418, N298, N1270, N406);
xor XOR2 (N1429, N1405, N231);
buf BUF1 (N1430, N1427);
and AND2 (N1431, N1425, N610);
xor XOR2 (N1432, N1431, N1141);
or OR2 (N1433, N1421, N562);
not NOT1 (N1434, N1423);
buf BUF1 (N1435, N1429);
or OR4 (N1436, N1419, N939, N923, N173);
buf BUF1 (N1437, N1432);
or OR3 (N1438, N1433, N303, N1402);
or OR2 (N1439, N1437, N849);
nand NAND2 (N1440, N1439, N934);
or OR4 (N1441, N1422, N333, N771, N1262);
nand NAND2 (N1442, N1426, N232);
nor NOR3 (N1443, N1435, N22, N179);
nor NOR4 (N1444, N1436, N846, N555, N693);
and AND2 (N1445, N1441, N466);
nor NOR4 (N1446, N1438, N469, N340, N411);
xor XOR2 (N1447, N1428, N7);
nor NOR3 (N1448, N1443, N482, N898);
nor NOR2 (N1449, N1424, N57);
nor NOR4 (N1450, N1430, N1236, N413, N382);
or OR3 (N1451, N1442, N791, N428);
or OR2 (N1452, N1434, N1198);
or OR2 (N1453, N1449, N212);
or OR4 (N1454, N1448, N1380, N651, N408);
nand NAND4 (N1455, N1444, N126, N420, N1314);
buf BUF1 (N1456, N1445);
not NOT1 (N1457, N1453);
nor NOR4 (N1458, N1457, N1456, N348, N1177);
nand NAND4 (N1459, N291, N11, N85, N214);
or OR4 (N1460, N1446, N461, N107, N1139);
nor NOR4 (N1461, N1459, N1180, N289, N579);
buf BUF1 (N1462, N1447);
nor NOR3 (N1463, N1455, N62, N1454);
xor XOR2 (N1464, N447, N360);
or OR3 (N1465, N1460, N786, N1144);
or OR4 (N1466, N1451, N993, N29, N7);
or OR2 (N1467, N1452, N730);
xor XOR2 (N1468, N1466, N325);
buf BUF1 (N1469, N1458);
not NOT1 (N1470, N1463);
and AND3 (N1471, N1440, N607, N973);
nor NOR4 (N1472, N1461, N695, N932, N742);
xor XOR2 (N1473, N1470, N801);
or OR4 (N1474, N1465, N87, N1194, N575);
xor XOR2 (N1475, N1467, N581);
or OR4 (N1476, N1472, N128, N1111, N291);
xor XOR2 (N1477, N1464, N1258);
or OR2 (N1478, N1462, N516);
not NOT1 (N1479, N1475);
nor NOR2 (N1480, N1476, N1034);
or OR3 (N1481, N1469, N1457, N755);
buf BUF1 (N1482, N1480);
buf BUF1 (N1483, N1478);
nand NAND3 (N1484, N1468, N846, N188);
xor XOR2 (N1485, N1479, N459);
nand NAND3 (N1486, N1482, N382, N234);
buf BUF1 (N1487, N1486);
xor XOR2 (N1488, N1471, N1414);
xor XOR2 (N1489, N1487, N622);
nor NOR3 (N1490, N1483, N453, N1249);
buf BUF1 (N1491, N1450);
buf BUF1 (N1492, N1484);
or OR2 (N1493, N1477, N577);
xor XOR2 (N1494, N1473, N570);
nor NOR2 (N1495, N1489, N1272);
or OR3 (N1496, N1481, N388, N977);
or OR4 (N1497, N1485, N1309, N1321, N355);
nor NOR3 (N1498, N1496, N1444, N1165);
buf BUF1 (N1499, N1491);
or OR4 (N1500, N1492, N1401, N372, N792);
buf BUF1 (N1501, N1500);
or OR3 (N1502, N1488, N97, N512);
nand NAND2 (N1503, N1493, N722);
buf BUF1 (N1504, N1502);
nor NOR3 (N1505, N1501, N719, N1283);
and AND3 (N1506, N1504, N1001, N339);
xor XOR2 (N1507, N1503, N699);
buf BUF1 (N1508, N1490);
xor XOR2 (N1509, N1494, N1141);
xor XOR2 (N1510, N1509, N1038);
nand NAND4 (N1511, N1508, N1286, N1443, N1060);
and AND4 (N1512, N1507, N770, N333, N503);
nor NOR2 (N1513, N1499, N1235);
nand NAND4 (N1514, N1474, N205, N565, N83);
xor XOR2 (N1515, N1510, N287);
and AND3 (N1516, N1498, N1358, N712);
buf BUF1 (N1517, N1497);
buf BUF1 (N1518, N1517);
and AND4 (N1519, N1495, N493, N686, N1279);
nor NOR3 (N1520, N1515, N839, N612);
or OR4 (N1521, N1512, N578, N157, N432);
and AND3 (N1522, N1519, N1181, N1233);
and AND3 (N1523, N1516, N238, N829);
or OR4 (N1524, N1522, N237, N1142, N1369);
and AND4 (N1525, N1506, N1468, N1414, N820);
nor NOR2 (N1526, N1513, N285);
and AND3 (N1527, N1505, N960, N314);
xor XOR2 (N1528, N1518, N725);
buf BUF1 (N1529, N1526);
not NOT1 (N1530, N1528);
buf BUF1 (N1531, N1530);
buf BUF1 (N1532, N1531);
and AND4 (N1533, N1511, N522, N1306, N1527);
nand NAND4 (N1534, N798, N675, N1385, N1420);
buf BUF1 (N1535, N1521);
or OR3 (N1536, N1532, N331, N158);
nor NOR2 (N1537, N1536, N1479);
nand NAND3 (N1538, N1535, N624, N97);
nor NOR3 (N1539, N1538, N1465, N1023);
xor XOR2 (N1540, N1537, N570);
or OR4 (N1541, N1529, N293, N673, N982);
nand NAND2 (N1542, N1520, N269);
or OR4 (N1543, N1534, N1381, N537, N1399);
nand NAND3 (N1544, N1533, N1518, N595);
buf BUF1 (N1545, N1523);
or OR3 (N1546, N1545, N1305, N264);
nand NAND3 (N1547, N1543, N1402, N1531);
and AND3 (N1548, N1525, N588, N467);
xor XOR2 (N1549, N1524, N1396);
xor XOR2 (N1550, N1547, N39);
not NOT1 (N1551, N1540);
and AND2 (N1552, N1548, N1091);
and AND3 (N1553, N1514, N99, N1058);
nand NAND2 (N1554, N1553, N561);
nor NOR3 (N1555, N1554, N803, N1436);
nand NAND3 (N1556, N1542, N310, N20);
nor NOR2 (N1557, N1552, N1449);
nor NOR4 (N1558, N1555, N778, N782, N190);
nor NOR3 (N1559, N1544, N1178, N1317);
and AND4 (N1560, N1546, N389, N1217, N103);
buf BUF1 (N1561, N1559);
nor NOR3 (N1562, N1557, N573, N719);
and AND4 (N1563, N1561, N648, N712, N1409);
nor NOR4 (N1564, N1550, N1518, N748, N371);
or OR4 (N1565, N1539, N1045, N245, N761);
or OR3 (N1566, N1560, N971, N939);
and AND4 (N1567, N1563, N679, N408, N1099);
nand NAND2 (N1568, N1541, N856);
buf BUF1 (N1569, N1551);
or OR2 (N1570, N1566, N196);
not NOT1 (N1571, N1564);
buf BUF1 (N1572, N1571);
xor XOR2 (N1573, N1568, N1295);
or OR4 (N1574, N1558, N1169, N1057, N178);
and AND3 (N1575, N1567, N741, N553);
nor NOR2 (N1576, N1573, N1203);
nand NAND3 (N1577, N1572, N714, N761);
not NOT1 (N1578, N1569);
nand NAND4 (N1579, N1562, N40, N171, N1424);
nor NOR2 (N1580, N1570, N1484);
and AND4 (N1581, N1578, N640, N720, N1283);
nand NAND4 (N1582, N1579, N389, N925, N638);
and AND4 (N1583, N1575, N1060, N531, N954);
nand NAND2 (N1584, N1580, N1446);
or OR2 (N1585, N1574, N1198);
not NOT1 (N1586, N1584);
and AND3 (N1587, N1577, N1498, N887);
not NOT1 (N1588, N1581);
or OR2 (N1589, N1556, N609);
nand NAND2 (N1590, N1589, N219);
or OR3 (N1591, N1586, N493, N1007);
nor NOR4 (N1592, N1587, N591, N1094, N22);
or OR4 (N1593, N1592, N1535, N812, N1297);
nor NOR3 (N1594, N1591, N1513, N971);
xor XOR2 (N1595, N1585, N973);
nand NAND4 (N1596, N1595, N273, N1122, N442);
or OR3 (N1597, N1565, N494, N203);
xor XOR2 (N1598, N1583, N1324);
or OR4 (N1599, N1590, N1578, N611, N27);
or OR2 (N1600, N1582, N1328);
or OR2 (N1601, N1596, N547);
nor NOR2 (N1602, N1599, N429);
xor XOR2 (N1603, N1601, N382);
or OR3 (N1604, N1602, N1237, N999);
nor NOR4 (N1605, N1598, N1464, N884, N1006);
buf BUF1 (N1606, N1588);
not NOT1 (N1607, N1597);
nand NAND4 (N1608, N1600, N803, N516, N314);
or OR4 (N1609, N1549, N880, N78, N565);
xor XOR2 (N1610, N1609, N523);
nand NAND2 (N1611, N1604, N674);
or OR2 (N1612, N1606, N326);
and AND4 (N1613, N1605, N1096, N1104, N942);
and AND4 (N1614, N1593, N1513, N963, N1061);
nand NAND3 (N1615, N1576, N389, N775);
buf BUF1 (N1616, N1594);
buf BUF1 (N1617, N1603);
nand NAND2 (N1618, N1614, N247);
not NOT1 (N1619, N1615);
xor XOR2 (N1620, N1617, N1406);
and AND2 (N1621, N1610, N1613);
and AND2 (N1622, N1593, N329);
or OR4 (N1623, N1620, N349, N1599, N1310);
buf BUF1 (N1624, N1623);
not NOT1 (N1625, N1618);
and AND2 (N1626, N1611, N812);
and AND4 (N1627, N1624, N253, N1539, N1078);
or OR3 (N1628, N1622, N1420, N353);
or OR2 (N1629, N1619, N382);
xor XOR2 (N1630, N1629, N290);
or OR2 (N1631, N1628, N303);
xor XOR2 (N1632, N1607, N22);
or OR2 (N1633, N1616, N771);
nand NAND2 (N1634, N1630, N1473);
xor XOR2 (N1635, N1626, N722);
or OR2 (N1636, N1625, N736);
and AND4 (N1637, N1632, N89, N916, N1482);
and AND4 (N1638, N1631, N862, N39, N1144);
or OR2 (N1639, N1637, N138);
and AND4 (N1640, N1627, N1336, N1405, N1544);
and AND2 (N1641, N1612, N206);
buf BUF1 (N1642, N1635);
and AND4 (N1643, N1642, N1540, N434, N1536);
buf BUF1 (N1644, N1639);
buf BUF1 (N1645, N1644);
or OR2 (N1646, N1641, N742);
nor NOR4 (N1647, N1643, N1286, N1278, N1229);
xor XOR2 (N1648, N1608, N998);
or OR2 (N1649, N1646, N1626);
and AND2 (N1650, N1647, N966);
buf BUF1 (N1651, N1636);
buf BUF1 (N1652, N1621);
and AND2 (N1653, N1649, N944);
nand NAND3 (N1654, N1633, N132, N445);
nor NOR4 (N1655, N1634, N307, N1273, N1520);
not NOT1 (N1656, N1638);
not NOT1 (N1657, N1648);
not NOT1 (N1658, N1656);
not NOT1 (N1659, N1645);
nand NAND2 (N1660, N1658, N1169);
nand NAND2 (N1661, N1652, N1180);
buf BUF1 (N1662, N1654);
nor NOR3 (N1663, N1662, N1219, N1421);
buf BUF1 (N1664, N1655);
or OR3 (N1665, N1661, N732, N803);
and AND3 (N1666, N1659, N364, N363);
buf BUF1 (N1667, N1653);
nor NOR2 (N1668, N1640, N1358);
buf BUF1 (N1669, N1668);
or OR4 (N1670, N1651, N933, N1024, N464);
or OR2 (N1671, N1657, N16);
xor XOR2 (N1672, N1665, N1138);
nor NOR2 (N1673, N1667, N1372);
nor NOR2 (N1674, N1666, N1052);
buf BUF1 (N1675, N1673);
xor XOR2 (N1676, N1675, N49);
or OR3 (N1677, N1669, N613, N499);
and AND4 (N1678, N1650, N800, N726, N618);
nand NAND4 (N1679, N1678, N310, N518, N316);
not NOT1 (N1680, N1679);
and AND3 (N1681, N1674, N1546, N1426);
nand NAND4 (N1682, N1676, N1662, N801, N610);
xor XOR2 (N1683, N1682, N1478);
not NOT1 (N1684, N1681);
buf BUF1 (N1685, N1677);
nor NOR4 (N1686, N1670, N586, N1611, N996);
xor XOR2 (N1687, N1664, N976);
not NOT1 (N1688, N1686);
not NOT1 (N1689, N1672);
nor NOR3 (N1690, N1684, N838, N905);
nand NAND4 (N1691, N1689, N1209, N53, N1307);
buf BUF1 (N1692, N1683);
xor XOR2 (N1693, N1663, N662);
not NOT1 (N1694, N1691);
nor NOR4 (N1695, N1693, N86, N788, N1022);
or OR2 (N1696, N1690, N1076);
not NOT1 (N1697, N1692);
or OR3 (N1698, N1697, N978, N856);
xor XOR2 (N1699, N1660, N439);
nor NOR2 (N1700, N1688, N821);
or OR4 (N1701, N1687, N539, N1193, N707);
and AND2 (N1702, N1700, N1617);
buf BUF1 (N1703, N1694);
xor XOR2 (N1704, N1671, N410);
buf BUF1 (N1705, N1680);
or OR4 (N1706, N1705, N663, N631, N353);
nor NOR3 (N1707, N1695, N593, N431);
nand NAND3 (N1708, N1704, N1259, N1295);
buf BUF1 (N1709, N1698);
and AND4 (N1710, N1685, N53, N207, N591);
xor XOR2 (N1711, N1701, N151);
nor NOR4 (N1712, N1699, N709, N1154, N591);
buf BUF1 (N1713, N1708);
nand NAND4 (N1714, N1706, N738, N394, N621);
xor XOR2 (N1715, N1703, N116);
nand NAND4 (N1716, N1712, N1632, N1611, N37);
xor XOR2 (N1717, N1713, N1270);
or OR3 (N1718, N1714, N9, N1544);
not NOT1 (N1719, N1696);
buf BUF1 (N1720, N1718);
nand NAND3 (N1721, N1719, N155, N795);
or OR2 (N1722, N1711, N1060);
or OR2 (N1723, N1710, N1226);
xor XOR2 (N1724, N1716, N1175);
and AND4 (N1725, N1721, N809, N76, N1701);
xor XOR2 (N1726, N1702, N1523);
not NOT1 (N1727, N1717);
xor XOR2 (N1728, N1715, N15);
nor NOR4 (N1729, N1709, N1361, N943, N336);
buf BUF1 (N1730, N1724);
not NOT1 (N1731, N1723);
xor XOR2 (N1732, N1707, N1715);
or OR4 (N1733, N1726, N1065, N11, N137);
not NOT1 (N1734, N1725);
and AND4 (N1735, N1722, N586, N964, N797);
buf BUF1 (N1736, N1730);
not NOT1 (N1737, N1732);
and AND2 (N1738, N1734, N1357);
nand NAND3 (N1739, N1729, N346, N968);
not NOT1 (N1740, N1737);
xor XOR2 (N1741, N1727, N1094);
nand NAND4 (N1742, N1731, N687, N557, N184);
nand NAND2 (N1743, N1728, N1083);
xor XOR2 (N1744, N1736, N645);
nand NAND3 (N1745, N1743, N828, N493);
not NOT1 (N1746, N1741);
nand NAND4 (N1747, N1744, N512, N1224, N1722);
not NOT1 (N1748, N1745);
or OR4 (N1749, N1739, N1165, N189, N284);
xor XOR2 (N1750, N1749, N315);
nor NOR2 (N1751, N1746, N159);
and AND3 (N1752, N1742, N1521, N275);
and AND2 (N1753, N1751, N1467);
nor NOR3 (N1754, N1735, N941, N798);
xor XOR2 (N1755, N1738, N361);
or OR2 (N1756, N1720, N159);
xor XOR2 (N1757, N1755, N1274);
nor NOR2 (N1758, N1754, N6);
or OR3 (N1759, N1733, N1317, N194);
xor XOR2 (N1760, N1740, N1506);
buf BUF1 (N1761, N1748);
and AND2 (N1762, N1750, N301);
xor XOR2 (N1763, N1760, N1105);
not NOT1 (N1764, N1761);
and AND3 (N1765, N1758, N531, N1578);
and AND2 (N1766, N1757, N886);
nand NAND4 (N1767, N1747, N1315, N661, N737);
xor XOR2 (N1768, N1766, N252);
not NOT1 (N1769, N1767);
xor XOR2 (N1770, N1756, N1121);
xor XOR2 (N1771, N1763, N1465);
xor XOR2 (N1772, N1762, N664);
nand NAND2 (N1773, N1764, N685);
and AND4 (N1774, N1773, N433, N1066, N1174);
not NOT1 (N1775, N1753);
or OR4 (N1776, N1775, N1559, N767, N526);
xor XOR2 (N1777, N1768, N916);
buf BUF1 (N1778, N1765);
buf BUF1 (N1779, N1771);
nor NOR3 (N1780, N1777, N1727, N910);
not NOT1 (N1781, N1780);
nand NAND4 (N1782, N1778, N1010, N606, N1631);
not NOT1 (N1783, N1782);
or OR4 (N1784, N1783, N1708, N743, N1630);
nor NOR3 (N1785, N1776, N515, N450);
or OR4 (N1786, N1770, N1365, N1038, N835);
not NOT1 (N1787, N1769);
not NOT1 (N1788, N1785);
or OR4 (N1789, N1786, N126, N1092, N1175);
xor XOR2 (N1790, N1774, N974);
and AND4 (N1791, N1772, N530, N941, N1695);
nand NAND4 (N1792, N1752, N600, N1440, N1130);
nor NOR2 (N1793, N1789, N1303);
nor NOR3 (N1794, N1790, N214, N1451);
not NOT1 (N1795, N1791);
and AND4 (N1796, N1793, N1599, N1265, N565);
xor XOR2 (N1797, N1788, N1020);
xor XOR2 (N1798, N1796, N241);
nor NOR3 (N1799, N1792, N1143, N397);
nor NOR3 (N1800, N1779, N639, N1780);
xor XOR2 (N1801, N1798, N1419);
nand NAND3 (N1802, N1794, N701, N706);
xor XOR2 (N1803, N1799, N1529);
buf BUF1 (N1804, N1803);
xor XOR2 (N1805, N1802, N580);
not NOT1 (N1806, N1804);
buf BUF1 (N1807, N1800);
and AND2 (N1808, N1784, N106);
nand NAND4 (N1809, N1806, N1497, N64, N1248);
or OR3 (N1810, N1805, N37, N270);
nor NOR2 (N1811, N1787, N1192);
not NOT1 (N1812, N1795);
or OR2 (N1813, N1810, N813);
or OR3 (N1814, N1797, N489, N1528);
xor XOR2 (N1815, N1759, N114);
buf BUF1 (N1816, N1812);
xor XOR2 (N1817, N1809, N928);
nor NOR3 (N1818, N1817, N139, N1128);
nor NOR4 (N1819, N1818, N888, N1102, N927);
nand NAND4 (N1820, N1814, N477, N439, N425);
nor NOR2 (N1821, N1781, N1529);
nand NAND2 (N1822, N1820, N1486);
nor NOR3 (N1823, N1801, N550, N883);
not NOT1 (N1824, N1822);
not NOT1 (N1825, N1813);
nand NAND3 (N1826, N1825, N937, N111);
buf BUF1 (N1827, N1823);
and AND2 (N1828, N1824, N1438);
not NOT1 (N1829, N1826);
not NOT1 (N1830, N1815);
and AND4 (N1831, N1829, N1731, N1464, N193);
not NOT1 (N1832, N1821);
not NOT1 (N1833, N1830);
not NOT1 (N1834, N1819);
and AND2 (N1835, N1807, N1088);
nand NAND3 (N1836, N1828, N988, N1033);
buf BUF1 (N1837, N1827);
buf BUF1 (N1838, N1816);
buf BUF1 (N1839, N1835);
not NOT1 (N1840, N1839);
nand NAND3 (N1841, N1831, N1171, N94);
nand NAND2 (N1842, N1837, N410);
buf BUF1 (N1843, N1842);
nand NAND4 (N1844, N1808, N182, N1211, N1416);
or OR4 (N1845, N1841, N1148, N1330, N987);
nand NAND2 (N1846, N1838, N997);
xor XOR2 (N1847, N1832, N739);
nand NAND2 (N1848, N1844, N412);
xor XOR2 (N1849, N1834, N970);
and AND3 (N1850, N1811, N844, N1718);
nand NAND3 (N1851, N1849, N179, N359);
not NOT1 (N1852, N1848);
nand NAND2 (N1853, N1846, N192);
nor NOR3 (N1854, N1850, N368, N1402);
and AND4 (N1855, N1833, N1158, N1359, N1071);
and AND3 (N1856, N1852, N182, N1032);
not NOT1 (N1857, N1854);
not NOT1 (N1858, N1855);
xor XOR2 (N1859, N1853, N1717);
or OR2 (N1860, N1845, N237);
xor XOR2 (N1861, N1847, N249);
xor XOR2 (N1862, N1856, N1020);
not NOT1 (N1863, N1858);
and AND3 (N1864, N1836, N1723, N1069);
nor NOR4 (N1865, N1859, N1093, N861, N973);
buf BUF1 (N1866, N1857);
not NOT1 (N1867, N1866);
or OR2 (N1868, N1851, N1424);
nor NOR3 (N1869, N1861, N749, N647);
not NOT1 (N1870, N1860);
buf BUF1 (N1871, N1862);
nand NAND4 (N1872, N1863, N1434, N708, N1113);
nand NAND2 (N1873, N1840, N1527);
xor XOR2 (N1874, N1865, N1448);
nor NOR3 (N1875, N1867, N1744, N1167);
not NOT1 (N1876, N1871);
xor XOR2 (N1877, N1874, N58);
nor NOR4 (N1878, N1873, N293, N1454, N1638);
and AND3 (N1879, N1843, N112, N1506);
or OR3 (N1880, N1864, N232, N1626);
not NOT1 (N1881, N1870);
buf BUF1 (N1882, N1878);
xor XOR2 (N1883, N1881, N608);
nand NAND2 (N1884, N1883, N1509);
nand NAND3 (N1885, N1882, N221, N1180);
xor XOR2 (N1886, N1876, N690);
xor XOR2 (N1887, N1885, N916);
not NOT1 (N1888, N1880);
nor NOR4 (N1889, N1888, N209, N891, N212);
nor NOR2 (N1890, N1887, N556);
xor XOR2 (N1891, N1879, N421);
buf BUF1 (N1892, N1890);
and AND2 (N1893, N1869, N377);
xor XOR2 (N1894, N1872, N781);
nor NOR2 (N1895, N1886, N474);
buf BUF1 (N1896, N1895);
not NOT1 (N1897, N1884);
not NOT1 (N1898, N1889);
or OR2 (N1899, N1875, N1804);
and AND3 (N1900, N1877, N99, N1505);
not NOT1 (N1901, N1899);
xor XOR2 (N1902, N1891, N1378);
xor XOR2 (N1903, N1902, N690);
nand NAND2 (N1904, N1893, N312);
nand NAND2 (N1905, N1898, N1398);
and AND2 (N1906, N1868, N295);
buf BUF1 (N1907, N1904);
xor XOR2 (N1908, N1903, N62);
nor NOR4 (N1909, N1908, N218, N876, N1345);
and AND4 (N1910, N1909, N1029, N1872, N62);
xor XOR2 (N1911, N1892, N844);
and AND2 (N1912, N1911, N977);
xor XOR2 (N1913, N1894, N1707);
nand NAND4 (N1914, N1906, N319, N1800, N1864);
nand NAND4 (N1915, N1913, N160, N1761, N1774);
or OR3 (N1916, N1914, N1341, N1158);
not NOT1 (N1917, N1900);
nand NAND3 (N1918, N1907, N1729, N1679);
nand NAND2 (N1919, N1910, N1367);
nand NAND2 (N1920, N1912, N391);
and AND2 (N1921, N1896, N165);
or OR4 (N1922, N1917, N876, N1756, N1307);
nand NAND4 (N1923, N1905, N1746, N1828, N621);
and AND4 (N1924, N1897, N538, N1025, N193);
and AND4 (N1925, N1901, N1374, N464, N1425);
buf BUF1 (N1926, N1919);
xor XOR2 (N1927, N1926, N1534);
or OR3 (N1928, N1923, N1339, N888);
or OR3 (N1929, N1927, N618, N782);
nor NOR2 (N1930, N1915, N723);
not NOT1 (N1931, N1922);
xor XOR2 (N1932, N1928, N1092);
nor NOR3 (N1933, N1925, N293, N1673);
buf BUF1 (N1934, N1929);
buf BUF1 (N1935, N1924);
nand NAND2 (N1936, N1921, N634);
xor XOR2 (N1937, N1930, N440);
or OR4 (N1938, N1920, N1040, N1517, N629);
not NOT1 (N1939, N1918);
and AND4 (N1940, N1935, N280, N919, N1748);
xor XOR2 (N1941, N1933, N605);
buf BUF1 (N1942, N1937);
buf BUF1 (N1943, N1936);
buf BUF1 (N1944, N1916);
xor XOR2 (N1945, N1932, N560);
or OR2 (N1946, N1943, N1858);
nand NAND4 (N1947, N1931, N814, N1796, N129);
buf BUF1 (N1948, N1947);
nand NAND4 (N1949, N1940, N1492, N1531, N1905);
nand NAND4 (N1950, N1945, N1753, N1908, N1875);
or OR3 (N1951, N1950, N403, N483);
nor NOR4 (N1952, N1939, N1061, N397, N694);
nor NOR3 (N1953, N1952, N1843, N475);
not NOT1 (N1954, N1941);
xor XOR2 (N1955, N1948, N673);
not NOT1 (N1956, N1946);
buf BUF1 (N1957, N1942);
nand NAND4 (N1958, N1954, N437, N305, N1445);
or OR2 (N1959, N1957, N1460);
and AND4 (N1960, N1955, N336, N1475, N1806);
not NOT1 (N1961, N1944);
or OR3 (N1962, N1956, N1528, N1070);
nor NOR2 (N1963, N1961, N562);
buf BUF1 (N1964, N1963);
xor XOR2 (N1965, N1960, N822);
xor XOR2 (N1966, N1934, N86);
nor NOR3 (N1967, N1964, N1578, N242);
or OR3 (N1968, N1953, N1945, N1751);
buf BUF1 (N1969, N1962);
not NOT1 (N1970, N1967);
not NOT1 (N1971, N1969);
not NOT1 (N1972, N1938);
buf BUF1 (N1973, N1968);
nor NOR2 (N1974, N1951, N246);
not NOT1 (N1975, N1958);
or OR4 (N1976, N1966, N923, N633, N1430);
nor NOR4 (N1977, N1965, N579, N578, N1237);
or OR3 (N1978, N1970, N65, N1852);
not NOT1 (N1979, N1972);
nand NAND4 (N1980, N1973, N1141, N329, N553);
nor NOR3 (N1981, N1975, N1079, N808);
buf BUF1 (N1982, N1979);
nor NOR4 (N1983, N1981, N1915, N196, N713);
not NOT1 (N1984, N1978);
and AND4 (N1985, N1971, N1682, N1726, N651);
xor XOR2 (N1986, N1974, N1448);
not NOT1 (N1987, N1959);
and AND2 (N1988, N1983, N1889);
nand NAND2 (N1989, N1984, N1281);
xor XOR2 (N1990, N1976, N282);
xor XOR2 (N1991, N1985, N974);
and AND4 (N1992, N1988, N909, N827, N83);
buf BUF1 (N1993, N1991);
not NOT1 (N1994, N1982);
or OR2 (N1995, N1980, N1369);
not NOT1 (N1996, N1986);
nor NOR2 (N1997, N1992, N1883);
nand NAND4 (N1998, N1989, N194, N562, N909);
xor XOR2 (N1999, N1993, N535);
and AND2 (N2000, N1990, N397);
and AND2 (N2001, N1994, N636);
buf BUF1 (N2002, N1999);
not NOT1 (N2003, N1987);
nand NAND2 (N2004, N2002, N966);
not NOT1 (N2005, N1998);
and AND3 (N2006, N1996, N1614, N917);
nor NOR4 (N2007, N2003, N1487, N5, N194);
not NOT1 (N2008, N1949);
not NOT1 (N2009, N1997);
and AND2 (N2010, N2006, N320);
xor XOR2 (N2011, N2000, N479);
buf BUF1 (N2012, N2001);
and AND2 (N2013, N2005, N1190);
and AND4 (N2014, N2008, N1761, N399, N41);
nand NAND3 (N2015, N2011, N895, N945);
and AND2 (N2016, N2007, N1242);
or OR3 (N2017, N2009, N1393, N522);
or OR3 (N2018, N1995, N1085, N1450);
nor NOR2 (N2019, N2018, N567);
xor XOR2 (N2020, N2016, N659);
nor NOR2 (N2021, N2004, N1709);
buf BUF1 (N2022, N2020);
nor NOR4 (N2023, N2017, N353, N1329, N381);
or OR3 (N2024, N2021, N381, N147);
xor XOR2 (N2025, N2019, N937);
nand NAND2 (N2026, N2015, N543);
not NOT1 (N2027, N2013);
buf BUF1 (N2028, N1977);
nand NAND2 (N2029, N2027, N1154);
nand NAND3 (N2030, N2026, N993, N1031);
not NOT1 (N2031, N2010);
nand NAND3 (N2032, N2028, N374, N241);
nor NOR3 (N2033, N2029, N1491, N1381);
or OR4 (N2034, N2023, N105, N82, N1840);
xor XOR2 (N2035, N2030, N987);
buf BUF1 (N2036, N2034);
nor NOR2 (N2037, N2025, N948);
or OR2 (N2038, N2033, N701);
buf BUF1 (N2039, N2012);
not NOT1 (N2040, N2037);
nor NOR3 (N2041, N2038, N1478, N1654);
not NOT1 (N2042, N2032);
nor NOR2 (N2043, N2024, N1455);
and AND2 (N2044, N2042, N832);
xor XOR2 (N2045, N2044, N1481);
and AND4 (N2046, N2036, N1006, N1586, N640);
or OR4 (N2047, N2031, N1966, N1103, N505);
not NOT1 (N2048, N2041);
nand NAND3 (N2049, N2045, N767, N1127);
buf BUF1 (N2050, N2040);
buf BUF1 (N2051, N2043);
or OR2 (N2052, N2049, N431);
and AND3 (N2053, N2047, N1566, N1082);
and AND3 (N2054, N2048, N1139, N1982);
or OR2 (N2055, N2050, N347);
and AND2 (N2056, N2052, N1890);
xor XOR2 (N2057, N2046, N1559);
nand NAND3 (N2058, N2056, N2027, N583);
nor NOR4 (N2059, N2014, N1317, N1212, N256);
buf BUF1 (N2060, N2059);
xor XOR2 (N2061, N2039, N395);
and AND2 (N2062, N2057, N1059);
nor NOR2 (N2063, N2054, N1925);
xor XOR2 (N2064, N2035, N209);
nand NAND2 (N2065, N2063, N1834);
and AND3 (N2066, N2022, N81, N1131);
nand NAND2 (N2067, N2064, N1345);
not NOT1 (N2068, N2065);
buf BUF1 (N2069, N2051);
or OR4 (N2070, N2066, N733, N1594, N1008);
nand NAND4 (N2071, N2067, N600, N402, N919);
buf BUF1 (N2072, N2060);
xor XOR2 (N2073, N2070, N1917);
and AND4 (N2074, N2055, N995, N727, N108);
nand NAND4 (N2075, N2053, N393, N1090, N92);
buf BUF1 (N2076, N2058);
and AND2 (N2077, N2069, N668);
not NOT1 (N2078, N2073);
not NOT1 (N2079, N2072);
xor XOR2 (N2080, N2071, N802);
nand NAND2 (N2081, N2075, N1856);
and AND2 (N2082, N2080, N1112);
not NOT1 (N2083, N2078);
nor NOR3 (N2084, N2081, N730, N431);
and AND2 (N2085, N2084, N1203);
and AND4 (N2086, N2082, N347, N1058, N972);
nor NOR4 (N2087, N2068, N596, N1406, N1470);
nor NOR3 (N2088, N2077, N729, N1953);
nor NOR2 (N2089, N2086, N831);
buf BUF1 (N2090, N2088);
xor XOR2 (N2091, N2062, N166);
and AND3 (N2092, N2076, N1676, N2070);
nor NOR3 (N2093, N2090, N1241, N1603);
nor NOR4 (N2094, N2089, N1478, N1757, N795);
or OR4 (N2095, N2091, N1069, N102, N450);
xor XOR2 (N2096, N2079, N1083);
and AND3 (N2097, N2085, N859, N995);
or OR2 (N2098, N2087, N198);
or OR4 (N2099, N2093, N1436, N1040, N1513);
and AND4 (N2100, N2097, N1695, N2041, N1979);
xor XOR2 (N2101, N2099, N1932);
xor XOR2 (N2102, N2061, N368);
not NOT1 (N2103, N2096);
buf BUF1 (N2104, N2100);
xor XOR2 (N2105, N2101, N120);
and AND2 (N2106, N2102, N373);
not NOT1 (N2107, N2103);
or OR4 (N2108, N2094, N1520, N1798, N1938);
not NOT1 (N2109, N2083);
and AND4 (N2110, N2092, N1313, N906, N967);
xor XOR2 (N2111, N2106, N1362);
not NOT1 (N2112, N2109);
or OR3 (N2113, N2074, N853, N1088);
nor NOR2 (N2114, N2113, N838);
buf BUF1 (N2115, N2095);
xor XOR2 (N2116, N2098, N1432);
buf BUF1 (N2117, N2107);
nor NOR4 (N2118, N2105, N591, N367, N1117);
nor NOR2 (N2119, N2108, N504);
nand NAND4 (N2120, N2116, N1819, N558, N1470);
xor XOR2 (N2121, N2110, N2031);
not NOT1 (N2122, N2115);
nor NOR2 (N2123, N2114, N684);
nand NAND3 (N2124, N2123, N1049, N788);
nor NOR2 (N2125, N2104, N1996);
and AND2 (N2126, N2121, N1898);
nor NOR2 (N2127, N2124, N814);
nor NOR3 (N2128, N2111, N1631, N101);
nor NOR2 (N2129, N2112, N1855);
nand NAND3 (N2130, N2120, N227, N568);
not NOT1 (N2131, N2122);
nor NOR4 (N2132, N2117, N948, N1799, N1422);
xor XOR2 (N2133, N2128, N1781);
buf BUF1 (N2134, N2131);
and AND4 (N2135, N2129, N90, N1472, N290);
or OR4 (N2136, N2133, N466, N52, N1790);
and AND4 (N2137, N2136, N106, N588, N1679);
nor NOR3 (N2138, N2134, N634, N583);
buf BUF1 (N2139, N2135);
nand NAND2 (N2140, N2139, N1532);
nor NOR2 (N2141, N2137, N275);
xor XOR2 (N2142, N2127, N1202);
not NOT1 (N2143, N2126);
buf BUF1 (N2144, N2142);
nand NAND4 (N2145, N2140, N129, N1658, N902);
nor NOR4 (N2146, N2130, N1921, N1729, N1679);
and AND3 (N2147, N2146, N1177, N1733);
or OR2 (N2148, N2141, N1241);
and AND3 (N2149, N2145, N232, N1267);
xor XOR2 (N2150, N2125, N719);
xor XOR2 (N2151, N2132, N300);
nand NAND4 (N2152, N2151, N1489, N1743, N970);
xor XOR2 (N2153, N2152, N1980);
nand NAND2 (N2154, N2143, N1826);
not NOT1 (N2155, N2144);
and AND4 (N2156, N2118, N627, N954, N624);
nand NAND4 (N2157, N2155, N1043, N33, N1339);
nor NOR3 (N2158, N2147, N937, N1090);
and AND4 (N2159, N2150, N975, N949, N2091);
buf BUF1 (N2160, N2158);
or OR3 (N2161, N2119, N141, N701);
nand NAND3 (N2162, N2148, N1822, N1849);
not NOT1 (N2163, N2156);
or OR3 (N2164, N2160, N1684, N473);
xor XOR2 (N2165, N2138, N431);
nor NOR3 (N2166, N2149, N1051, N841);
or OR4 (N2167, N2163, N351, N1272, N744);
not NOT1 (N2168, N2161);
or OR3 (N2169, N2157, N492, N2014);
xor XOR2 (N2170, N2159, N1511);
buf BUF1 (N2171, N2170);
xor XOR2 (N2172, N2164, N598);
nor NOR4 (N2173, N2168, N470, N1516, N959);
nor NOR4 (N2174, N2171, N1146, N1346, N1127);
not NOT1 (N2175, N2169);
nor NOR3 (N2176, N2165, N1591, N290);
xor XOR2 (N2177, N2166, N1674);
not NOT1 (N2178, N2172);
and AND3 (N2179, N2153, N1700, N1715);
nand NAND2 (N2180, N2179, N1384);
buf BUF1 (N2181, N2174);
and AND3 (N2182, N2154, N1702, N1297);
xor XOR2 (N2183, N2173, N1724);
and AND3 (N2184, N2167, N426, N893);
nor NOR4 (N2185, N2181, N1160, N1367, N62);
or OR2 (N2186, N2175, N493);
nand NAND4 (N2187, N2162, N1059, N1717, N1961);
nand NAND2 (N2188, N2180, N1556);
xor XOR2 (N2189, N2184, N1226);
buf BUF1 (N2190, N2185);
nor NOR2 (N2191, N2190, N1565);
xor XOR2 (N2192, N2189, N282);
buf BUF1 (N2193, N2183);
xor XOR2 (N2194, N2188, N919);
nor NOR3 (N2195, N2186, N479, N813);
not NOT1 (N2196, N2176);
not NOT1 (N2197, N2177);
not NOT1 (N2198, N2178);
not NOT1 (N2199, N2187);
or OR3 (N2200, N2196, N51, N609);
xor XOR2 (N2201, N2197, N355);
and AND4 (N2202, N2198, N147, N272, N28);
and AND2 (N2203, N2182, N1191);
xor XOR2 (N2204, N2192, N608);
buf BUF1 (N2205, N2201);
not NOT1 (N2206, N2199);
and AND2 (N2207, N2202, N511);
xor XOR2 (N2208, N2191, N698);
nand NAND4 (N2209, N2194, N663, N2052, N26);
and AND4 (N2210, N2209, N1250, N43, N954);
or OR3 (N2211, N2205, N1345, N65);
xor XOR2 (N2212, N2210, N1325);
nor NOR2 (N2213, N2208, N324);
not NOT1 (N2214, N2206);
or OR2 (N2215, N2214, N1578);
and AND2 (N2216, N2211, N1418);
buf BUF1 (N2217, N2204);
buf BUF1 (N2218, N2215);
buf BUF1 (N2219, N2193);
nand NAND2 (N2220, N2213, N1244);
nor NOR3 (N2221, N2200, N1058, N373);
nor NOR3 (N2222, N2207, N23, N195);
not NOT1 (N2223, N2221);
buf BUF1 (N2224, N2218);
nor NOR3 (N2225, N2220, N777, N1052);
or OR2 (N2226, N2216, N603);
not NOT1 (N2227, N2225);
or OR2 (N2228, N2226, N253);
buf BUF1 (N2229, N2217);
nor NOR2 (N2230, N2219, N446);
and AND2 (N2231, N2223, N1431);
buf BUF1 (N2232, N2230);
nor NOR3 (N2233, N2228, N250, N1101);
and AND4 (N2234, N2212, N775, N581, N654);
or OR2 (N2235, N2222, N2107);
and AND4 (N2236, N2229, N1006, N958, N1890);
xor XOR2 (N2237, N2235, N1332);
nand NAND4 (N2238, N2231, N1061, N1105, N2221);
nor NOR4 (N2239, N2233, N2213, N1529, N200);
not NOT1 (N2240, N2236);
and AND2 (N2241, N2237, N1282);
buf BUF1 (N2242, N2232);
nand NAND2 (N2243, N2203, N1221);
or OR2 (N2244, N2238, N577);
and AND3 (N2245, N2241, N240, N2072);
or OR2 (N2246, N2242, N1205);
xor XOR2 (N2247, N2227, N666);
xor XOR2 (N2248, N2224, N527);
nand NAND4 (N2249, N2244, N1046, N449, N2070);
nor NOR2 (N2250, N2195, N1028);
or OR3 (N2251, N2249, N712, N1151);
nor NOR2 (N2252, N2251, N1168);
nand NAND3 (N2253, N2240, N1519, N705);
and AND4 (N2254, N2239, N1119, N2060, N2146);
nand NAND4 (N2255, N2248, N140, N549, N149);
and AND2 (N2256, N2255, N1807);
xor XOR2 (N2257, N2247, N1867);
not NOT1 (N2258, N2243);
nor NOR3 (N2259, N2256, N1450, N293);
or OR4 (N2260, N2259, N1528, N771, N2079);
or OR4 (N2261, N2253, N538, N549, N725);
xor XOR2 (N2262, N2250, N1267);
buf BUF1 (N2263, N2246);
buf BUF1 (N2264, N2258);
and AND2 (N2265, N2260, N1431);
and AND4 (N2266, N2261, N1774, N1982, N1672);
and AND4 (N2267, N2262, N622, N794, N765);
nand NAND3 (N2268, N2265, N788, N522);
not NOT1 (N2269, N2268);
or OR4 (N2270, N2266, N676, N659, N56);
xor XOR2 (N2271, N2245, N1615);
xor XOR2 (N2272, N2252, N75);
or OR3 (N2273, N2234, N1890, N908);
buf BUF1 (N2274, N2271);
or OR3 (N2275, N2263, N1912, N538);
nor NOR3 (N2276, N2257, N83, N1992);
or OR2 (N2277, N2276, N169);
and AND3 (N2278, N2274, N1775, N240);
nand NAND2 (N2279, N2264, N1693);
or OR4 (N2280, N2267, N178, N1220, N1757);
not NOT1 (N2281, N2270);
nor NOR4 (N2282, N2280, N245, N2047, N320);
or OR4 (N2283, N2277, N1979, N1215, N1212);
xor XOR2 (N2284, N2254, N1784);
buf BUF1 (N2285, N2281);
nand NAND2 (N2286, N2282, N95);
nand NAND3 (N2287, N2286, N520, N874);
or OR4 (N2288, N2283, N63, N1851, N2059);
buf BUF1 (N2289, N2278);
nor NOR3 (N2290, N2289, N1535, N514);
nand NAND4 (N2291, N2290, N959, N62, N25);
and AND2 (N2292, N2284, N1882);
not NOT1 (N2293, N2285);
buf BUF1 (N2294, N2279);
nor NOR3 (N2295, N2294, N2224, N2278);
buf BUF1 (N2296, N2272);
not NOT1 (N2297, N2287);
buf BUF1 (N2298, N2269);
or OR3 (N2299, N2298, N1314, N1908);
not NOT1 (N2300, N2292);
nand NAND4 (N2301, N2296, N2110, N851, N1031);
nand NAND4 (N2302, N2275, N815, N1774, N80);
or OR3 (N2303, N2293, N43, N1203);
xor XOR2 (N2304, N2297, N1265);
or OR3 (N2305, N2303, N1217, N1287);
nand NAND3 (N2306, N2299, N673, N2039);
xor XOR2 (N2307, N2302, N1725);
xor XOR2 (N2308, N2304, N782);
or OR4 (N2309, N2300, N794, N1018, N1775);
nand NAND4 (N2310, N2291, N165, N2218, N1657);
nor NOR2 (N2311, N2288, N2270);
nand NAND3 (N2312, N2311, N870, N1965);
or OR4 (N2313, N2273, N1887, N711, N769);
or OR3 (N2314, N2305, N532, N405);
nand NAND2 (N2315, N2309, N1283);
xor XOR2 (N2316, N2307, N1574);
not NOT1 (N2317, N2308);
not NOT1 (N2318, N2295);
nand NAND4 (N2319, N2313, N161, N866, N1884);
nand NAND3 (N2320, N2317, N1551, N1390);
xor XOR2 (N2321, N2315, N274);
or OR4 (N2322, N2318, N1261, N2216, N2115);
not NOT1 (N2323, N2321);
nor NOR4 (N2324, N2301, N2234, N1269, N389);
and AND3 (N2325, N2319, N673, N1566);
buf BUF1 (N2326, N2314);
buf BUF1 (N2327, N2316);
xor XOR2 (N2328, N2326, N1571);
not NOT1 (N2329, N2323);
nand NAND3 (N2330, N2306, N59, N2161);
buf BUF1 (N2331, N2324);
and AND3 (N2332, N2328, N1816, N614);
or OR4 (N2333, N2327, N1390, N463, N2210);
xor XOR2 (N2334, N2320, N34);
buf BUF1 (N2335, N2334);
or OR2 (N2336, N2322, N903);
buf BUF1 (N2337, N2329);
not NOT1 (N2338, N2333);
xor XOR2 (N2339, N2330, N474);
buf BUF1 (N2340, N2336);
not NOT1 (N2341, N2325);
buf BUF1 (N2342, N2312);
not NOT1 (N2343, N2339);
and AND2 (N2344, N2343, N1480);
nor NOR4 (N2345, N2335, N1581, N587, N2219);
buf BUF1 (N2346, N2344);
and AND4 (N2347, N2340, N801, N882, N2292);
or OR3 (N2348, N2331, N2202, N1073);
and AND2 (N2349, N2342, N142);
or OR3 (N2350, N2346, N641, N605);
or OR3 (N2351, N2349, N1851, N540);
and AND4 (N2352, N2350, N1158, N1293, N1360);
nor NOR2 (N2353, N2332, N498);
buf BUF1 (N2354, N2353);
not NOT1 (N2355, N2341);
nand NAND2 (N2356, N2348, N1353);
buf BUF1 (N2357, N2337);
or OR4 (N2358, N2351, N1325, N1546, N2256);
not NOT1 (N2359, N2352);
nand NAND2 (N2360, N2347, N953);
and AND2 (N2361, N2354, N316);
or OR4 (N2362, N2355, N1710, N330, N2217);
and AND3 (N2363, N2362, N1231, N787);
nand NAND2 (N2364, N2310, N174);
and AND2 (N2365, N2357, N375);
xor XOR2 (N2366, N2363, N428);
buf BUF1 (N2367, N2364);
and AND4 (N2368, N2358, N1163, N441, N364);
buf BUF1 (N2369, N2360);
xor XOR2 (N2370, N2367, N199);
buf BUF1 (N2371, N2361);
buf BUF1 (N2372, N2369);
not NOT1 (N2373, N2366);
or OR4 (N2374, N2371, N789, N623, N1070);
xor XOR2 (N2375, N2359, N117);
and AND4 (N2376, N2375, N2047, N1728, N1135);
buf BUF1 (N2377, N2372);
or OR4 (N2378, N2370, N1080, N2162, N1562);
nor NOR2 (N2379, N2376, N246);
buf BUF1 (N2380, N2345);
xor XOR2 (N2381, N2356, N199);
and AND2 (N2382, N2338, N1951);
or OR3 (N2383, N2374, N505, N481);
and AND3 (N2384, N2377, N455, N2353);
and AND3 (N2385, N2373, N1342, N2016);
xor XOR2 (N2386, N2379, N1036);
nand NAND2 (N2387, N2368, N1151);
or OR2 (N2388, N2381, N206);
nor NOR2 (N2389, N2387, N337);
xor XOR2 (N2390, N2365, N2015);
nor NOR2 (N2391, N2385, N1609);
nor NOR4 (N2392, N2389, N1729, N798, N1795);
buf BUF1 (N2393, N2392);
nor NOR3 (N2394, N2393, N579, N1377);
buf BUF1 (N2395, N2384);
buf BUF1 (N2396, N2391);
buf BUF1 (N2397, N2386);
nor NOR2 (N2398, N2378, N1953);
or OR4 (N2399, N2380, N227, N1034, N1761);
and AND4 (N2400, N2394, N24, N521, N1926);
nand NAND4 (N2401, N2388, N56, N458, N1703);
buf BUF1 (N2402, N2383);
not NOT1 (N2403, N2382);
nor NOR2 (N2404, N2400, N38);
nand NAND2 (N2405, N2398, N1894);
nand NAND4 (N2406, N2402, N487, N965, N1121);
nor NOR4 (N2407, N2397, N1059, N1031, N1363);
or OR3 (N2408, N2405, N2122, N411);
or OR2 (N2409, N2407, N1806);
xor XOR2 (N2410, N2409, N316);
or OR3 (N2411, N2408, N1443, N485);
nor NOR4 (N2412, N2406, N1322, N870, N2047);
xor XOR2 (N2413, N2410, N2000);
or OR2 (N2414, N2411, N484);
xor XOR2 (N2415, N2399, N805);
nand NAND4 (N2416, N2395, N687, N1940, N2315);
not NOT1 (N2417, N2414);
and AND4 (N2418, N2415, N1315, N2264, N1891);
or OR2 (N2419, N2396, N2150);
and AND4 (N2420, N2416, N404, N1564, N279);
xor XOR2 (N2421, N2417, N631);
or OR3 (N2422, N2390, N423, N2292);
or OR4 (N2423, N2422, N1761, N946, N158);
nor NOR3 (N2424, N2420, N2308, N550);
and AND2 (N2425, N2401, N1290);
nand NAND3 (N2426, N2413, N1676, N18);
xor XOR2 (N2427, N2426, N610);
or OR4 (N2428, N2423, N2124, N1626, N1141);
and AND3 (N2429, N2403, N1457, N355);
nand NAND4 (N2430, N2424, N2372, N1813, N1387);
xor XOR2 (N2431, N2428, N92);
and AND3 (N2432, N2430, N1542, N574);
not NOT1 (N2433, N2425);
xor XOR2 (N2434, N2421, N1151);
and AND3 (N2435, N2429, N1558, N707);
and AND4 (N2436, N2434, N280, N2165, N1972);
nor NOR3 (N2437, N2435, N1489, N1829);
buf BUF1 (N2438, N2436);
xor XOR2 (N2439, N2431, N1051);
not NOT1 (N2440, N2427);
xor XOR2 (N2441, N2412, N325);
not NOT1 (N2442, N2437);
or OR2 (N2443, N2419, N438);
nor NOR4 (N2444, N2432, N81, N1078, N515);
buf BUF1 (N2445, N2441);
buf BUF1 (N2446, N2439);
and AND2 (N2447, N2418, N1717);
and AND2 (N2448, N2442, N232);
and AND3 (N2449, N2440, N952, N2121);
xor XOR2 (N2450, N2433, N1276);
and AND2 (N2451, N2446, N1693);
buf BUF1 (N2452, N2443);
or OR4 (N2453, N2447, N282, N922, N2444);
nand NAND2 (N2454, N1788, N365);
and AND3 (N2455, N2404, N457, N271);
or OR2 (N2456, N2453, N1679);
buf BUF1 (N2457, N2448);
nand NAND2 (N2458, N2457, N79);
xor XOR2 (N2459, N2454, N1387);
not NOT1 (N2460, N2445);
not NOT1 (N2461, N2455);
or OR3 (N2462, N2451, N691, N475);
not NOT1 (N2463, N2459);
nor NOR3 (N2464, N2449, N1308, N1598);
buf BUF1 (N2465, N2456);
buf BUF1 (N2466, N2465);
and AND2 (N2467, N2450, N1524);
not NOT1 (N2468, N2460);
or OR2 (N2469, N2461, N282);
or OR4 (N2470, N2464, N218, N1582, N487);
nor NOR4 (N2471, N2469, N229, N1103, N503);
nor NOR3 (N2472, N2471, N2165, N1384);
buf BUF1 (N2473, N2467);
nand NAND2 (N2474, N2466, N702);
not NOT1 (N2475, N2473);
nand NAND3 (N2476, N2463, N1557, N1565);
and AND3 (N2477, N2470, N879, N993);
buf BUF1 (N2478, N2438);
and AND2 (N2479, N2477, N1529);
and AND3 (N2480, N2476, N1551, N2421);
nor NOR2 (N2481, N2462, N761);
and AND3 (N2482, N2480, N1918, N1500);
nor NOR2 (N2483, N2468, N1248);
not NOT1 (N2484, N2452);
nand NAND2 (N2485, N2472, N735);
xor XOR2 (N2486, N2482, N2443);
not NOT1 (N2487, N2458);
nor NOR3 (N2488, N2475, N1329, N1104);
and AND4 (N2489, N2486, N1340, N1662, N2314);
xor XOR2 (N2490, N2478, N19);
not NOT1 (N2491, N2487);
xor XOR2 (N2492, N2481, N1258);
not NOT1 (N2493, N2479);
xor XOR2 (N2494, N2492, N405);
xor XOR2 (N2495, N2484, N1025);
and AND4 (N2496, N2494, N1187, N1166, N2224);
xor XOR2 (N2497, N2485, N628);
nor NOR2 (N2498, N2493, N391);
nand NAND3 (N2499, N2474, N1060, N1613);
nand NAND4 (N2500, N2490, N2035, N2352, N1158);
nand NAND2 (N2501, N2497, N1155);
nor NOR2 (N2502, N2496, N562);
xor XOR2 (N2503, N2498, N1006);
not NOT1 (N2504, N2502);
not NOT1 (N2505, N2483);
xor XOR2 (N2506, N2489, N2298);
nand NAND4 (N2507, N2504, N1170, N1427, N595);
and AND2 (N2508, N2491, N1346);
or OR4 (N2509, N2488, N1923, N1892, N314);
not NOT1 (N2510, N2495);
xor XOR2 (N2511, N2505, N2289);
and AND3 (N2512, N2506, N472, N2085);
or OR4 (N2513, N2501, N2135, N42, N2060);
xor XOR2 (N2514, N2512, N1093);
xor XOR2 (N2515, N2514, N628);
xor XOR2 (N2516, N2499, N1613);
nand NAND2 (N2517, N2515, N167);
and AND3 (N2518, N2508, N38, N144);
not NOT1 (N2519, N2517);
not NOT1 (N2520, N2510);
buf BUF1 (N2521, N2511);
and AND3 (N2522, N2521, N2465, N2391);
not NOT1 (N2523, N2503);
nor NOR3 (N2524, N2518, N185, N2138);
buf BUF1 (N2525, N2524);
buf BUF1 (N2526, N2500);
not NOT1 (N2527, N2509);
and AND4 (N2528, N2525, N2450, N2412, N2516);
nor NOR4 (N2529, N1055, N810, N1826, N2067);
not NOT1 (N2530, N2523);
nor NOR2 (N2531, N2513, N2242);
not NOT1 (N2532, N2529);
nor NOR2 (N2533, N2530, N1296);
buf BUF1 (N2534, N2519);
nand NAND3 (N2535, N2528, N870, N231);
not NOT1 (N2536, N2532);
and AND4 (N2537, N2507, N1500, N967, N1427);
nor NOR2 (N2538, N2533, N489);
xor XOR2 (N2539, N2531, N664);
not NOT1 (N2540, N2539);
or OR4 (N2541, N2526, N1829, N1205, N975);
and AND2 (N2542, N2538, N2506);
buf BUF1 (N2543, N2537);
and AND3 (N2544, N2543, N2097, N159);
nor NOR4 (N2545, N2535, N134, N1043, N592);
or OR4 (N2546, N2545, N65, N1434, N1850);
xor XOR2 (N2547, N2544, N1694);
buf BUF1 (N2548, N2520);
buf BUF1 (N2549, N2546);
nand NAND2 (N2550, N2522, N1507);
and AND3 (N2551, N2548, N408, N1423);
not NOT1 (N2552, N2547);
or OR3 (N2553, N2550, N1845, N1660);
or OR3 (N2554, N2540, N1750, N1415);
xor XOR2 (N2555, N2551, N1838);
not NOT1 (N2556, N2555);
or OR3 (N2557, N2534, N2419, N2448);
nand NAND2 (N2558, N2552, N1756);
not NOT1 (N2559, N2536);
or OR2 (N2560, N2542, N1596);
xor XOR2 (N2561, N2560, N1900);
or OR3 (N2562, N2559, N1043, N33);
nand NAND4 (N2563, N2554, N1594, N452, N1455);
buf BUF1 (N2564, N2556);
xor XOR2 (N2565, N2558, N230);
xor XOR2 (N2566, N2527, N521);
nor NOR3 (N2567, N2565, N2142, N714);
or OR4 (N2568, N2553, N1495, N2502, N139);
nor NOR2 (N2569, N2557, N2243);
and AND2 (N2570, N2566, N1228);
not NOT1 (N2571, N2561);
xor XOR2 (N2572, N2568, N135);
and AND2 (N2573, N2541, N1);
or OR3 (N2574, N2563, N45, N1417);
not NOT1 (N2575, N2569);
xor XOR2 (N2576, N2549, N1308);
buf BUF1 (N2577, N2576);
xor XOR2 (N2578, N2570, N2319);
and AND2 (N2579, N2578, N326);
buf BUF1 (N2580, N2577);
or OR2 (N2581, N2580, N1661);
not NOT1 (N2582, N2579);
and AND4 (N2583, N2567, N2184, N147, N1106);
buf BUF1 (N2584, N2575);
or OR4 (N2585, N2581, N2355, N526, N294);
or OR3 (N2586, N2584, N567, N1943);
xor XOR2 (N2587, N2571, N1689);
xor XOR2 (N2588, N2572, N1662);
xor XOR2 (N2589, N2564, N1186);
not NOT1 (N2590, N2574);
xor XOR2 (N2591, N2573, N667);
buf BUF1 (N2592, N2562);
or OR2 (N2593, N2585, N644);
not NOT1 (N2594, N2592);
buf BUF1 (N2595, N2594);
and AND2 (N2596, N2586, N802);
nor NOR2 (N2597, N2595, N43);
nand NAND3 (N2598, N2582, N1838, N2371);
nand NAND3 (N2599, N2588, N1261, N699);
nand NAND4 (N2600, N2599, N846, N1654, N755);
not NOT1 (N2601, N2597);
nor NOR2 (N2602, N2601, N2418);
nand NAND2 (N2603, N2598, N1236);
nor NOR4 (N2604, N2591, N11, N33, N2547);
buf BUF1 (N2605, N2593);
xor XOR2 (N2606, N2602, N2335);
nor NOR3 (N2607, N2590, N1223, N382);
xor XOR2 (N2608, N2607, N2429);
buf BUF1 (N2609, N2608);
not NOT1 (N2610, N2596);
nand NAND3 (N2611, N2600, N2352, N1254);
not NOT1 (N2612, N2609);
not NOT1 (N2613, N2589);
and AND2 (N2614, N2587, N70);
and AND3 (N2615, N2611, N1801, N1427);
nor NOR4 (N2616, N2612, N2425, N41, N1578);
not NOT1 (N2617, N2616);
not NOT1 (N2618, N2614);
xor XOR2 (N2619, N2613, N94);
or OR2 (N2620, N2617, N811);
buf BUF1 (N2621, N2605);
or OR2 (N2622, N2621, N1242);
nor NOR4 (N2623, N2606, N460, N1736, N1726);
buf BUF1 (N2624, N2604);
and AND4 (N2625, N2622, N2288, N582, N576);
xor XOR2 (N2626, N2603, N1655);
not NOT1 (N2627, N2610);
buf BUF1 (N2628, N2583);
and AND2 (N2629, N2628, N372);
xor XOR2 (N2630, N2618, N1100);
not NOT1 (N2631, N2627);
nor NOR4 (N2632, N2623, N546, N627, N1923);
xor XOR2 (N2633, N2629, N2472);
nor NOR2 (N2634, N2633, N2552);
not NOT1 (N2635, N2626);
nor NOR2 (N2636, N2615, N2598);
xor XOR2 (N2637, N2631, N1857);
nor NOR4 (N2638, N2637, N1480, N655, N1163);
xor XOR2 (N2639, N2630, N2096);
xor XOR2 (N2640, N2635, N552);
or OR2 (N2641, N2639, N645);
nand NAND2 (N2642, N2640, N1409);
xor XOR2 (N2643, N2634, N664);
xor XOR2 (N2644, N2620, N1706);
xor XOR2 (N2645, N2638, N105);
and AND4 (N2646, N2625, N333, N1126, N894);
nand NAND4 (N2647, N2619, N5, N1133, N604);
or OR2 (N2648, N2642, N673);
and AND4 (N2649, N2644, N2445, N1912, N460);
buf BUF1 (N2650, N2647);
not NOT1 (N2651, N2636);
buf BUF1 (N2652, N2649);
nand NAND4 (N2653, N2645, N2100, N2241, N1943);
buf BUF1 (N2654, N2632);
xor XOR2 (N2655, N2654, N920);
nand NAND2 (N2656, N2624, N2069);
buf BUF1 (N2657, N2641);
nor NOR2 (N2658, N2657, N1008);
nor NOR4 (N2659, N2655, N1899, N1784, N143);
nor NOR4 (N2660, N2651, N1495, N548, N1477);
and AND2 (N2661, N2646, N1686);
nor NOR2 (N2662, N2661, N251);
nor NOR4 (N2663, N2659, N650, N1170, N2299);
nand NAND2 (N2664, N2648, N1968);
and AND4 (N2665, N2652, N746, N835, N1077);
nor NOR3 (N2666, N2643, N693, N1918);
or OR4 (N2667, N2663, N1911, N1513, N2628);
nor NOR2 (N2668, N2650, N1349);
xor XOR2 (N2669, N2656, N1183);
or OR4 (N2670, N2666, N80, N2056, N2581);
nor NOR3 (N2671, N2665, N647, N477);
and AND2 (N2672, N2662, N390);
buf BUF1 (N2673, N2671);
xor XOR2 (N2674, N2658, N1559);
nor NOR3 (N2675, N2664, N1581, N116);
nand NAND2 (N2676, N2674, N2585);
not NOT1 (N2677, N2673);
not NOT1 (N2678, N2672);
nand NAND4 (N2679, N2677, N2570, N1931, N805);
buf BUF1 (N2680, N2669);
nor NOR2 (N2681, N2678, N30);
nand NAND4 (N2682, N2670, N1275, N2256, N907);
not NOT1 (N2683, N2680);
and AND4 (N2684, N2667, N1240, N1846, N1715);
or OR4 (N2685, N2675, N2518, N1847, N1901);
xor XOR2 (N2686, N2682, N2513);
xor XOR2 (N2687, N2685, N1598);
not NOT1 (N2688, N2683);
xor XOR2 (N2689, N2668, N1027);
and AND2 (N2690, N2688, N454);
buf BUF1 (N2691, N2681);
xor XOR2 (N2692, N2653, N1722);
and AND4 (N2693, N2692, N1568, N1900, N136);
buf BUF1 (N2694, N2691);
or OR4 (N2695, N2689, N2296, N39, N299);
not NOT1 (N2696, N2690);
or OR2 (N2697, N2679, N105);
not NOT1 (N2698, N2660);
not NOT1 (N2699, N2693);
nor NOR3 (N2700, N2694, N2682, N1755);
buf BUF1 (N2701, N2696);
not NOT1 (N2702, N2676);
not NOT1 (N2703, N2695);
nand NAND4 (N2704, N2698, N2400, N2524, N1446);
or OR2 (N2705, N2704, N342);
xor XOR2 (N2706, N2686, N570);
nand NAND3 (N2707, N2700, N2661, N212);
xor XOR2 (N2708, N2684, N1494);
and AND4 (N2709, N2703, N1807, N2463, N2055);
nor NOR3 (N2710, N2699, N237, N600);
and AND4 (N2711, N2707, N2416, N526, N1108);
nor NOR4 (N2712, N2708, N2376, N1779, N1447);
not NOT1 (N2713, N2711);
or OR3 (N2714, N2709, N733, N1939);
xor XOR2 (N2715, N2714, N1047);
nand NAND2 (N2716, N2701, N1640);
nand NAND3 (N2717, N2716, N2508, N581);
nor NOR2 (N2718, N2705, N1250);
nor NOR4 (N2719, N2706, N1221, N1330, N1876);
buf BUF1 (N2720, N2717);
nand NAND3 (N2721, N2715, N1024, N45);
buf BUF1 (N2722, N2702);
xor XOR2 (N2723, N2697, N1086);
or OR2 (N2724, N2710, N1263);
xor XOR2 (N2725, N2723, N178);
not NOT1 (N2726, N2724);
buf BUF1 (N2727, N2687);
buf BUF1 (N2728, N2721);
and AND2 (N2729, N2725, N1439);
and AND4 (N2730, N2729, N357, N312, N937);
buf BUF1 (N2731, N2728);
and AND3 (N2732, N2726, N2571, N2173);
or OR4 (N2733, N2731, N2048, N1883, N867);
nand NAND2 (N2734, N2720, N356);
xor XOR2 (N2735, N2733, N2229);
and AND2 (N2736, N2732, N1447);
nand NAND2 (N2737, N2713, N2150);
nand NAND3 (N2738, N2730, N157, N1731);
buf BUF1 (N2739, N2738);
nand NAND3 (N2740, N2727, N2358, N2536);
or OR2 (N2741, N2719, N1341);
buf BUF1 (N2742, N2734);
buf BUF1 (N2743, N2742);
nor NOR4 (N2744, N2741, N193, N2420, N130);
xor XOR2 (N2745, N2744, N1796);
or OR3 (N2746, N2745, N2323, N695);
and AND3 (N2747, N2712, N1312, N1216);
xor XOR2 (N2748, N2722, N218);
not NOT1 (N2749, N2740);
or OR3 (N2750, N2739, N34, N2144);
not NOT1 (N2751, N2736);
not NOT1 (N2752, N2748);
or OR2 (N2753, N2718, N1994);
nand NAND3 (N2754, N2752, N1351, N1395);
nor NOR3 (N2755, N2749, N1151, N631);
and AND2 (N2756, N2751, N471);
nor NOR3 (N2757, N2750, N1001, N1206);
nor NOR2 (N2758, N2747, N1459);
not NOT1 (N2759, N2753);
or OR4 (N2760, N2757, N1827, N1249, N2624);
nand NAND3 (N2761, N2743, N150, N155);
buf BUF1 (N2762, N2755);
buf BUF1 (N2763, N2735);
and AND4 (N2764, N2758, N366, N2194, N188);
buf BUF1 (N2765, N2759);
xor XOR2 (N2766, N2764, N1234);
buf BUF1 (N2767, N2760);
not NOT1 (N2768, N2761);
and AND3 (N2769, N2763, N1054, N631);
nor NOR3 (N2770, N2756, N1034, N116);
nor NOR2 (N2771, N2754, N1783);
nand NAND4 (N2772, N2770, N2194, N52, N1540);
buf BUF1 (N2773, N2771);
nor NOR2 (N2774, N2768, N1674);
buf BUF1 (N2775, N2774);
xor XOR2 (N2776, N2767, N1780);
nor NOR3 (N2777, N2762, N1664, N1476);
nand NAND4 (N2778, N2772, N499, N2241, N2714);
buf BUF1 (N2779, N2776);
nor NOR3 (N2780, N2778, N591, N1597);
buf BUF1 (N2781, N2775);
buf BUF1 (N2782, N2769);
and AND2 (N2783, N2766, N2120);
or OR3 (N2784, N2781, N305, N2035);
xor XOR2 (N2785, N2784, N354);
and AND4 (N2786, N2773, N2662, N992, N896);
nor NOR3 (N2787, N2779, N1296, N2105);
nand NAND4 (N2788, N2765, N1828, N759, N682);
and AND4 (N2789, N2787, N1656, N2640, N2249);
or OR4 (N2790, N2786, N2597, N1371, N1620);
nor NOR3 (N2791, N2746, N2150, N986);
nand NAND3 (N2792, N2790, N2220, N1627);
xor XOR2 (N2793, N2785, N662);
nor NOR4 (N2794, N2788, N1946, N2559, N2556);
and AND3 (N2795, N2794, N372, N1929);
buf BUF1 (N2796, N2783);
buf BUF1 (N2797, N2782);
or OR3 (N2798, N2789, N1477, N1196);
and AND3 (N2799, N2798, N596, N2598);
or OR2 (N2800, N2777, N2699);
buf BUF1 (N2801, N2780);
nor NOR3 (N2802, N2796, N2392, N1097);
nand NAND3 (N2803, N2800, N2111, N2787);
buf BUF1 (N2804, N2793);
and AND2 (N2805, N2803, N2746);
or OR3 (N2806, N2737, N2678, N1026);
nand NAND4 (N2807, N2805, N1411, N804, N1625);
and AND2 (N2808, N2797, N583);
not NOT1 (N2809, N2799);
nand NAND2 (N2810, N2804, N544);
nor NOR3 (N2811, N2807, N1617, N1959);
not NOT1 (N2812, N2795);
nor NOR4 (N2813, N2791, N566, N1549, N2165);
not NOT1 (N2814, N2808);
and AND4 (N2815, N2802, N1729, N2037, N1504);
nor NOR4 (N2816, N2792, N1010, N1050, N235);
nor NOR3 (N2817, N2814, N1550, N1257);
xor XOR2 (N2818, N2817, N872);
xor XOR2 (N2819, N2801, N1156);
nor NOR3 (N2820, N2813, N2266, N2669);
not NOT1 (N2821, N2820);
xor XOR2 (N2822, N2815, N2783);
or OR3 (N2823, N2811, N2313, N2134);
nand NAND4 (N2824, N2810, N1524, N2037, N1198);
and AND3 (N2825, N2819, N261, N494);
nand NAND2 (N2826, N2816, N2674);
nand NAND2 (N2827, N2809, N1005);
buf BUF1 (N2828, N2822);
not NOT1 (N2829, N2827);
buf BUF1 (N2830, N2806);
nor NOR4 (N2831, N2829, N1677, N2578, N1931);
or OR3 (N2832, N2824, N2133, N666);
xor XOR2 (N2833, N2812, N271);
and AND2 (N2834, N2833, N710);
xor XOR2 (N2835, N2831, N1143);
not NOT1 (N2836, N2826);
nand NAND2 (N2837, N2835, N532);
xor XOR2 (N2838, N2821, N363);
buf BUF1 (N2839, N2823);
xor XOR2 (N2840, N2828, N2553);
not NOT1 (N2841, N2818);
not NOT1 (N2842, N2830);
nor NOR4 (N2843, N2841, N2386, N405, N2781);
and AND3 (N2844, N2837, N2652, N1575);
nor NOR2 (N2845, N2838, N2827);
not NOT1 (N2846, N2825);
buf BUF1 (N2847, N2844);
not NOT1 (N2848, N2839);
and AND3 (N2849, N2843, N1369, N331);
nor NOR2 (N2850, N2845, N2755);
nor NOR4 (N2851, N2834, N1151, N2706, N376);
or OR2 (N2852, N2849, N1614);
xor XOR2 (N2853, N2848, N978);
not NOT1 (N2854, N2846);
buf BUF1 (N2855, N2854);
or OR3 (N2856, N2847, N446, N2207);
nand NAND4 (N2857, N2840, N197, N1210, N1123);
xor XOR2 (N2858, N2857, N1832);
not NOT1 (N2859, N2832);
not NOT1 (N2860, N2850);
or OR4 (N2861, N2852, N1348, N1488, N1278);
nand NAND2 (N2862, N2836, N2560);
not NOT1 (N2863, N2851);
nor NOR4 (N2864, N2858, N2482, N1584, N1685);
nor NOR3 (N2865, N2863, N1959, N2800);
nor NOR3 (N2866, N2855, N1409, N1176);
xor XOR2 (N2867, N2856, N231);
nand NAND2 (N2868, N2859, N2565);
nor NOR3 (N2869, N2853, N907, N1469);
not NOT1 (N2870, N2862);
xor XOR2 (N2871, N2842, N596);
nand NAND3 (N2872, N2868, N2408, N373);
buf BUF1 (N2873, N2869);
not NOT1 (N2874, N2866);
buf BUF1 (N2875, N2870);
not NOT1 (N2876, N2867);
xor XOR2 (N2877, N2865, N2000);
xor XOR2 (N2878, N2871, N1230);
nor NOR2 (N2879, N2872, N32);
xor XOR2 (N2880, N2873, N380);
nand NAND4 (N2881, N2861, N2707, N2757, N1689);
buf BUF1 (N2882, N2878);
xor XOR2 (N2883, N2864, N2748);
or OR3 (N2884, N2882, N266, N2144);
buf BUF1 (N2885, N2860);
not NOT1 (N2886, N2885);
nand NAND2 (N2887, N2879, N2286);
or OR4 (N2888, N2880, N2696, N2473, N1140);
buf BUF1 (N2889, N2876);
xor XOR2 (N2890, N2877, N735);
xor XOR2 (N2891, N2875, N456);
or OR3 (N2892, N2881, N2863, N2822);
and AND4 (N2893, N2890, N1345, N1882, N2466);
or OR2 (N2894, N2891, N1775);
not NOT1 (N2895, N2888);
and AND2 (N2896, N2894, N2638);
xor XOR2 (N2897, N2887, N1734);
nand NAND2 (N2898, N2895, N2116);
nand NAND3 (N2899, N2884, N2800, N2518);
xor XOR2 (N2900, N2897, N1657);
not NOT1 (N2901, N2874);
nor NOR2 (N2902, N2898, N1050);
nand NAND4 (N2903, N2899, N2341, N2166, N1897);
and AND3 (N2904, N2903, N283, N1768);
buf BUF1 (N2905, N2904);
or OR3 (N2906, N2901, N2372, N1055);
xor XOR2 (N2907, N2896, N1721);
nor NOR2 (N2908, N2905, N1879);
or OR4 (N2909, N2892, N320, N847, N1996);
or OR2 (N2910, N2893, N340);
buf BUF1 (N2911, N2910);
nand NAND2 (N2912, N2886, N39);
or OR2 (N2913, N2902, N98);
and AND3 (N2914, N2908, N2303, N773);
xor XOR2 (N2915, N2883, N2282);
xor XOR2 (N2916, N2907, N2601);
nor NOR2 (N2917, N2909, N1756);
buf BUF1 (N2918, N2889);
nor NOR4 (N2919, N2900, N111, N2327, N1520);
xor XOR2 (N2920, N2918, N140);
and AND3 (N2921, N2916, N317, N2706);
or OR4 (N2922, N2915, N755, N1729, N1064);
xor XOR2 (N2923, N2922, N2385);
xor XOR2 (N2924, N2906, N1848);
or OR4 (N2925, N2914, N1598, N2453, N385);
xor XOR2 (N2926, N2917, N2682);
buf BUF1 (N2927, N2911);
or OR2 (N2928, N2924, N894);
nand NAND3 (N2929, N2927, N1039, N2864);
not NOT1 (N2930, N2928);
and AND4 (N2931, N2921, N1281, N2860, N2840);
nor NOR3 (N2932, N2923, N263, N2295);
buf BUF1 (N2933, N2931);
nor NOR4 (N2934, N2933, N65, N1765, N2573);
and AND4 (N2935, N2912, N2001, N1729, N1832);
and AND2 (N2936, N2920, N2181);
or OR2 (N2937, N2935, N977);
and AND4 (N2938, N2913, N528, N2713, N1187);
and AND4 (N2939, N2929, N21, N394, N457);
nor NOR4 (N2940, N2936, N1502, N1298, N1375);
nand NAND3 (N2941, N2925, N630, N1669);
not NOT1 (N2942, N2937);
nand NAND3 (N2943, N2930, N384, N1391);
xor XOR2 (N2944, N2943, N2151);
or OR3 (N2945, N2941, N905, N346);
nand NAND2 (N2946, N2934, N1549);
not NOT1 (N2947, N2932);
and AND3 (N2948, N2926, N2429, N1449);
xor XOR2 (N2949, N2940, N2757);
and AND4 (N2950, N2942, N1207, N2099, N2759);
nand NAND2 (N2951, N2949, N779);
and AND3 (N2952, N2938, N2116, N2031);
nor NOR3 (N2953, N2919, N2909, N207);
buf BUF1 (N2954, N2950);
nor NOR2 (N2955, N2954, N2031);
and AND4 (N2956, N2948, N923, N818, N444);
nand NAND4 (N2957, N2951, N1474, N1079, N2847);
buf BUF1 (N2958, N2946);
not NOT1 (N2959, N2958);
xor XOR2 (N2960, N2947, N431);
and AND3 (N2961, N2956, N2685, N1549);
xor XOR2 (N2962, N2955, N2546);
buf BUF1 (N2963, N2959);
buf BUF1 (N2964, N2952);
nor NOR3 (N2965, N2957, N306, N2413);
and AND4 (N2966, N2960, N760, N62, N864);
xor XOR2 (N2967, N2962, N2669);
and AND4 (N2968, N2967, N777, N438, N377);
and AND4 (N2969, N2939, N1387, N50, N35);
not NOT1 (N2970, N2968);
xor XOR2 (N2971, N2964, N1834);
nor NOR4 (N2972, N2961, N1893, N464, N2762);
and AND4 (N2973, N2971, N101, N2839, N101);
or OR3 (N2974, N2972, N54, N1085);
xor XOR2 (N2975, N2974, N147);
not NOT1 (N2976, N2969);
buf BUF1 (N2977, N2945);
and AND3 (N2978, N2977, N1998, N2680);
not NOT1 (N2979, N2953);
buf BUF1 (N2980, N2978);
or OR3 (N2981, N2963, N1774, N929);
buf BUF1 (N2982, N2979);
buf BUF1 (N2983, N2981);
nor NOR3 (N2984, N2975, N1544, N2356);
buf BUF1 (N2985, N2983);
not NOT1 (N2986, N2965);
not NOT1 (N2987, N2980);
not NOT1 (N2988, N2976);
nor NOR3 (N2989, N2987, N2141, N2502);
and AND2 (N2990, N2986, N502);
and AND3 (N2991, N2970, N2329, N1407);
buf BUF1 (N2992, N2984);
and AND3 (N2993, N2990, N138, N2407);
nor NOR2 (N2994, N2982, N681);
or OR2 (N2995, N2989, N46);
nand NAND3 (N2996, N2991, N902, N954);
buf BUF1 (N2997, N2995);
xor XOR2 (N2998, N2985, N2612);
buf BUF1 (N2999, N2994);
not NOT1 (N3000, N2944);
or OR3 (N3001, N2973, N2885, N2177);
not NOT1 (N3002, N2992);
or OR2 (N3003, N2988, N1572);
xor XOR2 (N3004, N2997, N550);
nand NAND2 (N3005, N3001, N360);
buf BUF1 (N3006, N2966);
xor XOR2 (N3007, N3005, N560);
nand NAND4 (N3008, N3006, N685, N165, N1620);
nand NAND2 (N3009, N3002, N1811);
buf BUF1 (N3010, N3000);
and AND3 (N3011, N3004, N1150, N2198);
or OR2 (N3012, N3011, N2417);
or OR2 (N3013, N2998, N2814);
buf BUF1 (N3014, N3012);
and AND3 (N3015, N3013, N2728, N1341);
not NOT1 (N3016, N2999);
nor NOR3 (N3017, N3014, N2626, N241);
not NOT1 (N3018, N3003);
xor XOR2 (N3019, N3017, N2710);
xor XOR2 (N3020, N2996, N1806);
xor XOR2 (N3021, N3010, N146);
or OR3 (N3022, N3019, N2067, N2431);
and AND3 (N3023, N3018, N2077, N1884);
and AND4 (N3024, N3021, N1785, N507, N1003);
and AND2 (N3025, N3015, N2319);
or OR3 (N3026, N3025, N308, N576);
or OR3 (N3027, N3009, N362, N2919);
and AND4 (N3028, N3016, N240, N2856, N2955);
nand NAND4 (N3029, N3024, N2086, N2236, N2261);
not NOT1 (N3030, N3008);
and AND2 (N3031, N3030, N1119);
xor XOR2 (N3032, N3031, N2238);
nor NOR2 (N3033, N3028, N1200);
and AND3 (N3034, N3032, N1026, N154);
not NOT1 (N3035, N3023);
nor NOR4 (N3036, N3026, N1839, N559, N268);
not NOT1 (N3037, N3033);
xor XOR2 (N3038, N3022, N899);
nor NOR2 (N3039, N3036, N1753);
nand NAND3 (N3040, N3007, N2969, N780);
or OR3 (N3041, N3040, N1753, N2758);
buf BUF1 (N3042, N3038);
nor NOR4 (N3043, N3041, N646, N1301, N1835);
not NOT1 (N3044, N3027);
not NOT1 (N3045, N3037);
or OR2 (N3046, N3039, N2629);
buf BUF1 (N3047, N3035);
and AND4 (N3048, N2993, N508, N917, N1585);
or OR4 (N3049, N3044, N2622, N1260, N999);
or OR4 (N3050, N3047, N1272, N1857, N2207);
or OR2 (N3051, N3034, N2709);
and AND4 (N3052, N3048, N2468, N338, N2257);
xor XOR2 (N3053, N3049, N346);
xor XOR2 (N3054, N3051, N135);
and AND2 (N3055, N3050, N879);
nor NOR2 (N3056, N3053, N429);
nor NOR2 (N3057, N3043, N2161);
xor XOR2 (N3058, N3029, N873);
xor XOR2 (N3059, N3054, N1508);
or OR3 (N3060, N3056, N792, N706);
buf BUF1 (N3061, N3020);
and AND4 (N3062, N3046, N1423, N2178, N872);
xor XOR2 (N3063, N3057, N1691);
nand NAND3 (N3064, N3052, N1524, N135);
xor XOR2 (N3065, N3042, N2817);
xor XOR2 (N3066, N3058, N1253);
nor NOR4 (N3067, N3055, N1133, N982, N1595);
or OR2 (N3068, N3059, N2828);
or OR4 (N3069, N3067, N1908, N2156, N1974);
nor NOR2 (N3070, N3066, N2020);
and AND2 (N3071, N3060, N2802);
not NOT1 (N3072, N3064);
buf BUF1 (N3073, N3063);
nor NOR2 (N3074, N3073, N809);
nand NAND4 (N3075, N3062, N569, N852, N821);
and AND4 (N3076, N3045, N2513, N2702, N1118);
not NOT1 (N3077, N3068);
and AND4 (N3078, N3061, N659, N607, N826);
nor NOR4 (N3079, N3070, N48, N1026, N2205);
nor NOR3 (N3080, N3072, N952, N956);
nand NAND3 (N3081, N3069, N2492, N2424);
nor NOR4 (N3082, N3071, N1363, N2841, N11);
and AND4 (N3083, N3082, N1825, N1990, N2378);
not NOT1 (N3084, N3083);
xor XOR2 (N3085, N3080, N1867);
xor XOR2 (N3086, N3076, N2089);
not NOT1 (N3087, N3074);
or OR4 (N3088, N3081, N213, N2486, N609);
and AND3 (N3089, N3075, N1227, N1677);
nand NAND2 (N3090, N3085, N430);
not NOT1 (N3091, N3084);
buf BUF1 (N3092, N3089);
nand NAND3 (N3093, N3086, N306, N2908);
not NOT1 (N3094, N3078);
xor XOR2 (N3095, N3079, N620);
and AND3 (N3096, N3091, N967, N844);
buf BUF1 (N3097, N3087);
xor XOR2 (N3098, N3092, N1144);
nand NAND3 (N3099, N3090, N646, N892);
and AND4 (N3100, N3097, N2094, N2494, N729);
buf BUF1 (N3101, N3095);
xor XOR2 (N3102, N3096, N1325);
buf BUF1 (N3103, N3099);
nor NOR4 (N3104, N3077, N265, N879, N527);
nor NOR2 (N3105, N3101, N2234);
or OR3 (N3106, N3100, N2180, N73);
xor XOR2 (N3107, N3103, N1477);
not NOT1 (N3108, N3093);
and AND3 (N3109, N3088, N915, N1310);
xor XOR2 (N3110, N3107, N260);
nor NOR3 (N3111, N3065, N980, N465);
and AND2 (N3112, N3106, N1237);
or OR4 (N3113, N3094, N1855, N40, N1838);
not NOT1 (N3114, N3104);
or OR4 (N3115, N3102, N1505, N929, N2301);
not NOT1 (N3116, N3110);
or OR3 (N3117, N3112, N1529, N124);
nor NOR2 (N3118, N3117, N1651);
not NOT1 (N3119, N3105);
xor XOR2 (N3120, N3114, N836);
not NOT1 (N3121, N3108);
not NOT1 (N3122, N3121);
buf BUF1 (N3123, N3120);
buf BUF1 (N3124, N3109);
or OR2 (N3125, N3122, N2994);
not NOT1 (N3126, N3123);
or OR2 (N3127, N3111, N2947);
nor NOR3 (N3128, N3118, N1523, N2040);
or OR4 (N3129, N3116, N2599, N1465, N2590);
nor NOR2 (N3130, N3126, N2371);
xor XOR2 (N3131, N3113, N2740);
nor NOR3 (N3132, N3115, N78, N1156);
not NOT1 (N3133, N3132);
buf BUF1 (N3134, N3127);
buf BUF1 (N3135, N3130);
not NOT1 (N3136, N3119);
or OR3 (N3137, N3128, N1733, N1293);
xor XOR2 (N3138, N3135, N2888);
nor NOR4 (N3139, N3137, N88, N718, N2184);
nor NOR3 (N3140, N3136, N1656, N684);
nor NOR4 (N3141, N3140, N649, N1275, N1642);
nand NAND3 (N3142, N3131, N234, N187);
xor XOR2 (N3143, N3133, N2858);
or OR3 (N3144, N3124, N3037, N2705);
buf BUF1 (N3145, N3098);
nor NOR3 (N3146, N3141, N732, N2504);
not NOT1 (N3147, N3146);
nand NAND2 (N3148, N3145, N988);
nor NOR4 (N3149, N3134, N2508, N906, N10);
nor NOR4 (N3150, N3138, N1902, N1119, N1129);
nand NAND4 (N3151, N3150, N1694, N68, N1606);
and AND3 (N3152, N3148, N835, N1940);
not NOT1 (N3153, N3125);
and AND2 (N3154, N3152, N920);
not NOT1 (N3155, N3139);
not NOT1 (N3156, N3144);
nor NOR3 (N3157, N3149, N1721, N229);
buf BUF1 (N3158, N3155);
not NOT1 (N3159, N3154);
nand NAND2 (N3160, N3158, N695);
buf BUF1 (N3161, N3160);
or OR3 (N3162, N3142, N2580, N400);
buf BUF1 (N3163, N3156);
and AND3 (N3164, N3161, N2816, N438);
nor NOR3 (N3165, N3143, N2891, N2015);
not NOT1 (N3166, N3151);
buf BUF1 (N3167, N3129);
or OR3 (N3168, N3153, N2643, N302);
and AND3 (N3169, N3165, N2218, N742);
buf BUF1 (N3170, N3163);
nor NOR2 (N3171, N3168, N2151);
buf BUF1 (N3172, N3162);
xor XOR2 (N3173, N3172, N3027);
xor XOR2 (N3174, N3147, N452);
buf BUF1 (N3175, N3174);
xor XOR2 (N3176, N3167, N436);
or OR2 (N3177, N3164, N1051);
nand NAND2 (N3178, N3166, N1389);
or OR2 (N3179, N3173, N1011);
or OR3 (N3180, N3175, N2346, N1212);
not NOT1 (N3181, N3171);
xor XOR2 (N3182, N3170, N3087);
and AND4 (N3183, N3182, N2732, N36, N1444);
buf BUF1 (N3184, N3157);
or OR3 (N3185, N3178, N473, N938);
xor XOR2 (N3186, N3183, N2600);
and AND3 (N3187, N3186, N1074, N2822);
buf BUF1 (N3188, N3179);
buf BUF1 (N3189, N3180);
xor XOR2 (N3190, N3176, N2428);
not NOT1 (N3191, N3177);
xor XOR2 (N3192, N3184, N3044);
nand NAND2 (N3193, N3192, N1357);
not NOT1 (N3194, N3169);
nor NOR3 (N3195, N3185, N2419, N1398);
nand NAND2 (N3196, N3195, N1220);
nand NAND2 (N3197, N3193, N1379);
nand NAND4 (N3198, N3190, N2292, N823, N1407);
buf BUF1 (N3199, N3196);
xor XOR2 (N3200, N3188, N3136);
nor NOR2 (N3201, N3181, N2781);
buf BUF1 (N3202, N3197);
nor NOR2 (N3203, N3202, N1089);
nand NAND4 (N3204, N3187, N1879, N608, N1847);
or OR3 (N3205, N3203, N2144, N441);
buf BUF1 (N3206, N3201);
xor XOR2 (N3207, N3200, N449);
buf BUF1 (N3208, N3205);
not NOT1 (N3209, N3194);
and AND2 (N3210, N3191, N1363);
nand NAND4 (N3211, N3208, N1324, N853, N3137);
nand NAND4 (N3212, N3204, N2249, N1024, N239);
buf BUF1 (N3213, N3206);
and AND3 (N3214, N3209, N136, N2195);
buf BUF1 (N3215, N3214);
buf BUF1 (N3216, N3199);
buf BUF1 (N3217, N3207);
or OR3 (N3218, N3216, N1351, N36);
and AND3 (N3219, N3189, N2478, N380);
nor NOR3 (N3220, N3217, N42, N660);
and AND4 (N3221, N3212, N2397, N1602, N3136);
nand NAND3 (N3222, N3220, N424, N2275);
nand NAND3 (N3223, N3219, N1624, N1173);
or OR2 (N3224, N3218, N2108);
and AND4 (N3225, N3159, N219, N223, N2511);
not NOT1 (N3226, N3198);
buf BUF1 (N3227, N3222);
and AND4 (N3228, N3224, N3005, N510, N1710);
not NOT1 (N3229, N3225);
or OR4 (N3230, N3210, N1744, N89, N3034);
nand NAND3 (N3231, N3230, N778, N2870);
buf BUF1 (N3232, N3213);
nand NAND3 (N3233, N3231, N2375, N2882);
nand NAND2 (N3234, N3228, N1300);
or OR3 (N3235, N3226, N619, N399);
buf BUF1 (N3236, N3233);
nor NOR3 (N3237, N3235, N620, N1326);
nand NAND2 (N3238, N3227, N2163);
not NOT1 (N3239, N3223);
not NOT1 (N3240, N3229);
nor NOR4 (N3241, N3240, N1740, N235, N3124);
not NOT1 (N3242, N3241);
buf BUF1 (N3243, N3215);
nand NAND2 (N3244, N3237, N3106);
or OR2 (N3245, N3239, N2812);
nor NOR4 (N3246, N3234, N2033, N168, N2271);
or OR3 (N3247, N3236, N2507, N2661);
or OR3 (N3248, N3232, N827, N3154);
buf BUF1 (N3249, N3243);
nand NAND4 (N3250, N3221, N806, N236, N488);
nor NOR4 (N3251, N3250, N3081, N2287, N1485);
not NOT1 (N3252, N3242);
buf BUF1 (N3253, N3238);
buf BUF1 (N3254, N3248);
nand NAND4 (N3255, N3254, N1828, N688, N1132);
or OR2 (N3256, N3244, N1300);
and AND2 (N3257, N3246, N1025);
buf BUF1 (N3258, N3255);
nor NOR3 (N3259, N3245, N1935, N1613);
or OR3 (N3260, N3259, N433, N1022);
nand NAND2 (N3261, N3257, N2766);
and AND2 (N3262, N3247, N103);
or OR4 (N3263, N3260, N3178, N726, N1603);
or OR3 (N3264, N3258, N3072, N1022);
not NOT1 (N3265, N3256);
nor NOR2 (N3266, N3253, N604);
buf BUF1 (N3267, N3249);
nand NAND2 (N3268, N3262, N2202);
or OR4 (N3269, N3266, N1041, N572, N1620);
not NOT1 (N3270, N3269);
and AND3 (N3271, N3211, N2594, N2503);
not NOT1 (N3272, N3252);
buf BUF1 (N3273, N3270);
or OR2 (N3274, N3273, N2);
xor XOR2 (N3275, N3272, N425);
not NOT1 (N3276, N3261);
not NOT1 (N3277, N3271);
not NOT1 (N3278, N3264);
buf BUF1 (N3279, N3251);
buf BUF1 (N3280, N3274);
or OR4 (N3281, N3263, N1609, N963, N1971);
or OR4 (N3282, N3265, N2145, N466, N124);
xor XOR2 (N3283, N3276, N2355);
or OR2 (N3284, N3280, N3281);
nand NAND3 (N3285, N402, N2366, N2328);
xor XOR2 (N3286, N3284, N3277);
or OR3 (N3287, N1642, N2860, N1014);
and AND4 (N3288, N3267, N2344, N3128, N1055);
or OR4 (N3289, N3279, N384, N101, N2065);
xor XOR2 (N3290, N3268, N2777);
or OR3 (N3291, N3282, N1917, N3010);
xor XOR2 (N3292, N3283, N2034);
nand NAND3 (N3293, N3289, N2244, N119);
nand NAND4 (N3294, N3290, N2227, N2360, N2832);
not NOT1 (N3295, N3291);
not NOT1 (N3296, N3295);
nand NAND3 (N3297, N3287, N3159, N214);
and AND4 (N3298, N3275, N1417, N1639, N2387);
or OR3 (N3299, N3285, N2106, N833);
and AND3 (N3300, N3297, N626, N1237);
not NOT1 (N3301, N3286);
and AND2 (N3302, N3301, N2172);
and AND4 (N3303, N3293, N334, N1122, N2627);
nor NOR3 (N3304, N3302, N1342, N2796);
and AND2 (N3305, N3296, N768);
buf BUF1 (N3306, N3294);
buf BUF1 (N3307, N3292);
buf BUF1 (N3308, N3306);
nand NAND3 (N3309, N3288, N896, N418);
nor NOR3 (N3310, N3304, N2847, N2065);
buf BUF1 (N3311, N3300);
not NOT1 (N3312, N3298);
nor NOR2 (N3313, N3309, N1242);
nand NAND3 (N3314, N3278, N3293, N1153);
or OR4 (N3315, N3303, N1752, N949, N2017);
and AND2 (N3316, N3315, N131);
nand NAND3 (N3317, N3314, N349, N1297);
not NOT1 (N3318, N3307);
or OR2 (N3319, N3316, N595);
nand NAND3 (N3320, N3313, N227, N998);
nand NAND3 (N3321, N3320, N210, N2135);
or OR3 (N3322, N3311, N2567, N1287);
nor NOR2 (N3323, N3319, N1918);
buf BUF1 (N3324, N3299);
xor XOR2 (N3325, N3310, N619);
and AND3 (N3326, N3312, N3115, N1045);
buf BUF1 (N3327, N3324);
nor NOR2 (N3328, N3317, N895);
and AND4 (N3329, N3322, N3282, N1762, N319);
and AND4 (N3330, N3323, N1210, N1373, N2102);
nand NAND4 (N3331, N3305, N2676, N807, N660);
nor NOR4 (N3332, N3330, N1330, N124, N2555);
not NOT1 (N3333, N3328);
buf BUF1 (N3334, N3308);
not NOT1 (N3335, N3333);
or OR2 (N3336, N3327, N3246);
or OR2 (N3337, N3329, N1843);
xor XOR2 (N3338, N3337, N94);
nor NOR2 (N3339, N3332, N1932);
or OR4 (N3340, N3335, N2736, N1997, N1138);
or OR4 (N3341, N3318, N374, N1978, N1704);
not NOT1 (N3342, N3338);
and AND2 (N3343, N3340, N822);
xor XOR2 (N3344, N3343, N931);
nand NAND2 (N3345, N3331, N1077);
nand NAND2 (N3346, N3321, N2380);
nand NAND2 (N3347, N3341, N2947);
nor NOR2 (N3348, N3326, N1297);
xor XOR2 (N3349, N3334, N110);
or OR4 (N3350, N3339, N2497, N2279, N2055);
and AND3 (N3351, N3346, N2604, N835);
and AND4 (N3352, N3342, N1587, N1499, N1110);
not NOT1 (N3353, N3347);
nand NAND3 (N3354, N3348, N62, N3268);
nor NOR3 (N3355, N3325, N719, N270);
not NOT1 (N3356, N3355);
not NOT1 (N3357, N3352);
nand NAND4 (N3358, N3345, N3217, N2725, N807);
or OR4 (N3359, N3358, N791, N556, N521);
not NOT1 (N3360, N3356);
not NOT1 (N3361, N3353);
xor XOR2 (N3362, N3360, N2779);
nor NOR3 (N3363, N3350, N3098, N1087);
xor XOR2 (N3364, N3363, N766);
nand NAND2 (N3365, N3349, N439);
nor NOR2 (N3366, N3364, N2737);
buf BUF1 (N3367, N3354);
nor NOR3 (N3368, N3359, N492, N1003);
and AND4 (N3369, N3336, N279, N518, N1116);
xor XOR2 (N3370, N3369, N3319);
or OR3 (N3371, N3366, N1715, N701);
buf BUF1 (N3372, N3368);
and AND3 (N3373, N3351, N3118, N506);
buf BUF1 (N3374, N3370);
not NOT1 (N3375, N3373);
nand NAND2 (N3376, N3372, N726);
buf BUF1 (N3377, N3344);
nor NOR3 (N3378, N3371, N2111, N2213);
nor NOR4 (N3379, N3357, N641, N2516, N2549);
buf BUF1 (N3380, N3379);
not NOT1 (N3381, N3380);
or OR2 (N3382, N3361, N977);
nand NAND4 (N3383, N3381, N2138, N2727, N964);
not NOT1 (N3384, N3362);
xor XOR2 (N3385, N3365, N1382);
xor XOR2 (N3386, N3374, N2512);
and AND3 (N3387, N3384, N1114, N1114);
not NOT1 (N3388, N3386);
nor NOR2 (N3389, N3387, N2461);
not NOT1 (N3390, N3367);
or OR2 (N3391, N3383, N1194);
nand NAND2 (N3392, N3375, N2632);
and AND2 (N3393, N3385, N2622);
and AND2 (N3394, N3376, N1084);
nor NOR3 (N3395, N3393, N2010, N1515);
nand NAND2 (N3396, N3389, N333);
buf BUF1 (N3397, N3382);
or OR3 (N3398, N3378, N1162, N2903);
nor NOR2 (N3399, N3398, N1322);
buf BUF1 (N3400, N3390);
and AND4 (N3401, N3377, N1633, N1799, N3309);
and AND3 (N3402, N3396, N2395, N3370);
xor XOR2 (N3403, N3401, N87);
xor XOR2 (N3404, N3391, N2057);
xor XOR2 (N3405, N3397, N2029);
or OR3 (N3406, N3394, N2209, N2104);
nand NAND2 (N3407, N3392, N3172);
not NOT1 (N3408, N3406);
nand NAND2 (N3409, N3407, N1065);
xor XOR2 (N3410, N3395, N1487);
nand NAND4 (N3411, N3408, N368, N2351, N3012);
or OR2 (N3412, N3411, N2708);
not NOT1 (N3413, N3402);
not NOT1 (N3414, N3388);
or OR2 (N3415, N3410, N37);
nor NOR2 (N3416, N3415, N1540);
xor XOR2 (N3417, N3403, N946);
not NOT1 (N3418, N3405);
buf BUF1 (N3419, N3413);
not NOT1 (N3420, N3414);
not NOT1 (N3421, N3416);
xor XOR2 (N3422, N3417, N2364);
nand NAND2 (N3423, N3409, N2831);
and AND4 (N3424, N3400, N461, N2336, N3368);
nor NOR4 (N3425, N3399, N31, N3169, N1999);
xor XOR2 (N3426, N3404, N1697);
xor XOR2 (N3427, N3412, N2582);
buf BUF1 (N3428, N3421);
nor NOR4 (N3429, N3425, N2740, N1283, N1027);
nor NOR3 (N3430, N3423, N1366, N1859);
buf BUF1 (N3431, N3419);
and AND2 (N3432, N3422, N2075);
nor NOR3 (N3433, N3424, N22, N1174);
not NOT1 (N3434, N3428);
xor XOR2 (N3435, N3432, N2430);
nand NAND3 (N3436, N3434, N1371, N1224);
nor NOR3 (N3437, N3436, N2840, N761);
nand NAND3 (N3438, N3433, N3123, N1756);
not NOT1 (N3439, N3418);
nand NAND3 (N3440, N3435, N1007, N349);
or OR3 (N3441, N3440, N2735, N1270);
nor NOR4 (N3442, N3427, N907, N2428, N123);
and AND3 (N3443, N3438, N2696, N456);
xor XOR2 (N3444, N3426, N1545);
and AND4 (N3445, N3431, N515, N480, N2515);
nor NOR3 (N3446, N3439, N2606, N3350);
buf BUF1 (N3447, N3430);
nor NOR3 (N3448, N3446, N1999, N1231);
nand NAND4 (N3449, N3445, N1278, N1278, N1330);
nand NAND4 (N3450, N3437, N3227, N3153, N2397);
nand NAND2 (N3451, N3420, N1796);
xor XOR2 (N3452, N3444, N2556);
and AND3 (N3453, N3448, N1201, N3232);
nand NAND3 (N3454, N3441, N2562, N502);
xor XOR2 (N3455, N3451, N1998);
nor NOR2 (N3456, N3442, N1960);
nor NOR2 (N3457, N3453, N2352);
or OR2 (N3458, N3447, N1571);
nand NAND3 (N3459, N3454, N3387, N1973);
buf BUF1 (N3460, N3456);
not NOT1 (N3461, N3459);
xor XOR2 (N3462, N3457, N857);
buf BUF1 (N3463, N3462);
buf BUF1 (N3464, N3458);
nor NOR3 (N3465, N3455, N1373, N2651);
and AND2 (N3466, N3461, N116);
and AND4 (N3467, N3449, N2509, N972, N1492);
xor XOR2 (N3468, N3467, N3442);
nor NOR2 (N3469, N3463, N1754);
not NOT1 (N3470, N3466);
and AND2 (N3471, N3465, N228);
nand NAND3 (N3472, N3468, N3356, N1440);
not NOT1 (N3473, N3470);
or OR3 (N3474, N3443, N1980, N2265);
nor NOR4 (N3475, N3464, N695, N2081, N2030);
not NOT1 (N3476, N3475);
or OR3 (N3477, N3469, N2539, N306);
or OR3 (N3478, N3429, N3407, N2755);
not NOT1 (N3479, N3460);
nor NOR3 (N3480, N3476, N3235, N1781);
not NOT1 (N3481, N3479);
nand NAND3 (N3482, N3471, N2939, N2678);
nor NOR4 (N3483, N3474, N515, N186, N2101);
nand NAND2 (N3484, N3452, N1757);
or OR2 (N3485, N3477, N3059);
xor XOR2 (N3486, N3481, N2539);
or OR3 (N3487, N3473, N3213, N27);
buf BUF1 (N3488, N3480);
buf BUF1 (N3489, N3478);
or OR3 (N3490, N3450, N443, N1377);
nor NOR3 (N3491, N3488, N2917, N2060);
and AND2 (N3492, N3482, N2091);
or OR2 (N3493, N3491, N206);
nor NOR3 (N3494, N3490, N320, N845);
nor NOR4 (N3495, N3486, N661, N2013, N3317);
xor XOR2 (N3496, N3492, N2590);
nand NAND3 (N3497, N3487, N2757, N708);
nor NOR2 (N3498, N3483, N2707);
buf BUF1 (N3499, N3493);
and AND2 (N3500, N3499, N2422);
nand NAND3 (N3501, N3472, N1604, N3401);
buf BUF1 (N3502, N3497);
xor XOR2 (N3503, N3500, N3098);
buf BUF1 (N3504, N3496);
buf BUF1 (N3505, N3503);
buf BUF1 (N3506, N3489);
nand NAND3 (N3507, N3494, N245, N2386);
xor XOR2 (N3508, N3507, N3311);
buf BUF1 (N3509, N3506);
buf BUF1 (N3510, N3505);
nor NOR2 (N3511, N3509, N2119);
or OR4 (N3512, N3502, N948, N2106, N605);
not NOT1 (N3513, N3508);
and AND2 (N3514, N3501, N2172);
nor NOR2 (N3515, N3513, N2331);
nor NOR3 (N3516, N3515, N553, N2393);
buf BUF1 (N3517, N3484);
nor NOR2 (N3518, N3511, N349);
nor NOR4 (N3519, N3485, N2534, N2428, N1036);
nand NAND4 (N3520, N3498, N1632, N3379, N463);
not NOT1 (N3521, N3520);
not NOT1 (N3522, N3521);
not NOT1 (N3523, N3495);
xor XOR2 (N3524, N3522, N1356);
not NOT1 (N3525, N3519);
and AND4 (N3526, N3525, N1639, N420, N1939);
or OR4 (N3527, N3504, N2343, N1262, N890);
not NOT1 (N3528, N3517);
and AND2 (N3529, N3524, N2696);
nor NOR2 (N3530, N3518, N1991);
nand NAND3 (N3531, N3530, N188, N2032);
and AND2 (N3532, N3512, N2455);
buf BUF1 (N3533, N3514);
or OR2 (N3534, N3529, N2093);
and AND4 (N3535, N3528, N345, N2868, N18);
not NOT1 (N3536, N3535);
buf BUF1 (N3537, N3523);
nor NOR2 (N3538, N3510, N2188);
not NOT1 (N3539, N3536);
xor XOR2 (N3540, N3538, N2299);
not NOT1 (N3541, N3526);
buf BUF1 (N3542, N3537);
buf BUF1 (N3543, N3527);
nor NOR3 (N3544, N3531, N2007, N47);
nor NOR2 (N3545, N3540, N2948);
buf BUF1 (N3546, N3545);
nor NOR3 (N3547, N3541, N1551, N1993);
nand NAND3 (N3548, N3534, N63, N1471);
nor NOR4 (N3549, N3542, N840, N1491, N2078);
xor XOR2 (N3550, N3546, N40);
xor XOR2 (N3551, N3533, N3467);
nand NAND2 (N3552, N3548, N1934);
buf BUF1 (N3553, N3532);
and AND4 (N3554, N3516, N2460, N3075, N1170);
xor XOR2 (N3555, N3543, N1377);
nand NAND4 (N3556, N3552, N2772, N652, N2991);
and AND4 (N3557, N3551, N3354, N1148, N39);
nand NAND2 (N3558, N3547, N2393);
and AND4 (N3559, N3554, N1349, N685, N3091);
not NOT1 (N3560, N3550);
nand NAND4 (N3561, N3539, N487, N3320, N2047);
nor NOR3 (N3562, N3559, N286, N679);
buf BUF1 (N3563, N3561);
and AND2 (N3564, N3562, N2916);
not NOT1 (N3565, N3544);
nor NOR3 (N3566, N3553, N431, N1540);
nor NOR2 (N3567, N3566, N2081);
xor XOR2 (N3568, N3555, N1319);
or OR3 (N3569, N3557, N1001, N432);
nand NAND4 (N3570, N3556, N2212, N1418, N1983);
nor NOR2 (N3571, N3565, N2143);
nor NOR4 (N3572, N3563, N2566, N2132, N2466);
xor XOR2 (N3573, N3572, N1216);
nand NAND2 (N3574, N3560, N2725);
xor XOR2 (N3575, N3571, N17);
xor XOR2 (N3576, N3569, N3061);
not NOT1 (N3577, N3576);
xor XOR2 (N3578, N3573, N2177);
or OR3 (N3579, N3564, N212, N1879);
nand NAND4 (N3580, N3558, N366, N548, N461);
nor NOR3 (N3581, N3580, N170, N937);
and AND2 (N3582, N3575, N2704);
or OR2 (N3583, N3574, N3290);
xor XOR2 (N3584, N3581, N265);
nor NOR4 (N3585, N3568, N1909, N789, N1720);
or OR2 (N3586, N3549, N2765);
buf BUF1 (N3587, N3570);
nor NOR2 (N3588, N3577, N1870);
and AND3 (N3589, N3567, N20, N1706);
xor XOR2 (N3590, N3586, N1184);
or OR4 (N3591, N3582, N1473, N3211, N2330);
nand NAND2 (N3592, N3590, N3300);
not NOT1 (N3593, N3584);
nor NOR4 (N3594, N3587, N864, N404, N2687);
xor XOR2 (N3595, N3588, N3465);
not NOT1 (N3596, N3583);
xor XOR2 (N3597, N3595, N2895);
xor XOR2 (N3598, N3578, N3283);
nand NAND2 (N3599, N3592, N3366);
xor XOR2 (N3600, N3591, N574);
buf BUF1 (N3601, N3599);
and AND4 (N3602, N3598, N811, N2280, N1604);
nand NAND3 (N3603, N3589, N2951, N3460);
and AND2 (N3604, N3585, N1988);
and AND3 (N3605, N3601, N2197, N1272);
xor XOR2 (N3606, N3600, N1600);
xor XOR2 (N3607, N3579, N1810);
or OR2 (N3608, N3594, N3232);
nand NAND4 (N3609, N3603, N1237, N98, N2307);
xor XOR2 (N3610, N3602, N1783);
nand NAND3 (N3611, N3596, N1628, N547);
and AND2 (N3612, N3593, N3330);
not NOT1 (N3613, N3608);
buf BUF1 (N3614, N3605);
buf BUF1 (N3615, N3607);
buf BUF1 (N3616, N3611);
xor XOR2 (N3617, N3614, N1058);
and AND4 (N3618, N3606, N1155, N2538, N3414);
buf BUF1 (N3619, N3604);
buf BUF1 (N3620, N3597);
buf BUF1 (N3621, N3620);
and AND3 (N3622, N3619, N1592, N1622);
xor XOR2 (N3623, N3613, N1576);
buf BUF1 (N3624, N3615);
nor NOR2 (N3625, N3617, N2715);
nand NAND4 (N3626, N3618, N3189, N2958, N974);
buf BUF1 (N3627, N3612);
and AND2 (N3628, N3627, N1141);
buf BUF1 (N3629, N3625);
or OR2 (N3630, N3626, N1060);
xor XOR2 (N3631, N3609, N240);
buf BUF1 (N3632, N3629);
and AND4 (N3633, N3632, N660, N2767, N93);
nor NOR4 (N3634, N3623, N2996, N956, N3386);
and AND3 (N3635, N3634, N3328, N3385);
buf BUF1 (N3636, N3628);
buf BUF1 (N3637, N3616);
buf BUF1 (N3638, N3631);
nor NOR4 (N3639, N3624, N2280, N1732, N1174);
xor XOR2 (N3640, N3630, N1650);
nand NAND2 (N3641, N3636, N984);
not NOT1 (N3642, N3640);
or OR3 (N3643, N3641, N2987, N669);
xor XOR2 (N3644, N3639, N2424);
nor NOR3 (N3645, N3643, N2421, N3245);
nand NAND3 (N3646, N3637, N1090, N2202);
and AND2 (N3647, N3644, N3556);
or OR4 (N3648, N3642, N3120, N504, N2041);
xor XOR2 (N3649, N3647, N2606);
and AND2 (N3650, N3649, N2938);
not NOT1 (N3651, N3648);
buf BUF1 (N3652, N3638);
or OR4 (N3653, N3645, N1489, N2497, N1074);
nor NOR2 (N3654, N3652, N683);
buf BUF1 (N3655, N3646);
nor NOR3 (N3656, N3651, N791, N1451);
not NOT1 (N3657, N3655);
nand NAND4 (N3658, N3656, N3073, N290, N2395);
buf BUF1 (N3659, N3621);
xor XOR2 (N3660, N3635, N64);
or OR2 (N3661, N3622, N760);
or OR2 (N3662, N3657, N8);
not NOT1 (N3663, N3633);
and AND3 (N3664, N3658, N119, N2807);
nand NAND2 (N3665, N3650, N1616);
buf BUF1 (N3666, N3660);
or OR3 (N3667, N3661, N3130, N681);
buf BUF1 (N3668, N3667);
nand NAND3 (N3669, N3663, N385, N1475);
xor XOR2 (N3670, N3665, N712);
nand NAND3 (N3671, N3670, N1351, N1313);
xor XOR2 (N3672, N3668, N69);
xor XOR2 (N3673, N3659, N295);
nand NAND4 (N3674, N3662, N3054, N2839, N1918);
buf BUF1 (N3675, N3666);
not NOT1 (N3676, N3654);
buf BUF1 (N3677, N3664);
and AND3 (N3678, N3671, N608, N597);
nand NAND3 (N3679, N3674, N131, N2546);
xor XOR2 (N3680, N3676, N2259);
or OR4 (N3681, N3678, N941, N180, N1689);
nor NOR4 (N3682, N3673, N3595, N589, N1093);
and AND3 (N3683, N3681, N1279, N2406);
and AND2 (N3684, N3679, N1760);
not NOT1 (N3685, N3684);
xor XOR2 (N3686, N3669, N2982);
and AND4 (N3687, N3682, N1513, N2534, N781);
nand NAND4 (N3688, N3675, N1021, N2628, N1211);
xor XOR2 (N3689, N3686, N1059);
and AND3 (N3690, N3680, N1971, N762);
nand NAND2 (N3691, N3685, N3550);
and AND2 (N3692, N3610, N805);
and AND2 (N3693, N3689, N3507);
not NOT1 (N3694, N3691);
and AND2 (N3695, N3688, N2935);
nor NOR2 (N3696, N3687, N366);
buf BUF1 (N3697, N3696);
and AND3 (N3698, N3653, N1682, N2138);
nand NAND4 (N3699, N3690, N136, N1058, N326);
nor NOR3 (N3700, N3694, N1258, N2418);
or OR4 (N3701, N3698, N599, N588, N2471);
and AND2 (N3702, N3699, N1087);
or OR2 (N3703, N3701, N993);
nor NOR3 (N3704, N3692, N1836, N814);
xor XOR2 (N3705, N3672, N849);
buf BUF1 (N3706, N3697);
not NOT1 (N3707, N3704);
buf BUF1 (N3708, N3706);
nor NOR4 (N3709, N3707, N2277, N2476, N3240);
and AND2 (N3710, N3695, N1268);
buf BUF1 (N3711, N3693);
or OR3 (N3712, N3708, N2160, N3528);
not NOT1 (N3713, N3712);
or OR2 (N3714, N3677, N624);
xor XOR2 (N3715, N3705, N2416);
nand NAND3 (N3716, N3715, N1426, N453);
or OR3 (N3717, N3714, N1001, N1280);
buf BUF1 (N3718, N3709);
nor NOR4 (N3719, N3713, N3000, N1654, N3134);
nand NAND2 (N3720, N3700, N2032);
and AND2 (N3721, N3703, N788);
not NOT1 (N3722, N3719);
buf BUF1 (N3723, N3683);
nand NAND2 (N3724, N3716, N1802);
nand NAND3 (N3725, N3721, N1994, N1098);
nor NOR2 (N3726, N3724, N1904);
or OR2 (N3727, N3702, N787);
nand NAND2 (N3728, N3723, N2205);
nand NAND2 (N3729, N3727, N1103);
nor NOR3 (N3730, N3725, N1706, N866);
nor NOR4 (N3731, N3730, N810, N1289, N3212);
xor XOR2 (N3732, N3731, N394);
buf BUF1 (N3733, N3710);
nand NAND2 (N3734, N3717, N2339);
xor XOR2 (N3735, N3728, N3115);
buf BUF1 (N3736, N3734);
xor XOR2 (N3737, N3733, N79);
not NOT1 (N3738, N3718);
nand NAND2 (N3739, N3720, N1559);
nor NOR4 (N3740, N3735, N3619, N3201, N750);
not NOT1 (N3741, N3738);
nor NOR2 (N3742, N3736, N2276);
nand NAND4 (N3743, N3726, N257, N425, N2428);
not NOT1 (N3744, N3739);
nand NAND3 (N3745, N3743, N2664, N1939);
nor NOR3 (N3746, N3742, N3017, N2901);
xor XOR2 (N3747, N3722, N1986);
or OR4 (N3748, N3741, N1606, N2760, N2118);
not NOT1 (N3749, N3737);
nand NAND2 (N3750, N3749, N691);
and AND2 (N3751, N3747, N2833);
xor XOR2 (N3752, N3744, N135);
nand NAND2 (N3753, N3750, N3491);
nand NAND3 (N3754, N3711, N867, N1763);
or OR2 (N3755, N3751, N2416);
buf BUF1 (N3756, N3752);
nand NAND2 (N3757, N3753, N2907);
buf BUF1 (N3758, N3740);
nor NOR3 (N3759, N3757, N2564, N701);
buf BUF1 (N3760, N3732);
nor NOR3 (N3761, N3760, N17, N2383);
nor NOR4 (N3762, N3756, N3730, N3755, N3251);
nor NOR2 (N3763, N1950, N1876);
not NOT1 (N3764, N3758);
or OR4 (N3765, N3729, N2272, N3551, N3066);
buf BUF1 (N3766, N3765);
and AND3 (N3767, N3746, N1640, N2164);
and AND4 (N3768, N3761, N48, N347, N2385);
buf BUF1 (N3769, N3767);
or OR4 (N3770, N3763, N3000, N1082, N619);
nand NAND4 (N3771, N3770, N1038, N554, N2072);
xor XOR2 (N3772, N3745, N1624);
nor NOR2 (N3773, N3754, N1984);
and AND3 (N3774, N3764, N2713, N964);
or OR3 (N3775, N3766, N257, N2526);
and AND2 (N3776, N3769, N2307);
nand NAND4 (N3777, N3762, N1857, N2141, N2067);
not NOT1 (N3778, N3773);
buf BUF1 (N3779, N3772);
nor NOR4 (N3780, N3771, N2932, N375, N177);
or OR4 (N3781, N3759, N1532, N1769, N1411);
nor NOR4 (N3782, N3775, N1324, N3521, N1042);
nor NOR4 (N3783, N3779, N2641, N82, N780);
nand NAND2 (N3784, N3748, N3332);
not NOT1 (N3785, N3783);
xor XOR2 (N3786, N3777, N1670);
or OR2 (N3787, N3785, N2392);
not NOT1 (N3788, N3768);
or OR2 (N3789, N3786, N1369);
buf BUF1 (N3790, N3778);
and AND4 (N3791, N3781, N2060, N2696, N24);
and AND2 (N3792, N3788, N658);
or OR3 (N3793, N3787, N2705, N3743);
not NOT1 (N3794, N3782);
nor NOR3 (N3795, N3793, N1015, N949);
nand NAND2 (N3796, N3776, N84);
and AND4 (N3797, N3792, N1028, N200, N1595);
or OR3 (N3798, N3774, N2400, N828);
nor NOR3 (N3799, N3795, N171, N894);
xor XOR2 (N3800, N3791, N2706);
or OR2 (N3801, N3796, N307);
not NOT1 (N3802, N3801);
xor XOR2 (N3803, N3789, N2062);
buf BUF1 (N3804, N3798);
nor NOR4 (N3805, N3803, N2474, N3107, N479);
nand NAND2 (N3806, N3802, N3535);
nand NAND3 (N3807, N3780, N2215, N3638);
nand NAND4 (N3808, N3806, N2481, N2244, N3318);
or OR4 (N3809, N3799, N2724, N2161, N652);
xor XOR2 (N3810, N3809, N2713);
nand NAND3 (N3811, N3797, N1450, N2220);
and AND3 (N3812, N3811, N2084, N2468);
or OR4 (N3813, N3790, N1028, N3528, N2035);
not NOT1 (N3814, N3813);
buf BUF1 (N3815, N3804);
nand NAND4 (N3816, N3794, N2103, N3780, N331);
and AND2 (N3817, N3784, N3035);
and AND4 (N3818, N3800, N972, N1697, N903);
nor NOR2 (N3819, N3818, N2877);
and AND3 (N3820, N3815, N2666, N3747);
xor XOR2 (N3821, N3820, N451);
buf BUF1 (N3822, N3816);
nand NAND2 (N3823, N3821, N762);
xor XOR2 (N3824, N3808, N3259);
buf BUF1 (N3825, N3823);
nor NOR2 (N3826, N3822, N796);
nand NAND3 (N3827, N3805, N572, N1571);
or OR2 (N3828, N3824, N2326);
buf BUF1 (N3829, N3819);
xor XOR2 (N3830, N3828, N3087);
nor NOR3 (N3831, N3812, N3786, N1419);
xor XOR2 (N3832, N3831, N1451);
buf BUF1 (N3833, N3817);
and AND3 (N3834, N3827, N649, N1532);
and AND3 (N3835, N3834, N1735, N1737);
xor XOR2 (N3836, N3825, N1978);
not NOT1 (N3837, N3832);
nand NAND3 (N3838, N3826, N2141, N2488);
nor NOR3 (N3839, N3833, N2471, N3024);
nor NOR3 (N3840, N3807, N1824, N2282);
and AND2 (N3841, N3835, N296);
nor NOR2 (N3842, N3841, N2855);
xor XOR2 (N3843, N3836, N3508);
xor XOR2 (N3844, N3810, N1259);
nand NAND3 (N3845, N3843, N2289, N356);
or OR2 (N3846, N3845, N3318);
or OR4 (N3847, N3830, N950, N2911, N1284);
not NOT1 (N3848, N3838);
or OR2 (N3849, N3848, N1999);
xor XOR2 (N3850, N3839, N937);
or OR3 (N3851, N3842, N1321, N935);
buf BUF1 (N3852, N3851);
not NOT1 (N3853, N3846);
nand NAND2 (N3854, N3847, N2021);
xor XOR2 (N3855, N3814, N3318);
nand NAND3 (N3856, N3849, N1259, N2255);
buf BUF1 (N3857, N3837);
and AND3 (N3858, N3854, N1153, N2197);
and AND4 (N3859, N3855, N3364, N1257, N2172);
buf BUF1 (N3860, N3857);
buf BUF1 (N3861, N3852);
not NOT1 (N3862, N3859);
nand NAND3 (N3863, N3858, N607, N964);
nor NOR3 (N3864, N3861, N404, N2310);
not NOT1 (N3865, N3850);
and AND2 (N3866, N3862, N3197);
and AND3 (N3867, N3863, N2591, N3558);
not NOT1 (N3868, N3853);
xor XOR2 (N3869, N3860, N95);
buf BUF1 (N3870, N3844);
buf BUF1 (N3871, N3864);
buf BUF1 (N3872, N3866);
buf BUF1 (N3873, N3856);
not NOT1 (N3874, N3867);
nor NOR4 (N3875, N3829, N2278, N184, N60);
xor XOR2 (N3876, N3865, N943);
xor XOR2 (N3877, N3840, N519);
buf BUF1 (N3878, N3873);
and AND2 (N3879, N3869, N3656);
nand NAND3 (N3880, N3878, N1385, N660);
or OR2 (N3881, N3870, N3854);
and AND2 (N3882, N3881, N2854);
not NOT1 (N3883, N3876);
xor XOR2 (N3884, N3871, N2349);
buf BUF1 (N3885, N3879);
or OR4 (N3886, N3875, N1406, N3795, N2095);
nor NOR3 (N3887, N3872, N2137, N1231);
or OR3 (N3888, N3884, N2863, N3422);
and AND4 (N3889, N3887, N3812, N1332, N2373);
buf BUF1 (N3890, N3880);
nor NOR4 (N3891, N3877, N3814, N3454, N1364);
xor XOR2 (N3892, N3883, N972);
and AND3 (N3893, N3891, N2889, N1128);
nor NOR2 (N3894, N3890, N2569);
nor NOR4 (N3895, N3868, N3031, N2642, N1881);
buf BUF1 (N3896, N3874);
buf BUF1 (N3897, N3889);
nor NOR3 (N3898, N3895, N1001, N2403);
not NOT1 (N3899, N3893);
or OR2 (N3900, N3897, N3517);
nand NAND3 (N3901, N3886, N1118, N281);
xor XOR2 (N3902, N3898, N2172);
not NOT1 (N3903, N3882);
nand NAND2 (N3904, N3900, N228);
nand NAND2 (N3905, N3902, N3138);
nand NAND3 (N3906, N3896, N3328, N676);
nor NOR3 (N3907, N3894, N2570, N3160);
not NOT1 (N3908, N3905);
or OR2 (N3909, N3892, N1938);
not NOT1 (N3910, N3899);
nand NAND3 (N3911, N3910, N2995, N1174);
or OR4 (N3912, N3907, N2075, N1224, N2775);
and AND4 (N3913, N3888, N3738, N1485, N1942);
xor XOR2 (N3914, N3885, N1457);
buf BUF1 (N3915, N3903);
nor NOR3 (N3916, N3909, N103, N1967);
buf BUF1 (N3917, N3904);
not NOT1 (N3918, N3915);
nor NOR3 (N3919, N3913, N3515, N645);
xor XOR2 (N3920, N3912, N3146);
not NOT1 (N3921, N3918);
nand NAND2 (N3922, N3917, N3212);
xor XOR2 (N3923, N3920, N1993);
xor XOR2 (N3924, N3919, N1166);
xor XOR2 (N3925, N3923, N2319);
nor NOR3 (N3926, N3921, N3338, N1744);
buf BUF1 (N3927, N3926);
and AND3 (N3928, N3908, N3778, N2354);
or OR4 (N3929, N3911, N3186, N2471, N899);
buf BUF1 (N3930, N3924);
and AND3 (N3931, N3929, N3550, N823);
and AND4 (N3932, N3914, N2027, N2873, N2279);
not NOT1 (N3933, N3922);
nand NAND3 (N3934, N3928, N2336, N1908);
or OR3 (N3935, N3916, N1604, N426);
nand NAND4 (N3936, N3901, N3319, N1081, N3653);
buf BUF1 (N3937, N3934);
not NOT1 (N3938, N3933);
buf BUF1 (N3939, N3906);
nand NAND3 (N3940, N3939, N3260, N3010);
buf BUF1 (N3941, N3935);
buf BUF1 (N3942, N3941);
buf BUF1 (N3943, N3930);
xor XOR2 (N3944, N3932, N3419);
xor XOR2 (N3945, N3931, N2313);
nor NOR2 (N3946, N3940, N2374);
or OR4 (N3947, N3946, N2853, N3547, N205);
nand NAND4 (N3948, N3943, N2849, N3849, N3148);
buf BUF1 (N3949, N3936);
or OR2 (N3950, N3947, N2954);
or OR3 (N3951, N3944, N1139, N3801);
buf BUF1 (N3952, N3945);
nand NAND2 (N3953, N3927, N1942);
nand NAND3 (N3954, N3948, N2262, N409);
nand NAND3 (N3955, N3951, N2147, N1745);
buf BUF1 (N3956, N3937);
or OR2 (N3957, N3955, N3930);
and AND3 (N3958, N3956, N1170, N1931);
not NOT1 (N3959, N3949);
and AND2 (N3960, N3942, N315);
and AND4 (N3961, N3958, N1161, N2843, N2551);
and AND2 (N3962, N3953, N1324);
and AND3 (N3963, N3959, N441, N202);
and AND2 (N3964, N3963, N3155);
and AND3 (N3965, N3964, N433, N1794);
and AND2 (N3966, N3938, N21);
and AND3 (N3967, N3966, N3928, N3840);
xor XOR2 (N3968, N3965, N1237);
nand NAND3 (N3969, N3968, N2498, N1389);
buf BUF1 (N3970, N3961);
nor NOR2 (N3971, N3950, N3508);
or OR2 (N3972, N3970, N463);
and AND4 (N3973, N3925, N1323, N1276, N3494);
nand NAND2 (N3974, N3971, N375);
nor NOR3 (N3975, N3952, N812, N3011);
xor XOR2 (N3976, N3960, N2910);
not NOT1 (N3977, N3962);
or OR3 (N3978, N3975, N886, N2436);
nor NOR4 (N3979, N3969, N461, N2303, N3851);
and AND2 (N3980, N3978, N3035);
nor NOR4 (N3981, N3967, N2085, N822, N3278);
buf BUF1 (N3982, N3977);
nor NOR2 (N3983, N3982, N1109);
and AND3 (N3984, N3954, N385, N3216);
and AND2 (N3985, N3981, N2439);
not NOT1 (N3986, N3976);
or OR2 (N3987, N3984, N2453);
xor XOR2 (N3988, N3980, N1192);
buf BUF1 (N3989, N3987);
not NOT1 (N3990, N3985);
buf BUF1 (N3991, N3983);
or OR3 (N3992, N3986, N2610, N633);
nand NAND4 (N3993, N3979, N2199, N2381, N2791);
nor NOR4 (N3994, N3988, N1758, N502, N3724);
nor NOR3 (N3995, N3994, N2340, N2788);
or OR2 (N3996, N3995, N3135);
buf BUF1 (N3997, N3990);
buf BUF1 (N3998, N3989);
nor NOR4 (N3999, N3998, N121, N279, N3767);
and AND3 (N4000, N3973, N629, N3468);
or OR2 (N4001, N3999, N1811);
buf BUF1 (N4002, N4001);
or OR2 (N4003, N3993, N3098);
not NOT1 (N4004, N3991);
nand NAND2 (N4005, N3997, N329);
or OR2 (N4006, N3974, N448);
xor XOR2 (N4007, N4004, N3991);
buf BUF1 (N4008, N3996);
nand NAND2 (N4009, N4008, N699);
xor XOR2 (N4010, N4006, N2236);
nor NOR3 (N4011, N4003, N3515, N2789);
or OR2 (N4012, N3992, N388);
xor XOR2 (N4013, N3972, N615);
xor XOR2 (N4014, N3957, N2185);
nand NAND3 (N4015, N4002, N1590, N195);
xor XOR2 (N4016, N4015, N781);
buf BUF1 (N4017, N4011);
nor NOR3 (N4018, N4010, N680, N3258);
nor NOR4 (N4019, N4000, N263, N2765, N2998);
and AND4 (N4020, N4009, N2263, N3935, N1453);
endmodule