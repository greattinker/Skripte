// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;

output N25620,N25615,N25612,N25621,N25616,N25614,N25617,N25589,N25618,N25622;

and AND2 (N23, N1, N19);
not NOT1 (N24, N17);
not NOT1 (N25, N19);
buf BUF1 (N26, N25);
buf BUF1 (N27, N19);
not NOT1 (N28, N10);
buf BUF1 (N29, N9);
xor XOR2 (N30, N5, N28);
nand NAND4 (N31, N28, N1, N25, N25);
or OR3 (N32, N28, N27, N17);
buf BUF1 (N33, N3);
buf BUF1 (N34, N21);
nor NOR3 (N35, N17, N19, N23);
and AND3 (N36, N11, N5, N10);
or OR2 (N37, N34, N13);
not NOT1 (N38, N36);
not NOT1 (N39, N32);
and AND4 (N40, N26, N36, N29, N7);
or OR3 (N41, N35, N14, N31);
and AND3 (N42, N16, N19, N21);
or OR3 (N43, N42, N9, N10);
and AND4 (N44, N6, N31, N28, N19);
nor NOR2 (N45, N39, N2);
nor NOR4 (N46, N43, N21, N27, N3);
nand NAND4 (N47, N40, N13, N41, N36);
or OR4 (N48, N47, N15, N14, N7);
or OR3 (N49, N10, N18, N6);
xor XOR2 (N50, N30, N46);
nand NAND4 (N51, N29, N1, N12, N16);
nor NOR4 (N52, N48, N39, N44, N46);
not NOT1 (N53, N44);
buf BUF1 (N54, N33);
xor XOR2 (N55, N51, N1);
nand NAND2 (N56, N45, N48);
xor XOR2 (N57, N56, N23);
and AND3 (N58, N53, N13, N38);
and AND4 (N59, N53, N25, N55, N56);
or OR2 (N60, N38, N2);
or OR2 (N61, N54, N25);
and AND4 (N62, N59, N22, N3, N3);
xor XOR2 (N63, N61, N50);
nand NAND3 (N64, N37, N53, N60);
not NOT1 (N65, N13);
nor NOR3 (N66, N48, N45, N8);
nand NAND4 (N67, N52, N22, N63, N60);
nor NOR4 (N68, N6, N45, N42, N22);
nand NAND3 (N69, N24, N28, N17);
or OR4 (N70, N65, N38, N27, N69);
or OR3 (N71, N1, N10, N51);
not NOT1 (N72, N62);
or OR3 (N73, N49, N4, N48);
xor XOR2 (N74, N64, N52);
or OR4 (N75, N72, N51, N13, N36);
or OR4 (N76, N73, N7, N66, N17);
nand NAND3 (N77, N26, N66, N36);
or OR4 (N78, N67, N1, N5, N43);
xor XOR2 (N79, N74, N10);
buf BUF1 (N80, N70);
xor XOR2 (N81, N58, N1);
and AND3 (N82, N77, N78, N46);
and AND3 (N83, N54, N23, N57);
nor NOR2 (N84, N36, N67);
nand NAND2 (N85, N71, N70);
nor NOR4 (N86, N81, N60, N31, N12);
nor NOR4 (N87, N68, N54, N78, N31);
or OR2 (N88, N79, N58);
xor XOR2 (N89, N84, N57);
buf BUF1 (N90, N76);
buf BUF1 (N91, N90);
and AND4 (N92, N75, N72, N59, N70);
not NOT1 (N93, N83);
not NOT1 (N94, N93);
xor XOR2 (N95, N94, N20);
or OR4 (N96, N88, N48, N86, N80);
buf BUF1 (N97, N20);
buf BUF1 (N98, N14);
xor XOR2 (N99, N82, N26);
xor XOR2 (N100, N89, N58);
or OR3 (N101, N95, N73, N7);
and AND4 (N102, N101, N54, N69, N33);
buf BUF1 (N103, N96);
or OR4 (N104, N103, N26, N45, N37);
and AND2 (N105, N104, N45);
not NOT1 (N106, N105);
and AND4 (N107, N87, N30, N89, N11);
or OR4 (N108, N98, N48, N104, N38);
and AND4 (N109, N106, N15, N50, N61);
nor NOR3 (N110, N99, N44, N97);
buf BUF1 (N111, N76);
or OR4 (N112, N111, N23, N110, N11);
buf BUF1 (N113, N92);
buf BUF1 (N114, N85);
nand NAND3 (N115, N8, N91, N43);
xor XOR2 (N116, N50, N12);
nor NOR4 (N117, N100, N36, N17, N42);
not NOT1 (N118, N112);
xor XOR2 (N119, N107, N39);
not NOT1 (N120, N117);
xor XOR2 (N121, N119, N60);
xor XOR2 (N122, N109, N119);
nor NOR4 (N123, N114, N13, N32, N90);
not NOT1 (N124, N123);
buf BUF1 (N125, N115);
not NOT1 (N126, N118);
xor XOR2 (N127, N102, N24);
xor XOR2 (N128, N122, N60);
buf BUF1 (N129, N128);
buf BUF1 (N130, N108);
nor NOR2 (N131, N120, N39);
and AND2 (N132, N125, N1);
buf BUF1 (N133, N113);
not NOT1 (N134, N130);
not NOT1 (N135, N134);
xor XOR2 (N136, N116, N26);
nand NAND3 (N137, N124, N1, N116);
or OR3 (N138, N137, N84, N92);
buf BUF1 (N139, N129);
not NOT1 (N140, N127);
not NOT1 (N141, N140);
nand NAND4 (N142, N132, N131, N76, N101);
not NOT1 (N143, N16);
or OR3 (N144, N126, N61, N67);
nand NAND2 (N145, N138, N131);
nand NAND2 (N146, N139, N145);
or OR2 (N147, N57, N6);
not NOT1 (N148, N135);
buf BUF1 (N149, N121);
xor XOR2 (N150, N143, N81);
xor XOR2 (N151, N149, N42);
xor XOR2 (N152, N141, N62);
not NOT1 (N153, N133);
xor XOR2 (N154, N152, N86);
nor NOR2 (N155, N144, N24);
nand NAND4 (N156, N148, N148, N142, N12);
buf BUF1 (N157, N27);
or OR3 (N158, N155, N99, N77);
buf BUF1 (N159, N147);
or OR2 (N160, N159, N3);
nand NAND2 (N161, N151, N64);
buf BUF1 (N162, N161);
not NOT1 (N163, N158);
buf BUF1 (N164, N153);
nand NAND3 (N165, N146, N155, N162);
buf BUF1 (N166, N45);
not NOT1 (N167, N150);
not NOT1 (N168, N165);
buf BUF1 (N169, N160);
buf BUF1 (N170, N164);
or OR2 (N171, N136, N41);
xor XOR2 (N172, N166, N170);
and AND4 (N173, N60, N60, N72, N41);
or OR4 (N174, N172, N148, N76, N100);
nand NAND3 (N175, N157, N17, N73);
buf BUF1 (N176, N154);
xor XOR2 (N177, N163, N6);
and AND4 (N178, N175, N151, N52, N12);
nor NOR2 (N179, N167, N158);
nand NAND4 (N180, N178, N143, N35, N143);
xor XOR2 (N181, N180, N164);
nor NOR2 (N182, N173, N61);
xor XOR2 (N183, N181, N20);
nor NOR3 (N184, N156, N62, N68);
nand NAND2 (N185, N168, N32);
and AND4 (N186, N185, N149, N126, N62);
nand NAND2 (N187, N177, N144);
buf BUF1 (N188, N176);
xor XOR2 (N189, N182, N88);
nand NAND3 (N190, N186, N178, N187);
or OR2 (N191, N161, N168);
or OR2 (N192, N174, N166);
nand NAND4 (N193, N169, N115, N141, N64);
xor XOR2 (N194, N171, N127);
and AND4 (N195, N192, N97, N95, N152);
buf BUF1 (N196, N195);
buf BUF1 (N197, N183);
buf BUF1 (N198, N179);
buf BUF1 (N199, N188);
and AND4 (N200, N198, N89, N120, N42);
and AND4 (N201, N184, N111, N163, N41);
nor NOR3 (N202, N199, N150, N192);
or OR2 (N203, N197, N192);
or OR3 (N204, N200, N124, N155);
not NOT1 (N205, N202);
not NOT1 (N206, N193);
nor NOR4 (N207, N203, N76, N111, N35);
not NOT1 (N208, N206);
xor XOR2 (N209, N205, N45);
xor XOR2 (N210, N208, N180);
buf BUF1 (N211, N209);
buf BUF1 (N212, N194);
xor XOR2 (N213, N212, N37);
buf BUF1 (N214, N189);
not NOT1 (N215, N204);
or OR3 (N216, N213, N133, N115);
not NOT1 (N217, N216);
nor NOR4 (N218, N196, N178, N123, N43);
nand NAND3 (N219, N214, N52, N180);
nand NAND4 (N220, N219, N171, N156, N188);
xor XOR2 (N221, N207, N12);
nand NAND3 (N222, N221, N114, N157);
xor XOR2 (N223, N190, N88);
nand NAND2 (N224, N220, N37);
nor NOR4 (N225, N191, N132, N189, N74);
nor NOR3 (N226, N201, N70, N161);
not NOT1 (N227, N217);
nor NOR2 (N228, N224, N96);
buf BUF1 (N229, N215);
buf BUF1 (N230, N223);
not NOT1 (N231, N218);
nand NAND2 (N232, N229, N57);
nand NAND2 (N233, N227, N78);
nand NAND3 (N234, N233, N72, N18);
xor XOR2 (N235, N226, N13);
buf BUF1 (N236, N231);
nor NOR4 (N237, N230, N10, N172, N57);
not NOT1 (N238, N235);
buf BUF1 (N239, N210);
not NOT1 (N240, N225);
or OR3 (N241, N232, N204, N229);
nor NOR4 (N242, N240, N8, N77, N94);
nor NOR4 (N243, N222, N229, N117, N33);
xor XOR2 (N244, N243, N63);
nand NAND3 (N245, N211, N126, N229);
not NOT1 (N246, N237);
buf BUF1 (N247, N238);
or OR2 (N248, N245, N64);
or OR2 (N249, N246, N89);
nor NOR3 (N250, N247, N179, N200);
and AND4 (N251, N248, N131, N55, N119);
nor NOR4 (N252, N250, N135, N145, N63);
nor NOR3 (N253, N249, N229, N166);
and AND2 (N254, N242, N111);
xor XOR2 (N255, N239, N248);
nor NOR3 (N256, N241, N196, N1);
nand NAND4 (N257, N234, N119, N146, N228);
nand NAND4 (N258, N112, N98, N177, N233);
nor NOR3 (N259, N256, N246, N209);
nand NAND2 (N260, N254, N36);
nand NAND2 (N261, N252, N260);
nor NOR4 (N262, N185, N99, N141, N182);
or OR2 (N263, N261, N33);
or OR2 (N264, N263, N46);
and AND2 (N265, N262, N14);
xor XOR2 (N266, N258, N145);
and AND2 (N267, N251, N101);
buf BUF1 (N268, N265);
xor XOR2 (N269, N257, N252);
or OR4 (N270, N259, N24, N134, N78);
xor XOR2 (N271, N253, N232);
xor XOR2 (N272, N271, N24);
not NOT1 (N273, N244);
and AND2 (N274, N236, N244);
nand NAND4 (N275, N274, N54, N236, N235);
not NOT1 (N276, N272);
buf BUF1 (N277, N276);
xor XOR2 (N278, N273, N209);
not NOT1 (N279, N268);
or OR2 (N280, N278, N167);
not NOT1 (N281, N266);
and AND3 (N282, N279, N146, N155);
nor NOR4 (N283, N281, N273, N263, N280);
or OR4 (N284, N64, N131, N20, N144);
or OR3 (N285, N282, N16, N248);
or OR2 (N286, N269, N155);
xor XOR2 (N287, N270, N173);
or OR3 (N288, N285, N68, N48);
or OR4 (N289, N275, N280, N269, N140);
nor NOR2 (N290, N277, N157);
not NOT1 (N291, N284);
xor XOR2 (N292, N267, N43);
or OR2 (N293, N289, N150);
nand NAND2 (N294, N264, N267);
or OR2 (N295, N293, N249);
and AND2 (N296, N287, N65);
buf BUF1 (N297, N292);
nand NAND3 (N298, N294, N105, N104);
and AND3 (N299, N298, N174, N191);
and AND3 (N300, N283, N115, N43);
nand NAND3 (N301, N295, N23, N217);
nand NAND3 (N302, N291, N130, N121);
and AND4 (N303, N255, N267, N223, N166);
or OR4 (N304, N303, N44, N178, N117);
and AND4 (N305, N300, N11, N131, N162);
buf BUF1 (N306, N301);
xor XOR2 (N307, N290, N31);
not NOT1 (N308, N306);
and AND3 (N309, N288, N57, N152);
not NOT1 (N310, N309);
xor XOR2 (N311, N297, N177);
nand NAND2 (N312, N304, N61);
buf BUF1 (N313, N310);
and AND4 (N314, N299, N101, N252, N206);
xor XOR2 (N315, N311, N146);
not NOT1 (N316, N305);
nand NAND2 (N317, N314, N41);
xor XOR2 (N318, N313, N241);
and AND3 (N319, N315, N41, N146);
or OR4 (N320, N312, N62, N99, N27);
and AND4 (N321, N316, N250, N109, N157);
buf BUF1 (N322, N320);
xor XOR2 (N323, N286, N264);
or OR3 (N324, N296, N29, N93);
not NOT1 (N325, N317);
and AND4 (N326, N302, N251, N41, N136);
nand NAND3 (N327, N308, N180, N226);
and AND3 (N328, N324, N126, N58);
nand NAND3 (N329, N326, N139, N273);
xor XOR2 (N330, N321, N298);
not NOT1 (N331, N330);
nor NOR4 (N332, N328, N286, N161, N115);
or OR4 (N333, N307, N219, N39, N232);
buf BUF1 (N334, N331);
buf BUF1 (N335, N323);
xor XOR2 (N336, N329, N194);
nand NAND4 (N337, N333, N149, N226, N119);
nor NOR4 (N338, N334, N257, N104, N236);
not NOT1 (N339, N337);
buf BUF1 (N340, N325);
and AND3 (N341, N327, N18, N226);
or OR2 (N342, N336, N152);
not NOT1 (N343, N338);
xor XOR2 (N344, N340, N26);
or OR4 (N345, N342, N275, N271, N120);
buf BUF1 (N346, N322);
nor NOR4 (N347, N343, N299, N213, N158);
not NOT1 (N348, N345);
nor NOR3 (N349, N348, N93, N178);
nand NAND2 (N350, N339, N149);
xor XOR2 (N351, N319, N58);
xor XOR2 (N352, N349, N308);
buf BUF1 (N353, N350);
not NOT1 (N354, N318);
xor XOR2 (N355, N344, N341);
buf BUF1 (N356, N302);
xor XOR2 (N357, N347, N147);
or OR3 (N358, N335, N145, N129);
nand NAND3 (N359, N355, N194, N253);
nand NAND2 (N360, N353, N106);
buf BUF1 (N361, N360);
or OR2 (N362, N352, N267);
not NOT1 (N363, N357);
or OR2 (N364, N346, N61);
not NOT1 (N365, N363);
nor NOR3 (N366, N332, N121, N281);
nand NAND3 (N367, N358, N331, N183);
and AND3 (N368, N356, N326, N182);
buf BUF1 (N369, N365);
xor XOR2 (N370, N364, N291);
buf BUF1 (N371, N351);
nor NOR2 (N372, N370, N104);
nand NAND2 (N373, N362, N67);
nor NOR4 (N374, N373, N35, N189, N320);
buf BUF1 (N375, N372);
buf BUF1 (N376, N371);
nor NOR2 (N377, N374, N123);
and AND2 (N378, N377, N117);
nand NAND3 (N379, N375, N115, N106);
and AND3 (N380, N376, N189, N227);
not NOT1 (N381, N359);
or OR4 (N382, N378, N232, N209, N35);
not NOT1 (N383, N368);
buf BUF1 (N384, N379);
nand NAND3 (N385, N354, N151, N177);
not NOT1 (N386, N367);
buf BUF1 (N387, N369);
and AND4 (N388, N384, N312, N18, N119);
not NOT1 (N389, N366);
buf BUF1 (N390, N389);
xor XOR2 (N391, N385, N102);
buf BUF1 (N392, N386);
buf BUF1 (N393, N380);
xor XOR2 (N394, N383, N125);
buf BUF1 (N395, N390);
buf BUF1 (N396, N361);
xor XOR2 (N397, N387, N80);
or OR4 (N398, N388, N320, N386, N330);
not NOT1 (N399, N391);
buf BUF1 (N400, N398);
or OR4 (N401, N399, N11, N182, N331);
nand NAND2 (N402, N395, N349);
xor XOR2 (N403, N397, N171);
nor NOR4 (N404, N403, N53, N156, N398);
xor XOR2 (N405, N400, N43);
buf BUF1 (N406, N402);
buf BUF1 (N407, N401);
nand NAND2 (N408, N393, N295);
nor NOR2 (N409, N408, N25);
xor XOR2 (N410, N406, N286);
nor NOR3 (N411, N407, N347, N8);
or OR2 (N412, N396, N270);
xor XOR2 (N413, N410, N334);
nand NAND2 (N414, N405, N304);
buf BUF1 (N415, N412);
nand NAND4 (N416, N382, N5, N251, N107);
nor NOR4 (N417, N381, N168, N64, N159);
not NOT1 (N418, N413);
not NOT1 (N419, N411);
or OR3 (N420, N414, N227, N321);
not NOT1 (N421, N416);
buf BUF1 (N422, N421);
nand NAND3 (N423, N417, N157, N250);
nand NAND2 (N424, N394, N53);
xor XOR2 (N425, N424, N411);
buf BUF1 (N426, N418);
and AND2 (N427, N415, N414);
and AND2 (N428, N392, N387);
buf BUF1 (N429, N428);
xor XOR2 (N430, N422, N370);
xor XOR2 (N431, N429, N210);
or OR2 (N432, N427, N66);
and AND2 (N433, N423, N131);
nor NOR4 (N434, N420, N76, N60, N370);
buf BUF1 (N435, N426);
or OR2 (N436, N419, N288);
buf BUF1 (N437, N404);
and AND3 (N438, N425, N434, N223);
xor XOR2 (N439, N180, N219);
xor XOR2 (N440, N409, N438);
nor NOR3 (N441, N268, N99, N42);
buf BUF1 (N442, N432);
not NOT1 (N443, N436);
nor NOR3 (N444, N433, N295, N161);
not NOT1 (N445, N444);
nand NAND4 (N446, N445, N191, N1, N257);
or OR2 (N447, N430, N169);
buf BUF1 (N448, N435);
or OR4 (N449, N437, N222, N94, N366);
and AND4 (N450, N443, N360, N170, N256);
not NOT1 (N451, N448);
nor NOR4 (N452, N447, N77, N334, N309);
buf BUF1 (N453, N440);
nand NAND3 (N454, N439, N296, N59);
buf BUF1 (N455, N450);
buf BUF1 (N456, N449);
nor NOR2 (N457, N455, N91);
or OR3 (N458, N456, N419, N119);
nor NOR4 (N459, N446, N288, N394, N214);
nor NOR3 (N460, N452, N229, N275);
nand NAND3 (N461, N442, N421, N55);
nor NOR4 (N462, N458, N57, N293, N128);
xor XOR2 (N463, N457, N399);
nor NOR3 (N464, N461, N69, N251);
nand NAND3 (N465, N463, N154, N225);
or OR4 (N466, N462, N184, N183, N359);
buf BUF1 (N467, N464);
or OR3 (N468, N441, N202, N142);
nand NAND4 (N469, N431, N26, N312, N460);
xor XOR2 (N470, N17, N403);
nand NAND4 (N471, N466, N309, N466, N209);
nand NAND2 (N472, N467, N432);
or OR4 (N473, N468, N448, N383, N316);
xor XOR2 (N474, N470, N151);
xor XOR2 (N475, N459, N145);
buf BUF1 (N476, N472);
not NOT1 (N477, N473);
buf BUF1 (N478, N474);
nor NOR2 (N479, N465, N127);
nand NAND2 (N480, N453, N406);
buf BUF1 (N481, N451);
not NOT1 (N482, N480);
xor XOR2 (N483, N477, N26);
nand NAND3 (N484, N483, N40, N366);
or OR4 (N485, N478, N345, N151, N249);
not NOT1 (N486, N484);
nor NOR4 (N487, N454, N9, N483, N322);
or OR4 (N488, N486, N348, N268, N101);
xor XOR2 (N489, N482, N260);
nand NAND3 (N490, N489, N235, N239);
or OR3 (N491, N481, N211, N215);
xor XOR2 (N492, N487, N436);
and AND2 (N493, N490, N454);
or OR3 (N494, N492, N413, N45);
xor XOR2 (N495, N494, N447);
not NOT1 (N496, N479);
and AND2 (N497, N496, N66);
and AND3 (N498, N491, N209, N409);
not NOT1 (N499, N475);
not NOT1 (N500, N499);
not NOT1 (N501, N495);
not NOT1 (N502, N501);
not NOT1 (N503, N471);
nand NAND4 (N504, N485, N418, N28, N396);
nor NOR3 (N505, N498, N481, N339);
buf BUF1 (N506, N493);
nor NOR2 (N507, N500, N409);
and AND2 (N508, N497, N236);
and AND4 (N509, N469, N149, N158, N226);
xor XOR2 (N510, N488, N127);
and AND3 (N511, N507, N418, N213);
nand NAND2 (N512, N476, N414);
and AND2 (N513, N504, N296);
xor XOR2 (N514, N502, N113);
nand NAND2 (N515, N506, N167);
or OR4 (N516, N511, N435, N400, N193);
or OR3 (N517, N510, N94, N241);
buf BUF1 (N518, N512);
buf BUF1 (N519, N508);
and AND4 (N520, N514, N132, N253, N514);
nor NOR4 (N521, N517, N90, N303, N206);
or OR3 (N522, N518, N435, N521);
buf BUF1 (N523, N379);
and AND2 (N524, N503, N134);
buf BUF1 (N525, N524);
xor XOR2 (N526, N519, N12);
nand NAND4 (N527, N523, N506, N40, N322);
not NOT1 (N528, N513);
or OR4 (N529, N505, N233, N368, N432);
nand NAND2 (N530, N525, N161);
nor NOR4 (N531, N522, N270, N466, N525);
and AND4 (N532, N520, N382, N489, N301);
or OR4 (N533, N509, N146, N396, N463);
and AND3 (N534, N515, N348, N365);
nand NAND3 (N535, N534, N310, N343);
xor XOR2 (N536, N530, N353);
buf BUF1 (N537, N529);
not NOT1 (N538, N532);
and AND3 (N539, N531, N202, N342);
not NOT1 (N540, N536);
nand NAND4 (N541, N538, N466, N160, N367);
nor NOR2 (N542, N533, N23);
buf BUF1 (N543, N537);
buf BUF1 (N544, N542);
buf BUF1 (N545, N539);
and AND3 (N546, N527, N166, N187);
and AND3 (N547, N543, N239, N303);
nand NAND2 (N548, N544, N178);
not NOT1 (N549, N535);
nor NOR3 (N550, N546, N534, N529);
buf BUF1 (N551, N516);
not NOT1 (N552, N550);
nand NAND3 (N553, N545, N266, N358);
xor XOR2 (N554, N547, N247);
xor XOR2 (N555, N548, N392);
nand NAND4 (N556, N528, N157, N234, N128);
and AND3 (N557, N552, N86, N337);
not NOT1 (N558, N554);
nand NAND2 (N559, N553, N557);
nor NOR4 (N560, N112, N424, N387, N251);
and AND3 (N561, N559, N73, N133);
and AND4 (N562, N541, N126, N520, N188);
not NOT1 (N563, N560);
xor XOR2 (N564, N563, N208);
buf BUF1 (N565, N556);
xor XOR2 (N566, N564, N97);
nor NOR4 (N567, N561, N92, N120, N396);
xor XOR2 (N568, N565, N507);
and AND2 (N569, N568, N73);
not NOT1 (N570, N558);
not NOT1 (N571, N567);
or OR3 (N572, N549, N189, N210);
and AND4 (N573, N569, N36, N16, N245);
buf BUF1 (N574, N573);
xor XOR2 (N575, N566, N447);
not NOT1 (N576, N551);
xor XOR2 (N577, N555, N510);
nor NOR4 (N578, N571, N401, N245, N475);
or OR3 (N579, N576, N360, N315);
xor XOR2 (N580, N526, N472);
not NOT1 (N581, N574);
nand NAND4 (N582, N540, N20, N101, N581);
buf BUF1 (N583, N456);
or OR2 (N584, N578, N338);
xor XOR2 (N585, N570, N515);
or OR4 (N586, N582, N94, N183, N300);
buf BUF1 (N587, N580);
or OR3 (N588, N575, N555, N485);
and AND3 (N589, N586, N456, N146);
or OR3 (N590, N562, N298, N66);
nor NOR3 (N591, N589, N512, N403);
or OR2 (N592, N590, N365);
or OR3 (N593, N584, N323, N6);
nor NOR4 (N594, N588, N557, N410, N495);
buf BUF1 (N595, N583);
nand NAND2 (N596, N594, N417);
not NOT1 (N597, N585);
buf BUF1 (N598, N591);
or OR4 (N599, N596, N467, N335, N130);
or OR3 (N600, N599, N153, N163);
nor NOR4 (N601, N597, N460, N480, N487);
nor NOR3 (N602, N579, N64, N380);
xor XOR2 (N603, N600, N473);
nand NAND3 (N604, N577, N471, N487);
and AND4 (N605, N587, N168, N546, N532);
and AND4 (N606, N602, N92, N435, N107);
buf BUF1 (N607, N593);
nor NOR3 (N608, N595, N531, N256);
not NOT1 (N609, N572);
xor XOR2 (N610, N605, N96);
not NOT1 (N611, N606);
nor NOR4 (N612, N603, N293, N512, N195);
not NOT1 (N613, N608);
nor NOR3 (N614, N611, N556, N54);
buf BUF1 (N615, N601);
not NOT1 (N616, N598);
not NOT1 (N617, N610);
buf BUF1 (N618, N609);
nand NAND4 (N619, N613, N8, N176, N156);
xor XOR2 (N620, N614, N191);
xor XOR2 (N621, N620, N609);
and AND2 (N622, N616, N100);
and AND4 (N623, N622, N316, N337, N601);
not NOT1 (N624, N617);
not NOT1 (N625, N612);
nand NAND4 (N626, N615, N413, N502, N118);
buf BUF1 (N627, N625);
nor NOR4 (N628, N623, N245, N185, N468);
buf BUF1 (N629, N607);
buf BUF1 (N630, N626);
nor NOR3 (N631, N619, N138, N318);
not NOT1 (N632, N592);
not NOT1 (N633, N618);
xor XOR2 (N634, N631, N171);
not NOT1 (N635, N628);
nor NOR2 (N636, N632, N567);
and AND3 (N637, N636, N489, N232);
not NOT1 (N638, N637);
xor XOR2 (N639, N604, N369);
or OR4 (N640, N634, N543, N246, N199);
nand NAND4 (N641, N621, N585, N424, N640);
and AND2 (N642, N495, N529);
nand NAND4 (N643, N641, N111, N641, N561);
nor NOR2 (N644, N627, N230);
not NOT1 (N645, N629);
buf BUF1 (N646, N633);
not NOT1 (N647, N639);
xor XOR2 (N648, N645, N480);
and AND2 (N649, N630, N555);
xor XOR2 (N650, N624, N29);
nor NOR3 (N651, N644, N50, N13);
nor NOR3 (N652, N651, N318, N642);
and AND3 (N653, N366, N380, N169);
or OR2 (N654, N643, N217);
and AND4 (N655, N638, N426, N3, N96);
nand NAND2 (N656, N652, N632);
nor NOR3 (N657, N648, N129, N368);
buf BUF1 (N658, N656);
nor NOR2 (N659, N646, N433);
not NOT1 (N660, N649);
nor NOR2 (N661, N650, N18);
or OR3 (N662, N654, N253, N470);
and AND3 (N663, N658, N243, N372);
or OR3 (N664, N660, N517, N458);
or OR2 (N665, N664, N543);
nor NOR2 (N666, N653, N71);
nor NOR4 (N667, N635, N268, N239, N435);
not NOT1 (N668, N659);
or OR2 (N669, N668, N114);
nor NOR3 (N670, N662, N457, N582);
xor XOR2 (N671, N669, N612);
buf BUF1 (N672, N657);
nand NAND4 (N673, N665, N435, N625, N190);
buf BUF1 (N674, N663);
and AND2 (N675, N666, N338);
nand NAND3 (N676, N671, N670, N642);
buf BUF1 (N677, N636);
xor XOR2 (N678, N661, N143);
not NOT1 (N679, N667);
nor NOR2 (N680, N655, N402);
or OR4 (N681, N675, N174, N478, N27);
nand NAND2 (N682, N676, N292);
xor XOR2 (N683, N678, N288);
or OR3 (N684, N674, N162, N71);
xor XOR2 (N685, N683, N150);
xor XOR2 (N686, N672, N341);
nand NAND2 (N687, N681, N24);
xor XOR2 (N688, N686, N432);
nor NOR2 (N689, N688, N362);
or OR4 (N690, N673, N626, N30, N262);
and AND4 (N691, N679, N90, N372, N613);
not NOT1 (N692, N687);
buf BUF1 (N693, N691);
and AND2 (N694, N680, N207);
nor NOR2 (N695, N689, N102);
or OR4 (N696, N695, N452, N661, N640);
and AND3 (N697, N690, N541, N686);
or OR3 (N698, N685, N246, N486);
and AND4 (N699, N697, N397, N335, N209);
or OR2 (N700, N693, N170);
buf BUF1 (N701, N698);
buf BUF1 (N702, N677);
nand NAND3 (N703, N702, N184, N524);
nor NOR3 (N704, N696, N519, N559);
nand NAND4 (N705, N692, N416, N6, N220);
not NOT1 (N706, N684);
nand NAND4 (N707, N701, N691, N285, N478);
and AND3 (N708, N705, N214, N399);
nand NAND4 (N709, N704, N602, N67, N627);
buf BUF1 (N710, N703);
not NOT1 (N711, N694);
and AND4 (N712, N682, N471, N169, N139);
not NOT1 (N713, N700);
xor XOR2 (N714, N709, N353);
buf BUF1 (N715, N711);
nand NAND4 (N716, N708, N128, N376, N189);
nand NAND3 (N717, N714, N370, N103);
buf BUF1 (N718, N707);
nand NAND4 (N719, N713, N99, N507, N486);
and AND2 (N720, N699, N709);
or OR4 (N721, N720, N279, N50, N354);
nor NOR3 (N722, N715, N4, N433);
and AND3 (N723, N710, N687, N415);
or OR2 (N724, N719, N664);
nor NOR4 (N725, N647, N661, N251, N24);
nand NAND4 (N726, N718, N441, N332, N163);
nor NOR2 (N727, N706, N444);
xor XOR2 (N728, N717, N615);
buf BUF1 (N729, N725);
or OR4 (N730, N716, N227, N518, N212);
xor XOR2 (N731, N726, N311);
not NOT1 (N732, N727);
xor XOR2 (N733, N728, N105);
and AND4 (N734, N723, N612, N228, N38);
buf BUF1 (N735, N712);
or OR4 (N736, N729, N624, N102, N304);
buf BUF1 (N737, N735);
xor XOR2 (N738, N736, N682);
not NOT1 (N739, N737);
and AND4 (N740, N730, N437, N285, N102);
xor XOR2 (N741, N740, N677);
nand NAND3 (N742, N724, N88, N119);
or OR3 (N743, N734, N318, N255);
nand NAND3 (N744, N739, N734, N137);
or OR2 (N745, N722, N34);
not NOT1 (N746, N733);
not NOT1 (N747, N742);
nand NAND2 (N748, N744, N531);
not NOT1 (N749, N721);
xor XOR2 (N750, N741, N150);
or OR4 (N751, N731, N316, N26, N256);
nor NOR4 (N752, N749, N224, N172, N664);
and AND4 (N753, N747, N246, N427, N187);
nand NAND3 (N754, N751, N107, N600);
or OR4 (N755, N748, N676, N593, N196);
nor NOR4 (N756, N743, N520, N96, N361);
or OR2 (N757, N732, N16);
buf BUF1 (N758, N757);
nor NOR2 (N759, N753, N660);
buf BUF1 (N760, N746);
buf BUF1 (N761, N750);
and AND4 (N762, N758, N654, N371, N719);
nor NOR3 (N763, N755, N84, N456);
and AND4 (N764, N761, N268, N161, N583);
nand NAND4 (N765, N738, N446, N330, N173);
or OR4 (N766, N760, N372, N452, N502);
and AND4 (N767, N759, N405, N495, N464);
not NOT1 (N768, N752);
nor NOR4 (N769, N768, N642, N343, N523);
buf BUF1 (N770, N765);
buf BUF1 (N771, N764);
nand NAND4 (N772, N745, N373, N296, N161);
xor XOR2 (N773, N772, N342);
not NOT1 (N774, N766);
nand NAND2 (N775, N756, N57);
and AND2 (N776, N771, N110);
not NOT1 (N777, N770);
nor NOR2 (N778, N754, N585);
xor XOR2 (N779, N774, N323);
nand NAND4 (N780, N763, N461, N622, N433);
and AND4 (N781, N769, N737, N704, N750);
or OR4 (N782, N776, N332, N278, N81);
xor XOR2 (N783, N775, N75);
buf BUF1 (N784, N780);
or OR3 (N785, N783, N721, N375);
and AND3 (N786, N778, N743, N178);
nor NOR4 (N787, N781, N69, N89, N499);
or OR4 (N788, N785, N532, N206, N109);
not NOT1 (N789, N762);
buf BUF1 (N790, N789);
nand NAND2 (N791, N788, N282);
buf BUF1 (N792, N784);
not NOT1 (N793, N787);
or OR2 (N794, N779, N117);
or OR3 (N795, N793, N246, N235);
buf BUF1 (N796, N777);
nor NOR4 (N797, N786, N621, N771, N45);
nor NOR2 (N798, N790, N20);
nor NOR3 (N799, N794, N241, N533);
and AND4 (N800, N792, N750, N463, N576);
or OR3 (N801, N767, N772, N384);
nand NAND2 (N802, N798, N733);
nor NOR3 (N803, N801, N701, N308);
nand NAND3 (N804, N773, N288, N634);
buf BUF1 (N805, N804);
nor NOR2 (N806, N796, N443);
nand NAND4 (N807, N805, N399, N765, N624);
xor XOR2 (N808, N799, N318);
and AND3 (N809, N795, N118, N682);
and AND3 (N810, N791, N568, N301);
or OR3 (N811, N807, N179, N714);
nor NOR2 (N812, N810, N464);
and AND3 (N813, N800, N781, N691);
buf BUF1 (N814, N806);
nor NOR3 (N815, N797, N724, N140);
nand NAND3 (N816, N815, N291, N258);
or OR2 (N817, N813, N36);
or OR2 (N818, N809, N459);
nor NOR4 (N819, N811, N124, N157, N610);
not NOT1 (N820, N816);
or OR3 (N821, N818, N116, N345);
not NOT1 (N822, N820);
and AND2 (N823, N803, N775);
and AND4 (N824, N817, N183, N508, N320);
not NOT1 (N825, N814);
not NOT1 (N826, N808);
xor XOR2 (N827, N824, N783);
and AND2 (N828, N827, N165);
buf BUF1 (N829, N802);
or OR2 (N830, N826, N269);
or OR4 (N831, N812, N342, N288, N206);
nand NAND2 (N832, N823, N657);
or OR3 (N833, N782, N804, N811);
or OR3 (N834, N829, N196, N246);
nor NOR2 (N835, N831, N609);
not NOT1 (N836, N822);
or OR2 (N837, N821, N530);
or OR2 (N838, N837, N30);
xor XOR2 (N839, N819, N737);
or OR4 (N840, N836, N471, N366, N303);
or OR3 (N841, N838, N211, N124);
nor NOR4 (N842, N828, N349, N188, N297);
xor XOR2 (N843, N840, N59);
buf BUF1 (N844, N839);
buf BUF1 (N845, N830);
or OR4 (N846, N833, N119, N728, N409);
xor XOR2 (N847, N843, N746);
buf BUF1 (N848, N845);
and AND2 (N849, N847, N571);
or OR4 (N850, N848, N577, N399, N789);
and AND4 (N851, N849, N379, N503, N651);
not NOT1 (N852, N825);
xor XOR2 (N853, N841, N367);
or OR4 (N854, N851, N799, N108, N1);
nor NOR4 (N855, N842, N102, N783, N664);
buf BUF1 (N856, N853);
not NOT1 (N857, N854);
nand NAND4 (N858, N855, N325, N457, N147);
xor XOR2 (N859, N852, N749);
nor NOR3 (N860, N858, N764, N586);
and AND3 (N861, N856, N614, N70);
nor NOR4 (N862, N859, N291, N59, N384);
nand NAND3 (N863, N835, N509, N755);
nor NOR2 (N864, N857, N487);
and AND4 (N865, N850, N684, N189, N403);
xor XOR2 (N866, N844, N493);
nand NAND3 (N867, N834, N194, N642);
xor XOR2 (N868, N866, N261);
or OR3 (N869, N865, N859, N807);
buf BUF1 (N870, N863);
nor NOR3 (N871, N870, N621, N741);
xor XOR2 (N872, N867, N836);
xor XOR2 (N873, N832, N456);
or OR3 (N874, N872, N756, N386);
buf BUF1 (N875, N864);
buf BUF1 (N876, N846);
or OR2 (N877, N875, N58);
nand NAND3 (N878, N869, N230, N373);
nor NOR3 (N879, N862, N390, N494);
nand NAND3 (N880, N877, N326, N623);
nand NAND4 (N881, N880, N39, N843, N765);
or OR4 (N882, N878, N843, N872, N389);
xor XOR2 (N883, N882, N376);
or OR4 (N884, N871, N310, N377, N134);
and AND2 (N885, N881, N298);
nand NAND3 (N886, N868, N599, N123);
not NOT1 (N887, N884);
or OR3 (N888, N879, N522, N551);
nand NAND2 (N889, N888, N187);
buf BUF1 (N890, N887);
buf BUF1 (N891, N876);
nor NOR4 (N892, N861, N674, N288, N416);
xor XOR2 (N893, N885, N826);
nor NOR3 (N894, N892, N2, N73);
xor XOR2 (N895, N886, N652);
and AND4 (N896, N860, N375, N399, N212);
nand NAND2 (N897, N873, N197);
nor NOR3 (N898, N883, N673, N262);
nor NOR3 (N899, N891, N304, N775);
xor XOR2 (N900, N893, N380);
or OR2 (N901, N896, N798);
nand NAND3 (N902, N889, N205, N886);
not NOT1 (N903, N894);
xor XOR2 (N904, N900, N716);
nand NAND3 (N905, N874, N512, N252);
xor XOR2 (N906, N904, N475);
not NOT1 (N907, N890);
xor XOR2 (N908, N902, N468);
buf BUF1 (N909, N895);
buf BUF1 (N910, N897);
and AND2 (N911, N909, N767);
and AND3 (N912, N905, N621, N113);
nor NOR4 (N913, N906, N865, N371, N777);
nor NOR3 (N914, N913, N260, N430);
or OR4 (N915, N899, N82, N91, N574);
and AND3 (N916, N898, N469, N645);
or OR2 (N917, N914, N464);
buf BUF1 (N918, N903);
nand NAND4 (N919, N910, N84, N174, N210);
buf BUF1 (N920, N916);
and AND3 (N921, N917, N879, N747);
nand NAND4 (N922, N912, N441, N857, N21);
nand NAND4 (N923, N907, N457, N140, N32);
not NOT1 (N924, N923);
or OR2 (N925, N908, N275);
nor NOR2 (N926, N918, N237);
and AND4 (N927, N924, N561, N20, N329);
buf BUF1 (N928, N915);
nand NAND2 (N929, N911, N690);
buf BUF1 (N930, N901);
and AND4 (N931, N927, N564, N909, N577);
xor XOR2 (N932, N929, N585);
and AND2 (N933, N925, N804);
nor NOR3 (N934, N926, N493, N612);
not NOT1 (N935, N919);
nand NAND4 (N936, N930, N641, N109, N448);
xor XOR2 (N937, N936, N438);
xor XOR2 (N938, N922, N835);
or OR4 (N939, N937, N649, N478, N705);
and AND4 (N940, N935, N435, N444, N134);
buf BUF1 (N941, N931);
buf BUF1 (N942, N921);
xor XOR2 (N943, N920, N792);
and AND3 (N944, N939, N114, N379);
xor XOR2 (N945, N932, N603);
nor NOR2 (N946, N944, N858);
xor XOR2 (N947, N946, N687);
not NOT1 (N948, N947);
xor XOR2 (N949, N948, N63);
nand NAND2 (N950, N934, N181);
nand NAND3 (N951, N933, N99, N425);
nand NAND2 (N952, N950, N949);
nor NOR4 (N953, N191, N375, N665, N320);
buf BUF1 (N954, N938);
xor XOR2 (N955, N945, N804);
or OR2 (N956, N954, N807);
xor XOR2 (N957, N941, N657);
nor NOR2 (N958, N953, N884);
nand NAND4 (N959, N958, N900, N191, N185);
buf BUF1 (N960, N940);
buf BUF1 (N961, N955);
or OR4 (N962, N956, N444, N200, N846);
and AND4 (N963, N943, N157, N657, N837);
not NOT1 (N964, N952);
buf BUF1 (N965, N962);
nor NOR2 (N966, N965, N327);
buf BUF1 (N967, N964);
nor NOR3 (N968, N959, N439, N490);
nand NAND2 (N969, N942, N841);
xor XOR2 (N970, N951, N803);
and AND3 (N971, N928, N305, N659);
not NOT1 (N972, N970);
xor XOR2 (N973, N966, N609);
nand NAND4 (N974, N971, N739, N551, N599);
nor NOR4 (N975, N957, N570, N195, N14);
or OR3 (N976, N973, N224, N543);
buf BUF1 (N977, N960);
buf BUF1 (N978, N972);
not NOT1 (N979, N978);
xor XOR2 (N980, N967, N503);
xor XOR2 (N981, N963, N105);
and AND3 (N982, N969, N516, N819);
nand NAND2 (N983, N979, N975);
nand NAND4 (N984, N163, N134, N779, N396);
xor XOR2 (N985, N977, N742);
not NOT1 (N986, N985);
not NOT1 (N987, N974);
nand NAND2 (N988, N984, N167);
xor XOR2 (N989, N982, N322);
nand NAND2 (N990, N980, N21);
nand NAND4 (N991, N961, N333, N381, N727);
nor NOR2 (N992, N991, N357);
nand NAND4 (N993, N976, N523, N954, N51);
or OR4 (N994, N981, N125, N325, N273);
buf BUF1 (N995, N989);
not NOT1 (N996, N993);
and AND2 (N997, N995, N982);
and AND3 (N998, N992, N232, N800);
buf BUF1 (N999, N998);
and AND4 (N1000, N988, N571, N557, N498);
xor XOR2 (N1001, N1000, N728);
xor XOR2 (N1002, N996, N938);
not NOT1 (N1003, N1001);
buf BUF1 (N1004, N1003);
and AND3 (N1005, N1002, N749, N545);
nand NAND4 (N1006, N999, N88, N682, N22);
nor NOR4 (N1007, N1005, N558, N709, N690);
not NOT1 (N1008, N983);
nand NAND4 (N1009, N990, N595, N152, N786);
xor XOR2 (N1010, N1007, N212);
buf BUF1 (N1011, N987);
xor XOR2 (N1012, N1008, N816);
or OR3 (N1013, N1009, N65, N796);
not NOT1 (N1014, N994);
xor XOR2 (N1015, N1006, N34);
and AND4 (N1016, N1015, N342, N22, N903);
xor XOR2 (N1017, N1004, N326);
or OR3 (N1018, N1011, N326, N717);
buf BUF1 (N1019, N1016);
nand NAND3 (N1020, N1012, N423, N668);
xor XOR2 (N1021, N1014, N707);
not NOT1 (N1022, N1020);
nand NAND3 (N1023, N1017, N902, N938);
and AND2 (N1024, N1010, N529);
nor NOR3 (N1025, N1019, N871, N629);
xor XOR2 (N1026, N1023, N851);
nand NAND2 (N1027, N1013, N634);
and AND3 (N1028, N968, N368, N1018);
or OR4 (N1029, N84, N702, N44, N1028);
or OR4 (N1030, N15, N523, N49, N221);
nor NOR3 (N1031, N997, N271, N694);
xor XOR2 (N1032, N1027, N1019);
nor NOR2 (N1033, N1029, N582);
and AND4 (N1034, N986, N546, N371, N93);
or OR4 (N1035, N1031, N992, N1033, N857);
not NOT1 (N1036, N71);
and AND2 (N1037, N1035, N584);
xor XOR2 (N1038, N1025, N227);
nor NOR4 (N1039, N1032, N40, N634, N107);
or OR4 (N1040, N1024, N975, N1005, N784);
xor XOR2 (N1041, N1030, N140);
xor XOR2 (N1042, N1036, N825);
not NOT1 (N1043, N1042);
buf BUF1 (N1044, N1040);
or OR3 (N1045, N1044, N580, N271);
and AND2 (N1046, N1039, N573);
or OR3 (N1047, N1021, N799, N940);
not NOT1 (N1048, N1046);
or OR2 (N1049, N1047, N308);
nor NOR4 (N1050, N1026, N671, N614, N309);
not NOT1 (N1051, N1041);
or OR2 (N1052, N1038, N433);
or OR3 (N1053, N1045, N595, N374);
not NOT1 (N1054, N1051);
or OR4 (N1055, N1034, N711, N859, N968);
not NOT1 (N1056, N1022);
and AND4 (N1057, N1048, N502, N702, N235);
nor NOR3 (N1058, N1037, N561, N149);
or OR3 (N1059, N1050, N921, N268);
nand NAND2 (N1060, N1056, N939);
nor NOR2 (N1061, N1055, N112);
nand NAND4 (N1062, N1059, N155, N846, N651);
nand NAND4 (N1063, N1061, N845, N305, N814);
buf BUF1 (N1064, N1049);
nor NOR3 (N1065, N1058, N453, N27);
nand NAND3 (N1066, N1053, N1040, N998);
nor NOR4 (N1067, N1054, N1033, N261, N24);
xor XOR2 (N1068, N1066, N299);
not NOT1 (N1069, N1057);
xor XOR2 (N1070, N1043, N970);
nor NOR2 (N1071, N1065, N251);
buf BUF1 (N1072, N1071);
nor NOR4 (N1073, N1068, N20, N106, N908);
and AND4 (N1074, N1060, N977, N986, N775);
xor XOR2 (N1075, N1072, N847);
nand NAND3 (N1076, N1069, N465, N473);
buf BUF1 (N1077, N1052);
buf BUF1 (N1078, N1062);
nand NAND3 (N1079, N1070, N523, N306);
or OR4 (N1080, N1078, N402, N947, N602);
nor NOR4 (N1081, N1080, N403, N830, N965);
xor XOR2 (N1082, N1074, N1012);
xor XOR2 (N1083, N1064, N932);
not NOT1 (N1084, N1077);
not NOT1 (N1085, N1076);
xor XOR2 (N1086, N1073, N636);
nor NOR4 (N1087, N1082, N908, N1070, N309);
nand NAND3 (N1088, N1063, N1074, N296);
or OR4 (N1089, N1075, N56, N745, N126);
buf BUF1 (N1090, N1081);
nand NAND4 (N1091, N1083, N989, N343, N1045);
buf BUF1 (N1092, N1084);
and AND4 (N1093, N1088, N238, N218, N374);
xor XOR2 (N1094, N1090, N734);
nor NOR2 (N1095, N1093, N1081);
nor NOR2 (N1096, N1092, N236);
nor NOR4 (N1097, N1079, N656, N402, N601);
and AND2 (N1098, N1087, N620);
nand NAND4 (N1099, N1094, N632, N742, N291);
xor XOR2 (N1100, N1097, N901);
nand NAND2 (N1101, N1091, N765);
buf BUF1 (N1102, N1099);
or OR3 (N1103, N1100, N880, N843);
or OR3 (N1104, N1103, N383, N4);
buf BUF1 (N1105, N1102);
nand NAND2 (N1106, N1104, N885);
and AND3 (N1107, N1096, N117, N1101);
or OR4 (N1108, N781, N117, N510, N536);
not NOT1 (N1109, N1085);
xor XOR2 (N1110, N1086, N471);
and AND3 (N1111, N1105, N743, N976);
buf BUF1 (N1112, N1089);
nand NAND4 (N1113, N1107, N1018, N538, N673);
not NOT1 (N1114, N1098);
not NOT1 (N1115, N1111);
nand NAND2 (N1116, N1108, N502);
buf BUF1 (N1117, N1067);
nor NOR4 (N1118, N1112, N890, N195, N1087);
nand NAND3 (N1119, N1095, N86, N32);
nand NAND4 (N1120, N1110, N120, N989, N470);
and AND3 (N1121, N1117, N693, N472);
buf BUF1 (N1122, N1115);
nor NOR3 (N1123, N1120, N1080, N405);
nand NAND2 (N1124, N1119, N1031);
or OR3 (N1125, N1114, N1065, N334);
and AND3 (N1126, N1106, N744, N343);
or OR2 (N1127, N1113, N490);
and AND2 (N1128, N1122, N1055);
not NOT1 (N1129, N1121);
nor NOR4 (N1130, N1124, N1048, N638, N449);
or OR3 (N1131, N1123, N650, N218);
or OR2 (N1132, N1130, N409);
nor NOR4 (N1133, N1127, N1072, N79, N650);
and AND3 (N1134, N1131, N528, N455);
buf BUF1 (N1135, N1125);
nand NAND4 (N1136, N1126, N122, N674, N720);
nor NOR2 (N1137, N1134, N613);
and AND2 (N1138, N1118, N742);
xor XOR2 (N1139, N1138, N991);
xor XOR2 (N1140, N1109, N359);
nor NOR3 (N1141, N1135, N30, N350);
nor NOR3 (N1142, N1136, N656, N160);
buf BUF1 (N1143, N1139);
buf BUF1 (N1144, N1142);
not NOT1 (N1145, N1132);
xor XOR2 (N1146, N1143, N89);
not NOT1 (N1147, N1128);
nor NOR3 (N1148, N1137, N1138, N231);
nor NOR4 (N1149, N1148, N857, N334, N457);
nor NOR4 (N1150, N1145, N144, N116, N282);
buf BUF1 (N1151, N1129);
and AND3 (N1152, N1151, N1093, N638);
not NOT1 (N1153, N1150);
buf BUF1 (N1154, N1152);
and AND3 (N1155, N1141, N929, N307);
or OR4 (N1156, N1146, N334, N719, N891);
and AND3 (N1157, N1149, N888, N998);
nand NAND4 (N1158, N1133, N933, N787, N559);
not NOT1 (N1159, N1157);
buf BUF1 (N1160, N1154);
not NOT1 (N1161, N1147);
nand NAND4 (N1162, N1161, N481, N630, N394);
buf BUF1 (N1163, N1156);
buf BUF1 (N1164, N1160);
nor NOR3 (N1165, N1116, N448, N368);
buf BUF1 (N1166, N1163);
buf BUF1 (N1167, N1165);
buf BUF1 (N1168, N1155);
xor XOR2 (N1169, N1159, N1007);
and AND4 (N1170, N1162, N680, N154, N817);
xor XOR2 (N1171, N1167, N173);
buf BUF1 (N1172, N1140);
or OR2 (N1173, N1170, N73);
or OR2 (N1174, N1153, N1036);
not NOT1 (N1175, N1144);
buf BUF1 (N1176, N1174);
or OR4 (N1177, N1175, N1170, N194, N684);
or OR2 (N1178, N1173, N1010);
buf BUF1 (N1179, N1168);
or OR3 (N1180, N1166, N772, N627);
or OR3 (N1181, N1178, N358, N999);
not NOT1 (N1182, N1164);
not NOT1 (N1183, N1176);
nor NOR3 (N1184, N1171, N1014, N118);
or OR2 (N1185, N1158, N863);
nor NOR2 (N1186, N1177, N366);
not NOT1 (N1187, N1183);
not NOT1 (N1188, N1185);
and AND4 (N1189, N1172, N676, N639, N482);
or OR3 (N1190, N1184, N715, N1181);
and AND4 (N1191, N1028, N124, N127, N753);
buf BUF1 (N1192, N1169);
xor XOR2 (N1193, N1191, N1030);
not NOT1 (N1194, N1193);
nor NOR3 (N1195, N1188, N510, N455);
or OR4 (N1196, N1180, N406, N687, N1030);
and AND4 (N1197, N1195, N627, N1151, N1024);
nor NOR4 (N1198, N1189, N556, N764, N257);
and AND3 (N1199, N1186, N1123, N151);
and AND2 (N1200, N1182, N392);
nor NOR2 (N1201, N1194, N886);
or OR2 (N1202, N1201, N351);
nor NOR4 (N1203, N1190, N978, N29, N500);
buf BUF1 (N1204, N1179);
buf BUF1 (N1205, N1199);
not NOT1 (N1206, N1196);
xor XOR2 (N1207, N1200, N834);
nand NAND3 (N1208, N1204, N665, N916);
buf BUF1 (N1209, N1207);
nand NAND4 (N1210, N1187, N507, N1013, N255);
or OR2 (N1211, N1206, N359);
nand NAND4 (N1212, N1211, N940, N425, N507);
and AND2 (N1213, N1210, N833);
and AND4 (N1214, N1208, N844, N1117, N445);
xor XOR2 (N1215, N1198, N244);
not NOT1 (N1216, N1209);
not NOT1 (N1217, N1214);
nand NAND3 (N1218, N1205, N217, N984);
nand NAND2 (N1219, N1203, N613);
and AND4 (N1220, N1197, N460, N462, N230);
and AND4 (N1221, N1216, N680, N21, N976);
buf BUF1 (N1222, N1221);
not NOT1 (N1223, N1219);
nand NAND2 (N1224, N1223, N664);
nand NAND2 (N1225, N1224, N49);
xor XOR2 (N1226, N1213, N827);
xor XOR2 (N1227, N1217, N1154);
xor XOR2 (N1228, N1225, N295);
buf BUF1 (N1229, N1215);
nand NAND4 (N1230, N1226, N972, N1109, N888);
or OR4 (N1231, N1220, N754, N162, N1085);
and AND4 (N1232, N1222, N739, N558, N316);
nor NOR4 (N1233, N1231, N118, N1198, N728);
buf BUF1 (N1234, N1192);
nor NOR4 (N1235, N1218, N728, N775, N283);
or OR2 (N1236, N1227, N228);
xor XOR2 (N1237, N1229, N335);
nand NAND2 (N1238, N1228, N1052);
xor XOR2 (N1239, N1236, N1048);
nor NOR3 (N1240, N1233, N514, N1107);
nand NAND4 (N1241, N1240, N393, N554, N1167);
or OR2 (N1242, N1237, N670);
buf BUF1 (N1243, N1241);
xor XOR2 (N1244, N1202, N1236);
or OR2 (N1245, N1234, N1212);
and AND2 (N1246, N969, N1003);
not NOT1 (N1247, N1243);
xor XOR2 (N1248, N1238, N781);
nand NAND4 (N1249, N1232, N747, N90, N1097);
nand NAND2 (N1250, N1230, N392);
nand NAND4 (N1251, N1247, N423, N686, N1059);
nor NOR4 (N1252, N1249, N36, N611, N156);
not NOT1 (N1253, N1248);
not NOT1 (N1254, N1253);
or OR2 (N1255, N1250, N410);
not NOT1 (N1256, N1245);
buf BUF1 (N1257, N1235);
not NOT1 (N1258, N1246);
not NOT1 (N1259, N1252);
buf BUF1 (N1260, N1255);
and AND4 (N1261, N1258, N581, N639, N586);
xor XOR2 (N1262, N1242, N233);
and AND3 (N1263, N1262, N1167, N955);
not NOT1 (N1264, N1259);
or OR3 (N1265, N1251, N1155, N85);
or OR4 (N1266, N1264, N1098, N187, N764);
xor XOR2 (N1267, N1263, N346);
nor NOR2 (N1268, N1260, N624);
and AND4 (N1269, N1244, N1153, N749, N1225);
not NOT1 (N1270, N1256);
nand NAND4 (N1271, N1268, N723, N746, N376);
xor XOR2 (N1272, N1254, N377);
and AND4 (N1273, N1261, N503, N639, N1043);
xor XOR2 (N1274, N1269, N49);
buf BUF1 (N1275, N1274);
or OR3 (N1276, N1271, N1141, N920);
not NOT1 (N1277, N1267);
nand NAND2 (N1278, N1266, N1158);
buf BUF1 (N1279, N1272);
xor XOR2 (N1280, N1257, N585);
nand NAND4 (N1281, N1280, N102, N782, N779);
nand NAND4 (N1282, N1239, N720, N325, N31);
nand NAND3 (N1283, N1281, N778, N979);
not NOT1 (N1284, N1275);
nand NAND3 (N1285, N1276, N1148, N1055);
nand NAND2 (N1286, N1273, N699);
not NOT1 (N1287, N1282);
or OR3 (N1288, N1283, N1073, N374);
nor NOR3 (N1289, N1287, N161, N811);
nor NOR4 (N1290, N1270, N23, N562, N526);
nand NAND3 (N1291, N1288, N533, N773);
or OR2 (N1292, N1290, N1110);
buf BUF1 (N1293, N1285);
xor XOR2 (N1294, N1293, N228);
xor XOR2 (N1295, N1286, N664);
nand NAND2 (N1296, N1294, N537);
nor NOR4 (N1297, N1279, N752, N299, N763);
or OR2 (N1298, N1292, N1218);
or OR3 (N1299, N1284, N310, N1013);
and AND4 (N1300, N1296, N192, N542, N659);
and AND3 (N1301, N1295, N544, N1127);
nand NAND4 (N1302, N1300, N219, N873, N1231);
or OR3 (N1303, N1277, N296, N470);
and AND4 (N1304, N1303, N494, N72, N559);
nor NOR3 (N1305, N1278, N945, N34);
not NOT1 (N1306, N1299);
buf BUF1 (N1307, N1302);
buf BUF1 (N1308, N1265);
or OR2 (N1309, N1304, N321);
nor NOR2 (N1310, N1309, N635);
not NOT1 (N1311, N1291);
nor NOR2 (N1312, N1298, N1258);
not NOT1 (N1313, N1307);
nor NOR3 (N1314, N1312, N764, N477);
xor XOR2 (N1315, N1305, N562);
and AND2 (N1316, N1310, N508);
and AND2 (N1317, N1313, N895);
nor NOR3 (N1318, N1301, N455, N1057);
and AND3 (N1319, N1314, N848, N21);
nand NAND2 (N1320, N1289, N256);
xor XOR2 (N1321, N1311, N49);
and AND3 (N1322, N1297, N734, N1137);
nand NAND4 (N1323, N1308, N383, N127, N1180);
nand NAND4 (N1324, N1319, N1315, N961, N229);
nor NOR4 (N1325, N251, N383, N739, N838);
nor NOR4 (N1326, N1306, N970, N397, N273);
and AND2 (N1327, N1316, N381);
nand NAND3 (N1328, N1320, N713, N112);
and AND2 (N1329, N1326, N280);
or OR2 (N1330, N1329, N587);
xor XOR2 (N1331, N1328, N860);
xor XOR2 (N1332, N1331, N961);
xor XOR2 (N1333, N1327, N170);
and AND4 (N1334, N1332, N770, N1083, N297);
not NOT1 (N1335, N1317);
or OR2 (N1336, N1334, N57);
xor XOR2 (N1337, N1318, N807);
nand NAND3 (N1338, N1321, N1087, N1003);
not NOT1 (N1339, N1323);
buf BUF1 (N1340, N1336);
and AND2 (N1341, N1333, N274);
or OR2 (N1342, N1330, N126);
xor XOR2 (N1343, N1324, N520);
buf BUF1 (N1344, N1337);
xor XOR2 (N1345, N1342, N683);
nor NOR3 (N1346, N1345, N625, N620);
xor XOR2 (N1347, N1325, N831);
nand NAND4 (N1348, N1340, N624, N78, N882);
and AND2 (N1349, N1341, N780);
and AND3 (N1350, N1347, N65, N670);
xor XOR2 (N1351, N1346, N529);
and AND3 (N1352, N1344, N107, N1114);
buf BUF1 (N1353, N1338);
not NOT1 (N1354, N1351);
nor NOR2 (N1355, N1352, N901);
nand NAND4 (N1356, N1353, N1179, N356, N541);
nor NOR2 (N1357, N1322, N611);
not NOT1 (N1358, N1355);
nand NAND2 (N1359, N1349, N107);
nand NAND3 (N1360, N1335, N863, N659);
or OR2 (N1361, N1357, N255);
nand NAND3 (N1362, N1350, N498, N7);
xor XOR2 (N1363, N1339, N654);
and AND4 (N1364, N1359, N884, N349, N820);
nand NAND2 (N1365, N1358, N35);
or OR3 (N1366, N1356, N886, N519);
not NOT1 (N1367, N1363);
nor NOR4 (N1368, N1354, N1315, N315, N633);
or OR2 (N1369, N1366, N394);
xor XOR2 (N1370, N1365, N984);
not NOT1 (N1371, N1360);
and AND3 (N1372, N1370, N230, N403);
and AND4 (N1373, N1362, N605, N1315, N116);
xor XOR2 (N1374, N1373, N1220);
not NOT1 (N1375, N1371);
xor XOR2 (N1376, N1361, N995);
buf BUF1 (N1377, N1367);
nor NOR4 (N1378, N1376, N304, N392, N859);
not NOT1 (N1379, N1368);
or OR3 (N1380, N1364, N285, N162);
nand NAND4 (N1381, N1348, N427, N693, N875);
nor NOR4 (N1382, N1343, N797, N1109, N585);
not NOT1 (N1383, N1381);
nand NAND3 (N1384, N1380, N813, N705);
or OR2 (N1385, N1372, N108);
nor NOR2 (N1386, N1379, N391);
not NOT1 (N1387, N1374);
buf BUF1 (N1388, N1377);
buf BUF1 (N1389, N1387);
buf BUF1 (N1390, N1386);
and AND2 (N1391, N1383, N607);
xor XOR2 (N1392, N1369, N459);
buf BUF1 (N1393, N1389);
nor NOR3 (N1394, N1385, N628, N1376);
xor XOR2 (N1395, N1375, N462);
or OR3 (N1396, N1394, N504, N1102);
and AND4 (N1397, N1393, N403, N778, N1345);
not NOT1 (N1398, N1382);
and AND2 (N1399, N1388, N222);
not NOT1 (N1400, N1398);
not NOT1 (N1401, N1399);
or OR4 (N1402, N1396, N1053, N925, N1182);
buf BUF1 (N1403, N1400);
xor XOR2 (N1404, N1397, N1129);
and AND4 (N1405, N1401, N983, N281, N371);
xor XOR2 (N1406, N1395, N93);
xor XOR2 (N1407, N1402, N801);
or OR2 (N1408, N1403, N1254);
xor XOR2 (N1409, N1405, N15);
and AND2 (N1410, N1391, N774);
and AND3 (N1411, N1390, N1064, N364);
or OR2 (N1412, N1406, N299);
xor XOR2 (N1413, N1409, N1359);
or OR3 (N1414, N1411, N1274, N1298);
nor NOR4 (N1415, N1412, N606, N467, N298);
xor XOR2 (N1416, N1392, N26);
or OR4 (N1417, N1408, N1105, N771, N957);
or OR3 (N1418, N1413, N1037, N220);
nor NOR3 (N1419, N1384, N605, N632);
xor XOR2 (N1420, N1410, N77);
nand NAND2 (N1421, N1404, N607);
xor XOR2 (N1422, N1420, N1399);
xor XOR2 (N1423, N1418, N58);
not NOT1 (N1424, N1378);
not NOT1 (N1425, N1424);
buf BUF1 (N1426, N1423);
or OR2 (N1427, N1407, N94);
nand NAND3 (N1428, N1425, N813, N805);
not NOT1 (N1429, N1422);
nand NAND2 (N1430, N1426, N382);
and AND4 (N1431, N1414, N1068, N1229, N743);
not NOT1 (N1432, N1419);
buf BUF1 (N1433, N1416);
nand NAND2 (N1434, N1415, N579);
and AND3 (N1435, N1430, N406, N423);
nand NAND4 (N1436, N1432, N68, N654, N1247);
nor NOR3 (N1437, N1431, N995, N439);
xor XOR2 (N1438, N1429, N1293);
or OR4 (N1439, N1435, N1211, N524, N1398);
nand NAND3 (N1440, N1433, N1237, N1360);
nor NOR2 (N1441, N1438, N712);
not NOT1 (N1442, N1428);
xor XOR2 (N1443, N1437, N626);
nand NAND3 (N1444, N1441, N82, N1247);
nand NAND2 (N1445, N1421, N448);
or OR2 (N1446, N1434, N1279);
nand NAND2 (N1447, N1427, N1081);
buf BUF1 (N1448, N1447);
or OR2 (N1449, N1448, N58);
nand NAND3 (N1450, N1440, N144, N446);
not NOT1 (N1451, N1442);
nor NOR3 (N1452, N1439, N380, N702);
not NOT1 (N1453, N1436);
not NOT1 (N1454, N1443);
and AND3 (N1455, N1445, N1292, N366);
and AND4 (N1456, N1455, N1131, N1430, N614);
xor XOR2 (N1457, N1452, N1129);
xor XOR2 (N1458, N1454, N1107);
nor NOR3 (N1459, N1451, N267, N524);
not NOT1 (N1460, N1444);
not NOT1 (N1461, N1446);
nand NAND3 (N1462, N1450, N848, N655);
nand NAND2 (N1463, N1458, N1029);
buf BUF1 (N1464, N1459);
xor XOR2 (N1465, N1463, N183);
or OR3 (N1466, N1449, N1463, N41);
nand NAND2 (N1467, N1460, N1249);
not NOT1 (N1468, N1464);
not NOT1 (N1469, N1465);
and AND2 (N1470, N1466, N247);
or OR4 (N1471, N1417, N1251, N977, N1417);
nor NOR2 (N1472, N1462, N1239);
buf BUF1 (N1473, N1457);
nand NAND2 (N1474, N1468, N577);
or OR3 (N1475, N1473, N1083, N134);
nand NAND4 (N1476, N1461, N30, N399, N317);
or OR2 (N1477, N1476, N1203);
and AND3 (N1478, N1474, N770, N12);
nor NOR3 (N1479, N1478, N1112, N781);
or OR4 (N1480, N1472, N1145, N419, N849);
or OR4 (N1481, N1453, N1031, N1108, N272);
nand NAND3 (N1482, N1479, N507, N499);
and AND2 (N1483, N1470, N495);
nand NAND3 (N1484, N1483, N696, N890);
nand NAND2 (N1485, N1475, N111);
nand NAND2 (N1486, N1480, N574);
xor XOR2 (N1487, N1485, N408);
xor XOR2 (N1488, N1477, N775);
buf BUF1 (N1489, N1471);
nor NOR3 (N1490, N1467, N270, N485);
or OR3 (N1491, N1490, N1240, N1217);
not NOT1 (N1492, N1484);
or OR3 (N1493, N1469, N520, N1405);
or OR2 (N1494, N1489, N705);
xor XOR2 (N1495, N1481, N1050);
xor XOR2 (N1496, N1482, N882);
not NOT1 (N1497, N1456);
and AND3 (N1498, N1488, N256, N1333);
and AND2 (N1499, N1486, N1063);
nand NAND3 (N1500, N1499, N244, N645);
nor NOR3 (N1501, N1497, N1204, N1291);
buf BUF1 (N1502, N1491);
xor XOR2 (N1503, N1495, N235);
nor NOR3 (N1504, N1502, N1314, N1097);
nor NOR3 (N1505, N1487, N789, N1093);
xor XOR2 (N1506, N1503, N1092);
xor XOR2 (N1507, N1498, N1336);
nand NAND3 (N1508, N1500, N613, N1420);
and AND4 (N1509, N1494, N602, N1353, N145);
not NOT1 (N1510, N1504);
not NOT1 (N1511, N1501);
xor XOR2 (N1512, N1507, N1244);
or OR2 (N1513, N1508, N43);
nor NOR4 (N1514, N1513, N18, N751, N766);
xor XOR2 (N1515, N1506, N171);
buf BUF1 (N1516, N1510);
not NOT1 (N1517, N1511);
nand NAND2 (N1518, N1505, N1484);
nor NOR4 (N1519, N1496, N1057, N1366, N109);
nand NAND4 (N1520, N1516, N697, N226, N582);
nand NAND2 (N1521, N1518, N1320);
or OR2 (N1522, N1512, N169);
not NOT1 (N1523, N1514);
not NOT1 (N1524, N1509);
buf BUF1 (N1525, N1492);
or OR4 (N1526, N1523, N994, N1021, N367);
xor XOR2 (N1527, N1522, N504);
and AND2 (N1528, N1527, N1179);
nand NAND2 (N1529, N1526, N980);
nand NAND2 (N1530, N1521, N1276);
or OR2 (N1531, N1528, N742);
or OR4 (N1532, N1529, N209, N1038, N1145);
not NOT1 (N1533, N1515);
and AND4 (N1534, N1520, N1264, N1064, N587);
xor XOR2 (N1535, N1533, N560);
not NOT1 (N1536, N1534);
not NOT1 (N1537, N1535);
nand NAND4 (N1538, N1493, N1464, N1319, N95);
nor NOR3 (N1539, N1517, N251, N1471);
buf BUF1 (N1540, N1532);
nor NOR2 (N1541, N1530, N85);
nor NOR3 (N1542, N1536, N232, N1303);
buf BUF1 (N1543, N1524);
and AND2 (N1544, N1543, N1278);
and AND2 (N1545, N1539, N763);
not NOT1 (N1546, N1540);
buf BUF1 (N1547, N1525);
nor NOR4 (N1548, N1546, N1383, N1071, N138);
not NOT1 (N1549, N1541);
nor NOR2 (N1550, N1531, N1260);
xor XOR2 (N1551, N1544, N1164);
nor NOR4 (N1552, N1548, N107, N1268, N1309);
or OR4 (N1553, N1551, N1509, N1396, N947);
nand NAND3 (N1554, N1547, N546, N1368);
nor NOR3 (N1555, N1545, N160, N315);
nand NAND2 (N1556, N1550, N1465);
or OR2 (N1557, N1556, N1470);
nand NAND3 (N1558, N1552, N339, N183);
nor NOR2 (N1559, N1519, N402);
buf BUF1 (N1560, N1537);
nand NAND2 (N1561, N1549, N1027);
nor NOR2 (N1562, N1558, N169);
or OR3 (N1563, N1562, N641, N1056);
nor NOR2 (N1564, N1560, N519);
not NOT1 (N1565, N1542);
and AND2 (N1566, N1555, N1316);
or OR2 (N1567, N1553, N840);
and AND2 (N1568, N1538, N280);
not NOT1 (N1569, N1554);
xor XOR2 (N1570, N1563, N19);
xor XOR2 (N1571, N1557, N1290);
and AND3 (N1572, N1565, N1090, N361);
not NOT1 (N1573, N1566);
xor XOR2 (N1574, N1573, N393);
buf BUF1 (N1575, N1561);
xor XOR2 (N1576, N1574, N841);
nor NOR2 (N1577, N1569, N497);
or OR3 (N1578, N1570, N612, N712);
or OR3 (N1579, N1576, N156, N594);
xor XOR2 (N1580, N1559, N1456);
not NOT1 (N1581, N1568);
nor NOR3 (N1582, N1572, N1191, N281);
nand NAND2 (N1583, N1567, N565);
nor NOR4 (N1584, N1577, N1280, N1441, N655);
buf BUF1 (N1585, N1584);
and AND4 (N1586, N1580, N49, N449, N92);
not NOT1 (N1587, N1586);
nand NAND2 (N1588, N1583, N641);
nor NOR4 (N1589, N1578, N569, N229, N399);
and AND4 (N1590, N1575, N648, N801, N924);
not NOT1 (N1591, N1581);
nor NOR2 (N1592, N1587, N1384);
not NOT1 (N1593, N1579);
buf BUF1 (N1594, N1591);
and AND4 (N1595, N1588, N743, N241, N1480);
or OR4 (N1596, N1590, N251, N1344, N1162);
nor NOR4 (N1597, N1582, N146, N681, N347);
not NOT1 (N1598, N1597);
xor XOR2 (N1599, N1596, N906);
nor NOR3 (N1600, N1598, N351, N142);
buf BUF1 (N1601, N1564);
nand NAND2 (N1602, N1571, N780);
xor XOR2 (N1603, N1592, N1211);
buf BUF1 (N1604, N1593);
nand NAND4 (N1605, N1599, N1164, N1493, N842);
nand NAND2 (N1606, N1602, N473);
buf BUF1 (N1607, N1600);
or OR3 (N1608, N1607, N1188, N65);
xor XOR2 (N1609, N1585, N135);
buf BUF1 (N1610, N1608);
buf BUF1 (N1611, N1595);
or OR3 (N1612, N1594, N700, N847);
nand NAND4 (N1613, N1606, N167, N957, N1137);
and AND4 (N1614, N1613, N720, N1280, N443);
buf BUF1 (N1615, N1604);
or OR3 (N1616, N1615, N1345, N1282);
buf BUF1 (N1617, N1611);
and AND2 (N1618, N1603, N1529);
xor XOR2 (N1619, N1609, N1493);
nor NOR2 (N1620, N1605, N1310);
not NOT1 (N1621, N1618);
not NOT1 (N1622, N1610);
not NOT1 (N1623, N1622);
and AND2 (N1624, N1614, N1263);
nand NAND2 (N1625, N1620, N664);
not NOT1 (N1626, N1616);
buf BUF1 (N1627, N1623);
nand NAND4 (N1628, N1589, N429, N415, N1520);
xor XOR2 (N1629, N1617, N1058);
buf BUF1 (N1630, N1625);
and AND3 (N1631, N1624, N1446, N1377);
and AND2 (N1632, N1630, N1031);
and AND3 (N1633, N1629, N635, N1520);
nand NAND4 (N1634, N1632, N1410, N1569, N1431);
buf BUF1 (N1635, N1601);
and AND2 (N1636, N1621, N1462);
nor NOR3 (N1637, N1636, N732, N492);
nor NOR4 (N1638, N1612, N376, N966, N920);
xor XOR2 (N1639, N1634, N1521);
not NOT1 (N1640, N1637);
or OR4 (N1641, N1633, N176, N106, N1428);
or OR2 (N1642, N1640, N840);
nand NAND4 (N1643, N1635, N1017, N1548, N135);
xor XOR2 (N1644, N1642, N407);
buf BUF1 (N1645, N1641);
buf BUF1 (N1646, N1619);
not NOT1 (N1647, N1646);
and AND2 (N1648, N1627, N922);
nor NOR2 (N1649, N1639, N874);
buf BUF1 (N1650, N1645);
or OR2 (N1651, N1631, N825);
and AND2 (N1652, N1643, N1289);
and AND4 (N1653, N1652, N1154, N727, N1607);
xor XOR2 (N1654, N1650, N386);
and AND3 (N1655, N1649, N1202, N30);
xor XOR2 (N1656, N1651, N1336);
nand NAND3 (N1657, N1638, N69, N1580);
or OR2 (N1658, N1657, N1171);
buf BUF1 (N1659, N1628);
or OR4 (N1660, N1644, N1630, N166, N1053);
and AND4 (N1661, N1653, N1596, N890, N98);
nor NOR2 (N1662, N1654, N1024);
nand NAND2 (N1663, N1659, N526);
nand NAND2 (N1664, N1662, N1575);
nand NAND4 (N1665, N1647, N554, N396, N798);
not NOT1 (N1666, N1648);
nor NOR4 (N1667, N1664, N762, N688, N107);
nand NAND3 (N1668, N1663, N1345, N830);
xor XOR2 (N1669, N1668, N860);
buf BUF1 (N1670, N1665);
and AND3 (N1671, N1626, N452, N1633);
buf BUF1 (N1672, N1655);
or OR3 (N1673, N1660, N466, N1522);
or OR4 (N1674, N1666, N1187, N172, N231);
or OR2 (N1675, N1661, N101);
nand NAND4 (N1676, N1673, N1007, N1272, N1522);
xor XOR2 (N1677, N1667, N302);
xor XOR2 (N1678, N1672, N530);
or OR2 (N1679, N1678, N642);
and AND4 (N1680, N1675, N190, N1596, N456);
nand NAND2 (N1681, N1671, N811);
and AND3 (N1682, N1680, N422, N1391);
nand NAND2 (N1683, N1679, N1474);
xor XOR2 (N1684, N1669, N882);
and AND3 (N1685, N1670, N1027, N958);
not NOT1 (N1686, N1681);
xor XOR2 (N1687, N1676, N485);
and AND4 (N1688, N1658, N218, N1045, N558);
nand NAND3 (N1689, N1685, N1203, N151);
nand NAND4 (N1690, N1686, N835, N1329, N775);
or OR3 (N1691, N1682, N1306, N201);
buf BUF1 (N1692, N1689);
nand NAND3 (N1693, N1690, N1602, N1238);
buf BUF1 (N1694, N1656);
nor NOR3 (N1695, N1684, N295, N1192);
nor NOR2 (N1696, N1694, N524);
and AND4 (N1697, N1691, N232, N765, N460);
xor XOR2 (N1698, N1677, N1165);
and AND3 (N1699, N1693, N1383, N629);
buf BUF1 (N1700, N1696);
and AND3 (N1701, N1698, N1264, N440);
nor NOR2 (N1702, N1700, N201);
or OR2 (N1703, N1695, N989);
and AND2 (N1704, N1674, N596);
buf BUF1 (N1705, N1692);
not NOT1 (N1706, N1687);
and AND3 (N1707, N1699, N1256, N461);
and AND2 (N1708, N1707, N185);
nor NOR2 (N1709, N1683, N709);
xor XOR2 (N1710, N1706, N342);
nand NAND4 (N1711, N1701, N545, N1555, N1047);
or OR4 (N1712, N1703, N1286, N648, N554);
nor NOR3 (N1713, N1712, N924, N1092);
or OR3 (N1714, N1711, N315, N782);
or OR4 (N1715, N1713, N1409, N485, N495);
buf BUF1 (N1716, N1710);
and AND4 (N1717, N1688, N18, N898, N891);
nor NOR3 (N1718, N1715, N1435, N1515);
nand NAND3 (N1719, N1697, N1689, N735);
or OR4 (N1720, N1709, N28, N400, N205);
buf BUF1 (N1721, N1717);
not NOT1 (N1722, N1714);
or OR4 (N1723, N1716, N1285, N1114, N1685);
nor NOR2 (N1724, N1719, N838);
nand NAND3 (N1725, N1724, N18, N1546);
nor NOR3 (N1726, N1723, N11, N493);
and AND2 (N1727, N1726, N1178);
buf BUF1 (N1728, N1720);
or OR4 (N1729, N1704, N1401, N1122, N1371);
or OR3 (N1730, N1721, N626, N484);
and AND3 (N1731, N1718, N723, N1198);
and AND4 (N1732, N1729, N1208, N227, N1529);
xor XOR2 (N1733, N1728, N181);
nand NAND4 (N1734, N1731, N475, N836, N1631);
xor XOR2 (N1735, N1705, N508);
and AND4 (N1736, N1708, N1195, N71, N1584);
not NOT1 (N1737, N1730);
not NOT1 (N1738, N1733);
or OR3 (N1739, N1727, N75, N420);
xor XOR2 (N1740, N1734, N1473);
xor XOR2 (N1741, N1739, N1381);
xor XOR2 (N1742, N1722, N1555);
or OR4 (N1743, N1736, N1008, N749, N1111);
or OR2 (N1744, N1743, N903);
not NOT1 (N1745, N1740);
nand NAND4 (N1746, N1702, N1391, N1236, N1426);
nor NOR4 (N1747, N1725, N525, N1346, N1274);
xor XOR2 (N1748, N1732, N1492);
nand NAND4 (N1749, N1745, N363, N1093, N834);
not NOT1 (N1750, N1735);
xor XOR2 (N1751, N1737, N694);
not NOT1 (N1752, N1741);
xor XOR2 (N1753, N1748, N1587);
buf BUF1 (N1754, N1744);
xor XOR2 (N1755, N1749, N312);
buf BUF1 (N1756, N1747);
and AND3 (N1757, N1746, N1601, N1420);
buf BUF1 (N1758, N1756);
nand NAND2 (N1759, N1758, N1085);
nand NAND4 (N1760, N1751, N1490, N846, N1146);
nand NAND2 (N1761, N1754, N768);
buf BUF1 (N1762, N1753);
not NOT1 (N1763, N1752);
nor NOR3 (N1764, N1755, N1322, N1438);
nor NOR3 (N1765, N1764, N1079, N389);
and AND4 (N1766, N1738, N1371, N1682, N1019);
and AND4 (N1767, N1750, N630, N1137, N729);
nand NAND2 (N1768, N1767, N687);
nand NAND3 (N1769, N1761, N660, N129);
buf BUF1 (N1770, N1768);
nor NOR4 (N1771, N1760, N269, N1663, N1645);
xor XOR2 (N1772, N1757, N1318);
and AND3 (N1773, N1762, N395, N45);
not NOT1 (N1774, N1772);
buf BUF1 (N1775, N1766);
nand NAND4 (N1776, N1759, N311, N598, N1258);
or OR3 (N1777, N1765, N297, N1050);
xor XOR2 (N1778, N1773, N310);
buf BUF1 (N1779, N1774);
xor XOR2 (N1780, N1771, N190);
not NOT1 (N1781, N1775);
and AND3 (N1782, N1779, N120, N1022);
not NOT1 (N1783, N1776);
buf BUF1 (N1784, N1780);
and AND4 (N1785, N1778, N374, N1086, N1127);
or OR2 (N1786, N1777, N751);
not NOT1 (N1787, N1781);
or OR2 (N1788, N1787, N1438);
nor NOR2 (N1789, N1763, N883);
nand NAND3 (N1790, N1770, N1117, N917);
buf BUF1 (N1791, N1789);
buf BUF1 (N1792, N1788);
xor XOR2 (N1793, N1791, N1489);
not NOT1 (N1794, N1784);
nor NOR3 (N1795, N1783, N941, N411);
xor XOR2 (N1796, N1793, N823);
xor XOR2 (N1797, N1796, N60);
and AND2 (N1798, N1785, N1362);
nand NAND3 (N1799, N1797, N504, N739);
nand NAND2 (N1800, N1790, N1630);
not NOT1 (N1801, N1769);
nor NOR2 (N1802, N1799, N478);
not NOT1 (N1803, N1798);
nor NOR3 (N1804, N1795, N1101, N89);
xor XOR2 (N1805, N1742, N216);
or OR3 (N1806, N1800, N537, N859);
xor XOR2 (N1807, N1794, N115);
buf BUF1 (N1808, N1803);
xor XOR2 (N1809, N1804, N1554);
buf BUF1 (N1810, N1782);
or OR3 (N1811, N1792, N1789, N970);
not NOT1 (N1812, N1808);
xor XOR2 (N1813, N1811, N1331);
or OR4 (N1814, N1810, N860, N430, N539);
and AND3 (N1815, N1801, N171, N1689);
and AND4 (N1816, N1815, N1681, N873, N360);
buf BUF1 (N1817, N1809);
or OR2 (N1818, N1807, N59);
xor XOR2 (N1819, N1806, N1743);
and AND4 (N1820, N1816, N1108, N1682, N821);
not NOT1 (N1821, N1820);
or OR4 (N1822, N1786, N671, N650, N540);
nand NAND3 (N1823, N1813, N705, N193);
nand NAND4 (N1824, N1802, N1168, N1638, N879);
nor NOR2 (N1825, N1814, N1535);
nor NOR3 (N1826, N1812, N1514, N1642);
buf BUF1 (N1827, N1818);
nand NAND3 (N1828, N1821, N1165, N464);
nor NOR3 (N1829, N1822, N56, N402);
nand NAND3 (N1830, N1826, N351, N947);
buf BUF1 (N1831, N1823);
and AND4 (N1832, N1817, N1249, N1632, N1355);
nand NAND2 (N1833, N1832, N1403);
nand NAND3 (N1834, N1830, N1781, N1004);
or OR4 (N1835, N1831, N1022, N256, N812);
nand NAND3 (N1836, N1819, N1699, N1607);
buf BUF1 (N1837, N1835);
xor XOR2 (N1838, N1834, N42);
nand NAND4 (N1839, N1837, N1319, N1403, N390);
nand NAND2 (N1840, N1805, N903);
buf BUF1 (N1841, N1827);
xor XOR2 (N1842, N1824, N136);
and AND3 (N1843, N1829, N713, N1031);
or OR3 (N1844, N1843, N789, N898);
nor NOR3 (N1845, N1838, N116, N1274);
and AND3 (N1846, N1840, N947, N738);
nand NAND4 (N1847, N1833, N298, N1666, N1528);
xor XOR2 (N1848, N1836, N445);
xor XOR2 (N1849, N1825, N1226);
nand NAND2 (N1850, N1848, N438);
or OR2 (N1851, N1846, N1812);
not NOT1 (N1852, N1847);
and AND3 (N1853, N1844, N1696, N1358);
xor XOR2 (N1854, N1851, N1119);
buf BUF1 (N1855, N1850);
or OR4 (N1856, N1849, N1203, N97, N316);
not NOT1 (N1857, N1855);
buf BUF1 (N1858, N1841);
or OR4 (N1859, N1852, N918, N463, N858);
nor NOR3 (N1860, N1859, N1298, N1361);
nand NAND3 (N1861, N1860, N1831, N94);
nor NOR2 (N1862, N1845, N1759);
and AND2 (N1863, N1853, N1538);
xor XOR2 (N1864, N1839, N1835);
nor NOR4 (N1865, N1864, N1824, N1091, N232);
nor NOR3 (N1866, N1865, N1266, N1446);
nand NAND4 (N1867, N1861, N1464, N1150, N1579);
and AND3 (N1868, N1854, N1032, N1788);
and AND4 (N1869, N1858, N572, N120, N1756);
or OR4 (N1870, N1842, N794, N1841, N1716);
not NOT1 (N1871, N1868);
and AND3 (N1872, N1863, N1622, N1394);
buf BUF1 (N1873, N1871);
nor NOR4 (N1874, N1869, N1746, N40, N1142);
or OR2 (N1875, N1870, N100);
and AND4 (N1876, N1873, N1700, N1770, N679);
and AND3 (N1877, N1872, N349, N1);
or OR4 (N1878, N1876, N1206, N1546, N1778);
nand NAND2 (N1879, N1857, N124);
nor NOR4 (N1880, N1867, N1847, N1774, N1212);
buf BUF1 (N1881, N1879);
nor NOR3 (N1882, N1877, N576, N531);
or OR3 (N1883, N1866, N156, N849);
not NOT1 (N1884, N1883);
not NOT1 (N1885, N1882);
or OR3 (N1886, N1881, N599, N763);
not NOT1 (N1887, N1878);
buf BUF1 (N1888, N1887);
nor NOR4 (N1889, N1888, N1006, N301, N64);
or OR4 (N1890, N1856, N628, N162, N1728);
buf BUF1 (N1891, N1828);
buf BUF1 (N1892, N1886);
not NOT1 (N1893, N1885);
xor XOR2 (N1894, N1890, N1841);
and AND4 (N1895, N1880, N1626, N1845, N1807);
or OR3 (N1896, N1894, N1753, N1256);
buf BUF1 (N1897, N1893);
and AND4 (N1898, N1862, N686, N1805, N1717);
not NOT1 (N1899, N1889);
buf BUF1 (N1900, N1875);
nor NOR4 (N1901, N1900, N845, N1639, N772);
not NOT1 (N1902, N1901);
and AND3 (N1903, N1902, N646, N449);
nand NAND4 (N1904, N1896, N1752, N1255, N904);
nand NAND3 (N1905, N1891, N1294, N1741);
buf BUF1 (N1906, N1905);
nand NAND4 (N1907, N1895, N1905, N1872, N1149);
or OR3 (N1908, N1884, N1235, N1505);
not NOT1 (N1909, N1892);
or OR2 (N1910, N1898, N1780);
or OR2 (N1911, N1910, N1438);
xor XOR2 (N1912, N1899, N1880);
and AND3 (N1913, N1906, N1043, N744);
or OR2 (N1914, N1907, N1208);
and AND3 (N1915, N1908, N1053, N601);
buf BUF1 (N1916, N1915);
not NOT1 (N1917, N1874);
xor XOR2 (N1918, N1917, N799);
or OR4 (N1919, N1912, N278, N1087, N1597);
or OR3 (N1920, N1911, N382, N1585);
buf BUF1 (N1921, N1919);
nor NOR2 (N1922, N1916, N1348);
xor XOR2 (N1923, N1909, N65);
and AND3 (N1924, N1921, N815, N767);
not NOT1 (N1925, N1918);
xor XOR2 (N1926, N1920, N1848);
buf BUF1 (N1927, N1913);
not NOT1 (N1928, N1903);
nand NAND2 (N1929, N1922, N122);
nor NOR2 (N1930, N1928, N1370);
xor XOR2 (N1931, N1897, N657);
buf BUF1 (N1932, N1931);
and AND2 (N1933, N1904, N1380);
and AND2 (N1934, N1924, N302);
and AND3 (N1935, N1923, N712, N328);
xor XOR2 (N1936, N1934, N947);
xor XOR2 (N1937, N1929, N780);
buf BUF1 (N1938, N1925);
nor NOR2 (N1939, N1926, N1879);
and AND4 (N1940, N1935, N1491, N681, N1325);
nand NAND4 (N1941, N1937, N1324, N1927, N1592);
and AND3 (N1942, N215, N626, N705);
and AND2 (N1943, N1936, N1421);
nor NOR4 (N1944, N1914, N1809, N1759, N1646);
nor NOR4 (N1945, N1940, N1397, N1159, N1721);
or OR2 (N1946, N1938, N945);
nand NAND4 (N1947, N1945, N138, N248, N716);
buf BUF1 (N1948, N1947);
not NOT1 (N1949, N1944);
or OR4 (N1950, N1932, N1348, N224, N1012);
nor NOR3 (N1951, N1949, N1736, N691);
or OR3 (N1952, N1939, N1919, N1519);
not NOT1 (N1953, N1941);
nand NAND3 (N1954, N1953, N1381, N528);
not NOT1 (N1955, N1948);
and AND4 (N1956, N1951, N1208, N855, N1253);
nor NOR2 (N1957, N1952, N72);
not NOT1 (N1958, N1954);
and AND3 (N1959, N1930, N1086, N631);
not NOT1 (N1960, N1933);
xor XOR2 (N1961, N1960, N661);
or OR2 (N1962, N1958, N963);
xor XOR2 (N1963, N1959, N1911);
buf BUF1 (N1964, N1957);
nand NAND3 (N1965, N1950, N1952, N1596);
or OR2 (N1966, N1942, N93);
xor XOR2 (N1967, N1946, N1881);
xor XOR2 (N1968, N1964, N323);
not NOT1 (N1969, N1943);
buf BUF1 (N1970, N1961);
buf BUF1 (N1971, N1966);
buf BUF1 (N1972, N1968);
or OR2 (N1973, N1969, N1652);
buf BUF1 (N1974, N1970);
and AND2 (N1975, N1972, N1332);
or OR3 (N1976, N1963, N1009, N1386);
and AND2 (N1977, N1971, N1234);
xor XOR2 (N1978, N1973, N1933);
xor XOR2 (N1979, N1956, N32);
xor XOR2 (N1980, N1955, N1232);
nand NAND3 (N1981, N1974, N1685, N1574);
nand NAND4 (N1982, N1977, N914, N1060, N800);
nand NAND2 (N1983, N1965, N676);
or OR3 (N1984, N1982, N637, N1799);
nand NAND2 (N1985, N1967, N526);
and AND2 (N1986, N1981, N70);
buf BUF1 (N1987, N1975);
not NOT1 (N1988, N1976);
buf BUF1 (N1989, N1980);
buf BUF1 (N1990, N1979);
or OR2 (N1991, N1983, N110);
or OR4 (N1992, N1991, N1797, N561, N1022);
buf BUF1 (N1993, N1985);
xor XOR2 (N1994, N1987, N1353);
and AND2 (N1995, N1986, N1975);
or OR4 (N1996, N1962, N304, N840, N1644);
not NOT1 (N1997, N1984);
nor NOR3 (N1998, N1978, N714, N1924);
xor XOR2 (N1999, N1996, N885);
not NOT1 (N2000, N1998);
or OR2 (N2001, N1992, N1586);
or OR4 (N2002, N2001, N418, N1071, N875);
nor NOR2 (N2003, N1989, N1832);
nor NOR2 (N2004, N1997, N225);
not NOT1 (N2005, N2004);
not NOT1 (N2006, N1994);
or OR4 (N2007, N2005, N981, N1425, N1026);
nor NOR2 (N2008, N2007, N649);
nor NOR2 (N2009, N2006, N841);
not NOT1 (N2010, N1999);
buf BUF1 (N2011, N1988);
nand NAND2 (N2012, N2010, N575);
or OR4 (N2013, N2011, N483, N824, N225);
xor XOR2 (N2014, N2002, N1252);
xor XOR2 (N2015, N2012, N877);
buf BUF1 (N2016, N2014);
nand NAND4 (N2017, N2016, N1879, N1965, N437);
nor NOR4 (N2018, N2009, N103, N1163, N402);
not NOT1 (N2019, N2003);
and AND4 (N2020, N2008, N1308, N1790, N1153);
not NOT1 (N2021, N1993);
and AND3 (N2022, N1990, N1046, N1742);
nor NOR3 (N2023, N2018, N198, N1019);
nand NAND2 (N2024, N2017, N1959);
not NOT1 (N2025, N2023);
nand NAND4 (N2026, N2013, N941, N257, N525);
and AND2 (N2027, N2015, N1920);
buf BUF1 (N2028, N2022);
not NOT1 (N2029, N2025);
not NOT1 (N2030, N2021);
and AND2 (N2031, N2029, N417);
not NOT1 (N2032, N2027);
nand NAND2 (N2033, N2020, N162);
xor XOR2 (N2034, N2030, N1736);
or OR3 (N2035, N1995, N191, N439);
or OR2 (N2036, N2033, N320);
not NOT1 (N2037, N2024);
not NOT1 (N2038, N2026);
and AND3 (N2039, N2028, N1052, N562);
not NOT1 (N2040, N2019);
not NOT1 (N2041, N2032);
nor NOR2 (N2042, N2034, N940);
and AND3 (N2043, N2039, N666, N641);
xor XOR2 (N2044, N2031, N713);
buf BUF1 (N2045, N2041);
and AND3 (N2046, N2040, N1971, N650);
not NOT1 (N2047, N2043);
nor NOR3 (N2048, N2000, N419, N1562);
not NOT1 (N2049, N2037);
or OR2 (N2050, N2045, N1612);
xor XOR2 (N2051, N2047, N661);
not NOT1 (N2052, N2042);
not NOT1 (N2053, N2048);
nand NAND4 (N2054, N2049, N624, N318, N1499);
buf BUF1 (N2055, N2044);
not NOT1 (N2056, N2046);
not NOT1 (N2057, N2054);
or OR4 (N2058, N2056, N1463, N1783, N284);
xor XOR2 (N2059, N2052, N1196);
buf BUF1 (N2060, N2050);
and AND3 (N2061, N2055, N1198, N281);
or OR3 (N2062, N2059, N1474, N469);
buf BUF1 (N2063, N2035);
nor NOR4 (N2064, N2051, N1844, N2060, N47);
not NOT1 (N2065, N1951);
nand NAND2 (N2066, N2064, N244);
or OR4 (N2067, N2063, N1913, N133, N578);
nor NOR3 (N2068, N2053, N453, N942);
not NOT1 (N2069, N2057);
and AND2 (N2070, N2061, N1069);
xor XOR2 (N2071, N2058, N1357);
and AND4 (N2072, N2067, N294, N301, N115);
or OR3 (N2073, N2072, N1315, N598);
xor XOR2 (N2074, N2069, N1116);
buf BUF1 (N2075, N2070);
or OR3 (N2076, N2071, N1400, N656);
and AND4 (N2077, N2074, N294, N2068, N1149);
buf BUF1 (N2078, N1162);
xor XOR2 (N2079, N2065, N111);
buf BUF1 (N2080, N2077);
not NOT1 (N2081, N2036);
nand NAND3 (N2082, N2080, N186, N938);
nor NOR2 (N2083, N2081, N551);
buf BUF1 (N2084, N2073);
buf BUF1 (N2085, N2075);
nand NAND2 (N2086, N2066, N1883);
nor NOR4 (N2087, N2078, N1089, N1052, N330);
and AND4 (N2088, N2076, N931, N93, N501);
not NOT1 (N2089, N2079);
nor NOR4 (N2090, N2038, N1003, N826, N28);
xor XOR2 (N2091, N2084, N988);
nor NOR3 (N2092, N2083, N1426, N1277);
xor XOR2 (N2093, N2082, N260);
and AND4 (N2094, N2087, N450, N1057, N1961);
nor NOR4 (N2095, N2093, N1985, N1747, N1777);
nor NOR4 (N2096, N2089, N1748, N1510, N500);
buf BUF1 (N2097, N2095);
and AND2 (N2098, N2085, N1933);
nand NAND4 (N2099, N2090, N105, N1672, N1664);
and AND4 (N2100, N2088, N630, N1376, N1729);
or OR4 (N2101, N2098, N1497, N1712, N1281);
nand NAND4 (N2102, N2091, N1040, N2074, N1170);
nand NAND3 (N2103, N2086, N2055, N340);
and AND2 (N2104, N2102, N223);
nand NAND3 (N2105, N2094, N1542, N1336);
xor XOR2 (N2106, N2097, N1520);
xor XOR2 (N2107, N2099, N1745);
xor XOR2 (N2108, N2105, N1390);
xor XOR2 (N2109, N2107, N628);
buf BUF1 (N2110, N2109);
nand NAND2 (N2111, N2104, N1272);
or OR3 (N2112, N2111, N1415, N47);
buf BUF1 (N2113, N2101);
not NOT1 (N2114, N2106);
nor NOR4 (N2115, N2113, N1547, N1738, N2101);
xor XOR2 (N2116, N2114, N465);
not NOT1 (N2117, N2108);
or OR2 (N2118, N2062, N235);
buf BUF1 (N2119, N2100);
buf BUF1 (N2120, N2096);
or OR2 (N2121, N2103, N2050);
buf BUF1 (N2122, N2117);
nand NAND3 (N2123, N2115, N2009, N209);
nor NOR4 (N2124, N2116, N1386, N1049, N362);
or OR2 (N2125, N2112, N1759);
not NOT1 (N2126, N2119);
and AND2 (N2127, N2118, N132);
nand NAND4 (N2128, N2123, N43, N1138, N137);
or OR3 (N2129, N2126, N397, N1684);
nor NOR4 (N2130, N2124, N933, N1792, N868);
xor XOR2 (N2131, N2127, N413);
nor NOR3 (N2132, N2121, N1842, N205);
or OR2 (N2133, N2131, N1618);
nand NAND2 (N2134, N2133, N286);
not NOT1 (N2135, N2120);
xor XOR2 (N2136, N2130, N1160);
nand NAND4 (N2137, N2122, N274, N731, N1167);
not NOT1 (N2138, N2125);
or OR4 (N2139, N2128, N778, N467, N1144);
nand NAND4 (N2140, N2132, N200, N60, N323);
nand NAND3 (N2141, N2140, N1360, N523);
nor NOR2 (N2142, N2110, N1170);
and AND4 (N2143, N2141, N470, N1372, N815);
nor NOR2 (N2144, N2137, N902);
and AND3 (N2145, N2143, N507, N1596);
or OR3 (N2146, N2134, N850, N1843);
buf BUF1 (N2147, N2139);
nor NOR4 (N2148, N2147, N960, N1251, N1540);
nor NOR3 (N2149, N2145, N1392, N383);
not NOT1 (N2150, N2129);
buf BUF1 (N2151, N2138);
nand NAND2 (N2152, N2142, N1253);
or OR4 (N2153, N2151, N553, N107, N248);
and AND4 (N2154, N2092, N139, N1352, N30);
not NOT1 (N2155, N2144);
xor XOR2 (N2156, N2149, N259);
nor NOR4 (N2157, N2136, N701, N828, N1207);
or OR3 (N2158, N2155, N875, N1549);
xor XOR2 (N2159, N2150, N2019);
not NOT1 (N2160, N2148);
nand NAND4 (N2161, N2157, N368, N2069, N1175);
not NOT1 (N2162, N2156);
nor NOR3 (N2163, N2162, N905, N1697);
xor XOR2 (N2164, N2161, N462);
xor XOR2 (N2165, N2135, N567);
buf BUF1 (N2166, N2153);
and AND4 (N2167, N2152, N739, N965, N23);
and AND2 (N2168, N2164, N67);
and AND2 (N2169, N2160, N168);
buf BUF1 (N2170, N2146);
or OR2 (N2171, N2166, N1919);
xor XOR2 (N2172, N2159, N967);
or OR2 (N2173, N2170, N1345);
or OR4 (N2174, N2165, N757, N1117, N1206);
and AND4 (N2175, N2172, N407, N169, N1423);
not NOT1 (N2176, N2154);
and AND2 (N2177, N2167, N1978);
nor NOR3 (N2178, N2175, N297, N925);
buf BUF1 (N2179, N2169);
not NOT1 (N2180, N2163);
or OR3 (N2181, N2180, N712, N1643);
not NOT1 (N2182, N2181);
nor NOR2 (N2183, N2176, N1005);
not NOT1 (N2184, N2158);
or OR3 (N2185, N2178, N940, N625);
xor XOR2 (N2186, N2184, N1208);
or OR4 (N2187, N2183, N33, N1936, N1149);
xor XOR2 (N2188, N2179, N287);
nand NAND4 (N2189, N2186, N163, N2076, N1112);
buf BUF1 (N2190, N2185);
buf BUF1 (N2191, N2171);
xor XOR2 (N2192, N2191, N516);
not NOT1 (N2193, N2177);
and AND2 (N2194, N2190, N462);
nor NOR2 (N2195, N2173, N894);
nand NAND3 (N2196, N2182, N1350, N1559);
or OR4 (N2197, N2196, N882, N1197, N770);
and AND4 (N2198, N2197, N922, N1294, N822);
xor XOR2 (N2199, N2198, N1258);
not NOT1 (N2200, N2189);
nor NOR2 (N2201, N2199, N43);
buf BUF1 (N2202, N2195);
or OR2 (N2203, N2201, N664);
xor XOR2 (N2204, N2168, N902);
nand NAND3 (N2205, N2188, N1140, N2134);
not NOT1 (N2206, N2204);
xor XOR2 (N2207, N2202, N1881);
or OR2 (N2208, N2187, N2160);
nand NAND3 (N2209, N2203, N704, N1890);
nor NOR4 (N2210, N2193, N1421, N1415, N665);
and AND2 (N2211, N2208, N87);
and AND2 (N2212, N2174, N1177);
nand NAND4 (N2213, N2212, N1787, N1563, N1184);
nand NAND4 (N2214, N2211, N1282, N2112, N836);
and AND4 (N2215, N2209, N1548, N768, N923);
nand NAND4 (N2216, N2210, N2186, N328, N452);
nor NOR2 (N2217, N2200, N840);
nand NAND4 (N2218, N2192, N2042, N1403, N1796);
or OR2 (N2219, N2217, N1004);
and AND4 (N2220, N2214, N519, N502, N647);
not NOT1 (N2221, N2207);
not NOT1 (N2222, N2221);
and AND3 (N2223, N2219, N1965, N1097);
xor XOR2 (N2224, N2216, N646);
and AND4 (N2225, N2213, N1793, N1970, N809);
nor NOR2 (N2226, N2224, N1335);
and AND2 (N2227, N2220, N2013);
xor XOR2 (N2228, N2194, N2121);
xor XOR2 (N2229, N2218, N291);
and AND3 (N2230, N2222, N71, N1296);
xor XOR2 (N2231, N2215, N1394);
nand NAND4 (N2232, N2231, N2074, N982, N1865);
buf BUF1 (N2233, N2225);
or OR2 (N2234, N2205, N1107);
not NOT1 (N2235, N2227);
nor NOR3 (N2236, N2234, N592, N1038);
nand NAND2 (N2237, N2228, N1295);
not NOT1 (N2238, N2226);
and AND3 (N2239, N2223, N947, N248);
nor NOR2 (N2240, N2236, N1348);
nor NOR3 (N2241, N2237, N807, N1713);
or OR3 (N2242, N2240, N204, N529);
and AND4 (N2243, N2232, N815, N789, N683);
nor NOR2 (N2244, N2242, N1275);
nor NOR2 (N2245, N2233, N1001);
or OR2 (N2246, N2229, N772);
nand NAND4 (N2247, N2243, N2210, N2137, N851);
buf BUF1 (N2248, N2245);
buf BUF1 (N2249, N2241);
xor XOR2 (N2250, N2247, N229);
nor NOR2 (N2251, N2238, N420);
xor XOR2 (N2252, N2249, N1322);
not NOT1 (N2253, N2206);
nor NOR4 (N2254, N2230, N1555, N785, N1744);
buf BUF1 (N2255, N2250);
nor NOR3 (N2256, N2246, N2096, N1099);
buf BUF1 (N2257, N2255);
not NOT1 (N2258, N2239);
nor NOR3 (N2259, N2253, N691, N1734);
or OR4 (N2260, N2248, N505, N1905, N371);
and AND4 (N2261, N2252, N508, N1063, N1432);
nand NAND4 (N2262, N2254, N2106, N277, N555);
nor NOR2 (N2263, N2244, N1123);
nand NAND4 (N2264, N2261, N1437, N2005, N1217);
not NOT1 (N2265, N2259);
xor XOR2 (N2266, N2235, N876);
nor NOR3 (N2267, N2251, N1647, N936);
not NOT1 (N2268, N2263);
not NOT1 (N2269, N2264);
or OR4 (N2270, N2260, N677, N2207, N2032);
or OR4 (N2271, N2270, N857, N2170, N1202);
not NOT1 (N2272, N2256);
or OR2 (N2273, N2267, N452);
xor XOR2 (N2274, N2266, N824);
xor XOR2 (N2275, N2271, N1786);
xor XOR2 (N2276, N2272, N2239);
not NOT1 (N2277, N2265);
or OR4 (N2278, N2275, N361, N1394, N1134);
not NOT1 (N2279, N2262);
or OR4 (N2280, N2273, N243, N915, N774);
not NOT1 (N2281, N2280);
not NOT1 (N2282, N2281);
xor XOR2 (N2283, N2274, N296);
not NOT1 (N2284, N2269);
and AND3 (N2285, N2258, N2051, N1398);
not NOT1 (N2286, N2276);
not NOT1 (N2287, N2279);
or OR2 (N2288, N2268, N166);
and AND4 (N2289, N2257, N1201, N572, N213);
and AND4 (N2290, N2286, N541, N633, N2100);
buf BUF1 (N2291, N2288);
nand NAND3 (N2292, N2291, N252, N1818);
xor XOR2 (N2293, N2285, N771);
nand NAND2 (N2294, N2282, N624);
or OR3 (N2295, N2277, N2080, N1806);
nand NAND3 (N2296, N2278, N1266, N1305);
xor XOR2 (N2297, N2294, N980);
nand NAND3 (N2298, N2284, N173, N1994);
nand NAND3 (N2299, N2296, N333, N1583);
and AND3 (N2300, N2287, N899, N1566);
and AND4 (N2301, N2295, N683, N1275, N1656);
nand NAND2 (N2302, N2297, N1523);
and AND3 (N2303, N2300, N1, N391);
buf BUF1 (N2304, N2293);
nand NAND2 (N2305, N2289, N1718);
or OR2 (N2306, N2302, N596);
or OR2 (N2307, N2301, N2196);
buf BUF1 (N2308, N2290);
nor NOR4 (N2309, N2305, N1845, N288, N1602);
or OR2 (N2310, N2299, N1605);
not NOT1 (N2311, N2310);
and AND4 (N2312, N2283, N1608, N1522, N853);
and AND4 (N2313, N2298, N878, N2256, N1452);
and AND2 (N2314, N2308, N2083);
or OR4 (N2315, N2303, N1827, N1824, N1300);
not NOT1 (N2316, N2292);
not NOT1 (N2317, N2316);
and AND3 (N2318, N2306, N681, N182);
not NOT1 (N2319, N2313);
nor NOR2 (N2320, N2311, N220);
nor NOR3 (N2321, N2307, N2320, N1278);
nand NAND3 (N2322, N2078, N368, N293);
nor NOR4 (N2323, N2312, N966, N2154, N2318);
xor XOR2 (N2324, N1639, N280);
nand NAND4 (N2325, N2323, N2268, N178, N233);
nand NAND3 (N2326, N2324, N1626, N1023);
and AND2 (N2327, N2325, N1645);
xor XOR2 (N2328, N2321, N1931);
buf BUF1 (N2329, N2314);
xor XOR2 (N2330, N2328, N208);
or OR2 (N2331, N2329, N1919);
buf BUF1 (N2332, N2304);
not NOT1 (N2333, N2331);
nand NAND4 (N2334, N2333, N503, N857, N1575);
not NOT1 (N2335, N2327);
xor XOR2 (N2336, N2332, N947);
and AND2 (N2337, N2317, N437);
nand NAND3 (N2338, N2322, N1288, N1906);
not NOT1 (N2339, N2330);
nand NAND2 (N2340, N2319, N216);
not NOT1 (N2341, N2336);
not NOT1 (N2342, N2334);
nor NOR2 (N2343, N2342, N1173);
nand NAND4 (N2344, N2343, N475, N637, N549);
not NOT1 (N2345, N2326);
xor XOR2 (N2346, N2315, N1708);
nor NOR3 (N2347, N2338, N1997, N622);
and AND3 (N2348, N2340, N2248, N1960);
nand NAND2 (N2349, N2339, N1546);
or OR2 (N2350, N2309, N2017);
buf BUF1 (N2351, N2335);
nor NOR2 (N2352, N2346, N860);
nand NAND3 (N2353, N2337, N1494, N719);
or OR2 (N2354, N2345, N1833);
or OR4 (N2355, N2353, N2290, N1868, N1345);
not NOT1 (N2356, N2349);
xor XOR2 (N2357, N2344, N2275);
not NOT1 (N2358, N2354);
not NOT1 (N2359, N2348);
or OR2 (N2360, N2355, N645);
or OR2 (N2361, N2360, N1035);
nand NAND3 (N2362, N2352, N134, N367);
or OR2 (N2363, N2356, N758);
not NOT1 (N2364, N2362);
not NOT1 (N2365, N2361);
or OR2 (N2366, N2358, N2230);
not NOT1 (N2367, N2365);
nor NOR4 (N2368, N2364, N976, N1172, N1035);
nor NOR2 (N2369, N2363, N751);
nand NAND3 (N2370, N2366, N1120, N740);
nand NAND4 (N2371, N2367, N2149, N727, N442);
not NOT1 (N2372, N2370);
nand NAND2 (N2373, N2372, N719);
buf BUF1 (N2374, N2359);
and AND4 (N2375, N2369, N540, N1075, N809);
or OR3 (N2376, N2357, N948, N387);
or OR3 (N2377, N2347, N567, N2202);
xor XOR2 (N2378, N2376, N901);
buf BUF1 (N2379, N2371);
or OR2 (N2380, N2375, N1958);
not NOT1 (N2381, N2341);
not NOT1 (N2382, N2374);
buf BUF1 (N2383, N2380);
not NOT1 (N2384, N2350);
xor XOR2 (N2385, N2384, N1541);
nor NOR3 (N2386, N2385, N117, N95);
buf BUF1 (N2387, N2383);
buf BUF1 (N2388, N2382);
buf BUF1 (N2389, N2377);
not NOT1 (N2390, N2379);
nand NAND4 (N2391, N2373, N798, N1462, N644);
nor NOR2 (N2392, N2389, N675);
xor XOR2 (N2393, N2387, N1730);
and AND4 (N2394, N2378, N1578, N557, N139);
buf BUF1 (N2395, N2381);
nand NAND4 (N2396, N2394, N647, N1001, N2122);
xor XOR2 (N2397, N2392, N733);
not NOT1 (N2398, N2391);
and AND3 (N2399, N2397, N1597, N671);
buf BUF1 (N2400, N2395);
or OR4 (N2401, N2400, N1549, N636, N1508);
nand NAND2 (N2402, N2351, N50);
nand NAND4 (N2403, N2368, N1560, N2107, N2334);
and AND3 (N2404, N2388, N1216, N2373);
or OR3 (N2405, N2386, N122, N30);
nor NOR2 (N2406, N2402, N351);
or OR3 (N2407, N2404, N980, N1747);
nor NOR2 (N2408, N2399, N2354);
or OR2 (N2409, N2408, N1035);
not NOT1 (N2410, N2393);
or OR4 (N2411, N2409, N2317, N2240, N744);
and AND4 (N2412, N2398, N841, N931, N2024);
or OR4 (N2413, N2403, N2144, N407, N1739);
or OR3 (N2414, N2412, N426, N1168);
and AND4 (N2415, N2413, N2045, N1738, N2020);
and AND2 (N2416, N2415, N2356);
nand NAND4 (N2417, N2396, N1234, N1670, N216);
and AND3 (N2418, N2406, N1960, N163);
and AND2 (N2419, N2414, N34);
nand NAND4 (N2420, N2411, N415, N1444, N1379);
and AND2 (N2421, N2410, N126);
or OR2 (N2422, N2419, N2417);
xor XOR2 (N2423, N1670, N828);
not NOT1 (N2424, N2418);
or OR4 (N2425, N2422, N1478, N1861, N1371);
buf BUF1 (N2426, N2407);
not NOT1 (N2427, N2426);
buf BUF1 (N2428, N2405);
xor XOR2 (N2429, N2425, N182);
not NOT1 (N2430, N2420);
buf BUF1 (N2431, N2423);
or OR3 (N2432, N2416, N2242, N1592);
or OR3 (N2433, N2421, N730, N1312);
and AND4 (N2434, N2431, N106, N292, N1239);
nor NOR2 (N2435, N2424, N191);
buf BUF1 (N2436, N2401);
or OR3 (N2437, N2435, N1549, N1286);
and AND4 (N2438, N2432, N1667, N336, N980);
and AND3 (N2439, N2433, N1514, N2403);
nand NAND2 (N2440, N2390, N1755);
buf BUF1 (N2441, N2428);
buf BUF1 (N2442, N2438);
or OR2 (N2443, N2442, N751);
and AND2 (N2444, N2434, N1591);
or OR2 (N2445, N2444, N1112);
not NOT1 (N2446, N2430);
or OR4 (N2447, N2446, N2319, N499, N2007);
nor NOR3 (N2448, N2427, N366, N994);
nand NAND3 (N2449, N2445, N921, N1737);
nand NAND3 (N2450, N2443, N1412, N2066);
buf BUF1 (N2451, N2429);
xor XOR2 (N2452, N2450, N1153);
and AND2 (N2453, N2449, N1979);
or OR4 (N2454, N2451, N1411, N1312, N2257);
buf BUF1 (N2455, N2440);
or OR3 (N2456, N2437, N642, N1715);
and AND2 (N2457, N2456, N6);
nand NAND2 (N2458, N2448, N2128);
not NOT1 (N2459, N2447);
not NOT1 (N2460, N2457);
not NOT1 (N2461, N2454);
nor NOR4 (N2462, N2458, N76, N1442, N356);
not NOT1 (N2463, N2436);
buf BUF1 (N2464, N2455);
nand NAND2 (N2465, N2453, N1790);
and AND4 (N2466, N2460, N920, N896, N451);
and AND3 (N2467, N2439, N41, N1198);
or OR4 (N2468, N2462, N343, N378, N1335);
not NOT1 (N2469, N2465);
buf BUF1 (N2470, N2467);
buf BUF1 (N2471, N2464);
not NOT1 (N2472, N2459);
not NOT1 (N2473, N2471);
nand NAND4 (N2474, N2463, N1034, N656, N1164);
not NOT1 (N2475, N2468);
xor XOR2 (N2476, N2466, N2385);
nor NOR2 (N2477, N2469, N2049);
and AND2 (N2478, N2441, N315);
buf BUF1 (N2479, N2478);
and AND4 (N2480, N2477, N1012, N866, N162);
xor XOR2 (N2481, N2479, N1432);
buf BUF1 (N2482, N2461);
nand NAND2 (N2483, N2475, N500);
nor NOR2 (N2484, N2452, N1874);
and AND2 (N2485, N2483, N811);
and AND3 (N2486, N2470, N1172, N206);
nand NAND4 (N2487, N2476, N1514, N289, N450);
buf BUF1 (N2488, N2482);
not NOT1 (N2489, N2474);
buf BUF1 (N2490, N2480);
and AND2 (N2491, N2473, N2308);
not NOT1 (N2492, N2487);
not NOT1 (N2493, N2485);
nor NOR4 (N2494, N2486, N1417, N1569, N333);
buf BUF1 (N2495, N2492);
nand NAND3 (N2496, N2494, N96, N787);
buf BUF1 (N2497, N2481);
buf BUF1 (N2498, N2496);
buf BUF1 (N2499, N2490);
nor NOR4 (N2500, N2499, N2446, N876, N2031);
nand NAND3 (N2501, N2489, N1773, N2427);
and AND4 (N2502, N2495, N470, N2207, N466);
nand NAND4 (N2503, N2497, N2047, N1703, N2111);
nor NOR2 (N2504, N2484, N1406);
xor XOR2 (N2505, N2472, N261);
xor XOR2 (N2506, N2505, N385);
buf BUF1 (N2507, N2501);
nor NOR2 (N2508, N2503, N2474);
and AND4 (N2509, N2502, N520, N532, N741);
or OR2 (N2510, N2508, N1155);
and AND4 (N2511, N2504, N2066, N1855, N1914);
nand NAND3 (N2512, N2498, N922, N2198);
nand NAND2 (N2513, N2507, N2431);
nor NOR3 (N2514, N2488, N1694, N982);
and AND2 (N2515, N2511, N2030);
or OR3 (N2516, N2491, N721, N180);
buf BUF1 (N2517, N2506);
or OR2 (N2518, N2513, N476);
and AND4 (N2519, N2512, N2335, N1946, N857);
not NOT1 (N2520, N2510);
nor NOR2 (N2521, N2516, N425);
not NOT1 (N2522, N2500);
not NOT1 (N2523, N2509);
xor XOR2 (N2524, N2518, N1982);
or OR4 (N2525, N2514, N703, N942, N2505);
and AND4 (N2526, N2515, N470, N1981, N736);
not NOT1 (N2527, N2526);
nor NOR4 (N2528, N2522, N2330, N695, N509);
or OR4 (N2529, N2524, N615, N1033, N2446);
buf BUF1 (N2530, N2520);
nand NAND2 (N2531, N2523, N1201);
and AND2 (N2532, N2531, N46);
and AND3 (N2533, N2493, N268, N1689);
not NOT1 (N2534, N2517);
or OR4 (N2535, N2519, N2452, N1266, N1705);
or OR2 (N2536, N2534, N2195);
not NOT1 (N2537, N2527);
xor XOR2 (N2538, N2528, N1304);
nand NAND4 (N2539, N2538, N2372, N550, N795);
not NOT1 (N2540, N2525);
or OR4 (N2541, N2539, N2189, N665, N2005);
or OR3 (N2542, N2540, N1361, N1378);
or OR3 (N2543, N2529, N1190, N1667);
or OR4 (N2544, N2533, N664, N1626, N382);
xor XOR2 (N2545, N2543, N20);
and AND3 (N2546, N2532, N1281, N9);
xor XOR2 (N2547, N2537, N545);
nor NOR3 (N2548, N2544, N614, N795);
xor XOR2 (N2549, N2542, N379);
or OR4 (N2550, N2548, N852, N783, N2430);
buf BUF1 (N2551, N2536);
or OR2 (N2552, N2545, N1120);
and AND3 (N2553, N2550, N472, N2215);
nand NAND3 (N2554, N2541, N743, N1494);
nand NAND4 (N2555, N2521, N2292, N954, N2353);
nand NAND4 (N2556, N2549, N742, N749, N1268);
not NOT1 (N2557, N2551);
nor NOR4 (N2558, N2546, N1936, N2166, N1620);
or OR3 (N2559, N2558, N8, N1525);
and AND4 (N2560, N2535, N210, N18, N279);
nor NOR4 (N2561, N2530, N2335, N2428, N142);
nor NOR4 (N2562, N2559, N440, N1725, N389);
not NOT1 (N2563, N2560);
not NOT1 (N2564, N2553);
nand NAND4 (N2565, N2556, N132, N1819, N1727);
xor XOR2 (N2566, N2562, N287);
xor XOR2 (N2567, N2566, N732);
nor NOR2 (N2568, N2547, N2110);
nor NOR4 (N2569, N2567, N1640, N2074, N440);
not NOT1 (N2570, N2554);
and AND4 (N2571, N2564, N589, N172, N1269);
nand NAND3 (N2572, N2555, N2220, N862);
not NOT1 (N2573, N2570);
xor XOR2 (N2574, N2561, N395);
xor XOR2 (N2575, N2565, N692);
or OR3 (N2576, N2552, N186, N1587);
not NOT1 (N2577, N2573);
nand NAND2 (N2578, N2563, N653);
and AND4 (N2579, N2557, N1620, N1789, N1091);
xor XOR2 (N2580, N2571, N56);
xor XOR2 (N2581, N2572, N965);
or OR4 (N2582, N2569, N441, N2326, N609);
xor XOR2 (N2583, N2579, N2053);
nor NOR2 (N2584, N2568, N19);
buf BUF1 (N2585, N2581);
nor NOR2 (N2586, N2578, N1233);
nand NAND4 (N2587, N2576, N2380, N125, N580);
and AND3 (N2588, N2586, N843, N586);
nand NAND2 (N2589, N2577, N2359);
and AND4 (N2590, N2575, N683, N895, N89);
and AND2 (N2591, N2574, N2142);
or OR2 (N2592, N2590, N113);
buf BUF1 (N2593, N2591);
not NOT1 (N2594, N2589);
not NOT1 (N2595, N2588);
or OR2 (N2596, N2585, N833);
or OR4 (N2597, N2584, N1663, N263, N733);
not NOT1 (N2598, N2593);
buf BUF1 (N2599, N2595);
or OR3 (N2600, N2598, N2350, N140);
nor NOR3 (N2601, N2583, N2229, N1348);
nor NOR2 (N2602, N2597, N43);
xor XOR2 (N2603, N2587, N1824);
or OR2 (N2604, N2580, N429);
nand NAND3 (N2605, N2599, N2075, N773);
and AND4 (N2606, N2600, N1593, N2003, N2108);
not NOT1 (N2607, N2596);
xor XOR2 (N2608, N2603, N716);
not NOT1 (N2609, N2582);
and AND2 (N2610, N2605, N1359);
and AND3 (N2611, N2592, N2544, N663);
not NOT1 (N2612, N2601);
buf BUF1 (N2613, N2604);
nor NOR4 (N2614, N2611, N2535, N2350, N2541);
or OR3 (N2615, N2606, N2478, N1693);
xor XOR2 (N2616, N2614, N1060);
or OR2 (N2617, N2612, N1405);
buf BUF1 (N2618, N2594);
nand NAND3 (N2619, N2609, N530, N988);
xor XOR2 (N2620, N2617, N79);
and AND3 (N2621, N2619, N2189, N2291);
nor NOR2 (N2622, N2608, N2234);
buf BUF1 (N2623, N2610);
nand NAND2 (N2624, N2621, N1165);
xor XOR2 (N2625, N2622, N1347);
nor NOR4 (N2626, N2616, N1380, N1045, N695);
not NOT1 (N2627, N2602);
nor NOR3 (N2628, N2607, N443, N626);
nand NAND3 (N2629, N2626, N686, N1890);
buf BUF1 (N2630, N2623);
or OR3 (N2631, N2624, N373, N2159);
or OR2 (N2632, N2628, N130);
and AND4 (N2633, N2631, N1597, N2459, N907);
nor NOR2 (N2634, N2618, N1785);
and AND3 (N2635, N2615, N22, N1099);
xor XOR2 (N2636, N2633, N1071);
not NOT1 (N2637, N2625);
not NOT1 (N2638, N2635);
xor XOR2 (N2639, N2613, N303);
or OR2 (N2640, N2627, N1910);
xor XOR2 (N2641, N2629, N1240);
or OR2 (N2642, N2634, N666);
buf BUF1 (N2643, N2642);
nor NOR4 (N2644, N2638, N1755, N972, N457);
xor XOR2 (N2645, N2639, N1931);
and AND3 (N2646, N2632, N1998, N582);
nor NOR4 (N2647, N2644, N2117, N2020, N1103);
nand NAND4 (N2648, N2637, N1224, N2229, N517);
or OR3 (N2649, N2646, N1645, N2446);
or OR2 (N2650, N2620, N601);
and AND4 (N2651, N2647, N809, N878, N2521);
nor NOR3 (N2652, N2636, N106, N545);
buf BUF1 (N2653, N2645);
and AND3 (N2654, N2651, N851, N1963);
buf BUF1 (N2655, N2643);
xor XOR2 (N2656, N2641, N2241);
buf BUF1 (N2657, N2650);
not NOT1 (N2658, N2648);
nor NOR3 (N2659, N2652, N1187, N1271);
buf BUF1 (N2660, N2658);
nand NAND3 (N2661, N2653, N2513, N1357);
or OR2 (N2662, N2649, N806);
buf BUF1 (N2663, N2661);
buf BUF1 (N2664, N2654);
xor XOR2 (N2665, N2660, N1665);
buf BUF1 (N2666, N2657);
or OR2 (N2667, N2664, N1787);
nand NAND4 (N2668, N2630, N1893, N838, N1595);
buf BUF1 (N2669, N2662);
nand NAND3 (N2670, N2655, N391, N1683);
nand NAND2 (N2671, N2666, N1466);
nand NAND4 (N2672, N2671, N1538, N1763, N1921);
xor XOR2 (N2673, N2668, N1493);
or OR4 (N2674, N2663, N377, N464, N1469);
not NOT1 (N2675, N2667);
xor XOR2 (N2676, N2659, N364);
nor NOR3 (N2677, N2670, N1273, N141);
not NOT1 (N2678, N2676);
buf BUF1 (N2679, N2675);
or OR2 (N2680, N2665, N359);
nand NAND3 (N2681, N2640, N2011, N2545);
nor NOR4 (N2682, N2681, N442, N2497, N2096);
and AND2 (N2683, N2656, N1567);
and AND4 (N2684, N2673, N1712, N1692, N1316);
xor XOR2 (N2685, N2669, N2209);
buf BUF1 (N2686, N2672);
nor NOR2 (N2687, N2674, N1798);
not NOT1 (N2688, N2677);
nand NAND4 (N2689, N2684, N1362, N2539, N2432);
not NOT1 (N2690, N2687);
nor NOR3 (N2691, N2686, N2555, N2117);
or OR4 (N2692, N2682, N1484, N943, N1653);
xor XOR2 (N2693, N2678, N1349);
xor XOR2 (N2694, N2691, N233);
nand NAND4 (N2695, N2683, N1642, N1521, N857);
not NOT1 (N2696, N2685);
or OR2 (N2697, N2692, N848);
or OR2 (N2698, N2693, N51);
nand NAND2 (N2699, N2697, N1358);
buf BUF1 (N2700, N2690);
nor NOR3 (N2701, N2695, N2611, N695);
not NOT1 (N2702, N2694);
nor NOR2 (N2703, N2701, N1343);
not NOT1 (N2704, N2679);
not NOT1 (N2705, N2680);
not NOT1 (N2706, N2699);
and AND2 (N2707, N2698, N463);
nor NOR4 (N2708, N2704, N2482, N945, N2704);
not NOT1 (N2709, N2708);
nor NOR4 (N2710, N2700, N489, N1865, N1684);
and AND3 (N2711, N2688, N2707, N1727);
and AND2 (N2712, N1409, N2229);
not NOT1 (N2713, N2702);
and AND3 (N2714, N2712, N1584, N814);
and AND3 (N2715, N2706, N2191, N2673);
not NOT1 (N2716, N2713);
or OR2 (N2717, N2715, N1903);
buf BUF1 (N2718, N2716);
or OR3 (N2719, N2714, N1438, N28);
xor XOR2 (N2720, N2718, N83);
nor NOR3 (N2721, N2696, N2596, N2532);
or OR2 (N2722, N2689, N1054);
not NOT1 (N2723, N2711);
buf BUF1 (N2724, N2705);
not NOT1 (N2725, N2709);
or OR4 (N2726, N2717, N2207, N1124, N1698);
xor XOR2 (N2727, N2725, N1640);
xor XOR2 (N2728, N2721, N2209);
and AND3 (N2729, N2722, N998, N2638);
xor XOR2 (N2730, N2729, N2033);
nand NAND4 (N2731, N2703, N2536, N2149, N2065);
nand NAND3 (N2732, N2720, N1127, N426);
nand NAND2 (N2733, N2728, N585);
nor NOR4 (N2734, N2731, N1791, N1869, N2154);
not NOT1 (N2735, N2733);
and AND3 (N2736, N2732, N1620, N844);
not NOT1 (N2737, N2730);
nand NAND2 (N2738, N2735, N441);
and AND3 (N2739, N2710, N2721, N623);
not NOT1 (N2740, N2738);
nor NOR3 (N2741, N2740, N2373, N699);
nor NOR2 (N2742, N2726, N2350);
nand NAND2 (N2743, N2736, N2424);
not NOT1 (N2744, N2741);
not NOT1 (N2745, N2727);
and AND2 (N2746, N2745, N1656);
nor NOR2 (N2747, N2737, N2041);
buf BUF1 (N2748, N2743);
nand NAND4 (N2749, N2742, N2219, N390, N907);
or OR4 (N2750, N2744, N647, N2241, N2120);
not NOT1 (N2751, N2739);
or OR2 (N2752, N2723, N61);
not NOT1 (N2753, N2749);
and AND3 (N2754, N2753, N2472, N2310);
or OR2 (N2755, N2750, N2257);
nor NOR4 (N2756, N2752, N157, N171, N1584);
and AND3 (N2757, N2734, N1156, N1791);
and AND2 (N2758, N2751, N1026);
buf BUF1 (N2759, N2756);
or OR3 (N2760, N2755, N2049, N119);
nor NOR4 (N2761, N2746, N163, N184, N612);
not NOT1 (N2762, N2747);
nand NAND4 (N2763, N2719, N61, N827, N2440);
not NOT1 (N2764, N2760);
xor XOR2 (N2765, N2759, N290);
buf BUF1 (N2766, N2762);
xor XOR2 (N2767, N2761, N1263);
xor XOR2 (N2768, N2748, N2689);
buf BUF1 (N2769, N2763);
not NOT1 (N2770, N2724);
not NOT1 (N2771, N2758);
not NOT1 (N2772, N2769);
nand NAND4 (N2773, N2757, N1672, N838, N738);
xor XOR2 (N2774, N2770, N480);
buf BUF1 (N2775, N2766);
nor NOR3 (N2776, N2768, N232, N2765);
not NOT1 (N2777, N2295);
nor NOR4 (N2778, N2775, N2237, N77, N427);
nor NOR4 (N2779, N2771, N765, N433, N419);
and AND2 (N2780, N2778, N2403);
nor NOR3 (N2781, N2779, N1794, N2433);
not NOT1 (N2782, N2767);
buf BUF1 (N2783, N2780);
nand NAND3 (N2784, N2782, N786, N2302);
or OR4 (N2785, N2764, N2385, N2106, N1283);
nor NOR3 (N2786, N2785, N321, N2062);
or OR3 (N2787, N2774, N656, N913);
nand NAND2 (N2788, N2787, N1842);
or OR3 (N2789, N2788, N749, N93);
buf BUF1 (N2790, N2777);
nand NAND3 (N2791, N2783, N2148, N2657);
nand NAND3 (N2792, N2786, N2724, N1100);
or OR3 (N2793, N2781, N1173, N1157);
and AND3 (N2794, N2773, N1923, N856);
nand NAND4 (N2795, N2784, N1974, N1642, N298);
nand NAND3 (N2796, N2794, N1749, N505);
or OR2 (N2797, N2795, N2644);
not NOT1 (N2798, N2793);
or OR3 (N2799, N2796, N2702, N2684);
or OR3 (N2800, N2791, N817, N2258);
or OR4 (N2801, N2789, N1557, N1457, N2628);
buf BUF1 (N2802, N2799);
nor NOR3 (N2803, N2797, N2596, N1282);
not NOT1 (N2804, N2798);
not NOT1 (N2805, N2754);
or OR4 (N2806, N2801, N1191, N274, N1745);
xor XOR2 (N2807, N2792, N413);
and AND3 (N2808, N2802, N327, N2542);
not NOT1 (N2809, N2804);
xor XOR2 (N2810, N2790, N261);
nor NOR2 (N2811, N2805, N2218);
nand NAND2 (N2812, N2810, N2810);
and AND4 (N2813, N2807, N2352, N2045, N2442);
not NOT1 (N2814, N2776);
or OR3 (N2815, N2800, N1535, N1099);
buf BUF1 (N2816, N2808);
xor XOR2 (N2817, N2814, N1251);
buf BUF1 (N2818, N2772);
nand NAND4 (N2819, N2815, N1435, N421, N2704);
buf BUF1 (N2820, N2813);
nand NAND4 (N2821, N2803, N570, N1058, N332);
or OR3 (N2822, N2819, N2209, N1462);
not NOT1 (N2823, N2812);
buf BUF1 (N2824, N2809);
not NOT1 (N2825, N2806);
buf BUF1 (N2826, N2822);
or OR4 (N2827, N2811, N395, N5, N699);
not NOT1 (N2828, N2824);
nor NOR4 (N2829, N2821, N901, N1902, N116);
and AND4 (N2830, N2818, N2699, N2500, N403);
buf BUF1 (N2831, N2823);
and AND3 (N2832, N2820, N2563, N148);
nand NAND2 (N2833, N2827, N2665);
xor XOR2 (N2834, N2816, N651);
or OR2 (N2835, N2830, N566);
nand NAND4 (N2836, N2828, N732, N2266, N1559);
or OR3 (N2837, N2834, N2122, N2025);
nor NOR3 (N2838, N2837, N2693, N279);
not NOT1 (N2839, N2831);
nor NOR2 (N2840, N2817, N567);
nand NAND2 (N2841, N2836, N2526);
xor XOR2 (N2842, N2825, N2497);
and AND2 (N2843, N2833, N1452);
nand NAND2 (N2844, N2832, N2399);
xor XOR2 (N2845, N2840, N1190);
nor NOR3 (N2846, N2841, N2809, N2422);
or OR3 (N2847, N2846, N462, N2725);
nor NOR3 (N2848, N2839, N933, N1598);
buf BUF1 (N2849, N2845);
nor NOR2 (N2850, N2848, N337);
nand NAND3 (N2851, N2849, N580, N610);
and AND3 (N2852, N2838, N374, N2338);
xor XOR2 (N2853, N2835, N2322);
and AND2 (N2854, N2844, N725);
buf BUF1 (N2855, N2854);
nor NOR2 (N2856, N2853, N2600);
nor NOR3 (N2857, N2855, N356, N1821);
nor NOR4 (N2858, N2843, N2696, N1223, N632);
nand NAND3 (N2859, N2856, N2401, N626);
not NOT1 (N2860, N2850);
nand NAND2 (N2861, N2860, N2699);
xor XOR2 (N2862, N2852, N800);
not NOT1 (N2863, N2862);
xor XOR2 (N2864, N2847, N2529);
xor XOR2 (N2865, N2857, N1880);
or OR4 (N2866, N2864, N2467, N2207, N65);
buf BUF1 (N2867, N2861);
or OR4 (N2868, N2826, N1641, N2707, N2343);
and AND2 (N2869, N2863, N1036);
nand NAND4 (N2870, N2865, N40, N1508, N1671);
xor XOR2 (N2871, N2842, N1364);
buf BUF1 (N2872, N2866);
not NOT1 (N2873, N2867);
and AND4 (N2874, N2871, N2013, N389, N507);
or OR4 (N2875, N2858, N890, N2466, N1257);
buf BUF1 (N2876, N2874);
nor NOR3 (N2877, N2872, N2212, N2374);
nor NOR3 (N2878, N2868, N2294, N2551);
buf BUF1 (N2879, N2851);
xor XOR2 (N2880, N2875, N2156);
not NOT1 (N2881, N2829);
or OR3 (N2882, N2881, N1358, N2812);
and AND4 (N2883, N2869, N1150, N1746, N2154);
not NOT1 (N2884, N2870);
nand NAND4 (N2885, N2882, N1006, N2646, N2019);
or OR3 (N2886, N2880, N1944, N2372);
buf BUF1 (N2887, N2876);
xor XOR2 (N2888, N2885, N2780);
and AND4 (N2889, N2873, N1551, N721, N420);
not NOT1 (N2890, N2886);
buf BUF1 (N2891, N2884);
nand NAND3 (N2892, N2891, N2825, N2533);
not NOT1 (N2893, N2888);
buf BUF1 (N2894, N2893);
and AND3 (N2895, N2883, N210, N637);
or OR3 (N2896, N2879, N173, N2376);
nor NOR3 (N2897, N2877, N199, N449);
or OR2 (N2898, N2859, N440);
not NOT1 (N2899, N2878);
and AND4 (N2900, N2887, N313, N1703, N2723);
and AND4 (N2901, N2898, N2407, N963, N672);
or OR2 (N2902, N2895, N441);
and AND2 (N2903, N2900, N120);
not NOT1 (N2904, N2896);
not NOT1 (N2905, N2894);
buf BUF1 (N2906, N2902);
nand NAND2 (N2907, N2905, N1813);
not NOT1 (N2908, N2889);
buf BUF1 (N2909, N2899);
nor NOR3 (N2910, N2892, N1434, N2492);
and AND4 (N2911, N2890, N2005, N2391, N2061);
and AND2 (N2912, N2903, N665);
buf BUF1 (N2913, N2912);
nor NOR3 (N2914, N2913, N1906, N2070);
nor NOR2 (N2915, N2908, N390);
nand NAND4 (N2916, N2901, N1000, N144, N2839);
nor NOR4 (N2917, N2915, N1872, N86, N905);
or OR3 (N2918, N2906, N2317, N222);
nand NAND2 (N2919, N2916, N2363);
xor XOR2 (N2920, N2918, N1177);
nand NAND2 (N2921, N2914, N1154);
buf BUF1 (N2922, N2907);
or OR3 (N2923, N2920, N695, N208);
nor NOR2 (N2924, N2904, N2129);
nand NAND2 (N2925, N2917, N2108);
nor NOR2 (N2926, N2909, N1388);
buf BUF1 (N2927, N2911);
not NOT1 (N2928, N2924);
buf BUF1 (N2929, N2897);
buf BUF1 (N2930, N2919);
not NOT1 (N2931, N2928);
and AND4 (N2932, N2923, N1244, N1493, N990);
buf BUF1 (N2933, N2922);
not NOT1 (N2934, N2910);
nand NAND4 (N2935, N2932, N81, N124, N1894);
xor XOR2 (N2936, N2925, N800);
nand NAND4 (N2937, N2921, N1868, N1219, N396);
nand NAND3 (N2938, N2926, N1117, N415);
and AND4 (N2939, N2931, N2407, N428, N1853);
not NOT1 (N2940, N2939);
nand NAND4 (N2941, N2927, N236, N1377, N21);
and AND2 (N2942, N2929, N688);
or OR2 (N2943, N2933, N933);
and AND3 (N2944, N2940, N2360, N2035);
nor NOR2 (N2945, N2941, N1153);
buf BUF1 (N2946, N2943);
nand NAND3 (N2947, N2935, N2665, N2781);
or OR4 (N2948, N2936, N1443, N1492, N2026);
buf BUF1 (N2949, N2948);
or OR3 (N2950, N2944, N628, N43);
buf BUF1 (N2951, N2950);
nor NOR3 (N2952, N2945, N1524, N218);
nand NAND3 (N2953, N2938, N518, N2873);
and AND4 (N2954, N2942, N1849, N1627, N2259);
buf BUF1 (N2955, N2934);
xor XOR2 (N2956, N2955, N1965);
not NOT1 (N2957, N2953);
or OR3 (N2958, N2954, N2684, N2573);
nand NAND3 (N2959, N2937, N1041, N1129);
and AND4 (N2960, N2951, N215, N2020, N80);
buf BUF1 (N2961, N2960);
and AND2 (N2962, N2959, N2341);
xor XOR2 (N2963, N2947, N1139);
nor NOR4 (N2964, N2961, N1888, N796, N1349);
nand NAND4 (N2965, N2952, N2160, N1293, N662);
nor NOR2 (N2966, N2949, N483);
and AND4 (N2967, N2963, N2596, N110, N2190);
nand NAND4 (N2968, N2957, N2864, N2365, N2355);
or OR2 (N2969, N2968, N2960);
nor NOR2 (N2970, N2966, N930);
or OR4 (N2971, N2930, N962, N2226, N1045);
buf BUF1 (N2972, N2958);
nand NAND4 (N2973, N2967, N2676, N1009, N2893);
and AND3 (N2974, N2970, N1576, N745);
not NOT1 (N2975, N2969);
buf BUF1 (N2976, N2974);
nor NOR4 (N2977, N2973, N527, N2237, N716);
and AND4 (N2978, N2971, N1782, N1263, N36);
xor XOR2 (N2979, N2964, N1203);
buf BUF1 (N2980, N2972);
buf BUF1 (N2981, N2975);
xor XOR2 (N2982, N2981, N2444);
not NOT1 (N2983, N2956);
buf BUF1 (N2984, N2982);
and AND2 (N2985, N2979, N1758);
or OR2 (N2986, N2946, N1838);
nor NOR2 (N2987, N2986, N2306);
or OR2 (N2988, N2976, N2835);
not NOT1 (N2989, N2984);
not NOT1 (N2990, N2988);
xor XOR2 (N2991, N2985, N2830);
not NOT1 (N2992, N2991);
nor NOR2 (N2993, N2983, N562);
xor XOR2 (N2994, N2992, N614);
nor NOR3 (N2995, N2993, N1893, N911);
nand NAND3 (N2996, N2987, N2208, N200);
not NOT1 (N2997, N2996);
not NOT1 (N2998, N2990);
xor XOR2 (N2999, N2997, N2318);
nand NAND4 (N3000, N2962, N1614, N1212, N1477);
xor XOR2 (N3001, N2977, N1042);
and AND3 (N3002, N2998, N2478, N2820);
nor NOR4 (N3003, N2989, N2386, N2381, N2435);
nor NOR2 (N3004, N2980, N375);
xor XOR2 (N3005, N3004, N2072);
not NOT1 (N3006, N2994);
nand NAND4 (N3007, N2999, N1549, N2853, N1314);
nor NOR2 (N3008, N2995, N1137);
nand NAND2 (N3009, N3006, N1360);
nor NOR3 (N3010, N2965, N1487, N2918);
buf BUF1 (N3011, N3001);
not NOT1 (N3012, N3011);
and AND4 (N3013, N3010, N1384, N639, N2088);
nor NOR2 (N3014, N3008, N2346);
nand NAND3 (N3015, N3013, N2810, N1337);
or OR2 (N3016, N2978, N1632);
not NOT1 (N3017, N3002);
nor NOR4 (N3018, N3007, N701, N1913, N2638);
xor XOR2 (N3019, N3005, N2493);
nor NOR2 (N3020, N3012, N1447);
and AND4 (N3021, N3020, N2645, N2597, N1591);
buf BUF1 (N3022, N3003);
not NOT1 (N3023, N3000);
xor XOR2 (N3024, N3019, N1161);
nor NOR2 (N3025, N3018, N1789);
nor NOR4 (N3026, N3024, N2161, N2702, N47);
and AND4 (N3027, N3009, N937, N2932, N1023);
buf BUF1 (N3028, N3025);
and AND2 (N3029, N3017, N2460);
or OR3 (N3030, N3028, N593, N1261);
nor NOR3 (N3031, N3016, N326, N606);
xor XOR2 (N3032, N3031, N1135);
buf BUF1 (N3033, N3015);
and AND2 (N3034, N3033, N2277);
not NOT1 (N3035, N3014);
nor NOR4 (N3036, N3022, N1753, N172, N2153);
nor NOR4 (N3037, N3034, N2737, N2649, N866);
buf BUF1 (N3038, N3030);
not NOT1 (N3039, N3029);
nand NAND2 (N3040, N3037, N2361);
xor XOR2 (N3041, N3032, N778);
not NOT1 (N3042, N3026);
nor NOR4 (N3043, N3039, N1656, N1201, N1839);
and AND3 (N3044, N3043, N1655, N1633);
nand NAND3 (N3045, N3023, N1797, N2077);
nand NAND4 (N3046, N3044, N2712, N1368, N6);
xor XOR2 (N3047, N3036, N1249);
nand NAND2 (N3048, N3041, N1358);
not NOT1 (N3049, N3047);
buf BUF1 (N3050, N3038);
buf BUF1 (N3051, N3021);
or OR2 (N3052, N3046, N2594);
buf BUF1 (N3053, N3050);
buf BUF1 (N3054, N3042);
buf BUF1 (N3055, N3051);
or OR4 (N3056, N3045, N723, N803, N2621);
nor NOR4 (N3057, N3056, N2956, N1982, N2214);
buf BUF1 (N3058, N3048);
nand NAND2 (N3059, N3054, N2419);
xor XOR2 (N3060, N3058, N2786);
buf BUF1 (N3061, N3060);
nor NOR4 (N3062, N3055, N197, N354, N712);
or OR2 (N3063, N3053, N566);
nand NAND4 (N3064, N3063, N1115, N169, N1034);
and AND2 (N3065, N3062, N967);
or OR4 (N3066, N3061, N511, N572, N2372);
and AND3 (N3067, N3064, N1183, N1667);
buf BUF1 (N3068, N3057);
buf BUF1 (N3069, N3067);
and AND4 (N3070, N3065, N2846, N1299, N136);
nand NAND4 (N3071, N3070, N418, N3066, N1455);
buf BUF1 (N3072, N392);
and AND4 (N3073, N3059, N2164, N1909, N69);
xor XOR2 (N3074, N3072, N92);
nor NOR2 (N3075, N3069, N1279);
xor XOR2 (N3076, N3073, N1666);
xor XOR2 (N3077, N3049, N1174);
nand NAND3 (N3078, N3075, N347, N378);
nand NAND4 (N3079, N3052, N653, N764, N1946);
xor XOR2 (N3080, N3040, N2626);
and AND4 (N3081, N3080, N2338, N624, N1147);
nor NOR3 (N3082, N3078, N2538, N2814);
and AND3 (N3083, N3076, N1586, N1035);
and AND4 (N3084, N3071, N1090, N2995, N1909);
not NOT1 (N3085, N3084);
nor NOR4 (N3086, N3077, N2032, N1841, N1069);
nand NAND2 (N3087, N3086, N2135);
or OR2 (N3088, N3079, N2639);
or OR4 (N3089, N3087, N1674, N2378, N1410);
nor NOR2 (N3090, N3074, N2347);
buf BUF1 (N3091, N3082);
xor XOR2 (N3092, N3027, N503);
xor XOR2 (N3093, N3081, N902);
and AND4 (N3094, N3083, N142, N321, N2254);
xor XOR2 (N3095, N3090, N1916);
xor XOR2 (N3096, N3068, N752);
not NOT1 (N3097, N3093);
xor XOR2 (N3098, N3088, N575);
or OR3 (N3099, N3091, N2630, N665);
nand NAND3 (N3100, N3035, N1357, N940);
nor NOR4 (N3101, N3100, N1572, N2690, N2483);
and AND2 (N3102, N3096, N2041);
buf BUF1 (N3103, N3094);
or OR2 (N3104, N3099, N1768);
nor NOR4 (N3105, N3085, N962, N12, N2835);
nor NOR3 (N3106, N3105, N1029, N2996);
nand NAND4 (N3107, N3106, N39, N2993, N2721);
buf BUF1 (N3108, N3101);
xor XOR2 (N3109, N3107, N2284);
xor XOR2 (N3110, N3095, N2123);
nand NAND3 (N3111, N3097, N441, N2811);
buf BUF1 (N3112, N3089);
and AND3 (N3113, N3112, N612, N1474);
not NOT1 (N3114, N3110);
and AND2 (N3115, N3109, N689);
xor XOR2 (N3116, N3114, N2237);
or OR4 (N3117, N3098, N1774, N2151, N490);
not NOT1 (N3118, N3117);
nand NAND3 (N3119, N3118, N2567, N2098);
nand NAND3 (N3120, N3103, N1220, N2617);
nor NOR3 (N3121, N3092, N1783, N1658);
and AND4 (N3122, N3116, N2252, N1423, N338);
buf BUF1 (N3123, N3120);
or OR2 (N3124, N3108, N2094);
xor XOR2 (N3125, N3122, N958);
not NOT1 (N3126, N3104);
buf BUF1 (N3127, N3125);
xor XOR2 (N3128, N3102, N1264);
or OR4 (N3129, N3127, N399, N485, N2703);
buf BUF1 (N3130, N3128);
buf BUF1 (N3131, N3119);
nor NOR4 (N3132, N3111, N2004, N1816, N921);
nand NAND2 (N3133, N3126, N1003);
not NOT1 (N3134, N3124);
or OR3 (N3135, N3131, N2119, N792);
not NOT1 (N3136, N3113);
and AND3 (N3137, N3130, N2253, N763);
or OR3 (N3138, N3123, N1268, N2418);
or OR3 (N3139, N3121, N2623, N1547);
not NOT1 (N3140, N3137);
nand NAND4 (N3141, N3132, N1962, N639, N1438);
not NOT1 (N3142, N3134);
not NOT1 (N3143, N3135);
not NOT1 (N3144, N3129);
nand NAND4 (N3145, N3139, N2871, N2788, N2444);
nand NAND2 (N3146, N3141, N959);
buf BUF1 (N3147, N3115);
nand NAND3 (N3148, N3136, N1960, N172);
nor NOR2 (N3149, N3146, N3097);
buf BUF1 (N3150, N3147);
buf BUF1 (N3151, N3145);
nor NOR3 (N3152, N3140, N2025, N2133);
nand NAND4 (N3153, N3133, N1398, N1556, N1494);
nand NAND4 (N3154, N3153, N97, N510, N432);
or OR4 (N3155, N3143, N1379, N1565, N807);
buf BUF1 (N3156, N3151);
buf BUF1 (N3157, N3152);
nor NOR3 (N3158, N3155, N1711, N1416);
not NOT1 (N3159, N3142);
nand NAND2 (N3160, N3158, N281);
nor NOR4 (N3161, N3149, N2397, N2401, N2979);
or OR4 (N3162, N3159, N2046, N736, N14);
or OR2 (N3163, N3138, N3136);
not NOT1 (N3164, N3162);
and AND2 (N3165, N3144, N1211);
not NOT1 (N3166, N3148);
xor XOR2 (N3167, N3165, N608);
or OR3 (N3168, N3167, N2160, N244);
not NOT1 (N3169, N3150);
not NOT1 (N3170, N3166);
and AND4 (N3171, N3169, N1265, N1945, N2370);
nand NAND3 (N3172, N3156, N2327, N400);
xor XOR2 (N3173, N3163, N2550);
or OR3 (N3174, N3154, N2109, N535);
and AND3 (N3175, N3164, N1611, N1900);
buf BUF1 (N3176, N3168);
and AND2 (N3177, N3170, N2057);
not NOT1 (N3178, N3160);
or OR4 (N3179, N3171, N1209, N1240, N135);
nand NAND2 (N3180, N3176, N1033);
buf BUF1 (N3181, N3179);
xor XOR2 (N3182, N3178, N677);
and AND2 (N3183, N3172, N1158);
not NOT1 (N3184, N3173);
not NOT1 (N3185, N3174);
xor XOR2 (N3186, N3183, N1951);
or OR2 (N3187, N3184, N580);
or OR2 (N3188, N3175, N1348);
buf BUF1 (N3189, N3187);
buf BUF1 (N3190, N3157);
xor XOR2 (N3191, N3180, N2092);
and AND4 (N3192, N3189, N698, N392, N179);
not NOT1 (N3193, N3190);
and AND2 (N3194, N3193, N294);
nand NAND4 (N3195, N3177, N1314, N2542, N1964);
or OR2 (N3196, N3194, N82);
buf BUF1 (N3197, N3186);
or OR3 (N3198, N3182, N2344, N2848);
nand NAND4 (N3199, N3188, N2038, N1382, N2850);
buf BUF1 (N3200, N3199);
buf BUF1 (N3201, N3195);
or OR2 (N3202, N3196, N2937);
and AND2 (N3203, N3201, N1722);
or OR4 (N3204, N3197, N2110, N92, N3137);
nor NOR3 (N3205, N3185, N1113, N984);
and AND2 (N3206, N3203, N2084);
not NOT1 (N3207, N3191);
or OR3 (N3208, N3192, N1143, N1674);
buf BUF1 (N3209, N3205);
or OR2 (N3210, N3208, N2094);
nand NAND2 (N3211, N3204, N1852);
buf BUF1 (N3212, N3161);
buf BUF1 (N3213, N3198);
not NOT1 (N3214, N3211);
or OR2 (N3215, N3207, N856);
nor NOR4 (N3216, N3200, N1941, N1113, N218);
nand NAND3 (N3217, N3216, N1564, N1516);
nor NOR4 (N3218, N3215, N1391, N613, N3144);
not NOT1 (N3219, N3214);
not NOT1 (N3220, N3181);
xor XOR2 (N3221, N3218, N483);
nor NOR3 (N3222, N3209, N1585, N781);
nand NAND4 (N3223, N3221, N1875, N2906, N887);
buf BUF1 (N3224, N3219);
buf BUF1 (N3225, N3224);
buf BUF1 (N3226, N3222);
nor NOR2 (N3227, N3210, N806);
xor XOR2 (N3228, N3225, N378);
and AND3 (N3229, N3223, N2224, N2331);
xor XOR2 (N3230, N3213, N1653);
not NOT1 (N3231, N3228);
or OR3 (N3232, N3212, N479, N411);
xor XOR2 (N3233, N3232, N2865);
nor NOR4 (N3234, N3206, N1934, N3119, N2135);
and AND3 (N3235, N3229, N3183, N114);
buf BUF1 (N3236, N3202);
nand NAND2 (N3237, N3227, N2789);
nand NAND4 (N3238, N3226, N3067, N208, N3090);
nor NOR4 (N3239, N3220, N2710, N478, N1940);
and AND2 (N3240, N3239, N1095);
and AND2 (N3241, N3230, N266);
buf BUF1 (N3242, N3237);
nor NOR2 (N3243, N3231, N2825);
nor NOR2 (N3244, N3241, N2407);
not NOT1 (N3245, N3235);
xor XOR2 (N3246, N3245, N2197);
or OR3 (N3247, N3243, N2737, N143);
nand NAND3 (N3248, N3242, N3094, N2010);
xor XOR2 (N3249, N3247, N1479);
nor NOR2 (N3250, N3233, N2384);
nor NOR4 (N3251, N3240, N2371, N3114, N2829);
or OR2 (N3252, N3249, N1571);
not NOT1 (N3253, N3238);
buf BUF1 (N3254, N3217);
or OR2 (N3255, N3251, N2735);
nand NAND2 (N3256, N3252, N615);
nand NAND3 (N3257, N3234, N2865, N5);
xor XOR2 (N3258, N3255, N2948);
nand NAND3 (N3259, N3257, N1784, N2517);
not NOT1 (N3260, N3246);
nand NAND2 (N3261, N3248, N1566);
nor NOR4 (N3262, N3260, N753, N1057, N1408);
not NOT1 (N3263, N3258);
nand NAND4 (N3264, N3261, N2601, N2327, N202);
not NOT1 (N3265, N3236);
not NOT1 (N3266, N3256);
xor XOR2 (N3267, N3264, N893);
not NOT1 (N3268, N3266);
xor XOR2 (N3269, N3253, N2178);
buf BUF1 (N3270, N3254);
buf BUF1 (N3271, N3269);
xor XOR2 (N3272, N3244, N3225);
nand NAND2 (N3273, N3267, N3123);
and AND2 (N3274, N3272, N931);
not NOT1 (N3275, N3271);
not NOT1 (N3276, N3259);
buf BUF1 (N3277, N3262);
or OR2 (N3278, N3250, N1490);
and AND3 (N3279, N3268, N2759, N738);
or OR4 (N3280, N3270, N143, N1842, N17);
and AND2 (N3281, N3277, N2893);
xor XOR2 (N3282, N3278, N1745);
nand NAND4 (N3283, N3273, N2622, N2017, N1424);
nor NOR3 (N3284, N3282, N1159, N897);
nand NAND2 (N3285, N3283, N2308);
nand NAND2 (N3286, N3281, N1165);
nor NOR4 (N3287, N3284, N1375, N1635, N2122);
not NOT1 (N3288, N3263);
nand NAND2 (N3289, N3265, N2080);
xor XOR2 (N3290, N3288, N1912);
nand NAND4 (N3291, N3290, N500, N1790, N773);
nor NOR4 (N3292, N3279, N2348, N2513, N1959);
xor XOR2 (N3293, N3289, N1849);
xor XOR2 (N3294, N3286, N588);
nor NOR4 (N3295, N3275, N2025, N2592, N1519);
nor NOR4 (N3296, N3274, N1096, N2764, N1447);
buf BUF1 (N3297, N3292);
and AND2 (N3298, N3295, N327);
nand NAND3 (N3299, N3276, N2980, N354);
not NOT1 (N3300, N3294);
xor XOR2 (N3301, N3297, N2308);
buf BUF1 (N3302, N3291);
and AND4 (N3303, N3280, N3091, N550, N2218);
not NOT1 (N3304, N3300);
or OR2 (N3305, N3302, N2082);
xor XOR2 (N3306, N3303, N1873);
buf BUF1 (N3307, N3306);
nand NAND2 (N3308, N3285, N3014);
nor NOR4 (N3309, N3308, N2473, N577, N2889);
or OR3 (N3310, N3299, N2502, N2987);
nor NOR3 (N3311, N3310, N2217, N2682);
nand NAND2 (N3312, N3293, N1843);
xor XOR2 (N3313, N3312, N1811);
and AND2 (N3314, N3301, N1112);
or OR4 (N3315, N3314, N1401, N939, N2956);
not NOT1 (N3316, N3304);
not NOT1 (N3317, N3309);
nor NOR3 (N3318, N3298, N389, N1264);
xor XOR2 (N3319, N3287, N1828);
or OR3 (N3320, N3319, N3183, N3138);
xor XOR2 (N3321, N3305, N1328);
not NOT1 (N3322, N3320);
or OR4 (N3323, N3296, N1612, N1464, N1195);
xor XOR2 (N3324, N3316, N2538);
not NOT1 (N3325, N3311);
nand NAND4 (N3326, N3318, N3131, N1177, N193);
and AND2 (N3327, N3313, N1189);
xor XOR2 (N3328, N3325, N1575);
or OR3 (N3329, N3324, N2990, N423);
nand NAND4 (N3330, N3326, N2730, N117, N125);
nor NOR2 (N3331, N3327, N2151);
and AND2 (N3332, N3315, N1845);
nand NAND4 (N3333, N3323, N1632, N1024, N1370);
xor XOR2 (N3334, N3328, N2918);
xor XOR2 (N3335, N3307, N1060);
buf BUF1 (N3336, N3331);
nor NOR4 (N3337, N3317, N1399, N2255, N2758);
and AND3 (N3338, N3322, N1655, N1574);
nor NOR2 (N3339, N3334, N9);
nand NAND4 (N3340, N3329, N2441, N795, N609);
nand NAND2 (N3341, N3330, N536);
not NOT1 (N3342, N3337);
not NOT1 (N3343, N3333);
and AND4 (N3344, N3340, N1399, N736, N1366);
nor NOR3 (N3345, N3321, N1443, N2619);
buf BUF1 (N3346, N3336);
buf BUF1 (N3347, N3335);
and AND4 (N3348, N3346, N815, N2813, N1672);
nor NOR4 (N3349, N3339, N1068, N908, N464);
and AND4 (N3350, N3332, N1240, N3336, N2469);
and AND3 (N3351, N3347, N2926, N1663);
buf BUF1 (N3352, N3350);
nand NAND3 (N3353, N3349, N3298, N1893);
not NOT1 (N3354, N3342);
buf BUF1 (N3355, N3344);
not NOT1 (N3356, N3351);
and AND2 (N3357, N3343, N1579);
buf BUF1 (N3358, N3352);
nand NAND2 (N3359, N3345, N806);
and AND2 (N3360, N3358, N2524);
not NOT1 (N3361, N3357);
nand NAND3 (N3362, N3360, N2260, N3176);
xor XOR2 (N3363, N3356, N1172);
nor NOR2 (N3364, N3363, N1752);
xor XOR2 (N3365, N3341, N2464);
nor NOR2 (N3366, N3338, N691);
or OR2 (N3367, N3364, N2917);
or OR3 (N3368, N3348, N813, N1421);
nand NAND3 (N3369, N3367, N1486, N1605);
xor XOR2 (N3370, N3368, N2178);
buf BUF1 (N3371, N3370);
nor NOR2 (N3372, N3354, N1896);
or OR3 (N3373, N3366, N1679, N434);
not NOT1 (N3374, N3371);
nand NAND2 (N3375, N3361, N3131);
and AND2 (N3376, N3375, N1806);
xor XOR2 (N3377, N3374, N2834);
nor NOR3 (N3378, N3373, N1033, N1582);
nand NAND2 (N3379, N3353, N1663);
or OR4 (N3380, N3376, N2410, N2612, N2997);
nand NAND3 (N3381, N3379, N2073, N3201);
buf BUF1 (N3382, N3362);
not NOT1 (N3383, N3377);
or OR3 (N3384, N3381, N2727, N557);
and AND3 (N3385, N3359, N2444, N1296);
nand NAND2 (N3386, N3382, N3311);
nor NOR4 (N3387, N3365, N2135, N1952, N3150);
xor XOR2 (N3388, N3380, N3002);
nand NAND3 (N3389, N3384, N3192, N711);
or OR3 (N3390, N3385, N296, N2517);
or OR2 (N3391, N3389, N2069);
nor NOR2 (N3392, N3378, N440);
not NOT1 (N3393, N3388);
or OR3 (N3394, N3393, N2766, N2694);
nor NOR4 (N3395, N3394, N1806, N1972, N2477);
nor NOR2 (N3396, N3387, N2239);
nor NOR4 (N3397, N3372, N761, N2414, N177);
or OR3 (N3398, N3383, N1286, N793);
or OR4 (N3399, N3397, N2999, N2174, N728);
or OR4 (N3400, N3398, N2646, N2366, N3377);
or OR2 (N3401, N3355, N528);
buf BUF1 (N3402, N3401);
and AND3 (N3403, N3395, N800, N1223);
buf BUF1 (N3404, N3386);
and AND4 (N3405, N3396, N778, N2892, N2928);
nor NOR2 (N3406, N3391, N1271);
not NOT1 (N3407, N3403);
and AND2 (N3408, N3400, N1373);
not NOT1 (N3409, N3407);
and AND2 (N3410, N3369, N2459);
or OR3 (N3411, N3399, N1269, N3265);
not NOT1 (N3412, N3402);
buf BUF1 (N3413, N3411);
nand NAND4 (N3414, N3390, N1165, N703, N3075);
xor XOR2 (N3415, N3408, N1346);
or OR4 (N3416, N3392, N2778, N3387, N599);
not NOT1 (N3417, N3409);
and AND4 (N3418, N3417, N332, N2417, N1717);
buf BUF1 (N3419, N3413);
and AND4 (N3420, N3416, N2922, N275, N798);
or OR2 (N3421, N3420, N3411);
nor NOR2 (N3422, N3410, N860);
and AND4 (N3423, N3418, N2848, N2474, N3106);
or OR2 (N3424, N3423, N1366);
nand NAND3 (N3425, N3415, N2256, N3189);
buf BUF1 (N3426, N3404);
buf BUF1 (N3427, N3406);
nand NAND3 (N3428, N3419, N3342, N2096);
not NOT1 (N3429, N3421);
not NOT1 (N3430, N3405);
and AND3 (N3431, N3414, N2176, N517);
not NOT1 (N3432, N3427);
buf BUF1 (N3433, N3429);
nor NOR4 (N3434, N3422, N1534, N3262, N1278);
xor XOR2 (N3435, N3433, N3226);
xor XOR2 (N3436, N3431, N2674);
or OR3 (N3437, N3428, N2814, N2253);
xor XOR2 (N3438, N3430, N3412);
or OR2 (N3439, N2289, N2090);
nor NOR2 (N3440, N3437, N3405);
or OR2 (N3441, N3439, N579);
not NOT1 (N3442, N3441);
or OR2 (N3443, N3436, N113);
and AND4 (N3444, N3434, N2580, N3065, N1948);
buf BUF1 (N3445, N3432);
buf BUF1 (N3446, N3442);
and AND2 (N3447, N3444, N269);
xor XOR2 (N3448, N3446, N596);
and AND3 (N3449, N3425, N2607, N1298);
and AND3 (N3450, N3447, N3358, N1469);
nor NOR2 (N3451, N3448, N1938);
or OR2 (N3452, N3426, N1149);
nor NOR3 (N3453, N3438, N1458, N760);
buf BUF1 (N3454, N3440);
or OR3 (N3455, N3452, N904, N728);
or OR3 (N3456, N3424, N2945, N938);
nor NOR3 (N3457, N3450, N2189, N3181);
nor NOR4 (N3458, N3453, N197, N1804, N929);
buf BUF1 (N3459, N3455);
nor NOR3 (N3460, N3443, N1939, N2080);
nor NOR4 (N3461, N3460, N2410, N3219, N2786);
xor XOR2 (N3462, N3457, N2766);
and AND4 (N3463, N3461, N1771, N1844, N777);
buf BUF1 (N3464, N3445);
nand NAND4 (N3465, N3462, N1687, N1188, N3370);
xor XOR2 (N3466, N3465, N1097);
xor XOR2 (N3467, N3435, N2288);
nor NOR3 (N3468, N3463, N1538, N3205);
or OR2 (N3469, N3458, N1473);
or OR2 (N3470, N3459, N1626);
and AND3 (N3471, N3466, N1564, N1187);
xor XOR2 (N3472, N3468, N2764);
xor XOR2 (N3473, N3469, N1436);
or OR2 (N3474, N3470, N2715);
and AND3 (N3475, N3454, N2487, N1821);
xor XOR2 (N3476, N3451, N2157);
xor XOR2 (N3477, N3456, N1471);
and AND4 (N3478, N3472, N2740, N1376, N1622);
and AND4 (N3479, N3471, N2175, N745, N616);
buf BUF1 (N3480, N3476);
nor NOR3 (N3481, N3449, N1905, N2812);
nand NAND3 (N3482, N3475, N2204, N551);
xor XOR2 (N3483, N3481, N2174);
xor XOR2 (N3484, N3479, N1818);
or OR3 (N3485, N3464, N2864, N766);
or OR3 (N3486, N3478, N144, N221);
buf BUF1 (N3487, N3482);
buf BUF1 (N3488, N3483);
nand NAND3 (N3489, N3488, N489, N1024);
not NOT1 (N3490, N3480);
nor NOR2 (N3491, N3490, N105);
buf BUF1 (N3492, N3491);
nand NAND2 (N3493, N3492, N1153);
xor XOR2 (N3494, N3485, N1191);
or OR3 (N3495, N3486, N2235, N1250);
or OR4 (N3496, N3473, N2247, N2400, N581);
nor NOR4 (N3497, N3493, N2714, N3062, N1885);
not NOT1 (N3498, N3477);
xor XOR2 (N3499, N3494, N2762);
buf BUF1 (N3500, N3467);
xor XOR2 (N3501, N3497, N1135);
not NOT1 (N3502, N3499);
nand NAND3 (N3503, N3489, N601, N3298);
nor NOR2 (N3504, N3503, N2993);
nor NOR2 (N3505, N3504, N2659);
buf BUF1 (N3506, N3474);
and AND2 (N3507, N3502, N1632);
or OR2 (N3508, N3500, N2601);
and AND2 (N3509, N3498, N2584);
not NOT1 (N3510, N3501);
not NOT1 (N3511, N3495);
nand NAND2 (N3512, N3487, N245);
or OR2 (N3513, N3507, N668);
and AND3 (N3514, N3484, N1653, N3166);
nor NOR3 (N3515, N3505, N2228, N653);
xor XOR2 (N3516, N3512, N2223);
not NOT1 (N3517, N3515);
and AND2 (N3518, N3509, N747);
nand NAND3 (N3519, N3518, N2455, N2048);
or OR4 (N3520, N3517, N2326, N346, N1562);
nand NAND3 (N3521, N3510, N2090, N1999);
xor XOR2 (N3522, N3506, N2310);
xor XOR2 (N3523, N3508, N948);
buf BUF1 (N3524, N3513);
buf BUF1 (N3525, N3523);
buf BUF1 (N3526, N3524);
and AND4 (N3527, N3521, N1008, N531, N149);
nor NOR3 (N3528, N3516, N1401, N2567);
and AND3 (N3529, N3514, N668, N1946);
not NOT1 (N3530, N3526);
nor NOR2 (N3531, N3530, N913);
nor NOR2 (N3532, N3531, N3164);
xor XOR2 (N3533, N3511, N862);
or OR3 (N3534, N3525, N1894, N495);
and AND2 (N3535, N3532, N3081);
and AND3 (N3536, N3529, N1229, N3448);
xor XOR2 (N3537, N3520, N22);
xor XOR2 (N3538, N3533, N1153);
xor XOR2 (N3539, N3527, N1458);
not NOT1 (N3540, N3536);
nor NOR3 (N3541, N3522, N2219, N861);
or OR4 (N3542, N3539, N3217, N3021, N2009);
nor NOR4 (N3543, N3496, N852, N2252, N1288);
and AND4 (N3544, N3543, N16, N3438, N2770);
nor NOR2 (N3545, N3542, N1849);
and AND4 (N3546, N3544, N2936, N521, N443);
nor NOR3 (N3547, N3537, N1319, N243);
not NOT1 (N3548, N3541);
nor NOR2 (N3549, N3545, N3519);
xor XOR2 (N3550, N3220, N3385);
not NOT1 (N3551, N3548);
nand NAND2 (N3552, N3547, N2213);
buf BUF1 (N3553, N3534);
not NOT1 (N3554, N3546);
not NOT1 (N3555, N3551);
nor NOR2 (N3556, N3552, N2015);
nor NOR2 (N3557, N3550, N3143);
nand NAND3 (N3558, N3555, N1566, N1512);
or OR3 (N3559, N3553, N511, N2075);
buf BUF1 (N3560, N3559);
xor XOR2 (N3561, N3560, N2445);
not NOT1 (N3562, N3549);
not NOT1 (N3563, N3558);
buf BUF1 (N3564, N3538);
or OR2 (N3565, N3535, N1020);
xor XOR2 (N3566, N3554, N1619);
xor XOR2 (N3567, N3528, N953);
nand NAND3 (N3568, N3557, N1708, N2300);
not NOT1 (N3569, N3568);
nand NAND4 (N3570, N3564, N922, N1534, N1759);
or OR4 (N3571, N3556, N3111, N586, N3534);
not NOT1 (N3572, N3566);
buf BUF1 (N3573, N3567);
xor XOR2 (N3574, N3563, N3190);
xor XOR2 (N3575, N3572, N331);
xor XOR2 (N3576, N3573, N947);
xor XOR2 (N3577, N3540, N1496);
buf BUF1 (N3578, N3575);
xor XOR2 (N3579, N3574, N2066);
buf BUF1 (N3580, N3577);
nor NOR2 (N3581, N3562, N2849);
nor NOR4 (N3582, N3565, N3501, N2539, N3325);
or OR2 (N3583, N3579, N257);
buf BUF1 (N3584, N3576);
buf BUF1 (N3585, N3570);
buf BUF1 (N3586, N3561);
and AND2 (N3587, N3581, N2816);
nor NOR2 (N3588, N3578, N2271);
buf BUF1 (N3589, N3586);
not NOT1 (N3590, N3587);
xor XOR2 (N3591, N3585, N1255);
buf BUF1 (N3592, N3584);
buf BUF1 (N3593, N3589);
nor NOR3 (N3594, N3571, N193, N3402);
buf BUF1 (N3595, N3590);
not NOT1 (N3596, N3588);
or OR4 (N3597, N3582, N2703, N158, N3101);
nor NOR3 (N3598, N3592, N1430, N3556);
and AND2 (N3599, N3597, N2905);
and AND3 (N3600, N3599, N3103, N2354);
nor NOR4 (N3601, N3598, N1761, N678, N1959);
nand NAND2 (N3602, N3580, N2486);
nand NAND3 (N3603, N3591, N3075, N2502);
xor XOR2 (N3604, N3601, N2229);
buf BUF1 (N3605, N3602);
buf BUF1 (N3606, N3604);
xor XOR2 (N3607, N3603, N1479);
xor XOR2 (N3608, N3596, N3184);
or OR3 (N3609, N3595, N388, N3331);
nand NAND2 (N3610, N3583, N3526);
buf BUF1 (N3611, N3609);
nand NAND4 (N3612, N3600, N207, N1738, N1412);
nand NAND2 (N3613, N3608, N2761);
xor XOR2 (N3614, N3610, N3499);
buf BUF1 (N3615, N3614);
nand NAND4 (N3616, N3611, N299, N3136, N3239);
and AND3 (N3617, N3616, N66, N1462);
nor NOR2 (N3618, N3569, N2905);
or OR3 (N3619, N3594, N3069, N2871);
nor NOR2 (N3620, N3593, N2245);
nor NOR3 (N3621, N3620, N2560, N1286);
xor XOR2 (N3622, N3613, N880);
or OR2 (N3623, N3606, N46);
and AND3 (N3624, N3621, N409, N791);
xor XOR2 (N3625, N3622, N2874);
and AND4 (N3626, N3605, N1185, N2681, N3195);
or OR4 (N3627, N3625, N2525, N2525, N264);
buf BUF1 (N3628, N3615);
not NOT1 (N3629, N3607);
not NOT1 (N3630, N3612);
nand NAND3 (N3631, N3628, N2632, N2555);
or OR2 (N3632, N3629, N1466);
and AND4 (N3633, N3624, N550, N140, N3586);
nand NAND3 (N3634, N3630, N2319, N2750);
xor XOR2 (N3635, N3633, N2617);
xor XOR2 (N3636, N3626, N3333);
nand NAND2 (N3637, N3617, N2785);
and AND4 (N3638, N3636, N329, N2903, N2254);
or OR2 (N3639, N3631, N373);
not NOT1 (N3640, N3637);
not NOT1 (N3641, N3640);
and AND2 (N3642, N3627, N650);
nor NOR2 (N3643, N3618, N2962);
xor XOR2 (N3644, N3634, N2730);
buf BUF1 (N3645, N3632);
xor XOR2 (N3646, N3644, N534);
nor NOR4 (N3647, N3623, N1946, N996, N483);
nor NOR3 (N3648, N3635, N2644, N1134);
xor XOR2 (N3649, N3642, N3506);
and AND3 (N3650, N3619, N1436, N1746);
xor XOR2 (N3651, N3646, N2520);
nor NOR4 (N3652, N3638, N1312, N2592, N817);
xor XOR2 (N3653, N3650, N3633);
not NOT1 (N3654, N3652);
and AND4 (N3655, N3654, N895, N676, N1477);
xor XOR2 (N3656, N3641, N303);
not NOT1 (N3657, N3648);
nand NAND4 (N3658, N3655, N585, N318, N818);
xor XOR2 (N3659, N3653, N3633);
nand NAND2 (N3660, N3658, N2554);
nand NAND3 (N3661, N3656, N336, N11);
nand NAND2 (N3662, N3659, N3472);
nand NAND2 (N3663, N3651, N1132);
nand NAND2 (N3664, N3657, N2998);
nor NOR2 (N3665, N3639, N1830);
or OR4 (N3666, N3664, N442, N519, N610);
not NOT1 (N3667, N3647);
nand NAND3 (N3668, N3665, N194, N1657);
not NOT1 (N3669, N3660);
nand NAND3 (N3670, N3649, N1272, N1052);
xor XOR2 (N3671, N3667, N3600);
buf BUF1 (N3672, N3661);
not NOT1 (N3673, N3643);
nor NOR2 (N3674, N3673, N2881);
xor XOR2 (N3675, N3645, N3632);
not NOT1 (N3676, N3666);
nor NOR3 (N3677, N3669, N2952, N1058);
not NOT1 (N3678, N3672);
or OR2 (N3679, N3677, N1641);
not NOT1 (N3680, N3670);
not NOT1 (N3681, N3674);
buf BUF1 (N3682, N3681);
or OR4 (N3683, N3662, N95, N2453, N588);
nand NAND2 (N3684, N3668, N1123);
xor XOR2 (N3685, N3671, N3011);
and AND3 (N3686, N3685, N3163, N1762);
not NOT1 (N3687, N3676);
not NOT1 (N3688, N3683);
xor XOR2 (N3689, N3663, N3134);
or OR2 (N3690, N3678, N3106);
and AND2 (N3691, N3675, N686);
xor XOR2 (N3692, N3691, N2731);
buf BUF1 (N3693, N3692);
and AND4 (N3694, N3687, N2935, N1118, N1563);
nand NAND3 (N3695, N3684, N1850, N506);
or OR2 (N3696, N3689, N922);
nand NAND3 (N3697, N3694, N161, N891);
or OR2 (N3698, N3679, N995);
and AND4 (N3699, N3690, N3445, N2509, N1518);
or OR3 (N3700, N3697, N2915, N3390);
buf BUF1 (N3701, N3696);
xor XOR2 (N3702, N3699, N2621);
buf BUF1 (N3703, N3701);
nand NAND3 (N3704, N3682, N864, N1262);
xor XOR2 (N3705, N3702, N58);
nor NOR4 (N3706, N3698, N1995, N1021, N340);
nand NAND4 (N3707, N3704, N646, N2116, N3339);
not NOT1 (N3708, N3707);
xor XOR2 (N3709, N3693, N1268);
nor NOR4 (N3710, N3700, N318, N907, N3345);
or OR4 (N3711, N3695, N1862, N2516, N588);
xor XOR2 (N3712, N3680, N2893);
or OR4 (N3713, N3712, N1223, N659, N2026);
buf BUF1 (N3714, N3705);
nand NAND2 (N3715, N3711, N2464);
or OR4 (N3716, N3709, N1897, N3507, N1738);
nor NOR3 (N3717, N3688, N195, N1203);
nand NAND4 (N3718, N3717, N3327, N1959, N3584);
nand NAND4 (N3719, N3714, N590, N3088, N685);
not NOT1 (N3720, N3708);
xor XOR2 (N3721, N3715, N1473);
buf BUF1 (N3722, N3721);
nor NOR4 (N3723, N3718, N2017, N2317, N833);
or OR4 (N3724, N3716, N2720, N3484, N408);
nor NOR3 (N3725, N3703, N3420, N2103);
or OR3 (N3726, N3722, N1060, N3570);
not NOT1 (N3727, N3725);
nand NAND2 (N3728, N3726, N3168);
buf BUF1 (N3729, N3723);
nor NOR3 (N3730, N3713, N2031, N1125);
buf BUF1 (N3731, N3686);
nand NAND2 (N3732, N3720, N2835);
xor XOR2 (N3733, N3719, N2736);
nor NOR3 (N3734, N3732, N1969, N430);
xor XOR2 (N3735, N3710, N3257);
not NOT1 (N3736, N3727);
nand NAND3 (N3737, N3706, N2874, N372);
and AND4 (N3738, N3731, N1101, N1250, N1372);
nor NOR3 (N3739, N3729, N2430, N2216);
xor XOR2 (N3740, N3735, N1015);
and AND2 (N3741, N3740, N2132);
not NOT1 (N3742, N3738);
xor XOR2 (N3743, N3739, N1867);
nor NOR4 (N3744, N3733, N1949, N34, N3317);
xor XOR2 (N3745, N3730, N3288);
or OR4 (N3746, N3741, N355, N1635, N2777);
xor XOR2 (N3747, N3734, N406);
nand NAND3 (N3748, N3745, N2218, N1928);
and AND3 (N3749, N3728, N2726, N2001);
xor XOR2 (N3750, N3724, N2081);
nand NAND3 (N3751, N3746, N1111, N1283);
nor NOR2 (N3752, N3744, N2338);
not NOT1 (N3753, N3743);
not NOT1 (N3754, N3749);
and AND4 (N3755, N3751, N796, N481, N3474);
not NOT1 (N3756, N3755);
or OR3 (N3757, N3753, N739, N3673);
nand NAND2 (N3758, N3754, N1855);
not NOT1 (N3759, N3757);
nand NAND2 (N3760, N3759, N578);
nand NAND3 (N3761, N3737, N590, N2262);
not NOT1 (N3762, N3760);
nand NAND3 (N3763, N3761, N2330, N814);
nand NAND2 (N3764, N3748, N2529);
and AND3 (N3765, N3758, N1658, N1482);
xor XOR2 (N3766, N3764, N404);
nor NOR4 (N3767, N3765, N2319, N1813, N3533);
or OR2 (N3768, N3736, N817);
buf BUF1 (N3769, N3752);
and AND4 (N3770, N3756, N1583, N568, N2461);
nand NAND3 (N3771, N3763, N1485, N3019);
buf BUF1 (N3772, N3747);
buf BUF1 (N3773, N3750);
or OR3 (N3774, N3742, N452, N675);
xor XOR2 (N3775, N3762, N2786);
buf BUF1 (N3776, N3766);
not NOT1 (N3777, N3770);
and AND3 (N3778, N3771, N682, N1199);
or OR4 (N3779, N3767, N1331, N3093, N212);
nand NAND2 (N3780, N3769, N1655);
and AND3 (N3781, N3776, N3020, N2127);
nand NAND2 (N3782, N3777, N2526);
or OR3 (N3783, N3773, N2588, N870);
and AND2 (N3784, N3778, N1195);
buf BUF1 (N3785, N3775);
nor NOR3 (N3786, N3781, N3405, N164);
not NOT1 (N3787, N3782);
nand NAND3 (N3788, N3786, N1376, N1753);
nor NOR3 (N3789, N3768, N2017, N2805);
nor NOR4 (N3790, N3779, N1337, N3594, N1353);
or OR2 (N3791, N3787, N2009);
and AND2 (N3792, N3791, N3494);
buf BUF1 (N3793, N3785);
and AND4 (N3794, N3783, N2170, N262, N1687);
nand NAND4 (N3795, N3794, N1699, N2451, N3435);
buf BUF1 (N3796, N3788);
nand NAND4 (N3797, N3793, N633, N3381, N3071);
or OR4 (N3798, N3784, N1773, N3699, N1249);
and AND3 (N3799, N3796, N3160, N2506);
or OR2 (N3800, N3789, N2567);
xor XOR2 (N3801, N3798, N947);
nand NAND4 (N3802, N3797, N1380, N1472, N3782);
buf BUF1 (N3803, N3772);
nand NAND2 (N3804, N3803, N518);
nor NOR3 (N3805, N3800, N1422, N1515);
not NOT1 (N3806, N3802);
not NOT1 (N3807, N3804);
nand NAND3 (N3808, N3805, N1017, N2470);
and AND2 (N3809, N3790, N1564);
and AND2 (N3810, N3780, N1920);
xor XOR2 (N3811, N3801, N2598);
nand NAND3 (N3812, N3795, N2753, N2519);
nand NAND3 (N3813, N3810, N3692, N2704);
not NOT1 (N3814, N3774);
xor XOR2 (N3815, N3812, N140);
xor XOR2 (N3816, N3809, N2305);
and AND3 (N3817, N3815, N3270, N3010);
buf BUF1 (N3818, N3799);
or OR3 (N3819, N3816, N2254, N3613);
buf BUF1 (N3820, N3806);
nand NAND4 (N3821, N3813, N1143, N594, N473);
and AND4 (N3822, N3818, N636, N653, N2607);
and AND2 (N3823, N3822, N3759);
buf BUF1 (N3824, N3823);
not NOT1 (N3825, N3819);
nor NOR4 (N3826, N3824, N2876, N156, N396);
buf BUF1 (N3827, N3821);
buf BUF1 (N3828, N3807);
nand NAND4 (N3829, N3814, N1025, N2133, N1211);
or OR4 (N3830, N3808, N912, N3525, N1217);
nor NOR2 (N3831, N3829, N1672);
buf BUF1 (N3832, N3825);
buf BUF1 (N3833, N3832);
not NOT1 (N3834, N3831);
buf BUF1 (N3835, N3834);
not NOT1 (N3836, N3792);
nand NAND4 (N3837, N3828, N752, N1068, N3819);
nor NOR3 (N3838, N3820, N2578, N2714);
nand NAND2 (N3839, N3835, N3113);
nor NOR4 (N3840, N3826, N3150, N1201, N2559);
nor NOR3 (N3841, N3827, N1938, N1123);
not NOT1 (N3842, N3840);
xor XOR2 (N3843, N3842, N102);
buf BUF1 (N3844, N3836);
or OR3 (N3845, N3843, N1153, N278);
not NOT1 (N3846, N3817);
or OR3 (N3847, N3838, N711, N1981);
or OR4 (N3848, N3847, N2109, N2218, N387);
nand NAND3 (N3849, N3811, N2586, N1445);
nor NOR4 (N3850, N3837, N2303, N1274, N1875);
buf BUF1 (N3851, N3848);
or OR3 (N3852, N3850, N1556, N3308);
xor XOR2 (N3853, N3830, N215);
or OR3 (N3854, N3849, N2751, N1363);
buf BUF1 (N3855, N3854);
and AND3 (N3856, N3845, N253, N1423);
or OR2 (N3857, N3841, N1312);
buf BUF1 (N3858, N3852);
not NOT1 (N3859, N3853);
xor XOR2 (N3860, N3833, N661);
not NOT1 (N3861, N3855);
buf BUF1 (N3862, N3839);
nand NAND2 (N3863, N3846, N462);
nor NOR3 (N3864, N3860, N1026, N1769);
nor NOR2 (N3865, N3856, N3501);
nand NAND2 (N3866, N3865, N2757);
buf BUF1 (N3867, N3844);
and AND2 (N3868, N3858, N2808);
nor NOR2 (N3869, N3862, N2982);
not NOT1 (N3870, N3861);
nor NOR4 (N3871, N3867, N1460, N848, N3394);
or OR3 (N3872, N3863, N1656, N2864);
xor XOR2 (N3873, N3857, N2746);
xor XOR2 (N3874, N3869, N2576);
buf BUF1 (N3875, N3874);
buf BUF1 (N3876, N3871);
xor XOR2 (N3877, N3851, N2064);
and AND3 (N3878, N3872, N1818, N277);
or OR2 (N3879, N3868, N989);
buf BUF1 (N3880, N3864);
or OR3 (N3881, N3875, N3700, N2382);
buf BUF1 (N3882, N3866);
nand NAND3 (N3883, N3882, N2928, N2279);
or OR4 (N3884, N3878, N2230, N3366, N2590);
xor XOR2 (N3885, N3870, N2010);
or OR3 (N3886, N3859, N1667, N1559);
and AND4 (N3887, N3886, N3522, N3331, N2564);
nor NOR3 (N3888, N3887, N394, N43);
buf BUF1 (N3889, N3873);
xor XOR2 (N3890, N3889, N3477);
nand NAND3 (N3891, N3883, N2789, N3783);
or OR4 (N3892, N3877, N3296, N2449, N460);
xor XOR2 (N3893, N3891, N736);
nor NOR4 (N3894, N3893, N3717, N407, N1760);
and AND4 (N3895, N3876, N914, N3264, N142);
not NOT1 (N3896, N3895);
nand NAND3 (N3897, N3881, N257, N2052);
and AND4 (N3898, N3890, N2447, N3659, N2517);
and AND3 (N3899, N3898, N2184, N1511);
and AND4 (N3900, N3884, N2558, N24, N1057);
nand NAND4 (N3901, N3897, N1570, N3016, N2132);
xor XOR2 (N3902, N3892, N3469);
not NOT1 (N3903, N3899);
xor XOR2 (N3904, N3888, N1946);
nand NAND2 (N3905, N3885, N2928);
not NOT1 (N3906, N3902);
xor XOR2 (N3907, N3894, N3616);
not NOT1 (N3908, N3879);
nand NAND2 (N3909, N3901, N2088);
nand NAND4 (N3910, N3880, N2324, N1326, N3171);
and AND4 (N3911, N3900, N3185, N2974, N1597);
and AND4 (N3912, N3907, N3601, N35, N2055);
nand NAND2 (N3913, N3896, N1254);
buf BUF1 (N3914, N3905);
xor XOR2 (N3915, N3910, N2379);
or OR4 (N3916, N3911, N3309, N3456, N2138);
buf BUF1 (N3917, N3909);
or OR2 (N3918, N3915, N824);
not NOT1 (N3919, N3913);
xor XOR2 (N3920, N3903, N875);
xor XOR2 (N3921, N3916, N1404);
or OR3 (N3922, N3912, N1888, N3588);
xor XOR2 (N3923, N3906, N1610);
buf BUF1 (N3924, N3908);
nand NAND3 (N3925, N3904, N3130, N3227);
xor XOR2 (N3926, N3919, N1050);
or OR2 (N3927, N3918, N91);
or OR2 (N3928, N3917, N848);
nor NOR4 (N3929, N3924, N409, N1122, N3470);
nor NOR3 (N3930, N3928, N2342, N1975);
not NOT1 (N3931, N3920);
xor XOR2 (N3932, N3930, N746);
nand NAND2 (N3933, N3929, N315);
xor XOR2 (N3934, N3923, N3435);
not NOT1 (N3935, N3921);
nor NOR2 (N3936, N3926, N3243);
xor XOR2 (N3937, N3935, N3803);
nand NAND2 (N3938, N3934, N474);
or OR2 (N3939, N3937, N1527);
nand NAND4 (N3940, N3914, N1187, N1857, N2603);
and AND2 (N3941, N3927, N1411);
not NOT1 (N3942, N3938);
not NOT1 (N3943, N3922);
nand NAND4 (N3944, N3940, N3605, N2204, N80);
xor XOR2 (N3945, N3931, N1412);
nand NAND2 (N3946, N3945, N3757);
xor XOR2 (N3947, N3944, N948);
not NOT1 (N3948, N3925);
or OR4 (N3949, N3942, N2330, N2382, N722);
or OR3 (N3950, N3932, N1872, N2173);
nor NOR2 (N3951, N3950, N3834);
buf BUF1 (N3952, N3933);
nand NAND4 (N3953, N3951, N2133, N71, N1368);
nand NAND4 (N3954, N3936, N437, N3435, N528);
nand NAND4 (N3955, N3954, N2699, N2740, N2505);
or OR4 (N3956, N3955, N772, N3134, N16);
not NOT1 (N3957, N3949);
buf BUF1 (N3958, N3939);
not NOT1 (N3959, N3946);
not NOT1 (N3960, N3952);
and AND2 (N3961, N3948, N789);
buf BUF1 (N3962, N3947);
nor NOR3 (N3963, N3962, N166, N1986);
xor XOR2 (N3964, N3959, N3358);
nand NAND2 (N3965, N3960, N3055);
nand NAND3 (N3966, N3956, N2503, N1951);
or OR2 (N3967, N3957, N3931);
nand NAND3 (N3968, N3967, N3931, N1669);
buf BUF1 (N3969, N3968);
nand NAND3 (N3970, N3943, N295, N2185);
and AND2 (N3971, N3941, N888);
nand NAND4 (N3972, N3963, N3565, N2434, N1931);
and AND2 (N3973, N3971, N1512);
nand NAND4 (N3974, N3972, N1327, N361, N2583);
and AND4 (N3975, N3966, N1236, N3559, N777);
nor NOR3 (N3976, N3975, N862, N3449);
or OR4 (N3977, N3976, N1429, N696, N2068);
xor XOR2 (N3978, N3953, N2721);
not NOT1 (N3979, N3974);
nand NAND2 (N3980, N3965, N3220);
and AND4 (N3981, N3958, N1789, N3530, N1728);
not NOT1 (N3982, N3970);
or OR4 (N3983, N3978, N1798, N919, N2562);
nand NAND2 (N3984, N3982, N2382);
or OR4 (N3985, N3980, N2724, N2896, N1918);
xor XOR2 (N3986, N3969, N1360);
nand NAND3 (N3987, N3986, N603, N424);
and AND4 (N3988, N3985, N325, N3716, N3226);
or OR3 (N3989, N3983, N2094, N3578);
nor NOR2 (N3990, N3964, N3487);
buf BUF1 (N3991, N3989);
and AND3 (N3992, N3988, N586, N714);
xor XOR2 (N3993, N3973, N2633);
xor XOR2 (N3994, N3992, N2957);
and AND4 (N3995, N3984, N2555, N2874, N2010);
not NOT1 (N3996, N3987);
nor NOR4 (N3997, N3995, N485, N3347, N800);
xor XOR2 (N3998, N3961, N2780);
xor XOR2 (N3999, N3977, N1741);
nand NAND2 (N4000, N3991, N681);
xor XOR2 (N4001, N3999, N1205);
not NOT1 (N4002, N3994);
and AND3 (N4003, N4002, N1377, N2631);
nand NAND4 (N4004, N3996, N3959, N1543, N1757);
nor NOR4 (N4005, N3997, N454, N1590, N2545);
and AND2 (N4006, N3981, N2407);
buf BUF1 (N4007, N4005);
not NOT1 (N4008, N3990);
not NOT1 (N4009, N4000);
or OR3 (N4010, N4008, N1724, N3071);
nand NAND2 (N4011, N4009, N1493);
or OR2 (N4012, N4007, N1607);
not NOT1 (N4013, N4006);
xor XOR2 (N4014, N4010, N3660);
nand NAND2 (N4015, N4011, N2398);
or OR2 (N4016, N4014, N1545);
nor NOR2 (N4017, N4013, N1722);
buf BUF1 (N4018, N3993);
or OR4 (N4019, N4004, N3873, N2337, N2495);
and AND4 (N4020, N4003, N3643, N3812, N3968);
buf BUF1 (N4021, N4016);
xor XOR2 (N4022, N4019, N3606);
or OR3 (N4023, N4021, N3659, N2361);
and AND2 (N4024, N3998, N1096);
xor XOR2 (N4025, N3979, N1439);
nor NOR4 (N4026, N4018, N1039, N1636, N1350);
and AND2 (N4027, N4026, N425);
nor NOR2 (N4028, N4020, N392);
not NOT1 (N4029, N4015);
and AND2 (N4030, N4012, N355);
not NOT1 (N4031, N4022);
or OR4 (N4032, N4028, N2810, N2914, N2567);
xor XOR2 (N4033, N4024, N28);
xor XOR2 (N4034, N4030, N1427);
buf BUF1 (N4035, N4027);
not NOT1 (N4036, N4017);
buf BUF1 (N4037, N4031);
xor XOR2 (N4038, N4023, N3183);
buf BUF1 (N4039, N4033);
and AND3 (N4040, N4025, N2034, N2445);
or OR4 (N4041, N4036, N754, N1020, N183);
and AND4 (N4042, N4040, N970, N962, N3695);
nor NOR2 (N4043, N4001, N2013);
nand NAND4 (N4044, N4037, N2081, N886, N4035);
or OR4 (N4045, N3539, N3798, N1467, N2647);
and AND3 (N4046, N4034, N2743, N1046);
not NOT1 (N4047, N4046);
xor XOR2 (N4048, N4038, N1202);
nand NAND4 (N4049, N4047, N3440, N3886, N2385);
or OR4 (N4050, N4045, N2783, N428, N2284);
or OR4 (N4051, N4049, N2912, N3471, N4032);
nand NAND2 (N4052, N1261, N1234);
buf BUF1 (N4053, N4048);
and AND2 (N4054, N4053, N376);
and AND4 (N4055, N4039, N1820, N2871, N3520);
buf BUF1 (N4056, N4051);
xor XOR2 (N4057, N4054, N784);
nor NOR3 (N4058, N4044, N2263, N1410);
xor XOR2 (N4059, N4058, N3335);
xor XOR2 (N4060, N4029, N594);
buf BUF1 (N4061, N4041);
buf BUF1 (N4062, N4056);
not NOT1 (N4063, N4055);
xor XOR2 (N4064, N4042, N2600);
nand NAND3 (N4065, N4061, N496, N2609);
xor XOR2 (N4066, N4062, N2866);
or OR3 (N4067, N4057, N2175, N2030);
or OR4 (N4068, N4065, N3201, N2342, N1023);
xor XOR2 (N4069, N4060, N2447);
xor XOR2 (N4070, N4063, N2950);
xor XOR2 (N4071, N4050, N3455);
nor NOR4 (N4072, N4069, N885, N53, N3588);
nor NOR4 (N4073, N4071, N2724, N109, N2114);
xor XOR2 (N4074, N4067, N3299);
buf BUF1 (N4075, N4070);
nand NAND2 (N4076, N4066, N3612);
buf BUF1 (N4077, N4074);
nand NAND4 (N4078, N4076, N3286, N2531, N3100);
and AND4 (N4079, N4075, N3641, N2058, N1492);
not NOT1 (N4080, N4064);
buf BUF1 (N4081, N4059);
not NOT1 (N4082, N4080);
nand NAND4 (N4083, N4077, N1588, N295, N1783);
nor NOR3 (N4084, N4052, N1279, N87);
nor NOR4 (N4085, N4079, N3874, N3009, N3210);
and AND2 (N4086, N4073, N3887);
nand NAND4 (N4087, N4083, N1760, N1500, N2182);
nor NOR4 (N4088, N4068, N964, N1268, N1337);
not NOT1 (N4089, N4082);
buf BUF1 (N4090, N4072);
not NOT1 (N4091, N4084);
not NOT1 (N4092, N4078);
xor XOR2 (N4093, N4043, N3788);
xor XOR2 (N4094, N4081, N844);
not NOT1 (N4095, N4090);
nand NAND2 (N4096, N4086, N2955);
or OR4 (N4097, N4091, N1496, N3371, N3324);
or OR4 (N4098, N4097, N650, N2070, N2040);
not NOT1 (N4099, N4098);
not NOT1 (N4100, N4087);
not NOT1 (N4101, N4088);
xor XOR2 (N4102, N4101, N3409);
xor XOR2 (N4103, N4094, N1765);
nor NOR4 (N4104, N4099, N1004, N368, N228);
or OR3 (N4105, N4096, N1984, N1720);
not NOT1 (N4106, N4095);
and AND3 (N4107, N4092, N114, N3206);
and AND3 (N4108, N4089, N4015, N1203);
nor NOR3 (N4109, N4103, N2200, N1934);
xor XOR2 (N4110, N4104, N3538);
not NOT1 (N4111, N4100);
nor NOR4 (N4112, N4106, N315, N1653, N3067);
and AND4 (N4113, N4093, N2196, N3410, N1764);
not NOT1 (N4114, N4113);
not NOT1 (N4115, N4102);
and AND2 (N4116, N4115, N2870);
not NOT1 (N4117, N4109);
nor NOR4 (N4118, N4108, N1860, N781, N937);
nand NAND3 (N4119, N4107, N2073, N56);
not NOT1 (N4120, N4111);
nor NOR3 (N4121, N4114, N3348, N457);
xor XOR2 (N4122, N4120, N398);
or OR4 (N4123, N4122, N10, N2742, N2539);
and AND4 (N4124, N4118, N2175, N1256, N1146);
or OR2 (N4125, N4105, N3461);
and AND3 (N4126, N4124, N1314, N2635);
nand NAND3 (N4127, N4116, N1425, N1117);
nor NOR2 (N4128, N4125, N1184);
or OR2 (N4129, N4085, N917);
or OR2 (N4130, N4117, N956);
or OR3 (N4131, N4127, N3684, N4110);
nand NAND3 (N4132, N4110, N2125, N3552);
or OR3 (N4133, N4129, N737, N12);
and AND2 (N4134, N4133, N4030);
and AND3 (N4135, N4134, N1661, N3138);
xor XOR2 (N4136, N4119, N564);
nand NAND2 (N4137, N4121, N536);
and AND4 (N4138, N4123, N1311, N1397, N3968);
and AND3 (N4139, N4126, N3072, N481);
not NOT1 (N4140, N4112);
not NOT1 (N4141, N4139);
xor XOR2 (N4142, N4138, N3485);
nor NOR3 (N4143, N4128, N1715, N2620);
nor NOR2 (N4144, N4143, N346);
not NOT1 (N4145, N4136);
xor XOR2 (N4146, N4130, N3478);
buf BUF1 (N4147, N4131);
not NOT1 (N4148, N4140);
not NOT1 (N4149, N4137);
nand NAND3 (N4150, N4147, N905, N3045);
or OR4 (N4151, N4146, N1736, N875, N1151);
or OR2 (N4152, N4151, N2646);
nand NAND3 (N4153, N4144, N750, N1914);
buf BUF1 (N4154, N4148);
not NOT1 (N4155, N4153);
xor XOR2 (N4156, N4152, N2707);
xor XOR2 (N4157, N4132, N2978);
nor NOR4 (N4158, N4141, N379, N839, N3325);
nand NAND4 (N4159, N4145, N3767, N3285, N3562);
and AND2 (N4160, N4135, N2802);
xor XOR2 (N4161, N4160, N3734);
xor XOR2 (N4162, N4150, N1596);
not NOT1 (N4163, N4156);
and AND3 (N4164, N4149, N3117, N238);
not NOT1 (N4165, N4164);
buf BUF1 (N4166, N4163);
nor NOR2 (N4167, N4155, N2426);
buf BUF1 (N4168, N4142);
nand NAND3 (N4169, N4167, N2001, N572);
or OR2 (N4170, N4154, N1306);
and AND3 (N4171, N4161, N3349, N3018);
or OR2 (N4172, N4157, N3023);
nor NOR2 (N4173, N4162, N2295);
not NOT1 (N4174, N4159);
and AND3 (N4175, N4171, N1982, N2148);
buf BUF1 (N4176, N4166);
xor XOR2 (N4177, N4158, N2404);
and AND3 (N4178, N4176, N3349, N2912);
xor XOR2 (N4179, N4168, N1094);
nor NOR3 (N4180, N4172, N3255, N50);
nor NOR3 (N4181, N4177, N60, N1509);
or OR2 (N4182, N4174, N2242);
xor XOR2 (N4183, N4175, N2350);
buf BUF1 (N4184, N4170);
nand NAND3 (N4185, N4173, N3980, N2374);
xor XOR2 (N4186, N4182, N2390);
xor XOR2 (N4187, N4180, N2035);
nand NAND2 (N4188, N4181, N1824);
or OR3 (N4189, N4183, N1644, N3312);
xor XOR2 (N4190, N4189, N2896);
nand NAND3 (N4191, N4178, N1969, N2225);
xor XOR2 (N4192, N4190, N3391);
not NOT1 (N4193, N4184);
xor XOR2 (N4194, N4193, N1629);
or OR4 (N4195, N4194, N4013, N4153, N3158);
xor XOR2 (N4196, N4192, N2574);
not NOT1 (N4197, N4186);
nand NAND3 (N4198, N4191, N1809, N2345);
xor XOR2 (N4199, N4198, N1553);
not NOT1 (N4200, N4196);
and AND4 (N4201, N4197, N1403, N2275, N469);
or OR2 (N4202, N4185, N1648);
xor XOR2 (N4203, N4165, N1875);
not NOT1 (N4204, N4199);
not NOT1 (N4205, N4195);
nor NOR4 (N4206, N4179, N2681, N499, N3844);
and AND4 (N4207, N4169, N1415, N816, N1719);
not NOT1 (N4208, N4205);
or OR2 (N4209, N4188, N43);
or OR4 (N4210, N4200, N1707, N2181, N1080);
nor NOR4 (N4211, N4209, N872, N3492, N1193);
and AND2 (N4212, N4203, N3421);
or OR2 (N4213, N4212, N742);
xor XOR2 (N4214, N4207, N2866);
nor NOR3 (N4215, N4211, N2827, N1985);
buf BUF1 (N4216, N4215);
nor NOR2 (N4217, N4201, N1566);
xor XOR2 (N4218, N4204, N721);
buf BUF1 (N4219, N4213);
xor XOR2 (N4220, N4214, N1522);
nor NOR3 (N4221, N4219, N645, N106);
and AND3 (N4222, N4208, N1925, N2767);
xor XOR2 (N4223, N4206, N4118);
or OR2 (N4224, N4210, N2992);
and AND3 (N4225, N4218, N2893, N1053);
buf BUF1 (N4226, N4221);
not NOT1 (N4227, N4224);
nand NAND4 (N4228, N4225, N1861, N3775, N3507);
nand NAND4 (N4229, N4226, N3213, N1279, N4143);
or OR2 (N4230, N4229, N2857);
nor NOR3 (N4231, N4217, N2434, N2794);
not NOT1 (N4232, N4187);
or OR3 (N4233, N4222, N2124, N2017);
xor XOR2 (N4234, N4232, N3594);
xor XOR2 (N4235, N4216, N3597);
not NOT1 (N4236, N4230);
and AND2 (N4237, N4233, N1100);
or OR3 (N4238, N4234, N1845, N3359);
and AND2 (N4239, N4223, N1104);
nand NAND2 (N4240, N4227, N124);
nor NOR4 (N4241, N4239, N827, N266, N4230);
not NOT1 (N4242, N4237);
or OR3 (N4243, N4235, N4081, N2410);
not NOT1 (N4244, N4242);
nand NAND3 (N4245, N4231, N174, N589);
xor XOR2 (N4246, N4228, N377);
not NOT1 (N4247, N4236);
and AND3 (N4248, N4202, N2335, N2150);
not NOT1 (N4249, N4241);
buf BUF1 (N4250, N4245);
not NOT1 (N4251, N4248);
buf BUF1 (N4252, N4220);
and AND2 (N4253, N4249, N3119);
buf BUF1 (N4254, N4250);
and AND2 (N4255, N4252, N1372);
buf BUF1 (N4256, N4244);
xor XOR2 (N4257, N4251, N2578);
or OR3 (N4258, N4257, N280, N568);
not NOT1 (N4259, N4256);
buf BUF1 (N4260, N4255);
and AND4 (N4261, N4253, N3688, N1543, N447);
buf BUF1 (N4262, N4238);
xor XOR2 (N4263, N4261, N1378);
or OR3 (N4264, N4247, N2358, N1845);
or OR2 (N4265, N4243, N3389);
or OR2 (N4266, N4265, N650);
or OR4 (N4267, N4264, N1211, N3755, N3598);
or OR2 (N4268, N4254, N1314);
and AND3 (N4269, N4267, N3938, N1212);
nand NAND2 (N4270, N4263, N3554);
not NOT1 (N4271, N4260);
nand NAND4 (N4272, N4262, N1366, N2230, N1368);
and AND2 (N4273, N4271, N2835);
xor XOR2 (N4274, N4270, N4090);
nor NOR3 (N4275, N4266, N3115, N24);
nor NOR2 (N4276, N4259, N3546);
nand NAND2 (N4277, N4240, N1568);
buf BUF1 (N4278, N4274);
not NOT1 (N4279, N4268);
nand NAND4 (N4280, N4246, N1670, N1794, N289);
and AND3 (N4281, N4279, N4268, N783);
nand NAND2 (N4282, N4277, N2201);
xor XOR2 (N4283, N4282, N954);
xor XOR2 (N4284, N4278, N3403);
buf BUF1 (N4285, N4284);
or OR3 (N4286, N4283, N2927, N4004);
and AND3 (N4287, N4269, N3012, N1414);
nor NOR4 (N4288, N4281, N775, N4246, N3415);
and AND3 (N4289, N4285, N1590, N1948);
buf BUF1 (N4290, N4289);
or OR4 (N4291, N4286, N3697, N4236, N1288);
nand NAND3 (N4292, N4273, N1622, N43);
or OR3 (N4293, N4292, N1359, N1170);
or OR4 (N4294, N4291, N514, N1032, N73);
and AND2 (N4295, N4287, N3611);
nor NOR3 (N4296, N4288, N40, N1003);
not NOT1 (N4297, N4276);
and AND4 (N4298, N4290, N240, N103, N2801);
not NOT1 (N4299, N4293);
not NOT1 (N4300, N4296);
nand NAND3 (N4301, N4258, N4065, N3824);
and AND3 (N4302, N4301, N3769, N2822);
nor NOR2 (N4303, N4297, N1532);
buf BUF1 (N4304, N4302);
nand NAND4 (N4305, N4300, N1491, N3646, N589);
buf BUF1 (N4306, N4280);
nor NOR4 (N4307, N4298, N1656, N1143, N613);
and AND2 (N4308, N4299, N553);
xor XOR2 (N4309, N4307, N3556);
buf BUF1 (N4310, N4309);
buf BUF1 (N4311, N4310);
buf BUF1 (N4312, N4308);
buf BUF1 (N4313, N4306);
xor XOR2 (N4314, N4312, N879);
and AND4 (N4315, N4275, N2721, N2773, N1687);
buf BUF1 (N4316, N4313);
nor NOR3 (N4317, N4316, N1046, N3994);
or OR4 (N4318, N4294, N2445, N2596, N3449);
nor NOR2 (N4319, N4317, N125);
and AND2 (N4320, N4272, N971);
nand NAND3 (N4321, N4304, N1343, N716);
nand NAND3 (N4322, N4314, N437, N2095);
buf BUF1 (N4323, N4311);
xor XOR2 (N4324, N4318, N3546);
and AND3 (N4325, N4319, N1056, N313);
nor NOR2 (N4326, N4324, N2037);
nand NAND4 (N4327, N4315, N1231, N4278, N2047);
xor XOR2 (N4328, N4295, N4097);
xor XOR2 (N4329, N4323, N1503);
nand NAND2 (N4330, N4329, N3376);
buf BUF1 (N4331, N4321);
not NOT1 (N4332, N4320);
nand NAND3 (N4333, N4303, N4075, N3079);
not NOT1 (N4334, N4325);
nor NOR3 (N4335, N4326, N2021, N340);
not NOT1 (N4336, N4332);
and AND3 (N4337, N4335, N2327, N2339);
and AND2 (N4338, N4327, N4137);
buf BUF1 (N4339, N4336);
and AND2 (N4340, N4334, N755);
nor NOR2 (N4341, N4322, N2326);
nand NAND4 (N4342, N4328, N1268, N2277, N1625);
and AND2 (N4343, N4341, N3307);
xor XOR2 (N4344, N4343, N739);
nor NOR2 (N4345, N4331, N3310);
nor NOR4 (N4346, N4342, N3531, N162, N2555);
and AND4 (N4347, N4337, N1016, N1377, N976);
nand NAND2 (N4348, N4346, N1757);
not NOT1 (N4349, N4344);
buf BUF1 (N4350, N4349);
nand NAND3 (N4351, N4345, N1280, N1224);
and AND2 (N4352, N4333, N2361);
not NOT1 (N4353, N4340);
or OR4 (N4354, N4353, N4348, N2815, N2141);
nor NOR3 (N4355, N461, N2503, N2961);
xor XOR2 (N4356, N4355, N3742);
xor XOR2 (N4357, N4305, N3068);
nand NAND4 (N4358, N4352, N1185, N1456, N1786);
buf BUF1 (N4359, N4338);
nor NOR2 (N4360, N4347, N2072);
not NOT1 (N4361, N4358);
buf BUF1 (N4362, N4359);
buf BUF1 (N4363, N4361);
not NOT1 (N4364, N4363);
nor NOR2 (N4365, N4354, N3010);
nor NOR2 (N4366, N4360, N3415);
buf BUF1 (N4367, N4330);
buf BUF1 (N4368, N4350);
buf BUF1 (N4369, N4356);
and AND2 (N4370, N4339, N3066);
nand NAND4 (N4371, N4367, N953, N2586, N1365);
nand NAND2 (N4372, N4351, N776);
xor XOR2 (N4373, N4357, N2634);
or OR4 (N4374, N4369, N1731, N3954, N220);
buf BUF1 (N4375, N4362);
nand NAND4 (N4376, N4371, N1259, N365, N4288);
xor XOR2 (N4377, N4370, N1742);
not NOT1 (N4378, N4377);
buf BUF1 (N4379, N4376);
xor XOR2 (N4380, N4368, N1846);
buf BUF1 (N4381, N4380);
nand NAND3 (N4382, N4378, N2136, N2825);
and AND4 (N4383, N4374, N3941, N1302, N2715);
nand NAND4 (N4384, N4372, N180, N3145, N3677);
nor NOR4 (N4385, N4381, N4084, N2798, N775);
not NOT1 (N4386, N4385);
nand NAND2 (N4387, N4365, N1304);
and AND3 (N4388, N4383, N3086, N2940);
nand NAND2 (N4389, N4384, N49);
nor NOR3 (N4390, N4387, N1446, N74);
nand NAND2 (N4391, N4373, N3044);
or OR2 (N4392, N4375, N2734);
xor XOR2 (N4393, N4388, N316);
buf BUF1 (N4394, N4390);
and AND2 (N4395, N4394, N1445);
nor NOR2 (N4396, N4364, N1624);
nand NAND3 (N4397, N4392, N2772, N2785);
not NOT1 (N4398, N4366);
xor XOR2 (N4399, N4397, N3568);
or OR3 (N4400, N4389, N1807, N4393);
not NOT1 (N4401, N3358);
nor NOR4 (N4402, N4395, N691, N169, N2244);
or OR2 (N4403, N4396, N3454);
not NOT1 (N4404, N4402);
buf BUF1 (N4405, N4382);
nor NOR2 (N4406, N4401, N3107);
buf BUF1 (N4407, N4399);
nand NAND2 (N4408, N4379, N2360);
xor XOR2 (N4409, N4386, N2390);
buf BUF1 (N4410, N4409);
and AND2 (N4411, N4404, N871);
nand NAND4 (N4412, N4406, N3760, N3478, N1357);
xor XOR2 (N4413, N4412, N1134);
nand NAND2 (N4414, N4413, N2737);
nor NOR2 (N4415, N4407, N2346);
nand NAND4 (N4416, N4411, N3831, N3874, N3358);
and AND3 (N4417, N4398, N3640, N1085);
and AND4 (N4418, N4408, N2071, N1153, N3202);
or OR3 (N4419, N4414, N3924, N212);
buf BUF1 (N4420, N4410);
and AND3 (N4421, N4417, N2846, N1781);
buf BUF1 (N4422, N4421);
nor NOR4 (N4423, N4422, N4272, N1938, N1850);
buf BUF1 (N4424, N4400);
nand NAND3 (N4425, N4416, N2819, N3073);
buf BUF1 (N4426, N4418);
or OR4 (N4427, N4426, N756, N3368, N470);
nand NAND2 (N4428, N4424, N1706);
or OR4 (N4429, N4391, N3384, N1171, N1095);
and AND3 (N4430, N4405, N3014, N675);
nand NAND3 (N4431, N4427, N3708, N928);
nand NAND4 (N4432, N4415, N4304, N1128, N704);
or OR3 (N4433, N4432, N1961, N3505);
or OR3 (N4434, N4433, N4335, N4093);
and AND3 (N4435, N4430, N1817, N4205);
not NOT1 (N4436, N4420);
not NOT1 (N4437, N4425);
nor NOR4 (N4438, N4437, N2628, N2475, N3874);
or OR2 (N4439, N4438, N1006);
xor XOR2 (N4440, N4419, N2518);
not NOT1 (N4441, N4429);
or OR4 (N4442, N4403, N2702, N1115, N1190);
nand NAND2 (N4443, N4441, N1851);
nor NOR3 (N4444, N4428, N873, N2166);
buf BUF1 (N4445, N4444);
nand NAND3 (N4446, N4445, N2904, N644);
buf BUF1 (N4447, N4439);
nand NAND3 (N4448, N4446, N1815, N2778);
or OR3 (N4449, N4435, N402, N1463);
buf BUF1 (N4450, N4434);
xor XOR2 (N4451, N4440, N426);
nand NAND2 (N4452, N4442, N3985);
nor NOR2 (N4453, N4431, N570);
or OR2 (N4454, N4448, N2831);
buf BUF1 (N4455, N4450);
nand NAND2 (N4456, N4455, N3412);
not NOT1 (N4457, N4449);
and AND4 (N4458, N4451, N1015, N3100, N1303);
or OR4 (N4459, N4436, N206, N1424, N116);
not NOT1 (N4460, N4459);
not NOT1 (N4461, N4447);
nor NOR3 (N4462, N4454, N4386, N1274);
nand NAND4 (N4463, N4452, N703, N3809, N536);
buf BUF1 (N4464, N4463);
nor NOR2 (N4465, N4443, N2700);
or OR4 (N4466, N4457, N1004, N3578, N3133);
buf BUF1 (N4467, N4461);
not NOT1 (N4468, N4466);
and AND3 (N4469, N4458, N2442, N1061);
nor NOR2 (N4470, N4464, N3884);
xor XOR2 (N4471, N4469, N387);
buf BUF1 (N4472, N4468);
or OR2 (N4473, N4471, N2498);
buf BUF1 (N4474, N4462);
nor NOR4 (N4475, N4465, N68, N2486, N1088);
nor NOR3 (N4476, N4423, N2664, N3366);
buf BUF1 (N4477, N4467);
xor XOR2 (N4478, N4472, N2573);
or OR4 (N4479, N4477, N2485, N1061, N4257);
xor XOR2 (N4480, N4476, N3130);
or OR2 (N4481, N4478, N508);
nand NAND2 (N4482, N4453, N1201);
and AND4 (N4483, N4481, N1837, N1215, N1017);
not NOT1 (N4484, N4474);
nand NAND4 (N4485, N4460, N3811, N3903, N3168);
or OR2 (N4486, N4483, N2157);
buf BUF1 (N4487, N4456);
and AND2 (N4488, N4485, N3948);
xor XOR2 (N4489, N4482, N638);
or OR2 (N4490, N4486, N1689);
nand NAND4 (N4491, N4480, N923, N958, N4097);
buf BUF1 (N4492, N4487);
not NOT1 (N4493, N4491);
nor NOR2 (N4494, N4473, N3088);
or OR4 (N4495, N4475, N4258, N1335, N2547);
and AND3 (N4496, N4479, N1452, N2128);
not NOT1 (N4497, N4470);
nand NAND3 (N4498, N4497, N2803, N3405);
or OR3 (N4499, N4488, N1308, N2313);
nor NOR3 (N4500, N4498, N4380, N2772);
not NOT1 (N4501, N4494);
nor NOR2 (N4502, N4489, N2578);
and AND3 (N4503, N4500, N1149, N3950);
and AND2 (N4504, N4499, N585);
nand NAND3 (N4505, N4490, N1294, N2101);
nor NOR2 (N4506, N4504, N2088);
and AND4 (N4507, N4495, N2859, N3859, N2482);
buf BUF1 (N4508, N4506);
buf BUF1 (N4509, N4507);
not NOT1 (N4510, N4503);
buf BUF1 (N4511, N4492);
and AND2 (N4512, N4501, N1628);
nor NOR2 (N4513, N4493, N554);
xor XOR2 (N4514, N4510, N4432);
nor NOR2 (N4515, N4496, N1403);
and AND4 (N4516, N4511, N517, N2357, N3978);
and AND2 (N4517, N4502, N3287);
nand NAND2 (N4518, N4514, N2833);
not NOT1 (N4519, N4508);
not NOT1 (N4520, N4505);
nand NAND2 (N4521, N4512, N3806);
or OR3 (N4522, N4509, N1945, N4356);
or OR3 (N4523, N4513, N1786, N3232);
xor XOR2 (N4524, N4521, N4369);
buf BUF1 (N4525, N4515);
nand NAND2 (N4526, N4516, N3052);
nor NOR2 (N4527, N4522, N52);
nor NOR3 (N4528, N4524, N1481, N3017);
not NOT1 (N4529, N4484);
or OR3 (N4530, N4527, N3209, N2484);
nand NAND3 (N4531, N4519, N4507, N3255);
xor XOR2 (N4532, N4520, N11);
and AND2 (N4533, N4530, N1322);
nor NOR3 (N4534, N4523, N2350, N3902);
nand NAND3 (N4535, N4533, N1141, N3882);
or OR2 (N4536, N4526, N623);
or OR4 (N4537, N4531, N2086, N2960, N765);
and AND4 (N4538, N4534, N2397, N2599, N4431);
and AND2 (N4539, N4538, N2835);
nor NOR2 (N4540, N4536, N3907);
not NOT1 (N4541, N4525);
buf BUF1 (N4542, N4535);
nand NAND4 (N4543, N4540, N1375, N4506, N4513);
nand NAND4 (N4544, N4532, N4301, N4264, N3470);
or OR4 (N4545, N4543, N1138, N3735, N3228);
or OR4 (N4546, N4541, N2245, N2356, N3532);
nand NAND2 (N4547, N4545, N433);
nand NAND3 (N4548, N4518, N1558, N2698);
buf BUF1 (N4549, N4529);
nor NOR2 (N4550, N4547, N3097);
and AND4 (N4551, N4544, N583, N99, N567);
buf BUF1 (N4552, N4549);
or OR4 (N4553, N4539, N2692, N2410, N2199);
not NOT1 (N4554, N4542);
buf BUF1 (N4555, N4517);
nor NOR3 (N4556, N4552, N4375, N3235);
not NOT1 (N4557, N4546);
xor XOR2 (N4558, N4555, N1047);
xor XOR2 (N4559, N4556, N3505);
nor NOR3 (N4560, N4537, N2479, N695);
nor NOR2 (N4561, N4548, N4303);
nand NAND4 (N4562, N4560, N1023, N4504, N2258);
buf BUF1 (N4563, N4551);
buf BUF1 (N4564, N4557);
not NOT1 (N4565, N4562);
nor NOR3 (N4566, N4563, N968, N3070);
xor XOR2 (N4567, N4554, N3760);
nor NOR2 (N4568, N4558, N2318);
xor XOR2 (N4569, N4568, N2736);
or OR4 (N4570, N4566, N3026, N2161, N2720);
xor XOR2 (N4571, N4528, N1963);
buf BUF1 (N4572, N4570);
nand NAND3 (N4573, N4550, N3860, N4492);
not NOT1 (N4574, N4559);
xor XOR2 (N4575, N4553, N534);
or OR4 (N4576, N4572, N3553, N134, N3824);
buf BUF1 (N4577, N4576);
or OR4 (N4578, N4569, N4123, N3917, N4349);
nand NAND4 (N4579, N4564, N637, N553, N4503);
and AND2 (N4580, N4574, N3447);
nor NOR3 (N4581, N4573, N30, N2971);
buf BUF1 (N4582, N4575);
and AND2 (N4583, N4580, N3397);
xor XOR2 (N4584, N4577, N851);
nor NOR2 (N4585, N4561, N480);
nor NOR4 (N4586, N4567, N3457, N140, N3834);
and AND4 (N4587, N4586, N3395, N3849, N3734);
not NOT1 (N4588, N4584);
or OR2 (N4589, N4583, N1270);
buf BUF1 (N4590, N4585);
or OR3 (N4591, N4578, N3831, N625);
nand NAND4 (N4592, N4582, N4591, N714, N1090);
buf BUF1 (N4593, N2329);
not NOT1 (N4594, N4579);
buf BUF1 (N4595, N4589);
buf BUF1 (N4596, N4595);
xor XOR2 (N4597, N4565, N4064);
nor NOR4 (N4598, N4587, N3492, N68, N1309);
xor XOR2 (N4599, N4581, N4045);
buf BUF1 (N4600, N4594);
xor XOR2 (N4601, N4590, N4389);
buf BUF1 (N4602, N4599);
nand NAND2 (N4603, N4602, N2913);
buf BUF1 (N4604, N4592);
or OR4 (N4605, N4598, N477, N965, N636);
not NOT1 (N4606, N4588);
or OR2 (N4607, N4605, N571);
and AND2 (N4608, N4597, N4206);
buf BUF1 (N4609, N4608);
xor XOR2 (N4610, N4601, N409);
or OR3 (N4611, N4600, N3359, N792);
xor XOR2 (N4612, N4593, N2116);
and AND2 (N4613, N4610, N1410);
xor XOR2 (N4614, N4613, N962);
not NOT1 (N4615, N4614);
not NOT1 (N4616, N4606);
nor NOR3 (N4617, N4607, N2967, N603);
nand NAND4 (N4618, N4603, N2756, N1885, N3370);
nor NOR2 (N4619, N4615, N2994);
and AND3 (N4620, N4609, N3484, N3766);
buf BUF1 (N4621, N4617);
nor NOR3 (N4622, N4571, N1180, N4030);
nor NOR4 (N4623, N4621, N4508, N1920, N4131);
nor NOR3 (N4624, N4612, N192, N2778);
and AND3 (N4625, N4596, N3115, N357);
and AND2 (N4626, N4625, N870);
not NOT1 (N4627, N4626);
not NOT1 (N4628, N4623);
nand NAND2 (N4629, N4628, N3008);
nor NOR4 (N4630, N4616, N3990, N501, N684);
xor XOR2 (N4631, N4630, N3537);
buf BUF1 (N4632, N4629);
buf BUF1 (N4633, N4619);
buf BUF1 (N4634, N4631);
buf BUF1 (N4635, N4633);
xor XOR2 (N4636, N4620, N3929);
and AND3 (N4637, N4636, N421, N2485);
nor NOR2 (N4638, N4634, N1828);
buf BUF1 (N4639, N4624);
xor XOR2 (N4640, N4618, N4059);
xor XOR2 (N4641, N4604, N3874);
nand NAND2 (N4642, N4611, N1162);
not NOT1 (N4643, N4640);
nor NOR3 (N4644, N4627, N3286, N3868);
buf BUF1 (N4645, N4643);
and AND2 (N4646, N4637, N3943);
or OR2 (N4647, N4641, N2355);
nor NOR4 (N4648, N4622, N3875, N2812, N2568);
nand NAND3 (N4649, N4639, N1403, N3469);
buf BUF1 (N4650, N4642);
xor XOR2 (N4651, N4635, N3695);
buf BUF1 (N4652, N4649);
not NOT1 (N4653, N4644);
xor XOR2 (N4654, N4651, N776);
buf BUF1 (N4655, N4638);
not NOT1 (N4656, N4650);
or OR3 (N4657, N4655, N2377, N591);
buf BUF1 (N4658, N4645);
not NOT1 (N4659, N4648);
buf BUF1 (N4660, N4632);
nor NOR4 (N4661, N4659, N4522, N2612, N3127);
not NOT1 (N4662, N4657);
nor NOR3 (N4663, N4660, N1596, N3835);
nor NOR4 (N4664, N4654, N2954, N1224, N1923);
and AND3 (N4665, N4656, N3605, N3936);
or OR2 (N4666, N4661, N566);
buf BUF1 (N4667, N4647);
buf BUF1 (N4668, N4658);
buf BUF1 (N4669, N4665);
nand NAND2 (N4670, N4668, N3917);
nand NAND4 (N4671, N4662, N3369, N3799, N715);
or OR2 (N4672, N4669, N2682);
or OR3 (N4673, N4663, N2790, N4532);
buf BUF1 (N4674, N4673);
not NOT1 (N4675, N4672);
xor XOR2 (N4676, N4666, N972);
not NOT1 (N4677, N4676);
not NOT1 (N4678, N4677);
buf BUF1 (N4679, N4652);
nor NOR4 (N4680, N4674, N2814, N354, N4120);
not NOT1 (N4681, N4646);
nand NAND2 (N4682, N4675, N2537);
xor XOR2 (N4683, N4681, N3077);
not NOT1 (N4684, N4664);
buf BUF1 (N4685, N4683);
and AND4 (N4686, N4679, N3645, N1091, N2666);
and AND2 (N4687, N4671, N434);
and AND4 (N4688, N4687, N3072, N668, N2321);
not NOT1 (N4689, N4688);
nand NAND3 (N4690, N4684, N3721, N1821);
and AND3 (N4691, N4667, N2079, N2784);
and AND2 (N4692, N4653, N558);
nor NOR3 (N4693, N4686, N4241, N2922);
xor XOR2 (N4694, N4691, N4457);
buf BUF1 (N4695, N4692);
and AND3 (N4696, N4693, N3378, N3124);
not NOT1 (N4697, N4695);
or OR4 (N4698, N4689, N2311, N2801, N1205);
and AND2 (N4699, N4682, N4476);
not NOT1 (N4700, N4694);
not NOT1 (N4701, N4697);
xor XOR2 (N4702, N4696, N2153);
nor NOR3 (N4703, N4690, N4213, N2452);
not NOT1 (N4704, N4698);
or OR2 (N4705, N4703, N4027);
not NOT1 (N4706, N4701);
nor NOR4 (N4707, N4705, N4526, N358, N3100);
or OR2 (N4708, N4706, N1852);
buf BUF1 (N4709, N4702);
not NOT1 (N4710, N4708);
or OR2 (N4711, N4699, N575);
nand NAND2 (N4712, N4700, N3361);
nand NAND4 (N4713, N4710, N4491, N974, N167);
nand NAND4 (N4714, N4678, N3042, N451, N2708);
buf BUF1 (N4715, N4707);
nor NOR2 (N4716, N4704, N977);
or OR3 (N4717, N4670, N4173, N3982);
nor NOR3 (N4718, N4712, N3192, N3282);
buf BUF1 (N4719, N4680);
not NOT1 (N4720, N4718);
nand NAND2 (N4721, N4716, N143);
nor NOR3 (N4722, N4713, N1390, N232);
not NOT1 (N4723, N4715);
and AND4 (N4724, N4717, N953, N3009, N1907);
nand NAND4 (N4725, N4722, N4437, N4450, N4086);
nor NOR2 (N4726, N4719, N3526);
nand NAND2 (N4727, N4723, N606);
nor NOR3 (N4728, N4685, N3512, N4681);
not NOT1 (N4729, N4714);
not NOT1 (N4730, N4728);
nor NOR4 (N4731, N4724, N3679, N4207, N2585);
not NOT1 (N4732, N4729);
not NOT1 (N4733, N4730);
nand NAND3 (N4734, N4709, N1537, N1296);
nand NAND4 (N4735, N4734, N4235, N3720, N4604);
not NOT1 (N4736, N4720);
not NOT1 (N4737, N4711);
and AND2 (N4738, N4735, N122);
nor NOR2 (N4739, N4727, N2314);
not NOT1 (N4740, N4726);
nand NAND3 (N4741, N4736, N3361, N3837);
nand NAND2 (N4742, N4721, N1557);
nor NOR2 (N4743, N4737, N1640);
xor XOR2 (N4744, N4741, N3282);
not NOT1 (N4745, N4725);
not NOT1 (N4746, N4745);
or OR2 (N4747, N4732, N3727);
buf BUF1 (N4748, N4746);
nand NAND3 (N4749, N4731, N1953, N5);
nand NAND3 (N4750, N4749, N990, N492);
buf BUF1 (N4751, N4733);
xor XOR2 (N4752, N4742, N1713);
not NOT1 (N4753, N4738);
not NOT1 (N4754, N4739);
or OR4 (N4755, N4750, N1058, N4111, N4162);
not NOT1 (N4756, N4752);
buf BUF1 (N4757, N4744);
xor XOR2 (N4758, N4743, N1824);
xor XOR2 (N4759, N4755, N4045);
nand NAND2 (N4760, N4747, N2124);
buf BUF1 (N4761, N4760);
nor NOR2 (N4762, N4754, N712);
or OR2 (N4763, N4748, N3733);
and AND4 (N4764, N4740, N3826, N560, N3091);
or OR3 (N4765, N4753, N1178, N3440);
buf BUF1 (N4766, N4761);
and AND3 (N4767, N4758, N925, N4400);
nor NOR4 (N4768, N4766, N4608, N4298, N4019);
not NOT1 (N4769, N4757);
or OR2 (N4770, N4765, N2512);
xor XOR2 (N4771, N4767, N2877);
nand NAND4 (N4772, N4759, N2208, N2119, N1582);
not NOT1 (N4773, N4762);
not NOT1 (N4774, N4771);
not NOT1 (N4775, N4763);
not NOT1 (N4776, N4756);
and AND2 (N4777, N4772, N1951);
buf BUF1 (N4778, N4776);
nand NAND4 (N4779, N4777, N2252, N2363, N2495);
nand NAND2 (N4780, N4768, N457);
nor NOR4 (N4781, N4764, N4735, N4107, N960);
nand NAND4 (N4782, N4751, N1447, N3078, N4262);
nand NAND3 (N4783, N4781, N828, N117);
buf BUF1 (N4784, N4782);
nand NAND3 (N4785, N4783, N2125, N1508);
and AND3 (N4786, N4785, N3126, N1994);
xor XOR2 (N4787, N4780, N111);
or OR2 (N4788, N4773, N4747);
nor NOR4 (N4789, N4786, N1645, N593, N4742);
buf BUF1 (N4790, N4784);
xor XOR2 (N4791, N4778, N2514);
xor XOR2 (N4792, N4774, N2157);
nor NOR4 (N4793, N4790, N2949, N1993, N2943);
or OR4 (N4794, N4770, N3764, N1965, N1526);
not NOT1 (N4795, N4775);
xor XOR2 (N4796, N4791, N4238);
nand NAND4 (N4797, N4787, N3987, N2524, N147);
nand NAND2 (N4798, N4788, N4707);
nor NOR2 (N4799, N4797, N154);
not NOT1 (N4800, N4779);
buf BUF1 (N4801, N4796);
xor XOR2 (N4802, N4793, N1424);
or OR4 (N4803, N4795, N247, N2743, N2766);
and AND4 (N4804, N4802, N3997, N4719, N1043);
or OR4 (N4805, N4789, N1130, N1659, N961);
buf BUF1 (N4806, N4803);
not NOT1 (N4807, N4798);
nor NOR3 (N4808, N4804, N3844, N411);
not NOT1 (N4809, N4800);
or OR4 (N4810, N4801, N3573, N2024, N3987);
xor XOR2 (N4811, N4808, N1017);
buf BUF1 (N4812, N4769);
nand NAND2 (N4813, N4812, N556);
buf BUF1 (N4814, N4806);
buf BUF1 (N4815, N4814);
and AND4 (N4816, N4809, N1502, N842, N3515);
or OR3 (N4817, N4816, N4429, N1920);
or OR3 (N4818, N4817, N1219, N4071);
not NOT1 (N4819, N4807);
xor XOR2 (N4820, N4810, N2970);
xor XOR2 (N4821, N4799, N3425);
or OR3 (N4822, N4818, N2703, N2471);
xor XOR2 (N4823, N4822, N4214);
buf BUF1 (N4824, N4805);
nor NOR2 (N4825, N4811, N2050);
not NOT1 (N4826, N4820);
and AND2 (N4827, N4826, N3033);
nand NAND3 (N4828, N4827, N1811, N2421);
buf BUF1 (N4829, N4815);
and AND2 (N4830, N4813, N1622);
not NOT1 (N4831, N4825);
nor NOR3 (N4832, N4830, N908, N760);
nor NOR3 (N4833, N4824, N298, N1880);
xor XOR2 (N4834, N4831, N1736);
and AND3 (N4835, N4819, N1202, N705);
buf BUF1 (N4836, N4794);
buf BUF1 (N4837, N4834);
not NOT1 (N4838, N4837);
buf BUF1 (N4839, N4836);
nor NOR2 (N4840, N4832, N255);
and AND4 (N4841, N4829, N4618, N878, N2856);
buf BUF1 (N4842, N4835);
nand NAND2 (N4843, N4840, N2688);
buf BUF1 (N4844, N4833);
nand NAND2 (N4845, N4842, N2226);
xor XOR2 (N4846, N4839, N4693);
or OR3 (N4847, N4838, N4148, N4703);
xor XOR2 (N4848, N4823, N2738);
nand NAND2 (N4849, N4828, N2685);
not NOT1 (N4850, N4845);
not NOT1 (N4851, N4843);
nor NOR4 (N4852, N4821, N3814, N3340, N338);
or OR3 (N4853, N4846, N2864, N32);
and AND4 (N4854, N4851, N4546, N2293, N2734);
or OR3 (N4855, N4852, N3337, N4536);
nor NOR4 (N4856, N4850, N4302, N2251, N781);
buf BUF1 (N4857, N4855);
nand NAND4 (N4858, N4857, N482, N2515, N1952);
xor XOR2 (N4859, N4854, N970);
xor XOR2 (N4860, N4858, N1670);
nand NAND4 (N4861, N4853, N3503, N4662, N2411);
nor NOR2 (N4862, N4841, N4804);
not NOT1 (N4863, N4856);
buf BUF1 (N4864, N4844);
nand NAND2 (N4865, N4860, N2859);
nand NAND4 (N4866, N4863, N2483, N1509, N345);
not NOT1 (N4867, N4859);
not NOT1 (N4868, N4862);
nand NAND4 (N4869, N4868, N4437, N4308, N4666);
xor XOR2 (N4870, N4792, N3029);
nand NAND2 (N4871, N4861, N766);
nor NOR2 (N4872, N4871, N2972);
nand NAND2 (N4873, N4869, N107);
xor XOR2 (N4874, N4872, N2768);
nor NOR3 (N4875, N4865, N3478, N1479);
or OR4 (N4876, N4866, N2728, N2608, N4797);
buf BUF1 (N4877, N4876);
buf BUF1 (N4878, N4873);
or OR2 (N4879, N4867, N1615);
nand NAND4 (N4880, N4849, N2688, N3795, N3502);
xor XOR2 (N4881, N4875, N1200);
not NOT1 (N4882, N4848);
and AND3 (N4883, N4880, N2725, N1478);
not NOT1 (N4884, N4864);
xor XOR2 (N4885, N4870, N191);
or OR4 (N4886, N4877, N1233, N2772, N2671);
nor NOR3 (N4887, N4882, N2919, N4362);
or OR4 (N4888, N4878, N3565, N3815, N4616);
and AND3 (N4889, N4887, N3692, N4169);
not NOT1 (N4890, N4879);
xor XOR2 (N4891, N4883, N2366);
not NOT1 (N4892, N4874);
buf BUF1 (N4893, N4890);
or OR2 (N4894, N4885, N3117);
not NOT1 (N4895, N4891);
nand NAND3 (N4896, N4894, N3211, N245);
nand NAND3 (N4897, N4886, N3855, N1750);
nor NOR2 (N4898, N4884, N2966);
not NOT1 (N4899, N4888);
buf BUF1 (N4900, N4893);
and AND2 (N4901, N4900, N3765);
xor XOR2 (N4902, N4898, N4660);
and AND3 (N4903, N4896, N3212, N183);
and AND2 (N4904, N4902, N4583);
buf BUF1 (N4905, N4892);
nand NAND4 (N4906, N4901, N1934, N146, N2825);
and AND4 (N4907, N4895, N4064, N3686, N2275);
buf BUF1 (N4908, N4906);
or OR4 (N4909, N4847, N1256, N437, N3223);
nand NAND4 (N4910, N4909, N4776, N1475, N2188);
and AND2 (N4911, N4904, N2);
nand NAND2 (N4912, N4907, N1897);
nand NAND4 (N4913, N4897, N4065, N4389, N130);
or OR2 (N4914, N4910, N2652);
not NOT1 (N4915, N4911);
or OR2 (N4916, N4889, N4547);
nand NAND3 (N4917, N4916, N1121, N1759);
and AND4 (N4918, N4899, N3249, N4822, N1279);
or OR4 (N4919, N4908, N490, N4461, N3293);
buf BUF1 (N4920, N4919);
buf BUF1 (N4921, N4913);
nand NAND2 (N4922, N4903, N3485);
and AND3 (N4923, N4920, N3419, N1129);
and AND4 (N4924, N4912, N515, N625, N4259);
and AND4 (N4925, N4917, N244, N4579, N535);
buf BUF1 (N4926, N4925);
nand NAND3 (N4927, N4921, N1840, N1149);
and AND3 (N4928, N4915, N2646, N3261);
buf BUF1 (N4929, N4924);
nand NAND4 (N4930, N4929, N2455, N1991, N213);
and AND3 (N4931, N4914, N179, N1775);
nor NOR4 (N4932, N4881, N268, N4322, N1309);
or OR4 (N4933, N4930, N4229, N2178, N1961);
not NOT1 (N4934, N4923);
xor XOR2 (N4935, N4933, N365);
or OR2 (N4936, N4927, N2023);
or OR2 (N4937, N4931, N4934);
buf BUF1 (N4938, N4015);
nor NOR4 (N4939, N4918, N591, N518, N2527);
or OR2 (N4940, N4928, N2477);
xor XOR2 (N4941, N4940, N4810);
nand NAND2 (N4942, N4941, N514);
nor NOR4 (N4943, N4942, N2841, N816, N4638);
xor XOR2 (N4944, N4936, N100);
not NOT1 (N4945, N4938);
not NOT1 (N4946, N4939);
nand NAND4 (N4947, N4926, N2009, N3723, N3713);
not NOT1 (N4948, N4947);
or OR3 (N4949, N4945, N4072, N3671);
nor NOR3 (N4950, N4948, N3202, N1971);
or OR2 (N4951, N4944, N1240);
nand NAND2 (N4952, N4951, N1501);
buf BUF1 (N4953, N4943);
buf BUF1 (N4954, N4935);
buf BUF1 (N4955, N4952);
buf BUF1 (N4956, N4922);
xor XOR2 (N4957, N4950, N2145);
xor XOR2 (N4958, N4946, N3677);
or OR4 (N4959, N4905, N1913, N79, N1201);
not NOT1 (N4960, N4957);
buf BUF1 (N4961, N4937);
nor NOR4 (N4962, N4932, N2856, N245, N1885);
buf BUF1 (N4963, N4954);
buf BUF1 (N4964, N4955);
or OR3 (N4965, N4963, N34, N4048);
xor XOR2 (N4966, N4958, N1412);
xor XOR2 (N4967, N4949, N2513);
nor NOR3 (N4968, N4962, N568, N1735);
xor XOR2 (N4969, N4959, N580);
buf BUF1 (N4970, N4956);
nor NOR2 (N4971, N4966, N2889);
nor NOR2 (N4972, N4967, N1798);
xor XOR2 (N4973, N4971, N3276);
buf BUF1 (N4974, N4960);
and AND2 (N4975, N4973, N3297);
xor XOR2 (N4976, N4972, N2961);
nor NOR2 (N4977, N4964, N2881);
and AND4 (N4978, N4961, N4646, N2188, N2380);
and AND4 (N4979, N4969, N2050, N2811, N431);
xor XOR2 (N4980, N4965, N1957);
or OR4 (N4981, N4953, N744, N677, N4690);
xor XOR2 (N4982, N4978, N1898);
buf BUF1 (N4983, N4979);
xor XOR2 (N4984, N4968, N1205);
xor XOR2 (N4985, N4981, N3050);
not NOT1 (N4986, N4985);
or OR2 (N4987, N4974, N4538);
buf BUF1 (N4988, N4984);
xor XOR2 (N4989, N4977, N3278);
nand NAND2 (N4990, N4980, N3147);
xor XOR2 (N4991, N4982, N4027);
nand NAND3 (N4992, N4990, N958, N4771);
or OR3 (N4993, N4988, N1236, N4629);
not NOT1 (N4994, N4989);
xor XOR2 (N4995, N4987, N941);
or OR4 (N4996, N4993, N3351, N360, N1682);
not NOT1 (N4997, N4994);
nand NAND2 (N4998, N4995, N121);
xor XOR2 (N4999, N4998, N3829);
nor NOR3 (N5000, N4976, N2787, N1426);
and AND2 (N5001, N4997, N2526);
nand NAND2 (N5002, N4991, N1871);
or OR2 (N5003, N5000, N2688);
buf BUF1 (N5004, N4999);
buf BUF1 (N5005, N4970);
xor XOR2 (N5006, N5002, N2819);
buf BUF1 (N5007, N5005);
or OR3 (N5008, N5001, N766, N2707);
buf BUF1 (N5009, N4983);
and AND4 (N5010, N5008, N1286, N3410, N3390);
and AND2 (N5011, N4975, N1935);
not NOT1 (N5012, N5011);
nor NOR3 (N5013, N5003, N2036, N4289);
or OR4 (N5014, N4996, N3943, N865, N1516);
xor XOR2 (N5015, N5010, N759);
and AND2 (N5016, N5004, N3740);
and AND3 (N5017, N5014, N218, N4153);
xor XOR2 (N5018, N5017, N4827);
and AND2 (N5019, N5006, N2209);
nand NAND3 (N5020, N5013, N4808, N2268);
xor XOR2 (N5021, N5018, N854);
or OR2 (N5022, N5021, N2149);
nor NOR2 (N5023, N5012, N4275);
buf BUF1 (N5024, N5007);
xor XOR2 (N5025, N5019, N4774);
nand NAND4 (N5026, N5016, N1721, N983, N1386);
buf BUF1 (N5027, N5026);
nand NAND2 (N5028, N5023, N830);
not NOT1 (N5029, N5020);
nor NOR3 (N5030, N4986, N1326, N3819);
xor XOR2 (N5031, N5029, N2424);
and AND4 (N5032, N5030, N4554, N2179, N903);
xor XOR2 (N5033, N5031, N2062);
not NOT1 (N5034, N5028);
nor NOR3 (N5035, N5024, N2315, N4781);
or OR2 (N5036, N5027, N4200);
nor NOR2 (N5037, N5022, N2726);
not NOT1 (N5038, N4992);
and AND3 (N5039, N5009, N3558, N196);
buf BUF1 (N5040, N5015);
and AND3 (N5041, N5039, N4259, N4712);
xor XOR2 (N5042, N5025, N3821);
xor XOR2 (N5043, N5036, N822);
not NOT1 (N5044, N5034);
or OR2 (N5045, N5037, N108);
or OR2 (N5046, N5038, N15);
buf BUF1 (N5047, N5041);
and AND2 (N5048, N5043, N4711);
nor NOR4 (N5049, N5048, N4694, N3374, N4432);
or OR2 (N5050, N5042, N513);
not NOT1 (N5051, N5047);
buf BUF1 (N5052, N5051);
not NOT1 (N5053, N5052);
nor NOR4 (N5054, N5049, N2879, N3455, N1627);
nand NAND2 (N5055, N5035, N2474);
not NOT1 (N5056, N5033);
or OR2 (N5057, N5045, N4220);
and AND3 (N5058, N5032, N4401, N3287);
xor XOR2 (N5059, N5055, N2181);
buf BUF1 (N5060, N5058);
xor XOR2 (N5061, N5040, N4664);
or OR2 (N5062, N5061, N2390);
xor XOR2 (N5063, N5057, N2139);
not NOT1 (N5064, N5060);
nor NOR3 (N5065, N5053, N2368, N1823);
xor XOR2 (N5066, N5056, N2209);
xor XOR2 (N5067, N5044, N1441);
buf BUF1 (N5068, N5065);
buf BUF1 (N5069, N5050);
and AND2 (N5070, N5054, N208);
not NOT1 (N5071, N5063);
xor XOR2 (N5072, N5062, N4567);
xor XOR2 (N5073, N5067, N4641);
nor NOR2 (N5074, N5071, N858);
nor NOR2 (N5075, N5064, N392);
or OR3 (N5076, N5066, N3579, N1482);
buf BUF1 (N5077, N5073);
nand NAND4 (N5078, N5072, N523, N599, N4250);
buf BUF1 (N5079, N5075);
buf BUF1 (N5080, N5070);
buf BUF1 (N5081, N5077);
not NOT1 (N5082, N5068);
buf BUF1 (N5083, N5046);
buf BUF1 (N5084, N5059);
nor NOR3 (N5085, N5079, N2261, N271);
and AND3 (N5086, N5080, N1394, N1828);
buf BUF1 (N5087, N5078);
or OR3 (N5088, N5069, N424, N4151);
nand NAND3 (N5089, N5084, N3170, N377);
nand NAND2 (N5090, N5076, N3380);
and AND2 (N5091, N5074, N4253);
nand NAND3 (N5092, N5087, N521, N2088);
nand NAND3 (N5093, N5086, N916, N59);
not NOT1 (N5094, N5085);
xor XOR2 (N5095, N5094, N1777);
or OR3 (N5096, N5091, N4571, N3959);
or OR4 (N5097, N5092, N2260, N3924, N3341);
buf BUF1 (N5098, N5096);
xor XOR2 (N5099, N5081, N1182);
buf BUF1 (N5100, N5093);
and AND4 (N5101, N5088, N4616, N2501, N2048);
and AND3 (N5102, N5090, N1770, N1122);
nand NAND4 (N5103, N5099, N967, N4852, N3309);
nand NAND3 (N5104, N5089, N3815, N4819);
nand NAND2 (N5105, N5104, N4400);
and AND2 (N5106, N5098, N1417);
and AND2 (N5107, N5103, N3994);
or OR2 (N5108, N5082, N4912);
or OR3 (N5109, N5106, N642, N3401);
xor XOR2 (N5110, N5100, N424);
and AND2 (N5111, N5083, N4734);
xor XOR2 (N5112, N5095, N3555);
not NOT1 (N5113, N5097);
and AND4 (N5114, N5105, N3657, N4908, N4737);
buf BUF1 (N5115, N5113);
not NOT1 (N5116, N5109);
nand NAND4 (N5117, N5108, N1979, N1130, N2326);
and AND2 (N5118, N5110, N2034);
buf BUF1 (N5119, N5107);
xor XOR2 (N5120, N5118, N1176);
not NOT1 (N5121, N5112);
xor XOR2 (N5122, N5121, N2372);
xor XOR2 (N5123, N5116, N4263);
nor NOR4 (N5124, N5120, N4762, N5051, N1229);
buf BUF1 (N5125, N5114);
nor NOR4 (N5126, N5101, N4242, N3348, N825);
buf BUF1 (N5127, N5125);
nand NAND3 (N5128, N5117, N1620, N777);
nor NOR4 (N5129, N5111, N630, N5015, N3887);
nor NOR2 (N5130, N5123, N533);
and AND2 (N5131, N5128, N2776);
xor XOR2 (N5132, N5124, N3527);
xor XOR2 (N5133, N5129, N2875);
nor NOR4 (N5134, N5127, N4167, N2392, N63);
not NOT1 (N5135, N5130);
or OR3 (N5136, N5135, N534, N3375);
xor XOR2 (N5137, N5132, N1171);
xor XOR2 (N5138, N5131, N2243);
buf BUF1 (N5139, N5115);
nor NOR2 (N5140, N5139, N1934);
and AND3 (N5141, N5133, N3274, N1612);
buf BUF1 (N5142, N5122);
xor XOR2 (N5143, N5138, N4488);
buf BUF1 (N5144, N5140);
and AND3 (N5145, N5134, N3070, N3004);
or OR2 (N5146, N5126, N4981);
nor NOR2 (N5147, N5119, N2014);
xor XOR2 (N5148, N5143, N2418);
not NOT1 (N5149, N5145);
and AND2 (N5150, N5136, N2045);
xor XOR2 (N5151, N5147, N3594);
buf BUF1 (N5152, N5141);
and AND2 (N5153, N5151, N4373);
or OR4 (N5154, N5150, N3398, N3781, N2838);
buf BUF1 (N5155, N5142);
and AND3 (N5156, N5137, N3569, N4556);
not NOT1 (N5157, N5144);
xor XOR2 (N5158, N5152, N2458);
buf BUF1 (N5159, N5148);
buf BUF1 (N5160, N5149);
and AND3 (N5161, N5102, N397, N3162);
nand NAND2 (N5162, N5157, N2673);
nor NOR2 (N5163, N5159, N2798);
not NOT1 (N5164, N5153);
buf BUF1 (N5165, N5163);
not NOT1 (N5166, N5158);
nand NAND2 (N5167, N5156, N4966);
or OR4 (N5168, N5161, N1189, N1382, N4328);
nor NOR4 (N5169, N5160, N4173, N3785, N2898);
and AND2 (N5170, N5167, N1547);
nand NAND4 (N5171, N5146, N3063, N2751, N2928);
buf BUF1 (N5172, N5169);
buf BUF1 (N5173, N5166);
or OR3 (N5174, N5173, N3672, N742);
or OR2 (N5175, N5164, N1374);
xor XOR2 (N5176, N5174, N1085);
not NOT1 (N5177, N5165);
and AND4 (N5178, N5168, N2920, N2181, N3607);
nor NOR3 (N5179, N5172, N125, N939);
nand NAND4 (N5180, N5178, N3611, N4530, N4985);
nand NAND2 (N5181, N5175, N3899);
not NOT1 (N5182, N5181);
nor NOR3 (N5183, N5180, N2031, N1456);
and AND2 (N5184, N5154, N1777);
not NOT1 (N5185, N5184);
nor NOR2 (N5186, N5170, N3002);
buf BUF1 (N5187, N5185);
nor NOR3 (N5188, N5171, N4728, N2308);
buf BUF1 (N5189, N5179);
and AND2 (N5190, N5177, N3105);
or OR3 (N5191, N5182, N1143, N1432);
nor NOR3 (N5192, N5190, N1856, N5063);
not NOT1 (N5193, N5162);
or OR4 (N5194, N5193, N2083, N2227, N794);
nor NOR3 (N5195, N5192, N3647, N4138);
xor XOR2 (N5196, N5176, N268);
and AND3 (N5197, N5196, N5072, N2175);
nand NAND2 (N5198, N5194, N3176);
buf BUF1 (N5199, N5197);
buf BUF1 (N5200, N5195);
not NOT1 (N5201, N5186);
nand NAND3 (N5202, N5198, N552, N4183);
xor XOR2 (N5203, N5201, N6);
and AND3 (N5204, N5155, N5124, N2583);
xor XOR2 (N5205, N5199, N3569);
xor XOR2 (N5206, N5203, N3951);
xor XOR2 (N5207, N5205, N2310);
xor XOR2 (N5208, N5188, N4262);
nor NOR4 (N5209, N5191, N3843, N3386, N2343);
buf BUF1 (N5210, N5208);
nand NAND3 (N5211, N5187, N2368, N4527);
and AND3 (N5212, N5210, N886, N3666);
not NOT1 (N5213, N5183);
nor NOR3 (N5214, N5202, N480, N3022);
xor XOR2 (N5215, N5189, N2719);
buf BUF1 (N5216, N5214);
nor NOR2 (N5217, N5204, N5040);
nand NAND3 (N5218, N5209, N4439, N3192);
xor XOR2 (N5219, N5206, N1195);
and AND4 (N5220, N5216, N2600, N661, N493);
and AND3 (N5221, N5220, N2207, N1803);
and AND4 (N5222, N5217, N1387, N3577, N3403);
not NOT1 (N5223, N5212);
buf BUF1 (N5224, N5200);
nor NOR4 (N5225, N5223, N4282, N3578, N5224);
buf BUF1 (N5226, N3024);
buf BUF1 (N5227, N5213);
xor XOR2 (N5228, N5222, N202);
nand NAND4 (N5229, N5221, N3661, N1726, N2795);
and AND2 (N5230, N5215, N4416);
not NOT1 (N5231, N5218);
nand NAND2 (N5232, N5226, N2122);
and AND4 (N5233, N5207, N269, N1044, N4799);
or OR4 (N5234, N5233, N4284, N3396, N3193);
or OR3 (N5235, N5232, N1183, N4406);
and AND2 (N5236, N5227, N1880);
nor NOR3 (N5237, N5234, N2081, N2001);
xor XOR2 (N5238, N5228, N3694);
not NOT1 (N5239, N5229);
xor XOR2 (N5240, N5237, N1498);
xor XOR2 (N5241, N5240, N489);
nor NOR4 (N5242, N5236, N5236, N2642, N1549);
xor XOR2 (N5243, N5238, N3482);
nand NAND4 (N5244, N5239, N2540, N641, N5013);
nand NAND4 (N5245, N5244, N3353, N4048, N1724);
and AND2 (N5246, N5225, N4520);
nand NAND4 (N5247, N5230, N1686, N1206, N2242);
xor XOR2 (N5248, N5247, N530);
nor NOR3 (N5249, N5245, N517, N4826);
and AND2 (N5250, N5235, N5162);
nor NOR3 (N5251, N5219, N4665, N1516);
and AND4 (N5252, N5241, N3986, N3646, N3230);
nor NOR2 (N5253, N5252, N1356);
nand NAND4 (N5254, N5250, N3633, N4845, N4669);
nor NOR3 (N5255, N5243, N3016, N2725);
not NOT1 (N5256, N5211);
nand NAND2 (N5257, N5255, N2472);
nor NOR4 (N5258, N5248, N1514, N1900, N270);
buf BUF1 (N5259, N5242);
or OR3 (N5260, N5246, N881, N2808);
nor NOR2 (N5261, N5249, N1886);
nor NOR2 (N5262, N5256, N414);
not NOT1 (N5263, N5259);
xor XOR2 (N5264, N5254, N4886);
or OR2 (N5265, N5260, N922);
and AND4 (N5266, N5264, N3957, N4032, N3636);
or OR2 (N5267, N5263, N2651);
or OR2 (N5268, N5261, N3995);
buf BUF1 (N5269, N5265);
or OR3 (N5270, N5266, N2803, N5086);
buf BUF1 (N5271, N5257);
nor NOR4 (N5272, N5269, N502, N1366, N2743);
not NOT1 (N5273, N5268);
buf BUF1 (N5274, N5272);
nand NAND3 (N5275, N5271, N4417, N870);
or OR3 (N5276, N5231, N839, N2521);
buf BUF1 (N5277, N5276);
xor XOR2 (N5278, N5258, N3839);
xor XOR2 (N5279, N5253, N1175);
not NOT1 (N5280, N5274);
and AND2 (N5281, N5270, N1449);
and AND3 (N5282, N5281, N811, N1710);
buf BUF1 (N5283, N5280);
nand NAND3 (N5284, N5267, N3769, N4512);
and AND3 (N5285, N5251, N3576, N2310);
nand NAND3 (N5286, N5282, N4854, N4716);
nor NOR2 (N5287, N5275, N1228);
nor NOR4 (N5288, N5279, N2254, N3075, N4867);
not NOT1 (N5289, N5277);
nor NOR3 (N5290, N5286, N4712, N2154);
or OR4 (N5291, N5284, N2674, N3998, N5186);
and AND3 (N5292, N5287, N3008, N2640);
xor XOR2 (N5293, N5289, N3534);
xor XOR2 (N5294, N5273, N812);
nand NAND2 (N5295, N5293, N4260);
or OR3 (N5296, N5288, N2273, N4631);
or OR2 (N5297, N5296, N2586);
not NOT1 (N5298, N5291);
xor XOR2 (N5299, N5295, N2670);
nand NAND2 (N5300, N5285, N5229);
not NOT1 (N5301, N5298);
nor NOR4 (N5302, N5290, N2324, N1281, N3916);
not NOT1 (N5303, N5292);
buf BUF1 (N5304, N5262);
nor NOR3 (N5305, N5302, N5237, N4389);
or OR3 (N5306, N5301, N398, N2752);
or OR4 (N5307, N5299, N805, N3165, N507);
nand NAND3 (N5308, N5304, N2797, N4533);
or OR4 (N5309, N5300, N2075, N4053, N1624);
and AND2 (N5310, N5297, N3683);
and AND3 (N5311, N5306, N2705, N1872);
and AND2 (N5312, N5309, N2775);
not NOT1 (N5313, N5278);
not NOT1 (N5314, N5313);
not NOT1 (N5315, N5303);
buf BUF1 (N5316, N5314);
and AND4 (N5317, N5294, N2182, N3451, N4330);
nor NOR2 (N5318, N5310, N2035);
buf BUF1 (N5319, N5318);
not NOT1 (N5320, N5307);
buf BUF1 (N5321, N5320);
nor NOR4 (N5322, N5315, N3074, N4793, N4323);
nor NOR4 (N5323, N5317, N2476, N2818, N3411);
nand NAND2 (N5324, N5322, N3500);
buf BUF1 (N5325, N5324);
xor XOR2 (N5326, N5312, N2827);
xor XOR2 (N5327, N5311, N1631);
buf BUF1 (N5328, N5319);
or OR3 (N5329, N5328, N199, N84);
not NOT1 (N5330, N5323);
nand NAND2 (N5331, N5330, N2680);
and AND2 (N5332, N5308, N779);
buf BUF1 (N5333, N5326);
or OR3 (N5334, N5331, N5, N2442);
buf BUF1 (N5335, N5334);
nand NAND4 (N5336, N5283, N1098, N1311, N2751);
xor XOR2 (N5337, N5329, N1538);
not NOT1 (N5338, N5337);
buf BUF1 (N5339, N5305);
not NOT1 (N5340, N5339);
or OR4 (N5341, N5336, N1525, N2124, N3185);
buf BUF1 (N5342, N5325);
nand NAND2 (N5343, N5333, N3526);
or OR4 (N5344, N5343, N3357, N1449, N4524);
nand NAND4 (N5345, N5338, N381, N288, N3029);
nor NOR2 (N5346, N5345, N627);
xor XOR2 (N5347, N5342, N2743);
nor NOR2 (N5348, N5335, N4819);
xor XOR2 (N5349, N5327, N4651);
nand NAND3 (N5350, N5347, N5091, N4658);
buf BUF1 (N5351, N5340);
nand NAND3 (N5352, N5341, N3283, N4246);
nand NAND2 (N5353, N5316, N1076);
or OR4 (N5354, N5349, N1218, N5145, N2902);
nand NAND4 (N5355, N5321, N4372, N1141, N55);
or OR2 (N5356, N5346, N548);
or OR3 (N5357, N5344, N3299, N1725);
nand NAND3 (N5358, N5352, N2896, N153);
not NOT1 (N5359, N5332);
buf BUF1 (N5360, N5348);
xor XOR2 (N5361, N5360, N673);
and AND2 (N5362, N5351, N2708);
not NOT1 (N5363, N5355);
or OR3 (N5364, N5354, N974, N985);
and AND2 (N5365, N5364, N894);
or OR4 (N5366, N5356, N478, N969, N1738);
xor XOR2 (N5367, N5358, N77);
xor XOR2 (N5368, N5359, N2669);
nor NOR3 (N5369, N5353, N5323, N3428);
buf BUF1 (N5370, N5362);
or OR4 (N5371, N5357, N4023, N4013, N329);
buf BUF1 (N5372, N5361);
or OR3 (N5373, N5369, N55, N1314);
nand NAND4 (N5374, N5372, N2516, N4254, N1491);
not NOT1 (N5375, N5365);
nor NOR2 (N5376, N5370, N387);
nand NAND4 (N5377, N5368, N1278, N4011, N163);
or OR4 (N5378, N5374, N405, N3651, N4645);
nor NOR3 (N5379, N5367, N2245, N1429);
nand NAND4 (N5380, N5375, N5085, N2359, N4856);
xor XOR2 (N5381, N5371, N493);
not NOT1 (N5382, N5376);
nor NOR3 (N5383, N5382, N2062, N2309);
not NOT1 (N5384, N5380);
nor NOR3 (N5385, N5373, N3071, N361);
buf BUF1 (N5386, N5363);
buf BUF1 (N5387, N5381);
and AND2 (N5388, N5386, N818);
nor NOR3 (N5389, N5385, N1646, N63);
nor NOR3 (N5390, N5366, N166, N2385);
nor NOR3 (N5391, N5389, N3577, N2714);
nand NAND3 (N5392, N5383, N993, N1689);
nor NOR2 (N5393, N5377, N2270);
not NOT1 (N5394, N5391);
and AND2 (N5395, N5350, N2044);
buf BUF1 (N5396, N5394);
nand NAND4 (N5397, N5379, N4834, N857, N3063);
nor NOR3 (N5398, N5387, N5258, N3554);
not NOT1 (N5399, N5397);
and AND2 (N5400, N5396, N1182);
nand NAND2 (N5401, N5398, N1365);
xor XOR2 (N5402, N5395, N380);
and AND4 (N5403, N5392, N1614, N145, N1344);
nand NAND3 (N5404, N5388, N3244, N1606);
not NOT1 (N5405, N5403);
xor XOR2 (N5406, N5399, N1317);
and AND3 (N5407, N5406, N3086, N1391);
buf BUF1 (N5408, N5407);
nand NAND4 (N5409, N5393, N2031, N5402, N1644);
xor XOR2 (N5410, N742, N3434);
xor XOR2 (N5411, N5378, N3376);
nand NAND3 (N5412, N5408, N3725, N2594);
not NOT1 (N5413, N5409);
buf BUF1 (N5414, N5413);
nand NAND4 (N5415, N5384, N3985, N3846, N3228);
or OR3 (N5416, N5390, N70, N4844);
buf BUF1 (N5417, N5405);
nor NOR4 (N5418, N5416, N5226, N1356, N1771);
buf BUF1 (N5419, N5417);
and AND3 (N5420, N5415, N2332, N72);
not NOT1 (N5421, N5418);
and AND3 (N5422, N5419, N1548, N2751);
buf BUF1 (N5423, N5410);
xor XOR2 (N5424, N5420, N1246);
not NOT1 (N5425, N5401);
or OR3 (N5426, N5424, N2269, N3735);
xor XOR2 (N5427, N5411, N5276);
nand NAND2 (N5428, N5426, N3498);
or OR3 (N5429, N5422, N1241, N3983);
or OR2 (N5430, N5421, N3868);
nor NOR2 (N5431, N5414, N1478);
xor XOR2 (N5432, N5412, N3459);
and AND3 (N5433, N5427, N5120, N5073);
xor XOR2 (N5434, N5425, N1481);
nor NOR2 (N5435, N5433, N3916);
xor XOR2 (N5436, N5423, N1408);
nor NOR3 (N5437, N5431, N3919, N3664);
nand NAND4 (N5438, N5434, N2729, N696, N3262);
and AND2 (N5439, N5435, N860);
buf BUF1 (N5440, N5436);
not NOT1 (N5441, N5404);
xor XOR2 (N5442, N5400, N4035);
not NOT1 (N5443, N5440);
nand NAND4 (N5444, N5430, N332, N5012, N5140);
or OR4 (N5445, N5432, N5068, N2904, N2921);
nor NOR4 (N5446, N5441, N2761, N1985, N3254);
buf BUF1 (N5447, N5439);
and AND3 (N5448, N5447, N3955, N4289);
not NOT1 (N5449, N5438);
nor NOR2 (N5450, N5442, N715);
not NOT1 (N5451, N5448);
nand NAND4 (N5452, N5443, N4108, N2260, N5412);
nor NOR4 (N5453, N5429, N3271, N2403, N1518);
nor NOR3 (N5454, N5452, N5413, N1511);
or OR2 (N5455, N5428, N3403);
and AND4 (N5456, N5437, N130, N4531, N3069);
nand NAND4 (N5457, N5450, N2422, N604, N265);
xor XOR2 (N5458, N5449, N4420);
not NOT1 (N5459, N5457);
not NOT1 (N5460, N5458);
buf BUF1 (N5461, N5460);
nand NAND2 (N5462, N5456, N3968);
xor XOR2 (N5463, N5446, N3564);
nand NAND4 (N5464, N5444, N1337, N4669, N4881);
or OR4 (N5465, N5464, N1879, N3263, N4914);
buf BUF1 (N5466, N5459);
and AND4 (N5467, N5451, N961, N644, N1564);
xor XOR2 (N5468, N5463, N4494);
not NOT1 (N5469, N5454);
buf BUF1 (N5470, N5465);
nand NAND4 (N5471, N5470, N4034, N5202, N3993);
or OR2 (N5472, N5462, N4832);
and AND3 (N5473, N5466, N4447, N1255);
nand NAND3 (N5474, N5469, N3961, N2101);
xor XOR2 (N5475, N5472, N5058);
not NOT1 (N5476, N5473);
nand NAND2 (N5477, N5475, N3607);
or OR2 (N5478, N5467, N2785);
nor NOR2 (N5479, N5453, N1895);
nand NAND3 (N5480, N5445, N1180, N2755);
nor NOR3 (N5481, N5468, N804, N114);
or OR2 (N5482, N5474, N1741);
buf BUF1 (N5483, N5476);
buf BUF1 (N5484, N5480);
nand NAND4 (N5485, N5461, N3116, N2771, N567);
or OR4 (N5486, N5483, N1452, N2314, N3137);
not NOT1 (N5487, N5471);
or OR4 (N5488, N5481, N369, N4315, N5432);
buf BUF1 (N5489, N5477);
or OR2 (N5490, N5484, N3206);
not NOT1 (N5491, N5486);
and AND3 (N5492, N5489, N2646, N3867);
nand NAND4 (N5493, N5488, N164, N1354, N3489);
xor XOR2 (N5494, N5491, N4713);
nand NAND4 (N5495, N5455, N142, N1359, N1645);
or OR4 (N5496, N5487, N3949, N616, N4445);
and AND2 (N5497, N5490, N1531);
buf BUF1 (N5498, N5493);
and AND4 (N5499, N5494, N5097, N2017, N5184);
buf BUF1 (N5500, N5498);
or OR3 (N5501, N5478, N2770, N4661);
not NOT1 (N5502, N5499);
nor NOR4 (N5503, N5496, N246, N5222, N3744);
nand NAND4 (N5504, N5503, N2715, N1974, N4983);
and AND4 (N5505, N5501, N5202, N1337, N81);
not NOT1 (N5506, N5495);
and AND2 (N5507, N5506, N735);
xor XOR2 (N5508, N5502, N4546);
nor NOR2 (N5509, N5505, N4240);
buf BUF1 (N5510, N5492);
nand NAND4 (N5511, N5497, N4350, N2408, N4986);
not NOT1 (N5512, N5508);
buf BUF1 (N5513, N5482);
buf BUF1 (N5514, N5511);
and AND4 (N5515, N5500, N265, N2776, N5181);
nor NOR4 (N5516, N5513, N3742, N3565, N5313);
nor NOR3 (N5517, N5515, N849, N1998);
buf BUF1 (N5518, N5510);
nand NAND2 (N5519, N5507, N5007);
not NOT1 (N5520, N5519);
not NOT1 (N5521, N5512);
xor XOR2 (N5522, N5518, N3136);
nor NOR2 (N5523, N5522, N4767);
and AND3 (N5524, N5514, N2060, N4774);
nand NAND3 (N5525, N5520, N4450, N2805);
buf BUF1 (N5526, N5504);
nor NOR3 (N5527, N5524, N939, N1210);
and AND4 (N5528, N5527, N3834, N1923, N5328);
not NOT1 (N5529, N5526);
or OR4 (N5530, N5517, N1729, N4909, N1219);
not NOT1 (N5531, N5530);
or OR2 (N5532, N5531, N4668);
xor XOR2 (N5533, N5532, N3551);
buf BUF1 (N5534, N5516);
nand NAND4 (N5535, N5479, N2855, N5031, N1517);
and AND3 (N5536, N5535, N1740, N1555);
nand NAND2 (N5537, N5523, N5075);
xor XOR2 (N5538, N5536, N940);
xor XOR2 (N5539, N5521, N2699);
xor XOR2 (N5540, N5534, N124);
nand NAND4 (N5541, N5525, N3545, N1376, N880);
nor NOR2 (N5542, N5485, N2692);
buf BUF1 (N5543, N5540);
nand NAND3 (N5544, N5509, N4548, N1838);
not NOT1 (N5545, N5529);
xor XOR2 (N5546, N5539, N1236);
not NOT1 (N5547, N5537);
nor NOR3 (N5548, N5542, N5403, N2910);
buf BUF1 (N5549, N5538);
buf BUF1 (N5550, N5548);
and AND4 (N5551, N5541, N4589, N722, N195);
nand NAND2 (N5552, N5550, N3002);
xor XOR2 (N5553, N5545, N4474);
and AND3 (N5554, N5533, N3089, N4859);
nor NOR2 (N5555, N5552, N2881);
buf BUF1 (N5556, N5543);
or OR3 (N5557, N5551, N3653, N3981);
not NOT1 (N5558, N5549);
nand NAND2 (N5559, N5553, N3816);
xor XOR2 (N5560, N5559, N1519);
not NOT1 (N5561, N5547);
nor NOR2 (N5562, N5560, N1151);
nand NAND3 (N5563, N5561, N4476, N1917);
or OR4 (N5564, N5562, N303, N5274, N4864);
buf BUF1 (N5565, N5528);
nand NAND3 (N5566, N5558, N5023, N5486);
and AND4 (N5567, N5544, N3901, N1305, N4721);
not NOT1 (N5568, N5567);
nor NOR2 (N5569, N5556, N2796);
xor XOR2 (N5570, N5568, N4608);
buf BUF1 (N5571, N5554);
nand NAND3 (N5572, N5565, N3544, N1128);
and AND2 (N5573, N5569, N4861);
and AND3 (N5574, N5555, N5325, N2390);
and AND4 (N5575, N5563, N3926, N4551, N2470);
or OR2 (N5576, N5575, N428);
xor XOR2 (N5577, N5566, N230);
and AND2 (N5578, N5574, N4701);
and AND2 (N5579, N5573, N3350);
nor NOR4 (N5580, N5570, N5576, N219, N353);
or OR4 (N5581, N5435, N906, N5569, N5351);
and AND2 (N5582, N5557, N3421);
not NOT1 (N5583, N5578);
xor XOR2 (N5584, N5571, N5300);
buf BUF1 (N5585, N5546);
nor NOR4 (N5586, N5572, N5301, N5502, N634);
xor XOR2 (N5587, N5584, N2537);
and AND2 (N5588, N5583, N5240);
not NOT1 (N5589, N5564);
nor NOR3 (N5590, N5580, N2945, N4054);
or OR4 (N5591, N5586, N2230, N2850, N3352);
nand NAND4 (N5592, N5588, N2277, N5231, N1941);
nor NOR2 (N5593, N5585, N899);
or OR2 (N5594, N5581, N2434);
not NOT1 (N5595, N5594);
xor XOR2 (N5596, N5582, N3698);
xor XOR2 (N5597, N5591, N3220);
not NOT1 (N5598, N5587);
not NOT1 (N5599, N5579);
buf BUF1 (N5600, N5596);
and AND3 (N5601, N5597, N5377, N1112);
xor XOR2 (N5602, N5593, N1236);
xor XOR2 (N5603, N5602, N3769);
or OR4 (N5604, N5603, N942, N2736, N2052);
or OR2 (N5605, N5590, N5099);
not NOT1 (N5606, N5600);
nand NAND3 (N5607, N5577, N327, N3173);
and AND4 (N5608, N5589, N3047, N2883, N635);
or OR3 (N5609, N5598, N3281, N3081);
and AND4 (N5610, N5595, N3078, N706, N5442);
nand NAND2 (N5611, N5607, N4524);
xor XOR2 (N5612, N5592, N4186);
nand NAND4 (N5613, N5606, N3547, N4193, N2516);
and AND4 (N5614, N5613, N2212, N267, N3645);
or OR2 (N5615, N5610, N4936);
or OR2 (N5616, N5608, N2973);
nand NAND3 (N5617, N5615, N1114, N1608);
or OR4 (N5618, N5612, N341, N745, N3094);
xor XOR2 (N5619, N5605, N3476);
nor NOR4 (N5620, N5609, N1721, N1412, N1204);
or OR2 (N5621, N5614, N5187);
buf BUF1 (N5622, N5619);
and AND2 (N5623, N5617, N235);
or OR4 (N5624, N5611, N3940, N1379, N2151);
not NOT1 (N5625, N5624);
nor NOR3 (N5626, N5618, N4409, N3946);
nand NAND4 (N5627, N5620, N553, N1017, N1545);
nor NOR2 (N5628, N5626, N5168);
nand NAND3 (N5629, N5621, N4574, N5324);
and AND3 (N5630, N5629, N389, N2757);
buf BUF1 (N5631, N5616);
xor XOR2 (N5632, N5625, N3335);
nor NOR3 (N5633, N5604, N194, N3001);
nor NOR3 (N5634, N5601, N3287, N1242);
and AND3 (N5635, N5628, N39, N832);
xor XOR2 (N5636, N5623, N4464);
nor NOR2 (N5637, N5633, N2336);
and AND2 (N5638, N5637, N1736);
not NOT1 (N5639, N5635);
and AND2 (N5640, N5627, N4131);
nand NAND4 (N5641, N5622, N706, N389, N4393);
and AND3 (N5642, N5639, N3547, N961);
nand NAND2 (N5643, N5640, N3832);
not NOT1 (N5644, N5643);
or OR4 (N5645, N5642, N4966, N911, N4397);
nor NOR2 (N5646, N5634, N627);
not NOT1 (N5647, N5636);
or OR2 (N5648, N5638, N2353);
nor NOR3 (N5649, N5632, N4788, N78);
xor XOR2 (N5650, N5641, N1217);
or OR4 (N5651, N5650, N2600, N3639, N633);
buf BUF1 (N5652, N5647);
nand NAND2 (N5653, N5644, N5635);
or OR2 (N5654, N5645, N776);
nor NOR2 (N5655, N5651, N2612);
xor XOR2 (N5656, N5631, N1550);
or OR4 (N5657, N5646, N3646, N5561, N1267);
xor XOR2 (N5658, N5657, N2510);
and AND2 (N5659, N5653, N2928);
nand NAND3 (N5660, N5630, N3915, N339);
or OR3 (N5661, N5652, N4931, N4720);
xor XOR2 (N5662, N5658, N726);
or OR3 (N5663, N5662, N1791, N4056);
and AND4 (N5664, N5655, N4421, N3129, N1156);
and AND2 (N5665, N5649, N58);
nand NAND4 (N5666, N5661, N4363, N1258, N947);
nand NAND2 (N5667, N5648, N3237);
or OR2 (N5668, N5654, N1101);
nand NAND3 (N5669, N5665, N438, N701);
nand NAND3 (N5670, N5659, N2993, N1982);
xor XOR2 (N5671, N5670, N1224);
or OR3 (N5672, N5599, N3475, N1726);
xor XOR2 (N5673, N5668, N665);
not NOT1 (N5674, N5667);
or OR4 (N5675, N5663, N199, N3216, N1699);
or OR4 (N5676, N5660, N1694, N4802, N4167);
xor XOR2 (N5677, N5675, N3809);
nor NOR4 (N5678, N5677, N824, N417, N261);
and AND4 (N5679, N5669, N277, N1133, N2664);
buf BUF1 (N5680, N5674);
or OR3 (N5681, N5664, N1582, N4493);
nand NAND2 (N5682, N5672, N1631);
not NOT1 (N5683, N5681);
not NOT1 (N5684, N5671);
or OR4 (N5685, N5656, N4349, N5663, N4675);
not NOT1 (N5686, N5684);
not NOT1 (N5687, N5673);
not NOT1 (N5688, N5686);
nor NOR4 (N5689, N5683, N979, N5376, N2334);
nand NAND4 (N5690, N5689, N5113, N4201, N2696);
or OR4 (N5691, N5679, N4588, N4076, N5241);
and AND3 (N5692, N5680, N2584, N1510);
nor NOR3 (N5693, N5682, N4183, N573);
nor NOR4 (N5694, N5666, N1727, N2297, N4204);
buf BUF1 (N5695, N5694);
not NOT1 (N5696, N5676);
xor XOR2 (N5697, N5691, N3721);
nor NOR3 (N5698, N5690, N4985, N4605);
nand NAND2 (N5699, N5693, N1136);
buf BUF1 (N5700, N5685);
nor NOR2 (N5701, N5700, N5513);
or OR3 (N5702, N5698, N4560, N2815);
not NOT1 (N5703, N5692);
nor NOR2 (N5704, N5687, N1105);
and AND4 (N5705, N5704, N5066, N3502, N5114);
and AND2 (N5706, N5696, N1686);
nor NOR2 (N5707, N5702, N177);
and AND4 (N5708, N5706, N3866, N5266, N5336);
nand NAND3 (N5709, N5697, N604, N5127);
and AND3 (N5710, N5709, N4271, N3495);
nor NOR4 (N5711, N5695, N2057, N1468, N1719);
and AND2 (N5712, N5705, N5285);
or OR4 (N5713, N5707, N4894, N5573, N30);
not NOT1 (N5714, N5712);
nor NOR2 (N5715, N5708, N5491);
not NOT1 (N5716, N5678);
buf BUF1 (N5717, N5699);
not NOT1 (N5718, N5717);
not NOT1 (N5719, N5703);
or OR4 (N5720, N5718, N707, N1960, N5152);
nand NAND4 (N5721, N5713, N3035, N4819, N2006);
and AND2 (N5722, N5721, N1709);
nor NOR3 (N5723, N5710, N231, N4103);
or OR4 (N5724, N5723, N4782, N3902, N2387);
nand NAND4 (N5725, N5722, N1142, N1141, N689);
nor NOR2 (N5726, N5711, N2420);
nor NOR2 (N5727, N5725, N4517);
and AND4 (N5728, N5715, N2407, N2461, N5280);
nor NOR3 (N5729, N5720, N1389, N4032);
buf BUF1 (N5730, N5726);
nand NAND2 (N5731, N5728, N1885);
and AND2 (N5732, N5731, N1278);
or OR2 (N5733, N5719, N1130);
or OR3 (N5734, N5714, N4973, N1100);
xor XOR2 (N5735, N5732, N5724);
nand NAND3 (N5736, N4605, N1511, N477);
xor XOR2 (N5737, N5729, N4182);
xor XOR2 (N5738, N5733, N156);
and AND3 (N5739, N5734, N5399, N869);
and AND4 (N5740, N5736, N71, N2561, N41);
or OR3 (N5741, N5688, N1586, N5480);
nand NAND3 (N5742, N5737, N2833, N331);
and AND2 (N5743, N5740, N2267);
and AND4 (N5744, N5743, N1494, N2504, N5405);
nand NAND2 (N5745, N5744, N4165);
buf BUF1 (N5746, N5745);
and AND4 (N5747, N5746, N4417, N4527, N2079);
and AND3 (N5748, N5747, N3072, N2303);
xor XOR2 (N5749, N5735, N4903);
not NOT1 (N5750, N5716);
xor XOR2 (N5751, N5730, N222);
nor NOR3 (N5752, N5738, N4669, N1654);
nand NAND3 (N5753, N5727, N1328, N3249);
not NOT1 (N5754, N5741);
nor NOR2 (N5755, N5754, N4157);
or OR3 (N5756, N5755, N3101, N2690);
buf BUF1 (N5757, N5753);
nand NAND2 (N5758, N5752, N2822);
not NOT1 (N5759, N5742);
and AND2 (N5760, N5759, N4528);
or OR2 (N5761, N5758, N2409);
nand NAND4 (N5762, N5756, N5749, N2997, N2793);
or OR2 (N5763, N2122, N1261);
or OR2 (N5764, N5701, N2714);
not NOT1 (N5765, N5760);
buf BUF1 (N5766, N5761);
nor NOR3 (N5767, N5762, N511, N4680);
or OR4 (N5768, N5748, N1288, N2831, N5080);
buf BUF1 (N5769, N5757);
not NOT1 (N5770, N5768);
buf BUF1 (N5771, N5769);
xor XOR2 (N5772, N5767, N3555);
nor NOR2 (N5773, N5751, N2297);
buf BUF1 (N5774, N5771);
xor XOR2 (N5775, N5750, N293);
buf BUF1 (N5776, N5739);
xor XOR2 (N5777, N5773, N3858);
not NOT1 (N5778, N5764);
or OR3 (N5779, N5772, N1121, N1899);
and AND4 (N5780, N5778, N1518, N2225, N3057);
or OR4 (N5781, N5776, N1907, N3920, N3787);
not NOT1 (N5782, N5777);
buf BUF1 (N5783, N5774);
nor NOR4 (N5784, N5766, N2453, N873, N5331);
not NOT1 (N5785, N5775);
nor NOR4 (N5786, N5779, N2648, N2621, N3015);
xor XOR2 (N5787, N5784, N4615);
xor XOR2 (N5788, N5785, N223);
or OR3 (N5789, N5782, N4139, N3514);
nor NOR3 (N5790, N5786, N4009, N4052);
xor XOR2 (N5791, N5780, N1945);
or OR2 (N5792, N5783, N4683);
not NOT1 (N5793, N5770);
nand NAND2 (N5794, N5790, N495);
nand NAND2 (N5795, N5787, N5505);
buf BUF1 (N5796, N5763);
xor XOR2 (N5797, N5795, N5352);
nand NAND3 (N5798, N5789, N110, N2984);
xor XOR2 (N5799, N5797, N96);
nor NOR2 (N5800, N5792, N1312);
buf BUF1 (N5801, N5765);
buf BUF1 (N5802, N5796);
or OR4 (N5803, N5788, N821, N2941, N4700);
and AND3 (N5804, N5794, N5380, N4750);
and AND2 (N5805, N5798, N1804);
xor XOR2 (N5806, N5804, N3305);
xor XOR2 (N5807, N5805, N1337);
buf BUF1 (N5808, N5803);
buf BUF1 (N5809, N5807);
buf BUF1 (N5810, N5793);
or OR3 (N5811, N5801, N11, N2877);
nand NAND2 (N5812, N5781, N5188);
not NOT1 (N5813, N5811);
not NOT1 (N5814, N5791);
nand NAND3 (N5815, N5802, N2407, N1445);
not NOT1 (N5816, N5815);
or OR2 (N5817, N5808, N1689);
nor NOR3 (N5818, N5816, N853, N246);
or OR3 (N5819, N5812, N542, N319);
not NOT1 (N5820, N5814);
or OR3 (N5821, N5799, N4456, N1757);
not NOT1 (N5822, N5809);
nor NOR3 (N5823, N5800, N4126, N3140);
and AND3 (N5824, N5817, N4712, N3579);
xor XOR2 (N5825, N5821, N4277);
or OR2 (N5826, N5813, N2853);
nor NOR2 (N5827, N5806, N2929);
xor XOR2 (N5828, N5824, N1511);
nand NAND4 (N5829, N5810, N1975, N1556, N5377);
not NOT1 (N5830, N5827);
buf BUF1 (N5831, N5819);
buf BUF1 (N5832, N5825);
not NOT1 (N5833, N5826);
or OR2 (N5834, N5818, N47);
xor XOR2 (N5835, N5823, N781);
or OR2 (N5836, N5829, N1817);
nor NOR4 (N5837, N5836, N5381, N3063, N1294);
xor XOR2 (N5838, N5831, N5728);
buf BUF1 (N5839, N5837);
or OR3 (N5840, N5830, N2790, N3000);
and AND2 (N5841, N5835, N2102);
not NOT1 (N5842, N5839);
xor XOR2 (N5843, N5838, N3690);
nor NOR2 (N5844, N5820, N773);
or OR4 (N5845, N5832, N2691, N147, N468);
nor NOR3 (N5846, N5833, N4352, N4050);
nand NAND3 (N5847, N5845, N3550, N5666);
and AND3 (N5848, N5828, N4943, N2022);
nand NAND4 (N5849, N5822, N2269, N1229, N4195);
xor XOR2 (N5850, N5849, N3629);
nor NOR4 (N5851, N5842, N4192, N2302, N3826);
and AND2 (N5852, N5840, N1639);
buf BUF1 (N5853, N5843);
or OR3 (N5854, N5852, N1153, N883);
xor XOR2 (N5855, N5851, N984);
nor NOR3 (N5856, N5848, N2598, N3766);
not NOT1 (N5857, N5850);
or OR4 (N5858, N5854, N602, N4700, N5375);
or OR2 (N5859, N5858, N1183);
or OR2 (N5860, N5857, N1620);
not NOT1 (N5861, N5841);
xor XOR2 (N5862, N5860, N2738);
buf BUF1 (N5863, N5861);
and AND4 (N5864, N5847, N2289, N978, N5452);
not NOT1 (N5865, N5859);
or OR3 (N5866, N5856, N489, N338);
buf BUF1 (N5867, N5853);
nand NAND2 (N5868, N5866, N438);
nor NOR2 (N5869, N5867, N824);
xor XOR2 (N5870, N5863, N3446);
not NOT1 (N5871, N5846);
xor XOR2 (N5872, N5855, N5457);
nor NOR4 (N5873, N5864, N4894, N2661, N888);
nor NOR2 (N5874, N5834, N2268);
nand NAND4 (N5875, N5870, N4211, N2461, N4786);
or OR3 (N5876, N5868, N3314, N2274);
nor NOR4 (N5877, N5872, N256, N3279, N3923);
nand NAND3 (N5878, N5876, N3949, N2905);
buf BUF1 (N5879, N5873);
or OR2 (N5880, N5869, N3126);
buf BUF1 (N5881, N5862);
buf BUF1 (N5882, N5877);
buf BUF1 (N5883, N5880);
nand NAND3 (N5884, N5875, N3333, N4891);
xor XOR2 (N5885, N5881, N1105);
nor NOR4 (N5886, N5882, N2325, N3950, N872);
xor XOR2 (N5887, N5879, N1430);
nor NOR4 (N5888, N5886, N5210, N4011, N3412);
or OR3 (N5889, N5844, N1218, N4652);
nor NOR4 (N5890, N5888, N3796, N909, N1514);
nand NAND4 (N5891, N5884, N3348, N3371, N2141);
xor XOR2 (N5892, N5891, N4789);
nor NOR3 (N5893, N5889, N2896, N124);
or OR4 (N5894, N5883, N5508, N3655, N3776);
nor NOR4 (N5895, N5871, N5288, N596, N4195);
and AND3 (N5896, N5887, N3755, N1621);
or OR2 (N5897, N5895, N897);
and AND2 (N5898, N5897, N1596);
or OR4 (N5899, N5874, N2961, N2911, N2524);
nor NOR3 (N5900, N5898, N1348, N4319);
xor XOR2 (N5901, N5890, N5739);
buf BUF1 (N5902, N5865);
or OR3 (N5903, N5896, N3445, N3914);
buf BUF1 (N5904, N5892);
xor XOR2 (N5905, N5900, N5676);
buf BUF1 (N5906, N5893);
nand NAND4 (N5907, N5878, N2296, N3251, N4469);
or OR3 (N5908, N5899, N4712, N384);
xor XOR2 (N5909, N5906, N5740);
not NOT1 (N5910, N5885);
buf BUF1 (N5911, N5904);
nor NOR2 (N5912, N5902, N2);
and AND3 (N5913, N5894, N65, N2389);
or OR4 (N5914, N5908, N5860, N3978, N4999);
buf BUF1 (N5915, N5907);
nand NAND3 (N5916, N5915, N3169, N3093);
nor NOR2 (N5917, N5901, N1246);
and AND3 (N5918, N5910, N4040, N1693);
and AND4 (N5919, N5916, N1289, N4875, N3284);
xor XOR2 (N5920, N5909, N5214);
and AND3 (N5921, N5912, N3020, N2648);
buf BUF1 (N5922, N5913);
not NOT1 (N5923, N5903);
and AND4 (N5924, N5923, N5278, N5057, N2354);
not NOT1 (N5925, N5917);
buf BUF1 (N5926, N5905);
xor XOR2 (N5927, N5924, N2866);
buf BUF1 (N5928, N5926);
and AND2 (N5929, N5918, N2730);
nor NOR4 (N5930, N5919, N3665, N2419, N2686);
or OR3 (N5931, N5920, N109, N3496);
and AND2 (N5932, N5922, N4297);
nand NAND4 (N5933, N5932, N702, N3437, N2606);
nand NAND3 (N5934, N5928, N5896, N1493);
or OR2 (N5935, N5921, N1255);
buf BUF1 (N5936, N5925);
and AND4 (N5937, N5934, N4722, N2792, N5812);
nand NAND4 (N5938, N5929, N769, N3542, N1250);
nand NAND4 (N5939, N5938, N607, N4195, N2020);
or OR4 (N5940, N5930, N832, N2385, N3199);
or OR2 (N5941, N5911, N2037);
xor XOR2 (N5942, N5940, N3301);
xor XOR2 (N5943, N5936, N3524);
or OR2 (N5944, N5931, N4310);
xor XOR2 (N5945, N5944, N1054);
or OR3 (N5946, N5943, N529, N965);
nand NAND3 (N5947, N5942, N1302, N2500);
not NOT1 (N5948, N5937);
not NOT1 (N5949, N5946);
and AND4 (N5950, N5933, N125, N4009, N3223);
or OR2 (N5951, N5914, N4678);
not NOT1 (N5952, N5941);
buf BUF1 (N5953, N5952);
nor NOR2 (N5954, N5949, N4775);
nor NOR3 (N5955, N5935, N2841, N4526);
nand NAND4 (N5956, N5954, N125, N3644, N3709);
nor NOR2 (N5957, N5951, N1563);
nor NOR2 (N5958, N5945, N3565);
xor XOR2 (N5959, N5939, N4085);
buf BUF1 (N5960, N5957);
nand NAND3 (N5961, N5955, N5350, N2225);
and AND4 (N5962, N5959, N486, N5920, N5762);
not NOT1 (N5963, N5956);
not NOT1 (N5964, N5948);
not NOT1 (N5965, N5958);
and AND2 (N5966, N5953, N1324);
buf BUF1 (N5967, N5965);
or OR3 (N5968, N5966, N4609, N2984);
not NOT1 (N5969, N5960);
xor XOR2 (N5970, N5969, N3280);
not NOT1 (N5971, N5950);
buf BUF1 (N5972, N5962);
nor NOR4 (N5973, N5968, N4374, N2408, N2810);
nor NOR4 (N5974, N5961, N234, N1902, N1023);
nor NOR3 (N5975, N5972, N3429, N2816);
or OR3 (N5976, N5970, N3925, N2082);
nand NAND3 (N5977, N5974, N3607, N1570);
xor XOR2 (N5978, N5967, N5207);
buf BUF1 (N5979, N5927);
and AND4 (N5980, N5976, N365, N2119, N4066);
nand NAND4 (N5981, N5963, N410, N451, N4535);
xor XOR2 (N5982, N5980, N5469);
nand NAND3 (N5983, N5978, N5936, N5724);
xor XOR2 (N5984, N5979, N4927);
or OR2 (N5985, N5977, N640);
xor XOR2 (N5986, N5975, N3748);
or OR3 (N5987, N5947, N3705, N3368);
xor XOR2 (N5988, N5983, N5010);
not NOT1 (N5989, N5973);
nor NOR3 (N5990, N5971, N938, N1874);
buf BUF1 (N5991, N5989);
and AND4 (N5992, N5985, N29, N5058, N1997);
and AND4 (N5993, N5986, N1899, N147, N3116);
nand NAND3 (N5994, N5993, N3767, N4536);
buf BUF1 (N5995, N5981);
not NOT1 (N5996, N5987);
not NOT1 (N5997, N5988);
nand NAND4 (N5998, N5991, N1114, N659, N2815);
nor NOR2 (N5999, N5982, N3641);
or OR2 (N6000, N5999, N809);
not NOT1 (N6001, N5995);
and AND2 (N6002, N6001, N533);
buf BUF1 (N6003, N5990);
not NOT1 (N6004, N5996);
and AND2 (N6005, N5992, N2238);
nor NOR2 (N6006, N6005, N4722);
nor NOR2 (N6007, N6000, N3315);
not NOT1 (N6008, N6007);
and AND3 (N6009, N6004, N3221, N4537);
and AND2 (N6010, N6008, N3133);
or OR3 (N6011, N6010, N4059, N3277);
nor NOR4 (N6012, N5964, N145, N697, N5661);
and AND3 (N6013, N5998, N3702, N5282);
buf BUF1 (N6014, N6012);
not NOT1 (N6015, N5994);
nor NOR3 (N6016, N6002, N3726, N1513);
and AND4 (N6017, N6013, N5703, N4582, N2043);
xor XOR2 (N6018, N6009, N2601);
or OR3 (N6019, N6015, N2036, N3591);
nand NAND4 (N6020, N6018, N5167, N2913, N3345);
xor XOR2 (N6021, N6020, N2145);
xor XOR2 (N6022, N6021, N4569);
not NOT1 (N6023, N6014);
nor NOR2 (N6024, N6011, N3993);
xor XOR2 (N6025, N6017, N2740);
not NOT1 (N6026, N6022);
or OR3 (N6027, N6003, N1767, N3591);
nand NAND3 (N6028, N6026, N134, N1969);
or OR2 (N6029, N6019, N3088);
buf BUF1 (N6030, N5984);
xor XOR2 (N6031, N6028, N3061);
and AND4 (N6032, N6016, N5980, N4903, N2308);
xor XOR2 (N6033, N6027, N1818);
buf BUF1 (N6034, N6023);
not NOT1 (N6035, N6032);
buf BUF1 (N6036, N6024);
not NOT1 (N6037, N6035);
nand NAND2 (N6038, N6033, N2236);
nand NAND4 (N6039, N6006, N817, N1590, N3569);
nand NAND3 (N6040, N6029, N2567, N3394);
buf BUF1 (N6041, N6031);
and AND3 (N6042, N6036, N3381, N1055);
nand NAND3 (N6043, N6034, N1847, N3546);
nor NOR4 (N6044, N6042, N4733, N5710, N706);
xor XOR2 (N6045, N6030, N4196);
not NOT1 (N6046, N6040);
buf BUF1 (N6047, N6046);
nor NOR4 (N6048, N6047, N4485, N5174, N17);
buf BUF1 (N6049, N6044);
nor NOR3 (N6050, N6049, N1902, N5223);
and AND4 (N6051, N6048, N3510, N5964, N3341);
nand NAND2 (N6052, N6050, N3801);
xor XOR2 (N6053, N6025, N2132);
or OR4 (N6054, N5997, N1782, N5298, N2256);
nor NOR3 (N6055, N6039, N5269, N4421);
xor XOR2 (N6056, N6053, N450);
not NOT1 (N6057, N6056);
not NOT1 (N6058, N6038);
xor XOR2 (N6059, N6045, N2343);
and AND4 (N6060, N6057, N2567, N3955, N5922);
not NOT1 (N6061, N6054);
not NOT1 (N6062, N6052);
nand NAND3 (N6063, N6037, N5579, N2029);
nand NAND3 (N6064, N6060, N46, N5157);
xor XOR2 (N6065, N6051, N1929);
nand NAND3 (N6066, N6063, N3351, N6062);
or OR4 (N6067, N3489, N3674, N1489, N858);
nand NAND4 (N6068, N6067, N5761, N3164, N4418);
and AND3 (N6069, N6041, N4310, N5764);
nor NOR4 (N6070, N6066, N23, N1918, N1452);
nand NAND3 (N6071, N6065, N4682, N2);
xor XOR2 (N6072, N6059, N5833);
or OR2 (N6073, N6072, N3975);
or OR2 (N6074, N6058, N368);
and AND4 (N6075, N6061, N3085, N340, N3966);
not NOT1 (N6076, N6043);
buf BUF1 (N6077, N6055);
or OR2 (N6078, N6070, N4340);
xor XOR2 (N6079, N6075, N2359);
and AND3 (N6080, N6074, N3906, N4949);
xor XOR2 (N6081, N6078, N2214);
nor NOR2 (N6082, N6073, N659);
not NOT1 (N6083, N6069);
nand NAND3 (N6084, N6076, N3433, N2251);
nand NAND4 (N6085, N6071, N2097, N2279, N6011);
or OR2 (N6086, N6077, N4209);
nor NOR2 (N6087, N6064, N3412);
or OR4 (N6088, N6079, N1734, N5441, N3592);
nand NAND3 (N6089, N6083, N2338, N790);
nor NOR2 (N6090, N6080, N5799);
xor XOR2 (N6091, N6086, N5848);
not NOT1 (N6092, N6082);
xor XOR2 (N6093, N6089, N281);
nand NAND2 (N6094, N6093, N5301);
or OR3 (N6095, N6094, N1243, N3440);
not NOT1 (N6096, N6085);
xor XOR2 (N6097, N6096, N3987);
xor XOR2 (N6098, N6095, N1300);
or OR2 (N6099, N6068, N4556);
and AND2 (N6100, N6090, N3404);
nand NAND2 (N6101, N6097, N3415);
or OR2 (N6102, N6081, N4515);
xor XOR2 (N6103, N6084, N4267);
not NOT1 (N6104, N6100);
or OR4 (N6105, N6091, N2100, N5833, N3585);
nand NAND2 (N6106, N6102, N3654);
or OR3 (N6107, N6101, N1897, N347);
and AND4 (N6108, N6104, N1701, N816, N455);
nor NOR2 (N6109, N6098, N5843);
and AND4 (N6110, N6103, N2463, N5539, N5250);
xor XOR2 (N6111, N6099, N2506);
not NOT1 (N6112, N6106);
xor XOR2 (N6113, N6112, N858);
or OR3 (N6114, N6108, N505, N3634);
not NOT1 (N6115, N6088);
not NOT1 (N6116, N6087);
xor XOR2 (N6117, N6109, N1359);
or OR3 (N6118, N6092, N1818, N2958);
or OR2 (N6119, N6117, N5207);
not NOT1 (N6120, N6118);
xor XOR2 (N6121, N6120, N2075);
not NOT1 (N6122, N6115);
buf BUF1 (N6123, N6113);
nor NOR3 (N6124, N6107, N3374, N2350);
not NOT1 (N6125, N6122);
or OR2 (N6126, N6121, N5760);
or OR2 (N6127, N6119, N1494);
nor NOR4 (N6128, N6127, N353, N6041, N2116);
and AND2 (N6129, N6116, N2158);
and AND3 (N6130, N6128, N1853, N567);
nor NOR2 (N6131, N6126, N1470);
nand NAND3 (N6132, N6105, N1783, N1052);
or OR4 (N6133, N6110, N1849, N1470, N3520);
nand NAND3 (N6134, N6130, N5659, N724);
nand NAND4 (N6135, N6134, N1495, N2362, N2712);
not NOT1 (N6136, N6129);
nor NOR3 (N6137, N6114, N2139, N3004);
or OR4 (N6138, N6133, N1691, N3680, N2197);
not NOT1 (N6139, N6136);
buf BUF1 (N6140, N6131);
not NOT1 (N6141, N6125);
buf BUF1 (N6142, N6123);
or OR2 (N6143, N6124, N5432);
not NOT1 (N6144, N6132);
or OR4 (N6145, N6141, N5845, N3274, N2419);
buf BUF1 (N6146, N6144);
nor NOR4 (N6147, N6145, N1694, N717, N4702);
not NOT1 (N6148, N6146);
or OR4 (N6149, N6111, N728, N5031, N4346);
buf BUF1 (N6150, N6143);
and AND2 (N6151, N6138, N4916);
nor NOR2 (N6152, N6137, N4994);
buf BUF1 (N6153, N6140);
nor NOR3 (N6154, N6150, N5295, N5966);
or OR2 (N6155, N6147, N1489);
buf BUF1 (N6156, N6155);
and AND3 (N6157, N6156, N1187, N2206);
xor XOR2 (N6158, N6152, N2338);
and AND4 (N6159, N6151, N568, N2734, N3240);
nand NAND4 (N6160, N6149, N4746, N2934, N4512);
nand NAND4 (N6161, N6159, N3892, N2962, N1846);
not NOT1 (N6162, N6148);
buf BUF1 (N6163, N6139);
not NOT1 (N6164, N6160);
nor NOR4 (N6165, N6163, N1068, N5816, N3783);
xor XOR2 (N6166, N6161, N3705);
and AND2 (N6167, N6164, N281);
nor NOR4 (N6168, N6135, N4100, N4324, N2951);
or OR3 (N6169, N6165, N1625, N6089);
xor XOR2 (N6170, N6154, N3447);
nand NAND3 (N6171, N6169, N577, N1557);
xor XOR2 (N6172, N6170, N4052);
and AND3 (N6173, N6162, N1071, N4169);
or OR3 (N6174, N6168, N1103, N5537);
xor XOR2 (N6175, N6171, N4373);
xor XOR2 (N6176, N6175, N4005);
and AND4 (N6177, N6157, N3551, N3859, N5026);
nand NAND4 (N6178, N6167, N1764, N2457, N809);
and AND2 (N6179, N6177, N4977);
not NOT1 (N6180, N6142);
nand NAND2 (N6181, N6166, N4157);
xor XOR2 (N6182, N6158, N4225);
not NOT1 (N6183, N6178);
not NOT1 (N6184, N6182);
or OR2 (N6185, N6181, N2028);
buf BUF1 (N6186, N6172);
nor NOR3 (N6187, N6183, N1882, N2130);
or OR4 (N6188, N6179, N2003, N4449, N3202);
and AND3 (N6189, N6173, N1891, N802);
not NOT1 (N6190, N6180);
nor NOR2 (N6191, N6188, N4564);
nand NAND4 (N6192, N6185, N5843, N3299, N5482);
or OR3 (N6193, N6192, N3891, N3242);
nor NOR3 (N6194, N6176, N4359, N1839);
xor XOR2 (N6195, N6191, N5750);
nand NAND3 (N6196, N6193, N6086, N1334);
or OR4 (N6197, N6196, N3276, N1392, N1709);
nand NAND4 (N6198, N6190, N3795, N4099, N53);
buf BUF1 (N6199, N6153);
or OR3 (N6200, N6194, N2083, N4813);
not NOT1 (N6201, N6200);
xor XOR2 (N6202, N6195, N2113);
and AND3 (N6203, N6198, N1260, N5087);
nor NOR3 (N6204, N6184, N5353, N3259);
and AND2 (N6205, N6199, N1511);
xor XOR2 (N6206, N6186, N542);
nand NAND4 (N6207, N6203, N6062, N832, N4702);
or OR2 (N6208, N6206, N3347);
nor NOR3 (N6209, N6187, N5223, N4489);
nor NOR3 (N6210, N6207, N3105, N6026);
and AND2 (N6211, N6204, N3835);
nand NAND3 (N6212, N6209, N2378, N3061);
not NOT1 (N6213, N6201);
nand NAND2 (N6214, N6205, N1120);
not NOT1 (N6215, N6214);
not NOT1 (N6216, N6202);
nand NAND3 (N6217, N6216, N5325, N753);
xor XOR2 (N6218, N6212, N5251);
nand NAND2 (N6219, N6218, N3491);
nor NOR4 (N6220, N6189, N5382, N3645, N5607);
xor XOR2 (N6221, N6220, N2852);
and AND4 (N6222, N6217, N3316, N4269, N1117);
nor NOR2 (N6223, N6221, N2600);
buf BUF1 (N6224, N6211);
not NOT1 (N6225, N6208);
buf BUF1 (N6226, N6210);
and AND4 (N6227, N6197, N5392, N3550, N1366);
buf BUF1 (N6228, N6223);
not NOT1 (N6229, N6174);
buf BUF1 (N6230, N6225);
buf BUF1 (N6231, N6215);
and AND2 (N6232, N6228, N1001);
or OR2 (N6233, N6213, N3014);
buf BUF1 (N6234, N6233);
nand NAND3 (N6235, N6219, N171, N1187);
or OR2 (N6236, N6229, N3216);
and AND2 (N6237, N6230, N5430);
buf BUF1 (N6238, N6236);
not NOT1 (N6239, N6226);
nand NAND2 (N6240, N6238, N2395);
buf BUF1 (N6241, N6224);
nand NAND3 (N6242, N6240, N1403, N4862);
not NOT1 (N6243, N6227);
and AND2 (N6244, N6235, N4191);
and AND2 (N6245, N6237, N5242);
not NOT1 (N6246, N6222);
nor NOR2 (N6247, N6241, N5401);
not NOT1 (N6248, N6242);
buf BUF1 (N6249, N6234);
nor NOR3 (N6250, N6248, N2523, N5030);
xor XOR2 (N6251, N6250, N1078);
buf BUF1 (N6252, N6251);
xor XOR2 (N6253, N6247, N2228);
not NOT1 (N6254, N6239);
nand NAND2 (N6255, N6252, N1523);
xor XOR2 (N6256, N6254, N1583);
or OR4 (N6257, N6246, N593, N5731, N1009);
and AND2 (N6258, N6256, N5701);
buf BUF1 (N6259, N6245);
and AND2 (N6260, N6253, N2491);
or OR2 (N6261, N6259, N769);
not NOT1 (N6262, N6243);
nand NAND3 (N6263, N6257, N1997, N3531);
and AND3 (N6264, N6244, N217, N5653);
or OR2 (N6265, N6231, N3480);
not NOT1 (N6266, N6255);
or OR3 (N6267, N6258, N5103, N169);
buf BUF1 (N6268, N6264);
xor XOR2 (N6269, N6263, N5401);
and AND2 (N6270, N6249, N5896);
not NOT1 (N6271, N6270);
or OR4 (N6272, N6262, N6049, N3530, N861);
or OR2 (N6273, N6268, N278);
and AND4 (N6274, N6232, N4129, N1662, N2249);
nand NAND4 (N6275, N6266, N1864, N5427, N3733);
or OR3 (N6276, N6260, N2055, N1536);
buf BUF1 (N6277, N6267);
or OR2 (N6278, N6274, N835);
and AND3 (N6279, N6265, N3182, N1952);
and AND4 (N6280, N6269, N1091, N855, N5243);
and AND4 (N6281, N6272, N4413, N4169, N6208);
and AND2 (N6282, N6281, N2577);
buf BUF1 (N6283, N6279);
nand NAND4 (N6284, N6273, N1347, N4191, N2506);
nor NOR2 (N6285, N6278, N3891);
or OR4 (N6286, N6283, N1683, N1391, N2427);
not NOT1 (N6287, N6275);
buf BUF1 (N6288, N6277);
xor XOR2 (N6289, N6280, N402);
buf BUF1 (N6290, N6287);
nand NAND3 (N6291, N6276, N1303, N128);
xor XOR2 (N6292, N6286, N136);
nand NAND4 (N6293, N6285, N2285, N4133, N3861);
nor NOR2 (N6294, N6284, N4116);
or OR4 (N6295, N6261, N5006, N2607, N171);
nor NOR2 (N6296, N6288, N5690);
not NOT1 (N6297, N6292);
xor XOR2 (N6298, N6297, N3144);
or OR2 (N6299, N6282, N3104);
or OR2 (N6300, N6298, N6201);
and AND4 (N6301, N6300, N2983, N5108, N999);
not NOT1 (N6302, N6301);
xor XOR2 (N6303, N6299, N3417);
nand NAND4 (N6304, N6295, N6099, N5715, N2699);
xor XOR2 (N6305, N6294, N1270);
buf BUF1 (N6306, N6304);
and AND2 (N6307, N6289, N1781);
not NOT1 (N6308, N6290);
and AND2 (N6309, N6271, N4016);
buf BUF1 (N6310, N6303);
nand NAND2 (N6311, N6309, N3643);
and AND4 (N6312, N6307, N4140, N535, N673);
and AND3 (N6313, N6311, N4097, N1888);
nand NAND3 (N6314, N6310, N202, N2089);
and AND3 (N6315, N6312, N5703, N1829);
nand NAND3 (N6316, N6313, N3776, N5319);
buf BUF1 (N6317, N6305);
not NOT1 (N6318, N6306);
not NOT1 (N6319, N6318);
buf BUF1 (N6320, N6317);
or OR2 (N6321, N6291, N6145);
nor NOR4 (N6322, N6308, N5071, N5800, N1373);
nand NAND4 (N6323, N6322, N2810, N81, N365);
xor XOR2 (N6324, N6321, N975);
nand NAND2 (N6325, N6323, N6147);
nand NAND2 (N6326, N6315, N367);
xor XOR2 (N6327, N6326, N2943);
and AND3 (N6328, N6327, N1621, N6044);
nand NAND4 (N6329, N6316, N1323, N2257, N1114);
nand NAND3 (N6330, N6329, N1459, N2219);
nand NAND3 (N6331, N6330, N1700, N2000);
and AND2 (N6332, N6319, N3316);
or OR2 (N6333, N6320, N232);
nand NAND4 (N6334, N6293, N4517, N3261, N597);
xor XOR2 (N6335, N6302, N866);
xor XOR2 (N6336, N6328, N4852);
nor NOR3 (N6337, N6333, N4425, N5037);
not NOT1 (N6338, N6324);
nor NOR2 (N6339, N6334, N2760);
buf BUF1 (N6340, N6331);
and AND2 (N6341, N6337, N1398);
xor XOR2 (N6342, N6325, N1473);
nand NAND4 (N6343, N6340, N2612, N5794, N4929);
and AND2 (N6344, N6342, N4276);
not NOT1 (N6345, N6314);
and AND4 (N6346, N6332, N3717, N4317, N5118);
and AND3 (N6347, N6335, N6235, N980);
nor NOR3 (N6348, N6341, N3798, N4613);
not NOT1 (N6349, N6296);
nor NOR3 (N6350, N6346, N1699, N2119);
nand NAND4 (N6351, N6345, N4202, N3623, N3099);
xor XOR2 (N6352, N6338, N5355);
nor NOR3 (N6353, N6352, N1654, N6343);
nand NAND4 (N6354, N2403, N5115, N6232, N1436);
and AND3 (N6355, N6339, N3306, N4857);
nand NAND3 (N6356, N6350, N2636, N6029);
not NOT1 (N6357, N6354);
or OR2 (N6358, N6347, N5771);
nand NAND4 (N6359, N6358, N6160, N5575, N4520);
not NOT1 (N6360, N6355);
nor NOR2 (N6361, N6360, N5052);
nor NOR3 (N6362, N6348, N427, N3184);
xor XOR2 (N6363, N6362, N2777);
xor XOR2 (N6364, N6359, N2899);
xor XOR2 (N6365, N6356, N1783);
nor NOR3 (N6366, N6353, N3928, N4286);
or OR3 (N6367, N6336, N1315, N639);
xor XOR2 (N6368, N6357, N617);
not NOT1 (N6369, N6361);
nand NAND4 (N6370, N6363, N2418, N5139, N4321);
not NOT1 (N6371, N6366);
nand NAND4 (N6372, N6368, N2423, N4746, N5751);
xor XOR2 (N6373, N6351, N5129);
and AND4 (N6374, N6372, N5762, N6049, N2429);
nand NAND3 (N6375, N6371, N3770, N4121);
and AND2 (N6376, N6365, N2618);
nor NOR4 (N6377, N6374, N457, N2150, N661);
xor XOR2 (N6378, N6370, N4546);
or OR4 (N6379, N6369, N557, N2279, N1819);
xor XOR2 (N6380, N6379, N476);
not NOT1 (N6381, N6378);
or OR4 (N6382, N6376, N1502, N2001, N2729);
nor NOR4 (N6383, N6375, N5140, N1780, N549);
buf BUF1 (N6384, N6377);
not NOT1 (N6385, N6380);
not NOT1 (N6386, N6344);
nor NOR3 (N6387, N6349, N1912, N1764);
buf BUF1 (N6388, N6382);
not NOT1 (N6389, N6367);
nor NOR4 (N6390, N6388, N4624, N3249, N5071);
xor XOR2 (N6391, N6386, N5454);
or OR2 (N6392, N6373, N3054);
nand NAND2 (N6393, N6383, N5111);
and AND4 (N6394, N6385, N1812, N3088, N4959);
xor XOR2 (N6395, N6384, N3893);
not NOT1 (N6396, N6364);
or OR2 (N6397, N6387, N5980);
or OR3 (N6398, N6390, N5426, N4156);
nand NAND3 (N6399, N6397, N3553, N2242);
nor NOR3 (N6400, N6399, N6063, N918);
xor XOR2 (N6401, N6398, N3120);
and AND2 (N6402, N6389, N2555);
nand NAND3 (N6403, N6393, N4481, N3667);
xor XOR2 (N6404, N6395, N2301);
or OR2 (N6405, N6400, N2213);
xor XOR2 (N6406, N6381, N808);
buf BUF1 (N6407, N6392);
or OR2 (N6408, N6405, N1952);
nand NAND2 (N6409, N6396, N4292);
nor NOR4 (N6410, N6403, N5176, N770, N3338);
nand NAND2 (N6411, N6402, N4022);
or OR4 (N6412, N6391, N4058, N1900, N5255);
xor XOR2 (N6413, N6412, N2599);
and AND4 (N6414, N6410, N5922, N1262, N2610);
and AND3 (N6415, N6404, N5850, N343);
or OR3 (N6416, N6409, N3125, N4723);
and AND4 (N6417, N6411, N4452, N5810, N1032);
nand NAND4 (N6418, N6401, N2859, N841, N5568);
nor NOR4 (N6419, N6415, N4264, N1360, N897);
and AND3 (N6420, N6406, N1151, N927);
buf BUF1 (N6421, N6420);
nand NAND2 (N6422, N6408, N4963);
nor NOR4 (N6423, N6414, N1443, N448, N4153);
xor XOR2 (N6424, N6417, N5422);
buf BUF1 (N6425, N6418);
nor NOR2 (N6426, N6421, N3164);
nand NAND3 (N6427, N6416, N6251, N5519);
not NOT1 (N6428, N6394);
and AND4 (N6429, N6422, N5295, N168, N4863);
and AND4 (N6430, N6423, N3121, N2512, N2046);
xor XOR2 (N6431, N6419, N3623);
and AND2 (N6432, N6430, N4111);
xor XOR2 (N6433, N6413, N1080);
buf BUF1 (N6434, N6426);
and AND4 (N6435, N6407, N2765, N2254, N3033);
not NOT1 (N6436, N6427);
nand NAND4 (N6437, N6424, N6411, N1532, N1070);
not NOT1 (N6438, N6435);
buf BUF1 (N6439, N6437);
nor NOR3 (N6440, N6433, N2646, N1571);
nor NOR3 (N6441, N6436, N2319, N4368);
not NOT1 (N6442, N6439);
or OR3 (N6443, N6440, N4517, N3315);
nor NOR4 (N6444, N6443, N1926, N1817, N4063);
and AND2 (N6445, N6428, N2794);
or OR4 (N6446, N6432, N1220, N870, N6061);
and AND3 (N6447, N6434, N3724, N141);
xor XOR2 (N6448, N6447, N4978);
or OR2 (N6449, N6445, N4499);
nand NAND4 (N6450, N6425, N2595, N3337, N4818);
or OR3 (N6451, N6431, N6158, N3161);
or OR4 (N6452, N6446, N4488, N3230, N5532);
and AND4 (N6453, N6438, N1070, N762, N5196);
and AND3 (N6454, N6452, N5829, N2011);
not NOT1 (N6455, N6444);
or OR4 (N6456, N6442, N4491, N5877, N1494);
buf BUF1 (N6457, N6429);
and AND2 (N6458, N6453, N3248);
nor NOR2 (N6459, N6457, N3626);
buf BUF1 (N6460, N6454);
not NOT1 (N6461, N6441);
buf BUF1 (N6462, N6459);
buf BUF1 (N6463, N6449);
nor NOR2 (N6464, N6455, N88);
nand NAND3 (N6465, N6460, N6221, N3542);
or OR2 (N6466, N6458, N653);
nor NOR2 (N6467, N6456, N6335);
and AND4 (N6468, N6466, N3559, N2092, N5166);
not NOT1 (N6469, N6465);
xor XOR2 (N6470, N6461, N1787);
nand NAND3 (N6471, N6467, N6411, N2561);
nor NOR3 (N6472, N6451, N3611, N6120);
xor XOR2 (N6473, N6469, N4733);
xor XOR2 (N6474, N6472, N3974);
and AND2 (N6475, N6468, N2526);
nand NAND2 (N6476, N6462, N5818);
not NOT1 (N6477, N6463);
or OR3 (N6478, N6477, N2554, N3274);
and AND3 (N6479, N6474, N3162, N4566);
buf BUF1 (N6480, N6475);
or OR3 (N6481, N6478, N1619, N3424);
nand NAND4 (N6482, N6480, N4699, N380, N5881);
or OR4 (N6483, N6481, N3208, N4968, N43);
or OR4 (N6484, N6450, N3614, N2614, N4487);
and AND2 (N6485, N6470, N861);
nand NAND4 (N6486, N6471, N4974, N426, N326);
and AND3 (N6487, N6476, N5970, N2510);
nor NOR4 (N6488, N6464, N627, N4308, N2587);
or OR4 (N6489, N6486, N2476, N4292, N1568);
nand NAND3 (N6490, N6487, N2121, N5672);
and AND2 (N6491, N6448, N4970);
nand NAND2 (N6492, N6490, N3504);
and AND2 (N6493, N6484, N6144);
and AND3 (N6494, N6473, N3330, N3196);
buf BUF1 (N6495, N6483);
or OR2 (N6496, N6488, N4789);
and AND2 (N6497, N6489, N6353);
nor NOR4 (N6498, N6479, N1985, N2332, N6391);
nand NAND4 (N6499, N6495, N1035, N2654, N1783);
nor NOR2 (N6500, N6497, N1373);
nor NOR3 (N6501, N6485, N3764, N6050);
nand NAND2 (N6502, N6499, N2647);
or OR3 (N6503, N6482, N4409, N2171);
xor XOR2 (N6504, N6494, N1350);
xor XOR2 (N6505, N6492, N2601);
or OR3 (N6506, N6504, N1101, N2701);
and AND2 (N6507, N6505, N3604);
buf BUF1 (N6508, N6496);
and AND2 (N6509, N6503, N5425);
and AND2 (N6510, N6506, N3952);
buf BUF1 (N6511, N6500);
not NOT1 (N6512, N6491);
or OR2 (N6513, N6508, N3109);
nor NOR4 (N6514, N6493, N5715, N284, N1214);
buf BUF1 (N6515, N6502);
and AND3 (N6516, N6509, N3069, N1365);
and AND2 (N6517, N6516, N883);
nand NAND3 (N6518, N6511, N6362, N4226);
buf BUF1 (N6519, N6501);
nor NOR3 (N6520, N6510, N1403, N530);
and AND3 (N6521, N6519, N6382, N3763);
nand NAND3 (N6522, N6515, N583, N2538);
and AND2 (N6523, N6513, N2437);
nand NAND2 (N6524, N6522, N356);
not NOT1 (N6525, N6517);
or OR2 (N6526, N6512, N4590);
not NOT1 (N6527, N6498);
xor XOR2 (N6528, N6514, N6220);
or OR2 (N6529, N6527, N4770);
or OR2 (N6530, N6507, N5113);
nand NAND4 (N6531, N6528, N5204, N552, N6012);
nor NOR4 (N6532, N6526, N5583, N3338, N3261);
not NOT1 (N6533, N6530);
and AND4 (N6534, N6533, N6149, N4354, N4506);
nor NOR3 (N6535, N6525, N2579, N2286);
xor XOR2 (N6536, N6529, N4623);
not NOT1 (N6537, N6521);
and AND4 (N6538, N6532, N4412, N4816, N2890);
xor XOR2 (N6539, N6537, N3841);
xor XOR2 (N6540, N6535, N3229);
nand NAND2 (N6541, N6538, N5377);
nand NAND3 (N6542, N6531, N4081, N6533);
and AND2 (N6543, N6524, N284);
xor XOR2 (N6544, N6536, N2366);
xor XOR2 (N6545, N6544, N6456);
not NOT1 (N6546, N6523);
buf BUF1 (N6547, N6539);
buf BUF1 (N6548, N6545);
buf BUF1 (N6549, N6518);
nor NOR3 (N6550, N6541, N4773, N6154);
buf BUF1 (N6551, N6549);
and AND2 (N6552, N6520, N5794);
nor NOR4 (N6553, N6551, N3723, N1161, N3609);
xor XOR2 (N6554, N6553, N1037);
not NOT1 (N6555, N6542);
not NOT1 (N6556, N6540);
nor NOR3 (N6557, N6556, N123, N5023);
nor NOR2 (N6558, N6546, N4053);
nand NAND3 (N6559, N6552, N5585, N2474);
or OR3 (N6560, N6543, N5804, N846);
and AND2 (N6561, N6550, N1120);
not NOT1 (N6562, N6560);
buf BUF1 (N6563, N6561);
not NOT1 (N6564, N6555);
nand NAND3 (N6565, N6562, N1468, N1518);
and AND2 (N6566, N6548, N3722);
buf BUF1 (N6567, N6566);
xor XOR2 (N6568, N6564, N4394);
not NOT1 (N6569, N6568);
or OR2 (N6570, N6547, N1736);
or OR2 (N6571, N6558, N1046);
not NOT1 (N6572, N6557);
nor NOR3 (N6573, N6563, N6483, N3111);
and AND2 (N6574, N6567, N2842);
xor XOR2 (N6575, N6565, N1073);
xor XOR2 (N6576, N6572, N814);
nand NAND2 (N6577, N6570, N3166);
buf BUF1 (N6578, N6559);
buf BUF1 (N6579, N6554);
nor NOR4 (N6580, N6575, N3028, N1639, N4686);
nor NOR4 (N6581, N6573, N11, N1430, N5919);
nor NOR4 (N6582, N6577, N1222, N773, N6386);
nor NOR4 (N6583, N6574, N3230, N5173, N5947);
xor XOR2 (N6584, N6571, N5822);
or OR3 (N6585, N6578, N6098, N5424);
or OR2 (N6586, N6576, N6536);
not NOT1 (N6587, N6584);
buf BUF1 (N6588, N6587);
or OR3 (N6589, N6569, N9, N4603);
xor XOR2 (N6590, N6579, N4128);
nor NOR4 (N6591, N6583, N2271, N1617, N5693);
xor XOR2 (N6592, N6588, N160);
nor NOR4 (N6593, N6581, N2493, N4494, N5615);
nor NOR2 (N6594, N6534, N6034);
and AND2 (N6595, N6591, N5988);
buf BUF1 (N6596, N6595);
xor XOR2 (N6597, N6585, N480);
not NOT1 (N6598, N6596);
buf BUF1 (N6599, N6580);
nand NAND3 (N6600, N6582, N224, N866);
or OR2 (N6601, N6597, N859);
nor NOR3 (N6602, N6598, N2455, N5498);
nor NOR4 (N6603, N6593, N1763, N5164, N3475);
and AND2 (N6604, N6589, N1091);
nand NAND4 (N6605, N6594, N1950, N3278, N1993);
nand NAND2 (N6606, N6586, N5957);
nand NAND2 (N6607, N6604, N5672);
nor NOR4 (N6608, N6603, N871, N4609, N5604);
not NOT1 (N6609, N6601);
buf BUF1 (N6610, N6599);
and AND2 (N6611, N6607, N5143);
not NOT1 (N6612, N6605);
nand NAND4 (N6613, N6608, N4503, N5866, N23);
and AND2 (N6614, N6610, N297);
not NOT1 (N6615, N6602);
buf BUF1 (N6616, N6592);
buf BUF1 (N6617, N6606);
buf BUF1 (N6618, N6616);
not NOT1 (N6619, N6615);
nand NAND3 (N6620, N6590, N4868, N6076);
buf BUF1 (N6621, N6619);
not NOT1 (N6622, N6612);
buf BUF1 (N6623, N6617);
and AND3 (N6624, N6620, N4514, N3144);
nor NOR4 (N6625, N6624, N330, N4630, N2491);
nor NOR3 (N6626, N6622, N6623, N3141);
not NOT1 (N6627, N242);
nor NOR3 (N6628, N6618, N333, N5540);
and AND2 (N6629, N6609, N1735);
xor XOR2 (N6630, N6627, N4551);
not NOT1 (N6631, N6629);
buf BUF1 (N6632, N6625);
xor XOR2 (N6633, N6614, N855);
not NOT1 (N6634, N6631);
and AND2 (N6635, N6632, N2818);
nor NOR2 (N6636, N6621, N2540);
buf BUF1 (N6637, N6611);
xor XOR2 (N6638, N6613, N407);
and AND4 (N6639, N6633, N3591, N2838, N1335);
and AND4 (N6640, N6634, N3109, N724, N646);
not NOT1 (N6641, N6628);
xor XOR2 (N6642, N6639, N1388);
not NOT1 (N6643, N6642);
buf BUF1 (N6644, N6635);
and AND3 (N6645, N6630, N819, N5419);
nor NOR4 (N6646, N6626, N1534, N3633, N1477);
nor NOR2 (N6647, N6646, N6257);
nor NOR2 (N6648, N6647, N4406);
and AND4 (N6649, N6637, N3636, N4136, N4522);
and AND2 (N6650, N6600, N6014);
nor NOR2 (N6651, N6650, N5992);
buf BUF1 (N6652, N6649);
xor XOR2 (N6653, N6644, N3170);
xor XOR2 (N6654, N6648, N3214);
not NOT1 (N6655, N6638);
xor XOR2 (N6656, N6643, N4878);
or OR2 (N6657, N6636, N1779);
nand NAND2 (N6658, N6655, N588);
nand NAND4 (N6659, N6653, N86, N4263, N6219);
and AND3 (N6660, N6645, N5553, N2947);
nor NOR2 (N6661, N6660, N4468);
nor NOR4 (N6662, N6640, N1561, N1315, N4685);
nand NAND2 (N6663, N6658, N4486);
buf BUF1 (N6664, N6654);
and AND4 (N6665, N6652, N2832, N2617, N172);
nor NOR2 (N6666, N6651, N4516);
xor XOR2 (N6667, N6659, N2709);
buf BUF1 (N6668, N6661);
xor XOR2 (N6669, N6665, N251);
not NOT1 (N6670, N6657);
or OR4 (N6671, N6662, N2835, N4836, N3840);
or OR3 (N6672, N6667, N345, N3976);
not NOT1 (N6673, N6672);
and AND4 (N6674, N6669, N5057, N2048, N968);
buf BUF1 (N6675, N6674);
xor XOR2 (N6676, N6673, N702);
buf BUF1 (N6677, N6663);
xor XOR2 (N6678, N6675, N2809);
and AND4 (N6679, N6641, N2434, N3534, N5066);
not NOT1 (N6680, N6666);
buf BUF1 (N6681, N6680);
xor XOR2 (N6682, N6681, N1620);
and AND3 (N6683, N6677, N572, N6155);
not NOT1 (N6684, N6671);
or OR4 (N6685, N6664, N664, N975, N1826);
nor NOR2 (N6686, N6670, N3712);
buf BUF1 (N6687, N6682);
xor XOR2 (N6688, N6684, N4871);
or OR2 (N6689, N6679, N942);
nand NAND3 (N6690, N6683, N1025, N910);
not NOT1 (N6691, N6690);
nand NAND2 (N6692, N6688, N634);
nor NOR3 (N6693, N6692, N3969, N6081);
or OR2 (N6694, N6685, N6394);
buf BUF1 (N6695, N6694);
not NOT1 (N6696, N6676);
nand NAND2 (N6697, N6696, N745);
not NOT1 (N6698, N6689);
not NOT1 (N6699, N6668);
xor XOR2 (N6700, N6699, N6525);
nor NOR2 (N6701, N6700, N2126);
or OR4 (N6702, N6697, N4175, N244, N2069);
and AND2 (N6703, N6701, N2797);
or OR3 (N6704, N6691, N99, N1845);
nand NAND2 (N6705, N6656, N4440);
or OR4 (N6706, N6703, N1533, N818, N4055);
not NOT1 (N6707, N6686);
nor NOR3 (N6708, N6705, N2407, N1657);
nor NOR2 (N6709, N6698, N1134);
and AND4 (N6710, N6695, N1423, N709, N5760);
and AND3 (N6711, N6706, N1555, N4585);
xor XOR2 (N6712, N6704, N5623);
not NOT1 (N6713, N6693);
nor NOR4 (N6714, N6678, N3981, N3746, N5111);
xor XOR2 (N6715, N6713, N1919);
xor XOR2 (N6716, N6709, N4653);
nand NAND2 (N6717, N6716, N281);
xor XOR2 (N6718, N6687, N2536);
nand NAND4 (N6719, N6711, N325, N1956, N2878);
buf BUF1 (N6720, N6715);
nor NOR2 (N6721, N6720, N3110);
buf BUF1 (N6722, N6707);
and AND2 (N6723, N6722, N2349);
xor XOR2 (N6724, N6719, N1954);
xor XOR2 (N6725, N6721, N4212);
or OR2 (N6726, N6714, N2301);
xor XOR2 (N6727, N6708, N1102);
xor XOR2 (N6728, N6718, N5765);
not NOT1 (N6729, N6723);
buf BUF1 (N6730, N6726);
and AND4 (N6731, N6729, N4418, N1198, N2703);
xor XOR2 (N6732, N6728, N6515);
not NOT1 (N6733, N6712);
nor NOR4 (N6734, N6727, N4500, N2572, N3158);
not NOT1 (N6735, N6710);
nor NOR3 (N6736, N6734, N6468, N1229);
or OR3 (N6737, N6717, N2770, N2333);
buf BUF1 (N6738, N6724);
buf BUF1 (N6739, N6735);
and AND2 (N6740, N6702, N4333);
not NOT1 (N6741, N6737);
nor NOR4 (N6742, N6733, N4755, N517, N1693);
or OR4 (N6743, N6739, N3192, N3877, N816);
nor NOR3 (N6744, N6736, N5233, N5585);
buf BUF1 (N6745, N6725);
and AND2 (N6746, N6740, N1074);
xor XOR2 (N6747, N6745, N4597);
xor XOR2 (N6748, N6741, N5517);
and AND4 (N6749, N6743, N3303, N273, N2125);
not NOT1 (N6750, N6732);
nand NAND4 (N6751, N6742, N3118, N3542, N1501);
and AND2 (N6752, N6751, N6749);
xor XOR2 (N6753, N3510, N4367);
and AND2 (N6754, N6750, N839);
not NOT1 (N6755, N6730);
not NOT1 (N6756, N6754);
or OR2 (N6757, N6747, N5732);
nor NOR3 (N6758, N6744, N4974, N5826);
xor XOR2 (N6759, N6731, N437);
xor XOR2 (N6760, N6753, N6590);
and AND4 (N6761, N6755, N4052, N1250, N5539);
xor XOR2 (N6762, N6746, N2431);
xor XOR2 (N6763, N6752, N5050);
and AND3 (N6764, N6763, N4855, N1674);
buf BUF1 (N6765, N6756);
buf BUF1 (N6766, N6757);
xor XOR2 (N6767, N6758, N3096);
not NOT1 (N6768, N6748);
not NOT1 (N6769, N6768);
xor XOR2 (N6770, N6761, N5593);
buf BUF1 (N6771, N6770);
or OR4 (N6772, N6767, N3018, N2954, N4793);
buf BUF1 (N6773, N6772);
and AND3 (N6774, N6762, N3385, N1537);
not NOT1 (N6775, N6760);
not NOT1 (N6776, N6759);
nand NAND2 (N6777, N6765, N391);
buf BUF1 (N6778, N6773);
nand NAND3 (N6779, N6771, N3140, N1101);
not NOT1 (N6780, N6777);
nand NAND4 (N6781, N6738, N322, N3184, N1903);
buf BUF1 (N6782, N6781);
or OR3 (N6783, N6769, N2483, N4179);
nand NAND3 (N6784, N6779, N185, N1262);
not NOT1 (N6785, N6774);
nand NAND2 (N6786, N6764, N1798);
or OR2 (N6787, N6778, N6339);
nand NAND3 (N6788, N6775, N3671, N1952);
or OR4 (N6789, N6788, N5472, N5943, N2640);
nand NAND3 (N6790, N6784, N6736, N5255);
not NOT1 (N6791, N6776);
or OR3 (N6792, N6780, N4702, N4566);
nor NOR4 (N6793, N6787, N1717, N1839, N3241);
and AND4 (N6794, N6786, N2569, N148, N4881);
and AND4 (N6795, N6792, N3631, N3461, N1448);
xor XOR2 (N6796, N6795, N1260);
nand NAND3 (N6797, N6785, N1943, N2559);
xor XOR2 (N6798, N6791, N95);
and AND2 (N6799, N6796, N39);
buf BUF1 (N6800, N6794);
and AND4 (N6801, N6782, N1517, N1625, N6641);
nand NAND4 (N6802, N6799, N2818, N6692, N3591);
xor XOR2 (N6803, N6766, N3244);
and AND3 (N6804, N6783, N3979, N6692);
nor NOR4 (N6805, N6802, N2070, N4420, N6668);
nand NAND2 (N6806, N6805, N4791);
not NOT1 (N6807, N6800);
and AND4 (N6808, N6798, N5508, N6242, N6311);
or OR2 (N6809, N6804, N879);
or OR3 (N6810, N6793, N1398, N5248);
not NOT1 (N6811, N6808);
or OR4 (N6812, N6790, N1060, N5470, N3576);
xor XOR2 (N6813, N6811, N1141);
nor NOR3 (N6814, N6807, N2269, N2380);
nand NAND2 (N6815, N6810, N3597);
xor XOR2 (N6816, N6803, N4691);
or OR2 (N6817, N6797, N3566);
xor XOR2 (N6818, N6814, N4219);
nor NOR2 (N6819, N6816, N622);
xor XOR2 (N6820, N6812, N1306);
or OR4 (N6821, N6817, N4153, N986, N3836);
buf BUF1 (N6822, N6806);
or OR2 (N6823, N6820, N1112);
nand NAND4 (N6824, N6815, N1046, N1940, N6103);
or OR2 (N6825, N6821, N4854);
nand NAND2 (N6826, N6824, N4252);
xor XOR2 (N6827, N6823, N3409);
nor NOR2 (N6828, N6822, N4980);
buf BUF1 (N6829, N6826);
not NOT1 (N6830, N6819);
buf BUF1 (N6831, N6789);
nand NAND3 (N6832, N6827, N4219, N390);
not NOT1 (N6833, N6829);
or OR2 (N6834, N6831, N739);
nor NOR4 (N6835, N6813, N1138, N2733, N946);
nand NAND3 (N6836, N6832, N3384, N2069);
xor XOR2 (N6837, N6830, N2771);
xor XOR2 (N6838, N6825, N6790);
nand NAND2 (N6839, N6809, N1856);
or OR3 (N6840, N6836, N569, N2516);
nor NOR3 (N6841, N6835, N6808, N1372);
buf BUF1 (N6842, N6801);
nand NAND3 (N6843, N6841, N2300, N4938);
nand NAND3 (N6844, N6833, N4765, N4909);
or OR2 (N6845, N6844, N5619);
not NOT1 (N6846, N6842);
nand NAND4 (N6847, N6845, N661, N1320, N723);
nor NOR4 (N6848, N6839, N3375, N1556, N5880);
nor NOR2 (N6849, N6847, N331);
buf BUF1 (N6850, N6828);
nand NAND3 (N6851, N6818, N4552, N6615);
not NOT1 (N6852, N6837);
xor XOR2 (N6853, N6851, N3765);
not NOT1 (N6854, N6850);
nand NAND3 (N6855, N6854, N683, N5313);
nor NOR2 (N6856, N6849, N1150);
xor XOR2 (N6857, N6856, N4619);
buf BUF1 (N6858, N6857);
and AND2 (N6859, N6840, N6355);
or OR2 (N6860, N6852, N5774);
buf BUF1 (N6861, N6843);
buf BUF1 (N6862, N6838);
nor NOR3 (N6863, N6859, N850, N118);
nor NOR4 (N6864, N6848, N598, N740, N6046);
xor XOR2 (N6865, N6855, N3017);
and AND4 (N6866, N6858, N805, N2279, N6545);
and AND3 (N6867, N6853, N2583, N1569);
or OR3 (N6868, N6867, N3154, N6666);
xor XOR2 (N6869, N6865, N6802);
buf BUF1 (N6870, N6866);
buf BUF1 (N6871, N6870);
and AND4 (N6872, N6871, N848, N3303, N5198);
nand NAND2 (N6873, N6834, N3160);
nor NOR3 (N6874, N6860, N5763, N2898);
and AND3 (N6875, N6869, N2620, N748);
nand NAND2 (N6876, N6875, N2704);
xor XOR2 (N6877, N6876, N4378);
or OR2 (N6878, N6864, N6067);
buf BUF1 (N6879, N6861);
and AND3 (N6880, N6877, N1759, N333);
not NOT1 (N6881, N6846);
nor NOR3 (N6882, N6874, N337, N3751);
buf BUF1 (N6883, N6879);
nand NAND4 (N6884, N6872, N1945, N1544, N582);
and AND2 (N6885, N6873, N3538);
or OR4 (N6886, N6884, N5952, N2839, N4399);
buf BUF1 (N6887, N6886);
nand NAND3 (N6888, N6880, N6587, N615);
and AND2 (N6889, N6881, N2247);
buf BUF1 (N6890, N6885);
or OR2 (N6891, N6888, N5385);
not NOT1 (N6892, N6890);
buf BUF1 (N6893, N6882);
buf BUF1 (N6894, N6883);
buf BUF1 (N6895, N6889);
and AND2 (N6896, N6878, N1282);
not NOT1 (N6897, N6863);
nor NOR4 (N6898, N6896, N3907, N392, N3400);
and AND2 (N6899, N6895, N5367);
buf BUF1 (N6900, N6897);
nand NAND4 (N6901, N6887, N4394, N4137, N1818);
not NOT1 (N6902, N6894);
buf BUF1 (N6903, N6868);
buf BUF1 (N6904, N6901);
xor XOR2 (N6905, N6898, N4430);
xor XOR2 (N6906, N6891, N1240);
or OR3 (N6907, N6904, N2014, N6821);
not NOT1 (N6908, N6907);
or OR3 (N6909, N6899, N3502, N1530);
not NOT1 (N6910, N6862);
buf BUF1 (N6911, N6909);
buf BUF1 (N6912, N6893);
and AND2 (N6913, N6892, N200);
buf BUF1 (N6914, N6913);
nor NOR2 (N6915, N6900, N4505);
xor XOR2 (N6916, N6910, N6420);
or OR2 (N6917, N6908, N3407);
nor NOR2 (N6918, N6903, N2914);
nor NOR4 (N6919, N6912, N2946, N595, N3116);
xor XOR2 (N6920, N6902, N6407);
nor NOR2 (N6921, N6916, N4390);
not NOT1 (N6922, N6919);
not NOT1 (N6923, N6920);
not NOT1 (N6924, N6921);
and AND4 (N6925, N6924, N4587, N6314, N6516);
xor XOR2 (N6926, N6905, N615);
nand NAND4 (N6927, N6911, N1996, N941, N6711);
not NOT1 (N6928, N6918);
or OR4 (N6929, N6927, N3505, N3061, N1149);
and AND4 (N6930, N6915, N2844, N761, N3907);
and AND3 (N6931, N6914, N172, N777);
nor NOR4 (N6932, N6906, N3444, N5038, N3325);
or OR3 (N6933, N6926, N2982, N667);
nor NOR2 (N6934, N6917, N3011);
not NOT1 (N6935, N6930);
and AND4 (N6936, N6928, N986, N3155, N5575);
buf BUF1 (N6937, N6932);
or OR3 (N6938, N6925, N6055, N2799);
nand NAND3 (N6939, N6934, N5554, N4968);
buf BUF1 (N6940, N6937);
buf BUF1 (N6941, N6933);
buf BUF1 (N6942, N6939);
buf BUF1 (N6943, N6935);
not NOT1 (N6944, N6942);
nor NOR4 (N6945, N6943, N808, N1844, N4011);
buf BUF1 (N6946, N6945);
xor XOR2 (N6947, N6938, N1127);
not NOT1 (N6948, N6946);
not NOT1 (N6949, N6941);
not NOT1 (N6950, N6947);
or OR2 (N6951, N6948, N2958);
nor NOR4 (N6952, N6949, N4546, N3626, N2089);
or OR2 (N6953, N6951, N2381);
nand NAND2 (N6954, N6929, N5926);
or OR2 (N6955, N6954, N1417);
xor XOR2 (N6956, N6923, N4846);
and AND3 (N6957, N6931, N5028, N6387);
not NOT1 (N6958, N6922);
not NOT1 (N6959, N6955);
or OR2 (N6960, N6950, N6051);
buf BUF1 (N6961, N6936);
buf BUF1 (N6962, N6940);
nand NAND4 (N6963, N6952, N2250, N5308, N684);
nor NOR2 (N6964, N6956, N5342);
nor NOR4 (N6965, N6953, N6937, N3115, N2593);
nor NOR2 (N6966, N6965, N281);
or OR2 (N6967, N6964, N889);
or OR4 (N6968, N6960, N6491, N3411, N2348);
and AND4 (N6969, N6967, N5278, N6689, N5183);
buf BUF1 (N6970, N6944);
and AND2 (N6971, N6969, N1061);
not NOT1 (N6972, N6962);
buf BUF1 (N6973, N6971);
not NOT1 (N6974, N6961);
or OR4 (N6975, N6970, N4271, N5402, N1878);
xor XOR2 (N6976, N6959, N709);
nand NAND2 (N6977, N6974, N3547);
and AND2 (N6978, N6958, N97);
buf BUF1 (N6979, N6963);
not NOT1 (N6980, N6977);
xor XOR2 (N6981, N6966, N5163);
nor NOR4 (N6982, N6978, N5286, N6664, N6750);
nand NAND3 (N6983, N6980, N5792, N3598);
nand NAND4 (N6984, N6957, N2944, N3518, N6488);
nand NAND3 (N6985, N6981, N5721, N2572);
nand NAND3 (N6986, N6972, N4970, N4818);
nor NOR4 (N6987, N6979, N3268, N1394, N2854);
or OR4 (N6988, N6985, N330, N4778, N5083);
not NOT1 (N6989, N6987);
buf BUF1 (N6990, N6988);
nand NAND3 (N6991, N6984, N340, N5558);
or OR4 (N6992, N6983, N6678, N1664, N6872);
nor NOR4 (N6993, N6976, N661, N3696, N1678);
or OR3 (N6994, N6990, N3673, N5561);
nor NOR3 (N6995, N6986, N2461, N3583);
xor XOR2 (N6996, N6975, N4394);
or OR3 (N6997, N6994, N5671, N3339);
buf BUF1 (N6998, N6991);
or OR4 (N6999, N6992, N6174, N2304, N6515);
not NOT1 (N7000, N6998);
and AND2 (N7001, N6996, N4997);
nand NAND4 (N7002, N6989, N4926, N2709, N3009);
buf BUF1 (N7003, N6997);
nor NOR4 (N7004, N6973, N2987, N2779, N3883);
buf BUF1 (N7005, N7001);
nor NOR3 (N7006, N6993, N1918, N284);
nor NOR4 (N7007, N6982, N5112, N5862, N2294);
nand NAND4 (N7008, N6999, N2826, N5518, N670);
nand NAND2 (N7009, N6968, N2390);
nor NOR2 (N7010, N7003, N4002);
xor XOR2 (N7011, N7002, N1117);
nand NAND4 (N7012, N7009, N3288, N4844, N4906);
and AND3 (N7013, N6995, N676, N2061);
nor NOR4 (N7014, N7005, N3300, N5189, N4975);
not NOT1 (N7015, N7000);
not NOT1 (N7016, N7015);
not NOT1 (N7017, N7006);
xor XOR2 (N7018, N7010, N1814);
nand NAND4 (N7019, N7016, N3085, N2747, N3099);
and AND4 (N7020, N7007, N2655, N6911, N3269);
buf BUF1 (N7021, N7011);
not NOT1 (N7022, N7020);
not NOT1 (N7023, N7008);
xor XOR2 (N7024, N7023, N5438);
xor XOR2 (N7025, N7012, N5240);
not NOT1 (N7026, N7024);
not NOT1 (N7027, N7022);
nor NOR3 (N7028, N7019, N6269, N5972);
buf BUF1 (N7029, N7004);
or OR2 (N7030, N7018, N2597);
and AND2 (N7031, N7013, N1470);
and AND4 (N7032, N7029, N5523, N919, N5892);
xor XOR2 (N7033, N7017, N454);
and AND3 (N7034, N7014, N3236, N4303);
nand NAND4 (N7035, N7033, N4257, N5389, N5490);
and AND4 (N7036, N7021, N799, N1235, N4705);
not NOT1 (N7037, N7027);
or OR2 (N7038, N7035, N3793);
nand NAND3 (N7039, N7034, N4556, N6855);
nand NAND3 (N7040, N7036, N443, N4856);
nor NOR4 (N7041, N7025, N301, N6162, N4558);
buf BUF1 (N7042, N7037);
or OR3 (N7043, N7041, N3564, N5994);
or OR4 (N7044, N7030, N883, N4585, N1782);
nand NAND3 (N7045, N7039, N15, N5482);
xor XOR2 (N7046, N7026, N4560);
or OR2 (N7047, N7032, N2428);
nand NAND2 (N7048, N7044, N4070);
buf BUF1 (N7049, N7045);
or OR3 (N7050, N7028, N2478, N6136);
nand NAND4 (N7051, N7042, N5691, N4445, N2267);
or OR2 (N7052, N7049, N5943);
nor NOR3 (N7053, N7046, N1928, N362);
and AND3 (N7054, N7043, N1376, N6864);
and AND2 (N7055, N7050, N3684);
nor NOR2 (N7056, N7048, N6644);
nand NAND4 (N7057, N7051, N1716, N4270, N161);
xor XOR2 (N7058, N7055, N1922);
not NOT1 (N7059, N7053);
and AND4 (N7060, N7031, N3856, N4962, N525);
or OR3 (N7061, N7047, N2826, N3035);
nor NOR2 (N7062, N7059, N677);
and AND3 (N7063, N7058, N1711, N6556);
nor NOR3 (N7064, N7054, N3066, N3102);
buf BUF1 (N7065, N7061);
nand NAND3 (N7066, N7062, N5939, N6110);
nand NAND2 (N7067, N7038, N4488);
and AND4 (N7068, N7065, N272, N2364, N1236);
nand NAND4 (N7069, N7060, N5912, N3439, N4441);
or OR4 (N7070, N7064, N1907, N3090, N6413);
nand NAND3 (N7071, N7067, N2424, N3779);
not NOT1 (N7072, N7069);
nor NOR3 (N7073, N7072, N2152, N5065);
nor NOR3 (N7074, N7063, N4598, N201);
not NOT1 (N7075, N7066);
not NOT1 (N7076, N7068);
or OR3 (N7077, N7040, N938, N6048);
nand NAND3 (N7078, N7075, N6577, N5639);
nor NOR3 (N7079, N7056, N622, N4693);
nor NOR3 (N7080, N7070, N4500, N5976);
and AND3 (N7081, N7074, N4596, N2983);
or OR2 (N7082, N7081, N3157);
nor NOR3 (N7083, N7080, N5429, N1052);
or OR3 (N7084, N7083, N2591, N893);
nand NAND2 (N7085, N7078, N4427);
not NOT1 (N7086, N7084);
or OR4 (N7087, N7079, N5668, N5787, N5099);
buf BUF1 (N7088, N7071);
not NOT1 (N7089, N7085);
nor NOR4 (N7090, N7057, N376, N6044, N5559);
buf BUF1 (N7091, N7073);
nand NAND4 (N7092, N7086, N1295, N6506, N2955);
buf BUF1 (N7093, N7091);
buf BUF1 (N7094, N7052);
xor XOR2 (N7095, N7088, N6996);
not NOT1 (N7096, N7087);
not NOT1 (N7097, N7077);
xor XOR2 (N7098, N7093, N4823);
nand NAND3 (N7099, N7096, N3525, N1545);
xor XOR2 (N7100, N7090, N1265);
not NOT1 (N7101, N7097);
buf BUF1 (N7102, N7100);
and AND2 (N7103, N7099, N5582);
xor XOR2 (N7104, N7101, N6109);
xor XOR2 (N7105, N7104, N305);
nand NAND2 (N7106, N7094, N1834);
buf BUF1 (N7107, N7089);
buf BUF1 (N7108, N7082);
nor NOR2 (N7109, N7092, N323);
xor XOR2 (N7110, N7106, N7077);
not NOT1 (N7111, N7105);
buf BUF1 (N7112, N7111);
and AND3 (N7113, N7108, N5801, N6821);
or OR4 (N7114, N7095, N7024, N1857, N552);
and AND4 (N7115, N7076, N5387, N3793, N6718);
or OR4 (N7116, N7103, N1261, N2885, N4257);
and AND2 (N7117, N7115, N3051);
nor NOR4 (N7118, N7113, N5098, N162, N2624);
nand NAND3 (N7119, N7110, N4509, N2840);
not NOT1 (N7120, N7109);
buf BUF1 (N7121, N7107);
buf BUF1 (N7122, N7119);
nor NOR3 (N7123, N7120, N5654, N3022);
nor NOR4 (N7124, N7116, N2044, N6715, N3338);
not NOT1 (N7125, N7122);
buf BUF1 (N7126, N7112);
xor XOR2 (N7127, N7125, N2747);
not NOT1 (N7128, N7117);
buf BUF1 (N7129, N7123);
nor NOR4 (N7130, N7127, N2485, N5660, N2505);
not NOT1 (N7131, N7098);
nor NOR3 (N7132, N7118, N4470, N1034);
nor NOR2 (N7133, N7121, N6862);
nor NOR3 (N7134, N7130, N2831, N2348);
or OR2 (N7135, N7114, N2217);
not NOT1 (N7136, N7132);
buf BUF1 (N7137, N7128);
or OR2 (N7138, N7102, N5482);
and AND2 (N7139, N7133, N6080);
or OR2 (N7140, N7136, N4410);
buf BUF1 (N7141, N7139);
xor XOR2 (N7142, N7138, N79);
and AND4 (N7143, N7141, N6683, N2842, N1029);
and AND3 (N7144, N7142, N1429, N4489);
not NOT1 (N7145, N7140);
not NOT1 (N7146, N7144);
buf BUF1 (N7147, N7129);
and AND4 (N7148, N7137, N3270, N6240, N1648);
not NOT1 (N7149, N7145);
not NOT1 (N7150, N7126);
buf BUF1 (N7151, N7147);
or OR3 (N7152, N7150, N4855, N3942);
nor NOR3 (N7153, N7148, N5541, N1617);
not NOT1 (N7154, N7124);
nor NOR3 (N7155, N7152, N3731, N6601);
nor NOR2 (N7156, N7153, N1022);
not NOT1 (N7157, N7134);
nand NAND2 (N7158, N7154, N3155);
buf BUF1 (N7159, N7143);
nor NOR4 (N7160, N7158, N6502, N6929, N2726);
xor XOR2 (N7161, N7157, N2128);
xor XOR2 (N7162, N7149, N3798);
nand NAND3 (N7163, N7131, N4788, N1257);
and AND3 (N7164, N7151, N201, N3101);
not NOT1 (N7165, N7135);
buf BUF1 (N7166, N7163);
xor XOR2 (N7167, N7165, N5090);
not NOT1 (N7168, N7167);
buf BUF1 (N7169, N7146);
and AND4 (N7170, N7161, N419, N5369, N4039);
nor NOR4 (N7171, N7159, N3694, N5467, N1987);
and AND4 (N7172, N7170, N579, N5190, N6011);
xor XOR2 (N7173, N7162, N800);
xor XOR2 (N7174, N7169, N2140);
or OR3 (N7175, N7174, N6958, N7006);
and AND4 (N7176, N7172, N1010, N1833, N3634);
xor XOR2 (N7177, N7164, N85);
buf BUF1 (N7178, N7155);
buf BUF1 (N7179, N7177);
and AND2 (N7180, N7176, N5828);
xor XOR2 (N7181, N7160, N6518);
or OR3 (N7182, N7178, N2039, N1077);
and AND3 (N7183, N7181, N5367, N666);
not NOT1 (N7184, N7171);
not NOT1 (N7185, N7180);
nor NOR3 (N7186, N7166, N82, N2113);
xor XOR2 (N7187, N7183, N3703);
buf BUF1 (N7188, N7187);
xor XOR2 (N7189, N7182, N1909);
xor XOR2 (N7190, N7168, N7097);
or OR3 (N7191, N7156, N276, N5184);
xor XOR2 (N7192, N7189, N640);
or OR3 (N7193, N7179, N7012, N225);
not NOT1 (N7194, N7191);
or OR2 (N7195, N7194, N6400);
nand NAND4 (N7196, N7195, N2319, N2040, N3589);
nand NAND3 (N7197, N7193, N4395, N345);
nor NOR2 (N7198, N7173, N1101);
or OR3 (N7199, N7197, N3979, N1454);
xor XOR2 (N7200, N7186, N4552);
not NOT1 (N7201, N7199);
buf BUF1 (N7202, N7184);
or OR4 (N7203, N7202, N3355, N147, N1982);
nand NAND3 (N7204, N7188, N2079, N558);
nor NOR4 (N7205, N7203, N6008, N7041, N5930);
or OR2 (N7206, N7185, N6979);
buf BUF1 (N7207, N7201);
or OR3 (N7208, N7198, N2579, N2778);
xor XOR2 (N7209, N7206, N5256);
xor XOR2 (N7210, N7192, N5816);
nand NAND2 (N7211, N7200, N4454);
or OR4 (N7212, N7210, N3133, N4204, N5007);
and AND3 (N7213, N7190, N2625, N2914);
nor NOR2 (N7214, N7209, N6814);
not NOT1 (N7215, N7205);
and AND3 (N7216, N7211, N1540, N831);
xor XOR2 (N7217, N7175, N3679);
not NOT1 (N7218, N7215);
buf BUF1 (N7219, N7196);
and AND4 (N7220, N7218, N1647, N224, N1982);
or OR2 (N7221, N7213, N2254);
and AND2 (N7222, N7204, N1793);
and AND2 (N7223, N7222, N104);
nand NAND4 (N7224, N7214, N6824, N663, N115);
buf BUF1 (N7225, N7223);
nand NAND2 (N7226, N7208, N2126);
nand NAND2 (N7227, N7219, N3591);
xor XOR2 (N7228, N7216, N6322);
not NOT1 (N7229, N7227);
not NOT1 (N7230, N7221);
nor NOR3 (N7231, N7212, N2647, N5486);
or OR3 (N7232, N7231, N5964, N3956);
nand NAND4 (N7233, N7224, N3093, N3687, N543);
xor XOR2 (N7234, N7220, N18);
buf BUF1 (N7235, N7234);
and AND4 (N7236, N7229, N318, N4350, N5978);
nand NAND4 (N7237, N7226, N1507, N3979, N3834);
and AND2 (N7238, N7235, N568);
nand NAND4 (N7239, N7207, N2284, N5298, N3791);
not NOT1 (N7240, N7217);
xor XOR2 (N7241, N7233, N1786);
buf BUF1 (N7242, N7228);
or OR4 (N7243, N7225, N749, N2876, N7097);
buf BUF1 (N7244, N7240);
buf BUF1 (N7245, N7242);
xor XOR2 (N7246, N7243, N3666);
nand NAND3 (N7247, N7238, N5568, N5898);
or OR2 (N7248, N7236, N1563);
or OR3 (N7249, N7237, N5134, N6712);
or OR2 (N7250, N7244, N4543);
buf BUF1 (N7251, N7241);
buf BUF1 (N7252, N7248);
and AND4 (N7253, N7249, N3217, N2602, N4985);
or OR3 (N7254, N7250, N512, N6050);
xor XOR2 (N7255, N7252, N576);
and AND3 (N7256, N7255, N5487, N3955);
xor XOR2 (N7257, N7254, N4363);
xor XOR2 (N7258, N7232, N5903);
and AND4 (N7259, N7256, N1837, N2026, N1007);
xor XOR2 (N7260, N7230, N469);
or OR2 (N7261, N7259, N4276);
xor XOR2 (N7262, N7261, N2602);
nand NAND4 (N7263, N7253, N718, N6021, N6868);
xor XOR2 (N7264, N7257, N428);
nor NOR3 (N7265, N7264, N5366, N971);
and AND4 (N7266, N7246, N3501, N1087, N648);
or OR4 (N7267, N7263, N4834, N432, N6079);
or OR4 (N7268, N7245, N2134, N3291, N5617);
or OR2 (N7269, N7251, N2715);
not NOT1 (N7270, N7269);
nand NAND2 (N7271, N7258, N4745);
or OR2 (N7272, N7265, N977);
and AND3 (N7273, N7267, N5736, N2357);
nor NOR3 (N7274, N7260, N5937, N374);
or OR2 (N7275, N7266, N6823);
xor XOR2 (N7276, N7273, N6435);
buf BUF1 (N7277, N7247);
nor NOR4 (N7278, N7277, N6776, N4932, N771);
or OR4 (N7279, N7272, N4663, N6151, N5709);
and AND3 (N7280, N7271, N6812, N3352);
not NOT1 (N7281, N7239);
xor XOR2 (N7282, N7276, N421);
nor NOR4 (N7283, N7268, N754, N3565, N709);
not NOT1 (N7284, N7283);
or OR3 (N7285, N7279, N2660, N5345);
or OR2 (N7286, N7280, N4231);
xor XOR2 (N7287, N7281, N4303);
nand NAND3 (N7288, N7270, N2546, N1961);
xor XOR2 (N7289, N7275, N5499);
nor NOR4 (N7290, N7282, N4793, N5322, N6659);
or OR3 (N7291, N7288, N4731, N4032);
and AND2 (N7292, N7286, N2058);
and AND3 (N7293, N7262, N196, N3236);
not NOT1 (N7294, N7292);
nor NOR2 (N7295, N7287, N84);
and AND2 (N7296, N7294, N659);
nor NOR3 (N7297, N7291, N4907, N3192);
and AND2 (N7298, N7290, N6664);
or OR3 (N7299, N7298, N4835, N2237);
nand NAND3 (N7300, N7284, N5855, N5240);
nor NOR4 (N7301, N7285, N5598, N899, N5532);
nor NOR4 (N7302, N7299, N4111, N6195, N1932);
and AND2 (N7303, N7296, N5897);
not NOT1 (N7304, N7300);
or OR4 (N7305, N7297, N5254, N7278, N7075);
buf BUF1 (N7306, N7156);
not NOT1 (N7307, N7293);
not NOT1 (N7308, N7301);
buf BUF1 (N7309, N7302);
or OR2 (N7310, N7308, N3736);
buf BUF1 (N7311, N7305);
xor XOR2 (N7312, N7304, N2431);
nor NOR3 (N7313, N7306, N2581, N6533);
buf BUF1 (N7314, N7309);
or OR3 (N7315, N7312, N3177, N6870);
buf BUF1 (N7316, N7303);
nand NAND3 (N7317, N7274, N3049, N6901);
xor XOR2 (N7318, N7315, N3632);
nand NAND3 (N7319, N7317, N6265, N310);
xor XOR2 (N7320, N7310, N6861);
and AND2 (N7321, N7289, N2124);
or OR2 (N7322, N7314, N4552);
nor NOR3 (N7323, N7313, N5835, N1435);
not NOT1 (N7324, N7316);
buf BUF1 (N7325, N7319);
nand NAND4 (N7326, N7324, N5450, N6597, N2156);
nor NOR3 (N7327, N7325, N187, N6207);
and AND2 (N7328, N7322, N2849);
xor XOR2 (N7329, N7327, N5209);
xor XOR2 (N7330, N7311, N186);
or OR4 (N7331, N7329, N4981, N3557, N5991);
nand NAND4 (N7332, N7330, N4926, N2939, N5581);
buf BUF1 (N7333, N7295);
nor NOR4 (N7334, N7331, N4052, N5363, N3025);
not NOT1 (N7335, N7332);
buf BUF1 (N7336, N7307);
xor XOR2 (N7337, N7326, N6600);
nor NOR2 (N7338, N7320, N3677);
and AND4 (N7339, N7321, N3513, N3540, N1972);
or OR4 (N7340, N7338, N6271, N3374, N2223);
not NOT1 (N7341, N7335);
xor XOR2 (N7342, N7336, N4604);
nand NAND3 (N7343, N7334, N2184, N5886);
buf BUF1 (N7344, N7318);
and AND2 (N7345, N7337, N1923);
and AND2 (N7346, N7328, N2785);
or OR4 (N7347, N7333, N6113, N6330, N226);
xor XOR2 (N7348, N7342, N4116);
buf BUF1 (N7349, N7343);
buf BUF1 (N7350, N7347);
xor XOR2 (N7351, N7345, N1198);
xor XOR2 (N7352, N7341, N6600);
not NOT1 (N7353, N7346);
nor NOR2 (N7354, N7350, N2862);
and AND4 (N7355, N7354, N3397, N1677, N2661);
and AND2 (N7356, N7355, N1060);
and AND3 (N7357, N7349, N3581, N507);
nor NOR3 (N7358, N7340, N5720, N5656);
not NOT1 (N7359, N7357);
or OR4 (N7360, N7351, N4092, N6612, N7029);
or OR4 (N7361, N7358, N3196, N3395, N6695);
or OR3 (N7362, N7323, N1474, N5122);
buf BUF1 (N7363, N7344);
nand NAND2 (N7364, N7353, N4773);
or OR4 (N7365, N7348, N2690, N6585, N3844);
nor NOR3 (N7366, N7352, N4849, N119);
nand NAND3 (N7367, N7365, N559, N1994);
nor NOR4 (N7368, N7364, N4343, N1106, N6539);
nor NOR3 (N7369, N7368, N5154, N7339);
nor NOR2 (N7370, N1706, N828);
nor NOR2 (N7371, N7356, N1105);
or OR2 (N7372, N7359, N2304);
and AND2 (N7373, N7367, N2053);
nor NOR3 (N7374, N7362, N5441, N5775);
xor XOR2 (N7375, N7366, N5047);
or OR4 (N7376, N7375, N922, N2245, N6922);
buf BUF1 (N7377, N7373);
nor NOR3 (N7378, N7371, N2433, N2206);
xor XOR2 (N7379, N7363, N1692);
not NOT1 (N7380, N7376);
not NOT1 (N7381, N7372);
or OR2 (N7382, N7369, N2470);
not NOT1 (N7383, N7377);
buf BUF1 (N7384, N7360);
nand NAND2 (N7385, N7370, N983);
xor XOR2 (N7386, N7384, N6761);
or OR2 (N7387, N7383, N3282);
nand NAND4 (N7388, N7386, N2245, N4556, N3978);
xor XOR2 (N7389, N7382, N3558);
nand NAND2 (N7390, N7387, N4454);
or OR2 (N7391, N7390, N6225);
nand NAND4 (N7392, N7378, N3443, N2251, N6423);
and AND2 (N7393, N7391, N4361);
buf BUF1 (N7394, N7361);
not NOT1 (N7395, N7374);
and AND2 (N7396, N7394, N1267);
not NOT1 (N7397, N7393);
and AND3 (N7398, N7385, N6603, N2100);
or OR4 (N7399, N7397, N3972, N3018, N4202);
not NOT1 (N7400, N7389);
not NOT1 (N7401, N7400);
xor XOR2 (N7402, N7379, N3001);
nor NOR3 (N7403, N7388, N5116, N3477);
nor NOR4 (N7404, N7395, N7144, N5853, N4966);
xor XOR2 (N7405, N7396, N6716);
and AND3 (N7406, N7401, N449, N5393);
nor NOR4 (N7407, N7392, N1946, N44, N4712);
not NOT1 (N7408, N7406);
or OR4 (N7409, N7403, N3419, N4848, N7259);
nor NOR3 (N7410, N7399, N1337, N5259);
not NOT1 (N7411, N7408);
or OR2 (N7412, N7398, N6339);
nand NAND4 (N7413, N7411, N5329, N1287, N1180);
nor NOR2 (N7414, N7381, N1954);
and AND3 (N7415, N7405, N6546, N1692);
or OR4 (N7416, N7410, N7246, N2064, N5157);
xor XOR2 (N7417, N7404, N201);
buf BUF1 (N7418, N7380);
nor NOR4 (N7419, N7416, N964, N6875, N1461);
and AND4 (N7420, N7413, N5874, N1943, N7130);
not NOT1 (N7421, N7417);
nor NOR2 (N7422, N7414, N4084);
and AND4 (N7423, N7419, N7251, N2098, N4337);
xor XOR2 (N7424, N7412, N286);
buf BUF1 (N7425, N7418);
nand NAND3 (N7426, N7425, N4661, N566);
or OR2 (N7427, N7424, N5271);
buf BUF1 (N7428, N7422);
nand NAND4 (N7429, N7415, N3740, N4468, N2789);
nor NOR3 (N7430, N7426, N6533, N1326);
or OR2 (N7431, N7427, N7329);
and AND4 (N7432, N7421, N4271, N889, N1584);
xor XOR2 (N7433, N7420, N388);
nand NAND2 (N7434, N7402, N566);
and AND2 (N7435, N7409, N4612);
buf BUF1 (N7436, N7432);
not NOT1 (N7437, N7428);
nor NOR3 (N7438, N7423, N7139, N5398);
and AND3 (N7439, N7431, N6173, N1670);
not NOT1 (N7440, N7437);
not NOT1 (N7441, N7434);
or OR3 (N7442, N7439, N2081, N1795);
nand NAND4 (N7443, N7407, N1593, N5853, N4569);
xor XOR2 (N7444, N7440, N6974);
not NOT1 (N7445, N7430);
or OR2 (N7446, N7441, N6690);
nor NOR2 (N7447, N7438, N231);
or OR2 (N7448, N7442, N1416);
nand NAND2 (N7449, N7435, N4772);
not NOT1 (N7450, N7429);
or OR2 (N7451, N7443, N878);
xor XOR2 (N7452, N7444, N1530);
nand NAND2 (N7453, N7449, N6223);
and AND3 (N7454, N7445, N1676, N2666);
buf BUF1 (N7455, N7450);
buf BUF1 (N7456, N7455);
buf BUF1 (N7457, N7448);
or OR2 (N7458, N7451, N1826);
not NOT1 (N7459, N7447);
or OR2 (N7460, N7452, N3605);
and AND2 (N7461, N7436, N2787);
or OR2 (N7462, N7458, N953);
not NOT1 (N7463, N7453);
buf BUF1 (N7464, N7459);
or OR3 (N7465, N7446, N2281, N7307);
buf BUF1 (N7466, N7465);
nand NAND2 (N7467, N7454, N4645);
and AND2 (N7468, N7457, N5258);
buf BUF1 (N7469, N7456);
nor NOR3 (N7470, N7467, N4346, N6773);
nand NAND4 (N7471, N7470, N3361, N1829, N1856);
nor NOR3 (N7472, N7461, N4891, N3288);
buf BUF1 (N7473, N7463);
buf BUF1 (N7474, N7473);
xor XOR2 (N7475, N7472, N7457);
xor XOR2 (N7476, N7469, N4749);
or OR2 (N7477, N7474, N4399);
or OR4 (N7478, N7433, N3048, N6263, N1339);
buf BUF1 (N7479, N7478);
and AND3 (N7480, N7471, N5959, N1074);
nand NAND2 (N7481, N7477, N4025);
and AND4 (N7482, N7480, N3440, N1527, N2499);
and AND3 (N7483, N7482, N717, N7421);
not NOT1 (N7484, N7479);
or OR4 (N7485, N7466, N2385, N7056, N1572);
nand NAND2 (N7486, N7468, N741);
nor NOR3 (N7487, N7462, N4578, N4667);
nand NAND2 (N7488, N7476, N7397);
not NOT1 (N7489, N7485);
or OR4 (N7490, N7460, N4651, N5376, N3218);
nand NAND4 (N7491, N7484, N1903, N1860, N5523);
nor NOR2 (N7492, N7481, N3184);
nand NAND2 (N7493, N7491, N152);
nand NAND2 (N7494, N7486, N1146);
nand NAND2 (N7495, N7490, N240);
or OR2 (N7496, N7495, N3325);
nor NOR2 (N7497, N7494, N699);
buf BUF1 (N7498, N7487);
nand NAND2 (N7499, N7493, N2623);
xor XOR2 (N7500, N7496, N3360);
nor NOR3 (N7501, N7499, N668, N733);
and AND3 (N7502, N7492, N6348, N200);
and AND3 (N7503, N7497, N6927, N1555);
buf BUF1 (N7504, N7489);
or OR2 (N7505, N7502, N89);
xor XOR2 (N7506, N7500, N4697);
nand NAND4 (N7507, N7506, N3052, N2525, N5242);
buf BUF1 (N7508, N7501);
nor NOR2 (N7509, N7464, N5608);
or OR3 (N7510, N7508, N4710, N6167);
xor XOR2 (N7511, N7507, N579);
or OR3 (N7512, N7511, N5050, N6425);
or OR3 (N7513, N7504, N5099, N3121);
or OR3 (N7514, N7475, N1717, N864);
buf BUF1 (N7515, N7509);
nand NAND2 (N7516, N7514, N3187);
and AND2 (N7517, N7513, N809);
not NOT1 (N7518, N7512);
or OR3 (N7519, N7518, N3223, N1404);
not NOT1 (N7520, N7515);
nand NAND3 (N7521, N7517, N5860, N2114);
xor XOR2 (N7522, N7510, N2501);
xor XOR2 (N7523, N7521, N6348);
or OR4 (N7524, N7516, N3878, N2990, N2669);
buf BUF1 (N7525, N7505);
and AND4 (N7526, N7483, N4337, N4546, N6413);
nand NAND4 (N7527, N7519, N6556, N7026, N6229);
not NOT1 (N7528, N7503);
and AND2 (N7529, N7528, N4780);
xor XOR2 (N7530, N7525, N396);
buf BUF1 (N7531, N7520);
nand NAND2 (N7532, N7529, N2312);
buf BUF1 (N7533, N7526);
or OR4 (N7534, N7523, N3905, N1094, N6016);
not NOT1 (N7535, N7530);
buf BUF1 (N7536, N7522);
not NOT1 (N7537, N7534);
and AND3 (N7538, N7498, N2891, N908);
xor XOR2 (N7539, N7531, N7050);
or OR2 (N7540, N7536, N4221);
xor XOR2 (N7541, N7537, N3996);
and AND4 (N7542, N7488, N5910, N5084, N358);
nor NOR2 (N7543, N7535, N6944);
or OR2 (N7544, N7533, N2132);
nor NOR3 (N7545, N7538, N7345, N4187);
xor XOR2 (N7546, N7541, N2365);
and AND2 (N7547, N7545, N2378);
xor XOR2 (N7548, N7540, N6174);
buf BUF1 (N7549, N7547);
and AND3 (N7550, N7527, N4629, N276);
nor NOR2 (N7551, N7542, N3127);
or OR3 (N7552, N7543, N1777, N3385);
or OR2 (N7553, N7532, N4698);
xor XOR2 (N7554, N7553, N3593);
nand NAND4 (N7555, N7524, N3830, N4450, N3258);
and AND2 (N7556, N7554, N6223);
not NOT1 (N7557, N7544);
and AND3 (N7558, N7551, N1516, N4369);
not NOT1 (N7559, N7550);
buf BUF1 (N7560, N7557);
nor NOR3 (N7561, N7560, N534, N6456);
and AND4 (N7562, N7548, N1711, N6948, N6291);
xor XOR2 (N7563, N7549, N3541);
or OR4 (N7564, N7558, N5743, N5397, N164);
buf BUF1 (N7565, N7555);
and AND3 (N7566, N7565, N1335, N5159);
or OR4 (N7567, N7564, N6262, N5855, N4462);
and AND4 (N7568, N7552, N1678, N5141, N5296);
buf BUF1 (N7569, N7561);
buf BUF1 (N7570, N7546);
nand NAND2 (N7571, N7556, N3249);
nand NAND3 (N7572, N7568, N5674, N3617);
xor XOR2 (N7573, N7571, N970);
xor XOR2 (N7574, N7539, N6428);
or OR3 (N7575, N7574, N2223, N3208);
not NOT1 (N7576, N7563);
or OR3 (N7577, N7576, N3243, N5674);
not NOT1 (N7578, N7566);
not NOT1 (N7579, N7567);
not NOT1 (N7580, N7579);
or OR2 (N7581, N7570, N6544);
xor XOR2 (N7582, N7559, N3854);
buf BUF1 (N7583, N7582);
and AND3 (N7584, N7583, N5526, N3154);
not NOT1 (N7585, N7581);
xor XOR2 (N7586, N7572, N4721);
buf BUF1 (N7587, N7584);
not NOT1 (N7588, N7578);
xor XOR2 (N7589, N7580, N1224);
buf BUF1 (N7590, N7577);
or OR4 (N7591, N7575, N157, N7562, N506);
nor NOR2 (N7592, N7205, N4711);
nor NOR2 (N7593, N7588, N1146);
nor NOR4 (N7594, N7591, N6069, N2468, N7412);
and AND4 (N7595, N7590, N3861, N3403, N3425);
or OR2 (N7596, N7595, N144);
not NOT1 (N7597, N7573);
or OR2 (N7598, N7587, N3461);
or OR2 (N7599, N7594, N3916);
nor NOR3 (N7600, N7598, N2295, N1715);
or OR4 (N7601, N7599, N1975, N1017, N5623);
not NOT1 (N7602, N7596);
or OR2 (N7603, N7597, N166);
xor XOR2 (N7604, N7602, N3110);
or OR3 (N7605, N7601, N3336, N1610);
xor XOR2 (N7606, N7569, N6338);
or OR2 (N7607, N7589, N6104);
buf BUF1 (N7608, N7604);
and AND4 (N7609, N7607, N2244, N2425, N1594);
and AND3 (N7610, N7600, N7108, N2948);
nand NAND4 (N7611, N7610, N2189, N7174, N1070);
or OR2 (N7612, N7608, N2904);
xor XOR2 (N7613, N7593, N5339);
or OR3 (N7614, N7605, N3485, N980);
nor NOR4 (N7615, N7606, N26, N2017, N1502);
not NOT1 (N7616, N7603);
and AND4 (N7617, N7614, N5580, N5183, N4125);
and AND3 (N7618, N7585, N5208, N5972);
or OR3 (N7619, N7618, N2058, N303);
or OR4 (N7620, N7613, N4387, N3313, N7227);
and AND4 (N7621, N7615, N3481, N5919, N2894);
nand NAND2 (N7622, N7620, N2850);
nand NAND3 (N7623, N7621, N2308, N1180);
nor NOR2 (N7624, N7617, N5376);
buf BUF1 (N7625, N7616);
not NOT1 (N7626, N7619);
or OR3 (N7627, N7611, N592, N7559);
or OR4 (N7628, N7624, N3037, N2546, N1851);
nand NAND2 (N7629, N7623, N6213);
nor NOR2 (N7630, N7612, N672);
xor XOR2 (N7631, N7630, N613);
nor NOR3 (N7632, N7609, N3482, N887);
nand NAND4 (N7633, N7628, N6307, N1573, N5073);
not NOT1 (N7634, N7627);
and AND2 (N7635, N7622, N7613);
nor NOR3 (N7636, N7635, N356, N4050);
nand NAND4 (N7637, N7631, N348, N5577, N2157);
buf BUF1 (N7638, N7637);
nor NOR3 (N7639, N7636, N1278, N342);
buf BUF1 (N7640, N7586);
nor NOR2 (N7641, N7633, N1065);
not NOT1 (N7642, N7639);
and AND2 (N7643, N7642, N2606);
or OR2 (N7644, N7638, N4334);
buf BUF1 (N7645, N7644);
buf BUF1 (N7646, N7592);
buf BUF1 (N7647, N7643);
or OR4 (N7648, N7634, N5042, N3011, N6577);
not NOT1 (N7649, N7647);
nand NAND4 (N7650, N7648, N1862, N2684, N506);
or OR3 (N7651, N7646, N7034, N7036);
nor NOR2 (N7652, N7651, N6587);
and AND4 (N7653, N7652, N333, N6613, N1458);
and AND4 (N7654, N7641, N3479, N6361, N893);
and AND4 (N7655, N7632, N7527, N4233, N6330);
nand NAND3 (N7656, N7655, N1672, N4408);
or OR3 (N7657, N7640, N5508, N316);
nand NAND4 (N7658, N7650, N1042, N1313, N689);
xor XOR2 (N7659, N7626, N4999);
or OR4 (N7660, N7657, N7190, N1467, N1945);
xor XOR2 (N7661, N7625, N1939);
not NOT1 (N7662, N7645);
not NOT1 (N7663, N7662);
and AND2 (N7664, N7658, N3048);
buf BUF1 (N7665, N7661);
nand NAND3 (N7666, N7649, N2915, N4145);
nand NAND3 (N7667, N7663, N7278, N2027);
nor NOR2 (N7668, N7666, N3899);
and AND3 (N7669, N7667, N3166, N5728);
or OR3 (N7670, N7659, N405, N5914);
xor XOR2 (N7671, N7669, N1900);
nor NOR4 (N7672, N7670, N6414, N2524, N5004);
nor NOR2 (N7673, N7656, N5942);
and AND3 (N7674, N7665, N7350, N2464);
buf BUF1 (N7675, N7660);
nor NOR4 (N7676, N7675, N386, N2656, N6622);
nor NOR3 (N7677, N7673, N6896, N2321);
xor XOR2 (N7678, N7671, N837);
not NOT1 (N7679, N7668);
buf BUF1 (N7680, N7674);
and AND4 (N7681, N7654, N3836, N5824, N5571);
and AND4 (N7682, N7672, N3255, N7021, N4777);
nor NOR2 (N7683, N7653, N3640);
or OR3 (N7684, N7683, N1062, N5769);
nor NOR4 (N7685, N7681, N6263, N7361, N1658);
nor NOR2 (N7686, N7678, N4013);
and AND4 (N7687, N7682, N4039, N3156, N1528);
nor NOR4 (N7688, N7629, N1365, N2733, N6797);
or OR2 (N7689, N7687, N7593);
nand NAND3 (N7690, N7679, N983, N451);
xor XOR2 (N7691, N7684, N2789);
or OR3 (N7692, N7664, N4813, N6775);
nand NAND2 (N7693, N7680, N2097);
xor XOR2 (N7694, N7676, N630);
nand NAND3 (N7695, N7689, N3620, N6545);
xor XOR2 (N7696, N7691, N4994);
nand NAND3 (N7697, N7677, N5390, N7661);
not NOT1 (N7698, N7695);
nand NAND2 (N7699, N7693, N7206);
nor NOR2 (N7700, N7696, N6585);
xor XOR2 (N7701, N7697, N68);
not NOT1 (N7702, N7701);
and AND3 (N7703, N7694, N5067, N3591);
nand NAND4 (N7704, N7700, N703, N4581, N4604);
or OR2 (N7705, N7704, N2620);
not NOT1 (N7706, N7692);
buf BUF1 (N7707, N7706);
and AND4 (N7708, N7703, N4436, N7604, N1086);
xor XOR2 (N7709, N7705, N1249);
and AND3 (N7710, N7690, N3024, N5016);
nand NAND4 (N7711, N7709, N316, N6544, N5677);
nand NAND3 (N7712, N7711, N6238, N567);
buf BUF1 (N7713, N7710);
or OR4 (N7714, N7685, N2314, N4659, N1829);
xor XOR2 (N7715, N7699, N2257);
and AND2 (N7716, N7713, N5642);
buf BUF1 (N7717, N7716);
not NOT1 (N7718, N7688);
or OR3 (N7719, N7718, N4713, N4842);
nor NOR3 (N7720, N7702, N6823, N3020);
not NOT1 (N7721, N7708);
nand NAND2 (N7722, N7717, N1659);
nor NOR3 (N7723, N7720, N7149, N5214);
nand NAND3 (N7724, N7698, N3987, N2951);
or OR4 (N7725, N7724, N982, N2938, N2586);
and AND4 (N7726, N7686, N1532, N621, N4330);
nor NOR2 (N7727, N7712, N4131);
and AND2 (N7728, N7707, N5971);
xor XOR2 (N7729, N7726, N4813);
nor NOR2 (N7730, N7725, N1065);
not NOT1 (N7731, N7728);
nand NAND3 (N7732, N7727, N1711, N1911);
not NOT1 (N7733, N7731);
xor XOR2 (N7734, N7723, N3223);
xor XOR2 (N7735, N7722, N3506);
or OR4 (N7736, N7714, N5857, N679, N6553);
nor NOR3 (N7737, N7721, N1066, N6085);
xor XOR2 (N7738, N7733, N7083);
not NOT1 (N7739, N7734);
xor XOR2 (N7740, N7739, N6320);
not NOT1 (N7741, N7736);
not NOT1 (N7742, N7740);
or OR4 (N7743, N7741, N772, N146, N744);
buf BUF1 (N7744, N7715);
and AND2 (N7745, N7744, N983);
not NOT1 (N7746, N7730);
nor NOR4 (N7747, N7732, N3219, N6041, N4280);
xor XOR2 (N7748, N7742, N2783);
buf BUF1 (N7749, N7735);
not NOT1 (N7750, N7747);
or OR3 (N7751, N7750, N410, N6607);
buf BUF1 (N7752, N7729);
or OR2 (N7753, N7752, N2031);
and AND4 (N7754, N7745, N199, N176, N6579);
nand NAND3 (N7755, N7743, N7632, N1265);
not NOT1 (N7756, N7754);
nor NOR3 (N7757, N7756, N7580, N7045);
and AND4 (N7758, N7738, N7202, N2667, N7001);
nand NAND4 (N7759, N7719, N99, N5734, N3296);
nand NAND2 (N7760, N7757, N2211);
buf BUF1 (N7761, N7749);
not NOT1 (N7762, N7748);
buf BUF1 (N7763, N7760);
nor NOR3 (N7764, N7758, N1609, N2882);
or OR2 (N7765, N7753, N6908);
and AND4 (N7766, N7751, N7413, N7157, N3263);
and AND4 (N7767, N7765, N5938, N2701, N752);
not NOT1 (N7768, N7763);
buf BUF1 (N7769, N7746);
not NOT1 (N7770, N7764);
and AND3 (N7771, N7767, N6393, N6469);
nor NOR4 (N7772, N7759, N7483, N123, N6881);
xor XOR2 (N7773, N7771, N4584);
nor NOR3 (N7774, N7755, N3689, N5072);
nand NAND2 (N7775, N7768, N6698);
xor XOR2 (N7776, N7737, N1684);
and AND3 (N7777, N7761, N5739, N1147);
nand NAND2 (N7778, N7770, N1377);
and AND2 (N7779, N7777, N4035);
buf BUF1 (N7780, N7778);
and AND3 (N7781, N7773, N2646, N1338);
or OR3 (N7782, N7769, N7698, N4213);
nand NAND3 (N7783, N7775, N3221, N2192);
not NOT1 (N7784, N7782);
nand NAND2 (N7785, N7781, N511);
buf BUF1 (N7786, N7785);
or OR3 (N7787, N7774, N7611, N6627);
buf BUF1 (N7788, N7783);
or OR3 (N7789, N7784, N1948, N5134);
buf BUF1 (N7790, N7789);
or OR4 (N7791, N7772, N4701, N4130, N1860);
nor NOR2 (N7792, N7766, N1853);
nor NOR4 (N7793, N7790, N4160, N2476, N6960);
buf BUF1 (N7794, N7786);
nor NOR3 (N7795, N7794, N1156, N5768);
nor NOR3 (N7796, N7776, N362, N5441);
buf BUF1 (N7797, N7779);
not NOT1 (N7798, N7797);
not NOT1 (N7799, N7795);
nand NAND2 (N7800, N7793, N2038);
nor NOR3 (N7801, N7791, N2092, N7295);
not NOT1 (N7802, N7796);
nand NAND4 (N7803, N7788, N3350, N2461, N1945);
and AND3 (N7804, N7801, N6897, N2401);
buf BUF1 (N7805, N7780);
buf BUF1 (N7806, N7802);
buf BUF1 (N7807, N7804);
not NOT1 (N7808, N7798);
xor XOR2 (N7809, N7806, N6315);
nand NAND2 (N7810, N7803, N5515);
or OR3 (N7811, N7810, N7421, N5934);
nor NOR3 (N7812, N7762, N6018, N3117);
not NOT1 (N7813, N7812);
nor NOR4 (N7814, N7807, N7414, N5893, N5534);
xor XOR2 (N7815, N7805, N3158);
buf BUF1 (N7816, N7814);
not NOT1 (N7817, N7799);
or OR3 (N7818, N7811, N5191, N7049);
nand NAND4 (N7819, N7787, N1747, N992, N2484);
buf BUF1 (N7820, N7813);
nor NOR3 (N7821, N7792, N7733, N1043);
and AND4 (N7822, N7816, N3723, N5948, N551);
not NOT1 (N7823, N7809);
not NOT1 (N7824, N7819);
nand NAND2 (N7825, N7808, N7777);
nor NOR2 (N7826, N7818, N3830);
not NOT1 (N7827, N7820);
or OR4 (N7828, N7815, N6434, N6558, N3798);
xor XOR2 (N7829, N7823, N7373);
and AND4 (N7830, N7824, N1335, N283, N474);
nand NAND3 (N7831, N7827, N6246, N1772);
and AND2 (N7832, N7817, N760);
xor XOR2 (N7833, N7821, N2390);
nand NAND2 (N7834, N7830, N6954);
buf BUF1 (N7835, N7834);
not NOT1 (N7836, N7835);
and AND2 (N7837, N7833, N6539);
and AND4 (N7838, N7831, N3607, N2145, N4949);
buf BUF1 (N7839, N7838);
and AND3 (N7840, N7837, N2128, N2746);
and AND3 (N7841, N7822, N7839, N6976);
nand NAND2 (N7842, N2109, N7191);
or OR3 (N7843, N7829, N2630, N2991);
buf BUF1 (N7844, N7828);
nand NAND2 (N7845, N7826, N6161);
xor XOR2 (N7846, N7836, N909);
nand NAND3 (N7847, N7832, N377, N2670);
xor XOR2 (N7848, N7846, N7390);
xor XOR2 (N7849, N7840, N6404);
or OR2 (N7850, N7847, N1104);
nand NAND4 (N7851, N7844, N6688, N4028, N5065);
nand NAND2 (N7852, N7849, N6072);
or OR2 (N7853, N7843, N5945);
nor NOR2 (N7854, N7848, N904);
nor NOR3 (N7855, N7854, N4338, N6874);
not NOT1 (N7856, N7845);
xor XOR2 (N7857, N7856, N6626);
and AND4 (N7858, N7850, N2975, N4020, N6090);
nor NOR4 (N7859, N7842, N1250, N5118, N7546);
nor NOR4 (N7860, N7855, N3792, N4597, N119);
xor XOR2 (N7861, N7857, N1609);
not NOT1 (N7862, N7852);
or OR2 (N7863, N7851, N2704);
or OR3 (N7864, N7861, N2219, N3764);
or OR3 (N7865, N7841, N7666, N4820);
or OR4 (N7866, N7800, N7281, N2882, N2887);
xor XOR2 (N7867, N7859, N6917);
nor NOR3 (N7868, N7865, N2144, N4268);
not NOT1 (N7869, N7863);
xor XOR2 (N7870, N7864, N12);
and AND4 (N7871, N7853, N3735, N2126, N219);
not NOT1 (N7872, N7868);
not NOT1 (N7873, N7825);
xor XOR2 (N7874, N7871, N5329);
buf BUF1 (N7875, N7874);
not NOT1 (N7876, N7872);
xor XOR2 (N7877, N7867, N5282);
nor NOR2 (N7878, N7873, N922);
not NOT1 (N7879, N7860);
nand NAND2 (N7880, N7862, N4346);
buf BUF1 (N7881, N7879);
and AND4 (N7882, N7866, N4099, N6816, N612);
not NOT1 (N7883, N7858);
nand NAND4 (N7884, N7870, N7726, N5388, N7570);
and AND4 (N7885, N7882, N2568, N843, N7103);
buf BUF1 (N7886, N7885);
not NOT1 (N7887, N7883);
nor NOR4 (N7888, N7884, N4247, N3841, N15);
nand NAND3 (N7889, N7876, N5326, N3164);
buf BUF1 (N7890, N7888);
not NOT1 (N7891, N7875);
xor XOR2 (N7892, N7890, N4699);
and AND4 (N7893, N7880, N5781, N6119, N2117);
nand NAND4 (N7894, N7893, N2813, N5075, N3759);
xor XOR2 (N7895, N7881, N660);
xor XOR2 (N7896, N7895, N5909);
and AND2 (N7897, N7869, N826);
and AND4 (N7898, N7889, N349, N2936, N3501);
and AND2 (N7899, N7891, N6886);
not NOT1 (N7900, N7877);
buf BUF1 (N7901, N7897);
xor XOR2 (N7902, N7886, N3171);
not NOT1 (N7903, N7901);
xor XOR2 (N7904, N7892, N4915);
not NOT1 (N7905, N7903);
buf BUF1 (N7906, N7905);
not NOT1 (N7907, N7898);
and AND2 (N7908, N7878, N3431);
xor XOR2 (N7909, N7900, N7617);
and AND3 (N7910, N7899, N921, N2858);
nand NAND3 (N7911, N7896, N7687, N7129);
xor XOR2 (N7912, N7910, N6523);
not NOT1 (N7913, N7904);
or OR4 (N7914, N7908, N3101, N6002, N6904);
nor NOR2 (N7915, N7911, N3054);
xor XOR2 (N7916, N7894, N6068);
not NOT1 (N7917, N7912);
nand NAND2 (N7918, N7902, N1798);
not NOT1 (N7919, N7914);
buf BUF1 (N7920, N7918);
nand NAND2 (N7921, N7915, N2848);
and AND3 (N7922, N7913, N3069, N5684);
nand NAND3 (N7923, N7917, N5603, N1162);
nand NAND2 (N7924, N7887, N2810);
not NOT1 (N7925, N7924);
nor NOR2 (N7926, N7920, N7870);
not NOT1 (N7927, N7919);
buf BUF1 (N7928, N7907);
nand NAND3 (N7929, N7925, N3541, N5455);
not NOT1 (N7930, N7906);
nor NOR2 (N7931, N7927, N7692);
xor XOR2 (N7932, N7928, N3341);
xor XOR2 (N7933, N7929, N2436);
xor XOR2 (N7934, N7930, N897);
nand NAND3 (N7935, N7933, N3767, N2132);
or OR2 (N7936, N7923, N3826);
nand NAND3 (N7937, N7926, N4655, N2950);
buf BUF1 (N7938, N7937);
and AND3 (N7939, N7931, N3220, N3470);
nand NAND3 (N7940, N7922, N231, N4757);
buf BUF1 (N7941, N7938);
and AND3 (N7942, N7935, N2160, N5201);
nand NAND2 (N7943, N7942, N6078);
nor NOR2 (N7944, N7943, N47);
xor XOR2 (N7945, N7934, N2742);
xor XOR2 (N7946, N7945, N385);
not NOT1 (N7947, N7939);
and AND4 (N7948, N7944, N879, N7612, N2952);
buf BUF1 (N7949, N7948);
buf BUF1 (N7950, N7940);
or OR2 (N7951, N7936, N2645);
xor XOR2 (N7952, N7916, N3633);
not NOT1 (N7953, N7950);
and AND2 (N7954, N7921, N7504);
nor NOR4 (N7955, N7941, N3506, N3901, N6593);
and AND4 (N7956, N7951, N3111, N6873, N5483);
and AND2 (N7957, N7947, N1698);
not NOT1 (N7958, N7946);
or OR3 (N7959, N7949, N3780, N1820);
or OR2 (N7960, N7956, N7125);
not NOT1 (N7961, N7953);
xor XOR2 (N7962, N7955, N5169);
xor XOR2 (N7963, N7962, N3807);
buf BUF1 (N7964, N7959);
buf BUF1 (N7965, N7961);
and AND4 (N7966, N7952, N4120, N7836, N4354);
or OR2 (N7967, N7964, N2191);
or OR2 (N7968, N7954, N35);
and AND3 (N7969, N7963, N1198, N7456);
or OR3 (N7970, N7967, N7501, N827);
nor NOR4 (N7971, N7958, N2639, N7512, N6584);
or OR4 (N7972, N7960, N5369, N1067, N6618);
xor XOR2 (N7973, N7932, N12);
and AND3 (N7974, N7970, N3471, N6776);
nor NOR4 (N7975, N7965, N1282, N1208, N7763);
and AND2 (N7976, N7975, N2032);
not NOT1 (N7977, N7974);
or OR2 (N7978, N7957, N2651);
and AND4 (N7979, N7969, N5775, N1923, N7004);
nor NOR3 (N7980, N7909, N3193, N3270);
nor NOR4 (N7981, N7968, N5084, N6653, N495);
or OR3 (N7982, N7978, N2755, N1045);
nand NAND4 (N7983, N7981, N3255, N5496, N959);
or OR4 (N7984, N7966, N7946, N6528, N5437);
and AND3 (N7985, N7979, N2874, N7080);
and AND3 (N7986, N7973, N708, N4058);
nor NOR2 (N7987, N7977, N1096);
and AND3 (N7988, N7972, N2290, N696);
not NOT1 (N7989, N7984);
nor NOR2 (N7990, N7988, N370);
and AND4 (N7991, N7982, N965, N1005, N6597);
xor XOR2 (N7992, N7983, N2256);
not NOT1 (N7993, N7976);
xor XOR2 (N7994, N7985, N7192);
not NOT1 (N7995, N7989);
nor NOR4 (N7996, N7980, N2832, N7414, N6400);
nand NAND2 (N7997, N7987, N1056);
or OR3 (N7998, N7991, N6755, N4525);
and AND2 (N7999, N7998, N5252);
buf BUF1 (N8000, N7995);
buf BUF1 (N8001, N7990);
nor NOR3 (N8002, N7997, N7621, N4694);
or OR4 (N8003, N7986, N7412, N7533, N6717);
xor XOR2 (N8004, N7994, N1638);
or OR3 (N8005, N8001, N459, N5774);
or OR3 (N8006, N7996, N1483, N1447);
not NOT1 (N8007, N7993);
xor XOR2 (N8008, N8002, N7972);
nand NAND3 (N8009, N8005, N7328, N4827);
or OR3 (N8010, N8000, N6519, N47);
xor XOR2 (N8011, N8007, N3401);
buf BUF1 (N8012, N8010);
nor NOR3 (N8013, N8008, N2347, N4848);
buf BUF1 (N8014, N7992);
nand NAND4 (N8015, N8004, N1305, N1890, N5029);
not NOT1 (N8016, N8011);
buf BUF1 (N8017, N7999);
not NOT1 (N8018, N8003);
or OR3 (N8019, N8013, N4063, N5470);
not NOT1 (N8020, N8018);
nand NAND4 (N8021, N8016, N6191, N5739, N322);
buf BUF1 (N8022, N8014);
nor NOR2 (N8023, N8006, N4170);
nand NAND4 (N8024, N8019, N6208, N186, N711);
not NOT1 (N8025, N8023);
nor NOR3 (N8026, N8017, N2824, N1219);
or OR4 (N8027, N7971, N1583, N6070, N170);
not NOT1 (N8028, N8025);
xor XOR2 (N8029, N8021, N4882);
or OR3 (N8030, N8022, N5769, N7387);
xor XOR2 (N8031, N8020, N6088);
buf BUF1 (N8032, N8028);
xor XOR2 (N8033, N8027, N4902);
not NOT1 (N8034, N8026);
nand NAND3 (N8035, N8029, N498, N3610);
xor XOR2 (N8036, N8012, N4912);
and AND4 (N8037, N8032, N5803, N3455, N1975);
nor NOR2 (N8038, N8037, N415);
not NOT1 (N8039, N8035);
nor NOR4 (N8040, N8031, N4210, N663, N4428);
or OR2 (N8041, N8030, N5388);
and AND2 (N8042, N8009, N3230);
nand NAND2 (N8043, N8040, N2141);
or OR4 (N8044, N8043, N989, N2866, N5215);
nand NAND4 (N8045, N8015, N2635, N5052, N3975);
xor XOR2 (N8046, N8024, N756);
nand NAND4 (N8047, N8044, N720, N425, N1435);
not NOT1 (N8048, N8033);
nor NOR3 (N8049, N8039, N2728, N5470);
buf BUF1 (N8050, N8047);
nand NAND4 (N8051, N8045, N2161, N857, N3529);
not NOT1 (N8052, N8046);
and AND4 (N8053, N8041, N1595, N2563, N7065);
buf BUF1 (N8054, N8051);
xor XOR2 (N8055, N8049, N3843);
or OR4 (N8056, N8038, N6349, N1177, N7185);
nand NAND4 (N8057, N8042, N5795, N3156, N4290);
and AND3 (N8058, N8056, N2581, N4924);
or OR4 (N8059, N8054, N1386, N1008, N7978);
or OR4 (N8060, N8053, N3333, N3151, N1507);
buf BUF1 (N8061, N8057);
xor XOR2 (N8062, N8058, N2591);
or OR4 (N8063, N8059, N93, N4969, N1661);
nand NAND2 (N8064, N8055, N4330);
nand NAND3 (N8065, N8060, N5763, N4706);
nand NAND2 (N8066, N8052, N4044);
nand NAND4 (N8067, N8061, N4533, N4421, N8029);
nor NOR3 (N8068, N8050, N5262, N4065);
xor XOR2 (N8069, N8062, N1451);
nand NAND2 (N8070, N8064, N4458);
nor NOR2 (N8071, N8069, N3665);
nand NAND2 (N8072, N8034, N5077);
xor XOR2 (N8073, N8067, N3505);
nand NAND2 (N8074, N8072, N4073);
and AND4 (N8075, N8066, N631, N1252, N1864);
xor XOR2 (N8076, N8036, N7609);
buf BUF1 (N8077, N8048);
not NOT1 (N8078, N8074);
or OR3 (N8079, N8073, N5531, N1229);
nand NAND3 (N8080, N8071, N797, N7504);
buf BUF1 (N8081, N8077);
not NOT1 (N8082, N8076);
or OR3 (N8083, N8063, N3837, N1949);
nor NOR4 (N8084, N8068, N3302, N2296, N4294);
nand NAND4 (N8085, N8075, N1107, N1798, N1142);
nand NAND4 (N8086, N8070, N6615, N3542, N5156);
xor XOR2 (N8087, N8086, N5845);
or OR3 (N8088, N8084, N360, N7013);
xor XOR2 (N8089, N8085, N6770);
or OR3 (N8090, N8083, N4832, N4460);
or OR3 (N8091, N8081, N5274, N2631);
xor XOR2 (N8092, N8091, N2488);
and AND4 (N8093, N8089, N6993, N932, N2758);
not NOT1 (N8094, N8090);
nor NOR3 (N8095, N8094, N7244, N2831);
xor XOR2 (N8096, N8093, N5631);
nand NAND4 (N8097, N8088, N4925, N6172, N3255);
buf BUF1 (N8098, N8095);
xor XOR2 (N8099, N8080, N1443);
or OR2 (N8100, N8097, N6797);
buf BUF1 (N8101, N8099);
xor XOR2 (N8102, N8079, N2028);
xor XOR2 (N8103, N8096, N6499);
or OR2 (N8104, N8098, N2586);
buf BUF1 (N8105, N8101);
buf BUF1 (N8106, N8100);
nor NOR3 (N8107, N8065, N2692, N2657);
not NOT1 (N8108, N8103);
nand NAND4 (N8109, N8105, N7787, N7239, N1285);
buf BUF1 (N8110, N8104);
and AND2 (N8111, N8078, N6622);
and AND3 (N8112, N8087, N4349, N1433);
nor NOR2 (N8113, N8112, N2428);
xor XOR2 (N8114, N8092, N7361);
or OR3 (N8115, N8114, N1630, N4066);
xor XOR2 (N8116, N8110, N2451);
nand NAND2 (N8117, N8106, N2316);
nor NOR4 (N8118, N8107, N7579, N1480, N3150);
and AND3 (N8119, N8115, N2364, N4570);
not NOT1 (N8120, N8108);
not NOT1 (N8121, N8109);
buf BUF1 (N8122, N8111);
nand NAND3 (N8123, N8121, N6065, N7680);
nor NOR3 (N8124, N8082, N664, N7342);
nor NOR4 (N8125, N8117, N4291, N7945, N5177);
nor NOR4 (N8126, N8124, N5711, N2763, N6064);
nor NOR4 (N8127, N8113, N2476, N7717, N7770);
nand NAND2 (N8128, N8102, N3746);
and AND3 (N8129, N8119, N4006, N4000);
xor XOR2 (N8130, N8126, N1926);
or OR3 (N8131, N8128, N5550, N2874);
nand NAND3 (N8132, N8125, N3676, N5725);
not NOT1 (N8133, N8132);
or OR2 (N8134, N8131, N7492);
and AND2 (N8135, N8116, N2398);
nand NAND4 (N8136, N8127, N2670, N4613, N5531);
and AND2 (N8137, N8136, N3052);
and AND3 (N8138, N8122, N7331, N4718);
nand NAND3 (N8139, N8134, N7906, N7196);
nand NAND4 (N8140, N8129, N4374, N5643, N8079);
buf BUF1 (N8141, N8123);
buf BUF1 (N8142, N8141);
nor NOR4 (N8143, N8118, N2345, N5368, N7808);
buf BUF1 (N8144, N8142);
nor NOR3 (N8145, N8137, N4571, N578);
or OR4 (N8146, N8144, N1857, N4618, N8069);
nand NAND3 (N8147, N8130, N532, N1320);
nand NAND3 (N8148, N8133, N1748, N7086);
xor XOR2 (N8149, N8145, N5239);
nor NOR3 (N8150, N8147, N1955, N7296);
and AND3 (N8151, N8140, N7916, N4165);
nor NOR4 (N8152, N8150, N4117, N6383, N5326);
xor XOR2 (N8153, N8143, N1617);
and AND3 (N8154, N8135, N7032, N733);
nor NOR3 (N8155, N8120, N6581, N7794);
xor XOR2 (N8156, N8149, N1471);
or OR2 (N8157, N8153, N2280);
nand NAND3 (N8158, N8139, N6187, N2148);
nand NAND4 (N8159, N8152, N5994, N3209, N506);
nand NAND3 (N8160, N8148, N1108, N1558);
xor XOR2 (N8161, N8151, N7799);
nand NAND3 (N8162, N8157, N107, N2067);
or OR2 (N8163, N8155, N6181);
not NOT1 (N8164, N8146);
or OR4 (N8165, N8164, N2443, N1843, N1344);
xor XOR2 (N8166, N8165, N4569);
nand NAND3 (N8167, N8162, N6906, N5258);
buf BUF1 (N8168, N8159);
nand NAND3 (N8169, N8138, N2183, N2568);
nor NOR2 (N8170, N8161, N2702);
and AND4 (N8171, N8163, N567, N3222, N4075);
or OR3 (N8172, N8160, N3249, N2291);
xor XOR2 (N8173, N8172, N4437);
xor XOR2 (N8174, N8158, N7397);
xor XOR2 (N8175, N8169, N1866);
not NOT1 (N8176, N8154);
nand NAND2 (N8177, N8166, N3604);
xor XOR2 (N8178, N8168, N3085);
xor XOR2 (N8179, N8170, N7163);
buf BUF1 (N8180, N8175);
nor NOR3 (N8181, N8171, N8019, N4266);
or OR3 (N8182, N8179, N5660, N1010);
and AND2 (N8183, N8178, N5622);
xor XOR2 (N8184, N8183, N2173);
buf BUF1 (N8185, N8173);
or OR2 (N8186, N8182, N6875);
nand NAND2 (N8187, N8184, N1767);
nor NOR3 (N8188, N8167, N4868, N5273);
buf BUF1 (N8189, N8174);
or OR2 (N8190, N8186, N6293);
nor NOR3 (N8191, N8185, N1518, N5729);
buf BUF1 (N8192, N8191);
xor XOR2 (N8193, N8180, N1234);
nand NAND4 (N8194, N8189, N7307, N6085, N5371);
nand NAND4 (N8195, N8176, N1448, N7402, N3074);
and AND4 (N8196, N8187, N1060, N8047, N1718);
or OR3 (N8197, N8193, N2951, N8028);
nand NAND2 (N8198, N8188, N1243);
not NOT1 (N8199, N8197);
nor NOR2 (N8200, N8192, N3483);
xor XOR2 (N8201, N8195, N5270);
or OR4 (N8202, N8194, N3670, N1517, N9);
xor XOR2 (N8203, N8181, N7509);
xor XOR2 (N8204, N8202, N3098);
not NOT1 (N8205, N8203);
and AND2 (N8206, N8200, N1782);
or OR3 (N8207, N8199, N4122, N352);
not NOT1 (N8208, N8196);
and AND3 (N8209, N8190, N5306, N5742);
and AND2 (N8210, N8198, N6137);
buf BUF1 (N8211, N8210);
and AND2 (N8212, N8177, N2694);
and AND2 (N8213, N8156, N8161);
or OR3 (N8214, N8205, N6532, N3464);
xor XOR2 (N8215, N8211, N6029);
nor NOR3 (N8216, N8206, N5947, N4171);
nand NAND3 (N8217, N8201, N4112, N6679);
nor NOR3 (N8218, N8209, N1236, N6969);
xor XOR2 (N8219, N8217, N3391);
buf BUF1 (N8220, N8215);
buf BUF1 (N8221, N8218);
nor NOR4 (N8222, N8219, N6745, N3201, N2648);
xor XOR2 (N8223, N8220, N1414);
not NOT1 (N8224, N8207);
buf BUF1 (N8225, N8223);
not NOT1 (N8226, N8214);
xor XOR2 (N8227, N8225, N6311);
nand NAND3 (N8228, N8222, N1882, N7518);
buf BUF1 (N8229, N8227);
not NOT1 (N8230, N8208);
nor NOR4 (N8231, N8216, N1833, N4631, N2503);
buf BUF1 (N8232, N8221);
not NOT1 (N8233, N8228);
xor XOR2 (N8234, N8230, N5879);
nand NAND4 (N8235, N8226, N2899, N7689, N305);
nor NOR2 (N8236, N8212, N6816);
or OR2 (N8237, N8235, N5352);
and AND3 (N8238, N8224, N4954, N5263);
buf BUF1 (N8239, N8232);
xor XOR2 (N8240, N8213, N5376);
xor XOR2 (N8241, N8240, N2091);
nor NOR2 (N8242, N8239, N3464);
buf BUF1 (N8243, N8237);
buf BUF1 (N8244, N8233);
xor XOR2 (N8245, N8238, N2209);
nand NAND4 (N8246, N8231, N6657, N4082, N3500);
not NOT1 (N8247, N8236);
not NOT1 (N8248, N8204);
nor NOR4 (N8249, N8245, N583, N3438, N3016);
xor XOR2 (N8250, N8234, N1707);
and AND2 (N8251, N8248, N6168);
or OR4 (N8252, N8244, N7271, N8227, N1674);
xor XOR2 (N8253, N8229, N3722);
xor XOR2 (N8254, N8253, N3317);
buf BUF1 (N8255, N8242);
nand NAND4 (N8256, N8255, N3361, N2696, N7694);
or OR2 (N8257, N8254, N3984);
nor NOR4 (N8258, N8257, N6960, N2359, N2521);
or OR3 (N8259, N8258, N754, N1076);
nand NAND3 (N8260, N8241, N914, N4881);
or OR4 (N8261, N8251, N7229, N1250, N6263);
and AND3 (N8262, N8261, N6955, N1385);
not NOT1 (N8263, N8247);
or OR2 (N8264, N8246, N4959);
nor NOR4 (N8265, N8256, N3813, N2552, N5722);
and AND3 (N8266, N8264, N5927, N6425);
buf BUF1 (N8267, N8259);
buf BUF1 (N8268, N8252);
and AND3 (N8269, N8263, N379, N6216);
and AND4 (N8270, N8269, N3066, N4172, N6257);
and AND2 (N8271, N8262, N2903);
and AND3 (N8272, N8249, N3349, N3218);
or OR2 (N8273, N8270, N6697);
or OR3 (N8274, N8268, N7604, N404);
nor NOR2 (N8275, N8271, N7064);
or OR2 (N8276, N8273, N2087);
nand NAND2 (N8277, N8260, N5567);
nor NOR3 (N8278, N8277, N7527, N5263);
xor XOR2 (N8279, N8276, N958);
not NOT1 (N8280, N8243);
nor NOR3 (N8281, N8272, N1902, N6909);
nor NOR3 (N8282, N8265, N7924, N6027);
nor NOR4 (N8283, N8266, N3085, N179, N487);
not NOT1 (N8284, N8279);
and AND4 (N8285, N8283, N6320, N7808, N4473);
nor NOR3 (N8286, N8285, N1324, N6015);
and AND2 (N8287, N8284, N3067);
buf BUF1 (N8288, N8287);
not NOT1 (N8289, N8274);
buf BUF1 (N8290, N8288);
not NOT1 (N8291, N8289);
or OR3 (N8292, N8282, N7511, N6887);
or OR3 (N8293, N8278, N6594, N1731);
and AND2 (N8294, N8290, N1093);
nor NOR3 (N8295, N8281, N8025, N6812);
nor NOR4 (N8296, N8286, N5630, N3677, N4695);
not NOT1 (N8297, N8275);
not NOT1 (N8298, N8297);
and AND3 (N8299, N8293, N4849, N3485);
nand NAND2 (N8300, N8250, N5599);
and AND4 (N8301, N8280, N317, N1208, N6531);
and AND4 (N8302, N8267, N764, N6047, N2327);
and AND3 (N8303, N8298, N177, N4118);
or OR2 (N8304, N8294, N6763);
nor NOR4 (N8305, N8304, N5299, N222, N3951);
buf BUF1 (N8306, N8291);
nand NAND4 (N8307, N8292, N4265, N3537, N7371);
nand NAND3 (N8308, N8306, N5786, N5755);
and AND4 (N8309, N8301, N7258, N1517, N953);
or OR3 (N8310, N8302, N2083, N6591);
and AND3 (N8311, N8300, N6032, N4273);
or OR4 (N8312, N8311, N4365, N464, N2563);
xor XOR2 (N8313, N8307, N2491);
nand NAND3 (N8314, N8308, N5386, N2179);
not NOT1 (N8315, N8313);
or OR3 (N8316, N8296, N5116, N7707);
nor NOR3 (N8317, N8315, N1112, N3731);
nand NAND2 (N8318, N8295, N1280);
and AND2 (N8319, N8312, N6845);
buf BUF1 (N8320, N8317);
and AND4 (N8321, N8303, N7588, N5348, N5729);
or OR3 (N8322, N8305, N4414, N5930);
nor NOR3 (N8323, N8299, N2608, N98);
nor NOR2 (N8324, N8321, N3142);
and AND4 (N8325, N8318, N3770, N6155, N2896);
buf BUF1 (N8326, N8325);
and AND2 (N8327, N8322, N675);
and AND3 (N8328, N8316, N1874, N3818);
nand NAND3 (N8329, N8327, N3635, N6028);
nor NOR4 (N8330, N8326, N4724, N180, N7004);
buf BUF1 (N8331, N8330);
and AND3 (N8332, N8320, N177, N7320);
buf BUF1 (N8333, N8319);
nor NOR2 (N8334, N8310, N8297);
nor NOR4 (N8335, N8314, N423, N2399, N4188);
or OR3 (N8336, N8323, N371, N4477);
not NOT1 (N8337, N8309);
not NOT1 (N8338, N8332);
xor XOR2 (N8339, N8329, N4159);
and AND4 (N8340, N8338, N2465, N281, N3291);
not NOT1 (N8341, N8334);
and AND3 (N8342, N8340, N1506, N3356);
nor NOR3 (N8343, N8341, N2277, N621);
or OR2 (N8344, N8336, N7339);
nor NOR2 (N8345, N8337, N5719);
nor NOR2 (N8346, N8324, N3639);
xor XOR2 (N8347, N8346, N5648);
and AND2 (N8348, N8335, N5799);
nand NAND2 (N8349, N8333, N4958);
not NOT1 (N8350, N8343);
xor XOR2 (N8351, N8347, N4654);
nand NAND2 (N8352, N8339, N3656);
xor XOR2 (N8353, N8349, N2297);
and AND3 (N8354, N8342, N2241, N6844);
not NOT1 (N8355, N8352);
or OR3 (N8356, N8348, N3484, N3849);
not NOT1 (N8357, N8350);
and AND3 (N8358, N8331, N3415, N5591);
and AND2 (N8359, N8358, N7826);
buf BUF1 (N8360, N8351);
buf BUF1 (N8361, N8357);
xor XOR2 (N8362, N8360, N2802);
nor NOR3 (N8363, N8353, N1304, N2641);
buf BUF1 (N8364, N8355);
xor XOR2 (N8365, N8344, N7249);
nor NOR3 (N8366, N8354, N4544, N4435);
xor XOR2 (N8367, N8366, N6888);
nand NAND4 (N8368, N8362, N2444, N3262, N6322);
nand NAND4 (N8369, N8356, N4548, N5232, N5824);
nor NOR2 (N8370, N8367, N29);
nand NAND3 (N8371, N8369, N2409, N5014);
and AND3 (N8372, N8359, N6250, N4462);
or OR2 (N8373, N8361, N2475);
buf BUF1 (N8374, N8345);
and AND3 (N8375, N8371, N7304, N6377);
or OR2 (N8376, N8364, N3784);
or OR3 (N8377, N8372, N2020, N6743);
nand NAND2 (N8378, N8370, N18);
buf BUF1 (N8379, N8363);
buf BUF1 (N8380, N8373);
not NOT1 (N8381, N8380);
and AND3 (N8382, N8365, N7306, N1806);
buf BUF1 (N8383, N8381);
or OR4 (N8384, N8382, N1926, N628, N1734);
buf BUF1 (N8385, N8378);
nand NAND4 (N8386, N8328, N2356, N4858, N354);
not NOT1 (N8387, N8386);
or OR4 (N8388, N8385, N6595, N7381, N136);
and AND2 (N8389, N8388, N5401);
and AND2 (N8390, N8376, N5104);
or OR4 (N8391, N8390, N7565, N7037, N3556);
not NOT1 (N8392, N8368);
or OR2 (N8393, N8379, N771);
not NOT1 (N8394, N8389);
and AND2 (N8395, N8383, N2496);
and AND3 (N8396, N8387, N1469, N8000);
xor XOR2 (N8397, N8377, N4339);
xor XOR2 (N8398, N8375, N608);
nand NAND3 (N8399, N8397, N947, N6122);
nor NOR4 (N8400, N8392, N7335, N8316, N3749);
nand NAND2 (N8401, N8394, N7532);
not NOT1 (N8402, N8391);
nor NOR2 (N8403, N8393, N5088);
not NOT1 (N8404, N8399);
or OR2 (N8405, N8401, N4866);
nor NOR2 (N8406, N8400, N580);
or OR3 (N8407, N8406, N7425, N4852);
xor XOR2 (N8408, N8403, N5789);
xor XOR2 (N8409, N8374, N1436);
nand NAND3 (N8410, N8395, N2625, N1676);
nand NAND3 (N8411, N8384, N1896, N2347);
or OR4 (N8412, N8405, N7070, N399, N238);
or OR2 (N8413, N8398, N3046);
nor NOR3 (N8414, N8413, N7086, N4841);
buf BUF1 (N8415, N8410);
not NOT1 (N8416, N8396);
xor XOR2 (N8417, N8411, N5323);
xor XOR2 (N8418, N8412, N1297);
nor NOR4 (N8419, N8409, N1993, N3362, N5857);
or OR4 (N8420, N8402, N8172, N463, N4182);
nor NOR4 (N8421, N8408, N3190, N2123, N958);
or OR4 (N8422, N8415, N8167, N3106, N7340);
buf BUF1 (N8423, N8417);
nand NAND2 (N8424, N8419, N6636);
buf BUF1 (N8425, N8416);
xor XOR2 (N8426, N8421, N2746);
nand NAND2 (N8427, N8422, N8292);
and AND2 (N8428, N8404, N6825);
and AND2 (N8429, N8428, N7025);
nand NAND4 (N8430, N8429, N790, N7817, N207);
nor NOR2 (N8431, N8427, N3258);
or OR3 (N8432, N8414, N2427, N1368);
nand NAND4 (N8433, N8418, N803, N2910, N5593);
buf BUF1 (N8434, N8424);
and AND3 (N8435, N8433, N1505, N7539);
or OR2 (N8436, N8435, N6519);
not NOT1 (N8437, N8420);
nor NOR4 (N8438, N8423, N3430, N6252, N2388);
buf BUF1 (N8439, N8434);
buf BUF1 (N8440, N8407);
xor XOR2 (N8441, N8432, N7917);
nand NAND2 (N8442, N8438, N7428);
and AND4 (N8443, N8440, N7589, N8036, N7244);
nand NAND2 (N8444, N8430, N4304);
not NOT1 (N8445, N8442);
nor NOR3 (N8446, N8445, N5068, N6182);
not NOT1 (N8447, N8446);
nor NOR3 (N8448, N8431, N7702, N5274);
not NOT1 (N8449, N8439);
or OR3 (N8450, N8449, N5562, N1720);
or OR4 (N8451, N8447, N1750, N6513, N7842);
xor XOR2 (N8452, N8436, N6106);
buf BUF1 (N8453, N8441);
or OR3 (N8454, N8452, N6270, N6792);
nand NAND3 (N8455, N8443, N2291, N7488);
and AND4 (N8456, N8425, N6542, N6103, N7705);
and AND2 (N8457, N8453, N3926);
nand NAND2 (N8458, N8450, N2253);
xor XOR2 (N8459, N8456, N993);
not NOT1 (N8460, N8458);
nor NOR2 (N8461, N8444, N3645);
xor XOR2 (N8462, N8455, N1882);
nand NAND2 (N8463, N8462, N1570);
nand NAND4 (N8464, N8426, N2116, N5367, N3587);
xor XOR2 (N8465, N8463, N7513);
nand NAND2 (N8466, N8465, N6827);
xor XOR2 (N8467, N8461, N7250);
or OR2 (N8468, N8451, N2840);
not NOT1 (N8469, N8437);
or OR3 (N8470, N8448, N7365, N2513);
or OR4 (N8471, N8460, N7290, N2320, N1468);
nor NOR4 (N8472, N8466, N5230, N817, N2559);
xor XOR2 (N8473, N8469, N2104);
and AND3 (N8474, N8457, N5746, N1953);
and AND3 (N8475, N8472, N670, N3838);
buf BUF1 (N8476, N8475);
or OR4 (N8477, N8473, N5246, N7774, N2479);
and AND3 (N8478, N8471, N7147, N8279);
nand NAND4 (N8479, N8468, N5888, N5522, N7322);
nand NAND2 (N8480, N8478, N8229);
nor NOR4 (N8481, N8467, N2205, N3866, N5369);
buf BUF1 (N8482, N8454);
or OR3 (N8483, N8474, N7386, N1906);
or OR4 (N8484, N8470, N2119, N2690, N3757);
not NOT1 (N8485, N8476);
and AND4 (N8486, N8459, N7082, N5919, N5611);
or OR4 (N8487, N8480, N2279, N1186, N1725);
buf BUF1 (N8488, N8481);
nand NAND4 (N8489, N8479, N519, N478, N3134);
xor XOR2 (N8490, N8488, N8464);
nand NAND3 (N8491, N3815, N5429, N6715);
or OR4 (N8492, N8489, N8026, N7285, N3282);
nor NOR3 (N8493, N8477, N1165, N2910);
nand NAND3 (N8494, N8485, N2402, N2666);
buf BUF1 (N8495, N8487);
nand NAND4 (N8496, N8493, N2125, N113, N73);
buf BUF1 (N8497, N8496);
nand NAND3 (N8498, N8490, N5060, N6658);
or OR3 (N8499, N8482, N4706, N1173);
or OR4 (N8500, N8486, N3211, N6182, N7526);
not NOT1 (N8501, N8499);
xor XOR2 (N8502, N8501, N1693);
and AND2 (N8503, N8497, N3377);
buf BUF1 (N8504, N8502);
not NOT1 (N8505, N8483);
buf BUF1 (N8506, N8492);
nand NAND4 (N8507, N8498, N4530, N3606, N4333);
buf BUF1 (N8508, N8495);
nand NAND2 (N8509, N8507, N7224);
nand NAND4 (N8510, N8505, N903, N4724, N4195);
nor NOR3 (N8511, N8510, N5071, N1202);
not NOT1 (N8512, N8504);
nor NOR3 (N8513, N8491, N7175, N539);
nand NAND2 (N8514, N8503, N477);
or OR4 (N8515, N8513, N3303, N1905, N5258);
not NOT1 (N8516, N8506);
xor XOR2 (N8517, N8484, N2744);
not NOT1 (N8518, N8500);
and AND3 (N8519, N8515, N8118, N5272);
or OR3 (N8520, N8519, N5550, N1771);
and AND3 (N8521, N8508, N1837, N2034);
not NOT1 (N8522, N8514);
not NOT1 (N8523, N8516);
not NOT1 (N8524, N8522);
not NOT1 (N8525, N8524);
nand NAND2 (N8526, N8517, N3918);
and AND2 (N8527, N8525, N2970);
buf BUF1 (N8528, N8521);
not NOT1 (N8529, N8528);
or OR2 (N8530, N8526, N2160);
nor NOR2 (N8531, N8523, N5245);
nor NOR3 (N8532, N8529, N2737, N687);
buf BUF1 (N8533, N8518);
not NOT1 (N8534, N8532);
not NOT1 (N8535, N8531);
buf BUF1 (N8536, N8509);
not NOT1 (N8537, N8535);
or OR4 (N8538, N8494, N8491, N774, N5254);
not NOT1 (N8539, N8533);
xor XOR2 (N8540, N8538, N2335);
nand NAND3 (N8541, N8536, N4972, N6133);
not NOT1 (N8542, N8541);
or OR3 (N8543, N8530, N3598, N331);
buf BUF1 (N8544, N8542);
nor NOR2 (N8545, N8537, N189);
xor XOR2 (N8546, N8527, N7336);
or OR2 (N8547, N8540, N5698);
or OR2 (N8548, N8511, N5561);
nor NOR3 (N8549, N8548, N5055, N3374);
or OR4 (N8550, N8545, N417, N1222, N7889);
not NOT1 (N8551, N8512);
and AND4 (N8552, N8550, N1168, N8510, N7366);
buf BUF1 (N8553, N8546);
buf BUF1 (N8554, N8543);
or OR4 (N8555, N8539, N4034, N7571, N4698);
or OR3 (N8556, N8534, N5776, N8396);
nor NOR4 (N8557, N8520, N6874, N4879, N2941);
xor XOR2 (N8558, N8551, N604);
buf BUF1 (N8559, N8544);
and AND3 (N8560, N8555, N2405, N6367);
buf BUF1 (N8561, N8558);
nand NAND3 (N8562, N8560, N4667, N5519);
not NOT1 (N8563, N8562);
and AND2 (N8564, N8556, N4594);
nand NAND2 (N8565, N8554, N8225);
and AND3 (N8566, N8565, N2004, N6156);
nor NOR2 (N8567, N8559, N3041);
or OR4 (N8568, N8547, N71, N2772, N8155);
not NOT1 (N8569, N8549);
buf BUF1 (N8570, N8557);
buf BUF1 (N8571, N8553);
not NOT1 (N8572, N8570);
and AND4 (N8573, N8563, N3678, N4216, N8194);
not NOT1 (N8574, N8572);
buf BUF1 (N8575, N8573);
and AND4 (N8576, N8552, N2220, N7712, N460);
nand NAND3 (N8577, N8566, N3303, N3756);
nor NOR3 (N8578, N8574, N5754, N5105);
and AND3 (N8579, N8569, N8311, N1194);
or OR4 (N8580, N8571, N6025, N2763, N3895);
nand NAND4 (N8581, N8577, N3105, N5634, N6688);
xor XOR2 (N8582, N8580, N4581);
buf BUF1 (N8583, N8575);
and AND3 (N8584, N8578, N2081, N8118);
not NOT1 (N8585, N8583);
nand NAND3 (N8586, N8585, N2967, N1324);
buf BUF1 (N8587, N8586);
buf BUF1 (N8588, N8582);
buf BUF1 (N8589, N8579);
xor XOR2 (N8590, N8581, N3976);
nand NAND4 (N8591, N8576, N8530, N8245, N4882);
and AND3 (N8592, N8590, N5750, N6415);
xor XOR2 (N8593, N8561, N1176);
and AND3 (N8594, N8568, N6734, N208);
nor NOR3 (N8595, N8567, N221, N442);
not NOT1 (N8596, N8588);
xor XOR2 (N8597, N8593, N3215);
and AND4 (N8598, N8594, N3984, N1271, N3942);
buf BUF1 (N8599, N8589);
or OR4 (N8600, N8595, N482, N6630, N4132);
xor XOR2 (N8601, N8584, N564);
or OR2 (N8602, N8599, N4088);
nor NOR3 (N8603, N8602, N8288, N4867);
xor XOR2 (N8604, N8597, N6863);
xor XOR2 (N8605, N8601, N1296);
and AND3 (N8606, N8591, N4461, N1876);
nor NOR2 (N8607, N8592, N3498);
or OR2 (N8608, N8606, N3912);
not NOT1 (N8609, N8598);
not NOT1 (N8610, N8564);
nor NOR4 (N8611, N8596, N7141, N6032, N5582);
buf BUF1 (N8612, N8603);
nand NAND4 (N8613, N8612, N4675, N6229, N7954);
nor NOR2 (N8614, N8611, N4579);
buf BUF1 (N8615, N8604);
nand NAND4 (N8616, N8587, N3050, N3193, N2445);
nand NAND4 (N8617, N8608, N2291, N116, N5423);
nor NOR4 (N8618, N8607, N6649, N5036, N6800);
nand NAND2 (N8619, N8609, N6713);
nand NAND4 (N8620, N8613, N8034, N1895, N5381);
or OR2 (N8621, N8617, N8598);
or OR4 (N8622, N8621, N7268, N3936, N5965);
nand NAND4 (N8623, N8622, N4839, N445, N4103);
and AND4 (N8624, N8615, N2135, N7789, N604);
nand NAND3 (N8625, N8619, N5788, N5781);
and AND2 (N8626, N8623, N8259);
or OR4 (N8627, N8625, N7660, N7351, N8089);
nor NOR3 (N8628, N8624, N7390, N5689);
buf BUF1 (N8629, N8614);
nand NAND4 (N8630, N8616, N1612, N3367, N7073);
nand NAND4 (N8631, N8618, N5832, N3808, N3136);
xor XOR2 (N8632, N8620, N2059);
nand NAND4 (N8633, N8631, N48, N4318, N4902);
and AND2 (N8634, N8610, N778);
or OR4 (N8635, N8629, N3246, N7314, N612);
not NOT1 (N8636, N8632);
buf BUF1 (N8637, N8600);
nor NOR3 (N8638, N8635, N686, N6394);
or OR4 (N8639, N8630, N4540, N1011, N1051);
and AND3 (N8640, N8605, N6464, N6147);
and AND2 (N8641, N8627, N3556);
buf BUF1 (N8642, N8628);
nor NOR2 (N8643, N8633, N4703);
nand NAND2 (N8644, N8626, N3681);
and AND2 (N8645, N8641, N5971);
and AND2 (N8646, N8636, N98);
xor XOR2 (N8647, N8640, N7117);
and AND4 (N8648, N8642, N1370, N5640, N6782);
or OR4 (N8649, N8648, N5240, N4511, N1260);
not NOT1 (N8650, N8638);
or OR2 (N8651, N8643, N7657);
nor NOR3 (N8652, N8637, N8625, N5081);
and AND4 (N8653, N8652, N5020, N2763, N54);
nand NAND4 (N8654, N8647, N4214, N3756, N7140);
not NOT1 (N8655, N8651);
not NOT1 (N8656, N8655);
nand NAND4 (N8657, N8634, N1404, N3312, N1295);
xor XOR2 (N8658, N8654, N1897);
and AND4 (N8659, N8650, N3704, N3954, N3987);
xor XOR2 (N8660, N8659, N5174);
nand NAND4 (N8661, N8649, N1371, N3282, N6410);
xor XOR2 (N8662, N8644, N7726);
buf BUF1 (N8663, N8646);
or OR4 (N8664, N8656, N2834, N5148, N175);
and AND3 (N8665, N8653, N5964, N2844);
or OR2 (N8666, N8657, N3491);
and AND4 (N8667, N8665, N2778, N1515, N7001);
nand NAND4 (N8668, N8666, N6406, N287, N4267);
xor XOR2 (N8669, N8662, N4057);
nor NOR3 (N8670, N8639, N4170, N6394);
and AND2 (N8671, N8667, N831);
or OR2 (N8672, N8658, N1562);
or OR2 (N8673, N8672, N2404);
not NOT1 (N8674, N8664);
xor XOR2 (N8675, N8674, N7692);
nand NAND2 (N8676, N8668, N2876);
and AND3 (N8677, N8669, N199, N5966);
and AND2 (N8678, N8676, N5800);
nor NOR2 (N8679, N8663, N594);
nor NOR2 (N8680, N8677, N7027);
or OR3 (N8681, N8661, N4015, N4403);
not NOT1 (N8682, N8673);
nand NAND4 (N8683, N8682, N215, N1965, N3663);
or OR2 (N8684, N8645, N3626);
xor XOR2 (N8685, N8680, N3286);
nor NOR2 (N8686, N8671, N4670);
or OR3 (N8687, N8675, N539, N226);
and AND2 (N8688, N8687, N513);
not NOT1 (N8689, N8679);
buf BUF1 (N8690, N8660);
xor XOR2 (N8691, N8683, N757);
and AND3 (N8692, N8689, N5809, N6166);
and AND3 (N8693, N8670, N7892, N95);
nand NAND3 (N8694, N8688, N6180, N5648);
not NOT1 (N8695, N8684);
and AND3 (N8696, N8678, N6244, N4650);
and AND4 (N8697, N8686, N8473, N1223, N1815);
not NOT1 (N8698, N8693);
buf BUF1 (N8699, N8690);
nand NAND4 (N8700, N8696, N1306, N2038, N2401);
nor NOR4 (N8701, N8699, N7166, N837, N7239);
buf BUF1 (N8702, N8698);
buf BUF1 (N8703, N8697);
nand NAND2 (N8704, N8685, N3615);
nor NOR4 (N8705, N8695, N578, N7578, N3384);
nor NOR4 (N8706, N8692, N181, N1962, N5876);
xor XOR2 (N8707, N8703, N7399);
nor NOR3 (N8708, N8705, N6518, N3993);
xor XOR2 (N8709, N8702, N6425);
and AND4 (N8710, N8694, N7277, N2502, N198);
nand NAND3 (N8711, N8710, N7822, N7247);
or OR4 (N8712, N8709, N343, N4987, N890);
and AND3 (N8713, N8691, N5074, N2980);
or OR4 (N8714, N8681, N7040, N2281, N864);
not NOT1 (N8715, N8707);
not NOT1 (N8716, N8711);
or OR2 (N8717, N8701, N7422);
and AND2 (N8718, N8714, N3461);
not NOT1 (N8719, N8706);
and AND4 (N8720, N8700, N5984, N2351, N7914);
nand NAND3 (N8721, N8712, N6735, N318);
not NOT1 (N8722, N8704);
and AND3 (N8723, N8719, N347, N5487);
buf BUF1 (N8724, N8721);
xor XOR2 (N8725, N8718, N6001);
buf BUF1 (N8726, N8723);
buf BUF1 (N8727, N8722);
nand NAND4 (N8728, N8727, N4045, N8461, N2610);
or OR3 (N8729, N8713, N4464, N4908);
xor XOR2 (N8730, N8726, N2192);
buf BUF1 (N8731, N8730);
and AND2 (N8732, N8725, N8301);
xor XOR2 (N8733, N8728, N5733);
and AND2 (N8734, N8717, N3846);
or OR2 (N8735, N8729, N934);
not NOT1 (N8736, N8720);
nand NAND2 (N8737, N8736, N3239);
nor NOR4 (N8738, N8735, N4520, N2925, N1612);
or OR4 (N8739, N8732, N3227, N200, N8419);
xor XOR2 (N8740, N8708, N6219);
or OR2 (N8741, N8731, N5093);
xor XOR2 (N8742, N8739, N2054);
nor NOR4 (N8743, N8715, N7935, N4370, N345);
and AND4 (N8744, N8737, N8729, N7540, N4113);
nor NOR2 (N8745, N8716, N8383);
and AND4 (N8746, N8745, N6745, N2992, N5161);
xor XOR2 (N8747, N8746, N8716);
nand NAND4 (N8748, N8741, N8495, N3375, N4332);
nor NOR2 (N8749, N8734, N6337);
not NOT1 (N8750, N8724);
and AND4 (N8751, N8740, N6440, N3097, N3112);
buf BUF1 (N8752, N8751);
xor XOR2 (N8753, N8738, N993);
nor NOR4 (N8754, N8748, N459, N7871, N4810);
or OR4 (N8755, N8750, N2512, N7002, N1996);
buf BUF1 (N8756, N8753);
xor XOR2 (N8757, N8744, N6239);
and AND4 (N8758, N8747, N8491, N7052, N3142);
nor NOR4 (N8759, N8752, N2939, N6347, N4997);
buf BUF1 (N8760, N8758);
buf BUF1 (N8761, N8760);
not NOT1 (N8762, N8756);
or OR3 (N8763, N8749, N6436, N3564);
nor NOR4 (N8764, N8757, N6827, N4213, N5398);
nor NOR3 (N8765, N8764, N7558, N180);
nor NOR3 (N8766, N8743, N8018, N237);
xor XOR2 (N8767, N8742, N5498);
nor NOR2 (N8768, N8766, N8733);
xor XOR2 (N8769, N4232, N7568);
nor NOR2 (N8770, N8759, N3988);
nand NAND3 (N8771, N8755, N1946, N4066);
not NOT1 (N8772, N8769);
xor XOR2 (N8773, N8762, N3631);
nor NOR3 (N8774, N8763, N8707, N7338);
xor XOR2 (N8775, N8772, N8554);
xor XOR2 (N8776, N8761, N6701);
nor NOR2 (N8777, N8768, N3029);
nand NAND4 (N8778, N8770, N3256, N4276, N6971);
or OR4 (N8779, N8774, N8022, N629, N643);
nor NOR2 (N8780, N8779, N1849);
nand NAND4 (N8781, N8777, N8647, N4953, N1411);
and AND2 (N8782, N8775, N3202);
and AND4 (N8783, N8778, N2315, N2050, N7765);
nor NOR2 (N8784, N8781, N1713);
nand NAND2 (N8785, N8765, N8453);
or OR4 (N8786, N8784, N3298, N1762, N7354);
nand NAND4 (N8787, N8773, N297, N4428, N7436);
or OR4 (N8788, N8783, N3427, N5807, N4008);
and AND4 (N8789, N8782, N3456, N1779, N4417);
or OR2 (N8790, N8776, N3175);
nand NAND4 (N8791, N8789, N6920, N3847, N2378);
nand NAND2 (N8792, N8785, N7002);
buf BUF1 (N8793, N8790);
and AND3 (N8794, N8788, N3881, N6844);
and AND4 (N8795, N8791, N6500, N351, N3710);
not NOT1 (N8796, N8793);
nor NOR2 (N8797, N8780, N7054);
nand NAND2 (N8798, N8796, N3389);
nand NAND2 (N8799, N8797, N8510);
buf BUF1 (N8800, N8787);
nand NAND4 (N8801, N8799, N7437, N4905, N3468);
and AND2 (N8802, N8754, N6998);
and AND3 (N8803, N8794, N7988, N3542);
nor NOR4 (N8804, N8800, N7225, N3826, N1751);
nor NOR4 (N8805, N8801, N8432, N649, N2429);
nor NOR3 (N8806, N8792, N3932, N5917);
or OR2 (N8807, N8771, N2359);
nand NAND4 (N8808, N8786, N6360, N7195, N5022);
nand NAND4 (N8809, N8802, N8501, N1110, N1823);
nor NOR4 (N8810, N8803, N5213, N5474, N4679);
or OR3 (N8811, N8806, N2285, N8035);
buf BUF1 (N8812, N8811);
not NOT1 (N8813, N8810);
nor NOR2 (N8814, N8807, N8657);
nand NAND2 (N8815, N8814, N3454);
nor NOR4 (N8816, N8798, N2572, N7306, N5000);
buf BUF1 (N8817, N8808);
buf BUF1 (N8818, N8809);
not NOT1 (N8819, N8805);
nand NAND2 (N8820, N8812, N3179);
or OR2 (N8821, N8813, N5427);
buf BUF1 (N8822, N8817);
nor NOR3 (N8823, N8820, N8310, N8107);
xor XOR2 (N8824, N8767, N3406);
not NOT1 (N8825, N8821);
or OR2 (N8826, N8815, N5261);
and AND3 (N8827, N8823, N263, N1390);
buf BUF1 (N8828, N8822);
and AND4 (N8829, N8819, N7964, N2865, N2384);
buf BUF1 (N8830, N8829);
not NOT1 (N8831, N8825);
buf BUF1 (N8832, N8818);
or OR4 (N8833, N8795, N1057, N157, N3698);
buf BUF1 (N8834, N8833);
xor XOR2 (N8835, N8832, N7362);
not NOT1 (N8836, N8824);
nand NAND4 (N8837, N8804, N1458, N8106, N4098);
nand NAND3 (N8838, N8828, N7714, N6165);
nor NOR3 (N8839, N8831, N2323, N7467);
and AND3 (N8840, N8826, N8747, N4212);
or OR2 (N8841, N8837, N8236);
xor XOR2 (N8842, N8841, N8493);
not NOT1 (N8843, N8816);
xor XOR2 (N8844, N8836, N6578);
nand NAND3 (N8845, N8827, N2744, N61);
xor XOR2 (N8846, N8834, N3139);
buf BUF1 (N8847, N8839);
or OR3 (N8848, N8840, N8241, N6609);
buf BUF1 (N8849, N8844);
nor NOR3 (N8850, N8846, N5977, N3789);
nor NOR3 (N8851, N8835, N7086, N5742);
and AND3 (N8852, N8847, N3959, N4875);
not NOT1 (N8853, N8848);
nand NAND2 (N8854, N8849, N7998);
not NOT1 (N8855, N8845);
and AND3 (N8856, N8850, N5807, N8643);
or OR2 (N8857, N8855, N5890);
xor XOR2 (N8858, N8830, N8774);
and AND3 (N8859, N8853, N8184, N8689);
xor XOR2 (N8860, N8838, N4229);
not NOT1 (N8861, N8858);
or OR3 (N8862, N8860, N8341, N5452);
nor NOR2 (N8863, N8856, N7948);
nand NAND4 (N8864, N8843, N3436, N5126, N3280);
nand NAND2 (N8865, N8859, N7768);
nor NOR3 (N8866, N8861, N5657, N540);
or OR3 (N8867, N8863, N441, N4344);
nor NOR4 (N8868, N8842, N4519, N7460, N6185);
buf BUF1 (N8869, N8851);
not NOT1 (N8870, N8857);
or OR2 (N8871, N8869, N954);
not NOT1 (N8872, N8854);
nand NAND3 (N8873, N8864, N1920, N7090);
xor XOR2 (N8874, N8873, N8827);
not NOT1 (N8875, N8866);
nand NAND3 (N8876, N8862, N4198, N2484);
not NOT1 (N8877, N8870);
nand NAND3 (N8878, N8875, N4297, N2791);
buf BUF1 (N8879, N8878);
nand NAND3 (N8880, N8852, N794, N8709);
xor XOR2 (N8881, N8868, N2669);
nor NOR3 (N8882, N8879, N2741, N4305);
or OR4 (N8883, N8872, N8004, N2940, N6012);
or OR3 (N8884, N8874, N7178, N3333);
nand NAND2 (N8885, N8880, N3014);
or OR2 (N8886, N8867, N4597);
not NOT1 (N8887, N8881);
nor NOR4 (N8888, N8885, N2082, N6947, N1793);
xor XOR2 (N8889, N8865, N1441);
buf BUF1 (N8890, N8888);
not NOT1 (N8891, N8884);
xor XOR2 (N8892, N8890, N8584);
and AND3 (N8893, N8883, N2345, N1187);
buf BUF1 (N8894, N8887);
xor XOR2 (N8895, N8893, N4668);
nor NOR3 (N8896, N8892, N2985, N7376);
nor NOR2 (N8897, N8889, N5736);
or OR4 (N8898, N8895, N4594, N7474, N8855);
nor NOR4 (N8899, N8876, N4278, N1042, N1961);
buf BUF1 (N8900, N8882);
and AND3 (N8901, N8894, N4348, N4806);
xor XOR2 (N8902, N8901, N6070);
buf BUF1 (N8903, N8900);
buf BUF1 (N8904, N8902);
buf BUF1 (N8905, N8896);
buf BUF1 (N8906, N8905);
xor XOR2 (N8907, N8877, N4639);
or OR4 (N8908, N8897, N2889, N1779, N193);
or OR2 (N8909, N8906, N3480);
nor NOR4 (N8910, N8908, N390, N2274, N8746);
and AND4 (N8911, N8909, N6849, N7940, N7658);
and AND3 (N8912, N8891, N7908, N5530);
buf BUF1 (N8913, N8899);
and AND4 (N8914, N8886, N2057, N1673, N1136);
buf BUF1 (N8915, N8910);
not NOT1 (N8916, N8898);
or OR3 (N8917, N8904, N172, N5033);
nor NOR3 (N8918, N8917, N8464, N8833);
nand NAND3 (N8919, N8913, N3407, N2453);
xor XOR2 (N8920, N8918, N113);
not NOT1 (N8921, N8919);
not NOT1 (N8922, N8914);
and AND2 (N8923, N8922, N8489);
buf BUF1 (N8924, N8916);
xor XOR2 (N8925, N8923, N7949);
nand NAND3 (N8926, N8907, N6130, N6435);
not NOT1 (N8927, N8915);
buf BUF1 (N8928, N8871);
buf BUF1 (N8929, N8912);
nand NAND3 (N8930, N8921, N7603, N7972);
and AND3 (N8931, N8930, N7426, N6118);
and AND4 (N8932, N8920, N1753, N2235, N1527);
nand NAND3 (N8933, N8911, N2994, N2540);
or OR3 (N8934, N8926, N1419, N6360);
not NOT1 (N8935, N8924);
xor XOR2 (N8936, N8931, N7969);
or OR4 (N8937, N8936, N8066, N199, N7125);
buf BUF1 (N8938, N8928);
xor XOR2 (N8939, N8934, N7360);
nand NAND4 (N8940, N8938, N6890, N568, N8819);
not NOT1 (N8941, N8925);
nor NOR4 (N8942, N8903, N4063, N4073, N2435);
nor NOR2 (N8943, N8935, N4118);
not NOT1 (N8944, N8941);
nand NAND2 (N8945, N8942, N6342);
and AND4 (N8946, N8937, N7522, N8315, N4865);
nor NOR3 (N8947, N8927, N5010, N8744);
and AND3 (N8948, N8945, N290, N6007);
nor NOR4 (N8949, N8939, N657, N3192, N270);
nand NAND2 (N8950, N8949, N2353);
xor XOR2 (N8951, N8932, N5596);
nor NOR2 (N8952, N8948, N2266);
nor NOR3 (N8953, N8944, N6592, N2351);
or OR4 (N8954, N8933, N4886, N1754, N1126);
not NOT1 (N8955, N8943);
nor NOR3 (N8956, N8953, N6056, N1779);
not NOT1 (N8957, N8956);
not NOT1 (N8958, N8954);
not NOT1 (N8959, N8952);
nand NAND3 (N8960, N8929, N2921, N1594);
or OR3 (N8961, N8940, N5885, N2959);
xor XOR2 (N8962, N8950, N8352);
nor NOR2 (N8963, N8955, N2617);
or OR2 (N8964, N8946, N5522);
buf BUF1 (N8965, N8963);
nand NAND4 (N8966, N8964, N6880, N8596, N5186);
and AND2 (N8967, N8960, N8213);
and AND4 (N8968, N8959, N4614, N1904, N1592);
nand NAND3 (N8969, N8968, N339, N5831);
nor NOR3 (N8970, N8966, N1945, N8329);
nand NAND4 (N8971, N8962, N5878, N8733, N645);
or OR3 (N8972, N8957, N3250, N2581);
or OR3 (N8973, N8947, N2987, N689);
buf BUF1 (N8974, N8972);
or OR2 (N8975, N8967, N2660);
nand NAND4 (N8976, N8958, N5330, N6717, N2871);
xor XOR2 (N8977, N8975, N4837);
or OR2 (N8978, N8961, N139);
buf BUF1 (N8979, N8977);
nor NOR2 (N8980, N8974, N4467);
buf BUF1 (N8981, N8978);
or OR2 (N8982, N8981, N8613);
and AND4 (N8983, N8982, N5296, N5594, N4885);
nand NAND4 (N8984, N8976, N5170, N3503, N4507);
and AND2 (N8985, N8984, N794);
nand NAND2 (N8986, N8973, N516);
or OR4 (N8987, N8983, N2924, N1202, N989);
and AND4 (N8988, N8986, N2914, N5829, N575);
nand NAND4 (N8989, N8951, N5456, N6065, N855);
nand NAND4 (N8990, N8979, N6037, N8965, N5008);
and AND3 (N8991, N655, N6384, N3059);
xor XOR2 (N8992, N8980, N6270);
buf BUF1 (N8993, N8991);
and AND4 (N8994, N8989, N3335, N1432, N7778);
nor NOR2 (N8995, N8985, N8985);
and AND3 (N8996, N8990, N5345, N4279);
not NOT1 (N8997, N8996);
buf BUF1 (N8998, N8995);
xor XOR2 (N8999, N8988, N3197);
xor XOR2 (N9000, N8969, N1872);
buf BUF1 (N9001, N8970);
and AND3 (N9002, N8971, N127, N3570);
and AND3 (N9003, N8997, N7316, N1595);
or OR2 (N9004, N8999, N7993);
and AND3 (N9005, N8987, N2749, N5712);
and AND2 (N9006, N9004, N3927);
nand NAND3 (N9007, N8992, N3801, N3548);
xor XOR2 (N9008, N9006, N8938);
not NOT1 (N9009, N9000);
and AND3 (N9010, N9001, N5660, N1499);
not NOT1 (N9011, N8994);
nor NOR3 (N9012, N9002, N2897, N7019);
xor XOR2 (N9013, N9003, N2009);
or OR4 (N9014, N9008, N7770, N8311, N5189);
xor XOR2 (N9015, N9014, N6717);
and AND4 (N9016, N9013, N747, N7441, N4500);
nand NAND4 (N9017, N9009, N6491, N6754, N4606);
or OR2 (N9018, N9017, N3434);
not NOT1 (N9019, N9011);
nand NAND3 (N9020, N8993, N8715, N3378);
buf BUF1 (N9021, N9016);
xor XOR2 (N9022, N8998, N5518);
buf BUF1 (N9023, N9020);
buf BUF1 (N9024, N9010);
and AND3 (N9025, N9021, N3625, N4244);
buf BUF1 (N9026, N9019);
buf BUF1 (N9027, N9005);
not NOT1 (N9028, N9023);
buf BUF1 (N9029, N9025);
not NOT1 (N9030, N9027);
nand NAND4 (N9031, N9029, N7691, N1054, N4458);
nand NAND4 (N9032, N9012, N3637, N7124, N3156);
nand NAND4 (N9033, N9032, N3127, N3882, N6660);
or OR3 (N9034, N9030, N1476, N7361);
buf BUF1 (N9035, N9022);
and AND2 (N9036, N9033, N5283);
not NOT1 (N9037, N9018);
and AND4 (N9038, N9036, N8711, N4426, N6655);
not NOT1 (N9039, N9028);
or OR4 (N9040, N9007, N8038, N8031, N1943);
not NOT1 (N9041, N9038);
not NOT1 (N9042, N9031);
not NOT1 (N9043, N9015);
nand NAND3 (N9044, N9040, N8581, N7768);
not NOT1 (N9045, N9037);
or OR2 (N9046, N9043, N8676);
not NOT1 (N9047, N9041);
xor XOR2 (N9048, N9047, N5065);
xor XOR2 (N9049, N9034, N8760);
not NOT1 (N9050, N9024);
nor NOR2 (N9051, N9045, N4308);
nand NAND4 (N9052, N9044, N771, N3412, N3371);
or OR4 (N9053, N9049, N5561, N6479, N5071);
nor NOR2 (N9054, N9051, N8568);
nand NAND4 (N9055, N9035, N503, N6326, N6271);
buf BUF1 (N9056, N9055);
and AND4 (N9057, N9026, N3704, N1952, N4591);
and AND4 (N9058, N9052, N8131, N6096, N1957);
nand NAND4 (N9059, N9046, N1470, N4065, N8402);
not NOT1 (N9060, N9058);
and AND4 (N9061, N9042, N164, N2711, N4663);
nor NOR3 (N9062, N9061, N463, N2136);
not NOT1 (N9063, N9057);
nor NOR3 (N9064, N9039, N3707, N4270);
or OR3 (N9065, N9054, N6744, N2263);
or OR3 (N9066, N9048, N8125, N2918);
and AND4 (N9067, N9063, N8308, N8971, N1351);
nor NOR4 (N9068, N9053, N6329, N971, N562);
nor NOR4 (N9069, N9050, N2208, N6698, N3551);
xor XOR2 (N9070, N9067, N7136);
or OR4 (N9071, N9065, N4227, N2630, N7136);
nand NAND2 (N9072, N9059, N4199);
not NOT1 (N9073, N9066);
nor NOR3 (N9074, N9072, N8717, N2078);
buf BUF1 (N9075, N9062);
or OR4 (N9076, N9070, N8146, N482, N7784);
buf BUF1 (N9077, N9071);
and AND3 (N9078, N9074, N4354, N3295);
xor XOR2 (N9079, N9068, N7367);
and AND4 (N9080, N9076, N3290, N7596, N3498);
or OR2 (N9081, N9060, N2868);
or OR3 (N9082, N9079, N3733, N7063);
not NOT1 (N9083, N9080);
xor XOR2 (N9084, N9078, N422);
xor XOR2 (N9085, N9056, N7571);
and AND3 (N9086, N9081, N6345, N1895);
buf BUF1 (N9087, N9082);
or OR2 (N9088, N9073, N2854);
xor XOR2 (N9089, N9064, N2262);
and AND2 (N9090, N9086, N3896);
nand NAND4 (N9091, N9087, N7470, N5695, N7244);
not NOT1 (N9092, N9084);
not NOT1 (N9093, N9090);
not NOT1 (N9094, N9069);
and AND3 (N9095, N9088, N8933, N5569);
and AND4 (N9096, N9091, N8468, N8422, N6980);
and AND2 (N9097, N9089, N3837);
nor NOR4 (N9098, N9092, N8831, N301, N1755);
nor NOR4 (N9099, N9097, N7133, N8630, N2856);
not NOT1 (N9100, N9094);
nand NAND3 (N9101, N9100, N7590, N6917);
buf BUF1 (N9102, N9093);
buf BUF1 (N9103, N9101);
nor NOR4 (N9104, N9099, N260, N2501, N8218);
xor XOR2 (N9105, N9083, N7679);
nand NAND2 (N9106, N9102, N1330);
nor NOR3 (N9107, N9103, N3510, N2437);
and AND3 (N9108, N9095, N1022, N4555);
buf BUF1 (N9109, N9106);
nand NAND4 (N9110, N9109, N4193, N4221, N8343);
xor XOR2 (N9111, N9085, N8087);
or OR2 (N9112, N9096, N2980);
not NOT1 (N9113, N9108);
nor NOR2 (N9114, N9104, N7827);
nand NAND4 (N9115, N9107, N3052, N4305, N6570);
nand NAND4 (N9116, N9075, N72, N3519, N8504);
buf BUF1 (N9117, N9112);
nor NOR3 (N9118, N9113, N8274, N5865);
and AND3 (N9119, N9077, N1890, N8391);
or OR2 (N9120, N9119, N6549);
nor NOR3 (N9121, N9116, N2227, N7868);
xor XOR2 (N9122, N9110, N8873);
xor XOR2 (N9123, N9118, N8275);
or OR2 (N9124, N9098, N5532);
not NOT1 (N9125, N9121);
buf BUF1 (N9126, N9125);
buf BUF1 (N9127, N9120);
not NOT1 (N9128, N9114);
and AND3 (N9129, N9126, N7865, N7500);
nor NOR4 (N9130, N9124, N6097, N8337, N2646);
and AND4 (N9131, N9128, N8064, N6280, N5333);
xor XOR2 (N9132, N9130, N442);
nor NOR3 (N9133, N9132, N6379, N7132);
or OR4 (N9134, N9122, N4330, N1484, N7714);
not NOT1 (N9135, N9134);
nor NOR3 (N9136, N9127, N1489, N6443);
not NOT1 (N9137, N9117);
and AND3 (N9138, N9115, N7926, N1276);
or OR4 (N9139, N9133, N6598, N7691, N7098);
and AND2 (N9140, N9129, N3332);
nor NOR3 (N9141, N9139, N3915, N3257);
or OR4 (N9142, N9105, N2020, N6705, N6202);
nand NAND3 (N9143, N9137, N1611, N5101);
xor XOR2 (N9144, N9136, N8390);
nor NOR2 (N9145, N9144, N841);
xor XOR2 (N9146, N9138, N6629);
and AND3 (N9147, N9141, N6167, N157);
xor XOR2 (N9148, N9147, N8178);
or OR3 (N9149, N9148, N6136, N3088);
nor NOR3 (N9150, N9123, N9144, N2406);
buf BUF1 (N9151, N9146);
xor XOR2 (N9152, N9143, N5804);
nand NAND2 (N9153, N9150, N4317);
not NOT1 (N9154, N9131);
xor XOR2 (N9155, N9145, N2249);
buf BUF1 (N9156, N9149);
nor NOR2 (N9157, N9152, N6502);
or OR4 (N9158, N9111, N7977, N669, N4641);
not NOT1 (N9159, N9153);
nand NAND4 (N9160, N9151, N7478, N2420, N8959);
xor XOR2 (N9161, N9140, N4686);
and AND3 (N9162, N9157, N6523, N1913);
buf BUF1 (N9163, N9158);
not NOT1 (N9164, N9160);
nand NAND4 (N9165, N9155, N7398, N6960, N6437);
nor NOR2 (N9166, N9154, N2567);
nor NOR3 (N9167, N9164, N4849, N3213);
not NOT1 (N9168, N9167);
xor XOR2 (N9169, N9165, N3589);
nor NOR2 (N9170, N9161, N8117);
nor NOR4 (N9171, N9156, N2329, N6711, N8464);
buf BUF1 (N9172, N9159);
or OR2 (N9173, N9166, N1181);
xor XOR2 (N9174, N9172, N3393);
not NOT1 (N9175, N9174);
buf BUF1 (N9176, N9170);
nand NAND3 (N9177, N9168, N7718, N8643);
xor XOR2 (N9178, N9176, N8605);
and AND3 (N9179, N9163, N6905, N8454);
or OR3 (N9180, N9173, N196, N5602);
nand NAND2 (N9181, N9175, N2280);
nand NAND2 (N9182, N9135, N6057);
buf BUF1 (N9183, N9171);
xor XOR2 (N9184, N9177, N4293);
nor NOR4 (N9185, N9142, N1911, N1667, N2021);
not NOT1 (N9186, N9169);
nand NAND4 (N9187, N9183, N8393, N1587, N2139);
buf BUF1 (N9188, N9186);
nor NOR4 (N9189, N9178, N9071, N3845, N2079);
nand NAND3 (N9190, N9180, N1835, N5471);
or OR2 (N9191, N9190, N133);
nor NOR2 (N9192, N9187, N3108);
nor NOR2 (N9193, N9185, N2887);
nor NOR2 (N9194, N9191, N3594);
nand NAND4 (N9195, N9179, N9139, N8587, N978);
nor NOR3 (N9196, N9189, N3761, N2296);
buf BUF1 (N9197, N9162);
nand NAND3 (N9198, N9193, N1721, N134);
xor XOR2 (N9199, N9184, N2425);
nand NAND4 (N9200, N9198, N7569, N5371, N8934);
nand NAND4 (N9201, N9181, N4277, N7143, N649);
xor XOR2 (N9202, N9201, N1778);
nand NAND4 (N9203, N9197, N3427, N1593, N6401);
not NOT1 (N9204, N9203);
nor NOR3 (N9205, N9199, N7520, N8424);
not NOT1 (N9206, N9205);
nand NAND3 (N9207, N9192, N6692, N623);
not NOT1 (N9208, N9182);
xor XOR2 (N9209, N9200, N3199);
buf BUF1 (N9210, N9206);
buf BUF1 (N9211, N9207);
xor XOR2 (N9212, N9204, N1730);
not NOT1 (N9213, N9211);
buf BUF1 (N9214, N9202);
or OR3 (N9215, N9188, N9085, N810);
buf BUF1 (N9216, N9208);
xor XOR2 (N9217, N9213, N3166);
xor XOR2 (N9218, N9195, N7319);
not NOT1 (N9219, N9212);
not NOT1 (N9220, N9215);
nand NAND2 (N9221, N9209, N605);
or OR2 (N9222, N9196, N1553);
not NOT1 (N9223, N9210);
and AND2 (N9224, N9214, N1841);
xor XOR2 (N9225, N9222, N7787);
buf BUF1 (N9226, N9220);
xor XOR2 (N9227, N9226, N5118);
nor NOR2 (N9228, N9225, N1081);
xor XOR2 (N9229, N9194, N3888);
not NOT1 (N9230, N9217);
and AND2 (N9231, N9223, N4255);
buf BUF1 (N9232, N9229);
buf BUF1 (N9233, N9232);
xor XOR2 (N9234, N9233, N255);
nand NAND4 (N9235, N9228, N7140, N6275, N569);
and AND4 (N9236, N9216, N3559, N4945, N7431);
xor XOR2 (N9237, N9236, N810);
not NOT1 (N9238, N9219);
not NOT1 (N9239, N9238);
nand NAND4 (N9240, N9230, N3164, N7809, N3734);
and AND4 (N9241, N9224, N8596, N5186, N9227);
xor XOR2 (N9242, N5016, N5435);
xor XOR2 (N9243, N9218, N5607);
or OR2 (N9244, N9243, N3561);
nor NOR2 (N9245, N9234, N564);
not NOT1 (N9246, N9221);
nor NOR2 (N9247, N9245, N137);
or OR4 (N9248, N9239, N5164, N1945, N4050);
not NOT1 (N9249, N9246);
nor NOR3 (N9250, N9237, N7551, N2522);
nor NOR2 (N9251, N9247, N8786);
buf BUF1 (N9252, N9235);
nand NAND4 (N9253, N9248, N3705, N5901, N3132);
buf BUF1 (N9254, N9251);
or OR4 (N9255, N9249, N3020, N3523, N5853);
and AND2 (N9256, N9244, N2701);
buf BUF1 (N9257, N9231);
nand NAND4 (N9258, N9241, N2409, N5500, N4211);
and AND4 (N9259, N9258, N20, N3845, N4738);
buf BUF1 (N9260, N9257);
nor NOR3 (N9261, N9252, N6776, N6778);
xor XOR2 (N9262, N9255, N1004);
nand NAND3 (N9263, N9253, N8643, N8737);
and AND4 (N9264, N9254, N1638, N5996, N1500);
not NOT1 (N9265, N9240);
xor XOR2 (N9266, N9260, N8520);
nor NOR3 (N9267, N9242, N1691, N1548);
nand NAND3 (N9268, N9267, N7367, N2005);
nand NAND4 (N9269, N9263, N2754, N8697, N4782);
nand NAND4 (N9270, N9262, N7834, N2507, N4647);
not NOT1 (N9271, N9270);
and AND3 (N9272, N9264, N7063, N9016);
not NOT1 (N9273, N9272);
xor XOR2 (N9274, N9259, N1);
or OR2 (N9275, N9273, N2302);
xor XOR2 (N9276, N9269, N786);
xor XOR2 (N9277, N9266, N2208);
buf BUF1 (N9278, N9268);
and AND4 (N9279, N9278, N3389, N44, N7566);
nand NAND2 (N9280, N9279, N4184);
xor XOR2 (N9281, N9274, N1547);
buf BUF1 (N9282, N9265);
nor NOR2 (N9283, N9256, N9078);
nor NOR4 (N9284, N9261, N849, N3696, N426);
nor NOR2 (N9285, N9271, N4909);
not NOT1 (N9286, N9250);
xor XOR2 (N9287, N9285, N64);
not NOT1 (N9288, N9275);
nand NAND3 (N9289, N9283, N162, N4268);
xor XOR2 (N9290, N9281, N7499);
not NOT1 (N9291, N9277);
xor XOR2 (N9292, N9287, N6310);
buf BUF1 (N9293, N9291);
or OR4 (N9294, N9286, N4333, N2308, N1132);
not NOT1 (N9295, N9292);
xor XOR2 (N9296, N9282, N7766);
nand NAND3 (N9297, N9293, N5593, N4428);
nor NOR3 (N9298, N9289, N6713, N5933);
not NOT1 (N9299, N9294);
not NOT1 (N9300, N9276);
nand NAND2 (N9301, N9297, N768);
or OR3 (N9302, N9298, N5469, N6130);
buf BUF1 (N9303, N9300);
nand NAND2 (N9304, N9288, N1864);
xor XOR2 (N9305, N9290, N2245);
xor XOR2 (N9306, N9280, N7857);
or OR2 (N9307, N9305, N8358);
nand NAND3 (N9308, N9306, N4559, N7259);
xor XOR2 (N9309, N9295, N8750);
and AND4 (N9310, N9303, N7785, N4759, N7759);
nor NOR4 (N9311, N9310, N8588, N8913, N4660);
or OR2 (N9312, N9296, N4673);
not NOT1 (N9313, N9309);
xor XOR2 (N9314, N9311, N5386);
and AND2 (N9315, N9302, N3036);
not NOT1 (N9316, N9307);
and AND2 (N9317, N9299, N4449);
not NOT1 (N9318, N9315);
nor NOR4 (N9319, N9316, N1614, N8684, N427);
nand NAND2 (N9320, N9312, N208);
and AND4 (N9321, N9314, N2706, N394, N2486);
buf BUF1 (N9322, N9304);
buf BUF1 (N9323, N9317);
nor NOR3 (N9324, N9308, N2057, N4216);
xor XOR2 (N9325, N9318, N2863);
xor XOR2 (N9326, N9319, N3053);
buf BUF1 (N9327, N9322);
not NOT1 (N9328, N9321);
xor XOR2 (N9329, N9301, N6540);
nand NAND4 (N9330, N9320, N3660, N8305, N346);
buf BUF1 (N9331, N9325);
xor XOR2 (N9332, N9326, N8558);
buf BUF1 (N9333, N9328);
or OR2 (N9334, N9327, N9240);
buf BUF1 (N9335, N9331);
nor NOR2 (N9336, N9324, N8098);
or OR3 (N9337, N9334, N9265, N1577);
xor XOR2 (N9338, N9336, N6815);
nand NAND3 (N9339, N9329, N7413, N6425);
not NOT1 (N9340, N9313);
xor XOR2 (N9341, N9340, N6162);
not NOT1 (N9342, N9339);
buf BUF1 (N9343, N9337);
and AND2 (N9344, N9335, N8404);
not NOT1 (N9345, N9333);
nand NAND2 (N9346, N9343, N8477);
buf BUF1 (N9347, N9323);
buf BUF1 (N9348, N9347);
xor XOR2 (N9349, N9284, N6752);
buf BUF1 (N9350, N9332);
not NOT1 (N9351, N9345);
xor XOR2 (N9352, N9348, N4435);
buf BUF1 (N9353, N9344);
nand NAND4 (N9354, N9338, N4207, N4587, N1426);
or OR3 (N9355, N9342, N2751, N5504);
buf BUF1 (N9356, N9353);
or OR2 (N9357, N9330, N2206);
nor NOR4 (N9358, N9354, N4602, N3219, N2077);
nand NAND2 (N9359, N9349, N7686);
or OR4 (N9360, N9358, N4732, N7193, N8597);
nand NAND4 (N9361, N9341, N5979, N6703, N3849);
or OR3 (N9362, N9356, N2743, N7422);
nor NOR4 (N9363, N9352, N3099, N7286, N586);
xor XOR2 (N9364, N9357, N7332);
buf BUF1 (N9365, N9350);
buf BUF1 (N9366, N9363);
nor NOR3 (N9367, N9361, N1265, N6867);
and AND4 (N9368, N9366, N7781, N5681, N5915);
xor XOR2 (N9369, N9362, N8870);
xor XOR2 (N9370, N9365, N3844);
and AND2 (N9371, N9360, N1074);
not NOT1 (N9372, N9359);
and AND3 (N9373, N9371, N2389, N6509);
xor XOR2 (N9374, N9367, N5010);
and AND3 (N9375, N9374, N8060, N5166);
buf BUF1 (N9376, N9370);
and AND2 (N9377, N9351, N5834);
nor NOR3 (N9378, N9376, N6827, N7532);
or OR2 (N9379, N9369, N2959);
and AND4 (N9380, N9346, N4897, N2260, N5885);
nand NAND2 (N9381, N9375, N8085);
nor NOR4 (N9382, N9379, N9291, N824, N3320);
not NOT1 (N9383, N9355);
xor XOR2 (N9384, N9381, N3607);
buf BUF1 (N9385, N9377);
buf BUF1 (N9386, N9372);
and AND2 (N9387, N9383, N6336);
and AND4 (N9388, N9387, N9250, N8697, N9178);
not NOT1 (N9389, N9380);
or OR3 (N9390, N9378, N1655, N3695);
buf BUF1 (N9391, N9364);
nor NOR3 (N9392, N9390, N2371, N3915);
nor NOR3 (N9393, N9388, N399, N4053);
and AND2 (N9394, N9391, N7610);
and AND4 (N9395, N9394, N7285, N708, N1757);
xor XOR2 (N9396, N9395, N6951);
buf BUF1 (N9397, N9384);
nor NOR2 (N9398, N9385, N7429);
not NOT1 (N9399, N9373);
not NOT1 (N9400, N9399);
buf BUF1 (N9401, N9400);
buf BUF1 (N9402, N9393);
nand NAND4 (N9403, N9401, N6754, N7619, N5807);
nand NAND4 (N9404, N9396, N3714, N2866, N321);
not NOT1 (N9405, N9368);
nand NAND4 (N9406, N9389, N4692, N4242, N3355);
nand NAND4 (N9407, N9403, N4289, N1303, N3817);
not NOT1 (N9408, N9397);
buf BUF1 (N9409, N9392);
or OR2 (N9410, N9386, N7376);
nor NOR4 (N9411, N9410, N8465, N5062, N1645);
buf BUF1 (N9412, N9406);
and AND4 (N9413, N9405, N7267, N3075, N8623);
buf BUF1 (N9414, N9413);
nor NOR4 (N9415, N9408, N5075, N5942, N9347);
buf BUF1 (N9416, N9402);
or OR4 (N9417, N9412, N2424, N4569, N6605);
or OR3 (N9418, N9415, N3865, N1666);
nor NOR4 (N9419, N9411, N9388, N8752, N41);
nand NAND3 (N9420, N9398, N6485, N2510);
xor XOR2 (N9421, N9407, N900);
or OR3 (N9422, N9418, N7458, N3896);
not NOT1 (N9423, N9409);
nand NAND3 (N9424, N9416, N1587, N5221);
and AND4 (N9425, N9424, N2954, N7499, N7479);
buf BUF1 (N9426, N9421);
not NOT1 (N9427, N9426);
nand NAND2 (N9428, N9427, N5978);
xor XOR2 (N9429, N9425, N2650);
not NOT1 (N9430, N9428);
buf BUF1 (N9431, N9382);
nor NOR4 (N9432, N9414, N7450, N7448, N7726);
nor NOR4 (N9433, N9423, N3369, N6794, N5141);
not NOT1 (N9434, N9432);
xor XOR2 (N9435, N9430, N8360);
nand NAND2 (N9436, N9431, N7619);
or OR4 (N9437, N9419, N5254, N8551, N7135);
nand NAND4 (N9438, N9422, N295, N5307, N9414);
buf BUF1 (N9439, N9429);
nor NOR4 (N9440, N9434, N5170, N1611, N6381);
xor XOR2 (N9441, N9435, N4326);
buf BUF1 (N9442, N9436);
xor XOR2 (N9443, N9420, N5600);
and AND3 (N9444, N9433, N6629, N1341);
buf BUF1 (N9445, N9439);
and AND2 (N9446, N9404, N1608);
nor NOR3 (N9447, N9437, N1835, N4219);
or OR4 (N9448, N9442, N2419, N2085, N6247);
nand NAND3 (N9449, N9446, N3359, N1136);
xor XOR2 (N9450, N9447, N6618);
or OR3 (N9451, N9448, N3887, N2316);
nand NAND4 (N9452, N9441, N2948, N348, N3896);
not NOT1 (N9453, N9443);
and AND3 (N9454, N9438, N8502, N4640);
xor XOR2 (N9455, N9453, N246);
and AND4 (N9456, N9445, N1695, N1431, N5190);
or OR3 (N9457, N9454, N348, N7538);
not NOT1 (N9458, N9452);
xor XOR2 (N9459, N9417, N8132);
not NOT1 (N9460, N9457);
and AND3 (N9461, N9458, N3152, N1331);
nand NAND2 (N9462, N9444, N5779);
and AND3 (N9463, N9462, N2205, N8138);
not NOT1 (N9464, N9463);
or OR4 (N9465, N9461, N2354, N1980, N5782);
and AND3 (N9466, N9450, N2471, N471);
xor XOR2 (N9467, N9455, N6224);
nand NAND3 (N9468, N9466, N8082, N5406);
or OR2 (N9469, N9449, N640);
nor NOR4 (N9470, N9469, N4900, N4345, N2546);
and AND4 (N9471, N9467, N5237, N5380, N2514);
and AND3 (N9472, N9440, N192, N248);
or OR3 (N9473, N9470, N3087, N1125);
or OR4 (N9474, N9459, N7148, N1168, N1951);
nor NOR2 (N9475, N9474, N4507);
nand NAND4 (N9476, N9456, N2746, N9430, N5255);
and AND3 (N9477, N9475, N5451, N3890);
not NOT1 (N9478, N9477);
xor XOR2 (N9479, N9464, N6603);
and AND4 (N9480, N9473, N5313, N3531, N5352);
nor NOR4 (N9481, N9472, N1997, N4168, N9225);
and AND2 (N9482, N9479, N6493);
and AND2 (N9483, N9481, N3007);
nor NOR4 (N9484, N9465, N8036, N7618, N6544);
and AND4 (N9485, N9471, N1763, N3707, N4619);
and AND2 (N9486, N9482, N7991);
not NOT1 (N9487, N9484);
xor XOR2 (N9488, N9476, N4788);
nand NAND2 (N9489, N9486, N3503);
buf BUF1 (N9490, N9487);
nand NAND2 (N9491, N9489, N3044);
or OR4 (N9492, N9460, N7975, N6341, N2167);
buf BUF1 (N9493, N9483);
not NOT1 (N9494, N9491);
buf BUF1 (N9495, N9480);
not NOT1 (N9496, N9492);
or OR3 (N9497, N9488, N247, N7097);
nand NAND4 (N9498, N9468, N4906, N3938, N6495);
not NOT1 (N9499, N9495);
xor XOR2 (N9500, N9496, N5394);
not NOT1 (N9501, N9497);
buf BUF1 (N9502, N9500);
nand NAND3 (N9503, N9502, N3100, N2786);
xor XOR2 (N9504, N9494, N1411);
buf BUF1 (N9505, N9504);
and AND2 (N9506, N9478, N8800);
xor XOR2 (N9507, N9485, N2051);
and AND3 (N9508, N9507, N2193, N6072);
not NOT1 (N9509, N9493);
xor XOR2 (N9510, N9509, N6974);
buf BUF1 (N9511, N9503);
nor NOR3 (N9512, N9499, N5272, N1241);
or OR4 (N9513, N9508, N2807, N392, N1672);
nand NAND2 (N9514, N9511, N7828);
not NOT1 (N9515, N9512);
xor XOR2 (N9516, N9501, N1557);
xor XOR2 (N9517, N9490, N7695);
buf BUF1 (N9518, N9506);
nor NOR2 (N9519, N9505, N1679);
buf BUF1 (N9520, N9519);
or OR4 (N9521, N9498, N4490, N8383, N3956);
nand NAND3 (N9522, N9518, N7775, N6647);
nor NOR2 (N9523, N9513, N5055);
and AND3 (N9524, N9520, N3488, N2106);
buf BUF1 (N9525, N9521);
nand NAND2 (N9526, N9515, N7455);
xor XOR2 (N9527, N9526, N2037);
not NOT1 (N9528, N9527);
and AND4 (N9529, N9451, N8856, N2256, N8554);
nand NAND2 (N9530, N9517, N8880);
and AND4 (N9531, N9516, N607, N4205, N4184);
not NOT1 (N9532, N9522);
buf BUF1 (N9533, N9524);
xor XOR2 (N9534, N9529, N5385);
or OR3 (N9535, N9531, N7331, N3810);
or OR4 (N9536, N9534, N6743, N3994, N4032);
xor XOR2 (N9537, N9523, N4827);
buf BUF1 (N9538, N9537);
and AND2 (N9539, N9514, N8980);
or OR3 (N9540, N9532, N170, N94);
nand NAND4 (N9541, N9530, N6124, N1201, N7148);
nand NAND2 (N9542, N9525, N7024);
and AND4 (N9543, N9533, N8789, N4505, N594);
and AND3 (N9544, N9540, N1414, N8364);
or OR3 (N9545, N9510, N3790, N8447);
and AND3 (N9546, N9542, N7106, N1621);
xor XOR2 (N9547, N9539, N1462);
xor XOR2 (N9548, N9547, N9226);
nor NOR2 (N9549, N9544, N9319);
nor NOR4 (N9550, N9545, N6518, N7782, N2344);
or OR4 (N9551, N9536, N7734, N5811, N5237);
xor XOR2 (N9552, N9543, N8198);
and AND4 (N9553, N9546, N1444, N607, N52);
xor XOR2 (N9554, N9552, N150);
or OR2 (N9555, N9549, N6904);
nand NAND3 (N9556, N9541, N5571, N6144);
not NOT1 (N9557, N9556);
nor NOR2 (N9558, N9557, N6407);
xor XOR2 (N9559, N9551, N675);
xor XOR2 (N9560, N9553, N8620);
or OR4 (N9561, N9555, N2832, N2652, N6621);
nand NAND4 (N9562, N9548, N6748, N3293, N9039);
not NOT1 (N9563, N9562);
not NOT1 (N9564, N9535);
and AND3 (N9565, N9559, N7254, N9137);
or OR2 (N9566, N9558, N1607);
not NOT1 (N9567, N9561);
nand NAND2 (N9568, N9528, N7378);
and AND4 (N9569, N9560, N4567, N5229, N6847);
not NOT1 (N9570, N9550);
buf BUF1 (N9571, N9565);
nor NOR4 (N9572, N9568, N2542, N9197, N4827);
buf BUF1 (N9573, N9566);
nor NOR3 (N9574, N9570, N1413, N8934);
or OR3 (N9575, N9569, N7294, N5144);
or OR3 (N9576, N9564, N5143, N7632);
buf BUF1 (N9577, N9575);
nor NOR2 (N9578, N9571, N2074);
xor XOR2 (N9579, N9578, N1226);
nand NAND3 (N9580, N9574, N173, N5432);
and AND3 (N9581, N9576, N5881, N7178);
and AND2 (N9582, N9579, N1358);
buf BUF1 (N9583, N9567);
xor XOR2 (N9584, N9573, N850);
nand NAND3 (N9585, N9538, N2485, N7582);
or OR2 (N9586, N9577, N2753);
or OR3 (N9587, N9581, N4271, N9407);
not NOT1 (N9588, N9583);
and AND3 (N9589, N9563, N2058, N4394);
or OR3 (N9590, N9588, N590, N8390);
xor XOR2 (N9591, N9589, N7169);
xor XOR2 (N9592, N9586, N4557);
nand NAND2 (N9593, N9554, N7301);
nand NAND4 (N9594, N9590, N6624, N3924, N4103);
nand NAND3 (N9595, N9584, N2573, N2019);
not NOT1 (N9596, N9572);
buf BUF1 (N9597, N9585);
or OR2 (N9598, N9593, N657);
not NOT1 (N9599, N9597);
not NOT1 (N9600, N9598);
or OR3 (N9601, N9600, N2085, N2544);
nand NAND4 (N9602, N9599, N2218, N7585, N5989);
or OR4 (N9603, N9582, N900, N1844, N3575);
buf BUF1 (N9604, N9594);
not NOT1 (N9605, N9601);
nor NOR2 (N9606, N9604, N2836);
nor NOR3 (N9607, N9606, N6231, N3077);
xor XOR2 (N9608, N9605, N375);
xor XOR2 (N9609, N9587, N2784);
and AND2 (N9610, N9596, N2999);
and AND3 (N9611, N9603, N4023, N3466);
and AND2 (N9612, N9607, N3580);
nor NOR3 (N9613, N9595, N8090, N3169);
xor XOR2 (N9614, N9591, N1791);
xor XOR2 (N9615, N9610, N6845);
nor NOR2 (N9616, N9612, N8498);
nand NAND2 (N9617, N9611, N2655);
xor XOR2 (N9618, N9617, N9317);
not NOT1 (N9619, N9616);
not NOT1 (N9620, N9619);
or OR2 (N9621, N9608, N162);
buf BUF1 (N9622, N9614);
and AND3 (N9623, N9620, N4781, N5488);
xor XOR2 (N9624, N9592, N1599);
buf BUF1 (N9625, N9623);
not NOT1 (N9626, N9625);
xor XOR2 (N9627, N9621, N6134);
or OR3 (N9628, N9622, N478, N2205);
and AND4 (N9629, N9618, N4041, N7628, N6585);
xor XOR2 (N9630, N9602, N1150);
not NOT1 (N9631, N9580);
not NOT1 (N9632, N9627);
buf BUF1 (N9633, N9630);
nand NAND4 (N9634, N9628, N7627, N7724, N7884);
or OR4 (N9635, N9613, N3958, N7770, N2014);
nor NOR3 (N9636, N9609, N8629, N8184);
nand NAND2 (N9637, N9624, N9232);
nor NOR4 (N9638, N9633, N6009, N7540, N7635);
nor NOR2 (N9639, N9629, N1381);
and AND4 (N9640, N9626, N6371, N2417, N7737);
and AND4 (N9641, N9636, N6870, N9375, N154);
not NOT1 (N9642, N9632);
not NOT1 (N9643, N9641);
buf BUF1 (N9644, N9640);
nor NOR3 (N9645, N9644, N5832, N7737);
or OR2 (N9646, N9645, N4847);
buf BUF1 (N9647, N9615);
not NOT1 (N9648, N9643);
buf BUF1 (N9649, N9634);
xor XOR2 (N9650, N9631, N3120);
xor XOR2 (N9651, N9650, N1112);
or OR3 (N9652, N9637, N5656, N874);
nand NAND3 (N9653, N9647, N2524, N1578);
not NOT1 (N9654, N9649);
or OR4 (N9655, N9639, N2612, N8828, N4019);
and AND3 (N9656, N9642, N8543, N5891);
nand NAND4 (N9657, N9638, N8138, N2656, N1878);
buf BUF1 (N9658, N9651);
xor XOR2 (N9659, N9657, N3901);
or OR3 (N9660, N9646, N5803, N4983);
not NOT1 (N9661, N9656);
not NOT1 (N9662, N9653);
nand NAND3 (N9663, N9661, N4282, N2055);
or OR4 (N9664, N9654, N1875, N2353, N3139);
or OR3 (N9665, N9648, N8960, N202);
or OR4 (N9666, N9660, N2822, N3327, N8664);
nor NOR4 (N9667, N9664, N5359, N668, N1335);
nor NOR4 (N9668, N9655, N177, N2897, N5972);
not NOT1 (N9669, N9659);
buf BUF1 (N9670, N9663);
buf BUF1 (N9671, N9658);
and AND4 (N9672, N9666, N8602, N3127, N3463);
nand NAND4 (N9673, N9652, N2677, N3524, N7533);
not NOT1 (N9674, N9669);
and AND2 (N9675, N9670, N796);
not NOT1 (N9676, N9665);
nand NAND4 (N9677, N9676, N1294, N6146, N5017);
and AND3 (N9678, N9668, N9572, N9650);
xor XOR2 (N9679, N9635, N7743);
not NOT1 (N9680, N9678);
or OR4 (N9681, N9667, N7604, N6960, N5457);
and AND3 (N9682, N9679, N5240, N519);
buf BUF1 (N9683, N9673);
xor XOR2 (N9684, N9672, N8753);
not NOT1 (N9685, N9682);
and AND4 (N9686, N9683, N2586, N4027, N1021);
and AND3 (N9687, N9685, N7919, N6964);
buf BUF1 (N9688, N9671);
xor XOR2 (N9689, N9686, N3292);
not NOT1 (N9690, N9674);
nor NOR4 (N9691, N9688, N3231, N8621, N4820);
xor XOR2 (N9692, N9681, N6199);
not NOT1 (N9693, N9690);
nor NOR3 (N9694, N9689, N1589, N8538);
xor XOR2 (N9695, N9692, N1968);
not NOT1 (N9696, N9662);
nor NOR4 (N9697, N9695, N601, N1780, N7566);
xor XOR2 (N9698, N9680, N3654);
or OR2 (N9699, N9675, N2897);
not NOT1 (N9700, N9697);
nand NAND3 (N9701, N9687, N1843, N8171);
buf BUF1 (N9702, N9691);
or OR2 (N9703, N9699, N7065);
or OR4 (N9704, N9696, N8299, N9601, N4269);
and AND2 (N9705, N9698, N3685);
not NOT1 (N9706, N9677);
and AND4 (N9707, N9705, N2918, N2184, N6956);
xor XOR2 (N9708, N9702, N3442);
nor NOR4 (N9709, N9708, N6506, N9155, N754);
nand NAND3 (N9710, N9693, N1332, N748);
and AND4 (N9711, N9701, N9259, N6316, N8175);
xor XOR2 (N9712, N9704, N2973);
nor NOR3 (N9713, N9709, N835, N7076);
nor NOR2 (N9714, N9700, N5212);
buf BUF1 (N9715, N9711);
and AND4 (N9716, N9684, N7896, N4942, N9055);
and AND4 (N9717, N9715, N8042, N8708, N185);
xor XOR2 (N9718, N9717, N9466);
nor NOR3 (N9719, N9712, N360, N5110);
xor XOR2 (N9720, N9718, N924);
and AND3 (N9721, N9713, N8921, N2913);
or OR2 (N9722, N9719, N9716);
and AND2 (N9723, N3454, N4586);
nor NOR3 (N9724, N9706, N4741, N6026);
or OR3 (N9725, N9703, N7132, N5321);
or OR4 (N9726, N9722, N7661, N8964, N7617);
xor XOR2 (N9727, N9720, N7575);
xor XOR2 (N9728, N9707, N6755);
nand NAND4 (N9729, N9694, N1847, N4489, N6500);
or OR4 (N9730, N9728, N8532, N5117, N2924);
nand NAND2 (N9731, N9724, N7293);
nand NAND4 (N9732, N9726, N4401, N8293, N1153);
buf BUF1 (N9733, N9732);
xor XOR2 (N9734, N9710, N3080);
nor NOR2 (N9735, N9721, N7057);
xor XOR2 (N9736, N9733, N603);
nor NOR2 (N9737, N9727, N691);
xor XOR2 (N9738, N9723, N3036);
not NOT1 (N9739, N9736);
not NOT1 (N9740, N9737);
xor XOR2 (N9741, N9730, N6980);
or OR4 (N9742, N9738, N2124, N4666, N8538);
not NOT1 (N9743, N9742);
not NOT1 (N9744, N9735);
nand NAND4 (N9745, N9740, N8227, N4483, N6982);
or OR3 (N9746, N9729, N117, N937);
not NOT1 (N9747, N9744);
nand NAND3 (N9748, N9714, N3248, N9153);
or OR3 (N9749, N9739, N9354, N442);
nand NAND4 (N9750, N9741, N4188, N141, N6473);
buf BUF1 (N9751, N9725);
or OR4 (N9752, N9731, N1310, N9329, N639);
not NOT1 (N9753, N9752);
nand NAND3 (N9754, N9743, N2282, N1293);
not NOT1 (N9755, N9754);
or OR3 (N9756, N9745, N5092, N3876);
buf BUF1 (N9757, N9753);
nor NOR4 (N9758, N9757, N4873, N4630, N797);
and AND4 (N9759, N9746, N2175, N870, N7452);
or OR4 (N9760, N9758, N7242, N9478, N6835);
and AND4 (N9761, N9747, N7836, N2170, N3022);
nand NAND4 (N9762, N9761, N7399, N2967, N855);
and AND3 (N9763, N9756, N3929, N275);
nand NAND3 (N9764, N9762, N4364, N3604);
or OR4 (N9765, N9734, N878, N8535, N7684);
or OR2 (N9766, N9749, N1767);
or OR4 (N9767, N9751, N7409, N5482, N3);
nor NOR4 (N9768, N9748, N657, N4231, N5582);
and AND3 (N9769, N9766, N9703, N2270);
nand NAND3 (N9770, N9763, N2200, N1318);
nand NAND2 (N9771, N9764, N2878);
xor XOR2 (N9772, N9769, N3210);
buf BUF1 (N9773, N9750);
nor NOR3 (N9774, N9760, N7189, N8949);
nand NAND2 (N9775, N9772, N5863);
and AND2 (N9776, N9773, N8905);
or OR3 (N9777, N9771, N3244, N4579);
not NOT1 (N9778, N9770);
xor XOR2 (N9779, N9777, N3976);
nand NAND3 (N9780, N9767, N665, N5290);
nand NAND4 (N9781, N9776, N2904, N3610, N5350);
xor XOR2 (N9782, N9759, N6411);
and AND2 (N9783, N9774, N5198);
not NOT1 (N9784, N9783);
not NOT1 (N9785, N9782);
or OR2 (N9786, N9768, N9764);
nor NOR4 (N9787, N9786, N6994, N8025, N3517);
nor NOR4 (N9788, N9780, N1645, N6650, N6451);
xor XOR2 (N9789, N9765, N2347);
nor NOR4 (N9790, N9775, N2532, N533, N1279);
and AND4 (N9791, N9787, N1787, N7074, N2464);
nor NOR2 (N9792, N9789, N3959);
or OR4 (N9793, N9779, N7230, N1166, N5435);
nand NAND3 (N9794, N9784, N6353, N2875);
nand NAND2 (N9795, N9781, N7570);
nor NOR2 (N9796, N9785, N914);
nand NAND2 (N9797, N9778, N7723);
xor XOR2 (N9798, N9796, N2706);
buf BUF1 (N9799, N9788);
buf BUF1 (N9800, N9798);
not NOT1 (N9801, N9799);
or OR4 (N9802, N9755, N8233, N985, N4483);
not NOT1 (N9803, N9794);
nor NOR4 (N9804, N9792, N4532, N5776, N90);
xor XOR2 (N9805, N9801, N2632);
and AND3 (N9806, N9790, N7484, N2817);
and AND4 (N9807, N9804, N452, N7322, N6403);
nand NAND3 (N9808, N9802, N5100, N4827);
xor XOR2 (N9809, N9793, N5029);
not NOT1 (N9810, N9797);
buf BUF1 (N9811, N9806);
nand NAND3 (N9812, N9808, N2689, N5464);
or OR3 (N9813, N9803, N8977, N6212);
not NOT1 (N9814, N9810);
nor NOR2 (N9815, N9807, N9196);
xor XOR2 (N9816, N9811, N6871);
nor NOR2 (N9817, N9795, N6296);
xor XOR2 (N9818, N9800, N7862);
buf BUF1 (N9819, N9809);
buf BUF1 (N9820, N9812);
nor NOR4 (N9821, N9816, N57, N1473, N2147);
nand NAND3 (N9822, N9791, N7806, N6965);
buf BUF1 (N9823, N9821);
xor XOR2 (N9824, N9815, N8611);
xor XOR2 (N9825, N9822, N6127);
and AND4 (N9826, N9817, N1349, N7302, N8308);
nor NOR4 (N9827, N9824, N1262, N5393, N4225);
xor XOR2 (N9828, N9818, N7032);
nand NAND3 (N9829, N9825, N4662, N6362);
buf BUF1 (N9830, N9819);
nand NAND2 (N9831, N9820, N3794);
buf BUF1 (N9832, N9827);
buf BUF1 (N9833, N9832);
or OR2 (N9834, N9828, N6179);
not NOT1 (N9835, N9805);
nand NAND2 (N9836, N9829, N7302);
xor XOR2 (N9837, N9833, N4955);
nand NAND2 (N9838, N9836, N3954);
and AND3 (N9839, N9823, N289, N7571);
nor NOR2 (N9840, N9835, N6016);
buf BUF1 (N9841, N9840);
nand NAND2 (N9842, N9813, N2286);
or OR4 (N9843, N9841, N8040, N5428, N2542);
or OR3 (N9844, N9843, N5397, N3937);
or OR3 (N9845, N9839, N8841, N7133);
buf BUF1 (N9846, N9837);
and AND3 (N9847, N9844, N6232, N3171);
nand NAND3 (N9848, N9830, N5842, N8751);
nor NOR3 (N9849, N9846, N527, N8691);
and AND3 (N9850, N9847, N1248, N3253);
not NOT1 (N9851, N9848);
buf BUF1 (N9852, N9838);
and AND2 (N9853, N9826, N6598);
xor XOR2 (N9854, N9853, N6325);
or OR4 (N9855, N9834, N5671, N6426, N8761);
not NOT1 (N9856, N9831);
xor XOR2 (N9857, N9845, N479);
buf BUF1 (N9858, N9849);
not NOT1 (N9859, N9855);
not NOT1 (N9860, N9858);
buf BUF1 (N9861, N9857);
and AND4 (N9862, N9851, N3156, N1186, N7638);
or OR2 (N9863, N9860, N4990);
buf BUF1 (N9864, N9814);
xor XOR2 (N9865, N9842, N7036);
nor NOR3 (N9866, N9859, N5215, N6469);
and AND4 (N9867, N9862, N2010, N5398, N12);
or OR4 (N9868, N9864, N6518, N4083, N2035);
or OR4 (N9869, N9852, N4221, N2635, N2946);
not NOT1 (N9870, N9865);
and AND2 (N9871, N9856, N5548);
nor NOR2 (N9872, N9868, N2188);
nor NOR2 (N9873, N9861, N9297);
or OR3 (N9874, N9866, N488, N6102);
xor XOR2 (N9875, N9874, N9668);
nor NOR3 (N9876, N9863, N2642, N833);
not NOT1 (N9877, N9871);
or OR4 (N9878, N9867, N4750, N9090, N2087);
nand NAND2 (N9879, N9850, N3556);
xor XOR2 (N9880, N9876, N568);
or OR4 (N9881, N9879, N8922, N4767, N1859);
or OR4 (N9882, N9870, N7120, N4288, N7167);
xor XOR2 (N9883, N9869, N8997);
buf BUF1 (N9884, N9875);
not NOT1 (N9885, N9878);
or OR2 (N9886, N9873, N5028);
nor NOR2 (N9887, N9854, N8633);
nand NAND3 (N9888, N9886, N9218, N7768);
nor NOR4 (N9889, N9888, N6616, N5474, N8679);
nor NOR4 (N9890, N9889, N7866, N1803, N5669);
not NOT1 (N9891, N9883);
and AND2 (N9892, N9882, N1063);
and AND4 (N9893, N9892, N7815, N8364, N2474);
buf BUF1 (N9894, N9887);
buf BUF1 (N9895, N9890);
not NOT1 (N9896, N9895);
nand NAND2 (N9897, N9877, N6728);
buf BUF1 (N9898, N9880);
and AND3 (N9899, N9896, N4268, N7582);
buf BUF1 (N9900, N9891);
not NOT1 (N9901, N9897);
buf BUF1 (N9902, N9894);
or OR2 (N9903, N9898, N4625);
nand NAND2 (N9904, N9902, N6503);
buf BUF1 (N9905, N9881);
buf BUF1 (N9906, N9899);
nand NAND2 (N9907, N9900, N2778);
nand NAND3 (N9908, N9885, N1092, N3199);
xor XOR2 (N9909, N9904, N9385);
and AND3 (N9910, N9909, N783, N4312);
nand NAND3 (N9911, N9906, N3812, N904);
or OR2 (N9912, N9907, N1146);
not NOT1 (N9913, N9893);
nor NOR3 (N9914, N9910, N866, N5658);
nor NOR3 (N9915, N9911, N5645, N1543);
and AND3 (N9916, N9901, N790, N9163);
and AND3 (N9917, N9913, N53, N7719);
nor NOR3 (N9918, N9917, N653, N1211);
buf BUF1 (N9919, N9872);
not NOT1 (N9920, N9903);
buf BUF1 (N9921, N9905);
nand NAND4 (N9922, N9919, N2326, N2290, N6736);
xor XOR2 (N9923, N9922, N7186);
or OR4 (N9924, N9908, N6483, N7681, N1733);
nor NOR4 (N9925, N9884, N9588, N4758, N1251);
nor NOR4 (N9926, N9925, N5549, N7348, N2409);
nand NAND2 (N9927, N9918, N5808);
buf BUF1 (N9928, N9915);
nand NAND3 (N9929, N9914, N5804, N221);
or OR4 (N9930, N9921, N8347, N4520, N8062);
and AND4 (N9931, N9920, N4272, N6549, N1945);
and AND3 (N9932, N9924, N7307, N6918);
nor NOR4 (N9933, N9916, N4043, N8744, N8010);
nand NAND4 (N9934, N9931, N8748, N8035, N9493);
nand NAND4 (N9935, N9928, N2195, N4293, N6961);
and AND2 (N9936, N9933, N6854);
buf BUF1 (N9937, N9926);
nor NOR2 (N9938, N9936, N7992);
nand NAND4 (N9939, N9929, N5568, N9413, N7458);
nor NOR4 (N9940, N9934, N1670, N3039, N8647);
not NOT1 (N9941, N9938);
and AND4 (N9942, N9940, N4963, N3177, N8498);
buf BUF1 (N9943, N9935);
or OR4 (N9944, N9942, N3709, N300, N5593);
nand NAND3 (N9945, N9941, N264, N6487);
and AND2 (N9946, N9912, N3661);
nor NOR4 (N9947, N9945, N7291, N5659, N5126);
nand NAND3 (N9948, N9932, N2727, N4146);
not NOT1 (N9949, N9947);
not NOT1 (N9950, N9937);
buf BUF1 (N9951, N9930);
or OR3 (N9952, N9943, N5495, N6200);
and AND2 (N9953, N9923, N5409);
buf BUF1 (N9954, N9948);
not NOT1 (N9955, N9952);
xor XOR2 (N9956, N9953, N305);
xor XOR2 (N9957, N9954, N2686);
nor NOR3 (N9958, N9956, N5882, N9821);
or OR4 (N9959, N9955, N1204, N5643, N5910);
xor XOR2 (N9960, N9946, N9631);
nor NOR4 (N9961, N9949, N6807, N8686, N4678);
or OR2 (N9962, N9961, N9304);
and AND2 (N9963, N9959, N7869);
buf BUF1 (N9964, N9927);
xor XOR2 (N9965, N9944, N8468);
or OR3 (N9966, N9963, N6832, N4620);
buf BUF1 (N9967, N9957);
nor NOR2 (N9968, N9966, N2046);
and AND4 (N9969, N9965, N8125, N1225, N7146);
not NOT1 (N9970, N9950);
xor XOR2 (N9971, N9939, N6436);
buf BUF1 (N9972, N9958);
xor XOR2 (N9973, N9962, N29);
nor NOR2 (N9974, N9967, N8797);
not NOT1 (N9975, N9970);
not NOT1 (N9976, N9964);
xor XOR2 (N9977, N9974, N4276);
xor XOR2 (N9978, N9960, N302);
xor XOR2 (N9979, N9968, N6688);
buf BUF1 (N9980, N9969);
nor NOR4 (N9981, N9979, N4747, N2184, N7150);
buf BUF1 (N9982, N9972);
xor XOR2 (N9983, N9982, N7827);
nor NOR4 (N9984, N9981, N6220, N1222, N6922);
nor NOR3 (N9985, N9980, N1353, N7058);
buf BUF1 (N9986, N9975);
or OR3 (N9987, N9983, N1296, N2105);
nand NAND4 (N9988, N9971, N6776, N9860, N7442);
not NOT1 (N9989, N9951);
nand NAND3 (N9990, N9986, N4579, N6237);
not NOT1 (N9991, N9988);
nor NOR4 (N9992, N9991, N9068, N8461, N1442);
or OR2 (N9993, N9977, N6551);
not NOT1 (N9994, N9989);
xor XOR2 (N9995, N9990, N5846);
and AND3 (N9996, N9987, N4075, N7865);
nor NOR3 (N9997, N9973, N9909, N7767);
or OR2 (N9998, N9993, N132);
buf BUF1 (N9999, N9992);
xor XOR2 (N10000, N9976, N3110);
and AND3 (N10001, N9985, N2363, N5024);
or OR4 (N10002, N9998, N418, N2666, N8061);
or OR4 (N10003, N9994, N4295, N1327, N9239);
and AND3 (N10004, N10003, N9518, N7279);
buf BUF1 (N10005, N9995);
nor NOR3 (N10006, N9984, N8279, N6939);
nor NOR2 (N10007, N10002, N3281);
or OR2 (N10008, N10001, N4175);
nand NAND4 (N10009, N9999, N7925, N7782, N4379);
or OR3 (N10010, N10004, N9466, N4226);
buf BUF1 (N10011, N9978);
xor XOR2 (N10012, N9996, N4880);
buf BUF1 (N10013, N10000);
and AND4 (N10014, N9997, N284, N8765, N2807);
buf BUF1 (N10015, N10006);
nor NOR3 (N10016, N10011, N8242, N994);
xor XOR2 (N10017, N10015, N9379);
xor XOR2 (N10018, N10016, N3499);
buf BUF1 (N10019, N10009);
and AND2 (N10020, N10012, N61);
xor XOR2 (N10021, N10020, N7611);
or OR4 (N10022, N10008, N6568, N7294, N8358);
buf BUF1 (N10023, N10019);
buf BUF1 (N10024, N10018);
buf BUF1 (N10025, N10017);
not NOT1 (N10026, N10024);
not NOT1 (N10027, N10026);
nor NOR3 (N10028, N10010, N3587, N7891);
not NOT1 (N10029, N10007);
xor XOR2 (N10030, N10025, N4745);
nor NOR3 (N10031, N10013, N7034, N1890);
not NOT1 (N10032, N10005);
not NOT1 (N10033, N10029);
and AND4 (N10034, N10023, N8684, N2276, N604);
nor NOR3 (N10035, N10031, N7210, N6532);
not NOT1 (N10036, N10035);
nand NAND2 (N10037, N10014, N1263);
or OR3 (N10038, N10036, N8397, N5281);
or OR4 (N10039, N10030, N8014, N5113, N10025);
nand NAND2 (N10040, N10032, N3946);
xor XOR2 (N10041, N10028, N9184);
nand NAND2 (N10042, N10039, N5253);
nor NOR2 (N10043, N10037, N8183);
or OR3 (N10044, N10022, N2994, N5505);
nor NOR2 (N10045, N10038, N4803);
nand NAND4 (N10046, N10040, N898, N6697, N3805);
not NOT1 (N10047, N10043);
not NOT1 (N10048, N10046);
and AND2 (N10049, N10027, N7806);
nor NOR3 (N10050, N10045, N7934, N7520);
nor NOR2 (N10051, N10021, N9546);
or OR3 (N10052, N10044, N4987, N4182);
not NOT1 (N10053, N10049);
buf BUF1 (N10054, N10050);
nor NOR4 (N10055, N10041, N9533, N7418, N7909);
buf BUF1 (N10056, N10034);
xor XOR2 (N10057, N10051, N8857);
or OR2 (N10058, N10052, N6549);
buf BUF1 (N10059, N10048);
nor NOR2 (N10060, N10033, N5276);
or OR3 (N10061, N10054, N7414, N2646);
nand NAND3 (N10062, N10060, N8690, N6094);
or OR2 (N10063, N10055, N3348);
nand NAND3 (N10064, N10059, N4259, N9590);
nand NAND3 (N10065, N10058, N6436, N1080);
and AND3 (N10066, N10047, N4164, N1602);
and AND3 (N10067, N10062, N1100, N1254);
and AND2 (N10068, N10063, N2401);
and AND2 (N10069, N10042, N7352);
nor NOR2 (N10070, N10061, N864);
xor XOR2 (N10071, N10069, N3786);
or OR4 (N10072, N10070, N7722, N9088, N6517);
xor XOR2 (N10073, N10065, N2545);
and AND4 (N10074, N10068, N2537, N5081, N9463);
or OR2 (N10075, N10057, N10015);
xor XOR2 (N10076, N10064, N4223);
and AND3 (N10077, N10076, N7929, N1446);
nor NOR4 (N10078, N10066, N9972, N3455, N7614);
not NOT1 (N10079, N10075);
not NOT1 (N10080, N10053);
and AND3 (N10081, N10074, N1344, N1965);
or OR3 (N10082, N10056, N4824, N6778);
xor XOR2 (N10083, N10071, N4074);
nor NOR4 (N10084, N10078, N8593, N7896, N4880);
nor NOR4 (N10085, N10083, N8584, N249, N3474);
and AND2 (N10086, N10084, N9165);
buf BUF1 (N10087, N10086);
xor XOR2 (N10088, N10077, N1235);
xor XOR2 (N10089, N10072, N7615);
buf BUF1 (N10090, N10067);
or OR4 (N10091, N10087, N6497, N4615, N1446);
or OR2 (N10092, N10089, N7466);
xor XOR2 (N10093, N10085, N4699);
and AND4 (N10094, N10080, N2685, N965, N1936);
buf BUF1 (N10095, N10073);
and AND4 (N10096, N10094, N139, N1515, N7589);
buf BUF1 (N10097, N10092);
buf BUF1 (N10098, N10095);
buf BUF1 (N10099, N10088);
not NOT1 (N10100, N10097);
xor XOR2 (N10101, N10099, N5965);
not NOT1 (N10102, N10081);
not NOT1 (N10103, N10093);
xor XOR2 (N10104, N10091, N1776);
xor XOR2 (N10105, N10101, N1873);
or OR4 (N10106, N10105, N2926, N7861, N6305);
or OR2 (N10107, N10090, N5283);
buf BUF1 (N10108, N10100);
or OR3 (N10109, N10108, N1184, N6464);
xor XOR2 (N10110, N10098, N6620);
or OR3 (N10111, N10110, N2672, N9493);
and AND3 (N10112, N10103, N6356, N1997);
and AND2 (N10113, N10096, N8027);
nor NOR2 (N10114, N10079, N369);
and AND3 (N10115, N10111, N5730, N5906);
nor NOR3 (N10116, N10106, N7590, N7079);
nor NOR2 (N10117, N10116, N6446);
xor XOR2 (N10118, N10109, N7784);
buf BUF1 (N10119, N10115);
nor NOR4 (N10120, N10107, N7540, N196, N9851);
nor NOR4 (N10121, N10120, N6675, N3364, N7140);
or OR4 (N10122, N10082, N6657, N4474, N1489);
xor XOR2 (N10123, N10117, N3136);
not NOT1 (N10124, N10104);
or OR3 (N10125, N10112, N7506, N1542);
or OR2 (N10126, N10118, N2865);
nand NAND4 (N10127, N10121, N2536, N9581, N10018);
nor NOR2 (N10128, N10122, N9673);
buf BUF1 (N10129, N10114);
nand NAND4 (N10130, N10129, N4058, N6544, N7267);
xor XOR2 (N10131, N10119, N9977);
not NOT1 (N10132, N10124);
buf BUF1 (N10133, N10113);
buf BUF1 (N10134, N10133);
or OR4 (N10135, N10132, N5203, N8463, N8597);
nand NAND4 (N10136, N10127, N7127, N982, N1829);
not NOT1 (N10137, N10125);
xor XOR2 (N10138, N10134, N4112);
xor XOR2 (N10139, N10126, N1504);
not NOT1 (N10140, N10131);
buf BUF1 (N10141, N10140);
nor NOR4 (N10142, N10141, N7954, N883, N6274);
xor XOR2 (N10143, N10139, N1147);
not NOT1 (N10144, N10102);
nand NAND4 (N10145, N10138, N3802, N1540, N4532);
xor XOR2 (N10146, N10128, N7426);
or OR4 (N10147, N10144, N8062, N8413, N4569);
buf BUF1 (N10148, N10137);
nand NAND4 (N10149, N10147, N9893, N9042, N8258);
xor XOR2 (N10150, N10142, N7387);
or OR4 (N10151, N10130, N9555, N8089, N4717);
or OR4 (N10152, N10136, N7499, N6529, N1912);
nand NAND3 (N10153, N10146, N1097, N2136);
not NOT1 (N10154, N10148);
nand NAND3 (N10155, N10152, N1057, N3068);
and AND4 (N10156, N10153, N1824, N9143, N1538);
buf BUF1 (N10157, N10156);
xor XOR2 (N10158, N10157, N1499);
nor NOR4 (N10159, N10150, N3829, N7281, N518);
not NOT1 (N10160, N10159);
not NOT1 (N10161, N10145);
nand NAND4 (N10162, N10158, N4309, N616, N3240);
and AND4 (N10163, N10161, N9681, N5630, N5824);
and AND4 (N10164, N10155, N7042, N6666, N2414);
xor XOR2 (N10165, N10149, N5032);
and AND3 (N10166, N10151, N3934, N5084);
and AND4 (N10167, N10166, N6527, N10052, N5155);
xor XOR2 (N10168, N10164, N4045);
nand NAND3 (N10169, N10160, N4203, N10071);
xor XOR2 (N10170, N10163, N5954);
buf BUF1 (N10171, N10154);
and AND4 (N10172, N10135, N4643, N9886, N6371);
nand NAND2 (N10173, N10171, N9239);
xor XOR2 (N10174, N10143, N4213);
nor NOR3 (N10175, N10173, N8230, N3148);
xor XOR2 (N10176, N10170, N6866);
not NOT1 (N10177, N10165);
xor XOR2 (N10178, N10174, N7558);
buf BUF1 (N10179, N10168);
or OR3 (N10180, N10167, N596, N2013);
nor NOR4 (N10181, N10162, N2134, N391, N6197);
not NOT1 (N10182, N10177);
xor XOR2 (N10183, N10179, N999);
and AND3 (N10184, N10181, N7884, N8176);
buf BUF1 (N10185, N10169);
buf BUF1 (N10186, N10183);
nor NOR2 (N10187, N10184, N4711);
not NOT1 (N10188, N10185);
buf BUF1 (N10189, N10186);
and AND4 (N10190, N10187, N4135, N9602, N177);
nand NAND4 (N10191, N10182, N8390, N4346, N5978);
buf BUF1 (N10192, N10178);
nor NOR2 (N10193, N10180, N7536);
not NOT1 (N10194, N10123);
xor XOR2 (N10195, N10193, N4099);
or OR3 (N10196, N10188, N1579, N4873);
or OR4 (N10197, N10189, N822, N452, N2734);
and AND4 (N10198, N10190, N645, N8782, N392);
and AND2 (N10199, N10176, N9648);
xor XOR2 (N10200, N10194, N7439);
nand NAND2 (N10201, N10172, N10172);
or OR2 (N10202, N10200, N3883);
buf BUF1 (N10203, N10192);
or OR3 (N10204, N10196, N4033, N6050);
nor NOR2 (N10205, N10201, N7805);
xor XOR2 (N10206, N10204, N2558);
nor NOR3 (N10207, N10198, N6733, N3365);
buf BUF1 (N10208, N10207);
nand NAND4 (N10209, N10199, N2174, N4057, N1368);
and AND2 (N10210, N10209, N669);
nand NAND3 (N10211, N10210, N4610, N2677);
nor NOR3 (N10212, N10203, N6207, N38);
not NOT1 (N10213, N10205);
xor XOR2 (N10214, N10202, N8338);
nand NAND2 (N10215, N10208, N7506);
buf BUF1 (N10216, N10212);
xor XOR2 (N10217, N10215, N8260);
or OR3 (N10218, N10175, N8162, N4342);
nor NOR3 (N10219, N10211, N5916, N4678);
xor XOR2 (N10220, N10216, N947);
or OR4 (N10221, N10219, N9068, N4027, N5324);
nand NAND4 (N10222, N10214, N4225, N828, N164);
nand NAND3 (N10223, N10206, N5725, N4182);
buf BUF1 (N10224, N10220);
xor XOR2 (N10225, N10195, N6611);
not NOT1 (N10226, N10197);
nor NOR2 (N10227, N10222, N5016);
buf BUF1 (N10228, N10191);
or OR2 (N10229, N10217, N8895);
and AND3 (N10230, N10223, N3996, N9275);
nor NOR4 (N10231, N10228, N471, N10149, N5263);
nor NOR3 (N10232, N10221, N2537, N288);
or OR2 (N10233, N10229, N4433);
xor XOR2 (N10234, N10225, N5033);
nor NOR2 (N10235, N10230, N3273);
or OR2 (N10236, N10218, N2942);
xor XOR2 (N10237, N10232, N3121);
nor NOR2 (N10238, N10235, N4522);
or OR3 (N10239, N10237, N3622, N3852);
xor XOR2 (N10240, N10224, N8654);
xor XOR2 (N10241, N10238, N287);
not NOT1 (N10242, N10233);
not NOT1 (N10243, N10231);
nand NAND4 (N10244, N10240, N3494, N5449, N493);
xor XOR2 (N10245, N10243, N1740);
and AND4 (N10246, N10213, N3640, N2146, N9369);
buf BUF1 (N10247, N10236);
nor NOR2 (N10248, N10227, N9668);
buf BUF1 (N10249, N10242);
or OR3 (N10250, N10246, N8878, N4963);
and AND3 (N10251, N10250, N8698, N996);
buf BUF1 (N10252, N10247);
xor XOR2 (N10253, N10244, N4565);
nor NOR3 (N10254, N10249, N1944, N9660);
nand NAND3 (N10255, N10248, N5943, N10112);
nor NOR3 (N10256, N10253, N4339, N8705);
and AND4 (N10257, N10239, N8481, N423, N2573);
xor XOR2 (N10258, N10251, N10004);
nand NAND3 (N10259, N10255, N7365, N4363);
and AND4 (N10260, N10241, N1365, N3972, N2551);
xor XOR2 (N10261, N10258, N9773);
buf BUF1 (N10262, N10259);
xor XOR2 (N10263, N10261, N162);
nor NOR3 (N10264, N10257, N9036, N4388);
or OR2 (N10265, N10262, N8513);
and AND4 (N10266, N10265, N9570, N8275, N3627);
xor XOR2 (N10267, N10260, N9176);
not NOT1 (N10268, N10245);
nand NAND4 (N10269, N10263, N760, N2213, N4602);
nor NOR3 (N10270, N10252, N543, N7202);
and AND2 (N10271, N10254, N1591);
not NOT1 (N10272, N10226);
and AND4 (N10273, N10269, N83, N10085, N3442);
xor XOR2 (N10274, N10234, N3254);
buf BUF1 (N10275, N10256);
nand NAND2 (N10276, N10273, N7486);
nor NOR4 (N10277, N10271, N7234, N573, N449);
nor NOR4 (N10278, N10272, N9815, N51, N4345);
xor XOR2 (N10279, N10275, N4084);
nor NOR2 (N10280, N10268, N5277);
nor NOR4 (N10281, N10277, N7912, N6432, N6776);
buf BUF1 (N10282, N10280);
nand NAND2 (N10283, N10266, N7018);
and AND2 (N10284, N10264, N4761);
nand NAND4 (N10285, N10281, N9555, N3454, N5658);
and AND4 (N10286, N10282, N1948, N9627, N1464);
nor NOR3 (N10287, N10285, N1017, N6173);
or OR2 (N10288, N10287, N6465);
or OR3 (N10289, N10274, N4803, N4975);
nand NAND2 (N10290, N10267, N101);
or OR4 (N10291, N10283, N9284, N3, N8428);
and AND2 (N10292, N10279, N9746);
or OR3 (N10293, N10278, N7380, N7696);
buf BUF1 (N10294, N10292);
or OR4 (N10295, N10284, N3792, N6154, N1503);
or OR2 (N10296, N10294, N5927);
nor NOR4 (N10297, N10290, N3188, N1053, N1793);
nor NOR4 (N10298, N10296, N8044, N4989, N1473);
and AND4 (N10299, N10298, N6073, N778, N6227);
nor NOR4 (N10300, N10293, N5962, N9331, N10056);
xor XOR2 (N10301, N10286, N9835);
and AND3 (N10302, N10288, N8085, N6176);
not NOT1 (N10303, N10295);
or OR2 (N10304, N10276, N4559);
and AND3 (N10305, N10304, N5377, N2033);
nor NOR3 (N10306, N10297, N5444, N5390);
xor XOR2 (N10307, N10270, N887);
nand NAND2 (N10308, N10302, N5114);
or OR3 (N10309, N10308, N1623, N4323);
nor NOR3 (N10310, N10291, N1317, N4458);
nand NAND2 (N10311, N10289, N5677);
nor NOR4 (N10312, N10311, N6665, N8974, N7076);
and AND4 (N10313, N10305, N3845, N9612, N8653);
not NOT1 (N10314, N10310);
and AND2 (N10315, N10299, N5897);
or OR4 (N10316, N10315, N2217, N295, N6420);
not NOT1 (N10317, N10303);
not NOT1 (N10318, N10307);
or OR2 (N10319, N10318, N2563);
xor XOR2 (N10320, N10314, N6707);
nand NAND2 (N10321, N10317, N4820);
and AND4 (N10322, N10312, N9438, N6108, N8308);
nor NOR3 (N10323, N10319, N1826, N5940);
nor NOR2 (N10324, N10323, N1776);
buf BUF1 (N10325, N10320);
not NOT1 (N10326, N10306);
not NOT1 (N10327, N10324);
or OR3 (N10328, N10313, N2457, N10076);
nand NAND3 (N10329, N10301, N4483, N6014);
xor XOR2 (N10330, N10328, N6942);
buf BUF1 (N10331, N10322);
nand NAND2 (N10332, N10309, N1691);
xor XOR2 (N10333, N10327, N9231);
nor NOR4 (N10334, N10331, N5106, N6567, N7291);
not NOT1 (N10335, N10334);
and AND4 (N10336, N10330, N8049, N7732, N7149);
nand NAND2 (N10337, N10335, N9135);
and AND3 (N10338, N10321, N1847, N859);
not NOT1 (N10339, N10338);
or OR4 (N10340, N10329, N1322, N9363, N6241);
buf BUF1 (N10341, N10340);
xor XOR2 (N10342, N10325, N3016);
xor XOR2 (N10343, N10336, N6120);
or OR3 (N10344, N10300, N7482, N3169);
and AND3 (N10345, N10342, N3994, N2637);
not NOT1 (N10346, N10332);
nand NAND4 (N10347, N10346, N1063, N5574, N4220);
not NOT1 (N10348, N10343);
nand NAND3 (N10349, N10339, N3988, N508);
buf BUF1 (N10350, N10326);
buf BUF1 (N10351, N10345);
or OR3 (N10352, N10350, N5165, N7235);
nand NAND4 (N10353, N10348, N1930, N8021, N8291);
or OR3 (N10354, N10352, N2161, N3553);
and AND2 (N10355, N10347, N2550);
nand NAND3 (N10356, N10353, N550, N3809);
nand NAND3 (N10357, N10333, N1121, N4599);
and AND3 (N10358, N10357, N180, N10122);
xor XOR2 (N10359, N10355, N2872);
buf BUF1 (N10360, N10316);
buf BUF1 (N10361, N10341);
buf BUF1 (N10362, N10349);
buf BUF1 (N10363, N10356);
nand NAND4 (N10364, N10361, N205, N2869, N2594);
or OR4 (N10365, N10337, N8148, N9877, N4831);
nand NAND3 (N10366, N10364, N535, N5104);
nor NOR2 (N10367, N10358, N5321);
buf BUF1 (N10368, N10354);
and AND2 (N10369, N10362, N647);
or OR4 (N10370, N10360, N8595, N1911, N1342);
nand NAND4 (N10371, N10359, N614, N3803, N1987);
xor XOR2 (N10372, N10370, N8304);
and AND3 (N10373, N10344, N6577, N507);
and AND2 (N10374, N10372, N1681);
buf BUF1 (N10375, N10374);
buf BUF1 (N10376, N10367);
and AND3 (N10377, N10369, N9094, N2533);
buf BUF1 (N10378, N10363);
and AND3 (N10379, N10371, N3037, N7882);
or OR4 (N10380, N10368, N10295, N2929, N5103);
not NOT1 (N10381, N10377);
or OR4 (N10382, N10381, N9718, N9100, N9591);
or OR4 (N10383, N10366, N1508, N5509, N4647);
or OR4 (N10384, N10382, N10166, N9961, N4293);
buf BUF1 (N10385, N10379);
or OR4 (N10386, N10373, N2889, N4195, N9627);
nor NOR2 (N10387, N10365, N3293);
nand NAND2 (N10388, N10351, N8815);
and AND4 (N10389, N10384, N3020, N3026, N6415);
buf BUF1 (N10390, N10387);
nand NAND4 (N10391, N10385, N8217, N3390, N8057);
buf BUF1 (N10392, N10376);
nand NAND3 (N10393, N10375, N7225, N9378);
nor NOR2 (N10394, N10380, N181);
nor NOR2 (N10395, N10388, N1297);
buf BUF1 (N10396, N10393);
and AND4 (N10397, N10383, N5579, N1544, N8811);
xor XOR2 (N10398, N10391, N1697);
or OR2 (N10399, N10389, N1912);
or OR3 (N10400, N10378, N10243, N2114);
and AND2 (N10401, N10396, N5283);
nor NOR2 (N10402, N10386, N3192);
xor XOR2 (N10403, N10390, N866);
xor XOR2 (N10404, N10402, N3710);
and AND4 (N10405, N10397, N9177, N3763, N8277);
and AND3 (N10406, N10395, N4942, N3746);
xor XOR2 (N10407, N10404, N8024);
nand NAND4 (N10408, N10403, N2803, N9125, N2835);
buf BUF1 (N10409, N10405);
nor NOR4 (N10410, N10409, N2506, N6772, N344);
nand NAND4 (N10411, N10399, N834, N9262, N2316);
xor XOR2 (N10412, N10398, N5449);
not NOT1 (N10413, N10406);
or OR3 (N10414, N10401, N8731, N2950);
xor XOR2 (N10415, N10410, N6973);
xor XOR2 (N10416, N10412, N1659);
nand NAND4 (N10417, N10416, N7485, N5814, N4961);
xor XOR2 (N10418, N10400, N4787);
xor XOR2 (N10419, N10408, N10360);
or OR4 (N10420, N10417, N4502, N9761, N9197);
xor XOR2 (N10421, N10414, N2529);
nor NOR3 (N10422, N10419, N520, N8653);
and AND3 (N10423, N10407, N4172, N9646);
xor XOR2 (N10424, N10420, N2159);
and AND3 (N10425, N10394, N3661, N7341);
and AND2 (N10426, N10415, N2573);
not NOT1 (N10427, N10421);
buf BUF1 (N10428, N10425);
nor NOR4 (N10429, N10422, N770, N7223, N2572);
or OR3 (N10430, N10411, N8, N9521);
and AND2 (N10431, N10427, N4113);
nand NAND2 (N10432, N10392, N8924);
or OR2 (N10433, N10424, N9483);
or OR4 (N10434, N10433, N8649, N7365, N6879);
buf BUF1 (N10435, N10434);
nor NOR3 (N10436, N10430, N9288, N6107);
buf BUF1 (N10437, N10432);
or OR2 (N10438, N10429, N8119);
buf BUF1 (N10439, N10413);
buf BUF1 (N10440, N10431);
buf BUF1 (N10441, N10426);
nor NOR4 (N10442, N10437, N7186, N5393, N3284);
nor NOR2 (N10443, N10428, N2538);
not NOT1 (N10444, N10418);
nand NAND3 (N10445, N10443, N8322, N10305);
buf BUF1 (N10446, N10438);
not NOT1 (N10447, N10423);
and AND2 (N10448, N10436, N6162);
or OR2 (N10449, N10439, N1495);
and AND2 (N10450, N10447, N4056);
nor NOR2 (N10451, N10448, N1737);
xor XOR2 (N10452, N10442, N2005);
nand NAND4 (N10453, N10452, N6911, N1932, N7863);
nor NOR3 (N10454, N10445, N1773, N6273);
buf BUF1 (N10455, N10435);
nor NOR4 (N10456, N10440, N9052, N180, N1423);
nand NAND2 (N10457, N10444, N1396);
nor NOR3 (N10458, N10450, N7098, N393);
buf BUF1 (N10459, N10458);
nor NOR4 (N10460, N10453, N6682, N2116, N10176);
or OR3 (N10461, N10441, N1540, N6385);
buf BUF1 (N10462, N10449);
not NOT1 (N10463, N10446);
buf BUF1 (N10464, N10456);
or OR2 (N10465, N10455, N8483);
buf BUF1 (N10466, N10465);
nand NAND4 (N10467, N10461, N6882, N9386, N2871);
or OR2 (N10468, N10466, N1327);
and AND3 (N10469, N10459, N5865, N6906);
nand NAND3 (N10470, N10460, N816, N6913);
or OR2 (N10471, N10469, N1166);
nor NOR4 (N10472, N10467, N3326, N2489, N972);
nand NAND3 (N10473, N10454, N224, N2963);
nand NAND4 (N10474, N10464, N7820, N7306, N479);
or OR2 (N10475, N10471, N7288);
and AND2 (N10476, N10474, N8676);
buf BUF1 (N10477, N10463);
not NOT1 (N10478, N10470);
buf BUF1 (N10479, N10473);
buf BUF1 (N10480, N10478);
and AND2 (N10481, N10476, N1735);
not NOT1 (N10482, N10477);
nand NAND3 (N10483, N10457, N10239, N799);
nand NAND2 (N10484, N10462, N6776);
not NOT1 (N10485, N10451);
xor XOR2 (N10486, N10483, N3196);
buf BUF1 (N10487, N10484);
and AND3 (N10488, N10482, N6172, N2955);
buf BUF1 (N10489, N10480);
nor NOR4 (N10490, N10475, N5526, N6273, N6806);
or OR4 (N10491, N10489, N3263, N8618, N8591);
xor XOR2 (N10492, N10486, N603);
or OR4 (N10493, N10487, N7754, N8066, N6514);
nand NAND3 (N10494, N10493, N5354, N2102);
nand NAND4 (N10495, N10481, N614, N7806, N6954);
nand NAND3 (N10496, N10479, N473, N8621);
or OR2 (N10497, N10494, N6129);
xor XOR2 (N10498, N10496, N6525);
and AND3 (N10499, N10490, N2589, N7381);
or OR2 (N10500, N10491, N6558);
buf BUF1 (N10501, N10495);
nor NOR2 (N10502, N10497, N9040);
xor XOR2 (N10503, N10499, N6533);
and AND3 (N10504, N10500, N7084, N2275);
nor NOR3 (N10505, N10503, N9133, N3974);
not NOT1 (N10506, N10472);
not NOT1 (N10507, N10501);
and AND4 (N10508, N10498, N8331, N9550, N2242);
not NOT1 (N10509, N10468);
nor NOR4 (N10510, N10488, N2128, N3099, N9871);
nor NOR4 (N10511, N10485, N2841, N7731, N9609);
and AND4 (N10512, N10511, N1346, N7994, N6563);
or OR3 (N10513, N10502, N1044, N9850);
not NOT1 (N10514, N10504);
or OR4 (N10515, N10513, N1760, N8094, N2844);
xor XOR2 (N10516, N10509, N9648);
nor NOR4 (N10517, N10492, N9285, N6111, N6419);
nand NAND4 (N10518, N10515, N5474, N420, N2243);
not NOT1 (N10519, N10516);
or OR2 (N10520, N10505, N1348);
buf BUF1 (N10521, N10519);
nor NOR4 (N10522, N10521, N5390, N2306, N7939);
nor NOR2 (N10523, N10517, N2890);
buf BUF1 (N10524, N10506);
nand NAND2 (N10525, N10520, N784);
xor XOR2 (N10526, N10508, N7425);
nor NOR3 (N10527, N10524, N4627, N690);
and AND4 (N10528, N10525, N795, N4473, N2450);
xor XOR2 (N10529, N10512, N2328);
or OR2 (N10530, N10518, N2064);
or OR3 (N10531, N10530, N3952, N611);
buf BUF1 (N10532, N10531);
buf BUF1 (N10533, N10532);
nor NOR2 (N10534, N10523, N3459);
buf BUF1 (N10535, N10522);
nand NAND2 (N10536, N10535, N9346);
xor XOR2 (N10537, N10510, N5396);
or OR4 (N10538, N10534, N9673, N7569, N476);
not NOT1 (N10539, N10533);
nor NOR3 (N10540, N10526, N796, N6710);
xor XOR2 (N10541, N10527, N2708);
buf BUF1 (N10542, N10536);
nor NOR3 (N10543, N10539, N4174, N5772);
not NOT1 (N10544, N10529);
or OR3 (N10545, N10544, N9953, N7231);
buf BUF1 (N10546, N10542);
xor XOR2 (N10547, N10507, N2974);
not NOT1 (N10548, N10528);
and AND3 (N10549, N10538, N4385, N2859);
not NOT1 (N10550, N10547);
or OR3 (N10551, N10550, N5488, N5820);
nand NAND4 (N10552, N10541, N2065, N9234, N3259);
xor XOR2 (N10553, N10551, N9788);
nor NOR2 (N10554, N10546, N9372);
xor XOR2 (N10555, N10514, N8235);
and AND4 (N10556, N10549, N204, N2399, N8816);
xor XOR2 (N10557, N10537, N567);
nand NAND4 (N10558, N10543, N3392, N2316, N1049);
not NOT1 (N10559, N10552);
or OR4 (N10560, N10557, N1391, N5150, N8332);
nand NAND2 (N10561, N10560, N9349);
nor NOR2 (N10562, N10558, N1742);
and AND2 (N10563, N10555, N171);
nor NOR3 (N10564, N10562, N10377, N3601);
nand NAND3 (N10565, N10564, N2103, N3642);
nor NOR4 (N10566, N10548, N7867, N1446, N10214);
xor XOR2 (N10567, N10545, N8238);
or OR3 (N10568, N10554, N6048, N9593);
and AND2 (N10569, N10566, N3705);
and AND2 (N10570, N10561, N2713);
not NOT1 (N10571, N10556);
not NOT1 (N10572, N10571);
or OR3 (N10573, N10565, N1163, N1127);
nand NAND4 (N10574, N10559, N5987, N9184, N10331);
and AND4 (N10575, N10572, N6453, N2480, N729);
or OR4 (N10576, N10575, N1738, N1514, N6517);
and AND3 (N10577, N10567, N9638, N3197);
buf BUF1 (N10578, N10573);
and AND4 (N10579, N10540, N6527, N9962, N7658);
buf BUF1 (N10580, N10576);
and AND4 (N10581, N10568, N1880, N1373, N1447);
and AND2 (N10582, N10553, N4264);
not NOT1 (N10583, N10582);
buf BUF1 (N10584, N10577);
or OR3 (N10585, N10570, N9574, N5311);
not NOT1 (N10586, N10585);
not NOT1 (N10587, N10583);
or OR2 (N10588, N10578, N2901);
not NOT1 (N10589, N10588);
nor NOR3 (N10590, N10569, N3669, N3201);
or OR4 (N10591, N10586, N5500, N96, N1050);
not NOT1 (N10592, N10563);
nor NOR3 (N10593, N10580, N1078, N10468);
nor NOR3 (N10594, N10579, N782, N239);
nor NOR2 (N10595, N10587, N6153);
xor XOR2 (N10596, N10574, N6918);
and AND4 (N10597, N10581, N7931, N6815, N10539);
buf BUF1 (N10598, N10594);
nor NOR2 (N10599, N10598, N7307);
not NOT1 (N10600, N10591);
or OR4 (N10601, N10595, N280, N8504, N2002);
nand NAND4 (N10602, N10592, N8678, N9644, N4694);
or OR4 (N10603, N10600, N10045, N9146, N98);
buf BUF1 (N10604, N10584);
or OR3 (N10605, N10590, N5129, N9335);
nand NAND3 (N10606, N10601, N8409, N1844);
or OR3 (N10607, N10604, N242, N427);
xor XOR2 (N10608, N10607, N10314);
buf BUF1 (N10609, N10605);
xor XOR2 (N10610, N10606, N5918);
buf BUF1 (N10611, N10608);
nand NAND3 (N10612, N10602, N6219, N1472);
nor NOR3 (N10613, N10603, N6276, N2942);
and AND4 (N10614, N10597, N4714, N10590, N4060);
xor XOR2 (N10615, N10610, N9059);
and AND4 (N10616, N10599, N8891, N2175, N5534);
not NOT1 (N10617, N10615);
nor NOR3 (N10618, N10616, N9396, N3322);
nor NOR4 (N10619, N10589, N8031, N6545, N597);
xor XOR2 (N10620, N10609, N9679);
or OR4 (N10621, N10617, N4325, N929, N10461);
nand NAND3 (N10622, N10596, N9014, N3528);
and AND2 (N10623, N10620, N5343);
not NOT1 (N10624, N10623);
not NOT1 (N10625, N10613);
nor NOR2 (N10626, N10612, N3174);
nand NAND2 (N10627, N10625, N6007);
xor XOR2 (N10628, N10621, N10458);
buf BUF1 (N10629, N10593);
and AND3 (N10630, N10622, N6544, N777);
xor XOR2 (N10631, N10614, N10475);
not NOT1 (N10632, N10629);
nor NOR4 (N10633, N10619, N6328, N1783, N1384);
nor NOR3 (N10634, N10633, N213, N3927);
xor XOR2 (N10635, N10626, N6206);
or OR3 (N10636, N10631, N7442, N1353);
buf BUF1 (N10637, N10634);
buf BUF1 (N10638, N10630);
nor NOR2 (N10639, N10637, N8810);
not NOT1 (N10640, N10636);
nor NOR4 (N10641, N10639, N427, N6500, N415);
not NOT1 (N10642, N10611);
buf BUF1 (N10643, N10641);
and AND3 (N10644, N10640, N2864, N641);
nor NOR4 (N10645, N10638, N10254, N10292, N8649);
nand NAND3 (N10646, N10645, N5717, N7097);
nor NOR2 (N10647, N10627, N7887);
xor XOR2 (N10648, N10647, N4491);
not NOT1 (N10649, N10643);
nor NOR2 (N10650, N10644, N1961);
nand NAND2 (N10651, N10642, N4780);
or OR4 (N10652, N10649, N1976, N7881, N9965);
or OR3 (N10653, N10652, N2197, N4332);
buf BUF1 (N10654, N10646);
buf BUF1 (N10655, N10624);
buf BUF1 (N10656, N10653);
xor XOR2 (N10657, N10648, N7596);
and AND4 (N10658, N10635, N5757, N2855, N6335);
not NOT1 (N10659, N10654);
xor XOR2 (N10660, N10659, N4785);
xor XOR2 (N10661, N10651, N9038);
or OR2 (N10662, N10656, N6210);
xor XOR2 (N10663, N10632, N522);
xor XOR2 (N10664, N10618, N4404);
xor XOR2 (N10665, N10650, N996);
xor XOR2 (N10666, N10661, N4519);
or OR4 (N10667, N10663, N2499, N532, N2425);
not NOT1 (N10668, N10664);
buf BUF1 (N10669, N10668);
nand NAND4 (N10670, N10665, N4892, N9935, N2581);
nor NOR4 (N10671, N10670, N1994, N721, N7156);
and AND4 (N10672, N10671, N2161, N6627, N7921);
nand NAND2 (N10673, N10657, N10164);
xor XOR2 (N10674, N10655, N1202);
nor NOR2 (N10675, N10628, N9727);
nand NAND4 (N10676, N10673, N1937, N5494, N7302);
or OR3 (N10677, N10675, N5848, N866);
or OR2 (N10678, N10669, N7748);
and AND3 (N10679, N10667, N4553, N8349);
or OR4 (N10680, N10672, N3080, N5278, N4307);
or OR3 (N10681, N10679, N453, N4826);
nor NOR2 (N10682, N10660, N259);
not NOT1 (N10683, N10678);
buf BUF1 (N10684, N10682);
xor XOR2 (N10685, N10681, N7558);
not NOT1 (N10686, N10662);
xor XOR2 (N10687, N10666, N7748);
buf BUF1 (N10688, N10658);
buf BUF1 (N10689, N10676);
buf BUF1 (N10690, N10689);
xor XOR2 (N10691, N10683, N3083);
not NOT1 (N10692, N10687);
and AND4 (N10693, N10685, N2245, N10562, N5951);
nor NOR2 (N10694, N10686, N4163);
nor NOR3 (N10695, N10680, N5812, N3266);
and AND3 (N10696, N10693, N5908, N2109);
nor NOR3 (N10697, N10692, N10401, N4519);
buf BUF1 (N10698, N10674);
not NOT1 (N10699, N10697);
or OR3 (N10700, N10696, N6241, N5702);
or OR2 (N10701, N10698, N9332);
nand NAND2 (N10702, N10700, N256);
or OR2 (N10703, N10690, N1606);
buf BUF1 (N10704, N10691);
and AND3 (N10705, N10688, N2613, N787);
nand NAND4 (N10706, N10695, N4148, N9340, N3112);
not NOT1 (N10707, N10705);
nor NOR3 (N10708, N10677, N2779, N4085);
nor NOR3 (N10709, N10707, N4469, N7110);
nand NAND4 (N10710, N10702, N905, N7822, N1479);
xor XOR2 (N10711, N10704, N2262);
buf BUF1 (N10712, N10709);
not NOT1 (N10713, N10710);
nor NOR2 (N10714, N10708, N4776);
xor XOR2 (N10715, N10701, N7866);
and AND2 (N10716, N10699, N8606);
nand NAND4 (N10717, N10714, N122, N419, N10028);
or OR2 (N10718, N10706, N4480);
or OR4 (N10719, N10717, N5276, N8806, N10148);
nor NOR2 (N10720, N10719, N4152);
and AND3 (N10721, N10713, N8085, N10367);
nand NAND2 (N10722, N10684, N1605);
buf BUF1 (N10723, N10721);
nand NAND3 (N10724, N10720, N4241, N1650);
not NOT1 (N10725, N10694);
buf BUF1 (N10726, N10722);
nor NOR2 (N10727, N10725, N10452);
nand NAND3 (N10728, N10718, N8286, N6524);
and AND3 (N10729, N10703, N7865, N3025);
nand NAND3 (N10730, N10715, N4453, N1632);
not NOT1 (N10731, N10728);
xor XOR2 (N10732, N10711, N8035);
or OR4 (N10733, N10732, N4254, N3758, N1715);
or OR2 (N10734, N10723, N10585);
nor NOR3 (N10735, N10733, N2138, N8603);
nand NAND4 (N10736, N10731, N7968, N1417, N753);
not NOT1 (N10737, N10716);
not NOT1 (N10738, N10726);
and AND2 (N10739, N10727, N5131);
not NOT1 (N10740, N10738);
or OR3 (N10741, N10712, N6334, N3353);
not NOT1 (N10742, N10729);
nand NAND2 (N10743, N10724, N7361);
nand NAND3 (N10744, N10737, N9890, N9333);
not NOT1 (N10745, N10739);
or OR3 (N10746, N10730, N10375, N1875);
not NOT1 (N10747, N10735);
not NOT1 (N10748, N10736);
and AND2 (N10749, N10743, N4685);
and AND3 (N10750, N10740, N8862, N2863);
buf BUF1 (N10751, N10749);
nand NAND2 (N10752, N10746, N7972);
nor NOR4 (N10753, N10745, N1639, N4707, N1867);
and AND4 (N10754, N10753, N7347, N1337, N7538);
or OR2 (N10755, N10754, N1621);
nor NOR4 (N10756, N10750, N7428, N434, N4233);
and AND2 (N10757, N10748, N9296);
or OR3 (N10758, N10747, N2613, N3386);
nand NAND3 (N10759, N10742, N8714, N845);
or OR3 (N10760, N10756, N1779, N8713);
or OR2 (N10761, N10759, N6572);
or OR4 (N10762, N10760, N7323, N6622, N3294);
nor NOR4 (N10763, N10752, N6696, N885, N2441);
and AND4 (N10764, N10758, N2958, N10675, N2628);
buf BUF1 (N10765, N10755);
and AND2 (N10766, N10734, N9399);
or OR4 (N10767, N10766, N6299, N5802, N9243);
not NOT1 (N10768, N10767);
and AND3 (N10769, N10741, N2742, N4966);
and AND2 (N10770, N10768, N4195);
xor XOR2 (N10771, N10769, N10615);
or OR2 (N10772, N10751, N1038);
not NOT1 (N10773, N10757);
nor NOR2 (N10774, N10764, N7117);
xor XOR2 (N10775, N10761, N5339);
nor NOR3 (N10776, N10773, N5146, N1303);
nor NOR3 (N10777, N10765, N5391, N7844);
buf BUF1 (N10778, N10775);
xor XOR2 (N10779, N10772, N3759);
xor XOR2 (N10780, N10770, N4081);
not NOT1 (N10781, N10774);
or OR4 (N10782, N10763, N4604, N386, N8891);
nand NAND3 (N10783, N10778, N9479, N2139);
and AND2 (N10784, N10780, N6494);
or OR2 (N10785, N10784, N7193);
nor NOR2 (N10786, N10783, N3401);
nor NOR3 (N10787, N10785, N3593, N10598);
nor NOR3 (N10788, N10744, N6109, N9131);
not NOT1 (N10789, N10788);
nor NOR4 (N10790, N10771, N3278, N9411, N6412);
not NOT1 (N10791, N10777);
not NOT1 (N10792, N10762);
or OR2 (N10793, N10787, N8904);
or OR2 (N10794, N10782, N5443);
and AND3 (N10795, N10791, N1273, N6123);
nand NAND4 (N10796, N10792, N9432, N154, N1561);
and AND3 (N10797, N10789, N3489, N6680);
nor NOR2 (N10798, N10794, N10213);
not NOT1 (N10799, N10795);
and AND4 (N10800, N10781, N2579, N2192, N6528);
and AND3 (N10801, N10798, N4655, N6935);
or OR4 (N10802, N10801, N2774, N10653, N1784);
and AND3 (N10803, N10797, N4499, N6697);
nand NAND2 (N10804, N10776, N10241);
xor XOR2 (N10805, N10790, N5921);
nor NOR2 (N10806, N10800, N1397);
not NOT1 (N10807, N10806);
or OR2 (N10808, N10779, N7095);
or OR3 (N10809, N10807, N5241, N1992);
and AND2 (N10810, N10803, N742);
and AND4 (N10811, N10808, N157, N5584, N5945);
xor XOR2 (N10812, N10810, N9356);
not NOT1 (N10813, N10811);
nand NAND3 (N10814, N10804, N3202, N4762);
and AND4 (N10815, N10813, N781, N4775, N10786);
xor XOR2 (N10816, N2411, N8314);
nand NAND2 (N10817, N10802, N6846);
and AND3 (N10818, N10814, N879, N143);
not NOT1 (N10819, N10817);
nand NAND2 (N10820, N10799, N6007);
nand NAND2 (N10821, N10818, N5237);
not NOT1 (N10822, N10805);
not NOT1 (N10823, N10793);
nor NOR2 (N10824, N10820, N7643);
and AND4 (N10825, N10823, N6665, N871, N10513);
xor XOR2 (N10826, N10809, N5994);
buf BUF1 (N10827, N10796);
or OR4 (N10828, N10819, N9935, N6447, N7753);
nand NAND3 (N10829, N10812, N3560, N815);
and AND4 (N10830, N10827, N10676, N3322, N5070);
not NOT1 (N10831, N10826);
not NOT1 (N10832, N10828);
nor NOR3 (N10833, N10824, N4345, N5005);
not NOT1 (N10834, N10832);
and AND3 (N10835, N10833, N2794, N1700);
not NOT1 (N10836, N10829);
xor XOR2 (N10837, N10834, N3025);
and AND3 (N10838, N10831, N4420, N3576);
and AND3 (N10839, N10836, N6098, N4633);
nor NOR2 (N10840, N10835, N237);
not NOT1 (N10841, N10839);
xor XOR2 (N10842, N10830, N5655);
and AND2 (N10843, N10842, N9442);
nand NAND2 (N10844, N10821, N8148);
xor XOR2 (N10845, N10837, N10034);
buf BUF1 (N10846, N10816);
buf BUF1 (N10847, N10822);
nand NAND3 (N10848, N10845, N9151, N5516);
nor NOR2 (N10849, N10840, N7595);
or OR4 (N10850, N10846, N10519, N5278, N1655);
or OR2 (N10851, N10850, N3558);
xor XOR2 (N10852, N10847, N7873);
and AND2 (N10853, N10843, N2256);
nor NOR3 (N10854, N10838, N5333, N5093);
buf BUF1 (N10855, N10852);
and AND2 (N10856, N10849, N8677);
nor NOR4 (N10857, N10825, N3501, N4460, N9953);
or OR2 (N10858, N10851, N3823);
or OR3 (N10859, N10815, N5605, N1643);
nand NAND2 (N10860, N10857, N1068);
not NOT1 (N10861, N10854);
or OR2 (N10862, N10853, N7196);
nor NOR3 (N10863, N10841, N1351, N10745);
and AND3 (N10864, N10844, N3835, N4420);
not NOT1 (N10865, N10860);
buf BUF1 (N10866, N10865);
or OR4 (N10867, N10848, N3871, N499, N1148);
nor NOR4 (N10868, N10855, N10184, N10382, N505);
or OR2 (N10869, N10866, N1553);
nand NAND3 (N10870, N10859, N10619, N2893);
nor NOR2 (N10871, N10867, N6533);
nor NOR4 (N10872, N10861, N2849, N5541, N10531);
and AND4 (N10873, N10872, N232, N9722, N8983);
nor NOR3 (N10874, N10869, N7507, N2963);
nand NAND2 (N10875, N10874, N1402);
nor NOR3 (N10876, N10858, N9498, N3639);
not NOT1 (N10877, N10873);
and AND2 (N10878, N10856, N3983);
and AND2 (N10879, N10871, N3174);
not NOT1 (N10880, N10878);
or OR3 (N10881, N10863, N4182, N2104);
nor NOR4 (N10882, N10877, N10637, N7506, N353);
not NOT1 (N10883, N10876);
nand NAND3 (N10884, N10881, N885, N4058);
or OR3 (N10885, N10883, N470, N1647);
or OR4 (N10886, N10885, N7470, N482, N9842);
or OR3 (N10887, N10884, N3875, N9297);
not NOT1 (N10888, N10862);
buf BUF1 (N10889, N10868);
not NOT1 (N10890, N10887);
buf BUF1 (N10891, N10882);
and AND4 (N10892, N10890, N4617, N1393, N9282);
and AND3 (N10893, N10889, N10641, N10193);
buf BUF1 (N10894, N10875);
nand NAND2 (N10895, N10864, N6467);
or OR2 (N10896, N10870, N7988);
nand NAND3 (N10897, N10891, N9559, N5329);
nor NOR3 (N10898, N10894, N4359, N10150);
nor NOR4 (N10899, N10886, N3774, N535, N1181);
and AND2 (N10900, N10892, N269);
and AND4 (N10901, N10899, N383, N5470, N3843);
nand NAND4 (N10902, N10896, N6322, N1468, N2288);
or OR4 (N10903, N10901, N6279, N10780, N9523);
nor NOR3 (N10904, N10898, N4339, N3738);
not NOT1 (N10905, N10880);
xor XOR2 (N10906, N10902, N5300);
or OR2 (N10907, N10879, N3182);
or OR4 (N10908, N10904, N2666, N39, N6873);
nor NOR2 (N10909, N10895, N2312);
nor NOR3 (N10910, N10909, N10554, N9154);
not NOT1 (N10911, N10893);
nor NOR3 (N10912, N10911, N6713, N9918);
nor NOR4 (N10913, N10905, N4903, N2683, N8672);
and AND2 (N10914, N10906, N4380);
nor NOR4 (N10915, N10903, N6549, N8048, N2255);
not NOT1 (N10916, N10908);
or OR3 (N10917, N10910, N3504, N5315);
not NOT1 (N10918, N10912);
not NOT1 (N10919, N10918);
nand NAND3 (N10920, N10919, N1963, N9137);
buf BUF1 (N10921, N10913);
not NOT1 (N10922, N10897);
nor NOR3 (N10923, N10907, N5133, N8768);
buf BUF1 (N10924, N10900);
nand NAND3 (N10925, N10917, N5442, N5350);
xor XOR2 (N10926, N10922, N1416);
not NOT1 (N10927, N10915);
not NOT1 (N10928, N10926);
xor XOR2 (N10929, N10923, N687);
or OR4 (N10930, N10888, N5273, N5237, N5053);
or OR3 (N10931, N10914, N333, N9906);
xor XOR2 (N10932, N10925, N6717);
or OR2 (N10933, N10929, N721);
buf BUF1 (N10934, N10921);
nor NOR4 (N10935, N10932, N6059, N2613, N556);
nor NOR4 (N10936, N10930, N2236, N896, N10048);
not NOT1 (N10937, N10928);
or OR4 (N10938, N10937, N5952, N4985, N10099);
nor NOR3 (N10939, N10927, N1149, N6148);
not NOT1 (N10940, N10933);
not NOT1 (N10941, N10924);
or OR4 (N10942, N10935, N7453, N7428, N2805);
xor XOR2 (N10943, N10942, N350);
or OR2 (N10944, N10920, N8670);
nand NAND4 (N10945, N10940, N6369, N8248, N587);
xor XOR2 (N10946, N10936, N853);
or OR4 (N10947, N10941, N6638, N7784, N7053);
or OR3 (N10948, N10947, N725, N2530);
buf BUF1 (N10949, N10946);
buf BUF1 (N10950, N10916);
xor XOR2 (N10951, N10944, N1404);
buf BUF1 (N10952, N10951);
xor XOR2 (N10953, N10938, N4734);
not NOT1 (N10954, N10949);
nand NAND3 (N10955, N10950, N941, N8644);
not NOT1 (N10956, N10952);
not NOT1 (N10957, N10956);
and AND2 (N10958, N10954, N2739);
xor XOR2 (N10959, N10945, N4710);
or OR4 (N10960, N10931, N3867, N3003, N3229);
or OR2 (N10961, N10957, N8203);
nor NOR3 (N10962, N10958, N1690, N8098);
nand NAND3 (N10963, N10955, N8890, N4474);
not NOT1 (N10964, N10943);
not NOT1 (N10965, N10963);
nor NOR3 (N10966, N10965, N5422, N6806);
nand NAND3 (N10967, N10960, N8476, N5541);
nor NOR3 (N10968, N10939, N4835, N6334);
or OR2 (N10969, N10968, N4302);
and AND2 (N10970, N10961, N3094);
or OR2 (N10971, N10959, N6887);
buf BUF1 (N10972, N10969);
not NOT1 (N10973, N10953);
not NOT1 (N10974, N10972);
xor XOR2 (N10975, N10971, N206);
and AND2 (N10976, N10975, N3862);
buf BUF1 (N10977, N10964);
buf BUF1 (N10978, N10973);
not NOT1 (N10979, N10962);
buf BUF1 (N10980, N10967);
xor XOR2 (N10981, N10966, N2612);
buf BUF1 (N10982, N10977);
not NOT1 (N10983, N10970);
nor NOR2 (N10984, N10979, N1215);
nor NOR3 (N10985, N10934, N5552, N9374);
or OR2 (N10986, N10984, N4749);
nor NOR2 (N10987, N10974, N9810);
and AND3 (N10988, N10985, N4896, N7797);
or OR3 (N10989, N10986, N1871, N7103);
nor NOR3 (N10990, N10988, N10506, N693);
buf BUF1 (N10991, N10983);
not NOT1 (N10992, N10987);
not NOT1 (N10993, N10981);
xor XOR2 (N10994, N10976, N10277);
and AND4 (N10995, N10980, N9173, N8976, N7520);
buf BUF1 (N10996, N10982);
not NOT1 (N10997, N10993);
and AND2 (N10998, N10994, N9856);
and AND2 (N10999, N10997, N5147);
xor XOR2 (N11000, N10999, N10926);
not NOT1 (N11001, N10989);
xor XOR2 (N11002, N10948, N2080);
or OR3 (N11003, N11000, N9100, N9825);
nand NAND3 (N11004, N10990, N6453, N4504);
and AND4 (N11005, N10992, N4479, N1852, N8151);
buf BUF1 (N11006, N10998);
buf BUF1 (N11007, N11005);
not NOT1 (N11008, N11003);
or OR4 (N11009, N11006, N1464, N1776, N9919);
xor XOR2 (N11010, N11008, N10870);
not NOT1 (N11011, N11010);
not NOT1 (N11012, N11004);
or OR4 (N11013, N10978, N400, N838, N7000);
not NOT1 (N11014, N10996);
and AND4 (N11015, N11012, N8980, N1769, N7221);
or OR4 (N11016, N11014, N8383, N4990, N3022);
and AND3 (N11017, N11016, N6136, N4471);
nor NOR3 (N11018, N11009, N3146, N4418);
nand NAND3 (N11019, N11007, N10077, N9264);
nor NOR3 (N11020, N10991, N6600, N10994);
or OR2 (N11021, N11013, N10516);
xor XOR2 (N11022, N11002, N6292);
not NOT1 (N11023, N11001);
not NOT1 (N11024, N11015);
xor XOR2 (N11025, N10995, N2009);
and AND3 (N11026, N11017, N7176, N764);
buf BUF1 (N11027, N11024);
nand NAND4 (N11028, N11021, N2565, N10720, N1748);
and AND2 (N11029, N11019, N8522);
nor NOR3 (N11030, N11018, N5817, N6410);
nor NOR4 (N11031, N11029, N7440, N10600, N8808);
nand NAND3 (N11032, N11011, N3211, N8914);
or OR3 (N11033, N11020, N1044, N10886);
nand NAND2 (N11034, N11027, N6430);
buf BUF1 (N11035, N11033);
xor XOR2 (N11036, N11035, N1939);
and AND3 (N11037, N11023, N4725, N7769);
and AND2 (N11038, N11036, N3909);
buf BUF1 (N11039, N11034);
not NOT1 (N11040, N11031);
or OR4 (N11041, N11032, N7393, N7543, N8439);
nand NAND3 (N11042, N11028, N213, N7101);
nor NOR3 (N11043, N11037, N396, N3744);
nor NOR2 (N11044, N11025, N204);
xor XOR2 (N11045, N11042, N5629);
not NOT1 (N11046, N11041);
xor XOR2 (N11047, N11022, N10050);
and AND4 (N11048, N11040, N6987, N10995, N2681);
not NOT1 (N11049, N11048);
nor NOR2 (N11050, N11047, N1986);
not NOT1 (N11051, N11026);
and AND4 (N11052, N11045, N8573, N1423, N1259);
or OR2 (N11053, N11043, N10678);
nor NOR3 (N11054, N11049, N3935, N10179);
not NOT1 (N11055, N11030);
xor XOR2 (N11056, N11053, N10334);
buf BUF1 (N11057, N11052);
nand NAND4 (N11058, N11055, N46, N5766, N6831);
nand NAND2 (N11059, N11058, N10034);
not NOT1 (N11060, N11051);
not NOT1 (N11061, N11060);
or OR2 (N11062, N11057, N1767);
buf BUF1 (N11063, N11056);
and AND4 (N11064, N11059, N3556, N9578, N460);
and AND3 (N11065, N11054, N8808, N3382);
buf BUF1 (N11066, N11050);
buf BUF1 (N11067, N11039);
nor NOR4 (N11068, N11038, N4458, N1409, N1216);
and AND4 (N11069, N11046, N130, N960, N6449);
or OR4 (N11070, N11065, N7568, N5889, N1226);
nor NOR3 (N11071, N11061, N6725, N3652);
and AND2 (N11072, N11068, N5227);
not NOT1 (N11073, N11069);
xor XOR2 (N11074, N11066, N2635);
and AND4 (N11075, N11072, N10468, N6473, N2457);
nor NOR4 (N11076, N11075, N2828, N2284, N7156);
nor NOR2 (N11077, N11070, N8633);
and AND2 (N11078, N11063, N10371);
nand NAND4 (N11079, N11071, N6612, N1123, N10714);
and AND4 (N11080, N11067, N1558, N5559, N10775);
or OR3 (N11081, N11076, N4148, N1059);
not NOT1 (N11082, N11074);
and AND4 (N11083, N11077, N6184, N9615, N6125);
or OR2 (N11084, N11044, N8784);
not NOT1 (N11085, N11078);
nand NAND4 (N11086, N11080, N7282, N6795, N10551);
xor XOR2 (N11087, N11084, N9016);
xor XOR2 (N11088, N11083, N9855);
nand NAND3 (N11089, N11062, N8712, N9966);
or OR2 (N11090, N11088, N8115);
nor NOR2 (N11091, N11079, N7075);
not NOT1 (N11092, N11090);
buf BUF1 (N11093, N11064);
nor NOR3 (N11094, N11087, N2355, N3707);
nand NAND4 (N11095, N11089, N1329, N892, N7591);
and AND3 (N11096, N11081, N2743, N2174);
not NOT1 (N11097, N11082);
and AND4 (N11098, N11096, N5584, N5188, N7228);
xor XOR2 (N11099, N11093, N3801);
and AND4 (N11100, N11097, N10984, N3022, N2375);
nand NAND2 (N11101, N11073, N8865);
buf BUF1 (N11102, N11092);
xor XOR2 (N11103, N11099, N1016);
nor NOR4 (N11104, N11103, N83, N2945, N10213);
nand NAND3 (N11105, N11100, N3440, N2377);
and AND3 (N11106, N11095, N5568, N3629);
buf BUF1 (N11107, N11106);
nand NAND4 (N11108, N11102, N9315, N634, N7958);
and AND2 (N11109, N11105, N1385);
xor XOR2 (N11110, N11109, N9715);
xor XOR2 (N11111, N11101, N5717);
nand NAND4 (N11112, N11091, N3536, N6467, N7852);
not NOT1 (N11113, N11112);
and AND3 (N11114, N11108, N3662, N1685);
not NOT1 (N11115, N11086);
xor XOR2 (N11116, N11098, N10133);
nor NOR2 (N11117, N11113, N8437);
xor XOR2 (N11118, N11116, N3117);
and AND3 (N11119, N11118, N3735, N9314);
nand NAND2 (N11120, N11104, N11045);
and AND2 (N11121, N11114, N5066);
xor XOR2 (N11122, N11094, N5348);
or OR3 (N11123, N11120, N3046, N5137);
nor NOR2 (N11124, N11122, N3322);
or OR4 (N11125, N11124, N3455, N1483, N8983);
buf BUF1 (N11126, N11085);
nand NAND2 (N11127, N11119, N11124);
nand NAND3 (N11128, N11125, N2649, N2049);
or OR4 (N11129, N11107, N8057, N1221, N1304);
and AND3 (N11130, N11129, N3792, N6217);
xor XOR2 (N11131, N11121, N4434);
buf BUF1 (N11132, N11123);
and AND3 (N11133, N11131, N7257, N3513);
nor NOR2 (N11134, N11111, N350);
nor NOR3 (N11135, N11134, N10647, N10369);
not NOT1 (N11136, N11117);
nor NOR4 (N11137, N11115, N3741, N4127, N6377);
not NOT1 (N11138, N11128);
xor XOR2 (N11139, N11133, N409);
and AND3 (N11140, N11136, N8518, N6144);
nor NOR3 (N11141, N11138, N2901, N8343);
not NOT1 (N11142, N11130);
and AND3 (N11143, N11137, N3335, N7745);
and AND2 (N11144, N11132, N8998);
or OR3 (N11145, N11144, N188, N9517);
not NOT1 (N11146, N11139);
not NOT1 (N11147, N11143);
or OR4 (N11148, N11126, N5991, N6085, N7353);
nor NOR3 (N11149, N11127, N10043, N4059);
nand NAND3 (N11150, N11141, N8392, N7793);
nand NAND4 (N11151, N11147, N3760, N7364, N5184);
nand NAND3 (N11152, N11145, N5332, N2372);
nor NOR2 (N11153, N11148, N1900);
nor NOR2 (N11154, N11149, N1690);
nor NOR3 (N11155, N11146, N7345, N9686);
not NOT1 (N11156, N11135);
and AND2 (N11157, N11152, N2298);
and AND2 (N11158, N11142, N6192);
or OR2 (N11159, N11150, N9823);
buf BUF1 (N11160, N11155);
xor XOR2 (N11161, N11140, N9262);
not NOT1 (N11162, N11159);
buf BUF1 (N11163, N11153);
and AND4 (N11164, N11151, N6123, N8833, N4367);
or OR4 (N11165, N11161, N7545, N10759, N3548);
nand NAND3 (N11166, N11157, N8262, N7848);
not NOT1 (N11167, N11158);
buf BUF1 (N11168, N11154);
and AND3 (N11169, N11168, N2236, N4474);
nand NAND3 (N11170, N11160, N732, N7225);
nand NAND4 (N11171, N11165, N9803, N4621, N9811);
buf BUF1 (N11172, N11170);
xor XOR2 (N11173, N11163, N9333);
nand NAND3 (N11174, N11156, N5324, N6346);
xor XOR2 (N11175, N11110, N5522);
xor XOR2 (N11176, N11162, N8107);
nand NAND2 (N11177, N11169, N5108);
xor XOR2 (N11178, N11167, N915);
nand NAND2 (N11179, N11176, N3366);
not NOT1 (N11180, N11171);
or OR2 (N11181, N11173, N5511);
or OR3 (N11182, N11175, N772, N2411);
nand NAND2 (N11183, N11178, N5580);
or OR4 (N11184, N11177, N9132, N885, N593);
or OR4 (N11185, N11166, N8844, N1119, N5740);
nand NAND3 (N11186, N11174, N6695, N6097);
and AND4 (N11187, N11182, N2200, N6508, N1417);
nor NOR4 (N11188, N11185, N5080, N7684, N10230);
and AND3 (N11189, N11164, N10984, N9705);
nand NAND2 (N11190, N11188, N3742);
buf BUF1 (N11191, N11184);
or OR2 (N11192, N11172, N11164);
nor NOR3 (N11193, N11189, N8263, N3465);
not NOT1 (N11194, N11183);
not NOT1 (N11195, N11180);
or OR3 (N11196, N11194, N4959, N7073);
buf BUF1 (N11197, N11179);
or OR3 (N11198, N11193, N4738, N29);
not NOT1 (N11199, N11192);
nor NOR2 (N11200, N11190, N5967);
or OR3 (N11201, N11181, N6386, N1804);
xor XOR2 (N11202, N11186, N5704);
nand NAND2 (N11203, N11195, N10848);
xor XOR2 (N11204, N11199, N473);
buf BUF1 (N11205, N11203);
and AND4 (N11206, N11200, N9762, N9670, N6627);
xor XOR2 (N11207, N11191, N1655);
and AND3 (N11208, N11197, N6510, N6247);
xor XOR2 (N11209, N11196, N8164);
buf BUF1 (N11210, N11207);
or OR3 (N11211, N11201, N3738, N10676);
buf BUF1 (N11212, N11211);
nor NOR3 (N11213, N11187, N2819, N6481);
or OR2 (N11214, N11206, N7733);
or OR4 (N11215, N11204, N10978, N1855, N3113);
not NOT1 (N11216, N11198);
not NOT1 (N11217, N11215);
and AND4 (N11218, N11208, N11002, N5118, N187);
and AND3 (N11219, N11202, N3560, N4786);
buf BUF1 (N11220, N11210);
xor XOR2 (N11221, N11205, N10077);
and AND4 (N11222, N11217, N8865, N11023, N8493);
or OR2 (N11223, N11214, N802);
and AND4 (N11224, N11221, N8750, N1782, N4851);
not NOT1 (N11225, N11209);
or OR4 (N11226, N11218, N5082, N1616, N5959);
xor XOR2 (N11227, N11225, N5794);
and AND2 (N11228, N11223, N6981);
not NOT1 (N11229, N11228);
and AND4 (N11230, N11222, N10512, N11060, N8936);
or OR4 (N11231, N11220, N7132, N6665, N7783);
or OR2 (N11232, N11216, N4772);
nor NOR4 (N11233, N11219, N9663, N8096, N7802);
buf BUF1 (N11234, N11231);
buf BUF1 (N11235, N11224);
not NOT1 (N11236, N11213);
and AND4 (N11237, N11212, N6768, N1556, N1096);
xor XOR2 (N11238, N11226, N7899);
not NOT1 (N11239, N11230);
nor NOR2 (N11240, N11233, N7263);
nand NAND2 (N11241, N11235, N5745);
or OR2 (N11242, N11234, N4540);
xor XOR2 (N11243, N11242, N4417);
not NOT1 (N11244, N11238);
xor XOR2 (N11245, N11236, N9448);
xor XOR2 (N11246, N11237, N9891);
xor XOR2 (N11247, N11246, N5932);
not NOT1 (N11248, N11227);
buf BUF1 (N11249, N11243);
nor NOR4 (N11250, N11249, N1740, N4968, N1655);
buf BUF1 (N11251, N11247);
not NOT1 (N11252, N11245);
xor XOR2 (N11253, N11252, N2440);
and AND4 (N11254, N11232, N879, N284, N6620);
or OR2 (N11255, N11250, N8502);
and AND3 (N11256, N11239, N9424, N10301);
nor NOR2 (N11257, N11255, N10898);
buf BUF1 (N11258, N11253);
xor XOR2 (N11259, N11240, N228);
nand NAND2 (N11260, N11259, N8961);
xor XOR2 (N11261, N11260, N2109);
not NOT1 (N11262, N11254);
nor NOR2 (N11263, N11248, N2711);
nand NAND4 (N11264, N11257, N9107, N10374, N3425);
not NOT1 (N11265, N11258);
xor XOR2 (N11266, N11262, N9457);
not NOT1 (N11267, N11264);
not NOT1 (N11268, N11263);
nand NAND2 (N11269, N11268, N4652);
nand NAND2 (N11270, N11229, N5939);
nand NAND2 (N11271, N11241, N801);
xor XOR2 (N11272, N11261, N7381);
or OR4 (N11273, N11271, N8043, N6322, N8816);
nor NOR2 (N11274, N11256, N9614);
nand NAND4 (N11275, N11269, N410, N574, N4505);
nand NAND4 (N11276, N11270, N4467, N1460, N2964);
buf BUF1 (N11277, N11275);
and AND2 (N11278, N11251, N3148);
nor NOR2 (N11279, N11244, N9232);
and AND2 (N11280, N11279, N5181);
not NOT1 (N11281, N11277);
and AND4 (N11282, N11274, N1125, N9140, N6137);
not NOT1 (N11283, N11273);
and AND3 (N11284, N11282, N878, N6948);
nor NOR4 (N11285, N11266, N5064, N8305, N7471);
and AND3 (N11286, N11265, N5270, N11270);
buf BUF1 (N11287, N11285);
nor NOR3 (N11288, N11276, N155, N2816);
not NOT1 (N11289, N11288);
and AND4 (N11290, N11278, N7288, N5214, N9085);
and AND4 (N11291, N11286, N3534, N7993, N2412);
or OR2 (N11292, N11290, N11115);
xor XOR2 (N11293, N11284, N4892);
or OR3 (N11294, N11291, N2835, N2477);
not NOT1 (N11295, N11283);
not NOT1 (N11296, N11272);
xor XOR2 (N11297, N11267, N5790);
not NOT1 (N11298, N11294);
nor NOR3 (N11299, N11289, N5563, N9717);
buf BUF1 (N11300, N11280);
nand NAND4 (N11301, N11299, N9115, N10795, N3115);
nand NAND2 (N11302, N11300, N669);
xor XOR2 (N11303, N11297, N6207);
and AND4 (N11304, N11281, N2444, N1108, N7268);
or OR3 (N11305, N11296, N2200, N10003);
nor NOR3 (N11306, N11292, N524, N4992);
nand NAND3 (N11307, N11304, N8123, N4115);
or OR4 (N11308, N11302, N9265, N7312, N10881);
nor NOR2 (N11309, N11307, N2571);
and AND2 (N11310, N11309, N8403);
buf BUF1 (N11311, N11303);
xor XOR2 (N11312, N11293, N1493);
and AND3 (N11313, N11287, N4259, N9428);
nand NAND4 (N11314, N11305, N10838, N10364, N6103);
not NOT1 (N11315, N11298);
and AND4 (N11316, N11313, N9046, N5228, N2099);
not NOT1 (N11317, N11306);
nand NAND2 (N11318, N11310, N1738);
or OR3 (N11319, N11317, N1591, N4615);
nand NAND3 (N11320, N11319, N7006, N7511);
nand NAND3 (N11321, N11295, N2261, N881);
and AND4 (N11322, N11321, N4015, N10306, N8300);
or OR3 (N11323, N11315, N421, N8918);
and AND2 (N11324, N11318, N1331);
buf BUF1 (N11325, N11314);
or OR3 (N11326, N11325, N7098, N6881);
and AND4 (N11327, N11326, N5583, N2989, N3047);
xor XOR2 (N11328, N11311, N7204);
or OR3 (N11329, N11327, N2977, N5212);
and AND2 (N11330, N11323, N5400);
not NOT1 (N11331, N11322);
nand NAND2 (N11332, N11330, N2581);
and AND4 (N11333, N11328, N3224, N6744, N5365);
or OR4 (N11334, N11329, N5124, N10416, N10598);
nand NAND4 (N11335, N11320, N860, N4957, N9195);
not NOT1 (N11336, N11324);
nand NAND3 (N11337, N11332, N8765, N7709);
and AND4 (N11338, N11337, N6751, N10337, N2998);
nand NAND3 (N11339, N11335, N2725, N4569);
nand NAND3 (N11340, N11336, N9680, N5415);
and AND4 (N11341, N11339, N1338, N2773, N782);
nand NAND4 (N11342, N11308, N1096, N4951, N926);
nor NOR4 (N11343, N11312, N70, N4263, N3687);
nand NAND4 (N11344, N11333, N7691, N933, N8870);
nor NOR3 (N11345, N11301, N3028, N4864);
nand NAND4 (N11346, N11342, N9895, N4924, N6789);
buf BUF1 (N11347, N11338);
buf BUF1 (N11348, N11331);
or OR2 (N11349, N11343, N1507);
xor XOR2 (N11350, N11345, N2718);
nor NOR4 (N11351, N11350, N8334, N9092, N5781);
or OR2 (N11352, N11351, N10681);
buf BUF1 (N11353, N11341);
and AND4 (N11354, N11340, N7415, N11167, N9909);
or OR2 (N11355, N11316, N1951);
xor XOR2 (N11356, N11352, N2924);
or OR4 (N11357, N11344, N7769, N464, N8449);
xor XOR2 (N11358, N11334, N3137);
and AND4 (N11359, N11357, N8581, N10257, N8898);
xor XOR2 (N11360, N11348, N10388);
xor XOR2 (N11361, N11360, N6137);
buf BUF1 (N11362, N11358);
nor NOR3 (N11363, N11347, N6144, N6145);
xor XOR2 (N11364, N11353, N572);
and AND3 (N11365, N11354, N7631, N7647);
nand NAND4 (N11366, N11362, N2919, N5453, N5838);
buf BUF1 (N11367, N11366);
and AND2 (N11368, N11356, N9865);
and AND4 (N11369, N11346, N523, N9788, N4601);
or OR3 (N11370, N11368, N102, N10304);
buf BUF1 (N11371, N11369);
nand NAND4 (N11372, N11359, N9694, N1012, N3047);
or OR3 (N11373, N11361, N4660, N7422);
nor NOR4 (N11374, N11364, N8240, N9501, N3314);
and AND2 (N11375, N11374, N9253);
buf BUF1 (N11376, N11363);
buf BUF1 (N11377, N11355);
buf BUF1 (N11378, N11370);
nand NAND4 (N11379, N11378, N1021, N3468, N6428);
nor NOR2 (N11380, N11372, N9798);
or OR4 (N11381, N11379, N5116, N5123, N8517);
not NOT1 (N11382, N11371);
not NOT1 (N11383, N11377);
buf BUF1 (N11384, N11383);
not NOT1 (N11385, N11380);
buf BUF1 (N11386, N11376);
and AND2 (N11387, N11382, N1580);
xor XOR2 (N11388, N11381, N1559);
or OR4 (N11389, N11384, N2517, N117, N9385);
xor XOR2 (N11390, N11373, N8964);
nand NAND2 (N11391, N11385, N9039);
and AND3 (N11392, N11387, N10444, N2747);
nand NAND2 (N11393, N11390, N7284);
buf BUF1 (N11394, N11349);
not NOT1 (N11395, N11392);
and AND4 (N11396, N11395, N1815, N7092, N2420);
nor NOR4 (N11397, N11391, N10325, N5129, N10654);
or OR4 (N11398, N11396, N8506, N11133, N7345);
nor NOR2 (N11399, N11397, N1912);
nor NOR4 (N11400, N11399, N8189, N841, N946);
buf BUF1 (N11401, N11375);
or OR3 (N11402, N11398, N8491, N977);
nand NAND3 (N11403, N11400, N954, N10342);
and AND3 (N11404, N11403, N4456, N9014);
or OR2 (N11405, N11404, N4237);
nor NOR3 (N11406, N11365, N6363, N1177);
or OR2 (N11407, N11367, N7703);
nor NOR3 (N11408, N11407, N3513, N8633);
and AND3 (N11409, N11389, N3504, N4997);
nor NOR4 (N11410, N11406, N3865, N10034, N2426);
xor XOR2 (N11411, N11401, N7740);
xor XOR2 (N11412, N11405, N11068);
nor NOR4 (N11413, N11394, N2501, N407, N10804);
and AND4 (N11414, N11412, N892, N4799, N126);
buf BUF1 (N11415, N11408);
buf BUF1 (N11416, N11386);
or OR2 (N11417, N11413, N3255);
and AND4 (N11418, N11411, N2862, N6047, N2559);
nor NOR2 (N11419, N11388, N10918);
buf BUF1 (N11420, N11414);
nor NOR2 (N11421, N11417, N1103);
not NOT1 (N11422, N11421);
not NOT1 (N11423, N11393);
nand NAND3 (N11424, N11418, N5688, N4323);
not NOT1 (N11425, N11420);
xor XOR2 (N11426, N11419, N5837);
buf BUF1 (N11427, N11402);
and AND3 (N11428, N11425, N3699, N3031);
xor XOR2 (N11429, N11428, N7476);
not NOT1 (N11430, N11422);
nand NAND2 (N11431, N11426, N5651);
or OR4 (N11432, N11415, N5305, N2659, N3833);
nand NAND3 (N11433, N11424, N10130, N121);
or OR3 (N11434, N11429, N3471, N590);
not NOT1 (N11435, N11434);
or OR3 (N11436, N11432, N5636, N8992);
buf BUF1 (N11437, N11427);
and AND2 (N11438, N11433, N8722);
nor NOR2 (N11439, N11410, N6960);
not NOT1 (N11440, N11430);
and AND4 (N11441, N11436, N6616, N7937, N2407);
nand NAND3 (N11442, N11423, N6910, N9622);
not NOT1 (N11443, N11442);
buf BUF1 (N11444, N11440);
not NOT1 (N11445, N11444);
not NOT1 (N11446, N11409);
or OR3 (N11447, N11416, N10723, N31);
nor NOR3 (N11448, N11431, N8854, N6358);
not NOT1 (N11449, N11448);
and AND4 (N11450, N11445, N761, N9962, N1349);
or OR3 (N11451, N11447, N9340, N9238);
buf BUF1 (N11452, N11435);
or OR4 (N11453, N11446, N816, N6435, N10281);
buf BUF1 (N11454, N11452);
xor XOR2 (N11455, N11450, N5232);
nor NOR2 (N11456, N11437, N8690);
or OR3 (N11457, N11449, N141, N9002);
or OR4 (N11458, N11439, N4270, N4454, N4219);
or OR2 (N11459, N11456, N4332);
xor XOR2 (N11460, N11455, N7149);
buf BUF1 (N11461, N11458);
or OR2 (N11462, N11454, N136);
nand NAND2 (N11463, N11451, N1824);
or OR2 (N11464, N11441, N1685);
nand NAND4 (N11465, N11453, N1279, N11132, N11034);
nand NAND3 (N11466, N11464, N6890, N11425);
and AND2 (N11467, N11463, N10027);
nand NAND3 (N11468, N11466, N4637, N3799);
nor NOR3 (N11469, N11461, N11156, N871);
nand NAND3 (N11470, N11460, N6456, N8186);
and AND3 (N11471, N11443, N1284, N1321);
or OR2 (N11472, N11470, N9696);
xor XOR2 (N11473, N11468, N7937);
or OR2 (N11474, N11462, N8113);
nor NOR3 (N11475, N11469, N3888, N11120);
nand NAND2 (N11476, N11475, N7037);
xor XOR2 (N11477, N11472, N6547);
or OR2 (N11478, N11474, N3635);
buf BUF1 (N11479, N11457);
xor XOR2 (N11480, N11471, N4203);
buf BUF1 (N11481, N11476);
nand NAND4 (N11482, N11459, N10284, N5736, N4593);
and AND4 (N11483, N11480, N994, N8722, N6799);
xor XOR2 (N11484, N11477, N8872);
nand NAND3 (N11485, N11482, N11113, N3260);
and AND2 (N11486, N11485, N3606);
nand NAND4 (N11487, N11481, N2291, N2405, N3931);
nor NOR4 (N11488, N11484, N146, N5603, N5072);
buf BUF1 (N11489, N11487);
or OR4 (N11490, N11486, N5599, N6069, N4769);
or OR3 (N11491, N11473, N3897, N3418);
and AND4 (N11492, N11478, N7720, N10637, N3461);
nand NAND3 (N11493, N11491, N10431, N7578);
nor NOR2 (N11494, N11493, N1612);
buf BUF1 (N11495, N11438);
xor XOR2 (N11496, N11488, N4488);
buf BUF1 (N11497, N11479);
nand NAND3 (N11498, N11490, N557, N10826);
xor XOR2 (N11499, N11498, N2120);
xor XOR2 (N11500, N11483, N9881);
or OR4 (N11501, N11465, N10760, N1680, N6000);
nor NOR2 (N11502, N11495, N4510);
buf BUF1 (N11503, N11501);
not NOT1 (N11504, N11500);
nor NOR2 (N11505, N11492, N9712);
buf BUF1 (N11506, N11502);
buf BUF1 (N11507, N11494);
or OR4 (N11508, N11497, N9434, N9405, N10140);
xor XOR2 (N11509, N11496, N5235);
nor NOR4 (N11510, N11505, N931, N4625, N6699);
and AND4 (N11511, N11503, N4483, N2732, N4102);
buf BUF1 (N11512, N11499);
or OR2 (N11513, N11504, N1288);
and AND3 (N11514, N11511, N7397, N6878);
xor XOR2 (N11515, N11512, N8305);
buf BUF1 (N11516, N11507);
nand NAND4 (N11517, N11489, N9213, N9903, N8707);
nor NOR4 (N11518, N11516, N8243, N1247, N9336);
nor NOR3 (N11519, N11510, N1225, N3011);
buf BUF1 (N11520, N11506);
xor XOR2 (N11521, N11519, N3679);
and AND2 (N11522, N11517, N7162);
or OR4 (N11523, N11518, N10132, N11320, N9423);
nor NOR3 (N11524, N11509, N4857, N11483);
nand NAND3 (N11525, N11467, N7539, N1090);
and AND3 (N11526, N11515, N792, N8585);
nand NAND3 (N11527, N11508, N833, N4578);
xor XOR2 (N11528, N11521, N9006);
xor XOR2 (N11529, N11524, N547);
and AND3 (N11530, N11522, N9456, N2209);
buf BUF1 (N11531, N11513);
or OR3 (N11532, N11530, N7463, N8551);
nor NOR3 (N11533, N11520, N2226, N5562);
xor XOR2 (N11534, N11523, N9420);
nor NOR4 (N11535, N11527, N6914, N3629, N3117);
or OR2 (N11536, N11535, N5373);
buf BUF1 (N11537, N11534);
xor XOR2 (N11538, N11531, N4610);
xor XOR2 (N11539, N11538, N2878);
xor XOR2 (N11540, N11537, N10250);
nand NAND2 (N11541, N11536, N2507);
nor NOR3 (N11542, N11514, N2373, N2300);
not NOT1 (N11543, N11532);
and AND4 (N11544, N11542, N11387, N6278, N3490);
or OR4 (N11545, N11541, N1933, N3633, N10589);
and AND4 (N11546, N11528, N1587, N8926, N3821);
nor NOR4 (N11547, N11533, N1101, N10591, N1650);
and AND4 (N11548, N11540, N9345, N6600, N2790);
xor XOR2 (N11549, N11525, N729);
not NOT1 (N11550, N11549);
not NOT1 (N11551, N11547);
nor NOR3 (N11552, N11548, N2346, N5875);
buf BUF1 (N11553, N11552);
nor NOR4 (N11554, N11545, N11341, N1781, N5864);
and AND3 (N11555, N11539, N2020, N5743);
not NOT1 (N11556, N11554);
not NOT1 (N11557, N11555);
buf BUF1 (N11558, N11544);
and AND4 (N11559, N11526, N3586, N2238, N10967);
or OR3 (N11560, N11556, N7407, N2820);
or OR2 (N11561, N11543, N3749);
xor XOR2 (N11562, N11546, N7398);
nor NOR3 (N11563, N11559, N3379, N4303);
nand NAND3 (N11564, N11557, N11044, N9604);
and AND3 (N11565, N11563, N7089, N11507);
or OR3 (N11566, N11561, N9788, N2456);
and AND2 (N11567, N11560, N3122);
and AND3 (N11568, N11558, N10373, N9720);
buf BUF1 (N11569, N11562);
nand NAND4 (N11570, N11566, N2511, N3239, N6830);
and AND3 (N11571, N11569, N8519, N6220);
not NOT1 (N11572, N11565);
nand NAND4 (N11573, N11550, N8405, N5661, N8743);
nand NAND4 (N11574, N11573, N3920, N10462, N8929);
nor NOR2 (N11575, N11568, N10164);
or OR3 (N11576, N11553, N1376, N7810);
and AND3 (N11577, N11575, N11269, N515);
and AND2 (N11578, N11564, N289);
xor XOR2 (N11579, N11529, N1046);
nand NAND4 (N11580, N11579, N5176, N6150, N9271);
nor NOR3 (N11581, N11571, N8603, N7643);
buf BUF1 (N11582, N11580);
xor XOR2 (N11583, N11576, N2442);
not NOT1 (N11584, N11551);
xor XOR2 (N11585, N11584, N8988);
nor NOR2 (N11586, N11567, N6400);
not NOT1 (N11587, N11572);
nand NAND4 (N11588, N11587, N5921, N8147, N7539);
not NOT1 (N11589, N11570);
xor XOR2 (N11590, N11577, N10229);
not NOT1 (N11591, N11582);
xor XOR2 (N11592, N11589, N2457);
xor XOR2 (N11593, N11583, N6778);
not NOT1 (N11594, N11586);
nand NAND4 (N11595, N11588, N3157, N4290, N5180);
nand NAND4 (N11596, N11593, N9055, N3077, N7841);
and AND4 (N11597, N11592, N3135, N7054, N7590);
or OR3 (N11598, N11595, N5517, N84);
nand NAND3 (N11599, N11591, N8765, N10817);
or OR4 (N11600, N11581, N10458, N11263, N5979);
xor XOR2 (N11601, N11596, N2900);
nor NOR2 (N11602, N11585, N8101);
not NOT1 (N11603, N11597);
or OR2 (N11604, N11594, N7314);
nor NOR3 (N11605, N11578, N6684, N766);
nor NOR2 (N11606, N11598, N8645);
or OR3 (N11607, N11574, N9510, N5570);
nor NOR3 (N11608, N11605, N5548, N3963);
and AND3 (N11609, N11600, N7120, N6202);
nand NAND3 (N11610, N11609, N8975, N4260);
and AND3 (N11611, N11604, N6489, N4756);
xor XOR2 (N11612, N11611, N3417);
nor NOR3 (N11613, N11601, N7134, N6266);
and AND3 (N11614, N11612, N1295, N10479);
xor XOR2 (N11615, N11603, N8918);
buf BUF1 (N11616, N11615);
xor XOR2 (N11617, N11613, N10736);
buf BUF1 (N11618, N11616);
nand NAND2 (N11619, N11608, N7373);
nand NAND4 (N11620, N11602, N3561, N1011, N10384);
nand NAND4 (N11621, N11620, N5910, N2390, N10150);
nand NAND4 (N11622, N11607, N7070, N10176, N11124);
nand NAND3 (N11623, N11590, N2576, N4311);
nand NAND4 (N11624, N11614, N9780, N822, N8202);
and AND3 (N11625, N11617, N9940, N1723);
buf BUF1 (N11626, N11625);
buf BUF1 (N11627, N11619);
buf BUF1 (N11628, N11626);
buf BUF1 (N11629, N11624);
or OR2 (N11630, N11628, N3474);
nor NOR3 (N11631, N11599, N1159, N7791);
buf BUF1 (N11632, N11621);
nand NAND2 (N11633, N11631, N11372);
buf BUF1 (N11634, N11610);
nor NOR3 (N11635, N11633, N8590, N2196);
nor NOR2 (N11636, N11630, N2096);
buf BUF1 (N11637, N11636);
or OR3 (N11638, N11635, N130, N5445);
buf BUF1 (N11639, N11637);
buf BUF1 (N11640, N11639);
not NOT1 (N11641, N11627);
not NOT1 (N11642, N11606);
not NOT1 (N11643, N11638);
and AND3 (N11644, N11623, N5673, N8675);
buf BUF1 (N11645, N11622);
nand NAND3 (N11646, N11642, N9763, N4904);
and AND3 (N11647, N11634, N2301, N8346);
nor NOR2 (N11648, N11643, N961);
buf BUF1 (N11649, N11645);
xor XOR2 (N11650, N11648, N11488);
nand NAND3 (N11651, N11650, N5114, N5441);
and AND4 (N11652, N11641, N8287, N11164, N10711);
nand NAND3 (N11653, N11640, N3549, N3657);
nor NOR4 (N11654, N11618, N3446, N10369, N9214);
nand NAND4 (N11655, N11651, N11333, N1435, N3085);
or OR2 (N11656, N11649, N7256);
nand NAND2 (N11657, N11644, N9914);
or OR4 (N11658, N11653, N2944, N4369, N2194);
and AND2 (N11659, N11647, N1085);
buf BUF1 (N11660, N11632);
xor XOR2 (N11661, N11652, N367);
not NOT1 (N11662, N11656);
nand NAND4 (N11663, N11659, N8789, N9940, N6323);
nor NOR4 (N11664, N11646, N5507, N3874, N6520);
and AND2 (N11665, N11663, N1849);
nor NOR2 (N11666, N11662, N575);
nand NAND4 (N11667, N11666, N8286, N10706, N5678);
buf BUF1 (N11668, N11654);
xor XOR2 (N11669, N11629, N11422);
buf BUF1 (N11670, N11661);
buf BUF1 (N11671, N11658);
xor XOR2 (N11672, N11660, N11027);
nor NOR2 (N11673, N11665, N2639);
not NOT1 (N11674, N11657);
nor NOR3 (N11675, N11667, N4809, N9944);
xor XOR2 (N11676, N11675, N10427);
not NOT1 (N11677, N11676);
not NOT1 (N11678, N11669);
buf BUF1 (N11679, N11655);
nor NOR2 (N11680, N11677, N4438);
nand NAND4 (N11681, N11671, N298, N4272, N7183);
or OR2 (N11682, N11668, N8769);
or OR3 (N11683, N11670, N3971, N6972);
nand NAND2 (N11684, N11679, N5449);
xor XOR2 (N11685, N11678, N163);
xor XOR2 (N11686, N11682, N1701);
and AND2 (N11687, N11686, N8741);
not NOT1 (N11688, N11674);
and AND2 (N11689, N11680, N6147);
xor XOR2 (N11690, N11664, N3426);
buf BUF1 (N11691, N11687);
nor NOR3 (N11692, N11685, N3585, N4073);
buf BUF1 (N11693, N11689);
or OR4 (N11694, N11693, N5283, N1831, N1967);
xor XOR2 (N11695, N11683, N9917);
buf BUF1 (N11696, N11673);
nor NOR4 (N11697, N11692, N11013, N2368, N10506);
not NOT1 (N11698, N11672);
not NOT1 (N11699, N11694);
not NOT1 (N11700, N11697);
xor XOR2 (N11701, N11688, N9474);
and AND4 (N11702, N11700, N105, N11521, N4717);
nand NAND2 (N11703, N11698, N6852);
not NOT1 (N11704, N11681);
nor NOR2 (N11705, N11703, N9905);
and AND3 (N11706, N11699, N4592, N8309);
buf BUF1 (N11707, N11690);
nor NOR4 (N11708, N11706, N2067, N2760, N151);
or OR3 (N11709, N11691, N3441, N6732);
nand NAND3 (N11710, N11701, N2068, N9801);
buf BUF1 (N11711, N11702);
nand NAND4 (N11712, N11704, N1321, N5497, N9371);
or OR2 (N11713, N11707, N10788);
buf BUF1 (N11714, N11708);
and AND4 (N11715, N11714, N9406, N10613, N1519);
or OR4 (N11716, N11715, N11414, N10383, N9889);
not NOT1 (N11717, N11716);
not NOT1 (N11718, N11705);
xor XOR2 (N11719, N11712, N2260);
and AND2 (N11720, N11696, N11105);
or OR3 (N11721, N11709, N145, N7392);
and AND3 (N11722, N11695, N10653, N1424);
buf BUF1 (N11723, N11720);
buf BUF1 (N11724, N11684);
nand NAND4 (N11725, N11718, N36, N6178, N11561);
or OR4 (N11726, N11717, N6715, N675, N2080);
nor NOR4 (N11727, N11713, N2693, N10447, N2372);
buf BUF1 (N11728, N11723);
xor XOR2 (N11729, N11726, N9585);
buf BUF1 (N11730, N11719);
nand NAND4 (N11731, N11724, N4746, N1923, N4969);
or OR4 (N11732, N11727, N11361, N6661, N9963);
buf BUF1 (N11733, N11711);
nand NAND3 (N11734, N11725, N11703, N1587);
nand NAND2 (N11735, N11721, N11193);
xor XOR2 (N11736, N11732, N8136);
not NOT1 (N11737, N11736);
nand NAND2 (N11738, N11733, N9299);
xor XOR2 (N11739, N11734, N3059);
buf BUF1 (N11740, N11731);
not NOT1 (N11741, N11730);
xor XOR2 (N11742, N11738, N1039);
or OR4 (N11743, N11742, N8734, N2536, N3000);
nand NAND4 (N11744, N11741, N11615, N8833, N4436);
xor XOR2 (N11745, N11710, N3674);
xor XOR2 (N11746, N11744, N8401);
xor XOR2 (N11747, N11728, N6362);
nor NOR4 (N11748, N11745, N4716, N953, N3033);
not NOT1 (N11749, N11748);
and AND2 (N11750, N11737, N1081);
buf BUF1 (N11751, N11722);
nand NAND2 (N11752, N11729, N6880);
nor NOR4 (N11753, N11743, N4516, N8736, N4598);
and AND3 (N11754, N11753, N6282, N9986);
nand NAND2 (N11755, N11739, N10020);
xor XOR2 (N11756, N11754, N669);
not NOT1 (N11757, N11755);
buf BUF1 (N11758, N11749);
nor NOR4 (N11759, N11757, N2482, N896, N11557);
nand NAND3 (N11760, N11747, N5365, N7583);
not NOT1 (N11761, N11740);
and AND2 (N11762, N11761, N1282);
buf BUF1 (N11763, N11751);
or OR3 (N11764, N11760, N9844, N7444);
and AND3 (N11765, N11735, N11202, N9103);
nand NAND3 (N11766, N11764, N54, N6830);
nand NAND2 (N11767, N11746, N9670);
and AND2 (N11768, N11762, N11711);
buf BUF1 (N11769, N11768);
xor XOR2 (N11770, N11763, N6517);
or OR3 (N11771, N11758, N4290, N10485);
and AND4 (N11772, N11750, N2365, N3088, N4800);
nand NAND3 (N11773, N11756, N8470, N6965);
or OR4 (N11774, N11752, N4838, N5359, N216);
or OR3 (N11775, N11770, N9458, N2907);
nand NAND3 (N11776, N11772, N2993, N8175);
nand NAND3 (N11777, N11769, N5309, N4095);
or OR4 (N11778, N11776, N3475, N848, N6954);
not NOT1 (N11779, N11778);
xor XOR2 (N11780, N11759, N3152);
or OR4 (N11781, N11767, N4788, N11444, N5907);
and AND3 (N11782, N11766, N1700, N4302);
xor XOR2 (N11783, N11774, N6918);
nor NOR4 (N11784, N11777, N1654, N402, N178);
not NOT1 (N11785, N11783);
or OR3 (N11786, N11780, N9302, N5987);
xor XOR2 (N11787, N11782, N10866);
xor XOR2 (N11788, N11786, N8954);
nor NOR2 (N11789, N11788, N1817);
nand NAND2 (N11790, N11787, N441);
and AND4 (N11791, N11775, N4440, N4255, N2395);
nor NOR4 (N11792, N11771, N10738, N2128, N10934);
not NOT1 (N11793, N11765);
not NOT1 (N11794, N11773);
nand NAND4 (N11795, N11785, N9467, N10546, N6405);
or OR3 (N11796, N11795, N2836, N7249);
xor XOR2 (N11797, N11790, N771);
and AND3 (N11798, N11797, N9918, N3347);
nor NOR3 (N11799, N11779, N1798, N11324);
nor NOR3 (N11800, N11799, N9750, N8729);
not NOT1 (N11801, N11791);
or OR2 (N11802, N11796, N10882);
and AND3 (N11803, N11798, N2077, N8150);
or OR3 (N11804, N11789, N11782, N5295);
and AND4 (N11805, N11803, N8060, N5396, N2372);
and AND4 (N11806, N11802, N6788, N6015, N5729);
and AND3 (N11807, N11781, N8209, N8960);
buf BUF1 (N11808, N11805);
buf BUF1 (N11809, N11807);
or OR4 (N11810, N11794, N46, N705, N10568);
nor NOR4 (N11811, N11808, N701, N3886, N8826);
or OR3 (N11812, N11784, N9922, N7777);
not NOT1 (N11813, N11793);
and AND2 (N11814, N11800, N9981);
xor XOR2 (N11815, N11801, N2545);
and AND3 (N11816, N11792, N7717, N11437);
not NOT1 (N11817, N11815);
buf BUF1 (N11818, N11812);
buf BUF1 (N11819, N11810);
nor NOR2 (N11820, N11818, N5064);
or OR4 (N11821, N11809, N5807, N8117, N1897);
nand NAND4 (N11822, N11804, N10200, N9423, N3667);
buf BUF1 (N11823, N11816);
or OR3 (N11824, N11813, N4167, N6667);
not NOT1 (N11825, N11823);
and AND4 (N11826, N11811, N8192, N3439, N5171);
or OR2 (N11827, N11814, N2614);
and AND3 (N11828, N11821, N256, N5114);
xor XOR2 (N11829, N11806, N10592);
not NOT1 (N11830, N11827);
buf BUF1 (N11831, N11822);
buf BUF1 (N11832, N11824);
nor NOR4 (N11833, N11825, N5013, N11445, N10383);
and AND4 (N11834, N11826, N6224, N227, N820);
and AND2 (N11835, N11820, N4320);
buf BUF1 (N11836, N11828);
not NOT1 (N11837, N11829);
and AND2 (N11838, N11835, N10706);
xor XOR2 (N11839, N11830, N5928);
nor NOR3 (N11840, N11832, N1654, N10710);
and AND3 (N11841, N11834, N6587, N7634);
nand NAND3 (N11842, N11831, N1017, N5072);
nor NOR4 (N11843, N11840, N6218, N2304, N11061);
nor NOR4 (N11844, N11819, N6388, N8272, N10579);
nor NOR2 (N11845, N11817, N418);
nor NOR4 (N11846, N11839, N4516, N5188, N1857);
not NOT1 (N11847, N11845);
and AND3 (N11848, N11842, N11703, N11113);
nor NOR4 (N11849, N11844, N7365, N5458, N151);
nor NOR3 (N11850, N11848, N2784, N4039);
buf BUF1 (N11851, N11838);
nand NAND4 (N11852, N11846, N4678, N3797, N6425);
and AND2 (N11853, N11837, N2539);
or OR3 (N11854, N11841, N1141, N9248);
buf BUF1 (N11855, N11850);
and AND4 (N11856, N11855, N8129, N7819, N10542);
and AND2 (N11857, N11843, N7324);
xor XOR2 (N11858, N11856, N6065);
and AND4 (N11859, N11853, N4393, N8387, N5810);
or OR2 (N11860, N11849, N11598);
xor XOR2 (N11861, N11833, N9568);
nand NAND2 (N11862, N11854, N8149);
not NOT1 (N11863, N11836);
buf BUF1 (N11864, N11863);
and AND2 (N11865, N11862, N11816);
buf BUF1 (N11866, N11857);
or OR4 (N11867, N11864, N3422, N178, N9391);
nor NOR4 (N11868, N11861, N11775, N9247, N1972);
not NOT1 (N11869, N11867);
nor NOR3 (N11870, N11865, N11550, N679);
nand NAND4 (N11871, N11860, N4333, N6531, N2604);
buf BUF1 (N11872, N11858);
nand NAND2 (N11873, N11852, N6535);
buf BUF1 (N11874, N11847);
nand NAND2 (N11875, N11871, N1266);
buf BUF1 (N11876, N11866);
nor NOR3 (N11877, N11851, N4952, N2851);
not NOT1 (N11878, N11869);
xor XOR2 (N11879, N11868, N8726);
or OR2 (N11880, N11873, N10728);
not NOT1 (N11881, N11875);
xor XOR2 (N11882, N11881, N8230);
xor XOR2 (N11883, N11879, N2178);
xor XOR2 (N11884, N11883, N181);
not NOT1 (N11885, N11884);
and AND3 (N11886, N11880, N10384, N1984);
and AND2 (N11887, N11859, N11201);
not NOT1 (N11888, N11886);
not NOT1 (N11889, N11872);
xor XOR2 (N11890, N11882, N1524);
buf BUF1 (N11891, N11885);
nand NAND4 (N11892, N11887, N1756, N5817, N3253);
nor NOR3 (N11893, N11891, N8241, N4856);
and AND2 (N11894, N11893, N8791);
nand NAND2 (N11895, N11878, N6667);
xor XOR2 (N11896, N11870, N2032);
and AND3 (N11897, N11890, N4652, N4915);
xor XOR2 (N11898, N11874, N6414);
nor NOR2 (N11899, N11897, N11601);
buf BUF1 (N11900, N11889);
or OR3 (N11901, N11899, N877, N8109);
not NOT1 (N11902, N11898);
and AND2 (N11903, N11876, N7281);
nor NOR2 (N11904, N11901, N11252);
nor NOR2 (N11905, N11903, N4575);
and AND2 (N11906, N11896, N8323);
buf BUF1 (N11907, N11906);
nor NOR2 (N11908, N11900, N9857);
xor XOR2 (N11909, N11905, N11720);
nand NAND4 (N11910, N11888, N4617, N8791, N11324);
buf BUF1 (N11911, N11902);
buf BUF1 (N11912, N11910);
nor NOR3 (N11913, N11907, N4794, N11777);
nand NAND3 (N11914, N11909, N4030, N5667);
nor NOR2 (N11915, N11913, N11742);
not NOT1 (N11916, N11912);
and AND3 (N11917, N11892, N8706, N6682);
nor NOR2 (N11918, N11877, N8723);
nand NAND3 (N11919, N11894, N4091, N8499);
nor NOR4 (N11920, N11915, N7716, N5305, N8108);
and AND3 (N11921, N11917, N5746, N7974);
not NOT1 (N11922, N11921);
and AND3 (N11923, N11914, N11324, N737);
and AND3 (N11924, N11920, N9071, N10253);
buf BUF1 (N11925, N11924);
buf BUF1 (N11926, N11908);
nand NAND4 (N11927, N11923, N7951, N519, N11497);
and AND2 (N11928, N11925, N6941);
nor NOR2 (N11929, N11926, N8507);
and AND4 (N11930, N11929, N10027, N580, N11365);
xor XOR2 (N11931, N11919, N8573);
not NOT1 (N11932, N11895);
and AND4 (N11933, N11918, N3629, N3308, N6752);
not NOT1 (N11934, N11904);
buf BUF1 (N11935, N11934);
buf BUF1 (N11936, N11922);
buf BUF1 (N11937, N11928);
xor XOR2 (N11938, N11935, N8367);
not NOT1 (N11939, N11911);
not NOT1 (N11940, N11937);
nand NAND2 (N11941, N11930, N9237);
or OR3 (N11942, N11941, N11145, N11530);
nand NAND2 (N11943, N11942, N11758);
and AND4 (N11944, N11916, N8388, N8927, N9873);
nor NOR2 (N11945, N11931, N10028);
or OR3 (N11946, N11940, N1433, N9202);
not NOT1 (N11947, N11946);
or OR4 (N11948, N11933, N11836, N8575, N6358);
and AND3 (N11949, N11943, N785, N8878);
buf BUF1 (N11950, N11932);
nor NOR3 (N11951, N11938, N7599, N5257);
nor NOR2 (N11952, N11951, N4004);
nor NOR2 (N11953, N11936, N9596);
nor NOR2 (N11954, N11947, N8589);
xor XOR2 (N11955, N11952, N5721);
xor XOR2 (N11956, N11949, N464);
nor NOR4 (N11957, N11954, N7728, N972, N8090);
not NOT1 (N11958, N11955);
nand NAND3 (N11959, N11945, N10342, N2049);
or OR2 (N11960, N11958, N1032);
and AND3 (N11961, N11948, N3019, N8375);
buf BUF1 (N11962, N11950);
or OR4 (N11963, N11962, N9057, N3416, N8106);
or OR4 (N11964, N11944, N1707, N5028, N6147);
not NOT1 (N11965, N11939);
not NOT1 (N11966, N11960);
xor XOR2 (N11967, N11965, N2325);
buf BUF1 (N11968, N11953);
nand NAND4 (N11969, N11956, N489, N4709, N11766);
nor NOR2 (N11970, N11964, N8655);
nor NOR2 (N11971, N11969, N4972);
buf BUF1 (N11972, N11927);
buf BUF1 (N11973, N11972);
buf BUF1 (N11974, N11971);
and AND3 (N11975, N11963, N7501, N3341);
xor XOR2 (N11976, N11966, N6215);
and AND3 (N11977, N11976, N2258, N6027);
or OR4 (N11978, N11961, N1558, N5837, N1867);
and AND3 (N11979, N11970, N1408, N1518);
buf BUF1 (N11980, N11979);
xor XOR2 (N11981, N11974, N3185);
buf BUF1 (N11982, N11980);
and AND2 (N11983, N11973, N10522);
nor NOR3 (N11984, N11983, N9946, N10566);
xor XOR2 (N11985, N11984, N8626);
and AND4 (N11986, N11977, N6859, N8942, N3234);
and AND2 (N11987, N11975, N8248);
nor NOR3 (N11988, N11978, N8255, N8571);
or OR3 (N11989, N11959, N7471, N6753);
nor NOR4 (N11990, N11957, N7444, N6847, N5191);
nor NOR2 (N11991, N11982, N1539);
nor NOR3 (N11992, N11986, N1547, N1015);
buf BUF1 (N11993, N11968);
xor XOR2 (N11994, N11988, N4190);
buf BUF1 (N11995, N11987);
or OR3 (N11996, N11967, N6681, N6648);
or OR4 (N11997, N11994, N8494, N1654, N1700);
nand NAND2 (N11998, N11989, N1020);
not NOT1 (N11999, N11981);
or OR2 (N12000, N11999, N11213);
not NOT1 (N12001, N11993);
not NOT1 (N12002, N11997);
not NOT1 (N12003, N12002);
not NOT1 (N12004, N12001);
and AND2 (N12005, N12003, N672);
and AND3 (N12006, N11990, N5249, N5616);
nand NAND3 (N12007, N11998, N6536, N10854);
nand NAND2 (N12008, N11992, N11781);
nor NOR3 (N12009, N12004, N8391, N6728);
and AND3 (N12010, N11995, N9953, N9964);
and AND3 (N12011, N12000, N6939, N11798);
xor XOR2 (N12012, N12008, N6991);
not NOT1 (N12013, N12010);
and AND3 (N12014, N12012, N1692, N7967);
xor XOR2 (N12015, N12009, N4577);
or OR2 (N12016, N12011, N9883);
buf BUF1 (N12017, N12005);
xor XOR2 (N12018, N12016, N7442);
or OR4 (N12019, N12017, N1813, N4163, N2568);
or OR2 (N12020, N12014, N9224);
not NOT1 (N12021, N12006);
nor NOR3 (N12022, N12021, N3590, N11762);
nand NAND2 (N12023, N12015, N2597);
nand NAND3 (N12024, N12007, N4418, N4636);
xor XOR2 (N12025, N12013, N175);
buf BUF1 (N12026, N12023);
nor NOR3 (N12027, N11991, N500, N374);
nand NAND3 (N12028, N12025, N1828, N7136);
or OR4 (N12029, N12018, N11337, N8012, N11596);
buf BUF1 (N12030, N12027);
xor XOR2 (N12031, N12024, N10928);
xor XOR2 (N12032, N11985, N25);
nand NAND4 (N12033, N12031, N5723, N9669, N7514);
nand NAND2 (N12034, N12028, N2750);
nand NAND2 (N12035, N12033, N5528);
and AND3 (N12036, N12032, N11759, N7250);
buf BUF1 (N12037, N12020);
nand NAND2 (N12038, N12029, N5350);
or OR4 (N12039, N12030, N7925, N10469, N9241);
and AND2 (N12040, N12026, N6708);
nor NOR4 (N12041, N12036, N1013, N3642, N7160);
not NOT1 (N12042, N12041);
buf BUF1 (N12043, N12022);
xor XOR2 (N12044, N12042, N9489);
nand NAND4 (N12045, N11996, N9981, N7513, N7840);
nor NOR2 (N12046, N12044, N2947);
not NOT1 (N12047, N12045);
and AND3 (N12048, N12047, N5317, N3536);
buf BUF1 (N12049, N12048);
and AND4 (N12050, N12043, N5415, N3427, N1648);
not NOT1 (N12051, N12037);
xor XOR2 (N12052, N12019, N9439);
xor XOR2 (N12053, N12052, N2372);
not NOT1 (N12054, N12039);
buf BUF1 (N12055, N12038);
nand NAND2 (N12056, N12040, N9471);
xor XOR2 (N12057, N12050, N9441);
nand NAND4 (N12058, N12054, N5827, N9018, N10763);
xor XOR2 (N12059, N12046, N8179);
or OR2 (N12060, N12034, N7797);
nand NAND2 (N12061, N12055, N2399);
nand NAND3 (N12062, N12035, N9528, N11540);
and AND2 (N12063, N12062, N10442);
not NOT1 (N12064, N12051);
and AND2 (N12065, N12056, N866);
or OR4 (N12066, N12053, N1114, N9887, N4416);
nand NAND4 (N12067, N12061, N9391, N3003, N6384);
or OR2 (N12068, N12067, N10370);
not NOT1 (N12069, N12058);
nor NOR2 (N12070, N12065, N3528);
nand NAND2 (N12071, N12059, N5047);
nand NAND2 (N12072, N12066, N6782);
nand NAND2 (N12073, N12068, N11393);
nand NAND2 (N12074, N12073, N11492);
buf BUF1 (N12075, N12057);
nor NOR2 (N12076, N12072, N1931);
and AND4 (N12077, N12064, N3149, N10370, N9704);
nor NOR2 (N12078, N12069, N1930);
xor XOR2 (N12079, N12063, N8418);
buf BUF1 (N12080, N12070);
or OR2 (N12081, N12076, N9004);
and AND3 (N12082, N12049, N1757, N8620);
not NOT1 (N12083, N12075);
xor XOR2 (N12084, N12077, N1578);
or OR4 (N12085, N12078, N10822, N8241, N8357);
or OR3 (N12086, N12074, N2007, N3126);
buf BUF1 (N12087, N12060);
nand NAND4 (N12088, N12083, N1457, N11710, N11368);
buf BUF1 (N12089, N12086);
and AND2 (N12090, N12084, N10276);
nor NOR2 (N12091, N12079, N7784);
nor NOR3 (N12092, N12085, N9615, N3753);
or OR4 (N12093, N12081, N4338, N11245, N5846);
xor XOR2 (N12094, N12093, N3381);
not NOT1 (N12095, N12080);
xor XOR2 (N12096, N12087, N4148);
or OR3 (N12097, N12090, N4534, N7213);
xor XOR2 (N12098, N12092, N7978);
xor XOR2 (N12099, N12096, N5617);
or OR4 (N12100, N12091, N9079, N8033, N6416);
buf BUF1 (N12101, N12098);
not NOT1 (N12102, N12094);
xor XOR2 (N12103, N12088, N107);
or OR3 (N12104, N12071, N3527, N5247);
buf BUF1 (N12105, N12095);
xor XOR2 (N12106, N12082, N7936);
nand NAND2 (N12107, N12104, N5238);
nor NOR3 (N12108, N12100, N10017, N6209);
and AND4 (N12109, N12097, N1634, N8791, N8092);
not NOT1 (N12110, N12106);
xor XOR2 (N12111, N12110, N2021);
nor NOR2 (N12112, N12089, N11668);
nor NOR3 (N12113, N12102, N4498, N5855);
nor NOR3 (N12114, N12105, N7651, N3554);
nand NAND3 (N12115, N12109, N1827, N11217);
or OR3 (N12116, N12108, N9281, N10543);
or OR2 (N12117, N12115, N6358);
not NOT1 (N12118, N12101);
not NOT1 (N12119, N12118);
nor NOR3 (N12120, N12113, N10493, N6768);
or OR3 (N12121, N12117, N4532, N672);
xor XOR2 (N12122, N12111, N4);
xor XOR2 (N12123, N12121, N10211);
and AND4 (N12124, N12123, N11539, N4731, N685);
and AND2 (N12125, N12107, N10110);
xor XOR2 (N12126, N12116, N4113);
buf BUF1 (N12127, N12103);
nor NOR2 (N12128, N12124, N9489);
xor XOR2 (N12129, N12127, N7962);
nor NOR2 (N12130, N12122, N6982);
buf BUF1 (N12131, N12125);
xor XOR2 (N12132, N12129, N11223);
xor XOR2 (N12133, N12099, N10707);
xor XOR2 (N12134, N12131, N7646);
or OR3 (N12135, N12128, N10954, N3666);
and AND2 (N12136, N12114, N8900);
and AND3 (N12137, N12130, N2667, N9320);
nor NOR4 (N12138, N12136, N1950, N6587, N8862);
nand NAND3 (N12139, N12132, N6925, N6185);
not NOT1 (N12140, N12120);
nor NOR4 (N12141, N12139, N1237, N194, N11906);
nor NOR3 (N12142, N12126, N10547, N10380);
nand NAND3 (N12143, N12135, N5615, N6869);
and AND2 (N12144, N12133, N2263);
buf BUF1 (N12145, N12143);
nand NAND3 (N12146, N12112, N11712, N9240);
nand NAND4 (N12147, N12138, N11367, N8127, N10869);
xor XOR2 (N12148, N12145, N11321);
or OR4 (N12149, N12148, N6824, N3916, N7546);
and AND2 (N12150, N12137, N5857);
not NOT1 (N12151, N12134);
not NOT1 (N12152, N12151);
not NOT1 (N12153, N12119);
and AND3 (N12154, N12152, N9607, N9914);
or OR2 (N12155, N12153, N10016);
not NOT1 (N12156, N12155);
buf BUF1 (N12157, N12140);
nor NOR4 (N12158, N12156, N4271, N5228, N5629);
and AND4 (N12159, N12150, N6976, N6433, N5661);
xor XOR2 (N12160, N12159, N449);
and AND2 (N12161, N12160, N3440);
not NOT1 (N12162, N12144);
not NOT1 (N12163, N12157);
or OR4 (N12164, N12162, N775, N1674, N9487);
nor NOR2 (N12165, N12163, N2100);
or OR2 (N12166, N12165, N4173);
nor NOR3 (N12167, N12142, N766, N3345);
or OR2 (N12168, N12161, N9714);
and AND2 (N12169, N12141, N5075);
or OR4 (N12170, N12164, N10691, N3933, N394);
not NOT1 (N12171, N12166);
nand NAND2 (N12172, N12167, N5698);
and AND2 (N12173, N12149, N6880);
and AND3 (N12174, N12169, N3560, N8209);
not NOT1 (N12175, N12174);
nor NOR2 (N12176, N12147, N6996);
nand NAND3 (N12177, N12175, N4892, N2584);
nor NOR2 (N12178, N12177, N9161);
not NOT1 (N12179, N12171);
buf BUF1 (N12180, N12170);
not NOT1 (N12181, N12179);
xor XOR2 (N12182, N12154, N5512);
nand NAND4 (N12183, N12158, N6406, N2738, N2236);
not NOT1 (N12184, N12172);
not NOT1 (N12185, N12184);
nor NOR2 (N12186, N12183, N8696);
nand NAND4 (N12187, N12168, N9068, N6811, N3541);
not NOT1 (N12188, N12180);
buf BUF1 (N12189, N12176);
not NOT1 (N12190, N12178);
or OR3 (N12191, N12187, N2736, N8904);
or OR4 (N12192, N12190, N8786, N6153, N4951);
not NOT1 (N12193, N12185);
xor XOR2 (N12194, N12191, N1318);
not NOT1 (N12195, N12173);
buf BUF1 (N12196, N12192);
not NOT1 (N12197, N12194);
buf BUF1 (N12198, N12186);
nand NAND2 (N12199, N12189, N5435);
nand NAND2 (N12200, N12198, N1751);
and AND2 (N12201, N12188, N9512);
not NOT1 (N12202, N12146);
or OR3 (N12203, N12199, N900, N8337);
nor NOR4 (N12204, N12200, N780, N6318, N191);
xor XOR2 (N12205, N12193, N874);
nor NOR4 (N12206, N12181, N8436, N8746, N2798);
and AND2 (N12207, N12206, N10956);
or OR2 (N12208, N12202, N1630);
nand NAND4 (N12209, N12182, N7260, N5274, N11542);
or OR2 (N12210, N12205, N8020);
not NOT1 (N12211, N12207);
and AND2 (N12212, N12209, N8791);
not NOT1 (N12213, N12196);
nor NOR4 (N12214, N12213, N1186, N6160, N2611);
buf BUF1 (N12215, N12212);
and AND4 (N12216, N12203, N9543, N11472, N9611);
or OR2 (N12217, N12195, N10395);
nand NAND2 (N12218, N12201, N2745);
and AND3 (N12219, N12211, N2331, N3215);
or OR3 (N12220, N12208, N6717, N4383);
and AND2 (N12221, N12219, N7695);
xor XOR2 (N12222, N12210, N2063);
nor NOR4 (N12223, N12216, N5284, N11463, N3367);
or OR4 (N12224, N12220, N10277, N12051, N1943);
xor XOR2 (N12225, N12221, N11682);
nand NAND3 (N12226, N12224, N3860, N3357);
buf BUF1 (N12227, N12215);
xor XOR2 (N12228, N12226, N345);
or OR4 (N12229, N12227, N9970, N2820, N10080);
nand NAND3 (N12230, N12217, N8582, N4299);
nor NOR2 (N12231, N12230, N2115);
not NOT1 (N12232, N12228);
nor NOR3 (N12233, N12223, N11090, N6102);
nor NOR3 (N12234, N12222, N6566, N8351);
or OR4 (N12235, N12204, N3792, N6028, N10819);
and AND3 (N12236, N12225, N10539, N2200);
xor XOR2 (N12237, N12231, N5233);
not NOT1 (N12238, N12197);
and AND3 (N12239, N12214, N7959, N2414);
xor XOR2 (N12240, N12237, N6106);
buf BUF1 (N12241, N12218);
nand NAND3 (N12242, N12240, N276, N10014);
and AND2 (N12243, N12239, N5728);
buf BUF1 (N12244, N12241);
and AND2 (N12245, N12244, N3105);
xor XOR2 (N12246, N12229, N1638);
nand NAND2 (N12247, N12243, N7914);
nand NAND2 (N12248, N12235, N8687);
xor XOR2 (N12249, N12247, N4446);
and AND4 (N12250, N12248, N1339, N4865, N1139);
buf BUF1 (N12251, N12246);
nor NOR3 (N12252, N12233, N8998, N10787);
nand NAND2 (N12253, N12252, N5034);
xor XOR2 (N12254, N12249, N9950);
or OR3 (N12255, N12242, N1621, N8949);
or OR2 (N12256, N12234, N8718);
nor NOR3 (N12257, N12256, N3469, N5471);
buf BUF1 (N12258, N12250);
buf BUF1 (N12259, N12232);
not NOT1 (N12260, N12245);
and AND2 (N12261, N12259, N459);
nor NOR4 (N12262, N12261, N538, N1237, N301);
or OR4 (N12263, N12236, N8083, N12002, N3996);
and AND4 (N12264, N12262, N2306, N6946, N10081);
nand NAND2 (N12265, N12255, N8502);
and AND4 (N12266, N12254, N4164, N2863, N4583);
and AND4 (N12267, N12253, N1401, N10672, N6357);
not NOT1 (N12268, N12264);
xor XOR2 (N12269, N12251, N8036);
and AND4 (N12270, N12267, N6235, N4635, N3833);
or OR4 (N12271, N12268, N4805, N7805, N7310);
not NOT1 (N12272, N12238);
nor NOR3 (N12273, N12260, N6051, N575);
xor XOR2 (N12274, N12270, N350);
and AND3 (N12275, N12269, N2877, N4031);
nand NAND2 (N12276, N12258, N162);
nor NOR2 (N12277, N12271, N10763);
nand NAND2 (N12278, N12275, N10934);
nor NOR2 (N12279, N12263, N6337);
not NOT1 (N12280, N12257);
nand NAND2 (N12281, N12273, N12274);
and AND3 (N12282, N575, N2216, N595);
nand NAND2 (N12283, N12276, N196);
or OR4 (N12284, N12272, N8696, N89, N7561);
not NOT1 (N12285, N12284);
and AND3 (N12286, N12277, N4807, N5999);
nand NAND2 (N12287, N12278, N548);
buf BUF1 (N12288, N12283);
or OR2 (N12289, N12286, N6016);
buf BUF1 (N12290, N12289);
nor NOR4 (N12291, N12287, N7837, N8308, N6303);
xor XOR2 (N12292, N12281, N8246);
buf BUF1 (N12293, N12291);
xor XOR2 (N12294, N12285, N11469);
xor XOR2 (N12295, N12265, N2717);
and AND3 (N12296, N12292, N8525, N5966);
nand NAND4 (N12297, N12266, N10254, N6318, N726);
or OR4 (N12298, N12282, N5565, N1216, N7737);
nor NOR3 (N12299, N12293, N1849, N9577);
buf BUF1 (N12300, N12279);
xor XOR2 (N12301, N12300, N8135);
and AND3 (N12302, N12290, N831, N7080);
xor XOR2 (N12303, N12301, N4610);
xor XOR2 (N12304, N12295, N913);
xor XOR2 (N12305, N12299, N8348);
or OR3 (N12306, N12298, N11793, N1708);
xor XOR2 (N12307, N12303, N11692);
and AND2 (N12308, N12280, N1717);
and AND2 (N12309, N12296, N664);
buf BUF1 (N12310, N12305);
buf BUF1 (N12311, N12308);
buf BUF1 (N12312, N12302);
xor XOR2 (N12313, N12297, N6275);
or OR2 (N12314, N12313, N1219);
or OR2 (N12315, N12304, N4298);
nand NAND4 (N12316, N12314, N2367, N6824, N9118);
buf BUF1 (N12317, N12316);
and AND3 (N12318, N12317, N11831, N5183);
and AND2 (N12319, N12309, N11014);
or OR2 (N12320, N12318, N12049);
or OR2 (N12321, N12315, N11338);
xor XOR2 (N12322, N12319, N11269);
or OR3 (N12323, N12311, N6862, N10090);
or OR2 (N12324, N12321, N1480);
not NOT1 (N12325, N12320);
xor XOR2 (N12326, N12288, N7963);
and AND4 (N12327, N12307, N7609, N1844, N3157);
and AND4 (N12328, N12327, N7105, N9364, N4584);
nand NAND2 (N12329, N12294, N5732);
not NOT1 (N12330, N12312);
nor NOR2 (N12331, N12328, N6339);
nand NAND2 (N12332, N12325, N4648);
and AND4 (N12333, N12329, N8678, N10812, N7247);
xor XOR2 (N12334, N12324, N872);
nand NAND3 (N12335, N12326, N4399, N2688);
nor NOR3 (N12336, N12330, N11769, N1423);
not NOT1 (N12337, N12322);
and AND4 (N12338, N12337, N9528, N9098, N475);
nand NAND4 (N12339, N12335, N5314, N1340, N6148);
and AND2 (N12340, N12338, N10100);
or OR4 (N12341, N12334, N6191, N8374, N1625);
nor NOR4 (N12342, N12331, N1941, N10477, N12139);
nor NOR2 (N12343, N12340, N8543);
xor XOR2 (N12344, N12306, N5780);
xor XOR2 (N12345, N12343, N590);
and AND3 (N12346, N12344, N8666, N5070);
nand NAND4 (N12347, N12345, N12197, N10828, N10091);
buf BUF1 (N12348, N12341);
or OR3 (N12349, N12323, N5901, N5201);
and AND4 (N12350, N12342, N8922, N9414, N11821);
buf BUF1 (N12351, N12336);
and AND2 (N12352, N12339, N5537);
buf BUF1 (N12353, N12310);
nor NOR4 (N12354, N12346, N1715, N5827, N11422);
xor XOR2 (N12355, N12350, N6025);
or OR4 (N12356, N12347, N5105, N12250, N9420);
not NOT1 (N12357, N12333);
xor XOR2 (N12358, N12348, N1415);
xor XOR2 (N12359, N12358, N10020);
not NOT1 (N12360, N12332);
buf BUF1 (N12361, N12355);
buf BUF1 (N12362, N12349);
xor XOR2 (N12363, N12351, N1480);
nand NAND4 (N12364, N12363, N8577, N11522, N5756);
and AND3 (N12365, N12360, N221, N8571);
buf BUF1 (N12366, N12352);
buf BUF1 (N12367, N12362);
and AND3 (N12368, N12354, N3804, N945);
or OR4 (N12369, N12353, N17, N7026, N12124);
not NOT1 (N12370, N12366);
and AND4 (N12371, N12357, N12223, N5132, N6777);
and AND3 (N12372, N12364, N11544, N973);
or OR2 (N12373, N12356, N8938);
nand NAND3 (N12374, N12361, N10298, N4888);
nor NOR3 (N12375, N12365, N11960, N10764);
xor XOR2 (N12376, N12370, N539);
or OR3 (N12377, N12372, N649, N4552);
nor NOR4 (N12378, N12359, N9969, N7649, N3917);
xor XOR2 (N12379, N12373, N7520);
nand NAND3 (N12380, N12379, N5425, N1281);
and AND3 (N12381, N12371, N9253, N6767);
not NOT1 (N12382, N12369);
xor XOR2 (N12383, N12375, N7454);
not NOT1 (N12384, N12368);
nor NOR3 (N12385, N12377, N8882, N3452);
xor XOR2 (N12386, N12381, N3582);
not NOT1 (N12387, N12382);
nand NAND2 (N12388, N12376, N11831);
and AND4 (N12389, N12386, N2085, N4731, N3702);
nor NOR4 (N12390, N12384, N9012, N4235, N6102);
xor XOR2 (N12391, N12390, N8757);
or OR4 (N12392, N12387, N4228, N5855, N10394);
or OR4 (N12393, N12367, N7326, N4751, N1728);
nor NOR4 (N12394, N12388, N1377, N3525, N11803);
nand NAND2 (N12395, N12393, N1049);
nor NOR3 (N12396, N12389, N10136, N11526);
or OR2 (N12397, N12374, N5996);
buf BUF1 (N12398, N12383);
nand NAND2 (N12399, N12392, N5000);
or OR4 (N12400, N12399, N9405, N10803, N3672);
nand NAND4 (N12401, N12394, N4715, N4088, N10195);
xor XOR2 (N12402, N12378, N3318);
or OR4 (N12403, N12395, N6798, N8663, N6869);
nor NOR2 (N12404, N12396, N2220);
not NOT1 (N12405, N12397);
xor XOR2 (N12406, N12403, N9470);
buf BUF1 (N12407, N12391);
nor NOR4 (N12408, N12398, N2503, N12202, N4645);
or OR3 (N12409, N12400, N12058, N12367);
not NOT1 (N12410, N12405);
and AND4 (N12411, N12410, N4354, N10679, N12046);
xor XOR2 (N12412, N12404, N6578);
and AND2 (N12413, N12412, N10040);
xor XOR2 (N12414, N12411, N2738);
nor NOR4 (N12415, N12406, N4898, N1945, N11896);
buf BUF1 (N12416, N12385);
nand NAND4 (N12417, N12380, N5547, N10073, N9557);
nor NOR4 (N12418, N12409, N6305, N4690, N422);
nor NOR3 (N12419, N12408, N1102, N2383);
not NOT1 (N12420, N12413);
or OR3 (N12421, N12419, N6296, N1911);
xor XOR2 (N12422, N12401, N763);
not NOT1 (N12423, N12417);
buf BUF1 (N12424, N12418);
nor NOR4 (N12425, N12424, N5096, N7009, N666);
not NOT1 (N12426, N12420);
or OR2 (N12427, N12423, N629);
nand NAND4 (N12428, N12416, N961, N2796, N9492);
or OR4 (N12429, N12402, N4765, N8446, N12257);
nor NOR3 (N12430, N12429, N6477, N3799);
and AND2 (N12431, N12414, N3899);
not NOT1 (N12432, N12430);
and AND4 (N12433, N12432, N227, N2008, N2525);
not NOT1 (N12434, N12421);
nor NOR2 (N12435, N12431, N2502);
nand NAND3 (N12436, N12433, N10493, N3838);
xor XOR2 (N12437, N12415, N355);
nand NAND2 (N12438, N12428, N11643);
xor XOR2 (N12439, N12434, N10018);
and AND2 (N12440, N12437, N6964);
and AND2 (N12441, N12426, N3534);
not NOT1 (N12442, N12438);
nor NOR2 (N12443, N12422, N5149);
buf BUF1 (N12444, N12407);
or OR2 (N12445, N12440, N8725);
nand NAND3 (N12446, N12435, N6647, N33);
and AND4 (N12447, N12446, N5392, N2487, N9060);
and AND4 (N12448, N12447, N6747, N10771, N7488);
nor NOR3 (N12449, N12441, N4186, N4384);
and AND2 (N12450, N12439, N9270);
nor NOR4 (N12451, N12445, N11184, N7926, N11406);
or OR2 (N12452, N12449, N10718);
buf BUF1 (N12453, N12448);
and AND3 (N12454, N12451, N5831, N2124);
not NOT1 (N12455, N12450);
nand NAND4 (N12456, N12425, N9841, N4845, N804);
and AND2 (N12457, N12444, N4485);
buf BUF1 (N12458, N12457);
nor NOR4 (N12459, N12453, N8305, N673, N3221);
nor NOR2 (N12460, N12459, N7304);
buf BUF1 (N12461, N12456);
not NOT1 (N12462, N12452);
nor NOR2 (N12463, N12454, N11544);
and AND3 (N12464, N12443, N11330, N3623);
nor NOR2 (N12465, N12460, N5469);
xor XOR2 (N12466, N12463, N1944);
or OR3 (N12467, N12427, N6418, N2118);
nand NAND3 (N12468, N12436, N5577, N2329);
nand NAND2 (N12469, N12442, N2138);
not NOT1 (N12470, N12465);
nand NAND3 (N12471, N12461, N3865, N374);
and AND2 (N12472, N12470, N9460);
nand NAND3 (N12473, N12468, N2155, N7818);
xor XOR2 (N12474, N12472, N11078);
nor NOR4 (N12475, N12464, N10137, N1944, N5029);
xor XOR2 (N12476, N12474, N2465);
or OR4 (N12477, N12471, N3851, N1397, N11164);
and AND3 (N12478, N12455, N5106, N9672);
or OR3 (N12479, N12473, N8472, N7678);
not NOT1 (N12480, N12462);
or OR4 (N12481, N12475, N11100, N12028, N2817);
nor NOR4 (N12482, N12467, N9487, N6328, N10893);
not NOT1 (N12483, N12466);
and AND2 (N12484, N12480, N11407);
not NOT1 (N12485, N12458);
and AND2 (N12486, N12478, N5263);
xor XOR2 (N12487, N12486, N6505);
nor NOR2 (N12488, N12484, N8041);
xor XOR2 (N12489, N12487, N8063);
not NOT1 (N12490, N12476);
and AND3 (N12491, N12485, N6451, N6420);
or OR2 (N12492, N12481, N3390);
not NOT1 (N12493, N12491);
or OR2 (N12494, N12490, N11682);
and AND2 (N12495, N12494, N6210);
buf BUF1 (N12496, N12479);
not NOT1 (N12497, N12483);
not NOT1 (N12498, N12489);
buf BUF1 (N12499, N12498);
buf BUF1 (N12500, N12496);
xor XOR2 (N12501, N12499, N2141);
or OR3 (N12502, N12469, N9716, N1347);
nor NOR4 (N12503, N12502, N475, N3778, N1065);
not NOT1 (N12504, N12497);
not NOT1 (N12505, N12477);
xor XOR2 (N12506, N12505, N3574);
or OR2 (N12507, N12501, N10562);
nor NOR3 (N12508, N12495, N10940, N8253);
or OR3 (N12509, N12500, N6059, N275);
and AND2 (N12510, N12488, N12392);
and AND2 (N12511, N12504, N3044);
nand NAND2 (N12512, N12482, N4474);
not NOT1 (N12513, N12508);
nor NOR4 (N12514, N12511, N10405, N9783, N9681);
and AND3 (N12515, N12492, N5882, N518);
nand NAND2 (N12516, N12513, N6498);
and AND3 (N12517, N12516, N7311, N5855);
or OR2 (N12518, N12514, N152);
xor XOR2 (N12519, N12507, N3091);
xor XOR2 (N12520, N12517, N6582);
nand NAND2 (N12521, N12506, N10055);
buf BUF1 (N12522, N12510);
nor NOR2 (N12523, N12515, N10989);
buf BUF1 (N12524, N12520);
not NOT1 (N12525, N12493);
xor XOR2 (N12526, N12512, N4954);
nor NOR3 (N12527, N12519, N1126, N8422);
not NOT1 (N12528, N12524);
xor XOR2 (N12529, N12521, N1522);
or OR3 (N12530, N12526, N11551, N4581);
or OR3 (N12531, N12523, N1403, N6621);
nor NOR3 (N12532, N12530, N11675, N2081);
nand NAND2 (N12533, N12531, N11598);
nor NOR4 (N12534, N12532, N1348, N7040, N4956);
xor XOR2 (N12535, N12534, N4548);
nor NOR2 (N12536, N12509, N1047);
or OR4 (N12537, N12533, N8355, N112, N136);
nand NAND2 (N12538, N12536, N1347);
nor NOR4 (N12539, N12537, N3930, N1612, N4169);
buf BUF1 (N12540, N12522);
nand NAND4 (N12541, N12535, N11991, N9869, N4693);
nor NOR3 (N12542, N12538, N1214, N3076);
and AND2 (N12543, N12542, N7535);
nand NAND4 (N12544, N12527, N640, N11036, N8827);
and AND2 (N12545, N12540, N6530);
buf BUF1 (N12546, N12528);
or OR3 (N12547, N12529, N3024, N8508);
buf BUF1 (N12548, N12503);
buf BUF1 (N12549, N12546);
buf BUF1 (N12550, N12544);
and AND3 (N12551, N12541, N5371, N2257);
nand NAND2 (N12552, N12548, N4567);
buf BUF1 (N12553, N12525);
nand NAND3 (N12554, N12553, N10174, N6972);
nand NAND4 (N12555, N12547, N9004, N6971, N1278);
xor XOR2 (N12556, N12539, N3700);
nand NAND2 (N12557, N12543, N2656);
nand NAND2 (N12558, N12549, N6554);
xor XOR2 (N12559, N12550, N9548);
nor NOR2 (N12560, N12518, N11031);
nor NOR2 (N12561, N12558, N528);
nand NAND2 (N12562, N12561, N4019);
or OR2 (N12563, N12559, N6241);
and AND3 (N12564, N12554, N129, N1280);
not NOT1 (N12565, N12545);
nor NOR3 (N12566, N12555, N7285, N5259);
nand NAND3 (N12567, N12565, N2996, N5974);
buf BUF1 (N12568, N12551);
nor NOR2 (N12569, N12568, N10620);
not NOT1 (N12570, N12566);
nor NOR4 (N12571, N12570, N1777, N5251, N6095);
buf BUF1 (N12572, N12571);
not NOT1 (N12573, N12567);
xor XOR2 (N12574, N12562, N7624);
or OR2 (N12575, N12560, N12023);
not NOT1 (N12576, N12573);
and AND3 (N12577, N12552, N11190, N625);
and AND4 (N12578, N12557, N3773, N1321, N2108);
nor NOR4 (N12579, N12556, N12083, N1024, N939);
buf BUF1 (N12580, N12569);
or OR4 (N12581, N12574, N2212, N4663, N7533);
nor NOR4 (N12582, N12577, N1030, N317, N2614);
not NOT1 (N12583, N12572);
buf BUF1 (N12584, N12578);
not NOT1 (N12585, N12575);
xor XOR2 (N12586, N12583, N8807);
nor NOR3 (N12587, N12579, N960, N6084);
nor NOR3 (N12588, N12581, N3448, N3253);
not NOT1 (N12589, N12584);
buf BUF1 (N12590, N12576);
and AND4 (N12591, N12582, N8101, N4523, N9902);
and AND3 (N12592, N12586, N5875, N1626);
or OR4 (N12593, N12591, N7154, N7426, N6845);
and AND2 (N12594, N12589, N3087);
xor XOR2 (N12595, N12590, N10206);
nand NAND4 (N12596, N12594, N7106, N10104, N6083);
buf BUF1 (N12597, N12580);
not NOT1 (N12598, N12587);
not NOT1 (N12599, N12597);
and AND3 (N12600, N12588, N12060, N5852);
buf BUF1 (N12601, N12598);
not NOT1 (N12602, N12564);
buf BUF1 (N12603, N12563);
and AND4 (N12604, N12601, N338, N5881, N12595);
or OR3 (N12605, N3120, N3356, N12084);
nor NOR4 (N12606, N12592, N7382, N4343, N8957);
buf BUF1 (N12607, N12585);
buf BUF1 (N12608, N12596);
buf BUF1 (N12609, N12600);
nand NAND3 (N12610, N12608, N952, N5900);
nor NOR4 (N12611, N12593, N3450, N8198, N10860);
nor NOR2 (N12612, N12606, N9772);
and AND4 (N12613, N12604, N283, N11933, N1367);
nand NAND3 (N12614, N12609, N791, N5785);
nor NOR4 (N12615, N12602, N10681, N6278, N3862);
nand NAND4 (N12616, N12605, N3779, N4978, N5259);
xor XOR2 (N12617, N12611, N5470);
buf BUF1 (N12618, N12599);
nor NOR2 (N12619, N12614, N8183);
nand NAND4 (N12620, N12613, N11879, N12465, N7730);
buf BUF1 (N12621, N12616);
buf BUF1 (N12622, N12607);
nor NOR4 (N12623, N12612, N5295, N9445, N7268);
or OR3 (N12624, N12620, N2098, N11144);
buf BUF1 (N12625, N12621);
not NOT1 (N12626, N12623);
and AND4 (N12627, N12618, N7334, N6408, N3257);
nand NAND4 (N12628, N12617, N1551, N10270, N4356);
not NOT1 (N12629, N12619);
nand NAND3 (N12630, N12628, N4279, N12473);
nand NAND3 (N12631, N12630, N12429, N5969);
or OR2 (N12632, N12626, N4422);
and AND4 (N12633, N12610, N7834, N8322, N53);
or OR3 (N12634, N12633, N6719, N4741);
not NOT1 (N12635, N12629);
buf BUF1 (N12636, N12622);
xor XOR2 (N12637, N12631, N10946);
nand NAND3 (N12638, N12625, N36, N7227);
or OR2 (N12639, N12632, N12456);
not NOT1 (N12640, N12638);
not NOT1 (N12641, N12640);
xor XOR2 (N12642, N12634, N714);
nand NAND4 (N12643, N12641, N1288, N9780, N11204);
nand NAND2 (N12644, N12636, N9495);
not NOT1 (N12645, N12637);
and AND3 (N12646, N12645, N10101, N5806);
not NOT1 (N12647, N12646);
xor XOR2 (N12648, N12647, N4573);
nand NAND4 (N12649, N12615, N6280, N5969, N10247);
buf BUF1 (N12650, N12642);
and AND4 (N12651, N12643, N5234, N4244, N10526);
xor XOR2 (N12652, N12644, N9854);
buf BUF1 (N12653, N12651);
nand NAND4 (N12654, N12603, N10209, N3837, N6269);
buf BUF1 (N12655, N12649);
xor XOR2 (N12656, N12627, N2100);
buf BUF1 (N12657, N12624);
or OR2 (N12658, N12657, N11601);
nand NAND4 (N12659, N12656, N1839, N8361, N8330);
or OR3 (N12660, N12659, N7478, N7105);
or OR4 (N12661, N12660, N6368, N9172, N4479);
xor XOR2 (N12662, N12648, N10968);
nand NAND2 (N12663, N12635, N3075);
nor NOR2 (N12664, N12653, N9131);
nor NOR3 (N12665, N12658, N7595, N5430);
or OR3 (N12666, N12655, N10255, N11933);
nor NOR3 (N12667, N12639, N4781, N7625);
or OR3 (N12668, N12652, N7100, N9200);
and AND4 (N12669, N12661, N6397, N6729, N12662);
nand NAND3 (N12670, N8155, N10096, N4412);
nor NOR2 (N12671, N12664, N9133);
xor XOR2 (N12672, N12666, N5394);
not NOT1 (N12673, N12671);
xor XOR2 (N12674, N12650, N3097);
xor XOR2 (N12675, N12668, N1528);
nor NOR2 (N12676, N12669, N10484);
xor XOR2 (N12677, N12663, N3305);
and AND4 (N12678, N12677, N303, N8849, N1039);
nand NAND4 (N12679, N12678, N5694, N329, N6820);
or OR2 (N12680, N12654, N3662);
xor XOR2 (N12681, N12673, N9927);
xor XOR2 (N12682, N12679, N9387);
nand NAND3 (N12683, N12672, N3515, N12243);
nand NAND2 (N12684, N12676, N2700);
or OR3 (N12685, N12670, N6386, N6899);
and AND3 (N12686, N12680, N731, N5442);
and AND2 (N12687, N12674, N10094);
and AND2 (N12688, N12686, N1939);
nand NAND4 (N12689, N12684, N2496, N8277, N9987);
not NOT1 (N12690, N12687);
and AND4 (N12691, N12683, N7284, N708, N7151);
buf BUF1 (N12692, N12688);
nand NAND3 (N12693, N12691, N9433, N2227);
not NOT1 (N12694, N12675);
not NOT1 (N12695, N12667);
nor NOR4 (N12696, N12685, N5159, N3976, N4368);
nand NAND2 (N12697, N12692, N4068);
not NOT1 (N12698, N12696);
nor NOR2 (N12699, N12694, N4676);
or OR4 (N12700, N12697, N4035, N187, N1150);
or OR3 (N12701, N12700, N5831, N4313);
xor XOR2 (N12702, N12695, N3446);
nor NOR3 (N12703, N12690, N7187, N7423);
or OR3 (N12704, N12698, N2629, N8554);
buf BUF1 (N12705, N12702);
nor NOR2 (N12706, N12689, N11511);
or OR2 (N12707, N12681, N3501);
nor NOR3 (N12708, N12706, N10746, N9728);
not NOT1 (N12709, N12682);
nand NAND3 (N12710, N12709, N9323, N1775);
xor XOR2 (N12711, N12699, N11537);
buf BUF1 (N12712, N12703);
not NOT1 (N12713, N12708);
not NOT1 (N12714, N12711);
nor NOR3 (N12715, N12701, N7086, N6715);
buf BUF1 (N12716, N12665);
not NOT1 (N12717, N12693);
not NOT1 (N12718, N12710);
not NOT1 (N12719, N12716);
buf BUF1 (N12720, N12713);
or OR4 (N12721, N12720, N10437, N10852, N1753);
nor NOR4 (N12722, N12717, N7916, N2463, N10003);
xor XOR2 (N12723, N12705, N10618);
nor NOR4 (N12724, N12723, N5742, N10402, N8470);
or OR3 (N12725, N12724, N5848, N8461);
nand NAND4 (N12726, N12721, N11530, N7858, N12443);
nand NAND2 (N12727, N12722, N3714);
nand NAND2 (N12728, N12712, N7044);
not NOT1 (N12729, N12704);
and AND2 (N12730, N12715, N6592);
or OR3 (N12731, N12726, N9790, N380);
nor NOR4 (N12732, N12729, N4301, N2881, N2453);
nor NOR3 (N12733, N12731, N4736, N7947);
nor NOR2 (N12734, N12730, N12284);
nor NOR4 (N12735, N12707, N1105, N10123, N432);
nor NOR2 (N12736, N12725, N11193);
buf BUF1 (N12737, N12719);
xor XOR2 (N12738, N12733, N2522);
xor XOR2 (N12739, N12718, N6483);
not NOT1 (N12740, N12735);
and AND4 (N12741, N12732, N11848, N1041, N1091);
not NOT1 (N12742, N12734);
nand NAND2 (N12743, N12740, N10541);
nand NAND3 (N12744, N12738, N11835, N7063);
and AND3 (N12745, N12741, N5017, N9228);
buf BUF1 (N12746, N12743);
buf BUF1 (N12747, N12737);
xor XOR2 (N12748, N12742, N6146);
not NOT1 (N12749, N12744);
not NOT1 (N12750, N12748);
not NOT1 (N12751, N12727);
nor NOR3 (N12752, N12736, N3483, N1053);
buf BUF1 (N12753, N12747);
or OR4 (N12754, N12752, N5644, N5731, N3417);
xor XOR2 (N12755, N12753, N4242);
and AND4 (N12756, N12728, N5728, N9466, N6628);
nor NOR2 (N12757, N12755, N685);
nand NAND4 (N12758, N12750, N9098, N11173, N8055);
buf BUF1 (N12759, N12739);
buf BUF1 (N12760, N12714);
nor NOR2 (N12761, N12749, N3960);
and AND3 (N12762, N12745, N7037, N9707);
or OR3 (N12763, N12757, N7575, N3996);
nor NOR3 (N12764, N12762, N12022, N12664);
not NOT1 (N12765, N12758);
nand NAND3 (N12766, N12765, N1293, N9534);
buf BUF1 (N12767, N12746);
and AND2 (N12768, N12763, N4133);
nor NOR2 (N12769, N12760, N905);
nor NOR3 (N12770, N12751, N4109, N2019);
or OR4 (N12771, N12768, N4350, N2703, N11158);
nor NOR2 (N12772, N12761, N7810);
xor XOR2 (N12773, N12766, N11180);
buf BUF1 (N12774, N12754);
buf BUF1 (N12775, N12756);
or OR2 (N12776, N12759, N4408);
or OR3 (N12777, N12771, N3060, N1687);
not NOT1 (N12778, N12770);
and AND2 (N12779, N12776, N2269);
buf BUF1 (N12780, N12767);
nor NOR3 (N12781, N12778, N2043, N973);
nor NOR3 (N12782, N12775, N7681, N8380);
and AND3 (N12783, N12780, N2049, N9377);
nor NOR4 (N12784, N12772, N9215, N3489, N2071);
xor XOR2 (N12785, N12781, N522);
buf BUF1 (N12786, N12769);
nor NOR4 (N12787, N12779, N7414, N2831, N10960);
or OR2 (N12788, N12787, N2024);
or OR2 (N12789, N12784, N8843);
not NOT1 (N12790, N12764);
nor NOR2 (N12791, N12777, N588);
xor XOR2 (N12792, N12785, N9394);
and AND4 (N12793, N12789, N11664, N10445, N2949);
not NOT1 (N12794, N12782);
or OR3 (N12795, N12788, N10728, N753);
or OR2 (N12796, N12774, N9077);
and AND4 (N12797, N12791, N1332, N5545, N4345);
or OR3 (N12798, N12793, N3145, N10087);
and AND2 (N12799, N12794, N1978);
nor NOR2 (N12800, N12792, N7531);
nand NAND3 (N12801, N12798, N533, N2095);
not NOT1 (N12802, N12790);
and AND4 (N12803, N12800, N6769, N8168, N1930);
xor XOR2 (N12804, N12795, N3824);
and AND4 (N12805, N12797, N6892, N11473, N3404);
xor XOR2 (N12806, N12804, N8493);
or OR2 (N12807, N12799, N8248);
nand NAND2 (N12808, N12805, N9670);
not NOT1 (N12809, N12786);
nand NAND3 (N12810, N12803, N4943, N9988);
xor XOR2 (N12811, N12810, N12669);
or OR3 (N12812, N12773, N9486, N9571);
and AND4 (N12813, N12808, N2854, N9982, N1809);
not NOT1 (N12814, N12811);
xor XOR2 (N12815, N12806, N3453);
not NOT1 (N12816, N12814);
and AND2 (N12817, N12813, N8522);
and AND4 (N12818, N12796, N12427, N7232, N12651);
and AND4 (N12819, N12816, N11754, N692, N5146);
buf BUF1 (N12820, N12801);
and AND3 (N12821, N12820, N2739, N3966);
buf BUF1 (N12822, N12809);
buf BUF1 (N12823, N12819);
xor XOR2 (N12824, N12822, N1126);
nor NOR4 (N12825, N12812, N6048, N10600, N2455);
nor NOR4 (N12826, N12783, N8488, N12624, N705);
buf BUF1 (N12827, N12821);
nor NOR2 (N12828, N12807, N12642);
buf BUF1 (N12829, N12828);
nor NOR4 (N12830, N12818, N7789, N11077, N8432);
and AND4 (N12831, N12802, N6863, N12353, N769);
not NOT1 (N12832, N12823);
not NOT1 (N12833, N12826);
or OR3 (N12834, N12815, N1498, N2258);
and AND3 (N12835, N12833, N11812, N3269);
and AND4 (N12836, N12831, N6675, N1264, N10260);
nand NAND2 (N12837, N12827, N1098);
xor XOR2 (N12838, N12825, N2780);
not NOT1 (N12839, N12829);
xor XOR2 (N12840, N12835, N1991);
nor NOR4 (N12841, N12834, N4544, N10604, N7582);
not NOT1 (N12842, N12839);
xor XOR2 (N12843, N12832, N3914);
nand NAND3 (N12844, N12843, N8995, N4403);
or OR4 (N12845, N12838, N7817, N2239, N7026);
nand NAND2 (N12846, N12844, N7177);
not NOT1 (N12847, N12841);
not NOT1 (N12848, N12817);
nor NOR3 (N12849, N12846, N7331, N3551);
xor XOR2 (N12850, N12837, N8660);
and AND4 (N12851, N12830, N8558, N6660, N2128);
xor XOR2 (N12852, N12851, N5246);
and AND3 (N12853, N12824, N1120, N3386);
not NOT1 (N12854, N12845);
or OR2 (N12855, N12854, N5437);
not NOT1 (N12856, N12848);
and AND2 (N12857, N12842, N420);
buf BUF1 (N12858, N12850);
nor NOR4 (N12859, N12857, N6857, N10566, N2565);
nand NAND3 (N12860, N12849, N10715, N5088);
not NOT1 (N12861, N12856);
or OR3 (N12862, N12858, N427, N3334);
not NOT1 (N12863, N12836);
nand NAND3 (N12864, N12840, N2248, N4985);
buf BUF1 (N12865, N12863);
and AND2 (N12866, N12855, N6875);
not NOT1 (N12867, N12865);
nand NAND2 (N12868, N12862, N3852);
nor NOR2 (N12869, N12868, N2037);
xor XOR2 (N12870, N12861, N819);
nor NOR4 (N12871, N12869, N8421, N9486, N6137);
nor NOR4 (N12872, N12853, N11498, N5001, N6270);
buf BUF1 (N12873, N12867);
and AND3 (N12874, N12866, N4107, N434);
buf BUF1 (N12875, N12852);
and AND3 (N12876, N12864, N8755, N9773);
nor NOR3 (N12877, N12874, N9673, N3715);
and AND3 (N12878, N12859, N5585, N2207);
not NOT1 (N12879, N12877);
nand NAND4 (N12880, N12860, N7880, N2775, N6455);
nor NOR3 (N12881, N12880, N5460, N5799);
nor NOR2 (N12882, N12878, N2130);
not NOT1 (N12883, N12876);
nor NOR2 (N12884, N12883, N5514);
nand NAND4 (N12885, N12875, N8934, N862, N5501);
nand NAND4 (N12886, N12871, N12864, N9428, N1030);
xor XOR2 (N12887, N12881, N3494);
or OR2 (N12888, N12847, N2306);
buf BUF1 (N12889, N12885);
nand NAND4 (N12890, N12870, N6197, N4493, N11036);
and AND4 (N12891, N12873, N974, N3550, N659);
xor XOR2 (N12892, N12888, N7200);
nand NAND2 (N12893, N12879, N3128);
nor NOR2 (N12894, N12893, N10089);
nor NOR2 (N12895, N12889, N12700);
or OR4 (N12896, N12892, N3979, N161, N932);
nor NOR2 (N12897, N12896, N1587);
nor NOR3 (N12898, N12882, N9496, N6437);
not NOT1 (N12899, N12897);
xor XOR2 (N12900, N12899, N6370);
nand NAND3 (N12901, N12894, N3283, N9918);
not NOT1 (N12902, N12895);
or OR3 (N12903, N12901, N7265, N6681);
nor NOR3 (N12904, N12898, N3745, N5117);
and AND2 (N12905, N12884, N7963);
not NOT1 (N12906, N12903);
buf BUF1 (N12907, N12900);
or OR3 (N12908, N12904, N8165, N9083);
xor XOR2 (N12909, N12887, N5000);
not NOT1 (N12910, N12891);
nand NAND4 (N12911, N12890, N4336, N2800, N6319);
and AND2 (N12912, N12872, N12090);
nand NAND4 (N12913, N12909, N7339, N8525, N6225);
xor XOR2 (N12914, N12911, N11504);
nor NOR3 (N12915, N12907, N1979, N2800);
or OR2 (N12916, N12908, N5628);
and AND2 (N12917, N12916, N4739);
buf BUF1 (N12918, N12910);
nor NOR3 (N12919, N12917, N12856, N12170);
buf BUF1 (N12920, N12919);
or OR4 (N12921, N12920, N6925, N159, N10416);
not NOT1 (N12922, N12915);
or OR3 (N12923, N12902, N7913, N2906);
buf BUF1 (N12924, N12886);
or OR2 (N12925, N12913, N7124);
buf BUF1 (N12926, N12914);
or OR3 (N12927, N12905, N5296, N10180);
nor NOR2 (N12928, N12927, N4551);
and AND3 (N12929, N12918, N6099, N9639);
nand NAND4 (N12930, N12912, N5181, N3820, N7538);
not NOT1 (N12931, N12928);
xor XOR2 (N12932, N12923, N180);
nand NAND3 (N12933, N12926, N1100, N2773);
buf BUF1 (N12934, N12921);
nor NOR4 (N12935, N12924, N1353, N1747, N8600);
or OR4 (N12936, N12922, N10186, N5350, N8481);
nor NOR4 (N12937, N12930, N10532, N1784, N838);
nor NOR2 (N12938, N12935, N8283);
and AND4 (N12939, N12931, N9461, N2349, N9724);
nor NOR3 (N12940, N12934, N979, N12799);
not NOT1 (N12941, N12929);
not NOT1 (N12942, N12936);
and AND4 (N12943, N12941, N10922, N273, N12893);
buf BUF1 (N12944, N12940);
and AND2 (N12945, N12944, N12636);
buf BUF1 (N12946, N12925);
or OR3 (N12947, N12938, N3214, N3831);
not NOT1 (N12948, N12943);
and AND4 (N12949, N12945, N12271, N6236, N12743);
buf BUF1 (N12950, N12949);
buf BUF1 (N12951, N12933);
not NOT1 (N12952, N12951);
or OR3 (N12953, N12942, N11305, N6909);
nand NAND4 (N12954, N12932, N10772, N7903, N10023);
not NOT1 (N12955, N12906);
or OR4 (N12956, N12947, N2525, N12143, N12871);
or OR3 (N12957, N12954, N7188, N7008);
xor XOR2 (N12958, N12953, N11409);
nor NOR2 (N12959, N12939, N8530);
and AND4 (N12960, N12950, N2084, N9638, N9776);
and AND2 (N12961, N12959, N2625);
buf BUF1 (N12962, N12957);
nor NOR2 (N12963, N12955, N35);
xor XOR2 (N12964, N12948, N1042);
not NOT1 (N12965, N12958);
and AND2 (N12966, N12961, N8360);
or OR2 (N12967, N12952, N1700);
buf BUF1 (N12968, N12967);
xor XOR2 (N12969, N12956, N9699);
xor XOR2 (N12970, N12968, N2295);
buf BUF1 (N12971, N12969);
nor NOR3 (N12972, N12970, N5206, N8589);
nand NAND4 (N12973, N12963, N3263, N12561, N934);
buf BUF1 (N12974, N12964);
nand NAND4 (N12975, N12973, N5443, N9941, N11783);
nand NAND4 (N12976, N12937, N4862, N9726, N12842);
nand NAND4 (N12977, N12946, N10863, N5077, N9566);
not NOT1 (N12978, N12975);
not NOT1 (N12979, N12977);
buf BUF1 (N12980, N12972);
nor NOR2 (N12981, N12974, N2210);
nor NOR2 (N12982, N12962, N7124);
not NOT1 (N12983, N12966);
nand NAND4 (N12984, N12980, N7863, N5198, N2560);
xor XOR2 (N12985, N12984, N1091);
or OR3 (N12986, N12983, N3870, N5077);
nor NOR3 (N12987, N12986, N9383, N1610);
nor NOR4 (N12988, N12965, N4875, N1483, N8185);
nand NAND4 (N12989, N12976, N2992, N9808, N7703);
and AND4 (N12990, N12960, N4907, N1228, N12151);
and AND3 (N12991, N12985, N3277, N12810);
nand NAND4 (N12992, N12989, N3368, N6252, N5785);
and AND3 (N12993, N12992, N5245, N424);
buf BUF1 (N12994, N12979);
and AND4 (N12995, N12982, N9156, N11862, N3933);
nand NAND4 (N12996, N12995, N4711, N12131, N6641);
nor NOR4 (N12997, N12988, N6412, N675, N2432);
buf BUF1 (N12998, N12997);
and AND4 (N12999, N12991, N8643, N8071, N12);
xor XOR2 (N13000, N12998, N10768);
xor XOR2 (N13001, N12987, N9283);
buf BUF1 (N13002, N12981);
buf BUF1 (N13003, N12996);
nor NOR2 (N13004, N12990, N6055);
nand NAND2 (N13005, N12993, N7938);
nand NAND2 (N13006, N13005, N9133);
and AND3 (N13007, N13001, N2817, N10510);
buf BUF1 (N13008, N13007);
and AND3 (N13009, N12994, N11026, N3623);
nor NOR3 (N13010, N12971, N8457, N10440);
not NOT1 (N13011, N12978);
not NOT1 (N13012, N13003);
not NOT1 (N13013, N12999);
or OR2 (N13014, N13012, N12776);
or OR4 (N13015, N13004, N3278, N9299, N4278);
nand NAND2 (N13016, N13009, N6927);
xor XOR2 (N13017, N13010, N8321);
buf BUF1 (N13018, N13013);
not NOT1 (N13019, N13008);
not NOT1 (N13020, N13018);
nor NOR4 (N13021, N13000, N12494, N1941, N12013);
or OR4 (N13022, N13002, N1869, N1201, N11009);
xor XOR2 (N13023, N13014, N12673);
nand NAND4 (N13024, N13019, N8271, N4017, N6058);
buf BUF1 (N13025, N13011);
buf BUF1 (N13026, N13022);
xor XOR2 (N13027, N13015, N4379);
and AND3 (N13028, N13017, N2921, N9408);
xor XOR2 (N13029, N13023, N332);
not NOT1 (N13030, N13006);
buf BUF1 (N13031, N13026);
and AND4 (N13032, N13031, N10841, N7820, N11759);
or OR2 (N13033, N13030, N8796);
or OR2 (N13034, N13027, N1308);
xor XOR2 (N13035, N13028, N4630);
nand NAND3 (N13036, N13032, N3596, N1067);
and AND3 (N13037, N13024, N11266, N6769);
nand NAND3 (N13038, N13016, N6614, N11883);
and AND4 (N13039, N13035, N11673, N10038, N1678);
and AND4 (N13040, N13037, N1306, N9314, N5718);
or OR3 (N13041, N13020, N9018, N7070);
buf BUF1 (N13042, N13040);
nand NAND4 (N13043, N13029, N3795, N3828, N11181);
not NOT1 (N13044, N13036);
xor XOR2 (N13045, N13033, N12234);
buf BUF1 (N13046, N13044);
nor NOR4 (N13047, N13025, N2833, N12107, N8631);
xor XOR2 (N13048, N13046, N6128);
not NOT1 (N13049, N13039);
buf BUF1 (N13050, N13043);
or OR2 (N13051, N13045, N3139);
buf BUF1 (N13052, N13021);
and AND3 (N13053, N13041, N11815, N4267);
or OR3 (N13054, N13047, N10434, N9433);
not NOT1 (N13055, N13053);
buf BUF1 (N13056, N13052);
or OR4 (N13057, N13050, N6945, N7460, N12551);
xor XOR2 (N13058, N13057, N2512);
xor XOR2 (N13059, N13051, N2954);
or OR3 (N13060, N13054, N11105, N1120);
or OR3 (N13061, N13049, N3083, N4885);
buf BUF1 (N13062, N13056);
buf BUF1 (N13063, N13058);
nor NOR2 (N13064, N13034, N9685);
xor XOR2 (N13065, N13061, N4296);
or OR2 (N13066, N13060, N7315);
not NOT1 (N13067, N13064);
xor XOR2 (N13068, N13048, N3488);
nor NOR2 (N13069, N13067, N7348);
buf BUF1 (N13070, N13062);
not NOT1 (N13071, N13066);
nand NAND3 (N13072, N13070, N12975, N12603);
buf BUF1 (N13073, N13038);
nor NOR3 (N13074, N13055, N10121, N2914);
or OR3 (N13075, N13042, N10230, N1880);
and AND4 (N13076, N13071, N3625, N11294, N11301);
and AND4 (N13077, N13068, N12693, N810, N6857);
nor NOR3 (N13078, N13077, N3534, N8837);
not NOT1 (N13079, N13072);
nand NAND3 (N13080, N13079, N8101, N3787);
not NOT1 (N13081, N13059);
nand NAND2 (N13082, N13073, N2059);
xor XOR2 (N13083, N13082, N3374);
and AND4 (N13084, N13078, N2536, N12524, N4117);
nor NOR3 (N13085, N13063, N10757, N4358);
xor XOR2 (N13086, N13076, N5582);
not NOT1 (N13087, N13081);
or OR3 (N13088, N13086, N9320, N12143);
nand NAND3 (N13089, N13084, N5405, N7311);
not NOT1 (N13090, N13083);
and AND3 (N13091, N13090, N7453, N5234);
nor NOR2 (N13092, N13085, N2845);
not NOT1 (N13093, N13074);
nor NOR3 (N13094, N13069, N4415, N1687);
nor NOR2 (N13095, N13093, N8687);
xor XOR2 (N13096, N13095, N3683);
or OR3 (N13097, N13091, N9968, N4079);
or OR4 (N13098, N13097, N6068, N1144, N2403);
xor XOR2 (N13099, N13092, N7484);
nand NAND2 (N13100, N13075, N11359);
nor NOR3 (N13101, N13099, N7291, N4405);
xor XOR2 (N13102, N13080, N5895);
or OR4 (N13103, N13100, N12772, N2113, N1002);
or OR3 (N13104, N13065, N6601, N4988);
and AND2 (N13105, N13103, N12839);
or OR3 (N13106, N13098, N9079, N9661);
buf BUF1 (N13107, N13106);
buf BUF1 (N13108, N13105);
and AND4 (N13109, N13102, N11921, N12748, N11885);
xor XOR2 (N13110, N13108, N4271);
nor NOR3 (N13111, N13104, N2804, N11450);
or OR4 (N13112, N13110, N780, N5395, N6343);
xor XOR2 (N13113, N13112, N2815);
buf BUF1 (N13114, N13113);
buf BUF1 (N13115, N13096);
or OR2 (N13116, N13087, N5505);
not NOT1 (N13117, N13089);
nor NOR4 (N13118, N13115, N12803, N6307, N6537);
xor XOR2 (N13119, N13116, N4418);
and AND3 (N13120, N13107, N5797, N1533);
nor NOR2 (N13121, N13119, N720);
nand NAND2 (N13122, N13094, N12962);
and AND2 (N13123, N13117, N9771);
nor NOR4 (N13124, N13088, N2946, N1014, N3908);
xor XOR2 (N13125, N13101, N905);
and AND2 (N13126, N13111, N5860);
and AND4 (N13127, N13123, N5155, N9569, N3770);
nor NOR3 (N13128, N13118, N3145, N1802);
not NOT1 (N13129, N13114);
or OR4 (N13130, N13120, N1128, N8925, N478);
not NOT1 (N13131, N13125);
nand NAND4 (N13132, N13127, N3405, N6687, N4815);
nand NAND2 (N13133, N13121, N7931);
nor NOR3 (N13134, N13126, N7661, N11299);
nor NOR3 (N13135, N13122, N5615, N12038);
and AND2 (N13136, N13133, N4198);
not NOT1 (N13137, N13128);
or OR3 (N13138, N13131, N5103, N10633);
nand NAND2 (N13139, N13124, N11400);
buf BUF1 (N13140, N13136);
xor XOR2 (N13141, N13132, N11251);
xor XOR2 (N13142, N13140, N3939);
or OR4 (N13143, N13139, N9, N6310, N5368);
xor XOR2 (N13144, N13129, N11271);
or OR4 (N13145, N13143, N163, N24, N3485);
xor XOR2 (N13146, N13144, N3952);
and AND3 (N13147, N13109, N4230, N851);
or OR3 (N13148, N13146, N10922, N8102);
and AND3 (N13149, N13145, N4590, N10534);
nor NOR4 (N13150, N13147, N6965, N9589, N2538);
nand NAND4 (N13151, N13135, N4303, N2225, N6960);
xor XOR2 (N13152, N13149, N7504);
or OR2 (N13153, N13152, N3999);
nor NOR2 (N13154, N13142, N11522);
and AND4 (N13155, N13153, N3266, N4436, N8605);
nand NAND3 (N13156, N13130, N12278, N1179);
or OR2 (N13157, N13148, N2046);
not NOT1 (N13158, N13138);
not NOT1 (N13159, N13156);
nand NAND3 (N13160, N13151, N9846, N12058);
and AND3 (N13161, N13158, N1423, N12491);
xor XOR2 (N13162, N13161, N2675);
nor NOR4 (N13163, N13155, N5746, N4739, N12793);
nand NAND2 (N13164, N13150, N2298);
xor XOR2 (N13165, N13141, N1141);
nor NOR2 (N13166, N13134, N11787);
nand NAND4 (N13167, N13137, N1048, N1606, N8880);
nor NOR2 (N13168, N13167, N8829);
and AND2 (N13169, N13157, N9621);
and AND4 (N13170, N13163, N882, N4654, N1385);
xor XOR2 (N13171, N13165, N9920);
buf BUF1 (N13172, N13170);
xor XOR2 (N13173, N13162, N2766);
not NOT1 (N13174, N13154);
xor XOR2 (N13175, N13169, N9249);
not NOT1 (N13176, N13164);
or OR3 (N13177, N13175, N7643, N439);
nor NOR3 (N13178, N13160, N11191, N10183);
nand NAND2 (N13179, N13168, N7145);
or OR3 (N13180, N13172, N2054, N2102);
nand NAND4 (N13181, N13177, N8556, N3398, N3017);
xor XOR2 (N13182, N13180, N5632);
and AND3 (N13183, N13182, N12401, N4091);
nor NOR3 (N13184, N13176, N6814, N348);
xor XOR2 (N13185, N13178, N5430);
and AND4 (N13186, N13183, N2791, N3513, N6207);
xor XOR2 (N13187, N13159, N10075);
nor NOR3 (N13188, N13186, N945, N11034);
xor XOR2 (N13189, N13187, N358);
and AND2 (N13190, N13171, N11036);
buf BUF1 (N13191, N13174);
or OR2 (N13192, N13188, N420);
or OR3 (N13193, N13166, N5820, N1930);
and AND4 (N13194, N13184, N6864, N12746, N4580);
not NOT1 (N13195, N13185);
nor NOR4 (N13196, N13179, N8197, N12203, N5794);
nand NAND2 (N13197, N13195, N6864);
nand NAND2 (N13198, N13189, N8444);
xor XOR2 (N13199, N13194, N8210);
buf BUF1 (N13200, N13199);
buf BUF1 (N13201, N13200);
not NOT1 (N13202, N13193);
xor XOR2 (N13203, N13201, N6480);
nand NAND2 (N13204, N13197, N8945);
nand NAND2 (N13205, N13191, N5350);
nor NOR4 (N13206, N13181, N6810, N10002, N7318);
or OR2 (N13207, N13206, N5127);
or OR3 (N13208, N13202, N5671, N8555);
or OR3 (N13209, N13173, N7570, N3038);
and AND3 (N13210, N13196, N12459, N12330);
nor NOR3 (N13211, N13205, N7635, N10369);
not NOT1 (N13212, N13210);
buf BUF1 (N13213, N13192);
not NOT1 (N13214, N13203);
not NOT1 (N13215, N13198);
xor XOR2 (N13216, N13209, N8550);
and AND4 (N13217, N13207, N6927, N8591, N7740);
and AND3 (N13218, N13217, N4142, N11613);
nor NOR2 (N13219, N13216, N2705);
nor NOR4 (N13220, N13214, N6819, N11156, N9218);
or OR4 (N13221, N13212, N3433, N10322, N11566);
buf BUF1 (N13222, N13221);
and AND2 (N13223, N13208, N9175);
nand NAND4 (N13224, N13213, N4107, N4420, N10444);
buf BUF1 (N13225, N13224);
and AND3 (N13226, N13190, N7882, N654);
nor NOR4 (N13227, N13218, N812, N3102, N7395);
buf BUF1 (N13228, N13204);
buf BUF1 (N13229, N13225);
xor XOR2 (N13230, N13219, N6760);
nor NOR3 (N13231, N13222, N7301, N1003);
buf BUF1 (N13232, N13228);
nand NAND2 (N13233, N13211, N12332);
buf BUF1 (N13234, N13229);
nor NOR4 (N13235, N13215, N6802, N12792, N10971);
nor NOR3 (N13236, N13230, N3824, N4146);
xor XOR2 (N13237, N13234, N7651);
or OR4 (N13238, N13236, N5803, N5733, N10431);
buf BUF1 (N13239, N13233);
and AND4 (N13240, N13226, N8375, N4350, N12907);
nor NOR3 (N13241, N13220, N10016, N8608);
and AND2 (N13242, N13237, N13128);
and AND3 (N13243, N13235, N3857, N11181);
or OR2 (N13244, N13241, N12410);
or OR3 (N13245, N13227, N3313, N3508);
nand NAND4 (N13246, N13231, N10451, N2436, N9734);
and AND2 (N13247, N13243, N10174);
and AND4 (N13248, N13245, N275, N1920, N12135);
or OR4 (N13249, N13238, N5083, N12014, N185);
or OR3 (N13250, N13248, N13003, N2199);
not NOT1 (N13251, N13244);
nor NOR2 (N13252, N13247, N9335);
nand NAND4 (N13253, N13249, N5432, N6461, N10524);
nor NOR3 (N13254, N13242, N12108, N4154);
or OR2 (N13255, N13253, N6640);
xor XOR2 (N13256, N13251, N2832);
or OR3 (N13257, N13239, N5387, N11783);
or OR2 (N13258, N13255, N13224);
xor XOR2 (N13259, N13223, N4813);
and AND4 (N13260, N13256, N7505, N4016, N10029);
not NOT1 (N13261, N13232);
or OR2 (N13262, N13259, N2078);
nor NOR2 (N13263, N13262, N6925);
buf BUF1 (N13264, N13260);
nand NAND3 (N13265, N13264, N9278, N3509);
or OR3 (N13266, N13257, N7576, N4706);
nand NAND2 (N13267, N13250, N2980);
and AND4 (N13268, N13254, N8052, N1337, N11252);
xor XOR2 (N13269, N13263, N6637);
or OR2 (N13270, N13265, N9189);
nor NOR3 (N13271, N13261, N5385, N11495);
not NOT1 (N13272, N13270);
buf BUF1 (N13273, N13240);
buf BUF1 (N13274, N13273);
and AND4 (N13275, N13266, N4104, N10956, N1840);
nor NOR2 (N13276, N13268, N876);
xor XOR2 (N13277, N13267, N6326);
and AND2 (N13278, N13274, N5313);
or OR3 (N13279, N13275, N10300, N2252);
and AND2 (N13280, N13246, N7477);
or OR4 (N13281, N13280, N4136, N10167, N904);
or OR3 (N13282, N13252, N10568, N8265);
xor XOR2 (N13283, N13279, N13115);
or OR4 (N13284, N13258, N1208, N4259, N2322);
nand NAND2 (N13285, N13276, N4559);
and AND3 (N13286, N13284, N2698, N11372);
not NOT1 (N13287, N13271);
nand NAND4 (N13288, N13278, N168, N8091, N1242);
nor NOR4 (N13289, N13286, N3823, N10399, N8538);
not NOT1 (N13290, N13285);
buf BUF1 (N13291, N13272);
nor NOR3 (N13292, N13281, N695, N3935);
buf BUF1 (N13293, N13282);
not NOT1 (N13294, N13283);
nand NAND4 (N13295, N13292, N7389, N5597, N5290);
or OR4 (N13296, N13269, N7537, N13131, N3966);
not NOT1 (N13297, N13289);
nor NOR4 (N13298, N13296, N11293, N7169, N4388);
and AND2 (N13299, N13298, N11603);
or OR4 (N13300, N13291, N1200, N2259, N5168);
or OR3 (N13301, N13294, N1935, N11661);
not NOT1 (N13302, N13288);
not NOT1 (N13303, N13297);
not NOT1 (N13304, N13290);
buf BUF1 (N13305, N13293);
and AND2 (N13306, N13304, N2707);
not NOT1 (N13307, N13302);
nor NOR3 (N13308, N13307, N13024, N11313);
buf BUF1 (N13309, N13306);
and AND3 (N13310, N13299, N1179, N665);
or OR4 (N13311, N13295, N1741, N3668, N5152);
not NOT1 (N13312, N13311);
or OR3 (N13313, N13300, N1806, N3469);
xor XOR2 (N13314, N13313, N3568);
nand NAND2 (N13315, N13314, N1825);
nand NAND3 (N13316, N13312, N7237, N12969);
xor XOR2 (N13317, N13301, N4353);
not NOT1 (N13318, N13303);
and AND2 (N13319, N13310, N8760);
or OR4 (N13320, N13308, N5110, N1806, N8304);
not NOT1 (N13321, N13277);
buf BUF1 (N13322, N13319);
xor XOR2 (N13323, N13316, N4166);
xor XOR2 (N13324, N13305, N8159);
buf BUF1 (N13325, N13315);
xor XOR2 (N13326, N13325, N10704);
nand NAND3 (N13327, N13320, N7330, N3865);
not NOT1 (N13328, N13287);
xor XOR2 (N13329, N13323, N5435);
not NOT1 (N13330, N13329);
nand NAND4 (N13331, N13321, N11094, N3861, N4478);
xor XOR2 (N13332, N13327, N465);
nand NAND2 (N13333, N13317, N11988);
nand NAND2 (N13334, N13332, N3377);
not NOT1 (N13335, N13309);
nand NAND4 (N13336, N13335, N3734, N8901, N268);
and AND2 (N13337, N13324, N8337);
and AND3 (N13338, N13331, N355, N8998);
nand NAND2 (N13339, N13333, N6439);
not NOT1 (N13340, N13326);
buf BUF1 (N13341, N13337);
or OR4 (N13342, N13334, N3957, N9508, N10572);
nor NOR4 (N13343, N13339, N5381, N10303, N1661);
nand NAND4 (N13344, N13322, N8969, N5440, N6626);
nand NAND4 (N13345, N13336, N10268, N1484, N3023);
buf BUF1 (N13346, N13340);
nor NOR2 (N13347, N13328, N12776);
nand NAND2 (N13348, N13346, N10164);
buf BUF1 (N13349, N13330);
nand NAND3 (N13350, N13348, N774, N10365);
and AND2 (N13351, N13342, N6674);
nor NOR2 (N13352, N13351, N145);
xor XOR2 (N13353, N13345, N13326);
buf BUF1 (N13354, N13350);
not NOT1 (N13355, N13344);
xor XOR2 (N13356, N13347, N2516);
xor XOR2 (N13357, N13343, N3942);
nor NOR4 (N13358, N13341, N8932, N7745, N10293);
and AND4 (N13359, N13349, N11264, N2926, N3775);
not NOT1 (N13360, N13355);
xor XOR2 (N13361, N13354, N7478);
buf BUF1 (N13362, N13318);
buf BUF1 (N13363, N13358);
nand NAND3 (N13364, N13338, N6222, N6209);
nand NAND4 (N13365, N13363, N13129, N11923, N788);
xor XOR2 (N13366, N13365, N7123);
not NOT1 (N13367, N13359);
buf BUF1 (N13368, N13366);
nor NOR4 (N13369, N13357, N9933, N10753, N120);
buf BUF1 (N13370, N13353);
or OR2 (N13371, N13360, N8594);
buf BUF1 (N13372, N13361);
buf BUF1 (N13373, N13372);
nor NOR2 (N13374, N13362, N1238);
nor NOR2 (N13375, N13369, N9886);
or OR2 (N13376, N13375, N7932);
xor XOR2 (N13377, N13373, N1933);
and AND4 (N13378, N13364, N6209, N6688, N11050);
buf BUF1 (N13379, N13378);
xor XOR2 (N13380, N13367, N7270);
buf BUF1 (N13381, N13370);
nor NOR2 (N13382, N13374, N295);
not NOT1 (N13383, N13368);
xor XOR2 (N13384, N13380, N4633);
not NOT1 (N13385, N13379);
xor XOR2 (N13386, N13371, N9323);
nor NOR2 (N13387, N13382, N12824);
nand NAND4 (N13388, N13381, N2535, N6814, N7714);
nand NAND4 (N13389, N13388, N11840, N2044, N1426);
buf BUF1 (N13390, N13352);
or OR2 (N13391, N13385, N4522);
and AND3 (N13392, N13376, N10601, N10447);
not NOT1 (N13393, N13383);
nand NAND3 (N13394, N13393, N10396, N10993);
buf BUF1 (N13395, N13386);
and AND2 (N13396, N13395, N2255);
or OR3 (N13397, N13396, N10204, N8196);
nand NAND2 (N13398, N13356, N12616);
nand NAND2 (N13399, N13391, N5408);
nand NAND4 (N13400, N13397, N6287, N11428, N7779);
and AND4 (N13401, N13392, N8105, N1736, N12297);
buf BUF1 (N13402, N13377);
nor NOR3 (N13403, N13401, N9184, N12917);
not NOT1 (N13404, N13387);
xor XOR2 (N13405, N13390, N6676);
nand NAND4 (N13406, N13402, N3133, N6388, N4696);
nand NAND2 (N13407, N13399, N8801);
nor NOR4 (N13408, N13406, N407, N6195, N9480);
buf BUF1 (N13409, N13400);
nand NAND2 (N13410, N13403, N8196);
and AND3 (N13411, N13408, N716, N11343);
buf BUF1 (N13412, N13398);
nand NAND4 (N13413, N13411, N12518, N10466, N12239);
and AND3 (N13414, N13412, N7983, N10560);
nor NOR2 (N13415, N13404, N11790);
and AND2 (N13416, N13414, N7716);
nor NOR3 (N13417, N13384, N9285, N2790);
xor XOR2 (N13418, N13407, N3109);
nand NAND3 (N13419, N13389, N10681, N315);
not NOT1 (N13420, N13410);
or OR4 (N13421, N13419, N4366, N7104, N11092);
nand NAND2 (N13422, N13394, N1064);
or OR3 (N13423, N13409, N5842, N1280);
and AND4 (N13424, N13421, N10158, N12708, N6610);
buf BUF1 (N13425, N13420);
or OR4 (N13426, N13416, N3458, N9072, N8330);
or OR3 (N13427, N13426, N3885, N8939);
or OR3 (N13428, N13424, N2309, N3909);
nor NOR2 (N13429, N13428, N11370);
nor NOR2 (N13430, N13417, N9);
and AND2 (N13431, N13422, N2449);
nor NOR3 (N13432, N13423, N13036, N9095);
buf BUF1 (N13433, N13425);
nor NOR2 (N13434, N13427, N12703);
and AND2 (N13435, N13433, N3146);
and AND4 (N13436, N13418, N2981, N9875, N7743);
xor XOR2 (N13437, N13431, N7477);
nand NAND4 (N13438, N13405, N8579, N2143, N8096);
not NOT1 (N13439, N13430);
nor NOR4 (N13440, N13437, N12126, N5520, N11692);
or OR2 (N13441, N13440, N5369);
xor XOR2 (N13442, N13439, N2976);
buf BUF1 (N13443, N13436);
nand NAND3 (N13444, N13415, N5539, N12637);
and AND2 (N13445, N13432, N12769);
nand NAND4 (N13446, N13444, N1171, N6776, N8833);
nor NOR4 (N13447, N13413, N2238, N7170, N8154);
buf BUF1 (N13448, N13443);
and AND3 (N13449, N13448, N10517, N3234);
not NOT1 (N13450, N13447);
xor XOR2 (N13451, N13450, N8856);
nor NOR2 (N13452, N13445, N2748);
nor NOR2 (N13453, N13429, N9077);
xor XOR2 (N13454, N13442, N10796);
nand NAND2 (N13455, N13435, N9898);
nand NAND4 (N13456, N13438, N12132, N12009, N8414);
xor XOR2 (N13457, N13454, N2822);
and AND4 (N13458, N13446, N12384, N3634, N6657);
not NOT1 (N13459, N13455);
xor XOR2 (N13460, N13456, N6367);
or OR4 (N13461, N13449, N6744, N4084, N12135);
xor XOR2 (N13462, N13460, N7445);
xor XOR2 (N13463, N13458, N4871);
not NOT1 (N13464, N13452);
not NOT1 (N13465, N13464);
or OR2 (N13466, N13434, N9585);
nor NOR3 (N13467, N13459, N11696, N4564);
xor XOR2 (N13468, N13467, N859);
and AND4 (N13469, N13457, N9547, N13384, N13116);
buf BUF1 (N13470, N13463);
nand NAND4 (N13471, N13469, N10738, N6192, N8227);
buf BUF1 (N13472, N13451);
and AND3 (N13473, N13470, N2593, N7839);
not NOT1 (N13474, N13468);
xor XOR2 (N13475, N13474, N9769);
not NOT1 (N13476, N13466);
not NOT1 (N13477, N13461);
nor NOR3 (N13478, N13477, N6576, N11360);
not NOT1 (N13479, N13453);
or OR3 (N13480, N13479, N13460, N6305);
nor NOR3 (N13481, N13480, N1398, N12155);
nor NOR2 (N13482, N13471, N7585);
xor XOR2 (N13483, N13482, N8690);
not NOT1 (N13484, N13478);
not NOT1 (N13485, N13465);
and AND3 (N13486, N13441, N7353, N2490);
xor XOR2 (N13487, N13476, N12886);
nand NAND4 (N13488, N13462, N37, N10213, N12266);
not NOT1 (N13489, N13488);
or OR4 (N13490, N13485, N3772, N13438, N5386);
xor XOR2 (N13491, N13481, N2260);
not NOT1 (N13492, N13484);
xor XOR2 (N13493, N13489, N8855);
buf BUF1 (N13494, N13473);
or OR3 (N13495, N13472, N7503, N6724);
and AND4 (N13496, N13494, N9776, N12674, N9745);
and AND3 (N13497, N13496, N3159, N11109);
nor NOR3 (N13498, N13475, N11111, N8988);
nor NOR3 (N13499, N13497, N573, N986);
not NOT1 (N13500, N13493);
nor NOR4 (N13501, N13498, N8838, N8294, N3114);
or OR4 (N13502, N13500, N4498, N958, N117);
nand NAND3 (N13503, N13483, N7262, N1815);
nand NAND2 (N13504, N13492, N9346);
nand NAND2 (N13505, N13491, N7072);
buf BUF1 (N13506, N13490);
buf BUF1 (N13507, N13486);
nand NAND3 (N13508, N13505, N286, N781);
nand NAND2 (N13509, N13503, N10115);
or OR3 (N13510, N13499, N1230, N6635);
or OR4 (N13511, N13510, N9438, N11370, N7161);
nand NAND2 (N13512, N13501, N11534);
nand NAND3 (N13513, N13509, N1398, N2563);
not NOT1 (N13514, N13512);
xor XOR2 (N13515, N13506, N5627);
or OR4 (N13516, N13487, N3816, N12809, N10960);
buf BUF1 (N13517, N13513);
nor NOR3 (N13518, N13516, N6662, N6932);
nor NOR2 (N13519, N13502, N9103);
or OR4 (N13520, N13507, N8701, N1925, N5779);
nand NAND4 (N13521, N13508, N4312, N1494, N10000);
not NOT1 (N13522, N13504);
and AND2 (N13523, N13522, N6958);
nor NOR2 (N13524, N13518, N9455);
or OR3 (N13525, N13511, N7431, N4305);
nand NAND2 (N13526, N13524, N11319);
buf BUF1 (N13527, N13520);
xor XOR2 (N13528, N13523, N6732);
nand NAND2 (N13529, N13521, N1057);
buf BUF1 (N13530, N13527);
nor NOR4 (N13531, N13526, N3028, N1403, N13096);
and AND3 (N13532, N13517, N5452, N3314);
and AND4 (N13533, N13531, N4738, N10470, N729);
not NOT1 (N13534, N13528);
buf BUF1 (N13535, N13525);
not NOT1 (N13536, N13535);
not NOT1 (N13537, N13515);
nor NOR4 (N13538, N13534, N3563, N9257, N13415);
nor NOR2 (N13539, N13533, N7827);
nand NAND3 (N13540, N13529, N6242, N8780);
or OR2 (N13541, N13519, N10413);
or OR4 (N13542, N13514, N12120, N12809, N5712);
xor XOR2 (N13543, N13538, N13227);
and AND3 (N13544, N13537, N5272, N1245);
nand NAND2 (N13545, N13542, N12637);
or OR3 (N13546, N13532, N11896, N5048);
not NOT1 (N13547, N13495);
xor XOR2 (N13548, N13540, N9751);
xor XOR2 (N13549, N13547, N9347);
nor NOR2 (N13550, N13541, N514);
not NOT1 (N13551, N13543);
and AND3 (N13552, N13539, N1990, N8885);
not NOT1 (N13553, N13548);
nand NAND2 (N13554, N13551, N8514);
or OR2 (N13555, N13544, N3124);
nand NAND3 (N13556, N13530, N2485, N10063);
not NOT1 (N13557, N13549);
buf BUF1 (N13558, N13553);
nand NAND3 (N13559, N13555, N11725, N1308);
xor XOR2 (N13560, N13550, N3657);
xor XOR2 (N13561, N13546, N1819);
or OR2 (N13562, N13561, N340);
nand NAND4 (N13563, N13545, N7514, N111, N6696);
or OR2 (N13564, N13558, N12909);
nand NAND4 (N13565, N13536, N10877, N2773, N765);
and AND4 (N13566, N13562, N10031, N2035, N8450);
nand NAND2 (N13567, N13565, N7703);
nor NOR4 (N13568, N13559, N28, N6786, N1441);
xor XOR2 (N13569, N13568, N10844);
nand NAND2 (N13570, N13567, N5870);
nand NAND2 (N13571, N13556, N6305);
nor NOR3 (N13572, N13557, N12605, N11394);
buf BUF1 (N13573, N13552);
or OR3 (N13574, N13572, N9395, N3539);
or OR4 (N13575, N13563, N12384, N1793, N6535);
not NOT1 (N13576, N13571);
or OR2 (N13577, N13573, N3177);
or OR3 (N13578, N13564, N2047, N3936);
buf BUF1 (N13579, N13575);
and AND3 (N13580, N13574, N6462, N8181);
nor NOR4 (N13581, N13579, N6016, N7749, N679);
xor XOR2 (N13582, N13570, N9846);
and AND3 (N13583, N13577, N12733, N3950);
nor NOR2 (N13584, N13580, N7533);
xor XOR2 (N13585, N13566, N10908);
and AND2 (N13586, N13554, N1144);
xor XOR2 (N13587, N13560, N785);
or OR3 (N13588, N13585, N4773, N2798);
not NOT1 (N13589, N13584);
or OR2 (N13590, N13581, N2103);
and AND3 (N13591, N13586, N10928, N534);
nand NAND4 (N13592, N13569, N10798, N7561, N9073);
nand NAND4 (N13593, N13592, N5669, N12932, N8574);
not NOT1 (N13594, N13589);
nand NAND2 (N13595, N13593, N11436);
and AND4 (N13596, N13582, N8700, N5441, N10023);
or OR3 (N13597, N13576, N9438, N4926);
xor XOR2 (N13598, N13583, N7202);
or OR2 (N13599, N13597, N3920);
nand NAND3 (N13600, N13595, N2815, N9345);
and AND3 (N13601, N13587, N11737, N13571);
nor NOR3 (N13602, N13590, N5826, N8671);
or OR4 (N13603, N13600, N6531, N8036, N4095);
or OR4 (N13604, N13588, N12856, N2577, N12255);
nand NAND4 (N13605, N13601, N8562, N67, N9216);
nor NOR2 (N13606, N13596, N1985);
not NOT1 (N13607, N13599);
or OR2 (N13608, N13591, N6636);
not NOT1 (N13609, N13578);
and AND2 (N13610, N13605, N8622);
nand NAND3 (N13611, N13610, N11669, N7702);
buf BUF1 (N13612, N13604);
and AND4 (N13613, N13608, N6728, N1514, N3225);
xor XOR2 (N13614, N13611, N5807);
nand NAND3 (N13615, N13594, N7995, N10296);
nand NAND2 (N13616, N13607, N9516);
and AND2 (N13617, N13613, N12569);
xor XOR2 (N13618, N13615, N7693);
xor XOR2 (N13619, N13616, N2688);
not NOT1 (N13620, N13618);
nor NOR3 (N13621, N13619, N7746, N3849);
nand NAND3 (N13622, N13603, N8744, N13473);
xor XOR2 (N13623, N13612, N10164);
and AND2 (N13624, N13598, N6907);
xor XOR2 (N13625, N13624, N11448);
nor NOR4 (N13626, N13622, N11178, N12425, N2764);
xor XOR2 (N13627, N13625, N10144);
or OR4 (N13628, N13626, N5715, N1435, N2688);
buf BUF1 (N13629, N13621);
nor NOR2 (N13630, N13617, N7078);
nand NAND4 (N13631, N13630, N7610, N7854, N12757);
buf BUF1 (N13632, N13629);
xor XOR2 (N13633, N13620, N8849);
xor XOR2 (N13634, N13614, N5186);
nand NAND3 (N13635, N13628, N5627, N8728);
not NOT1 (N13636, N13633);
buf BUF1 (N13637, N13631);
or OR2 (N13638, N13606, N12459);
buf BUF1 (N13639, N13636);
and AND4 (N13640, N13632, N6325, N4461, N8405);
nor NOR3 (N13641, N13602, N11405, N4415);
buf BUF1 (N13642, N13641);
and AND4 (N13643, N13640, N13261, N5821, N5363);
nand NAND2 (N13644, N13635, N238);
nor NOR3 (N13645, N13644, N4359, N2479);
nor NOR2 (N13646, N13638, N3440);
not NOT1 (N13647, N13645);
not NOT1 (N13648, N13643);
not NOT1 (N13649, N13637);
or OR2 (N13650, N13634, N10384);
xor XOR2 (N13651, N13639, N11888);
and AND4 (N13652, N13642, N7363, N5432, N4842);
and AND3 (N13653, N13646, N5194, N10094);
xor XOR2 (N13654, N13653, N6100);
buf BUF1 (N13655, N13623);
nor NOR3 (N13656, N13627, N2997, N1312);
buf BUF1 (N13657, N13652);
and AND3 (N13658, N13657, N13376, N3051);
not NOT1 (N13659, N13650);
and AND2 (N13660, N13648, N7419);
and AND2 (N13661, N13647, N11471);
and AND3 (N13662, N13661, N12181, N12030);
nand NAND4 (N13663, N13649, N960, N613, N10159);
buf BUF1 (N13664, N13655);
not NOT1 (N13665, N13659);
and AND3 (N13666, N13665, N1106, N10514);
nor NOR2 (N13667, N13658, N233);
nand NAND4 (N13668, N13663, N2170, N10459, N4011);
or OR2 (N13669, N13667, N2797);
buf BUF1 (N13670, N13609);
or OR2 (N13671, N13669, N7460);
nand NAND3 (N13672, N13668, N2903, N4987);
nor NOR2 (N13673, N13666, N10671);
nand NAND3 (N13674, N13672, N5576, N13320);
xor XOR2 (N13675, N13662, N11177);
buf BUF1 (N13676, N13654);
not NOT1 (N13677, N13670);
xor XOR2 (N13678, N13651, N185);
xor XOR2 (N13679, N13677, N8268);
xor XOR2 (N13680, N13675, N709);
xor XOR2 (N13681, N13671, N6092);
buf BUF1 (N13682, N13673);
xor XOR2 (N13683, N13656, N5477);
buf BUF1 (N13684, N13664);
buf BUF1 (N13685, N13682);
nand NAND3 (N13686, N13680, N11051, N4560);
and AND3 (N13687, N13685, N12250, N10729);
and AND2 (N13688, N13684, N9069);
buf BUF1 (N13689, N13678);
not NOT1 (N13690, N13679);
or OR3 (N13691, N13687, N11720, N3312);
nor NOR2 (N13692, N13674, N5622);
nand NAND2 (N13693, N13690, N8141);
buf BUF1 (N13694, N13688);
buf BUF1 (N13695, N13689);
buf BUF1 (N13696, N13693);
buf BUF1 (N13697, N13686);
buf BUF1 (N13698, N13692);
or OR2 (N13699, N13697, N3749);
nand NAND4 (N13700, N13683, N11425, N5974, N405);
nand NAND2 (N13701, N13681, N3537);
or OR4 (N13702, N13694, N4123, N13009, N6020);
or OR4 (N13703, N13700, N5784, N10011, N10143);
nor NOR2 (N13704, N13701, N3656);
not NOT1 (N13705, N13698);
buf BUF1 (N13706, N13660);
buf BUF1 (N13707, N13704);
nor NOR4 (N13708, N13705, N5171, N4779, N257);
xor XOR2 (N13709, N13691, N5844);
xor XOR2 (N13710, N13676, N12126);
buf BUF1 (N13711, N13696);
not NOT1 (N13712, N13702);
nor NOR3 (N13713, N13695, N7153, N9615);
xor XOR2 (N13714, N13710, N5598);
and AND2 (N13715, N13712, N7363);
nor NOR3 (N13716, N13714, N1370, N12667);
or OR4 (N13717, N13716, N762, N9738, N647);
buf BUF1 (N13718, N13699);
not NOT1 (N13719, N13715);
buf BUF1 (N13720, N13708);
or OR4 (N13721, N13709, N6291, N8984, N5104);
or OR2 (N13722, N13706, N11221);
and AND3 (N13723, N13711, N11410, N7358);
nand NAND4 (N13724, N13718, N5388, N9085, N2641);
or OR4 (N13725, N13723, N1961, N8190, N10415);
nor NOR3 (N13726, N13707, N10820, N4520);
nand NAND2 (N13727, N13719, N7240);
nand NAND4 (N13728, N13720, N1445, N12886, N10461);
xor XOR2 (N13729, N13725, N3085);
nor NOR3 (N13730, N13724, N8730, N9098);
buf BUF1 (N13731, N13722);
xor XOR2 (N13732, N13730, N5917);
nand NAND2 (N13733, N13717, N12374);
nand NAND4 (N13734, N13728, N7190, N13472, N9992);
buf BUF1 (N13735, N13703);
not NOT1 (N13736, N13731);
and AND2 (N13737, N13733, N8459);
and AND2 (N13738, N13732, N9045);
buf BUF1 (N13739, N13735);
xor XOR2 (N13740, N13734, N8444);
nor NOR4 (N13741, N13738, N1095, N11931, N10941);
nor NOR3 (N13742, N13741, N4511, N2436);
and AND2 (N13743, N13726, N907);
xor XOR2 (N13744, N13740, N12027);
buf BUF1 (N13745, N13713);
nor NOR3 (N13746, N13739, N984, N8110);
nand NAND2 (N13747, N13727, N6210);
nand NAND2 (N13748, N13729, N10853);
or OR4 (N13749, N13747, N133, N5367, N11477);
nand NAND3 (N13750, N13746, N3080, N11655);
nand NAND4 (N13751, N13749, N4742, N5918, N7999);
or OR4 (N13752, N13721, N1974, N10056, N2297);
and AND3 (N13753, N13752, N765, N5845);
and AND4 (N13754, N13745, N6901, N6271, N8330);
not NOT1 (N13755, N13750);
xor XOR2 (N13756, N13743, N1032);
or OR3 (N13757, N13753, N4707, N2151);
not NOT1 (N13758, N13742);
nor NOR3 (N13759, N13755, N13665, N429);
buf BUF1 (N13760, N13737);
nand NAND2 (N13761, N13754, N690);
nor NOR3 (N13762, N13759, N9709, N10819);
and AND4 (N13763, N13758, N10305, N6822, N7447);
not NOT1 (N13764, N13744);
nand NAND3 (N13765, N13764, N12496, N10534);
nor NOR4 (N13766, N13760, N7226, N1181, N93);
nor NOR3 (N13767, N13757, N2815, N9338);
nand NAND4 (N13768, N13761, N7950, N13171, N9105);
or OR2 (N13769, N13767, N10295);
and AND4 (N13770, N13765, N1557, N6307, N12400);
buf BUF1 (N13771, N13770);
or OR3 (N13772, N13771, N9217, N8276);
and AND3 (N13773, N13756, N5893, N9637);
and AND4 (N13774, N13772, N10710, N9589, N7634);
and AND3 (N13775, N13751, N2104, N5657);
xor XOR2 (N13776, N13775, N2109);
or OR3 (N13777, N13736, N9354, N5767);
nand NAND2 (N13778, N13762, N2769);
nor NOR4 (N13779, N13778, N13029, N6940, N6851);
and AND4 (N13780, N13774, N13108, N12129, N11580);
xor XOR2 (N13781, N13773, N6760);
buf BUF1 (N13782, N13766);
buf BUF1 (N13783, N13768);
not NOT1 (N13784, N13777);
and AND3 (N13785, N13782, N2473, N795);
nand NAND2 (N13786, N13784, N1398);
or OR3 (N13787, N13786, N8872, N4270);
xor XOR2 (N13788, N13748, N13274);
not NOT1 (N13789, N13779);
nor NOR2 (N13790, N13789, N7780);
nand NAND2 (N13791, N13776, N6020);
not NOT1 (N13792, N13785);
not NOT1 (N13793, N13787);
nor NOR4 (N13794, N13792, N7550, N4302, N6768);
not NOT1 (N13795, N13769);
nand NAND4 (N13796, N13791, N6609, N2496, N11842);
nor NOR2 (N13797, N13794, N6512);
nand NAND4 (N13798, N13790, N1839, N10528, N7288);
and AND4 (N13799, N13783, N2471, N5129, N2694);
not NOT1 (N13800, N13781);
or OR2 (N13801, N13799, N10934);
or OR4 (N13802, N13780, N6269, N9813, N11051);
not NOT1 (N13803, N13797);
nand NAND3 (N13804, N13788, N12328, N5393);
nand NAND3 (N13805, N13795, N1080, N11149);
buf BUF1 (N13806, N13804);
nor NOR3 (N13807, N13803, N13223, N2830);
and AND2 (N13808, N13796, N13690);
not NOT1 (N13809, N13805);
nand NAND2 (N13810, N13807, N839);
and AND4 (N13811, N13798, N9174, N6882, N2122);
nor NOR4 (N13812, N13800, N7497, N11247, N6146);
buf BUF1 (N13813, N13811);
and AND3 (N13814, N13802, N11296, N9807);
not NOT1 (N13815, N13763);
and AND2 (N13816, N13801, N3646);
not NOT1 (N13817, N13812);
buf BUF1 (N13818, N13793);
xor XOR2 (N13819, N13808, N3989);
xor XOR2 (N13820, N13815, N12115);
not NOT1 (N13821, N13818);
and AND3 (N13822, N13806, N11203, N2467);
nand NAND3 (N13823, N13814, N10087, N9369);
nor NOR4 (N13824, N13813, N2275, N323, N11215);
not NOT1 (N13825, N13823);
and AND3 (N13826, N13820, N5431, N174);
and AND2 (N13827, N13809, N6063);
and AND3 (N13828, N13810, N5620, N12296);
not NOT1 (N13829, N13819);
buf BUF1 (N13830, N13828);
buf BUF1 (N13831, N13827);
buf BUF1 (N13832, N13831);
nand NAND2 (N13833, N13830, N2521);
or OR3 (N13834, N13821, N7934, N4029);
and AND2 (N13835, N13817, N1133);
and AND2 (N13836, N13816, N10789);
and AND2 (N13837, N13834, N13502);
and AND4 (N13838, N13833, N13447, N5254, N4824);
or OR3 (N13839, N13832, N4074, N10568);
not NOT1 (N13840, N13826);
buf BUF1 (N13841, N13824);
or OR2 (N13842, N13822, N9913);
or OR4 (N13843, N13836, N10952, N2178, N13163);
buf BUF1 (N13844, N13837);
not NOT1 (N13845, N13841);
or OR2 (N13846, N13843, N1817);
nand NAND3 (N13847, N13839, N8369, N4325);
and AND4 (N13848, N13846, N441, N10144, N9160);
and AND2 (N13849, N13825, N5999);
buf BUF1 (N13850, N13848);
nand NAND2 (N13851, N13838, N4520);
xor XOR2 (N13852, N13844, N5044);
buf BUF1 (N13853, N13840);
and AND3 (N13854, N13850, N1913, N8794);
not NOT1 (N13855, N13853);
not NOT1 (N13856, N13835);
and AND3 (N13857, N13856, N10372, N2476);
nor NOR2 (N13858, N13855, N11396);
xor XOR2 (N13859, N13842, N7311);
not NOT1 (N13860, N13849);
buf BUF1 (N13861, N13854);
not NOT1 (N13862, N13858);
and AND3 (N13863, N13851, N13387, N8583);
xor XOR2 (N13864, N13852, N2565);
nand NAND2 (N13865, N13847, N9010);
buf BUF1 (N13866, N13862);
xor XOR2 (N13867, N13829, N227);
nand NAND3 (N13868, N13861, N1356, N7229);
not NOT1 (N13869, N13857);
or OR4 (N13870, N13859, N4671, N4490, N5588);
nor NOR4 (N13871, N13866, N12438, N8771, N1009);
xor XOR2 (N13872, N13865, N13174);
and AND3 (N13873, N13869, N6168, N4599);
or OR2 (N13874, N13873, N4765);
and AND3 (N13875, N13863, N6335, N3359);
or OR2 (N13876, N13874, N3398);
nand NAND3 (N13877, N13871, N5352, N7020);
not NOT1 (N13878, N13870);
nor NOR4 (N13879, N13878, N5400, N1183, N4511);
or OR3 (N13880, N13868, N8806, N1767);
buf BUF1 (N13881, N13880);
nand NAND4 (N13882, N13881, N12015, N5389, N170);
xor XOR2 (N13883, N13882, N6349);
or OR2 (N13884, N13879, N649);
nor NOR2 (N13885, N13864, N13411);
nand NAND3 (N13886, N13883, N10553, N6953);
and AND3 (N13887, N13872, N6056, N9155);
nor NOR2 (N13888, N13875, N2194);
or OR3 (N13889, N13887, N9692, N6331);
xor XOR2 (N13890, N13876, N11997);
not NOT1 (N13891, N13889);
nor NOR3 (N13892, N13888, N2064, N2818);
nand NAND3 (N13893, N13891, N11184, N7847);
and AND3 (N13894, N13860, N167, N4066);
nor NOR2 (N13895, N13884, N8797);
or OR4 (N13896, N13893, N5186, N13545, N13608);
buf BUF1 (N13897, N13886);
not NOT1 (N13898, N13877);
not NOT1 (N13899, N13897);
nor NOR2 (N13900, N13867, N7262);
buf BUF1 (N13901, N13900);
nor NOR3 (N13902, N13896, N5623, N4209);
nand NAND4 (N13903, N13894, N7355, N7396, N7673);
not NOT1 (N13904, N13898);
and AND3 (N13905, N13895, N6019, N1528);
and AND3 (N13906, N13885, N8227, N10150);
xor XOR2 (N13907, N13845, N9841);
nor NOR2 (N13908, N13890, N10198);
not NOT1 (N13909, N13907);
or OR2 (N13910, N13903, N2284);
xor XOR2 (N13911, N13909, N601);
or OR2 (N13912, N13911, N13491);
and AND3 (N13913, N13892, N12956, N13141);
xor XOR2 (N13914, N13908, N7826);
nor NOR3 (N13915, N13906, N8472, N2615);
nand NAND4 (N13916, N13914, N408, N4418, N3370);
nand NAND4 (N13917, N13913, N7476, N10842, N11377);
not NOT1 (N13918, N13905);
nand NAND2 (N13919, N13904, N9533);
and AND4 (N13920, N13910, N1978, N3169, N8282);
or OR2 (N13921, N13912, N8586);
or OR4 (N13922, N13916, N5417, N8643, N10101);
not NOT1 (N13923, N13920);
xor XOR2 (N13924, N13902, N7996);
buf BUF1 (N13925, N13923);
not NOT1 (N13926, N13924);
buf BUF1 (N13927, N13925);
not NOT1 (N13928, N13918);
buf BUF1 (N13929, N13927);
or OR4 (N13930, N13901, N8270, N291, N7425);
or OR3 (N13931, N13926, N8700, N3598);
nor NOR4 (N13932, N13931, N9009, N8915, N814);
and AND2 (N13933, N13899, N3343);
and AND4 (N13934, N13917, N742, N6432, N13809);
nand NAND2 (N13935, N13933, N1777);
nand NAND4 (N13936, N13929, N9943, N2446, N12077);
not NOT1 (N13937, N13935);
and AND2 (N13938, N13934, N3782);
buf BUF1 (N13939, N13932);
or OR3 (N13940, N13921, N9003, N1276);
and AND2 (N13941, N13915, N10267);
nand NAND3 (N13942, N13936, N9781, N5415);
nand NAND4 (N13943, N13941, N10730, N4128, N9035);
buf BUF1 (N13944, N13930);
buf BUF1 (N13945, N13943);
not NOT1 (N13946, N13940);
not NOT1 (N13947, N13946);
nand NAND4 (N13948, N13937, N13738, N4345, N13300);
buf BUF1 (N13949, N13947);
nor NOR2 (N13950, N13939, N1209);
and AND3 (N13951, N13945, N5901, N2143);
nand NAND4 (N13952, N13928, N9335, N4125, N7008);
buf BUF1 (N13953, N13952);
xor XOR2 (N13954, N13922, N4360);
nand NAND4 (N13955, N13944, N9083, N13370, N3042);
xor XOR2 (N13956, N13954, N2633);
or OR4 (N13957, N13942, N5575, N225, N4816);
not NOT1 (N13958, N13948);
xor XOR2 (N13959, N13957, N6108);
and AND4 (N13960, N13956, N5326, N4930, N7550);
not NOT1 (N13961, N13949);
nor NOR2 (N13962, N13960, N2621);
nor NOR2 (N13963, N13950, N2057);
buf BUF1 (N13964, N13963);
or OR3 (N13965, N13961, N8595, N2143);
nand NAND2 (N13966, N13953, N6059);
buf BUF1 (N13967, N13938);
and AND4 (N13968, N13962, N10890, N1632, N1198);
nand NAND4 (N13969, N13968, N2047, N12321, N12432);
or OR3 (N13970, N13966, N4445, N174);
or OR4 (N13971, N13958, N13570, N1933, N2957);
buf BUF1 (N13972, N13919);
nand NAND2 (N13973, N13965, N8093);
nor NOR3 (N13974, N13971, N7665, N10441);
buf BUF1 (N13975, N13970);
and AND4 (N13976, N13973, N8757, N6680, N10896);
buf BUF1 (N13977, N13951);
xor XOR2 (N13978, N13974, N8292);
and AND3 (N13979, N13959, N3237, N12657);
buf BUF1 (N13980, N13972);
not NOT1 (N13981, N13977);
xor XOR2 (N13982, N13978, N4136);
buf BUF1 (N13983, N13982);
nor NOR3 (N13984, N13967, N6592, N12152);
not NOT1 (N13985, N13964);
not NOT1 (N13986, N13955);
buf BUF1 (N13987, N13975);
buf BUF1 (N13988, N13981);
or OR4 (N13989, N13988, N2050, N4503, N9211);
and AND3 (N13990, N13980, N2918, N10825);
nor NOR2 (N13991, N13989, N11835);
xor XOR2 (N13992, N13985, N4188);
xor XOR2 (N13993, N13986, N11478);
buf BUF1 (N13994, N13983);
or OR2 (N13995, N13991, N1978);
and AND4 (N13996, N13987, N7918, N11545, N1128);
xor XOR2 (N13997, N13984, N5398);
xor XOR2 (N13998, N13979, N5592);
xor XOR2 (N13999, N13996, N7087);
xor XOR2 (N14000, N13994, N2573);
xor XOR2 (N14001, N13969, N1492);
or OR2 (N14002, N14000, N8060);
nor NOR4 (N14003, N13992, N8593, N7972, N4976);
nor NOR4 (N14004, N13990, N5406, N4585, N2397);
or OR3 (N14005, N14002, N10716, N363);
buf BUF1 (N14006, N14001);
or OR4 (N14007, N14006, N9623, N1871, N2017);
xor XOR2 (N14008, N13998, N5565);
and AND2 (N14009, N14007, N1293);
nand NAND4 (N14010, N13976, N9701, N2557, N2949);
not NOT1 (N14011, N13995);
nor NOR4 (N14012, N14009, N6042, N1425, N13771);
and AND2 (N14013, N14012, N8009);
or OR2 (N14014, N13999, N6997);
nor NOR2 (N14015, N14014, N8622);
or OR4 (N14016, N14015, N8095, N8751, N5676);
xor XOR2 (N14017, N13993, N10300);
buf BUF1 (N14018, N14010);
nor NOR3 (N14019, N14013, N9082, N9133);
or OR4 (N14020, N14003, N725, N563, N4809);
nand NAND3 (N14021, N14005, N5341, N9076);
buf BUF1 (N14022, N14008);
or OR2 (N14023, N14020, N9538);
xor XOR2 (N14024, N14018, N12485);
and AND4 (N14025, N14019, N2900, N13546, N7046);
not NOT1 (N14026, N14023);
and AND2 (N14027, N14017, N3876);
or OR2 (N14028, N14011, N5869);
and AND2 (N14029, N14022, N264);
or OR2 (N14030, N14026, N2371);
nand NAND2 (N14031, N13997, N555);
and AND4 (N14032, N14029, N13646, N828, N10844);
nor NOR3 (N14033, N14004, N7338, N2845);
nor NOR2 (N14034, N14027, N12802);
buf BUF1 (N14035, N14032);
not NOT1 (N14036, N14025);
not NOT1 (N14037, N14034);
nand NAND2 (N14038, N14024, N13933);
or OR4 (N14039, N14021, N2416, N10511, N1654);
nand NAND4 (N14040, N14035, N9976, N4810, N5241);
not NOT1 (N14041, N14037);
and AND2 (N14042, N14039, N6027);
or OR2 (N14043, N14031, N8822);
nor NOR2 (N14044, N14036, N9886);
nand NAND3 (N14045, N14038, N12849, N12362);
buf BUF1 (N14046, N14041);
or OR2 (N14047, N14040, N4953);
nand NAND2 (N14048, N14028, N14008);
not NOT1 (N14049, N14042);
or OR3 (N14050, N14043, N8574, N11179);
nand NAND2 (N14051, N14048, N4881);
and AND4 (N14052, N14033, N5681, N5955, N12360);
xor XOR2 (N14053, N14045, N8510);
nor NOR2 (N14054, N14049, N9005);
buf BUF1 (N14055, N14054);
nor NOR2 (N14056, N14046, N6891);
not NOT1 (N14057, N14052);
buf BUF1 (N14058, N14050);
xor XOR2 (N14059, N14058, N2924);
or OR4 (N14060, N14055, N8407, N13122, N12616);
nand NAND3 (N14061, N14059, N12807, N9756);
nor NOR3 (N14062, N14053, N9261, N12343);
xor XOR2 (N14063, N14051, N2299);
xor XOR2 (N14064, N14060, N9631);
nand NAND3 (N14065, N14061, N921, N4235);
nand NAND2 (N14066, N14057, N9537);
xor XOR2 (N14067, N14066, N11027);
or OR2 (N14068, N14016, N12574);
nor NOR2 (N14069, N14030, N10366);
not NOT1 (N14070, N14067);
not NOT1 (N14071, N14047);
nand NAND4 (N14072, N14071, N13661, N7298, N9202);
or OR3 (N14073, N14062, N3759, N7227);
not NOT1 (N14074, N14064);
xor XOR2 (N14075, N14068, N10358);
buf BUF1 (N14076, N14044);
nand NAND3 (N14077, N14063, N9563, N5185);
and AND4 (N14078, N14076, N12700, N9347, N10060);
not NOT1 (N14079, N14077);
not NOT1 (N14080, N14070);
not NOT1 (N14081, N14075);
or OR4 (N14082, N14078, N11849, N14018, N11891);
or OR2 (N14083, N14056, N8794);
xor XOR2 (N14084, N14082, N3448);
or OR3 (N14085, N14072, N8422, N12383);
nand NAND4 (N14086, N14074, N13171, N6323, N12516);
nor NOR3 (N14087, N14080, N5311, N14033);
and AND2 (N14088, N14085, N10967);
or OR2 (N14089, N14065, N2453);
or OR3 (N14090, N14069, N6129, N13921);
and AND2 (N14091, N14083, N6678);
xor XOR2 (N14092, N14073, N13420);
nor NOR2 (N14093, N14088, N13586);
not NOT1 (N14094, N14091);
nand NAND3 (N14095, N14092, N7284, N10135);
or OR3 (N14096, N14094, N13470, N12601);
nor NOR2 (N14097, N14079, N12130);
nand NAND2 (N14098, N14093, N3486);
not NOT1 (N14099, N14086);
nor NOR4 (N14100, N14084, N10617, N5158, N7815);
not NOT1 (N14101, N14089);
not NOT1 (N14102, N14090);
nor NOR4 (N14103, N14099, N5161, N9956, N3286);
buf BUF1 (N14104, N14100);
or OR2 (N14105, N14087, N12878);
nand NAND4 (N14106, N14105, N3857, N7117, N4383);
buf BUF1 (N14107, N14104);
xor XOR2 (N14108, N14081, N11066);
buf BUF1 (N14109, N14098);
and AND3 (N14110, N14103, N12315, N954);
or OR2 (N14111, N14097, N11934);
nand NAND4 (N14112, N14109, N12949, N11232, N1779);
or OR4 (N14113, N14107, N288, N6799, N6434);
or OR2 (N14114, N14106, N701);
not NOT1 (N14115, N14113);
or OR3 (N14116, N14096, N1935, N11539);
xor XOR2 (N14117, N14108, N2196);
buf BUF1 (N14118, N14114);
and AND2 (N14119, N14102, N425);
xor XOR2 (N14120, N14117, N5992);
not NOT1 (N14121, N14101);
nand NAND4 (N14122, N14118, N13054, N12162, N4618);
not NOT1 (N14123, N14110);
and AND2 (N14124, N14123, N4);
xor XOR2 (N14125, N14116, N7371);
or OR3 (N14126, N14124, N584, N5825);
or OR3 (N14127, N14122, N12981, N6121);
nand NAND4 (N14128, N14112, N11908, N756, N12998);
xor XOR2 (N14129, N14119, N13089);
xor XOR2 (N14130, N14111, N7456);
not NOT1 (N14131, N14129);
nand NAND4 (N14132, N14130, N10762, N7731, N7251);
nor NOR2 (N14133, N14131, N1363);
nand NAND4 (N14134, N14127, N10163, N3761, N11882);
xor XOR2 (N14135, N14115, N2935);
nand NAND2 (N14136, N14133, N4857);
not NOT1 (N14137, N14125);
or OR4 (N14138, N14121, N12539, N12424, N10530);
nor NOR4 (N14139, N14138, N7133, N11409, N5614);
nor NOR4 (N14140, N14136, N12893, N14080, N3207);
and AND3 (N14141, N14132, N1547, N3169);
xor XOR2 (N14142, N14139, N12548);
xor XOR2 (N14143, N14142, N5014);
or OR3 (N14144, N14095, N12304, N1225);
xor XOR2 (N14145, N14134, N690);
buf BUF1 (N14146, N14135);
nor NOR3 (N14147, N14145, N5030, N1602);
not NOT1 (N14148, N14144);
and AND4 (N14149, N14120, N2068, N3255, N12175);
xor XOR2 (N14150, N14126, N6008);
nand NAND3 (N14151, N14150, N11263, N716);
nand NAND4 (N14152, N14141, N1223, N10860, N10099);
and AND2 (N14153, N14147, N13582);
nand NAND2 (N14154, N14149, N11751);
buf BUF1 (N14155, N14140);
and AND2 (N14156, N14137, N5479);
or OR2 (N14157, N14151, N9772);
nor NOR2 (N14158, N14128, N13367);
nand NAND2 (N14159, N14156, N12999);
or OR2 (N14160, N14158, N415);
xor XOR2 (N14161, N14157, N6347);
and AND3 (N14162, N14155, N423, N3936);
and AND3 (N14163, N14146, N13772, N8680);
not NOT1 (N14164, N14143);
and AND2 (N14165, N14162, N3897);
xor XOR2 (N14166, N14161, N7158);
or OR3 (N14167, N14152, N9447, N6676);
not NOT1 (N14168, N14148);
not NOT1 (N14169, N14166);
buf BUF1 (N14170, N14160);
xor XOR2 (N14171, N14159, N7545);
nand NAND2 (N14172, N14171, N14120);
nor NOR2 (N14173, N14153, N8828);
nor NOR3 (N14174, N14168, N982, N6424);
or OR3 (N14175, N14174, N11894, N893);
not NOT1 (N14176, N14175);
not NOT1 (N14177, N14163);
not NOT1 (N14178, N14176);
and AND4 (N14179, N14167, N3841, N6571, N1917);
nand NAND2 (N14180, N14170, N5833);
nand NAND4 (N14181, N14180, N5234, N14020, N7321);
not NOT1 (N14182, N14164);
not NOT1 (N14183, N14169);
buf BUF1 (N14184, N14172);
nor NOR3 (N14185, N14183, N2613, N5234);
nor NOR2 (N14186, N14165, N5081);
xor XOR2 (N14187, N14173, N13071);
and AND2 (N14188, N14187, N188);
buf BUF1 (N14189, N14185);
xor XOR2 (N14190, N14182, N3606);
xor XOR2 (N14191, N14190, N11712);
or OR3 (N14192, N14177, N10540, N1198);
and AND3 (N14193, N14188, N1125, N10685);
nor NOR3 (N14194, N14193, N1255, N4398);
buf BUF1 (N14195, N14186);
or OR3 (N14196, N14192, N10503, N7295);
nand NAND4 (N14197, N14189, N4271, N3607, N3761);
nor NOR2 (N14198, N14178, N8586);
xor XOR2 (N14199, N14196, N13415);
xor XOR2 (N14200, N14199, N4611);
or OR4 (N14201, N14179, N10340, N9998, N7463);
xor XOR2 (N14202, N14181, N11322);
not NOT1 (N14203, N14201);
not NOT1 (N14204, N14197);
nand NAND3 (N14205, N14203, N240, N7246);
or OR3 (N14206, N14200, N1612, N3102);
and AND3 (N14207, N14194, N1953, N7132);
buf BUF1 (N14208, N14198);
xor XOR2 (N14209, N14154, N2347);
buf BUF1 (N14210, N14202);
not NOT1 (N14211, N14204);
xor XOR2 (N14212, N14211, N4227);
nand NAND3 (N14213, N14195, N4770, N9348);
or OR3 (N14214, N14213, N6407, N1726);
and AND2 (N14215, N14212, N6100);
nor NOR3 (N14216, N14207, N751, N13102);
buf BUF1 (N14217, N14210);
not NOT1 (N14218, N14217);
not NOT1 (N14219, N14206);
nand NAND4 (N14220, N14214, N13426, N2975, N8353);
not NOT1 (N14221, N14216);
buf BUF1 (N14222, N14220);
nand NAND2 (N14223, N14208, N5803);
xor XOR2 (N14224, N14184, N4838);
nand NAND3 (N14225, N14215, N11928, N13412);
or OR4 (N14226, N14209, N1834, N4485, N2637);
xor XOR2 (N14227, N14205, N10625);
and AND3 (N14228, N14226, N5063, N9142);
or OR4 (N14229, N14228, N12200, N13151, N14046);
nor NOR3 (N14230, N14225, N41, N526);
nand NAND4 (N14231, N14222, N3556, N4610, N3435);
or OR2 (N14232, N14223, N11368);
not NOT1 (N14233, N14219);
buf BUF1 (N14234, N14218);
or OR2 (N14235, N14230, N5468);
nand NAND3 (N14236, N14231, N9359, N8033);
not NOT1 (N14237, N14236);
buf BUF1 (N14238, N14227);
xor XOR2 (N14239, N14237, N12830);
or OR3 (N14240, N14234, N5755, N5563);
nand NAND2 (N14241, N14221, N11525);
xor XOR2 (N14242, N14239, N2368);
nand NAND2 (N14243, N14238, N7275);
buf BUF1 (N14244, N14240);
or OR4 (N14245, N14244, N11519, N10384, N7141);
xor XOR2 (N14246, N14229, N3815);
xor XOR2 (N14247, N14233, N2248);
not NOT1 (N14248, N14246);
and AND2 (N14249, N14224, N9114);
and AND3 (N14250, N14235, N13849, N9440);
not NOT1 (N14251, N14245);
not NOT1 (N14252, N14232);
xor XOR2 (N14253, N14250, N12421);
and AND2 (N14254, N14247, N14053);
or OR4 (N14255, N14254, N3490, N241, N11630);
buf BUF1 (N14256, N14242);
or OR2 (N14257, N14248, N5308);
nand NAND4 (N14258, N14252, N11545, N13030, N11455);
xor XOR2 (N14259, N14251, N12584);
not NOT1 (N14260, N14241);
and AND3 (N14261, N14260, N3590, N9746);
and AND4 (N14262, N14259, N10689, N290, N6370);
buf BUF1 (N14263, N14262);
not NOT1 (N14264, N14253);
xor XOR2 (N14265, N14258, N5247);
and AND4 (N14266, N14265, N8844, N12891, N11215);
xor XOR2 (N14267, N14257, N6665);
nand NAND2 (N14268, N14264, N9718);
and AND4 (N14269, N14255, N5785, N1756, N9889);
nor NOR2 (N14270, N14267, N6180);
xor XOR2 (N14271, N14261, N3990);
nor NOR2 (N14272, N14243, N12088);
xor XOR2 (N14273, N14263, N10884);
or OR2 (N14274, N14272, N13655);
buf BUF1 (N14275, N14191);
or OR4 (N14276, N14274, N6281, N6900, N103);
or OR2 (N14277, N14273, N14144);
and AND3 (N14278, N14249, N2524, N3048);
nor NOR3 (N14279, N14275, N10051, N9162);
and AND3 (N14280, N14279, N6771, N3708);
xor XOR2 (N14281, N14270, N8877);
and AND2 (N14282, N14280, N8015);
and AND3 (N14283, N14256, N8775, N1109);
xor XOR2 (N14284, N14276, N4129);
nor NOR2 (N14285, N14277, N7688);
nor NOR4 (N14286, N14278, N11053, N11412, N3059);
and AND2 (N14287, N14282, N7820);
nand NAND4 (N14288, N14271, N13310, N4565, N6203);
buf BUF1 (N14289, N14288);
nor NOR4 (N14290, N14286, N5674, N2890, N14148);
nor NOR3 (N14291, N14266, N12253, N9966);
nand NAND2 (N14292, N14285, N13170);
nand NAND3 (N14293, N14289, N2070, N32);
buf BUF1 (N14294, N14284);
nor NOR3 (N14295, N14269, N804, N12782);
nand NAND4 (N14296, N14290, N13271, N7239, N11582);
nor NOR4 (N14297, N14296, N6809, N8207, N13128);
or OR3 (N14298, N14295, N11502, N11365);
not NOT1 (N14299, N14294);
or OR4 (N14300, N14293, N14207, N3604, N4801);
xor XOR2 (N14301, N14283, N712);
or OR3 (N14302, N14297, N1795, N2891);
nand NAND4 (N14303, N14268, N5214, N703, N6650);
not NOT1 (N14304, N14301);
not NOT1 (N14305, N14298);
not NOT1 (N14306, N14287);
xor XOR2 (N14307, N14303, N10964);
nand NAND4 (N14308, N14299, N5772, N58, N147);
nor NOR4 (N14309, N14304, N5042, N1237, N3798);
or OR2 (N14310, N14305, N11241);
nand NAND3 (N14311, N14300, N4188, N12596);
or OR4 (N14312, N14311, N2817, N3792, N6012);
xor XOR2 (N14313, N14306, N8892);
nand NAND3 (N14314, N14312, N542, N3913);
and AND4 (N14315, N14307, N3832, N7397, N3000);
not NOT1 (N14316, N14281);
buf BUF1 (N14317, N14314);
nand NAND4 (N14318, N14308, N11825, N2971, N2591);
not NOT1 (N14319, N14291);
and AND4 (N14320, N14302, N3896, N10257, N11019);
nor NOR4 (N14321, N14318, N7088, N1859, N9317);
not NOT1 (N14322, N14321);
buf BUF1 (N14323, N14320);
nand NAND4 (N14324, N14317, N13607, N2255, N1266);
or OR4 (N14325, N14322, N1887, N13237, N12636);
nand NAND2 (N14326, N14315, N6019);
nand NAND2 (N14327, N14326, N2863);
buf BUF1 (N14328, N14309);
and AND2 (N14329, N14313, N6479);
buf BUF1 (N14330, N14327);
nand NAND4 (N14331, N14324, N5504, N8190, N1414);
not NOT1 (N14332, N14292);
or OR3 (N14333, N14332, N5615, N2875);
buf BUF1 (N14334, N14319);
nand NAND3 (N14335, N14334, N6632, N7290);
buf BUF1 (N14336, N14325);
nand NAND2 (N14337, N14310, N1997);
and AND4 (N14338, N14335, N3763, N5820, N11657);
and AND4 (N14339, N14333, N13444, N11894, N12101);
nor NOR3 (N14340, N14329, N1374, N2782);
and AND2 (N14341, N14338, N946);
nand NAND4 (N14342, N14336, N10928, N12685, N7872);
or OR3 (N14343, N14340, N2534, N8112);
nand NAND4 (N14344, N14331, N13775, N2117, N799);
xor XOR2 (N14345, N14342, N5649);
nor NOR4 (N14346, N14330, N7294, N1102, N13851);
not NOT1 (N14347, N14316);
nand NAND3 (N14348, N14344, N8329, N10677);
xor XOR2 (N14349, N14341, N6884);
nand NAND4 (N14350, N14347, N5105, N175, N4707);
and AND3 (N14351, N14337, N3831, N4496);
and AND3 (N14352, N14343, N3527, N11159);
nor NOR2 (N14353, N14349, N10776);
buf BUF1 (N14354, N14345);
or OR2 (N14355, N14323, N1163);
not NOT1 (N14356, N14348);
xor XOR2 (N14357, N14328, N8437);
buf BUF1 (N14358, N14346);
nand NAND3 (N14359, N14355, N752, N12827);
nor NOR4 (N14360, N14359, N7429, N10687, N4246);
nand NAND4 (N14361, N14358, N5207, N1333, N9633);
nor NOR2 (N14362, N14351, N14355);
nand NAND2 (N14363, N14361, N10220);
nor NOR4 (N14364, N14362, N2226, N9792, N5057);
not NOT1 (N14365, N14350);
nand NAND2 (N14366, N14352, N2222);
and AND3 (N14367, N14356, N8542, N5520);
and AND2 (N14368, N14367, N2310);
and AND2 (N14369, N14357, N4569);
nor NOR2 (N14370, N14369, N12655);
xor XOR2 (N14371, N14363, N6987);
nor NOR3 (N14372, N14366, N1286, N6083);
not NOT1 (N14373, N14364);
xor XOR2 (N14374, N14353, N5830);
xor XOR2 (N14375, N14365, N7564);
nand NAND4 (N14376, N14370, N5482, N7251, N2679);
or OR2 (N14377, N14368, N1320);
and AND2 (N14378, N14375, N2160);
nand NAND4 (N14379, N14374, N968, N2488, N9050);
xor XOR2 (N14380, N14377, N6396);
xor XOR2 (N14381, N14379, N11772);
nand NAND3 (N14382, N14380, N13849, N415);
not NOT1 (N14383, N14378);
nor NOR2 (N14384, N14373, N3948);
xor XOR2 (N14385, N14384, N11350);
not NOT1 (N14386, N14372);
and AND4 (N14387, N14376, N5780, N8843, N12615);
xor XOR2 (N14388, N14339, N7896);
xor XOR2 (N14389, N14387, N13742);
and AND2 (N14390, N14371, N3912);
nand NAND4 (N14391, N14389, N13998, N7128, N12514);
nand NAND4 (N14392, N14388, N10796, N7746, N14374);
not NOT1 (N14393, N14385);
and AND4 (N14394, N14381, N12050, N14126, N4322);
nor NOR3 (N14395, N14392, N11814, N7063);
or OR2 (N14396, N14390, N9361);
nand NAND3 (N14397, N14391, N457, N14031);
nand NAND2 (N14398, N14383, N13798);
or OR2 (N14399, N14382, N10008);
xor XOR2 (N14400, N14399, N7381);
nand NAND3 (N14401, N14396, N13368, N870);
not NOT1 (N14402, N14401);
buf BUF1 (N14403, N14395);
not NOT1 (N14404, N14393);
buf BUF1 (N14405, N14398);
not NOT1 (N14406, N14394);
or OR2 (N14407, N14397, N13410);
xor XOR2 (N14408, N14400, N12105);
nor NOR3 (N14409, N14408, N13543, N11830);
buf BUF1 (N14410, N14405);
xor XOR2 (N14411, N14404, N3419);
and AND2 (N14412, N14410, N11903);
and AND4 (N14413, N14406, N7629, N13559, N8016);
or OR2 (N14414, N14411, N781);
buf BUF1 (N14415, N14403);
or OR4 (N14416, N14360, N12212, N13013, N2054);
not NOT1 (N14417, N14354);
or OR4 (N14418, N14417, N9547, N10108, N13021);
xor XOR2 (N14419, N14402, N9889);
not NOT1 (N14420, N14407);
or OR4 (N14421, N14420, N7531, N7017, N3112);
not NOT1 (N14422, N14409);
nand NAND4 (N14423, N14386, N10991, N10696, N1338);
nor NOR3 (N14424, N14415, N5307, N14331);
nor NOR4 (N14425, N14422, N14073, N7783, N3776);
nand NAND3 (N14426, N14419, N5344, N13588);
buf BUF1 (N14427, N14423);
not NOT1 (N14428, N14425);
and AND3 (N14429, N14421, N1625, N10808);
not NOT1 (N14430, N14429);
or OR4 (N14431, N14418, N2462, N5094, N8262);
xor XOR2 (N14432, N14413, N1063);
buf BUF1 (N14433, N14424);
and AND4 (N14434, N14430, N11843, N4803, N2840);
buf BUF1 (N14435, N14414);
not NOT1 (N14436, N14428);
nor NOR2 (N14437, N14435, N859);
buf BUF1 (N14438, N14434);
not NOT1 (N14439, N14431);
and AND3 (N14440, N14432, N691, N10285);
not NOT1 (N14441, N14426);
nor NOR2 (N14442, N14427, N3836);
or OR2 (N14443, N14441, N3164);
nand NAND3 (N14444, N14436, N12386, N13213);
nand NAND2 (N14445, N14440, N12165);
and AND4 (N14446, N14445, N13378, N9027, N11125);
and AND4 (N14447, N14438, N11620, N9382, N4124);
buf BUF1 (N14448, N14439);
nand NAND2 (N14449, N14412, N5266);
buf BUF1 (N14450, N14447);
buf BUF1 (N14451, N14450);
nor NOR3 (N14452, N14433, N11544, N2816);
buf BUF1 (N14453, N14443);
buf BUF1 (N14454, N14452);
xor XOR2 (N14455, N14451, N2532);
or OR3 (N14456, N14437, N9797, N4013);
nor NOR2 (N14457, N14448, N10314);
not NOT1 (N14458, N14442);
buf BUF1 (N14459, N14449);
not NOT1 (N14460, N14453);
nor NOR3 (N14461, N14455, N10564, N5097);
nand NAND4 (N14462, N14454, N7422, N2163, N12175);
nor NOR3 (N14463, N14444, N4895, N12959);
nor NOR2 (N14464, N14457, N9052);
and AND3 (N14465, N14464, N257, N13571);
buf BUF1 (N14466, N14459);
nand NAND3 (N14467, N14466, N2105, N7682);
buf BUF1 (N14468, N14446);
not NOT1 (N14469, N14458);
buf BUF1 (N14470, N14465);
or OR4 (N14471, N14467, N13767, N6891, N4059);
or OR4 (N14472, N14456, N7852, N3048, N3028);
or OR4 (N14473, N14471, N10896, N11610, N1849);
and AND2 (N14474, N14463, N5663);
and AND2 (N14475, N14470, N4789);
xor XOR2 (N14476, N14460, N6182);
buf BUF1 (N14477, N14416);
not NOT1 (N14478, N14462);
nor NOR3 (N14479, N14468, N4588, N573);
or OR3 (N14480, N14476, N12199, N12838);
or OR2 (N14481, N14479, N9529);
or OR2 (N14482, N14461, N2468);
not NOT1 (N14483, N14478);
buf BUF1 (N14484, N14472);
nor NOR4 (N14485, N14475, N4984, N9982, N7066);
nor NOR2 (N14486, N14469, N11826);
nor NOR4 (N14487, N14483, N10370, N2267, N10313);
buf BUF1 (N14488, N14481);
or OR4 (N14489, N14487, N1499, N7593, N1997);
nor NOR3 (N14490, N14474, N4395, N6376);
and AND3 (N14491, N14488, N1444, N8421);
nor NOR2 (N14492, N14485, N3320);
not NOT1 (N14493, N14477);
xor XOR2 (N14494, N14482, N4590);
buf BUF1 (N14495, N14491);
not NOT1 (N14496, N14484);
buf BUF1 (N14497, N14489);
buf BUF1 (N14498, N14480);
nor NOR2 (N14499, N14493, N13243);
xor XOR2 (N14500, N14498, N13060);
or OR3 (N14501, N14473, N328, N1424);
not NOT1 (N14502, N14492);
not NOT1 (N14503, N14502);
buf BUF1 (N14504, N14503);
xor XOR2 (N14505, N14497, N3698);
nor NOR4 (N14506, N14495, N3514, N11713, N820);
or OR2 (N14507, N14501, N11631);
buf BUF1 (N14508, N14486);
or OR3 (N14509, N14496, N2250, N6441);
and AND2 (N14510, N14506, N13961);
or OR4 (N14511, N14499, N3421, N9105, N12274);
or OR4 (N14512, N14507, N9659, N8057, N11621);
nor NOR3 (N14513, N14494, N179, N3362);
buf BUF1 (N14514, N14512);
nand NAND4 (N14515, N14508, N11855, N12633, N10131);
nand NAND2 (N14516, N14500, N3059);
xor XOR2 (N14517, N14490, N11538);
buf BUF1 (N14518, N14515);
and AND4 (N14519, N14504, N9539, N5303, N9056);
nand NAND4 (N14520, N14509, N12656, N5772, N7747);
buf BUF1 (N14521, N14511);
xor XOR2 (N14522, N14514, N10876);
buf BUF1 (N14523, N14518);
buf BUF1 (N14524, N14521);
xor XOR2 (N14525, N14510, N13768);
or OR2 (N14526, N14505, N3123);
nor NOR3 (N14527, N14520, N1583, N12677);
xor XOR2 (N14528, N14517, N9836);
and AND3 (N14529, N14525, N8587, N10726);
and AND4 (N14530, N14524, N12529, N1333, N3549);
nor NOR4 (N14531, N14523, N10568, N6778, N3435);
not NOT1 (N14532, N14526);
nor NOR2 (N14533, N14529, N1590);
or OR4 (N14534, N14531, N5859, N11320, N10079);
xor XOR2 (N14535, N14533, N1845);
or OR3 (N14536, N14522, N2994, N9701);
nor NOR3 (N14537, N14530, N4344, N3692);
or OR3 (N14538, N14537, N5254, N10256);
or OR2 (N14539, N14535, N3959);
buf BUF1 (N14540, N14536);
buf BUF1 (N14541, N14516);
xor XOR2 (N14542, N14539, N7905);
or OR4 (N14543, N14540, N11149, N12644, N6881);
nor NOR2 (N14544, N14541, N71);
xor XOR2 (N14545, N14513, N4253);
not NOT1 (N14546, N14545);
buf BUF1 (N14547, N14528);
buf BUF1 (N14548, N14527);
nand NAND3 (N14549, N14543, N16, N10319);
buf BUF1 (N14550, N14519);
xor XOR2 (N14551, N14548, N12531);
and AND2 (N14552, N14534, N13192);
nand NAND3 (N14553, N14550, N5135, N9385);
nor NOR2 (N14554, N14551, N1219);
nand NAND4 (N14555, N14532, N9181, N9482, N6306);
and AND3 (N14556, N14542, N6875, N2755);
not NOT1 (N14557, N14552);
or OR4 (N14558, N14557, N3294, N12546, N5822);
not NOT1 (N14559, N14547);
or OR2 (N14560, N14556, N10709);
buf BUF1 (N14561, N14544);
and AND2 (N14562, N14560, N6974);
xor XOR2 (N14563, N14561, N4329);
or OR4 (N14564, N14559, N5576, N14336, N10267);
and AND4 (N14565, N14546, N14438, N7428, N181);
not NOT1 (N14566, N14563);
or OR4 (N14567, N14564, N13872, N4904, N3648);
or OR2 (N14568, N14566, N6512);
nor NOR2 (N14569, N14565, N3596);
or OR3 (N14570, N14558, N12047, N3700);
nand NAND3 (N14571, N14568, N6050, N11100);
nor NOR3 (N14572, N14555, N7382, N10589);
xor XOR2 (N14573, N14567, N11982);
and AND2 (N14574, N14553, N6969);
nand NAND3 (N14575, N14573, N8405, N3614);
nand NAND2 (N14576, N14571, N790);
nand NAND4 (N14577, N14574, N6018, N5219, N13035);
nand NAND4 (N14578, N14554, N7392, N11180, N3431);
buf BUF1 (N14579, N14562);
xor XOR2 (N14580, N14576, N7178);
nor NOR3 (N14581, N14575, N10531, N13542);
buf BUF1 (N14582, N14549);
and AND4 (N14583, N14582, N6785, N5564, N3759);
and AND3 (N14584, N14577, N12616, N4548);
nor NOR4 (N14585, N14570, N3273, N11570, N1398);
or OR3 (N14586, N14583, N14530, N4823);
nand NAND3 (N14587, N14584, N2975, N9835);
nor NOR3 (N14588, N14587, N7717, N1167);
not NOT1 (N14589, N14585);
and AND3 (N14590, N14588, N10517, N1997);
or OR3 (N14591, N14578, N7912, N3211);
nand NAND4 (N14592, N14589, N9627, N2339, N2602);
or OR4 (N14593, N14580, N4313, N13545, N5696);
nand NAND3 (N14594, N14581, N11779, N3220);
nor NOR4 (N14595, N14594, N13089, N13849, N256);
or OR3 (N14596, N14572, N7123, N2309);
nand NAND4 (N14597, N14593, N10760, N12886, N1968);
buf BUF1 (N14598, N14591);
not NOT1 (N14599, N14586);
buf BUF1 (N14600, N14538);
nand NAND4 (N14601, N14600, N14098, N11171, N10210);
and AND3 (N14602, N14590, N11976, N12083);
xor XOR2 (N14603, N14592, N11850);
xor XOR2 (N14604, N14601, N2764);
buf BUF1 (N14605, N14598);
or OR4 (N14606, N14602, N11473, N10706, N14284);
nor NOR2 (N14607, N14606, N13730);
nor NOR2 (N14608, N14569, N94);
and AND4 (N14609, N14595, N14477, N508, N5846);
and AND3 (N14610, N14607, N9460, N5178);
xor XOR2 (N14611, N14579, N3020);
not NOT1 (N14612, N14611);
nor NOR4 (N14613, N14604, N13742, N13109, N1265);
buf BUF1 (N14614, N14609);
buf BUF1 (N14615, N14612);
xor XOR2 (N14616, N14605, N9457);
not NOT1 (N14617, N14614);
nand NAND2 (N14618, N14613, N324);
nor NOR3 (N14619, N14610, N9958, N2371);
buf BUF1 (N14620, N14616);
nand NAND3 (N14621, N14615, N1073, N2361);
not NOT1 (N14622, N14620);
and AND3 (N14623, N14621, N8557, N5567);
or OR2 (N14624, N14623, N2812);
and AND4 (N14625, N14596, N12437, N8598, N11206);
or OR4 (N14626, N14603, N5710, N4981, N1292);
nor NOR4 (N14627, N14626, N13567, N10342, N11780);
xor XOR2 (N14628, N14622, N556);
not NOT1 (N14629, N14599);
or OR3 (N14630, N14619, N7502, N523);
nand NAND3 (N14631, N14618, N1366, N9130);
not NOT1 (N14632, N14631);
nand NAND4 (N14633, N14608, N10904, N9893, N2973);
not NOT1 (N14634, N14597);
xor XOR2 (N14635, N14633, N4994);
buf BUF1 (N14636, N14628);
nand NAND4 (N14637, N14634, N2344, N3409, N5648);
xor XOR2 (N14638, N14637, N4668);
nor NOR2 (N14639, N14627, N3142);
buf BUF1 (N14640, N14635);
buf BUF1 (N14641, N14638);
or OR3 (N14642, N14629, N14125, N7143);
and AND3 (N14643, N14640, N7323, N7264);
xor XOR2 (N14644, N14617, N14010);
nand NAND2 (N14645, N14630, N13489);
buf BUF1 (N14646, N14636);
not NOT1 (N14647, N14624);
nor NOR3 (N14648, N14644, N4552, N4628);
nand NAND3 (N14649, N14642, N10392, N7211);
nor NOR2 (N14650, N14643, N9774);
and AND3 (N14651, N14641, N11151, N8667);
nor NOR3 (N14652, N14646, N3195, N2256);
buf BUF1 (N14653, N14648);
and AND2 (N14654, N14650, N11530);
not NOT1 (N14655, N14645);
nor NOR3 (N14656, N14652, N6647, N9659);
xor XOR2 (N14657, N14651, N8817);
buf BUF1 (N14658, N14655);
nand NAND3 (N14659, N14654, N5425, N1637);
buf BUF1 (N14660, N14625);
nand NAND4 (N14661, N14660, N5995, N732, N13409);
xor XOR2 (N14662, N14659, N13625);
nand NAND2 (N14663, N14647, N7791);
xor XOR2 (N14664, N14656, N14194);
or OR3 (N14665, N14661, N12295, N9691);
not NOT1 (N14666, N14632);
buf BUF1 (N14667, N14649);
nand NAND4 (N14668, N14666, N4098, N12967, N2261);
nor NOR3 (N14669, N14664, N2159, N6505);
xor XOR2 (N14670, N14663, N601);
or OR4 (N14671, N14639, N6491, N1995, N341);
buf BUF1 (N14672, N14665);
nand NAND2 (N14673, N14671, N10905);
not NOT1 (N14674, N14658);
and AND3 (N14675, N14669, N5050, N13120);
or OR4 (N14676, N14672, N1459, N14548, N9259);
not NOT1 (N14677, N14667);
not NOT1 (N14678, N14662);
or OR4 (N14679, N14653, N270, N13234, N12138);
not NOT1 (N14680, N14678);
nor NOR4 (N14681, N14680, N3822, N741, N11143);
xor XOR2 (N14682, N14676, N10512);
not NOT1 (N14683, N14673);
not NOT1 (N14684, N14657);
buf BUF1 (N14685, N14675);
xor XOR2 (N14686, N14674, N6313);
nand NAND3 (N14687, N14684, N6924, N9780);
nand NAND4 (N14688, N14687, N11675, N5042, N13134);
xor XOR2 (N14689, N14668, N13940);
nor NOR2 (N14690, N14681, N9464);
nor NOR3 (N14691, N14682, N8131, N6861);
and AND2 (N14692, N14691, N8676);
and AND4 (N14693, N14688, N7364, N2784, N10356);
nand NAND2 (N14694, N14683, N5012);
nand NAND4 (N14695, N14677, N6161, N3495, N13509);
buf BUF1 (N14696, N14685);
buf BUF1 (N14697, N14689);
and AND4 (N14698, N14693, N1793, N5195, N988);
nor NOR3 (N14699, N14692, N371, N9581);
nand NAND4 (N14700, N14686, N4664, N10505, N7109);
and AND3 (N14701, N14697, N5470, N11506);
or OR3 (N14702, N14690, N10427, N14008);
and AND3 (N14703, N14698, N2708, N7966);
nand NAND2 (N14704, N14700, N3027);
nor NOR2 (N14705, N14696, N48);
and AND4 (N14706, N14670, N13693, N5478, N10516);
xor XOR2 (N14707, N14694, N13456);
nand NAND4 (N14708, N14707, N4039, N14673, N272);
not NOT1 (N14709, N14706);
xor XOR2 (N14710, N14709, N6057);
xor XOR2 (N14711, N14699, N5917);
xor XOR2 (N14712, N14708, N9924);
or OR4 (N14713, N14679, N2991, N7742, N3105);
buf BUF1 (N14714, N14710);
not NOT1 (N14715, N14712);
nor NOR2 (N14716, N14703, N8639);
and AND2 (N14717, N14714, N10880);
nand NAND4 (N14718, N14702, N14215, N14574, N7365);
xor XOR2 (N14719, N14711, N2388);
xor XOR2 (N14720, N14713, N13781);
nor NOR4 (N14721, N14701, N11038, N7019, N7833);
xor XOR2 (N14722, N14705, N5035);
buf BUF1 (N14723, N14716);
xor XOR2 (N14724, N14723, N13762);
xor XOR2 (N14725, N14724, N12255);
xor XOR2 (N14726, N14717, N9648);
and AND4 (N14727, N14722, N366, N1090, N9676);
not NOT1 (N14728, N14726);
or OR3 (N14729, N14718, N1891, N9044);
xor XOR2 (N14730, N14719, N4259);
or OR3 (N14731, N14730, N10685, N3504);
nor NOR3 (N14732, N14727, N13597, N6834);
nor NOR4 (N14733, N14721, N14140, N13760, N8504);
or OR4 (N14734, N14733, N13937, N6220, N11968);
xor XOR2 (N14735, N14704, N4920);
or OR2 (N14736, N14734, N5708);
and AND3 (N14737, N14720, N5237, N5495);
or OR2 (N14738, N14737, N14553);
or OR4 (N14739, N14735, N13857, N9291, N1342);
or OR2 (N14740, N14739, N5682);
and AND4 (N14741, N14731, N12392, N11843, N1084);
and AND4 (N14742, N14695, N3375, N9790, N6514);
not NOT1 (N14743, N14741);
not NOT1 (N14744, N14729);
buf BUF1 (N14745, N14732);
or OR4 (N14746, N14715, N8835, N13287, N4576);
buf BUF1 (N14747, N14740);
nand NAND4 (N14748, N14725, N8044, N10250, N726);
buf BUF1 (N14749, N14748);
or OR2 (N14750, N14745, N12143);
xor XOR2 (N14751, N14750, N8372);
nand NAND2 (N14752, N14728, N4572);
nor NOR3 (N14753, N14736, N2756, N325);
nor NOR2 (N14754, N14738, N3193);
buf BUF1 (N14755, N14754);
not NOT1 (N14756, N14746);
nor NOR4 (N14757, N14743, N7959, N5747, N6648);
not NOT1 (N14758, N14752);
nand NAND3 (N14759, N14758, N6687, N11142);
nand NAND4 (N14760, N14755, N11237, N13173, N3138);
nand NAND2 (N14761, N14744, N324);
and AND3 (N14762, N14742, N7526, N9943);
and AND2 (N14763, N14747, N4476);
nand NAND4 (N14764, N14753, N8940, N9117, N5054);
xor XOR2 (N14765, N14764, N7635);
xor XOR2 (N14766, N14756, N8982);
nand NAND4 (N14767, N14749, N10554, N742, N4474);
buf BUF1 (N14768, N14766);
nand NAND3 (N14769, N14760, N917, N1968);
and AND4 (N14770, N14761, N9756, N6438, N11595);
nand NAND3 (N14771, N14759, N14165, N2311);
nor NOR2 (N14772, N14770, N6785);
not NOT1 (N14773, N14767);
and AND2 (N14774, N14772, N9141);
not NOT1 (N14775, N14751);
nand NAND2 (N14776, N14775, N2655);
nand NAND2 (N14777, N14774, N178);
not NOT1 (N14778, N14763);
buf BUF1 (N14779, N14778);
not NOT1 (N14780, N14762);
nand NAND2 (N14781, N14771, N4139);
and AND2 (N14782, N14757, N4539);
and AND2 (N14783, N14777, N2913);
nand NAND4 (N14784, N14779, N1977, N5756, N6210);
nand NAND2 (N14785, N14782, N11932);
nand NAND4 (N14786, N14781, N9179, N13551, N3186);
xor XOR2 (N14787, N14780, N6368);
buf BUF1 (N14788, N14768);
or OR4 (N14789, N14788, N2820, N12658, N644);
or OR4 (N14790, N14783, N7001, N13894, N1138);
xor XOR2 (N14791, N14773, N11220);
nand NAND2 (N14792, N14765, N10374);
not NOT1 (N14793, N14785);
buf BUF1 (N14794, N14776);
buf BUF1 (N14795, N14789);
xor XOR2 (N14796, N14792, N14342);
nand NAND4 (N14797, N14790, N2417, N6631, N6063);
and AND2 (N14798, N14769, N5088);
or OR3 (N14799, N14786, N748, N13942);
nand NAND2 (N14800, N14796, N3808);
and AND2 (N14801, N14787, N5354);
nor NOR4 (N14802, N14800, N4630, N1169, N9166);
or OR3 (N14803, N14793, N10869, N6747);
and AND4 (N14804, N14802, N3933, N3114, N10623);
nor NOR4 (N14805, N14795, N4087, N13615, N3211);
nand NAND4 (N14806, N14803, N10342, N1932, N7506);
nand NAND4 (N14807, N14804, N5851, N4512, N7650);
or OR4 (N14808, N14799, N13659, N13626, N8215);
or OR3 (N14809, N14807, N12605, N12515);
nor NOR4 (N14810, N14798, N8716, N4242, N13441);
and AND2 (N14811, N14809, N13944);
buf BUF1 (N14812, N14784);
not NOT1 (N14813, N14810);
nand NAND4 (N14814, N14797, N1960, N5150, N11823);
and AND3 (N14815, N14806, N13146, N2114);
nand NAND3 (N14816, N14815, N11902, N12274);
buf BUF1 (N14817, N14808);
or OR3 (N14818, N14817, N4950, N13535);
xor XOR2 (N14819, N14794, N4410);
xor XOR2 (N14820, N14801, N8948);
or OR3 (N14821, N14816, N14674, N8370);
nor NOR2 (N14822, N14818, N1922);
xor XOR2 (N14823, N14811, N13867);
nor NOR4 (N14824, N14791, N4778, N12663, N14780);
or OR2 (N14825, N14823, N13833);
or OR2 (N14826, N14822, N11956);
buf BUF1 (N14827, N14813);
and AND2 (N14828, N14805, N1908);
nand NAND2 (N14829, N14820, N20);
xor XOR2 (N14830, N14824, N9123);
nand NAND2 (N14831, N14825, N5712);
not NOT1 (N14832, N14819);
nor NOR3 (N14833, N14821, N8244, N6644);
nor NOR4 (N14834, N14827, N7899, N4601, N1431);
buf BUF1 (N14835, N14826);
nor NOR4 (N14836, N14833, N8774, N10088, N12054);
nand NAND4 (N14837, N14834, N12341, N14677, N10331);
nor NOR3 (N14838, N14829, N12366, N10465);
nand NAND3 (N14839, N14838, N1091, N13851);
and AND4 (N14840, N14836, N5106, N11696, N10233);
or OR2 (N14841, N14828, N11767);
or OR4 (N14842, N14831, N13511, N14454, N14424);
nand NAND3 (N14843, N14830, N11019, N9702);
not NOT1 (N14844, N14812);
and AND4 (N14845, N14839, N8902, N11020, N2308);
not NOT1 (N14846, N14843);
and AND3 (N14847, N14842, N271, N9931);
nand NAND4 (N14848, N14840, N6611, N13882, N13582);
not NOT1 (N14849, N14845);
buf BUF1 (N14850, N14847);
not NOT1 (N14851, N14844);
buf BUF1 (N14852, N14851);
xor XOR2 (N14853, N14848, N1242);
or OR2 (N14854, N14853, N11176);
nor NOR2 (N14855, N14814, N928);
nor NOR2 (N14856, N14849, N11667);
nand NAND3 (N14857, N14835, N9883, N6584);
nand NAND4 (N14858, N14852, N12764, N7772, N755);
buf BUF1 (N14859, N14832);
buf BUF1 (N14860, N14855);
buf BUF1 (N14861, N14837);
and AND2 (N14862, N14860, N9646);
buf BUF1 (N14863, N14850);
and AND3 (N14864, N14854, N6327, N14090);
and AND2 (N14865, N14862, N4931);
nor NOR3 (N14866, N14858, N2389, N10656);
not NOT1 (N14867, N14856);
nand NAND3 (N14868, N14866, N4981, N10526);
and AND2 (N14869, N14846, N11709);
and AND3 (N14870, N14861, N9738, N11765);
or OR2 (N14871, N14870, N3748);
not NOT1 (N14872, N14864);
and AND3 (N14873, N14872, N7823, N9889);
nor NOR2 (N14874, N14859, N363);
nor NOR4 (N14875, N14874, N12892, N3141, N1222);
xor XOR2 (N14876, N14865, N12218);
and AND2 (N14877, N14868, N14532);
nand NAND4 (N14878, N14877, N14612, N8209, N5151);
nor NOR3 (N14879, N14863, N4724, N9936);
not NOT1 (N14880, N14873);
nor NOR3 (N14881, N14841, N8892, N11962);
not NOT1 (N14882, N14875);
not NOT1 (N14883, N14878);
nand NAND4 (N14884, N14882, N6372, N11237, N7771);
not NOT1 (N14885, N14884);
buf BUF1 (N14886, N14883);
not NOT1 (N14887, N14876);
buf BUF1 (N14888, N14885);
nor NOR3 (N14889, N14886, N614, N6648);
or OR2 (N14890, N14888, N8233);
buf BUF1 (N14891, N14890);
not NOT1 (N14892, N14869);
nand NAND3 (N14893, N14880, N7405, N2176);
or OR3 (N14894, N14892, N934, N1601);
nor NOR2 (N14895, N14879, N4759);
or OR3 (N14896, N14893, N6332, N9929);
xor XOR2 (N14897, N14895, N11927);
buf BUF1 (N14898, N14891);
not NOT1 (N14899, N14867);
nor NOR3 (N14900, N14894, N1100, N7017);
buf BUF1 (N14901, N14871);
and AND2 (N14902, N14889, N10709);
buf BUF1 (N14903, N14857);
nand NAND3 (N14904, N14881, N775, N11928);
not NOT1 (N14905, N14898);
and AND4 (N14906, N14887, N9554, N6507, N10207);
or OR3 (N14907, N14904, N11918, N3089);
buf BUF1 (N14908, N14902);
not NOT1 (N14909, N14899);
and AND2 (N14910, N14909, N10218);
buf BUF1 (N14911, N14896);
nor NOR2 (N14912, N14906, N1914);
xor XOR2 (N14913, N14912, N7015);
and AND2 (N14914, N14901, N11341);
not NOT1 (N14915, N14900);
not NOT1 (N14916, N14910);
nor NOR2 (N14917, N14897, N11668);
and AND4 (N14918, N14908, N8770, N3966, N6953);
nand NAND2 (N14919, N14915, N8247);
nand NAND3 (N14920, N14905, N11356, N5666);
xor XOR2 (N14921, N14917, N12616);
nand NAND2 (N14922, N14903, N3665);
not NOT1 (N14923, N14907);
buf BUF1 (N14924, N14920);
or OR4 (N14925, N14913, N3831, N9264, N6974);
xor XOR2 (N14926, N14916, N12731);
nor NOR3 (N14927, N14921, N5261, N13331);
buf BUF1 (N14928, N14911);
nand NAND4 (N14929, N14922, N5919, N13446, N13113);
not NOT1 (N14930, N14928);
and AND2 (N14931, N14924, N6466);
or OR2 (N14932, N14914, N174);
or OR3 (N14933, N14930, N4161, N10129);
and AND3 (N14934, N14925, N12352, N13068);
nand NAND3 (N14935, N14923, N4531, N8017);
and AND3 (N14936, N14931, N4762, N1210);
and AND3 (N14937, N14919, N2398, N969);
buf BUF1 (N14938, N14933);
not NOT1 (N14939, N14935);
buf BUF1 (N14940, N14926);
or OR4 (N14941, N14940, N14225, N10341, N8142);
nor NOR3 (N14942, N14939, N1627, N13035);
and AND2 (N14943, N14934, N3186);
buf BUF1 (N14944, N14927);
buf BUF1 (N14945, N14941);
not NOT1 (N14946, N14944);
nand NAND2 (N14947, N14943, N7857);
nand NAND4 (N14948, N14942, N5181, N11981, N5761);
nand NAND2 (N14949, N14937, N8216);
not NOT1 (N14950, N14948);
xor XOR2 (N14951, N14936, N10711);
nor NOR3 (N14952, N14951, N2493, N850);
buf BUF1 (N14953, N14947);
buf BUF1 (N14954, N14946);
nand NAND2 (N14955, N14938, N4893);
nor NOR2 (N14956, N14945, N10530);
nor NOR4 (N14957, N14918, N7833, N2622, N644);
not NOT1 (N14958, N14949);
and AND2 (N14959, N14955, N4086);
and AND2 (N14960, N14957, N4675);
or OR2 (N14961, N14958, N331);
nand NAND3 (N14962, N14953, N12712, N2322);
nor NOR4 (N14963, N14959, N5914, N13734, N4050);
or OR4 (N14964, N14956, N7421, N13131, N4670);
and AND4 (N14965, N14963, N9798, N9198, N9422);
nand NAND2 (N14966, N14950, N11359);
xor XOR2 (N14967, N14961, N3997);
or OR2 (N14968, N14954, N11085);
xor XOR2 (N14969, N14929, N11020);
nand NAND2 (N14970, N14969, N4955);
or OR2 (N14971, N14968, N6183);
xor XOR2 (N14972, N14960, N13095);
nand NAND2 (N14973, N14967, N12452);
buf BUF1 (N14974, N14972);
xor XOR2 (N14975, N14971, N9231);
or OR3 (N14976, N14973, N3456, N13283);
nor NOR3 (N14977, N14932, N202, N2948);
and AND4 (N14978, N14952, N4340, N3240, N14206);
not NOT1 (N14979, N14978);
nand NAND3 (N14980, N14964, N940, N908);
xor XOR2 (N14981, N14974, N3901);
buf BUF1 (N14982, N14970);
xor XOR2 (N14983, N14982, N11992);
or OR3 (N14984, N14975, N14727, N3918);
nand NAND3 (N14985, N14984, N4276, N13384);
and AND2 (N14986, N14966, N11325);
and AND3 (N14987, N14985, N4727, N14275);
xor XOR2 (N14988, N14976, N2261);
and AND2 (N14989, N14980, N947);
xor XOR2 (N14990, N14962, N14503);
nor NOR3 (N14991, N14977, N14063, N7944);
not NOT1 (N14992, N14983);
nor NOR3 (N14993, N14965, N1463, N11999);
buf BUF1 (N14994, N14979);
buf BUF1 (N14995, N14988);
buf BUF1 (N14996, N14992);
or OR4 (N14997, N14990, N8836, N4276, N3117);
not NOT1 (N14998, N14997);
and AND4 (N14999, N14989, N10156, N2918, N6858);
not NOT1 (N15000, N14995);
xor XOR2 (N15001, N14994, N541);
not NOT1 (N15002, N14987);
buf BUF1 (N15003, N14996);
not NOT1 (N15004, N14993);
or OR2 (N15005, N15002, N11984);
not NOT1 (N15006, N14981);
buf BUF1 (N15007, N15000);
nand NAND3 (N15008, N15005, N11052, N7033);
or OR4 (N15009, N15004, N4118, N14867, N1158);
xor XOR2 (N15010, N14991, N8911);
xor XOR2 (N15011, N15008, N2763);
nor NOR3 (N15012, N15011, N12898, N8784);
nor NOR3 (N15013, N15007, N10729, N8144);
not NOT1 (N15014, N15003);
xor XOR2 (N15015, N15013, N13646);
nand NAND3 (N15016, N14986, N13867, N5447);
nor NOR4 (N15017, N15016, N6115, N10170, N10052);
not NOT1 (N15018, N15014);
or OR2 (N15019, N15015, N3118);
and AND2 (N15020, N15018, N8769);
not NOT1 (N15021, N15019);
and AND3 (N15022, N15009, N6815, N11040);
buf BUF1 (N15023, N15012);
nor NOR3 (N15024, N15010, N1766, N14440);
nand NAND4 (N15025, N15022, N10728, N3966, N8996);
and AND4 (N15026, N15001, N8967, N9066, N12770);
buf BUF1 (N15027, N15023);
buf BUF1 (N15028, N15006);
nand NAND3 (N15029, N15026, N13078, N3064);
nand NAND2 (N15030, N15025, N11600);
not NOT1 (N15031, N15020);
or OR3 (N15032, N15027, N720, N7141);
not NOT1 (N15033, N15021);
or OR2 (N15034, N15024, N12143);
xor XOR2 (N15035, N15034, N3874);
or OR2 (N15036, N15029, N14846);
or OR3 (N15037, N14999, N13637, N11365);
and AND2 (N15038, N15033, N13480);
nor NOR3 (N15039, N15038, N11374, N6462);
nand NAND2 (N15040, N15036, N857);
and AND3 (N15041, N15030, N14159, N1010);
and AND3 (N15042, N15031, N14200, N9739);
buf BUF1 (N15043, N15039);
nand NAND4 (N15044, N14998, N7740, N9503, N3249);
xor XOR2 (N15045, N15043, N11365);
buf BUF1 (N15046, N15028);
and AND3 (N15047, N15017, N239, N9620);
or OR2 (N15048, N15035, N12030);
or OR3 (N15049, N15047, N4587, N1819);
not NOT1 (N15050, N15037);
buf BUF1 (N15051, N15044);
nor NOR3 (N15052, N15041, N14712, N13429);
or OR2 (N15053, N15045, N5022);
nor NOR3 (N15054, N15046, N4188, N14634);
and AND4 (N15055, N15053, N10158, N861, N651);
nand NAND2 (N15056, N15050, N11960);
and AND2 (N15057, N15056, N4861);
nor NOR2 (N15058, N15048, N6630);
and AND2 (N15059, N15040, N6806);
or OR4 (N15060, N15058, N9610, N5096, N10962);
nor NOR2 (N15061, N15032, N9898);
not NOT1 (N15062, N15060);
or OR4 (N15063, N15057, N8449, N8719, N3169);
and AND2 (N15064, N15042, N13742);
nor NOR3 (N15065, N15054, N11419, N2825);
and AND2 (N15066, N15055, N14410);
nor NOR3 (N15067, N15061, N11989, N11153);
buf BUF1 (N15068, N15049);
nand NAND2 (N15069, N15059, N685);
xor XOR2 (N15070, N15066, N12766);
nand NAND4 (N15071, N15062, N4462, N5893, N14242);
or OR3 (N15072, N15071, N13949, N10193);
xor XOR2 (N15073, N15067, N5624);
nor NOR3 (N15074, N15069, N13686, N5009);
nor NOR2 (N15075, N15064, N4725);
buf BUF1 (N15076, N15065);
xor XOR2 (N15077, N15073, N4009);
xor XOR2 (N15078, N15070, N5747);
xor XOR2 (N15079, N15072, N13404);
nand NAND2 (N15080, N15052, N8148);
nand NAND3 (N15081, N15075, N14691, N11298);
and AND4 (N15082, N15074, N5930, N14179, N14204);
buf BUF1 (N15083, N15077);
nand NAND4 (N15084, N15083, N4529, N10895, N2050);
or OR4 (N15085, N15063, N6471, N4713, N6874);
or OR4 (N15086, N15079, N2051, N1338, N12415);
xor XOR2 (N15087, N15078, N13111);
or OR4 (N15088, N15087, N1192, N10539, N5716);
nor NOR2 (N15089, N15076, N7191);
not NOT1 (N15090, N15080);
not NOT1 (N15091, N15089);
xor XOR2 (N15092, N15081, N6625);
xor XOR2 (N15093, N15068, N2886);
nor NOR3 (N15094, N15092, N10535, N11200);
nand NAND2 (N15095, N15094, N11354);
or OR4 (N15096, N15082, N457, N2381, N14797);
nor NOR4 (N15097, N15084, N4786, N11552, N8370);
or OR4 (N15098, N15096, N13587, N9342, N11180);
nor NOR4 (N15099, N15093, N6713, N10053, N8864);
nand NAND3 (N15100, N15098, N7440, N5171);
buf BUF1 (N15101, N15085);
nor NOR2 (N15102, N15097, N11491);
and AND2 (N15103, N15088, N5520);
nor NOR3 (N15104, N15090, N6183, N10259);
buf BUF1 (N15105, N15101);
and AND3 (N15106, N15103, N3841, N14574);
and AND2 (N15107, N15100, N6052);
buf BUF1 (N15108, N15106);
or OR2 (N15109, N15051, N7903);
or OR2 (N15110, N15091, N9945);
xor XOR2 (N15111, N15107, N8253);
nor NOR4 (N15112, N15102, N6243, N1493, N14656);
xor XOR2 (N15113, N15095, N5621);
or OR4 (N15114, N15099, N11277, N6722, N4712);
and AND3 (N15115, N15109, N7866, N716);
buf BUF1 (N15116, N15113);
and AND2 (N15117, N15110, N6212);
xor XOR2 (N15118, N15116, N759);
xor XOR2 (N15119, N15115, N11308);
buf BUF1 (N15120, N15118);
or OR2 (N15121, N15111, N9232);
buf BUF1 (N15122, N15117);
xor XOR2 (N15123, N15112, N6918);
and AND2 (N15124, N15105, N13498);
nor NOR4 (N15125, N15124, N13388, N10474, N11670);
nand NAND2 (N15126, N15125, N5279);
nor NOR2 (N15127, N15123, N2449);
nor NOR4 (N15128, N15122, N12938, N4242, N7397);
nor NOR2 (N15129, N15120, N7509);
or OR3 (N15130, N15128, N9667, N9542);
buf BUF1 (N15131, N15130);
nor NOR3 (N15132, N15129, N2428, N2313);
nor NOR2 (N15133, N15114, N4625);
nand NAND2 (N15134, N15121, N10481);
nor NOR2 (N15135, N15104, N1713);
nor NOR4 (N15136, N15133, N13194, N12153, N7364);
not NOT1 (N15137, N15108);
and AND4 (N15138, N15126, N14511, N7329, N12556);
or OR2 (N15139, N15134, N3359);
not NOT1 (N15140, N15135);
or OR4 (N15141, N15132, N2848, N11366, N5361);
not NOT1 (N15142, N15119);
buf BUF1 (N15143, N15086);
and AND2 (N15144, N15137, N9974);
nor NOR3 (N15145, N15136, N8508, N13481);
or OR3 (N15146, N15140, N3464, N5523);
nor NOR2 (N15147, N15139, N13683);
nand NAND3 (N15148, N15145, N4129, N5402);
not NOT1 (N15149, N15143);
not NOT1 (N15150, N15138);
and AND2 (N15151, N15131, N9938);
nand NAND2 (N15152, N15150, N458);
or OR2 (N15153, N15141, N12654);
not NOT1 (N15154, N15142);
buf BUF1 (N15155, N15147);
xor XOR2 (N15156, N15127, N8679);
and AND2 (N15157, N15156, N3991);
not NOT1 (N15158, N15154);
not NOT1 (N15159, N15155);
or OR3 (N15160, N15159, N9754, N9516);
not NOT1 (N15161, N15144);
not NOT1 (N15162, N15149);
or OR2 (N15163, N15160, N5544);
nor NOR3 (N15164, N15153, N10399, N1462);
and AND4 (N15165, N15152, N7531, N4082, N9211);
nor NOR3 (N15166, N15146, N6127, N11749);
or OR2 (N15167, N15157, N12591);
xor XOR2 (N15168, N15161, N1150);
buf BUF1 (N15169, N15167);
xor XOR2 (N15170, N15164, N2902);
or OR2 (N15171, N15166, N3248);
xor XOR2 (N15172, N15162, N8013);
nand NAND2 (N15173, N15163, N7190);
nor NOR2 (N15174, N15171, N10686);
buf BUF1 (N15175, N15168);
or OR4 (N15176, N15175, N8403, N3624, N14598);
or OR4 (N15177, N15174, N11240, N8536, N13643);
and AND2 (N15178, N15148, N4855);
not NOT1 (N15179, N15158);
nor NOR2 (N15180, N15176, N5799);
xor XOR2 (N15181, N15178, N6061);
and AND3 (N15182, N15181, N8708, N982);
or OR4 (N15183, N15170, N7706, N14380, N3993);
nor NOR4 (N15184, N15151, N4396, N2390, N14689);
or OR4 (N15185, N15169, N6332, N10950, N5918);
or OR3 (N15186, N15184, N3648, N10503);
or OR4 (N15187, N15179, N1671, N12664, N10129);
buf BUF1 (N15188, N15182);
xor XOR2 (N15189, N15180, N12110);
buf BUF1 (N15190, N15173);
nand NAND3 (N15191, N15190, N11276, N13949);
or OR4 (N15192, N15191, N2114, N13583, N7512);
buf BUF1 (N15193, N15185);
nor NOR4 (N15194, N15183, N2590, N7390, N3895);
nor NOR3 (N15195, N15165, N12520, N14413);
and AND3 (N15196, N15195, N213, N3897);
or OR4 (N15197, N15193, N11644, N9568, N14490);
buf BUF1 (N15198, N15196);
nor NOR3 (N15199, N15172, N2286, N3868);
not NOT1 (N15200, N15197);
xor XOR2 (N15201, N15186, N2644);
not NOT1 (N15202, N15177);
buf BUF1 (N15203, N15192);
or OR3 (N15204, N15198, N4221, N1383);
not NOT1 (N15205, N15204);
nor NOR4 (N15206, N15187, N10521, N6080, N4820);
xor XOR2 (N15207, N15200, N3215);
buf BUF1 (N15208, N15202);
or OR3 (N15209, N15189, N14142, N100);
or OR3 (N15210, N15203, N8863, N12543);
or OR4 (N15211, N15205, N1361, N2733, N14923);
or OR3 (N15212, N15201, N14380, N7074);
buf BUF1 (N15213, N15206);
xor XOR2 (N15214, N15199, N7576);
not NOT1 (N15215, N15188);
buf BUF1 (N15216, N15209);
and AND3 (N15217, N15216, N6819, N10615);
nor NOR4 (N15218, N15208, N7327, N13673, N7596);
nor NOR2 (N15219, N15214, N1612);
nor NOR2 (N15220, N15207, N743);
nand NAND2 (N15221, N15220, N2191);
or OR2 (N15222, N15217, N2856);
buf BUF1 (N15223, N15211);
and AND4 (N15224, N15221, N11089, N9918, N8665);
and AND2 (N15225, N15194, N1572);
nand NAND2 (N15226, N15212, N10085);
not NOT1 (N15227, N15219);
nand NAND2 (N15228, N15218, N12795);
nand NAND4 (N15229, N15215, N8714, N5821, N215);
nor NOR2 (N15230, N15210, N8761);
or OR4 (N15231, N15230, N6785, N8432, N3194);
xor XOR2 (N15232, N15226, N6163);
buf BUF1 (N15233, N15232);
nor NOR4 (N15234, N15222, N441, N967, N2258);
and AND3 (N15235, N15213, N9626, N2822);
nand NAND2 (N15236, N15231, N9051);
nor NOR4 (N15237, N15227, N14995, N12409, N11449);
and AND4 (N15238, N15236, N14559, N8531, N6329);
and AND2 (N15239, N15237, N9642);
and AND2 (N15240, N15223, N3133);
and AND2 (N15241, N15225, N3518);
nor NOR4 (N15242, N15239, N6780, N13395, N7818);
and AND3 (N15243, N15242, N10461, N7652);
nand NAND4 (N15244, N15238, N2058, N8016, N9);
xor XOR2 (N15245, N15241, N6601);
or OR4 (N15246, N15245, N13621, N11488, N14297);
buf BUF1 (N15247, N15240);
not NOT1 (N15248, N15233);
not NOT1 (N15249, N15228);
nor NOR3 (N15250, N15246, N11126, N1334);
not NOT1 (N15251, N15248);
or OR3 (N15252, N15247, N2546, N12304);
xor XOR2 (N15253, N15249, N5141);
and AND2 (N15254, N15250, N6435);
xor XOR2 (N15255, N15234, N12479);
buf BUF1 (N15256, N15253);
not NOT1 (N15257, N15254);
nor NOR2 (N15258, N15235, N4472);
or OR2 (N15259, N15244, N6656);
xor XOR2 (N15260, N15257, N5401);
or OR2 (N15261, N15260, N8644);
and AND4 (N15262, N15256, N14459, N10941, N1979);
nand NAND2 (N15263, N15262, N5616);
buf BUF1 (N15264, N15251);
xor XOR2 (N15265, N15258, N216);
nand NAND4 (N15266, N15255, N4067, N2506, N8588);
or OR3 (N15267, N15263, N13745, N3035);
not NOT1 (N15268, N15252);
or OR2 (N15269, N15267, N3567);
and AND4 (N15270, N15261, N7390, N12935, N58);
not NOT1 (N15271, N15270);
nor NOR2 (N15272, N15259, N619);
buf BUF1 (N15273, N15224);
not NOT1 (N15274, N15265);
xor XOR2 (N15275, N15273, N2715);
buf BUF1 (N15276, N15271);
not NOT1 (N15277, N15268);
nand NAND4 (N15278, N15272, N14411, N10533, N11106);
or OR3 (N15279, N15274, N762, N12538);
or OR2 (N15280, N15264, N356);
and AND4 (N15281, N15266, N5216, N6332, N6283);
and AND2 (N15282, N15229, N2867);
and AND4 (N15283, N15269, N3733, N7152, N5914);
nand NAND2 (N15284, N15276, N6083);
and AND3 (N15285, N15275, N943, N13224);
nor NOR2 (N15286, N15277, N12147);
or OR3 (N15287, N15281, N5920, N9204);
or OR3 (N15288, N15286, N1460, N8269);
nand NAND2 (N15289, N15279, N11784);
buf BUF1 (N15290, N15289);
or OR3 (N15291, N15280, N13484, N6107);
xor XOR2 (N15292, N15282, N10009);
xor XOR2 (N15293, N15288, N6937);
xor XOR2 (N15294, N15293, N13111);
buf BUF1 (N15295, N15290);
xor XOR2 (N15296, N15292, N13899);
xor XOR2 (N15297, N15283, N12519);
xor XOR2 (N15298, N15296, N11477);
or OR4 (N15299, N15284, N3239, N4878, N11286);
buf BUF1 (N15300, N15287);
buf BUF1 (N15301, N15291);
xor XOR2 (N15302, N15295, N9656);
and AND2 (N15303, N15298, N7033);
buf BUF1 (N15304, N15297);
and AND2 (N15305, N15278, N5754);
xor XOR2 (N15306, N15285, N15049);
not NOT1 (N15307, N15243);
nor NOR4 (N15308, N15303, N13231, N3760, N9317);
buf BUF1 (N15309, N15307);
xor XOR2 (N15310, N15309, N7537);
xor XOR2 (N15311, N15294, N5679);
nand NAND3 (N15312, N15305, N7052, N3861);
and AND3 (N15313, N15299, N8139, N501);
nor NOR4 (N15314, N15313, N5458, N4717, N6065);
not NOT1 (N15315, N15311);
buf BUF1 (N15316, N15310);
not NOT1 (N15317, N15314);
and AND2 (N15318, N15302, N5837);
buf BUF1 (N15319, N15306);
nand NAND4 (N15320, N15316, N12308, N2501, N2394);
buf BUF1 (N15321, N15315);
xor XOR2 (N15322, N15321, N5657);
nand NAND2 (N15323, N15312, N374);
and AND2 (N15324, N15323, N1708);
and AND4 (N15325, N15317, N11376, N11682, N11423);
not NOT1 (N15326, N15320);
and AND3 (N15327, N15322, N2448, N7697);
xor XOR2 (N15328, N15326, N7508);
buf BUF1 (N15329, N15327);
xor XOR2 (N15330, N15324, N3329);
xor XOR2 (N15331, N15319, N9869);
buf BUF1 (N15332, N15304);
nand NAND3 (N15333, N15332, N15201, N3642);
not NOT1 (N15334, N15300);
not NOT1 (N15335, N15333);
buf BUF1 (N15336, N15328);
not NOT1 (N15337, N15330);
nand NAND3 (N15338, N15325, N5368, N4168);
and AND4 (N15339, N15331, N12889, N12653, N1221);
nand NAND3 (N15340, N15318, N6054, N14032);
nor NOR3 (N15341, N15301, N5952, N11900);
or OR3 (N15342, N15308, N11258, N13597);
buf BUF1 (N15343, N15335);
not NOT1 (N15344, N15336);
not NOT1 (N15345, N15334);
and AND3 (N15346, N15337, N2442, N7554);
buf BUF1 (N15347, N15344);
nor NOR3 (N15348, N15338, N3044, N2995);
xor XOR2 (N15349, N15345, N13026);
nand NAND2 (N15350, N15348, N8025);
xor XOR2 (N15351, N15347, N3595);
nand NAND4 (N15352, N15346, N1863, N7458, N9322);
xor XOR2 (N15353, N15342, N8085);
nor NOR3 (N15354, N15341, N14475, N1979);
or OR4 (N15355, N15351, N14095, N12403, N3848);
buf BUF1 (N15356, N15339);
nor NOR2 (N15357, N15356, N147);
nor NOR4 (N15358, N15355, N5391, N5308, N762);
not NOT1 (N15359, N15354);
and AND4 (N15360, N15353, N6632, N8810, N12817);
nor NOR4 (N15361, N15349, N12498, N10443, N1297);
xor XOR2 (N15362, N15357, N4335);
nor NOR4 (N15363, N15340, N1420, N11853, N109);
nor NOR4 (N15364, N15352, N11408, N10969, N974);
nor NOR4 (N15365, N15364, N11306, N13131, N9731);
buf BUF1 (N15366, N15329);
or OR4 (N15367, N15343, N10887, N2508, N401);
buf BUF1 (N15368, N15366);
and AND2 (N15369, N15359, N8639);
and AND3 (N15370, N15363, N13588, N15312);
not NOT1 (N15371, N15370);
buf BUF1 (N15372, N15365);
xor XOR2 (N15373, N15362, N8164);
or OR4 (N15374, N15367, N2718, N7420, N3532);
xor XOR2 (N15375, N15358, N12270);
not NOT1 (N15376, N15374);
nor NOR3 (N15377, N15375, N12807, N12276);
nor NOR4 (N15378, N15361, N4662, N14802, N11583);
and AND4 (N15379, N15372, N13224, N2101, N15085);
nand NAND4 (N15380, N15371, N719, N4249, N11920);
or OR4 (N15381, N15369, N4364, N2615, N5594);
nor NOR2 (N15382, N15377, N8986);
xor XOR2 (N15383, N15381, N2610);
and AND4 (N15384, N15379, N5444, N4641, N11285);
buf BUF1 (N15385, N15360);
xor XOR2 (N15386, N15383, N13634);
or OR4 (N15387, N15376, N6254, N15029, N7400);
or OR4 (N15388, N15385, N11494, N10684, N1429);
buf BUF1 (N15389, N15387);
not NOT1 (N15390, N15368);
and AND4 (N15391, N15380, N1282, N1641, N9470);
nor NOR3 (N15392, N15390, N8718, N9689);
and AND2 (N15393, N15378, N3732);
or OR2 (N15394, N15350, N11927);
not NOT1 (N15395, N15388);
buf BUF1 (N15396, N15393);
or OR4 (N15397, N15391, N3854, N7928, N7011);
buf BUF1 (N15398, N15395);
nor NOR2 (N15399, N15396, N12511);
nand NAND2 (N15400, N15397, N10219);
xor XOR2 (N15401, N15399, N9025);
not NOT1 (N15402, N15400);
nand NAND3 (N15403, N15373, N129, N13188);
or OR3 (N15404, N15382, N2552, N1220);
nand NAND4 (N15405, N15389, N11627, N195, N4739);
nand NAND3 (N15406, N15404, N4536, N2329);
and AND4 (N15407, N15401, N121, N2903, N13318);
xor XOR2 (N15408, N15384, N13482);
or OR2 (N15409, N15394, N8129);
buf BUF1 (N15410, N15402);
xor XOR2 (N15411, N15406, N589);
and AND3 (N15412, N15405, N1657, N9136);
buf BUF1 (N15413, N15392);
and AND3 (N15414, N15412, N7184, N9909);
and AND2 (N15415, N15403, N468);
buf BUF1 (N15416, N15410);
or OR4 (N15417, N15413, N2997, N1119, N446);
buf BUF1 (N15418, N15415);
buf BUF1 (N15419, N15414);
or OR2 (N15420, N15409, N12307);
and AND4 (N15421, N15420, N2476, N3571, N5055);
buf BUF1 (N15422, N15386);
not NOT1 (N15423, N15419);
and AND3 (N15424, N15408, N1762, N6391);
nor NOR2 (N15425, N15421, N10765);
buf BUF1 (N15426, N15423);
or OR4 (N15427, N15416, N13721, N1598, N11041);
buf BUF1 (N15428, N15418);
or OR2 (N15429, N15427, N1940);
buf BUF1 (N15430, N15398);
buf BUF1 (N15431, N15428);
xor XOR2 (N15432, N15424, N7135);
xor XOR2 (N15433, N15430, N2286);
nor NOR4 (N15434, N15417, N2906, N14526, N8872);
not NOT1 (N15435, N15422);
nor NOR3 (N15436, N15411, N12418, N9242);
buf BUF1 (N15437, N15426);
not NOT1 (N15438, N15433);
not NOT1 (N15439, N15438);
not NOT1 (N15440, N15407);
xor XOR2 (N15441, N15434, N5840);
or OR3 (N15442, N15432, N8852, N9956);
or OR4 (N15443, N15431, N8792, N11582, N5778);
or OR3 (N15444, N15440, N2457, N13179);
nor NOR4 (N15445, N15425, N5795, N7050, N2868);
xor XOR2 (N15446, N15436, N8865);
not NOT1 (N15447, N15443);
xor XOR2 (N15448, N15429, N13546);
nand NAND2 (N15449, N15446, N2908);
xor XOR2 (N15450, N15441, N13757);
xor XOR2 (N15451, N15447, N1131);
nand NAND3 (N15452, N15449, N2705, N4811);
nand NAND3 (N15453, N15448, N2919, N8437);
nand NAND3 (N15454, N15453, N1421, N6610);
and AND2 (N15455, N15452, N5980);
or OR2 (N15456, N15442, N4022);
nand NAND3 (N15457, N15450, N4838, N5001);
or OR3 (N15458, N15444, N1601, N11492);
not NOT1 (N15459, N15457);
xor XOR2 (N15460, N15454, N9533);
xor XOR2 (N15461, N15456, N10611);
and AND3 (N15462, N15437, N2039, N477);
and AND2 (N15463, N15445, N8498);
or OR4 (N15464, N15451, N3129, N10672, N9591);
nand NAND2 (N15465, N15459, N2197);
buf BUF1 (N15466, N15458);
xor XOR2 (N15467, N15460, N13844);
or OR3 (N15468, N15466, N8419, N3227);
nand NAND4 (N15469, N15463, N6519, N12406, N10570);
xor XOR2 (N15470, N15469, N7748);
nand NAND3 (N15471, N15464, N9286, N11141);
nor NOR2 (N15472, N15471, N7538);
buf BUF1 (N15473, N15468);
nor NOR2 (N15474, N15435, N14698);
nand NAND3 (N15475, N15465, N9204, N13137);
and AND3 (N15476, N15474, N6244, N13375);
buf BUF1 (N15477, N15475);
nand NAND2 (N15478, N15467, N1624);
and AND3 (N15479, N15455, N10867, N13895);
or OR4 (N15480, N15479, N4238, N5087, N4238);
not NOT1 (N15481, N15473);
and AND2 (N15482, N15476, N15268);
not NOT1 (N15483, N15478);
xor XOR2 (N15484, N15477, N11532);
nor NOR3 (N15485, N15439, N5877, N13567);
nor NOR3 (N15486, N15480, N8413, N1601);
buf BUF1 (N15487, N15486);
and AND3 (N15488, N15484, N7060, N4970);
xor XOR2 (N15489, N15470, N11074);
or OR3 (N15490, N15487, N6332, N7409);
nor NOR2 (N15491, N15461, N11703);
buf BUF1 (N15492, N15472);
nor NOR3 (N15493, N15489, N6702, N12323);
xor XOR2 (N15494, N15462, N8577);
nor NOR4 (N15495, N15490, N127, N13324, N8627);
or OR3 (N15496, N15492, N920, N7413);
not NOT1 (N15497, N15481);
or OR4 (N15498, N15491, N7028, N12636, N10825);
xor XOR2 (N15499, N15493, N10332);
not NOT1 (N15500, N15495);
and AND3 (N15501, N15496, N2632, N7091);
and AND2 (N15502, N15483, N7685);
buf BUF1 (N15503, N15488);
buf BUF1 (N15504, N15482);
not NOT1 (N15505, N15499);
buf BUF1 (N15506, N15485);
and AND2 (N15507, N15504, N13904);
nor NOR3 (N15508, N15507, N4719, N12502);
nand NAND2 (N15509, N15503, N9817);
buf BUF1 (N15510, N15501);
buf BUF1 (N15511, N15502);
xor XOR2 (N15512, N15509, N2030);
xor XOR2 (N15513, N15506, N8075);
xor XOR2 (N15514, N15500, N4197);
or OR4 (N15515, N15511, N11378, N6054, N1169);
or OR3 (N15516, N15514, N10608, N3448);
not NOT1 (N15517, N15512);
not NOT1 (N15518, N15517);
or OR4 (N15519, N15510, N6030, N10348, N12501);
nor NOR2 (N15520, N15516, N3819);
or OR2 (N15521, N15498, N7477);
or OR2 (N15522, N15497, N14245);
nand NAND3 (N15523, N15520, N464, N4875);
and AND4 (N15524, N15494, N3519, N3606, N3709);
or OR2 (N15525, N15518, N14442);
and AND3 (N15526, N15524, N12547, N3767);
not NOT1 (N15527, N15525);
xor XOR2 (N15528, N15523, N6868);
not NOT1 (N15529, N15526);
and AND4 (N15530, N15528, N14303, N9232, N5503);
not NOT1 (N15531, N15521);
or OR4 (N15532, N15529, N15375, N2424, N12853);
or OR4 (N15533, N15515, N9389, N703, N9671);
or OR4 (N15534, N15532, N14030, N5793, N56);
buf BUF1 (N15535, N15531);
nor NOR2 (N15536, N15505, N2695);
or OR3 (N15537, N15530, N1395, N94);
nor NOR4 (N15538, N15508, N5316, N7485, N6456);
nand NAND3 (N15539, N15533, N12556, N14029);
not NOT1 (N15540, N15513);
and AND2 (N15541, N15539, N14024);
xor XOR2 (N15542, N15541, N4775);
not NOT1 (N15543, N15519);
nor NOR4 (N15544, N15527, N13451, N1630, N8435);
and AND4 (N15545, N15543, N1323, N13028, N4696);
nand NAND3 (N15546, N15544, N2838, N1081);
not NOT1 (N15547, N15545);
and AND2 (N15548, N15538, N8913);
nand NAND2 (N15549, N15542, N13355);
buf BUF1 (N15550, N15535);
not NOT1 (N15551, N15537);
nand NAND3 (N15552, N15522, N2782, N6185);
nand NAND4 (N15553, N15550, N3957, N8459, N9851);
buf BUF1 (N15554, N15552);
nand NAND2 (N15555, N15553, N3053);
xor XOR2 (N15556, N15549, N15316);
not NOT1 (N15557, N15540);
nand NAND3 (N15558, N15547, N941, N12585);
nor NOR2 (N15559, N15551, N4342);
and AND4 (N15560, N15536, N2840, N872, N11593);
buf BUF1 (N15561, N15554);
nand NAND2 (N15562, N15561, N1752);
and AND4 (N15563, N15555, N15397, N5179, N2759);
nor NOR4 (N15564, N15558, N4949, N12706, N4396);
not NOT1 (N15565, N15548);
xor XOR2 (N15566, N15564, N13224);
or OR3 (N15567, N15546, N10191, N12306);
not NOT1 (N15568, N15565);
and AND4 (N15569, N15534, N6218, N5571, N7246);
or OR2 (N15570, N15556, N9669);
nor NOR3 (N15571, N15569, N14288, N11432);
buf BUF1 (N15572, N15570);
and AND2 (N15573, N15571, N8096);
not NOT1 (N15574, N15566);
nor NOR4 (N15575, N15568, N1201, N443, N5938);
not NOT1 (N15576, N15572);
and AND4 (N15577, N15567, N12160, N13873, N2225);
or OR2 (N15578, N15576, N2159);
not NOT1 (N15579, N15578);
and AND2 (N15580, N15563, N13615);
nand NAND3 (N15581, N15574, N3674, N12153);
and AND4 (N15582, N15581, N7832, N10389, N8434);
or OR4 (N15583, N15577, N6512, N4529, N14260);
not NOT1 (N15584, N15573);
or OR3 (N15585, N15575, N5770, N424);
or OR2 (N15586, N15582, N11825);
or OR3 (N15587, N15559, N4163, N13935);
and AND4 (N15588, N15580, N1003, N7144, N5052);
buf BUF1 (N15589, N15579);
xor XOR2 (N15590, N15560, N114);
nor NOR2 (N15591, N15562, N7216);
nor NOR3 (N15592, N15591, N13709, N6326);
nor NOR3 (N15593, N15583, N13430, N1224);
nand NAND2 (N15594, N15590, N6107);
nand NAND2 (N15595, N15588, N10005);
and AND2 (N15596, N15585, N2415);
xor XOR2 (N15597, N15584, N6360);
buf BUF1 (N15598, N15557);
nand NAND2 (N15599, N15589, N5706);
and AND3 (N15600, N15592, N2396, N10319);
or OR4 (N15601, N15586, N1144, N8255, N5756);
and AND3 (N15602, N15587, N1493, N9373);
nand NAND3 (N15603, N15597, N4224, N5162);
xor XOR2 (N15604, N15600, N10833);
nor NOR3 (N15605, N15603, N14720, N11683);
and AND3 (N15606, N15605, N7498, N7402);
or OR3 (N15607, N15593, N15206, N9517);
xor XOR2 (N15608, N15599, N2519);
not NOT1 (N15609, N15595);
buf BUF1 (N15610, N15596);
and AND4 (N15611, N15609, N13074, N941, N4246);
nand NAND2 (N15612, N15601, N14731);
and AND4 (N15613, N15607, N9617, N15148, N3532);
buf BUF1 (N15614, N15594);
buf BUF1 (N15615, N15598);
xor XOR2 (N15616, N15604, N5614);
and AND4 (N15617, N15616, N5157, N1787, N12196);
or OR4 (N15618, N15617, N5395, N11063, N15398);
or OR2 (N15619, N15614, N5903);
xor XOR2 (N15620, N15611, N10605);
not NOT1 (N15621, N15619);
nand NAND3 (N15622, N15618, N8945, N2765);
nor NOR2 (N15623, N15602, N9211);
nor NOR4 (N15624, N15621, N15013, N1655, N2013);
nand NAND2 (N15625, N15623, N14235);
nor NOR2 (N15626, N15612, N5748);
or OR4 (N15627, N15622, N4077, N14887, N8254);
not NOT1 (N15628, N15615);
and AND2 (N15629, N15620, N10984);
buf BUF1 (N15630, N15625);
buf BUF1 (N15631, N15610);
or OR3 (N15632, N15613, N5896, N1295);
or OR3 (N15633, N15630, N2878, N12937);
xor XOR2 (N15634, N15633, N2795);
nand NAND4 (N15635, N15631, N10002, N12726, N7860);
nor NOR2 (N15636, N15629, N6611);
xor XOR2 (N15637, N15624, N15622);
buf BUF1 (N15638, N15632);
xor XOR2 (N15639, N15637, N251);
buf BUF1 (N15640, N15635);
and AND2 (N15641, N15626, N11588);
nor NOR4 (N15642, N15640, N7061, N10558, N2515);
nor NOR2 (N15643, N15636, N5469);
and AND3 (N15644, N15639, N1682, N761);
xor XOR2 (N15645, N15638, N12571);
xor XOR2 (N15646, N15641, N3112);
nand NAND4 (N15647, N15646, N15331, N310, N14395);
nand NAND2 (N15648, N15628, N11436);
and AND4 (N15649, N15627, N818, N15367, N6594);
or OR3 (N15650, N15648, N1726, N12933);
not NOT1 (N15651, N15606);
and AND4 (N15652, N15608, N209, N5681, N11689);
not NOT1 (N15653, N15642);
xor XOR2 (N15654, N15645, N7939);
buf BUF1 (N15655, N15634);
nor NOR3 (N15656, N15644, N12537, N1874);
or OR3 (N15657, N15653, N9992, N7566);
buf BUF1 (N15658, N15647);
and AND4 (N15659, N15649, N9464, N12424, N1027);
nor NOR4 (N15660, N15654, N13069, N9263, N2670);
xor XOR2 (N15661, N15652, N9483);
nor NOR4 (N15662, N15658, N1949, N9196, N9166);
nor NOR3 (N15663, N15661, N638, N3742);
not NOT1 (N15664, N15657);
and AND3 (N15665, N15663, N1888, N2048);
xor XOR2 (N15666, N15660, N11169);
xor XOR2 (N15667, N15662, N10637);
and AND2 (N15668, N15665, N1196);
buf BUF1 (N15669, N15650);
buf BUF1 (N15670, N15651);
nor NOR3 (N15671, N15669, N10551, N8059);
xor XOR2 (N15672, N15666, N6951);
xor XOR2 (N15673, N15643, N3466);
xor XOR2 (N15674, N15656, N13285);
and AND3 (N15675, N15673, N12657, N8340);
nand NAND2 (N15676, N15671, N4411);
xor XOR2 (N15677, N15675, N2997);
nand NAND3 (N15678, N15670, N13657, N4434);
nand NAND2 (N15679, N15664, N7570);
buf BUF1 (N15680, N15668);
and AND4 (N15681, N15679, N12799, N9659, N15663);
nor NOR2 (N15682, N15678, N10630);
not NOT1 (N15683, N15682);
not NOT1 (N15684, N15655);
nand NAND3 (N15685, N15667, N2214, N758);
nor NOR3 (N15686, N15683, N15380, N7737);
nor NOR2 (N15687, N15684, N9554);
nor NOR3 (N15688, N15681, N10349, N10913);
not NOT1 (N15689, N15680);
nor NOR4 (N15690, N15686, N9269, N4443, N14748);
or OR3 (N15691, N15688, N14895, N5552);
and AND3 (N15692, N15691, N11932, N8145);
and AND2 (N15693, N15689, N4363);
and AND2 (N15694, N15687, N5016);
buf BUF1 (N15695, N15685);
xor XOR2 (N15696, N15676, N2582);
and AND4 (N15697, N15696, N1532, N6027, N7302);
buf BUF1 (N15698, N15693);
buf BUF1 (N15699, N15674);
buf BUF1 (N15700, N15672);
and AND2 (N15701, N15659, N4735);
nor NOR3 (N15702, N15692, N1808, N13125);
or OR2 (N15703, N15699, N2800);
not NOT1 (N15704, N15697);
nor NOR3 (N15705, N15695, N4047, N13238);
or OR4 (N15706, N15690, N15629, N14888, N5550);
buf BUF1 (N15707, N15698);
nand NAND3 (N15708, N15706, N4769, N1977);
and AND2 (N15709, N15708, N9834);
or OR3 (N15710, N15704, N14152, N6019);
nand NAND3 (N15711, N15703, N613, N7164);
or OR2 (N15712, N15702, N12110);
xor XOR2 (N15713, N15705, N8516);
and AND4 (N15714, N15700, N6953, N14887, N7726);
nand NAND3 (N15715, N15713, N12353, N3638);
nor NOR4 (N15716, N15714, N9509, N5827, N5376);
not NOT1 (N15717, N15715);
and AND3 (N15718, N15707, N1754, N11973);
nand NAND3 (N15719, N15718, N2517, N10251);
nor NOR2 (N15720, N15677, N857);
buf BUF1 (N15721, N15709);
or OR4 (N15722, N15721, N5740, N12548, N1857);
buf BUF1 (N15723, N15711);
nand NAND3 (N15724, N15717, N414, N3532);
or OR4 (N15725, N15723, N15355, N2092, N8578);
nor NOR4 (N15726, N15719, N9745, N15177, N13684);
xor XOR2 (N15727, N15724, N12871);
xor XOR2 (N15728, N15701, N14340);
or OR3 (N15729, N15710, N8771, N14812);
or OR4 (N15730, N15726, N9358, N9754, N2008);
xor XOR2 (N15731, N15716, N6962);
or OR2 (N15732, N15720, N13079);
buf BUF1 (N15733, N15725);
nor NOR4 (N15734, N15732, N1661, N13005, N2212);
nand NAND2 (N15735, N15730, N3004);
and AND3 (N15736, N15735, N9804, N488);
nand NAND4 (N15737, N15694, N9030, N2159, N871);
nand NAND3 (N15738, N15737, N9611, N8977);
and AND3 (N15739, N15734, N1158, N8407);
and AND3 (N15740, N15739, N13133, N2701);
not NOT1 (N15741, N15722);
and AND2 (N15742, N15731, N8690);
and AND3 (N15743, N15729, N7775, N1907);
xor XOR2 (N15744, N15741, N11428);
nand NAND2 (N15745, N15736, N3499);
nand NAND4 (N15746, N15742, N13691, N11472, N276);
nand NAND3 (N15747, N15743, N9741, N5646);
buf BUF1 (N15748, N15733);
nor NOR3 (N15749, N15748, N8024, N14165);
xor XOR2 (N15750, N15746, N13071);
or OR2 (N15751, N15712, N3933);
and AND4 (N15752, N15749, N5046, N5584, N2208);
xor XOR2 (N15753, N15745, N1816);
nor NOR3 (N15754, N15738, N8717, N5492);
buf BUF1 (N15755, N15744);
buf BUF1 (N15756, N15750);
buf BUF1 (N15757, N15754);
buf BUF1 (N15758, N15727);
and AND4 (N15759, N15756, N13843, N14825, N699);
and AND3 (N15760, N15752, N5390, N14519);
nand NAND2 (N15761, N15759, N1679);
buf BUF1 (N15762, N15751);
nand NAND4 (N15763, N15753, N1634, N4048, N6743);
or OR4 (N15764, N15761, N15673, N8878, N11077);
nand NAND2 (N15765, N15760, N952);
or OR3 (N15766, N15763, N14537, N4197);
nand NAND4 (N15767, N15728, N11658, N9042, N10813);
buf BUF1 (N15768, N15755);
nand NAND2 (N15769, N15740, N9879);
nor NOR3 (N15770, N15767, N13266, N4734);
and AND3 (N15771, N15764, N6220, N15470);
buf BUF1 (N15772, N15758);
xor XOR2 (N15773, N15766, N5668);
nand NAND4 (N15774, N15771, N2779, N8347, N8231);
nor NOR3 (N15775, N15769, N1151, N2023);
nand NAND3 (N15776, N15757, N7100, N10887);
or OR3 (N15777, N15776, N5279, N1297);
or OR2 (N15778, N15770, N1260);
buf BUF1 (N15779, N15762);
xor XOR2 (N15780, N15777, N14800);
nor NOR2 (N15781, N15775, N5480);
and AND2 (N15782, N15768, N13189);
buf BUF1 (N15783, N15780);
xor XOR2 (N15784, N15782, N9081);
nor NOR2 (N15785, N15781, N5641);
nor NOR2 (N15786, N15779, N12574);
nor NOR3 (N15787, N15772, N14555, N11633);
buf BUF1 (N15788, N15747);
not NOT1 (N15789, N15787);
or OR4 (N15790, N15765, N6542, N11623, N11038);
nand NAND2 (N15791, N15783, N10631);
xor XOR2 (N15792, N15790, N8182);
nand NAND2 (N15793, N15788, N8328);
not NOT1 (N15794, N15791);
nor NOR4 (N15795, N15778, N2445, N7462, N12352);
and AND3 (N15796, N15789, N6061, N2049);
xor XOR2 (N15797, N15795, N2897);
not NOT1 (N15798, N15784);
xor XOR2 (N15799, N15798, N696);
and AND2 (N15800, N15785, N10525);
or OR4 (N15801, N15794, N14971, N1146, N11972);
not NOT1 (N15802, N15801);
or OR2 (N15803, N15796, N12485);
not NOT1 (N15804, N15774);
buf BUF1 (N15805, N15786);
not NOT1 (N15806, N15792);
or OR3 (N15807, N15806, N13286, N14248);
buf BUF1 (N15808, N15793);
nor NOR3 (N15809, N15799, N8191, N418);
buf BUF1 (N15810, N15804);
buf BUF1 (N15811, N15809);
or OR3 (N15812, N15811, N1384, N670);
nand NAND3 (N15813, N15810, N11328, N4870);
or OR3 (N15814, N15805, N11331, N5668);
nand NAND4 (N15815, N15813, N14326, N15125, N11398);
not NOT1 (N15816, N15807);
nand NAND2 (N15817, N15812, N5857);
and AND4 (N15818, N15816, N3785, N4032, N171);
not NOT1 (N15819, N15817);
buf BUF1 (N15820, N15808);
xor XOR2 (N15821, N15814, N8466);
xor XOR2 (N15822, N15820, N14596);
xor XOR2 (N15823, N15773, N4423);
not NOT1 (N15824, N15818);
buf BUF1 (N15825, N15821);
nor NOR4 (N15826, N15823, N4375, N7482, N9816);
buf BUF1 (N15827, N15819);
or OR3 (N15828, N15827, N5636, N14778);
nand NAND4 (N15829, N15828, N14499, N15660, N1582);
buf BUF1 (N15830, N15824);
nand NAND3 (N15831, N15815, N14627, N13794);
and AND4 (N15832, N15825, N2093, N7060, N3990);
and AND3 (N15833, N15832, N10746, N6572);
nand NAND3 (N15834, N15826, N9434, N1425);
not NOT1 (N15835, N15833);
and AND4 (N15836, N15800, N3216, N10073, N164);
nor NOR4 (N15837, N15831, N12460, N13243, N8832);
nand NAND3 (N15838, N15836, N411, N11113);
buf BUF1 (N15839, N15835);
xor XOR2 (N15840, N15829, N11435);
nor NOR3 (N15841, N15830, N6234, N14777);
nor NOR2 (N15842, N15802, N15217);
nor NOR3 (N15843, N15797, N13677, N4495);
or OR3 (N15844, N15843, N13494, N11924);
nor NOR3 (N15845, N15838, N1818, N14085);
or OR4 (N15846, N15839, N231, N12943, N14686);
nor NOR2 (N15847, N15842, N12804);
and AND4 (N15848, N15845, N6340, N5640, N11444);
or OR3 (N15849, N15834, N9362, N12435);
nand NAND4 (N15850, N15846, N2242, N11782, N9484);
buf BUF1 (N15851, N15847);
or OR3 (N15852, N15851, N6950, N2256);
buf BUF1 (N15853, N15840);
xor XOR2 (N15854, N15837, N6761);
buf BUF1 (N15855, N15844);
buf BUF1 (N15856, N15855);
and AND4 (N15857, N15822, N90, N12455, N10387);
and AND3 (N15858, N15803, N8374, N11365);
not NOT1 (N15859, N15858);
xor XOR2 (N15860, N15857, N9105);
buf BUF1 (N15861, N15853);
and AND2 (N15862, N15860, N2494);
nor NOR2 (N15863, N15862, N2803);
buf BUF1 (N15864, N15841);
nand NAND4 (N15865, N15848, N10609, N3599, N6461);
buf BUF1 (N15866, N15864);
nand NAND3 (N15867, N15863, N12556, N15084);
buf BUF1 (N15868, N15865);
or OR4 (N15869, N15852, N7923, N8231, N1509);
or OR3 (N15870, N15849, N14144, N3757);
or OR2 (N15871, N15868, N12564);
and AND3 (N15872, N15867, N9844, N12079);
not NOT1 (N15873, N15856);
nand NAND3 (N15874, N15870, N1118, N11114);
buf BUF1 (N15875, N15866);
nand NAND2 (N15876, N15854, N4876);
and AND2 (N15877, N15872, N13429);
and AND2 (N15878, N15859, N3033);
nand NAND2 (N15879, N15871, N5615);
nand NAND4 (N15880, N15878, N9776, N7155, N9349);
and AND3 (N15881, N15879, N6064, N13912);
xor XOR2 (N15882, N15881, N13203);
or OR4 (N15883, N15882, N1075, N2975, N7029);
xor XOR2 (N15884, N15883, N14290);
and AND2 (N15885, N15877, N9884);
or OR3 (N15886, N15850, N5271, N2330);
buf BUF1 (N15887, N15880);
and AND4 (N15888, N15886, N10059, N904, N1845);
nand NAND2 (N15889, N15869, N15797);
nor NOR4 (N15890, N15888, N10517, N125, N12723);
and AND2 (N15891, N15876, N11538);
buf BUF1 (N15892, N15874);
buf BUF1 (N15893, N15884);
nand NAND4 (N15894, N15889, N11860, N7897, N12402);
nor NOR4 (N15895, N15890, N11753, N5971, N11456);
nor NOR2 (N15896, N15894, N4435);
or OR2 (N15897, N15861, N6450);
nand NAND3 (N15898, N15891, N10510, N8220);
nor NOR3 (N15899, N15885, N3868, N15322);
buf BUF1 (N15900, N15895);
or OR3 (N15901, N15893, N9342, N6073);
or OR2 (N15902, N15901, N14543);
and AND2 (N15903, N15896, N4318);
nand NAND4 (N15904, N15903, N923, N4372, N12747);
nor NOR2 (N15905, N15875, N6623);
buf BUF1 (N15906, N15873);
and AND2 (N15907, N15887, N9272);
and AND4 (N15908, N15904, N7594, N14890, N15271);
nand NAND2 (N15909, N15900, N3781);
nand NAND2 (N15910, N15909, N1628);
or OR3 (N15911, N15906, N15850, N13971);
buf BUF1 (N15912, N15897);
not NOT1 (N15913, N15908);
and AND3 (N15914, N15912, N1877, N10282);
nor NOR2 (N15915, N15898, N3239);
xor XOR2 (N15916, N15910, N5336);
and AND3 (N15917, N15913, N513, N14541);
nor NOR2 (N15918, N15916, N8005);
nor NOR2 (N15919, N15911, N9255);
nand NAND4 (N15920, N15914, N945, N12712, N7858);
xor XOR2 (N15921, N15907, N7897);
xor XOR2 (N15922, N15892, N4408);
xor XOR2 (N15923, N15918, N9894);
or OR3 (N15924, N15921, N5821, N7113);
not NOT1 (N15925, N15922);
nor NOR2 (N15926, N15925, N12917);
not NOT1 (N15927, N15926);
or OR4 (N15928, N15905, N13222, N11479, N12493);
or OR2 (N15929, N15902, N15182);
nor NOR4 (N15930, N15924, N3020, N10847, N12242);
buf BUF1 (N15931, N15927);
xor XOR2 (N15932, N15919, N13823);
nand NAND4 (N15933, N15928, N4080, N12575, N1818);
buf BUF1 (N15934, N15929);
nor NOR2 (N15935, N15932, N5688);
or OR3 (N15936, N15917, N14793, N14296);
nand NAND3 (N15937, N15899, N15827, N2813);
nand NAND3 (N15938, N15937, N5591, N15319);
or OR2 (N15939, N15930, N164);
or OR3 (N15940, N15934, N357, N473);
not NOT1 (N15941, N15920);
buf BUF1 (N15942, N15923);
buf BUF1 (N15943, N15915);
nand NAND4 (N15944, N15938, N7478, N503, N15543);
nor NOR4 (N15945, N15931, N10070, N13689, N13472);
nand NAND4 (N15946, N15935, N12646, N7780, N10426);
xor XOR2 (N15947, N15942, N624);
or OR4 (N15948, N15945, N7778, N5276, N10254);
not NOT1 (N15949, N15947);
not NOT1 (N15950, N15939);
nand NAND4 (N15951, N15950, N1576, N4809, N11493);
and AND3 (N15952, N15949, N8728, N5168);
or OR4 (N15953, N15952, N6188, N9466, N327);
xor XOR2 (N15954, N15946, N11395);
xor XOR2 (N15955, N15944, N6984);
buf BUF1 (N15956, N15941);
buf BUF1 (N15957, N15948);
nand NAND3 (N15958, N15954, N4433, N3388);
not NOT1 (N15959, N15936);
and AND4 (N15960, N15951, N4451, N2891, N3684);
xor XOR2 (N15961, N15958, N4081);
or OR2 (N15962, N15953, N7652);
or OR2 (N15963, N15955, N4584);
nor NOR3 (N15964, N15961, N1100, N11621);
nor NOR3 (N15965, N15940, N2904, N9847);
xor XOR2 (N15966, N15963, N14319);
or OR3 (N15967, N15956, N12220, N6502);
buf BUF1 (N15968, N15965);
nand NAND4 (N15969, N15966, N12898, N1113, N4483);
nor NOR2 (N15970, N15968, N13926);
and AND4 (N15971, N15960, N5630, N11845, N4858);
or OR2 (N15972, N15964, N10132);
nor NOR3 (N15973, N15967, N15777, N4659);
buf BUF1 (N15974, N15969);
nand NAND2 (N15975, N15971, N7506);
nor NOR3 (N15976, N15970, N5295, N15973);
nor NOR4 (N15977, N13984, N14291, N8925, N427);
and AND2 (N15978, N15974, N7516);
nand NAND3 (N15979, N15962, N8287, N15304);
buf BUF1 (N15980, N15943);
or OR2 (N15981, N15972, N7222);
and AND4 (N15982, N15957, N7373, N4072, N11367);
or OR4 (N15983, N15980, N2607, N5390, N9193);
xor XOR2 (N15984, N15982, N6922);
nor NOR4 (N15985, N15975, N12570, N13791, N9594);
nor NOR2 (N15986, N15983, N7556);
nand NAND4 (N15987, N15984, N12539, N8999, N10667);
buf BUF1 (N15988, N15959);
nand NAND4 (N15989, N15985, N2585, N9703, N5276);
and AND4 (N15990, N15988, N14425, N1326, N15777);
xor XOR2 (N15991, N15976, N8593);
nand NAND2 (N15992, N15981, N8231);
nand NAND2 (N15993, N15987, N14855);
and AND2 (N15994, N15989, N10556);
or OR2 (N15995, N15994, N1751);
nor NOR4 (N15996, N15993, N2779, N7249, N14421);
not NOT1 (N15997, N15990);
xor XOR2 (N15998, N15978, N3486);
and AND2 (N15999, N15995, N9204);
buf BUF1 (N16000, N15991);
and AND3 (N16001, N15933, N14707, N154);
nor NOR4 (N16002, N15998, N7421, N9350, N14228);
or OR4 (N16003, N15999, N8440, N6860, N10037);
nand NAND4 (N16004, N15997, N9650, N3722, N15387);
nand NAND3 (N16005, N15977, N5795, N13396);
nor NOR2 (N16006, N15996, N13287);
buf BUF1 (N16007, N16003);
xor XOR2 (N16008, N16000, N8812);
buf BUF1 (N16009, N16001);
xor XOR2 (N16010, N16005, N4242);
or OR3 (N16011, N16006, N4289, N7287);
not NOT1 (N16012, N16007);
and AND4 (N16013, N15986, N589, N6673, N4413);
not NOT1 (N16014, N16002);
and AND4 (N16015, N16004, N2189, N7866, N4369);
buf BUF1 (N16016, N16013);
and AND2 (N16017, N16009, N4925);
and AND2 (N16018, N16017, N2227);
buf BUF1 (N16019, N15979);
not NOT1 (N16020, N16018);
nor NOR4 (N16021, N16008, N8302, N15777, N6046);
and AND4 (N16022, N16014, N171, N15985, N13687);
or OR3 (N16023, N16015, N780, N9217);
not NOT1 (N16024, N16023);
nand NAND4 (N16025, N16022, N7526, N10680, N1688);
nand NAND4 (N16026, N16024, N6487, N1227, N13409);
xor XOR2 (N16027, N16012, N13345);
xor XOR2 (N16028, N16019, N5458);
not NOT1 (N16029, N16026);
buf BUF1 (N16030, N16016);
xor XOR2 (N16031, N16027, N382);
and AND3 (N16032, N16010, N14984, N13843);
or OR4 (N16033, N16028, N5819, N6852, N2033);
xor XOR2 (N16034, N16021, N8522);
buf BUF1 (N16035, N16029);
nand NAND2 (N16036, N16011, N15225);
nand NAND3 (N16037, N16025, N10077, N13219);
buf BUF1 (N16038, N16032);
nand NAND2 (N16039, N15992, N14236);
or OR3 (N16040, N16033, N3050, N1883);
or OR4 (N16041, N16030, N8092, N5494, N15787);
buf BUF1 (N16042, N16041);
not NOT1 (N16043, N16038);
not NOT1 (N16044, N16036);
nor NOR3 (N16045, N16043, N4613, N12857);
not NOT1 (N16046, N16034);
xor XOR2 (N16047, N16035, N13386);
and AND2 (N16048, N16047, N9249);
and AND3 (N16049, N16045, N3621, N6218);
xor XOR2 (N16050, N16048, N6847);
xor XOR2 (N16051, N16020, N224);
or OR2 (N16052, N16046, N8962);
and AND3 (N16053, N16040, N997, N14964);
nand NAND3 (N16054, N16044, N13428, N3717);
not NOT1 (N16055, N16049);
and AND3 (N16056, N16031, N1232, N8847);
and AND4 (N16057, N16052, N4492, N6059, N7269);
or OR3 (N16058, N16055, N11614, N8005);
not NOT1 (N16059, N16058);
and AND3 (N16060, N16042, N7824, N3429);
not NOT1 (N16061, N16051);
nand NAND2 (N16062, N16037, N424);
nand NAND3 (N16063, N16062, N2038, N7316);
xor XOR2 (N16064, N16054, N4254);
nor NOR3 (N16065, N16060, N12517, N4741);
nor NOR3 (N16066, N16059, N11071, N2143);
or OR2 (N16067, N16065, N5423);
buf BUF1 (N16068, N16056);
nor NOR4 (N16069, N16057, N4287, N2751, N8634);
nand NAND2 (N16070, N16039, N10673);
not NOT1 (N16071, N16070);
buf BUF1 (N16072, N16050);
nor NOR2 (N16073, N16069, N4758);
not NOT1 (N16074, N16067);
buf BUF1 (N16075, N16071);
nand NAND3 (N16076, N16074, N12255, N9346);
or OR4 (N16077, N16063, N7434, N4766, N12214);
xor XOR2 (N16078, N16075, N10547);
xor XOR2 (N16079, N16077, N4826);
or OR2 (N16080, N16061, N8148);
nand NAND3 (N16081, N16076, N4026, N5188);
nand NAND3 (N16082, N16078, N8612, N14671);
nor NOR2 (N16083, N16068, N9037);
buf BUF1 (N16084, N16066);
nor NOR2 (N16085, N16079, N1863);
buf BUF1 (N16086, N16064);
or OR3 (N16087, N16082, N2494, N4064);
xor XOR2 (N16088, N16081, N3671);
xor XOR2 (N16089, N16088, N2703);
xor XOR2 (N16090, N16085, N4945);
nand NAND3 (N16091, N16084, N9326, N11783);
nor NOR3 (N16092, N16080, N7171, N15592);
buf BUF1 (N16093, N16072);
buf BUF1 (N16094, N16083);
nor NOR3 (N16095, N16091, N10796, N2739);
nand NAND2 (N16096, N16053, N6963);
xor XOR2 (N16097, N16073, N3951);
nand NAND2 (N16098, N16096, N4420);
xor XOR2 (N16099, N16089, N15188);
or OR4 (N16100, N16092, N13910, N2721, N13943);
buf BUF1 (N16101, N16090);
or OR3 (N16102, N16101, N3860, N2057);
and AND4 (N16103, N16086, N5269, N4156, N2947);
nor NOR3 (N16104, N16099, N3190, N7348);
or OR4 (N16105, N16100, N11251, N9583, N13622);
or OR2 (N16106, N16093, N8321);
buf BUF1 (N16107, N16104);
buf BUF1 (N16108, N16097);
xor XOR2 (N16109, N16098, N14448);
buf BUF1 (N16110, N16102);
or OR4 (N16111, N16105, N8031, N5188, N12841);
not NOT1 (N16112, N16108);
and AND2 (N16113, N16111, N7889);
nor NOR4 (N16114, N16095, N1723, N6684, N15329);
not NOT1 (N16115, N16106);
nand NAND3 (N16116, N16110, N3452, N12009);
xor XOR2 (N16117, N16103, N3371);
nor NOR3 (N16118, N16114, N1379, N12261);
xor XOR2 (N16119, N16109, N2138);
or OR3 (N16120, N16115, N6185, N7502);
nand NAND2 (N16121, N16117, N13531);
not NOT1 (N16122, N16112);
buf BUF1 (N16123, N16122);
or OR4 (N16124, N16113, N8829, N11541, N200);
buf BUF1 (N16125, N16116);
and AND4 (N16126, N16120, N3607, N6759, N3646);
buf BUF1 (N16127, N16124);
buf BUF1 (N16128, N16125);
nand NAND4 (N16129, N16128, N15163, N2312, N8358);
xor XOR2 (N16130, N16126, N15825);
nor NOR4 (N16131, N16094, N10361, N3867, N9487);
and AND3 (N16132, N16107, N14171, N14881);
and AND3 (N16133, N16118, N9010, N7961);
or OR3 (N16134, N16133, N6508, N11420);
or OR4 (N16135, N16131, N10026, N12825, N14524);
nor NOR3 (N16136, N16087, N864, N9575);
not NOT1 (N16137, N16121);
nor NOR2 (N16138, N16129, N5354);
buf BUF1 (N16139, N16136);
nand NAND3 (N16140, N16139, N8441, N11460);
xor XOR2 (N16141, N16130, N9741);
and AND2 (N16142, N16137, N8603);
and AND2 (N16143, N16134, N13684);
and AND2 (N16144, N16143, N5951);
nor NOR4 (N16145, N16140, N10163, N5280, N3569);
nor NOR2 (N16146, N16132, N12041);
nand NAND2 (N16147, N16123, N1576);
xor XOR2 (N16148, N16147, N11967);
nor NOR2 (N16149, N16135, N1938);
or OR3 (N16150, N16145, N8922, N9981);
and AND4 (N16151, N16141, N12059, N9854, N7814);
nand NAND2 (N16152, N16146, N3335);
nor NOR4 (N16153, N16152, N2549, N11508, N14577);
nand NAND4 (N16154, N16149, N6746, N6871, N2141);
xor XOR2 (N16155, N16148, N5998);
not NOT1 (N16156, N16119);
not NOT1 (N16157, N16127);
not NOT1 (N16158, N16142);
xor XOR2 (N16159, N16154, N7884);
not NOT1 (N16160, N16157);
nor NOR4 (N16161, N16153, N4523, N9534, N4041);
and AND3 (N16162, N16161, N1823, N7575);
nor NOR4 (N16163, N16159, N7592, N2066, N13925);
nor NOR3 (N16164, N16156, N11353, N8006);
nand NAND3 (N16165, N16158, N12936, N5127);
nor NOR3 (N16166, N16163, N9716, N8741);
and AND3 (N16167, N16164, N11022, N6361);
nor NOR4 (N16168, N16160, N12953, N12601, N9202);
not NOT1 (N16169, N16150);
nor NOR3 (N16170, N16144, N15559, N3412);
buf BUF1 (N16171, N16151);
or OR4 (N16172, N16162, N8460, N1071, N7484);
not NOT1 (N16173, N16171);
nor NOR4 (N16174, N16172, N12596, N13529, N2675);
or OR2 (N16175, N16155, N702);
not NOT1 (N16176, N16169);
buf BUF1 (N16177, N16173);
or OR4 (N16178, N16165, N2440, N4087, N2051);
not NOT1 (N16179, N16178);
or OR4 (N16180, N16170, N3318, N908, N4982);
or OR2 (N16181, N16138, N2493);
nand NAND2 (N16182, N16179, N11327);
or OR4 (N16183, N16177, N789, N10477, N3930);
or OR3 (N16184, N16181, N11781, N13368);
xor XOR2 (N16185, N16168, N15143);
nand NAND4 (N16186, N16174, N12667, N4746, N341);
nand NAND4 (N16187, N16167, N7201, N6432, N12009);
not NOT1 (N16188, N16187);
and AND4 (N16189, N16184, N11377, N7231, N13467);
not NOT1 (N16190, N16188);
or OR3 (N16191, N16189, N12326, N3746);
and AND2 (N16192, N16183, N8865);
nand NAND4 (N16193, N16180, N15322, N14257, N7637);
or OR2 (N16194, N16166, N14073);
and AND3 (N16195, N16182, N8543, N2221);
xor XOR2 (N16196, N16185, N7784);
nor NOR4 (N16197, N16176, N1465, N3803, N4949);
not NOT1 (N16198, N16192);
or OR3 (N16199, N16191, N1582, N11969);
or OR4 (N16200, N16175, N16144, N795, N1241);
and AND3 (N16201, N16186, N7474, N5251);
nor NOR4 (N16202, N16200, N13640, N8511, N6212);
or OR4 (N16203, N16194, N5935, N8430, N9940);
nand NAND2 (N16204, N16190, N10533);
and AND4 (N16205, N16198, N6969, N14918, N8813);
xor XOR2 (N16206, N16202, N12808);
buf BUF1 (N16207, N16196);
buf BUF1 (N16208, N16206);
or OR3 (N16209, N16195, N8576, N471);
nor NOR3 (N16210, N16204, N8991, N4772);
or OR3 (N16211, N16205, N4226, N11495);
and AND3 (N16212, N16207, N5187, N2323);
or OR2 (N16213, N16201, N3427);
and AND3 (N16214, N16208, N1499, N1609);
nand NAND4 (N16215, N16212, N1423, N23, N93);
or OR3 (N16216, N16199, N5999, N11005);
nor NOR4 (N16217, N16216, N8078, N7879, N11226);
and AND3 (N16218, N16211, N8736, N8168);
nor NOR3 (N16219, N16209, N2606, N12344);
and AND3 (N16220, N16193, N11441, N13807);
xor XOR2 (N16221, N16218, N8289);
nor NOR2 (N16222, N16214, N14373);
nand NAND4 (N16223, N16222, N13834, N16114, N4489);
xor XOR2 (N16224, N16221, N360);
nand NAND3 (N16225, N16224, N15545, N7056);
or OR4 (N16226, N16197, N8238, N4485, N14078);
and AND3 (N16227, N16220, N4953, N12490);
xor XOR2 (N16228, N16215, N7304);
nand NAND4 (N16229, N16225, N801, N4373, N1039);
nor NOR2 (N16230, N16210, N9010);
not NOT1 (N16231, N16213);
nor NOR4 (N16232, N16203, N10751, N279, N4761);
not NOT1 (N16233, N16217);
nand NAND3 (N16234, N16223, N3381, N14960);
not NOT1 (N16235, N16230);
or OR3 (N16236, N16229, N6971, N9807);
and AND4 (N16237, N16226, N9591, N7706, N4402);
or OR4 (N16238, N16231, N15572, N5282, N4155);
and AND3 (N16239, N16232, N706, N492);
nor NOR3 (N16240, N16237, N7445, N12276);
xor XOR2 (N16241, N16234, N206);
or OR2 (N16242, N16219, N15951);
xor XOR2 (N16243, N16227, N8194);
not NOT1 (N16244, N16243);
or OR3 (N16245, N16228, N15340, N13469);
or OR2 (N16246, N16242, N11812);
nand NAND2 (N16247, N16235, N6617);
nor NOR3 (N16248, N16233, N842, N1593);
nor NOR4 (N16249, N16238, N13715, N15022, N2885);
not NOT1 (N16250, N16249);
not NOT1 (N16251, N16244);
xor XOR2 (N16252, N16246, N15233);
buf BUF1 (N16253, N16236);
xor XOR2 (N16254, N16253, N6270);
nor NOR2 (N16255, N16252, N1734);
or OR3 (N16256, N16241, N14265, N7633);
nor NOR3 (N16257, N16245, N9209, N10626);
xor XOR2 (N16258, N16255, N5759);
xor XOR2 (N16259, N16248, N1615);
nand NAND3 (N16260, N16250, N15085, N13794);
buf BUF1 (N16261, N16254);
xor XOR2 (N16262, N16256, N10645);
not NOT1 (N16263, N16259);
buf BUF1 (N16264, N16260);
nand NAND3 (N16265, N16247, N7327, N4505);
not NOT1 (N16266, N16264);
nand NAND4 (N16267, N16239, N1817, N3368, N6240);
nand NAND2 (N16268, N16257, N10137);
buf BUF1 (N16269, N16266);
not NOT1 (N16270, N16258);
and AND2 (N16271, N16263, N3334);
nand NAND2 (N16272, N16251, N13266);
and AND4 (N16273, N16261, N3168, N10042, N14781);
and AND3 (N16274, N16272, N6614, N15638);
buf BUF1 (N16275, N16265);
nor NOR2 (N16276, N16273, N1446);
and AND3 (N16277, N16240, N420, N9062);
or OR2 (N16278, N16270, N4183);
or OR3 (N16279, N16267, N7305, N14213);
xor XOR2 (N16280, N16274, N2724);
or OR3 (N16281, N16262, N4986, N2895);
nor NOR3 (N16282, N16278, N12109, N3928);
not NOT1 (N16283, N16271);
xor XOR2 (N16284, N16268, N6228);
buf BUF1 (N16285, N16284);
nor NOR3 (N16286, N16281, N4572, N13551);
or OR3 (N16287, N16275, N12574, N10590);
not NOT1 (N16288, N16286);
buf BUF1 (N16289, N16277);
or OR4 (N16290, N16285, N7701, N6899, N1159);
not NOT1 (N16291, N16276);
xor XOR2 (N16292, N16290, N8460);
nand NAND3 (N16293, N16279, N5417, N12696);
and AND3 (N16294, N16283, N7220, N626);
nand NAND3 (N16295, N16289, N6633, N12292);
buf BUF1 (N16296, N16295);
not NOT1 (N16297, N16269);
or OR3 (N16298, N16288, N1557, N7376);
nor NOR4 (N16299, N16297, N9961, N12294, N13577);
nand NAND3 (N16300, N16299, N3012, N14019);
xor XOR2 (N16301, N16296, N2261);
and AND2 (N16302, N16292, N10211);
nor NOR4 (N16303, N16282, N14351, N11918, N3688);
nand NAND3 (N16304, N16300, N8394, N11195);
not NOT1 (N16305, N16303);
or OR2 (N16306, N16280, N4618);
nand NAND2 (N16307, N16305, N7508);
buf BUF1 (N16308, N16293);
nor NOR2 (N16309, N16304, N4221);
and AND4 (N16310, N16298, N12118, N6422, N16297);
nor NOR3 (N16311, N16310, N3997, N740);
or OR3 (N16312, N16302, N7816, N1054);
nand NAND3 (N16313, N16291, N4508, N7355);
nand NAND2 (N16314, N16308, N9106);
nor NOR3 (N16315, N16307, N9182, N4635);
or OR2 (N16316, N16313, N606);
or OR2 (N16317, N16316, N16230);
and AND4 (N16318, N16306, N6552, N7001, N4293);
not NOT1 (N16319, N16312);
nand NAND2 (N16320, N16301, N13202);
nand NAND2 (N16321, N16318, N2554);
not NOT1 (N16322, N16314);
not NOT1 (N16323, N16315);
nor NOR3 (N16324, N16319, N10501, N10357);
or OR2 (N16325, N16320, N3093);
not NOT1 (N16326, N16322);
and AND4 (N16327, N16294, N11025, N12129, N6864);
xor XOR2 (N16328, N16326, N12413);
or OR3 (N16329, N16287, N11332, N15670);
nand NAND3 (N16330, N16311, N3801, N12711);
nand NAND3 (N16331, N16323, N1762, N13842);
nor NOR4 (N16332, N16327, N1863, N350, N11031);
buf BUF1 (N16333, N16321);
nor NOR2 (N16334, N16324, N14395);
or OR3 (N16335, N16331, N11099, N866);
or OR2 (N16336, N16317, N16103);
and AND2 (N16337, N16325, N8654);
nand NAND2 (N16338, N16330, N2560);
or OR4 (N16339, N16309, N8140, N9363, N1004);
and AND2 (N16340, N16337, N16152);
xor XOR2 (N16341, N16328, N14291);
not NOT1 (N16342, N16332);
nor NOR4 (N16343, N16338, N15146, N15878, N9406);
and AND4 (N16344, N16343, N14799, N14231, N12602);
nor NOR3 (N16345, N16340, N5453, N1829);
and AND3 (N16346, N16333, N15054, N12443);
nand NAND3 (N16347, N16345, N14728, N12299);
xor XOR2 (N16348, N16344, N7425);
buf BUF1 (N16349, N16348);
xor XOR2 (N16350, N16349, N3041);
xor XOR2 (N16351, N16342, N10742);
nor NOR3 (N16352, N16341, N13337, N14344);
nor NOR4 (N16353, N16346, N15816, N5067, N7793);
xor XOR2 (N16354, N16334, N237);
nor NOR3 (N16355, N16354, N12984, N14401);
nand NAND3 (N16356, N16329, N5644, N7947);
nand NAND3 (N16357, N16335, N6778, N12883);
and AND4 (N16358, N16355, N1027, N9388, N6037);
nand NAND3 (N16359, N16350, N9306, N7885);
nand NAND2 (N16360, N16359, N14219);
buf BUF1 (N16361, N16357);
or OR3 (N16362, N16358, N12169, N15900);
buf BUF1 (N16363, N16360);
xor XOR2 (N16364, N16361, N9888);
nand NAND4 (N16365, N16363, N7845, N11463, N12788);
or OR2 (N16366, N16351, N5717);
or OR4 (N16367, N16364, N15268, N11870, N10542);
nor NOR4 (N16368, N16336, N10956, N12069, N9752);
nand NAND2 (N16369, N16368, N2724);
buf BUF1 (N16370, N16356);
or OR3 (N16371, N16365, N14120, N6286);
nor NOR2 (N16372, N16362, N8418);
nand NAND4 (N16373, N16353, N3510, N7507, N8638);
xor XOR2 (N16374, N16371, N14769);
and AND2 (N16375, N16352, N14035);
xor XOR2 (N16376, N16374, N14468);
nor NOR3 (N16377, N16367, N6713, N16097);
or OR2 (N16378, N16377, N11413);
xor XOR2 (N16379, N16372, N2507);
not NOT1 (N16380, N16339);
nand NAND3 (N16381, N16376, N4205, N10088);
nand NAND3 (N16382, N16375, N9546, N10085);
nand NAND3 (N16383, N16380, N15517, N14892);
not NOT1 (N16384, N16347);
xor XOR2 (N16385, N16369, N15257);
nand NAND3 (N16386, N16379, N3622, N2025);
buf BUF1 (N16387, N16382);
and AND2 (N16388, N16373, N13906);
not NOT1 (N16389, N16383);
not NOT1 (N16390, N16378);
not NOT1 (N16391, N16370);
not NOT1 (N16392, N16386);
buf BUF1 (N16393, N16391);
and AND4 (N16394, N16392, N11278, N2572, N10405);
or OR2 (N16395, N16393, N50);
nand NAND2 (N16396, N16381, N327);
or OR2 (N16397, N16387, N8363);
buf BUF1 (N16398, N16384);
xor XOR2 (N16399, N16366, N5968);
buf BUF1 (N16400, N16397);
nand NAND3 (N16401, N16388, N7305, N11680);
xor XOR2 (N16402, N16398, N8751);
and AND4 (N16403, N16394, N7525, N15684, N8609);
buf BUF1 (N16404, N16403);
nor NOR3 (N16405, N16389, N10603, N11949);
nor NOR4 (N16406, N16404, N1291, N3788, N4333);
nor NOR3 (N16407, N16400, N16171, N14733);
nor NOR2 (N16408, N16401, N8603);
not NOT1 (N16409, N16408);
or OR4 (N16410, N16406, N13401, N2450, N6334);
and AND3 (N16411, N16409, N13790, N8448);
buf BUF1 (N16412, N16395);
nand NAND4 (N16413, N16410, N113, N4235, N12085);
nor NOR3 (N16414, N16412, N8405, N10730);
buf BUF1 (N16415, N16411);
nor NOR3 (N16416, N16402, N5067, N16175);
nor NOR2 (N16417, N16407, N10371);
not NOT1 (N16418, N16415);
xor XOR2 (N16419, N16417, N13478);
nand NAND4 (N16420, N16413, N11104, N10215, N2192);
and AND2 (N16421, N16418, N3493);
nor NOR3 (N16422, N16416, N11841, N4406);
not NOT1 (N16423, N16420);
buf BUF1 (N16424, N16422);
buf BUF1 (N16425, N16405);
buf BUF1 (N16426, N16425);
or OR2 (N16427, N16385, N13712);
or OR3 (N16428, N16426, N489, N9427);
xor XOR2 (N16429, N16428, N4793);
not NOT1 (N16430, N16423);
nand NAND4 (N16431, N16427, N2947, N11697, N10820);
nor NOR2 (N16432, N16390, N10764);
nor NOR4 (N16433, N16419, N14613, N5840, N15884);
nand NAND2 (N16434, N16433, N14082);
xor XOR2 (N16435, N16430, N6421);
nor NOR3 (N16436, N16399, N16174, N14478);
xor XOR2 (N16437, N16414, N10219);
not NOT1 (N16438, N16434);
or OR2 (N16439, N16436, N7163);
nor NOR3 (N16440, N16421, N12540, N12125);
not NOT1 (N16441, N16424);
not NOT1 (N16442, N16437);
and AND3 (N16443, N16429, N4264, N892);
xor XOR2 (N16444, N16432, N4175);
or OR2 (N16445, N16440, N6936);
nand NAND4 (N16446, N16445, N10199, N4781, N8430);
and AND3 (N16447, N16439, N7831, N9321);
or OR4 (N16448, N16441, N11567, N15389, N11051);
and AND2 (N16449, N16444, N899);
xor XOR2 (N16450, N16431, N3074);
not NOT1 (N16451, N16450);
buf BUF1 (N16452, N16442);
xor XOR2 (N16453, N16435, N8488);
not NOT1 (N16454, N16443);
and AND3 (N16455, N16449, N2576, N11152);
not NOT1 (N16456, N16438);
or OR4 (N16457, N16452, N1607, N8962, N5572);
nand NAND3 (N16458, N16396, N6047, N6919);
or OR3 (N16459, N16458, N340, N5024);
buf BUF1 (N16460, N16457);
nor NOR2 (N16461, N16455, N15334);
nand NAND2 (N16462, N16461, N7030);
buf BUF1 (N16463, N16460);
not NOT1 (N16464, N16446);
nor NOR2 (N16465, N16447, N2696);
and AND2 (N16466, N16463, N7757);
buf BUF1 (N16467, N16465);
or OR3 (N16468, N16453, N14192, N9591);
xor XOR2 (N16469, N16456, N1788);
buf BUF1 (N16470, N16466);
nor NOR4 (N16471, N16469, N13089, N15842, N14627);
or OR4 (N16472, N16470, N545, N11838, N8870);
xor XOR2 (N16473, N16468, N1599);
and AND3 (N16474, N16454, N4723, N3360);
or OR3 (N16475, N16472, N5136, N11734);
buf BUF1 (N16476, N16464);
nand NAND2 (N16477, N16475, N7793);
buf BUF1 (N16478, N16476);
and AND3 (N16479, N16467, N15907, N12469);
and AND3 (N16480, N16471, N8442, N1056);
xor XOR2 (N16481, N16451, N8503);
nand NAND2 (N16482, N16474, N13904);
or OR4 (N16483, N16480, N6052, N4405, N13183);
nor NOR3 (N16484, N16459, N13146, N12765);
nand NAND2 (N16485, N16462, N9628);
nand NAND2 (N16486, N16478, N9914);
xor XOR2 (N16487, N16484, N6939);
not NOT1 (N16488, N16481);
buf BUF1 (N16489, N16482);
not NOT1 (N16490, N16488);
or OR3 (N16491, N16486, N2471, N9036);
nor NOR2 (N16492, N16473, N2709);
xor XOR2 (N16493, N16492, N12195);
nand NAND3 (N16494, N16489, N2363, N12925);
xor XOR2 (N16495, N16483, N7075);
nor NOR2 (N16496, N16487, N6644);
and AND2 (N16497, N16496, N4466);
or OR3 (N16498, N16477, N14224, N1762);
buf BUF1 (N16499, N16494);
buf BUF1 (N16500, N16490);
nor NOR2 (N16501, N16493, N14534);
buf BUF1 (N16502, N16501);
and AND4 (N16503, N16502, N13033, N9347, N1541);
not NOT1 (N16504, N16497);
not NOT1 (N16505, N16479);
buf BUF1 (N16506, N16498);
buf BUF1 (N16507, N16491);
nor NOR2 (N16508, N16504, N5482);
nor NOR2 (N16509, N16499, N7480);
or OR3 (N16510, N16506, N5750, N7685);
and AND2 (N16511, N16507, N12567);
nand NAND4 (N16512, N16508, N2590, N9285, N6002);
nor NOR3 (N16513, N16512, N14646, N14018);
or OR3 (N16514, N16513, N7778, N10421);
or OR3 (N16515, N16495, N5593, N7952);
and AND4 (N16516, N16514, N11413, N16371, N10539);
nor NOR2 (N16517, N16503, N10931);
nor NOR3 (N16518, N16511, N13469, N5845);
buf BUF1 (N16519, N16448);
nand NAND4 (N16520, N16510, N5291, N3620, N12393);
not NOT1 (N16521, N16515);
nor NOR3 (N16522, N16505, N2199, N13637);
or OR4 (N16523, N16522, N9565, N13802, N4780);
not NOT1 (N16524, N16518);
not NOT1 (N16525, N16517);
nand NAND4 (N16526, N16509, N2875, N10519, N5786);
buf BUF1 (N16527, N16519);
xor XOR2 (N16528, N16521, N7911);
nor NOR2 (N16529, N16524, N2573);
and AND3 (N16530, N16500, N6762, N6024);
xor XOR2 (N16531, N16529, N4742);
buf BUF1 (N16532, N16526);
nand NAND2 (N16533, N16527, N8193);
nor NOR4 (N16534, N16533, N9773, N10611, N6468);
buf BUF1 (N16535, N16530);
nand NAND2 (N16536, N16516, N6466);
nor NOR2 (N16537, N16536, N1732);
nor NOR2 (N16538, N16531, N13416);
nor NOR3 (N16539, N16532, N2560, N10802);
nand NAND4 (N16540, N16538, N12758, N12568, N2322);
nand NAND4 (N16541, N16520, N14775, N2871, N4348);
nor NOR3 (N16542, N16541, N6445, N962);
nand NAND3 (N16543, N16539, N772, N4798);
buf BUF1 (N16544, N16537);
nand NAND3 (N16545, N16528, N10175, N16246);
buf BUF1 (N16546, N16540);
not NOT1 (N16547, N16525);
xor XOR2 (N16548, N16545, N5241);
not NOT1 (N16549, N16547);
xor XOR2 (N16550, N16549, N8936);
or OR3 (N16551, N16548, N15256, N7003);
and AND3 (N16552, N16542, N9292, N6020);
xor XOR2 (N16553, N16535, N5382);
and AND3 (N16554, N16543, N209, N9665);
not NOT1 (N16555, N16523);
not NOT1 (N16556, N16553);
xor XOR2 (N16557, N16556, N15193);
and AND4 (N16558, N16552, N3521, N4503, N2164);
and AND2 (N16559, N16558, N9349);
xor XOR2 (N16560, N16551, N12491);
and AND2 (N16561, N16560, N6415);
buf BUF1 (N16562, N16544);
and AND2 (N16563, N16485, N2754);
not NOT1 (N16564, N16555);
not NOT1 (N16565, N16564);
xor XOR2 (N16566, N16563, N12192);
xor XOR2 (N16567, N16550, N5453);
xor XOR2 (N16568, N16567, N14923);
xor XOR2 (N16569, N16559, N6035);
xor XOR2 (N16570, N16557, N9458);
or OR3 (N16571, N16569, N9418, N12685);
xor XOR2 (N16572, N16554, N6421);
nor NOR4 (N16573, N16561, N6440, N8942, N3053);
nand NAND4 (N16574, N16565, N6328, N5573, N14391);
nand NAND2 (N16575, N16570, N6051);
and AND2 (N16576, N16575, N7835);
not NOT1 (N16577, N16571);
and AND4 (N16578, N16562, N13707, N12318, N5853);
or OR4 (N16579, N16573, N13171, N2594, N1083);
and AND4 (N16580, N16579, N4414, N433, N4775);
nand NAND2 (N16581, N16574, N1800);
nor NOR2 (N16582, N16566, N10208);
and AND4 (N16583, N16572, N4769, N4732, N8505);
buf BUF1 (N16584, N16577);
nand NAND4 (N16585, N16576, N16482, N15237, N10195);
xor XOR2 (N16586, N16580, N2228);
buf BUF1 (N16587, N16582);
nor NOR2 (N16588, N16587, N10023);
xor XOR2 (N16589, N16568, N739);
not NOT1 (N16590, N16586);
nor NOR3 (N16591, N16578, N5158, N4690);
xor XOR2 (N16592, N16546, N11134);
nor NOR2 (N16593, N16588, N8031);
or OR3 (N16594, N16591, N3900, N10406);
or OR2 (N16595, N16593, N6131);
or OR4 (N16596, N16581, N11720, N11510, N5781);
buf BUF1 (N16597, N16595);
buf BUF1 (N16598, N16590);
nor NOR2 (N16599, N16584, N9309);
xor XOR2 (N16600, N16589, N3386);
buf BUF1 (N16601, N16594);
and AND2 (N16602, N16601, N16332);
and AND3 (N16603, N16534, N11285, N1923);
buf BUF1 (N16604, N16583);
not NOT1 (N16605, N16603);
nor NOR3 (N16606, N16599, N10137, N8383);
buf BUF1 (N16607, N16606);
or OR2 (N16608, N16605, N1934);
not NOT1 (N16609, N16592);
and AND2 (N16610, N16597, N7072);
nand NAND4 (N16611, N16610, N11842, N2346, N12991);
not NOT1 (N16612, N16609);
xor XOR2 (N16613, N16612, N11392);
and AND2 (N16614, N16598, N7364);
not NOT1 (N16615, N16600);
or OR4 (N16616, N16607, N1179, N523, N7208);
nor NOR3 (N16617, N16604, N11056, N2827);
buf BUF1 (N16618, N16614);
not NOT1 (N16619, N16602);
xor XOR2 (N16620, N16608, N13310);
not NOT1 (N16621, N16617);
and AND3 (N16622, N16585, N1565, N6015);
buf BUF1 (N16623, N16620);
nand NAND3 (N16624, N16613, N10062, N6968);
not NOT1 (N16625, N16618);
nand NAND2 (N16626, N16611, N11727);
or OR2 (N16627, N16596, N11487);
buf BUF1 (N16628, N16622);
buf BUF1 (N16629, N16619);
xor XOR2 (N16630, N16626, N13026);
and AND3 (N16631, N16630, N3312, N12255);
or OR3 (N16632, N16627, N14337, N367);
not NOT1 (N16633, N16616);
buf BUF1 (N16634, N16632);
or OR4 (N16635, N16629, N2698, N8406, N5959);
buf BUF1 (N16636, N16623);
buf BUF1 (N16637, N16635);
nand NAND3 (N16638, N16633, N7317, N3391);
not NOT1 (N16639, N16637);
nand NAND2 (N16640, N16628, N7704);
not NOT1 (N16641, N16639);
xor XOR2 (N16642, N16615, N5059);
nand NAND4 (N16643, N16624, N7751, N5297, N6622);
or OR4 (N16644, N16640, N8617, N2022, N7136);
nor NOR2 (N16645, N16621, N14254);
or OR3 (N16646, N16631, N6684, N781);
nand NAND4 (N16647, N16643, N13401, N10852, N11600);
buf BUF1 (N16648, N16647);
not NOT1 (N16649, N16634);
or OR3 (N16650, N16649, N12937, N3520);
nand NAND4 (N16651, N16625, N5468, N9078, N979);
xor XOR2 (N16652, N16651, N4630);
nor NOR3 (N16653, N16646, N12433, N2718);
not NOT1 (N16654, N16645);
not NOT1 (N16655, N16654);
buf BUF1 (N16656, N16644);
or OR2 (N16657, N16641, N7613);
buf BUF1 (N16658, N16642);
nor NOR3 (N16659, N16638, N3798, N302);
not NOT1 (N16660, N16656);
xor XOR2 (N16661, N16650, N4896);
and AND4 (N16662, N16636, N10278, N688, N804);
nand NAND2 (N16663, N16658, N16410);
nand NAND3 (N16664, N16660, N2914, N7361);
xor XOR2 (N16665, N16657, N2588);
not NOT1 (N16666, N16652);
nand NAND2 (N16667, N16664, N9146);
xor XOR2 (N16668, N16655, N9237);
nand NAND2 (N16669, N16661, N11821);
xor XOR2 (N16670, N16648, N14904);
buf BUF1 (N16671, N16662);
and AND2 (N16672, N16671, N9245);
or OR2 (N16673, N16669, N7824);
buf BUF1 (N16674, N16673);
buf BUF1 (N16675, N16659);
xor XOR2 (N16676, N16668, N12482);
nand NAND2 (N16677, N16670, N2421);
buf BUF1 (N16678, N16677);
or OR2 (N16679, N16653, N5668);
xor XOR2 (N16680, N16665, N9058);
not NOT1 (N16681, N16679);
nor NOR2 (N16682, N16672, N7591);
nand NAND3 (N16683, N16676, N15037, N3725);
xor XOR2 (N16684, N16682, N14093);
xor XOR2 (N16685, N16666, N16112);
xor XOR2 (N16686, N16681, N5800);
buf BUF1 (N16687, N16663);
xor XOR2 (N16688, N16685, N14520);
nor NOR3 (N16689, N16683, N1103, N10192);
not NOT1 (N16690, N16675);
and AND2 (N16691, N16690, N2466);
nor NOR2 (N16692, N16667, N2171);
xor XOR2 (N16693, N16687, N15774);
xor XOR2 (N16694, N16691, N8629);
nor NOR3 (N16695, N16688, N16617, N7241);
nand NAND4 (N16696, N16694, N16131, N13386, N1128);
buf BUF1 (N16697, N16696);
and AND3 (N16698, N16680, N11334, N803);
xor XOR2 (N16699, N16674, N686);
and AND3 (N16700, N16699, N2568, N8250);
or OR3 (N16701, N16686, N1052, N15508);
not NOT1 (N16702, N16693);
not NOT1 (N16703, N16697);
not NOT1 (N16704, N16678);
xor XOR2 (N16705, N16692, N8992);
or OR4 (N16706, N16689, N730, N13189, N7422);
buf BUF1 (N16707, N16706);
or OR2 (N16708, N16698, N179);
not NOT1 (N16709, N16702);
and AND2 (N16710, N16709, N5631);
or OR4 (N16711, N16707, N6632, N10036, N16416);
not NOT1 (N16712, N16703);
xor XOR2 (N16713, N16701, N4954);
nor NOR4 (N16714, N16708, N7083, N3185, N16650);
and AND2 (N16715, N16704, N13668);
or OR2 (N16716, N16700, N6060);
nor NOR3 (N16717, N16705, N14778, N7894);
buf BUF1 (N16718, N16710);
xor XOR2 (N16719, N16718, N11894);
nand NAND4 (N16720, N16695, N10607, N14749, N14659);
or OR4 (N16721, N16714, N6126, N5915, N12294);
or OR2 (N16722, N16717, N5080);
buf BUF1 (N16723, N16719);
nand NAND2 (N16724, N16711, N7197);
nand NAND2 (N16725, N16716, N6504);
buf BUF1 (N16726, N16721);
nand NAND3 (N16727, N16720, N13289, N2699);
nor NOR2 (N16728, N16713, N3797);
xor XOR2 (N16729, N16722, N2303);
nand NAND2 (N16730, N16725, N3142);
nor NOR3 (N16731, N16684, N16233, N4617);
or OR2 (N16732, N16724, N15472);
nor NOR4 (N16733, N16730, N4809, N12021, N8679);
buf BUF1 (N16734, N16733);
buf BUF1 (N16735, N16734);
xor XOR2 (N16736, N16728, N13461);
nor NOR4 (N16737, N16729, N2205, N16239, N3271);
not NOT1 (N16738, N16735);
nand NAND3 (N16739, N16712, N778, N12470);
not NOT1 (N16740, N16726);
nor NOR2 (N16741, N16737, N6244);
or OR4 (N16742, N16727, N8696, N9891, N12413);
buf BUF1 (N16743, N16738);
and AND3 (N16744, N16731, N2599, N12091);
nor NOR3 (N16745, N16740, N6551, N1667);
or OR3 (N16746, N16715, N1349, N14632);
not NOT1 (N16747, N16745);
xor XOR2 (N16748, N16743, N5898);
nand NAND3 (N16749, N16744, N13674, N15375);
buf BUF1 (N16750, N16736);
nand NAND4 (N16751, N16742, N15123, N5194, N4499);
nor NOR4 (N16752, N16732, N11803, N15978, N7785);
nor NOR4 (N16753, N16750, N1589, N1898, N8723);
buf BUF1 (N16754, N16753);
nand NAND2 (N16755, N16748, N12488);
nand NAND3 (N16756, N16754, N2587, N16754);
buf BUF1 (N16757, N16755);
buf BUF1 (N16758, N16756);
not NOT1 (N16759, N16758);
buf BUF1 (N16760, N16746);
and AND3 (N16761, N16723, N13223, N11005);
buf BUF1 (N16762, N16739);
and AND3 (N16763, N16757, N7770, N67);
or OR2 (N16764, N16761, N1860);
xor XOR2 (N16765, N16752, N2129);
buf BUF1 (N16766, N16749);
and AND3 (N16767, N16765, N13685, N7072);
not NOT1 (N16768, N16747);
and AND3 (N16769, N16767, N3632, N3953);
not NOT1 (N16770, N16759);
or OR3 (N16771, N16751, N9702, N13809);
nor NOR2 (N16772, N16770, N10906);
not NOT1 (N16773, N16763);
buf BUF1 (N16774, N16760);
nand NAND4 (N16775, N16766, N4601, N16198, N7075);
nand NAND3 (N16776, N16774, N13261, N7312);
buf BUF1 (N16777, N16773);
xor XOR2 (N16778, N16772, N219);
or OR4 (N16779, N16771, N15995, N12463, N9745);
or OR3 (N16780, N16778, N12640, N8647);
buf BUF1 (N16781, N16764);
nand NAND3 (N16782, N16775, N15844, N8931);
nand NAND3 (N16783, N16741, N11316, N12963);
or OR3 (N16784, N16777, N5159, N16262);
buf BUF1 (N16785, N16769);
not NOT1 (N16786, N16783);
nand NAND4 (N16787, N16782, N549, N14163, N14620);
nor NOR3 (N16788, N16779, N7348, N2567);
and AND4 (N16789, N16787, N11529, N2873, N11219);
xor XOR2 (N16790, N16785, N9372);
nor NOR2 (N16791, N16780, N4649);
nand NAND3 (N16792, N16762, N2688, N9894);
nor NOR4 (N16793, N16791, N9686, N5748, N3663);
xor XOR2 (N16794, N16781, N16049);
nor NOR4 (N16795, N16768, N16159, N7697, N7236);
nor NOR3 (N16796, N16784, N3234, N1483);
nand NAND2 (N16797, N16786, N993);
nand NAND3 (N16798, N16789, N16087, N6671);
or OR2 (N16799, N16776, N4517);
and AND3 (N16800, N16794, N5199, N5242);
or OR2 (N16801, N16790, N5570);
and AND3 (N16802, N16798, N3119, N15409);
and AND3 (N16803, N16799, N7200, N15482);
buf BUF1 (N16804, N16801);
xor XOR2 (N16805, N16803, N2819);
nor NOR3 (N16806, N16788, N8546, N801);
or OR3 (N16807, N16793, N11130, N1576);
nand NAND3 (N16808, N16807, N3008, N9426);
buf BUF1 (N16809, N16795);
xor XOR2 (N16810, N16792, N1999);
not NOT1 (N16811, N16808);
xor XOR2 (N16812, N16809, N11803);
buf BUF1 (N16813, N16797);
xor XOR2 (N16814, N16806, N16536);
and AND2 (N16815, N16805, N2445);
not NOT1 (N16816, N16811);
and AND4 (N16817, N16800, N10860, N5659, N15639);
and AND4 (N16818, N16804, N9851, N13362, N10288);
not NOT1 (N16819, N16796);
and AND4 (N16820, N16819, N5989, N6894, N12088);
nand NAND4 (N16821, N16814, N11841, N3274, N8425);
nor NOR4 (N16822, N16812, N14005, N5074, N14396);
buf BUF1 (N16823, N16821);
nor NOR3 (N16824, N16820, N2805, N14242);
and AND3 (N16825, N16817, N15484, N12588);
nor NOR2 (N16826, N16825, N8431);
nor NOR2 (N16827, N16810, N9485);
buf BUF1 (N16828, N16802);
buf BUF1 (N16829, N16822);
nand NAND4 (N16830, N16827, N14316, N12849, N13167);
not NOT1 (N16831, N16815);
nand NAND2 (N16832, N16824, N6999);
nand NAND3 (N16833, N16832, N11958, N4933);
buf BUF1 (N16834, N16813);
buf BUF1 (N16835, N16826);
xor XOR2 (N16836, N16831, N11143);
not NOT1 (N16837, N16835);
or OR3 (N16838, N16823, N13378, N3585);
and AND4 (N16839, N16834, N5162, N3128, N14726);
nand NAND2 (N16840, N16828, N648);
and AND2 (N16841, N16818, N9506);
buf BUF1 (N16842, N16838);
or OR4 (N16843, N16842, N3196, N14686, N441);
not NOT1 (N16844, N16830);
nand NAND3 (N16845, N16844, N9652, N15969);
nand NAND4 (N16846, N16840, N10470, N16148, N9727);
not NOT1 (N16847, N16837);
xor XOR2 (N16848, N16845, N9557);
xor XOR2 (N16849, N16816, N3737);
nor NOR2 (N16850, N16833, N11304);
or OR2 (N16851, N16829, N7338);
nand NAND4 (N16852, N16847, N14452, N1483, N6537);
or OR3 (N16853, N16851, N4474, N2833);
nand NAND2 (N16854, N16836, N13860);
and AND2 (N16855, N16841, N4106);
buf BUF1 (N16856, N16853);
xor XOR2 (N16857, N16839, N7965);
buf BUF1 (N16858, N16848);
nand NAND3 (N16859, N16856, N6760, N4865);
xor XOR2 (N16860, N16855, N6593);
not NOT1 (N16861, N16858);
buf BUF1 (N16862, N16849);
and AND2 (N16863, N16854, N500);
or OR2 (N16864, N16846, N9978);
xor XOR2 (N16865, N16864, N5495);
and AND3 (N16866, N16857, N1813, N2641);
and AND2 (N16867, N16863, N14875);
buf BUF1 (N16868, N16867);
and AND4 (N16869, N16861, N11744, N9423, N15271);
not NOT1 (N16870, N16852);
nor NOR2 (N16871, N16859, N1597);
xor XOR2 (N16872, N16871, N483);
not NOT1 (N16873, N16843);
and AND4 (N16874, N16860, N6614, N2523, N11195);
and AND4 (N16875, N16873, N4696, N9131, N7780);
and AND2 (N16876, N16862, N14);
or OR3 (N16877, N16865, N14780, N2351);
nor NOR2 (N16878, N16866, N14937);
not NOT1 (N16879, N16850);
and AND4 (N16880, N16878, N15275, N2514, N11669);
nor NOR3 (N16881, N16879, N10430, N2535);
buf BUF1 (N16882, N16880);
not NOT1 (N16883, N16876);
not NOT1 (N16884, N16875);
xor XOR2 (N16885, N16881, N12397);
xor XOR2 (N16886, N16869, N6669);
buf BUF1 (N16887, N16870);
xor XOR2 (N16888, N16877, N16721);
and AND4 (N16889, N16884, N16040, N14915, N11714);
nand NAND2 (N16890, N16874, N4304);
xor XOR2 (N16891, N16890, N14667);
and AND2 (N16892, N16868, N5554);
not NOT1 (N16893, N16892);
xor XOR2 (N16894, N16885, N133);
and AND4 (N16895, N16882, N11016, N11646, N16163);
not NOT1 (N16896, N16888);
or OR2 (N16897, N16886, N7867);
xor XOR2 (N16898, N16896, N1333);
or OR4 (N16899, N16895, N9927, N16650, N11564);
nor NOR4 (N16900, N16883, N8817, N16105, N2814);
buf BUF1 (N16901, N16899);
and AND3 (N16902, N16887, N10253, N6763);
buf BUF1 (N16903, N16872);
buf BUF1 (N16904, N16900);
or OR2 (N16905, N16891, N16309);
or OR4 (N16906, N16894, N4100, N14485, N4371);
and AND2 (N16907, N16901, N16750);
xor XOR2 (N16908, N16897, N7725);
nor NOR3 (N16909, N16902, N15745, N7215);
nor NOR3 (N16910, N16893, N4608, N12015);
not NOT1 (N16911, N16909);
nor NOR2 (N16912, N16907, N4371);
buf BUF1 (N16913, N16908);
or OR4 (N16914, N16889, N10820, N2589, N4587);
and AND2 (N16915, N16905, N16558);
nor NOR3 (N16916, N16903, N12545, N15109);
and AND3 (N16917, N16916, N1219, N15960);
or OR2 (N16918, N16914, N9299);
xor XOR2 (N16919, N16915, N11246);
buf BUF1 (N16920, N16919);
nor NOR2 (N16921, N16898, N10900);
nand NAND2 (N16922, N16920, N9580);
and AND3 (N16923, N16913, N5436, N2471);
nand NAND3 (N16924, N16922, N7586, N12336);
and AND4 (N16925, N16904, N11233, N16010, N11413);
not NOT1 (N16926, N16918);
nor NOR4 (N16927, N16921, N10076, N5009, N4172);
nor NOR2 (N16928, N16923, N10108);
xor XOR2 (N16929, N16911, N2917);
not NOT1 (N16930, N16906);
nand NAND2 (N16931, N16927, N3391);
and AND4 (N16932, N16926, N13947, N4718, N1601);
nor NOR3 (N16933, N16929, N9912, N11066);
or OR2 (N16934, N16931, N5022);
not NOT1 (N16935, N16933);
or OR3 (N16936, N16928, N8516, N3898);
xor XOR2 (N16937, N16910, N4274);
buf BUF1 (N16938, N16936);
nor NOR4 (N16939, N16925, N10042, N4928, N12069);
xor XOR2 (N16940, N16935, N15316);
not NOT1 (N16941, N16912);
buf BUF1 (N16942, N16930);
buf BUF1 (N16943, N16924);
or OR3 (N16944, N16932, N3314, N3891);
and AND2 (N16945, N16944, N6042);
not NOT1 (N16946, N16942);
xor XOR2 (N16947, N16946, N11636);
buf BUF1 (N16948, N16934);
and AND2 (N16949, N16943, N6275);
and AND2 (N16950, N16917, N4871);
buf BUF1 (N16951, N16939);
or OR4 (N16952, N16948, N10879, N13602, N7199);
and AND3 (N16953, N16938, N9608, N15085);
nor NOR3 (N16954, N16949, N9253, N6947);
nand NAND2 (N16955, N16954, N4803);
and AND2 (N16956, N16940, N10492);
nor NOR4 (N16957, N16941, N4328, N5879, N6625);
or OR4 (N16958, N16945, N8735, N11840, N3145);
nor NOR2 (N16959, N16958, N13460);
or OR3 (N16960, N16959, N7040, N12475);
nor NOR3 (N16961, N16951, N15357, N2560);
xor XOR2 (N16962, N16950, N15279);
xor XOR2 (N16963, N16937, N14135);
buf BUF1 (N16964, N16960);
and AND4 (N16965, N16953, N5463, N6573, N1011);
nand NAND2 (N16966, N16957, N13800);
nor NOR4 (N16967, N16966, N1917, N6262, N14720);
nor NOR3 (N16968, N16947, N14321, N9650);
buf BUF1 (N16969, N16964);
nor NOR2 (N16970, N16965, N14573);
nand NAND4 (N16971, N16967, N12753, N13594, N13767);
nand NAND4 (N16972, N16961, N7433, N7080, N14672);
nand NAND3 (N16973, N16955, N10081, N191);
buf BUF1 (N16974, N16971);
buf BUF1 (N16975, N16970);
nand NAND3 (N16976, N16969, N8364, N15258);
xor XOR2 (N16977, N16974, N6604);
and AND4 (N16978, N16976, N2702, N8333, N2449);
or OR3 (N16979, N16977, N10298, N1314);
nand NAND2 (N16980, N16973, N8145);
and AND2 (N16981, N16972, N4790);
or OR4 (N16982, N16956, N2425, N252, N3346);
not NOT1 (N16983, N16982);
nor NOR4 (N16984, N16963, N14055, N6349, N12001);
buf BUF1 (N16985, N16978);
xor XOR2 (N16986, N16975, N13544);
nor NOR4 (N16987, N16952, N7282, N4865, N8815);
nor NOR2 (N16988, N16962, N10522);
nand NAND4 (N16989, N16979, N6282, N515, N15908);
buf BUF1 (N16990, N16986);
nand NAND3 (N16991, N16985, N11638, N16054);
not NOT1 (N16992, N16991);
nor NOR3 (N16993, N16988, N15360, N1925);
nand NAND2 (N16994, N16993, N12056);
nor NOR4 (N16995, N16981, N7769, N5233, N14834);
nor NOR2 (N16996, N16984, N16991);
or OR3 (N16997, N16989, N8124, N6286);
nand NAND2 (N16998, N16980, N15079);
buf BUF1 (N16999, N16998);
or OR4 (N17000, N16997, N4431, N4445, N1813);
nand NAND4 (N17001, N16995, N5319, N12931, N9531);
xor XOR2 (N17002, N17001, N3001);
xor XOR2 (N17003, N16994, N7498);
nor NOR4 (N17004, N16992, N14948, N2266, N7);
nor NOR3 (N17005, N16990, N2663, N5512);
nor NOR3 (N17006, N17003, N6669, N5213);
not NOT1 (N17007, N17006);
nor NOR4 (N17008, N16968, N2163, N11169, N6520);
nand NAND4 (N17009, N17005, N6888, N15424, N16811);
xor XOR2 (N17010, N16996, N10041);
or OR2 (N17011, N16983, N3154);
nand NAND2 (N17012, N16987, N8469);
nand NAND4 (N17013, N17010, N514, N4140, N1096);
xor XOR2 (N17014, N17009, N11024);
xor XOR2 (N17015, N17011, N9467);
buf BUF1 (N17016, N17008);
xor XOR2 (N17017, N17004, N16648);
or OR4 (N17018, N17007, N8906, N1947, N8501);
nand NAND2 (N17019, N17000, N5596);
buf BUF1 (N17020, N17015);
buf BUF1 (N17021, N16999);
xor XOR2 (N17022, N17019, N15913);
buf BUF1 (N17023, N17014);
or OR3 (N17024, N17018, N15846, N13530);
xor XOR2 (N17025, N17020, N12481);
nor NOR3 (N17026, N17024, N418, N12472);
nor NOR2 (N17027, N17022, N12872);
buf BUF1 (N17028, N17021);
buf BUF1 (N17029, N17025);
xor XOR2 (N17030, N17002, N10660);
xor XOR2 (N17031, N17026, N2639);
nand NAND4 (N17032, N17017, N15822, N8199, N2728);
or OR3 (N17033, N17013, N9633, N16377);
buf BUF1 (N17034, N17030);
not NOT1 (N17035, N17012);
xor XOR2 (N17036, N17034, N3289);
nand NAND4 (N17037, N17027, N4433, N13813, N10247);
and AND4 (N17038, N17016, N8283, N470, N12293);
not NOT1 (N17039, N17028);
buf BUF1 (N17040, N17029);
xor XOR2 (N17041, N17039, N10796);
nand NAND3 (N17042, N17037, N7757, N11113);
nand NAND2 (N17043, N17023, N16004);
or OR3 (N17044, N17036, N12203, N13496);
nand NAND2 (N17045, N17033, N6888);
xor XOR2 (N17046, N17040, N12914);
and AND4 (N17047, N17046, N4319, N16047, N16504);
buf BUF1 (N17048, N17041);
and AND3 (N17049, N17042, N419, N8130);
nor NOR3 (N17050, N17035, N14693, N11025);
nor NOR4 (N17051, N17045, N3328, N893, N16803);
and AND3 (N17052, N17047, N13589, N7849);
xor XOR2 (N17053, N17049, N6226);
and AND2 (N17054, N17031, N5688);
nor NOR3 (N17055, N17050, N7514, N16555);
and AND3 (N17056, N17048, N9564, N11180);
and AND4 (N17057, N17043, N6959, N1891, N3207);
nand NAND2 (N17058, N17052, N15104);
buf BUF1 (N17059, N17058);
buf BUF1 (N17060, N17032);
not NOT1 (N17061, N17038);
nand NAND4 (N17062, N17053, N5572, N2974, N3775);
nand NAND4 (N17063, N17062, N12096, N4376, N4804);
or OR4 (N17064, N17054, N921, N3691, N11163);
or OR2 (N17065, N17063, N13227);
or OR4 (N17066, N17060, N4158, N5961, N12237);
nand NAND3 (N17067, N17064, N15356, N12977);
xor XOR2 (N17068, N17057, N12723);
and AND2 (N17069, N17067, N7802);
nor NOR3 (N17070, N17051, N15886, N16241);
not NOT1 (N17071, N17066);
nand NAND2 (N17072, N17061, N13510);
not NOT1 (N17073, N17065);
or OR4 (N17074, N17056, N1833, N8405, N12272);
buf BUF1 (N17075, N17068);
xor XOR2 (N17076, N17069, N6167);
or OR2 (N17077, N17075, N11141);
buf BUF1 (N17078, N17076);
xor XOR2 (N17079, N17059, N8559);
buf BUF1 (N17080, N17074);
xor XOR2 (N17081, N17044, N7067);
xor XOR2 (N17082, N17079, N6722);
not NOT1 (N17083, N17072);
buf BUF1 (N17084, N17077);
nor NOR4 (N17085, N17084, N2061, N5287, N9326);
nand NAND3 (N17086, N17071, N6512, N880);
or OR3 (N17087, N17070, N3855, N5847);
and AND3 (N17088, N17086, N16290, N15554);
and AND4 (N17089, N17083, N8214, N108, N9868);
or OR4 (N17090, N17082, N13733, N9245, N9270);
nand NAND4 (N17091, N17089, N15231, N319, N889);
and AND2 (N17092, N17087, N16692);
nand NAND4 (N17093, N17085, N5606, N7593, N16597);
nor NOR4 (N17094, N17093, N12811, N66, N16128);
xor XOR2 (N17095, N17088, N14569);
nor NOR3 (N17096, N17090, N8690, N9963);
buf BUF1 (N17097, N17091);
nand NAND2 (N17098, N17078, N5788);
or OR4 (N17099, N17081, N17015, N2517, N15329);
xor XOR2 (N17100, N17073, N6190);
or OR4 (N17101, N17099, N8930, N9726, N4546);
nand NAND2 (N17102, N17092, N4882);
xor XOR2 (N17103, N17100, N10705);
and AND3 (N17104, N17097, N6150, N13189);
xor XOR2 (N17105, N17103, N16523);
nor NOR4 (N17106, N17094, N3050, N16363, N14443);
xor XOR2 (N17107, N17104, N15910);
nor NOR3 (N17108, N17096, N9080, N14630);
buf BUF1 (N17109, N17105);
or OR3 (N17110, N17107, N10427, N4412);
or OR4 (N17111, N17055, N14382, N7285, N13751);
nor NOR3 (N17112, N17095, N4999, N8742);
nand NAND2 (N17113, N17110, N2968);
buf BUF1 (N17114, N17106);
or OR4 (N17115, N17109, N7763, N13905, N13092);
nor NOR2 (N17116, N17115, N12847);
and AND4 (N17117, N17112, N14462, N354, N15181);
not NOT1 (N17118, N17117);
and AND4 (N17119, N17116, N15237, N154, N15074);
nor NOR4 (N17120, N17102, N11970, N5131, N3171);
or OR2 (N17121, N17080, N588);
xor XOR2 (N17122, N17119, N9706);
xor XOR2 (N17123, N17122, N16804);
not NOT1 (N17124, N17123);
not NOT1 (N17125, N17108);
or OR3 (N17126, N17098, N5039, N5804);
buf BUF1 (N17127, N17118);
nand NAND4 (N17128, N17114, N12930, N13707, N7631);
buf BUF1 (N17129, N17128);
xor XOR2 (N17130, N17125, N11040);
nor NOR3 (N17131, N17101, N2958, N16657);
nor NOR2 (N17132, N17129, N9658);
buf BUF1 (N17133, N17132);
buf BUF1 (N17134, N17121);
nand NAND2 (N17135, N17126, N14992);
and AND4 (N17136, N17120, N16480, N1493, N4044);
not NOT1 (N17137, N17134);
buf BUF1 (N17138, N17136);
xor XOR2 (N17139, N17127, N2980);
or OR2 (N17140, N17135, N6734);
buf BUF1 (N17141, N17138);
buf BUF1 (N17142, N17124);
or OR3 (N17143, N17133, N10120, N1595);
not NOT1 (N17144, N17140);
or OR2 (N17145, N17139, N5567);
nand NAND3 (N17146, N17130, N14466, N4235);
xor XOR2 (N17147, N17146, N11146);
buf BUF1 (N17148, N17147);
not NOT1 (N17149, N17143);
xor XOR2 (N17150, N17149, N2743);
nor NOR4 (N17151, N17141, N3174, N14743, N7139);
nand NAND2 (N17152, N17151, N5703);
buf BUF1 (N17153, N17142);
nand NAND3 (N17154, N17150, N891, N14389);
not NOT1 (N17155, N17111);
nand NAND4 (N17156, N17145, N3186, N2311, N13511);
and AND3 (N17157, N17137, N14441, N9775);
xor XOR2 (N17158, N17153, N4647);
or OR4 (N17159, N17152, N11915, N8611, N15864);
nand NAND4 (N17160, N17156, N4710, N3257, N5751);
not NOT1 (N17161, N17160);
nand NAND3 (N17162, N17113, N12330, N16457);
buf BUF1 (N17163, N17155);
and AND3 (N17164, N17162, N7169, N13200);
nor NOR3 (N17165, N17148, N194, N2351);
nor NOR4 (N17166, N17158, N7261, N1226, N4600);
buf BUF1 (N17167, N17164);
xor XOR2 (N17168, N17159, N8641);
nand NAND4 (N17169, N17144, N12708, N7430, N9237);
or OR4 (N17170, N17131, N15101, N9434, N16798);
nor NOR3 (N17171, N17157, N8418, N53);
buf BUF1 (N17172, N17171);
xor XOR2 (N17173, N17169, N4278);
or OR3 (N17174, N17154, N15447, N1391);
or OR4 (N17175, N17163, N9091, N13252, N16918);
not NOT1 (N17176, N17167);
xor XOR2 (N17177, N17168, N2818);
or OR2 (N17178, N17161, N4854);
nor NOR3 (N17179, N17178, N13351, N10248);
nand NAND4 (N17180, N17172, N5155, N4399, N1280);
xor XOR2 (N17181, N17180, N293);
or OR2 (N17182, N17177, N7551);
not NOT1 (N17183, N17170);
xor XOR2 (N17184, N17173, N2117);
buf BUF1 (N17185, N17165);
and AND2 (N17186, N17184, N3443);
nor NOR3 (N17187, N17186, N5630, N14205);
not NOT1 (N17188, N17176);
nand NAND4 (N17189, N17182, N11323, N5413, N12057);
nor NOR4 (N17190, N17189, N13315, N5897, N9075);
xor XOR2 (N17191, N17175, N10221);
and AND3 (N17192, N17187, N6049, N7111);
xor XOR2 (N17193, N17188, N6807);
not NOT1 (N17194, N17192);
or OR3 (N17195, N17181, N3093, N12247);
buf BUF1 (N17196, N17179);
nand NAND2 (N17197, N17166, N11900);
nand NAND4 (N17198, N17196, N13374, N12586, N3638);
not NOT1 (N17199, N17193);
nor NOR4 (N17200, N17190, N2541, N10479, N8566);
xor XOR2 (N17201, N17200, N4252);
xor XOR2 (N17202, N17174, N14770);
xor XOR2 (N17203, N17194, N13714);
or OR3 (N17204, N17185, N4471, N5129);
or OR4 (N17205, N17195, N3817, N10579, N11401);
or OR2 (N17206, N17199, N4356);
buf BUF1 (N17207, N17201);
nand NAND3 (N17208, N17183, N4458, N15391);
not NOT1 (N17209, N17205);
buf BUF1 (N17210, N17209);
not NOT1 (N17211, N17210);
and AND3 (N17212, N17207, N8851, N1065);
nor NOR3 (N17213, N17203, N13401, N8838);
xor XOR2 (N17214, N17211, N16333);
nor NOR4 (N17215, N17214, N8008, N9802, N12085);
or OR2 (N17216, N17191, N9779);
nor NOR3 (N17217, N17202, N15811, N13127);
buf BUF1 (N17218, N17213);
and AND3 (N17219, N17197, N2104, N13296);
nand NAND4 (N17220, N17215, N10966, N4225, N7814);
nor NOR4 (N17221, N17198, N15647, N6408, N7653);
buf BUF1 (N17222, N17221);
nand NAND2 (N17223, N17220, N7176);
xor XOR2 (N17224, N17218, N8164);
or OR4 (N17225, N17216, N5581, N10601, N1176);
xor XOR2 (N17226, N17212, N8325);
nor NOR4 (N17227, N17206, N7085, N8004, N11998);
nand NAND3 (N17228, N17223, N9672, N7858);
buf BUF1 (N17229, N17225);
buf BUF1 (N17230, N17204);
buf BUF1 (N17231, N17226);
not NOT1 (N17232, N17222);
nor NOR4 (N17233, N17224, N9945, N16083, N13235);
xor XOR2 (N17234, N17231, N6110);
nand NAND2 (N17235, N17233, N9497);
nand NAND2 (N17236, N17217, N3161);
not NOT1 (N17237, N17236);
nand NAND2 (N17238, N17232, N10266);
nor NOR4 (N17239, N17234, N6042, N9816, N12429);
xor XOR2 (N17240, N17238, N10285);
buf BUF1 (N17241, N17227);
nor NOR3 (N17242, N17237, N6621, N17123);
nor NOR3 (N17243, N17228, N16234, N14493);
or OR2 (N17244, N17230, N13473);
nand NAND3 (N17245, N17229, N7452, N4858);
and AND3 (N17246, N17240, N895, N8697);
nor NOR2 (N17247, N17235, N8693);
nand NAND4 (N17248, N17244, N8417, N5375, N2340);
not NOT1 (N17249, N17242);
or OR2 (N17250, N17249, N12785);
not NOT1 (N17251, N17241);
or OR2 (N17252, N17219, N12458);
xor XOR2 (N17253, N17245, N14952);
nor NOR3 (N17254, N17251, N15705, N16717);
xor XOR2 (N17255, N17253, N14909);
not NOT1 (N17256, N17239);
not NOT1 (N17257, N17256);
and AND4 (N17258, N17254, N181, N15295, N16984);
xor XOR2 (N17259, N17250, N2795);
and AND4 (N17260, N17247, N1151, N15258, N5384);
not NOT1 (N17261, N17258);
buf BUF1 (N17262, N17248);
not NOT1 (N17263, N17262);
or OR3 (N17264, N17208, N3837, N8292);
nor NOR4 (N17265, N17243, N13988, N7651, N9798);
nand NAND2 (N17266, N17259, N6626);
xor XOR2 (N17267, N17266, N16387);
nand NAND3 (N17268, N17261, N10117, N4503);
nand NAND2 (N17269, N17257, N11108);
not NOT1 (N17270, N17265);
and AND4 (N17271, N17252, N1764, N10590, N15224);
and AND3 (N17272, N17267, N16920, N75);
or OR2 (N17273, N17246, N7389);
buf BUF1 (N17274, N17269);
nor NOR2 (N17275, N17271, N16424);
not NOT1 (N17276, N17255);
xor XOR2 (N17277, N17263, N7193);
not NOT1 (N17278, N17268);
xor XOR2 (N17279, N17274, N7296);
nand NAND2 (N17280, N17264, N11361);
xor XOR2 (N17281, N17270, N2685);
nor NOR4 (N17282, N17276, N5366, N9247, N4758);
and AND4 (N17283, N17272, N10264, N10185, N15747);
and AND4 (N17284, N17273, N6070, N10993, N13165);
buf BUF1 (N17285, N17282);
nand NAND2 (N17286, N17285, N14343);
xor XOR2 (N17287, N17284, N12806);
nand NAND3 (N17288, N17286, N7890, N16879);
not NOT1 (N17289, N17277);
xor XOR2 (N17290, N17260, N13189);
not NOT1 (N17291, N17281);
or OR3 (N17292, N17280, N11750, N13551);
nor NOR4 (N17293, N17279, N1890, N6808, N646);
buf BUF1 (N17294, N17278);
buf BUF1 (N17295, N17292);
xor XOR2 (N17296, N17293, N8911);
buf BUF1 (N17297, N17289);
not NOT1 (N17298, N17283);
and AND4 (N17299, N17291, N9705, N9495, N573);
buf BUF1 (N17300, N17299);
and AND3 (N17301, N17300, N573, N11437);
xor XOR2 (N17302, N17301, N16568);
nand NAND2 (N17303, N17290, N3272);
not NOT1 (N17304, N17275);
buf BUF1 (N17305, N17294);
nor NOR4 (N17306, N17288, N13572, N2807, N16186);
and AND4 (N17307, N17303, N12374, N1371, N10164);
nand NAND2 (N17308, N17287, N10105);
buf BUF1 (N17309, N17308);
xor XOR2 (N17310, N17305, N2576);
buf BUF1 (N17311, N17302);
nor NOR2 (N17312, N17295, N3252);
and AND2 (N17313, N17307, N13027);
nor NOR4 (N17314, N17296, N4904, N2435, N16384);
and AND2 (N17315, N17313, N8179);
or OR2 (N17316, N17311, N13159);
nand NAND4 (N17317, N17316, N7017, N2830, N17261);
nor NOR4 (N17318, N17309, N13320, N10488, N10264);
xor XOR2 (N17319, N17315, N5616);
and AND4 (N17320, N17298, N13635, N10602, N4138);
buf BUF1 (N17321, N17314);
and AND3 (N17322, N17318, N11019, N16769);
or OR2 (N17323, N17320, N1868);
buf BUF1 (N17324, N17321);
nor NOR3 (N17325, N17306, N3362, N15841);
nor NOR3 (N17326, N17317, N1711, N6515);
nor NOR3 (N17327, N17323, N17223, N13982);
nor NOR3 (N17328, N17325, N6448, N2900);
xor XOR2 (N17329, N17312, N12527);
and AND3 (N17330, N17327, N5417, N16470);
not NOT1 (N17331, N17329);
nand NAND3 (N17332, N17326, N5937, N4296);
nor NOR2 (N17333, N17322, N5542);
nand NAND4 (N17334, N17333, N679, N12988, N10412);
or OR3 (N17335, N17319, N9362, N13430);
xor XOR2 (N17336, N17297, N9533);
nand NAND3 (N17337, N17335, N11683, N15477);
not NOT1 (N17338, N17324);
not NOT1 (N17339, N17328);
buf BUF1 (N17340, N17339);
or OR3 (N17341, N17330, N16842, N12186);
nand NAND3 (N17342, N17340, N9421, N11665);
buf BUF1 (N17343, N17334);
and AND2 (N17344, N17341, N9857);
not NOT1 (N17345, N17304);
not NOT1 (N17346, N17344);
or OR3 (N17347, N17310, N11012, N5624);
nor NOR3 (N17348, N17345, N9022, N15087);
xor XOR2 (N17349, N17337, N10089);
nor NOR2 (N17350, N17336, N9414);
nor NOR2 (N17351, N17343, N16162);
nor NOR3 (N17352, N17349, N10482, N4767);
nand NAND2 (N17353, N17347, N5481);
nand NAND3 (N17354, N17352, N5954, N1891);
buf BUF1 (N17355, N17346);
nand NAND4 (N17356, N17348, N1407, N10459, N5880);
and AND4 (N17357, N17353, N4825, N8423, N15833);
and AND3 (N17358, N17351, N10150, N279);
nor NOR3 (N17359, N17355, N14042, N10729);
nand NAND2 (N17360, N17331, N10325);
xor XOR2 (N17361, N17359, N1202);
and AND3 (N17362, N17338, N14609, N11356);
nor NOR2 (N17363, N17361, N16830);
not NOT1 (N17364, N17362);
nand NAND2 (N17365, N17342, N9026);
xor XOR2 (N17366, N17360, N7423);
or OR2 (N17367, N17356, N12533);
nand NAND3 (N17368, N17358, N5360, N615);
xor XOR2 (N17369, N17363, N11669);
buf BUF1 (N17370, N17367);
or OR2 (N17371, N17332, N6301);
and AND4 (N17372, N17368, N4361, N9299, N14392);
buf BUF1 (N17373, N17364);
xor XOR2 (N17374, N17371, N5079);
xor XOR2 (N17375, N17365, N640);
xor XOR2 (N17376, N17366, N1683);
nand NAND3 (N17377, N17350, N6288, N8721);
or OR3 (N17378, N17374, N5321, N11350);
xor XOR2 (N17379, N17369, N15202);
or OR3 (N17380, N17377, N17048, N373);
nand NAND2 (N17381, N17372, N16978);
buf BUF1 (N17382, N17357);
xor XOR2 (N17383, N17373, N16679);
nor NOR4 (N17384, N17375, N15995, N15798, N8677);
nand NAND2 (N17385, N17380, N2039);
xor XOR2 (N17386, N17381, N7766);
nand NAND3 (N17387, N17378, N5468, N4839);
not NOT1 (N17388, N17385);
not NOT1 (N17389, N17387);
buf BUF1 (N17390, N17376);
xor XOR2 (N17391, N17379, N16724);
or OR3 (N17392, N17386, N4427, N8258);
buf BUF1 (N17393, N17391);
xor XOR2 (N17394, N17393, N16287);
nor NOR3 (N17395, N17389, N15585, N16672);
or OR3 (N17396, N17354, N4958, N15116);
nor NOR2 (N17397, N17370, N11510);
not NOT1 (N17398, N17383);
or OR2 (N17399, N17392, N11842);
nand NAND2 (N17400, N17398, N16942);
buf BUF1 (N17401, N17400);
nor NOR2 (N17402, N17390, N17123);
not NOT1 (N17403, N17384);
nand NAND3 (N17404, N17396, N5378, N17176);
not NOT1 (N17405, N17382);
or OR3 (N17406, N17395, N12853, N3203);
or OR2 (N17407, N17402, N9639);
and AND2 (N17408, N17388, N16226);
not NOT1 (N17409, N17401);
nand NAND2 (N17410, N17409, N6627);
and AND2 (N17411, N17397, N2847);
and AND4 (N17412, N17406, N2051, N13418, N6055);
and AND3 (N17413, N17403, N12112, N2707);
and AND4 (N17414, N17408, N9581, N2899, N444);
and AND2 (N17415, N17405, N695);
buf BUF1 (N17416, N17414);
nor NOR4 (N17417, N17415, N12372, N12498, N10490);
nor NOR4 (N17418, N17416, N12152, N10807, N9412);
or OR2 (N17419, N17404, N12518);
not NOT1 (N17420, N17407);
and AND3 (N17421, N17410, N2485, N8045);
or OR4 (N17422, N17421, N7351, N10862, N12721);
not NOT1 (N17423, N17394);
not NOT1 (N17424, N17413);
not NOT1 (N17425, N17412);
and AND2 (N17426, N17419, N10675);
buf BUF1 (N17427, N17424);
and AND2 (N17428, N17423, N7203);
and AND2 (N17429, N17427, N6484);
or OR3 (N17430, N17417, N3876, N7277);
nand NAND3 (N17431, N17428, N17004, N10370);
not NOT1 (N17432, N17429);
buf BUF1 (N17433, N17426);
or OR3 (N17434, N17430, N1466, N5175);
nand NAND2 (N17435, N17411, N9823);
and AND2 (N17436, N17418, N1853);
nor NOR3 (N17437, N17431, N3223, N9576);
nand NAND4 (N17438, N17399, N4726, N7611, N6492);
and AND2 (N17439, N17422, N12920);
nor NOR3 (N17440, N17438, N2650, N12282);
nor NOR3 (N17441, N17420, N13358, N10090);
and AND4 (N17442, N17425, N736, N12392, N6838);
buf BUF1 (N17443, N17434);
buf BUF1 (N17444, N17433);
xor XOR2 (N17445, N17435, N13561);
not NOT1 (N17446, N17442);
not NOT1 (N17447, N17432);
buf BUF1 (N17448, N17444);
or OR2 (N17449, N17446, N14886);
not NOT1 (N17450, N17447);
buf BUF1 (N17451, N17437);
nor NOR3 (N17452, N17443, N8053, N12698);
not NOT1 (N17453, N17449);
nand NAND4 (N17454, N17448, N2386, N5291, N13755);
nand NAND4 (N17455, N17453, N14255, N13721, N6449);
xor XOR2 (N17456, N17436, N10856);
xor XOR2 (N17457, N17439, N15150);
or OR4 (N17458, N17440, N3587, N3580, N13778);
nand NAND3 (N17459, N17455, N16805, N4330);
buf BUF1 (N17460, N17454);
nor NOR4 (N17461, N17459, N4886, N17275, N9914);
not NOT1 (N17462, N17450);
not NOT1 (N17463, N17457);
nand NAND2 (N17464, N17452, N2038);
or OR4 (N17465, N17458, N13821, N15955, N2459);
xor XOR2 (N17466, N17463, N8838);
buf BUF1 (N17467, N17464);
buf BUF1 (N17468, N17461);
or OR3 (N17469, N17467, N6055, N7616);
buf BUF1 (N17470, N17465);
not NOT1 (N17471, N17468);
nand NAND2 (N17472, N17470, N16406);
xor XOR2 (N17473, N17445, N5513);
xor XOR2 (N17474, N17441, N12293);
or OR2 (N17475, N17471, N4573);
xor XOR2 (N17476, N17469, N15882);
not NOT1 (N17477, N17462);
buf BUF1 (N17478, N17451);
or OR4 (N17479, N17473, N2911, N4993, N2293);
not NOT1 (N17480, N17466);
or OR3 (N17481, N17476, N15332, N15188);
xor XOR2 (N17482, N17475, N7494);
and AND2 (N17483, N17474, N3133);
nor NOR2 (N17484, N17483, N1755);
nor NOR4 (N17485, N17484, N16026, N6953, N11228);
nand NAND3 (N17486, N17477, N8329, N3036);
nor NOR4 (N17487, N17481, N1178, N2920, N3858);
not NOT1 (N17488, N17478);
nor NOR3 (N17489, N17486, N564, N2110);
or OR2 (N17490, N17456, N3298);
buf BUF1 (N17491, N17487);
and AND2 (N17492, N17482, N16069);
not NOT1 (N17493, N17488);
xor XOR2 (N17494, N17491, N1600);
nand NAND3 (N17495, N17490, N8072, N16456);
xor XOR2 (N17496, N17495, N13264);
xor XOR2 (N17497, N17496, N16950);
not NOT1 (N17498, N17480);
xor XOR2 (N17499, N17460, N9115);
xor XOR2 (N17500, N17498, N12755);
xor XOR2 (N17501, N17485, N16844);
buf BUF1 (N17502, N17497);
xor XOR2 (N17503, N17493, N2889);
nor NOR2 (N17504, N17489, N4879);
or OR4 (N17505, N17492, N13755, N12451, N13520);
not NOT1 (N17506, N17499);
and AND3 (N17507, N17500, N11412, N17073);
nand NAND2 (N17508, N17472, N1847);
buf BUF1 (N17509, N17504);
or OR4 (N17510, N17502, N1667, N12476, N10162);
nor NOR2 (N17511, N17503, N9022);
not NOT1 (N17512, N17509);
nor NOR2 (N17513, N17505, N11470);
xor XOR2 (N17514, N17512, N14922);
nor NOR2 (N17515, N17479, N14767);
not NOT1 (N17516, N17514);
or OR4 (N17517, N17511, N2156, N4512, N12099);
or OR2 (N17518, N17517, N2022);
buf BUF1 (N17519, N17513);
buf BUF1 (N17520, N17519);
nor NOR2 (N17521, N17516, N11843);
and AND4 (N17522, N17510, N12618, N12418, N7729);
buf BUF1 (N17523, N17515);
buf BUF1 (N17524, N17522);
nand NAND3 (N17525, N17507, N4042, N10148);
or OR2 (N17526, N17524, N3243);
nor NOR2 (N17527, N17521, N16804);
and AND3 (N17528, N17494, N12087, N10782);
nand NAND3 (N17529, N17523, N14140, N13737);
buf BUF1 (N17530, N17518);
or OR3 (N17531, N17520, N8310, N16137);
buf BUF1 (N17532, N17526);
nand NAND2 (N17533, N17530, N651);
nand NAND4 (N17534, N17531, N12271, N3249, N11417);
buf BUF1 (N17535, N17534);
xor XOR2 (N17536, N17529, N399);
nand NAND3 (N17537, N17525, N13041, N11193);
not NOT1 (N17538, N17501);
nor NOR4 (N17539, N17527, N14514, N2545, N12398);
nor NOR2 (N17540, N17506, N14733);
nand NAND3 (N17541, N17532, N16063, N15860);
not NOT1 (N17542, N17541);
nor NOR4 (N17543, N17533, N17236, N1657, N1540);
and AND3 (N17544, N17535, N13166, N10774);
not NOT1 (N17545, N17508);
xor XOR2 (N17546, N17538, N16014);
nand NAND4 (N17547, N17528, N251, N5929, N15424);
xor XOR2 (N17548, N17540, N15022);
or OR4 (N17549, N17536, N6038, N17180, N13700);
xor XOR2 (N17550, N17548, N14263);
xor XOR2 (N17551, N17539, N10433);
nor NOR3 (N17552, N17544, N3050, N4514);
xor XOR2 (N17553, N17551, N6300);
buf BUF1 (N17554, N17543);
xor XOR2 (N17555, N17545, N4149);
and AND2 (N17556, N17546, N8009);
not NOT1 (N17557, N17555);
and AND4 (N17558, N17550, N2331, N12915, N1855);
and AND4 (N17559, N17556, N886, N10604, N4816);
and AND2 (N17560, N17537, N13111);
nor NOR4 (N17561, N17542, N8091, N16792, N14503);
not NOT1 (N17562, N17553);
xor XOR2 (N17563, N17549, N16094);
nand NAND3 (N17564, N17547, N9493, N12854);
nor NOR2 (N17565, N17557, N1930);
buf BUF1 (N17566, N17558);
or OR3 (N17567, N17563, N10712, N6607);
nand NAND3 (N17568, N17559, N4280, N9368);
or OR2 (N17569, N17560, N12578);
not NOT1 (N17570, N17568);
buf BUF1 (N17571, N17562);
xor XOR2 (N17572, N17566, N6212);
nor NOR3 (N17573, N17564, N5668, N1517);
nand NAND4 (N17574, N17570, N13436, N16065, N12737);
nor NOR4 (N17575, N17554, N14211, N13433, N15060);
xor XOR2 (N17576, N17561, N5618);
xor XOR2 (N17577, N17571, N15059);
nor NOR4 (N17578, N17573, N14502, N15404, N16905);
xor XOR2 (N17579, N17578, N8322);
nor NOR4 (N17580, N17552, N11220, N2440, N7693);
buf BUF1 (N17581, N17577);
and AND3 (N17582, N17565, N575, N16912);
nand NAND2 (N17583, N17581, N4631);
nor NOR2 (N17584, N17582, N12341);
buf BUF1 (N17585, N17574);
nor NOR4 (N17586, N17584, N6243, N17016, N7995);
not NOT1 (N17587, N17585);
buf BUF1 (N17588, N17579);
buf BUF1 (N17589, N17583);
not NOT1 (N17590, N17589);
not NOT1 (N17591, N17575);
or OR3 (N17592, N17580, N6596, N15621);
buf BUF1 (N17593, N17569);
nand NAND2 (N17594, N17587, N15459);
nor NOR3 (N17595, N17572, N3040, N15953);
xor XOR2 (N17596, N17594, N16955);
nor NOR3 (N17597, N17593, N1096, N14830);
nand NAND4 (N17598, N17567, N1696, N16133, N4757);
nor NOR4 (N17599, N17595, N8329, N15044, N1125);
and AND4 (N17600, N17596, N308, N14168, N17067);
and AND2 (N17601, N17591, N15140);
or OR2 (N17602, N17601, N8776);
buf BUF1 (N17603, N17590);
or OR4 (N17604, N17597, N10800, N9964, N14523);
or OR2 (N17605, N17599, N280);
nand NAND2 (N17606, N17603, N11392);
or OR4 (N17607, N17592, N6256, N9464, N3572);
buf BUF1 (N17608, N17606);
nor NOR2 (N17609, N17600, N3766);
or OR2 (N17610, N17588, N14528);
nor NOR4 (N17611, N17604, N12714, N9878, N3852);
nand NAND4 (N17612, N17609, N3211, N15410, N68);
buf BUF1 (N17613, N17602);
or OR3 (N17614, N17605, N13295, N2093);
and AND2 (N17615, N17611, N17129);
and AND2 (N17616, N17607, N7866);
nand NAND2 (N17617, N17613, N11678);
nand NAND2 (N17618, N17612, N15262);
not NOT1 (N17619, N17576);
and AND3 (N17620, N17586, N3080, N13520);
xor XOR2 (N17621, N17615, N5188);
or OR2 (N17622, N17620, N17146);
and AND4 (N17623, N17622, N13045, N5555, N13264);
or OR3 (N17624, N17618, N12055, N5247);
nor NOR2 (N17625, N17623, N4799);
not NOT1 (N17626, N17614);
nand NAND3 (N17627, N17598, N17480, N7644);
nor NOR2 (N17628, N17608, N401);
xor XOR2 (N17629, N17619, N3930);
nand NAND4 (N17630, N17629, N2041, N1570, N4593);
and AND3 (N17631, N17630, N17000, N1124);
nor NOR3 (N17632, N17624, N6239, N1069);
and AND4 (N17633, N17625, N1164, N2716, N14024);
xor XOR2 (N17634, N17628, N11537);
nand NAND4 (N17635, N17627, N7229, N11300, N300);
nand NAND3 (N17636, N17635, N10515, N1236);
or OR4 (N17637, N17634, N10581, N6685, N10684);
buf BUF1 (N17638, N17636);
nand NAND2 (N17639, N17637, N9954);
not NOT1 (N17640, N17610);
nor NOR3 (N17641, N17616, N17278, N4031);
nor NOR2 (N17642, N17633, N15280);
or OR4 (N17643, N17621, N1187, N5323, N12122);
not NOT1 (N17644, N17642);
xor XOR2 (N17645, N17631, N390);
or OR4 (N17646, N17639, N4119, N14718, N11655);
buf BUF1 (N17647, N17644);
and AND3 (N17648, N17638, N9824, N10370);
nand NAND4 (N17649, N17646, N6238, N6714, N6270);
xor XOR2 (N17650, N17617, N8785);
buf BUF1 (N17651, N17643);
xor XOR2 (N17652, N17650, N2560);
xor XOR2 (N17653, N17651, N866);
and AND3 (N17654, N17648, N1770, N17326);
not NOT1 (N17655, N17649);
xor XOR2 (N17656, N17640, N1428);
or OR4 (N17657, N17647, N559, N15218, N3282);
not NOT1 (N17658, N17653);
buf BUF1 (N17659, N17656);
nand NAND2 (N17660, N17657, N7393);
buf BUF1 (N17661, N17641);
buf BUF1 (N17662, N17660);
not NOT1 (N17663, N17626);
or OR2 (N17664, N17645, N3814);
nand NAND3 (N17665, N17662, N15562, N8700);
not NOT1 (N17666, N17664);
buf BUF1 (N17667, N17666);
not NOT1 (N17668, N17654);
xor XOR2 (N17669, N17652, N5195);
not NOT1 (N17670, N17665);
and AND4 (N17671, N17655, N12877, N5789, N9478);
not NOT1 (N17672, N17667);
nand NAND3 (N17673, N17672, N13706, N13605);
buf BUF1 (N17674, N17668);
or OR3 (N17675, N17659, N11647, N2740);
nor NOR3 (N17676, N17658, N6876, N9647);
xor XOR2 (N17677, N17661, N14856);
nor NOR2 (N17678, N17673, N5022);
or OR4 (N17679, N17675, N11763, N1602, N215);
nor NOR3 (N17680, N17669, N17314, N11732);
or OR4 (N17681, N17676, N6034, N669, N16758);
xor XOR2 (N17682, N17671, N1219);
nand NAND4 (N17683, N17663, N16115, N1645, N4013);
xor XOR2 (N17684, N17670, N10668);
or OR2 (N17685, N17684, N15281);
or OR3 (N17686, N17685, N8192, N16438);
and AND4 (N17687, N17686, N3983, N15933, N5492);
not NOT1 (N17688, N17687);
nor NOR4 (N17689, N17674, N16279, N1574, N2646);
and AND2 (N17690, N17679, N16117);
buf BUF1 (N17691, N17681);
nand NAND2 (N17692, N17677, N5806);
xor XOR2 (N17693, N17680, N13206);
not NOT1 (N17694, N17691);
not NOT1 (N17695, N17690);
buf BUF1 (N17696, N17694);
or OR4 (N17697, N17689, N12152, N8191, N8511);
or OR4 (N17698, N17683, N846, N4134, N15010);
buf BUF1 (N17699, N17693);
or OR4 (N17700, N17697, N15200, N3077, N12237);
xor XOR2 (N17701, N17688, N12149);
nand NAND3 (N17702, N17701, N5381, N4414);
and AND3 (N17703, N17696, N17157, N12393);
buf BUF1 (N17704, N17702);
nand NAND3 (N17705, N17632, N1752, N2109);
or OR4 (N17706, N17682, N17224, N6061, N16675);
nor NOR3 (N17707, N17704, N14758, N5451);
and AND2 (N17708, N17703, N3746);
xor XOR2 (N17709, N17706, N16064);
not NOT1 (N17710, N17709);
nor NOR4 (N17711, N17692, N15597, N12632, N15593);
nand NAND4 (N17712, N17710, N3899, N7021, N6950);
not NOT1 (N17713, N17700);
and AND3 (N17714, N17698, N10308, N8861);
not NOT1 (N17715, N17699);
and AND2 (N17716, N17715, N15193);
or OR4 (N17717, N17716, N5839, N5069, N5604);
xor XOR2 (N17718, N17711, N4711);
nand NAND3 (N17719, N17695, N13469, N2264);
not NOT1 (N17720, N17712);
xor XOR2 (N17721, N17707, N2645);
buf BUF1 (N17722, N17720);
xor XOR2 (N17723, N17722, N6677);
nor NOR3 (N17724, N17717, N15478, N17158);
and AND3 (N17725, N17678, N1868, N4330);
nand NAND2 (N17726, N17708, N9955);
nor NOR4 (N17727, N17718, N15055, N13022, N13277);
or OR2 (N17728, N17719, N533);
buf BUF1 (N17729, N17705);
nor NOR3 (N17730, N17728, N8225, N1683);
buf BUF1 (N17731, N17713);
and AND2 (N17732, N17721, N1963);
nand NAND4 (N17733, N17723, N1283, N2094, N14082);
nor NOR2 (N17734, N17724, N9095);
or OR2 (N17735, N17734, N8366);
xor XOR2 (N17736, N17732, N1790);
buf BUF1 (N17737, N17733);
and AND3 (N17738, N17714, N16247, N3791);
xor XOR2 (N17739, N17726, N9394);
buf BUF1 (N17740, N17736);
nand NAND3 (N17741, N17739, N12445, N5288);
xor XOR2 (N17742, N17737, N3558);
buf BUF1 (N17743, N17730);
nor NOR4 (N17744, N17735, N7184, N12171, N15845);
nor NOR4 (N17745, N17727, N5846, N6864, N990);
nand NAND2 (N17746, N17741, N14567);
and AND3 (N17747, N17731, N1435, N16570);
not NOT1 (N17748, N17743);
or OR4 (N17749, N17747, N10045, N11544, N12715);
nor NOR4 (N17750, N17729, N9938, N4694, N11875);
xor XOR2 (N17751, N17748, N8596);
nand NAND3 (N17752, N17750, N14595, N6042);
nand NAND4 (N17753, N17725, N5780, N10255, N4907);
buf BUF1 (N17754, N17752);
not NOT1 (N17755, N17742);
not NOT1 (N17756, N17755);
buf BUF1 (N17757, N17738);
nor NOR4 (N17758, N17751, N9460, N13875, N11908);
and AND4 (N17759, N17753, N15933, N11489, N6380);
xor XOR2 (N17760, N17756, N10564);
buf BUF1 (N17761, N17760);
xor XOR2 (N17762, N17746, N5642);
or OR3 (N17763, N17740, N7420, N4444);
or OR2 (N17764, N17745, N6392);
nand NAND4 (N17765, N17749, N3371, N7718, N7917);
and AND2 (N17766, N17744, N6190);
nor NOR4 (N17767, N17761, N15891, N15348, N5887);
or OR2 (N17768, N17763, N6686);
xor XOR2 (N17769, N17759, N602);
xor XOR2 (N17770, N17754, N6465);
buf BUF1 (N17771, N17767);
buf BUF1 (N17772, N17770);
not NOT1 (N17773, N17768);
not NOT1 (N17774, N17765);
and AND2 (N17775, N17774, N17204);
and AND4 (N17776, N17757, N5982, N6882, N3680);
not NOT1 (N17777, N17758);
nor NOR2 (N17778, N17762, N10823);
not NOT1 (N17779, N17766);
nor NOR4 (N17780, N17772, N9133, N16768, N16919);
nor NOR4 (N17781, N17778, N8083, N12946, N7782);
or OR3 (N17782, N17764, N2481, N9192);
buf BUF1 (N17783, N17782);
nor NOR2 (N17784, N17771, N4742);
and AND3 (N17785, N17773, N15111, N33);
xor XOR2 (N17786, N17780, N16816);
nor NOR4 (N17787, N17785, N10666, N14068, N9698);
xor XOR2 (N17788, N17779, N14120);
and AND4 (N17789, N17783, N1355, N7853, N13319);
or OR4 (N17790, N17776, N14507, N12033, N1861);
or OR2 (N17791, N17789, N17166);
nand NAND3 (N17792, N17788, N11843, N1360);
buf BUF1 (N17793, N17775);
not NOT1 (N17794, N17793);
not NOT1 (N17795, N17792);
not NOT1 (N17796, N17786);
xor XOR2 (N17797, N17794, N13880);
not NOT1 (N17798, N17787);
xor XOR2 (N17799, N17798, N15353);
xor XOR2 (N17800, N17781, N4967);
not NOT1 (N17801, N17791);
xor XOR2 (N17802, N17784, N16013);
buf BUF1 (N17803, N17769);
or OR2 (N17804, N17799, N5486);
buf BUF1 (N17805, N17795);
buf BUF1 (N17806, N17802);
and AND3 (N17807, N17777, N7195, N13646);
xor XOR2 (N17808, N17803, N11181);
nor NOR3 (N17809, N17801, N9223, N4952);
xor XOR2 (N17810, N17805, N4640);
and AND3 (N17811, N17797, N3374, N6898);
not NOT1 (N17812, N17808);
and AND4 (N17813, N17812, N2914, N7667, N7412);
and AND4 (N17814, N17809, N10796, N10479, N16753);
and AND2 (N17815, N17790, N11863);
or OR4 (N17816, N17807, N5124, N6668, N879);
xor XOR2 (N17817, N17815, N7670);
buf BUF1 (N17818, N17814);
xor XOR2 (N17819, N17796, N8066);
not NOT1 (N17820, N17800);
or OR2 (N17821, N17804, N4939);
not NOT1 (N17822, N17817);
nor NOR3 (N17823, N17819, N4834, N54);
xor XOR2 (N17824, N17818, N16612);
buf BUF1 (N17825, N17822);
and AND4 (N17826, N17824, N2139, N7658, N4682);
buf BUF1 (N17827, N17813);
buf BUF1 (N17828, N17823);
or OR3 (N17829, N17820, N9363, N5862);
not NOT1 (N17830, N17825);
or OR3 (N17831, N17806, N8024, N7707);
buf BUF1 (N17832, N17829);
nand NAND3 (N17833, N17826, N16969, N16898);
xor XOR2 (N17834, N17832, N15327);
and AND3 (N17835, N17821, N16748, N16785);
nand NAND4 (N17836, N17816, N4886, N3185, N17547);
xor XOR2 (N17837, N17835, N17653);
nand NAND3 (N17838, N17836, N14230, N12058);
xor XOR2 (N17839, N17834, N9349);
nand NAND4 (N17840, N17811, N11817, N7964, N1976);
buf BUF1 (N17841, N17837);
or OR4 (N17842, N17828, N7727, N7663, N4866);
xor XOR2 (N17843, N17838, N16697);
not NOT1 (N17844, N17831);
nand NAND3 (N17845, N17839, N5810, N8388);
and AND3 (N17846, N17844, N9346, N11436);
or OR4 (N17847, N17827, N15787, N14602, N11597);
xor XOR2 (N17848, N17840, N13635);
not NOT1 (N17849, N17846);
not NOT1 (N17850, N17847);
not NOT1 (N17851, N17843);
and AND2 (N17852, N17845, N537);
not NOT1 (N17853, N17830);
not NOT1 (N17854, N17810);
and AND2 (N17855, N17854, N7487);
and AND4 (N17856, N17855, N7563, N6979, N1587);
buf BUF1 (N17857, N17842);
nand NAND3 (N17858, N17852, N15412, N11458);
not NOT1 (N17859, N17849);
xor XOR2 (N17860, N17856, N12691);
not NOT1 (N17861, N17833);
not NOT1 (N17862, N17850);
not NOT1 (N17863, N17848);
buf BUF1 (N17864, N17861);
nor NOR4 (N17865, N17851, N3670, N874, N5008);
nand NAND2 (N17866, N17857, N7078);
and AND4 (N17867, N17865, N210, N127, N11123);
not NOT1 (N17868, N17862);
not NOT1 (N17869, N17864);
not NOT1 (N17870, N17866);
xor XOR2 (N17871, N17858, N10793);
and AND2 (N17872, N17853, N17482);
or OR4 (N17873, N17841, N8945, N13899, N9507);
nor NOR3 (N17874, N17859, N10602, N17291);
xor XOR2 (N17875, N17867, N5536);
xor XOR2 (N17876, N17868, N11725);
or OR3 (N17877, N17860, N5893, N501);
or OR2 (N17878, N17874, N15545);
or OR2 (N17879, N17877, N3836);
or OR3 (N17880, N17869, N2040, N15868);
nand NAND4 (N17881, N17875, N14678, N14469, N4342);
not NOT1 (N17882, N17878);
buf BUF1 (N17883, N17881);
and AND4 (N17884, N17870, N17419, N12365, N16931);
nand NAND2 (N17885, N17872, N9548);
buf BUF1 (N17886, N17884);
and AND4 (N17887, N17879, N10803, N2726, N10325);
nand NAND2 (N17888, N17885, N15556);
buf BUF1 (N17889, N17876);
or OR2 (N17890, N17888, N1106);
or OR4 (N17891, N17887, N3592, N11176, N4719);
and AND3 (N17892, N17889, N7800, N16274);
nor NOR3 (N17893, N17891, N17126, N6193);
and AND4 (N17894, N17873, N13122, N11051, N14004);
buf BUF1 (N17895, N17893);
and AND4 (N17896, N17871, N7551, N12481, N957);
not NOT1 (N17897, N17882);
or OR4 (N17898, N17897, N12337, N13963, N5301);
not NOT1 (N17899, N17898);
xor XOR2 (N17900, N17886, N3617);
not NOT1 (N17901, N17883);
or OR4 (N17902, N17896, N14165, N14707, N2633);
and AND3 (N17903, N17880, N6418, N16862);
buf BUF1 (N17904, N17895);
buf BUF1 (N17905, N17903);
buf BUF1 (N17906, N17901);
buf BUF1 (N17907, N17863);
nand NAND3 (N17908, N17894, N15104, N7287);
or OR4 (N17909, N17906, N14251, N4033, N3533);
nand NAND4 (N17910, N17905, N16103, N12579, N7990);
nand NAND3 (N17911, N17904, N14341, N14389);
nor NOR3 (N17912, N17908, N5154, N14153);
nor NOR3 (N17913, N17907, N15607, N959);
nor NOR3 (N17914, N17902, N11647, N7071);
xor XOR2 (N17915, N17913, N16157);
not NOT1 (N17916, N17915);
nor NOR2 (N17917, N17914, N767);
or OR2 (N17918, N17899, N12417);
xor XOR2 (N17919, N17917, N1826);
nor NOR2 (N17920, N17909, N10708);
and AND4 (N17921, N17892, N2274, N8339, N5702);
xor XOR2 (N17922, N17900, N16466);
buf BUF1 (N17923, N17918);
and AND2 (N17924, N17916, N932);
nor NOR2 (N17925, N17922, N352);
nand NAND4 (N17926, N17920, N10163, N4161, N14967);
xor XOR2 (N17927, N17912, N12016);
not NOT1 (N17928, N17919);
xor XOR2 (N17929, N17927, N16066);
or OR2 (N17930, N17911, N16578);
nor NOR3 (N17931, N17929, N17461, N13736);
not NOT1 (N17932, N17924);
and AND4 (N17933, N17928, N9794, N1232, N6092);
nand NAND4 (N17934, N17932, N2440, N5245, N12091);
nand NAND4 (N17935, N17890, N16076, N13449, N16782);
not NOT1 (N17936, N17935);
and AND3 (N17937, N17936, N366, N11211);
and AND3 (N17938, N17923, N3921, N14280);
xor XOR2 (N17939, N17926, N4910);
and AND3 (N17940, N17921, N11008, N17201);
and AND3 (N17941, N17934, N2768, N6233);
nand NAND3 (N17942, N17930, N1056, N936);
nor NOR3 (N17943, N17910, N9352, N1223);
nand NAND4 (N17944, N17933, N5925, N1736, N17475);
nand NAND3 (N17945, N17943, N13912, N16352);
not NOT1 (N17946, N17942);
buf BUF1 (N17947, N17941);
not NOT1 (N17948, N17939);
nor NOR4 (N17949, N17945, N5133, N7789, N16937);
buf BUF1 (N17950, N17948);
buf BUF1 (N17951, N17937);
or OR3 (N17952, N17940, N15436, N1302);
buf BUF1 (N17953, N17952);
nor NOR4 (N17954, N17949, N13673, N13675, N9283);
or OR2 (N17955, N17938, N4975);
xor XOR2 (N17956, N17947, N8413);
buf BUF1 (N17957, N17925);
and AND4 (N17958, N17956, N472, N12741, N6418);
nand NAND4 (N17959, N17955, N17633, N7452, N3304);
or OR4 (N17960, N17946, N13414, N2930, N10539);
and AND3 (N17961, N17958, N6732, N14244);
and AND4 (N17962, N17951, N4561, N2007, N3617);
not NOT1 (N17963, N17961);
buf BUF1 (N17964, N17953);
nand NAND2 (N17965, N17959, N10905);
xor XOR2 (N17966, N17964, N3456);
nor NOR4 (N17967, N17950, N17747, N8291, N4117);
buf BUF1 (N17968, N17966);
not NOT1 (N17969, N17968);
nand NAND3 (N17970, N17963, N8283, N16466);
buf BUF1 (N17971, N17970);
xor XOR2 (N17972, N17967, N5746);
not NOT1 (N17973, N17962);
and AND2 (N17974, N17972, N15769);
nor NOR4 (N17975, N17969, N14431, N6148, N6913);
buf BUF1 (N17976, N17965);
xor XOR2 (N17977, N17975, N6845);
nand NAND4 (N17978, N17973, N13261, N11710, N4984);
and AND4 (N17979, N17944, N14809, N385, N2833);
and AND3 (N17980, N17960, N5208, N12065);
xor XOR2 (N17981, N17954, N6472);
buf BUF1 (N17982, N17978);
nor NOR2 (N17983, N17979, N15836);
or OR4 (N17984, N17983, N13281, N5140, N15368);
nand NAND2 (N17985, N17982, N14170);
xor XOR2 (N17986, N17985, N10928);
not NOT1 (N17987, N17977);
not NOT1 (N17988, N17980);
xor XOR2 (N17989, N17988, N4513);
not NOT1 (N17990, N17981);
buf BUF1 (N17991, N17971);
nand NAND3 (N17992, N17989, N4650, N9307);
buf BUF1 (N17993, N17986);
xor XOR2 (N17994, N17974, N8526);
nand NAND4 (N17995, N17957, N15548, N3085, N16186);
nor NOR3 (N17996, N17931, N16916, N11350);
nor NOR3 (N17997, N17994, N740, N16595);
nand NAND4 (N17998, N17992, N16722, N9163, N13746);
buf BUF1 (N17999, N17996);
nand NAND2 (N18000, N17976, N16121);
or OR3 (N18001, N17993, N6607, N7882);
and AND3 (N18002, N17998, N6552, N11621);
or OR3 (N18003, N17984, N4250, N9039);
not NOT1 (N18004, N17990);
xor XOR2 (N18005, N18003, N927);
xor XOR2 (N18006, N18004, N17127);
not NOT1 (N18007, N18006);
nand NAND2 (N18008, N17987, N3232);
nor NOR4 (N18009, N18005, N572, N1192, N1799);
nand NAND2 (N18010, N18000, N62);
nand NAND2 (N18011, N18008, N7511);
buf BUF1 (N18012, N18011);
nand NAND2 (N18013, N18010, N11260);
nand NAND2 (N18014, N17995, N7872);
nor NOR2 (N18015, N18007, N10351);
or OR4 (N18016, N18015, N7357, N1429, N4997);
xor XOR2 (N18017, N18016, N8105);
nand NAND4 (N18018, N18017, N7932, N14796, N7572);
or OR4 (N18019, N17999, N14710, N3254, N8380);
or OR2 (N18020, N18002, N15468);
xor XOR2 (N18021, N17997, N1600);
nor NOR2 (N18022, N18009, N16753);
xor XOR2 (N18023, N17991, N16631);
xor XOR2 (N18024, N18022, N15710);
not NOT1 (N18025, N18024);
xor XOR2 (N18026, N18020, N7150);
or OR4 (N18027, N18021, N10474, N1893, N2707);
xor XOR2 (N18028, N18026, N3704);
xor XOR2 (N18029, N18025, N11990);
or OR3 (N18030, N18028, N4807, N14431);
buf BUF1 (N18031, N18014);
xor XOR2 (N18032, N18030, N3466);
nand NAND2 (N18033, N18013, N14154);
nor NOR4 (N18034, N18023, N17411, N3445, N11752);
buf BUF1 (N18035, N18012);
or OR3 (N18036, N18018, N17354, N1092);
not NOT1 (N18037, N18001);
nor NOR4 (N18038, N18027, N14332, N10197, N8980);
or OR2 (N18039, N18036, N13420);
or OR2 (N18040, N18037, N4319);
not NOT1 (N18041, N18032);
or OR3 (N18042, N18040, N15632, N13627);
and AND3 (N18043, N18039, N2915, N1047);
xor XOR2 (N18044, N18034, N16714);
or OR3 (N18045, N18019, N11573, N6839);
nand NAND2 (N18046, N18031, N1077);
and AND2 (N18047, N18043, N14081);
xor XOR2 (N18048, N18042, N15299);
buf BUF1 (N18049, N18033);
nor NOR2 (N18050, N18038, N1599);
or OR3 (N18051, N18041, N13161, N13121);
nand NAND3 (N18052, N18045, N869, N9130);
nand NAND3 (N18053, N18048, N60, N11408);
buf BUF1 (N18054, N18047);
xor XOR2 (N18055, N18029, N17993);
and AND3 (N18056, N18044, N5841, N1085);
nand NAND2 (N18057, N18050, N8575);
nor NOR2 (N18058, N18055, N926);
or OR4 (N18059, N18046, N1877, N1882, N2270);
nor NOR4 (N18060, N18056, N8842, N15443, N8787);
buf BUF1 (N18061, N18060);
nand NAND2 (N18062, N18061, N9848);
xor XOR2 (N18063, N18053, N10917);
nand NAND2 (N18064, N18051, N9092);
xor XOR2 (N18065, N18052, N15506);
buf BUF1 (N18066, N18063);
and AND4 (N18067, N18062, N2439, N8531, N5951);
or OR4 (N18068, N18059, N1474, N10879, N8170);
buf BUF1 (N18069, N18065);
or OR3 (N18070, N18049, N10591, N12573);
xor XOR2 (N18071, N18070, N5871);
and AND3 (N18072, N18068, N11545, N12830);
nor NOR3 (N18073, N18054, N4863, N191);
or OR2 (N18074, N18072, N3998);
nor NOR2 (N18075, N18064, N3293);
not NOT1 (N18076, N18069);
xor XOR2 (N18077, N18067, N11117);
nand NAND4 (N18078, N18035, N15646, N15080, N11766);
not NOT1 (N18079, N18076);
not NOT1 (N18080, N18078);
nor NOR2 (N18081, N18057, N7862);
and AND2 (N18082, N18077, N4069);
xor XOR2 (N18083, N18066, N10297);
nand NAND3 (N18084, N18079, N12041, N8522);
xor XOR2 (N18085, N18074, N7210);
nor NOR4 (N18086, N18084, N3900, N9090, N282);
and AND3 (N18087, N18080, N13373, N10794);
buf BUF1 (N18088, N18082);
nand NAND4 (N18089, N18081, N12410, N5833, N859);
or OR3 (N18090, N18083, N1105, N17288);
nand NAND4 (N18091, N18058, N10997, N3350, N1633);
nor NOR2 (N18092, N18087, N7589);
nand NAND4 (N18093, N18092, N12444, N1579, N17273);
nor NOR3 (N18094, N18085, N14678, N445);
or OR3 (N18095, N18090, N5826, N10756);
not NOT1 (N18096, N18071);
and AND2 (N18097, N18088, N12665);
xor XOR2 (N18098, N18093, N372);
nand NAND3 (N18099, N18095, N13818, N6394);
nor NOR3 (N18100, N18086, N11056, N11407);
nand NAND2 (N18101, N18097, N16860);
and AND2 (N18102, N18100, N8596);
nand NAND4 (N18103, N18094, N13063, N8793, N16262);
nand NAND3 (N18104, N18102, N10611, N13008);
nor NOR2 (N18105, N18098, N15562);
or OR4 (N18106, N18105, N3894, N6179, N15935);
xor XOR2 (N18107, N18104, N15632);
xor XOR2 (N18108, N18091, N4526);
nand NAND3 (N18109, N18106, N2575, N18085);
or OR2 (N18110, N18103, N13046);
not NOT1 (N18111, N18110);
or OR2 (N18112, N18107, N17031);
and AND2 (N18113, N18112, N2015);
buf BUF1 (N18114, N18089);
or OR2 (N18115, N18101, N4542);
nand NAND2 (N18116, N18114, N17629);
nand NAND4 (N18117, N18116, N564, N1277, N6693);
and AND3 (N18118, N18111, N14937, N11435);
or OR3 (N18119, N18118, N17464, N8378);
nor NOR3 (N18120, N18096, N1126, N14037);
xor XOR2 (N18121, N18113, N14619);
or OR3 (N18122, N18121, N8607, N11415);
xor XOR2 (N18123, N18120, N2534);
xor XOR2 (N18124, N18099, N17828);
buf BUF1 (N18125, N18123);
or OR2 (N18126, N18108, N12690);
buf BUF1 (N18127, N18117);
xor XOR2 (N18128, N18119, N7109);
buf BUF1 (N18129, N18109);
not NOT1 (N18130, N18129);
or OR3 (N18131, N18115, N13062, N9398);
xor XOR2 (N18132, N18075, N14272);
not NOT1 (N18133, N18124);
and AND4 (N18134, N18128, N2800, N567, N12644);
nand NAND2 (N18135, N18126, N4072);
nor NOR4 (N18136, N18135, N698, N1510, N2874);
xor XOR2 (N18137, N18122, N9219);
xor XOR2 (N18138, N18133, N3155);
not NOT1 (N18139, N18127);
nor NOR2 (N18140, N18125, N9248);
nor NOR4 (N18141, N18073, N8979, N14563, N102);
or OR2 (N18142, N18137, N7733);
or OR4 (N18143, N18134, N6947, N11904, N3318);
nand NAND2 (N18144, N18140, N2813);
or OR3 (N18145, N18141, N15470, N16737);
buf BUF1 (N18146, N18130);
not NOT1 (N18147, N18144);
not NOT1 (N18148, N18132);
or OR4 (N18149, N18147, N16962, N9059, N14243);
and AND2 (N18150, N18148, N16828);
and AND2 (N18151, N18145, N17578);
buf BUF1 (N18152, N18139);
nor NOR2 (N18153, N18146, N14470);
and AND4 (N18154, N18131, N14727, N6342, N7722);
or OR3 (N18155, N18150, N17964, N14850);
or OR3 (N18156, N18151, N11744, N9806);
nand NAND2 (N18157, N18142, N5684);
not NOT1 (N18158, N18153);
not NOT1 (N18159, N18156);
nor NOR3 (N18160, N18159, N13240, N16922);
nor NOR3 (N18161, N18155, N7513, N8015);
or OR3 (N18162, N18154, N14173, N4180);
or OR2 (N18163, N18162, N15914);
xor XOR2 (N18164, N18149, N11131);
nand NAND2 (N18165, N18136, N11193);
not NOT1 (N18166, N18158);
or OR3 (N18167, N18161, N10575, N14033);
or OR3 (N18168, N18166, N628, N689);
nand NAND3 (N18169, N18165, N4538, N9348);
nor NOR4 (N18170, N18152, N1693, N7906, N15347);
or OR4 (N18171, N18138, N8482, N9213, N7599);
not NOT1 (N18172, N18170);
buf BUF1 (N18173, N18172);
and AND4 (N18174, N18169, N7995, N15980, N9713);
xor XOR2 (N18175, N18164, N1522);
nor NOR3 (N18176, N18171, N812, N1258);
or OR3 (N18177, N18174, N17070, N104);
not NOT1 (N18178, N18168);
buf BUF1 (N18179, N18176);
and AND2 (N18180, N18173, N10085);
or OR4 (N18181, N18179, N8095, N8237, N15861);
nand NAND4 (N18182, N18177, N7822, N11624, N6160);
nor NOR4 (N18183, N18175, N15205, N9001, N11784);
and AND2 (N18184, N18178, N11040);
nor NOR2 (N18185, N18182, N524);
or OR3 (N18186, N18183, N13613, N14786);
and AND2 (N18187, N18143, N6024);
nor NOR2 (N18188, N18187, N16218);
and AND2 (N18189, N18163, N2529);
nand NAND2 (N18190, N18180, N15297);
buf BUF1 (N18191, N18190);
and AND4 (N18192, N18188, N7339, N16803, N9061);
not NOT1 (N18193, N18185);
and AND3 (N18194, N18191, N8586, N12711);
nand NAND3 (N18195, N18186, N6990, N5622);
nand NAND4 (N18196, N18167, N1292, N10091, N12933);
not NOT1 (N18197, N18192);
nand NAND2 (N18198, N18194, N15444);
nor NOR3 (N18199, N18181, N7574, N10697);
nor NOR2 (N18200, N18199, N5023);
not NOT1 (N18201, N18193);
and AND3 (N18202, N18196, N8409, N2769);
xor XOR2 (N18203, N18198, N16979);
nand NAND2 (N18204, N18184, N3102);
buf BUF1 (N18205, N18200);
not NOT1 (N18206, N18160);
not NOT1 (N18207, N18206);
and AND4 (N18208, N18195, N16069, N857, N5888);
xor XOR2 (N18209, N18157, N12294);
and AND2 (N18210, N18209, N734);
not NOT1 (N18211, N18201);
or OR2 (N18212, N18202, N388);
nor NOR3 (N18213, N18210, N9789, N8745);
nor NOR4 (N18214, N18212, N16415, N15767, N3572);
nor NOR4 (N18215, N18213, N3211, N15404, N1847);
nand NAND4 (N18216, N18197, N10465, N5568, N18001);
nand NAND2 (N18217, N18214, N6302);
nor NOR2 (N18218, N18215, N356);
buf BUF1 (N18219, N18216);
and AND2 (N18220, N18211, N16554);
nand NAND3 (N18221, N18218, N11262, N6840);
not NOT1 (N18222, N18204);
or OR3 (N18223, N18221, N4489, N16654);
or OR2 (N18224, N18217, N14920);
nor NOR4 (N18225, N18203, N16579, N12063, N12185);
xor XOR2 (N18226, N18219, N9660);
not NOT1 (N18227, N18224);
buf BUF1 (N18228, N18207);
and AND4 (N18229, N18208, N18139, N1017, N14801);
and AND3 (N18230, N18223, N13663, N10504);
nor NOR4 (N18231, N18189, N4634, N12609, N9866);
nor NOR4 (N18232, N18231, N10961, N11282, N6397);
or OR2 (N18233, N18232, N393);
not NOT1 (N18234, N18228);
xor XOR2 (N18235, N18222, N10996);
buf BUF1 (N18236, N18230);
and AND2 (N18237, N18226, N9507);
not NOT1 (N18238, N18229);
buf BUF1 (N18239, N18238);
xor XOR2 (N18240, N18234, N17068);
nor NOR2 (N18241, N18239, N8032);
buf BUF1 (N18242, N18240);
buf BUF1 (N18243, N18237);
nor NOR2 (N18244, N18243, N12894);
not NOT1 (N18245, N18242);
buf BUF1 (N18246, N18205);
or OR4 (N18247, N18220, N16598, N2534, N12782);
not NOT1 (N18248, N18247);
and AND4 (N18249, N18227, N1790, N6470, N1490);
xor XOR2 (N18250, N18246, N15123);
buf BUF1 (N18251, N18233);
nand NAND4 (N18252, N18251, N1733, N8888, N418);
xor XOR2 (N18253, N18244, N18221);
not NOT1 (N18254, N18235);
xor XOR2 (N18255, N18245, N10671);
nand NAND4 (N18256, N18241, N4610, N1855, N6256);
buf BUF1 (N18257, N18249);
not NOT1 (N18258, N18253);
xor XOR2 (N18259, N18255, N10497);
buf BUF1 (N18260, N18259);
buf BUF1 (N18261, N18258);
nand NAND2 (N18262, N18257, N8055);
nor NOR2 (N18263, N18261, N9300);
or OR4 (N18264, N18263, N16820, N9408, N17352);
not NOT1 (N18265, N18252);
or OR4 (N18266, N18265, N1629, N5926, N10239);
xor XOR2 (N18267, N18256, N15277);
not NOT1 (N18268, N18254);
nand NAND2 (N18269, N18248, N13760);
not NOT1 (N18270, N18236);
or OR2 (N18271, N18268, N636);
nand NAND3 (N18272, N18225, N7938, N11069);
buf BUF1 (N18273, N18264);
xor XOR2 (N18274, N18260, N4249);
xor XOR2 (N18275, N18274, N12551);
nor NOR3 (N18276, N18273, N9390, N4180);
xor XOR2 (N18277, N18275, N3887);
xor XOR2 (N18278, N18276, N15818);
and AND3 (N18279, N18266, N2698, N7795);
buf BUF1 (N18280, N18270);
xor XOR2 (N18281, N18271, N16147);
or OR2 (N18282, N18267, N11915);
not NOT1 (N18283, N18272);
and AND3 (N18284, N18280, N8538, N671);
nor NOR3 (N18285, N18281, N3263, N13548);
nand NAND4 (N18286, N18283, N18049, N13294, N15445);
and AND2 (N18287, N18277, N2954);
or OR3 (N18288, N18279, N2780, N12401);
nor NOR3 (N18289, N18288, N9647, N11781);
and AND3 (N18290, N18285, N14956, N4222);
and AND2 (N18291, N18287, N14565);
nor NOR2 (N18292, N18278, N120);
nand NAND2 (N18293, N18269, N6820);
or OR2 (N18294, N18289, N9401);
not NOT1 (N18295, N18293);
buf BUF1 (N18296, N18295);
xor XOR2 (N18297, N18291, N1986);
xor XOR2 (N18298, N18284, N3575);
or OR2 (N18299, N18290, N15207);
xor XOR2 (N18300, N18294, N14223);
nand NAND3 (N18301, N18299, N12924, N18255);
buf BUF1 (N18302, N18301);
not NOT1 (N18303, N18297);
and AND2 (N18304, N18262, N12975);
xor XOR2 (N18305, N18302, N17467);
xor XOR2 (N18306, N18300, N12487);
or OR4 (N18307, N18306, N4117, N16605, N531);
buf BUF1 (N18308, N18286);
and AND4 (N18309, N18250, N13961, N13217, N18135);
nand NAND2 (N18310, N18296, N16955);
nand NAND4 (N18311, N18307, N8846, N14540, N3152);
nand NAND4 (N18312, N18308, N11649, N5988, N15488);
nor NOR4 (N18313, N18298, N9441, N8547, N15708);
not NOT1 (N18314, N18310);
nand NAND3 (N18315, N18311, N5055, N10065);
and AND3 (N18316, N18314, N10935, N15736);
xor XOR2 (N18317, N18309, N3326);
and AND2 (N18318, N18315, N12467);
or OR4 (N18319, N18305, N13227, N4763, N1931);
and AND3 (N18320, N18304, N15363, N14068);
nor NOR4 (N18321, N18319, N15987, N3203, N13518);
not NOT1 (N18322, N18321);
not NOT1 (N18323, N18317);
nor NOR2 (N18324, N18322, N16556);
or OR4 (N18325, N18316, N11733, N4224, N4627);
nand NAND4 (N18326, N18312, N11197, N9764, N9173);
xor XOR2 (N18327, N18320, N5477);
or OR2 (N18328, N18313, N16385);
nor NOR3 (N18329, N18324, N9122, N13668);
not NOT1 (N18330, N18326);
and AND4 (N18331, N18329, N10141, N17114, N9052);
xor XOR2 (N18332, N18292, N611);
not NOT1 (N18333, N18330);
nand NAND3 (N18334, N18325, N7589, N12569);
xor XOR2 (N18335, N18333, N9469);
xor XOR2 (N18336, N18335, N10791);
xor XOR2 (N18337, N18334, N1336);
buf BUF1 (N18338, N18337);
and AND4 (N18339, N18318, N535, N9056, N10686);
buf BUF1 (N18340, N18328);
nor NOR2 (N18341, N18282, N13983);
and AND2 (N18342, N18303, N3225);
nor NOR4 (N18343, N18323, N6737, N1862, N7042);
nand NAND3 (N18344, N18343, N1166, N15463);
or OR4 (N18345, N18339, N8116, N16760, N7671);
xor XOR2 (N18346, N18327, N10281);
not NOT1 (N18347, N18332);
buf BUF1 (N18348, N18340);
nor NOR3 (N18349, N18338, N706, N13058);
not NOT1 (N18350, N18349);
not NOT1 (N18351, N18345);
or OR3 (N18352, N18350, N7723, N679);
nand NAND4 (N18353, N18344, N2059, N4714, N10749);
nor NOR3 (N18354, N18341, N14426, N3484);
buf BUF1 (N18355, N18342);
and AND2 (N18356, N18346, N13393);
nand NAND4 (N18357, N18336, N7330, N12524, N7912);
xor XOR2 (N18358, N18351, N5849);
and AND4 (N18359, N18356, N1203, N5889, N8795);
and AND4 (N18360, N18352, N17183, N14607, N17661);
not NOT1 (N18361, N18348);
and AND2 (N18362, N18354, N14387);
xor XOR2 (N18363, N18360, N13335);
nor NOR4 (N18364, N18359, N13377, N6818, N11484);
buf BUF1 (N18365, N18362);
buf BUF1 (N18366, N18364);
nand NAND2 (N18367, N18365, N15068);
xor XOR2 (N18368, N18361, N17957);
not NOT1 (N18369, N18347);
or OR4 (N18370, N18367, N10660, N12919, N16556);
nand NAND4 (N18371, N18355, N6676, N10079, N16381);
xor XOR2 (N18372, N18357, N17151);
nand NAND3 (N18373, N18366, N9110, N1389);
xor XOR2 (N18374, N18372, N15988);
buf BUF1 (N18375, N18363);
not NOT1 (N18376, N18374);
nor NOR4 (N18377, N18331, N5553, N9457, N13184);
nand NAND2 (N18378, N18373, N14520);
nand NAND4 (N18379, N18371, N3359, N3142, N3311);
or OR2 (N18380, N18370, N15432);
nand NAND4 (N18381, N18358, N14444, N4487, N4440);
xor XOR2 (N18382, N18377, N6488);
xor XOR2 (N18383, N18369, N3212);
nor NOR4 (N18384, N18383, N6191, N6946, N18160);
nor NOR4 (N18385, N18353, N7821, N12033, N1428);
xor XOR2 (N18386, N18376, N435);
not NOT1 (N18387, N18381);
and AND3 (N18388, N18387, N12515, N2309);
or OR4 (N18389, N18368, N12, N1438, N4670);
nor NOR3 (N18390, N18384, N12455, N10882);
not NOT1 (N18391, N18386);
nand NAND3 (N18392, N18378, N9722, N17366);
or OR3 (N18393, N18389, N12138, N17607);
not NOT1 (N18394, N18375);
nand NAND2 (N18395, N18394, N16014);
not NOT1 (N18396, N18385);
or OR3 (N18397, N18391, N15200, N811);
xor XOR2 (N18398, N18380, N8606);
nor NOR2 (N18399, N18379, N3803);
nand NAND2 (N18400, N18392, N4525);
nor NOR3 (N18401, N18398, N11164, N13262);
nand NAND4 (N18402, N18393, N7994, N17450, N17363);
xor XOR2 (N18403, N18399, N12813);
not NOT1 (N18404, N18382);
nand NAND2 (N18405, N18388, N12953);
xor XOR2 (N18406, N18395, N13501);
nor NOR3 (N18407, N18396, N15588, N6470);
or OR4 (N18408, N18403, N15755, N14793, N15146);
nor NOR4 (N18409, N18405, N6047, N12300, N12065);
or OR4 (N18410, N18397, N15462, N12802, N3144);
nor NOR4 (N18411, N18402, N1542, N5487, N4753);
nand NAND4 (N18412, N18400, N17247, N11110, N8881);
not NOT1 (N18413, N18406);
xor XOR2 (N18414, N18411, N16221);
nand NAND3 (N18415, N18414, N4239, N2040);
or OR2 (N18416, N18413, N1588);
or OR4 (N18417, N18416, N2524, N155, N18327);
nand NAND4 (N18418, N18409, N607, N10089, N3201);
nand NAND4 (N18419, N18390, N15821, N635, N2872);
nor NOR2 (N18420, N18419, N12327);
not NOT1 (N18421, N18408);
xor XOR2 (N18422, N18410, N12057);
buf BUF1 (N18423, N18404);
nand NAND4 (N18424, N18420, N15168, N3850, N11760);
nor NOR4 (N18425, N18418, N7162, N4551, N15295);
buf BUF1 (N18426, N18424);
xor XOR2 (N18427, N18407, N470);
and AND3 (N18428, N18426, N10744, N13635);
and AND3 (N18429, N18421, N3373, N3274);
nor NOR2 (N18430, N18401, N10644);
and AND3 (N18431, N18417, N11515, N6009);
not NOT1 (N18432, N18431);
xor XOR2 (N18433, N18428, N17950);
or OR4 (N18434, N18412, N6353, N3052, N15808);
buf BUF1 (N18435, N18434);
nand NAND3 (N18436, N18422, N14620, N11629);
nand NAND3 (N18437, N18415, N18080, N7485);
nand NAND3 (N18438, N18423, N8269, N7676);
nor NOR2 (N18439, N18432, N15958);
nand NAND2 (N18440, N18433, N9388);
nor NOR3 (N18441, N18429, N10187, N17196);
xor XOR2 (N18442, N18435, N14915);
not NOT1 (N18443, N18439);
buf BUF1 (N18444, N18436);
nor NOR2 (N18445, N18443, N7948);
not NOT1 (N18446, N18442);
xor XOR2 (N18447, N18437, N14173);
nor NOR3 (N18448, N18445, N16411, N12763);
xor XOR2 (N18449, N18441, N4367);
or OR3 (N18450, N18447, N4020, N11516);
not NOT1 (N18451, N18450);
nor NOR3 (N18452, N18438, N12568, N888);
or OR2 (N18453, N18440, N15611);
xor XOR2 (N18454, N18444, N2147);
nand NAND3 (N18455, N18454, N3811, N1291);
nand NAND3 (N18456, N18449, N4575, N6100);
buf BUF1 (N18457, N18427);
nor NOR2 (N18458, N18457, N10528);
buf BUF1 (N18459, N18448);
nor NOR4 (N18460, N18455, N1896, N1149, N9664);
buf BUF1 (N18461, N18430);
xor XOR2 (N18462, N18425, N8309);
and AND3 (N18463, N18458, N14290, N15194);
buf BUF1 (N18464, N18453);
nand NAND3 (N18465, N18446, N16499, N16234);
not NOT1 (N18466, N18464);
or OR4 (N18467, N18461, N2236, N9001, N10763);
or OR3 (N18468, N18459, N15939, N11392);
xor XOR2 (N18469, N18466, N10897);
and AND3 (N18470, N18465, N4747, N12062);
nand NAND2 (N18471, N18460, N13442);
nor NOR4 (N18472, N18469, N4719, N10376, N5790);
xor XOR2 (N18473, N18452, N9207);
nor NOR3 (N18474, N18470, N5217, N13561);
xor XOR2 (N18475, N18462, N15656);
buf BUF1 (N18476, N18451);
nand NAND4 (N18477, N18467, N15493, N13284, N3299);
nand NAND2 (N18478, N18474, N9940);
and AND2 (N18479, N18456, N13959);
not NOT1 (N18480, N18475);
xor XOR2 (N18481, N18471, N3738);
nand NAND3 (N18482, N18478, N15920, N9861);
xor XOR2 (N18483, N18468, N7094);
xor XOR2 (N18484, N18477, N2881);
and AND3 (N18485, N18463, N1543, N7022);
buf BUF1 (N18486, N18483);
nand NAND3 (N18487, N18472, N4160, N14050);
nand NAND4 (N18488, N18473, N15186, N11447, N3451);
buf BUF1 (N18489, N18480);
buf BUF1 (N18490, N18488);
and AND4 (N18491, N18486, N3102, N7182, N871);
xor XOR2 (N18492, N18476, N11824);
xor XOR2 (N18493, N18485, N6029);
or OR2 (N18494, N18479, N16070);
buf BUF1 (N18495, N18484);
nor NOR4 (N18496, N18487, N14966, N5877, N302);
and AND3 (N18497, N18482, N3547, N14106);
and AND4 (N18498, N18495, N11687, N10562, N11025);
and AND2 (N18499, N18493, N11755);
nand NAND4 (N18500, N18498, N17331, N4223, N10311);
xor XOR2 (N18501, N18497, N9041);
buf BUF1 (N18502, N18501);
nor NOR2 (N18503, N18481, N9425);
and AND2 (N18504, N18489, N7420);
buf BUF1 (N18505, N18500);
and AND4 (N18506, N18499, N4083, N2245, N9333);
buf BUF1 (N18507, N18502);
nand NAND3 (N18508, N18504, N14890, N10721);
and AND3 (N18509, N18494, N12459, N10647);
nor NOR2 (N18510, N18507, N5105);
not NOT1 (N18511, N18509);
nor NOR2 (N18512, N18492, N7828);
xor XOR2 (N18513, N18508, N14039);
nor NOR3 (N18514, N18510, N12094, N11576);
nand NAND2 (N18515, N18503, N6206);
and AND4 (N18516, N18505, N18123, N10125, N9782);
nor NOR2 (N18517, N18516, N17404);
not NOT1 (N18518, N18490);
buf BUF1 (N18519, N18514);
or OR4 (N18520, N18506, N14409, N5002, N757);
not NOT1 (N18521, N18512);
nand NAND4 (N18522, N18521, N1620, N17366, N7398);
buf BUF1 (N18523, N18511);
nand NAND3 (N18524, N18519, N16391, N1217);
nor NOR2 (N18525, N18491, N2739);
or OR3 (N18526, N18518, N3231, N5781);
nand NAND3 (N18527, N18517, N9631, N16244);
not NOT1 (N18528, N18522);
and AND3 (N18529, N18513, N8517, N12230);
and AND3 (N18530, N18515, N7383, N1384);
buf BUF1 (N18531, N18527);
and AND4 (N18532, N18525, N17645, N188, N3905);
nor NOR3 (N18533, N18532, N546, N4124);
and AND3 (N18534, N18524, N11569, N13137);
and AND4 (N18535, N18496, N6261, N995, N7477);
xor XOR2 (N18536, N18531, N4691);
nor NOR4 (N18537, N18520, N4204, N17570, N10548);
buf BUF1 (N18538, N18523);
buf BUF1 (N18539, N18526);
nor NOR3 (N18540, N18536, N18358, N9031);
not NOT1 (N18541, N18539);
nand NAND4 (N18542, N18533, N15014, N7194, N6579);
and AND2 (N18543, N18540, N11530);
nor NOR2 (N18544, N18534, N77);
xor XOR2 (N18545, N18537, N5399);
buf BUF1 (N18546, N18530);
nor NOR4 (N18547, N18546, N12162, N17002, N13905);
nand NAND4 (N18548, N18538, N9836, N5391, N18118);
nand NAND2 (N18549, N18548, N15795);
nand NAND2 (N18550, N18535, N1754);
xor XOR2 (N18551, N18542, N12221);
not NOT1 (N18552, N18545);
and AND2 (N18553, N18550, N1842);
or OR3 (N18554, N18529, N18034, N17319);
nor NOR4 (N18555, N18549, N12007, N15909, N13189);
or OR4 (N18556, N18541, N6620, N14608, N9624);
buf BUF1 (N18557, N18544);
and AND2 (N18558, N18543, N3421);
or OR3 (N18559, N18558, N3712, N3382);
not NOT1 (N18560, N18552);
not NOT1 (N18561, N18554);
nor NOR3 (N18562, N18557, N16062, N11784);
buf BUF1 (N18563, N18559);
xor XOR2 (N18564, N18553, N8207);
or OR2 (N18565, N18562, N9325);
nor NOR4 (N18566, N18564, N16664, N11527, N1214);
nor NOR4 (N18567, N18563, N16564, N1114, N18453);
nor NOR3 (N18568, N18566, N10588, N9937);
and AND4 (N18569, N18567, N2003, N15274, N8682);
not NOT1 (N18570, N18565);
or OR3 (N18571, N18528, N117, N13770);
not NOT1 (N18572, N18556);
nand NAND2 (N18573, N18555, N5131);
nand NAND2 (N18574, N18561, N16701);
nor NOR2 (N18575, N18551, N10852);
xor XOR2 (N18576, N18575, N9392);
nor NOR2 (N18577, N18572, N8861);
nand NAND2 (N18578, N18574, N12483);
xor XOR2 (N18579, N18570, N1014);
nand NAND4 (N18580, N18560, N1405, N664, N2625);
nand NAND2 (N18581, N18578, N3527);
or OR4 (N18582, N18569, N16896, N11583, N10050);
nor NOR4 (N18583, N18573, N3118, N8702, N3231);
or OR3 (N18584, N18576, N11724, N12798);
xor XOR2 (N18585, N18584, N14876);
or OR4 (N18586, N18547, N17328, N11789, N17593);
and AND3 (N18587, N18571, N17606, N16439);
and AND2 (N18588, N18568, N17736);
not NOT1 (N18589, N18585);
and AND4 (N18590, N18579, N2994, N563, N14160);
nand NAND3 (N18591, N18589, N1241, N15502);
buf BUF1 (N18592, N18581);
nand NAND4 (N18593, N18577, N11073, N7760, N16519);
xor XOR2 (N18594, N18587, N17488);
not NOT1 (N18595, N18580);
or OR3 (N18596, N18595, N4845, N13784);
and AND2 (N18597, N18588, N964);
buf BUF1 (N18598, N18593);
nor NOR3 (N18599, N18583, N17484, N16315);
xor XOR2 (N18600, N18599, N3651);
buf BUF1 (N18601, N18598);
not NOT1 (N18602, N18590);
buf BUF1 (N18603, N18596);
or OR3 (N18604, N18600, N12168, N12998);
xor XOR2 (N18605, N18602, N10869);
nor NOR2 (N18606, N18603, N11576);
nand NAND2 (N18607, N18604, N17532);
or OR4 (N18608, N18607, N14674, N2800, N3006);
or OR3 (N18609, N18601, N4156, N4115);
xor XOR2 (N18610, N18609, N12359);
xor XOR2 (N18611, N18592, N14315);
buf BUF1 (N18612, N18610);
nand NAND3 (N18613, N18597, N16020, N6325);
nand NAND3 (N18614, N18611, N7576, N5856);
nand NAND2 (N18615, N18614, N4662);
not NOT1 (N18616, N18606);
and AND3 (N18617, N18615, N8543, N7658);
xor XOR2 (N18618, N18594, N8684);
buf BUF1 (N18619, N18613);
not NOT1 (N18620, N18586);
xor XOR2 (N18621, N18616, N18377);
buf BUF1 (N18622, N18591);
xor XOR2 (N18623, N18617, N390);
not NOT1 (N18624, N18618);
nand NAND3 (N18625, N18605, N14228, N2776);
and AND2 (N18626, N18624, N16239);
or OR2 (N18627, N18626, N13170);
not NOT1 (N18628, N18620);
nor NOR4 (N18629, N18621, N8338, N2462, N2715);
nand NAND3 (N18630, N18622, N6823, N10315);
or OR4 (N18631, N18627, N3843, N12207, N813);
xor XOR2 (N18632, N18629, N15431);
nor NOR3 (N18633, N18628, N3369, N8822);
nor NOR3 (N18634, N18625, N15950, N6890);
xor XOR2 (N18635, N18634, N342);
and AND3 (N18636, N18623, N4404, N2419);
not NOT1 (N18637, N18619);
or OR4 (N18638, N18633, N4986, N10589, N9387);
or OR2 (N18639, N18638, N473);
buf BUF1 (N18640, N18639);
nand NAND2 (N18641, N18632, N5432);
buf BUF1 (N18642, N18635);
and AND3 (N18643, N18640, N12399, N17742);
xor XOR2 (N18644, N18612, N8745);
buf BUF1 (N18645, N18636);
and AND4 (N18646, N18637, N2287, N18495, N14732);
xor XOR2 (N18647, N18646, N7700);
nor NOR2 (N18648, N18630, N3961);
nand NAND3 (N18649, N18641, N11780, N3696);
not NOT1 (N18650, N18644);
or OR2 (N18651, N18608, N16221);
nor NOR3 (N18652, N18650, N16172, N9298);
xor XOR2 (N18653, N18649, N14411);
or OR2 (N18654, N18642, N3811);
nand NAND4 (N18655, N18651, N13272, N2316, N11167);
or OR2 (N18656, N18643, N1134);
buf BUF1 (N18657, N18648);
xor XOR2 (N18658, N18657, N5890);
nand NAND2 (N18659, N18654, N5258);
or OR3 (N18660, N18645, N15970, N11653);
and AND2 (N18661, N18647, N10825);
buf BUF1 (N18662, N18656);
xor XOR2 (N18663, N18655, N12815);
or OR3 (N18664, N18653, N3000, N7815);
or OR2 (N18665, N18660, N13886);
buf BUF1 (N18666, N18661);
buf BUF1 (N18667, N18582);
buf BUF1 (N18668, N18664);
nand NAND4 (N18669, N18658, N11274, N3288, N8731);
or OR2 (N18670, N18659, N1395);
not NOT1 (N18671, N18668);
nor NOR4 (N18672, N18671, N153, N4853, N12632);
not NOT1 (N18673, N18665);
not NOT1 (N18674, N18652);
nor NOR4 (N18675, N18674, N1658, N9529, N10340);
or OR2 (N18676, N18675, N6919);
nand NAND4 (N18677, N18672, N10626, N15508, N6017);
buf BUF1 (N18678, N18669);
or OR2 (N18679, N18670, N1613);
xor XOR2 (N18680, N18631, N11558);
not NOT1 (N18681, N18677);
not NOT1 (N18682, N18663);
nand NAND2 (N18683, N18667, N3195);
xor XOR2 (N18684, N18678, N9540);
nand NAND4 (N18685, N18681, N11742, N1469, N14908);
nand NAND4 (N18686, N18676, N4406, N3074, N15044);
buf BUF1 (N18687, N18682);
xor XOR2 (N18688, N18662, N11104);
nand NAND2 (N18689, N18687, N450);
not NOT1 (N18690, N18673);
not NOT1 (N18691, N18689);
buf BUF1 (N18692, N18691);
buf BUF1 (N18693, N18679);
and AND2 (N18694, N18666, N8420);
buf BUF1 (N18695, N18692);
or OR3 (N18696, N18685, N5840, N11048);
and AND3 (N18697, N18696, N455, N9275);
or OR3 (N18698, N18683, N12054, N2124);
nand NAND3 (N18699, N18690, N1285, N13492);
buf BUF1 (N18700, N18688);
nand NAND3 (N18701, N18698, N1422, N16061);
and AND2 (N18702, N18700, N15103);
xor XOR2 (N18703, N18702, N3092);
or OR4 (N18704, N18695, N12393, N5303, N14961);
xor XOR2 (N18705, N18701, N10859);
xor XOR2 (N18706, N18704, N12844);
nor NOR4 (N18707, N18703, N17250, N13792, N18069);
xor XOR2 (N18708, N18686, N11402);
and AND2 (N18709, N18680, N4590);
or OR2 (N18710, N18705, N11074);
and AND4 (N18711, N18709, N17597, N622, N1504);
xor XOR2 (N18712, N18694, N1733);
nor NOR2 (N18713, N18693, N15717);
buf BUF1 (N18714, N18699);
buf BUF1 (N18715, N18684);
xor XOR2 (N18716, N18713, N16919);
not NOT1 (N18717, N18715);
nor NOR3 (N18718, N18706, N5887, N14554);
not NOT1 (N18719, N18710);
nand NAND4 (N18720, N18712, N10700, N4389, N16207);
or OR4 (N18721, N18720, N6038, N3500, N14344);
nand NAND3 (N18722, N18717, N13375, N2119);
and AND2 (N18723, N18708, N2957);
nand NAND4 (N18724, N18718, N17443, N13985, N85);
buf BUF1 (N18725, N18724);
xor XOR2 (N18726, N18714, N8320);
or OR3 (N18727, N18711, N6115, N3995);
nand NAND2 (N18728, N18725, N5164);
nand NAND4 (N18729, N18726, N11040, N4617, N6369);
not NOT1 (N18730, N18728);
nand NAND2 (N18731, N18730, N4822);
nor NOR3 (N18732, N18721, N12300, N16516);
nand NAND2 (N18733, N18729, N6706);
xor XOR2 (N18734, N18732, N2579);
not NOT1 (N18735, N18734);
xor XOR2 (N18736, N18733, N14339);
nor NOR3 (N18737, N18731, N6341, N6001);
or OR4 (N18738, N18736, N11202, N4160, N13477);
or OR3 (N18739, N18723, N16077, N11268);
and AND2 (N18740, N18737, N5672);
nand NAND2 (N18741, N18707, N8717);
nand NAND3 (N18742, N18697, N2365, N3400);
not NOT1 (N18743, N18740);
nor NOR3 (N18744, N18727, N11334, N16406);
buf BUF1 (N18745, N18743);
not NOT1 (N18746, N18735);
nor NOR4 (N18747, N18742, N13719, N7222, N355);
nand NAND4 (N18748, N18716, N11122, N1407, N17814);
and AND3 (N18749, N18722, N5930, N11581);
not NOT1 (N18750, N18738);
buf BUF1 (N18751, N18719);
buf BUF1 (N18752, N18748);
and AND3 (N18753, N18750, N1540, N2498);
not NOT1 (N18754, N18745);
buf BUF1 (N18755, N18749);
nor NOR4 (N18756, N18739, N10231, N9515, N5754);
nand NAND4 (N18757, N18741, N18345, N15744, N15057);
and AND4 (N18758, N18756, N16200, N18614, N12871);
nor NOR2 (N18759, N18755, N16156);
nor NOR3 (N18760, N18751, N951, N16241);
xor XOR2 (N18761, N18754, N2592);
nand NAND3 (N18762, N18757, N10990, N12044);
nor NOR4 (N18763, N18747, N2248, N229, N11875);
not NOT1 (N18764, N18752);
xor XOR2 (N18765, N18761, N8089);
and AND3 (N18766, N18762, N5717, N11964);
nand NAND3 (N18767, N18765, N18133, N12704);
nand NAND2 (N18768, N18760, N14743);
buf BUF1 (N18769, N18767);
buf BUF1 (N18770, N18769);
nand NAND3 (N18771, N18763, N1050, N11236);
nor NOR2 (N18772, N18744, N13484);
not NOT1 (N18773, N18764);
and AND3 (N18774, N18753, N13485, N7977);
buf BUF1 (N18775, N18766);
and AND2 (N18776, N18758, N17027);
nand NAND2 (N18777, N18759, N16620);
nand NAND3 (N18778, N18777, N8527, N5178);
not NOT1 (N18779, N18768);
xor XOR2 (N18780, N18774, N16848);
not NOT1 (N18781, N18770);
buf BUF1 (N18782, N18772);
xor XOR2 (N18783, N18776, N9086);
not NOT1 (N18784, N18779);
not NOT1 (N18785, N18780);
nand NAND3 (N18786, N18785, N3464, N15947);
nor NOR2 (N18787, N18773, N13790);
nor NOR3 (N18788, N18784, N14934, N365);
not NOT1 (N18789, N18771);
not NOT1 (N18790, N18746);
nand NAND2 (N18791, N18783, N18523);
nor NOR4 (N18792, N18775, N10638, N11204, N2995);
not NOT1 (N18793, N18782);
and AND2 (N18794, N18786, N895);
or OR3 (N18795, N18787, N17795, N17675);
buf BUF1 (N18796, N18789);
not NOT1 (N18797, N18794);
xor XOR2 (N18798, N18795, N17712);
nor NOR3 (N18799, N18792, N6689, N3199);
and AND4 (N18800, N18781, N4947, N16130, N14069);
nor NOR2 (N18801, N18791, N17327);
and AND2 (N18802, N18788, N8112);
not NOT1 (N18803, N18797);
or OR4 (N18804, N18799, N16485, N9023, N12585);
nand NAND4 (N18805, N18778, N954, N10891, N18093);
and AND4 (N18806, N18802, N16594, N1777, N8036);
and AND4 (N18807, N18800, N9034, N8208, N18618);
and AND3 (N18808, N18804, N7623, N16640);
xor XOR2 (N18809, N18803, N15272);
and AND2 (N18810, N18798, N17601);
nor NOR2 (N18811, N18808, N7245);
buf BUF1 (N18812, N18809);
xor XOR2 (N18813, N18810, N9759);
not NOT1 (N18814, N18806);
or OR4 (N18815, N18796, N14446, N16697, N16538);
not NOT1 (N18816, N18811);
nand NAND2 (N18817, N18790, N9019);
nand NAND2 (N18818, N18815, N11033);
buf BUF1 (N18819, N18812);
buf BUF1 (N18820, N18801);
nor NOR3 (N18821, N18819, N15167, N4953);
buf BUF1 (N18822, N18820);
nand NAND3 (N18823, N18816, N7338, N17760);
not NOT1 (N18824, N18814);
not NOT1 (N18825, N18821);
xor XOR2 (N18826, N18817, N1687);
buf BUF1 (N18827, N18818);
buf BUF1 (N18828, N18824);
nand NAND4 (N18829, N18823, N15382, N6723, N9200);
nor NOR2 (N18830, N18813, N9949);
xor XOR2 (N18831, N18826, N90);
or OR4 (N18832, N18830, N2472, N8279, N16709);
nor NOR2 (N18833, N18827, N17760);
buf BUF1 (N18834, N18807);
buf BUF1 (N18835, N18833);
buf BUF1 (N18836, N18793);
not NOT1 (N18837, N18825);
or OR4 (N18838, N18831, N2336, N5015, N1876);
nand NAND4 (N18839, N18829, N9079, N12095, N8612);
xor XOR2 (N18840, N18834, N8157);
nand NAND4 (N18841, N18805, N15701, N13464, N4425);
or OR3 (N18842, N18832, N3091, N3266);
xor XOR2 (N18843, N18841, N13265);
nand NAND2 (N18844, N18835, N10296);
not NOT1 (N18845, N18840);
and AND4 (N18846, N18838, N4768, N8857, N9841);
or OR4 (N18847, N18839, N14767, N11062, N5195);
or OR4 (N18848, N18822, N9604, N16930, N4325);
and AND3 (N18849, N18844, N1538, N18117);
buf BUF1 (N18850, N18843);
not NOT1 (N18851, N18849);
and AND3 (N18852, N18850, N16814, N5764);
nand NAND2 (N18853, N18847, N4595);
nor NOR2 (N18854, N18842, N6525);
nor NOR2 (N18855, N18852, N2052);
and AND3 (N18856, N18836, N17431, N6859);
nand NAND4 (N18857, N18845, N12472, N5181, N12254);
nand NAND4 (N18858, N18848, N12574, N312, N6485);
nand NAND4 (N18859, N18851, N5034, N15875, N18645);
nor NOR4 (N18860, N18854, N983, N15168, N8485);
buf BUF1 (N18861, N18856);
and AND4 (N18862, N18853, N3671, N14768, N7791);
buf BUF1 (N18863, N18837);
or OR2 (N18864, N18846, N12465);
nor NOR2 (N18865, N18828, N13782);
xor XOR2 (N18866, N18858, N7107);
buf BUF1 (N18867, N18864);
xor XOR2 (N18868, N18855, N18214);
xor XOR2 (N18869, N18867, N7733);
buf BUF1 (N18870, N18860);
or OR2 (N18871, N18859, N9051);
or OR4 (N18872, N18862, N9902, N12889, N1174);
or OR4 (N18873, N18863, N18659, N6305, N10698);
or OR4 (N18874, N18857, N5242, N5949, N3069);
and AND3 (N18875, N18870, N4572, N10107);
and AND4 (N18876, N18872, N16419, N16175, N3615);
nand NAND4 (N18877, N18876, N16848, N12042, N3171);
and AND4 (N18878, N18877, N11391, N9039, N6223);
and AND4 (N18879, N18873, N14317, N384, N11270);
not NOT1 (N18880, N18871);
nand NAND3 (N18881, N18861, N5840, N7601);
xor XOR2 (N18882, N18880, N10145);
not NOT1 (N18883, N18882);
xor XOR2 (N18884, N18869, N13403);
or OR4 (N18885, N18875, N7377, N9833, N10275);
nand NAND3 (N18886, N18874, N6347, N15955);
nor NOR4 (N18887, N18879, N7413, N18021, N17765);
buf BUF1 (N18888, N18866);
or OR2 (N18889, N18878, N3557);
nor NOR3 (N18890, N18888, N17987, N5751);
buf BUF1 (N18891, N18881);
not NOT1 (N18892, N18885);
and AND3 (N18893, N18889, N7525, N2071);
or OR3 (N18894, N18868, N4929, N9577);
nand NAND3 (N18895, N18884, N8048, N17510);
nor NOR4 (N18896, N18891, N2573, N1471, N14410);
xor XOR2 (N18897, N18883, N13905);
nand NAND2 (N18898, N18892, N13090);
buf BUF1 (N18899, N18886);
or OR4 (N18900, N18893, N5397, N9199, N9307);
and AND3 (N18901, N18890, N16880, N13846);
nand NAND2 (N18902, N18897, N18545);
nor NOR4 (N18903, N18900, N13364, N12338, N5122);
or OR3 (N18904, N18894, N18654, N6572);
buf BUF1 (N18905, N18896);
not NOT1 (N18906, N18899);
not NOT1 (N18907, N18905);
nor NOR2 (N18908, N18902, N2899);
buf BUF1 (N18909, N18898);
and AND4 (N18910, N18865, N203, N12152, N4172);
xor XOR2 (N18911, N18908, N1766);
and AND4 (N18912, N18911, N9566, N14791, N459);
xor XOR2 (N18913, N18912, N11258);
and AND3 (N18914, N18909, N7715, N14335);
and AND2 (N18915, N18906, N5630);
xor XOR2 (N18916, N18904, N7833);
xor XOR2 (N18917, N18915, N9128);
not NOT1 (N18918, N18914);
xor XOR2 (N18919, N18907, N12382);
buf BUF1 (N18920, N18887);
and AND2 (N18921, N18895, N8566);
not NOT1 (N18922, N18913);
or OR3 (N18923, N18917, N2545, N6622);
nor NOR3 (N18924, N18919, N9396, N17921);
nor NOR3 (N18925, N18916, N12947, N8248);
not NOT1 (N18926, N18925);
not NOT1 (N18927, N18924);
or OR4 (N18928, N18922, N3942, N18420, N11931);
nand NAND4 (N18929, N18901, N6389, N3616, N17397);
nand NAND3 (N18930, N18918, N16228, N14927);
or OR3 (N18931, N18921, N16240, N16230);
or OR3 (N18932, N18903, N8393, N10934);
nor NOR2 (N18933, N18928, N14539);
or OR2 (N18934, N18931, N13971);
or OR3 (N18935, N18920, N12260, N18439);
nor NOR3 (N18936, N18935, N3916, N17216);
and AND2 (N18937, N18927, N234);
xor XOR2 (N18938, N18929, N14889);
not NOT1 (N18939, N18937);
or OR4 (N18940, N18930, N14642, N4850, N6059);
nor NOR2 (N18941, N18932, N16878);
nand NAND4 (N18942, N18936, N5823, N15665, N15288);
nor NOR4 (N18943, N18910, N7839, N608, N10397);
buf BUF1 (N18944, N18940);
buf BUF1 (N18945, N18941);
buf BUF1 (N18946, N18938);
xor XOR2 (N18947, N18942, N5545);
nand NAND4 (N18948, N18943, N1426, N6760, N3393);
not NOT1 (N18949, N18923);
not NOT1 (N18950, N18939);
and AND4 (N18951, N18934, N18577, N16373, N7141);
xor XOR2 (N18952, N18948, N9441);
nor NOR2 (N18953, N18946, N1497);
buf BUF1 (N18954, N18933);
xor XOR2 (N18955, N18926, N3071);
and AND3 (N18956, N18952, N8586, N7665);
or OR4 (N18957, N18955, N15678, N10371, N2460);
and AND4 (N18958, N18944, N1826, N5123, N14470);
buf BUF1 (N18959, N18951);
nor NOR3 (N18960, N18957, N3826, N9241);
xor XOR2 (N18961, N18950, N16405);
or OR2 (N18962, N18949, N4865);
xor XOR2 (N18963, N18953, N9952);
xor XOR2 (N18964, N18945, N11849);
nor NOR4 (N18965, N18954, N11935, N16274, N2118);
buf BUF1 (N18966, N18962);
or OR2 (N18967, N18960, N461);
not NOT1 (N18968, N18966);
not NOT1 (N18969, N18956);
nand NAND4 (N18970, N18969, N15914, N3138, N4525);
or OR2 (N18971, N18964, N14726);
nand NAND4 (N18972, N18961, N11451, N5113, N16757);
nor NOR3 (N18973, N18959, N6940, N7957);
or OR2 (N18974, N18963, N12000);
nor NOR2 (N18975, N18968, N15855);
or OR4 (N18976, N18971, N15030, N4595, N7372);
nand NAND3 (N18977, N18947, N10215, N16767);
or OR2 (N18978, N18976, N8848);
or OR2 (N18979, N18977, N9041);
and AND4 (N18980, N18979, N8921, N15520, N15924);
nor NOR3 (N18981, N18974, N10028, N18436);
or OR2 (N18982, N18965, N8558);
nand NAND2 (N18983, N18973, N620);
nor NOR4 (N18984, N18967, N6408, N262, N9701);
xor XOR2 (N18985, N18972, N11898);
or OR4 (N18986, N18982, N18223, N16841, N17912);
buf BUF1 (N18987, N18970);
nor NOR3 (N18988, N18983, N11645, N10747);
not NOT1 (N18989, N18985);
nor NOR2 (N18990, N18984, N1496);
nand NAND3 (N18991, N18989, N11187, N6281);
nand NAND3 (N18992, N18980, N2924, N2697);
nor NOR3 (N18993, N18981, N11959, N7305);
not NOT1 (N18994, N18990);
xor XOR2 (N18995, N18992, N1776);
buf BUF1 (N18996, N18988);
not NOT1 (N18997, N18991);
buf BUF1 (N18998, N18994);
buf BUF1 (N18999, N18997);
or OR3 (N19000, N18986, N3575, N12438);
buf BUF1 (N19001, N18958);
xor XOR2 (N19002, N19001, N6628);
not NOT1 (N19003, N18999);
buf BUF1 (N19004, N18995);
xor XOR2 (N19005, N19003, N1025);
and AND4 (N19006, N19002, N16214, N15995, N16142);
xor XOR2 (N19007, N18998, N7724);
nor NOR2 (N19008, N18996, N18399);
or OR3 (N19009, N19008, N6694, N16137);
buf BUF1 (N19010, N19009);
not NOT1 (N19011, N19004);
and AND2 (N19012, N18978, N14264);
nor NOR4 (N19013, N19010, N15488, N4898, N10018);
nor NOR3 (N19014, N19013, N5971, N9589);
and AND2 (N19015, N19011, N7509);
xor XOR2 (N19016, N19000, N2142);
or OR2 (N19017, N19012, N12945);
xor XOR2 (N19018, N18993, N9295);
nor NOR4 (N19019, N19006, N15494, N7740, N8706);
or OR3 (N19020, N19007, N10338, N10827);
buf BUF1 (N19021, N19020);
nand NAND3 (N19022, N19015, N16197, N12488);
xor XOR2 (N19023, N19017, N15250);
xor XOR2 (N19024, N19022, N14929);
not NOT1 (N19025, N19023);
not NOT1 (N19026, N19024);
buf BUF1 (N19027, N19021);
buf BUF1 (N19028, N18975);
nor NOR2 (N19029, N19027, N5356);
nand NAND3 (N19030, N19005, N8180, N15090);
buf BUF1 (N19031, N19025);
nor NOR4 (N19032, N19026, N6598, N14553, N9700);
nand NAND4 (N19033, N19028, N11331, N1757, N6762);
not NOT1 (N19034, N19018);
not NOT1 (N19035, N19016);
nor NOR3 (N19036, N19035, N9662, N8605);
or OR4 (N19037, N19029, N15066, N10643, N16937);
buf BUF1 (N19038, N19031);
xor XOR2 (N19039, N19019, N1322);
and AND2 (N19040, N19039, N924);
nand NAND3 (N19041, N18987, N15189, N6070);
nand NAND2 (N19042, N19037, N15395);
and AND3 (N19043, N19030, N14158, N3357);
xor XOR2 (N19044, N19038, N10450);
not NOT1 (N19045, N19041);
not NOT1 (N19046, N19045);
or OR2 (N19047, N19036, N2538);
or OR3 (N19048, N19043, N4928, N18071);
not NOT1 (N19049, N19046);
and AND2 (N19050, N19014, N17146);
buf BUF1 (N19051, N19049);
nand NAND3 (N19052, N19033, N2090, N13259);
not NOT1 (N19053, N19032);
nand NAND2 (N19054, N19052, N15917);
not NOT1 (N19055, N19042);
nor NOR3 (N19056, N19044, N7886, N564);
nor NOR2 (N19057, N19056, N3977);
xor XOR2 (N19058, N19053, N8081);
and AND2 (N19059, N19040, N4460);
nor NOR3 (N19060, N19057, N11711, N4605);
buf BUF1 (N19061, N19055);
xor XOR2 (N19062, N19059, N13863);
not NOT1 (N19063, N19061);
not NOT1 (N19064, N19050);
or OR4 (N19065, N19054, N12274, N13220, N16064);
xor XOR2 (N19066, N19060, N15386);
nor NOR3 (N19067, N19058, N4582, N16303);
not NOT1 (N19068, N19034);
buf BUF1 (N19069, N19067);
buf BUF1 (N19070, N19064);
not NOT1 (N19071, N19051);
xor XOR2 (N19072, N19070, N14522);
or OR3 (N19073, N19063, N7950, N18159);
or OR3 (N19074, N19062, N12978, N9934);
xor XOR2 (N19075, N19071, N9568);
and AND3 (N19076, N19048, N12205, N5932);
xor XOR2 (N19077, N19074, N8680);
or OR3 (N19078, N19077, N13568, N8461);
nand NAND3 (N19079, N19078, N13135, N11760);
or OR2 (N19080, N19068, N152);
xor XOR2 (N19081, N19065, N1641);
xor XOR2 (N19082, N19047, N3130);
buf BUF1 (N19083, N19069);
and AND3 (N19084, N19079, N17790, N5623);
not NOT1 (N19085, N19072);
or OR4 (N19086, N19083, N3844, N8987, N17363);
not NOT1 (N19087, N19076);
buf BUF1 (N19088, N19081);
nand NAND4 (N19089, N19084, N12222, N1114, N2142);
nand NAND4 (N19090, N19086, N1017, N11788, N3338);
and AND3 (N19091, N19085, N15139, N16982);
and AND4 (N19092, N19066, N15495, N7998, N9979);
and AND3 (N19093, N19091, N18533, N2637);
xor XOR2 (N19094, N19093, N14163);
or OR2 (N19095, N19087, N16851);
buf BUF1 (N19096, N19089);
xor XOR2 (N19097, N19090, N1386);
nand NAND4 (N19098, N19096, N7729, N17211, N15547);
not NOT1 (N19099, N19075);
or OR3 (N19100, N19095, N7998, N250);
nand NAND4 (N19101, N19073, N16505, N9455, N7901);
nand NAND3 (N19102, N19094, N7566, N8666);
not NOT1 (N19103, N19102);
nand NAND4 (N19104, N19099, N18784, N8348, N12679);
buf BUF1 (N19105, N19097);
buf BUF1 (N19106, N19088);
or OR4 (N19107, N19103, N10008, N2411, N167);
xor XOR2 (N19108, N19092, N16979);
buf BUF1 (N19109, N19100);
nor NOR2 (N19110, N19080, N2766);
not NOT1 (N19111, N19105);
buf BUF1 (N19112, N19107);
nand NAND2 (N19113, N19109, N5660);
buf BUF1 (N19114, N19082);
not NOT1 (N19115, N19098);
and AND4 (N19116, N19115, N14561, N9286, N2060);
nand NAND4 (N19117, N19101, N1550, N9942, N2627);
xor XOR2 (N19118, N19112, N13007);
and AND4 (N19119, N19110, N8012, N1236, N7172);
or OR4 (N19120, N19119, N14218, N8933, N7573);
xor XOR2 (N19121, N19113, N16445);
and AND3 (N19122, N19114, N10865, N7051);
xor XOR2 (N19123, N19106, N5662);
and AND2 (N19124, N19104, N11919);
nand NAND4 (N19125, N19122, N10811, N12003, N8674);
or OR4 (N19126, N19120, N17962, N9412, N13847);
nand NAND4 (N19127, N19126, N18892, N373, N2471);
nand NAND2 (N19128, N19123, N14210);
xor XOR2 (N19129, N19116, N480);
buf BUF1 (N19130, N19108);
xor XOR2 (N19131, N19121, N6954);
nor NOR2 (N19132, N19130, N8690);
xor XOR2 (N19133, N19131, N18682);
nor NOR3 (N19134, N19111, N16842, N4651);
buf BUF1 (N19135, N19117);
nor NOR2 (N19136, N19129, N14049);
and AND4 (N19137, N19133, N1239, N277, N14304);
xor XOR2 (N19138, N19125, N12396);
xor XOR2 (N19139, N19127, N2098);
buf BUF1 (N19140, N19135);
xor XOR2 (N19141, N19140, N3037);
xor XOR2 (N19142, N19134, N9944);
not NOT1 (N19143, N19128);
xor XOR2 (N19144, N19142, N15973);
not NOT1 (N19145, N19139);
and AND3 (N19146, N19136, N2489, N5763);
or OR4 (N19147, N19141, N3834, N10227, N9422);
nand NAND2 (N19148, N19132, N15202);
or OR3 (N19149, N19137, N14540, N5401);
or OR4 (N19150, N19118, N898, N8575, N1388);
or OR4 (N19151, N19150, N3268, N13075, N1361);
and AND2 (N19152, N19147, N251);
xor XOR2 (N19153, N19124, N16465);
not NOT1 (N19154, N19146);
or OR4 (N19155, N19153, N1204, N4458, N8459);
xor XOR2 (N19156, N19149, N798);
xor XOR2 (N19157, N19145, N13393);
nand NAND2 (N19158, N19154, N5562);
nor NOR2 (N19159, N19155, N18360);
buf BUF1 (N19160, N19152);
and AND4 (N19161, N19148, N6925, N9512, N13243);
or OR3 (N19162, N19158, N5598, N10919);
buf BUF1 (N19163, N19157);
and AND4 (N19164, N19162, N4387, N18373, N17566);
buf BUF1 (N19165, N19161);
buf BUF1 (N19166, N19156);
nand NAND4 (N19167, N19143, N8598, N18731, N1356);
buf BUF1 (N19168, N19167);
nand NAND2 (N19169, N19166, N2590);
nand NAND2 (N19170, N19168, N2447);
or OR2 (N19171, N19163, N7022);
nand NAND4 (N19172, N19144, N4199, N14647, N14603);
xor XOR2 (N19173, N19160, N17386);
and AND2 (N19174, N19169, N2559);
and AND4 (N19175, N19164, N17434, N3571, N16858);
buf BUF1 (N19176, N19151);
or OR4 (N19177, N19176, N16834, N17777, N12522);
xor XOR2 (N19178, N19138, N3994);
or OR4 (N19179, N19175, N8204, N2361, N15067);
and AND3 (N19180, N19170, N13867, N13687);
not NOT1 (N19181, N19165);
or OR2 (N19182, N19178, N8726);
buf BUF1 (N19183, N19181);
or OR3 (N19184, N19179, N19071, N5400);
nand NAND4 (N19185, N19173, N18439, N8506, N10708);
buf BUF1 (N19186, N19184);
nand NAND4 (N19187, N19180, N9980, N9469, N18982);
xor XOR2 (N19188, N19182, N11543);
xor XOR2 (N19189, N19188, N15133);
not NOT1 (N19190, N19172);
buf BUF1 (N19191, N19189);
and AND3 (N19192, N19187, N15586, N16852);
nor NOR3 (N19193, N19177, N3399, N13744);
and AND4 (N19194, N19192, N8367, N3842, N18272);
not NOT1 (N19195, N19190);
or OR2 (N19196, N19186, N11300);
not NOT1 (N19197, N19174);
not NOT1 (N19198, N19194);
xor XOR2 (N19199, N19195, N7310);
buf BUF1 (N19200, N19199);
or OR4 (N19201, N19183, N4944, N12427, N8170);
nand NAND3 (N19202, N19197, N12110, N1627);
and AND4 (N19203, N19185, N7234, N13740, N11030);
or OR2 (N19204, N19201, N11050);
or OR4 (N19205, N19193, N4096, N7475, N17847);
buf BUF1 (N19206, N19191);
not NOT1 (N19207, N19159);
nor NOR3 (N19208, N19203, N6205, N6614);
xor XOR2 (N19209, N19204, N8565);
or OR3 (N19210, N19209, N9862, N8937);
nor NOR3 (N19211, N19198, N4954, N10892);
xor XOR2 (N19212, N19211, N4142);
not NOT1 (N19213, N19196);
buf BUF1 (N19214, N19206);
not NOT1 (N19215, N19208);
or OR2 (N19216, N19210, N4169);
nor NOR3 (N19217, N19202, N18316, N10454);
xor XOR2 (N19218, N19205, N15327);
nand NAND2 (N19219, N19200, N16235);
not NOT1 (N19220, N19207);
or OR4 (N19221, N19212, N7242, N3834, N10118);
xor XOR2 (N19222, N19221, N2856);
not NOT1 (N19223, N19171);
buf BUF1 (N19224, N19215);
xor XOR2 (N19225, N19218, N5687);
nor NOR4 (N19226, N19223, N8298, N2073, N14617);
and AND4 (N19227, N19217, N8167, N3408, N18489);
or OR2 (N19228, N19224, N13018);
xor XOR2 (N19229, N19214, N15085);
xor XOR2 (N19230, N19225, N15940);
and AND2 (N19231, N19230, N10694);
nor NOR2 (N19232, N19226, N15553);
or OR3 (N19233, N19232, N7564, N12030);
not NOT1 (N19234, N19229);
nand NAND4 (N19235, N19227, N19213, N1411, N19208);
buf BUF1 (N19236, N2792);
nand NAND4 (N19237, N19220, N7753, N18494, N12403);
xor XOR2 (N19238, N19219, N15443);
or OR4 (N19239, N19238, N3963, N17244, N11850);
nand NAND2 (N19240, N19233, N770);
or OR4 (N19241, N19240, N15315, N18134, N13699);
not NOT1 (N19242, N19231);
buf BUF1 (N19243, N19216);
not NOT1 (N19244, N19243);
buf BUF1 (N19245, N19222);
nor NOR2 (N19246, N19236, N3107);
or OR4 (N19247, N19237, N18361, N14506, N4497);
nand NAND2 (N19248, N19235, N2779);
or OR3 (N19249, N19242, N5714, N16266);
and AND2 (N19250, N19247, N16834);
xor XOR2 (N19251, N19248, N120);
buf BUF1 (N19252, N19250);
not NOT1 (N19253, N19241);
nand NAND2 (N19254, N19246, N16705);
or OR2 (N19255, N19249, N1712);
or OR2 (N19256, N19255, N9571);
and AND2 (N19257, N19245, N4942);
buf BUF1 (N19258, N19234);
nor NOR2 (N19259, N19251, N15965);
and AND4 (N19260, N19253, N18087, N17032, N1830);
not NOT1 (N19261, N19257);
nor NOR2 (N19262, N19261, N9481);
xor XOR2 (N19263, N19262, N18500);
and AND3 (N19264, N19252, N8864, N14736);
not NOT1 (N19265, N19239);
xor XOR2 (N19266, N19264, N1879);
not NOT1 (N19267, N19265);
buf BUF1 (N19268, N19263);
and AND3 (N19269, N19228, N7333, N16246);
buf BUF1 (N19270, N19268);
buf BUF1 (N19271, N19260);
buf BUF1 (N19272, N19254);
nor NOR4 (N19273, N19269, N5651, N3973, N16458);
xor XOR2 (N19274, N19266, N3277);
xor XOR2 (N19275, N19259, N173);
nand NAND2 (N19276, N19272, N15678);
nor NOR3 (N19277, N19244, N7232, N18333);
and AND3 (N19278, N19274, N1011, N17139);
not NOT1 (N19279, N19273);
and AND4 (N19280, N19256, N17444, N17622, N15727);
nand NAND2 (N19281, N19267, N267);
buf BUF1 (N19282, N19276);
nand NAND2 (N19283, N19258, N18799);
nor NOR3 (N19284, N19279, N7102, N15248);
nand NAND4 (N19285, N19277, N17307, N8353, N334);
or OR3 (N19286, N19280, N11933, N6993);
nor NOR4 (N19287, N19271, N12722, N18703, N2704);
and AND3 (N19288, N19287, N14987, N14174);
buf BUF1 (N19289, N19275);
nor NOR4 (N19290, N19284, N16421, N10389, N15096);
nor NOR3 (N19291, N19278, N16134, N5087);
not NOT1 (N19292, N19285);
buf BUF1 (N19293, N19292);
xor XOR2 (N19294, N19288, N1927);
nor NOR3 (N19295, N19281, N5186, N16005);
or OR4 (N19296, N19286, N15600, N8332, N10670);
xor XOR2 (N19297, N19270, N952);
or OR2 (N19298, N19295, N9514);
and AND4 (N19299, N19291, N12403, N8866, N8415);
nor NOR4 (N19300, N19282, N12774, N3177, N10225);
xor XOR2 (N19301, N19299, N8710);
nor NOR4 (N19302, N19301, N4869, N10529, N2254);
xor XOR2 (N19303, N19298, N12920);
nand NAND4 (N19304, N19289, N12544, N10531, N6958);
or OR4 (N19305, N19303, N15101, N1657, N3222);
buf BUF1 (N19306, N19290);
xor XOR2 (N19307, N19283, N2331);
xor XOR2 (N19308, N19306, N9704);
or OR4 (N19309, N19300, N12401, N17041, N5246);
buf BUF1 (N19310, N19293);
or OR2 (N19311, N19309, N6851);
and AND2 (N19312, N19307, N4511);
not NOT1 (N19313, N19304);
or OR4 (N19314, N19310, N2925, N15750, N3611);
nand NAND2 (N19315, N19297, N613);
or OR3 (N19316, N19315, N12210, N11889);
xor XOR2 (N19317, N19308, N14195);
nor NOR3 (N19318, N19296, N2036, N105);
or OR2 (N19319, N19317, N478);
nand NAND4 (N19320, N19312, N6389, N11938, N7047);
nand NAND2 (N19321, N19313, N4671);
buf BUF1 (N19322, N19314);
nor NOR2 (N19323, N19305, N12170);
xor XOR2 (N19324, N19323, N13224);
not NOT1 (N19325, N19319);
nand NAND4 (N19326, N19324, N13771, N324, N9082);
xor XOR2 (N19327, N19321, N2838);
xor XOR2 (N19328, N19322, N844);
xor XOR2 (N19329, N19325, N15727);
xor XOR2 (N19330, N19318, N10939);
buf BUF1 (N19331, N19326);
or OR2 (N19332, N19316, N18648);
nand NAND4 (N19333, N19330, N8159, N12171, N5581);
and AND3 (N19334, N19332, N7520, N12444);
or OR4 (N19335, N19328, N1749, N12770, N11188);
xor XOR2 (N19336, N19334, N17038);
or OR2 (N19337, N19311, N911);
and AND4 (N19338, N19336, N1277, N3277, N17080);
nand NAND3 (N19339, N19302, N2735, N5007);
and AND2 (N19340, N19338, N9416);
or OR3 (N19341, N19320, N13726, N6980);
not NOT1 (N19342, N19329);
and AND4 (N19343, N19327, N7768, N13542, N10283);
nand NAND4 (N19344, N19337, N10818, N14889, N11200);
buf BUF1 (N19345, N19335);
nor NOR2 (N19346, N19343, N9827);
nand NAND4 (N19347, N19339, N16336, N14140, N14555);
nor NOR2 (N19348, N19344, N7418);
nand NAND4 (N19349, N19345, N14102, N9699, N3311);
or OR4 (N19350, N19349, N6859, N8464, N12240);
or OR2 (N19351, N19340, N13989);
nand NAND2 (N19352, N19348, N11162);
and AND2 (N19353, N19331, N7042);
nand NAND3 (N19354, N19346, N19199, N12608);
buf BUF1 (N19355, N19341);
nor NOR4 (N19356, N19342, N9250, N7536, N2506);
buf BUF1 (N19357, N19350);
nor NOR2 (N19358, N19353, N8138);
nor NOR4 (N19359, N19351, N868, N881, N4447);
xor XOR2 (N19360, N19356, N2504);
and AND2 (N19361, N19354, N9905);
nand NAND3 (N19362, N19361, N8488, N12025);
and AND2 (N19363, N19362, N12092);
nand NAND4 (N19364, N19347, N483, N11243, N11838);
nand NAND4 (N19365, N19357, N17662, N18475, N4253);
nor NOR3 (N19366, N19359, N3365, N8165);
and AND4 (N19367, N19364, N14781, N10776, N5068);
buf BUF1 (N19368, N19360);
xor XOR2 (N19369, N19365, N12561);
xor XOR2 (N19370, N19368, N6681);
nor NOR3 (N19371, N19370, N8597, N19173);
not NOT1 (N19372, N19366);
and AND3 (N19373, N19363, N8525, N17489);
buf BUF1 (N19374, N19333);
not NOT1 (N19375, N19369);
nand NAND2 (N19376, N19375, N12290);
and AND2 (N19377, N19371, N11443);
and AND2 (N19378, N19374, N13201);
or OR3 (N19379, N19372, N1451, N2946);
nand NAND4 (N19380, N19379, N7544, N7238, N15614);
nand NAND3 (N19381, N19358, N9491, N15419);
not NOT1 (N19382, N19355);
and AND2 (N19383, N19381, N16334);
nand NAND3 (N19384, N19352, N14639, N3779);
nor NOR3 (N19385, N19377, N4542, N130);
and AND4 (N19386, N19378, N16800, N672, N536);
xor XOR2 (N19387, N19383, N8961);
or OR3 (N19388, N19387, N7236, N7657);
nand NAND4 (N19389, N19384, N4922, N7193, N6182);
nor NOR3 (N19390, N19294, N2376, N6070);
xor XOR2 (N19391, N19385, N5670);
and AND3 (N19392, N19391, N2133, N5788);
nand NAND2 (N19393, N19388, N2379);
nand NAND4 (N19394, N19373, N15335, N17415, N1468);
xor XOR2 (N19395, N19376, N17820);
nor NOR3 (N19396, N19382, N7310, N5559);
or OR2 (N19397, N19392, N17121);
nand NAND3 (N19398, N19396, N11666, N12441);
nor NOR3 (N19399, N19380, N7333, N18798);
nor NOR3 (N19400, N19389, N8104, N8772);
nor NOR4 (N19401, N19400, N14397, N4337, N14945);
nand NAND2 (N19402, N19393, N3342);
nor NOR4 (N19403, N19397, N14225, N2250, N14891);
xor XOR2 (N19404, N19401, N14734);
nor NOR2 (N19405, N19399, N16149);
buf BUF1 (N19406, N19390);
xor XOR2 (N19407, N19405, N14963);
not NOT1 (N19408, N19398);
and AND4 (N19409, N19367, N768, N12042, N11410);
nor NOR2 (N19410, N19404, N2796);
xor XOR2 (N19411, N19402, N16310);
nand NAND2 (N19412, N19408, N3352);
and AND2 (N19413, N19409, N17691);
or OR2 (N19414, N19413, N927);
nor NOR2 (N19415, N19386, N6552);
xor XOR2 (N19416, N19406, N10273);
or OR2 (N19417, N19414, N2156);
not NOT1 (N19418, N19395);
nand NAND2 (N19419, N19407, N9667);
nor NOR4 (N19420, N19415, N10261, N3483, N7679);
nor NOR2 (N19421, N19394, N1364);
buf BUF1 (N19422, N19418);
buf BUF1 (N19423, N19419);
and AND2 (N19424, N19412, N10940);
nand NAND4 (N19425, N19416, N906, N14230, N19398);
xor XOR2 (N19426, N19422, N18769);
buf BUF1 (N19427, N19421);
and AND4 (N19428, N19424, N3895, N15804, N16366);
xor XOR2 (N19429, N19428, N19329);
nor NOR2 (N19430, N19411, N17672);
nor NOR2 (N19431, N19403, N3667);
nor NOR4 (N19432, N19423, N8778, N12014, N5633);
not NOT1 (N19433, N19432);
nor NOR2 (N19434, N19430, N1062);
xor XOR2 (N19435, N19426, N11728);
nor NOR2 (N19436, N19427, N4862);
nand NAND4 (N19437, N19425, N10848, N17812, N4073);
or OR2 (N19438, N19417, N11812);
not NOT1 (N19439, N19438);
nor NOR3 (N19440, N19437, N8677, N7566);
or OR3 (N19441, N19435, N14379, N8366);
nand NAND2 (N19442, N19434, N12504);
nor NOR4 (N19443, N19410, N3046, N4524, N3859);
or OR2 (N19444, N19433, N8572);
buf BUF1 (N19445, N19440);
and AND3 (N19446, N19420, N17419, N13900);
buf BUF1 (N19447, N19439);
buf BUF1 (N19448, N19447);
not NOT1 (N19449, N19436);
nand NAND4 (N19450, N19443, N13470, N11627, N18289);
nor NOR3 (N19451, N19446, N5829, N6362);
not NOT1 (N19452, N19445);
xor XOR2 (N19453, N19444, N5155);
nand NAND2 (N19454, N19453, N16543);
nand NAND2 (N19455, N19454, N3444);
xor XOR2 (N19456, N19429, N8858);
and AND4 (N19457, N19448, N4002, N9406, N18240);
nor NOR2 (N19458, N19451, N2699);
not NOT1 (N19459, N19441);
or OR2 (N19460, N19455, N9956);
or OR2 (N19461, N19442, N4894);
nand NAND2 (N19462, N19452, N4585);
not NOT1 (N19463, N19459);
xor XOR2 (N19464, N19450, N19058);
nor NOR3 (N19465, N19431, N9925, N3505);
not NOT1 (N19466, N19461);
nor NOR2 (N19467, N19464, N10457);
not NOT1 (N19468, N19458);
or OR4 (N19469, N19460, N9445, N2102, N3076);
and AND3 (N19470, N19463, N14324, N11395);
nor NOR2 (N19471, N19462, N14912);
buf BUF1 (N19472, N19457);
and AND2 (N19473, N19472, N418);
buf BUF1 (N19474, N19473);
or OR3 (N19475, N19467, N12419, N9752);
nand NAND3 (N19476, N19471, N19076, N13481);
and AND3 (N19477, N19474, N15720, N17929);
xor XOR2 (N19478, N19470, N18491);
buf BUF1 (N19479, N19465);
and AND2 (N19480, N19475, N1596);
nor NOR3 (N19481, N19466, N11753, N12076);
xor XOR2 (N19482, N19469, N9149);
or OR3 (N19483, N19468, N7202, N3189);
and AND2 (N19484, N19478, N3467);
or OR4 (N19485, N19479, N13167, N14591, N12497);
or OR4 (N19486, N19477, N18312, N10560, N4639);
not NOT1 (N19487, N19483);
nand NAND3 (N19488, N19456, N1449, N3665);
not NOT1 (N19489, N19476);
or OR4 (N19490, N19449, N15877, N13494, N12503);
and AND4 (N19491, N19480, N7698, N3459, N11230);
xor XOR2 (N19492, N19487, N15497);
buf BUF1 (N19493, N19492);
not NOT1 (N19494, N19482);
and AND2 (N19495, N19485, N6854);
nor NOR3 (N19496, N19490, N296, N14768);
xor XOR2 (N19497, N19495, N4998);
xor XOR2 (N19498, N19494, N12614);
nand NAND3 (N19499, N19484, N13516, N6087);
and AND2 (N19500, N19496, N5933);
xor XOR2 (N19501, N19500, N13563);
buf BUF1 (N19502, N19493);
nand NAND2 (N19503, N19502, N4754);
and AND4 (N19504, N19503, N8723, N5471, N7725);
nor NOR2 (N19505, N19488, N11537);
nor NOR3 (N19506, N19499, N8196, N10902);
or OR3 (N19507, N19481, N8138, N17167);
nand NAND3 (N19508, N19486, N5361, N14009);
xor XOR2 (N19509, N19497, N12343);
xor XOR2 (N19510, N19498, N12960);
or OR4 (N19511, N19491, N11329, N1625, N18902);
buf BUF1 (N19512, N19509);
nand NAND2 (N19513, N19504, N2474);
not NOT1 (N19514, N19501);
nand NAND2 (N19515, N19513, N9506);
nor NOR4 (N19516, N19507, N16987, N2423, N6597);
xor XOR2 (N19517, N19505, N12852);
or OR2 (N19518, N19517, N16936);
or OR4 (N19519, N19508, N362, N19074, N4451);
or OR3 (N19520, N19510, N1702, N2180);
not NOT1 (N19521, N19520);
not NOT1 (N19522, N19516);
xor XOR2 (N19523, N19511, N1129);
nor NOR3 (N19524, N19518, N11596, N14879);
buf BUF1 (N19525, N19522);
xor XOR2 (N19526, N19506, N9706);
and AND2 (N19527, N19512, N18444);
not NOT1 (N19528, N19526);
or OR3 (N19529, N19528, N13146, N9892);
nor NOR3 (N19530, N19525, N2442, N14342);
xor XOR2 (N19531, N19519, N16647);
nand NAND3 (N19532, N19529, N10511, N19058);
not NOT1 (N19533, N19530);
nor NOR3 (N19534, N19489, N8309, N5180);
nor NOR2 (N19535, N19533, N14431);
not NOT1 (N19536, N19514);
xor XOR2 (N19537, N19535, N8304);
nor NOR2 (N19538, N19532, N17467);
buf BUF1 (N19539, N19523);
xor XOR2 (N19540, N19524, N2056);
xor XOR2 (N19541, N19538, N15179);
nor NOR3 (N19542, N19536, N14381, N17387);
not NOT1 (N19543, N19540);
buf BUF1 (N19544, N19541);
nand NAND3 (N19545, N19544, N15886, N17391);
not NOT1 (N19546, N19521);
nor NOR4 (N19547, N19546, N8542, N3429, N18771);
or OR4 (N19548, N19534, N2555, N9486, N12268);
nand NAND3 (N19549, N19545, N13608, N8789);
and AND4 (N19550, N19549, N7720, N4720, N12903);
not NOT1 (N19551, N19548);
not NOT1 (N19552, N19531);
or OR2 (N19553, N19552, N16014);
or OR2 (N19554, N19515, N14740);
nand NAND4 (N19555, N19537, N13392, N12030, N7293);
nor NOR4 (N19556, N19551, N16833, N11473, N17625);
xor XOR2 (N19557, N19543, N9193);
nor NOR4 (N19558, N19553, N15172, N11202, N10092);
buf BUF1 (N19559, N19555);
xor XOR2 (N19560, N19527, N19445);
buf BUF1 (N19561, N19539);
xor XOR2 (N19562, N19560, N8220);
buf BUF1 (N19563, N19554);
and AND3 (N19564, N19561, N18327, N7367);
not NOT1 (N19565, N19557);
buf BUF1 (N19566, N19559);
nand NAND3 (N19567, N19542, N1011, N9622);
buf BUF1 (N19568, N19563);
xor XOR2 (N19569, N19566, N9902);
not NOT1 (N19570, N19567);
or OR2 (N19571, N19547, N17741);
not NOT1 (N19572, N19568);
nor NOR4 (N19573, N19550, N19435, N3041, N17578);
buf BUF1 (N19574, N19564);
and AND4 (N19575, N19558, N6105, N11656, N6434);
not NOT1 (N19576, N19574);
xor XOR2 (N19577, N19562, N5077);
buf BUF1 (N19578, N19573);
nand NAND2 (N19579, N19571, N812);
nand NAND3 (N19580, N19575, N7930, N7054);
not NOT1 (N19581, N19577);
not NOT1 (N19582, N19579);
nand NAND3 (N19583, N19572, N14150, N17544);
or OR4 (N19584, N19565, N16122, N19241, N8243);
buf BUF1 (N19585, N19570);
xor XOR2 (N19586, N19585, N8197);
nand NAND3 (N19587, N19584, N18875, N972);
nor NOR2 (N19588, N19582, N18906);
or OR2 (N19589, N19586, N10835);
nor NOR3 (N19590, N19581, N13539, N18431);
buf BUF1 (N19591, N19556);
xor XOR2 (N19592, N19588, N15409);
and AND3 (N19593, N19590, N8219, N17809);
buf BUF1 (N19594, N19583);
xor XOR2 (N19595, N19578, N5947);
or OR4 (N19596, N19589, N14492, N3471, N13355);
nor NOR2 (N19597, N19569, N7358);
and AND4 (N19598, N19592, N10813, N15641, N13123);
nand NAND2 (N19599, N19576, N7994);
xor XOR2 (N19600, N19596, N6082);
nand NAND2 (N19601, N19594, N3314);
buf BUF1 (N19602, N19587);
or OR3 (N19603, N19599, N12476, N18982);
buf BUF1 (N19604, N19600);
nand NAND2 (N19605, N19602, N9719);
xor XOR2 (N19606, N19603, N19360);
or OR4 (N19607, N19593, N5194, N12398, N18006);
xor XOR2 (N19608, N19597, N10376);
xor XOR2 (N19609, N19607, N11249);
and AND4 (N19610, N19604, N9003, N3139, N2840);
and AND2 (N19611, N19609, N2893);
buf BUF1 (N19612, N19605);
xor XOR2 (N19613, N19606, N6849);
and AND2 (N19614, N19601, N8427);
buf BUF1 (N19615, N19598);
nand NAND3 (N19616, N19595, N3373, N949);
buf BUF1 (N19617, N19616);
and AND4 (N19618, N19580, N1268, N18869, N3696);
or OR2 (N19619, N19613, N7169);
not NOT1 (N19620, N19614);
nand NAND3 (N19621, N19618, N14248, N3354);
or OR2 (N19622, N19610, N10295);
and AND3 (N19623, N19620, N6619, N10880);
xor XOR2 (N19624, N19619, N12170);
not NOT1 (N19625, N19617);
xor XOR2 (N19626, N19624, N10768);
not NOT1 (N19627, N19591);
nor NOR3 (N19628, N19622, N11262, N14866);
or OR4 (N19629, N19621, N18805, N15695, N5340);
nand NAND4 (N19630, N19608, N13671, N18725, N6831);
or OR3 (N19631, N19623, N8989, N11700);
nor NOR2 (N19632, N19630, N14367);
and AND3 (N19633, N19632, N11068, N7168);
nor NOR2 (N19634, N19633, N399);
nand NAND4 (N19635, N19625, N11087, N726, N920);
not NOT1 (N19636, N19612);
not NOT1 (N19637, N19634);
nor NOR4 (N19638, N19629, N8079, N1772, N3945);
nand NAND4 (N19639, N19636, N10473, N12703, N9069);
xor XOR2 (N19640, N19635, N11051);
nand NAND3 (N19641, N19627, N6752, N8744);
nand NAND3 (N19642, N19638, N15724, N7860);
nor NOR4 (N19643, N19626, N6247, N6551, N2807);
buf BUF1 (N19644, N19640);
buf BUF1 (N19645, N19631);
xor XOR2 (N19646, N19645, N7744);
buf BUF1 (N19647, N19628);
nand NAND3 (N19648, N19646, N17526, N18876);
xor XOR2 (N19649, N19611, N7300);
not NOT1 (N19650, N19643);
not NOT1 (N19651, N19648);
buf BUF1 (N19652, N19649);
not NOT1 (N19653, N19647);
not NOT1 (N19654, N19615);
nor NOR2 (N19655, N19652, N1919);
and AND2 (N19656, N19637, N14807);
and AND4 (N19657, N19654, N15861, N3443, N10412);
not NOT1 (N19658, N19641);
nor NOR4 (N19659, N19653, N5271, N3635, N13310);
xor XOR2 (N19660, N19642, N15504);
xor XOR2 (N19661, N19644, N17936);
or OR3 (N19662, N19661, N4348, N14295);
xor XOR2 (N19663, N19658, N4797);
nor NOR3 (N19664, N19655, N6478, N18375);
and AND4 (N19665, N19657, N9333, N16115, N16042);
and AND2 (N19666, N19650, N19233);
nor NOR3 (N19667, N19659, N14666, N4817);
or OR4 (N19668, N19665, N3066, N10629, N10502);
nand NAND4 (N19669, N19656, N6652, N9112, N16325);
or OR2 (N19670, N19669, N17356);
nor NOR2 (N19671, N19651, N9775);
not NOT1 (N19672, N19667);
nand NAND3 (N19673, N19666, N1701, N9100);
or OR4 (N19674, N19668, N3947, N1367, N12162);
buf BUF1 (N19675, N19660);
not NOT1 (N19676, N19675);
and AND2 (N19677, N19676, N18800);
and AND2 (N19678, N19671, N4417);
not NOT1 (N19679, N19677);
or OR3 (N19680, N19672, N4652, N657);
nand NAND2 (N19681, N19670, N11787);
nand NAND3 (N19682, N19680, N13909, N4184);
buf BUF1 (N19683, N19639);
or OR4 (N19684, N19682, N7225, N5350, N679);
xor XOR2 (N19685, N19681, N8318);
and AND4 (N19686, N19673, N5391, N483, N5511);
and AND3 (N19687, N19685, N5554, N13732);
nand NAND3 (N19688, N19674, N515, N8711);
nor NOR4 (N19689, N19684, N805, N6082, N11324);
buf BUF1 (N19690, N19689);
not NOT1 (N19691, N19662);
nand NAND3 (N19692, N19690, N5758, N2275);
nand NAND4 (N19693, N19692, N4726, N7952, N7099);
nand NAND2 (N19694, N19691, N5680);
and AND2 (N19695, N19686, N12146);
nor NOR4 (N19696, N19664, N2096, N19195, N3951);
or OR2 (N19697, N19688, N2946);
nand NAND4 (N19698, N19687, N11603, N11169, N12214);
nor NOR3 (N19699, N19697, N8026, N2747);
nand NAND2 (N19700, N19683, N6200);
buf BUF1 (N19701, N19694);
or OR4 (N19702, N19679, N10, N15511, N795);
buf BUF1 (N19703, N19701);
buf BUF1 (N19704, N19699);
buf BUF1 (N19705, N19704);
xor XOR2 (N19706, N19702, N19326);
nand NAND4 (N19707, N19698, N5646, N10237, N17525);
xor XOR2 (N19708, N19707, N1234);
nor NOR2 (N19709, N19703, N8196);
nor NOR4 (N19710, N19706, N15460, N9290, N3185);
or OR2 (N19711, N19696, N13514);
nor NOR3 (N19712, N19710, N5030, N19094);
xor XOR2 (N19713, N19708, N18473);
not NOT1 (N19714, N19712);
not NOT1 (N19715, N19705);
nand NAND2 (N19716, N19709, N18186);
and AND4 (N19717, N19714, N11887, N4742, N10186);
xor XOR2 (N19718, N19716, N4447);
or OR3 (N19719, N19713, N4503, N15384);
or OR3 (N19720, N19693, N9021, N5026);
or OR2 (N19721, N19720, N11689);
nor NOR3 (N19722, N19718, N11378, N7850);
not NOT1 (N19723, N19711);
or OR4 (N19724, N19678, N4468, N7176, N14731);
or OR4 (N19725, N19721, N17039, N8506, N8949);
or OR4 (N19726, N19725, N3282, N9504, N13135);
and AND4 (N19727, N19717, N19394, N12681, N4326);
xor XOR2 (N19728, N19722, N8112);
nand NAND4 (N19729, N19695, N18759, N16169, N7621);
nand NAND3 (N19730, N19724, N15797, N19625);
nand NAND3 (N19731, N19730, N14309, N6227);
not NOT1 (N19732, N19700);
nand NAND4 (N19733, N19726, N11042, N18091, N8328);
and AND4 (N19734, N19728, N3864, N652, N11602);
not NOT1 (N19735, N19715);
xor XOR2 (N19736, N19719, N5538);
or OR3 (N19737, N19736, N5857, N8645);
nor NOR2 (N19738, N19737, N12669);
nor NOR4 (N19739, N19729, N3955, N12730, N19259);
and AND3 (N19740, N19733, N2866, N12309);
nand NAND3 (N19741, N19738, N10612, N14936);
nand NAND4 (N19742, N19735, N12256, N11428, N394);
xor XOR2 (N19743, N19739, N291);
nand NAND3 (N19744, N19723, N16355, N19522);
not NOT1 (N19745, N19743);
and AND3 (N19746, N19734, N4692, N16240);
buf BUF1 (N19747, N19742);
buf BUF1 (N19748, N19747);
nor NOR3 (N19749, N19744, N18555, N5273);
nand NAND4 (N19750, N19740, N1723, N2282, N7811);
not NOT1 (N19751, N19749);
and AND2 (N19752, N19727, N12009);
xor XOR2 (N19753, N19750, N18904);
and AND2 (N19754, N19752, N10819);
nor NOR2 (N19755, N19753, N2077);
nor NOR4 (N19756, N19755, N8999, N14908, N19624);
not NOT1 (N19757, N19756);
or OR4 (N19758, N19751, N19640, N11929, N15627);
nor NOR2 (N19759, N19731, N13436);
not NOT1 (N19760, N19754);
xor XOR2 (N19761, N19663, N12618);
xor XOR2 (N19762, N19746, N16472);
or OR2 (N19763, N19759, N17796);
and AND2 (N19764, N19758, N19010);
nand NAND2 (N19765, N19757, N18838);
nand NAND3 (N19766, N19760, N19492, N5009);
buf BUF1 (N19767, N19741);
not NOT1 (N19768, N19732);
xor XOR2 (N19769, N19764, N12525);
nor NOR4 (N19770, N19768, N3111, N4039, N18814);
buf BUF1 (N19771, N19745);
not NOT1 (N19772, N19770);
and AND3 (N19773, N19769, N19246, N849);
buf BUF1 (N19774, N19761);
xor XOR2 (N19775, N19767, N13969);
and AND3 (N19776, N19762, N2458, N12930);
nand NAND3 (N19777, N19774, N10015, N13203);
and AND4 (N19778, N19773, N15171, N15824, N16456);
buf BUF1 (N19779, N19763);
and AND4 (N19780, N19772, N16545, N4861, N5820);
not NOT1 (N19781, N19779);
buf BUF1 (N19782, N19775);
xor XOR2 (N19783, N19776, N12005);
or OR2 (N19784, N19766, N11752);
not NOT1 (N19785, N19783);
xor XOR2 (N19786, N19780, N11505);
not NOT1 (N19787, N19765);
nor NOR4 (N19788, N19778, N6782, N11929, N4649);
buf BUF1 (N19789, N19748);
and AND3 (N19790, N19782, N16522, N14136);
and AND3 (N19791, N19771, N19122, N1299);
or OR2 (N19792, N19791, N3753);
or OR4 (N19793, N19784, N17788, N16137, N14401);
not NOT1 (N19794, N19790);
or OR2 (N19795, N19781, N9789);
not NOT1 (N19796, N19788);
buf BUF1 (N19797, N19785);
buf BUF1 (N19798, N19777);
nand NAND3 (N19799, N19798, N8374, N12294);
nand NAND4 (N19800, N19796, N18024, N5400, N16366);
nand NAND3 (N19801, N19794, N9773, N13344);
and AND2 (N19802, N19789, N11792);
and AND2 (N19803, N19800, N12245);
and AND3 (N19804, N19787, N13056, N2662);
nor NOR2 (N19805, N19793, N12450);
not NOT1 (N19806, N19792);
nor NOR2 (N19807, N19804, N17242);
xor XOR2 (N19808, N19799, N876);
and AND2 (N19809, N19795, N10778);
and AND2 (N19810, N19809, N14428);
not NOT1 (N19811, N19801);
nand NAND4 (N19812, N19786, N17081, N10809, N15343);
nand NAND4 (N19813, N19803, N18817, N11314, N6451);
nor NOR3 (N19814, N19797, N6055, N19023);
nand NAND3 (N19815, N19805, N4520, N731);
or OR2 (N19816, N19808, N1847);
or OR2 (N19817, N19813, N15469);
nor NOR3 (N19818, N19806, N14839, N18054);
and AND2 (N19819, N19811, N15162);
or OR2 (N19820, N19815, N3295);
nand NAND2 (N19821, N19810, N11568);
or OR4 (N19822, N19802, N1151, N18769, N13775);
and AND3 (N19823, N19807, N2711, N11721);
nand NAND4 (N19824, N19816, N7217, N10591, N8798);
not NOT1 (N19825, N19818);
not NOT1 (N19826, N19824);
or OR2 (N19827, N19814, N9470);
or OR3 (N19828, N19826, N3803, N5528);
and AND3 (N19829, N19825, N13909, N11973);
nand NAND4 (N19830, N19821, N2455, N11230, N13936);
xor XOR2 (N19831, N19817, N15301);
or OR3 (N19832, N19831, N9051, N5264);
or OR2 (N19833, N19822, N2460);
xor XOR2 (N19834, N19823, N18320);
and AND2 (N19835, N19827, N16043);
or OR2 (N19836, N19832, N3530);
nor NOR3 (N19837, N19834, N8408, N18337);
not NOT1 (N19838, N19836);
nor NOR3 (N19839, N19829, N4370, N12034);
xor XOR2 (N19840, N19837, N8142);
or OR2 (N19841, N19839, N15776);
buf BUF1 (N19842, N19828);
buf BUF1 (N19843, N19841);
and AND3 (N19844, N19812, N3215, N5016);
nor NOR4 (N19845, N19819, N4952, N6872, N9178);
xor XOR2 (N19846, N19835, N16563);
not NOT1 (N19847, N19830);
or OR2 (N19848, N19820, N14970);
or OR3 (N19849, N19833, N6517, N12651);
not NOT1 (N19850, N19849);
not NOT1 (N19851, N19847);
xor XOR2 (N19852, N19851, N9760);
buf BUF1 (N19853, N19848);
not NOT1 (N19854, N19846);
and AND3 (N19855, N19843, N15712, N19566);
nand NAND4 (N19856, N19850, N6377, N4448, N2509);
xor XOR2 (N19857, N19840, N10045);
xor XOR2 (N19858, N19854, N18520);
nor NOR2 (N19859, N19845, N14363);
buf BUF1 (N19860, N19852);
nand NAND3 (N19861, N19857, N1674, N9376);
xor XOR2 (N19862, N19860, N9117);
nor NOR2 (N19863, N19844, N3482);
and AND2 (N19864, N19858, N13267);
not NOT1 (N19865, N19855);
xor XOR2 (N19866, N19838, N2535);
and AND4 (N19867, N19853, N17863, N13852, N1922);
nor NOR3 (N19868, N19864, N4756, N9432);
xor XOR2 (N19869, N19865, N1131);
and AND3 (N19870, N19863, N6523, N8544);
and AND2 (N19871, N19861, N9776);
buf BUF1 (N19872, N19856);
not NOT1 (N19873, N19859);
nand NAND4 (N19874, N19868, N16951, N19862, N5015);
nand NAND3 (N19875, N8401, N15553, N15093);
or OR3 (N19876, N19873, N18651, N12385);
and AND3 (N19877, N19842, N1799, N7582);
xor XOR2 (N19878, N19870, N14907);
or OR3 (N19879, N19872, N8660, N8950);
nand NAND2 (N19880, N19879, N18533);
or OR2 (N19881, N19880, N13476);
and AND4 (N19882, N19871, N16643, N7811, N758);
nor NOR4 (N19883, N19881, N17870, N120, N19762);
nand NAND3 (N19884, N19876, N2758, N19289);
not NOT1 (N19885, N19884);
buf BUF1 (N19886, N19875);
or OR2 (N19887, N19874, N8277);
not NOT1 (N19888, N19867);
and AND4 (N19889, N19883, N17441, N7754, N10424);
nor NOR4 (N19890, N19882, N19536, N6998, N16960);
nor NOR2 (N19891, N19888, N18440);
nor NOR2 (N19892, N19890, N580);
nor NOR3 (N19893, N19892, N3522, N5132);
and AND4 (N19894, N19886, N8481, N16551, N268);
and AND3 (N19895, N19885, N3253, N14463);
nor NOR3 (N19896, N19894, N18135, N1908);
not NOT1 (N19897, N19891);
not NOT1 (N19898, N19895);
and AND3 (N19899, N19869, N12390, N6261);
not NOT1 (N19900, N19887);
nor NOR3 (N19901, N19900, N19268, N1018);
nor NOR2 (N19902, N19896, N9175);
or OR2 (N19903, N19877, N12372);
or OR4 (N19904, N19903, N18333, N11646, N4201);
buf BUF1 (N19905, N19902);
nand NAND4 (N19906, N19899, N14475, N14196, N3461);
xor XOR2 (N19907, N19904, N4695);
or OR4 (N19908, N19901, N10259, N13834, N6495);
nand NAND4 (N19909, N19866, N6041, N14559, N219);
and AND2 (N19910, N19898, N10124);
xor XOR2 (N19911, N19893, N12551);
or OR2 (N19912, N19906, N16849);
or OR2 (N19913, N19889, N15963);
nand NAND4 (N19914, N19897, N18449, N19099, N12782);
or OR2 (N19915, N19914, N17986);
and AND3 (N19916, N19905, N5765, N3222);
and AND3 (N19917, N19909, N14857, N5097);
xor XOR2 (N19918, N19916, N8337);
nand NAND4 (N19919, N19917, N8341, N5005, N9618);
buf BUF1 (N19920, N19918);
or OR4 (N19921, N19912, N3498, N19385, N14930);
and AND4 (N19922, N19921, N8542, N14579, N530);
or OR4 (N19923, N19878, N6641, N6126, N7582);
buf BUF1 (N19924, N19920);
buf BUF1 (N19925, N19915);
or OR2 (N19926, N19923, N17181);
nor NOR2 (N19927, N19925, N15934);
nand NAND4 (N19928, N19922, N4027, N17358, N14111);
nor NOR3 (N19929, N19907, N4541, N16344);
xor XOR2 (N19930, N19929, N8948);
not NOT1 (N19931, N19919);
not NOT1 (N19932, N19931);
nand NAND4 (N19933, N19924, N13182, N7, N2319);
nand NAND4 (N19934, N19910, N817, N12654, N18845);
not NOT1 (N19935, N19911);
not NOT1 (N19936, N19928);
nand NAND4 (N19937, N19934, N18129, N3280, N17788);
nand NAND2 (N19938, N19937, N10489);
buf BUF1 (N19939, N19933);
and AND2 (N19940, N19908, N14840);
nand NAND3 (N19941, N19940, N3325, N288);
nand NAND4 (N19942, N19941, N11219, N10678, N9942);
nor NOR3 (N19943, N19936, N13997, N11827);
nand NAND4 (N19944, N19939, N12854, N19499, N11334);
buf BUF1 (N19945, N19927);
xor XOR2 (N19946, N19943, N5932);
not NOT1 (N19947, N19945);
nand NAND2 (N19948, N19947, N14470);
or OR2 (N19949, N19946, N19697);
or OR4 (N19950, N19938, N17238, N11832, N19185);
or OR3 (N19951, N19949, N2649, N17248);
or OR2 (N19952, N19926, N12498);
nor NOR2 (N19953, N19935, N4723);
buf BUF1 (N19954, N19942);
nand NAND2 (N19955, N19953, N11655);
and AND3 (N19956, N19944, N3021, N12900);
xor XOR2 (N19957, N19952, N9846);
not NOT1 (N19958, N19954);
xor XOR2 (N19959, N19948, N4596);
nand NAND3 (N19960, N19958, N11206, N12752);
and AND3 (N19961, N19960, N7436, N9708);
or OR3 (N19962, N19950, N2477, N3546);
nor NOR3 (N19963, N19913, N12005, N11799);
xor XOR2 (N19964, N19956, N7890);
and AND2 (N19965, N19959, N6508);
or OR2 (N19966, N19951, N5759);
not NOT1 (N19967, N19961);
nand NAND4 (N19968, N19932, N10416, N9696, N16593);
and AND4 (N19969, N19964, N343, N18493, N1486);
not NOT1 (N19970, N19968);
and AND3 (N19971, N19963, N12060, N18575);
buf BUF1 (N19972, N19955);
nand NAND2 (N19973, N19930, N15567);
or OR2 (N19974, N19965, N5377);
nand NAND3 (N19975, N19962, N17267, N3918);
or OR4 (N19976, N19967, N16185, N13830, N5409);
or OR3 (N19977, N19975, N6326, N11162);
nand NAND2 (N19978, N19977, N958);
nor NOR3 (N19979, N19966, N16069, N12648);
buf BUF1 (N19980, N19979);
xor XOR2 (N19981, N19971, N8211);
nor NOR2 (N19982, N19980, N9762);
nor NOR3 (N19983, N19973, N4254, N8268);
and AND4 (N19984, N19982, N17518, N3239, N9657);
not NOT1 (N19985, N19983);
nor NOR3 (N19986, N19972, N15520, N14966);
xor XOR2 (N19987, N19957, N10415);
not NOT1 (N19988, N19986);
or OR4 (N19989, N19981, N7601, N13355, N12705);
buf BUF1 (N19990, N19985);
not NOT1 (N19991, N19974);
and AND2 (N19992, N19990, N18213);
buf BUF1 (N19993, N19991);
not NOT1 (N19994, N19987);
or OR3 (N19995, N19994, N6052, N19214);
nand NAND3 (N19996, N19992, N14740, N6737);
nand NAND2 (N19997, N19969, N11917);
or OR4 (N19998, N19995, N13539, N13042, N3092);
and AND3 (N19999, N19970, N13687, N11172);
or OR3 (N20000, N19993, N7779, N11565);
or OR3 (N20001, N19999, N2497, N4439);
nand NAND3 (N20002, N19996, N392, N2586);
xor XOR2 (N20003, N19997, N16230);
or OR3 (N20004, N20002, N2116, N5840);
or OR4 (N20005, N20003, N19498, N10173, N12946);
not NOT1 (N20006, N19984);
nand NAND2 (N20007, N20004, N9702);
not NOT1 (N20008, N20005);
and AND3 (N20009, N20007, N10072, N3050);
nand NAND4 (N20010, N20008, N2361, N14805, N18300);
nor NOR3 (N20011, N19978, N7788, N1444);
nor NOR3 (N20012, N20000, N17195, N10985);
or OR2 (N20013, N20011, N13201);
buf BUF1 (N20014, N20010);
nand NAND3 (N20015, N20001, N1596, N9772);
nor NOR3 (N20016, N19976, N8843, N15499);
xor XOR2 (N20017, N20009, N10858);
xor XOR2 (N20018, N20017, N19644);
or OR3 (N20019, N20013, N8151, N1407);
and AND3 (N20020, N20014, N5532, N17976);
nand NAND2 (N20021, N20019, N18385);
nor NOR2 (N20022, N20018, N15865);
or OR3 (N20023, N20021, N3512, N8772);
not NOT1 (N20024, N20022);
nor NOR4 (N20025, N20016, N6675, N17241, N6786);
and AND3 (N20026, N20024, N11318, N18462);
nand NAND4 (N20027, N20020, N8579, N13770, N6287);
or OR2 (N20028, N20023, N12836);
buf BUF1 (N20029, N19998);
nor NOR3 (N20030, N20012, N10880, N12064);
not NOT1 (N20031, N20029);
nor NOR4 (N20032, N20027, N18485, N16090, N11280);
buf BUF1 (N20033, N19989);
nor NOR2 (N20034, N20015, N18275);
nor NOR4 (N20035, N19988, N17527, N3351, N9695);
or OR4 (N20036, N20006, N3304, N8958, N17031);
and AND4 (N20037, N20030, N13933, N4674, N991);
xor XOR2 (N20038, N20037, N2239);
buf BUF1 (N20039, N20033);
buf BUF1 (N20040, N20034);
nand NAND3 (N20041, N20032, N19091, N14776);
buf BUF1 (N20042, N20031);
and AND4 (N20043, N20025, N4410, N12590, N18737);
not NOT1 (N20044, N20042);
or OR3 (N20045, N20040, N18958, N1014);
nand NAND3 (N20046, N20043, N15604, N19159);
nor NOR4 (N20047, N20028, N16424, N9338, N18679);
and AND4 (N20048, N20036, N17783, N7287, N5217);
xor XOR2 (N20049, N20048, N6776);
not NOT1 (N20050, N20039);
or OR3 (N20051, N20041, N9535, N13633);
xor XOR2 (N20052, N20045, N7428);
nand NAND3 (N20053, N20049, N5205, N7090);
not NOT1 (N20054, N20044);
nor NOR2 (N20055, N20054, N9843);
and AND4 (N20056, N20035, N14911, N7453, N13810);
nand NAND3 (N20057, N20046, N18158, N17508);
or OR4 (N20058, N20051, N19807, N12094, N478);
not NOT1 (N20059, N20058);
buf BUF1 (N20060, N20026);
not NOT1 (N20061, N20056);
and AND2 (N20062, N20061, N2837);
xor XOR2 (N20063, N20053, N1469);
buf BUF1 (N20064, N20062);
or OR4 (N20065, N20060, N18509, N1641, N4981);
nor NOR3 (N20066, N20047, N4234, N14916);
or OR3 (N20067, N20063, N12637, N5847);
xor XOR2 (N20068, N20064, N4763);
nand NAND3 (N20069, N20067, N19738, N17315);
buf BUF1 (N20070, N20068);
or OR3 (N20071, N20057, N3682, N16295);
nand NAND2 (N20072, N20052, N1900);
nand NAND3 (N20073, N20071, N13223, N12481);
or OR3 (N20074, N20065, N17490, N15890);
and AND3 (N20075, N20050, N354, N4409);
nand NAND4 (N20076, N20072, N17173, N17344, N17068);
nor NOR3 (N20077, N20070, N2205, N6345);
not NOT1 (N20078, N20055);
xor XOR2 (N20079, N20074, N4701);
nand NAND2 (N20080, N20073, N14836);
nand NAND3 (N20081, N20080, N11333, N1199);
and AND4 (N20082, N20081, N369, N16164, N6821);
xor XOR2 (N20083, N20066, N9768);
and AND2 (N20084, N20078, N13922);
and AND2 (N20085, N20076, N11673);
not NOT1 (N20086, N20059);
not NOT1 (N20087, N20082);
nand NAND4 (N20088, N20038, N6858, N5318, N19760);
buf BUF1 (N20089, N20069);
nor NOR3 (N20090, N20087, N18722, N15870);
and AND4 (N20091, N20083, N237, N8578, N4206);
and AND2 (N20092, N20089, N12276);
and AND3 (N20093, N20086, N19767, N2202);
or OR3 (N20094, N20093, N9889, N8187);
buf BUF1 (N20095, N20091);
nand NAND3 (N20096, N20077, N981, N7231);
buf BUF1 (N20097, N20096);
not NOT1 (N20098, N20092);
buf BUF1 (N20099, N20094);
nor NOR4 (N20100, N20084, N12886, N188, N18725);
buf BUF1 (N20101, N20079);
not NOT1 (N20102, N20098);
and AND2 (N20103, N20097, N12334);
and AND3 (N20104, N20095, N2424, N18850);
xor XOR2 (N20105, N20090, N6348);
or OR3 (N20106, N20101, N18380, N16683);
xor XOR2 (N20107, N20106, N985);
or OR2 (N20108, N20088, N13252);
buf BUF1 (N20109, N20102);
buf BUF1 (N20110, N20108);
buf BUF1 (N20111, N20104);
or OR3 (N20112, N20111, N13755, N11599);
and AND2 (N20113, N20075, N6640);
and AND2 (N20114, N20085, N3856);
and AND4 (N20115, N20114, N19452, N7907, N10320);
and AND3 (N20116, N20112, N16689, N11357);
nor NOR4 (N20117, N20107, N6132, N2128, N5365);
or OR4 (N20118, N20110, N3940, N8485, N19051);
nor NOR2 (N20119, N20103, N10377);
buf BUF1 (N20120, N20118);
or OR3 (N20121, N20115, N2583, N12436);
not NOT1 (N20122, N20120);
or OR2 (N20123, N20099, N18645);
not NOT1 (N20124, N20100);
nand NAND2 (N20125, N20109, N17891);
nor NOR2 (N20126, N20125, N17924);
and AND3 (N20127, N20116, N15736, N2992);
nor NOR3 (N20128, N20119, N13336, N8378);
buf BUF1 (N20129, N20117);
or OR3 (N20130, N20129, N6697, N9166);
xor XOR2 (N20131, N20113, N7610);
xor XOR2 (N20132, N20122, N18970);
not NOT1 (N20133, N20123);
and AND4 (N20134, N20128, N2146, N18579, N17097);
buf BUF1 (N20135, N20131);
nor NOR3 (N20136, N20133, N7471, N1071);
nand NAND4 (N20137, N20134, N13149, N12192, N13240);
nor NOR2 (N20138, N20130, N4647);
nor NOR2 (N20139, N20124, N18834);
not NOT1 (N20140, N20136);
and AND2 (N20141, N20121, N7984);
and AND4 (N20142, N20127, N17894, N10652, N4554);
xor XOR2 (N20143, N20126, N14330);
nor NOR2 (N20144, N20143, N3626);
nor NOR4 (N20145, N20135, N10543, N3357, N16031);
xor XOR2 (N20146, N20139, N6718);
and AND4 (N20147, N20138, N16167, N2371, N10223);
buf BUF1 (N20148, N20142);
not NOT1 (N20149, N20137);
nand NAND3 (N20150, N20141, N8237, N3606);
xor XOR2 (N20151, N20147, N11752);
nor NOR3 (N20152, N20150, N17370, N12764);
nor NOR4 (N20153, N20132, N11885, N9344, N15307);
nor NOR3 (N20154, N20151, N15505, N19606);
nor NOR3 (N20155, N20145, N8026, N8678);
not NOT1 (N20156, N20152);
or OR3 (N20157, N20144, N12290, N1548);
xor XOR2 (N20158, N20153, N3839);
nor NOR4 (N20159, N20148, N11295, N18070, N7764);
not NOT1 (N20160, N20157);
nor NOR4 (N20161, N20160, N7395, N17749, N1728);
nor NOR2 (N20162, N20140, N3411);
xor XOR2 (N20163, N20156, N4555);
xor XOR2 (N20164, N20149, N680);
nor NOR3 (N20165, N20164, N15842, N5920);
xor XOR2 (N20166, N20162, N15280);
nand NAND3 (N20167, N20158, N10123, N12539);
nor NOR4 (N20168, N20146, N15581, N15778, N10141);
xor XOR2 (N20169, N20167, N971);
and AND3 (N20170, N20154, N13208, N16677);
buf BUF1 (N20171, N20159);
xor XOR2 (N20172, N20155, N841);
not NOT1 (N20173, N20163);
or OR2 (N20174, N20105, N6733);
buf BUF1 (N20175, N20170);
xor XOR2 (N20176, N20172, N12801);
not NOT1 (N20177, N20161);
and AND2 (N20178, N20173, N6094);
xor XOR2 (N20179, N20168, N13753);
buf BUF1 (N20180, N20176);
buf BUF1 (N20181, N20171);
nand NAND3 (N20182, N20177, N17307, N6132);
nor NOR4 (N20183, N20179, N2804, N13152, N18573);
nand NAND4 (N20184, N20180, N6090, N18541, N15142);
xor XOR2 (N20185, N20183, N19781);
xor XOR2 (N20186, N20174, N13138);
or OR3 (N20187, N20175, N10445, N8534);
xor XOR2 (N20188, N20182, N14837);
buf BUF1 (N20189, N20188);
xor XOR2 (N20190, N20187, N1085);
xor XOR2 (N20191, N20184, N12093);
buf BUF1 (N20192, N20166);
nor NOR3 (N20193, N20189, N1474, N19939);
and AND3 (N20194, N20186, N10483, N10965);
buf BUF1 (N20195, N20169);
not NOT1 (N20196, N20193);
buf BUF1 (N20197, N20185);
xor XOR2 (N20198, N20190, N9474);
nand NAND4 (N20199, N20198, N15445, N13302, N445);
nand NAND4 (N20200, N20197, N918, N16673, N13004);
xor XOR2 (N20201, N20181, N901);
or OR3 (N20202, N20200, N17516, N13157);
buf BUF1 (N20203, N20195);
nand NAND3 (N20204, N20202, N7483, N5911);
not NOT1 (N20205, N20201);
buf BUF1 (N20206, N20191);
xor XOR2 (N20207, N20194, N649);
or OR3 (N20208, N20165, N15233, N19785);
or OR4 (N20209, N20203, N7358, N14298, N1232);
buf BUF1 (N20210, N20192);
or OR2 (N20211, N20207, N18363);
nand NAND2 (N20212, N20210, N12194);
nand NAND4 (N20213, N20209, N9269, N2241, N1709);
xor XOR2 (N20214, N20199, N5290);
xor XOR2 (N20215, N20196, N18747);
and AND2 (N20216, N20215, N14961);
buf BUF1 (N20217, N20216);
xor XOR2 (N20218, N20211, N19590);
xor XOR2 (N20219, N20208, N17193);
and AND2 (N20220, N20218, N10914);
nor NOR4 (N20221, N20212, N2285, N7494, N13173);
and AND2 (N20222, N20206, N6487);
and AND3 (N20223, N20204, N6066, N16585);
buf BUF1 (N20224, N20178);
and AND2 (N20225, N20219, N6796);
nand NAND3 (N20226, N20214, N3895, N6490);
not NOT1 (N20227, N20222);
xor XOR2 (N20228, N20217, N5164);
and AND4 (N20229, N20213, N12086, N19705, N16713);
nand NAND3 (N20230, N20227, N9010, N5432);
nand NAND4 (N20231, N20221, N16736, N628, N11485);
nand NAND3 (N20232, N20228, N104, N10353);
or OR4 (N20233, N20230, N8159, N16575, N5293);
xor XOR2 (N20234, N20226, N11554);
nand NAND2 (N20235, N20232, N4780);
buf BUF1 (N20236, N20223);
not NOT1 (N20237, N20224);
xor XOR2 (N20238, N20234, N5106);
nor NOR4 (N20239, N20220, N13487, N9916, N7202);
or OR3 (N20240, N20236, N8100, N13699);
and AND3 (N20241, N20205, N3464, N4969);
nor NOR2 (N20242, N20231, N12400);
and AND2 (N20243, N20241, N15728);
not NOT1 (N20244, N20243);
nand NAND4 (N20245, N20225, N8373, N15453, N12192);
or OR2 (N20246, N20233, N16004);
nand NAND4 (N20247, N20237, N5369, N13172, N4322);
xor XOR2 (N20248, N20247, N13163);
xor XOR2 (N20249, N20238, N15184);
and AND3 (N20250, N20235, N19723, N6719);
and AND3 (N20251, N20229, N1236, N20145);
xor XOR2 (N20252, N20249, N5174);
xor XOR2 (N20253, N20251, N5703);
nor NOR4 (N20254, N20246, N10770, N12560, N14459);
nand NAND4 (N20255, N20242, N11236, N660, N12417);
and AND3 (N20256, N20244, N16635, N12219);
buf BUF1 (N20257, N20245);
xor XOR2 (N20258, N20253, N1963);
and AND2 (N20259, N20255, N1465);
buf BUF1 (N20260, N20252);
and AND4 (N20261, N20254, N9673, N4618, N5998);
not NOT1 (N20262, N20261);
and AND2 (N20263, N20250, N3744);
xor XOR2 (N20264, N20240, N4516);
buf BUF1 (N20265, N20264);
nor NOR3 (N20266, N20259, N10359, N9232);
and AND2 (N20267, N20256, N6405);
xor XOR2 (N20268, N20258, N12987);
xor XOR2 (N20269, N20265, N18389);
not NOT1 (N20270, N20239);
nor NOR4 (N20271, N20260, N13406, N1993, N11928);
nand NAND3 (N20272, N20263, N14888, N17136);
nand NAND4 (N20273, N20266, N17680, N14376, N11134);
or OR4 (N20274, N20273, N9455, N8317, N6848);
buf BUF1 (N20275, N20274);
xor XOR2 (N20276, N20248, N11670);
xor XOR2 (N20277, N20269, N20226);
buf BUF1 (N20278, N20267);
nand NAND3 (N20279, N20278, N15997, N19536);
or OR3 (N20280, N20276, N8623, N1386);
or OR3 (N20281, N20262, N6202, N18461);
nor NOR3 (N20282, N20271, N12522, N10232);
not NOT1 (N20283, N20257);
buf BUF1 (N20284, N20272);
nor NOR4 (N20285, N20284, N11642, N10737, N5433);
and AND2 (N20286, N20285, N19029);
or OR4 (N20287, N20280, N3230, N4295, N13918);
nand NAND4 (N20288, N20275, N1118, N4452, N13406);
nand NAND2 (N20289, N20287, N5561);
or OR4 (N20290, N20288, N3316, N10112, N18113);
nor NOR3 (N20291, N20282, N8339, N6680);
xor XOR2 (N20292, N20291, N18909);
nor NOR2 (N20293, N20279, N5546);
or OR4 (N20294, N20270, N4067, N6182, N19595);
and AND4 (N20295, N20293, N3230, N12856, N15325);
nand NAND4 (N20296, N20294, N12795, N1200, N7508);
xor XOR2 (N20297, N20295, N5492);
not NOT1 (N20298, N20281);
or OR3 (N20299, N20292, N6928, N7982);
xor XOR2 (N20300, N20268, N17952);
and AND4 (N20301, N20296, N9552, N9932, N253);
and AND3 (N20302, N20301, N19184, N11107);
nand NAND4 (N20303, N20283, N11712, N20124, N15910);
or OR2 (N20304, N20298, N11324);
buf BUF1 (N20305, N20303);
buf BUF1 (N20306, N20299);
and AND2 (N20307, N20290, N14800);
buf BUF1 (N20308, N20307);
nor NOR2 (N20309, N20306, N6298);
not NOT1 (N20310, N20289);
buf BUF1 (N20311, N20304);
and AND4 (N20312, N20310, N5420, N480, N14329);
xor XOR2 (N20313, N20312, N11831);
or OR2 (N20314, N20300, N9241);
xor XOR2 (N20315, N20314, N1913);
nor NOR3 (N20316, N20313, N16827, N1763);
buf BUF1 (N20317, N20316);
xor XOR2 (N20318, N20297, N131);
and AND2 (N20319, N20302, N18007);
xor XOR2 (N20320, N20319, N40);
and AND4 (N20321, N20318, N10573, N8934, N1735);
or OR3 (N20322, N20321, N18274, N17270);
or OR4 (N20323, N20277, N15885, N2130, N2293);
xor XOR2 (N20324, N20322, N7940);
xor XOR2 (N20325, N20324, N5672);
xor XOR2 (N20326, N20305, N8437);
xor XOR2 (N20327, N20317, N17812);
and AND3 (N20328, N20327, N1026, N6000);
nand NAND3 (N20329, N20323, N17310, N2504);
nand NAND3 (N20330, N20315, N12148, N3170);
or OR3 (N20331, N20286, N19712, N14197);
or OR2 (N20332, N20331, N3491);
xor XOR2 (N20333, N20328, N3445);
not NOT1 (N20334, N20311);
nand NAND3 (N20335, N20329, N10173, N2627);
buf BUF1 (N20336, N20332);
and AND4 (N20337, N20309, N8862, N14060, N16802);
nand NAND2 (N20338, N20325, N7093);
not NOT1 (N20339, N20320);
xor XOR2 (N20340, N20326, N2811);
and AND2 (N20341, N20335, N16041);
xor XOR2 (N20342, N20337, N18924);
xor XOR2 (N20343, N20339, N8980);
nor NOR3 (N20344, N20343, N4132, N3778);
nor NOR3 (N20345, N20344, N9539, N15239);
and AND4 (N20346, N20341, N13034, N130, N18591);
not NOT1 (N20347, N20334);
nand NAND3 (N20348, N20347, N15951, N7512);
nor NOR3 (N20349, N20342, N11634, N16937);
and AND3 (N20350, N20346, N8465, N16139);
and AND3 (N20351, N20345, N10232, N8839);
nor NOR4 (N20352, N20351, N7892, N5703, N15184);
nand NAND2 (N20353, N20340, N19754);
or OR2 (N20354, N20348, N14989);
nor NOR2 (N20355, N20354, N5437);
and AND4 (N20356, N20336, N17109, N18343, N15690);
buf BUF1 (N20357, N20333);
not NOT1 (N20358, N20350);
nand NAND2 (N20359, N20330, N2638);
not NOT1 (N20360, N20357);
nand NAND2 (N20361, N20359, N6184);
nor NOR4 (N20362, N20356, N1756, N17718, N1458);
and AND2 (N20363, N20349, N20201);
nand NAND3 (N20364, N20363, N15331, N8029);
and AND3 (N20365, N20352, N996, N8212);
xor XOR2 (N20366, N20361, N13881);
nand NAND3 (N20367, N20364, N18609, N7588);
xor XOR2 (N20368, N20358, N9152);
xor XOR2 (N20369, N20367, N17671);
buf BUF1 (N20370, N20365);
not NOT1 (N20371, N20308);
nor NOR4 (N20372, N20338, N8855, N11435, N8947);
xor XOR2 (N20373, N20353, N20064);
xor XOR2 (N20374, N20370, N19349);
and AND2 (N20375, N20374, N6401);
nand NAND2 (N20376, N20371, N16341);
and AND2 (N20377, N20376, N15316);
and AND3 (N20378, N20368, N19100, N20206);
nand NAND4 (N20379, N20375, N7871, N12526, N2843);
not NOT1 (N20380, N20377);
nand NAND2 (N20381, N20362, N16036);
xor XOR2 (N20382, N20369, N8779);
nor NOR4 (N20383, N20355, N5723, N14233, N17704);
nor NOR3 (N20384, N20372, N15236, N7525);
nor NOR3 (N20385, N20383, N866, N91);
and AND2 (N20386, N20380, N18678);
or OR3 (N20387, N20384, N10904, N19014);
nor NOR2 (N20388, N20382, N1864);
and AND2 (N20389, N20378, N9834);
not NOT1 (N20390, N20379);
buf BUF1 (N20391, N20387);
xor XOR2 (N20392, N20366, N13252);
xor XOR2 (N20393, N20388, N7509);
xor XOR2 (N20394, N20385, N4365);
and AND4 (N20395, N20360, N6597, N19317, N20313);
xor XOR2 (N20396, N20392, N15273);
or OR4 (N20397, N20389, N16346, N18397, N19234);
buf BUF1 (N20398, N20391);
nand NAND4 (N20399, N20393, N14665, N795, N1136);
and AND2 (N20400, N20395, N11706);
not NOT1 (N20401, N20400);
nand NAND2 (N20402, N20399, N17375);
buf BUF1 (N20403, N20397);
and AND4 (N20404, N20403, N13366, N2258, N3084);
xor XOR2 (N20405, N20398, N6354);
nor NOR3 (N20406, N20394, N18136, N2636);
xor XOR2 (N20407, N20402, N6802);
not NOT1 (N20408, N20386);
buf BUF1 (N20409, N20404);
buf BUF1 (N20410, N20390);
or OR4 (N20411, N20396, N5049, N14183, N19551);
buf BUF1 (N20412, N20406);
not NOT1 (N20413, N20401);
xor XOR2 (N20414, N20412, N11984);
or OR2 (N20415, N20408, N10584);
xor XOR2 (N20416, N20405, N19411);
and AND2 (N20417, N20409, N17562);
or OR3 (N20418, N20415, N8465, N10151);
xor XOR2 (N20419, N20416, N9735);
xor XOR2 (N20420, N20419, N3632);
not NOT1 (N20421, N20414);
buf BUF1 (N20422, N20373);
not NOT1 (N20423, N20417);
nor NOR4 (N20424, N20418, N4781, N18982, N2425);
nand NAND4 (N20425, N20424, N14477, N12072, N17364);
and AND4 (N20426, N20381, N5488, N2565, N9612);
and AND3 (N20427, N20421, N5027, N16018);
not NOT1 (N20428, N20426);
and AND3 (N20429, N20420, N1001, N8929);
nor NOR3 (N20430, N20413, N18546, N2797);
and AND2 (N20431, N20410, N4802);
nor NOR4 (N20432, N20411, N16495, N9541, N13217);
nand NAND2 (N20433, N20428, N2283);
nor NOR2 (N20434, N20433, N3350);
xor XOR2 (N20435, N20432, N11151);
nand NAND2 (N20436, N20430, N1687);
and AND3 (N20437, N20425, N819, N14823);
nor NOR3 (N20438, N20436, N14054, N7376);
xor XOR2 (N20439, N20437, N12325);
buf BUF1 (N20440, N20438);
nor NOR4 (N20441, N20439, N2707, N13686, N5507);
nand NAND3 (N20442, N20431, N12074, N18224);
nand NAND3 (N20443, N20435, N8852, N11876);
nand NAND2 (N20444, N20423, N17215);
not NOT1 (N20445, N20442);
or OR4 (N20446, N20429, N12168, N9018, N6349);
or OR3 (N20447, N20445, N13924, N3320);
nor NOR4 (N20448, N20434, N10305, N10329, N11142);
nand NAND4 (N20449, N20447, N4416, N3754, N19841);
and AND2 (N20450, N20448, N535);
buf BUF1 (N20451, N20446);
nand NAND4 (N20452, N20441, N7737, N15308, N4795);
nand NAND2 (N20453, N20451, N6962);
nor NOR4 (N20454, N20427, N20010, N12474, N1594);
and AND4 (N20455, N20453, N12518, N260, N7356);
or OR4 (N20456, N20452, N14026, N1250, N9411);
buf BUF1 (N20457, N20440);
nor NOR2 (N20458, N20454, N7715);
not NOT1 (N20459, N20444);
and AND3 (N20460, N20459, N712, N20141);
xor XOR2 (N20461, N20456, N18435);
nand NAND2 (N20462, N20458, N9154);
xor XOR2 (N20463, N20450, N16591);
nand NAND3 (N20464, N20455, N3822, N19486);
buf BUF1 (N20465, N20460);
not NOT1 (N20466, N20465);
xor XOR2 (N20467, N20463, N10328);
xor XOR2 (N20468, N20462, N96);
nand NAND3 (N20469, N20468, N7496, N19622);
not NOT1 (N20470, N20407);
nor NOR3 (N20471, N20422, N18393, N19080);
nor NOR3 (N20472, N20457, N14293, N20060);
nor NOR3 (N20473, N20469, N16845, N17968);
nand NAND3 (N20474, N20449, N3152, N11899);
nor NOR2 (N20475, N20466, N15560);
nor NOR3 (N20476, N20474, N18768, N3480);
or OR2 (N20477, N20461, N1432);
xor XOR2 (N20478, N20476, N8617);
or OR3 (N20479, N20475, N9475, N14571);
nor NOR4 (N20480, N20471, N12281, N3638, N15072);
xor XOR2 (N20481, N20470, N12443);
nor NOR4 (N20482, N20467, N5647, N1033, N11847);
not NOT1 (N20483, N20480);
and AND3 (N20484, N20478, N3539, N13108);
nor NOR3 (N20485, N20482, N8885, N5882);
xor XOR2 (N20486, N20477, N11644);
and AND3 (N20487, N20484, N11830, N490);
nor NOR2 (N20488, N20486, N5123);
or OR4 (N20489, N20485, N15107, N19510, N17608);
or OR3 (N20490, N20473, N3344, N13464);
nor NOR2 (N20491, N20464, N3506);
buf BUF1 (N20492, N20491);
or OR3 (N20493, N20487, N3677, N17301);
xor XOR2 (N20494, N20492, N5124);
or OR2 (N20495, N20483, N8930);
and AND2 (N20496, N20479, N10269);
nor NOR2 (N20497, N20488, N12525);
buf BUF1 (N20498, N20481);
nor NOR3 (N20499, N20498, N8728, N284);
buf BUF1 (N20500, N20489);
nor NOR4 (N20501, N20497, N2940, N11892, N9507);
nand NAND2 (N20502, N20493, N5939);
xor XOR2 (N20503, N20502, N7418);
or OR4 (N20504, N20503, N1731, N17705, N13432);
and AND4 (N20505, N20496, N16356, N2356, N9511);
or OR2 (N20506, N20499, N2994);
or OR4 (N20507, N20495, N19287, N13852, N2375);
and AND2 (N20508, N20494, N18550);
xor XOR2 (N20509, N20500, N11902);
and AND3 (N20510, N20490, N1115, N9291);
nor NOR2 (N20511, N20472, N11618);
xor XOR2 (N20512, N20443, N9518);
not NOT1 (N20513, N20507);
xor XOR2 (N20514, N20505, N5468);
and AND4 (N20515, N20504, N14243, N2960, N14981);
not NOT1 (N20516, N20515);
buf BUF1 (N20517, N20513);
and AND3 (N20518, N20516, N10978, N19041);
xor XOR2 (N20519, N20518, N1280);
or OR3 (N20520, N20517, N12976, N17528);
buf BUF1 (N20521, N20501);
xor XOR2 (N20522, N20508, N5012);
nor NOR3 (N20523, N20522, N12369, N10754);
or OR3 (N20524, N20523, N795, N19102);
buf BUF1 (N20525, N20509);
or OR2 (N20526, N20521, N4303);
buf BUF1 (N20527, N20510);
buf BUF1 (N20528, N20506);
not NOT1 (N20529, N20519);
nor NOR4 (N20530, N20526, N8863, N5109, N13532);
xor XOR2 (N20531, N20527, N11133);
buf BUF1 (N20532, N20531);
not NOT1 (N20533, N20524);
xor XOR2 (N20534, N20530, N930);
nand NAND2 (N20535, N20514, N233);
nand NAND2 (N20536, N20511, N19205);
not NOT1 (N20537, N20528);
xor XOR2 (N20538, N20533, N202);
nor NOR4 (N20539, N20532, N3244, N6516, N7586);
xor XOR2 (N20540, N20538, N16619);
and AND3 (N20541, N20536, N12128, N13646);
not NOT1 (N20542, N20520);
and AND4 (N20543, N20512, N8482, N17071, N347);
nand NAND4 (N20544, N20540, N11828, N13864, N17484);
nand NAND3 (N20545, N20544, N20132, N15699);
nand NAND4 (N20546, N20539, N14950, N19914, N1488);
xor XOR2 (N20547, N20541, N3784);
buf BUF1 (N20548, N20542);
or OR4 (N20549, N20546, N4660, N1756, N3356);
not NOT1 (N20550, N20534);
and AND3 (N20551, N20547, N19887, N10470);
or OR2 (N20552, N20535, N3668);
nand NAND4 (N20553, N20529, N5128, N15194, N5399);
and AND2 (N20554, N20537, N16388);
not NOT1 (N20555, N20525);
xor XOR2 (N20556, N20548, N6924);
nand NAND4 (N20557, N20550, N6544, N3143, N5940);
or OR3 (N20558, N20543, N11638, N13704);
buf BUF1 (N20559, N20545);
or OR4 (N20560, N20551, N5385, N15608, N2105);
not NOT1 (N20561, N20555);
not NOT1 (N20562, N20556);
xor XOR2 (N20563, N20552, N18459);
and AND4 (N20564, N20562, N19980, N14150, N3684);
nor NOR2 (N20565, N20557, N9277);
nor NOR4 (N20566, N20559, N13478, N1779, N9597);
and AND2 (N20567, N20554, N2142);
nor NOR2 (N20568, N20558, N9529);
nand NAND4 (N20569, N20561, N15685, N10924, N6276);
nor NOR2 (N20570, N20549, N8738);
nand NAND4 (N20571, N20553, N18729, N2500, N16118);
or OR2 (N20572, N20564, N7721);
and AND3 (N20573, N20566, N7107, N20517);
buf BUF1 (N20574, N20568);
not NOT1 (N20575, N20569);
and AND3 (N20576, N20563, N2729, N15222);
nor NOR2 (N20577, N20570, N17768);
nand NAND3 (N20578, N20577, N2360, N3105);
xor XOR2 (N20579, N20572, N10661);
buf BUF1 (N20580, N20574);
not NOT1 (N20581, N20571);
not NOT1 (N20582, N20575);
nand NAND3 (N20583, N20560, N8054, N11451);
nand NAND3 (N20584, N20576, N10206, N17977);
nand NAND2 (N20585, N20580, N16761);
xor XOR2 (N20586, N20582, N4407);
or OR3 (N20587, N20567, N16923, N20295);
and AND4 (N20588, N20581, N14357, N12391, N8165);
nand NAND2 (N20589, N20588, N4798);
not NOT1 (N20590, N20589);
buf BUF1 (N20591, N20579);
nor NOR3 (N20592, N20584, N11326, N20530);
and AND3 (N20593, N20586, N2483, N16437);
xor XOR2 (N20594, N20587, N18165);
not NOT1 (N20595, N20565);
buf BUF1 (N20596, N20593);
nor NOR4 (N20597, N20578, N5818, N12161, N15852);
or OR4 (N20598, N20591, N6904, N16168, N18203);
or OR2 (N20599, N20597, N4241);
nor NOR3 (N20600, N20585, N16660, N9940);
xor XOR2 (N20601, N20599, N16590);
buf BUF1 (N20602, N20600);
not NOT1 (N20603, N20598);
not NOT1 (N20604, N20583);
and AND3 (N20605, N20601, N11474, N15900);
or OR2 (N20606, N20594, N624);
nand NAND2 (N20607, N20590, N13981);
not NOT1 (N20608, N20592);
nand NAND2 (N20609, N20604, N10205);
nor NOR4 (N20610, N20573, N14385, N3736, N9889);
or OR2 (N20611, N20605, N6832);
and AND3 (N20612, N20606, N14347, N17905);
xor XOR2 (N20613, N20609, N5471);
xor XOR2 (N20614, N20603, N15536);
or OR2 (N20615, N20611, N16707);
nor NOR2 (N20616, N20612, N271);
buf BUF1 (N20617, N20613);
and AND4 (N20618, N20607, N18539, N10644, N13627);
nor NOR4 (N20619, N20608, N4405, N7827, N20334);
or OR4 (N20620, N20595, N9113, N4593, N3434);
buf BUF1 (N20621, N20615);
and AND4 (N20622, N20616, N1008, N8614, N483);
xor XOR2 (N20623, N20610, N12411);
xor XOR2 (N20624, N20622, N5824);
or OR4 (N20625, N20596, N12702, N19278, N18593);
buf BUF1 (N20626, N20621);
buf BUF1 (N20627, N20624);
or OR4 (N20628, N20618, N5693, N4054, N3110);
and AND4 (N20629, N20623, N11183, N15651, N9256);
xor XOR2 (N20630, N20614, N15188);
or OR2 (N20631, N20619, N18479);
nor NOR2 (N20632, N20602, N3083);
not NOT1 (N20633, N20630);
nor NOR3 (N20634, N20632, N12004, N290);
nor NOR3 (N20635, N20625, N19948, N2355);
buf BUF1 (N20636, N20627);
nand NAND3 (N20637, N20617, N3750, N844);
not NOT1 (N20638, N20636);
xor XOR2 (N20639, N20628, N6116);
nor NOR3 (N20640, N20634, N16362, N17041);
and AND4 (N20641, N20637, N8970, N13106, N9744);
nor NOR3 (N20642, N20620, N18590, N3430);
buf BUF1 (N20643, N20638);
nand NAND2 (N20644, N20642, N19022);
nor NOR3 (N20645, N20626, N17749, N1720);
and AND4 (N20646, N20641, N20064, N19097, N20156);
xor XOR2 (N20647, N20644, N17056);
not NOT1 (N20648, N20646);
and AND4 (N20649, N20635, N11117, N6231, N5487);
xor XOR2 (N20650, N20649, N5839);
or OR4 (N20651, N20633, N9918, N17481, N15272);
buf BUF1 (N20652, N20645);
buf BUF1 (N20653, N20643);
buf BUF1 (N20654, N20650);
buf BUF1 (N20655, N20639);
nand NAND3 (N20656, N20653, N14572, N12535);
xor XOR2 (N20657, N20640, N4753);
buf BUF1 (N20658, N20656);
buf BUF1 (N20659, N20629);
xor XOR2 (N20660, N20659, N13023);
not NOT1 (N20661, N20657);
or OR3 (N20662, N20655, N19264, N837);
not NOT1 (N20663, N20651);
not NOT1 (N20664, N20652);
xor XOR2 (N20665, N20664, N12659);
nand NAND4 (N20666, N20662, N7551, N6156, N3916);
buf BUF1 (N20667, N20654);
buf BUF1 (N20668, N20663);
xor XOR2 (N20669, N20668, N5167);
or OR3 (N20670, N20660, N8094, N9400);
and AND2 (N20671, N20658, N6879);
or OR4 (N20672, N20661, N10183, N14126, N20573);
and AND3 (N20673, N20647, N17176, N2374);
or OR4 (N20674, N20648, N17066, N12988, N20134);
and AND2 (N20675, N20674, N1587);
and AND2 (N20676, N20631, N10843);
or OR4 (N20677, N20667, N683, N267, N18557);
buf BUF1 (N20678, N20676);
nand NAND3 (N20679, N20673, N18625, N14379);
nand NAND2 (N20680, N20672, N6320);
xor XOR2 (N20681, N20679, N14871);
xor XOR2 (N20682, N20666, N3580);
not NOT1 (N20683, N20677);
nor NOR3 (N20684, N20680, N6517, N12877);
buf BUF1 (N20685, N20684);
nor NOR4 (N20686, N20678, N16982, N1189, N6702);
nand NAND3 (N20687, N20682, N20428, N9079);
and AND2 (N20688, N20685, N4629);
buf BUF1 (N20689, N20671);
and AND2 (N20690, N20687, N4373);
buf BUF1 (N20691, N20683);
nor NOR2 (N20692, N20675, N4427);
not NOT1 (N20693, N20686);
or OR2 (N20694, N20693, N7848);
not NOT1 (N20695, N20691);
nand NAND2 (N20696, N20665, N19782);
or OR2 (N20697, N20694, N15412);
or OR2 (N20698, N20690, N11771);
nand NAND3 (N20699, N20696, N559, N16149);
xor XOR2 (N20700, N20688, N7481);
and AND4 (N20701, N20697, N11867, N11919, N13896);
nor NOR3 (N20702, N20698, N19399, N2593);
xor XOR2 (N20703, N20701, N889);
nor NOR3 (N20704, N20703, N11365, N3657);
and AND3 (N20705, N20704, N5003, N5310);
nor NOR4 (N20706, N20669, N18361, N6743, N3051);
xor XOR2 (N20707, N20670, N4348);
buf BUF1 (N20708, N20689);
and AND2 (N20709, N20702, N3054);
not NOT1 (N20710, N20695);
buf BUF1 (N20711, N20706);
nor NOR3 (N20712, N20705, N17577, N15166);
xor XOR2 (N20713, N20708, N7929);
xor XOR2 (N20714, N20709, N1540);
xor XOR2 (N20715, N20707, N18014);
xor XOR2 (N20716, N20692, N9035);
nor NOR4 (N20717, N20681, N1510, N4620, N99);
buf BUF1 (N20718, N20715);
and AND3 (N20719, N20711, N14606, N6921);
xor XOR2 (N20720, N20718, N18638);
or OR2 (N20721, N20700, N18646);
nand NAND4 (N20722, N20716, N16306, N2203, N13976);
and AND4 (N20723, N20714, N13337, N12933, N11368);
not NOT1 (N20724, N20699);
and AND4 (N20725, N20713, N18275, N8082, N7712);
nor NOR4 (N20726, N20723, N6112, N446, N10354);
nand NAND2 (N20727, N20724, N15264);
buf BUF1 (N20728, N20727);
nor NOR4 (N20729, N20722, N14139, N17218, N2201);
or OR2 (N20730, N20717, N17656);
or OR2 (N20731, N20725, N15385);
nand NAND4 (N20732, N20712, N17195, N14664, N16930);
buf BUF1 (N20733, N20719);
not NOT1 (N20734, N20732);
and AND3 (N20735, N20720, N8076, N16163);
or OR2 (N20736, N20726, N7);
buf BUF1 (N20737, N20730);
and AND4 (N20738, N20736, N3006, N11975, N2035);
not NOT1 (N20739, N20710);
xor XOR2 (N20740, N20721, N16023);
or OR4 (N20741, N20733, N16766, N5534, N14219);
not NOT1 (N20742, N20741);
buf BUF1 (N20743, N20728);
and AND4 (N20744, N20742, N20579, N19590, N16290);
buf BUF1 (N20745, N20731);
nor NOR4 (N20746, N20734, N10439, N5847, N18503);
xor XOR2 (N20747, N20735, N950);
buf BUF1 (N20748, N20747);
nand NAND3 (N20749, N20739, N20425, N9841);
xor XOR2 (N20750, N20737, N4469);
buf BUF1 (N20751, N20729);
nor NOR2 (N20752, N20749, N14913);
xor XOR2 (N20753, N20740, N1675);
or OR2 (N20754, N20748, N19184);
xor XOR2 (N20755, N20743, N8713);
and AND3 (N20756, N20738, N19914, N10681);
or OR3 (N20757, N20753, N8438, N4123);
or OR3 (N20758, N20755, N8044, N2687);
and AND2 (N20759, N20751, N12550);
xor XOR2 (N20760, N20759, N7047);
nand NAND3 (N20761, N20760, N14598, N7945);
xor XOR2 (N20762, N20746, N20214);
nand NAND4 (N20763, N20762, N3134, N6041, N10858);
nor NOR2 (N20764, N20763, N12376);
not NOT1 (N20765, N20745);
nor NOR4 (N20766, N20757, N11488, N15060, N369);
and AND2 (N20767, N20754, N2240);
or OR2 (N20768, N20744, N10573);
nand NAND4 (N20769, N20765, N20073, N7046, N10698);
or OR2 (N20770, N20758, N14760);
or OR2 (N20771, N20766, N15161);
nand NAND3 (N20772, N20771, N10134, N500);
and AND2 (N20773, N20750, N16649);
and AND2 (N20774, N20768, N16031);
nor NOR3 (N20775, N20770, N19367, N12929);
nand NAND3 (N20776, N20774, N11746, N7862);
buf BUF1 (N20777, N20767);
not NOT1 (N20778, N20775);
nand NAND3 (N20779, N20761, N8148, N3135);
buf BUF1 (N20780, N20779);
nand NAND4 (N20781, N20769, N13730, N9616, N7350);
nand NAND3 (N20782, N20780, N13043, N13631);
nand NAND3 (N20783, N20773, N18551, N15511);
not NOT1 (N20784, N20777);
and AND3 (N20785, N20756, N15392, N9532);
xor XOR2 (N20786, N20778, N12373);
xor XOR2 (N20787, N20783, N16105);
xor XOR2 (N20788, N20776, N6528);
buf BUF1 (N20789, N20764);
nand NAND3 (N20790, N20752, N19557, N12142);
nor NOR4 (N20791, N20785, N11370, N13586, N14752);
or OR2 (N20792, N20790, N14213);
buf BUF1 (N20793, N20792);
buf BUF1 (N20794, N20782);
and AND4 (N20795, N20772, N14241, N12479, N3138);
xor XOR2 (N20796, N20784, N12636);
nor NOR4 (N20797, N20787, N3057, N17746, N17181);
xor XOR2 (N20798, N20796, N7388);
or OR3 (N20799, N20781, N12006, N16451);
or OR2 (N20800, N20797, N15599);
buf BUF1 (N20801, N20791);
not NOT1 (N20802, N20801);
nor NOR4 (N20803, N20793, N6121, N1015, N4941);
or OR3 (N20804, N20799, N3752, N13063);
nand NAND2 (N20805, N20794, N15824);
nand NAND2 (N20806, N20786, N12189);
and AND4 (N20807, N20802, N8534, N8449, N15325);
nand NAND4 (N20808, N20795, N12365, N12849, N10257);
xor XOR2 (N20809, N20803, N17749);
nand NAND4 (N20810, N20789, N8383, N14904, N2579);
not NOT1 (N20811, N20809);
xor XOR2 (N20812, N20800, N11120);
not NOT1 (N20813, N20788);
nand NAND3 (N20814, N20811, N8693, N1169);
buf BUF1 (N20815, N20805);
not NOT1 (N20816, N20813);
nor NOR4 (N20817, N20816, N8986, N4105, N19332);
xor XOR2 (N20818, N20814, N11108);
not NOT1 (N20819, N20808);
buf BUF1 (N20820, N20798);
or OR3 (N20821, N20806, N20646, N3312);
not NOT1 (N20822, N20815);
buf BUF1 (N20823, N20818);
nand NAND4 (N20824, N20804, N11267, N4621, N1817);
nor NOR2 (N20825, N20807, N3146);
nor NOR2 (N20826, N20822, N19127);
and AND4 (N20827, N20819, N6102, N2501, N853);
buf BUF1 (N20828, N20823);
or OR2 (N20829, N20820, N10231);
not NOT1 (N20830, N20821);
nand NAND4 (N20831, N20810, N3263, N15755, N2636);
xor XOR2 (N20832, N20817, N14731);
xor XOR2 (N20833, N20826, N10053);
nand NAND3 (N20834, N20831, N223, N17885);
not NOT1 (N20835, N20829);
xor XOR2 (N20836, N20825, N10545);
nand NAND3 (N20837, N20828, N12624, N4909);
nand NAND4 (N20838, N20830, N16445, N18476, N3625);
nor NOR3 (N20839, N20812, N10020, N12561);
nor NOR2 (N20840, N20824, N1130);
and AND2 (N20841, N20839, N4672);
nor NOR4 (N20842, N20833, N9771, N9560, N16714);
nand NAND2 (N20843, N20834, N11328);
buf BUF1 (N20844, N20840);
buf BUF1 (N20845, N20827);
or OR3 (N20846, N20842, N992, N4765);
and AND3 (N20847, N20832, N9392, N20286);
and AND4 (N20848, N20838, N5474, N20497, N19271);
nand NAND4 (N20849, N20843, N12447, N5290, N2493);
nand NAND2 (N20850, N20841, N13954);
nand NAND4 (N20851, N20850, N8733, N14443, N2317);
nor NOR4 (N20852, N20847, N15794, N6429, N1563);
or OR3 (N20853, N20836, N432, N6973);
buf BUF1 (N20854, N20845);
buf BUF1 (N20855, N20848);
buf BUF1 (N20856, N20851);
or OR4 (N20857, N20854, N16889, N13724, N4065);
and AND3 (N20858, N20856, N14489, N20618);
xor XOR2 (N20859, N20846, N17983);
buf BUF1 (N20860, N20852);
and AND2 (N20861, N20844, N14835);
xor XOR2 (N20862, N20853, N7200);
not NOT1 (N20863, N20861);
buf BUF1 (N20864, N20849);
and AND2 (N20865, N20859, N9806);
and AND2 (N20866, N20862, N11646);
and AND3 (N20867, N20835, N20572, N4598);
nand NAND2 (N20868, N20857, N1546);
not NOT1 (N20869, N20863);
buf BUF1 (N20870, N20869);
and AND2 (N20871, N20858, N10337);
or OR4 (N20872, N20871, N11213, N932, N12981);
buf BUF1 (N20873, N20865);
nand NAND3 (N20874, N20872, N2543, N4669);
or OR2 (N20875, N20873, N4265);
nand NAND3 (N20876, N20870, N4833, N11525);
xor XOR2 (N20877, N20860, N6572);
nand NAND4 (N20878, N20876, N6856, N6543, N1361);
xor XOR2 (N20879, N20867, N14047);
nand NAND4 (N20880, N20875, N20212, N19719, N14055);
xor XOR2 (N20881, N20879, N13939);
or OR2 (N20882, N20864, N8555);
and AND2 (N20883, N20878, N19886);
xor XOR2 (N20884, N20868, N11291);
not NOT1 (N20885, N20883);
nand NAND3 (N20886, N20884, N15967, N19525);
nand NAND2 (N20887, N20877, N4943);
nand NAND3 (N20888, N20881, N9532, N2756);
nor NOR3 (N20889, N20885, N9656, N11485);
not NOT1 (N20890, N20837);
or OR2 (N20891, N20882, N351);
nand NAND4 (N20892, N20887, N14620, N9763, N7767);
buf BUF1 (N20893, N20886);
or OR2 (N20894, N20890, N20356);
not NOT1 (N20895, N20892);
nand NAND3 (N20896, N20874, N3210, N19468);
nand NAND3 (N20897, N20893, N18718, N503);
nor NOR4 (N20898, N20896, N6090, N6579, N20862);
and AND3 (N20899, N20897, N3178, N678);
nor NOR4 (N20900, N20898, N10003, N2918, N8481);
xor XOR2 (N20901, N20866, N10495);
xor XOR2 (N20902, N20899, N6447);
or OR2 (N20903, N20901, N12087);
nand NAND2 (N20904, N20855, N823);
or OR2 (N20905, N20895, N13328);
or OR2 (N20906, N20891, N6381);
nor NOR4 (N20907, N20906, N11436, N7140, N1886);
nand NAND2 (N20908, N20900, N10325);
or OR2 (N20909, N20905, N15570);
or OR2 (N20910, N20904, N20433);
not NOT1 (N20911, N20902);
not NOT1 (N20912, N20908);
xor XOR2 (N20913, N20911, N16523);
or OR2 (N20914, N20909, N19790);
or OR3 (N20915, N20888, N19643, N14737);
xor XOR2 (N20916, N20915, N2441);
buf BUF1 (N20917, N20903);
buf BUF1 (N20918, N20914);
nor NOR3 (N20919, N20894, N3428, N13160);
not NOT1 (N20920, N20910);
nor NOR4 (N20921, N20913, N20249, N13365, N20514);
or OR4 (N20922, N20907, N13306, N11761, N11437);
buf BUF1 (N20923, N20922);
nor NOR4 (N20924, N20920, N12577, N1673, N8201);
nand NAND2 (N20925, N20921, N9305);
and AND3 (N20926, N20918, N3317, N3275);
nor NOR3 (N20927, N20925, N5884, N15882);
xor XOR2 (N20928, N20917, N15883);
and AND2 (N20929, N20880, N6031);
buf BUF1 (N20930, N20928);
xor XOR2 (N20931, N20927, N18731);
and AND4 (N20932, N20926, N20559, N7864, N20558);
nand NAND4 (N20933, N20932, N15746, N14397, N272);
and AND4 (N20934, N20889, N1386, N15606, N123);
not NOT1 (N20935, N20924);
nor NOR4 (N20936, N20934, N911, N7637, N1426);
buf BUF1 (N20937, N20936);
buf BUF1 (N20938, N20916);
not NOT1 (N20939, N20929);
and AND4 (N20940, N20939, N1839, N9914, N16352);
and AND2 (N20941, N20912, N16897);
nand NAND2 (N20942, N20923, N6806);
nor NOR3 (N20943, N20935, N901, N11762);
xor XOR2 (N20944, N20943, N13605);
or OR3 (N20945, N20938, N6922, N4434);
xor XOR2 (N20946, N20933, N19924);
nand NAND4 (N20947, N20930, N11275, N15409, N16817);
xor XOR2 (N20948, N20941, N18711);
or OR3 (N20949, N20940, N19848, N3210);
or OR4 (N20950, N20948, N9441, N19232, N551);
xor XOR2 (N20951, N20931, N5284);
buf BUF1 (N20952, N20942);
xor XOR2 (N20953, N20951, N19848);
nand NAND3 (N20954, N20937, N11986, N10436);
and AND3 (N20955, N20950, N18252, N12267);
nand NAND2 (N20956, N20919, N13952);
or OR3 (N20957, N20945, N16056, N14715);
not NOT1 (N20958, N20954);
nor NOR3 (N20959, N20946, N9622, N19179);
and AND2 (N20960, N20959, N10416);
nand NAND4 (N20961, N20949, N20607, N468, N20598);
buf BUF1 (N20962, N20953);
buf BUF1 (N20963, N20961);
and AND4 (N20964, N20962, N1385, N11181, N10346);
nand NAND2 (N20965, N20960, N10692);
or OR2 (N20966, N20957, N5622);
xor XOR2 (N20967, N20955, N6490);
not NOT1 (N20968, N20967);
buf BUF1 (N20969, N20965);
not NOT1 (N20970, N20964);
or OR2 (N20971, N20966, N15356);
not NOT1 (N20972, N20963);
nor NOR3 (N20973, N20956, N9070, N2584);
or OR4 (N20974, N20971, N6692, N149, N9276);
or OR2 (N20975, N20958, N20145);
not NOT1 (N20976, N20947);
nor NOR2 (N20977, N20976, N1280);
xor XOR2 (N20978, N20952, N15297);
or OR2 (N20979, N20978, N10669);
nor NOR2 (N20980, N20970, N1197);
xor XOR2 (N20981, N20979, N9918);
nor NOR4 (N20982, N20981, N4279, N12817, N5475);
xor XOR2 (N20983, N20980, N7682);
nand NAND2 (N20984, N20973, N18558);
nand NAND2 (N20985, N20944, N5675);
nor NOR4 (N20986, N20968, N2627, N1246, N3682);
xor XOR2 (N20987, N20969, N8833);
not NOT1 (N20988, N20972);
nand NAND3 (N20989, N20982, N18263, N11685);
nand NAND2 (N20990, N20975, N4654);
buf BUF1 (N20991, N20988);
nor NOR3 (N20992, N20991, N286, N6336);
buf BUF1 (N20993, N20984);
or OR2 (N20994, N20992, N12425);
xor XOR2 (N20995, N20987, N19729);
xor XOR2 (N20996, N20990, N2828);
nand NAND2 (N20997, N20977, N13321);
xor XOR2 (N20998, N20989, N5761);
nor NOR4 (N20999, N20996, N2865, N8060, N3372);
not NOT1 (N21000, N20985);
nor NOR4 (N21001, N20983, N19249, N13413, N11985);
not NOT1 (N21002, N20986);
and AND2 (N21003, N20995, N13276);
nand NAND4 (N21004, N21003, N2270, N19171, N14092);
and AND2 (N21005, N21004, N9463);
or OR3 (N21006, N20999, N3715, N13927);
buf BUF1 (N21007, N21006);
not NOT1 (N21008, N20974);
or OR3 (N21009, N20994, N20041, N19939);
buf BUF1 (N21010, N21001);
and AND2 (N21011, N20997, N20125);
xor XOR2 (N21012, N21002, N15637);
xor XOR2 (N21013, N21005, N14643);
xor XOR2 (N21014, N21010, N16462);
nand NAND4 (N21015, N21014, N8244, N15217, N13325);
or OR3 (N21016, N21015, N4769, N15410);
nand NAND4 (N21017, N21000, N14814, N9375, N5399);
nand NAND3 (N21018, N21011, N20632, N4402);
not NOT1 (N21019, N21007);
or OR3 (N21020, N21008, N17482, N1181);
xor XOR2 (N21021, N21012, N16488);
xor XOR2 (N21022, N21018, N11488);
or OR2 (N21023, N21013, N19723);
not NOT1 (N21024, N20993);
not NOT1 (N21025, N21016);
nor NOR4 (N21026, N21021, N9540, N7696, N17430);
or OR3 (N21027, N21024, N18777, N10175);
xor XOR2 (N21028, N21027, N1194);
or OR2 (N21029, N21028, N12434);
xor XOR2 (N21030, N21009, N15770);
nand NAND2 (N21031, N21023, N10646);
or OR3 (N21032, N21030, N5797, N16488);
buf BUF1 (N21033, N21022);
nor NOR3 (N21034, N21020, N8601, N6411);
not NOT1 (N21035, N21026);
and AND2 (N21036, N21025, N6324);
nor NOR2 (N21037, N21036, N13110);
or OR4 (N21038, N21019, N19330, N15205, N1598);
nor NOR3 (N21039, N21032, N5217, N20619);
nand NAND3 (N21040, N21035, N13950, N20077);
nor NOR3 (N21041, N21039, N212, N18210);
xor XOR2 (N21042, N21017, N18253);
and AND4 (N21043, N21037, N12642, N13245, N8226);
xor XOR2 (N21044, N21029, N17795);
nor NOR4 (N21045, N21043, N7192, N2432, N16338);
not NOT1 (N21046, N21044);
or OR3 (N21047, N21033, N18201, N12634);
buf BUF1 (N21048, N21031);
not NOT1 (N21049, N21038);
nor NOR3 (N21050, N21041, N19888, N3203);
buf BUF1 (N21051, N21048);
and AND2 (N21052, N21046, N11412);
not NOT1 (N21053, N21051);
not NOT1 (N21054, N21053);
and AND2 (N21055, N21042, N9820);
and AND2 (N21056, N21047, N6098);
nor NOR3 (N21057, N21049, N15950, N5193);
buf BUF1 (N21058, N21050);
or OR4 (N21059, N21057, N14889, N8859, N10493);
xor XOR2 (N21060, N21059, N1747);
not NOT1 (N21061, N21052);
buf BUF1 (N21062, N21054);
nand NAND2 (N21063, N21055, N8184);
buf BUF1 (N21064, N21058);
nand NAND4 (N21065, N21040, N19372, N16537, N9938);
xor XOR2 (N21066, N21045, N19300);
not NOT1 (N21067, N21061);
nand NAND2 (N21068, N21065, N19646);
buf BUF1 (N21069, N21056);
nor NOR2 (N21070, N20998, N11807);
xor XOR2 (N21071, N21063, N18822);
or OR2 (N21072, N21034, N5026);
buf BUF1 (N21073, N21060);
nand NAND2 (N21074, N21071, N11908);
not NOT1 (N21075, N21068);
not NOT1 (N21076, N21073);
buf BUF1 (N21077, N21074);
or OR3 (N21078, N21069, N14078, N11554);
and AND4 (N21079, N21062, N9547, N9938, N935);
nand NAND4 (N21080, N21076, N17167, N16057, N6426);
or OR2 (N21081, N21067, N5146);
xor XOR2 (N21082, N21080, N18120);
and AND2 (N21083, N21082, N12340);
nor NOR3 (N21084, N21079, N5990, N20893);
buf BUF1 (N21085, N21084);
xor XOR2 (N21086, N21085, N18246);
xor XOR2 (N21087, N21066, N13503);
and AND2 (N21088, N21083, N11085);
xor XOR2 (N21089, N21078, N10591);
nand NAND3 (N21090, N21087, N8608, N15644);
xor XOR2 (N21091, N21075, N6228);
nor NOR4 (N21092, N21064, N3740, N16394, N19728);
nor NOR2 (N21093, N21092, N16921);
or OR3 (N21094, N21081, N6618, N8190);
or OR2 (N21095, N21086, N9744);
buf BUF1 (N21096, N21093);
not NOT1 (N21097, N21072);
xor XOR2 (N21098, N21089, N5811);
xor XOR2 (N21099, N21070, N3262);
nand NAND2 (N21100, N21090, N16002);
buf BUF1 (N21101, N21095);
xor XOR2 (N21102, N21091, N10476);
nor NOR2 (N21103, N21100, N14820);
nand NAND4 (N21104, N21103, N2413, N16964, N7203);
buf BUF1 (N21105, N21077);
nand NAND4 (N21106, N21102, N16825, N13713, N3629);
nor NOR3 (N21107, N21088, N4268, N16589);
xor XOR2 (N21108, N21094, N10229);
and AND2 (N21109, N21107, N12478);
or OR4 (N21110, N21108, N15583, N19643, N5983);
buf BUF1 (N21111, N21096);
and AND4 (N21112, N21109, N10979, N7445, N13869);
and AND4 (N21113, N21104, N5979, N14746, N6025);
nor NOR2 (N21114, N21105, N15246);
buf BUF1 (N21115, N21110);
not NOT1 (N21116, N21101);
buf BUF1 (N21117, N21098);
xor XOR2 (N21118, N21114, N10135);
nand NAND3 (N21119, N21106, N12760, N13924);
nor NOR4 (N21120, N21097, N2487, N2077, N17628);
or OR3 (N21121, N21116, N18217, N17221);
buf BUF1 (N21122, N21099);
buf BUF1 (N21123, N21122);
nand NAND4 (N21124, N21112, N9344, N17215, N20427);
and AND4 (N21125, N21118, N7409, N7454, N15073);
nand NAND3 (N21126, N21111, N9422, N6771);
nand NAND4 (N21127, N21113, N19176, N14701, N12187);
and AND2 (N21128, N21124, N1139);
not NOT1 (N21129, N21126);
nand NAND3 (N21130, N21120, N6794, N11934);
and AND3 (N21131, N21129, N2638, N3746);
nor NOR2 (N21132, N21123, N19134);
nor NOR4 (N21133, N21131, N10735, N19690, N9066);
buf BUF1 (N21134, N21121);
nand NAND4 (N21135, N21125, N4661, N2596, N13424);
not NOT1 (N21136, N21127);
nand NAND4 (N21137, N21135, N4352, N4867, N17523);
nand NAND2 (N21138, N21115, N13925);
buf BUF1 (N21139, N21133);
or OR2 (N21140, N21139, N3882);
xor XOR2 (N21141, N21137, N12806);
or OR2 (N21142, N21138, N8652);
xor XOR2 (N21143, N21119, N2134);
or OR3 (N21144, N21141, N20342, N21097);
not NOT1 (N21145, N21132);
buf BUF1 (N21146, N21128);
not NOT1 (N21147, N21117);
or OR4 (N21148, N21140, N12690, N8300, N9160);
or OR4 (N21149, N21146, N7554, N14105, N8484);
not NOT1 (N21150, N21148);
nand NAND3 (N21151, N21130, N8126, N20872);
nand NAND4 (N21152, N21136, N18823, N7512, N14176);
nand NAND3 (N21153, N21142, N8069, N908);
nor NOR2 (N21154, N21145, N10179);
nand NAND4 (N21155, N21150, N7153, N17388, N5950);
nand NAND2 (N21156, N21155, N1969);
nand NAND2 (N21157, N21151, N7220);
and AND2 (N21158, N21153, N18797);
buf BUF1 (N21159, N21143);
and AND3 (N21160, N21157, N12811, N5684);
or OR3 (N21161, N21134, N10629, N3391);
not NOT1 (N21162, N21154);
nand NAND3 (N21163, N21156, N243, N7184);
nor NOR3 (N21164, N21162, N17295, N9968);
nand NAND4 (N21165, N21152, N12012, N9790, N14342);
or OR2 (N21166, N21149, N20461);
buf BUF1 (N21167, N21165);
xor XOR2 (N21168, N21164, N4913);
nand NAND2 (N21169, N21144, N10611);
xor XOR2 (N21170, N21168, N859);
nand NAND2 (N21171, N21167, N4532);
or OR3 (N21172, N21169, N18470, N18061);
xor XOR2 (N21173, N21161, N10467);
and AND3 (N21174, N21159, N6747, N8888);
buf BUF1 (N21175, N21147);
not NOT1 (N21176, N21175);
buf BUF1 (N21177, N21163);
and AND2 (N21178, N21170, N19975);
nand NAND4 (N21179, N21173, N13589, N5921, N2328);
nand NAND2 (N21180, N21177, N2192);
and AND3 (N21181, N21179, N11699, N19602);
not NOT1 (N21182, N21178);
and AND2 (N21183, N21171, N9696);
and AND3 (N21184, N21181, N3826, N11572);
buf BUF1 (N21185, N21172);
or OR4 (N21186, N21183, N11399, N18718, N1604);
nor NOR4 (N21187, N21182, N20619, N1201, N10194);
nand NAND4 (N21188, N21186, N14063, N17265, N19504);
xor XOR2 (N21189, N21174, N9986);
nand NAND4 (N21190, N21180, N10586, N17914, N4402);
or OR2 (N21191, N21188, N906);
not NOT1 (N21192, N21176);
nand NAND3 (N21193, N21166, N8888, N19663);
xor XOR2 (N21194, N21189, N4408);
nand NAND4 (N21195, N21191, N14729, N11077, N20164);
and AND2 (N21196, N21192, N12512);
buf BUF1 (N21197, N21190);
not NOT1 (N21198, N21196);
xor XOR2 (N21199, N21194, N2660);
and AND4 (N21200, N21193, N5031, N21174, N15525);
not NOT1 (N21201, N21160);
buf BUF1 (N21202, N21199);
nor NOR4 (N21203, N21158, N8780, N5277, N19029);
not NOT1 (N21204, N21185);
and AND4 (N21205, N21197, N11661, N11973, N16934);
and AND4 (N21206, N21202, N14038, N15763, N11482);
and AND4 (N21207, N21201, N11825, N7420, N6080);
buf BUF1 (N21208, N21195);
or OR2 (N21209, N21184, N9554);
and AND4 (N21210, N21200, N20663, N19912, N16233);
xor XOR2 (N21211, N21210, N10456);
nor NOR3 (N21212, N21187, N20889, N1044);
xor XOR2 (N21213, N21205, N7979);
nor NOR3 (N21214, N21198, N14607, N13643);
nand NAND3 (N21215, N21212, N10221, N6092);
nor NOR4 (N21216, N21208, N2345, N15370, N3452);
not NOT1 (N21217, N21203);
nand NAND4 (N21218, N21207, N2231, N12685, N6957);
xor XOR2 (N21219, N21215, N5846);
nand NAND4 (N21220, N21214, N8627, N19896, N3541);
and AND2 (N21221, N21211, N14927);
buf BUF1 (N21222, N21219);
or OR3 (N21223, N21218, N2802, N10145);
nand NAND4 (N21224, N21221, N16455, N2092, N17540);
and AND3 (N21225, N21224, N6179, N16477);
nand NAND2 (N21226, N21220, N2505);
and AND3 (N21227, N21216, N9275, N20821);
xor XOR2 (N21228, N21223, N12892);
buf BUF1 (N21229, N21222);
nor NOR2 (N21230, N21228, N2355);
and AND3 (N21231, N21225, N14649, N20004);
xor XOR2 (N21232, N21209, N9318);
and AND4 (N21233, N21230, N14072, N17957, N6690);
nand NAND4 (N21234, N21231, N2298, N19175, N12562);
not NOT1 (N21235, N21226);
buf BUF1 (N21236, N21227);
xor XOR2 (N21237, N21213, N6125);
nand NAND2 (N21238, N21235, N20649);
nand NAND2 (N21239, N21229, N14022);
buf BUF1 (N21240, N21233);
xor XOR2 (N21241, N21217, N915);
xor XOR2 (N21242, N21241, N18557);
and AND2 (N21243, N21242, N3253);
or OR2 (N21244, N21239, N18722);
nand NAND2 (N21245, N21240, N20688);
or OR4 (N21246, N21236, N3822, N6176, N8114);
not NOT1 (N21247, N21245);
nor NOR4 (N21248, N21232, N10186, N17144, N963);
not NOT1 (N21249, N21206);
not NOT1 (N21250, N21237);
nand NAND4 (N21251, N21249, N8426, N19773, N3411);
and AND3 (N21252, N21234, N17541, N783);
nor NOR4 (N21253, N21246, N21067, N1401, N18570);
not NOT1 (N21254, N21252);
and AND2 (N21255, N21253, N5484);
nand NAND4 (N21256, N21244, N15796, N153, N15553);
nor NOR2 (N21257, N21254, N14016);
buf BUF1 (N21258, N21257);
xor XOR2 (N21259, N21251, N12326);
nand NAND2 (N21260, N21256, N3074);
and AND2 (N21261, N21238, N2783);
and AND2 (N21262, N21255, N17426);
and AND3 (N21263, N21261, N17765, N16513);
and AND2 (N21264, N21263, N10164);
buf BUF1 (N21265, N21204);
nor NOR3 (N21266, N21243, N8277, N20425);
nand NAND2 (N21267, N21259, N3490);
not NOT1 (N21268, N21247);
and AND2 (N21269, N21264, N10470);
xor XOR2 (N21270, N21265, N13090);
or OR2 (N21271, N21269, N3543);
nand NAND2 (N21272, N21271, N17634);
buf BUF1 (N21273, N21266);
xor XOR2 (N21274, N21267, N21113);
or OR4 (N21275, N21273, N14081, N19451, N17284);
buf BUF1 (N21276, N21270);
or OR2 (N21277, N21274, N4999);
not NOT1 (N21278, N21277);
nor NOR3 (N21279, N21260, N6009, N14402);
and AND3 (N21280, N21272, N19386, N1520);
nor NOR2 (N21281, N21278, N219);
buf BUF1 (N21282, N21262);
or OR3 (N21283, N21268, N7525, N16986);
xor XOR2 (N21284, N21283, N1317);
buf BUF1 (N21285, N21275);
nor NOR2 (N21286, N21285, N19110);
xor XOR2 (N21287, N21258, N10443);
or OR3 (N21288, N21284, N9604, N20530);
nand NAND4 (N21289, N21250, N14844, N2956, N8403);
buf BUF1 (N21290, N21282);
or OR2 (N21291, N21289, N11083);
nor NOR2 (N21292, N21281, N7626);
not NOT1 (N21293, N21280);
xor XOR2 (N21294, N21293, N17986);
not NOT1 (N21295, N21292);
or OR3 (N21296, N21287, N7567, N1946);
nand NAND4 (N21297, N21294, N12712, N3839, N15747);
nand NAND4 (N21298, N21286, N192, N7930, N10865);
nand NAND3 (N21299, N21290, N3199, N12172);
or OR3 (N21300, N21291, N8895, N18377);
nand NAND3 (N21301, N21276, N1810, N9685);
buf BUF1 (N21302, N21248);
buf BUF1 (N21303, N21298);
nand NAND3 (N21304, N21302, N2722, N21289);
xor XOR2 (N21305, N21299, N19058);
and AND3 (N21306, N21295, N12852, N10060);
not NOT1 (N21307, N21300);
and AND4 (N21308, N21306, N11425, N8504, N11780);
or OR4 (N21309, N21288, N14874, N14037, N15780);
nor NOR4 (N21310, N21307, N16237, N16387, N4983);
xor XOR2 (N21311, N21309, N2362);
or OR4 (N21312, N21279, N3706, N14097, N15942);
nor NOR3 (N21313, N21311, N651, N3282);
not NOT1 (N21314, N21303);
nor NOR4 (N21315, N21305, N145, N6523, N14847);
not NOT1 (N21316, N21297);
nor NOR3 (N21317, N21310, N8291, N5696);
buf BUF1 (N21318, N21315);
nand NAND2 (N21319, N21313, N7178);
and AND4 (N21320, N21312, N6527, N5821, N18879);
nor NOR3 (N21321, N21314, N11118, N10044);
or OR3 (N21322, N21317, N15946, N7173);
not NOT1 (N21323, N21296);
nand NAND3 (N21324, N21316, N306, N10937);
xor XOR2 (N21325, N21304, N16912);
xor XOR2 (N21326, N21318, N8530);
or OR4 (N21327, N21324, N744, N4311, N5046);
nor NOR4 (N21328, N21319, N12636, N11411, N16464);
and AND4 (N21329, N21320, N2444, N9952, N20912);
xor XOR2 (N21330, N21328, N18976);
nand NAND3 (N21331, N21301, N13718, N15068);
nand NAND3 (N21332, N21329, N7017, N6783);
nand NAND3 (N21333, N21331, N17794, N18824);
buf BUF1 (N21334, N21327);
buf BUF1 (N21335, N21308);
xor XOR2 (N21336, N21321, N21319);
xor XOR2 (N21337, N21333, N16987);
or OR3 (N21338, N21334, N13747, N7105);
and AND2 (N21339, N21330, N3501);
nand NAND3 (N21340, N21335, N12411, N12485);
not NOT1 (N21341, N21337);
nand NAND3 (N21342, N21332, N7531, N16002);
nor NOR4 (N21343, N21342, N5556, N20891, N17497);
xor XOR2 (N21344, N21343, N14818);
buf BUF1 (N21345, N21323);
and AND2 (N21346, N21345, N3862);
xor XOR2 (N21347, N21341, N4964);
not NOT1 (N21348, N21346);
xor XOR2 (N21349, N21325, N14739);
or OR4 (N21350, N21322, N922, N4728, N9933);
nand NAND4 (N21351, N21347, N14967, N8022, N7893);
nand NAND3 (N21352, N21326, N1173, N9649);
nor NOR4 (N21353, N21348, N19036, N15675, N15621);
or OR3 (N21354, N21338, N17180, N2986);
xor XOR2 (N21355, N21352, N19050);
not NOT1 (N21356, N21339);
or OR4 (N21357, N21349, N857, N3471, N16861);
not NOT1 (N21358, N21357);
and AND4 (N21359, N21350, N8300, N14575, N17970);
not NOT1 (N21360, N21340);
and AND2 (N21361, N21353, N15421);
or OR3 (N21362, N21355, N10140, N2282);
and AND4 (N21363, N21361, N20242, N8696, N5515);
nor NOR4 (N21364, N21356, N10333, N7148, N4491);
not NOT1 (N21365, N21360);
and AND2 (N21366, N21354, N12865);
nand NAND2 (N21367, N21362, N11640);
or OR4 (N21368, N21366, N20261, N10626, N17660);
xor XOR2 (N21369, N21365, N14721);
nor NOR2 (N21370, N21358, N4416);
or OR2 (N21371, N21367, N1601);
or OR3 (N21372, N21336, N1477, N8450);
not NOT1 (N21373, N21351);
nor NOR2 (N21374, N21369, N4764);
not NOT1 (N21375, N21374);
nor NOR3 (N21376, N21370, N13771, N14677);
xor XOR2 (N21377, N21363, N13208);
nor NOR4 (N21378, N21368, N5682, N20469, N7160);
nand NAND4 (N21379, N21364, N17907, N12957, N3233);
and AND2 (N21380, N21344, N1860);
nand NAND4 (N21381, N21359, N14306, N5297, N9412);
buf BUF1 (N21382, N21380);
not NOT1 (N21383, N21381);
or OR4 (N21384, N21377, N5226, N8404, N17220);
buf BUF1 (N21385, N21378);
not NOT1 (N21386, N21379);
not NOT1 (N21387, N21373);
or OR2 (N21388, N21376, N9847);
not NOT1 (N21389, N21384);
buf BUF1 (N21390, N21382);
buf BUF1 (N21391, N21387);
buf BUF1 (N21392, N21389);
buf BUF1 (N21393, N21375);
xor XOR2 (N21394, N21386, N15596);
not NOT1 (N21395, N21388);
not NOT1 (N21396, N21372);
nand NAND4 (N21397, N21393, N9892, N9250, N19110);
or OR2 (N21398, N21395, N2163);
not NOT1 (N21399, N21383);
buf BUF1 (N21400, N21394);
not NOT1 (N21401, N21400);
nand NAND4 (N21402, N21401, N11662, N13448, N8083);
or OR4 (N21403, N21385, N19321, N13863, N12223);
nor NOR3 (N21404, N21396, N10292, N7834);
and AND2 (N21405, N21391, N8961);
nor NOR3 (N21406, N21390, N8494, N9651);
not NOT1 (N21407, N21397);
xor XOR2 (N21408, N21402, N3579);
not NOT1 (N21409, N21371);
xor XOR2 (N21410, N21406, N9051);
nor NOR4 (N21411, N21398, N11579, N2025, N7605);
nor NOR4 (N21412, N21392, N17004, N18399, N12664);
and AND3 (N21413, N21408, N19653, N20681);
buf BUF1 (N21414, N21410);
xor XOR2 (N21415, N21403, N1671);
not NOT1 (N21416, N21407);
nor NOR4 (N21417, N21414, N15311, N317, N3373);
buf BUF1 (N21418, N21415);
nor NOR3 (N21419, N21413, N13740, N16803);
xor XOR2 (N21420, N21405, N1169);
or OR4 (N21421, N21404, N19439, N7158, N12854);
or OR3 (N21422, N21411, N19870, N18601);
not NOT1 (N21423, N21421);
nor NOR3 (N21424, N21423, N21277, N10249);
and AND4 (N21425, N21409, N4325, N113, N4733);
nand NAND2 (N21426, N21419, N12316);
nand NAND3 (N21427, N21424, N16384, N19272);
not NOT1 (N21428, N21417);
or OR3 (N21429, N21428, N17537, N6497);
and AND4 (N21430, N21425, N1673, N2214, N18696);
nand NAND2 (N21431, N21426, N6693);
xor XOR2 (N21432, N21416, N2748);
nand NAND4 (N21433, N21422, N19415, N20751, N8194);
nor NOR4 (N21434, N21418, N6506, N13980, N6826);
nor NOR3 (N21435, N21420, N5417, N11686);
xor XOR2 (N21436, N21433, N2940);
nand NAND3 (N21437, N21429, N14681, N16073);
nor NOR4 (N21438, N21399, N14114, N6970, N9716);
not NOT1 (N21439, N21435);
xor XOR2 (N21440, N21412, N1214);
nand NAND3 (N21441, N21430, N3006, N18802);
nand NAND3 (N21442, N21440, N9394, N8186);
or OR3 (N21443, N21436, N7996, N15883);
nand NAND3 (N21444, N21441, N15659, N12638);
nand NAND2 (N21445, N21427, N1310);
nand NAND4 (N21446, N21431, N3821, N13291, N2505);
buf BUF1 (N21447, N21432);
nand NAND4 (N21448, N21446, N17772, N15965, N9672);
not NOT1 (N21449, N21445);
or OR4 (N21450, N21437, N11782, N194, N8738);
and AND3 (N21451, N21447, N6343, N7650);
and AND2 (N21452, N21448, N9897);
nand NAND4 (N21453, N21434, N11554, N6175, N12846);
nor NOR2 (N21454, N21439, N11541);
buf BUF1 (N21455, N21451);
not NOT1 (N21456, N21442);
nor NOR3 (N21457, N21449, N3167, N1766);
buf BUF1 (N21458, N21438);
buf BUF1 (N21459, N21452);
or OR4 (N21460, N21455, N1957, N74, N6635);
not NOT1 (N21461, N21454);
nand NAND4 (N21462, N21458, N9148, N7983, N1847);
nor NOR3 (N21463, N21459, N19059, N8775);
nand NAND2 (N21464, N21462, N16740);
not NOT1 (N21465, N21443);
and AND3 (N21466, N21453, N18924, N7319);
xor XOR2 (N21467, N21460, N17906);
nor NOR4 (N21468, N21457, N21382, N1063, N16598);
nor NOR4 (N21469, N21450, N5989, N4185, N11660);
and AND4 (N21470, N21464, N16125, N2536, N10827);
not NOT1 (N21471, N21466);
nand NAND3 (N21472, N21465, N5435, N13994);
and AND4 (N21473, N21468, N19497, N2450, N11431);
not NOT1 (N21474, N21473);
xor XOR2 (N21475, N21463, N19607);
nor NOR4 (N21476, N21470, N19407, N10972, N1616);
nor NOR4 (N21477, N21456, N3870, N1529, N7113);
xor XOR2 (N21478, N21472, N12542);
buf BUF1 (N21479, N21474);
and AND2 (N21480, N21467, N3337);
not NOT1 (N21481, N21471);
and AND2 (N21482, N21479, N13132);
buf BUF1 (N21483, N21478);
nand NAND4 (N21484, N21481, N10913, N17551, N17772);
and AND3 (N21485, N21482, N2425, N4388);
xor XOR2 (N21486, N21469, N3779);
not NOT1 (N21487, N21444);
not NOT1 (N21488, N21461);
buf BUF1 (N21489, N21484);
not NOT1 (N21490, N21485);
and AND2 (N21491, N21488, N19179);
nor NOR2 (N21492, N21475, N13115);
or OR2 (N21493, N21480, N18948);
and AND2 (N21494, N21492, N3134);
xor XOR2 (N21495, N21483, N8712);
nand NAND2 (N21496, N21486, N21316);
or OR3 (N21497, N21493, N9747, N11812);
or OR4 (N21498, N21496, N1539, N4653, N102);
and AND2 (N21499, N21491, N2560);
or OR2 (N21500, N21494, N19946);
buf BUF1 (N21501, N21498);
not NOT1 (N21502, N21487);
buf BUF1 (N21503, N21500);
and AND4 (N21504, N21503, N13369, N5879, N3073);
nand NAND2 (N21505, N21477, N15058);
buf BUF1 (N21506, N21497);
nand NAND2 (N21507, N21476, N4772);
nand NAND3 (N21508, N21507, N9386, N10742);
nand NAND4 (N21509, N21489, N18106, N7295, N19980);
xor XOR2 (N21510, N21506, N19659);
buf BUF1 (N21511, N21504);
xor XOR2 (N21512, N21511, N42);
nor NOR3 (N21513, N21512, N3872, N5567);
or OR4 (N21514, N21509, N3873, N13172, N18446);
nand NAND3 (N21515, N21505, N19331, N20733);
or OR3 (N21516, N21510, N11709, N19905);
buf BUF1 (N21517, N21501);
not NOT1 (N21518, N21502);
buf BUF1 (N21519, N21508);
nand NAND3 (N21520, N21490, N6590, N9125);
nor NOR3 (N21521, N21513, N9951, N13212);
not NOT1 (N21522, N21520);
xor XOR2 (N21523, N21495, N874);
xor XOR2 (N21524, N21522, N281);
buf BUF1 (N21525, N21524);
and AND4 (N21526, N21516, N11452, N5591, N6276);
xor XOR2 (N21527, N21517, N16352);
nor NOR4 (N21528, N21514, N2722, N9281, N1502);
nand NAND4 (N21529, N21527, N1126, N17775, N12436);
or OR4 (N21530, N21519, N18237, N10893, N2719);
not NOT1 (N21531, N21526);
and AND3 (N21532, N21528, N147, N3926);
xor XOR2 (N21533, N21499, N13321);
buf BUF1 (N21534, N21533);
nor NOR2 (N21535, N21532, N19002);
buf BUF1 (N21536, N21525);
nor NOR4 (N21537, N21521, N11629, N5866, N13228);
and AND2 (N21538, N21523, N10239);
or OR2 (N21539, N21530, N3380);
xor XOR2 (N21540, N21539, N3931);
buf BUF1 (N21541, N21515);
xor XOR2 (N21542, N21540, N10652);
not NOT1 (N21543, N21529);
buf BUF1 (N21544, N21543);
not NOT1 (N21545, N21531);
and AND3 (N21546, N21535, N18537, N16989);
and AND4 (N21547, N21537, N20531, N19586, N20228);
and AND2 (N21548, N21518, N6583);
buf BUF1 (N21549, N21548);
not NOT1 (N21550, N21541);
nand NAND3 (N21551, N21550, N15631, N11043);
buf BUF1 (N21552, N21544);
and AND2 (N21553, N21551, N20040);
xor XOR2 (N21554, N21538, N365);
nor NOR4 (N21555, N21552, N2916, N7556, N15226);
nand NAND4 (N21556, N21534, N1252, N2310, N8879);
nor NOR2 (N21557, N21542, N7845);
not NOT1 (N21558, N21546);
or OR3 (N21559, N21545, N19913, N20017);
or OR3 (N21560, N21557, N15868, N14847);
nand NAND4 (N21561, N21559, N10756, N16742, N16896);
not NOT1 (N21562, N21555);
and AND2 (N21563, N21536, N16426);
xor XOR2 (N21564, N21562, N4798);
nor NOR4 (N21565, N21549, N9869, N19816, N12406);
nor NOR3 (N21566, N21564, N1055, N7742);
nor NOR3 (N21567, N21553, N20423, N14392);
buf BUF1 (N21568, N21554);
not NOT1 (N21569, N21561);
nor NOR3 (N21570, N21560, N16324, N17147);
xor XOR2 (N21571, N21570, N4354);
nand NAND4 (N21572, N21558, N13313, N13052, N10277);
buf BUF1 (N21573, N21563);
or OR4 (N21574, N21547, N18008, N9125, N14454);
nand NAND2 (N21575, N21565, N3458);
xor XOR2 (N21576, N21566, N11481);
and AND4 (N21577, N21556, N7415, N963, N13494);
buf BUF1 (N21578, N21576);
nand NAND3 (N21579, N21574, N746, N13106);
buf BUF1 (N21580, N21579);
buf BUF1 (N21581, N21568);
not NOT1 (N21582, N21567);
or OR2 (N21583, N21575, N11333);
and AND4 (N21584, N21572, N2867, N11004, N11326);
not NOT1 (N21585, N21584);
xor XOR2 (N21586, N21571, N9856);
buf BUF1 (N21587, N21580);
and AND2 (N21588, N21569, N6518);
not NOT1 (N21589, N21585);
not NOT1 (N21590, N21578);
buf BUF1 (N21591, N21589);
xor XOR2 (N21592, N21581, N482);
nor NOR2 (N21593, N21577, N1988);
buf BUF1 (N21594, N21573);
or OR2 (N21595, N21588, N18488);
or OR2 (N21596, N21590, N20679);
xor XOR2 (N21597, N21591, N5343);
and AND3 (N21598, N21596, N17268, N16516);
nor NOR2 (N21599, N21586, N5263);
not NOT1 (N21600, N21595);
not NOT1 (N21601, N21600);
nand NAND2 (N21602, N21592, N14366);
not NOT1 (N21603, N21598);
and AND2 (N21604, N21587, N2488);
not NOT1 (N21605, N21583);
or OR3 (N21606, N21594, N9735, N2501);
nand NAND3 (N21607, N21605, N20777, N11533);
nand NAND4 (N21608, N21607, N18839, N8431, N7929);
nor NOR3 (N21609, N21603, N7300, N19236);
nand NAND2 (N21610, N21604, N356);
not NOT1 (N21611, N21602);
xor XOR2 (N21612, N21582, N6836);
nand NAND4 (N21613, N21608, N4122, N11989, N6532);
not NOT1 (N21614, N21613);
and AND3 (N21615, N21612, N16517, N14964);
xor XOR2 (N21616, N21609, N12400);
xor XOR2 (N21617, N21610, N12115);
and AND2 (N21618, N21616, N6827);
or OR3 (N21619, N21601, N19124, N12067);
and AND3 (N21620, N21611, N17280, N7378);
nor NOR4 (N21621, N21597, N2289, N10352, N8837);
and AND2 (N21622, N21615, N4073);
and AND4 (N21623, N21614, N21608, N2346, N17638);
xor XOR2 (N21624, N21622, N7007);
buf BUF1 (N21625, N21606);
nand NAND4 (N21626, N21593, N15860, N18276, N21579);
xor XOR2 (N21627, N21599, N13622);
or OR2 (N21628, N21625, N17500);
not NOT1 (N21629, N21627);
nand NAND3 (N21630, N21620, N20960, N20898);
buf BUF1 (N21631, N21618);
xor XOR2 (N21632, N21630, N11427);
nor NOR2 (N21633, N21619, N8515);
and AND3 (N21634, N21626, N10530, N18824);
nor NOR2 (N21635, N21632, N11386);
or OR3 (N21636, N21623, N19929, N58);
nor NOR4 (N21637, N21633, N11982, N11981, N8618);
and AND2 (N21638, N21621, N17857);
nand NAND2 (N21639, N21628, N4768);
nand NAND2 (N21640, N21637, N18601);
and AND3 (N21641, N21624, N19215, N10430);
or OR3 (N21642, N21636, N3695, N5651);
and AND3 (N21643, N21629, N19290, N20192);
not NOT1 (N21644, N21641);
not NOT1 (N21645, N21640);
and AND3 (N21646, N21638, N8511, N18763);
nor NOR3 (N21647, N21634, N18191, N19986);
or OR3 (N21648, N21644, N13831, N16176);
not NOT1 (N21649, N21645);
nor NOR2 (N21650, N21643, N5006);
not NOT1 (N21651, N21617);
buf BUF1 (N21652, N21642);
not NOT1 (N21653, N21652);
or OR3 (N21654, N21646, N19687, N8035);
not NOT1 (N21655, N21648);
not NOT1 (N21656, N21635);
xor XOR2 (N21657, N21649, N6988);
or OR2 (N21658, N21654, N12662);
nor NOR3 (N21659, N21651, N13192, N12233);
buf BUF1 (N21660, N21658);
not NOT1 (N21661, N21660);
nand NAND2 (N21662, N21659, N2902);
buf BUF1 (N21663, N21662);
or OR2 (N21664, N21655, N7247);
buf BUF1 (N21665, N21653);
nor NOR4 (N21666, N21661, N1310, N2735, N19018);
and AND2 (N21667, N21666, N20372);
nor NOR4 (N21668, N21631, N4023, N71, N21609);
buf BUF1 (N21669, N21639);
buf BUF1 (N21670, N21665);
or OR3 (N21671, N21650, N991, N3696);
and AND4 (N21672, N21668, N8003, N230, N16972);
xor XOR2 (N21673, N21647, N14745);
and AND4 (N21674, N21656, N7192, N19437, N8349);
nand NAND3 (N21675, N21663, N9145, N1541);
buf BUF1 (N21676, N21669);
buf BUF1 (N21677, N21675);
xor XOR2 (N21678, N21657, N15715);
nor NOR4 (N21679, N21674, N5939, N10960, N18433);
buf BUF1 (N21680, N21672);
buf BUF1 (N21681, N21676);
and AND2 (N21682, N21671, N20780);
nor NOR4 (N21683, N21680, N15315, N12307, N4131);
nand NAND2 (N21684, N21673, N19986);
buf BUF1 (N21685, N21683);
not NOT1 (N21686, N21677);
nand NAND2 (N21687, N21682, N8175);
xor XOR2 (N21688, N21681, N15274);
or OR3 (N21689, N21667, N3322, N6838);
and AND2 (N21690, N21664, N2082);
nor NOR3 (N21691, N21684, N17556, N15345);
buf BUF1 (N21692, N21688);
nor NOR2 (N21693, N21687, N16878);
nand NAND3 (N21694, N21693, N4640, N4869);
buf BUF1 (N21695, N21689);
buf BUF1 (N21696, N21692);
not NOT1 (N21697, N21670);
buf BUF1 (N21698, N21685);
nand NAND4 (N21699, N21697, N17677, N6715, N21654);
xor XOR2 (N21700, N21698, N5607);
buf BUF1 (N21701, N21699);
nor NOR4 (N21702, N21690, N8570, N4964, N20151);
nor NOR3 (N21703, N21686, N3504, N17770);
buf BUF1 (N21704, N21678);
buf BUF1 (N21705, N21702);
and AND3 (N21706, N21701, N2019, N1949);
or OR3 (N21707, N21696, N16460, N17821);
buf BUF1 (N21708, N21700);
nand NAND4 (N21709, N21679, N1504, N5983, N1546);
nand NAND4 (N21710, N21695, N14999, N11876, N13703);
buf BUF1 (N21711, N21691);
and AND3 (N21712, N21711, N20335, N7333);
xor XOR2 (N21713, N21710, N880);
or OR3 (N21714, N21703, N6613, N19161);
and AND3 (N21715, N21704, N19529, N13784);
and AND2 (N21716, N21706, N6810);
buf BUF1 (N21717, N21714);
and AND4 (N21718, N21694, N10695, N21131, N13153);
or OR2 (N21719, N21717, N21377);
not NOT1 (N21720, N21716);
xor XOR2 (N21721, N21720, N19528);
nand NAND2 (N21722, N21705, N3667);
not NOT1 (N21723, N21708);
not NOT1 (N21724, N21709);
and AND3 (N21725, N21718, N11688, N126);
or OR2 (N21726, N21719, N7330);
and AND3 (N21727, N21721, N3751, N6204);
and AND4 (N21728, N21726, N16659, N12850, N12950);
buf BUF1 (N21729, N21712);
nand NAND2 (N21730, N21707, N18919);
nand NAND3 (N21731, N21722, N17972, N18136);
or OR3 (N21732, N21731, N993, N2851);
nor NOR4 (N21733, N21713, N2682, N2983, N2462);
not NOT1 (N21734, N21730);
or OR3 (N21735, N21734, N3723, N4140);
nor NOR2 (N21736, N21723, N8093);
and AND2 (N21737, N21735, N4541);
nor NOR2 (N21738, N21727, N19773);
nand NAND2 (N21739, N21732, N11494);
nand NAND3 (N21740, N21724, N17383, N19500);
buf BUF1 (N21741, N21737);
buf BUF1 (N21742, N21728);
xor XOR2 (N21743, N21741, N5311);
or OR3 (N21744, N21725, N5550, N11685);
nand NAND3 (N21745, N21742, N5042, N12450);
buf BUF1 (N21746, N21745);
nor NOR4 (N21747, N21733, N16991, N18508, N494);
or OR3 (N21748, N21739, N21223, N11430);
nand NAND4 (N21749, N21715, N15985, N4777, N9364);
and AND2 (N21750, N21738, N15559);
or OR2 (N21751, N21736, N15737);
nand NAND2 (N21752, N21729, N10134);
nand NAND2 (N21753, N21744, N3551);
buf BUF1 (N21754, N21748);
nand NAND3 (N21755, N21750, N11017, N15737);
and AND2 (N21756, N21751, N7953);
buf BUF1 (N21757, N21740);
and AND4 (N21758, N21754, N15899, N16325, N16787);
not NOT1 (N21759, N21749);
nor NOR3 (N21760, N21752, N9409, N19594);
and AND2 (N21761, N21743, N655);
and AND4 (N21762, N21760, N2622, N3019, N5456);
and AND3 (N21763, N21761, N15757, N10667);
not NOT1 (N21764, N21762);
and AND4 (N21765, N21764, N15918, N19348, N14129);
nand NAND3 (N21766, N21746, N9156, N6711);
xor XOR2 (N21767, N21759, N9448);
buf BUF1 (N21768, N21765);
buf BUF1 (N21769, N21767);
or OR2 (N21770, N21766, N17087);
not NOT1 (N21771, N21768);
not NOT1 (N21772, N21756);
buf BUF1 (N21773, N21770);
xor XOR2 (N21774, N21755, N10495);
nor NOR3 (N21775, N21747, N5008, N8232);
nand NAND2 (N21776, N21758, N19565);
xor XOR2 (N21777, N21773, N2513);
not NOT1 (N21778, N21775);
nand NAND2 (N21779, N21778, N8864);
or OR3 (N21780, N21774, N9868, N12053);
or OR2 (N21781, N21771, N1355);
buf BUF1 (N21782, N21779);
and AND2 (N21783, N21757, N2264);
xor XOR2 (N21784, N21753, N9290);
buf BUF1 (N21785, N21763);
and AND2 (N21786, N21769, N719);
nor NOR2 (N21787, N21782, N18354);
or OR4 (N21788, N21781, N2491, N659, N18307);
buf BUF1 (N21789, N21784);
xor XOR2 (N21790, N21785, N5491);
nand NAND4 (N21791, N21786, N7702, N9072, N14961);
nor NOR3 (N21792, N21780, N20210, N13103);
xor XOR2 (N21793, N21777, N7715);
nand NAND3 (N21794, N21790, N16800, N397);
xor XOR2 (N21795, N21783, N20862);
xor XOR2 (N21796, N21788, N18766);
not NOT1 (N21797, N21789);
and AND3 (N21798, N21787, N3707, N10829);
buf BUF1 (N21799, N21797);
xor XOR2 (N21800, N21796, N17148);
nor NOR3 (N21801, N21791, N21451, N14626);
nand NAND4 (N21802, N21776, N18958, N16954, N7899);
buf BUF1 (N21803, N21793);
nand NAND3 (N21804, N21802, N14055, N21654);
buf BUF1 (N21805, N21772);
and AND2 (N21806, N21803, N14572);
buf BUF1 (N21807, N21801);
or OR2 (N21808, N21807, N12060);
nand NAND4 (N21809, N21795, N6206, N4015, N15453);
xor XOR2 (N21810, N21800, N7005);
nand NAND4 (N21811, N21806, N18386, N15567, N7870);
nand NAND4 (N21812, N21792, N12147, N9035, N5450);
not NOT1 (N21813, N21804);
or OR3 (N21814, N21808, N19056, N7685);
not NOT1 (N21815, N21810);
buf BUF1 (N21816, N21799);
buf BUF1 (N21817, N21812);
and AND3 (N21818, N21813, N19401, N4419);
not NOT1 (N21819, N21815);
and AND2 (N21820, N21818, N2990);
nand NAND2 (N21821, N21811, N18484);
not NOT1 (N21822, N21819);
xor XOR2 (N21823, N21820, N2921);
or OR4 (N21824, N21814, N1659, N10116, N8225);
nor NOR4 (N21825, N21798, N10661, N9097, N4645);
nand NAND3 (N21826, N21816, N12381, N11513);
xor XOR2 (N21827, N21817, N18165);
xor XOR2 (N21828, N21822, N7536);
not NOT1 (N21829, N21828);
buf BUF1 (N21830, N21794);
and AND3 (N21831, N21823, N7585, N14058);
nand NAND3 (N21832, N21829, N16889, N18293);
and AND3 (N21833, N21831, N5886, N125);
nor NOR3 (N21834, N21833, N13532, N7231);
or OR3 (N21835, N21830, N9402, N8663);
and AND4 (N21836, N21827, N1456, N17607, N14002);
nand NAND4 (N21837, N21824, N11048, N14744, N2863);
not NOT1 (N21838, N21826);
or OR4 (N21839, N21821, N13855, N9653, N7250);
nor NOR2 (N21840, N21809, N11076);
and AND3 (N21841, N21838, N3207, N14396);
nor NOR3 (N21842, N21840, N17349, N13768);
nand NAND2 (N21843, N21825, N19061);
not NOT1 (N21844, N21805);
nand NAND3 (N21845, N21843, N1467, N5203);
buf BUF1 (N21846, N21835);
nor NOR4 (N21847, N21836, N4479, N6569, N8894);
or OR3 (N21848, N21844, N5203, N7651);
and AND3 (N21849, N21834, N15276, N15517);
not NOT1 (N21850, N21847);
xor XOR2 (N21851, N21839, N12936);
buf BUF1 (N21852, N21846);
buf BUF1 (N21853, N21841);
and AND4 (N21854, N21853, N5479, N12186, N16434);
xor XOR2 (N21855, N21842, N6416);
or OR3 (N21856, N21851, N8521, N8138);
and AND3 (N21857, N21855, N4907, N19179);
or OR3 (N21858, N21856, N6707, N13005);
xor XOR2 (N21859, N21854, N6411);
nand NAND4 (N21860, N21845, N2180, N11894, N1939);
nor NOR4 (N21861, N21857, N16911, N4653, N11691);
nor NOR2 (N21862, N21852, N20192);
nor NOR3 (N21863, N21849, N6855, N17491);
and AND3 (N21864, N21832, N21400, N15243);
nand NAND3 (N21865, N21859, N2007, N11297);
not NOT1 (N21866, N21864);
not NOT1 (N21867, N21837);
and AND3 (N21868, N21858, N12248, N18189);
xor XOR2 (N21869, N21861, N7335);
xor XOR2 (N21870, N21866, N10279);
not NOT1 (N21871, N21863);
nor NOR4 (N21872, N21850, N19616, N9604, N15737);
not NOT1 (N21873, N21860);
nand NAND3 (N21874, N21868, N135, N8194);
xor XOR2 (N21875, N21871, N12527);
nand NAND3 (N21876, N21865, N227, N5997);
not NOT1 (N21877, N21848);
or OR2 (N21878, N21873, N13739);
or OR4 (N21879, N21862, N20582, N106, N13258);
xor XOR2 (N21880, N21876, N7182);
xor XOR2 (N21881, N21878, N15253);
buf BUF1 (N21882, N21874);
buf BUF1 (N21883, N21875);
and AND3 (N21884, N21870, N1433, N7915);
xor XOR2 (N21885, N21867, N3747);
xor XOR2 (N21886, N21872, N13875);
buf BUF1 (N21887, N21886);
nor NOR3 (N21888, N21877, N10006, N8157);
xor XOR2 (N21889, N21881, N8326);
nand NAND3 (N21890, N21880, N15409, N9126);
nor NOR4 (N21891, N21869, N9854, N16601, N5904);
xor XOR2 (N21892, N21885, N21372);
buf BUF1 (N21893, N21891);
or OR2 (N21894, N21893, N12450);
nor NOR4 (N21895, N21889, N19399, N20139, N2910);
and AND3 (N21896, N21895, N5767, N17296);
buf BUF1 (N21897, N21879);
nand NAND4 (N21898, N21883, N9205, N19286, N9823);
and AND4 (N21899, N21898, N7290, N11457, N2707);
xor XOR2 (N21900, N21890, N8854);
not NOT1 (N21901, N21888);
nand NAND4 (N21902, N21894, N5079, N21406, N10955);
not NOT1 (N21903, N21882);
xor XOR2 (N21904, N21897, N801);
or OR4 (N21905, N21903, N6984, N23, N17322);
buf BUF1 (N21906, N21896);
or OR3 (N21907, N21887, N5497, N12755);
not NOT1 (N21908, N21884);
not NOT1 (N21909, N21906);
buf BUF1 (N21910, N21909);
nor NOR2 (N21911, N21892, N19685);
not NOT1 (N21912, N21901);
not NOT1 (N21913, N21900);
not NOT1 (N21914, N21913);
xor XOR2 (N21915, N21912, N15021);
and AND2 (N21916, N21902, N20959);
or OR3 (N21917, N21915, N9729, N4538);
and AND3 (N21918, N21904, N8423, N7750);
xor XOR2 (N21919, N21908, N95);
buf BUF1 (N21920, N21917);
not NOT1 (N21921, N21911);
and AND3 (N21922, N21910, N8082, N13766);
or OR4 (N21923, N21921, N6393, N2617, N19075);
or OR3 (N21924, N21914, N6949, N15362);
not NOT1 (N21925, N21919);
not NOT1 (N21926, N21907);
not NOT1 (N21927, N21925);
xor XOR2 (N21928, N21918, N21663);
xor XOR2 (N21929, N21916, N6295);
xor XOR2 (N21930, N21928, N9578);
buf BUF1 (N21931, N21920);
buf BUF1 (N21932, N21905);
xor XOR2 (N21933, N21932, N16365);
nand NAND4 (N21934, N21930, N21168, N3176, N4929);
nand NAND2 (N21935, N21929, N13288);
nor NOR3 (N21936, N21931, N16479, N7831);
nand NAND4 (N21937, N21924, N14373, N7308, N12);
nor NOR3 (N21938, N21933, N6636, N6310);
or OR3 (N21939, N21935, N14208, N789);
nor NOR3 (N21940, N21926, N18979, N5414);
and AND2 (N21941, N21922, N6068);
or OR4 (N21942, N21899, N13102, N17887, N18784);
nor NOR4 (N21943, N21941, N12255, N21005, N5402);
not NOT1 (N21944, N21943);
or OR2 (N21945, N21934, N18811);
buf BUF1 (N21946, N21939);
buf BUF1 (N21947, N21936);
xor XOR2 (N21948, N21938, N16971);
not NOT1 (N21949, N21923);
or OR2 (N21950, N21940, N7438);
not NOT1 (N21951, N21944);
or OR4 (N21952, N21927, N16183, N12768, N2129);
buf BUF1 (N21953, N21942);
nor NOR4 (N21954, N21946, N665, N20884, N18644);
nor NOR4 (N21955, N21954, N8643, N3677, N4892);
xor XOR2 (N21956, N21952, N15842);
nand NAND2 (N21957, N21955, N2009);
and AND3 (N21958, N21947, N10633, N6951);
or OR2 (N21959, N21957, N17445);
nor NOR4 (N21960, N21948, N8730, N14390, N15645);
and AND4 (N21961, N21956, N3164, N3889, N6698);
nor NOR2 (N21962, N21951, N6523);
and AND4 (N21963, N21953, N13012, N28, N21763);
or OR4 (N21964, N21937, N18067, N14411, N7910);
nand NAND2 (N21965, N21962, N21572);
or OR2 (N21966, N21965, N8695);
nor NOR4 (N21967, N21963, N20154, N10065, N16861);
buf BUF1 (N21968, N21959);
and AND4 (N21969, N21950, N19643, N11872, N4990);
buf BUF1 (N21970, N21967);
not NOT1 (N21971, N21961);
nor NOR2 (N21972, N21970, N18375);
xor XOR2 (N21973, N21949, N9681);
not NOT1 (N21974, N21960);
nand NAND3 (N21975, N21969, N12560, N9162);
xor XOR2 (N21976, N21945, N16);
nor NOR2 (N21977, N21973, N9958);
buf BUF1 (N21978, N21958);
not NOT1 (N21979, N21966);
or OR4 (N21980, N21964, N20964, N19662, N12417);
buf BUF1 (N21981, N21980);
nor NOR4 (N21982, N21972, N8525, N19737, N18844);
and AND4 (N21983, N21977, N12066, N13796, N18758);
not NOT1 (N21984, N21971);
not NOT1 (N21985, N21968);
and AND4 (N21986, N21974, N8285, N17876, N217);
not NOT1 (N21987, N21976);
or OR2 (N21988, N21983, N7785);
nand NAND4 (N21989, N21982, N19644, N3231, N7081);
nor NOR2 (N21990, N21987, N9829);
and AND4 (N21991, N21981, N17893, N17508, N5735);
and AND4 (N21992, N21989, N21500, N182, N8256);
xor XOR2 (N21993, N21988, N14248);
xor XOR2 (N21994, N21975, N11044);
nor NOR4 (N21995, N21992, N21213, N20309, N18513);
xor XOR2 (N21996, N21994, N3081);
xor XOR2 (N21997, N21984, N723);
or OR2 (N21998, N21991, N13328);
or OR4 (N21999, N21985, N20420, N8951, N1000);
or OR2 (N22000, N21995, N5103);
nor NOR2 (N22001, N21997, N15114);
or OR3 (N22002, N21978, N10255, N6451);
buf BUF1 (N22003, N22001);
buf BUF1 (N22004, N21986);
nor NOR4 (N22005, N21979, N12471, N5381, N10098);
xor XOR2 (N22006, N22005, N19744);
xor XOR2 (N22007, N22003, N18799);
nand NAND2 (N22008, N22004, N20514);
and AND2 (N22009, N22002, N4811);
buf BUF1 (N22010, N21998);
xor XOR2 (N22011, N21990, N19925);
not NOT1 (N22012, N21996);
xor XOR2 (N22013, N22010, N15672);
nor NOR4 (N22014, N22007, N4331, N3041, N9094);
or OR2 (N22015, N22000, N17737);
or OR2 (N22016, N22006, N325);
buf BUF1 (N22017, N22009);
nor NOR2 (N22018, N21993, N13427);
xor XOR2 (N22019, N22016, N12247);
buf BUF1 (N22020, N22017);
xor XOR2 (N22021, N22019, N21402);
xor XOR2 (N22022, N22008, N9433);
not NOT1 (N22023, N22012);
buf BUF1 (N22024, N22018);
not NOT1 (N22025, N22024);
not NOT1 (N22026, N22013);
xor XOR2 (N22027, N22026, N17912);
xor XOR2 (N22028, N22023, N8649);
not NOT1 (N22029, N21999);
not NOT1 (N22030, N22014);
buf BUF1 (N22031, N22029);
buf BUF1 (N22032, N22028);
nand NAND3 (N22033, N22020, N11105, N3686);
buf BUF1 (N22034, N22033);
not NOT1 (N22035, N22022);
nand NAND3 (N22036, N22030, N16275, N21544);
xor XOR2 (N22037, N22031, N11006);
and AND2 (N22038, N22035, N115);
nand NAND2 (N22039, N22034, N628);
buf BUF1 (N22040, N22032);
and AND2 (N22041, N22040, N11171);
nor NOR3 (N22042, N22015, N9239, N21771);
not NOT1 (N22043, N22039);
xor XOR2 (N22044, N22037, N12439);
not NOT1 (N22045, N22044);
nor NOR3 (N22046, N22011, N17456, N7283);
buf BUF1 (N22047, N22027);
not NOT1 (N22048, N22036);
xor XOR2 (N22049, N22038, N18082);
nor NOR4 (N22050, N22047, N17043, N14654, N21613);
not NOT1 (N22051, N22043);
buf BUF1 (N22052, N22045);
not NOT1 (N22053, N22052);
nand NAND3 (N22054, N22053, N11651, N8276);
xor XOR2 (N22055, N22046, N2638);
or OR3 (N22056, N22021, N7259, N1957);
not NOT1 (N22057, N22041);
buf BUF1 (N22058, N22054);
or OR2 (N22059, N22051, N10877);
nor NOR2 (N22060, N22058, N11966);
buf BUF1 (N22061, N22060);
nor NOR2 (N22062, N22042, N11633);
xor XOR2 (N22063, N22055, N16598);
or OR2 (N22064, N22063, N2210);
xor XOR2 (N22065, N22057, N20708);
xor XOR2 (N22066, N22025, N10988);
or OR2 (N22067, N22064, N8337);
buf BUF1 (N22068, N22062);
buf BUF1 (N22069, N22048);
xor XOR2 (N22070, N22068, N2406);
nand NAND4 (N22071, N22050, N17568, N1620, N5462);
xor XOR2 (N22072, N22056, N19995);
and AND4 (N22073, N22066, N1320, N18264, N1109);
and AND4 (N22074, N22073, N5252, N19695, N10069);
or OR2 (N22075, N22071, N19529);
not NOT1 (N22076, N22072);
or OR2 (N22077, N22065, N9470);
nand NAND3 (N22078, N22075, N9401, N9531);
and AND4 (N22079, N22069, N2389, N13699, N13045);
buf BUF1 (N22080, N22078);
xor XOR2 (N22081, N22077, N17008);
not NOT1 (N22082, N22080);
xor XOR2 (N22083, N22076, N8944);
nor NOR2 (N22084, N22083, N5677);
not NOT1 (N22085, N22059);
and AND4 (N22086, N22067, N8461, N19901, N2223);
not NOT1 (N22087, N22070);
not NOT1 (N22088, N22074);
and AND2 (N22089, N22084, N14800);
not NOT1 (N22090, N22049);
and AND3 (N22091, N22061, N17604, N21820);
nor NOR2 (N22092, N22089, N10355);
buf BUF1 (N22093, N22088);
nor NOR4 (N22094, N22085, N22060, N19093, N2389);
xor XOR2 (N22095, N22091, N14866);
nor NOR4 (N22096, N22087, N9976, N4526, N6608);
nor NOR3 (N22097, N22094, N18309, N12636);
xor XOR2 (N22098, N22096, N19873);
buf BUF1 (N22099, N22098);
nand NAND3 (N22100, N22093, N11962, N9282);
nand NAND3 (N22101, N22090, N8041, N7223);
nor NOR3 (N22102, N22079, N11007, N2099);
and AND4 (N22103, N22101, N8033, N19823, N2996);
not NOT1 (N22104, N22081);
buf BUF1 (N22105, N22099);
buf BUF1 (N22106, N22105);
or OR4 (N22107, N22106, N12460, N11306, N5271);
not NOT1 (N22108, N22104);
and AND4 (N22109, N22095, N8349, N6689, N10486);
nor NOR2 (N22110, N22100, N10043);
buf BUF1 (N22111, N22103);
nor NOR2 (N22112, N22111, N10434);
buf BUF1 (N22113, N22086);
or OR4 (N22114, N22102, N5074, N14646, N10127);
not NOT1 (N22115, N22109);
and AND4 (N22116, N22108, N17981, N16884, N10653);
and AND3 (N22117, N22110, N6482, N14524);
xor XOR2 (N22118, N22097, N17031);
xor XOR2 (N22119, N22118, N16957);
buf BUF1 (N22120, N22082);
and AND4 (N22121, N22112, N21674, N7190, N7156);
or OR4 (N22122, N22114, N14360, N19083, N15767);
nor NOR4 (N22123, N22121, N14445, N13614, N5647);
and AND2 (N22124, N22092, N8913);
xor XOR2 (N22125, N22115, N5536);
buf BUF1 (N22126, N22124);
nor NOR4 (N22127, N22107, N16260, N2121, N4279);
nand NAND3 (N22128, N22113, N2242, N13779);
nand NAND2 (N22129, N22125, N1791);
or OR4 (N22130, N22126, N5582, N333, N9634);
and AND2 (N22131, N22123, N346);
xor XOR2 (N22132, N22129, N11834);
and AND3 (N22133, N22127, N3731, N10973);
nor NOR4 (N22134, N22128, N1557, N2357, N2469);
and AND2 (N22135, N22122, N2677);
or OR2 (N22136, N22135, N20410);
nand NAND2 (N22137, N22117, N1830);
or OR2 (N22138, N22119, N8582);
and AND3 (N22139, N22133, N14095, N21662);
nor NOR2 (N22140, N22138, N12828);
and AND2 (N22141, N22131, N15614);
xor XOR2 (N22142, N22120, N18933);
nand NAND4 (N22143, N22132, N4532, N21493, N17026);
buf BUF1 (N22144, N22116);
not NOT1 (N22145, N22136);
xor XOR2 (N22146, N22142, N8492);
nor NOR3 (N22147, N22144, N9306, N4398);
xor XOR2 (N22148, N22143, N20812);
nor NOR4 (N22149, N22145, N14240, N4840, N9334);
xor XOR2 (N22150, N22130, N18516);
nand NAND3 (N22151, N22139, N7243, N6336);
xor XOR2 (N22152, N22147, N18280);
and AND4 (N22153, N22140, N5570, N4331, N5680);
not NOT1 (N22154, N22151);
nand NAND4 (N22155, N22146, N1425, N10465, N7900);
buf BUF1 (N22156, N22150);
xor XOR2 (N22157, N22152, N5706);
not NOT1 (N22158, N22155);
nand NAND4 (N22159, N22134, N9810, N9464, N13479);
buf BUF1 (N22160, N22156);
or OR3 (N22161, N22141, N2730, N9014);
nor NOR2 (N22162, N22158, N6792);
nand NAND4 (N22163, N22149, N22122, N13826, N14291);
and AND4 (N22164, N22163, N54, N3006, N186);
xor XOR2 (N22165, N22164, N16304);
nand NAND2 (N22166, N22162, N3986);
nor NOR4 (N22167, N22137, N17655, N4847, N21480);
nor NOR3 (N22168, N22160, N17453, N9126);
xor XOR2 (N22169, N22165, N10277);
and AND2 (N22170, N22167, N12014);
and AND2 (N22171, N22168, N7999);
and AND4 (N22172, N22157, N19450, N4763, N15863);
not NOT1 (N22173, N22170);
buf BUF1 (N22174, N22161);
not NOT1 (N22175, N22174);
or OR3 (N22176, N22154, N9722, N21957);
nand NAND3 (N22177, N22169, N20381, N12461);
xor XOR2 (N22178, N22153, N4630);
buf BUF1 (N22179, N22171);
xor XOR2 (N22180, N22172, N15126);
not NOT1 (N22181, N22159);
nor NOR2 (N22182, N22166, N19922);
nor NOR3 (N22183, N22180, N5291, N696);
buf BUF1 (N22184, N22177);
nor NOR2 (N22185, N22148, N19748);
or OR3 (N22186, N22178, N18860, N8186);
buf BUF1 (N22187, N22176);
and AND4 (N22188, N22185, N9929, N10708, N7337);
not NOT1 (N22189, N22188);
nor NOR4 (N22190, N22182, N17870, N3426, N11495);
not NOT1 (N22191, N22175);
xor XOR2 (N22192, N22183, N12896);
xor XOR2 (N22193, N22181, N13128);
xor XOR2 (N22194, N22190, N10948);
buf BUF1 (N22195, N22187);
nor NOR3 (N22196, N22195, N12187, N13444);
nor NOR2 (N22197, N22196, N14183);
xor XOR2 (N22198, N22189, N15160);
xor XOR2 (N22199, N22191, N1534);
and AND4 (N22200, N22184, N6052, N3643, N15758);
xor XOR2 (N22201, N22186, N3465);
and AND2 (N22202, N22173, N21369);
xor XOR2 (N22203, N22202, N15246);
and AND2 (N22204, N22193, N13680);
or OR2 (N22205, N22203, N19427);
and AND3 (N22206, N22194, N15882, N20475);
and AND3 (N22207, N22179, N1376, N9709);
nand NAND3 (N22208, N22205, N3555, N9611);
nor NOR3 (N22209, N22206, N20160, N13254);
nand NAND2 (N22210, N22207, N11561);
xor XOR2 (N22211, N22201, N5290);
not NOT1 (N22212, N22210);
and AND4 (N22213, N22198, N1048, N12828, N13709);
or OR2 (N22214, N22204, N18503);
or OR4 (N22215, N22214, N9903, N13268, N5222);
or OR4 (N22216, N22197, N8292, N18685, N9809);
or OR3 (N22217, N22199, N9895, N9402);
buf BUF1 (N22218, N22208);
not NOT1 (N22219, N22200);
and AND4 (N22220, N22211, N9204, N18903, N21149);
not NOT1 (N22221, N22209);
not NOT1 (N22222, N22215);
or OR2 (N22223, N22219, N1736);
nor NOR3 (N22224, N22218, N4229, N14346);
nand NAND4 (N22225, N22212, N14114, N13806, N20289);
or OR4 (N22226, N22224, N10568, N16832, N1508);
nor NOR3 (N22227, N22217, N4933, N5957);
or OR4 (N22228, N22226, N17399, N4941, N1753);
nor NOR4 (N22229, N22228, N19792, N13481, N4523);
nand NAND2 (N22230, N22223, N15104);
buf BUF1 (N22231, N22222);
xor XOR2 (N22232, N22192, N4275);
buf BUF1 (N22233, N22220);
buf BUF1 (N22234, N22213);
nor NOR4 (N22235, N22216, N14005, N19952, N4156);
nand NAND2 (N22236, N22230, N21156);
xor XOR2 (N22237, N22235, N2020);
not NOT1 (N22238, N22229);
nand NAND4 (N22239, N22238, N7524, N8885, N9889);
nor NOR2 (N22240, N22227, N17680);
and AND3 (N22241, N22236, N20622, N17241);
not NOT1 (N22242, N22225);
buf BUF1 (N22243, N22237);
nand NAND2 (N22244, N22240, N8098);
and AND2 (N22245, N22221, N15821);
xor XOR2 (N22246, N22243, N17313);
nor NOR3 (N22247, N22231, N9914, N18779);
or OR4 (N22248, N22239, N10853, N22085, N6013);
buf BUF1 (N22249, N22246);
not NOT1 (N22250, N22242);
nand NAND3 (N22251, N22232, N4301, N10055);
xor XOR2 (N22252, N22251, N14199);
nor NOR3 (N22253, N22248, N16818, N13960);
and AND4 (N22254, N22249, N18249, N10410, N4218);
buf BUF1 (N22255, N22234);
buf BUF1 (N22256, N22252);
and AND3 (N22257, N22244, N17876, N8629);
xor XOR2 (N22258, N22233, N17333);
xor XOR2 (N22259, N22255, N21248);
not NOT1 (N22260, N22245);
or OR4 (N22261, N22256, N22086, N347, N8930);
nand NAND4 (N22262, N22253, N16940, N10273, N8716);
buf BUF1 (N22263, N22247);
nand NAND3 (N22264, N22254, N18849, N22078);
not NOT1 (N22265, N22258);
xor XOR2 (N22266, N22261, N3596);
not NOT1 (N22267, N22262);
xor XOR2 (N22268, N22250, N2781);
not NOT1 (N22269, N22264);
nor NOR4 (N22270, N22263, N12168, N7156, N11515);
nand NAND2 (N22271, N22257, N21888);
buf BUF1 (N22272, N22241);
buf BUF1 (N22273, N22270);
not NOT1 (N22274, N22268);
xor XOR2 (N22275, N22260, N14408);
nand NAND3 (N22276, N22274, N13669, N12646);
buf BUF1 (N22277, N22269);
nand NAND2 (N22278, N22275, N15263);
nor NOR3 (N22279, N22272, N8077, N13242);
not NOT1 (N22280, N22277);
xor XOR2 (N22281, N22280, N15304);
nor NOR3 (N22282, N22271, N22240, N17091);
or OR3 (N22283, N22282, N20024, N15795);
or OR4 (N22284, N22267, N14227, N3572, N12954);
and AND3 (N22285, N22276, N13758, N1982);
or OR4 (N22286, N22281, N21410, N20602, N18496);
xor XOR2 (N22287, N22283, N14406);
buf BUF1 (N22288, N22287);
and AND2 (N22289, N22279, N39);
buf BUF1 (N22290, N22286);
and AND3 (N22291, N22289, N11973, N4552);
nor NOR4 (N22292, N22273, N15750, N21419, N17878);
buf BUF1 (N22293, N22278);
and AND3 (N22294, N22266, N6185, N12264);
or OR3 (N22295, N22285, N9990, N9072);
buf BUF1 (N22296, N22293);
and AND4 (N22297, N22290, N2403, N8024, N19624);
buf BUF1 (N22298, N22296);
buf BUF1 (N22299, N22298);
or OR4 (N22300, N22259, N4399, N12431, N5217);
xor XOR2 (N22301, N22288, N22004);
and AND2 (N22302, N22297, N11746);
nand NAND3 (N22303, N22299, N22278, N18155);
nor NOR4 (N22304, N22291, N14953, N11020, N14161);
not NOT1 (N22305, N22265);
nand NAND3 (N22306, N22303, N7037, N20459);
nor NOR3 (N22307, N22306, N16883, N2079);
xor XOR2 (N22308, N22300, N6997);
xor XOR2 (N22309, N22292, N3670);
nand NAND2 (N22310, N22309, N13743);
nor NOR4 (N22311, N22294, N21413, N21711, N8234);
or OR4 (N22312, N22284, N8003, N10956, N1553);
xor XOR2 (N22313, N22310, N11711);
nand NAND3 (N22314, N22308, N22200, N17342);
nor NOR2 (N22315, N22301, N18576);
or OR3 (N22316, N22295, N16447, N21031);
buf BUF1 (N22317, N22314);
not NOT1 (N22318, N22307);
nand NAND4 (N22319, N22311, N18771, N11772, N10285);
and AND2 (N22320, N22302, N17479);
xor XOR2 (N22321, N22318, N8805);
buf BUF1 (N22322, N22317);
and AND2 (N22323, N22312, N14556);
buf BUF1 (N22324, N22320);
or OR3 (N22325, N22319, N16393, N19723);
buf BUF1 (N22326, N22313);
or OR4 (N22327, N22325, N4364, N10332, N14736);
nand NAND2 (N22328, N22327, N12092);
and AND3 (N22329, N22321, N12765, N11907);
and AND3 (N22330, N22329, N17403, N19462);
and AND2 (N22331, N22316, N19512);
nand NAND2 (N22332, N22328, N17674);
and AND3 (N22333, N22332, N2804, N12682);
buf BUF1 (N22334, N22324);
or OR3 (N22335, N22331, N11794, N6615);
or OR2 (N22336, N22322, N16499);
nand NAND4 (N22337, N22335, N17580, N15147, N20324);
and AND4 (N22338, N22330, N19592, N18745, N6653);
nand NAND2 (N22339, N22336, N10249);
or OR4 (N22340, N22323, N21520, N5411, N5848);
xor XOR2 (N22341, N22338, N8209);
and AND3 (N22342, N22304, N16019, N15610);
or OR3 (N22343, N22334, N6449, N6715);
buf BUF1 (N22344, N22339);
not NOT1 (N22345, N22315);
and AND2 (N22346, N22326, N8456);
or OR2 (N22347, N22342, N17059);
and AND3 (N22348, N22347, N2085, N19380);
or OR4 (N22349, N22344, N17497, N2981, N8980);
and AND3 (N22350, N22305, N21234, N20905);
nor NOR2 (N22351, N22346, N15783);
buf BUF1 (N22352, N22341);
buf BUF1 (N22353, N22333);
xor XOR2 (N22354, N22350, N17676);
and AND4 (N22355, N22343, N963, N10196, N602);
not NOT1 (N22356, N22352);
nand NAND4 (N22357, N22340, N10075, N242, N660);
nor NOR3 (N22358, N22349, N21453, N11921);
or OR3 (N22359, N22345, N17916, N491);
xor XOR2 (N22360, N22358, N10772);
nand NAND4 (N22361, N22357, N5068, N9926, N8635);
not NOT1 (N22362, N22351);
nor NOR4 (N22363, N22355, N11656, N16067, N21382);
xor XOR2 (N22364, N22337, N651);
nor NOR4 (N22365, N22348, N21269, N1934, N9748);
or OR3 (N22366, N22365, N13601, N7718);
or OR3 (N22367, N22362, N18775, N21317);
not NOT1 (N22368, N22354);
or OR3 (N22369, N22366, N11785, N6537);
and AND2 (N22370, N22369, N12664);
and AND3 (N22371, N22367, N14200, N16283);
nand NAND2 (N22372, N22364, N9189);
not NOT1 (N22373, N22359);
xor XOR2 (N22374, N22353, N18931);
or OR3 (N22375, N22374, N18124, N4820);
xor XOR2 (N22376, N22372, N4886);
not NOT1 (N22377, N22371);
nand NAND2 (N22378, N22360, N19309);
nand NAND3 (N22379, N22370, N11120, N12264);
or OR3 (N22380, N22356, N12799, N6063);
xor XOR2 (N22381, N22380, N17502);
or OR2 (N22382, N22361, N14529);
not NOT1 (N22383, N22368);
nand NAND3 (N22384, N22363, N17460, N21245);
nor NOR4 (N22385, N22379, N4864, N16505, N22238);
buf BUF1 (N22386, N22376);
and AND4 (N22387, N22375, N8379, N13137, N20354);
or OR4 (N22388, N22385, N11538, N12962, N318);
or OR4 (N22389, N22383, N13850, N15016, N21648);
and AND3 (N22390, N22388, N16829, N11488);
nand NAND2 (N22391, N22389, N11828);
or OR4 (N22392, N22387, N16351, N15898, N1563);
buf BUF1 (N22393, N22386);
xor XOR2 (N22394, N22384, N13069);
buf BUF1 (N22395, N22394);
buf BUF1 (N22396, N22391);
buf BUF1 (N22397, N22377);
xor XOR2 (N22398, N22378, N13265);
nand NAND2 (N22399, N22393, N6562);
nor NOR4 (N22400, N22396, N18344, N11748, N17602);
nor NOR4 (N22401, N22399, N6819, N7621, N19794);
nand NAND2 (N22402, N22373, N10040);
not NOT1 (N22403, N22397);
or OR2 (N22404, N22400, N9729);
nor NOR4 (N22405, N22404, N21385, N7770, N7005);
nor NOR2 (N22406, N22395, N12084);
or OR4 (N22407, N22392, N3207, N9383, N4955);
or OR4 (N22408, N22390, N11963, N406, N14155);
or OR4 (N22409, N22401, N6669, N8026, N9007);
not NOT1 (N22410, N22407);
and AND3 (N22411, N22381, N12292, N9201);
and AND4 (N22412, N22410, N14985, N10032, N12332);
nor NOR3 (N22413, N22408, N15446, N13231);
xor XOR2 (N22414, N22411, N20366);
and AND4 (N22415, N22382, N21279, N291, N1227);
nand NAND2 (N22416, N22402, N13938);
nand NAND3 (N22417, N22414, N12918, N9034);
nand NAND3 (N22418, N22406, N13616, N17342);
buf BUF1 (N22419, N22415);
nand NAND2 (N22420, N22413, N3980);
nor NOR2 (N22421, N22417, N16249);
nor NOR3 (N22422, N22409, N10444, N9005);
nand NAND2 (N22423, N22412, N17523);
not NOT1 (N22424, N22419);
and AND4 (N22425, N22424, N20583, N22010, N20661);
xor XOR2 (N22426, N22425, N20572);
or OR3 (N22427, N22398, N21529, N14367);
buf BUF1 (N22428, N22423);
not NOT1 (N22429, N22403);
or OR4 (N22430, N22421, N5123, N5708, N6554);
nor NOR2 (N22431, N22420, N1195);
not NOT1 (N22432, N22430);
and AND4 (N22433, N22428, N11616, N16069, N12109);
not NOT1 (N22434, N22433);
buf BUF1 (N22435, N22431);
buf BUF1 (N22436, N22405);
buf BUF1 (N22437, N22432);
not NOT1 (N22438, N22427);
or OR2 (N22439, N22429, N9987);
and AND3 (N22440, N22426, N1822, N3388);
buf BUF1 (N22441, N22435);
nand NAND2 (N22442, N22418, N1888);
xor XOR2 (N22443, N22439, N21678);
not NOT1 (N22444, N22442);
xor XOR2 (N22445, N22436, N20147);
and AND3 (N22446, N22441, N19936, N2198);
xor XOR2 (N22447, N22422, N1609);
nand NAND3 (N22448, N22437, N4250, N9325);
nor NOR4 (N22449, N22448, N11365, N20377, N5586);
buf BUF1 (N22450, N22444);
and AND4 (N22451, N22440, N2188, N17142, N14890);
nand NAND4 (N22452, N22449, N19765, N11185, N5635);
nand NAND3 (N22453, N22450, N8640, N19251);
buf BUF1 (N22454, N22416);
buf BUF1 (N22455, N22454);
not NOT1 (N22456, N22445);
xor XOR2 (N22457, N22456, N17456);
and AND3 (N22458, N22438, N2968, N4606);
or OR3 (N22459, N22434, N5034, N13724);
nand NAND4 (N22460, N22443, N13099, N18498, N740);
xor XOR2 (N22461, N22459, N19470);
nor NOR4 (N22462, N22446, N12071, N19122, N2003);
xor XOR2 (N22463, N22458, N11502);
nand NAND4 (N22464, N22447, N6799, N11934, N14718);
and AND4 (N22465, N22451, N6720, N784, N1046);
and AND3 (N22466, N22455, N17204, N20312);
or OR4 (N22467, N22457, N17322, N10034, N3760);
buf BUF1 (N22468, N22464);
or OR4 (N22469, N22468, N15403, N14537, N11073);
not NOT1 (N22470, N22460);
buf BUF1 (N22471, N22466);
nor NOR3 (N22472, N22462, N19142, N11694);
not NOT1 (N22473, N22471);
not NOT1 (N22474, N22461);
nand NAND3 (N22475, N22453, N11576, N18727);
nand NAND3 (N22476, N22465, N12428, N15788);
nand NAND4 (N22477, N22476, N1610, N21710, N20059);
and AND2 (N22478, N22475, N13735);
nor NOR4 (N22479, N22474, N11516, N10051, N8462);
not NOT1 (N22480, N22479);
and AND3 (N22481, N22469, N4354, N21094);
xor XOR2 (N22482, N22472, N21945);
buf BUF1 (N22483, N22477);
not NOT1 (N22484, N22463);
and AND4 (N22485, N22473, N4976, N19366, N5339);
nand NAND3 (N22486, N22485, N6162, N21022);
not NOT1 (N22487, N22481);
or OR3 (N22488, N22470, N22317, N17013);
nor NOR4 (N22489, N22486, N13835, N22336, N3109);
nor NOR2 (N22490, N22480, N9598);
buf BUF1 (N22491, N22488);
or OR2 (N22492, N22487, N17368);
buf BUF1 (N22493, N22467);
not NOT1 (N22494, N22478);
not NOT1 (N22495, N22494);
not NOT1 (N22496, N22495);
not NOT1 (N22497, N22491);
buf BUF1 (N22498, N22497);
nor NOR4 (N22499, N22490, N18694, N13536, N16279);
buf BUF1 (N22500, N22499);
xor XOR2 (N22501, N22496, N14501);
buf BUF1 (N22502, N22484);
xor XOR2 (N22503, N22501, N12362);
buf BUF1 (N22504, N22452);
nand NAND3 (N22505, N22498, N19121, N16338);
buf BUF1 (N22506, N22493);
xor XOR2 (N22507, N22500, N21636);
nor NOR4 (N22508, N22507, N10654, N15454, N15419);
nor NOR3 (N22509, N22506, N10511, N16605);
xor XOR2 (N22510, N22508, N18933);
or OR2 (N22511, N22510, N14583);
xor XOR2 (N22512, N22483, N20038);
or OR3 (N22513, N22509, N19804, N20120);
not NOT1 (N22514, N22502);
and AND2 (N22515, N22514, N1822);
or OR3 (N22516, N22489, N9151, N5741);
nand NAND2 (N22517, N22511, N2458);
nand NAND4 (N22518, N22503, N11512, N13548, N13256);
nor NOR2 (N22519, N22515, N18263);
or OR3 (N22520, N22513, N713, N10074);
and AND2 (N22521, N22505, N4995);
nand NAND2 (N22522, N22482, N5316);
and AND2 (N22523, N22520, N20293);
buf BUF1 (N22524, N22521);
nor NOR2 (N22525, N22519, N16771);
nand NAND4 (N22526, N22518, N16537, N9346, N2174);
xor XOR2 (N22527, N22512, N19505);
buf BUF1 (N22528, N22526);
or OR4 (N22529, N22504, N9778, N21974, N14942);
nor NOR2 (N22530, N22522, N14757);
buf BUF1 (N22531, N22527);
xor XOR2 (N22532, N22525, N2094);
and AND4 (N22533, N22517, N14514, N22318, N1510);
not NOT1 (N22534, N22531);
xor XOR2 (N22535, N22530, N3042);
nor NOR4 (N22536, N22529, N14234, N17287, N19910);
nor NOR4 (N22537, N22516, N12836, N6333, N20316);
xor XOR2 (N22538, N22528, N14688);
nand NAND3 (N22539, N22492, N19207, N2128);
nand NAND4 (N22540, N22535, N6557, N9470, N13051);
nor NOR3 (N22541, N22523, N2991, N20779);
buf BUF1 (N22542, N22540);
and AND3 (N22543, N22536, N22157, N8804);
buf BUF1 (N22544, N22537);
buf BUF1 (N22545, N22533);
nand NAND4 (N22546, N22545, N21999, N9773, N5576);
or OR2 (N22547, N22539, N21882);
xor XOR2 (N22548, N22538, N4389);
buf BUF1 (N22549, N22547);
nor NOR2 (N22550, N22534, N8258);
xor XOR2 (N22551, N22550, N20343);
xor XOR2 (N22552, N22548, N903);
buf BUF1 (N22553, N22552);
and AND4 (N22554, N22549, N12211, N10235, N2678);
nand NAND3 (N22555, N22551, N281, N1743);
nor NOR3 (N22556, N22554, N21473, N19286);
nor NOR3 (N22557, N22546, N19788, N3569);
xor XOR2 (N22558, N22544, N12504);
and AND3 (N22559, N22556, N4220, N11001);
buf BUF1 (N22560, N22524);
and AND4 (N22561, N22553, N16720, N17098, N3236);
xor XOR2 (N22562, N22532, N16161);
not NOT1 (N22563, N22557);
xor XOR2 (N22564, N22543, N21907);
or OR2 (N22565, N22562, N8773);
and AND4 (N22566, N22559, N16566, N2002, N4070);
or OR3 (N22567, N22563, N11790, N18364);
buf BUF1 (N22568, N22565);
buf BUF1 (N22569, N22541);
buf BUF1 (N22570, N22555);
nand NAND4 (N22571, N22568, N3574, N11701, N6112);
or OR2 (N22572, N22564, N6373);
nand NAND3 (N22573, N22570, N21531, N18430);
nor NOR2 (N22574, N22567, N12021);
not NOT1 (N22575, N22572);
or OR3 (N22576, N22558, N21969, N3253);
or OR3 (N22577, N22573, N17678, N3321);
xor XOR2 (N22578, N22574, N3718);
nor NOR2 (N22579, N22561, N15563);
nor NOR2 (N22580, N22571, N15369);
or OR2 (N22581, N22578, N8057);
or OR4 (N22582, N22581, N8176, N21058, N4111);
not NOT1 (N22583, N22579);
nor NOR3 (N22584, N22566, N10585, N2913);
and AND4 (N22585, N22542, N20493, N19613, N19816);
or OR3 (N22586, N22560, N15094, N12320);
or OR2 (N22587, N22585, N10911);
nand NAND3 (N22588, N22580, N12808, N16116);
and AND2 (N22589, N22583, N19461);
not NOT1 (N22590, N22569);
not NOT1 (N22591, N22582);
nor NOR2 (N22592, N22577, N1277);
buf BUF1 (N22593, N22588);
nor NOR4 (N22594, N22576, N20579, N22004, N20224);
xor XOR2 (N22595, N22593, N16988);
not NOT1 (N22596, N22584);
nand NAND2 (N22597, N22589, N2478);
buf BUF1 (N22598, N22596);
nand NAND4 (N22599, N22575, N5394, N13820, N10144);
and AND4 (N22600, N22587, N4579, N1232, N21840);
and AND2 (N22601, N22592, N15611);
nor NOR4 (N22602, N22597, N1512, N6971, N3677);
xor XOR2 (N22603, N22602, N4135);
and AND2 (N22604, N22595, N22287);
not NOT1 (N22605, N22591);
or OR2 (N22606, N22600, N21981);
nand NAND2 (N22607, N22598, N9378);
nor NOR2 (N22608, N22594, N12346);
buf BUF1 (N22609, N22605);
buf BUF1 (N22610, N22606);
nand NAND3 (N22611, N22590, N15751, N8379);
xor XOR2 (N22612, N22611, N2024);
nand NAND2 (N22613, N22608, N4118);
nand NAND2 (N22614, N22586, N6571);
nor NOR2 (N22615, N22614, N8795);
and AND2 (N22616, N22609, N12742);
buf BUF1 (N22617, N22615);
nand NAND3 (N22618, N22617, N15153, N8944);
buf BUF1 (N22619, N22604);
nand NAND3 (N22620, N22607, N9399, N9229);
xor XOR2 (N22621, N22613, N21066);
not NOT1 (N22622, N22618);
not NOT1 (N22623, N22620);
nand NAND4 (N22624, N22619, N17268, N9867, N18380);
nor NOR4 (N22625, N22599, N21762, N8681, N14533);
xor XOR2 (N22626, N22601, N345);
xor XOR2 (N22627, N22610, N3774);
or OR2 (N22628, N22623, N22543);
nor NOR4 (N22629, N22626, N8348, N10887, N17377);
and AND4 (N22630, N22628, N18364, N5578, N17869);
not NOT1 (N22631, N22630);
and AND2 (N22632, N22603, N20271);
and AND4 (N22633, N22625, N6385, N16933, N12445);
xor XOR2 (N22634, N22624, N13012);
not NOT1 (N22635, N22622);
and AND3 (N22636, N22631, N21114, N21477);
and AND3 (N22637, N22629, N7017, N2145);
nand NAND2 (N22638, N22632, N17430);
xor XOR2 (N22639, N22637, N18232);
buf BUF1 (N22640, N22636);
nor NOR2 (N22641, N22621, N3526);
or OR3 (N22642, N22627, N18256, N10194);
buf BUF1 (N22643, N22612);
buf BUF1 (N22644, N22638);
and AND4 (N22645, N22635, N17024, N13439, N11723);
buf BUF1 (N22646, N22642);
and AND3 (N22647, N22643, N17189, N3759);
nand NAND3 (N22648, N22633, N4578, N16371);
not NOT1 (N22649, N22644);
buf BUF1 (N22650, N22647);
xor XOR2 (N22651, N22648, N3233);
buf BUF1 (N22652, N22645);
nor NOR2 (N22653, N22651, N19027);
nor NOR3 (N22654, N22639, N9675, N17751);
or OR4 (N22655, N22653, N15162, N16247, N7564);
nor NOR2 (N22656, N22654, N21156);
nor NOR2 (N22657, N22652, N7922);
nor NOR4 (N22658, N22634, N8534, N3875, N22305);
and AND3 (N22659, N22656, N13370, N5502);
xor XOR2 (N22660, N22659, N11572);
not NOT1 (N22661, N22649);
not NOT1 (N22662, N22646);
xor XOR2 (N22663, N22616, N20810);
and AND4 (N22664, N22641, N9436, N12786, N5568);
xor XOR2 (N22665, N22650, N8368);
xor XOR2 (N22666, N22661, N6218);
buf BUF1 (N22667, N22660);
buf BUF1 (N22668, N22657);
not NOT1 (N22669, N22665);
nor NOR3 (N22670, N22658, N10566, N16689);
nor NOR4 (N22671, N22662, N13512, N6480, N20602);
xor XOR2 (N22672, N22667, N5577);
nand NAND2 (N22673, N22666, N6041);
or OR3 (N22674, N22640, N101, N910);
nand NAND4 (N22675, N22655, N17648, N11954, N19916);
buf BUF1 (N22676, N22674);
or OR3 (N22677, N22672, N11548, N3515);
buf BUF1 (N22678, N22664);
nand NAND3 (N22679, N22670, N18481, N8073);
xor XOR2 (N22680, N22677, N18699);
xor XOR2 (N22681, N22679, N2449);
and AND3 (N22682, N22671, N10394, N18228);
or OR2 (N22683, N22675, N1645);
and AND4 (N22684, N22669, N3535, N7456, N19554);
buf BUF1 (N22685, N22684);
xor XOR2 (N22686, N22680, N17657);
nand NAND4 (N22687, N22673, N13769, N462, N19564);
nand NAND4 (N22688, N22678, N10463, N10065, N388);
nand NAND2 (N22689, N22682, N2096);
or OR2 (N22690, N22687, N4421);
nand NAND4 (N22691, N22686, N18477, N825, N16236);
nand NAND2 (N22692, N22691, N2126);
nand NAND4 (N22693, N22692, N16393, N8069, N1859);
nand NAND2 (N22694, N22689, N787);
nor NOR2 (N22695, N22676, N12945);
and AND2 (N22696, N22693, N4344);
or OR2 (N22697, N22690, N13855);
and AND3 (N22698, N22688, N7884, N17317);
xor XOR2 (N22699, N22694, N13769);
not NOT1 (N22700, N22699);
nor NOR2 (N22701, N22697, N8957);
not NOT1 (N22702, N22685);
buf BUF1 (N22703, N22696);
and AND3 (N22704, N22668, N12707, N2591);
or OR2 (N22705, N22702, N11655);
and AND4 (N22706, N22681, N13276, N3176, N19457);
xor XOR2 (N22707, N22703, N3772);
xor XOR2 (N22708, N22700, N2851);
not NOT1 (N22709, N22695);
buf BUF1 (N22710, N22707);
buf BUF1 (N22711, N22708);
nor NOR4 (N22712, N22709, N13706, N15380, N1745);
not NOT1 (N22713, N22711);
xor XOR2 (N22714, N22683, N8130);
or OR2 (N22715, N22705, N1318);
and AND4 (N22716, N22663, N18163, N19225, N14556);
nand NAND3 (N22717, N22715, N2207, N8571);
buf BUF1 (N22718, N22706);
nor NOR2 (N22719, N22698, N13181);
and AND4 (N22720, N22718, N21860, N158, N1279);
nor NOR3 (N22721, N22716, N14402, N8348);
nor NOR2 (N22722, N22719, N2856);
and AND3 (N22723, N22722, N17364, N6454);
xor XOR2 (N22724, N22721, N17543);
buf BUF1 (N22725, N22704);
nand NAND2 (N22726, N22712, N3868);
not NOT1 (N22727, N22713);
nand NAND2 (N22728, N22714, N5372);
not NOT1 (N22729, N22727);
nand NAND3 (N22730, N22717, N210, N13595);
not NOT1 (N22731, N22730);
not NOT1 (N22732, N22701);
xor XOR2 (N22733, N22732, N21200);
nor NOR4 (N22734, N22728, N7186, N970, N7704);
buf BUF1 (N22735, N22731);
nand NAND4 (N22736, N22733, N1245, N1574, N16825);
or OR4 (N22737, N22736, N18195, N17442, N16331);
not NOT1 (N22738, N22737);
xor XOR2 (N22739, N22723, N10867);
and AND4 (N22740, N22726, N15635, N17327, N5558);
nor NOR3 (N22741, N22740, N6071, N16800);
buf BUF1 (N22742, N22734);
xor XOR2 (N22743, N22729, N5293);
not NOT1 (N22744, N22724);
xor XOR2 (N22745, N22744, N7896);
and AND2 (N22746, N22725, N14612);
not NOT1 (N22747, N22720);
buf BUF1 (N22748, N22739);
not NOT1 (N22749, N22745);
and AND2 (N22750, N22738, N20427);
nor NOR3 (N22751, N22741, N3816, N922);
or OR2 (N22752, N22748, N10306);
buf BUF1 (N22753, N22752);
nor NOR3 (N22754, N22747, N6913, N9519);
buf BUF1 (N22755, N22735);
or OR2 (N22756, N22750, N5552);
or OR2 (N22757, N22749, N11746);
and AND4 (N22758, N22753, N14015, N10353, N19242);
buf BUF1 (N22759, N22756);
buf BUF1 (N22760, N22758);
not NOT1 (N22761, N22757);
or OR4 (N22762, N22761, N8402, N17271, N10387);
or OR2 (N22763, N22742, N6107);
xor XOR2 (N22764, N22754, N12102);
not NOT1 (N22765, N22746);
nor NOR2 (N22766, N22765, N10758);
buf BUF1 (N22767, N22755);
not NOT1 (N22768, N22751);
nor NOR2 (N22769, N22710, N11034);
buf BUF1 (N22770, N22760);
and AND4 (N22771, N22743, N8260, N22038, N2693);
buf BUF1 (N22772, N22770);
not NOT1 (N22773, N22762);
buf BUF1 (N22774, N22759);
buf BUF1 (N22775, N22763);
nor NOR4 (N22776, N22766, N3961, N4632, N3835);
nor NOR3 (N22777, N22776, N6736, N21079);
nand NAND4 (N22778, N22767, N19950, N15795, N9394);
or OR2 (N22779, N22777, N15444);
and AND3 (N22780, N22773, N9619, N22185);
and AND3 (N22781, N22771, N15523, N19365);
or OR4 (N22782, N22772, N2531, N7989, N19332);
not NOT1 (N22783, N22764);
nor NOR3 (N22784, N22782, N14670, N20862);
not NOT1 (N22785, N22769);
xor XOR2 (N22786, N22785, N4415);
nand NAND3 (N22787, N22779, N20480, N18047);
not NOT1 (N22788, N22768);
not NOT1 (N22789, N22783);
and AND2 (N22790, N22784, N22010);
and AND3 (N22791, N22786, N8735, N13189);
nand NAND4 (N22792, N22788, N14522, N8392, N17346);
not NOT1 (N22793, N22789);
not NOT1 (N22794, N22793);
nor NOR2 (N22795, N22790, N16976);
not NOT1 (N22796, N22778);
or OR3 (N22797, N22774, N21726, N20411);
buf BUF1 (N22798, N22787);
nor NOR4 (N22799, N22791, N8723, N8302, N4307);
nor NOR2 (N22800, N22797, N14795);
xor XOR2 (N22801, N22800, N12125);
and AND4 (N22802, N22792, N21225, N8657, N766);
and AND4 (N22803, N22802, N3932, N15630, N18118);
and AND4 (N22804, N22803, N15251, N19851, N19712);
nor NOR4 (N22805, N22799, N7591, N12809, N16923);
nor NOR2 (N22806, N22796, N6576);
nand NAND3 (N22807, N22775, N19754, N7210);
not NOT1 (N22808, N22798);
or OR4 (N22809, N22807, N17498, N5603, N6704);
and AND4 (N22810, N22806, N5692, N17307, N20300);
buf BUF1 (N22811, N22794);
xor XOR2 (N22812, N22795, N6998);
or OR2 (N22813, N22811, N21944);
nand NAND4 (N22814, N22805, N11436, N20853, N1456);
xor XOR2 (N22815, N22804, N1038);
buf BUF1 (N22816, N22812);
buf BUF1 (N22817, N22813);
not NOT1 (N22818, N22809);
nand NAND2 (N22819, N22816, N5288);
not NOT1 (N22820, N22818);
and AND2 (N22821, N22810, N9726);
and AND4 (N22822, N22781, N16877, N10837, N2718);
not NOT1 (N22823, N22819);
or OR4 (N22824, N22814, N2592, N12097, N13282);
buf BUF1 (N22825, N22815);
nand NAND4 (N22826, N22823, N21520, N19409, N13117);
xor XOR2 (N22827, N22821, N462);
xor XOR2 (N22828, N22824, N16222);
and AND4 (N22829, N22780, N9503, N2136, N9265);
or OR2 (N22830, N22808, N22362);
xor XOR2 (N22831, N22827, N22676);
nor NOR4 (N22832, N22830, N6114, N20178, N2544);
not NOT1 (N22833, N22826);
xor XOR2 (N22834, N22832, N10750);
not NOT1 (N22835, N22833);
not NOT1 (N22836, N22828);
buf BUF1 (N22837, N22835);
buf BUF1 (N22838, N22820);
nand NAND4 (N22839, N22829, N21459, N18902, N16808);
xor XOR2 (N22840, N22837, N5946);
nor NOR4 (N22841, N22822, N11284, N1260, N8759);
or OR2 (N22842, N22840, N22252);
buf BUF1 (N22843, N22825);
or OR3 (N22844, N22801, N1836, N8710);
buf BUF1 (N22845, N22838);
xor XOR2 (N22846, N22836, N10002);
and AND3 (N22847, N22841, N16061, N20521);
nand NAND2 (N22848, N22846, N995);
not NOT1 (N22849, N22842);
xor XOR2 (N22850, N22843, N6595);
nand NAND3 (N22851, N22850, N4820, N13267);
xor XOR2 (N22852, N22834, N359);
or OR2 (N22853, N22844, N21042);
xor XOR2 (N22854, N22845, N8940);
not NOT1 (N22855, N22853);
and AND3 (N22856, N22852, N7033, N15068);
or OR4 (N22857, N22849, N7411, N15953, N15917);
buf BUF1 (N22858, N22854);
nor NOR2 (N22859, N22858, N20400);
or OR2 (N22860, N22831, N642);
xor XOR2 (N22861, N22851, N5146);
xor XOR2 (N22862, N22859, N19485);
nand NAND2 (N22863, N22839, N12557);
or OR4 (N22864, N22855, N10662, N7428, N6638);
nor NOR3 (N22865, N22847, N5965, N18573);
buf BUF1 (N22866, N22856);
and AND2 (N22867, N22860, N11154);
buf BUF1 (N22868, N22862);
xor XOR2 (N22869, N22863, N18052);
xor XOR2 (N22870, N22868, N7344);
nor NOR3 (N22871, N22857, N13656, N21287);
xor XOR2 (N22872, N22871, N4141);
or OR2 (N22873, N22864, N8501);
xor XOR2 (N22874, N22867, N8235);
nor NOR3 (N22875, N22873, N11145, N6123);
or OR4 (N22876, N22866, N2854, N17508, N4656);
and AND4 (N22877, N22865, N12909, N14848, N16983);
or OR2 (N22878, N22861, N4861);
or OR3 (N22879, N22872, N3529, N950);
nand NAND3 (N22880, N22875, N7837, N22517);
nor NOR2 (N22881, N22848, N2018);
or OR2 (N22882, N22877, N8220);
nor NOR3 (N22883, N22869, N16306, N21510);
buf BUF1 (N22884, N22876);
xor XOR2 (N22885, N22817, N19804);
nand NAND3 (N22886, N22882, N17945, N15487);
and AND2 (N22887, N22874, N1944);
buf BUF1 (N22888, N22880);
or OR2 (N22889, N22879, N842);
buf BUF1 (N22890, N22878);
or OR4 (N22891, N22887, N16471, N10867, N7182);
not NOT1 (N22892, N22886);
not NOT1 (N22893, N22870);
or OR3 (N22894, N22893, N13121, N13002);
nand NAND2 (N22895, N22894, N21761);
nor NOR3 (N22896, N22890, N1033, N7434);
xor XOR2 (N22897, N22896, N13698);
and AND3 (N22898, N22888, N16057, N10381);
nor NOR4 (N22899, N22889, N9948, N21466, N4905);
or OR2 (N22900, N22881, N9792);
nand NAND3 (N22901, N22897, N1780, N21886);
buf BUF1 (N22902, N22884);
nor NOR3 (N22903, N22891, N3017, N5021);
or OR2 (N22904, N22895, N19049);
buf BUF1 (N22905, N22901);
nor NOR4 (N22906, N22885, N22514, N12221, N14173);
or OR2 (N22907, N22903, N10486);
not NOT1 (N22908, N22892);
nand NAND3 (N22909, N22900, N2688, N3710);
nand NAND2 (N22910, N22899, N18581);
buf BUF1 (N22911, N22909);
and AND4 (N22912, N22908, N6753, N19715, N5235);
xor XOR2 (N22913, N22902, N14464);
not NOT1 (N22914, N22907);
nand NAND3 (N22915, N22898, N21618, N3393);
or OR4 (N22916, N22883, N16595, N10398, N12022);
and AND3 (N22917, N22910, N20161, N22797);
nor NOR4 (N22918, N22914, N19965, N3576, N11949);
nor NOR4 (N22919, N22904, N14419, N15513, N3324);
or OR3 (N22920, N22912, N4083, N10158);
or OR2 (N22921, N22913, N6079);
buf BUF1 (N22922, N22921);
nor NOR4 (N22923, N22915, N22220, N1733, N8994);
and AND4 (N22924, N22920, N10346, N3676, N9376);
xor XOR2 (N22925, N22917, N12904);
nand NAND2 (N22926, N22916, N16715);
buf BUF1 (N22927, N22905);
nor NOR4 (N22928, N22911, N7134, N10681, N17349);
nor NOR4 (N22929, N22925, N2248, N12727, N17144);
nor NOR3 (N22930, N22924, N12597, N22414);
or OR4 (N22931, N22927, N22321, N18543, N12750);
and AND4 (N22932, N22906, N20653, N15022, N20342);
buf BUF1 (N22933, N22932);
and AND4 (N22934, N22931, N17100, N19262, N10450);
or OR3 (N22935, N22934, N16975, N21341);
buf BUF1 (N22936, N22935);
or OR3 (N22937, N22933, N15041, N4543);
xor XOR2 (N22938, N22918, N17355);
or OR4 (N22939, N22922, N18183, N21738, N7359);
buf BUF1 (N22940, N22930);
and AND2 (N22941, N22937, N7701);
nor NOR2 (N22942, N22939, N12698);
nor NOR4 (N22943, N22940, N17536, N3156, N4970);
not NOT1 (N22944, N22923);
and AND3 (N22945, N22941, N8353, N20610);
not NOT1 (N22946, N22942);
or OR4 (N22947, N22936, N9075, N5918, N3058);
or OR3 (N22948, N22919, N9582, N4252);
nand NAND4 (N22949, N22944, N7200, N455, N12686);
nor NOR3 (N22950, N22948, N14710, N11759);
xor XOR2 (N22951, N22949, N20464);
xor XOR2 (N22952, N22950, N9893);
and AND3 (N22953, N22946, N13581, N15097);
and AND4 (N22954, N22928, N5616, N3188, N20316);
nor NOR4 (N22955, N22943, N1875, N12009, N18474);
xor XOR2 (N22956, N22945, N22552);
not NOT1 (N22957, N22951);
or OR3 (N22958, N22947, N21865, N2917);
and AND2 (N22959, N22955, N7045);
buf BUF1 (N22960, N22956);
or OR2 (N22961, N22952, N7070);
or OR4 (N22962, N22957, N14064, N3001, N14378);
not NOT1 (N22963, N22953);
or OR4 (N22964, N22960, N9566, N14620, N15595);
and AND2 (N22965, N22938, N8040);
nand NAND4 (N22966, N22963, N17199, N230, N22738);
xor XOR2 (N22967, N22929, N16592);
not NOT1 (N22968, N22966);
not NOT1 (N22969, N22954);
buf BUF1 (N22970, N22959);
nand NAND4 (N22971, N22958, N13353, N2943, N3271);
and AND4 (N22972, N22968, N15419, N18119, N2998);
and AND2 (N22973, N22971, N735);
not NOT1 (N22974, N22970);
and AND4 (N22975, N22969, N15834, N7567, N19086);
not NOT1 (N22976, N22965);
nor NOR2 (N22977, N22972, N17494);
or OR3 (N22978, N22974, N14680, N19769);
and AND2 (N22979, N22964, N7360);
xor XOR2 (N22980, N22979, N13986);
not NOT1 (N22981, N22962);
buf BUF1 (N22982, N22961);
nand NAND2 (N22983, N22980, N8984);
nand NAND3 (N22984, N22926, N6254, N5209);
or OR4 (N22985, N22983, N9701, N2431, N10668);
or OR2 (N22986, N22976, N6463);
nand NAND4 (N22987, N22975, N109, N1029, N21394);
nor NOR2 (N22988, N22981, N13073);
nand NAND4 (N22989, N22988, N15142, N14073, N18894);
or OR4 (N22990, N22978, N18732, N22435, N16125);
or OR2 (N22991, N22987, N14387);
nand NAND4 (N22992, N22991, N20861, N8835, N21966);
and AND2 (N22993, N22986, N3102);
not NOT1 (N22994, N22993);
not NOT1 (N22995, N22967);
xor XOR2 (N22996, N22985, N9465);
and AND3 (N22997, N22996, N13636, N11719);
not NOT1 (N22998, N22994);
and AND2 (N22999, N22982, N12756);
or OR4 (N23000, N22973, N2498, N21747, N14853);
or OR2 (N23001, N22990, N13672);
and AND4 (N23002, N23000, N6754, N3631, N17748);
xor XOR2 (N23003, N22995, N11654);
xor XOR2 (N23004, N22989, N13769);
buf BUF1 (N23005, N23002);
and AND4 (N23006, N22998, N4992, N22436, N830);
not NOT1 (N23007, N23006);
nand NAND2 (N23008, N23007, N21176);
nor NOR3 (N23009, N23005, N17034, N8920);
nor NOR4 (N23010, N22999, N20477, N12226, N15032);
and AND2 (N23011, N22997, N858);
nand NAND4 (N23012, N23001, N9003, N1939, N9920);
xor XOR2 (N23013, N23010, N17070);
not NOT1 (N23014, N23008);
nor NOR3 (N23015, N22984, N3992, N1660);
not NOT1 (N23016, N23013);
xor XOR2 (N23017, N23012, N18984);
buf BUF1 (N23018, N23011);
not NOT1 (N23019, N22992);
not NOT1 (N23020, N23018);
nor NOR3 (N23021, N23009, N9395, N20275);
buf BUF1 (N23022, N23004);
nor NOR2 (N23023, N23017, N9745);
nand NAND4 (N23024, N23003, N17445, N7323, N16739);
and AND3 (N23025, N23021, N1061, N10338);
buf BUF1 (N23026, N22977);
or OR4 (N23027, N23026, N2382, N21392, N17083);
not NOT1 (N23028, N23024);
nor NOR4 (N23029, N23027, N21127, N16806, N7381);
or OR2 (N23030, N23020, N1616);
nand NAND4 (N23031, N23028, N10138, N3064, N5964);
nand NAND3 (N23032, N23029, N921, N2881);
nand NAND2 (N23033, N23025, N14087);
or OR2 (N23034, N23030, N15610);
nor NOR4 (N23035, N23022, N14463, N740, N15938);
or OR2 (N23036, N23015, N21332);
nand NAND4 (N23037, N23014, N4582, N21609, N8116);
not NOT1 (N23038, N23031);
buf BUF1 (N23039, N23033);
nand NAND4 (N23040, N23035, N14822, N20747, N4428);
nand NAND4 (N23041, N23034, N20334, N11609, N5033);
nor NOR4 (N23042, N23032, N9559, N3715, N14761);
buf BUF1 (N23043, N23019);
nor NOR3 (N23044, N23043, N14530, N1926);
or OR4 (N23045, N23041, N7669, N3349, N3646);
xor XOR2 (N23046, N23039, N14526);
not NOT1 (N23047, N23036);
nand NAND2 (N23048, N23037, N21633);
nand NAND3 (N23049, N23016, N1086, N8503);
not NOT1 (N23050, N23038);
nor NOR3 (N23051, N23040, N5000, N13947);
or OR4 (N23052, N23044, N6867, N19496, N14079);
nand NAND2 (N23053, N23023, N15845);
nor NOR4 (N23054, N23047, N19136, N18714, N17550);
xor XOR2 (N23055, N23050, N18768);
not NOT1 (N23056, N23042);
or OR2 (N23057, N23048, N1328);
buf BUF1 (N23058, N23051);
nor NOR4 (N23059, N23055, N11125, N21657, N21676);
nor NOR4 (N23060, N23049, N3930, N10806, N19753);
nand NAND3 (N23061, N23046, N19127, N120);
nand NAND3 (N23062, N23057, N4526, N21785);
or OR2 (N23063, N23059, N10940);
buf BUF1 (N23064, N23045);
not NOT1 (N23065, N23053);
nor NOR3 (N23066, N23052, N21511, N1412);
buf BUF1 (N23067, N23061);
nor NOR4 (N23068, N23058, N3084, N14535, N17611);
and AND3 (N23069, N23065, N13853, N3071);
not NOT1 (N23070, N23067);
xor XOR2 (N23071, N23056, N17649);
buf BUF1 (N23072, N23068);
not NOT1 (N23073, N23062);
nor NOR2 (N23074, N23060, N63);
or OR3 (N23075, N23074, N1918, N6117);
or OR3 (N23076, N23070, N7807, N2925);
nor NOR4 (N23077, N23076, N17599, N10371, N22721);
nor NOR3 (N23078, N23077, N2629, N10774);
or OR2 (N23079, N23054, N9297);
buf BUF1 (N23080, N23069);
nor NOR2 (N23081, N23080, N21551);
nand NAND4 (N23082, N23078, N20311, N17028, N10348);
not NOT1 (N23083, N23081);
nand NAND2 (N23084, N23083, N6627);
nor NOR2 (N23085, N23082, N11254);
and AND3 (N23086, N23073, N16364, N20724);
buf BUF1 (N23087, N23064);
nor NOR4 (N23088, N23087, N1134, N19068, N14695);
not NOT1 (N23089, N23088);
and AND2 (N23090, N23084, N10697);
nor NOR3 (N23091, N23086, N6467, N17063);
buf BUF1 (N23092, N23091);
nor NOR3 (N23093, N23090, N18463, N19773);
not NOT1 (N23094, N23079);
nand NAND3 (N23095, N23071, N21689, N526);
nand NAND2 (N23096, N23085, N7488);
xor XOR2 (N23097, N23093, N3638);
and AND4 (N23098, N23075, N10925, N18394, N1608);
nand NAND2 (N23099, N23063, N18429);
buf BUF1 (N23100, N23096);
or OR3 (N23101, N23094, N999, N17241);
xor XOR2 (N23102, N23100, N2090);
or OR4 (N23103, N23097, N12811, N10051, N9727);
nand NAND4 (N23104, N23095, N4865, N5281, N5697);
nor NOR4 (N23105, N23098, N13115, N8945, N11945);
buf BUF1 (N23106, N23105);
or OR2 (N23107, N23099, N15215);
nor NOR2 (N23108, N23072, N9820);
buf BUF1 (N23109, N23108);
buf BUF1 (N23110, N23106);
nor NOR2 (N23111, N23092, N12748);
nand NAND2 (N23112, N23109, N11585);
and AND3 (N23113, N23111, N11468, N407);
not NOT1 (N23114, N23113);
buf BUF1 (N23115, N23110);
not NOT1 (N23116, N23101);
nand NAND3 (N23117, N23112, N8938, N21026);
and AND2 (N23118, N23103, N13876);
or OR3 (N23119, N23107, N22520, N9049);
xor XOR2 (N23120, N23115, N11577);
nand NAND4 (N23121, N23066, N8019, N6734, N17171);
xor XOR2 (N23122, N23121, N17331);
not NOT1 (N23123, N23114);
not NOT1 (N23124, N23118);
not NOT1 (N23125, N23123);
buf BUF1 (N23126, N23119);
or OR3 (N23127, N23122, N16336, N7775);
or OR4 (N23128, N23102, N14041, N11456, N14701);
not NOT1 (N23129, N23104);
not NOT1 (N23130, N23117);
nor NOR3 (N23131, N23124, N18397, N19425);
nor NOR4 (N23132, N23131, N22650, N10995, N16875);
nand NAND4 (N23133, N23116, N22708, N17122, N5346);
buf BUF1 (N23134, N23130);
nor NOR4 (N23135, N23127, N5332, N6472, N13009);
and AND3 (N23136, N23135, N11405, N22073);
not NOT1 (N23137, N23129);
and AND2 (N23138, N23137, N7330);
or OR2 (N23139, N23089, N8643);
xor XOR2 (N23140, N23128, N14718);
not NOT1 (N23141, N23120);
not NOT1 (N23142, N23132);
or OR2 (N23143, N23142, N22684);
and AND3 (N23144, N23138, N19237, N19754);
and AND2 (N23145, N23139, N18956);
and AND4 (N23146, N23136, N13122, N20323, N403);
and AND4 (N23147, N23145, N15006, N465, N22764);
not NOT1 (N23148, N23143);
not NOT1 (N23149, N23133);
and AND3 (N23150, N23126, N4140, N22991);
not NOT1 (N23151, N23150);
and AND4 (N23152, N23146, N8399, N8959, N9688);
nor NOR2 (N23153, N23125, N21586);
buf BUF1 (N23154, N23147);
and AND3 (N23155, N23144, N18822, N10077);
not NOT1 (N23156, N23148);
and AND3 (N23157, N23155, N9793, N2115);
xor XOR2 (N23158, N23156, N17081);
nor NOR3 (N23159, N23149, N16834, N18414);
buf BUF1 (N23160, N23159);
and AND4 (N23161, N23153, N11452, N12806, N1835);
buf BUF1 (N23162, N23154);
and AND4 (N23163, N23140, N4859, N15120, N7334);
nor NOR2 (N23164, N23157, N19021);
xor XOR2 (N23165, N23151, N105);
xor XOR2 (N23166, N23162, N1419);
buf BUF1 (N23167, N23141);
nor NOR2 (N23168, N23158, N19971);
nor NOR3 (N23169, N23134, N13569, N15739);
xor XOR2 (N23170, N23163, N6988);
xor XOR2 (N23171, N23161, N15680);
buf BUF1 (N23172, N23169);
and AND3 (N23173, N23160, N16777, N16944);
nand NAND2 (N23174, N23164, N11357);
not NOT1 (N23175, N23172);
nor NOR4 (N23176, N23170, N3473, N20967, N21160);
nor NOR3 (N23177, N23174, N15420, N6972);
buf BUF1 (N23178, N23173);
nand NAND2 (N23179, N23171, N5911);
buf BUF1 (N23180, N23175);
or OR3 (N23181, N23165, N1234, N2129);
or OR4 (N23182, N23152, N3376, N18632, N20106);
not NOT1 (N23183, N23177);
and AND4 (N23184, N23179, N15027, N18093, N17896);
not NOT1 (N23185, N23178);
nor NOR3 (N23186, N23180, N17330, N2712);
and AND4 (N23187, N23181, N14227, N20935, N19378);
nand NAND3 (N23188, N23167, N13427, N15921);
nor NOR2 (N23189, N23188, N18454);
nand NAND2 (N23190, N23189, N3284);
not NOT1 (N23191, N23186);
and AND3 (N23192, N23191, N16866, N7957);
nand NAND3 (N23193, N23182, N5655, N855);
buf BUF1 (N23194, N23184);
nor NOR3 (N23195, N23190, N11475, N9944);
buf BUF1 (N23196, N23195);
nor NOR3 (N23197, N23194, N9250, N4117);
and AND4 (N23198, N23197, N645, N18379, N3112);
and AND3 (N23199, N23176, N9340, N5362);
not NOT1 (N23200, N23193);
buf BUF1 (N23201, N23187);
and AND4 (N23202, N23198, N19597, N14920, N10319);
nand NAND4 (N23203, N23200, N21942, N4008, N11779);
nand NAND3 (N23204, N23183, N2904, N4797);
and AND2 (N23205, N23166, N19023);
xor XOR2 (N23206, N23192, N21988);
buf BUF1 (N23207, N23202);
not NOT1 (N23208, N23206);
buf BUF1 (N23209, N23203);
or OR3 (N23210, N23196, N16214, N7420);
buf BUF1 (N23211, N23208);
buf BUF1 (N23212, N23209);
and AND4 (N23213, N23207, N13016, N723, N14425);
xor XOR2 (N23214, N23185, N13681);
xor XOR2 (N23215, N23211, N12065);
nor NOR3 (N23216, N23201, N13842, N6181);
xor XOR2 (N23217, N23199, N22987);
or OR4 (N23218, N23215, N5369, N14540, N1804);
nor NOR3 (N23219, N23218, N16359, N20332);
buf BUF1 (N23220, N23214);
not NOT1 (N23221, N23212);
nor NOR4 (N23222, N23220, N2361, N5965, N8264);
or OR4 (N23223, N23222, N1826, N8980, N857);
nand NAND3 (N23224, N23217, N9903, N257);
nand NAND2 (N23225, N23224, N1209);
not NOT1 (N23226, N23219);
buf BUF1 (N23227, N23205);
nand NAND2 (N23228, N23210, N18116);
not NOT1 (N23229, N23213);
xor XOR2 (N23230, N23227, N144);
and AND4 (N23231, N23230, N10191, N7165, N22255);
xor XOR2 (N23232, N23226, N11594);
or OR2 (N23233, N23228, N16521);
or OR4 (N23234, N23223, N10648, N22382, N7738);
buf BUF1 (N23235, N23225);
buf BUF1 (N23236, N23229);
nor NOR2 (N23237, N23236, N14225);
xor XOR2 (N23238, N23231, N21114);
not NOT1 (N23239, N23234);
nand NAND4 (N23240, N23221, N17258, N15635, N20771);
nand NAND3 (N23241, N23235, N18068, N17907);
buf BUF1 (N23242, N23239);
and AND3 (N23243, N23241, N18074, N19118);
xor XOR2 (N23244, N23233, N4326);
nor NOR4 (N23245, N23204, N21335, N15683, N20493);
and AND3 (N23246, N23237, N3310, N6766);
nand NAND2 (N23247, N23242, N2351);
nand NAND2 (N23248, N23243, N14027);
and AND3 (N23249, N23238, N10745, N18931);
and AND2 (N23250, N23244, N17357);
buf BUF1 (N23251, N23232);
xor XOR2 (N23252, N23246, N14061);
and AND2 (N23253, N23252, N137);
or OR2 (N23254, N23240, N3638);
and AND4 (N23255, N23168, N16866, N19961, N17424);
xor XOR2 (N23256, N23254, N6591);
buf BUF1 (N23257, N23216);
nor NOR4 (N23258, N23247, N18256, N16717, N12249);
or OR2 (N23259, N23250, N17413);
or OR3 (N23260, N23251, N1555, N19878);
nor NOR3 (N23261, N23253, N2127, N1518);
buf BUF1 (N23262, N23245);
nand NAND2 (N23263, N23248, N7111);
not NOT1 (N23264, N23257);
buf BUF1 (N23265, N23259);
buf BUF1 (N23266, N23256);
xor XOR2 (N23267, N23265, N21353);
not NOT1 (N23268, N23260);
not NOT1 (N23269, N23262);
not NOT1 (N23270, N23268);
and AND3 (N23271, N23269, N20800, N20900);
nand NAND2 (N23272, N23258, N16553);
xor XOR2 (N23273, N23264, N14765);
and AND2 (N23274, N23271, N19347);
and AND4 (N23275, N23274, N21116, N20593, N11991);
nand NAND3 (N23276, N23272, N13441, N9692);
and AND3 (N23277, N23276, N18504, N9118);
xor XOR2 (N23278, N23273, N17200);
or OR3 (N23279, N23270, N20957, N16067);
xor XOR2 (N23280, N23278, N11131);
nor NOR2 (N23281, N23249, N11207);
nor NOR2 (N23282, N23281, N22789);
and AND4 (N23283, N23263, N13044, N9622, N20221);
nor NOR3 (N23284, N23280, N3524, N12558);
not NOT1 (N23285, N23267);
buf BUF1 (N23286, N23277);
nand NAND2 (N23287, N23284, N17287);
buf BUF1 (N23288, N23285);
not NOT1 (N23289, N23286);
buf BUF1 (N23290, N23287);
nor NOR3 (N23291, N23266, N6068, N17313);
or OR2 (N23292, N23288, N11107);
or OR3 (N23293, N23289, N21996, N4675);
nor NOR2 (N23294, N23293, N10844);
xor XOR2 (N23295, N23290, N4550);
and AND2 (N23296, N23282, N3200);
nand NAND3 (N23297, N23261, N15875, N19987);
nor NOR2 (N23298, N23297, N9566);
xor XOR2 (N23299, N23292, N6718);
or OR2 (N23300, N23295, N6036);
nor NOR4 (N23301, N23300, N6204, N1462, N22664);
or OR2 (N23302, N23301, N19364);
not NOT1 (N23303, N23298);
or OR4 (N23304, N23275, N4397, N9532, N7727);
nand NAND4 (N23305, N23294, N11229, N22335, N2333);
xor XOR2 (N23306, N23291, N20953);
or OR2 (N23307, N23299, N7706);
nor NOR2 (N23308, N23283, N7116);
and AND3 (N23309, N23308, N11123, N5471);
buf BUF1 (N23310, N23304);
and AND3 (N23311, N23302, N13207, N11270);
and AND3 (N23312, N23255, N22832, N11042);
or OR2 (N23313, N23311, N10482);
xor XOR2 (N23314, N23306, N14393);
buf BUF1 (N23315, N23309);
nor NOR4 (N23316, N23315, N20714, N21558, N11600);
buf BUF1 (N23317, N23307);
and AND3 (N23318, N23313, N19867, N624);
xor XOR2 (N23319, N23316, N16398);
buf BUF1 (N23320, N23303);
nand NAND2 (N23321, N23310, N9144);
not NOT1 (N23322, N23279);
or OR4 (N23323, N23312, N21832, N4759, N661);
nand NAND3 (N23324, N23320, N3882, N7441);
not NOT1 (N23325, N23318);
nor NOR3 (N23326, N23325, N23059, N1894);
buf BUF1 (N23327, N23305);
nor NOR2 (N23328, N23317, N363);
and AND4 (N23329, N23323, N18369, N6497, N8298);
nand NAND4 (N23330, N23327, N3617, N22234, N15646);
and AND4 (N23331, N23328, N12595, N893, N18958);
nor NOR3 (N23332, N23322, N11048, N1524);
nand NAND2 (N23333, N23329, N20373);
and AND4 (N23334, N23321, N5176, N2865, N10599);
nand NAND3 (N23335, N23333, N18364, N8266);
buf BUF1 (N23336, N23330);
nor NOR4 (N23337, N23336, N18490, N22490, N19832);
xor XOR2 (N23338, N23331, N9154);
nand NAND3 (N23339, N23314, N2684, N23154);
nor NOR3 (N23340, N23334, N4309, N11899);
not NOT1 (N23341, N23339);
or OR2 (N23342, N23324, N7107);
and AND4 (N23343, N23319, N3989, N238, N20374);
or OR2 (N23344, N23338, N18988);
xor XOR2 (N23345, N23344, N17114);
nand NAND2 (N23346, N23345, N495);
nand NAND3 (N23347, N23342, N7365, N14097);
nor NOR3 (N23348, N23347, N703, N22103);
nand NAND4 (N23349, N23337, N8525, N12226, N18744);
nand NAND2 (N23350, N23332, N19648);
nor NOR4 (N23351, N23346, N18365, N9224, N3405);
xor XOR2 (N23352, N23341, N5179);
xor XOR2 (N23353, N23343, N4978);
buf BUF1 (N23354, N23349);
or OR4 (N23355, N23353, N22116, N22022, N10128);
buf BUF1 (N23356, N23340);
nand NAND4 (N23357, N23351, N10150, N22385, N13049);
xor XOR2 (N23358, N23356, N1132);
nand NAND4 (N23359, N23350, N7692, N7825, N15258);
or OR3 (N23360, N23348, N4496, N9531);
nand NAND3 (N23361, N23355, N9128, N19950);
nand NAND2 (N23362, N23354, N8971);
not NOT1 (N23363, N23359);
not NOT1 (N23364, N23360);
and AND3 (N23365, N23296, N4275, N3031);
not NOT1 (N23366, N23364);
nor NOR2 (N23367, N23365, N21630);
nor NOR3 (N23368, N23363, N38, N14718);
xor XOR2 (N23369, N23335, N9757);
nand NAND4 (N23370, N23357, N18508, N6006, N22932);
nor NOR2 (N23371, N23370, N16182);
nor NOR4 (N23372, N23358, N20512, N12017, N2894);
buf BUF1 (N23373, N23361);
buf BUF1 (N23374, N23366);
or OR2 (N23375, N23326, N1653);
xor XOR2 (N23376, N23374, N19376);
nor NOR3 (N23377, N23371, N13503, N20038);
nor NOR2 (N23378, N23368, N22339);
and AND4 (N23379, N23352, N4120, N15198, N249);
nor NOR2 (N23380, N23379, N11930);
buf BUF1 (N23381, N23369);
nor NOR2 (N23382, N23378, N17894);
not NOT1 (N23383, N23362);
buf BUF1 (N23384, N23381);
nand NAND4 (N23385, N23382, N8934, N6034, N12313);
xor XOR2 (N23386, N23377, N2898);
not NOT1 (N23387, N23380);
nor NOR2 (N23388, N23385, N22756);
nor NOR2 (N23389, N23384, N20374);
xor XOR2 (N23390, N23367, N19968);
and AND2 (N23391, N23387, N23217);
buf BUF1 (N23392, N23373);
and AND4 (N23393, N23388, N5240, N12471, N19492);
or OR4 (N23394, N23375, N5074, N542, N15088);
or OR2 (N23395, N23390, N19264);
nor NOR3 (N23396, N23393, N20780, N17468);
nor NOR2 (N23397, N23396, N20506);
not NOT1 (N23398, N23376);
and AND2 (N23399, N23372, N15696);
and AND2 (N23400, N23392, N15352);
xor XOR2 (N23401, N23397, N21829);
not NOT1 (N23402, N23386);
nand NAND3 (N23403, N23391, N8524, N5312);
not NOT1 (N23404, N23401);
not NOT1 (N23405, N23395);
nand NAND3 (N23406, N23394, N20263, N9981);
and AND4 (N23407, N23402, N15127, N9006, N19110);
xor XOR2 (N23408, N23403, N12268);
not NOT1 (N23409, N23408);
nand NAND4 (N23410, N23405, N21076, N758, N6950);
xor XOR2 (N23411, N23409, N21391);
nor NOR3 (N23412, N23407, N2977, N18296);
buf BUF1 (N23413, N23400);
buf BUF1 (N23414, N23383);
and AND3 (N23415, N23410, N17936, N609);
nor NOR2 (N23416, N23389, N9210);
xor XOR2 (N23417, N23399, N19313);
or OR3 (N23418, N23414, N22815, N4926);
nor NOR2 (N23419, N23406, N17474);
or OR4 (N23420, N23398, N11340, N16776, N18959);
and AND4 (N23421, N23415, N2883, N19311, N16635);
not NOT1 (N23422, N23417);
buf BUF1 (N23423, N23422);
not NOT1 (N23424, N23420);
not NOT1 (N23425, N23418);
not NOT1 (N23426, N23412);
nand NAND4 (N23427, N23426, N17180, N11033, N6164);
or OR4 (N23428, N23416, N6025, N15593, N7372);
buf BUF1 (N23429, N23423);
or OR2 (N23430, N23421, N6023);
xor XOR2 (N23431, N23404, N16579);
buf BUF1 (N23432, N23413);
and AND4 (N23433, N23432, N7844, N19466, N8791);
buf BUF1 (N23434, N23411);
xor XOR2 (N23435, N23429, N10432);
or OR4 (N23436, N23435, N6019, N8036, N9975);
nand NAND2 (N23437, N23431, N13782);
and AND4 (N23438, N23428, N13906, N5950, N16991);
and AND3 (N23439, N23430, N11765, N9211);
buf BUF1 (N23440, N23439);
xor XOR2 (N23441, N23434, N2725);
or OR2 (N23442, N23440, N7894);
not NOT1 (N23443, N23419);
and AND3 (N23444, N23443, N16019, N2071);
not NOT1 (N23445, N23427);
and AND3 (N23446, N23438, N8615, N7937);
nor NOR2 (N23447, N23425, N3579);
nand NAND3 (N23448, N23446, N8934, N15421);
nand NAND3 (N23449, N23447, N15295, N17529);
or OR3 (N23450, N23424, N6251, N12109);
not NOT1 (N23451, N23437);
not NOT1 (N23452, N23449);
xor XOR2 (N23453, N23450, N14305);
or OR4 (N23454, N23433, N16121, N15194, N556);
or OR3 (N23455, N23453, N5364, N21474);
xor XOR2 (N23456, N23445, N3104);
buf BUF1 (N23457, N23455);
not NOT1 (N23458, N23441);
buf BUF1 (N23459, N23456);
xor XOR2 (N23460, N23452, N12394);
xor XOR2 (N23461, N23457, N21232);
xor XOR2 (N23462, N23444, N18662);
or OR3 (N23463, N23462, N15856, N22335);
buf BUF1 (N23464, N23458);
buf BUF1 (N23465, N23463);
xor XOR2 (N23466, N23454, N15659);
buf BUF1 (N23467, N23436);
xor XOR2 (N23468, N23459, N1623);
nand NAND3 (N23469, N23468, N15177, N2819);
xor XOR2 (N23470, N23461, N20599);
nor NOR3 (N23471, N23448, N14602, N9630);
nor NOR2 (N23472, N23464, N5991);
not NOT1 (N23473, N23465);
and AND4 (N23474, N23451, N22194, N17949, N5946);
nand NAND3 (N23475, N23442, N3797, N4916);
nand NAND2 (N23476, N23469, N6109);
or OR4 (N23477, N23467, N6785, N7033, N14383);
buf BUF1 (N23478, N23472);
and AND3 (N23479, N23460, N12637, N2128);
or OR2 (N23480, N23477, N18662);
and AND4 (N23481, N23466, N7020, N5111, N21672);
and AND3 (N23482, N23474, N22035, N11088);
nor NOR2 (N23483, N23478, N8931);
nor NOR3 (N23484, N23479, N5286, N20156);
buf BUF1 (N23485, N23470);
nand NAND4 (N23486, N23473, N21393, N11566, N11076);
nor NOR2 (N23487, N23485, N9720);
nor NOR4 (N23488, N23482, N18072, N4533, N2271);
or OR3 (N23489, N23483, N23073, N2470);
not NOT1 (N23490, N23487);
and AND4 (N23491, N23489, N13228, N15220, N5471);
nand NAND4 (N23492, N23486, N17351, N3688, N18374);
or OR3 (N23493, N23476, N16329, N12466);
not NOT1 (N23494, N23480);
or OR2 (N23495, N23491, N1969);
not NOT1 (N23496, N23490);
and AND3 (N23497, N23496, N14483, N9907);
and AND3 (N23498, N23493, N14826, N21697);
nor NOR3 (N23499, N23492, N20329, N13111);
and AND3 (N23500, N23494, N14982, N8015);
buf BUF1 (N23501, N23500);
nand NAND3 (N23502, N23475, N10673, N18306);
buf BUF1 (N23503, N23481);
not NOT1 (N23504, N23495);
xor XOR2 (N23505, N23484, N1485);
xor XOR2 (N23506, N23503, N4959);
nand NAND4 (N23507, N23506, N19990, N171, N1031);
and AND4 (N23508, N23505, N10831, N14919, N19316);
buf BUF1 (N23509, N23471);
not NOT1 (N23510, N23498);
or OR2 (N23511, N23510, N1340);
xor XOR2 (N23512, N23497, N12310);
buf BUF1 (N23513, N23509);
nand NAND4 (N23514, N23513, N10233, N8766, N6182);
and AND3 (N23515, N23514, N7321, N16329);
xor XOR2 (N23516, N23511, N2275);
not NOT1 (N23517, N23508);
nor NOR4 (N23518, N23501, N4397, N6690, N21473);
nor NOR2 (N23519, N23515, N14);
xor XOR2 (N23520, N23499, N5582);
nand NAND4 (N23521, N23519, N11551, N2697, N20289);
nand NAND2 (N23522, N23518, N18324);
buf BUF1 (N23523, N23516);
xor XOR2 (N23524, N23517, N5702);
or OR4 (N23525, N23504, N7724, N21059, N5581);
or OR3 (N23526, N23525, N3263, N22683);
nand NAND3 (N23527, N23507, N11697, N6062);
nand NAND4 (N23528, N23520, N570, N11198, N8702);
xor XOR2 (N23529, N23522, N20978);
or OR2 (N23530, N23488, N19730);
and AND2 (N23531, N23502, N4746);
buf BUF1 (N23532, N23512);
not NOT1 (N23533, N23524);
xor XOR2 (N23534, N23526, N10215);
or OR2 (N23535, N23530, N23265);
nand NAND2 (N23536, N23533, N2268);
and AND3 (N23537, N23529, N6993, N14917);
xor XOR2 (N23538, N23535, N3623);
or OR3 (N23539, N23531, N23018, N3157);
and AND4 (N23540, N23523, N3195, N19359, N23060);
buf BUF1 (N23541, N23537);
nand NAND4 (N23542, N23539, N3442, N14042, N9518);
nor NOR3 (N23543, N23527, N284, N2710);
xor XOR2 (N23544, N23528, N22904);
not NOT1 (N23545, N23521);
nor NOR2 (N23546, N23538, N16073);
buf BUF1 (N23547, N23542);
not NOT1 (N23548, N23536);
and AND2 (N23549, N23532, N12334);
buf BUF1 (N23550, N23540);
or OR4 (N23551, N23547, N157, N21238, N15446);
not NOT1 (N23552, N23543);
not NOT1 (N23553, N23550);
buf BUF1 (N23554, N23548);
nor NOR2 (N23555, N23541, N16722);
nor NOR2 (N23556, N23552, N12098);
and AND3 (N23557, N23556, N8972, N23308);
buf BUF1 (N23558, N23557);
and AND3 (N23559, N23534, N6852, N21753);
or OR2 (N23560, N23555, N8308);
xor XOR2 (N23561, N23544, N12348);
buf BUF1 (N23562, N23561);
buf BUF1 (N23563, N23562);
buf BUF1 (N23564, N23553);
buf BUF1 (N23565, N23563);
and AND3 (N23566, N23560, N6451, N21265);
buf BUF1 (N23567, N23549);
nand NAND2 (N23568, N23546, N18697);
or OR4 (N23569, N23554, N23177, N3552, N10492);
xor XOR2 (N23570, N23567, N17884);
or OR4 (N23571, N23545, N12978, N19362, N13718);
buf BUF1 (N23572, N23568);
not NOT1 (N23573, N23565);
and AND3 (N23574, N23558, N18759, N23158);
buf BUF1 (N23575, N23551);
nor NOR3 (N23576, N23571, N21112, N6825);
xor XOR2 (N23577, N23575, N7735);
nand NAND2 (N23578, N23569, N9622);
xor XOR2 (N23579, N23577, N19397);
nand NAND2 (N23580, N23572, N10732);
not NOT1 (N23581, N23559);
not NOT1 (N23582, N23566);
nand NAND2 (N23583, N23576, N17376);
nor NOR2 (N23584, N23574, N15826);
nor NOR4 (N23585, N23573, N14692, N15754, N3233);
or OR2 (N23586, N23585, N4802);
or OR3 (N23587, N23586, N17423, N23183);
buf BUF1 (N23588, N23570);
xor XOR2 (N23589, N23581, N687);
nor NOR3 (N23590, N23587, N11642, N2646);
buf BUF1 (N23591, N23583);
nand NAND3 (N23592, N23579, N14909, N12190);
nand NAND4 (N23593, N23584, N13740, N20406, N5693);
nand NAND4 (N23594, N23591, N14476, N937, N18348);
nor NOR4 (N23595, N23582, N11234, N18848, N9299);
xor XOR2 (N23596, N23590, N23563);
and AND4 (N23597, N23594, N12338, N23176, N15988);
xor XOR2 (N23598, N23564, N4926);
not NOT1 (N23599, N23589);
or OR4 (N23600, N23592, N22248, N22604, N17846);
buf BUF1 (N23601, N23580);
not NOT1 (N23602, N23588);
nor NOR2 (N23603, N23578, N1526);
nand NAND4 (N23604, N23602, N6266, N17500, N4197);
nor NOR3 (N23605, N23593, N11563, N4444);
buf BUF1 (N23606, N23599);
and AND3 (N23607, N23598, N4549, N5168);
not NOT1 (N23608, N23600);
buf BUF1 (N23609, N23595);
nor NOR3 (N23610, N23606, N16847, N10855);
nor NOR4 (N23611, N23601, N7814, N15305, N18208);
xor XOR2 (N23612, N23609, N23041);
and AND2 (N23613, N23597, N22670);
buf BUF1 (N23614, N23596);
nor NOR2 (N23615, N23613, N14459);
nand NAND3 (N23616, N23614, N1055, N8078);
nor NOR3 (N23617, N23604, N14113, N2087);
and AND3 (N23618, N23615, N16666, N22420);
not NOT1 (N23619, N23605);
or OR2 (N23620, N23618, N20733);
or OR2 (N23621, N23617, N5230);
not NOT1 (N23622, N23608);
buf BUF1 (N23623, N23622);
nor NOR2 (N23624, N23619, N4239);
not NOT1 (N23625, N23624);
not NOT1 (N23626, N23612);
buf BUF1 (N23627, N23616);
not NOT1 (N23628, N23603);
xor XOR2 (N23629, N23626, N10150);
or OR3 (N23630, N23625, N19283, N9575);
nor NOR2 (N23631, N23620, N7418);
and AND3 (N23632, N23630, N8429, N15061);
and AND3 (N23633, N23629, N4525, N17919);
or OR2 (N23634, N23623, N3750);
not NOT1 (N23635, N23632);
and AND4 (N23636, N23610, N12300, N6886, N10922);
xor XOR2 (N23637, N23627, N22952);
or OR3 (N23638, N23633, N17820, N23462);
and AND2 (N23639, N23634, N3306);
not NOT1 (N23640, N23607);
xor XOR2 (N23641, N23631, N11222);
buf BUF1 (N23642, N23635);
not NOT1 (N23643, N23639);
not NOT1 (N23644, N23642);
nor NOR2 (N23645, N23621, N22568);
and AND4 (N23646, N23636, N4263, N23029, N21797);
buf BUF1 (N23647, N23644);
or OR3 (N23648, N23640, N21803, N10069);
or OR2 (N23649, N23643, N18184);
nor NOR4 (N23650, N23641, N20468, N4501, N724);
xor XOR2 (N23651, N23648, N17196);
not NOT1 (N23652, N23638);
nand NAND4 (N23653, N23628, N5333, N1308, N16880);
and AND4 (N23654, N23647, N741, N2758, N22197);
and AND2 (N23655, N23611, N8497);
or OR4 (N23656, N23637, N17815, N23356, N5839);
nand NAND4 (N23657, N23652, N9786, N4009, N20794);
nand NAND4 (N23658, N23646, N13469, N12637, N22160);
buf BUF1 (N23659, N23655);
nand NAND4 (N23660, N23653, N19615, N23148, N248);
or OR4 (N23661, N23657, N2026, N10028, N17617);
and AND4 (N23662, N23650, N16725, N19882, N14339);
buf BUF1 (N23663, N23660);
and AND2 (N23664, N23663, N18423);
and AND2 (N23665, N23649, N14393);
nand NAND2 (N23666, N23661, N9866);
not NOT1 (N23667, N23664);
not NOT1 (N23668, N23662);
or OR2 (N23669, N23667, N21333);
nor NOR2 (N23670, N23651, N12587);
xor XOR2 (N23671, N23656, N18443);
or OR2 (N23672, N23654, N5256);
not NOT1 (N23673, N23659);
nand NAND4 (N23674, N23671, N18293, N2407, N8066);
or OR2 (N23675, N23658, N4162);
not NOT1 (N23676, N23674);
xor XOR2 (N23677, N23676, N16418);
xor XOR2 (N23678, N23677, N8120);
not NOT1 (N23679, N23669);
and AND4 (N23680, N23675, N21621, N10902, N12150);
and AND3 (N23681, N23672, N11548, N3862);
and AND4 (N23682, N23678, N11553, N13547, N834);
nor NOR2 (N23683, N23666, N3511);
xor XOR2 (N23684, N23645, N23528);
or OR2 (N23685, N23683, N18515);
or OR4 (N23686, N23665, N3560, N11638, N13562);
not NOT1 (N23687, N23685);
not NOT1 (N23688, N23684);
or OR3 (N23689, N23668, N13440, N21119);
buf BUF1 (N23690, N23681);
buf BUF1 (N23691, N23679);
not NOT1 (N23692, N23680);
buf BUF1 (N23693, N23692);
and AND4 (N23694, N23673, N6468, N3477, N2812);
buf BUF1 (N23695, N23686);
and AND2 (N23696, N23682, N14434);
nor NOR3 (N23697, N23689, N1255, N16391);
xor XOR2 (N23698, N23691, N271);
or OR3 (N23699, N23698, N9938, N5322);
or OR4 (N23700, N23688, N1998, N4728, N17177);
not NOT1 (N23701, N23699);
buf BUF1 (N23702, N23693);
nand NAND3 (N23703, N23702, N14821, N3711);
not NOT1 (N23704, N23696);
or OR4 (N23705, N23670, N15447, N18241, N19499);
nor NOR3 (N23706, N23687, N15280, N22260);
xor XOR2 (N23707, N23701, N3398);
and AND3 (N23708, N23703, N23706, N11043);
or OR3 (N23709, N11060, N16772, N22383);
nand NAND3 (N23710, N23695, N6455, N14709);
buf BUF1 (N23711, N23708);
xor XOR2 (N23712, N23707, N10867);
xor XOR2 (N23713, N23710, N6177);
xor XOR2 (N23714, N23712, N984);
or OR2 (N23715, N23711, N16491);
or OR2 (N23716, N23713, N4968);
nor NOR4 (N23717, N23694, N21325, N23325, N22053);
not NOT1 (N23718, N23714);
xor XOR2 (N23719, N23704, N2266);
and AND3 (N23720, N23717, N23299, N8720);
xor XOR2 (N23721, N23720, N789);
xor XOR2 (N23722, N23709, N22701);
buf BUF1 (N23723, N23722);
not NOT1 (N23724, N23721);
and AND4 (N23725, N23700, N12457, N231, N22142);
not NOT1 (N23726, N23705);
not NOT1 (N23727, N23697);
xor XOR2 (N23728, N23726, N13626);
or OR2 (N23729, N23716, N22762);
xor XOR2 (N23730, N23724, N20808);
and AND2 (N23731, N23725, N23657);
and AND4 (N23732, N23719, N4894, N19770, N11673);
nor NOR3 (N23733, N23729, N16565, N531);
buf BUF1 (N23734, N23723);
nor NOR2 (N23735, N23715, N20949);
buf BUF1 (N23736, N23731);
buf BUF1 (N23737, N23727);
nor NOR2 (N23738, N23718, N13100);
and AND3 (N23739, N23737, N15225, N19083);
nor NOR2 (N23740, N23730, N20867);
nor NOR3 (N23741, N23728, N3789, N11897);
nor NOR4 (N23742, N23690, N6162, N20853, N20114);
nand NAND3 (N23743, N23735, N15331, N9833);
and AND3 (N23744, N23736, N618, N1771);
or OR3 (N23745, N23734, N3251, N23574);
buf BUF1 (N23746, N23732);
xor XOR2 (N23747, N23745, N23470);
not NOT1 (N23748, N23744);
not NOT1 (N23749, N23741);
nand NAND4 (N23750, N23739, N6241, N2103, N13995);
buf BUF1 (N23751, N23748);
buf BUF1 (N23752, N23749);
nor NOR3 (N23753, N23751, N22209, N19253);
and AND2 (N23754, N23753, N19501);
not NOT1 (N23755, N23743);
and AND2 (N23756, N23747, N12274);
nor NOR4 (N23757, N23742, N23744, N19379, N1122);
buf BUF1 (N23758, N23757);
and AND3 (N23759, N23738, N9908, N9178);
or OR3 (N23760, N23740, N14609, N6584);
not NOT1 (N23761, N23756);
buf BUF1 (N23762, N23733);
not NOT1 (N23763, N23746);
xor XOR2 (N23764, N23760, N22605);
nand NAND3 (N23765, N23755, N9410, N22578);
buf BUF1 (N23766, N23763);
or OR3 (N23767, N23759, N19269, N9579);
buf BUF1 (N23768, N23764);
xor XOR2 (N23769, N23750, N8333);
xor XOR2 (N23770, N23752, N13872);
not NOT1 (N23771, N23754);
or OR3 (N23772, N23771, N5439, N1502);
nor NOR2 (N23773, N23758, N23694);
xor XOR2 (N23774, N23773, N15462);
nor NOR4 (N23775, N23770, N11412, N11614, N16635);
or OR4 (N23776, N23766, N4973, N14127, N22260);
buf BUF1 (N23777, N23768);
xor XOR2 (N23778, N23762, N16098);
nor NOR4 (N23779, N23772, N17477, N1712, N13332);
xor XOR2 (N23780, N23769, N1902);
nand NAND4 (N23781, N23767, N12381, N16522, N9838);
and AND4 (N23782, N23761, N7615, N12798, N1560);
or OR2 (N23783, N23781, N1658);
not NOT1 (N23784, N23765);
buf BUF1 (N23785, N23777);
xor XOR2 (N23786, N23775, N475);
and AND3 (N23787, N23784, N4713, N18348);
xor XOR2 (N23788, N23778, N12576);
buf BUF1 (N23789, N23774);
not NOT1 (N23790, N23776);
nor NOR4 (N23791, N23790, N10193, N8168, N13569);
nand NAND4 (N23792, N23783, N5664, N15286, N10001);
and AND3 (N23793, N23787, N17787, N21492);
and AND2 (N23794, N23786, N6271);
and AND2 (N23795, N23793, N23463);
not NOT1 (N23796, N23794);
nand NAND4 (N23797, N23789, N8156, N18246, N16820);
not NOT1 (N23798, N23779);
xor XOR2 (N23799, N23792, N15916);
and AND4 (N23800, N23782, N17975, N17500, N14425);
nand NAND2 (N23801, N23798, N4947);
or OR3 (N23802, N23788, N5677, N17763);
and AND3 (N23803, N23780, N20303, N17731);
buf BUF1 (N23804, N23785);
and AND2 (N23805, N23796, N22110);
or OR4 (N23806, N23802, N9668, N2828, N6166);
and AND2 (N23807, N23804, N23798);
or OR3 (N23808, N23797, N1952, N1373);
nor NOR2 (N23809, N23800, N9421);
nor NOR2 (N23810, N23803, N20324);
not NOT1 (N23811, N23808);
or OR4 (N23812, N23805, N8180, N23451, N144);
not NOT1 (N23813, N23807);
nand NAND3 (N23814, N23795, N820, N18436);
xor XOR2 (N23815, N23810, N23390);
and AND4 (N23816, N23811, N18963, N4113, N3056);
buf BUF1 (N23817, N23813);
buf BUF1 (N23818, N23806);
buf BUF1 (N23819, N23817);
not NOT1 (N23820, N23815);
or OR3 (N23821, N23814, N21542, N274);
or OR4 (N23822, N23816, N12223, N799, N14902);
or OR4 (N23823, N23812, N21332, N550, N22182);
nor NOR3 (N23824, N23791, N19012, N18763);
nor NOR2 (N23825, N23809, N2818);
nor NOR4 (N23826, N23823, N17564, N10904, N3705);
or OR4 (N23827, N23801, N8362, N14189, N7315);
and AND4 (N23828, N23818, N915, N21526, N20898);
xor XOR2 (N23829, N23820, N18000);
nand NAND2 (N23830, N23829, N5015);
not NOT1 (N23831, N23799);
buf BUF1 (N23832, N23819);
not NOT1 (N23833, N23825);
xor XOR2 (N23834, N23826, N19618);
and AND2 (N23835, N23834, N3754);
or OR2 (N23836, N23828, N21820);
nor NOR4 (N23837, N23830, N22471, N21271, N10418);
xor XOR2 (N23838, N23822, N18573);
nor NOR3 (N23839, N23836, N11309, N21962);
nor NOR2 (N23840, N23839, N16318);
or OR2 (N23841, N23821, N7138);
xor XOR2 (N23842, N23824, N13461);
nor NOR2 (N23843, N23831, N6551);
buf BUF1 (N23844, N23842);
buf BUF1 (N23845, N23838);
nor NOR4 (N23846, N23832, N10139, N9509, N5734);
and AND2 (N23847, N23845, N14585);
nor NOR2 (N23848, N23840, N3948);
not NOT1 (N23849, N23843);
and AND2 (N23850, N23827, N7750);
not NOT1 (N23851, N23847);
and AND4 (N23852, N23837, N527, N10512, N16258);
or OR4 (N23853, N23848, N22587, N2637, N5095);
and AND2 (N23854, N23850, N10913);
nor NOR3 (N23855, N23849, N23561, N4373);
not NOT1 (N23856, N23853);
buf BUF1 (N23857, N23856);
or OR2 (N23858, N23835, N9840);
or OR3 (N23859, N23833, N23445, N7505);
buf BUF1 (N23860, N23841);
nand NAND2 (N23861, N23852, N12255);
nor NOR3 (N23862, N23844, N12391, N23406);
nor NOR4 (N23863, N23861, N6973, N5436, N3164);
xor XOR2 (N23864, N23863, N8356);
or OR4 (N23865, N23857, N18895, N6434, N18577);
and AND4 (N23866, N23859, N3858, N21468, N22511);
nor NOR3 (N23867, N23866, N21699, N9016);
and AND3 (N23868, N23865, N4638, N18318);
buf BUF1 (N23869, N23867);
xor XOR2 (N23870, N23860, N6530);
nand NAND2 (N23871, N23851, N14500);
or OR4 (N23872, N23846, N691, N1378, N8911);
buf BUF1 (N23873, N23862);
xor XOR2 (N23874, N23858, N20411);
or OR2 (N23875, N23873, N19410);
nor NOR2 (N23876, N23855, N13803);
nand NAND4 (N23877, N23872, N9416, N1039, N10867);
or OR3 (N23878, N23869, N12691, N2146);
nand NAND4 (N23879, N23876, N15193, N7241, N10811);
nand NAND3 (N23880, N23875, N22068, N19939);
or OR3 (N23881, N23877, N15037, N7379);
buf BUF1 (N23882, N23879);
not NOT1 (N23883, N23881);
nor NOR2 (N23884, N23868, N4767);
and AND2 (N23885, N23880, N16646);
not NOT1 (N23886, N23854);
and AND3 (N23887, N23878, N13657, N20000);
xor XOR2 (N23888, N23871, N20759);
nor NOR3 (N23889, N23888, N12905, N18895);
or OR2 (N23890, N23887, N17042);
nand NAND2 (N23891, N23884, N2501);
xor XOR2 (N23892, N23890, N2526);
not NOT1 (N23893, N23864);
nand NAND2 (N23894, N23889, N7819);
and AND4 (N23895, N23882, N556, N21807, N20216);
and AND3 (N23896, N23885, N496, N8536);
and AND3 (N23897, N23896, N12001, N17052);
or OR3 (N23898, N23893, N15669, N6826);
not NOT1 (N23899, N23883);
xor XOR2 (N23900, N23870, N9385);
buf BUF1 (N23901, N23874);
and AND4 (N23902, N23897, N14114, N11591, N18903);
and AND3 (N23903, N23902, N19833, N15680);
or OR2 (N23904, N23903, N2615);
not NOT1 (N23905, N23904);
nand NAND4 (N23906, N23901, N12744, N887, N22519);
nor NOR3 (N23907, N23900, N11977, N13183);
not NOT1 (N23908, N23886);
and AND2 (N23909, N23898, N15529);
xor XOR2 (N23910, N23906, N16907);
and AND4 (N23911, N23891, N7022, N2564, N8302);
or OR2 (N23912, N23909, N14801);
and AND3 (N23913, N23907, N14358, N1989);
not NOT1 (N23914, N23912);
nand NAND4 (N23915, N23908, N17822, N21410, N22626);
and AND4 (N23916, N23911, N13366, N12623, N9115);
or OR4 (N23917, N23899, N2670, N9597, N18784);
buf BUF1 (N23918, N23913);
nand NAND3 (N23919, N23914, N17254, N3272);
or OR3 (N23920, N23919, N20117, N20011);
buf BUF1 (N23921, N23892);
or OR3 (N23922, N23920, N22055, N11794);
nor NOR2 (N23923, N23905, N14757);
buf BUF1 (N23924, N23916);
and AND4 (N23925, N23923, N12459, N9713, N7952);
not NOT1 (N23926, N23894);
nor NOR4 (N23927, N23926, N7651, N6594, N17037);
nor NOR2 (N23928, N23921, N2692);
not NOT1 (N23929, N23924);
buf BUF1 (N23930, N23917);
nor NOR4 (N23931, N23895, N499, N14368, N20295);
buf BUF1 (N23932, N23930);
xor XOR2 (N23933, N23928, N6800);
nor NOR4 (N23934, N23929, N10087, N20559, N12558);
and AND3 (N23935, N23915, N4014, N20237);
buf BUF1 (N23936, N23918);
and AND3 (N23937, N23922, N7288, N17345);
not NOT1 (N23938, N23936);
buf BUF1 (N23939, N23934);
xor XOR2 (N23940, N23927, N5027);
or OR2 (N23941, N23933, N5779);
not NOT1 (N23942, N23931);
and AND2 (N23943, N23925, N21790);
and AND2 (N23944, N23938, N15994);
or OR3 (N23945, N23932, N18463, N1816);
xor XOR2 (N23946, N23943, N14684);
or OR4 (N23947, N23939, N4118, N4159, N9044);
xor XOR2 (N23948, N23942, N22052);
xor XOR2 (N23949, N23945, N14071);
or OR4 (N23950, N23941, N20488, N23937, N8873);
or OR4 (N23951, N561, N22022, N10174, N11628);
xor XOR2 (N23952, N23951, N2578);
and AND2 (N23953, N23948, N11178);
and AND2 (N23954, N23949, N10320);
buf BUF1 (N23955, N23910);
or OR3 (N23956, N23944, N22571, N21726);
not NOT1 (N23957, N23954);
nor NOR2 (N23958, N23953, N7900);
not NOT1 (N23959, N23935);
or OR4 (N23960, N23958, N15749, N1094, N7060);
nor NOR4 (N23961, N23959, N8403, N3510, N12892);
buf BUF1 (N23962, N23957);
not NOT1 (N23963, N23956);
or OR2 (N23964, N23960, N8639);
and AND4 (N23965, N23955, N7764, N22857, N22463);
xor XOR2 (N23966, N23962, N19894);
buf BUF1 (N23967, N23963);
buf BUF1 (N23968, N23965);
nor NOR2 (N23969, N23966, N16544);
nand NAND2 (N23970, N23952, N20172);
nand NAND3 (N23971, N23940, N19133, N7108);
or OR3 (N23972, N23967, N17905, N2960);
or OR4 (N23973, N23964, N13103, N11869, N12212);
nand NAND4 (N23974, N23946, N12632, N4141, N2491);
buf BUF1 (N23975, N23950);
xor XOR2 (N23976, N23974, N9825);
or OR3 (N23977, N23947, N12056, N12458);
xor XOR2 (N23978, N23971, N16855);
nor NOR4 (N23979, N23976, N16617, N22237, N11538);
not NOT1 (N23980, N23972);
nor NOR2 (N23981, N23979, N19923);
nor NOR3 (N23982, N23973, N12780, N17176);
xor XOR2 (N23983, N23969, N7236);
xor XOR2 (N23984, N23978, N20013);
or OR4 (N23985, N23977, N20244, N13263, N12594);
and AND4 (N23986, N23975, N5939, N1838, N22288);
and AND2 (N23987, N23981, N15419);
xor XOR2 (N23988, N23987, N7246);
nor NOR4 (N23989, N23970, N6282, N22191, N12236);
nor NOR2 (N23990, N23988, N372);
and AND2 (N23991, N23986, N19923);
and AND4 (N23992, N23980, N7089, N3640, N8445);
buf BUF1 (N23993, N23990);
buf BUF1 (N23994, N23968);
nor NOR3 (N23995, N23994, N8936, N17594);
not NOT1 (N23996, N23993);
not NOT1 (N23997, N23991);
not NOT1 (N23998, N23961);
nor NOR4 (N23999, N23982, N10494, N8268, N14646);
not NOT1 (N24000, N23999);
and AND4 (N24001, N23995, N1382, N19806, N16886);
not NOT1 (N24002, N23997);
xor XOR2 (N24003, N23998, N13842);
or OR4 (N24004, N23983, N10931, N22462, N8786);
or OR3 (N24005, N24004, N23352, N2636);
and AND3 (N24006, N23984, N22894, N8385);
or OR4 (N24007, N23996, N22330, N17868, N9718);
or OR2 (N24008, N24007, N915);
nand NAND4 (N24009, N24008, N2813, N552, N8787);
and AND4 (N24010, N24000, N5984, N22266, N11407);
xor XOR2 (N24011, N24002, N20766);
and AND2 (N24012, N24003, N10428);
buf BUF1 (N24013, N23985);
not NOT1 (N24014, N24013);
and AND2 (N24015, N24014, N20888);
and AND2 (N24016, N23992, N11162);
and AND4 (N24017, N24006, N1607, N16735, N3899);
nand NAND3 (N24018, N24001, N10990, N21160);
or OR3 (N24019, N24015, N5289, N18422);
and AND2 (N24020, N24019, N10708);
nand NAND4 (N24021, N24010, N23244, N2936, N18029);
nand NAND4 (N24022, N24005, N9014, N3814, N18831);
not NOT1 (N24023, N24011);
nor NOR4 (N24024, N24020, N7843, N2434, N10332);
or OR2 (N24025, N24012, N1154);
nand NAND3 (N24026, N24023, N20180, N557);
buf BUF1 (N24027, N23989);
buf BUF1 (N24028, N24024);
not NOT1 (N24029, N24027);
and AND3 (N24030, N24016, N12805, N21365);
or OR4 (N24031, N24009, N5061, N15321, N19741);
not NOT1 (N24032, N24031);
or OR3 (N24033, N24030, N883, N14745);
buf BUF1 (N24034, N24018);
nor NOR4 (N24035, N24021, N24021, N17749, N12667);
nand NAND4 (N24036, N24034, N13440, N20697, N10051);
nand NAND2 (N24037, N24036, N5134);
nor NOR3 (N24038, N24029, N10993, N11852);
xor XOR2 (N24039, N24032, N10504);
nand NAND2 (N24040, N24028, N22560);
or OR3 (N24041, N24017, N6047, N14034);
nand NAND3 (N24042, N24037, N3292, N3381);
xor XOR2 (N24043, N24026, N48);
or OR2 (N24044, N24042, N1975);
nand NAND2 (N24045, N24035, N14950);
nand NAND3 (N24046, N24033, N11513, N23489);
nor NOR2 (N24047, N24044, N22656);
xor XOR2 (N24048, N24038, N16965);
not NOT1 (N24049, N24040);
and AND2 (N24050, N24047, N4802);
and AND4 (N24051, N24025, N17169, N9066, N14469);
and AND3 (N24052, N24049, N13878, N13893);
and AND4 (N24053, N24041, N23802, N23454, N11405);
xor XOR2 (N24054, N24048, N3537);
nand NAND3 (N24055, N24039, N13120, N17823);
buf BUF1 (N24056, N24022);
nor NOR4 (N24057, N24053, N20773, N21264, N23849);
xor XOR2 (N24058, N24056, N22895);
xor XOR2 (N24059, N24058, N1524);
and AND4 (N24060, N24050, N9530, N579, N3616);
and AND2 (N24061, N24045, N10856);
buf BUF1 (N24062, N24060);
xor XOR2 (N24063, N24043, N6926);
not NOT1 (N24064, N24061);
nand NAND3 (N24065, N24062, N3467, N669);
buf BUF1 (N24066, N24065);
not NOT1 (N24067, N24046);
nand NAND3 (N24068, N24055, N19304, N10071);
xor XOR2 (N24069, N24064, N10543);
xor XOR2 (N24070, N24063, N3206);
not NOT1 (N24071, N24066);
not NOT1 (N24072, N24057);
not NOT1 (N24073, N24067);
xor XOR2 (N24074, N24071, N20080);
buf BUF1 (N24075, N24059);
not NOT1 (N24076, N24074);
and AND3 (N24077, N24070, N15027, N14108);
not NOT1 (N24078, N24068);
xor XOR2 (N24079, N24072, N22215);
xor XOR2 (N24080, N24052, N13950);
or OR4 (N24081, N24077, N1981, N578, N5022);
not NOT1 (N24082, N24081);
or OR2 (N24083, N24075, N16545);
nand NAND4 (N24084, N24069, N2327, N17658, N16308);
nand NAND2 (N24085, N24080, N609);
or OR3 (N24086, N24054, N16888, N9088);
or OR3 (N24087, N24085, N21437, N11751);
nand NAND2 (N24088, N24087, N17292);
buf BUF1 (N24089, N24079);
buf BUF1 (N24090, N24051);
or OR4 (N24091, N24090, N13864, N9156, N16774);
buf BUF1 (N24092, N24088);
or OR4 (N24093, N24073, N19750, N23247, N14354);
nor NOR2 (N24094, N24076, N13550);
or OR4 (N24095, N24092, N2756, N3049, N11599);
and AND3 (N24096, N24089, N5212, N94);
and AND4 (N24097, N24086, N7901, N8017, N5619);
or OR4 (N24098, N24095, N12017, N8667, N3978);
nor NOR2 (N24099, N24091, N10582);
buf BUF1 (N24100, N24097);
nor NOR2 (N24101, N24083, N10626);
and AND3 (N24102, N24094, N12592, N17194);
buf BUF1 (N24103, N24098);
xor XOR2 (N24104, N24078, N19404);
nand NAND2 (N24105, N24102, N5944);
or OR3 (N24106, N24084, N10605, N15722);
nand NAND4 (N24107, N24099, N170, N8763, N5452);
xor XOR2 (N24108, N24106, N14502);
nand NAND4 (N24109, N24107, N10765, N15401, N17199);
nand NAND4 (N24110, N24104, N14682, N3675, N21648);
not NOT1 (N24111, N24082);
and AND3 (N24112, N24093, N23770, N2877);
xor XOR2 (N24113, N24101, N6021);
xor XOR2 (N24114, N24113, N18268);
nand NAND3 (N24115, N24096, N3668, N11289);
and AND2 (N24116, N24100, N5065);
buf BUF1 (N24117, N24116);
and AND2 (N24118, N24103, N14088);
and AND2 (N24119, N24108, N16407);
not NOT1 (N24120, N24105);
buf BUF1 (N24121, N24115);
not NOT1 (N24122, N24119);
nor NOR4 (N24123, N24120, N2014, N16171, N5898);
and AND4 (N24124, N24110, N8882, N1626, N9748);
and AND4 (N24125, N24121, N17687, N9485, N1398);
or OR2 (N24126, N24112, N12945);
xor XOR2 (N24127, N24117, N20273);
not NOT1 (N24128, N24127);
and AND3 (N24129, N24128, N14687, N8602);
nor NOR3 (N24130, N24114, N22064, N18769);
nand NAND3 (N24131, N24130, N2011, N9218);
nand NAND3 (N24132, N24111, N17101, N22151);
and AND3 (N24133, N24122, N3137, N112);
nand NAND2 (N24134, N24118, N11920);
nand NAND3 (N24135, N24131, N9808, N20843);
nor NOR3 (N24136, N24125, N4899, N5588);
or OR4 (N24137, N24129, N628, N12816, N306);
and AND3 (N24138, N24137, N22467, N12520);
not NOT1 (N24139, N24138);
xor XOR2 (N24140, N24136, N3760);
buf BUF1 (N24141, N24123);
nand NAND4 (N24142, N24133, N11027, N9096, N4723);
not NOT1 (N24143, N24109);
nand NAND4 (N24144, N24142, N12885, N15225, N3378);
buf BUF1 (N24145, N24126);
nor NOR4 (N24146, N24139, N12391, N1056, N14711);
and AND2 (N24147, N24144, N21639);
nand NAND2 (N24148, N24134, N23306);
not NOT1 (N24149, N24145);
buf BUF1 (N24150, N24148);
and AND2 (N24151, N24146, N20140);
and AND4 (N24152, N24143, N924, N22523, N16922);
xor XOR2 (N24153, N24140, N3979);
xor XOR2 (N24154, N24124, N9287);
xor XOR2 (N24155, N24149, N18124);
and AND3 (N24156, N24150, N2937, N12116);
not NOT1 (N24157, N24132);
and AND4 (N24158, N24157, N20581, N11508, N15077);
or OR3 (N24159, N24152, N3352, N20970);
xor XOR2 (N24160, N24135, N18795);
nor NOR2 (N24161, N24156, N11234);
not NOT1 (N24162, N24153);
buf BUF1 (N24163, N24162);
nand NAND3 (N24164, N24141, N10739, N6862);
or OR2 (N24165, N24164, N13446);
nand NAND4 (N24166, N24154, N3665, N3840, N10577);
nand NAND2 (N24167, N24147, N4654);
xor XOR2 (N24168, N24155, N1728);
or OR2 (N24169, N24166, N23652);
or OR4 (N24170, N24160, N21704, N14466, N15505);
nor NOR4 (N24171, N24158, N22947, N19725, N23988);
or OR4 (N24172, N24167, N13520, N1661, N11568);
buf BUF1 (N24173, N24165);
nor NOR4 (N24174, N24163, N12849, N14654, N18548);
nand NAND2 (N24175, N24168, N5608);
not NOT1 (N24176, N24174);
not NOT1 (N24177, N24176);
buf BUF1 (N24178, N24177);
and AND4 (N24179, N24169, N22100, N639, N15569);
xor XOR2 (N24180, N24161, N20361);
xor XOR2 (N24181, N24170, N16927);
buf BUF1 (N24182, N24171);
nor NOR4 (N24183, N24159, N18541, N18345, N22113);
nand NAND2 (N24184, N24175, N16326);
nor NOR4 (N24185, N24178, N13158, N7754, N11951);
not NOT1 (N24186, N24183);
or OR4 (N24187, N24180, N20483, N17646, N12432);
buf BUF1 (N24188, N24187);
and AND2 (N24189, N24181, N20724);
and AND4 (N24190, N24186, N22515, N7235, N17747);
nand NAND4 (N24191, N24190, N5682, N23841, N16423);
buf BUF1 (N24192, N24188);
xor XOR2 (N24193, N24184, N18977);
xor XOR2 (N24194, N24191, N18834);
nand NAND4 (N24195, N24192, N12986, N5952, N9017);
and AND3 (N24196, N24193, N254, N22489);
nand NAND3 (N24197, N24195, N4296, N5585);
nand NAND4 (N24198, N24196, N11878, N22536, N22419);
nor NOR2 (N24199, N24198, N12318);
not NOT1 (N24200, N24197);
xor XOR2 (N24201, N24182, N15599);
buf BUF1 (N24202, N24173);
xor XOR2 (N24203, N24201, N5794);
not NOT1 (N24204, N24189);
and AND4 (N24205, N24185, N23013, N9290, N14377);
and AND2 (N24206, N24151, N15179);
and AND2 (N24207, N24203, N6691);
nand NAND2 (N24208, N24199, N12540);
buf BUF1 (N24209, N24200);
xor XOR2 (N24210, N24205, N10954);
or OR4 (N24211, N24202, N22603, N10140, N16088);
xor XOR2 (N24212, N24194, N20335);
and AND2 (N24213, N24208, N17922);
not NOT1 (N24214, N24209);
or OR4 (N24215, N24206, N2433, N23874, N8408);
nor NOR4 (N24216, N24213, N13211, N7170, N13729);
not NOT1 (N24217, N24172);
not NOT1 (N24218, N24215);
buf BUF1 (N24219, N24214);
or OR2 (N24220, N24211, N23346);
not NOT1 (N24221, N24218);
and AND3 (N24222, N24221, N5887, N17942);
nand NAND3 (N24223, N24210, N7831, N3333);
xor XOR2 (N24224, N24217, N2333);
and AND2 (N24225, N24223, N18044);
nand NAND3 (N24226, N24207, N4652, N22536);
xor XOR2 (N24227, N24224, N12498);
xor XOR2 (N24228, N24204, N5235);
not NOT1 (N24229, N24222);
nand NAND2 (N24230, N24212, N1568);
xor XOR2 (N24231, N24220, N1653);
nor NOR4 (N24232, N24229, N10088, N5338, N19855);
nand NAND3 (N24233, N24179, N11854, N15652);
or OR3 (N24234, N24230, N12287, N9430);
not NOT1 (N24235, N24231);
xor XOR2 (N24236, N24216, N12545);
buf BUF1 (N24237, N24228);
buf BUF1 (N24238, N24232);
nor NOR2 (N24239, N24225, N598);
nor NOR3 (N24240, N24227, N9082, N19168);
nor NOR2 (N24241, N24226, N21954);
or OR3 (N24242, N24240, N5501, N12857);
nor NOR3 (N24243, N24237, N610, N22571);
nand NAND2 (N24244, N24233, N12817);
and AND4 (N24245, N24236, N14220, N20830, N22691);
nand NAND2 (N24246, N24219, N11209);
xor XOR2 (N24247, N24238, N7790);
or OR2 (N24248, N24235, N9239);
and AND2 (N24249, N24244, N8614);
nand NAND2 (N24250, N24246, N3402);
nor NOR2 (N24251, N24242, N22676);
and AND2 (N24252, N24250, N16113);
buf BUF1 (N24253, N24241);
and AND4 (N24254, N24248, N1637, N15228, N7187);
or OR3 (N24255, N24239, N10554, N12459);
buf BUF1 (N24256, N24234);
nand NAND3 (N24257, N24245, N20288, N10);
buf BUF1 (N24258, N24253);
xor XOR2 (N24259, N24258, N660);
xor XOR2 (N24260, N24251, N13252);
and AND4 (N24261, N24257, N701, N16295, N4177);
buf BUF1 (N24262, N24261);
or OR3 (N24263, N24247, N4490, N13625);
or OR2 (N24264, N24252, N4365);
nand NAND4 (N24265, N24263, N8022, N6542, N23728);
buf BUF1 (N24266, N24260);
xor XOR2 (N24267, N24264, N15771);
nand NAND4 (N24268, N24265, N3224, N4123, N6244);
buf BUF1 (N24269, N24262);
and AND3 (N24270, N24266, N21839, N484);
nand NAND4 (N24271, N24254, N378, N20320, N16072);
and AND4 (N24272, N24256, N20746, N18325, N24159);
not NOT1 (N24273, N24249);
xor XOR2 (N24274, N24267, N9036);
or OR2 (N24275, N24243, N18538);
or OR4 (N24276, N24269, N4421, N17144, N15926);
xor XOR2 (N24277, N24275, N1968);
nand NAND3 (N24278, N24259, N5801, N21946);
nor NOR3 (N24279, N24278, N570, N14407);
xor XOR2 (N24280, N24268, N24078);
and AND4 (N24281, N24279, N5863, N17205, N19540);
and AND2 (N24282, N24276, N19524);
nand NAND2 (N24283, N24277, N5135);
nand NAND2 (N24284, N24282, N20088);
or OR4 (N24285, N24255, N22089, N6501, N23850);
not NOT1 (N24286, N24281);
or OR2 (N24287, N24284, N15381);
buf BUF1 (N24288, N24270);
buf BUF1 (N24289, N24283);
xor XOR2 (N24290, N24287, N24227);
nand NAND2 (N24291, N24289, N7662);
not NOT1 (N24292, N24272);
and AND3 (N24293, N24271, N2625, N4706);
not NOT1 (N24294, N24280);
and AND3 (N24295, N24274, N19127, N7476);
nand NAND4 (N24296, N24293, N12041, N1454, N13200);
buf BUF1 (N24297, N24285);
buf BUF1 (N24298, N24290);
or OR3 (N24299, N24297, N9933, N972);
buf BUF1 (N24300, N24299);
and AND3 (N24301, N24296, N23660, N15504);
not NOT1 (N24302, N24301);
nand NAND4 (N24303, N24291, N12597, N23434, N9899);
or OR2 (N24304, N24303, N12379);
not NOT1 (N24305, N24298);
nor NOR3 (N24306, N24286, N11174, N7616);
not NOT1 (N24307, N24288);
buf BUF1 (N24308, N24295);
nor NOR4 (N24309, N24306, N17580, N2432, N18140);
nand NAND4 (N24310, N24307, N15571, N16609, N9951);
buf BUF1 (N24311, N24302);
xor XOR2 (N24312, N24308, N33);
or OR4 (N24313, N24294, N6330, N10934, N15413);
not NOT1 (N24314, N24305);
buf BUF1 (N24315, N24311);
xor XOR2 (N24316, N24309, N18423);
or OR2 (N24317, N24313, N13570);
and AND4 (N24318, N24316, N6275, N18862, N20780);
and AND4 (N24319, N24304, N4336, N15188, N22753);
nor NOR2 (N24320, N24310, N3944);
and AND4 (N24321, N24319, N18738, N6993, N19968);
xor XOR2 (N24322, N24320, N6821);
and AND3 (N24323, N24321, N10178, N499);
buf BUF1 (N24324, N24273);
nor NOR4 (N24325, N24315, N14165, N4424, N20279);
or OR4 (N24326, N24318, N14108, N22857, N10216);
buf BUF1 (N24327, N24324);
not NOT1 (N24328, N24300);
not NOT1 (N24329, N24292);
not NOT1 (N24330, N24317);
nor NOR3 (N24331, N24325, N12256, N21278);
and AND3 (N24332, N24330, N10432, N15501);
or OR3 (N24333, N24328, N18123, N8339);
nand NAND4 (N24334, N24314, N4486, N5702, N12492);
xor XOR2 (N24335, N24327, N11346);
not NOT1 (N24336, N24326);
buf BUF1 (N24337, N24334);
nand NAND4 (N24338, N24335, N11313, N17447, N16408);
not NOT1 (N24339, N24336);
or OR2 (N24340, N24333, N7279);
xor XOR2 (N24341, N24337, N7025);
not NOT1 (N24342, N24339);
nor NOR3 (N24343, N24312, N9147, N21709);
or OR4 (N24344, N24343, N12128, N3594, N10870);
nor NOR2 (N24345, N24323, N18604);
not NOT1 (N24346, N24345);
xor XOR2 (N24347, N24342, N18552);
nand NAND3 (N24348, N24341, N4813, N18026);
nor NOR2 (N24349, N24340, N23514);
not NOT1 (N24350, N24322);
not NOT1 (N24351, N24348);
buf BUF1 (N24352, N24346);
not NOT1 (N24353, N24347);
buf BUF1 (N24354, N24331);
buf BUF1 (N24355, N24349);
and AND2 (N24356, N24338, N19084);
nand NAND4 (N24357, N24350, N15192, N8441, N15093);
buf BUF1 (N24358, N24356);
xor XOR2 (N24359, N24354, N21999);
not NOT1 (N24360, N24355);
not NOT1 (N24361, N24332);
nand NAND4 (N24362, N24352, N14145, N3045, N12825);
not NOT1 (N24363, N24353);
not NOT1 (N24364, N24361);
nor NOR2 (N24365, N24357, N6550);
and AND3 (N24366, N24351, N19222, N3651);
not NOT1 (N24367, N24359);
nor NOR3 (N24368, N24329, N13136, N19703);
or OR2 (N24369, N24366, N14024);
buf BUF1 (N24370, N24362);
buf BUF1 (N24371, N24360);
xor XOR2 (N24372, N24363, N22704);
nand NAND4 (N24373, N24372, N8573, N22342, N16209);
not NOT1 (N24374, N24364);
xor XOR2 (N24375, N24365, N18923);
xor XOR2 (N24376, N24368, N18301);
nor NOR4 (N24377, N24376, N9997, N14667, N3938);
xor XOR2 (N24378, N24371, N24153);
and AND3 (N24379, N24344, N10015, N72);
xor XOR2 (N24380, N24369, N10280);
xor XOR2 (N24381, N24367, N2829);
buf BUF1 (N24382, N24377);
not NOT1 (N24383, N24370);
xor XOR2 (N24384, N24382, N8208);
and AND3 (N24385, N24379, N7196, N23154);
not NOT1 (N24386, N24383);
nor NOR2 (N24387, N24373, N1125);
nor NOR4 (N24388, N24385, N5806, N11958, N13538);
buf BUF1 (N24389, N24374);
xor XOR2 (N24390, N24387, N19401);
or OR3 (N24391, N24380, N11836, N11000);
nor NOR3 (N24392, N24391, N12590, N6823);
not NOT1 (N24393, N24378);
nand NAND2 (N24394, N24393, N21569);
nand NAND2 (N24395, N24389, N24121);
nor NOR3 (N24396, N24384, N4713, N181);
xor XOR2 (N24397, N24390, N4575);
nand NAND2 (N24398, N24358, N15936);
or OR3 (N24399, N24395, N2436, N13007);
nand NAND2 (N24400, N24375, N6017);
and AND3 (N24401, N24397, N11222, N6212);
nand NAND3 (N24402, N24400, N2877, N22264);
nand NAND2 (N24403, N24386, N20886);
buf BUF1 (N24404, N24399);
nor NOR4 (N24405, N24404, N16528, N4013, N11992);
xor XOR2 (N24406, N24398, N21772);
nand NAND3 (N24407, N24388, N5220, N11572);
xor XOR2 (N24408, N24392, N20865);
buf BUF1 (N24409, N24381);
buf BUF1 (N24410, N24408);
and AND3 (N24411, N24406, N21255, N19537);
and AND2 (N24412, N24410, N19566);
or OR3 (N24413, N24407, N24016, N7476);
buf BUF1 (N24414, N24405);
nor NOR3 (N24415, N24413, N24051, N15387);
nor NOR2 (N24416, N24401, N18841);
or OR3 (N24417, N24394, N1068, N9919);
or OR3 (N24418, N24409, N12490, N23388);
nor NOR3 (N24419, N24403, N4033, N994);
and AND2 (N24420, N24418, N7383);
nor NOR3 (N24421, N24420, N16773, N6157);
or OR3 (N24422, N24412, N20888, N15643);
and AND2 (N24423, N24396, N15056);
or OR2 (N24424, N24402, N10095);
nor NOR3 (N24425, N24419, N10646, N16220);
and AND2 (N24426, N24414, N19732);
nor NOR2 (N24427, N24411, N18933);
xor XOR2 (N24428, N24422, N6834);
or OR4 (N24429, N24417, N20427, N13204, N12936);
nor NOR3 (N24430, N24416, N19815, N14330);
nand NAND4 (N24431, N24415, N22897, N10140, N22014);
and AND4 (N24432, N24424, N18605, N1942, N8671);
not NOT1 (N24433, N24425);
nand NAND3 (N24434, N24426, N8843, N10916);
nand NAND2 (N24435, N24429, N9892);
not NOT1 (N24436, N24433);
and AND2 (N24437, N24421, N15008);
or OR3 (N24438, N24432, N2791, N1859);
buf BUF1 (N24439, N24430);
not NOT1 (N24440, N24427);
not NOT1 (N24441, N24440);
nand NAND2 (N24442, N24441, N18346);
buf BUF1 (N24443, N24442);
and AND2 (N24444, N24438, N3469);
nor NOR4 (N24445, N24436, N12072, N3292, N6797);
and AND4 (N24446, N24444, N4845, N11382, N13307);
xor XOR2 (N24447, N24423, N3342);
or OR3 (N24448, N24446, N2534, N6330);
or OR2 (N24449, N24443, N8017);
buf BUF1 (N24450, N24445);
or OR3 (N24451, N24448, N10579, N19523);
xor XOR2 (N24452, N24437, N15315);
or OR4 (N24453, N24451, N13373, N22210, N8898);
and AND4 (N24454, N24449, N24012, N1986, N12657);
not NOT1 (N24455, N24434);
nand NAND4 (N24456, N24428, N16153, N7479, N21846);
nor NOR3 (N24457, N24453, N17569, N8477);
not NOT1 (N24458, N24456);
xor XOR2 (N24459, N24431, N4709);
and AND3 (N24460, N24457, N11465, N8156);
or OR2 (N24461, N24458, N10991);
xor XOR2 (N24462, N24435, N3395);
nand NAND4 (N24463, N24455, N457, N15862, N9903);
xor XOR2 (N24464, N24454, N11767);
xor XOR2 (N24465, N24450, N4422);
not NOT1 (N24466, N24439);
nand NAND4 (N24467, N24452, N1105, N8014, N21569);
not NOT1 (N24468, N24464);
buf BUF1 (N24469, N24468);
not NOT1 (N24470, N24467);
buf BUF1 (N24471, N24470);
not NOT1 (N24472, N24465);
nand NAND2 (N24473, N24466, N17049);
and AND4 (N24474, N24461, N10765, N2611, N3745);
and AND2 (N24475, N24462, N18009);
buf BUF1 (N24476, N24463);
and AND2 (N24477, N24459, N20715);
nand NAND2 (N24478, N24476, N16913);
and AND4 (N24479, N24475, N22770, N2472, N15951);
and AND3 (N24480, N24447, N2402, N19319);
xor XOR2 (N24481, N24473, N23839);
or OR3 (N24482, N24474, N5602, N2448);
nor NOR2 (N24483, N24472, N4899);
not NOT1 (N24484, N24481);
nor NOR2 (N24485, N24482, N7697);
nand NAND4 (N24486, N24460, N21536, N16611, N4181);
nand NAND3 (N24487, N24483, N21360, N13168);
and AND3 (N24488, N24480, N11400, N8630);
or OR3 (N24489, N24477, N20323, N5250);
xor XOR2 (N24490, N24484, N6443);
xor XOR2 (N24491, N24478, N22272);
buf BUF1 (N24492, N24486);
xor XOR2 (N24493, N24492, N7699);
not NOT1 (N24494, N24485);
buf BUF1 (N24495, N24491);
nand NAND3 (N24496, N24471, N10868, N22276);
or OR2 (N24497, N24494, N1689);
nand NAND3 (N24498, N24479, N15252, N23057);
or OR3 (N24499, N24488, N4940, N6879);
xor XOR2 (N24500, N24498, N15853);
xor XOR2 (N24501, N24496, N21579);
and AND4 (N24502, N24500, N508, N2911, N12361);
and AND3 (N24503, N24497, N17545, N15822);
or OR4 (N24504, N24503, N9877, N535, N7414);
nand NAND4 (N24505, N24487, N13034, N13979, N13329);
and AND4 (N24506, N24469, N1319, N8463, N21587);
xor XOR2 (N24507, N24506, N17736);
nand NAND4 (N24508, N24504, N1733, N11097, N22936);
not NOT1 (N24509, N24502);
nor NOR3 (N24510, N24508, N8349, N1409);
buf BUF1 (N24511, N24505);
xor XOR2 (N24512, N24495, N12902);
not NOT1 (N24513, N24509);
and AND2 (N24514, N24512, N11680);
and AND2 (N24515, N24490, N3146);
or OR2 (N24516, N24499, N2286);
nor NOR4 (N24517, N24507, N11161, N3524, N15370);
buf BUF1 (N24518, N24516);
buf BUF1 (N24519, N24518);
or OR3 (N24520, N24501, N7936, N12889);
nand NAND4 (N24521, N24520, N17038, N9074, N23518);
and AND2 (N24522, N24493, N23612);
buf BUF1 (N24523, N24514);
nor NOR3 (N24524, N24521, N18226, N9569);
or OR4 (N24525, N24519, N21035, N20123, N4888);
or OR2 (N24526, N24510, N7773);
nor NOR3 (N24527, N24511, N15572, N3759);
xor XOR2 (N24528, N24523, N18729);
and AND4 (N24529, N24525, N17409, N6929, N24238);
not NOT1 (N24530, N24529);
nand NAND3 (N24531, N24515, N9409, N6264);
nand NAND2 (N24532, N24531, N733);
nand NAND3 (N24533, N24489, N21448, N14388);
nor NOR2 (N24534, N24532, N20554);
not NOT1 (N24535, N24517);
nand NAND4 (N24536, N24527, N19210, N20840, N22306);
and AND4 (N24537, N24533, N16282, N14570, N8782);
nand NAND4 (N24538, N24528, N787, N3446, N13892);
and AND2 (N24539, N24524, N14948);
or OR2 (N24540, N24536, N14518);
or OR3 (N24541, N24513, N915, N3767);
and AND3 (N24542, N24537, N19964, N22189);
not NOT1 (N24543, N24535);
and AND3 (N24544, N24538, N16964, N13574);
buf BUF1 (N24545, N24542);
or OR4 (N24546, N24534, N381, N19068, N24267);
xor XOR2 (N24547, N24545, N4640);
buf BUF1 (N24548, N24530);
nand NAND3 (N24549, N24548, N17739, N12123);
buf BUF1 (N24550, N24522);
nor NOR4 (N24551, N24547, N12992, N21980, N19637);
not NOT1 (N24552, N24546);
buf BUF1 (N24553, N24541);
not NOT1 (N24554, N24526);
buf BUF1 (N24555, N24550);
nor NOR4 (N24556, N24552, N23925, N21263, N15391);
not NOT1 (N24557, N24551);
nand NAND4 (N24558, N24549, N20434, N23386, N1910);
not NOT1 (N24559, N24557);
nand NAND2 (N24560, N24540, N19468);
xor XOR2 (N24561, N24560, N10910);
xor XOR2 (N24562, N24555, N10699);
and AND4 (N24563, N24543, N22035, N20749, N20556);
nand NAND4 (N24564, N24563, N23056, N11713, N14547);
buf BUF1 (N24565, N24556);
or OR2 (N24566, N24561, N4973);
buf BUF1 (N24567, N24554);
nor NOR2 (N24568, N24562, N19806);
xor XOR2 (N24569, N24565, N14231);
nor NOR3 (N24570, N24553, N5767, N13978);
not NOT1 (N24571, N24559);
not NOT1 (N24572, N24544);
not NOT1 (N24573, N24572);
nand NAND3 (N24574, N24573, N17450, N23871);
and AND4 (N24575, N24574, N5984, N3720, N8544);
nand NAND2 (N24576, N24539, N8764);
nor NOR3 (N24577, N24567, N11204, N23632);
and AND3 (N24578, N24571, N15072, N8137);
nand NAND2 (N24579, N24577, N8858);
xor XOR2 (N24580, N24575, N14215);
nor NOR2 (N24581, N24580, N14643);
xor XOR2 (N24582, N24569, N7674);
or OR2 (N24583, N24568, N2846);
xor XOR2 (N24584, N24579, N13851);
nor NOR2 (N24585, N24584, N4882);
and AND3 (N24586, N24582, N18517, N9008);
nor NOR4 (N24587, N24570, N21078, N23388, N19488);
nand NAND4 (N24588, N24558, N1876, N19296, N9715);
buf BUF1 (N24589, N24588);
or OR3 (N24590, N24587, N16113, N5517);
nor NOR3 (N24591, N24583, N11154, N12398);
nor NOR2 (N24592, N24589, N13815);
nand NAND3 (N24593, N24581, N24002, N19466);
or OR3 (N24594, N24564, N18700, N1063);
not NOT1 (N24595, N24590);
buf BUF1 (N24596, N24586);
xor XOR2 (N24597, N24596, N15347);
and AND4 (N24598, N24592, N14582, N7730, N2733);
nand NAND3 (N24599, N24598, N3269, N9344);
xor XOR2 (N24600, N24591, N23506);
nor NOR3 (N24601, N24585, N3415, N16757);
nand NAND4 (N24602, N24597, N11438, N5532, N22192);
nor NOR3 (N24603, N24576, N7744, N7503);
and AND3 (N24604, N24602, N4683, N20466);
and AND2 (N24605, N24593, N4151);
nor NOR2 (N24606, N24600, N23225);
nor NOR3 (N24607, N24594, N20727, N20305);
nand NAND2 (N24608, N24606, N12632);
and AND2 (N24609, N24601, N19689);
nand NAND3 (N24610, N24578, N7991, N9740);
xor XOR2 (N24611, N24604, N6454);
nor NOR3 (N24612, N24609, N3756, N2299);
not NOT1 (N24613, N24566);
not NOT1 (N24614, N24611);
xor XOR2 (N24615, N24595, N10825);
not NOT1 (N24616, N24599);
buf BUF1 (N24617, N24603);
nor NOR2 (N24618, N24612, N207);
buf BUF1 (N24619, N24610);
nor NOR3 (N24620, N24617, N17600, N23093);
nand NAND4 (N24621, N24618, N22464, N23115, N17542);
xor XOR2 (N24622, N24605, N24501);
buf BUF1 (N24623, N24608);
not NOT1 (N24624, N24613);
not NOT1 (N24625, N24607);
nand NAND3 (N24626, N24615, N11152, N10203);
or OR3 (N24627, N24621, N3682, N11139);
not NOT1 (N24628, N24623);
or OR3 (N24629, N24614, N7185, N21821);
buf BUF1 (N24630, N24624);
xor XOR2 (N24631, N24616, N6922);
nor NOR2 (N24632, N24628, N5243);
xor XOR2 (N24633, N24631, N8177);
and AND3 (N24634, N24633, N2098, N6852);
nor NOR2 (N24635, N24632, N1505);
buf BUF1 (N24636, N24627);
and AND3 (N24637, N24636, N10665, N16740);
nor NOR3 (N24638, N24634, N19804, N10905);
or OR4 (N24639, N24625, N17710, N12035, N17815);
xor XOR2 (N24640, N24620, N1679);
or OR3 (N24641, N24629, N6376, N12235);
xor XOR2 (N24642, N24630, N6557);
nor NOR4 (N24643, N24622, N1543, N15469, N7377);
buf BUF1 (N24644, N24626);
nand NAND2 (N24645, N24637, N11769);
nor NOR3 (N24646, N24640, N1598, N1154);
nand NAND2 (N24647, N24646, N22766);
not NOT1 (N24648, N24644);
or OR3 (N24649, N24643, N19297, N2227);
and AND4 (N24650, N24648, N10193, N16325, N10207);
or OR4 (N24651, N24649, N17054, N16398, N1435);
buf BUF1 (N24652, N24638);
nor NOR3 (N24653, N24650, N18552, N7513);
or OR2 (N24654, N24635, N9506);
xor XOR2 (N24655, N24647, N13944);
not NOT1 (N24656, N24654);
nor NOR3 (N24657, N24655, N23132, N186);
nand NAND4 (N24658, N24653, N16914, N13618, N4905);
nand NAND4 (N24659, N24656, N2879, N22287, N5058);
or OR2 (N24660, N24652, N11733);
buf BUF1 (N24661, N24642);
not NOT1 (N24662, N24661);
not NOT1 (N24663, N24662);
and AND2 (N24664, N24657, N18440);
and AND4 (N24665, N24658, N7741, N18734, N8590);
buf BUF1 (N24666, N24663);
nor NOR2 (N24667, N24645, N14541);
xor XOR2 (N24668, N24641, N12174);
not NOT1 (N24669, N24667);
xor XOR2 (N24670, N24659, N13752);
nor NOR3 (N24671, N24668, N5522, N19346);
not NOT1 (N24672, N24664);
xor XOR2 (N24673, N24666, N15803);
nor NOR4 (N24674, N24673, N8470, N8884, N2449);
xor XOR2 (N24675, N24674, N2359);
not NOT1 (N24676, N24665);
and AND2 (N24677, N24651, N5991);
not NOT1 (N24678, N24669);
nand NAND3 (N24679, N24671, N17991, N15844);
buf BUF1 (N24680, N24679);
nor NOR2 (N24681, N24619, N9232);
nand NAND2 (N24682, N24660, N21608);
nor NOR3 (N24683, N24639, N8819, N5221);
not NOT1 (N24684, N24670);
nor NOR2 (N24685, N24678, N4665);
not NOT1 (N24686, N24677);
buf BUF1 (N24687, N24675);
not NOT1 (N24688, N24672);
or OR2 (N24689, N24684, N2888);
and AND3 (N24690, N24681, N10101, N22475);
not NOT1 (N24691, N24689);
nor NOR3 (N24692, N24687, N2770, N10040);
buf BUF1 (N24693, N24690);
xor XOR2 (N24694, N24688, N13436);
buf BUF1 (N24695, N24686);
xor XOR2 (N24696, N24683, N12771);
or OR2 (N24697, N24691, N3036);
or OR3 (N24698, N24685, N18972, N3875);
nand NAND3 (N24699, N24696, N10936, N20951);
nor NOR3 (N24700, N24692, N23254, N1443);
and AND3 (N24701, N24682, N12949, N8477);
nand NAND2 (N24702, N24700, N21667);
and AND2 (N24703, N24680, N15278);
not NOT1 (N24704, N24703);
nor NOR3 (N24705, N24704, N3995, N844);
nor NOR4 (N24706, N24702, N8055, N14160, N17227);
not NOT1 (N24707, N24693);
nor NOR2 (N24708, N24697, N11892);
xor XOR2 (N24709, N24708, N23192);
not NOT1 (N24710, N24701);
nand NAND4 (N24711, N24699, N5957, N11602, N13907);
nand NAND3 (N24712, N24695, N16236, N15247);
or OR4 (N24713, N24694, N5250, N3248, N1854);
nor NOR4 (N24714, N24707, N18872, N7526, N12654);
nor NOR3 (N24715, N24698, N10938, N24282);
or OR2 (N24716, N24706, N1308);
buf BUF1 (N24717, N24676);
nand NAND3 (N24718, N24715, N22571, N7466);
not NOT1 (N24719, N24718);
and AND3 (N24720, N24705, N14663, N10397);
nand NAND3 (N24721, N24712, N1943, N4804);
not NOT1 (N24722, N24709);
or OR2 (N24723, N24713, N20670);
nand NAND2 (N24724, N24716, N15191);
and AND4 (N24725, N24719, N12045, N23120, N8517);
or OR2 (N24726, N24722, N23713);
nor NOR3 (N24727, N24724, N5553, N4324);
or OR4 (N24728, N24725, N7015, N5632, N2161);
and AND3 (N24729, N24720, N11155, N1686);
nor NOR3 (N24730, N24727, N14036, N3877);
buf BUF1 (N24731, N24726);
buf BUF1 (N24732, N24711);
or OR2 (N24733, N24728, N520);
nor NOR3 (N24734, N24714, N2707, N19342);
not NOT1 (N24735, N24729);
and AND2 (N24736, N24733, N14314);
nand NAND4 (N24737, N24730, N1814, N22784, N6482);
buf BUF1 (N24738, N24717);
buf BUF1 (N24739, N24732);
nor NOR4 (N24740, N24737, N20913, N2920, N2876);
nand NAND2 (N24741, N24740, N2834);
nand NAND4 (N24742, N24731, N13665, N19118, N890);
or OR3 (N24743, N24723, N9531, N10086);
not NOT1 (N24744, N24739);
not NOT1 (N24745, N24743);
or OR2 (N24746, N24735, N17728);
not NOT1 (N24747, N24746);
or OR2 (N24748, N24710, N20020);
or OR4 (N24749, N24741, N9285, N13597, N16977);
nor NOR4 (N24750, N24742, N10733, N1441, N21553);
nand NAND4 (N24751, N24744, N9460, N20187, N1979);
not NOT1 (N24752, N24747);
xor XOR2 (N24753, N24751, N23949);
xor XOR2 (N24754, N24749, N19159);
xor XOR2 (N24755, N24734, N21113);
nor NOR4 (N24756, N24721, N11068, N4452, N16465);
and AND2 (N24757, N24754, N4290);
not NOT1 (N24758, N24753);
not NOT1 (N24759, N24757);
nand NAND4 (N24760, N24756, N4397, N17826, N10994);
buf BUF1 (N24761, N24759);
and AND3 (N24762, N24761, N3883, N15561);
not NOT1 (N24763, N24745);
nand NAND4 (N24764, N24758, N17748, N12095, N13949);
xor XOR2 (N24765, N24755, N1694);
xor XOR2 (N24766, N24736, N42);
not NOT1 (N24767, N24760);
nand NAND4 (N24768, N24752, N13229, N8752, N17309);
nand NAND3 (N24769, N24764, N17355, N22070);
not NOT1 (N24770, N24762);
not NOT1 (N24771, N24763);
nor NOR4 (N24772, N24767, N2740, N22417, N15710);
nand NAND4 (N24773, N24738, N6212, N6221, N6008);
buf BUF1 (N24774, N24748);
nor NOR3 (N24775, N24770, N1175, N22236);
xor XOR2 (N24776, N24771, N9188);
xor XOR2 (N24777, N24774, N15114);
nand NAND2 (N24778, N24775, N10311);
and AND4 (N24779, N24768, N19339, N17914, N16856);
buf BUF1 (N24780, N24772);
xor XOR2 (N24781, N24765, N3434);
buf BUF1 (N24782, N24773);
and AND2 (N24783, N24776, N9836);
xor XOR2 (N24784, N24778, N3216);
buf BUF1 (N24785, N24779);
xor XOR2 (N24786, N24766, N6761);
buf BUF1 (N24787, N24769);
nand NAND2 (N24788, N24777, N13511);
xor XOR2 (N24789, N24786, N12699);
xor XOR2 (N24790, N24784, N7161);
xor XOR2 (N24791, N24785, N6909);
xor XOR2 (N24792, N24787, N7441);
nand NAND2 (N24793, N24782, N5553);
nand NAND2 (N24794, N24781, N16704);
xor XOR2 (N24795, N24794, N11724);
nor NOR4 (N24796, N24791, N11311, N22243, N14929);
nand NAND4 (N24797, N24788, N22153, N16607, N7230);
buf BUF1 (N24798, N24780);
nand NAND2 (N24799, N24798, N4952);
not NOT1 (N24800, N24790);
not NOT1 (N24801, N24797);
xor XOR2 (N24802, N24792, N1729);
or OR2 (N24803, N24796, N950);
and AND3 (N24804, N24789, N17746, N9796);
xor XOR2 (N24805, N24802, N15803);
buf BUF1 (N24806, N24750);
nor NOR2 (N24807, N24805, N6732);
nor NOR3 (N24808, N24806, N4308, N4864);
nor NOR3 (N24809, N24804, N10625, N9921);
nand NAND4 (N24810, N24809, N10658, N24687, N567);
and AND3 (N24811, N24808, N24301, N18213);
xor XOR2 (N24812, N24795, N10090);
not NOT1 (N24813, N24793);
not NOT1 (N24814, N24799);
or OR2 (N24815, N24810, N1695);
nand NAND4 (N24816, N24801, N3889, N9456, N21320);
nand NAND3 (N24817, N24815, N21193, N6989);
buf BUF1 (N24818, N24812);
buf BUF1 (N24819, N24811);
nand NAND2 (N24820, N24816, N23137);
or OR2 (N24821, N24820, N10570);
nand NAND4 (N24822, N24817, N8693, N5314, N16405);
nor NOR4 (N24823, N24821, N21161, N19552, N10182);
or OR2 (N24824, N24814, N9352);
xor XOR2 (N24825, N24818, N9988);
nor NOR2 (N24826, N24823, N2912);
buf BUF1 (N24827, N24822);
and AND2 (N24828, N24803, N5450);
buf BUF1 (N24829, N24800);
or OR3 (N24830, N24783, N17798, N8970);
xor XOR2 (N24831, N24829, N11448);
and AND2 (N24832, N24825, N17039);
xor XOR2 (N24833, N24824, N12496);
or OR4 (N24834, N24826, N20272, N7915, N16880);
or OR2 (N24835, N24832, N11319);
or OR4 (N24836, N24831, N10596, N3376, N897);
xor XOR2 (N24837, N24835, N7487);
nor NOR2 (N24838, N24807, N15468);
buf BUF1 (N24839, N24838);
nand NAND3 (N24840, N24839, N14491, N3907);
nand NAND4 (N24841, N24837, N15477, N4879, N18462);
not NOT1 (N24842, N24836);
and AND2 (N24843, N24833, N7762);
xor XOR2 (N24844, N24841, N10799);
nand NAND2 (N24845, N24843, N10707);
nand NAND3 (N24846, N24827, N20734, N13565);
nor NOR4 (N24847, N24844, N7117, N5409, N8542);
nor NOR2 (N24848, N24842, N12381);
nor NOR2 (N24849, N24830, N24072);
nor NOR4 (N24850, N24847, N2967, N12167, N12246);
or OR2 (N24851, N24849, N13456);
or OR3 (N24852, N24846, N21541, N1330);
xor XOR2 (N24853, N24828, N12658);
nand NAND3 (N24854, N24851, N4049, N8388);
not NOT1 (N24855, N24848);
buf BUF1 (N24856, N24850);
or OR3 (N24857, N24834, N9848, N19360);
xor XOR2 (N24858, N24840, N17330);
buf BUF1 (N24859, N24857);
xor XOR2 (N24860, N24845, N17999);
and AND2 (N24861, N24858, N8695);
or OR2 (N24862, N24855, N13112);
nand NAND3 (N24863, N24819, N16241, N8877);
xor XOR2 (N24864, N24856, N16581);
xor XOR2 (N24865, N24854, N5222);
not NOT1 (N24866, N24813);
and AND4 (N24867, N24860, N20081, N21920, N3114);
and AND3 (N24868, N24867, N14757, N4106);
or OR4 (N24869, N24863, N18505, N19918, N23098);
not NOT1 (N24870, N24859);
xor XOR2 (N24871, N24868, N5870);
and AND3 (N24872, N24862, N1595, N19516);
nand NAND3 (N24873, N24866, N2665, N23037);
xor XOR2 (N24874, N24872, N13523);
or OR3 (N24875, N24874, N14987, N18238);
or OR3 (N24876, N24865, N428, N8658);
nand NAND2 (N24877, N24869, N6675);
xor XOR2 (N24878, N24871, N2412);
not NOT1 (N24879, N24878);
nor NOR2 (N24880, N24852, N15377);
or OR4 (N24881, N24853, N9238, N17609, N9524);
or OR4 (N24882, N24861, N2142, N5124, N7980);
nand NAND2 (N24883, N24875, N9082);
not NOT1 (N24884, N24877);
nor NOR3 (N24885, N24884, N12988, N2188);
buf BUF1 (N24886, N24873);
and AND2 (N24887, N24883, N21957);
not NOT1 (N24888, N24870);
buf BUF1 (N24889, N24879);
and AND2 (N24890, N24887, N7633);
not NOT1 (N24891, N24882);
nand NAND3 (N24892, N24881, N11766, N22543);
nand NAND2 (N24893, N24891, N6683);
and AND4 (N24894, N24892, N24342, N9798, N5073);
nand NAND3 (N24895, N24876, N6688, N19316);
buf BUF1 (N24896, N24895);
buf BUF1 (N24897, N24864);
buf BUF1 (N24898, N24889);
or OR3 (N24899, N24885, N16238, N10766);
xor XOR2 (N24900, N24899, N11545);
nand NAND4 (N24901, N24897, N11251, N2731, N13779);
buf BUF1 (N24902, N24896);
nor NOR3 (N24903, N24901, N817, N18465);
buf BUF1 (N24904, N24898);
nor NOR4 (N24905, N24890, N20000, N17121, N14759);
not NOT1 (N24906, N24902);
buf BUF1 (N24907, N24880);
xor XOR2 (N24908, N24907, N12313);
nand NAND3 (N24909, N24900, N8344, N19129);
or OR2 (N24910, N24893, N796);
buf BUF1 (N24911, N24906);
and AND3 (N24912, N24888, N450, N2048);
nand NAND4 (N24913, N24908, N18205, N9796, N14695);
or OR2 (N24914, N24912, N333);
not NOT1 (N24915, N24911);
or OR3 (N24916, N24915, N10793, N24);
xor XOR2 (N24917, N24914, N4489);
not NOT1 (N24918, N24913);
nor NOR3 (N24919, N24903, N7613, N8367);
and AND4 (N24920, N24905, N4626, N14967, N5333);
nor NOR3 (N24921, N24904, N10284, N22177);
xor XOR2 (N24922, N24920, N22531);
or OR3 (N24923, N24894, N20572, N9467);
nand NAND4 (N24924, N24917, N22687, N6981, N22804);
nand NAND3 (N24925, N24922, N8008, N11378);
nor NOR2 (N24926, N24886, N7681);
buf BUF1 (N24927, N24923);
not NOT1 (N24928, N24919);
nand NAND4 (N24929, N24916, N12982, N21118, N15558);
or OR4 (N24930, N24924, N11109, N1993, N16560);
nand NAND3 (N24931, N24910, N9915, N1563);
not NOT1 (N24932, N24929);
nor NOR4 (N24933, N24925, N5859, N11137, N23192);
and AND4 (N24934, N24926, N19549, N20085, N12099);
xor XOR2 (N24935, N24930, N12676);
buf BUF1 (N24936, N24909);
xor XOR2 (N24937, N24933, N6091);
not NOT1 (N24938, N24932);
or OR2 (N24939, N24937, N22897);
nand NAND2 (N24940, N24927, N13124);
not NOT1 (N24941, N24935);
buf BUF1 (N24942, N24939);
or OR3 (N24943, N24918, N15708, N5361);
xor XOR2 (N24944, N24931, N20099);
not NOT1 (N24945, N24940);
or OR4 (N24946, N24921, N6692, N6446, N17043);
buf BUF1 (N24947, N24941);
and AND4 (N24948, N24938, N15660, N23519, N9330);
or OR2 (N24949, N24944, N20811);
or OR4 (N24950, N24948, N3270, N14880, N23143);
or OR3 (N24951, N24928, N11648, N9560);
or OR2 (N24952, N24949, N10892);
and AND2 (N24953, N24950, N13564);
nand NAND3 (N24954, N24952, N5002, N12265);
and AND3 (N24955, N24951, N15990, N24282);
buf BUF1 (N24956, N24942);
or OR3 (N24957, N24954, N19572, N7248);
xor XOR2 (N24958, N24943, N636);
nor NOR4 (N24959, N24946, N19454, N15722, N7553);
nand NAND2 (N24960, N24958, N22414);
or OR2 (N24961, N24959, N9123);
not NOT1 (N24962, N24936);
and AND2 (N24963, N24947, N3185);
buf BUF1 (N24964, N24934);
not NOT1 (N24965, N24955);
not NOT1 (N24966, N24964);
buf BUF1 (N24967, N24953);
not NOT1 (N24968, N24961);
and AND4 (N24969, N24968, N9489, N5172, N2316);
nand NAND4 (N24970, N24945, N16360, N22640, N11542);
nand NAND2 (N24971, N24956, N17246);
or OR2 (N24972, N24962, N2722);
nand NAND3 (N24973, N24971, N2095, N11187);
nand NAND4 (N24974, N24966, N4201, N22338, N13480);
buf BUF1 (N24975, N24972);
xor XOR2 (N24976, N24973, N1492);
nor NOR2 (N24977, N24976, N2473);
xor XOR2 (N24978, N24970, N3341);
or OR4 (N24979, N24960, N7688, N9292, N3343);
not NOT1 (N24980, N24963);
or OR3 (N24981, N24975, N15430, N4216);
xor XOR2 (N24982, N24979, N8402);
or OR4 (N24983, N24982, N20245, N13651, N2573);
or OR4 (N24984, N24977, N3404, N24662, N11116);
buf BUF1 (N24985, N24980);
and AND2 (N24986, N24981, N2474);
nor NOR2 (N24987, N24985, N2965);
nand NAND2 (N24988, N24957, N22400);
or OR2 (N24989, N24983, N15659);
buf BUF1 (N24990, N24969);
or OR2 (N24991, N24978, N24057);
nand NAND2 (N24992, N24987, N19543);
or OR4 (N24993, N24984, N9877, N10828, N23394);
xor XOR2 (N24994, N24989, N12719);
xor XOR2 (N24995, N24991, N9941);
and AND3 (N24996, N24967, N5878, N265);
nand NAND2 (N24997, N24995, N12876);
nor NOR3 (N24998, N24996, N19778, N22041);
xor XOR2 (N24999, N24988, N20492);
nand NAND3 (N25000, N24997, N4081, N9836);
nand NAND3 (N25001, N24986, N19136, N16200);
nor NOR4 (N25002, N24994, N4143, N1006, N9139);
not NOT1 (N25003, N25002);
or OR3 (N25004, N24993, N16453, N16540);
buf BUF1 (N25005, N25004);
nor NOR4 (N25006, N24990, N11132, N15454, N18521);
xor XOR2 (N25007, N24992, N6585);
xor XOR2 (N25008, N24974, N2526);
buf BUF1 (N25009, N25005);
buf BUF1 (N25010, N24998);
buf BUF1 (N25011, N25006);
xor XOR2 (N25012, N25007, N10321);
xor XOR2 (N25013, N25009, N13632);
xor XOR2 (N25014, N25012, N16664);
not NOT1 (N25015, N25011);
nor NOR4 (N25016, N25015, N11246, N19771, N23267);
nor NOR4 (N25017, N25003, N19950, N22278, N7870);
nand NAND4 (N25018, N25017, N2564, N14640, N1131);
buf BUF1 (N25019, N24999);
not NOT1 (N25020, N25010);
and AND3 (N25021, N25008, N19251, N8748);
or OR2 (N25022, N25016, N20375);
and AND3 (N25023, N25000, N10631, N14739);
xor XOR2 (N25024, N25019, N4731);
buf BUF1 (N25025, N25001);
nand NAND3 (N25026, N24965, N6427, N19552);
not NOT1 (N25027, N25025);
xor XOR2 (N25028, N25027, N19012);
xor XOR2 (N25029, N25020, N5489);
xor XOR2 (N25030, N25014, N18857);
buf BUF1 (N25031, N25018);
or OR3 (N25032, N25024, N22444, N17430);
nor NOR2 (N25033, N25030, N7906);
or OR4 (N25034, N25026, N21745, N23488, N5925);
xor XOR2 (N25035, N25034, N8192);
nand NAND3 (N25036, N25035, N14553, N1122);
buf BUF1 (N25037, N25023);
nor NOR3 (N25038, N25022, N9099, N16820);
or OR4 (N25039, N25028, N17365, N4517, N5332);
and AND3 (N25040, N25039, N6175, N15591);
buf BUF1 (N25041, N25031);
nor NOR4 (N25042, N25037, N11107, N1207, N8804);
and AND2 (N25043, N25032, N22506);
or OR3 (N25044, N25021, N18861, N9883);
or OR3 (N25045, N25029, N4310, N22921);
nand NAND4 (N25046, N25044, N19187, N15875, N11228);
buf BUF1 (N25047, N25043);
buf BUF1 (N25048, N25036);
nor NOR4 (N25049, N25046, N16679, N7744, N11989);
or OR2 (N25050, N25048, N5756);
or OR4 (N25051, N25040, N24150, N9454, N1758);
and AND2 (N25052, N25041, N4629);
or OR2 (N25053, N25051, N17128);
nand NAND4 (N25054, N25013, N13518, N22588, N15216);
or OR3 (N25055, N25053, N10662, N5021);
and AND2 (N25056, N25052, N15117);
and AND3 (N25057, N25049, N6315, N12583);
nor NOR3 (N25058, N25045, N18843, N18663);
buf BUF1 (N25059, N25050);
nor NOR3 (N25060, N25047, N16886, N24308);
or OR4 (N25061, N25056, N22675, N19155, N6734);
not NOT1 (N25062, N25042);
nor NOR3 (N25063, N25061, N19040, N10872);
xor XOR2 (N25064, N25063, N18456);
nor NOR4 (N25065, N25033, N16163, N3619, N12980);
buf BUF1 (N25066, N25055);
or OR3 (N25067, N25064, N16290, N25010);
not NOT1 (N25068, N25058);
or OR3 (N25069, N25067, N21849, N18123);
xor XOR2 (N25070, N25057, N20303);
or OR2 (N25071, N25059, N6833);
nand NAND2 (N25072, N25071, N19654);
nand NAND4 (N25073, N25062, N11693, N5399, N20561);
and AND3 (N25074, N25060, N19251, N4261);
nor NOR3 (N25075, N25072, N12372, N21611);
not NOT1 (N25076, N25074);
and AND3 (N25077, N25054, N11089, N17605);
or OR3 (N25078, N25075, N19461, N14102);
nand NAND4 (N25079, N25065, N5061, N14423, N23780);
xor XOR2 (N25080, N25077, N19284);
or OR3 (N25081, N25070, N3515, N7624);
nand NAND4 (N25082, N25066, N24046, N22269, N9684);
not NOT1 (N25083, N25078);
buf BUF1 (N25084, N25080);
and AND4 (N25085, N25068, N6283, N4820, N3256);
buf BUF1 (N25086, N25073);
buf BUF1 (N25087, N25086);
and AND4 (N25088, N25083, N9609, N2856, N20736);
nor NOR2 (N25089, N25069, N21535);
xor XOR2 (N25090, N25089, N19074);
or OR3 (N25091, N25088, N16005, N21263);
xor XOR2 (N25092, N25085, N11252);
nand NAND3 (N25093, N25082, N4889, N5988);
not NOT1 (N25094, N25091);
not NOT1 (N25095, N25084);
xor XOR2 (N25096, N25092, N10599);
not NOT1 (N25097, N25081);
xor XOR2 (N25098, N25090, N1165);
xor XOR2 (N25099, N25076, N14636);
and AND2 (N25100, N25079, N16119);
or OR2 (N25101, N25097, N6638);
nand NAND4 (N25102, N25087, N12819, N17359, N24474);
buf BUF1 (N25103, N25038);
buf BUF1 (N25104, N25100);
nor NOR2 (N25105, N25102, N17590);
buf BUF1 (N25106, N25094);
buf BUF1 (N25107, N25101);
nand NAND3 (N25108, N25103, N13745, N16959);
nor NOR2 (N25109, N25095, N21903);
nor NOR2 (N25110, N25109, N23211);
buf BUF1 (N25111, N25106);
nand NAND3 (N25112, N25104, N16472, N17481);
xor XOR2 (N25113, N25099, N12931);
buf BUF1 (N25114, N25108);
and AND3 (N25115, N25111, N22335, N10288);
not NOT1 (N25116, N25107);
nand NAND2 (N25117, N25105, N23143);
not NOT1 (N25118, N25098);
nand NAND2 (N25119, N25110, N6301);
nor NOR2 (N25120, N25116, N20990);
not NOT1 (N25121, N25115);
nor NOR2 (N25122, N25117, N11288);
xor XOR2 (N25123, N25118, N5975);
nand NAND3 (N25124, N25120, N22621, N18968);
not NOT1 (N25125, N25124);
buf BUF1 (N25126, N25122);
nor NOR4 (N25127, N25112, N20084, N2377, N19915);
not NOT1 (N25128, N25113);
or OR4 (N25129, N25121, N23975, N14715, N24118);
and AND4 (N25130, N25125, N20111, N9475, N5301);
and AND3 (N25131, N25093, N2658, N17246);
buf BUF1 (N25132, N25096);
and AND2 (N25133, N25129, N24112);
or OR4 (N25134, N25133, N18394, N8749, N3868);
xor XOR2 (N25135, N25130, N13479);
or OR3 (N25136, N25126, N12928, N19422);
and AND2 (N25137, N25131, N602);
and AND3 (N25138, N25132, N24954, N8749);
or OR2 (N25139, N25136, N4351);
nor NOR2 (N25140, N25119, N21463);
nand NAND4 (N25141, N25128, N172, N7106, N7299);
xor XOR2 (N25142, N25140, N7326);
not NOT1 (N25143, N25127);
buf BUF1 (N25144, N25141);
xor XOR2 (N25145, N25142, N5414);
xor XOR2 (N25146, N25144, N12372);
not NOT1 (N25147, N25143);
buf BUF1 (N25148, N25145);
not NOT1 (N25149, N25123);
buf BUF1 (N25150, N25149);
xor XOR2 (N25151, N25137, N14747);
nor NOR2 (N25152, N25146, N12117);
buf BUF1 (N25153, N25150);
and AND3 (N25154, N25148, N16093, N24980);
nand NAND4 (N25155, N25114, N12036, N2514, N5792);
not NOT1 (N25156, N25151);
not NOT1 (N25157, N25147);
nor NOR2 (N25158, N25157, N8694);
not NOT1 (N25159, N25158);
or OR4 (N25160, N25154, N11362, N23726, N796);
buf BUF1 (N25161, N25153);
nor NOR4 (N25162, N25156, N11117, N8707, N1902);
buf BUF1 (N25163, N25162);
or OR3 (N25164, N25135, N14059, N17154);
not NOT1 (N25165, N25164);
and AND3 (N25166, N25134, N24862, N21137);
not NOT1 (N25167, N25163);
xor XOR2 (N25168, N25159, N20183);
and AND3 (N25169, N25152, N7403, N6880);
and AND2 (N25170, N25168, N16922);
buf BUF1 (N25171, N25160);
and AND2 (N25172, N25167, N13842);
buf BUF1 (N25173, N25139);
xor XOR2 (N25174, N25171, N7618);
nor NOR2 (N25175, N25169, N20700);
xor XOR2 (N25176, N25170, N15612);
and AND3 (N25177, N25173, N5829, N15868);
buf BUF1 (N25178, N25175);
xor XOR2 (N25179, N25177, N24701);
or OR3 (N25180, N25176, N17339, N17828);
and AND3 (N25181, N25172, N21296, N9468);
xor XOR2 (N25182, N25179, N20005);
not NOT1 (N25183, N25178);
nand NAND3 (N25184, N25180, N3259, N14703);
nor NOR3 (N25185, N25181, N23294, N10135);
not NOT1 (N25186, N25174);
nand NAND2 (N25187, N25185, N12573);
or OR4 (N25188, N25182, N2070, N223, N21504);
and AND4 (N25189, N25155, N3846, N21109, N18468);
or OR2 (N25190, N25166, N23858);
buf BUF1 (N25191, N25183);
not NOT1 (N25192, N25165);
nor NOR4 (N25193, N25187, N18057, N2511, N1803);
buf BUF1 (N25194, N25161);
xor XOR2 (N25195, N25138, N13466);
not NOT1 (N25196, N25184);
nor NOR3 (N25197, N25189, N1947, N21698);
nor NOR2 (N25198, N25192, N16757);
not NOT1 (N25199, N25191);
nor NOR2 (N25200, N25195, N2311);
not NOT1 (N25201, N25186);
nor NOR4 (N25202, N25194, N14663, N2327, N2822);
nand NAND3 (N25203, N25202, N15710, N2150);
or OR3 (N25204, N25198, N16704, N10739);
and AND3 (N25205, N25197, N8737, N21720);
not NOT1 (N25206, N25199);
nor NOR3 (N25207, N25193, N6877, N4478);
not NOT1 (N25208, N25200);
nand NAND2 (N25209, N25204, N7215);
nand NAND4 (N25210, N25209, N23765, N21624, N4934);
xor XOR2 (N25211, N25201, N21918);
nand NAND3 (N25212, N25205, N7851, N9326);
not NOT1 (N25213, N25206);
and AND2 (N25214, N25212, N24201);
xor XOR2 (N25215, N25207, N11333);
xor XOR2 (N25216, N25214, N17802);
or OR3 (N25217, N25213, N10677, N15264);
nand NAND3 (N25218, N25203, N20189, N8350);
or OR4 (N25219, N25217, N5649, N15536, N15148);
and AND3 (N25220, N25219, N6395, N8140);
not NOT1 (N25221, N25218);
xor XOR2 (N25222, N25216, N23921);
and AND3 (N25223, N25188, N14067, N9580);
or OR4 (N25224, N25210, N18584, N24541, N10362);
and AND2 (N25225, N25220, N16463);
and AND2 (N25226, N25208, N23229);
nor NOR4 (N25227, N25211, N7114, N7422, N7548);
nand NAND4 (N25228, N25227, N13157, N14758, N4309);
xor XOR2 (N25229, N25222, N12469);
nor NOR3 (N25230, N25229, N517, N14014);
not NOT1 (N25231, N25196);
and AND4 (N25232, N25230, N22021, N21135, N10385);
nor NOR2 (N25233, N25231, N8441);
or OR4 (N25234, N25233, N22958, N12951, N23338);
or OR4 (N25235, N25190, N18219, N4325, N11736);
not NOT1 (N25236, N25228);
and AND2 (N25237, N25223, N15982);
and AND3 (N25238, N25221, N1390, N19716);
nand NAND2 (N25239, N25215, N13149);
or OR2 (N25240, N25234, N19961);
nand NAND3 (N25241, N25236, N21526, N18875);
nand NAND2 (N25242, N25241, N12978);
not NOT1 (N25243, N25240);
or OR3 (N25244, N25235, N20398, N7953);
not NOT1 (N25245, N25224);
xor XOR2 (N25246, N25237, N22327);
buf BUF1 (N25247, N25232);
nand NAND3 (N25248, N25246, N22863, N22386);
not NOT1 (N25249, N25244);
and AND2 (N25250, N25225, N4232);
and AND3 (N25251, N25248, N3251, N14818);
and AND3 (N25252, N25247, N10968, N18149);
and AND2 (N25253, N25242, N11247);
and AND2 (N25254, N25251, N13116);
not NOT1 (N25255, N25250);
nor NOR4 (N25256, N25226, N455, N21330, N24790);
xor XOR2 (N25257, N25252, N3981);
or OR3 (N25258, N25249, N20067, N4698);
or OR2 (N25259, N25245, N18417);
not NOT1 (N25260, N25239);
and AND2 (N25261, N25257, N415);
xor XOR2 (N25262, N25255, N19105);
nand NAND4 (N25263, N25256, N12322, N6456, N14952);
not NOT1 (N25264, N25258);
nand NAND4 (N25265, N25259, N21512, N8354, N13522);
xor XOR2 (N25266, N25253, N14444);
buf BUF1 (N25267, N25264);
or OR2 (N25268, N25266, N11894);
buf BUF1 (N25269, N25265);
xor XOR2 (N25270, N25263, N13514);
or OR2 (N25271, N25260, N22060);
nand NAND3 (N25272, N25261, N17396, N7178);
or OR3 (N25273, N25254, N803, N1772);
buf BUF1 (N25274, N25267);
not NOT1 (N25275, N25270);
or OR2 (N25276, N25238, N6473);
not NOT1 (N25277, N25268);
not NOT1 (N25278, N25276);
xor XOR2 (N25279, N25273, N6016);
not NOT1 (N25280, N25272);
buf BUF1 (N25281, N25271);
buf BUF1 (N25282, N25269);
nor NOR4 (N25283, N25279, N15465, N19765, N10939);
xor XOR2 (N25284, N25243, N15453);
or OR3 (N25285, N25274, N9280, N18605);
nor NOR4 (N25286, N25284, N22222, N448, N3276);
buf BUF1 (N25287, N25281);
nand NAND4 (N25288, N25280, N973, N20674, N7066);
xor XOR2 (N25289, N25288, N24776);
or OR3 (N25290, N25287, N14498, N22545);
xor XOR2 (N25291, N25289, N2258);
buf BUF1 (N25292, N25286);
nand NAND4 (N25293, N25262, N18499, N22713, N4471);
buf BUF1 (N25294, N25293);
not NOT1 (N25295, N25277);
buf BUF1 (N25296, N25278);
not NOT1 (N25297, N25282);
or OR3 (N25298, N25285, N12543, N12800);
xor XOR2 (N25299, N25294, N24888);
nor NOR3 (N25300, N25283, N5046, N8356);
not NOT1 (N25301, N25296);
nor NOR3 (N25302, N25301, N12678, N89);
xor XOR2 (N25303, N25291, N14160);
not NOT1 (N25304, N25295);
nor NOR4 (N25305, N25303, N3253, N843, N15335);
or OR4 (N25306, N25302, N7879, N11463, N10119);
buf BUF1 (N25307, N25306);
nor NOR2 (N25308, N25299, N7239);
or OR2 (N25309, N25300, N15878);
nand NAND3 (N25310, N25307, N17623, N22301);
nor NOR3 (N25311, N25305, N19805, N6177);
xor XOR2 (N25312, N25308, N9516);
nor NOR3 (N25313, N25310, N1502, N15033);
nand NAND3 (N25314, N25298, N438, N20273);
not NOT1 (N25315, N25304);
or OR4 (N25316, N25297, N1714, N7379, N12026);
buf BUF1 (N25317, N25292);
and AND4 (N25318, N25290, N22216, N21832, N24434);
or OR2 (N25319, N25313, N3326);
not NOT1 (N25320, N25312);
not NOT1 (N25321, N25309);
nor NOR3 (N25322, N25320, N2536, N16868);
and AND2 (N25323, N25317, N4055);
xor XOR2 (N25324, N25316, N23427);
not NOT1 (N25325, N25323);
nor NOR2 (N25326, N25315, N8320);
or OR4 (N25327, N25314, N14777, N24798, N3863);
nand NAND2 (N25328, N25325, N17432);
nor NOR3 (N25329, N25318, N23380, N23454);
xor XOR2 (N25330, N25321, N24667);
buf BUF1 (N25331, N25329);
and AND2 (N25332, N25324, N2677);
and AND2 (N25333, N25311, N19779);
nand NAND3 (N25334, N25319, N6583, N20314);
nand NAND2 (N25335, N25330, N7287);
buf BUF1 (N25336, N25327);
not NOT1 (N25337, N25334);
and AND4 (N25338, N25333, N3736, N2988, N10885);
and AND4 (N25339, N25332, N23265, N11587, N9189);
nand NAND4 (N25340, N25275, N16805, N13542, N17321);
not NOT1 (N25341, N25326);
not NOT1 (N25342, N25331);
or OR4 (N25343, N25340, N18787, N13092, N12056);
buf BUF1 (N25344, N25343);
or OR3 (N25345, N25341, N8066, N15347);
nand NAND3 (N25346, N25336, N23169, N22841);
xor XOR2 (N25347, N25345, N11796);
nor NOR2 (N25348, N25342, N6221);
buf BUF1 (N25349, N25339);
nor NOR2 (N25350, N25322, N10689);
xor XOR2 (N25351, N25335, N2376);
nand NAND2 (N25352, N25346, N11130);
and AND4 (N25353, N25328, N221, N4059, N1185);
or OR4 (N25354, N25337, N2446, N20488, N13567);
buf BUF1 (N25355, N25353);
nand NAND4 (N25356, N25352, N8302, N9209, N16954);
or OR4 (N25357, N25356, N17644, N8257, N9201);
buf BUF1 (N25358, N25350);
xor XOR2 (N25359, N25348, N15893);
nor NOR3 (N25360, N25354, N20405, N4351);
xor XOR2 (N25361, N25347, N24401);
not NOT1 (N25362, N25359);
or OR2 (N25363, N25361, N18086);
nand NAND4 (N25364, N25358, N324, N7782, N23311);
xor XOR2 (N25365, N25355, N11454);
and AND3 (N25366, N25351, N6972, N23942);
xor XOR2 (N25367, N25365, N13055);
buf BUF1 (N25368, N25364);
or OR4 (N25369, N25362, N25013, N13870, N21582);
nand NAND4 (N25370, N25360, N13253, N9310, N12070);
and AND2 (N25371, N25367, N10884);
or OR3 (N25372, N25368, N13784, N2892);
buf BUF1 (N25373, N25357);
or OR3 (N25374, N25344, N22788, N17842);
or OR4 (N25375, N25363, N3029, N13597, N16722);
not NOT1 (N25376, N25370);
nor NOR3 (N25377, N25376, N11167, N16004);
and AND2 (N25378, N25349, N23734);
xor XOR2 (N25379, N25373, N8981);
nor NOR4 (N25380, N25369, N9436, N13641, N793);
and AND2 (N25381, N25372, N3527);
xor XOR2 (N25382, N25381, N3808);
nand NAND2 (N25383, N25379, N12680);
not NOT1 (N25384, N25338);
nand NAND3 (N25385, N25375, N12955, N18336);
not NOT1 (N25386, N25366);
xor XOR2 (N25387, N25384, N20808);
or OR2 (N25388, N25380, N6112);
buf BUF1 (N25389, N25371);
or OR4 (N25390, N25387, N4913, N12708, N12704);
nor NOR2 (N25391, N25377, N9762);
nand NAND3 (N25392, N25382, N17565, N20327);
nor NOR4 (N25393, N25389, N11761, N23279, N1620);
buf BUF1 (N25394, N25386);
xor XOR2 (N25395, N25378, N24781);
nor NOR2 (N25396, N25385, N14011);
or OR3 (N25397, N25390, N21086, N17968);
buf BUF1 (N25398, N25395);
nor NOR4 (N25399, N25397, N20398, N7909, N20085);
or OR3 (N25400, N25391, N58, N7119);
and AND2 (N25401, N25396, N25304);
nand NAND4 (N25402, N25383, N20649, N12384, N19404);
not NOT1 (N25403, N25392);
nor NOR2 (N25404, N25400, N5880);
and AND2 (N25405, N25393, N20362);
nor NOR4 (N25406, N25398, N3766, N8961, N10156);
xor XOR2 (N25407, N25402, N9356);
not NOT1 (N25408, N25404);
not NOT1 (N25409, N25399);
not NOT1 (N25410, N25408);
and AND4 (N25411, N25394, N4981, N8827, N10454);
not NOT1 (N25412, N25406);
buf BUF1 (N25413, N25401);
nor NOR2 (N25414, N25409, N6984);
buf BUF1 (N25415, N25412);
nand NAND4 (N25416, N25411, N14748, N24712, N5690);
nand NAND4 (N25417, N25405, N8260, N24091, N19140);
or OR3 (N25418, N25414, N24213, N4728);
nand NAND2 (N25419, N25410, N11882);
xor XOR2 (N25420, N25388, N6888);
or OR4 (N25421, N25418, N2895, N2513, N2011);
and AND2 (N25422, N25419, N2389);
and AND4 (N25423, N25417, N5105, N9976, N8523);
and AND3 (N25424, N25415, N17333, N23784);
not NOT1 (N25425, N25421);
and AND4 (N25426, N25407, N8232, N14109, N22708);
not NOT1 (N25427, N25416);
xor XOR2 (N25428, N25422, N3263);
xor XOR2 (N25429, N25413, N8256);
and AND4 (N25430, N25429, N11892, N4782, N25339);
or OR2 (N25431, N25425, N12784);
and AND3 (N25432, N25427, N12459, N4020);
and AND3 (N25433, N25428, N23767, N6060);
buf BUF1 (N25434, N25432);
or OR2 (N25435, N25420, N4472);
xor XOR2 (N25436, N25423, N12300);
and AND4 (N25437, N25424, N19784, N6826, N23778);
not NOT1 (N25438, N25434);
nor NOR3 (N25439, N25433, N12844, N7320);
not NOT1 (N25440, N25431);
nor NOR4 (N25441, N25437, N19930, N5176, N6867);
not NOT1 (N25442, N25441);
nor NOR2 (N25443, N25435, N23841);
nand NAND2 (N25444, N25403, N16342);
or OR4 (N25445, N25439, N832, N23181, N14391);
buf BUF1 (N25446, N25442);
nor NOR4 (N25447, N25438, N394, N5793, N18461);
xor XOR2 (N25448, N25447, N9660);
xor XOR2 (N25449, N25440, N2995);
nor NOR2 (N25450, N25445, N4640);
buf BUF1 (N25451, N25449);
and AND3 (N25452, N25430, N23245, N11327);
not NOT1 (N25453, N25450);
buf BUF1 (N25454, N25452);
nand NAND4 (N25455, N25443, N25061, N11849, N20583);
nand NAND3 (N25456, N25446, N14599, N16853);
and AND3 (N25457, N25436, N14419, N10341);
xor XOR2 (N25458, N25456, N5032);
nand NAND3 (N25459, N25457, N13958, N25013);
or OR3 (N25460, N25455, N20502, N20437);
not NOT1 (N25461, N25459);
or OR2 (N25462, N25444, N2477);
nand NAND2 (N25463, N25448, N9133);
not NOT1 (N25464, N25374);
and AND3 (N25465, N25454, N1692, N21393);
nor NOR4 (N25466, N25453, N20419, N6866, N20822);
and AND4 (N25467, N25466, N21795, N13639, N15983);
not NOT1 (N25468, N25460);
nor NOR4 (N25469, N25461, N13884, N12517, N12769);
or OR2 (N25470, N25465, N17117);
nand NAND4 (N25471, N25469, N18940, N20844, N8453);
or OR3 (N25472, N25470, N19375, N24888);
not NOT1 (N25473, N25458);
nand NAND4 (N25474, N25472, N1802, N2252, N20860);
and AND2 (N25475, N25451, N10518);
not NOT1 (N25476, N25468);
not NOT1 (N25477, N25474);
nor NOR4 (N25478, N25476, N16288, N14145, N12982);
buf BUF1 (N25479, N25478);
nand NAND4 (N25480, N25463, N5145, N25185, N21561);
xor XOR2 (N25481, N25475, N12187);
or OR3 (N25482, N25467, N17465, N19740);
xor XOR2 (N25483, N25477, N8622);
nor NOR4 (N25484, N25482, N7327, N2837, N11498);
or OR2 (N25485, N25473, N4834);
xor XOR2 (N25486, N25426, N17773);
buf BUF1 (N25487, N25485);
xor XOR2 (N25488, N25480, N25179);
and AND3 (N25489, N25483, N21192, N13830);
xor XOR2 (N25490, N25484, N6906);
nor NOR3 (N25491, N25487, N7111, N17568);
and AND3 (N25492, N25489, N3012, N24712);
nor NOR3 (N25493, N25481, N24842, N21229);
buf BUF1 (N25494, N25491);
buf BUF1 (N25495, N25493);
not NOT1 (N25496, N25494);
xor XOR2 (N25497, N25496, N2118);
and AND4 (N25498, N25462, N4856, N21022, N1815);
nor NOR4 (N25499, N25497, N8863, N14049, N5267);
or OR2 (N25500, N25498, N5655);
not NOT1 (N25501, N25492);
xor XOR2 (N25502, N25490, N13700);
and AND2 (N25503, N25502, N20923);
nand NAND3 (N25504, N25486, N10950, N8522);
xor XOR2 (N25505, N25495, N13703);
or OR3 (N25506, N25503, N7212, N13943);
nor NOR3 (N25507, N25464, N12113, N4928);
xor XOR2 (N25508, N25499, N23029);
nand NAND2 (N25509, N25471, N12558);
and AND3 (N25510, N25500, N16998, N22928);
buf BUF1 (N25511, N25504);
or OR2 (N25512, N25505, N18575);
buf BUF1 (N25513, N25506);
buf BUF1 (N25514, N25488);
not NOT1 (N25515, N25513);
or OR2 (N25516, N25509, N12047);
or OR4 (N25517, N25514, N9095, N13888, N25053);
nor NOR3 (N25518, N25508, N8947, N11706);
buf BUF1 (N25519, N25518);
nor NOR3 (N25520, N25507, N8285, N7748);
xor XOR2 (N25521, N25516, N5040);
nor NOR4 (N25522, N25510, N18903, N14996, N8029);
xor XOR2 (N25523, N25522, N3402);
buf BUF1 (N25524, N25521);
not NOT1 (N25525, N25524);
or OR2 (N25526, N25523, N15051);
xor XOR2 (N25527, N25520, N24709);
xor XOR2 (N25528, N25519, N17712);
and AND4 (N25529, N25528, N9179, N21281, N14610);
not NOT1 (N25530, N25529);
xor XOR2 (N25531, N25479, N15168);
buf BUF1 (N25532, N25501);
and AND3 (N25533, N25517, N5027, N491);
and AND4 (N25534, N25511, N7211, N7264, N21936);
buf BUF1 (N25535, N25531);
nor NOR4 (N25536, N25525, N22495, N20168, N6776);
nor NOR4 (N25537, N25527, N9501, N8578, N4189);
not NOT1 (N25538, N25532);
or OR3 (N25539, N25512, N17500, N24559);
buf BUF1 (N25540, N25537);
nand NAND3 (N25541, N25530, N10795, N9709);
and AND2 (N25542, N25540, N5209);
or OR2 (N25543, N25533, N25162);
buf BUF1 (N25544, N25515);
nor NOR2 (N25545, N25535, N19080);
nor NOR3 (N25546, N25544, N78, N19968);
nor NOR2 (N25547, N25534, N11826);
or OR3 (N25548, N25539, N19647, N17061);
xor XOR2 (N25549, N25546, N7477);
and AND2 (N25550, N25526, N103);
not NOT1 (N25551, N25547);
and AND4 (N25552, N25542, N21617, N8788, N8384);
and AND2 (N25553, N25538, N9498);
nor NOR2 (N25554, N25545, N10435);
and AND2 (N25555, N25551, N13999);
and AND3 (N25556, N25548, N5150, N3702);
not NOT1 (N25557, N25552);
not NOT1 (N25558, N25556);
nand NAND4 (N25559, N25536, N4372, N19713, N18347);
xor XOR2 (N25560, N25550, N2751);
not NOT1 (N25561, N25554);
xor XOR2 (N25562, N25558, N6442);
or OR2 (N25563, N25560, N2082);
and AND2 (N25564, N25557, N24679);
and AND3 (N25565, N25549, N11256, N225);
and AND2 (N25566, N25562, N20146);
and AND3 (N25567, N25559, N4080, N4862);
or OR4 (N25568, N25555, N5951, N984, N11960);
buf BUF1 (N25569, N25561);
nand NAND4 (N25570, N25541, N13432, N10738, N13914);
nand NAND2 (N25571, N25566, N8674);
buf BUF1 (N25572, N25570);
or OR3 (N25573, N25553, N19422, N8914);
not NOT1 (N25574, N25563);
and AND4 (N25575, N25543, N1610, N6654, N16806);
not NOT1 (N25576, N25564);
or OR3 (N25577, N25569, N15986, N20488);
and AND4 (N25578, N25573, N9084, N8214, N3478);
and AND4 (N25579, N25571, N7422, N2105, N22266);
not NOT1 (N25580, N25577);
buf BUF1 (N25581, N25574);
nand NAND2 (N25582, N25572, N18118);
xor XOR2 (N25583, N25576, N12864);
xor XOR2 (N25584, N25565, N4799);
nand NAND3 (N25585, N25584, N9405, N24792);
xor XOR2 (N25586, N25578, N16883);
buf BUF1 (N25587, N25568);
xor XOR2 (N25588, N25587, N12592);
nand NAND4 (N25589, N25575, N136, N17510, N14069);
not NOT1 (N25590, N25580);
nand NAND3 (N25591, N25567, N12905, N17655);
xor XOR2 (N25592, N25582, N5803);
nand NAND4 (N25593, N25591, N6167, N16144, N19196);
xor XOR2 (N25594, N25583, N23688);
not NOT1 (N25595, N25585);
nor NOR4 (N25596, N25590, N22362, N11162, N12296);
xor XOR2 (N25597, N25588, N20016);
not NOT1 (N25598, N25593);
or OR2 (N25599, N25598, N21312);
and AND3 (N25600, N25581, N19326, N7899);
buf BUF1 (N25601, N25592);
not NOT1 (N25602, N25586);
or OR4 (N25603, N25602, N12455, N13252, N6366);
xor XOR2 (N25604, N25600, N18884);
xor XOR2 (N25605, N25597, N10630);
nor NOR3 (N25606, N25596, N1950, N13684);
nand NAND4 (N25607, N25595, N5981, N16672, N19235);
buf BUF1 (N25608, N25607);
xor XOR2 (N25609, N25603, N12958);
or OR3 (N25610, N25605, N7948, N25450);
or OR2 (N25611, N25606, N21876);
not NOT1 (N25612, N25604);
buf BUF1 (N25613, N25608);
or OR4 (N25614, N25613, N6266, N18446, N16179);
buf BUF1 (N25615, N25599);
xor XOR2 (N25616, N25611, N7367);
and AND2 (N25617, N25579, N21096);
and AND4 (N25618, N25609, N24033, N3582, N22611);
nor NOR3 (N25619, N25610, N16458, N5465);
nor NOR2 (N25620, N25594, N20808);
buf BUF1 (N25621, N25619);
buf BUF1 (N25622, N25601);
endmodule