// Verilog Setup

module GateModel (N1);

input N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21;

output N720,N718,N667,N717,N719,N707,N689,N713,N696,N721;

nand NAND4 (N22, N21, N3, N17, N2);
and AND4 (N23, N18, N4, N10, N15);
buf BUF1 (N24, N20);
and AND4 (N25, N8, N22, N7, N11);
or OR4 (N26, N4, N23, N17, N4);
xor XOR2 (N27, N12, N20);
and AND4 (N28, N2, N14, N21, N10);
nand NAND2 (N29, N26, N27);
or OR3 (N30, N20, N1, N2);
and AND2 (N31, N26, N1);
and AND3 (N32, N1, N25, N22);
buf BUF1 (N33, N30);
or OR2 (N34, N7, N13);
not NOT1 (N35, N7);
not NOT1 (N36, N7);
nand NAND2 (N37, N31, N34);
nand NAND3 (N38, N34, N32, N9);
buf BUF1 (N39, N7);
or OR3 (N40, N16, N11, N15);
nor NOR3 (N41, N35, N3, N25);
nand NAND3 (N42, N29, N41, N40);
or OR3 (N43, N11, N5, N36);
nand NAND4 (N44, N17, N10, N20, N43);
not NOT1 (N45, N11);
or OR4 (N46, N27, N7, N21, N11);
or OR2 (N47, N39, N46);
and AND2 (N48, N10, N13);
nand NAND3 (N49, N24, N28, N15);
or OR3 (N50, N43, N3, N3);
not NOT1 (N51, N42);
and AND2 (N52, N38, N27);
or OR2 (N53, N48, N20);
nand NAND4 (N54, N50, N46, N26, N39);
buf BUF1 (N55, N45);
not NOT1 (N56, N33);
xor XOR2 (N57, N53, N1);
nand NAND2 (N58, N47, N27);
nor NOR4 (N59, N49, N10, N14, N42);
xor XOR2 (N60, N44, N1);
nand NAND2 (N61, N60, N31);
nor NOR3 (N62, N37, N32, N60);
not NOT1 (N63, N62);
or OR4 (N64, N61, N22, N26, N57);
or OR2 (N65, N6, N12);
and AND2 (N66, N59, N3);
and AND4 (N67, N55, N39, N34, N20);
xor XOR2 (N68, N54, N7);
buf BUF1 (N69, N63);
and AND3 (N70, N65, N21, N44);
nand NAND4 (N71, N56, N10, N11, N13);
not NOT1 (N72, N52);
nand NAND4 (N73, N58, N65, N46, N1);
nor NOR4 (N74, N72, N27, N53, N34);
nor NOR4 (N75, N74, N11, N30, N6);
not NOT1 (N76, N67);
not NOT1 (N77, N70);
buf BUF1 (N78, N64);
xor XOR2 (N79, N71, N57);
or OR4 (N80, N78, N71, N71, N3);
nand NAND2 (N81, N73, N70);
nand NAND2 (N82, N76, N52);
nand NAND2 (N83, N77, N15);
nand NAND2 (N84, N75, N62);
or OR3 (N85, N69, N45, N48);
xor XOR2 (N86, N51, N43);
or OR4 (N87, N84, N83, N18, N43);
and AND3 (N88, N29, N27, N22);
and AND4 (N89, N82, N71, N48, N51);
xor XOR2 (N90, N66, N76);
or OR2 (N91, N87, N72);
not NOT1 (N92, N85);
not NOT1 (N93, N80);
nor NOR2 (N94, N89, N79);
nand NAND2 (N95, N74, N14);
nand NAND4 (N96, N94, N47, N42, N67);
and AND4 (N97, N95, N72, N56, N71);
nand NAND3 (N98, N96, N48, N60);
xor XOR2 (N99, N91, N93);
not NOT1 (N100, N79);
nor NOR3 (N101, N92, N75, N84);
buf BUF1 (N102, N97);
xor XOR2 (N103, N81, N1);
or OR2 (N104, N90, N74);
or OR4 (N105, N102, N22, N6, N80);
and AND4 (N106, N100, N103, N3, N54);
nand NAND3 (N107, N98, N84, N95);
xor XOR2 (N108, N41, N21);
nor NOR2 (N109, N68, N40);
xor XOR2 (N110, N109, N31);
not NOT1 (N111, N108);
not NOT1 (N112, N86);
nand NAND3 (N113, N105, N33, N48);
buf BUF1 (N114, N111);
nor NOR4 (N115, N88, N37, N66, N39);
nand NAND2 (N116, N99, N72);
xor XOR2 (N117, N114, N77);
not NOT1 (N118, N101);
buf BUF1 (N119, N116);
or OR3 (N120, N119, N76, N84);
not NOT1 (N121, N120);
or OR2 (N122, N104, N49);
not NOT1 (N123, N115);
not NOT1 (N124, N112);
nand NAND3 (N125, N121, N124, N1);
buf BUF1 (N126, N93);
buf BUF1 (N127, N113);
nor NOR4 (N128, N118, N56, N87, N64);
or OR3 (N129, N125, N77, N63);
buf BUF1 (N130, N127);
nor NOR2 (N131, N117, N75);
not NOT1 (N132, N130);
xor XOR2 (N133, N131, N115);
xor XOR2 (N134, N126, N45);
nor NOR2 (N135, N134, N106);
xor XOR2 (N136, N63, N60);
nand NAND2 (N137, N132, N98);
xor XOR2 (N138, N123, N108);
xor XOR2 (N139, N136, N121);
xor XOR2 (N140, N128, N65);
and AND2 (N141, N122, N1);
not NOT1 (N142, N135);
not NOT1 (N143, N137);
xor XOR2 (N144, N133, N99);
or OR4 (N145, N110, N5, N96, N104);
xor XOR2 (N146, N142, N13);
xor XOR2 (N147, N145, N123);
not NOT1 (N148, N144);
not NOT1 (N149, N107);
xor XOR2 (N150, N138, N31);
not NOT1 (N151, N148);
not NOT1 (N152, N149);
and AND4 (N153, N140, N120, N139, N104);
xor XOR2 (N154, N61, N92);
nor NOR2 (N155, N151, N58);
nand NAND3 (N156, N155, N19, N108);
not NOT1 (N157, N154);
xor XOR2 (N158, N141, N26);
nor NOR3 (N159, N153, N155, N39);
and AND3 (N160, N147, N95, N130);
or OR2 (N161, N157, N5);
not NOT1 (N162, N143);
xor XOR2 (N163, N161, N109);
xor XOR2 (N164, N162, N107);
nor NOR3 (N165, N150, N88, N58);
xor XOR2 (N166, N163, N146);
xor XOR2 (N167, N80, N25);
nor NOR4 (N168, N167, N18, N114, N4);
or OR2 (N169, N160, N151);
nor NOR4 (N170, N166, N148, N103, N20);
nor NOR3 (N171, N156, N104, N168);
and AND2 (N172, N26, N105);
buf BUF1 (N173, N170);
xor XOR2 (N174, N164, N139);
buf BUF1 (N175, N172);
not NOT1 (N176, N158);
and AND4 (N177, N173, N33, N79, N109);
buf BUF1 (N178, N175);
or OR2 (N179, N178, N102);
not NOT1 (N180, N169);
nor NOR4 (N181, N152, N169, N128, N152);
nor NOR2 (N182, N171, N173);
nor NOR4 (N183, N180, N109, N82, N126);
buf BUF1 (N184, N183);
or OR2 (N185, N165, N50);
and AND3 (N186, N182, N52, N1);
buf BUF1 (N187, N176);
buf BUF1 (N188, N159);
not NOT1 (N189, N185);
and AND3 (N190, N189, N143, N132);
and AND3 (N191, N177, N69, N70);
and AND3 (N192, N191, N160, N49);
buf BUF1 (N193, N174);
not NOT1 (N194, N186);
nand NAND4 (N195, N188, N186, N35, N149);
buf BUF1 (N196, N179);
xor XOR2 (N197, N190, N60);
not NOT1 (N198, N129);
nor NOR3 (N199, N194, N161, N190);
xor XOR2 (N200, N181, N68);
or OR2 (N201, N192, N55);
not NOT1 (N202, N187);
not NOT1 (N203, N195);
buf BUF1 (N204, N202);
nand NAND3 (N205, N197, N30, N84);
nand NAND2 (N206, N205, N99);
buf BUF1 (N207, N198);
nor NOR3 (N208, N196, N58, N173);
nand NAND2 (N209, N200, N85);
buf BUF1 (N210, N201);
nor NOR4 (N211, N207, N144, N162, N182);
not NOT1 (N212, N199);
nand NAND3 (N213, N203, N165, N100);
xor XOR2 (N214, N213, N8);
not NOT1 (N215, N214);
nand NAND3 (N216, N204, N119, N38);
and AND4 (N217, N210, N133, N79, N107);
nand NAND2 (N218, N215, N175);
xor XOR2 (N219, N206, N34);
not NOT1 (N220, N211);
nand NAND4 (N221, N218, N187, N207, N22);
xor XOR2 (N222, N184, N11);
nor NOR2 (N223, N219, N149);
nand NAND2 (N224, N208, N21);
xor XOR2 (N225, N193, N27);
nor NOR2 (N226, N221, N56);
buf BUF1 (N227, N226);
or OR3 (N228, N222, N185, N17);
nand NAND2 (N229, N225, N180);
nor NOR3 (N230, N209, N7, N89);
and AND3 (N231, N224, N228, N155);
or OR4 (N232, N150, N203, N113, N171);
and AND2 (N233, N229, N143);
buf BUF1 (N234, N233);
xor XOR2 (N235, N216, N64);
or OR4 (N236, N220, N144, N187, N43);
xor XOR2 (N237, N227, N41);
and AND4 (N238, N231, N202, N150, N190);
buf BUF1 (N239, N238);
nor NOR2 (N240, N217, N223);
xor XOR2 (N241, N6, N109);
or OR4 (N242, N236, N112, N67, N43);
nor NOR2 (N243, N240, N119);
not NOT1 (N244, N239);
or OR3 (N245, N242, N212, N193);
or OR3 (N246, N65, N194, N203);
nand NAND2 (N247, N243, N54);
nor NOR3 (N248, N232, N109, N33);
buf BUF1 (N249, N248);
nor NOR2 (N250, N244, N93);
nand NAND4 (N251, N247, N79, N92, N211);
and AND4 (N252, N250, N129, N186, N182);
and AND3 (N253, N235, N74, N243);
not NOT1 (N254, N253);
buf BUF1 (N255, N245);
or OR3 (N256, N237, N239, N203);
nor NOR4 (N257, N230, N131, N144, N128);
and AND3 (N258, N249, N96, N92);
buf BUF1 (N259, N241);
not NOT1 (N260, N251);
and AND2 (N261, N259, N251);
and AND3 (N262, N257, N252, N143);
xor XOR2 (N263, N256, N97);
or OR3 (N264, N18, N103, N169);
nand NAND2 (N265, N234, N165);
or OR2 (N266, N263, N139);
nand NAND3 (N267, N265, N115, N65);
and AND4 (N268, N262, N214, N252, N239);
and AND2 (N269, N255, N80);
or OR3 (N270, N261, N59, N116);
xor XOR2 (N271, N258, N169);
buf BUF1 (N272, N270);
buf BUF1 (N273, N254);
buf BUF1 (N274, N269);
and AND2 (N275, N264, N206);
or OR3 (N276, N274, N169, N266);
or OR2 (N277, N256, N91);
nand NAND2 (N278, N277, N45);
and AND4 (N279, N272, N169, N240, N172);
and AND3 (N280, N273, N142, N47);
buf BUF1 (N281, N246);
and AND4 (N282, N278, N49, N179, N255);
xor XOR2 (N283, N279, N234);
nor NOR3 (N284, N276, N270, N280);
not NOT1 (N285, N90);
and AND2 (N286, N275, N51);
nor NOR2 (N287, N286, N30);
buf BUF1 (N288, N268);
buf BUF1 (N289, N284);
nor NOR4 (N290, N288, N277, N177, N205);
not NOT1 (N291, N260);
xor XOR2 (N292, N281, N171);
nand NAND3 (N293, N267, N73, N75);
nand NAND3 (N294, N282, N252, N173);
nand NAND2 (N295, N285, N235);
nand NAND4 (N296, N294, N46, N264, N237);
buf BUF1 (N297, N283);
nand NAND4 (N298, N295, N68, N167, N38);
nor NOR4 (N299, N291, N73, N93, N106);
not NOT1 (N300, N296);
or OR4 (N301, N298, N263, N144, N56);
nand NAND2 (N302, N287, N208);
nand NAND2 (N303, N299, N182);
not NOT1 (N304, N289);
and AND4 (N305, N297, N57, N167, N100);
nand NAND2 (N306, N301, N195);
xor XOR2 (N307, N302, N198);
not NOT1 (N308, N292);
or OR4 (N309, N271, N166, N39, N7);
nand NAND2 (N310, N305, N51);
and AND4 (N311, N310, N135, N235, N174);
not NOT1 (N312, N307);
not NOT1 (N313, N290);
and AND2 (N314, N306, N231);
buf BUF1 (N315, N303);
and AND3 (N316, N300, N294, N96);
or OR3 (N317, N314, N69, N92);
or OR3 (N318, N312, N210, N202);
buf BUF1 (N319, N316);
xor XOR2 (N320, N319, N121);
buf BUF1 (N321, N309);
buf BUF1 (N322, N308);
and AND4 (N323, N318, N291, N226, N240);
or OR4 (N324, N317, N258, N113, N162);
and AND3 (N325, N321, N206, N279);
nor NOR3 (N326, N325, N284, N79);
buf BUF1 (N327, N304);
and AND4 (N328, N323, N208, N5, N51);
or OR4 (N329, N320, N53, N103, N86);
nand NAND4 (N330, N328, N97, N209, N184);
buf BUF1 (N331, N329);
nor NOR2 (N332, N313, N191);
buf BUF1 (N333, N311);
or OR2 (N334, N327, N278);
not NOT1 (N335, N324);
and AND3 (N336, N335, N251, N35);
buf BUF1 (N337, N334);
buf BUF1 (N338, N315);
or OR3 (N339, N293, N255, N232);
xor XOR2 (N340, N338, N314);
and AND3 (N341, N331, N137, N285);
not NOT1 (N342, N340);
and AND2 (N343, N336, N25);
xor XOR2 (N344, N330, N333);
and AND2 (N345, N115, N86);
not NOT1 (N346, N342);
nor NOR3 (N347, N345, N191, N42);
nor NOR2 (N348, N347, N36);
buf BUF1 (N349, N322);
or OR2 (N350, N337, N28);
xor XOR2 (N351, N326, N119);
nand NAND3 (N352, N351, N174, N320);
and AND4 (N353, N344, N29, N36, N207);
and AND2 (N354, N346, N32);
nor NOR2 (N355, N341, N242);
xor XOR2 (N356, N349, N125);
xor XOR2 (N357, N356, N185);
and AND4 (N358, N350, N117, N339, N211);
buf BUF1 (N359, N350);
nor NOR2 (N360, N352, N151);
and AND2 (N361, N357, N269);
buf BUF1 (N362, N332);
not NOT1 (N363, N343);
buf BUF1 (N364, N358);
xor XOR2 (N365, N354, N38);
nand NAND3 (N366, N362, N139, N148);
xor XOR2 (N367, N359, N70);
not NOT1 (N368, N364);
and AND2 (N369, N355, N213);
buf BUF1 (N370, N348);
xor XOR2 (N371, N353, N86);
not NOT1 (N372, N360);
nor NOR4 (N373, N366, N319, N154, N106);
or OR3 (N374, N368, N162, N146);
xor XOR2 (N375, N367, N38);
or OR3 (N376, N361, N302, N81);
nand NAND3 (N377, N372, N27, N217);
nor NOR3 (N378, N365, N126, N291);
nand NAND4 (N379, N376, N371, N82, N301);
buf BUF1 (N380, N87);
xor XOR2 (N381, N378, N52);
buf BUF1 (N382, N380);
buf BUF1 (N383, N369);
or OR2 (N384, N373, N170);
buf BUF1 (N385, N382);
or OR4 (N386, N384, N260, N322, N131);
nand NAND2 (N387, N375, N134);
buf BUF1 (N388, N383);
nand NAND4 (N389, N379, N328, N95, N22);
or OR4 (N390, N370, N287, N381, N376);
and AND2 (N391, N271, N129);
and AND2 (N392, N377, N297);
xor XOR2 (N393, N392, N23);
buf BUF1 (N394, N385);
not NOT1 (N395, N388);
buf BUF1 (N396, N395);
nand NAND4 (N397, N374, N338, N232, N194);
buf BUF1 (N398, N363);
buf BUF1 (N399, N386);
nor NOR3 (N400, N399, N202, N124);
buf BUF1 (N401, N400);
nor NOR3 (N402, N389, N221, N158);
nand NAND4 (N403, N402, N224, N367, N213);
or OR4 (N404, N397, N75, N271, N382);
nand NAND4 (N405, N404, N1, N180, N38);
xor XOR2 (N406, N405, N97);
xor XOR2 (N407, N403, N183);
or OR2 (N408, N407, N407);
nor NOR2 (N409, N401, N232);
not NOT1 (N410, N394);
or OR3 (N411, N398, N11, N152);
not NOT1 (N412, N387);
buf BUF1 (N413, N408);
or OR3 (N414, N412, N265, N247);
not NOT1 (N415, N414);
buf BUF1 (N416, N406);
or OR2 (N417, N411, N75);
xor XOR2 (N418, N416, N1);
and AND2 (N419, N393, N235);
not NOT1 (N420, N391);
buf BUF1 (N421, N420);
buf BUF1 (N422, N409);
nand NAND2 (N423, N419, N394);
nand NAND3 (N424, N415, N43, N136);
not NOT1 (N425, N423);
nand NAND4 (N426, N417, N142, N183, N48);
buf BUF1 (N427, N426);
and AND2 (N428, N422, N106);
or OR3 (N429, N413, N165, N169);
xor XOR2 (N430, N427, N414);
xor XOR2 (N431, N425, N255);
or OR3 (N432, N396, N380, N232);
nor NOR3 (N433, N418, N159, N415);
nand NAND3 (N434, N431, N261, N277);
or OR3 (N435, N410, N238, N5);
and AND2 (N436, N390, N107);
not NOT1 (N437, N432);
not NOT1 (N438, N436);
and AND3 (N439, N435, N402, N367);
nor NOR4 (N440, N430, N408, N297, N391);
xor XOR2 (N441, N438, N331);
buf BUF1 (N442, N429);
not NOT1 (N443, N433);
not NOT1 (N444, N439);
or OR2 (N445, N424, N100);
or OR2 (N446, N444, N293);
nor NOR2 (N447, N434, N244);
and AND3 (N448, N437, N352, N95);
and AND2 (N449, N445, N363);
or OR4 (N450, N428, N109, N384, N177);
or OR2 (N451, N448, N90);
nor NOR3 (N452, N449, N390, N141);
nor NOR3 (N453, N452, N386, N213);
buf BUF1 (N454, N453);
nor NOR2 (N455, N454, N284);
xor XOR2 (N456, N450, N95);
or OR4 (N457, N443, N183, N325, N221);
or OR4 (N458, N447, N113, N284, N176);
nor NOR3 (N459, N455, N257, N113);
and AND2 (N460, N446, N145);
not NOT1 (N461, N440);
nor NOR2 (N462, N456, N56);
or OR2 (N463, N421, N318);
and AND3 (N464, N461, N137, N356);
buf BUF1 (N465, N464);
buf BUF1 (N466, N460);
xor XOR2 (N467, N465, N159);
not NOT1 (N468, N463);
nand NAND4 (N469, N441, N92, N174, N177);
xor XOR2 (N470, N451, N269);
or OR4 (N471, N462, N127, N449, N310);
xor XOR2 (N472, N459, N414);
xor XOR2 (N473, N467, N166);
not NOT1 (N474, N469);
and AND4 (N475, N457, N246, N63, N239);
and AND4 (N476, N474, N161, N82, N423);
nand NAND2 (N477, N472, N325);
or OR2 (N478, N477, N422);
not NOT1 (N479, N471);
nor NOR2 (N480, N478, N333);
not NOT1 (N481, N480);
and AND2 (N482, N479, N312);
nand NAND3 (N483, N468, N361, N165);
not NOT1 (N484, N470);
xor XOR2 (N485, N475, N158);
nand NAND4 (N486, N458, N77, N127, N84);
or OR3 (N487, N485, N460, N325);
nand NAND3 (N488, N483, N443, N272);
nor NOR3 (N489, N476, N61, N94);
nand NAND4 (N490, N486, N390, N423, N30);
nor NOR2 (N491, N490, N54);
nand NAND2 (N492, N484, N306);
nand NAND4 (N493, N466, N334, N243, N32);
xor XOR2 (N494, N492, N489);
and AND2 (N495, N412, N407);
or OR3 (N496, N482, N453, N206);
and AND3 (N497, N487, N182, N163);
nand NAND4 (N498, N497, N129, N424, N33);
xor XOR2 (N499, N488, N491);
not NOT1 (N500, N66);
not NOT1 (N501, N494);
xor XOR2 (N502, N496, N328);
and AND4 (N503, N501, N304, N136, N26);
xor XOR2 (N504, N481, N274);
nand NAND4 (N505, N495, N128, N28, N480);
nor NOR3 (N506, N442, N461, N160);
or OR3 (N507, N499, N90, N378);
or OR4 (N508, N498, N405, N419, N432);
not NOT1 (N509, N507);
buf BUF1 (N510, N503);
nand NAND4 (N511, N473, N472, N374, N199);
buf BUF1 (N512, N510);
nand NAND3 (N513, N493, N154, N261);
and AND4 (N514, N504, N62, N60, N251);
buf BUF1 (N515, N506);
buf BUF1 (N516, N514);
or OR4 (N517, N513, N290, N159, N50);
and AND3 (N518, N502, N453, N369);
and AND3 (N519, N518, N415, N118);
buf BUF1 (N520, N512);
nor NOR4 (N521, N509, N469, N144, N70);
nand NAND3 (N522, N517, N428, N84);
nor NOR2 (N523, N500, N237);
nand NAND2 (N524, N505, N196);
xor XOR2 (N525, N522, N317);
not NOT1 (N526, N515);
nor NOR4 (N527, N526, N386, N152, N266);
nor NOR2 (N528, N527, N458);
nand NAND2 (N529, N519, N35);
xor XOR2 (N530, N516, N524);
xor XOR2 (N531, N349, N15);
buf BUF1 (N532, N511);
nand NAND4 (N533, N525, N497, N8, N493);
nand NAND3 (N534, N528, N2, N332);
nand NAND4 (N535, N531, N460, N398, N474);
not NOT1 (N536, N532);
and AND2 (N537, N529, N361);
nand NAND4 (N538, N533, N146, N85, N135);
nor NOR3 (N539, N534, N319, N172);
nand NAND3 (N540, N530, N185, N78);
and AND3 (N541, N536, N311, N538);
buf BUF1 (N542, N409);
buf BUF1 (N543, N540);
buf BUF1 (N544, N537);
nor NOR4 (N545, N520, N129, N328, N126);
xor XOR2 (N546, N542, N397);
nor NOR2 (N547, N539, N5);
and AND2 (N548, N543, N516);
or OR2 (N549, N508, N110);
or OR3 (N550, N544, N99, N203);
or OR3 (N551, N521, N267, N331);
buf BUF1 (N552, N549);
buf BUF1 (N553, N552);
xor XOR2 (N554, N523, N165);
or OR4 (N555, N541, N422, N111, N5);
buf BUF1 (N556, N550);
not NOT1 (N557, N535);
nand NAND2 (N558, N557, N77);
xor XOR2 (N559, N556, N306);
and AND2 (N560, N551, N146);
or OR4 (N561, N558, N421, N276, N439);
nand NAND4 (N562, N559, N158, N546, N222);
not NOT1 (N563, N60);
not NOT1 (N564, N560);
nand NAND3 (N565, N561, N36, N202);
or OR4 (N566, N563, N521, N463, N225);
nand NAND2 (N567, N565, N475);
buf BUF1 (N568, N562);
and AND4 (N569, N554, N130, N442, N88);
nor NOR2 (N570, N555, N566);
or OR2 (N571, N447, N361);
and AND3 (N572, N568, N90, N356);
buf BUF1 (N573, N547);
not NOT1 (N574, N564);
buf BUF1 (N575, N572);
buf BUF1 (N576, N553);
xor XOR2 (N577, N569, N213);
not NOT1 (N578, N545);
not NOT1 (N579, N573);
xor XOR2 (N580, N574, N363);
buf BUF1 (N581, N570);
and AND4 (N582, N580, N230, N335, N394);
nor NOR3 (N583, N581, N248, N224);
xor XOR2 (N584, N577, N106);
xor XOR2 (N585, N579, N127);
and AND2 (N586, N575, N408);
and AND2 (N587, N576, N285);
and AND2 (N588, N578, N267);
or OR4 (N589, N585, N368, N428, N176);
not NOT1 (N590, N588);
and AND3 (N591, N548, N432, N94);
not NOT1 (N592, N586);
xor XOR2 (N593, N583, N205);
nand NAND3 (N594, N587, N36, N217);
buf BUF1 (N595, N593);
xor XOR2 (N596, N589, N544);
and AND3 (N597, N595, N517, N388);
buf BUF1 (N598, N567);
not NOT1 (N599, N590);
not NOT1 (N600, N571);
xor XOR2 (N601, N592, N539);
buf BUF1 (N602, N596);
buf BUF1 (N603, N599);
buf BUF1 (N604, N594);
nand NAND3 (N605, N602, N220, N101);
and AND3 (N606, N605, N203, N93);
buf BUF1 (N607, N597);
and AND2 (N608, N601, N226);
nor NOR2 (N609, N607, N484);
and AND4 (N610, N604, N537, N85, N367);
nand NAND3 (N611, N584, N353, N264);
nand NAND2 (N612, N582, N327);
and AND4 (N613, N591, N213, N531, N273);
not NOT1 (N614, N600);
buf BUF1 (N615, N612);
or OR4 (N616, N611, N533, N449, N280);
or OR4 (N617, N616, N246, N439, N322);
xor XOR2 (N618, N613, N113);
buf BUF1 (N619, N618);
xor XOR2 (N620, N603, N295);
not NOT1 (N621, N608);
buf BUF1 (N622, N598);
and AND2 (N623, N609, N46);
or OR4 (N624, N619, N346, N224, N460);
nand NAND4 (N625, N610, N296, N357, N107);
buf BUF1 (N626, N617);
nand NAND4 (N627, N624, N460, N363, N269);
buf BUF1 (N628, N621);
buf BUF1 (N629, N620);
nor NOR4 (N630, N623, N348, N285, N113);
xor XOR2 (N631, N627, N114);
buf BUF1 (N632, N625);
and AND4 (N633, N631, N102, N241, N124);
nor NOR2 (N634, N626, N357);
xor XOR2 (N635, N632, N620);
nand NAND4 (N636, N635, N459, N86, N89);
xor XOR2 (N637, N633, N598);
xor XOR2 (N638, N614, N318);
and AND4 (N639, N622, N110, N305, N260);
and AND3 (N640, N606, N480, N71);
xor XOR2 (N641, N640, N401);
nand NAND3 (N642, N628, N95, N380);
not NOT1 (N643, N638);
and AND2 (N644, N630, N631);
buf BUF1 (N645, N636);
xor XOR2 (N646, N642, N179);
nor NOR3 (N647, N645, N159, N249);
nor NOR2 (N648, N646, N241);
nand NAND3 (N649, N639, N104, N141);
not NOT1 (N650, N649);
xor XOR2 (N651, N647, N650);
buf BUF1 (N652, N171);
or OR3 (N653, N644, N213, N397);
nand NAND4 (N654, N634, N84, N572, N165);
and AND2 (N655, N643, N392);
nand NAND3 (N656, N641, N129, N448);
and AND4 (N657, N656, N60, N472, N228);
xor XOR2 (N658, N653, N523);
or OR4 (N659, N648, N364, N359, N356);
and AND3 (N660, N658, N17, N622);
not NOT1 (N661, N654);
not NOT1 (N662, N657);
and AND4 (N663, N651, N383, N644, N651);
or OR3 (N664, N661, N469, N355);
not NOT1 (N665, N662);
buf BUF1 (N666, N655);
buf BUF1 (N667, N652);
buf BUF1 (N668, N663);
nor NOR4 (N669, N659, N537, N344, N39);
nor NOR3 (N670, N665, N299, N175);
or OR3 (N671, N668, N62, N59);
nand NAND4 (N672, N629, N543, N494, N62);
and AND3 (N673, N615, N191, N290);
or OR2 (N674, N637, N521);
nand NAND2 (N675, N664, N491);
or OR4 (N676, N675, N410, N300, N291);
or OR4 (N677, N669, N75, N382, N74);
not NOT1 (N678, N660);
or OR3 (N679, N666, N1, N641);
and AND3 (N680, N673, N51, N326);
or OR2 (N681, N670, N100);
buf BUF1 (N682, N678);
and AND2 (N683, N672, N401);
nand NAND4 (N684, N674, N379, N587, N100);
or OR2 (N685, N683, N515);
and AND2 (N686, N681, N614);
or OR2 (N687, N685, N164);
not NOT1 (N688, N684);
or OR4 (N689, N688, N47, N158, N140);
nand NAND3 (N690, N680, N439, N133);
or OR4 (N691, N687, N320, N276, N87);
or OR3 (N692, N686, N541, N81);
xor XOR2 (N693, N682, N426);
nand NAND4 (N694, N693, N540, N280, N392);
nand NAND2 (N695, N671, N528);
nor NOR2 (N696, N691, N384);
xor XOR2 (N697, N677, N125);
buf BUF1 (N698, N697);
or OR3 (N699, N694, N371, N498);
xor XOR2 (N700, N690, N195);
nor NOR3 (N701, N698, N3, N693);
xor XOR2 (N702, N676, N179);
xor XOR2 (N703, N679, N130);
nand NAND3 (N704, N700, N7, N477);
nand NAND2 (N705, N703, N38);
or OR2 (N706, N702, N371);
and AND4 (N707, N699, N115, N429, N179);
buf BUF1 (N708, N692);
not NOT1 (N709, N705);
not NOT1 (N710, N708);
or OR4 (N711, N695, N507, N457, N289);
xor XOR2 (N712, N706, N632);
and AND3 (N713, N712, N48, N490);
nand NAND3 (N714, N711, N112, N247);
nand NAND3 (N715, N704, N208, N19);
nand NAND3 (N716, N714, N98, N99);
xor XOR2 (N717, N716, N372);
not NOT1 (N718, N701);
nand NAND2 (N719, N710, N480);
buf BUF1 (N720, N709);
or OR3 (N721, N715, N650, N363);
endmodule